* NGSPICE file created from opamp444.ext - technology: sky130A

.subckt opamp444 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n7636_8799.t28 plus.t5 a_n2903_n3924.t40 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X1 CSoutput.t179 a_n7636_8799.t36 vdd.t293 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X2 CSoutput.t16 commonsourceibias.t48 gnd.t181 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X3 a_n1808_13878.t19 a_n2408_n452.t48 vdd.t295 vdd.t294 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 a_n1808_13878.t11 a_n2408_n452.t31 a_n2408_n452.t32 vdd.t30 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 gnd.t133 gnd.t131 gnd.t132 gnd.t80 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X6 vdd.t292 a_n7636_8799.t37 CSoutput.t178 vdd.t227 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X7 CSoutput.t177 a_n7636_8799.t38 vdd.t291 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X8 gnd.t198 commonsourceibias.t49 CSoutput.t25 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 gnd.t130 gnd.t128 minus.t4 gnd.t129 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X10 CSoutput.t57 commonsourceibias.t50 gnd.t288 gnd.t287 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 CSoutput.t24 commonsourceibias.t51 gnd.t196 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X12 CSoutput.t176 a_n7636_8799.t39 vdd.t290 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X13 a_n2903_n3924.t33 plus.t6 a_n7636_8799.t27 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X14 output.t19 outputibias.t8 gnd.t221 gnd.t220 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X15 vdd.t129 vdd.t127 vdd.t128 vdd.t81 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X16 a_n2903_n3924.t14 minus.t5 a_n2408_n452.t34 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X17 a_n1986_8322.t19 a_n2408_n452.t49 a_n7636_8799.t35 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X18 vdd.t2 CSoutput.t192 output.t15 gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X19 CSoutput.t175 a_n7636_8799.t40 vdd.t289 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X20 gnd.t274 commonsourceibias.t52 CSoutput.t51 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X21 CSoutput.t56 commonsourceibias.t53 gnd.t286 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 gnd.t195 commonsourceibias.t54 CSoutput.t23 gnd.t151 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X23 vdd.t288 a_n7636_8799.t41 CSoutput.t174 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X24 CSoutput.t50 commonsourceibias.t55 gnd.t273 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 CSoutput.t55 commonsourceibias.t56 gnd.t285 gnd.t155 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 a_n2408_n452.t42 minus.t6 a_n2903_n3924.t49 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X27 gnd.t127 gnd.t124 gnd.t126 gnd.t125 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X28 CSoutput.t187 commonsourceibias.t57 gnd.t308 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X29 vdd.t287 a_n7636_8799.t42 CSoutput.t173 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X30 a_n2408_n452.t35 minus.t7 a_n2903_n3924.t15 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X31 CSoutput.t172 a_n7636_8799.t43 vdd.t286 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X32 vdd.t285 a_n7636_8799.t44 CSoutput.t171 vdd.t245 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X33 vdd.t284 a_n7636_8799.t45 CSoutput.t170 vdd.t271 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X34 a_n7636_8799.t33 a_n2408_n452.t50 a_n1986_8322.t18 vdd.t50 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X35 CSoutput.t9 commonsourceibias.t58 gnd.t163 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 gnd.t9 commonsourceibias.t59 CSoutput.t1 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 CSoutput.t169 a_n7636_8799.t46 vdd.t283 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X38 gnd.t123 gnd.t121 gnd.t122 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X39 CSoutput.t21 commonsourceibias.t60 gnd.t187 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 CSoutput.t193 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X41 a_n2903_n3924.t20 minus.t8 a_n2408_n452.t39 gnd.t232 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X42 CSoutput.t190 commonsourceibias.t61 gnd.t316 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 CSoutput.t168 a_n7636_8799.t47 vdd.t282 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X44 vdd.t126 vdd.t124 vdd.t125 vdd.t59 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X45 a_n2903_n3924.t12 diffpairibias.t16 gnd.t212 gnd.t211 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X46 CSoutput.t167 a_n7636_8799.t48 vdd.t281 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X47 gnd.t158 commonsourceibias.t62 CSoutput.t7 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X48 gnd.t120 gnd.t117 gnd.t119 gnd.t118 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X49 CSoutput.t45 commonsourceibias.t63 gnd.t268 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X50 gnd.t207 commonsourceibias.t46 commonsourceibias.t47 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 CSoutput.t29 commonsourceibias.t64 gnd.t216 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 CSoutput.t166 a_n7636_8799.t49 vdd.t280 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 a_n2903_n3924.t28 plus.t7 a_n7636_8799.t26 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X54 a_n1808_13878.t10 a_n2408_n452.t13 a_n2408_n452.t14 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X55 CSoutput.t59 commonsourceibias.t65 gnd.t296 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 vdd.t279 a_n7636_8799.t50 CSoutput.t165 vdd.t271 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X57 vdd.t123 vdd.t121 vdd.t122 vdd.t81 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X58 a_n7636_8799.t25 plus.t8 a_n2903_n3924.t37 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X59 CSoutput.t164 a_n7636_8799.t51 vdd.t278 vdd.t225 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X60 a_n2408_n452.t24 a_n2408_n452.t23 a_n1808_13878.t9 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X61 outputibias.t7 outputibias.t6 gnd.t323 gnd.t322 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X62 gnd.t272 commonsourceibias.t66 CSoutput.t49 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X63 a_n7636_8799.t24 plus.t9 a_n2903_n3924.t39 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X64 CSoutput.t163 a_n7636_8799.t52 vdd.t277 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X65 gnd.t208 commonsourceibias.t44 commonsourceibias.t45 gnd.t153 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X66 vdd.t120 vdd.t118 vdd.t119 vdd.t94 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X67 CSoutput.t4 commonsourceibias.t67 gnd.t139 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 vdd.t276 a_n7636_8799.t53 CSoutput.t162 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X69 gnd.t116 gnd.t114 gnd.t115 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X70 gnd.t113 gnd.t111 gnd.t112 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X71 CSoutput.t48 commonsourceibias.t68 gnd.t271 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X72 diffpairibias.t15 diffpairibias.t14 gnd.t223 gnd.t222 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X73 a_n2903_n3924.t26 plus.t10 a_n7636_8799.t23 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X74 a_n2408_n452.t47 minus.t9 a_n2903_n3924.t54 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X75 CSoutput.t8 commonsourceibias.t69 gnd.t161 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X76 CSoutput.t0 commonsourceibias.t70 gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X77 gnd.t291 commonsourceibias.t71 CSoutput.t58 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 CSoutput.t161 a_n7636_8799.t54 vdd.t275 vdd.t229 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X79 gnd.t240 commonsourceibias.t72 CSoutput.t37 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 gnd.t110 gnd.t108 plus.t1 gnd.t109 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X81 vdd.t274 a_n7636_8799.t55 CSoutput.t160 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 vdd.t273 a_n7636_8799.t56 CSoutput.t159 vdd.t245 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 vdd.t272 a_n7636_8799.t57 CSoutput.t158 vdd.t271 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X84 vdd.t270 a_n7636_8799.t58 CSoutput.t157 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X85 CSoutput.t189 commonsourceibias.t73 gnd.t315 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X86 diffpairibias.t13 diffpairibias.t12 gnd.t148 gnd.t147 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X87 CSoutput.t156 a_n7636_8799.t59 vdd.t269 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X88 CSoutput.t155 a_n7636_8799.t60 vdd.t268 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X89 gnd.t279 commonsourceibias.t42 commonsourceibias.t43 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 CSoutput.t6 commonsourceibias.t74 gnd.t156 gnd.t155 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 gnd.t267 commonsourceibias.t75 CSoutput.t44 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X92 output.t14 CSoutput.t194 vdd.t3 gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X93 CSoutput.t28 commonsourceibias.t76 gnd.t215 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 vdd.t267 a_n7636_8799.t61 CSoutput.t154 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X95 CSoutput.t153 a_n7636_8799.t62 vdd.t266 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 gnd.t239 commonsourceibias.t77 CSoutput.t36 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X97 CSoutput.t152 a_n7636_8799.t63 vdd.t265 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X98 CSoutput.t151 a_n7636_8799.t64 vdd.t263 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X99 CSoutput.t150 a_n7636_8799.t65 vdd.t264 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X100 vdd.t262 a_n7636_8799.t66 CSoutput.t149 vdd.t250 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X101 gnd.t107 gnd.t105 gnd.t106 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X102 gnd.t104 gnd.t102 plus.t0 gnd.t103 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X103 output.t13 CSoutput.t195 vdd.t16 gnd.t217 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X104 a_n2903_n3924.t24 plus.t11 a_n7636_8799.t22 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X105 gnd.t270 commonsourceibias.t78 CSoutput.t47 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X106 a_n2903_n3924.t48 diffpairibias.t17 gnd.t276 gnd.t275 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X107 vdd.t261 a_n7636_8799.t67 CSoutput.t148 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X108 gnd.t101 gnd.t99 gnd.t100 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X109 a_n2408_n452.t26 a_n2408_n452.t25 a_n1808_13878.t8 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X110 vdd.t260 a_n7636_8799.t68 CSoutput.t147 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X111 gnd.t269 commonsourceibias.t79 CSoutput.t46 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X112 a_n7636_8799.t34 a_n2408_n452.t51 a_n1986_8322.t17 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X113 vdd.t259 a_n7636_8799.t69 CSoutput.t146 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X114 a_n2408_n452.t30 a_n2408_n452.t29 a_n1808_13878.t7 vdd.t10 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X115 gnd.t98 gnd.t96 gnd.t97 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X116 vdd.t258 a_n7636_8799.t70 CSoutput.t145 vdd.t250 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X117 vdd.t232 a_n7636_8799.t71 CSoutput.t144 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X118 CSoutput.t143 a_n7636_8799.t72 vdd.t257 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X119 gnd.t238 commonsourceibias.t80 CSoutput.t35 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 a_n2408_n452.t8 minus.t10 a_n2903_n3924.t8 gnd.t142 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X121 output.t12 CSoutput.t196 vdd.t17 gnd.t218 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X122 vdd.t117 vdd.t115 vdd.t116 vdd.t102 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X123 vdd.t256 a_n7636_8799.t73 CSoutput.t142 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X124 gnd.t209 commonsourceibias.t40 commonsourceibias.t41 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X125 gnd.t237 commonsourceibias.t81 CSoutput.t34 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X126 CSoutput.t141 a_n7636_8799.t74 vdd.t255 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X127 vdd.t114 vdd.t111 vdd.t113 vdd.t112 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X128 output.t18 outputibias.t9 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X129 CSoutput.t197 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X130 a_n2903_n3924.t47 minus.t11 a_n2408_n452.t41 gnd.t256 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X131 vdd.t110 vdd.t108 vdd.t109 vdd.t55 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X132 gnd.t95 gnd.t92 gnd.t94 gnd.t93 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X133 vdd.t107 vdd.t105 vdd.t106 vdd.t98 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X134 vdd.t36 a_n2408_n452.t52 a_n1986_8322.t7 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X135 a_n1986_8322.t6 a_n2408_n452.t53 vdd.t38 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X136 a_n2903_n3924.t11 diffpairibias.t18 gnd.t202 gnd.t201 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X137 CSoutput.t140 a_n7636_8799.t75 vdd.t254 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X138 CSoutput.t139 a_n7636_8799.t76 vdd.t252 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X139 outputibias.t5 outputibias.t4 gnd.t144 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X140 vdd.t18 CSoutput.t198 output.t11 gnd.t219 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X141 CSoutput.t33 commonsourceibias.t82 gnd.t236 gnd.t155 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X142 CSoutput.t32 commonsourceibias.t83 gnd.t235 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X143 gnd.t91 gnd.t89 gnd.t90 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X144 vdd.t251 a_n7636_8799.t77 CSoutput.t138 vdd.t250 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X145 a_n2903_n3924.t2 minus.t12 a_n2408_n452.t2 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X146 a_n2903_n3924.t52 minus.t13 a_n2408_n452.t45 gnd.t258 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X147 vdd.t32 a_n2408_n452.t54 a_n1808_13878.t18 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X148 a_n2408_n452.t38 minus.t14 a_n2903_n3924.t19 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X149 a_n2903_n3924.t34 plus.t12 a_n7636_8799.t21 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X150 outputibias.t3 outputibias.t2 gnd.t325 gnd.t324 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X151 a_n2903_n3924.t27 plus.t13 a_n7636_8799.t20 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X152 vdd.t104 vdd.t101 vdd.t103 vdd.t102 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X153 a_n2408_n452.t3 minus.t15 a_n2903_n3924.t3 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X154 gnd.t88 gnd.t86 gnd.t87 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X155 vdd.t100 vdd.t97 vdd.t99 vdd.t98 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X156 vdd.t249 a_n7636_8799.t78 CSoutput.t137 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X157 gnd.t85 gnd.t83 plus.t2 gnd.t84 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X158 a_n7636_8799.t19 plus.t14 a_n2903_n3924.t29 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X159 a_n7636_8799.t18 plus.t15 a_n2903_n3924.t38 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X160 vdd.t96 vdd.t93 vdd.t95 vdd.t94 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X161 a_n1986_8322.t5 a_n2408_n452.t55 vdd.t34 vdd.t33 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X162 a_n7636_8799.t3 a_n2408_n452.t56 a_n1986_8322.t16 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X163 CSoutput.t136 a_n7636_8799.t79 vdd.t247 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X164 diffpairibias.t11 diffpairibias.t10 gnd.t300 gnd.t299 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X165 vdd.t246 a_n7636_8799.t80 CSoutput.t135 vdd.t245 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X166 a_n2408_n452.t33 minus.t16 a_n2903_n3924.t13 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X167 a_n2408_n452.t10 a_n2408_n452.t9 a_n1808_13878.t6 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X168 vdd.t244 a_n7636_8799.t81 CSoutput.t134 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X169 CSoutput.t186 commonsourceibias.t84 gnd.t307 gnd.t287 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X170 vdd.t51 CSoutput.t199 output.t10 gnd.t292 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X171 a_n7636_8799.t4 a_n2408_n452.t57 a_n1986_8322.t15 vdd.t30 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X172 CSoutput.t133 a_n7636_8799.t82 vdd.t243 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X173 commonsourceibias.t39 commonsourceibias.t38 gnd.t280 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X174 output.t9 CSoutput.t200 vdd.t52 gnd.t293 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X175 gnd.t306 commonsourceibias.t85 CSoutput.t185 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X176 a_n1808_13878.t5 a_n2408_n452.t27 a_n2408_n452.t28 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X177 a_n2903_n3924.t51 minus.t17 a_n2408_n452.t44 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X178 CSoutput.t201 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X179 output.t8 CSoutput.t202 vdd.t53 gnd.t294 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X180 CSoutput.t132 a_n7636_8799.t83 vdd.t233 vdd.t229 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X181 gnd.t82 gnd.t79 gnd.t81 gnd.t80 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X182 CSoutput.t184 commonsourceibias.t86 gnd.t305 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 vdd.t131 a_n2408_n452.t58 a_n1986_8322.t4 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X184 CSoutput.t203 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X185 vdd.t242 a_n7636_8799.t84 CSoutput.t131 vdd.t227 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X186 gnd.t301 commonsourceibias.t87 CSoutput.t180 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 gnd.t304 commonsourceibias.t88 CSoutput.t183 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 commonsourceibias.t37 commonsourceibias.t36 gnd.t241 gnd.t155 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 minus.t3 gnd.t76 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X190 CSoutput.t130 a_n7636_8799.t85 vdd.t241 vdd.t225 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X191 gnd.t303 commonsourceibias.t89 CSoutput.t182 gnd.t151 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X192 vdd.t240 a_n7636_8799.t86 CSoutput.t129 vdd.t140 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X193 outputibias.t1 outputibias.t0 gnd.t327 gnd.t326 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X194 a_n2903_n3924.t35 plus.t16 a_n7636_8799.t17 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X195 vdd.t239 a_n7636_8799.t87 CSoutput.t128 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X196 CSoutput.t40 commonsourceibias.t90 gnd.t253 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X197 a_n2903_n3924.t10 diffpairibias.t19 gnd.t200 gnd.t199 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X198 gnd.t75 gnd.t72 gnd.t74 gnd.t73 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X199 a_n2903_n3924.t9 diffpairibias.t20 gnd.t146 gnd.t145 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X200 commonsourceibias.t35 commonsourceibias.t34 gnd.t242 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 output.t17 outputibias.t10 gnd.t311 gnd.t310 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X202 vdd.t238 a_n7636_8799.t88 CSoutput.t127 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X203 vdd.t237 a_n7636_8799.t89 CSoutput.t126 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X204 a_n7636_8799.t16 plus.t17 a_n2903_n3924.t41 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X205 gnd.t71 gnd.t69 gnd.t70 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X206 vdd.t7 CSoutput.t204 output.t7 gnd.t172 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X207 CSoutput.t181 commonsourceibias.t91 gnd.t302 gnd.t287 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X208 CSoutput.t20 commonsourceibias.t92 gnd.t186 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X209 gnd.t68 gnd.t66 gnd.t67 gnd.t18 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X210 CSoutput.t125 a_n7636_8799.t90 vdd.t236 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X211 CSoutput.t124 a_n7636_8799.t91 vdd.t235 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X212 commonsourceibias.t33 commonsourceibias.t32 gnd.t210 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 CSoutput.t123 a_n7636_8799.t92 vdd.t231 vdd.t209 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X214 diffpairibias.t9 diffpairibias.t8 gnd.t230 gnd.t229 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X215 a_n1808_13878.t17 a_n2408_n452.t59 vdd.t133 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X216 vdd.t45 a_n2408_n452.t60 a_n1808_13878.t16 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X217 vdd.t92 vdd.t90 vdd.t91 vdd.t66 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X218 CSoutput.t15 commonsourceibias.t93 gnd.t180 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X219 CSoutput.t19 commonsourceibias.t94 gnd.t184 gnd.t134 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 vdd.t89 vdd.t87 vdd.t88 vdd.t74 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X221 CSoutput.t122 a_n7636_8799.t93 vdd.t230 vdd.t229 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X222 gnd.t243 commonsourceibias.t30 commonsourceibias.t31 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X223 vdd.t228 a_n7636_8799.t94 CSoutput.t121 vdd.t227 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X224 vdd.t86 vdd.t84 vdd.t85 vdd.t74 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X225 commonsourceibias.t29 commonsourceibias.t28 gnd.t281 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 plus.t3 gnd.t63 gnd.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X227 a_n2903_n3924.t5 minus.t18 a_n2408_n452.t5 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X228 gnd.t178 commonsourceibias.t95 CSoutput.t14 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X229 CSoutput.t120 a_n7636_8799.t95 vdd.t226 vdd.t225 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X230 commonsourceibias.t27 commonsourceibias.t26 gnd.t244 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X231 vdd.t224 a_n7636_8799.t96 CSoutput.t119 vdd.t140 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X232 vdd.t223 a_n7636_8799.t97 CSoutput.t118 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X233 a_n2408_n452.t7 minus.t19 a_n2903_n3924.t7 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X234 gnd.t245 commonsourceibias.t24 commonsourceibias.t25 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 a_n1986_8322.t14 a_n2408_n452.t61 a_n7636_8799.t31 vdd.t46 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X236 CSoutput.t117 a_n7636_8799.t98 vdd.t222 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X237 gnd.t62 gnd.t59 gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X238 diffpairibias.t7 diffpairibias.t6 gnd.t320 gnd.t319 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X239 gnd.t58 gnd.t56 gnd.t57 gnd.t18 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X240 vdd.t221 a_n7636_8799.t99 CSoutput.t116 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X241 commonsourceibias.t23 commonsourceibias.t22 gnd.t164 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X242 a_n2408_n452.t1 minus.t20 a_n2903_n3924.t1 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X243 CSoutput.t115 a_n7636_8799.t100 vdd.t219 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X244 a_n2408_n452.t43 minus.t21 a_n2903_n3924.t50 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X245 vdd.t218 a_n7636_8799.t101 CSoutput.t114 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X246 vdd.t27 a_n2408_n452.t62 a_n1986_8322.t3 vdd.t26 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X247 output.t6 CSoutput.t205 vdd.t8 gnd.t173 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X248 vdd.t216 a_n7636_8799.t102 CSoutput.t113 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X249 vdd.t215 a_n7636_8799.t103 CSoutput.t112 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X250 a_n2903_n3924.t53 minus.t22 a_n2408_n452.t46 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X251 a_n7636_8799.t15 plus.t18 a_n2903_n3924.t30 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X252 gnd.t183 commonsourceibias.t96 CSoutput.t18 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 output.t16 outputibias.t11 gnd.t290 gnd.t289 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X254 a_n2903_n3924.t22 minus.t23 a_n2408_n452.t40 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X255 gnd.t252 commonsourceibias.t20 commonsourceibias.t21 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X256 a_n1808_13878.t15 a_n2408_n452.t63 vdd.t29 vdd.t28 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X257 output.t5 CSoutput.t206 vdd.t9 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X258 vdd.t213 a_n7636_8799.t104 CSoutput.t111 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X259 CSoutput.t110 a_n7636_8799.t105 vdd.t212 vdd.t209 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X260 CSoutput.t109 a_n7636_8799.t106 vdd.t211 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X261 gnd.t55 gnd.t53 minus.t2 gnd.t54 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X262 vdd.t83 vdd.t80 vdd.t82 vdd.t81 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X263 gnd.t52 gnd.t49 gnd.t51 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X264 vdd.t79 vdd.t77 vdd.t78 vdd.t66 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X265 a_n2903_n3924.t21 diffpairibias.t21 gnd.t247 gnd.t246 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X266 vdd.t76 vdd.t73 vdd.t75 vdd.t74 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X267 vdd.t40 a_n2408_n452.t64 a_n1986_8322.t2 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X268 a_n1986_8322.t13 a_n2408_n452.t65 a_n7636_8799.t29 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X269 CSoutput.t108 a_n7636_8799.t107 vdd.t210 vdd.t209 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X270 gnd.t251 commonsourceibias.t18 commonsourceibias.t19 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X271 vdd.t208 a_n7636_8799.t108 CSoutput.t107 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X272 CSoutput.t106 a_n7636_8799.t109 vdd.t207 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 CSoutput.t207 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X274 vdd.t206 a_n7636_8799.t110 CSoutput.t105 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X275 vdd.t205 a_n7636_8799.t111 CSoutput.t104 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X276 a_n7636_8799.t14 plus.t19 a_n2903_n3924.t25 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X277 gnd.t160 commonsourceibias.t16 commonsourceibias.t17 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 vdd.t72 vdd.t69 vdd.t71 vdd.t70 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X279 a_n2903_n3924.t36 plus.t20 a_n7636_8799.t13 gnd.t232 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X280 vdd.t4 CSoutput.t208 output.t4 gnd.t165 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X281 vdd.t204 a_n7636_8799.t112 CSoutput.t103 vdd.t148 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X282 vdd.t5 CSoutput.t209 output.t3 gnd.t166 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X283 CSoutput.t102 a_n7636_8799.t113 vdd.t203 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X284 CSoutput.t13 commonsourceibias.t97 gnd.t176 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X285 a_n1808_13878.t4 a_n2408_n452.t19 a_n2408_n452.t20 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X286 CSoutput.t101 a_n7636_8799.t114 vdd.t201 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X287 a_n1986_8322.t12 a_n2408_n452.t66 a_n7636_8799.t2 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X288 diffpairibias.t5 diffpairibias.t4 gnd.t278 gnd.t277 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X289 gnd.t48 gnd.t45 gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X290 CSoutput.t100 a_n7636_8799.t115 vdd.t200 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X291 CSoutput.t99 a_n7636_8799.t116 vdd.t198 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X292 vdd.t197 a_n7636_8799.t117 CSoutput.t98 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 CSoutput.t41 commonsourceibias.t98 gnd.t254 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X294 vdd.t196 a_n7636_8799.t118 CSoutput.t97 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X295 a_n1986_8322.t1 a_n2408_n452.t67 vdd.t21 vdd.t20 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X296 CSoutput.t96 a_n7636_8799.t119 vdd.t194 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X297 gnd.t44 gnd.t42 gnd.t43 gnd.t18 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X298 gnd.t255 commonsourceibias.t99 CSoutput.t42 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X299 vdd.t42 a_n2408_n452.t68 a_n1808_13878.t14 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X300 plus.t4 gnd.t39 gnd.t41 gnd.t40 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X301 CSoutput.t95 a_n7636_8799.t120 vdd.t192 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X302 CSoutput.t94 a_n7636_8799.t121 vdd.t190 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X303 a_n2903_n3924.t46 plus.t21 a_n7636_8799.t12 gnd.t258 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X304 vdd.t137 a_n7636_8799.t122 CSoutput.t93 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X305 vdd.t189 a_n7636_8799.t123 CSoutput.t92 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X306 vdd.t68 vdd.t65 vdd.t67 vdd.t66 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X307 gnd.t249 commonsourceibias.t100 CSoutput.t38 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X308 gnd.t284 commonsourceibias.t101 CSoutput.t54 gnd.t153 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X309 output.t2 CSoutput.t210 vdd.t6 gnd.t167 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X310 a_n2903_n3924.t6 minus.t24 a_n2408_n452.t6 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X311 gnd.t38 gnd.t36 gnd.t37 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X312 a_n1986_8322.t11 a_n2408_n452.t69 a_n7636_8799.t30 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X313 vdd.t64 vdd.t62 vdd.t63 vdd.t59 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X314 commonsourceibias.t15 commonsourceibias.t14 gnd.t298 gnd.t287 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 vdd.t0 CSoutput.t211 output.t1 gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X316 CSoutput.t91 a_n7636_8799.t124 vdd.t188 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X317 a_n7636_8799.t32 a_n2408_n452.t70 a_n1986_8322.t10 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X318 a_n7636_8799.t11 plus.t22 a_n2903_n3924.t32 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X319 vdd.t186 a_n7636_8799.t125 CSoutput.t90 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X320 a_n1808_13878.t13 a_n2408_n452.t71 vdd.t49 vdd.t48 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X321 gnd.t283 commonsourceibias.t102 CSoutput.t53 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X322 vdd.t184 a_n7636_8799.t126 CSoutput.t89 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X323 a_n2408_n452.t4 minus.t25 a_n2903_n3924.t4 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X324 CSoutput.t88 a_n7636_8799.t127 vdd.t183 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 gnd.t282 commonsourceibias.t103 CSoutput.t52 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 commonsourceibias.t13 commonsourceibias.t12 gnd.t150 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X327 a_n7636_8799.t10 plus.t23 a_n2903_n3924.t31 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X328 gnd.t35 gnd.t32 gnd.t34 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X329 gnd.t31 gnd.t29 minus.t1 gnd.t30 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X330 gnd.t314 commonsourceibias.t104 CSoutput.t188 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X331 a_n2903_n3924.t17 minus.t26 a_n2408_n452.t37 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X332 vdd.t181 a_n7636_8799.t128 CSoutput.t87 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X333 gnd.t189 commonsourceibias.t10 commonsourceibias.t11 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X334 CSoutput.t86 a_n7636_8799.t129 vdd.t179 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X335 CSoutput.t85 a_n7636_8799.t130 vdd.t177 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X336 CSoutput.t84 a_n7636_8799.t131 vdd.t176 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X337 a_n1808_13878.t3 a_n2408_n452.t11 a_n2408_n452.t12 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X338 CSoutput.t83 a_n7636_8799.t132 vdd.t175 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 a_n2903_n3924.t23 plus.t24 a_n7636_8799.t9 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X340 vdd.t174 a_n7636_8799.t133 CSoutput.t82 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X341 gnd.t152 commonsourceibias.t8 commonsourceibias.t9 gnd.t151 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X342 commonsourceibias.t7 commonsourceibias.t6 gnd.t295 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X343 CSoutput.t81 a_n7636_8799.t134 vdd.t173 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X344 gnd.t321 commonsourceibias.t105 CSoutput.t191 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X345 a_n2903_n3924.t55 diffpairibias.t22 gnd.t318 gnd.t317 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X346 CSoutput.t43 commonsourceibias.t106 gnd.t265 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X347 vdd.t172 a_n7636_8799.t135 CSoutput.t80 vdd.t148 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X348 vdd.t171 a_n7636_8799.t136 CSoutput.t79 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X349 gnd.t250 commonsourceibias.t107 CSoutput.t39 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X350 CSoutput.t78 a_n7636_8799.t137 vdd.t170 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X351 a_n2408_n452.t22 a_n2408_n452.t21 a_n1808_13878.t2 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X352 gnd.t28 gnd.t25 gnd.t27 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X353 a_n7636_8799.t1 a_n2408_n452.t72 a_n1986_8322.t9 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X354 vdd.t1 CSoutput.t212 output.t0 gnd.t11 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X355 gnd.t24 gnd.t21 gnd.t23 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X356 vdd.t139 a_n7636_8799.t138 CSoutput.t77 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X357 CSoutput.t76 a_n7636_8799.t139 vdd.t169 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X358 a_n7636_8799.t8 plus.t25 a_n2903_n3924.t42 gnd.t142 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X359 vdd.t167 a_n7636_8799.t140 CSoutput.t75 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X360 CSoutput.t31 commonsourceibias.t108 gnd.t234 gnd.t134 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X361 gnd.t171 commonsourceibias.t109 CSoutput.t12 gnd.t151 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X362 commonsourceibias.t5 commonsourceibias.t4 gnd.t309 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X363 diffpairibias.t3 diffpairibias.t2 gnd.t264 gnd.t263 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X364 gnd.t20 gnd.t17 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X365 vdd.t166 a_n7636_8799.t141 CSoutput.t74 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X366 vdd.t61 vdd.t58 vdd.t60 vdd.t59 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X367 CSoutput.t73 a_n7636_8799.t142 vdd.t164 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X368 gnd.t233 commonsourceibias.t110 CSoutput.t30 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X369 a_n2903_n3924.t44 plus.t26 a_n7636_8799.t7 gnd.t256 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X370 vdd.t162 a_n7636_8799.t143 CSoutput.t72 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X371 CSoutput.t213 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X372 diffpairibias.t1 diffpairibias.t0 gnd.t313 gnd.t312 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X373 commonsourceibias.t3 commonsourceibias.t2 gnd.t194 gnd.t134 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X374 gnd.t205 commonsourceibias.t111 CSoutput.t27 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X375 a_n2903_n3924.t45 plus.t27 a_n7636_8799.t6 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X376 CSoutput.t3 commonsourceibias.t112 gnd.t137 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X377 vdd.t15 a_n2408_n452.t73 a_n1808_13878.t12 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X378 a_n7636_8799.t5 plus.t28 a_n2903_n3924.t43 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X379 CSoutput.t71 a_n7636_8799.t144 vdd.t160 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X380 a_n2903_n3924.t0 minus.t27 a_n2408_n452.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X381 CSoutput.t70 a_n7636_8799.t145 vdd.t158 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X382 vdd.t156 a_n7636_8799.t146 CSoutput.t69 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X383 vdd.t154 a_n7636_8799.t147 CSoutput.t68 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X384 gnd.t297 commonsourceibias.t0 commonsourceibias.t1 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X385 CSoutput.t67 a_n7636_8799.t148 vdd.t153 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X386 a_n2408_n452.t36 minus.t28 a_n2903_n3924.t16 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X387 CSoutput.t66 a_n7636_8799.t149 vdd.t151 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X388 gnd.t170 commonsourceibias.t113 CSoutput.t11 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X389 gnd.t204 commonsourceibias.t114 CSoutput.t26 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X390 a_n1986_8322.t8 a_n2408_n452.t74 a_n7636_8799.t0 vdd.t10 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X391 vdd.t149 a_n7636_8799.t150 CSoutput.t65 vdd.t148 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X392 vdd.t147 a_n7636_8799.t151 CSoutput.t64 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X393 CSoutput.t63 a_n7636_8799.t152 vdd.t145 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X394 CSoutput.t62 a_n7636_8799.t153 vdd.t143 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X395 vdd.t141 a_n7636_8799.t154 CSoutput.t61 vdd.t140 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X396 gnd.t154 commonsourceibias.t115 CSoutput.t5 gnd.t153 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X397 a_n1986_8322.t0 a_n2408_n452.t75 vdd.t12 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X398 gnd.t182 commonsourceibias.t116 CSoutput.t17 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X399 a_n1808_13878.t1 a_n2408_n452.t17 a_n2408_n452.t18 vdd.t50 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X400 gnd.t168 commonsourceibias.t117 CSoutput.t10 gnd.t153 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X401 CSoutput.t2 commonsourceibias.t118 gnd.t135 gnd.t134 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X402 vdd.t135 a_n7636_8799.t155 CSoutput.t60 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X403 CSoutput.t22 commonsourceibias.t119 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X404 minus.t0 gnd.t14 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X405 a_n2903_n3924.t18 diffpairibias.t23 gnd.t228 gnd.t227 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X406 a_n2408_n452.t16 a_n2408_n452.t15 a_n1808_13878.t0 vdd.t46 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X407 vdd.t57 vdd.t54 vdd.t56 vdd.t55 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
R0 plus.n53 plus.t20 323.478
R1 plus.n11 plus.t15 323.478
R2 plus.n52 plus.t19 297.12
R3 plus.n56 plus.t26 297.12
R4 plus.n58 plus.t25 297.12
R5 plus.n62 plus.t27 297.12
R6 plus.n64 plus.t9 297.12
R7 plus.n68 plus.t7 297.12
R8 plus.n70 plus.t14 297.12
R9 plus.n74 plus.t12 297.12
R10 plus.n76 plus.t28 297.12
R11 plus.n80 plus.t10 297.12
R12 plus.n82 plus.t8 297.12
R13 plus.n40 plus.t21 297.12
R14 plus.n38 plus.t22 297.12
R15 plus.n2 plus.t16 297.12
R16 plus.n32 plus.t17 297.12
R17 plus.n4 plus.t11 297.12
R18 plus.n26 plus.t5 297.12
R19 plus.n6 plus.t6 297.12
R20 plus.n20 plus.t23 297.12
R21 plus.n8 plus.t24 297.12
R22 plus.n14 plus.t18 297.12
R23 plus.n10 plus.t13 297.12
R24 plus.n86 plus.t2 243.97
R25 plus.n86 plus.n85 223.454
R26 plus.n88 plus.n87 223.454
R27 plus.n83 plus.n82 161.3
R28 plus.n81 plus.n42 161.3
R29 plus.n80 plus.n79 161.3
R30 plus.n78 plus.n43 161.3
R31 plus.n77 plus.n76 161.3
R32 plus.n75 plus.n44 161.3
R33 plus.n74 plus.n73 161.3
R34 plus.n72 plus.n45 161.3
R35 plus.n71 plus.n70 161.3
R36 plus.n69 plus.n46 161.3
R37 plus.n68 plus.n67 161.3
R38 plus.n66 plus.n47 161.3
R39 plus.n65 plus.n64 161.3
R40 plus.n63 plus.n48 161.3
R41 plus.n62 plus.n61 161.3
R42 plus.n60 plus.n49 161.3
R43 plus.n59 plus.n58 161.3
R44 plus.n57 plus.n50 161.3
R45 plus.n56 plus.n55 161.3
R46 plus.n54 plus.n51 161.3
R47 plus.n13 plus.n12 161.3
R48 plus.n14 plus.n9 161.3
R49 plus.n16 plus.n15 161.3
R50 plus.n17 plus.n8 161.3
R51 plus.n19 plus.n18 161.3
R52 plus.n20 plus.n7 161.3
R53 plus.n22 plus.n21 161.3
R54 plus.n23 plus.n6 161.3
R55 plus.n25 plus.n24 161.3
R56 plus.n26 plus.n5 161.3
R57 plus.n28 plus.n27 161.3
R58 plus.n29 plus.n4 161.3
R59 plus.n31 plus.n30 161.3
R60 plus.n32 plus.n3 161.3
R61 plus.n34 plus.n33 161.3
R62 plus.n35 plus.n2 161.3
R63 plus.n37 plus.n36 161.3
R64 plus.n38 plus.n1 161.3
R65 plus.n39 plus.n0 161.3
R66 plus.n41 plus.n40 161.3
R67 plus.n82 plus.n81 46.0096
R68 plus.n40 plus.n39 46.0096
R69 plus.n54 plus.n53 45.0871
R70 plus.n12 plus.n11 45.0871
R71 plus.n52 plus.n51 41.6278
R72 plus.n80 plus.n43 41.6278
R73 plus.n38 plus.n37 41.6278
R74 plus.n13 plus.n10 41.6278
R75 plus.n57 plus.n56 37.246
R76 plus.n76 plus.n75 37.246
R77 plus.n33 plus.n2 37.246
R78 plus.n15 plus.n14 37.246
R79 plus.n84 plus.n83 33.1766
R80 plus.n58 plus.n49 32.8641
R81 plus.n74 plus.n45 32.8641
R82 plus.n32 plus.n31 32.8641
R83 plus.n19 plus.n8 32.8641
R84 plus.n63 plus.n62 28.4823
R85 plus.n70 plus.n69 28.4823
R86 plus.n27 plus.n4 28.4823
R87 plus.n21 plus.n20 28.4823
R88 plus.n64 plus.n47 24.1005
R89 plus.n68 plus.n47 24.1005
R90 plus.n26 plus.n25 24.1005
R91 plus.n25 plus.n6 24.1005
R92 plus.n85 plus.t0 19.8005
R93 plus.n85 plus.t3 19.8005
R94 plus.n87 plus.t1 19.8005
R95 plus.n87 plus.t4 19.8005
R96 plus.n64 plus.n63 19.7187
R97 plus.n69 plus.n68 19.7187
R98 plus.n27 plus.n26 19.7187
R99 plus.n21 plus.n6 19.7187
R100 plus.n62 plus.n49 15.3369
R101 plus.n70 plus.n45 15.3369
R102 plus.n31 plus.n4 15.3369
R103 plus.n20 plus.n19 15.3369
R104 plus plus.n89 14.2409
R105 plus.n53 plus.n52 14.1472
R106 plus.n11 plus.n10 14.1472
R107 plus.n84 plus.n41 11.8774
R108 plus.n58 plus.n57 10.955
R109 plus.n75 plus.n74 10.955
R110 plus.n33 plus.n32 10.955
R111 plus.n15 plus.n8 10.955
R112 plus.n56 plus.n51 6.57323
R113 plus.n76 plus.n43 6.57323
R114 plus.n37 plus.n2 6.57323
R115 plus.n14 plus.n13 6.57323
R116 plus.n89 plus.n88 5.40567
R117 plus.n81 plus.n80 2.19141
R118 plus.n39 plus.n38 2.19141
R119 plus.n89 plus.n84 1.188
R120 plus.n88 plus.n86 0.716017
R121 plus.n55 plus.n54 0.189894
R122 plus.n55 plus.n50 0.189894
R123 plus.n59 plus.n50 0.189894
R124 plus.n60 plus.n59 0.189894
R125 plus.n61 plus.n60 0.189894
R126 plus.n61 plus.n48 0.189894
R127 plus.n65 plus.n48 0.189894
R128 plus.n66 plus.n65 0.189894
R129 plus.n67 plus.n66 0.189894
R130 plus.n67 plus.n46 0.189894
R131 plus.n71 plus.n46 0.189894
R132 plus.n72 plus.n71 0.189894
R133 plus.n73 plus.n72 0.189894
R134 plus.n73 plus.n44 0.189894
R135 plus.n77 plus.n44 0.189894
R136 plus.n78 plus.n77 0.189894
R137 plus.n79 plus.n78 0.189894
R138 plus.n79 plus.n42 0.189894
R139 plus.n83 plus.n42 0.189894
R140 plus.n41 plus.n0 0.189894
R141 plus.n1 plus.n0 0.189894
R142 plus.n36 plus.n1 0.189894
R143 plus.n36 plus.n35 0.189894
R144 plus.n35 plus.n34 0.189894
R145 plus.n34 plus.n3 0.189894
R146 plus.n30 plus.n3 0.189894
R147 plus.n30 plus.n29 0.189894
R148 plus.n29 plus.n28 0.189894
R149 plus.n28 plus.n5 0.189894
R150 plus.n24 plus.n5 0.189894
R151 plus.n24 plus.n23 0.189894
R152 plus.n23 plus.n22 0.189894
R153 plus.n22 plus.n7 0.189894
R154 plus.n18 plus.n7 0.189894
R155 plus.n18 plus.n17 0.189894
R156 plus.n17 plus.n16 0.189894
R157 plus.n16 plus.n9 0.189894
R158 plus.n12 plus.n9 0.189894
R159 a_n2903_n3924.n11 a_n2903_n3924.t21 214.643
R160 a_n2903_n3924.n7 a_n2903_n3924.t11 214.321
R161 a_n2903_n3924.n7 a_n2903_n3924.t55 214.321
R162 a_n2903_n3924.n5 a_n2903_n3924.t9 214.321
R163 a_n2903_n3924.n5 a_n2903_n3924.t18 214.321
R164 a_n2903_n3924.n6 a_n2903_n3924.t10 214.321
R165 a_n2903_n3924.n6 a_n2903_n3924.t12 214.321
R166 a_n2903_n3924.n11 a_n2903_n3924.t48 214.321
R167 a_n2903_n3924.n1 a_n2903_n3924.t36 55.8337
R168 a_n2903_n3924.n1 a_n2903_n3924.t16 55.8337
R169 a_n2903_n3924.n10 a_n2903_n3924.t52 55.8337
R170 a_n2903_n3924.n0 a_n2903_n3924.t37 55.8335
R171 a_n2903_n3924.n8 a_n2903_n3924.t7 55.8335
R172 a_n2903_n3924.n4 a_n2903_n3924.t20 55.8335
R173 a_n2903_n3924.n4 a_n2903_n3924.t38 55.8335
R174 a_n2903_n3924.n3 a_n2903_n3924.t46 55.8335
R175 a_n2903_n3924.n0 a_n2903_n3924.n28 53.0052
R176 a_n2903_n3924.n0 a_n2903_n3924.n29 53.0052
R177 a_n2903_n3924.n0 a_n2903_n3924.n30 53.0052
R178 a_n2903_n3924.n1 a_n2903_n3924.n31 53.0052
R179 a_n2903_n3924.n1 a_n2903_n3924.n32 53.0052
R180 a_n2903_n3924.n1 a_n2903_n3924.n12 53.0052
R181 a_n2903_n3924.n9 a_n2903_n3924.n13 53.0052
R182 a_n2903_n3924.n9 a_n2903_n3924.n14 53.0052
R183 a_n2903_n3924.n10 a_n2903_n3924.n15 53.0052
R184 a_n2903_n3924.n8 a_n2903_n3924.n26 53.0051
R185 a_n2903_n3924.n2 a_n2903_n3924.n25 53.0051
R186 a_n2903_n3924.n2 a_n2903_n3924.n24 53.0051
R187 a_n2903_n3924.n2 a_n2903_n3924.n23 53.0051
R188 a_n2903_n3924.n2 a_n2903_n3924.n22 53.0051
R189 a_n2903_n3924.n4 a_n2903_n3924.n21 53.0051
R190 a_n2903_n3924.n4 a_n2903_n3924.n20 53.0051
R191 a_n2903_n3924.n4 a_n2903_n3924.n19 53.0051
R192 a_n2903_n3924.n3 a_n2903_n3924.n18 53.0051
R193 a_n2903_n3924.n3 a_n2903_n3924.n17 53.0051
R194 a_n2903_n3924.n33 a_n2903_n3924.n1 53.0051
R195 a_n2903_n3924.n16 a_n2903_n3924.n10 12.1986
R196 a_n2903_n3924.n0 a_n2903_n3924.n27 12.1986
R197 a_n2903_n3924.n3 a_n2903_n3924.n16 5.11903
R198 a_n2903_n3924.n27 a_n2903_n3924.n8 5.11903
R199 a_n2903_n3924.n28 a_n2903_n3924.t43 2.82907
R200 a_n2903_n3924.n28 a_n2903_n3924.t26 2.82907
R201 a_n2903_n3924.n29 a_n2903_n3924.t29 2.82907
R202 a_n2903_n3924.n29 a_n2903_n3924.t34 2.82907
R203 a_n2903_n3924.n30 a_n2903_n3924.t39 2.82907
R204 a_n2903_n3924.n30 a_n2903_n3924.t28 2.82907
R205 a_n2903_n3924.n31 a_n2903_n3924.t42 2.82907
R206 a_n2903_n3924.n31 a_n2903_n3924.t45 2.82907
R207 a_n2903_n3924.n32 a_n2903_n3924.t25 2.82907
R208 a_n2903_n3924.n32 a_n2903_n3924.t44 2.82907
R209 a_n2903_n3924.n12 a_n2903_n3924.t13 2.82907
R210 a_n2903_n3924.n12 a_n2903_n3924.t51 2.82907
R211 a_n2903_n3924.n13 a_n2903_n3924.t50 2.82907
R212 a_n2903_n3924.n13 a_n2903_n3924.t22 2.82907
R213 a_n2903_n3924.n14 a_n2903_n3924.t49 2.82907
R214 a_n2903_n3924.n14 a_n2903_n3924.t17 2.82907
R215 a_n2903_n3924.n15 a_n2903_n3924.t3 2.82907
R216 a_n2903_n3924.n15 a_n2903_n3924.t14 2.82907
R217 a_n2903_n3924.n26 a_n2903_n3924.t19 2.82907
R218 a_n2903_n3924.n26 a_n2903_n3924.t53 2.82907
R219 a_n2903_n3924.n25 a_n2903_n3924.t4 2.82907
R220 a_n2903_n3924.n25 a_n2903_n3924.t6 2.82907
R221 a_n2903_n3924.n24 a_n2903_n3924.t1 2.82907
R222 a_n2903_n3924.n24 a_n2903_n3924.t5 2.82907
R223 a_n2903_n3924.n23 a_n2903_n3924.t8 2.82907
R224 a_n2903_n3924.n23 a_n2903_n3924.t2 2.82907
R225 a_n2903_n3924.n22 a_n2903_n3924.t15 2.82907
R226 a_n2903_n3924.n22 a_n2903_n3924.t47 2.82907
R227 a_n2903_n3924.n21 a_n2903_n3924.t30 2.82907
R228 a_n2903_n3924.n21 a_n2903_n3924.t27 2.82907
R229 a_n2903_n3924.n20 a_n2903_n3924.t31 2.82907
R230 a_n2903_n3924.n20 a_n2903_n3924.t23 2.82907
R231 a_n2903_n3924.n19 a_n2903_n3924.t40 2.82907
R232 a_n2903_n3924.n19 a_n2903_n3924.t33 2.82907
R233 a_n2903_n3924.n18 a_n2903_n3924.t41 2.82907
R234 a_n2903_n3924.n18 a_n2903_n3924.t24 2.82907
R235 a_n2903_n3924.n17 a_n2903_n3924.t32 2.82907
R236 a_n2903_n3924.n17 a_n2903_n3924.t35 2.82907
R237 a_n2903_n3924.n33 a_n2903_n3924.t54 2.82907
R238 a_n2903_n3924.t0 a_n2903_n3924.n33 2.82907
R239 a_n2903_n3924.n1 a_n2903_n3924.n0 2.66429
R240 a_n2903_n3924.n27 a_n2903_n3924.n7 2.16406
R241 a_n2903_n3924.n2 a_n2903_n3924.n4 2.01128
R242 a_n2903_n3924.n16 a_n2903_n3924.n11 1.95694
R243 a_n2903_n3924.n4 a_n2903_n3924.n3 1.77636
R244 a_n2903_n3924.n8 a_n2903_n3924.n2 1.77636
R245 a_n2903_n3924.n11 a_n2903_n3924.n6 1.69309
R246 a_n2903_n3924.n9 a_n2903_n3924.n1 1.56731
R247 a_n2903_n3924.n5 a_n2903_n3924.n7 1.34352
R248 a_n2903_n3924.n6 a_n2903_n3924.n5 1.34352
R249 a_n2903_n3924.n10 a_n2903_n3924.n9 1.3324
R250 a_n7636_8799.n219 a_n7636_8799.t64 485.149
R251 a_n7636_8799.n281 a_n7636_8799.t76 485.149
R252 a_n7636_8799.n344 a_n7636_8799.t113 485.149
R253 a_n7636_8799.n29 a_n7636_8799.t135 485.149
R254 a_n7636_8799.n91 a_n7636_8799.t150 485.149
R255 a_n7636_8799.n154 a_n7636_8799.t112 485.149
R256 a_n7636_8799.n262 a_n7636_8799.t86 464.166
R257 a_n7636_8799.n261 a_n7636_8799.t85 464.166
R258 a_n7636_8799.n203 a_n7636_8799.t58 464.166
R259 a_n7636_8799.n255 a_n7636_8799.t134 464.166
R260 a_n7636_8799.n254 a_n7636_8799.t89 464.166
R261 a_n7636_8799.n206 a_n7636_8799.t65 464.166
R262 a_n7636_8799.n248 a_n7636_8799.t140 464.166
R263 a_n7636_8799.n247 a_n7636_8799.t106 464.166
R264 a_n7636_8799.n209 a_n7636_8799.t104 464.166
R265 a_n7636_8799.n241 a_n7636_8799.t39 464.166
R266 a_n7636_8799.n240 a_n7636_8799.t110 464.166
R267 a_n7636_8799.n212 a_n7636_8799.t109 464.166
R268 a_n7636_8799.n234 a_n7636_8799.t41 464.166
R269 a_n7636_8799.n233 a_n7636_8799.t40 464.166
R270 a_n7636_8799.n215 a_n7636_8799.t126 464.166
R271 a_n7636_8799.n227 a_n7636_8799.t60 464.166
R272 a_n7636_8799.n226 a_n7636_8799.t44 464.166
R273 a_n7636_8799.n218 a_n7636_8799.t130 464.166
R274 a_n7636_8799.n220 a_n7636_8799.t88 464.166
R275 a_n7636_8799.n324 a_n7636_8799.t96 464.166
R276 a_n7636_8799.n323 a_n7636_8799.t95 464.166
R277 a_n7636_8799.n265 a_n7636_8799.t73 464.166
R278 a_n7636_8799.n317 a_n7636_8799.t149 464.166
R279 a_n7636_8799.n316 a_n7636_8799.t102 464.166
R280 a_n7636_8799.n268 a_n7636_8799.t75 464.166
R281 a_n7636_8799.n310 a_n7636_8799.t155 464.166
R282 a_n7636_8799.n309 a_n7636_8799.t119 464.166
R283 a_n7636_8799.n271 a_n7636_8799.t118 464.166
R284 a_n7636_8799.n303 a_n7636_8799.t49 464.166
R285 a_n7636_8799.n302 a_n7636_8799.t122 464.166
R286 a_n7636_8799.n274 a_n7636_8799.t121 464.166
R287 a_n7636_8799.n296 a_n7636_8799.t53 464.166
R288 a_n7636_8799.n295 a_n7636_8799.t52 464.166
R289 a_n7636_8799.n277 a_n7636_8799.t143 464.166
R290 a_n7636_8799.n289 a_n7636_8799.t74 464.166
R291 a_n7636_8799.n288 a_n7636_8799.t56 464.166
R292 a_n7636_8799.n280 a_n7636_8799.t144 464.166
R293 a_n7636_8799.n282 a_n7636_8799.t103 464.166
R294 a_n7636_8799.n387 a_n7636_8799.t154 464.166
R295 a_n7636_8799.n386 a_n7636_8799.t51 464.166
R296 a_n7636_8799.n328 a_n7636_8799.t101 464.166
R297 a_n7636_8799.n380 a_n7636_8799.t38 464.166
R298 a_n7636_8799.n379 a_n7636_8799.t125 464.166
R299 a_n7636_8799.n331 a_n7636_8799.t62 464.166
R300 a_n7636_8799.n373 a_n7636_8799.t108 464.166
R301 a_n7636_8799.n372 a_n7636_8799.t43 464.166
R302 a_n7636_8799.n334 a_n7636_8799.t68 464.166
R303 a_n7636_8799.n366 a_n7636_8799.t148 464.166
R304 a_n7636_8799.n365 a_n7636_8799.t117 464.166
R305 a_n7636_8799.n337 a_n7636_8799.t142 464.166
R306 a_n7636_8799.n359 a_n7636_8799.t99 464.166
R307 a_n7636_8799.n358 a_n7636_8799.t120 464.166
R308 a_n7636_8799.n340 a_n7636_8799.t55 464.166
R309 a_n7636_8799.n352 a_n7636_8799.t139 464.166
R310 a_n7636_8799.n351 a_n7636_8799.t80 464.166
R311 a_n7636_8799.n343 a_n7636_8799.t131 464.166
R312 a_n7636_8799.n345 a_n7636_8799.t67 464.166
R313 a_n7636_8799.n30 a_n7636_8799.t137 464.166
R314 a_n7636_8799.n32 a_n7636_8799.t87 464.166
R315 a_n7636_8799.n36 a_n7636_8799.t116 464.166
R316 a_n7636_8799.n37 a_n7636_8799.t133 464.166
R317 a_n7636_8799.n25 a_n7636_8799.t83 464.166
R318 a_n7636_8799.n43 a_n7636_8799.t84 464.166
R319 a_n7636_8799.n44 a_n7636_8799.t114 464.166
R320 a_n7636_8799.n48 a_n7636_8799.t71 464.166
R321 a_n7636_8799.n50 a_n7636_8799.t72 464.166
R322 a_n7636_8799.n21 a_n7636_8799.t111 464.166
R323 a_n7636_8799.n55 a_n7636_8799.t36 464.166
R324 a_n7636_8799.n19 a_n7636_8799.t69 464.166
R325 a_n7636_8799.n60 a_n7636_8799.t92 464.166
R326 a_n7636_8799.n62 a_n7636_8799.t136 464.166
R327 a_n7636_8799.n66 a_n7636_8799.t48 464.166
R328 a_n7636_8799.n67 a_n7636_8799.t66 464.166
R329 a_n7636_8799.n15 a_n7636_8799.t132 464.166
R330 a_n7636_8799.n73 a_n7636_8799.t45 464.166
R331 a_n7636_8799.n74 a_n7636_8799.t46 464.166
R332 a_n7636_8799.n92 a_n7636_8799.t153 464.166
R333 a_n7636_8799.n94 a_n7636_8799.t97 464.166
R334 a_n7636_8799.n98 a_n7636_8799.t129 464.166
R335 a_n7636_8799.n99 a_n7636_8799.t147 464.166
R336 a_n7636_8799.n87 a_n7636_8799.t93 464.166
R337 a_n7636_8799.n105 a_n7636_8799.t94 464.166
R338 a_n7636_8799.n106 a_n7636_8799.t127 464.166
R339 a_n7636_8799.n110 a_n7636_8799.t81 464.166
R340 a_n7636_8799.n112 a_n7636_8799.t82 464.166
R341 a_n7636_8799.n83 a_n7636_8799.t123 464.166
R342 a_n7636_8799.n117 a_n7636_8799.t47 464.166
R343 a_n7636_8799.n81 a_n7636_8799.t78 464.166
R344 a_n7636_8799.n122 a_n7636_8799.t105 464.166
R345 a_n7636_8799.n124 a_n7636_8799.t151 464.166
R346 a_n7636_8799.n128 a_n7636_8799.t63 464.166
R347 a_n7636_8799.n129 a_n7636_8799.t77 464.166
R348 a_n7636_8799.n77 a_n7636_8799.t145 464.166
R349 a_n7636_8799.n135 a_n7636_8799.t57 464.166
R350 a_n7636_8799.n136 a_n7636_8799.t59 464.166
R351 a_n7636_8799.n155 a_n7636_8799.t90 464.166
R352 a_n7636_8799.n157 a_n7636_8799.t128 464.166
R353 a_n7636_8799.n161 a_n7636_8799.t79 464.166
R354 a_n7636_8799.n162 a_n7636_8799.t138 464.166
R355 a_n7636_8799.n150 a_n7636_8799.t54 464.166
R356 a_n7636_8799.n168 a_n7636_8799.t37 464.166
R357 a_n7636_8799.n169 a_n7636_8799.t98 464.166
R358 a_n7636_8799.n173 a_n7636_8799.t141 464.166
R359 a_n7636_8799.n175 a_n7636_8799.t115 464.166
R360 a_n7636_8799.n146 a_n7636_8799.t146 464.166
R361 a_n7636_8799.n180 a_n7636_8799.t91 464.166
R362 a_n7636_8799.n144 a_n7636_8799.t42 464.166
R363 a_n7636_8799.n185 a_n7636_8799.t107 464.166
R364 a_n7636_8799.n187 a_n7636_8799.t61 464.166
R365 a_n7636_8799.n191 a_n7636_8799.t124 464.166
R366 a_n7636_8799.n192 a_n7636_8799.t70 464.166
R367 a_n7636_8799.n140 a_n7636_8799.t100 464.166
R368 a_n7636_8799.n198 a_n7636_8799.t50 464.166
R369 a_n7636_8799.n199 a_n7636_8799.t152 464.166
R370 a_n7636_8799.n222 a_n7636_8799.n221 161.3
R371 a_n7636_8799.n223 a_n7636_8799.n218 161.3
R372 a_n7636_8799.n225 a_n7636_8799.n224 161.3
R373 a_n7636_8799.n226 a_n7636_8799.n217 161.3
R374 a_n7636_8799.n227 a_n7636_8799.n216 161.3
R375 a_n7636_8799.n229 a_n7636_8799.n228 161.3
R376 a_n7636_8799.n230 a_n7636_8799.n215 161.3
R377 a_n7636_8799.n232 a_n7636_8799.n231 161.3
R378 a_n7636_8799.n233 a_n7636_8799.n214 161.3
R379 a_n7636_8799.n234 a_n7636_8799.n213 161.3
R380 a_n7636_8799.n236 a_n7636_8799.n235 161.3
R381 a_n7636_8799.n237 a_n7636_8799.n212 161.3
R382 a_n7636_8799.n239 a_n7636_8799.n238 161.3
R383 a_n7636_8799.n240 a_n7636_8799.n211 161.3
R384 a_n7636_8799.n241 a_n7636_8799.n210 161.3
R385 a_n7636_8799.n243 a_n7636_8799.n242 161.3
R386 a_n7636_8799.n244 a_n7636_8799.n209 161.3
R387 a_n7636_8799.n246 a_n7636_8799.n245 161.3
R388 a_n7636_8799.n247 a_n7636_8799.n208 161.3
R389 a_n7636_8799.n248 a_n7636_8799.n207 161.3
R390 a_n7636_8799.n250 a_n7636_8799.n249 161.3
R391 a_n7636_8799.n251 a_n7636_8799.n206 161.3
R392 a_n7636_8799.n253 a_n7636_8799.n252 161.3
R393 a_n7636_8799.n254 a_n7636_8799.n205 161.3
R394 a_n7636_8799.n255 a_n7636_8799.n204 161.3
R395 a_n7636_8799.n257 a_n7636_8799.n256 161.3
R396 a_n7636_8799.n258 a_n7636_8799.n203 161.3
R397 a_n7636_8799.n260 a_n7636_8799.n259 161.3
R398 a_n7636_8799.n261 a_n7636_8799.n202 161.3
R399 a_n7636_8799.n263 a_n7636_8799.n262 161.3
R400 a_n7636_8799.n284 a_n7636_8799.n283 161.3
R401 a_n7636_8799.n285 a_n7636_8799.n280 161.3
R402 a_n7636_8799.n287 a_n7636_8799.n286 161.3
R403 a_n7636_8799.n288 a_n7636_8799.n279 161.3
R404 a_n7636_8799.n289 a_n7636_8799.n278 161.3
R405 a_n7636_8799.n291 a_n7636_8799.n290 161.3
R406 a_n7636_8799.n292 a_n7636_8799.n277 161.3
R407 a_n7636_8799.n294 a_n7636_8799.n293 161.3
R408 a_n7636_8799.n295 a_n7636_8799.n276 161.3
R409 a_n7636_8799.n296 a_n7636_8799.n275 161.3
R410 a_n7636_8799.n298 a_n7636_8799.n297 161.3
R411 a_n7636_8799.n299 a_n7636_8799.n274 161.3
R412 a_n7636_8799.n301 a_n7636_8799.n300 161.3
R413 a_n7636_8799.n302 a_n7636_8799.n273 161.3
R414 a_n7636_8799.n303 a_n7636_8799.n272 161.3
R415 a_n7636_8799.n305 a_n7636_8799.n304 161.3
R416 a_n7636_8799.n306 a_n7636_8799.n271 161.3
R417 a_n7636_8799.n308 a_n7636_8799.n307 161.3
R418 a_n7636_8799.n309 a_n7636_8799.n270 161.3
R419 a_n7636_8799.n310 a_n7636_8799.n269 161.3
R420 a_n7636_8799.n312 a_n7636_8799.n311 161.3
R421 a_n7636_8799.n313 a_n7636_8799.n268 161.3
R422 a_n7636_8799.n315 a_n7636_8799.n314 161.3
R423 a_n7636_8799.n316 a_n7636_8799.n267 161.3
R424 a_n7636_8799.n317 a_n7636_8799.n266 161.3
R425 a_n7636_8799.n319 a_n7636_8799.n318 161.3
R426 a_n7636_8799.n320 a_n7636_8799.n265 161.3
R427 a_n7636_8799.n322 a_n7636_8799.n321 161.3
R428 a_n7636_8799.n323 a_n7636_8799.n264 161.3
R429 a_n7636_8799.n325 a_n7636_8799.n324 161.3
R430 a_n7636_8799.n347 a_n7636_8799.n346 161.3
R431 a_n7636_8799.n348 a_n7636_8799.n343 161.3
R432 a_n7636_8799.n350 a_n7636_8799.n349 161.3
R433 a_n7636_8799.n351 a_n7636_8799.n342 161.3
R434 a_n7636_8799.n352 a_n7636_8799.n341 161.3
R435 a_n7636_8799.n354 a_n7636_8799.n353 161.3
R436 a_n7636_8799.n355 a_n7636_8799.n340 161.3
R437 a_n7636_8799.n357 a_n7636_8799.n356 161.3
R438 a_n7636_8799.n358 a_n7636_8799.n339 161.3
R439 a_n7636_8799.n359 a_n7636_8799.n338 161.3
R440 a_n7636_8799.n361 a_n7636_8799.n360 161.3
R441 a_n7636_8799.n362 a_n7636_8799.n337 161.3
R442 a_n7636_8799.n364 a_n7636_8799.n363 161.3
R443 a_n7636_8799.n365 a_n7636_8799.n336 161.3
R444 a_n7636_8799.n366 a_n7636_8799.n335 161.3
R445 a_n7636_8799.n368 a_n7636_8799.n367 161.3
R446 a_n7636_8799.n369 a_n7636_8799.n334 161.3
R447 a_n7636_8799.n371 a_n7636_8799.n370 161.3
R448 a_n7636_8799.n372 a_n7636_8799.n333 161.3
R449 a_n7636_8799.n373 a_n7636_8799.n332 161.3
R450 a_n7636_8799.n375 a_n7636_8799.n374 161.3
R451 a_n7636_8799.n376 a_n7636_8799.n331 161.3
R452 a_n7636_8799.n378 a_n7636_8799.n377 161.3
R453 a_n7636_8799.n379 a_n7636_8799.n330 161.3
R454 a_n7636_8799.n380 a_n7636_8799.n329 161.3
R455 a_n7636_8799.n382 a_n7636_8799.n381 161.3
R456 a_n7636_8799.n383 a_n7636_8799.n328 161.3
R457 a_n7636_8799.n385 a_n7636_8799.n384 161.3
R458 a_n7636_8799.n386 a_n7636_8799.n327 161.3
R459 a_n7636_8799.n388 a_n7636_8799.n387 161.3
R460 a_n7636_8799.n75 a_n7636_8799.n74 161.3
R461 a_n7636_8799.n73 a_n7636_8799.n14 161.3
R462 a_n7636_8799.n72 a_n7636_8799.n71 161.3
R463 a_n7636_8799.n70 a_n7636_8799.n15 161.3
R464 a_n7636_8799.n69 a_n7636_8799.n68 161.3
R465 a_n7636_8799.n67 a_n7636_8799.n16 161.3
R466 a_n7636_8799.n66 a_n7636_8799.n65 161.3
R467 a_n7636_8799.n64 a_n7636_8799.n17 161.3
R468 a_n7636_8799.n63 a_n7636_8799.n62 161.3
R469 a_n7636_8799.n61 a_n7636_8799.n18 161.3
R470 a_n7636_8799.n60 a_n7636_8799.n59 161.3
R471 a_n7636_8799.n58 a_n7636_8799.n19 161.3
R472 a_n7636_8799.n57 a_n7636_8799.n56 161.3
R473 a_n7636_8799.n55 a_n7636_8799.n20 161.3
R474 a_n7636_8799.n54 a_n7636_8799.n53 161.3
R475 a_n7636_8799.n52 a_n7636_8799.n21 161.3
R476 a_n7636_8799.n51 a_n7636_8799.n50 161.3
R477 a_n7636_8799.n49 a_n7636_8799.n22 161.3
R478 a_n7636_8799.n48 a_n7636_8799.n47 161.3
R479 a_n7636_8799.n46 a_n7636_8799.n23 161.3
R480 a_n7636_8799.n45 a_n7636_8799.n44 161.3
R481 a_n7636_8799.n43 a_n7636_8799.n24 161.3
R482 a_n7636_8799.n42 a_n7636_8799.n41 161.3
R483 a_n7636_8799.n40 a_n7636_8799.n25 161.3
R484 a_n7636_8799.n39 a_n7636_8799.n38 161.3
R485 a_n7636_8799.n37 a_n7636_8799.n26 161.3
R486 a_n7636_8799.n36 a_n7636_8799.n35 161.3
R487 a_n7636_8799.n34 a_n7636_8799.n27 161.3
R488 a_n7636_8799.n33 a_n7636_8799.n32 161.3
R489 a_n7636_8799.n31 a_n7636_8799.n28 161.3
R490 a_n7636_8799.n137 a_n7636_8799.n136 161.3
R491 a_n7636_8799.n135 a_n7636_8799.n76 161.3
R492 a_n7636_8799.n134 a_n7636_8799.n133 161.3
R493 a_n7636_8799.n132 a_n7636_8799.n77 161.3
R494 a_n7636_8799.n131 a_n7636_8799.n130 161.3
R495 a_n7636_8799.n129 a_n7636_8799.n78 161.3
R496 a_n7636_8799.n128 a_n7636_8799.n127 161.3
R497 a_n7636_8799.n126 a_n7636_8799.n79 161.3
R498 a_n7636_8799.n125 a_n7636_8799.n124 161.3
R499 a_n7636_8799.n123 a_n7636_8799.n80 161.3
R500 a_n7636_8799.n122 a_n7636_8799.n121 161.3
R501 a_n7636_8799.n120 a_n7636_8799.n81 161.3
R502 a_n7636_8799.n119 a_n7636_8799.n118 161.3
R503 a_n7636_8799.n117 a_n7636_8799.n82 161.3
R504 a_n7636_8799.n116 a_n7636_8799.n115 161.3
R505 a_n7636_8799.n114 a_n7636_8799.n83 161.3
R506 a_n7636_8799.n113 a_n7636_8799.n112 161.3
R507 a_n7636_8799.n111 a_n7636_8799.n84 161.3
R508 a_n7636_8799.n110 a_n7636_8799.n109 161.3
R509 a_n7636_8799.n108 a_n7636_8799.n85 161.3
R510 a_n7636_8799.n107 a_n7636_8799.n106 161.3
R511 a_n7636_8799.n105 a_n7636_8799.n86 161.3
R512 a_n7636_8799.n104 a_n7636_8799.n103 161.3
R513 a_n7636_8799.n102 a_n7636_8799.n87 161.3
R514 a_n7636_8799.n101 a_n7636_8799.n100 161.3
R515 a_n7636_8799.n99 a_n7636_8799.n88 161.3
R516 a_n7636_8799.n98 a_n7636_8799.n97 161.3
R517 a_n7636_8799.n96 a_n7636_8799.n89 161.3
R518 a_n7636_8799.n95 a_n7636_8799.n94 161.3
R519 a_n7636_8799.n93 a_n7636_8799.n90 161.3
R520 a_n7636_8799.n200 a_n7636_8799.n199 161.3
R521 a_n7636_8799.n198 a_n7636_8799.n139 161.3
R522 a_n7636_8799.n197 a_n7636_8799.n196 161.3
R523 a_n7636_8799.n195 a_n7636_8799.n140 161.3
R524 a_n7636_8799.n194 a_n7636_8799.n193 161.3
R525 a_n7636_8799.n192 a_n7636_8799.n141 161.3
R526 a_n7636_8799.n191 a_n7636_8799.n190 161.3
R527 a_n7636_8799.n189 a_n7636_8799.n142 161.3
R528 a_n7636_8799.n188 a_n7636_8799.n187 161.3
R529 a_n7636_8799.n186 a_n7636_8799.n143 161.3
R530 a_n7636_8799.n185 a_n7636_8799.n184 161.3
R531 a_n7636_8799.n183 a_n7636_8799.n144 161.3
R532 a_n7636_8799.n182 a_n7636_8799.n181 161.3
R533 a_n7636_8799.n180 a_n7636_8799.n145 161.3
R534 a_n7636_8799.n179 a_n7636_8799.n178 161.3
R535 a_n7636_8799.n177 a_n7636_8799.n146 161.3
R536 a_n7636_8799.n176 a_n7636_8799.n175 161.3
R537 a_n7636_8799.n174 a_n7636_8799.n147 161.3
R538 a_n7636_8799.n173 a_n7636_8799.n172 161.3
R539 a_n7636_8799.n171 a_n7636_8799.n148 161.3
R540 a_n7636_8799.n170 a_n7636_8799.n169 161.3
R541 a_n7636_8799.n168 a_n7636_8799.n149 161.3
R542 a_n7636_8799.n167 a_n7636_8799.n166 161.3
R543 a_n7636_8799.n165 a_n7636_8799.n150 161.3
R544 a_n7636_8799.n164 a_n7636_8799.n163 161.3
R545 a_n7636_8799.n162 a_n7636_8799.n151 161.3
R546 a_n7636_8799.n161 a_n7636_8799.n160 161.3
R547 a_n7636_8799.n159 a_n7636_8799.n152 161.3
R548 a_n7636_8799.n158 a_n7636_8799.n157 161.3
R549 a_n7636_8799.n156 a_n7636_8799.n153 161.3
R550 a_n7636_8799.n10 a_n7636_8799.n8 98.9633
R551 a_n7636_8799.n5 a_n7636_8799.n3 98.9631
R552 a_n7636_8799.n12 a_n7636_8799.n11 98.6055
R553 a_n7636_8799.n10 a_n7636_8799.n9 98.6055
R554 a_n7636_8799.n5 a_n7636_8799.n4 98.6055
R555 a_n7636_8799.n7 a_n7636_8799.n6 98.6055
R556 a_n7636_8799.n394 a_n7636_8799.n392 81.3764
R557 a_n7636_8799.n406 a_n7636_8799.n404 81.3764
R558 a_n7636_8799.n2 a_n7636_8799.n0 81.3764
R559 a_n7636_8799.n411 a_n7636_8799.n410 80.9326
R560 a_n7636_8799.n403 a_n7636_8799.n402 80.9324
R561 a_n7636_8799.n401 a_n7636_8799.n400 80.9324
R562 a_n7636_8799.n399 a_n7636_8799.n398 80.9324
R563 a_n7636_8799.n396 a_n7636_8799.n395 80.9324
R564 a_n7636_8799.n394 a_n7636_8799.n393 80.9324
R565 a_n7636_8799.n406 a_n7636_8799.n405 80.9324
R566 a_n7636_8799.n408 a_n7636_8799.n407 80.9324
R567 a_n7636_8799.n2 a_n7636_8799.n1 80.9324
R568 a_n7636_8799.n222 a_n7636_8799.n219 70.4033
R569 a_n7636_8799.n284 a_n7636_8799.n281 70.4033
R570 a_n7636_8799.n347 a_n7636_8799.n344 70.4033
R571 a_n7636_8799.n29 a_n7636_8799.n28 70.4033
R572 a_n7636_8799.n91 a_n7636_8799.n90 70.4033
R573 a_n7636_8799.n154 a_n7636_8799.n153 70.4033
R574 a_n7636_8799.n262 a_n7636_8799.n261 48.2005
R575 a_n7636_8799.n255 a_n7636_8799.n254 48.2005
R576 a_n7636_8799.n248 a_n7636_8799.n247 48.2005
R577 a_n7636_8799.n241 a_n7636_8799.n240 48.2005
R578 a_n7636_8799.n234 a_n7636_8799.n233 48.2005
R579 a_n7636_8799.n227 a_n7636_8799.n226 48.2005
R580 a_n7636_8799.n324 a_n7636_8799.n323 48.2005
R581 a_n7636_8799.n317 a_n7636_8799.n316 48.2005
R582 a_n7636_8799.n310 a_n7636_8799.n309 48.2005
R583 a_n7636_8799.n303 a_n7636_8799.n302 48.2005
R584 a_n7636_8799.n296 a_n7636_8799.n295 48.2005
R585 a_n7636_8799.n289 a_n7636_8799.n288 48.2005
R586 a_n7636_8799.n387 a_n7636_8799.n386 48.2005
R587 a_n7636_8799.n380 a_n7636_8799.n379 48.2005
R588 a_n7636_8799.n373 a_n7636_8799.n372 48.2005
R589 a_n7636_8799.n366 a_n7636_8799.n365 48.2005
R590 a_n7636_8799.n359 a_n7636_8799.n358 48.2005
R591 a_n7636_8799.n352 a_n7636_8799.n351 48.2005
R592 a_n7636_8799.n37 a_n7636_8799.n36 48.2005
R593 a_n7636_8799.n44 a_n7636_8799.n43 48.2005
R594 a_n7636_8799.n50 a_n7636_8799.n21 48.2005
R595 a_n7636_8799.n60 a_n7636_8799.n19 48.2005
R596 a_n7636_8799.n67 a_n7636_8799.n66 48.2005
R597 a_n7636_8799.n74 a_n7636_8799.n73 48.2005
R598 a_n7636_8799.n99 a_n7636_8799.n98 48.2005
R599 a_n7636_8799.n106 a_n7636_8799.n105 48.2005
R600 a_n7636_8799.n112 a_n7636_8799.n83 48.2005
R601 a_n7636_8799.n122 a_n7636_8799.n81 48.2005
R602 a_n7636_8799.n129 a_n7636_8799.n128 48.2005
R603 a_n7636_8799.n136 a_n7636_8799.n135 48.2005
R604 a_n7636_8799.n162 a_n7636_8799.n161 48.2005
R605 a_n7636_8799.n169 a_n7636_8799.n168 48.2005
R606 a_n7636_8799.n175 a_n7636_8799.n146 48.2005
R607 a_n7636_8799.n185 a_n7636_8799.n144 48.2005
R608 a_n7636_8799.n192 a_n7636_8799.n191 48.2005
R609 a_n7636_8799.n199 a_n7636_8799.n198 48.2005
R610 a_n7636_8799.n260 a_n7636_8799.n203 40.1672
R611 a_n7636_8799.n221 a_n7636_8799.n218 40.1672
R612 a_n7636_8799.n322 a_n7636_8799.n265 40.1672
R613 a_n7636_8799.n283 a_n7636_8799.n280 40.1672
R614 a_n7636_8799.n385 a_n7636_8799.n328 40.1672
R615 a_n7636_8799.n346 a_n7636_8799.n343 40.1672
R616 a_n7636_8799.n32 a_n7636_8799.n31 40.1672
R617 a_n7636_8799.n72 a_n7636_8799.n15 40.1672
R618 a_n7636_8799.n94 a_n7636_8799.n93 40.1672
R619 a_n7636_8799.n134 a_n7636_8799.n77 40.1672
R620 a_n7636_8799.n157 a_n7636_8799.n156 40.1672
R621 a_n7636_8799.n197 a_n7636_8799.n140 40.1672
R622 a_n7636_8799.n253 a_n7636_8799.n206 38.7066
R623 a_n7636_8799.n228 a_n7636_8799.n215 38.7066
R624 a_n7636_8799.n315 a_n7636_8799.n268 38.7066
R625 a_n7636_8799.n290 a_n7636_8799.n277 38.7066
R626 a_n7636_8799.n378 a_n7636_8799.n331 38.7066
R627 a_n7636_8799.n353 a_n7636_8799.n340 38.7066
R628 a_n7636_8799.n38 a_n7636_8799.n25 38.7066
R629 a_n7636_8799.n62 a_n7636_8799.n17 38.7066
R630 a_n7636_8799.n100 a_n7636_8799.n87 38.7066
R631 a_n7636_8799.n124 a_n7636_8799.n79 38.7066
R632 a_n7636_8799.n163 a_n7636_8799.n150 38.7066
R633 a_n7636_8799.n187 a_n7636_8799.n142 38.7066
R634 a_n7636_8799.n246 a_n7636_8799.n209 37.246
R635 a_n7636_8799.n235 a_n7636_8799.n212 37.246
R636 a_n7636_8799.n308 a_n7636_8799.n271 37.246
R637 a_n7636_8799.n297 a_n7636_8799.n274 37.246
R638 a_n7636_8799.n371 a_n7636_8799.n334 37.246
R639 a_n7636_8799.n360 a_n7636_8799.n337 37.246
R640 a_n7636_8799.n48 a_n7636_8799.n23 37.246
R641 a_n7636_8799.n56 a_n7636_8799.n55 37.246
R642 a_n7636_8799.n110 a_n7636_8799.n85 37.246
R643 a_n7636_8799.n118 a_n7636_8799.n117 37.246
R644 a_n7636_8799.n173 a_n7636_8799.n148 37.246
R645 a_n7636_8799.n181 a_n7636_8799.n180 37.246
R646 a_n7636_8799.n242 a_n7636_8799.n209 35.7853
R647 a_n7636_8799.n239 a_n7636_8799.n212 35.7853
R648 a_n7636_8799.n304 a_n7636_8799.n271 35.7853
R649 a_n7636_8799.n301 a_n7636_8799.n274 35.7853
R650 a_n7636_8799.n367 a_n7636_8799.n334 35.7853
R651 a_n7636_8799.n364 a_n7636_8799.n337 35.7853
R652 a_n7636_8799.n49 a_n7636_8799.n48 35.7853
R653 a_n7636_8799.n55 a_n7636_8799.n54 35.7853
R654 a_n7636_8799.n111 a_n7636_8799.n110 35.7853
R655 a_n7636_8799.n117 a_n7636_8799.n116 35.7853
R656 a_n7636_8799.n174 a_n7636_8799.n173 35.7853
R657 a_n7636_8799.n180 a_n7636_8799.n179 35.7853
R658 a_n7636_8799.n249 a_n7636_8799.n206 34.3247
R659 a_n7636_8799.n232 a_n7636_8799.n215 34.3247
R660 a_n7636_8799.n311 a_n7636_8799.n268 34.3247
R661 a_n7636_8799.n294 a_n7636_8799.n277 34.3247
R662 a_n7636_8799.n374 a_n7636_8799.n331 34.3247
R663 a_n7636_8799.n357 a_n7636_8799.n340 34.3247
R664 a_n7636_8799.n42 a_n7636_8799.n25 34.3247
R665 a_n7636_8799.n62 a_n7636_8799.n61 34.3247
R666 a_n7636_8799.n104 a_n7636_8799.n87 34.3247
R667 a_n7636_8799.n124 a_n7636_8799.n123 34.3247
R668 a_n7636_8799.n167 a_n7636_8799.n150 34.3247
R669 a_n7636_8799.n187 a_n7636_8799.n186 34.3247
R670 a_n7636_8799.n409 a_n7636_8799.n403 33.4185
R671 a_n7636_8799.n256 a_n7636_8799.n203 32.8641
R672 a_n7636_8799.n225 a_n7636_8799.n218 32.8641
R673 a_n7636_8799.n318 a_n7636_8799.n265 32.8641
R674 a_n7636_8799.n287 a_n7636_8799.n280 32.8641
R675 a_n7636_8799.n381 a_n7636_8799.n328 32.8641
R676 a_n7636_8799.n350 a_n7636_8799.n343 32.8641
R677 a_n7636_8799.n32 a_n7636_8799.n27 32.8641
R678 a_n7636_8799.n68 a_n7636_8799.n15 32.8641
R679 a_n7636_8799.n94 a_n7636_8799.n89 32.8641
R680 a_n7636_8799.n130 a_n7636_8799.n77 32.8641
R681 a_n7636_8799.n157 a_n7636_8799.n152 32.8641
R682 a_n7636_8799.n193 a_n7636_8799.n140 32.8641
R683 a_n7636_8799.n13 a_n7636_8799.n7 30.9355
R684 a_n7636_8799.n220 a_n7636_8799.n219 20.9576
R685 a_n7636_8799.n282 a_n7636_8799.n281 20.9576
R686 a_n7636_8799.n345 a_n7636_8799.n344 20.9576
R687 a_n7636_8799.n30 a_n7636_8799.n29 20.9576
R688 a_n7636_8799.n92 a_n7636_8799.n91 20.9576
R689 a_n7636_8799.n155 a_n7636_8799.n154 20.9576
R690 a_n7636_8799.n13 a_n7636_8799.n12 17.5141
R691 a_n7636_8799.n256 a_n7636_8799.n255 15.3369
R692 a_n7636_8799.n226 a_n7636_8799.n225 15.3369
R693 a_n7636_8799.n318 a_n7636_8799.n317 15.3369
R694 a_n7636_8799.n288 a_n7636_8799.n287 15.3369
R695 a_n7636_8799.n381 a_n7636_8799.n380 15.3369
R696 a_n7636_8799.n351 a_n7636_8799.n350 15.3369
R697 a_n7636_8799.n36 a_n7636_8799.n27 15.3369
R698 a_n7636_8799.n68 a_n7636_8799.n67 15.3369
R699 a_n7636_8799.n98 a_n7636_8799.n89 15.3369
R700 a_n7636_8799.n130 a_n7636_8799.n129 15.3369
R701 a_n7636_8799.n161 a_n7636_8799.n152 15.3369
R702 a_n7636_8799.n193 a_n7636_8799.n192 15.3369
R703 a_n7636_8799.n249 a_n7636_8799.n248 13.8763
R704 a_n7636_8799.n233 a_n7636_8799.n232 13.8763
R705 a_n7636_8799.n311 a_n7636_8799.n310 13.8763
R706 a_n7636_8799.n295 a_n7636_8799.n294 13.8763
R707 a_n7636_8799.n374 a_n7636_8799.n373 13.8763
R708 a_n7636_8799.n358 a_n7636_8799.n357 13.8763
R709 a_n7636_8799.n43 a_n7636_8799.n42 13.8763
R710 a_n7636_8799.n61 a_n7636_8799.n60 13.8763
R711 a_n7636_8799.n105 a_n7636_8799.n104 13.8763
R712 a_n7636_8799.n123 a_n7636_8799.n122 13.8763
R713 a_n7636_8799.n168 a_n7636_8799.n167 13.8763
R714 a_n7636_8799.n186 a_n7636_8799.n185 13.8763
R715 a_n7636_8799.n242 a_n7636_8799.n241 12.4157
R716 a_n7636_8799.n240 a_n7636_8799.n239 12.4157
R717 a_n7636_8799.n304 a_n7636_8799.n303 12.4157
R718 a_n7636_8799.n302 a_n7636_8799.n301 12.4157
R719 a_n7636_8799.n367 a_n7636_8799.n366 12.4157
R720 a_n7636_8799.n365 a_n7636_8799.n364 12.4157
R721 a_n7636_8799.n50 a_n7636_8799.n49 12.4157
R722 a_n7636_8799.n54 a_n7636_8799.n21 12.4157
R723 a_n7636_8799.n112 a_n7636_8799.n111 12.4157
R724 a_n7636_8799.n116 a_n7636_8799.n83 12.4157
R725 a_n7636_8799.n175 a_n7636_8799.n174 12.4157
R726 a_n7636_8799.n179 a_n7636_8799.n146 12.4157
R727 a_n7636_8799.n397 a_n7636_8799.n391 12.3339
R728 a_n7636_8799.n391 a_n7636_8799.n13 11.4887
R729 a_n7636_8799.n247 a_n7636_8799.n246 10.955
R730 a_n7636_8799.n235 a_n7636_8799.n234 10.955
R731 a_n7636_8799.n309 a_n7636_8799.n308 10.955
R732 a_n7636_8799.n297 a_n7636_8799.n296 10.955
R733 a_n7636_8799.n372 a_n7636_8799.n371 10.955
R734 a_n7636_8799.n360 a_n7636_8799.n359 10.955
R735 a_n7636_8799.n44 a_n7636_8799.n23 10.955
R736 a_n7636_8799.n56 a_n7636_8799.n19 10.955
R737 a_n7636_8799.n106 a_n7636_8799.n85 10.955
R738 a_n7636_8799.n118 a_n7636_8799.n81 10.955
R739 a_n7636_8799.n169 a_n7636_8799.n148 10.955
R740 a_n7636_8799.n181 a_n7636_8799.n144 10.955
R741 a_n7636_8799.n254 a_n7636_8799.n253 9.49444
R742 a_n7636_8799.n228 a_n7636_8799.n227 9.49444
R743 a_n7636_8799.n316 a_n7636_8799.n315 9.49444
R744 a_n7636_8799.n290 a_n7636_8799.n289 9.49444
R745 a_n7636_8799.n379 a_n7636_8799.n378 9.49444
R746 a_n7636_8799.n353 a_n7636_8799.n352 9.49444
R747 a_n7636_8799.n38 a_n7636_8799.n37 9.49444
R748 a_n7636_8799.n66 a_n7636_8799.n17 9.49444
R749 a_n7636_8799.n100 a_n7636_8799.n99 9.49444
R750 a_n7636_8799.n128 a_n7636_8799.n79 9.49444
R751 a_n7636_8799.n163 a_n7636_8799.n162 9.49444
R752 a_n7636_8799.n191 a_n7636_8799.n142 9.49444
R753 a_n7636_8799.n326 a_n7636_8799.n263 9.04406
R754 a_n7636_8799.n138 a_n7636_8799.n75 9.04406
R755 a_n7636_8799.n261 a_n7636_8799.n260 8.03383
R756 a_n7636_8799.n221 a_n7636_8799.n220 8.03383
R757 a_n7636_8799.n323 a_n7636_8799.n322 8.03383
R758 a_n7636_8799.n283 a_n7636_8799.n282 8.03383
R759 a_n7636_8799.n386 a_n7636_8799.n385 8.03383
R760 a_n7636_8799.n346 a_n7636_8799.n345 8.03383
R761 a_n7636_8799.n31 a_n7636_8799.n30 8.03383
R762 a_n7636_8799.n73 a_n7636_8799.n72 8.03383
R763 a_n7636_8799.n93 a_n7636_8799.n92 8.03383
R764 a_n7636_8799.n135 a_n7636_8799.n134 8.03383
R765 a_n7636_8799.n156 a_n7636_8799.n155 8.03383
R766 a_n7636_8799.n198 a_n7636_8799.n197 8.03383
R767 a_n7636_8799.n390 a_n7636_8799.n201 6.90212
R768 a_n7636_8799.n390 a_n7636_8799.n389 6.48069
R769 a_n7636_8799.n326 a_n7636_8799.n325 4.93611
R770 a_n7636_8799.n389 a_n7636_8799.n388 4.93611
R771 a_n7636_8799.n138 a_n7636_8799.n137 4.93611
R772 a_n7636_8799.n201 a_n7636_8799.n200 4.93611
R773 a_n7636_8799.n389 a_n7636_8799.n326 4.10845
R774 a_n7636_8799.n201 a_n7636_8799.n138 4.10845
R775 a_n7636_8799.n11 a_n7636_8799.t2 3.61217
R776 a_n7636_8799.n11 a_n7636_8799.t1 3.61217
R777 a_n7636_8799.n9 a_n7636_8799.t31 3.61217
R778 a_n7636_8799.n9 a_n7636_8799.t34 3.61217
R779 a_n7636_8799.n8 a_n7636_8799.t0 3.61217
R780 a_n7636_8799.n8 a_n7636_8799.t4 3.61217
R781 a_n7636_8799.n3 a_n7636_8799.t29 3.61217
R782 a_n7636_8799.n3 a_n7636_8799.t33 3.61217
R783 a_n7636_8799.n4 a_n7636_8799.t35 3.61217
R784 a_n7636_8799.n4 a_n7636_8799.t3 3.61217
R785 a_n7636_8799.n6 a_n7636_8799.t30 3.61217
R786 a_n7636_8799.n6 a_n7636_8799.t32 3.61217
R787 a_n7636_8799.n391 a_n7636_8799.n390 3.4105
R788 a_n7636_8799.n404 a_n7636_8799.t20 2.82907
R789 a_n7636_8799.n404 a_n7636_8799.t18 2.82907
R790 a_n7636_8799.n405 a_n7636_8799.t9 2.82907
R791 a_n7636_8799.n405 a_n7636_8799.t15 2.82907
R792 a_n7636_8799.n407 a_n7636_8799.t27 2.82907
R793 a_n7636_8799.n407 a_n7636_8799.t10 2.82907
R794 a_n7636_8799.n1 a_n7636_8799.t17 2.82907
R795 a_n7636_8799.n1 a_n7636_8799.t16 2.82907
R796 a_n7636_8799.n0 a_n7636_8799.t12 2.82907
R797 a_n7636_8799.n0 a_n7636_8799.t11 2.82907
R798 a_n7636_8799.n402 a_n7636_8799.t23 2.82907
R799 a_n7636_8799.n402 a_n7636_8799.t25 2.82907
R800 a_n7636_8799.n400 a_n7636_8799.t21 2.82907
R801 a_n7636_8799.n400 a_n7636_8799.t5 2.82907
R802 a_n7636_8799.n398 a_n7636_8799.t26 2.82907
R803 a_n7636_8799.n398 a_n7636_8799.t19 2.82907
R804 a_n7636_8799.n395 a_n7636_8799.t6 2.82907
R805 a_n7636_8799.n395 a_n7636_8799.t24 2.82907
R806 a_n7636_8799.n393 a_n7636_8799.t7 2.82907
R807 a_n7636_8799.n393 a_n7636_8799.t8 2.82907
R808 a_n7636_8799.n392 a_n7636_8799.t13 2.82907
R809 a_n7636_8799.n392 a_n7636_8799.t14 2.82907
R810 a_n7636_8799.n411 a_n7636_8799.t22 2.82907
R811 a_n7636_8799.t28 a_n7636_8799.n411 2.82907
R812 a_n7636_8799.n396 a_n7636_8799.n394 0.444466
R813 a_n7636_8799.n401 a_n7636_8799.n399 0.444466
R814 a_n7636_8799.n403 a_n7636_8799.n401 0.444466
R815 a_n7636_8799.n410 a_n7636_8799.n2 0.444466
R816 a_n7636_8799.n408 a_n7636_8799.n406 0.444466
R817 a_n7636_8799.n12 a_n7636_8799.n10 0.358259
R818 a_n7636_8799.n7 a_n7636_8799.n5 0.358259
R819 a_n7636_8799.n397 a_n7636_8799.n396 0.222483
R820 a_n7636_8799.n399 a_n7636_8799.n397 0.222483
R821 a_n7636_8799.n410 a_n7636_8799.n409 0.222483
R822 a_n7636_8799.n409 a_n7636_8799.n408 0.222483
R823 a_n7636_8799.n263 a_n7636_8799.n202 0.189894
R824 a_n7636_8799.n259 a_n7636_8799.n202 0.189894
R825 a_n7636_8799.n259 a_n7636_8799.n258 0.189894
R826 a_n7636_8799.n258 a_n7636_8799.n257 0.189894
R827 a_n7636_8799.n257 a_n7636_8799.n204 0.189894
R828 a_n7636_8799.n205 a_n7636_8799.n204 0.189894
R829 a_n7636_8799.n252 a_n7636_8799.n205 0.189894
R830 a_n7636_8799.n252 a_n7636_8799.n251 0.189894
R831 a_n7636_8799.n251 a_n7636_8799.n250 0.189894
R832 a_n7636_8799.n250 a_n7636_8799.n207 0.189894
R833 a_n7636_8799.n208 a_n7636_8799.n207 0.189894
R834 a_n7636_8799.n245 a_n7636_8799.n208 0.189894
R835 a_n7636_8799.n245 a_n7636_8799.n244 0.189894
R836 a_n7636_8799.n244 a_n7636_8799.n243 0.189894
R837 a_n7636_8799.n243 a_n7636_8799.n210 0.189894
R838 a_n7636_8799.n211 a_n7636_8799.n210 0.189894
R839 a_n7636_8799.n238 a_n7636_8799.n211 0.189894
R840 a_n7636_8799.n238 a_n7636_8799.n237 0.189894
R841 a_n7636_8799.n237 a_n7636_8799.n236 0.189894
R842 a_n7636_8799.n236 a_n7636_8799.n213 0.189894
R843 a_n7636_8799.n214 a_n7636_8799.n213 0.189894
R844 a_n7636_8799.n231 a_n7636_8799.n214 0.189894
R845 a_n7636_8799.n231 a_n7636_8799.n230 0.189894
R846 a_n7636_8799.n230 a_n7636_8799.n229 0.189894
R847 a_n7636_8799.n229 a_n7636_8799.n216 0.189894
R848 a_n7636_8799.n217 a_n7636_8799.n216 0.189894
R849 a_n7636_8799.n224 a_n7636_8799.n217 0.189894
R850 a_n7636_8799.n224 a_n7636_8799.n223 0.189894
R851 a_n7636_8799.n223 a_n7636_8799.n222 0.189894
R852 a_n7636_8799.n325 a_n7636_8799.n264 0.189894
R853 a_n7636_8799.n321 a_n7636_8799.n264 0.189894
R854 a_n7636_8799.n321 a_n7636_8799.n320 0.189894
R855 a_n7636_8799.n320 a_n7636_8799.n319 0.189894
R856 a_n7636_8799.n319 a_n7636_8799.n266 0.189894
R857 a_n7636_8799.n267 a_n7636_8799.n266 0.189894
R858 a_n7636_8799.n314 a_n7636_8799.n267 0.189894
R859 a_n7636_8799.n314 a_n7636_8799.n313 0.189894
R860 a_n7636_8799.n313 a_n7636_8799.n312 0.189894
R861 a_n7636_8799.n312 a_n7636_8799.n269 0.189894
R862 a_n7636_8799.n270 a_n7636_8799.n269 0.189894
R863 a_n7636_8799.n307 a_n7636_8799.n270 0.189894
R864 a_n7636_8799.n307 a_n7636_8799.n306 0.189894
R865 a_n7636_8799.n306 a_n7636_8799.n305 0.189894
R866 a_n7636_8799.n305 a_n7636_8799.n272 0.189894
R867 a_n7636_8799.n273 a_n7636_8799.n272 0.189894
R868 a_n7636_8799.n300 a_n7636_8799.n273 0.189894
R869 a_n7636_8799.n300 a_n7636_8799.n299 0.189894
R870 a_n7636_8799.n299 a_n7636_8799.n298 0.189894
R871 a_n7636_8799.n298 a_n7636_8799.n275 0.189894
R872 a_n7636_8799.n276 a_n7636_8799.n275 0.189894
R873 a_n7636_8799.n293 a_n7636_8799.n276 0.189894
R874 a_n7636_8799.n293 a_n7636_8799.n292 0.189894
R875 a_n7636_8799.n292 a_n7636_8799.n291 0.189894
R876 a_n7636_8799.n291 a_n7636_8799.n278 0.189894
R877 a_n7636_8799.n279 a_n7636_8799.n278 0.189894
R878 a_n7636_8799.n286 a_n7636_8799.n279 0.189894
R879 a_n7636_8799.n286 a_n7636_8799.n285 0.189894
R880 a_n7636_8799.n285 a_n7636_8799.n284 0.189894
R881 a_n7636_8799.n388 a_n7636_8799.n327 0.189894
R882 a_n7636_8799.n384 a_n7636_8799.n327 0.189894
R883 a_n7636_8799.n384 a_n7636_8799.n383 0.189894
R884 a_n7636_8799.n383 a_n7636_8799.n382 0.189894
R885 a_n7636_8799.n382 a_n7636_8799.n329 0.189894
R886 a_n7636_8799.n330 a_n7636_8799.n329 0.189894
R887 a_n7636_8799.n377 a_n7636_8799.n330 0.189894
R888 a_n7636_8799.n377 a_n7636_8799.n376 0.189894
R889 a_n7636_8799.n376 a_n7636_8799.n375 0.189894
R890 a_n7636_8799.n375 a_n7636_8799.n332 0.189894
R891 a_n7636_8799.n333 a_n7636_8799.n332 0.189894
R892 a_n7636_8799.n370 a_n7636_8799.n333 0.189894
R893 a_n7636_8799.n370 a_n7636_8799.n369 0.189894
R894 a_n7636_8799.n369 a_n7636_8799.n368 0.189894
R895 a_n7636_8799.n368 a_n7636_8799.n335 0.189894
R896 a_n7636_8799.n336 a_n7636_8799.n335 0.189894
R897 a_n7636_8799.n363 a_n7636_8799.n336 0.189894
R898 a_n7636_8799.n363 a_n7636_8799.n362 0.189894
R899 a_n7636_8799.n362 a_n7636_8799.n361 0.189894
R900 a_n7636_8799.n361 a_n7636_8799.n338 0.189894
R901 a_n7636_8799.n339 a_n7636_8799.n338 0.189894
R902 a_n7636_8799.n356 a_n7636_8799.n339 0.189894
R903 a_n7636_8799.n356 a_n7636_8799.n355 0.189894
R904 a_n7636_8799.n355 a_n7636_8799.n354 0.189894
R905 a_n7636_8799.n354 a_n7636_8799.n341 0.189894
R906 a_n7636_8799.n342 a_n7636_8799.n341 0.189894
R907 a_n7636_8799.n349 a_n7636_8799.n342 0.189894
R908 a_n7636_8799.n349 a_n7636_8799.n348 0.189894
R909 a_n7636_8799.n348 a_n7636_8799.n347 0.189894
R910 a_n7636_8799.n33 a_n7636_8799.n28 0.189894
R911 a_n7636_8799.n34 a_n7636_8799.n33 0.189894
R912 a_n7636_8799.n35 a_n7636_8799.n34 0.189894
R913 a_n7636_8799.n35 a_n7636_8799.n26 0.189894
R914 a_n7636_8799.n39 a_n7636_8799.n26 0.189894
R915 a_n7636_8799.n40 a_n7636_8799.n39 0.189894
R916 a_n7636_8799.n41 a_n7636_8799.n40 0.189894
R917 a_n7636_8799.n41 a_n7636_8799.n24 0.189894
R918 a_n7636_8799.n45 a_n7636_8799.n24 0.189894
R919 a_n7636_8799.n46 a_n7636_8799.n45 0.189894
R920 a_n7636_8799.n47 a_n7636_8799.n46 0.189894
R921 a_n7636_8799.n47 a_n7636_8799.n22 0.189894
R922 a_n7636_8799.n51 a_n7636_8799.n22 0.189894
R923 a_n7636_8799.n52 a_n7636_8799.n51 0.189894
R924 a_n7636_8799.n53 a_n7636_8799.n52 0.189894
R925 a_n7636_8799.n53 a_n7636_8799.n20 0.189894
R926 a_n7636_8799.n57 a_n7636_8799.n20 0.189894
R927 a_n7636_8799.n58 a_n7636_8799.n57 0.189894
R928 a_n7636_8799.n59 a_n7636_8799.n58 0.189894
R929 a_n7636_8799.n59 a_n7636_8799.n18 0.189894
R930 a_n7636_8799.n63 a_n7636_8799.n18 0.189894
R931 a_n7636_8799.n64 a_n7636_8799.n63 0.189894
R932 a_n7636_8799.n65 a_n7636_8799.n64 0.189894
R933 a_n7636_8799.n65 a_n7636_8799.n16 0.189894
R934 a_n7636_8799.n69 a_n7636_8799.n16 0.189894
R935 a_n7636_8799.n70 a_n7636_8799.n69 0.189894
R936 a_n7636_8799.n71 a_n7636_8799.n70 0.189894
R937 a_n7636_8799.n71 a_n7636_8799.n14 0.189894
R938 a_n7636_8799.n75 a_n7636_8799.n14 0.189894
R939 a_n7636_8799.n95 a_n7636_8799.n90 0.189894
R940 a_n7636_8799.n96 a_n7636_8799.n95 0.189894
R941 a_n7636_8799.n97 a_n7636_8799.n96 0.189894
R942 a_n7636_8799.n97 a_n7636_8799.n88 0.189894
R943 a_n7636_8799.n101 a_n7636_8799.n88 0.189894
R944 a_n7636_8799.n102 a_n7636_8799.n101 0.189894
R945 a_n7636_8799.n103 a_n7636_8799.n102 0.189894
R946 a_n7636_8799.n103 a_n7636_8799.n86 0.189894
R947 a_n7636_8799.n107 a_n7636_8799.n86 0.189894
R948 a_n7636_8799.n108 a_n7636_8799.n107 0.189894
R949 a_n7636_8799.n109 a_n7636_8799.n108 0.189894
R950 a_n7636_8799.n109 a_n7636_8799.n84 0.189894
R951 a_n7636_8799.n113 a_n7636_8799.n84 0.189894
R952 a_n7636_8799.n114 a_n7636_8799.n113 0.189894
R953 a_n7636_8799.n115 a_n7636_8799.n114 0.189894
R954 a_n7636_8799.n115 a_n7636_8799.n82 0.189894
R955 a_n7636_8799.n119 a_n7636_8799.n82 0.189894
R956 a_n7636_8799.n120 a_n7636_8799.n119 0.189894
R957 a_n7636_8799.n121 a_n7636_8799.n120 0.189894
R958 a_n7636_8799.n121 a_n7636_8799.n80 0.189894
R959 a_n7636_8799.n125 a_n7636_8799.n80 0.189894
R960 a_n7636_8799.n126 a_n7636_8799.n125 0.189894
R961 a_n7636_8799.n127 a_n7636_8799.n126 0.189894
R962 a_n7636_8799.n127 a_n7636_8799.n78 0.189894
R963 a_n7636_8799.n131 a_n7636_8799.n78 0.189894
R964 a_n7636_8799.n132 a_n7636_8799.n131 0.189894
R965 a_n7636_8799.n133 a_n7636_8799.n132 0.189894
R966 a_n7636_8799.n133 a_n7636_8799.n76 0.189894
R967 a_n7636_8799.n137 a_n7636_8799.n76 0.189894
R968 a_n7636_8799.n158 a_n7636_8799.n153 0.189894
R969 a_n7636_8799.n159 a_n7636_8799.n158 0.189894
R970 a_n7636_8799.n160 a_n7636_8799.n159 0.189894
R971 a_n7636_8799.n160 a_n7636_8799.n151 0.189894
R972 a_n7636_8799.n164 a_n7636_8799.n151 0.189894
R973 a_n7636_8799.n165 a_n7636_8799.n164 0.189894
R974 a_n7636_8799.n166 a_n7636_8799.n165 0.189894
R975 a_n7636_8799.n166 a_n7636_8799.n149 0.189894
R976 a_n7636_8799.n170 a_n7636_8799.n149 0.189894
R977 a_n7636_8799.n171 a_n7636_8799.n170 0.189894
R978 a_n7636_8799.n172 a_n7636_8799.n171 0.189894
R979 a_n7636_8799.n172 a_n7636_8799.n147 0.189894
R980 a_n7636_8799.n176 a_n7636_8799.n147 0.189894
R981 a_n7636_8799.n177 a_n7636_8799.n176 0.189894
R982 a_n7636_8799.n178 a_n7636_8799.n177 0.189894
R983 a_n7636_8799.n178 a_n7636_8799.n145 0.189894
R984 a_n7636_8799.n182 a_n7636_8799.n145 0.189894
R985 a_n7636_8799.n183 a_n7636_8799.n182 0.189894
R986 a_n7636_8799.n184 a_n7636_8799.n183 0.189894
R987 a_n7636_8799.n184 a_n7636_8799.n143 0.189894
R988 a_n7636_8799.n188 a_n7636_8799.n143 0.189894
R989 a_n7636_8799.n189 a_n7636_8799.n188 0.189894
R990 a_n7636_8799.n190 a_n7636_8799.n189 0.189894
R991 a_n7636_8799.n190 a_n7636_8799.n141 0.189894
R992 a_n7636_8799.n194 a_n7636_8799.n141 0.189894
R993 a_n7636_8799.n195 a_n7636_8799.n194 0.189894
R994 a_n7636_8799.n196 a_n7636_8799.n195 0.189894
R995 a_n7636_8799.n196 a_n7636_8799.n139 0.189894
R996 a_n7636_8799.n200 a_n7636_8799.n139 0.189894
R997 gnd.n6905 gnd.n544 2174.34
R998 gnd.n4211 gnd.n3911 939.716
R999 gnd.n7282 gnd.n171 838.452
R1000 gnd.n7250 gnd.n169 838.452
R1001 gnd.n5138 gnd.n1608 838.452
R1002 gnd.n5206 gnd.n1610 838.452
R1003 gnd.n6198 gnd.n1142 838.452
R1004 gnd.n6118 gnd.n1140 838.452
R1005 gnd.n4049 gnd.n3949 838.452
R1006 gnd.n4090 gnd.n4089 838.452
R1007 gnd.n7284 gnd.n166 783.196
R1008 gnd.n382 gnd.n168 783.196
R1009 gnd.n5658 gnd.n1607 783.196
R1010 gnd.n5857 gnd.n1611 783.196
R1011 gnd.n6200 gnd.n1137 783.196
R1012 gnd.n1347 gnd.n1139 783.196
R1013 gnd.n4010 gnd.n2441 783.196
R1014 gnd.n4213 gnd.n2445 783.196
R1015 gnd.n6179 gnd.n1171 771.183
R1016 gnd.n5875 gnd.n1585 771.183
R1017 gnd.n6183 gnd.n1153 771.183
R1018 gnd.n5294 gnd.n1587 771.183
R1019 gnd.n3819 gnd.n2451 766.379
R1020 gnd.n3822 gnd.n3821 766.379
R1021 gnd.n3061 gnd.n2964 766.379
R1022 gnd.n3057 gnd.n2962 766.379
R1023 gnd.n3910 gnd.n2473 756.769
R1024 gnd.n3813 gnd.n3812 756.769
R1025 gnd.n3154 gnd.n2871 756.769
R1026 gnd.n3152 gnd.n2874 756.769
R1027 gnd.n6483 gnd.n796 756.769
R1028 gnd.n6904 gnd.n545 756.769
R1029 gnd.n7117 gnd.n7116 756.769
R1030 gnd.n6307 gnd.n961 756.769
R1031 gnd.n6479 gnd.n796 585
R1032 gnd.n796 gnd.n795 585
R1033 gnd.n6478 gnd.n6477 585
R1034 gnd.n6477 gnd.n6476 585
R1035 gnd.n799 gnd.n798 585
R1036 gnd.n6475 gnd.n799 585
R1037 gnd.n6473 gnd.n6472 585
R1038 gnd.n6474 gnd.n6473 585
R1039 gnd.n6471 gnd.n801 585
R1040 gnd.n801 gnd.n800 585
R1041 gnd.n6470 gnd.n6469 585
R1042 gnd.n6469 gnd.n6468 585
R1043 gnd.n807 gnd.n806 585
R1044 gnd.n6467 gnd.n807 585
R1045 gnd.n6465 gnd.n6464 585
R1046 gnd.n6466 gnd.n6465 585
R1047 gnd.n6463 gnd.n809 585
R1048 gnd.n809 gnd.n808 585
R1049 gnd.n6462 gnd.n6461 585
R1050 gnd.n6461 gnd.n6460 585
R1051 gnd.n815 gnd.n814 585
R1052 gnd.n6459 gnd.n815 585
R1053 gnd.n6457 gnd.n6456 585
R1054 gnd.n6458 gnd.n6457 585
R1055 gnd.n6455 gnd.n817 585
R1056 gnd.n817 gnd.n816 585
R1057 gnd.n6454 gnd.n6453 585
R1058 gnd.n6453 gnd.n6452 585
R1059 gnd.n823 gnd.n822 585
R1060 gnd.n6451 gnd.n823 585
R1061 gnd.n6449 gnd.n6448 585
R1062 gnd.n6450 gnd.n6449 585
R1063 gnd.n6447 gnd.n825 585
R1064 gnd.n825 gnd.n824 585
R1065 gnd.n6446 gnd.n6445 585
R1066 gnd.n6445 gnd.n6444 585
R1067 gnd.n831 gnd.n830 585
R1068 gnd.n6443 gnd.n831 585
R1069 gnd.n6441 gnd.n6440 585
R1070 gnd.n6442 gnd.n6441 585
R1071 gnd.n6439 gnd.n833 585
R1072 gnd.n833 gnd.n832 585
R1073 gnd.n6438 gnd.n6437 585
R1074 gnd.n6437 gnd.n6436 585
R1075 gnd.n839 gnd.n838 585
R1076 gnd.n6435 gnd.n839 585
R1077 gnd.n6433 gnd.n6432 585
R1078 gnd.n6434 gnd.n6433 585
R1079 gnd.n6431 gnd.n841 585
R1080 gnd.n841 gnd.n840 585
R1081 gnd.n6430 gnd.n6429 585
R1082 gnd.n6429 gnd.n6428 585
R1083 gnd.n847 gnd.n846 585
R1084 gnd.n6427 gnd.n847 585
R1085 gnd.n6425 gnd.n6424 585
R1086 gnd.n6426 gnd.n6425 585
R1087 gnd.n6423 gnd.n849 585
R1088 gnd.n849 gnd.n848 585
R1089 gnd.n6422 gnd.n6421 585
R1090 gnd.n6421 gnd.n6420 585
R1091 gnd.n855 gnd.n854 585
R1092 gnd.n6419 gnd.n855 585
R1093 gnd.n6417 gnd.n6416 585
R1094 gnd.n6418 gnd.n6417 585
R1095 gnd.n6415 gnd.n857 585
R1096 gnd.n857 gnd.n856 585
R1097 gnd.n6414 gnd.n6413 585
R1098 gnd.n6413 gnd.n6412 585
R1099 gnd.n863 gnd.n862 585
R1100 gnd.n6411 gnd.n863 585
R1101 gnd.n6409 gnd.n6408 585
R1102 gnd.n6410 gnd.n6409 585
R1103 gnd.n6407 gnd.n865 585
R1104 gnd.n865 gnd.n864 585
R1105 gnd.n6406 gnd.n6405 585
R1106 gnd.n6405 gnd.n6404 585
R1107 gnd.n871 gnd.n870 585
R1108 gnd.n6403 gnd.n871 585
R1109 gnd.n6401 gnd.n6400 585
R1110 gnd.n6402 gnd.n6401 585
R1111 gnd.n6399 gnd.n873 585
R1112 gnd.n873 gnd.n872 585
R1113 gnd.n6398 gnd.n6397 585
R1114 gnd.n6397 gnd.n6396 585
R1115 gnd.n879 gnd.n878 585
R1116 gnd.n6395 gnd.n879 585
R1117 gnd.n6393 gnd.n6392 585
R1118 gnd.n6394 gnd.n6393 585
R1119 gnd.n6391 gnd.n881 585
R1120 gnd.n881 gnd.n880 585
R1121 gnd.n6390 gnd.n6389 585
R1122 gnd.n6389 gnd.n6388 585
R1123 gnd.n887 gnd.n886 585
R1124 gnd.n6387 gnd.n887 585
R1125 gnd.n6385 gnd.n6384 585
R1126 gnd.n6386 gnd.n6385 585
R1127 gnd.n6383 gnd.n889 585
R1128 gnd.n889 gnd.n888 585
R1129 gnd.n6382 gnd.n6381 585
R1130 gnd.n6381 gnd.n6380 585
R1131 gnd.n895 gnd.n894 585
R1132 gnd.n6379 gnd.n895 585
R1133 gnd.n6377 gnd.n6376 585
R1134 gnd.n6378 gnd.n6377 585
R1135 gnd.n6375 gnd.n897 585
R1136 gnd.n897 gnd.n896 585
R1137 gnd.n6374 gnd.n6373 585
R1138 gnd.n6373 gnd.n6372 585
R1139 gnd.n903 gnd.n902 585
R1140 gnd.n6371 gnd.n903 585
R1141 gnd.n6369 gnd.n6368 585
R1142 gnd.n6370 gnd.n6369 585
R1143 gnd.n6367 gnd.n905 585
R1144 gnd.n905 gnd.n904 585
R1145 gnd.n6366 gnd.n6365 585
R1146 gnd.n6365 gnd.n6364 585
R1147 gnd.n911 gnd.n910 585
R1148 gnd.n6363 gnd.n911 585
R1149 gnd.n6361 gnd.n6360 585
R1150 gnd.n6362 gnd.n6361 585
R1151 gnd.n6359 gnd.n913 585
R1152 gnd.n913 gnd.n912 585
R1153 gnd.n6358 gnd.n6357 585
R1154 gnd.n6357 gnd.n6356 585
R1155 gnd.n919 gnd.n918 585
R1156 gnd.n6355 gnd.n919 585
R1157 gnd.n6353 gnd.n6352 585
R1158 gnd.n6354 gnd.n6353 585
R1159 gnd.n6351 gnd.n921 585
R1160 gnd.n921 gnd.n920 585
R1161 gnd.n6350 gnd.n6349 585
R1162 gnd.n6349 gnd.n6348 585
R1163 gnd.n927 gnd.n926 585
R1164 gnd.n6347 gnd.n927 585
R1165 gnd.n6345 gnd.n6344 585
R1166 gnd.n6346 gnd.n6345 585
R1167 gnd.n6343 gnd.n929 585
R1168 gnd.n929 gnd.n928 585
R1169 gnd.n6342 gnd.n6341 585
R1170 gnd.n6341 gnd.n6340 585
R1171 gnd.n935 gnd.n934 585
R1172 gnd.n6339 gnd.n935 585
R1173 gnd.n6337 gnd.n6336 585
R1174 gnd.n6338 gnd.n6337 585
R1175 gnd.n6335 gnd.n937 585
R1176 gnd.n937 gnd.n936 585
R1177 gnd.n6334 gnd.n6333 585
R1178 gnd.n6333 gnd.n6332 585
R1179 gnd.n943 gnd.n942 585
R1180 gnd.n6331 gnd.n943 585
R1181 gnd.n6329 gnd.n6328 585
R1182 gnd.n6330 gnd.n6329 585
R1183 gnd.n6327 gnd.n945 585
R1184 gnd.n945 gnd.n944 585
R1185 gnd.n6326 gnd.n6325 585
R1186 gnd.n6325 gnd.n6324 585
R1187 gnd.n951 gnd.n950 585
R1188 gnd.n6323 gnd.n951 585
R1189 gnd.n6321 gnd.n6320 585
R1190 gnd.n6322 gnd.n6321 585
R1191 gnd.n6319 gnd.n953 585
R1192 gnd.n953 gnd.n952 585
R1193 gnd.n6318 gnd.n6317 585
R1194 gnd.n6317 gnd.n6316 585
R1195 gnd.n959 gnd.n958 585
R1196 gnd.n6315 gnd.n959 585
R1197 gnd.n6313 gnd.n6312 585
R1198 gnd.n6314 gnd.n6313 585
R1199 gnd.n6483 gnd.n6482 585
R1200 gnd.n6484 gnd.n6483 585
R1201 gnd.n794 gnd.n793 585
R1202 gnd.n6485 gnd.n794 585
R1203 gnd.n6488 gnd.n6487 585
R1204 gnd.n6487 gnd.n6486 585
R1205 gnd.n791 gnd.n790 585
R1206 gnd.n790 gnd.n789 585
R1207 gnd.n6493 gnd.n6492 585
R1208 gnd.n6494 gnd.n6493 585
R1209 gnd.n788 gnd.n787 585
R1210 gnd.n6495 gnd.n788 585
R1211 gnd.n6498 gnd.n6497 585
R1212 gnd.n6497 gnd.n6496 585
R1213 gnd.n785 gnd.n784 585
R1214 gnd.n784 gnd.n783 585
R1215 gnd.n6503 gnd.n6502 585
R1216 gnd.n6504 gnd.n6503 585
R1217 gnd.n782 gnd.n781 585
R1218 gnd.n6505 gnd.n782 585
R1219 gnd.n6508 gnd.n6507 585
R1220 gnd.n6507 gnd.n6506 585
R1221 gnd.n779 gnd.n778 585
R1222 gnd.n778 gnd.n777 585
R1223 gnd.n6513 gnd.n6512 585
R1224 gnd.n6514 gnd.n6513 585
R1225 gnd.n776 gnd.n775 585
R1226 gnd.n6515 gnd.n776 585
R1227 gnd.n6518 gnd.n6517 585
R1228 gnd.n6517 gnd.n6516 585
R1229 gnd.n773 gnd.n772 585
R1230 gnd.n772 gnd.n771 585
R1231 gnd.n6523 gnd.n6522 585
R1232 gnd.n6524 gnd.n6523 585
R1233 gnd.n770 gnd.n769 585
R1234 gnd.n6525 gnd.n770 585
R1235 gnd.n6528 gnd.n6527 585
R1236 gnd.n6527 gnd.n6526 585
R1237 gnd.n767 gnd.n766 585
R1238 gnd.n766 gnd.n765 585
R1239 gnd.n6533 gnd.n6532 585
R1240 gnd.n6534 gnd.n6533 585
R1241 gnd.n764 gnd.n763 585
R1242 gnd.n6535 gnd.n764 585
R1243 gnd.n6538 gnd.n6537 585
R1244 gnd.n6537 gnd.n6536 585
R1245 gnd.n761 gnd.n760 585
R1246 gnd.n760 gnd.n759 585
R1247 gnd.n6543 gnd.n6542 585
R1248 gnd.n6544 gnd.n6543 585
R1249 gnd.n758 gnd.n757 585
R1250 gnd.n6545 gnd.n758 585
R1251 gnd.n6548 gnd.n6547 585
R1252 gnd.n6547 gnd.n6546 585
R1253 gnd.n755 gnd.n754 585
R1254 gnd.n754 gnd.n753 585
R1255 gnd.n6553 gnd.n6552 585
R1256 gnd.n6554 gnd.n6553 585
R1257 gnd.n752 gnd.n751 585
R1258 gnd.n6555 gnd.n752 585
R1259 gnd.n6558 gnd.n6557 585
R1260 gnd.n6557 gnd.n6556 585
R1261 gnd.n749 gnd.n748 585
R1262 gnd.n748 gnd.n747 585
R1263 gnd.n6563 gnd.n6562 585
R1264 gnd.n6564 gnd.n6563 585
R1265 gnd.n746 gnd.n745 585
R1266 gnd.n6565 gnd.n746 585
R1267 gnd.n6568 gnd.n6567 585
R1268 gnd.n6567 gnd.n6566 585
R1269 gnd.n743 gnd.n742 585
R1270 gnd.n742 gnd.n741 585
R1271 gnd.n6573 gnd.n6572 585
R1272 gnd.n6574 gnd.n6573 585
R1273 gnd.n740 gnd.n739 585
R1274 gnd.n6575 gnd.n740 585
R1275 gnd.n6578 gnd.n6577 585
R1276 gnd.n6577 gnd.n6576 585
R1277 gnd.n737 gnd.n736 585
R1278 gnd.n736 gnd.n735 585
R1279 gnd.n6583 gnd.n6582 585
R1280 gnd.n6584 gnd.n6583 585
R1281 gnd.n734 gnd.n733 585
R1282 gnd.n6585 gnd.n734 585
R1283 gnd.n6588 gnd.n6587 585
R1284 gnd.n6587 gnd.n6586 585
R1285 gnd.n731 gnd.n730 585
R1286 gnd.n730 gnd.n729 585
R1287 gnd.n6593 gnd.n6592 585
R1288 gnd.n6594 gnd.n6593 585
R1289 gnd.n728 gnd.n727 585
R1290 gnd.n6595 gnd.n728 585
R1291 gnd.n6598 gnd.n6597 585
R1292 gnd.n6597 gnd.n6596 585
R1293 gnd.n725 gnd.n724 585
R1294 gnd.n724 gnd.n723 585
R1295 gnd.n6603 gnd.n6602 585
R1296 gnd.n6604 gnd.n6603 585
R1297 gnd.n722 gnd.n721 585
R1298 gnd.n6605 gnd.n722 585
R1299 gnd.n6608 gnd.n6607 585
R1300 gnd.n6607 gnd.n6606 585
R1301 gnd.n719 gnd.n718 585
R1302 gnd.n718 gnd.n717 585
R1303 gnd.n6613 gnd.n6612 585
R1304 gnd.n6614 gnd.n6613 585
R1305 gnd.n716 gnd.n715 585
R1306 gnd.n6615 gnd.n716 585
R1307 gnd.n6618 gnd.n6617 585
R1308 gnd.n6617 gnd.n6616 585
R1309 gnd.n713 gnd.n712 585
R1310 gnd.n712 gnd.n711 585
R1311 gnd.n6623 gnd.n6622 585
R1312 gnd.n6624 gnd.n6623 585
R1313 gnd.n710 gnd.n709 585
R1314 gnd.n6625 gnd.n710 585
R1315 gnd.n6628 gnd.n6627 585
R1316 gnd.n6627 gnd.n6626 585
R1317 gnd.n707 gnd.n706 585
R1318 gnd.n706 gnd.n705 585
R1319 gnd.n6633 gnd.n6632 585
R1320 gnd.n6634 gnd.n6633 585
R1321 gnd.n704 gnd.n703 585
R1322 gnd.n6635 gnd.n704 585
R1323 gnd.n6638 gnd.n6637 585
R1324 gnd.n6637 gnd.n6636 585
R1325 gnd.n701 gnd.n700 585
R1326 gnd.n700 gnd.n699 585
R1327 gnd.n6643 gnd.n6642 585
R1328 gnd.n6644 gnd.n6643 585
R1329 gnd.n698 gnd.n697 585
R1330 gnd.n6645 gnd.n698 585
R1331 gnd.n6648 gnd.n6647 585
R1332 gnd.n6647 gnd.n6646 585
R1333 gnd.n695 gnd.n694 585
R1334 gnd.n694 gnd.n693 585
R1335 gnd.n6653 gnd.n6652 585
R1336 gnd.n6654 gnd.n6653 585
R1337 gnd.n692 gnd.n691 585
R1338 gnd.n6655 gnd.n692 585
R1339 gnd.n6658 gnd.n6657 585
R1340 gnd.n6657 gnd.n6656 585
R1341 gnd.n689 gnd.n688 585
R1342 gnd.n688 gnd.n687 585
R1343 gnd.n6663 gnd.n6662 585
R1344 gnd.n6664 gnd.n6663 585
R1345 gnd.n686 gnd.n685 585
R1346 gnd.n6665 gnd.n686 585
R1347 gnd.n6668 gnd.n6667 585
R1348 gnd.n6667 gnd.n6666 585
R1349 gnd.n683 gnd.n682 585
R1350 gnd.n682 gnd.n681 585
R1351 gnd.n6673 gnd.n6672 585
R1352 gnd.n6674 gnd.n6673 585
R1353 gnd.n680 gnd.n679 585
R1354 gnd.n6675 gnd.n680 585
R1355 gnd.n6678 gnd.n6677 585
R1356 gnd.n6677 gnd.n6676 585
R1357 gnd.n677 gnd.n676 585
R1358 gnd.n676 gnd.n675 585
R1359 gnd.n6683 gnd.n6682 585
R1360 gnd.n6684 gnd.n6683 585
R1361 gnd.n674 gnd.n673 585
R1362 gnd.n6685 gnd.n674 585
R1363 gnd.n6688 gnd.n6687 585
R1364 gnd.n6687 gnd.n6686 585
R1365 gnd.n671 gnd.n670 585
R1366 gnd.n670 gnd.n669 585
R1367 gnd.n6693 gnd.n6692 585
R1368 gnd.n6694 gnd.n6693 585
R1369 gnd.n668 gnd.n667 585
R1370 gnd.n6695 gnd.n668 585
R1371 gnd.n6698 gnd.n6697 585
R1372 gnd.n6697 gnd.n6696 585
R1373 gnd.n665 gnd.n664 585
R1374 gnd.n664 gnd.n663 585
R1375 gnd.n6703 gnd.n6702 585
R1376 gnd.n6704 gnd.n6703 585
R1377 gnd.n662 gnd.n661 585
R1378 gnd.n6705 gnd.n662 585
R1379 gnd.n6708 gnd.n6707 585
R1380 gnd.n6707 gnd.n6706 585
R1381 gnd.n659 gnd.n658 585
R1382 gnd.n658 gnd.n657 585
R1383 gnd.n6713 gnd.n6712 585
R1384 gnd.n6714 gnd.n6713 585
R1385 gnd.n656 gnd.n655 585
R1386 gnd.n6715 gnd.n656 585
R1387 gnd.n6718 gnd.n6717 585
R1388 gnd.n6717 gnd.n6716 585
R1389 gnd.n653 gnd.n652 585
R1390 gnd.n652 gnd.n651 585
R1391 gnd.n6723 gnd.n6722 585
R1392 gnd.n6724 gnd.n6723 585
R1393 gnd.n650 gnd.n649 585
R1394 gnd.n6725 gnd.n650 585
R1395 gnd.n6728 gnd.n6727 585
R1396 gnd.n6727 gnd.n6726 585
R1397 gnd.n647 gnd.n646 585
R1398 gnd.n646 gnd.n645 585
R1399 gnd.n6733 gnd.n6732 585
R1400 gnd.n6734 gnd.n6733 585
R1401 gnd.n644 gnd.n643 585
R1402 gnd.n6735 gnd.n644 585
R1403 gnd.n6738 gnd.n6737 585
R1404 gnd.n6737 gnd.n6736 585
R1405 gnd.n641 gnd.n640 585
R1406 gnd.n640 gnd.n639 585
R1407 gnd.n6743 gnd.n6742 585
R1408 gnd.n6744 gnd.n6743 585
R1409 gnd.n638 gnd.n637 585
R1410 gnd.n6745 gnd.n638 585
R1411 gnd.n6748 gnd.n6747 585
R1412 gnd.n6747 gnd.n6746 585
R1413 gnd.n635 gnd.n634 585
R1414 gnd.n634 gnd.n633 585
R1415 gnd.n6753 gnd.n6752 585
R1416 gnd.n6754 gnd.n6753 585
R1417 gnd.n632 gnd.n631 585
R1418 gnd.n6755 gnd.n632 585
R1419 gnd.n6758 gnd.n6757 585
R1420 gnd.n6757 gnd.n6756 585
R1421 gnd.n629 gnd.n628 585
R1422 gnd.n628 gnd.n627 585
R1423 gnd.n6763 gnd.n6762 585
R1424 gnd.n6764 gnd.n6763 585
R1425 gnd.n626 gnd.n625 585
R1426 gnd.n6765 gnd.n626 585
R1427 gnd.n6768 gnd.n6767 585
R1428 gnd.n6767 gnd.n6766 585
R1429 gnd.n623 gnd.n622 585
R1430 gnd.n622 gnd.n621 585
R1431 gnd.n6773 gnd.n6772 585
R1432 gnd.n6774 gnd.n6773 585
R1433 gnd.n620 gnd.n619 585
R1434 gnd.n6775 gnd.n620 585
R1435 gnd.n6778 gnd.n6777 585
R1436 gnd.n6777 gnd.n6776 585
R1437 gnd.n617 gnd.n616 585
R1438 gnd.n616 gnd.n615 585
R1439 gnd.n6783 gnd.n6782 585
R1440 gnd.n6784 gnd.n6783 585
R1441 gnd.n614 gnd.n613 585
R1442 gnd.n6785 gnd.n614 585
R1443 gnd.n6788 gnd.n6787 585
R1444 gnd.n6787 gnd.n6786 585
R1445 gnd.n611 gnd.n610 585
R1446 gnd.n610 gnd.n609 585
R1447 gnd.n6793 gnd.n6792 585
R1448 gnd.n6794 gnd.n6793 585
R1449 gnd.n608 gnd.n607 585
R1450 gnd.n6795 gnd.n608 585
R1451 gnd.n6798 gnd.n6797 585
R1452 gnd.n6797 gnd.n6796 585
R1453 gnd.n605 gnd.n604 585
R1454 gnd.n604 gnd.n603 585
R1455 gnd.n6803 gnd.n6802 585
R1456 gnd.n6804 gnd.n6803 585
R1457 gnd.n602 gnd.n601 585
R1458 gnd.n6805 gnd.n602 585
R1459 gnd.n6808 gnd.n6807 585
R1460 gnd.n6807 gnd.n6806 585
R1461 gnd.n599 gnd.n598 585
R1462 gnd.n598 gnd.n597 585
R1463 gnd.n6813 gnd.n6812 585
R1464 gnd.n6814 gnd.n6813 585
R1465 gnd.n596 gnd.n595 585
R1466 gnd.n6815 gnd.n596 585
R1467 gnd.n6818 gnd.n6817 585
R1468 gnd.n6817 gnd.n6816 585
R1469 gnd.n593 gnd.n592 585
R1470 gnd.n592 gnd.n591 585
R1471 gnd.n6823 gnd.n6822 585
R1472 gnd.n6824 gnd.n6823 585
R1473 gnd.n590 gnd.n589 585
R1474 gnd.n6825 gnd.n590 585
R1475 gnd.n6828 gnd.n6827 585
R1476 gnd.n6827 gnd.n6826 585
R1477 gnd.n587 gnd.n586 585
R1478 gnd.n586 gnd.n585 585
R1479 gnd.n6833 gnd.n6832 585
R1480 gnd.n6834 gnd.n6833 585
R1481 gnd.n584 gnd.n583 585
R1482 gnd.n6835 gnd.n584 585
R1483 gnd.n6838 gnd.n6837 585
R1484 gnd.n6837 gnd.n6836 585
R1485 gnd.n581 gnd.n580 585
R1486 gnd.n580 gnd.n579 585
R1487 gnd.n6843 gnd.n6842 585
R1488 gnd.n6844 gnd.n6843 585
R1489 gnd.n578 gnd.n577 585
R1490 gnd.n6845 gnd.n578 585
R1491 gnd.n6848 gnd.n6847 585
R1492 gnd.n6847 gnd.n6846 585
R1493 gnd.n575 gnd.n574 585
R1494 gnd.n574 gnd.n573 585
R1495 gnd.n6853 gnd.n6852 585
R1496 gnd.n6854 gnd.n6853 585
R1497 gnd.n572 gnd.n571 585
R1498 gnd.n6855 gnd.n572 585
R1499 gnd.n6858 gnd.n6857 585
R1500 gnd.n6857 gnd.n6856 585
R1501 gnd.n569 gnd.n568 585
R1502 gnd.n568 gnd.n567 585
R1503 gnd.n6863 gnd.n6862 585
R1504 gnd.n6864 gnd.n6863 585
R1505 gnd.n566 gnd.n565 585
R1506 gnd.n6865 gnd.n566 585
R1507 gnd.n6868 gnd.n6867 585
R1508 gnd.n6867 gnd.n6866 585
R1509 gnd.n563 gnd.n562 585
R1510 gnd.n562 gnd.n561 585
R1511 gnd.n6873 gnd.n6872 585
R1512 gnd.n6874 gnd.n6873 585
R1513 gnd.n560 gnd.n559 585
R1514 gnd.n6875 gnd.n560 585
R1515 gnd.n6878 gnd.n6877 585
R1516 gnd.n6877 gnd.n6876 585
R1517 gnd.n557 gnd.n556 585
R1518 gnd.n556 gnd.n555 585
R1519 gnd.n6883 gnd.n6882 585
R1520 gnd.n6884 gnd.n6883 585
R1521 gnd.n554 gnd.n553 585
R1522 gnd.n6885 gnd.n554 585
R1523 gnd.n6888 gnd.n6887 585
R1524 gnd.n6887 gnd.n6886 585
R1525 gnd.n551 gnd.n550 585
R1526 gnd.n550 gnd.n549 585
R1527 gnd.n6894 gnd.n6893 585
R1528 gnd.n6895 gnd.n6894 585
R1529 gnd.n548 gnd.n547 585
R1530 gnd.n6896 gnd.n548 585
R1531 gnd.n6899 gnd.n6898 585
R1532 gnd.n6898 gnd.n6897 585
R1533 gnd.n6900 gnd.n545 585
R1534 gnd.n545 gnd.n544 585
R1535 gnd.n420 gnd.n419 585
R1536 gnd.n7107 gnd.n419 585
R1537 gnd.n7110 gnd.n7109 585
R1538 gnd.n7109 gnd.n7108 585
R1539 gnd.n423 gnd.n422 585
R1540 gnd.n7106 gnd.n423 585
R1541 gnd.n7104 gnd.n7103 585
R1542 gnd.n7105 gnd.n7104 585
R1543 gnd.n426 gnd.n425 585
R1544 gnd.n425 gnd.n424 585
R1545 gnd.n7099 gnd.n7098 585
R1546 gnd.n7098 gnd.n7097 585
R1547 gnd.n429 gnd.n428 585
R1548 gnd.n7096 gnd.n429 585
R1549 gnd.n7094 gnd.n7093 585
R1550 gnd.n7095 gnd.n7094 585
R1551 gnd.n432 gnd.n431 585
R1552 gnd.n431 gnd.n430 585
R1553 gnd.n7089 gnd.n7088 585
R1554 gnd.n7088 gnd.n7087 585
R1555 gnd.n435 gnd.n434 585
R1556 gnd.n7086 gnd.n435 585
R1557 gnd.n7084 gnd.n7083 585
R1558 gnd.n7085 gnd.n7084 585
R1559 gnd.n438 gnd.n437 585
R1560 gnd.n437 gnd.n436 585
R1561 gnd.n7079 gnd.n7078 585
R1562 gnd.n7078 gnd.n7077 585
R1563 gnd.n441 gnd.n440 585
R1564 gnd.n7076 gnd.n441 585
R1565 gnd.n7074 gnd.n7073 585
R1566 gnd.n7075 gnd.n7074 585
R1567 gnd.n444 gnd.n443 585
R1568 gnd.n443 gnd.n442 585
R1569 gnd.n7069 gnd.n7068 585
R1570 gnd.n7068 gnd.n7067 585
R1571 gnd.n447 gnd.n446 585
R1572 gnd.n7066 gnd.n447 585
R1573 gnd.n7064 gnd.n7063 585
R1574 gnd.n7065 gnd.n7064 585
R1575 gnd.n450 gnd.n449 585
R1576 gnd.n449 gnd.n448 585
R1577 gnd.n7059 gnd.n7058 585
R1578 gnd.n7058 gnd.n7057 585
R1579 gnd.n453 gnd.n452 585
R1580 gnd.n7056 gnd.n453 585
R1581 gnd.n7054 gnd.n7053 585
R1582 gnd.n7055 gnd.n7054 585
R1583 gnd.n456 gnd.n455 585
R1584 gnd.n455 gnd.n454 585
R1585 gnd.n7049 gnd.n7048 585
R1586 gnd.n7048 gnd.n7047 585
R1587 gnd.n459 gnd.n458 585
R1588 gnd.n7046 gnd.n459 585
R1589 gnd.n7044 gnd.n7043 585
R1590 gnd.n7045 gnd.n7044 585
R1591 gnd.n462 gnd.n461 585
R1592 gnd.n461 gnd.n460 585
R1593 gnd.n7039 gnd.n7038 585
R1594 gnd.n7038 gnd.n7037 585
R1595 gnd.n465 gnd.n464 585
R1596 gnd.n7036 gnd.n465 585
R1597 gnd.n7034 gnd.n7033 585
R1598 gnd.n7035 gnd.n7034 585
R1599 gnd.n468 gnd.n467 585
R1600 gnd.n467 gnd.n466 585
R1601 gnd.n7029 gnd.n7028 585
R1602 gnd.n7028 gnd.n7027 585
R1603 gnd.n471 gnd.n470 585
R1604 gnd.n7026 gnd.n471 585
R1605 gnd.n7024 gnd.n7023 585
R1606 gnd.n7025 gnd.n7024 585
R1607 gnd.n474 gnd.n473 585
R1608 gnd.n473 gnd.n472 585
R1609 gnd.n7019 gnd.n7018 585
R1610 gnd.n7018 gnd.n7017 585
R1611 gnd.n477 gnd.n476 585
R1612 gnd.n7016 gnd.n477 585
R1613 gnd.n7014 gnd.n7013 585
R1614 gnd.n7015 gnd.n7014 585
R1615 gnd.n480 gnd.n479 585
R1616 gnd.n479 gnd.n478 585
R1617 gnd.n7009 gnd.n7008 585
R1618 gnd.n7008 gnd.n7007 585
R1619 gnd.n483 gnd.n482 585
R1620 gnd.n7006 gnd.n483 585
R1621 gnd.n7004 gnd.n7003 585
R1622 gnd.n7005 gnd.n7004 585
R1623 gnd.n486 gnd.n485 585
R1624 gnd.n485 gnd.n484 585
R1625 gnd.n6999 gnd.n6998 585
R1626 gnd.n6998 gnd.n6997 585
R1627 gnd.n489 gnd.n488 585
R1628 gnd.n6996 gnd.n489 585
R1629 gnd.n6994 gnd.n6993 585
R1630 gnd.n6995 gnd.n6994 585
R1631 gnd.n492 gnd.n491 585
R1632 gnd.n491 gnd.n490 585
R1633 gnd.n6989 gnd.n6988 585
R1634 gnd.n6988 gnd.n6987 585
R1635 gnd.n495 gnd.n494 585
R1636 gnd.n6986 gnd.n495 585
R1637 gnd.n6984 gnd.n6983 585
R1638 gnd.n6985 gnd.n6984 585
R1639 gnd.n498 gnd.n497 585
R1640 gnd.n497 gnd.n496 585
R1641 gnd.n6979 gnd.n6978 585
R1642 gnd.n6978 gnd.n6977 585
R1643 gnd.n501 gnd.n500 585
R1644 gnd.n6976 gnd.n501 585
R1645 gnd.n6974 gnd.n6973 585
R1646 gnd.n6975 gnd.n6974 585
R1647 gnd.n504 gnd.n503 585
R1648 gnd.n503 gnd.n502 585
R1649 gnd.n6969 gnd.n6968 585
R1650 gnd.n6968 gnd.n6967 585
R1651 gnd.n507 gnd.n506 585
R1652 gnd.n6966 gnd.n507 585
R1653 gnd.n6964 gnd.n6963 585
R1654 gnd.n6965 gnd.n6964 585
R1655 gnd.n510 gnd.n509 585
R1656 gnd.n509 gnd.n508 585
R1657 gnd.n6959 gnd.n6958 585
R1658 gnd.n6958 gnd.n6957 585
R1659 gnd.n513 gnd.n512 585
R1660 gnd.n6956 gnd.n513 585
R1661 gnd.n6954 gnd.n6953 585
R1662 gnd.n6955 gnd.n6954 585
R1663 gnd.n516 gnd.n515 585
R1664 gnd.n515 gnd.n514 585
R1665 gnd.n6949 gnd.n6948 585
R1666 gnd.n6948 gnd.n6947 585
R1667 gnd.n519 gnd.n518 585
R1668 gnd.n6946 gnd.n519 585
R1669 gnd.n6944 gnd.n6943 585
R1670 gnd.n6945 gnd.n6944 585
R1671 gnd.n522 gnd.n521 585
R1672 gnd.n521 gnd.n520 585
R1673 gnd.n6939 gnd.n6938 585
R1674 gnd.n6938 gnd.n6937 585
R1675 gnd.n525 gnd.n524 585
R1676 gnd.n6936 gnd.n525 585
R1677 gnd.n6934 gnd.n6933 585
R1678 gnd.n6935 gnd.n6934 585
R1679 gnd.n528 gnd.n527 585
R1680 gnd.n527 gnd.n526 585
R1681 gnd.n6929 gnd.n6928 585
R1682 gnd.n6928 gnd.n6927 585
R1683 gnd.n531 gnd.n530 585
R1684 gnd.n6926 gnd.n531 585
R1685 gnd.n6924 gnd.n6923 585
R1686 gnd.n6925 gnd.n6924 585
R1687 gnd.n534 gnd.n533 585
R1688 gnd.n533 gnd.n532 585
R1689 gnd.n6919 gnd.n6918 585
R1690 gnd.n6918 gnd.n6917 585
R1691 gnd.n537 gnd.n536 585
R1692 gnd.n6916 gnd.n537 585
R1693 gnd.n6914 gnd.n6913 585
R1694 gnd.n6915 gnd.n6914 585
R1695 gnd.n540 gnd.n539 585
R1696 gnd.n539 gnd.n538 585
R1697 gnd.n6909 gnd.n6908 585
R1698 gnd.n6908 gnd.n6907 585
R1699 gnd.n543 gnd.n542 585
R1700 gnd.n6906 gnd.n543 585
R1701 gnd.n6904 gnd.n6903 585
R1702 gnd.n6905 gnd.n6904 585
R1703 gnd.n6198 gnd.n6197 585
R1704 gnd.n6199 gnd.n6198 585
R1705 gnd.n1127 gnd.n1126 585
R1706 gnd.n6192 gnd.n1127 585
R1707 gnd.n6207 gnd.n6206 585
R1708 gnd.n6206 gnd.n6205 585
R1709 gnd.n6208 gnd.n1122 585
R1710 gnd.n4398 gnd.n1122 585
R1711 gnd.n6210 gnd.n6209 585
R1712 gnd.n6211 gnd.n6210 585
R1713 gnd.n1107 gnd.n1106 585
R1714 gnd.n4392 gnd.n1107 585
R1715 gnd.n6219 gnd.n6218 585
R1716 gnd.n6218 gnd.n6217 585
R1717 gnd.n6220 gnd.n1102 585
R1718 gnd.n4409 gnd.n1102 585
R1719 gnd.n6222 gnd.n6221 585
R1720 gnd.n6223 gnd.n6222 585
R1721 gnd.n1086 gnd.n1085 585
R1722 gnd.n4385 gnd.n1086 585
R1723 gnd.n6231 gnd.n6230 585
R1724 gnd.n6230 gnd.n6229 585
R1725 gnd.n6232 gnd.n1081 585
R1726 gnd.n4377 gnd.n1081 585
R1727 gnd.n6234 gnd.n6233 585
R1728 gnd.n6235 gnd.n6234 585
R1729 gnd.n1067 gnd.n1066 585
R1730 gnd.n4371 gnd.n1067 585
R1731 gnd.n6243 gnd.n6242 585
R1732 gnd.n6242 gnd.n6241 585
R1733 gnd.n6244 gnd.n1062 585
R1734 gnd.n4363 gnd.n1062 585
R1735 gnd.n6246 gnd.n6245 585
R1736 gnd.n6247 gnd.n6246 585
R1737 gnd.n1049 gnd.n1048 585
R1738 gnd.n4307 gnd.n1049 585
R1739 gnd.n6256 gnd.n6255 585
R1740 gnd.n6255 gnd.n6254 585
R1741 gnd.n6257 gnd.n1044 585
R1742 gnd.n4315 gnd.n1044 585
R1743 gnd.n6259 gnd.n6258 585
R1744 gnd.n6260 gnd.n6259 585
R1745 gnd.n1033 gnd.n1032 585
R1746 gnd.n4296 gnd.n1033 585
R1747 gnd.n6269 gnd.n6268 585
R1748 gnd.n6268 gnd.n6267 585
R1749 gnd.n6270 gnd.n1027 585
R1750 gnd.n4326 gnd.n1027 585
R1751 gnd.n6272 gnd.n6271 585
R1752 gnd.n6273 gnd.n6272 585
R1753 gnd.n1028 gnd.n1026 585
R1754 gnd.n4332 gnd.n1026 585
R1755 gnd.n1011 gnd.n1010 585
R1756 gnd.n2370 gnd.n1011 585
R1757 gnd.n6283 gnd.n6282 585
R1758 gnd.n6282 gnd.n6281 585
R1759 gnd.n6284 gnd.n1006 585
R1760 gnd.n4279 gnd.n1006 585
R1761 gnd.n6286 gnd.n6285 585
R1762 gnd.n6287 gnd.n6286 585
R1763 gnd.n990 gnd.n989 585
R1764 gnd.n4267 gnd.n990 585
R1765 gnd.n6295 gnd.n6294 585
R1766 gnd.n6294 gnd.n6293 585
R1767 gnd.n6296 gnd.n984 585
R1768 gnd.n4260 gnd.n984 585
R1769 gnd.n6298 gnd.n6297 585
R1770 gnd.n6299 gnd.n6298 585
R1771 gnd.n985 gnd.n983 585
R1772 gnd.n4252 gnd.n983 585
R1773 gnd.n4247 gnd.n971 585
R1774 gnd.n6305 gnd.n971 585
R1775 gnd.n4246 gnd.n4245 585
R1776 gnd.n4245 gnd.n967 585
R1777 gnd.n4244 gnd.n2421 585
R1778 gnd.n4244 gnd.n4243 585
R1779 gnd.n4231 gnd.n2422 585
R1780 gnd.n2434 gnd.n2422 585
R1781 gnd.n4233 gnd.n4232 585
R1782 gnd.n4234 gnd.n4233 585
R1783 gnd.n2436 gnd.n2435 585
R1784 gnd.n2435 gnd.n2431 585
R1785 gnd.n4092 gnd.n2444 585
R1786 gnd.n4220 gnd.n2444 585
R1787 gnd.n4091 gnd.n4090 585
R1788 gnd.n4090 gnd.n2442 585
R1789 gnd.n4089 gnd.n4088 585
R1790 gnd.n4087 gnd.n4086 585
R1791 gnd.n4085 gnd.n4084 585
R1792 gnd.n4083 gnd.n4082 585
R1793 gnd.n4081 gnd.n4080 585
R1794 gnd.n4079 gnd.n4078 585
R1795 gnd.n4077 gnd.n4076 585
R1796 gnd.n4075 gnd.n4074 585
R1797 gnd.n4073 gnd.n4072 585
R1798 gnd.n4071 gnd.n4070 585
R1799 gnd.n4069 gnd.n4068 585
R1800 gnd.n4067 gnd.n4066 585
R1801 gnd.n4065 gnd.n4064 585
R1802 gnd.n4063 gnd.n4062 585
R1803 gnd.n4061 gnd.n4060 585
R1804 gnd.n4059 gnd.n4058 585
R1805 gnd.n4057 gnd.n4056 585
R1806 gnd.n4033 gnd.n4030 585
R1807 gnd.n4052 gnd.n3949 585
R1808 gnd.n4211 gnd.n3949 585
R1809 gnd.n6119 gnd.n6118 585
R1810 gnd.n6120 gnd.n1242 585
R1811 gnd.n6121 gnd.n1237 585
R1812 gnd.n1255 gnd.n1226 585
R1813 gnd.n6128 gnd.n1225 585
R1814 gnd.n6129 gnd.n1224 585
R1815 gnd.n1252 gnd.n1218 585
R1816 gnd.n6136 gnd.n1217 585
R1817 gnd.n6137 gnd.n1216 585
R1818 gnd.n1250 gnd.n1208 585
R1819 gnd.n6144 gnd.n1207 585
R1820 gnd.n6145 gnd.n1206 585
R1821 gnd.n1247 gnd.n1200 585
R1822 gnd.n6152 gnd.n1199 585
R1823 gnd.n6153 gnd.n1198 585
R1824 gnd.n1245 gnd.n1190 585
R1825 gnd.n6160 gnd.n1189 585
R1826 gnd.n6161 gnd.n1188 585
R1827 gnd.n1187 gnd.n1142 585
R1828 gnd.n6116 gnd.n1142 585
R1829 gnd.n1147 gnd.n1140 585
R1830 gnd.n6199 gnd.n1140 585
R1831 gnd.n6191 gnd.n6190 585
R1832 gnd.n6192 gnd.n6191 585
R1833 gnd.n1146 gnd.n1130 585
R1834 gnd.n6205 gnd.n1130 585
R1835 gnd.n4401 gnd.n4399 585
R1836 gnd.n4399 gnd.n4398 585
R1837 gnd.n4402 gnd.n1120 585
R1838 gnd.n6211 gnd.n1120 585
R1839 gnd.n4403 gnd.n2344 585
R1840 gnd.n4392 gnd.n2344 585
R1841 gnd.n2341 gnd.n1109 585
R1842 gnd.n6217 gnd.n1109 585
R1843 gnd.n4408 gnd.n4407 585
R1844 gnd.n4409 gnd.n4408 585
R1845 gnd.n2340 gnd.n1100 585
R1846 gnd.n6223 gnd.n1100 585
R1847 gnd.n4384 gnd.n4383 585
R1848 gnd.n4385 gnd.n4384 585
R1849 gnd.n2347 gnd.n1089 585
R1850 gnd.n6229 gnd.n1089 585
R1851 gnd.n4379 gnd.n4378 585
R1852 gnd.n4378 gnd.n4377 585
R1853 gnd.n2349 gnd.n1080 585
R1854 gnd.n6235 gnd.n1080 585
R1855 gnd.n4370 gnd.n4369 585
R1856 gnd.n4371 gnd.n4370 585
R1857 gnd.n2353 gnd.n1069 585
R1858 gnd.n6241 gnd.n1069 585
R1859 gnd.n4365 gnd.n4364 585
R1860 gnd.n4364 gnd.n4363 585
R1861 gnd.n2355 gnd.n1060 585
R1862 gnd.n6247 gnd.n1060 585
R1863 gnd.n4309 gnd.n4308 585
R1864 gnd.n4308 gnd.n4307 585
R1865 gnd.n2390 gnd.n1052 585
R1866 gnd.n6254 gnd.n1052 585
R1867 gnd.n4314 gnd.n4313 585
R1868 gnd.n4315 gnd.n4314 585
R1869 gnd.n2389 gnd.n1043 585
R1870 gnd.n6260 gnd.n1043 585
R1871 gnd.n4295 gnd.n4294 585
R1872 gnd.n4296 gnd.n4295 585
R1873 gnd.n2377 gnd.n1035 585
R1874 gnd.n6267 gnd.n1035 585
R1875 gnd.n4328 gnd.n4327 585
R1876 gnd.n4327 gnd.n4326 585
R1877 gnd.n4329 gnd.n1024 585
R1878 gnd.n6273 gnd.n1024 585
R1879 gnd.n4331 gnd.n4330 585
R1880 gnd.n4332 gnd.n4331 585
R1881 gnd.n2373 gnd.n2372 585
R1882 gnd.n2372 gnd.n2370 585
R1883 gnd.n4275 gnd.n1013 585
R1884 gnd.n6281 gnd.n1013 585
R1885 gnd.n4277 gnd.n4276 585
R1886 gnd.n4279 gnd.n4277 585
R1887 gnd.n2393 gnd.n1004 585
R1888 gnd.n6287 gnd.n1004 585
R1889 gnd.n4269 gnd.n4268 585
R1890 gnd.n4268 gnd.n4267 585
R1891 gnd.n2395 gnd.n993 585
R1892 gnd.n6293 gnd.n993 585
R1893 gnd.n4259 gnd.n4258 585
R1894 gnd.n4260 gnd.n4259 585
R1895 gnd.n2416 gnd.n982 585
R1896 gnd.n6299 gnd.n982 585
R1897 gnd.n4254 gnd.n4253 585
R1898 gnd.n4253 gnd.n4252 585
R1899 gnd.n2418 gnd.n969 585
R1900 gnd.n6305 gnd.n969 585
R1901 gnd.n4041 gnd.n4040 585
R1902 gnd.n4040 gnd.n967 585
R1903 gnd.n4042 gnd.n2425 585
R1904 gnd.n4243 gnd.n2425 585
R1905 gnd.n4044 gnd.n4043 585
R1906 gnd.n4043 gnd.n2434 585
R1907 gnd.n4045 gnd.n2433 585
R1908 gnd.n4234 gnd.n2433 585
R1909 gnd.n4047 gnd.n4046 585
R1910 gnd.n4046 gnd.n2431 585
R1911 gnd.n4048 gnd.n2443 585
R1912 gnd.n4220 gnd.n2443 585
R1913 gnd.n4050 gnd.n4049 585
R1914 gnd.n4049 gnd.n2442 585
R1915 gnd.n3819 gnd.n3818 585
R1916 gnd.n3820 gnd.n3819 585
R1917 gnd.n2526 gnd.n2525 585
R1918 gnd.n2532 gnd.n2525 585
R1919 gnd.n3794 gnd.n2544 585
R1920 gnd.n2544 gnd.n2531 585
R1921 gnd.n3796 gnd.n3795 585
R1922 gnd.n3797 gnd.n3796 585
R1923 gnd.n2545 gnd.n2543 585
R1924 gnd.n2543 gnd.n2539 585
R1925 gnd.n3528 gnd.n3527 585
R1926 gnd.n3527 gnd.n3526 585
R1927 gnd.n2550 gnd.n2549 585
R1928 gnd.n3497 gnd.n2550 585
R1929 gnd.n3517 gnd.n3516 585
R1930 gnd.n3516 gnd.n3515 585
R1931 gnd.n2557 gnd.n2556 585
R1932 gnd.n3503 gnd.n2557 585
R1933 gnd.n3473 gnd.n2577 585
R1934 gnd.n2577 gnd.n2576 585
R1935 gnd.n3475 gnd.n3474 585
R1936 gnd.n3476 gnd.n3475 585
R1937 gnd.n2578 gnd.n2575 585
R1938 gnd.n2586 gnd.n2575 585
R1939 gnd.n3451 gnd.n2598 585
R1940 gnd.n2598 gnd.n2585 585
R1941 gnd.n3453 gnd.n3452 585
R1942 gnd.n3454 gnd.n3453 585
R1943 gnd.n2599 gnd.n2597 585
R1944 gnd.n2597 gnd.n2593 585
R1945 gnd.n3439 gnd.n3438 585
R1946 gnd.n3438 gnd.n3437 585
R1947 gnd.n2604 gnd.n2603 585
R1948 gnd.n2614 gnd.n2604 585
R1949 gnd.n3428 gnd.n3427 585
R1950 gnd.n3427 gnd.n3426 585
R1951 gnd.n2611 gnd.n2610 585
R1952 gnd.n3414 gnd.n2611 585
R1953 gnd.n3388 gnd.n2632 585
R1954 gnd.n2632 gnd.n2621 585
R1955 gnd.n3390 gnd.n3389 585
R1956 gnd.n3391 gnd.n3390 585
R1957 gnd.n2633 gnd.n2631 585
R1958 gnd.n2641 gnd.n2631 585
R1959 gnd.n3366 gnd.n2653 585
R1960 gnd.n2653 gnd.n2640 585
R1961 gnd.n3368 gnd.n3367 585
R1962 gnd.n3369 gnd.n3368 585
R1963 gnd.n2654 gnd.n2652 585
R1964 gnd.n2652 gnd.n2648 585
R1965 gnd.n3354 gnd.n3353 585
R1966 gnd.n3353 gnd.n3352 585
R1967 gnd.n2659 gnd.n2658 585
R1968 gnd.n2668 gnd.n2659 585
R1969 gnd.n3343 gnd.n3342 585
R1970 gnd.n3342 gnd.n3341 585
R1971 gnd.n2666 gnd.n2665 585
R1972 gnd.n3329 gnd.n2666 585
R1973 gnd.n2767 gnd.n2766 585
R1974 gnd.n2767 gnd.n2675 585
R1975 gnd.n3286 gnd.n3285 585
R1976 gnd.n3285 gnd.n3284 585
R1977 gnd.n3287 gnd.n2761 585
R1978 gnd.n2772 gnd.n2761 585
R1979 gnd.n3289 gnd.n3288 585
R1980 gnd.n3290 gnd.n3289 585
R1981 gnd.n2762 gnd.n2760 585
R1982 gnd.n2785 gnd.n2760 585
R1983 gnd.n2745 gnd.n2744 585
R1984 gnd.n2748 gnd.n2745 585
R1985 gnd.n3300 gnd.n3299 585
R1986 gnd.n3299 gnd.n3298 585
R1987 gnd.n3301 gnd.n2739 585
R1988 gnd.n3260 gnd.n2739 585
R1989 gnd.n3303 gnd.n3302 585
R1990 gnd.n3304 gnd.n3303 585
R1991 gnd.n2740 gnd.n2738 585
R1992 gnd.n2799 gnd.n2738 585
R1993 gnd.n3252 gnd.n3251 585
R1994 gnd.n3251 gnd.n3250 585
R1995 gnd.n2796 gnd.n2795 585
R1996 gnd.n3234 gnd.n2796 585
R1997 gnd.n3221 gnd.n2815 585
R1998 gnd.n2815 gnd.n2814 585
R1999 gnd.n3223 gnd.n3222 585
R2000 gnd.n3224 gnd.n3223 585
R2001 gnd.n2816 gnd.n2813 585
R2002 gnd.n2822 gnd.n2813 585
R2003 gnd.n3202 gnd.n3201 585
R2004 gnd.n3203 gnd.n3202 585
R2005 gnd.n2833 gnd.n2832 585
R2006 gnd.n2832 gnd.n2828 585
R2007 gnd.n3192 gnd.n3191 585
R2008 gnd.n3193 gnd.n3192 585
R2009 gnd.n2843 gnd.n2842 585
R2010 gnd.n2848 gnd.n2842 585
R2011 gnd.n3170 gnd.n2861 585
R2012 gnd.n2861 gnd.n2847 585
R2013 gnd.n3172 gnd.n3171 585
R2014 gnd.n3173 gnd.n3172 585
R2015 gnd.n2862 gnd.n2860 585
R2016 gnd.n2860 gnd.n2856 585
R2017 gnd.n3161 gnd.n3160 585
R2018 gnd.n3162 gnd.n3161 585
R2019 gnd.n2869 gnd.n2868 585
R2020 gnd.n2873 gnd.n2868 585
R2021 gnd.n3138 gnd.n2890 585
R2022 gnd.n2890 gnd.n2872 585
R2023 gnd.n3140 gnd.n3139 585
R2024 gnd.n3141 gnd.n3140 585
R2025 gnd.n2891 gnd.n2889 585
R2026 gnd.n2889 gnd.n2880 585
R2027 gnd.n3133 gnd.n3132 585
R2028 gnd.n3132 gnd.n3131 585
R2029 gnd.n2938 gnd.n2937 585
R2030 gnd.n2939 gnd.n2938 585
R2031 gnd.n3092 gnd.n3091 585
R2032 gnd.n3093 gnd.n3092 585
R2033 gnd.n2948 gnd.n2947 585
R2034 gnd.n2947 gnd.n2946 585
R2035 gnd.n3087 gnd.n3086 585
R2036 gnd.n3086 gnd.n3085 585
R2037 gnd.n2951 gnd.n2950 585
R2038 gnd.n2952 gnd.n2951 585
R2039 gnd.n3076 gnd.n3075 585
R2040 gnd.n3077 gnd.n3076 585
R2041 gnd.n2959 gnd.n2958 585
R2042 gnd.n3068 gnd.n2958 585
R2043 gnd.n3071 gnd.n3070 585
R2044 gnd.n3070 gnd.n3069 585
R2045 gnd.n2962 gnd.n2961 585
R2046 gnd.n2963 gnd.n2962 585
R2047 gnd.n3057 gnd.n3056 585
R2048 gnd.n3055 gnd.n2981 585
R2049 gnd.n3054 gnd.n2980 585
R2050 gnd.n3059 gnd.n2980 585
R2051 gnd.n3053 gnd.n3052 585
R2052 gnd.n3051 gnd.n3050 585
R2053 gnd.n3049 gnd.n3048 585
R2054 gnd.n3047 gnd.n3046 585
R2055 gnd.n3045 gnd.n3044 585
R2056 gnd.n3043 gnd.n3042 585
R2057 gnd.n3041 gnd.n3040 585
R2058 gnd.n3039 gnd.n3038 585
R2059 gnd.n3037 gnd.n3036 585
R2060 gnd.n3035 gnd.n3034 585
R2061 gnd.n3033 gnd.n3032 585
R2062 gnd.n3031 gnd.n3030 585
R2063 gnd.n3029 gnd.n3028 585
R2064 gnd.n3027 gnd.n3026 585
R2065 gnd.n3025 gnd.n3024 585
R2066 gnd.n3023 gnd.n3022 585
R2067 gnd.n3021 gnd.n3020 585
R2068 gnd.n3019 gnd.n3018 585
R2069 gnd.n3017 gnd.n3016 585
R2070 gnd.n3015 gnd.n3014 585
R2071 gnd.n3013 gnd.n3012 585
R2072 gnd.n3011 gnd.n3010 585
R2073 gnd.n2968 gnd.n2967 585
R2074 gnd.n3062 gnd.n3061 585
R2075 gnd.n3823 gnd.n3822 585
R2076 gnd.n3825 gnd.n3824 585
R2077 gnd.n3827 gnd.n3826 585
R2078 gnd.n3829 gnd.n3828 585
R2079 gnd.n3831 gnd.n3830 585
R2080 gnd.n3833 gnd.n3832 585
R2081 gnd.n3835 gnd.n3834 585
R2082 gnd.n3837 gnd.n3836 585
R2083 gnd.n3839 gnd.n3838 585
R2084 gnd.n3841 gnd.n3840 585
R2085 gnd.n3843 gnd.n3842 585
R2086 gnd.n3845 gnd.n3844 585
R2087 gnd.n3847 gnd.n3846 585
R2088 gnd.n3849 gnd.n3848 585
R2089 gnd.n3851 gnd.n3850 585
R2090 gnd.n3853 gnd.n3852 585
R2091 gnd.n3855 gnd.n3854 585
R2092 gnd.n3857 gnd.n3856 585
R2093 gnd.n3859 gnd.n3858 585
R2094 gnd.n3861 gnd.n3860 585
R2095 gnd.n3863 gnd.n3862 585
R2096 gnd.n3865 gnd.n3864 585
R2097 gnd.n3867 gnd.n3866 585
R2098 gnd.n3869 gnd.n3868 585
R2099 gnd.n3871 gnd.n3870 585
R2100 gnd.n3872 gnd.n2493 585
R2101 gnd.n3873 gnd.n2451 585
R2102 gnd.n3911 gnd.n2451 585
R2103 gnd.n3821 gnd.n2523 585
R2104 gnd.n3821 gnd.n3820 585
R2105 gnd.n3490 gnd.n2522 585
R2106 gnd.n2532 gnd.n2522 585
R2107 gnd.n3492 gnd.n3491 585
R2108 gnd.n3491 gnd.n2531 585
R2109 gnd.n3493 gnd.n2541 585
R2110 gnd.n3797 gnd.n2541 585
R2111 gnd.n3495 gnd.n3494 585
R2112 gnd.n3494 gnd.n2539 585
R2113 gnd.n3496 gnd.n2552 585
R2114 gnd.n3526 gnd.n2552 585
R2115 gnd.n3499 gnd.n3498 585
R2116 gnd.n3498 gnd.n3497 585
R2117 gnd.n3500 gnd.n2559 585
R2118 gnd.n3515 gnd.n2559 585
R2119 gnd.n3502 gnd.n3501 585
R2120 gnd.n3503 gnd.n3502 585
R2121 gnd.n2569 gnd.n2568 585
R2122 gnd.n2576 gnd.n2568 585
R2123 gnd.n3478 gnd.n3477 585
R2124 gnd.n3477 gnd.n3476 585
R2125 gnd.n2572 gnd.n2571 585
R2126 gnd.n2586 gnd.n2572 585
R2127 gnd.n3404 gnd.n3403 585
R2128 gnd.n3403 gnd.n2585 585
R2129 gnd.n3405 gnd.n2595 585
R2130 gnd.n3454 gnd.n2595 585
R2131 gnd.n3407 gnd.n3406 585
R2132 gnd.n3406 gnd.n2593 585
R2133 gnd.n3408 gnd.n2606 585
R2134 gnd.n3437 gnd.n2606 585
R2135 gnd.n3410 gnd.n3409 585
R2136 gnd.n3409 gnd.n2614 585
R2137 gnd.n3411 gnd.n2613 585
R2138 gnd.n3426 gnd.n2613 585
R2139 gnd.n3413 gnd.n3412 585
R2140 gnd.n3414 gnd.n3413 585
R2141 gnd.n2625 gnd.n2624 585
R2142 gnd.n2624 gnd.n2621 585
R2143 gnd.n3393 gnd.n3392 585
R2144 gnd.n3392 gnd.n3391 585
R2145 gnd.n2628 gnd.n2627 585
R2146 gnd.n2641 gnd.n2628 585
R2147 gnd.n3317 gnd.n3316 585
R2148 gnd.n3316 gnd.n2640 585
R2149 gnd.n3318 gnd.n2650 585
R2150 gnd.n3369 gnd.n2650 585
R2151 gnd.n3320 gnd.n3319 585
R2152 gnd.n3319 gnd.n2648 585
R2153 gnd.n3321 gnd.n2661 585
R2154 gnd.n3352 gnd.n2661 585
R2155 gnd.n3323 gnd.n3322 585
R2156 gnd.n3322 gnd.n2668 585
R2157 gnd.n3324 gnd.n2667 585
R2158 gnd.n3341 gnd.n2667 585
R2159 gnd.n3326 gnd.n3325 585
R2160 gnd.n3329 gnd.n3326 585
R2161 gnd.n2678 gnd.n2677 585
R2162 gnd.n2677 gnd.n2675 585
R2163 gnd.n2769 gnd.n2768 585
R2164 gnd.n3284 gnd.n2768 585
R2165 gnd.n2771 gnd.n2770 585
R2166 gnd.n2772 gnd.n2771 585
R2167 gnd.n2782 gnd.n2758 585
R2168 gnd.n3290 gnd.n2758 585
R2169 gnd.n2784 gnd.n2783 585
R2170 gnd.n2785 gnd.n2784 585
R2171 gnd.n2781 gnd.n2780 585
R2172 gnd.n2781 gnd.n2748 585
R2173 gnd.n2779 gnd.n2746 585
R2174 gnd.n3298 gnd.n2746 585
R2175 gnd.n2735 gnd.n2733 585
R2176 gnd.n3260 gnd.n2735 585
R2177 gnd.n3306 gnd.n3305 585
R2178 gnd.n3305 gnd.n3304 585
R2179 gnd.n2734 gnd.n2732 585
R2180 gnd.n2799 gnd.n2734 585
R2181 gnd.n3231 gnd.n2798 585
R2182 gnd.n3250 gnd.n2798 585
R2183 gnd.n3233 gnd.n3232 585
R2184 gnd.n3234 gnd.n3233 585
R2185 gnd.n2808 gnd.n2807 585
R2186 gnd.n2814 gnd.n2807 585
R2187 gnd.n3226 gnd.n3225 585
R2188 gnd.n3225 gnd.n3224 585
R2189 gnd.n2811 gnd.n2810 585
R2190 gnd.n2822 gnd.n2811 585
R2191 gnd.n3111 gnd.n2830 585
R2192 gnd.n3203 gnd.n2830 585
R2193 gnd.n3113 gnd.n3112 585
R2194 gnd.n3112 gnd.n2828 585
R2195 gnd.n3114 gnd.n2841 585
R2196 gnd.n3193 gnd.n2841 585
R2197 gnd.n3116 gnd.n3115 585
R2198 gnd.n3116 gnd.n2848 585
R2199 gnd.n3118 gnd.n3117 585
R2200 gnd.n3117 gnd.n2847 585
R2201 gnd.n3119 gnd.n2858 585
R2202 gnd.n3173 gnd.n2858 585
R2203 gnd.n3121 gnd.n3120 585
R2204 gnd.n3120 gnd.n2856 585
R2205 gnd.n3122 gnd.n2867 585
R2206 gnd.n3162 gnd.n2867 585
R2207 gnd.n3124 gnd.n3123 585
R2208 gnd.n3124 gnd.n2873 585
R2209 gnd.n3126 gnd.n3125 585
R2210 gnd.n3125 gnd.n2872 585
R2211 gnd.n3127 gnd.n2888 585
R2212 gnd.n3141 gnd.n2888 585
R2213 gnd.n3128 gnd.n2941 585
R2214 gnd.n2941 gnd.n2880 585
R2215 gnd.n3130 gnd.n3129 585
R2216 gnd.n3131 gnd.n3130 585
R2217 gnd.n2942 gnd.n2940 585
R2218 gnd.n2940 gnd.n2939 585
R2219 gnd.n3095 gnd.n3094 585
R2220 gnd.n3094 gnd.n3093 585
R2221 gnd.n2945 gnd.n2944 585
R2222 gnd.n2946 gnd.n2945 585
R2223 gnd.n3084 gnd.n3083 585
R2224 gnd.n3085 gnd.n3084 585
R2225 gnd.n2954 gnd.n2953 585
R2226 gnd.n2953 gnd.n2952 585
R2227 gnd.n3079 gnd.n3078 585
R2228 gnd.n3078 gnd.n3077 585
R2229 gnd.n2957 gnd.n2956 585
R2230 gnd.n3068 gnd.n2957 585
R2231 gnd.n3067 gnd.n3066 585
R2232 gnd.n3069 gnd.n3067 585
R2233 gnd.n2965 gnd.n2964 585
R2234 gnd.n2964 gnd.n2963 585
R2235 gnd.n7282 gnd.n7281 585
R2236 gnd.n7283 gnd.n7282 585
R2237 gnd.n158 gnd.n157 585
R2238 gnd.n167 gnd.n158 585
R2239 gnd.n7291 gnd.n7290 585
R2240 gnd.n7290 gnd.n7289 585
R2241 gnd.n7292 gnd.n153 585
R2242 gnd.n153 gnd.n152 585
R2243 gnd.n7294 gnd.n7293 585
R2244 gnd.n7295 gnd.n7294 585
R2245 gnd.n137 gnd.n136 585
R2246 gnd.n141 gnd.n137 585
R2247 gnd.n7303 gnd.n7302 585
R2248 gnd.n7302 gnd.n7301 585
R2249 gnd.n7304 gnd.n132 585
R2250 gnd.n7266 gnd.n132 585
R2251 gnd.n7306 gnd.n7305 585
R2252 gnd.n7307 gnd.n7306 585
R2253 gnd.n116 gnd.n115 585
R2254 gnd.n7174 gnd.n116 585
R2255 gnd.n7315 gnd.n7314 585
R2256 gnd.n7314 gnd.n7313 585
R2257 gnd.n7316 gnd.n111 585
R2258 gnd.n7167 gnd.n111 585
R2259 gnd.n7318 gnd.n7317 585
R2260 gnd.n7319 gnd.n7318 585
R2261 gnd.n97 gnd.n96 585
R2262 gnd.n7159 gnd.n97 585
R2263 gnd.n7327 gnd.n7326 585
R2264 gnd.n7326 gnd.n7325 585
R2265 gnd.n7328 gnd.n91 585
R2266 gnd.n7152 gnd.n91 585
R2267 gnd.n7330 gnd.n7329 585
R2268 gnd.n7331 gnd.n7330 585
R2269 gnd.n92 gnd.n90 585
R2270 gnd.n7144 gnd.n90 585
R2271 gnd.n7139 gnd.n7138 585
R2272 gnd.n7138 gnd.n7137 585
R2273 gnd.n401 gnd.n72 585
R2274 gnd.n7339 gnd.n72 585
R2275 gnd.n5789 gnd.n1723 585
R2276 gnd.n5785 gnd.n1723 585
R2277 gnd.n5791 gnd.n5790 585
R2278 gnd.n5792 gnd.n5791 585
R2279 gnd.n1724 gnd.n1710 585
R2280 gnd.n5797 gnd.n1710 585
R2281 gnd.n5779 gnd.n5778 585
R2282 gnd.n5778 gnd.n1706 585
R2283 gnd.n5777 gnd.n5776 585
R2284 gnd.n5777 gnd.n1699 585
R2285 gnd.n1689 gnd.n1688 585
R2286 gnd.n5806 gnd.n1689 585
R2287 gnd.n5812 gnd.n5811 585
R2288 gnd.n5811 gnd.n5810 585
R2289 gnd.n5813 gnd.n1684 585
R2290 gnd.n5767 gnd.n1684 585
R2291 gnd.n5815 gnd.n5814 585
R2292 gnd.n5816 gnd.n5815 585
R2293 gnd.n1670 gnd.n1669 585
R2294 gnd.n5749 gnd.n1670 585
R2295 gnd.n5824 gnd.n5823 585
R2296 gnd.n5823 gnd.n5822 585
R2297 gnd.n5825 gnd.n1665 585
R2298 gnd.n5742 gnd.n1665 585
R2299 gnd.n5827 gnd.n5826 585
R2300 gnd.n5828 gnd.n5827 585
R2301 gnd.n1649 gnd.n1648 585
R2302 gnd.n5686 gnd.n1649 585
R2303 gnd.n5836 gnd.n5835 585
R2304 gnd.n5835 gnd.n5834 585
R2305 gnd.n5837 gnd.n1644 585
R2306 gnd.n5697 gnd.n1644 585
R2307 gnd.n5839 gnd.n5838 585
R2308 gnd.n5840 gnd.n5839 585
R2309 gnd.n1629 gnd.n1628 585
R2310 gnd.n5677 gnd.n1629 585
R2311 gnd.n5848 gnd.n5847 585
R2312 gnd.n5847 gnd.n5846 585
R2313 gnd.n5849 gnd.n1623 585
R2314 gnd.n5669 gnd.n1623 585
R2315 gnd.n5851 gnd.n5850 585
R2316 gnd.n5852 gnd.n5851 585
R2317 gnd.n1624 gnd.n1622 585
R2318 gnd.n5121 gnd.n1622 585
R2319 gnd.n5662 gnd.n1610 585
R2320 gnd.n5858 gnd.n1610 585
R2321 gnd.n5207 gnd.n5206 585
R2322 gnd.n5171 gnd.n5170 585
R2323 gnd.n5221 gnd.n5220 585
R2324 gnd.n5223 gnd.n5169 585
R2325 gnd.n5226 gnd.n5225 585
R2326 gnd.n5162 gnd.n5161 585
R2327 gnd.n5240 gnd.n5239 585
R2328 gnd.n5242 gnd.n5160 585
R2329 gnd.n5245 gnd.n5244 585
R2330 gnd.n5153 gnd.n5152 585
R2331 gnd.n5259 gnd.n5258 585
R2332 gnd.n5261 gnd.n5151 585
R2333 gnd.n5264 gnd.n5263 585
R2334 gnd.n5144 gnd.n5143 585
R2335 gnd.n5279 gnd.n5278 585
R2336 gnd.n5281 gnd.n5142 585
R2337 gnd.n5284 gnd.n5283 585
R2338 gnd.n5285 gnd.n5139 585
R2339 gnd.n5138 gnd.n5137 585
R2340 gnd.n5138 gnd.n1598 585
R2341 gnd.n7251 gnd.n7250 585
R2342 gnd.n7248 gnd.n7189 585
R2343 gnd.n7247 gnd.n7246 585
R2344 gnd.n7240 gnd.n7191 585
R2345 gnd.n7242 gnd.n7241 585
R2346 gnd.n7238 gnd.n7193 585
R2347 gnd.n7237 gnd.n7236 585
R2348 gnd.n7230 gnd.n7195 585
R2349 gnd.n7232 gnd.n7231 585
R2350 gnd.n7228 gnd.n7197 585
R2351 gnd.n7227 gnd.n7226 585
R2352 gnd.n7220 gnd.n7199 585
R2353 gnd.n7222 gnd.n7221 585
R2354 gnd.n7218 gnd.n7201 585
R2355 gnd.n7217 gnd.n7216 585
R2356 gnd.n7210 gnd.n7203 585
R2357 gnd.n7212 gnd.n7211 585
R2358 gnd.n7208 gnd.n7207 585
R2359 gnd.n7206 gnd.n171 585
R2360 gnd.n171 gnd.n170 585
R2361 gnd.n7254 gnd.n169 585
R2362 gnd.n7283 gnd.n169 585
R2363 gnd.n7256 gnd.n7255 585
R2364 gnd.n7255 gnd.n167 585
R2365 gnd.n7257 gnd.n160 585
R2366 gnd.n7289 gnd.n160 585
R2367 gnd.n7259 gnd.n7258 585
R2368 gnd.n7258 gnd.n152 585
R2369 gnd.n7260 gnd.n151 585
R2370 gnd.n7295 gnd.n151 585
R2371 gnd.n7262 gnd.n7261 585
R2372 gnd.n7261 gnd.n141 585
R2373 gnd.n7263 gnd.n140 585
R2374 gnd.n7301 gnd.n140 585
R2375 gnd.n7265 gnd.n7264 585
R2376 gnd.n7266 gnd.n7265 585
R2377 gnd.n387 gnd.n130 585
R2378 gnd.n7307 gnd.n130 585
R2379 gnd.n7176 gnd.n7175 585
R2380 gnd.n7175 gnd.n7174 585
R2381 gnd.n389 gnd.n119 585
R2382 gnd.n7313 gnd.n119 585
R2383 gnd.n7166 gnd.n7165 585
R2384 gnd.n7167 gnd.n7166 585
R2385 gnd.n392 gnd.n110 585
R2386 gnd.n7319 gnd.n110 585
R2387 gnd.n7161 gnd.n7160 585
R2388 gnd.n7160 gnd.n7159 585
R2389 gnd.n394 gnd.n100 585
R2390 gnd.n7325 gnd.n100 585
R2391 gnd.n7151 gnd.n7150 585
R2392 gnd.n7152 gnd.n7151 585
R2393 gnd.n396 gnd.n88 585
R2394 gnd.n7331 gnd.n88 585
R2395 gnd.n7146 gnd.n7145 585
R2396 gnd.n7145 gnd.n7144 585
R2397 gnd.n68 gnd.n67 585
R2398 gnd.n7137 gnd.n68 585
R2399 gnd.n7341 gnd.n7340 585
R2400 gnd.n7340 gnd.n7339 585
R2401 gnd.n7342 gnd.n66 585
R2402 gnd.n5785 gnd.n66 585
R2403 gnd.n1715 gnd.n64 585
R2404 gnd.n5792 gnd.n1715 585
R2405 gnd.n5757 gnd.n1708 585
R2406 gnd.n5797 gnd.n1708 585
R2407 gnd.n5759 gnd.n5756 585
R2408 gnd.n5756 gnd.n1706 585
R2409 gnd.n5760 gnd.n5755 585
R2410 gnd.n5755 gnd.n1699 585
R2411 gnd.n5761 gnd.n1698 585
R2412 gnd.n5806 gnd.n1698 585
R2413 gnd.n1731 gnd.n1692 585
R2414 gnd.n5810 gnd.n1692 585
R2415 gnd.n5766 gnd.n5765 585
R2416 gnd.n5767 gnd.n5766 585
R2417 gnd.n1730 gnd.n1683 585
R2418 gnd.n5816 gnd.n1683 585
R2419 gnd.n5751 gnd.n5750 585
R2420 gnd.n5750 gnd.n5749 585
R2421 gnd.n1733 gnd.n1672 585
R2422 gnd.n5822 gnd.n1672 585
R2423 gnd.n5689 gnd.n1735 585
R2424 gnd.n5742 gnd.n1735 585
R2425 gnd.n5690 gnd.n1663 585
R2426 gnd.n5828 gnd.n1663 585
R2427 gnd.n5691 gnd.n5687 585
R2428 gnd.n5687 gnd.n5686 585
R2429 gnd.n1743 gnd.n1652 585
R2430 gnd.n5834 gnd.n1652 585
R2431 gnd.n5696 gnd.n5695 585
R2432 gnd.n5697 gnd.n5696 585
R2433 gnd.n1742 gnd.n1643 585
R2434 gnd.n5840 gnd.n1643 585
R2435 gnd.n5676 gnd.n5675 585
R2436 gnd.n5677 gnd.n5676 585
R2437 gnd.n1748 gnd.n1632 585
R2438 gnd.n5846 gnd.n1632 585
R2439 gnd.n5671 gnd.n5670 585
R2440 gnd.n5670 gnd.n5669 585
R2441 gnd.n1750 gnd.n1620 585
R2442 gnd.n5852 gnd.n1620 585
R2443 gnd.n5123 gnd.n5122 585
R2444 gnd.n5122 gnd.n5121 585
R2445 gnd.n5124 gnd.n1608 585
R2446 gnd.n5858 gnd.n1608 585
R2447 gnd.n3806 gnd.n2473 585
R2448 gnd.n2473 gnd.n2450 585
R2449 gnd.n3807 gnd.n2534 585
R2450 gnd.n2534 gnd.n2524 585
R2451 gnd.n3809 gnd.n3808 585
R2452 gnd.n3810 gnd.n3809 585
R2453 gnd.n2535 gnd.n2533 585
R2454 gnd.n2542 gnd.n2533 585
R2455 gnd.n3800 gnd.n3799 585
R2456 gnd.n3799 gnd.n3798 585
R2457 gnd.n2538 gnd.n2537 585
R2458 gnd.n3525 gnd.n2538 585
R2459 gnd.n3511 gnd.n2561 585
R2460 gnd.n2561 gnd.n2551 585
R2461 gnd.n3513 gnd.n3512 585
R2462 gnd.n3514 gnd.n3513 585
R2463 gnd.n2562 gnd.n2560 585
R2464 gnd.n2560 gnd.n2558 585
R2465 gnd.n3506 gnd.n3505 585
R2466 gnd.n3505 gnd.n3504 585
R2467 gnd.n2565 gnd.n2564 585
R2468 gnd.n2574 gnd.n2565 585
R2469 gnd.n3462 gnd.n2588 585
R2470 gnd.n2588 gnd.n2573 585
R2471 gnd.n3464 gnd.n3463 585
R2472 gnd.n3465 gnd.n3464 585
R2473 gnd.n2589 gnd.n2587 585
R2474 gnd.n2596 gnd.n2587 585
R2475 gnd.n3457 gnd.n3456 585
R2476 gnd.n3456 gnd.n3455 585
R2477 gnd.n2592 gnd.n2591 585
R2478 gnd.n3436 gnd.n2592 585
R2479 gnd.n3422 gnd.n2616 585
R2480 gnd.n2616 gnd.n2605 585
R2481 gnd.n3424 gnd.n3423 585
R2482 gnd.n3425 gnd.n3424 585
R2483 gnd.n2617 gnd.n2615 585
R2484 gnd.n2615 gnd.n2612 585
R2485 gnd.n3417 gnd.n3416 585
R2486 gnd.n3416 gnd.n3415 585
R2487 gnd.n2620 gnd.n2619 585
R2488 gnd.n2630 gnd.n2620 585
R2489 gnd.n3377 gnd.n2643 585
R2490 gnd.n2643 gnd.n2629 585
R2491 gnd.n3379 gnd.n3378 585
R2492 gnd.n3380 gnd.n3379 585
R2493 gnd.n2644 gnd.n2642 585
R2494 gnd.n2651 gnd.n2642 585
R2495 gnd.n3372 gnd.n3371 585
R2496 gnd.n3371 gnd.n3370 585
R2497 gnd.n2647 gnd.n2646 585
R2498 gnd.n3351 gnd.n2647 585
R2499 gnd.n3337 gnd.n2670 585
R2500 gnd.n2670 gnd.n2660 585
R2501 gnd.n3339 gnd.n3338 585
R2502 gnd.n3340 gnd.n3339 585
R2503 gnd.n2671 gnd.n2669 585
R2504 gnd.n3328 gnd.n2669 585
R2505 gnd.n3332 gnd.n3331 585
R2506 gnd.n3331 gnd.n3330 585
R2507 gnd.n2674 gnd.n2673 585
R2508 gnd.n3283 gnd.n2674 585
R2509 gnd.n2776 gnd.n2775 585
R2510 gnd.n2777 gnd.n2776 585
R2511 gnd.n2756 gnd.n2755 585
R2512 gnd.n2759 gnd.n2756 585
R2513 gnd.n3293 gnd.n3292 585
R2514 gnd.n3292 gnd.n3291 585
R2515 gnd.n3294 gnd.n2750 585
R2516 gnd.n2786 gnd.n2750 585
R2517 gnd.n3296 gnd.n3295 585
R2518 gnd.n3297 gnd.n3296 585
R2519 gnd.n2751 gnd.n2749 585
R2520 gnd.n3261 gnd.n2749 585
R2521 gnd.n3245 gnd.n3244 585
R2522 gnd.n3244 gnd.n2737 585
R2523 gnd.n3246 gnd.n2801 585
R2524 gnd.n2801 gnd.n2736 585
R2525 gnd.n3248 gnd.n3247 585
R2526 gnd.n3249 gnd.n3248 585
R2527 gnd.n2802 gnd.n2800 585
R2528 gnd.n2800 gnd.n2797 585
R2529 gnd.n3237 gnd.n3236 585
R2530 gnd.n3236 gnd.n3235 585
R2531 gnd.n2805 gnd.n2804 585
R2532 gnd.n2812 gnd.n2805 585
R2533 gnd.n3211 gnd.n3210 585
R2534 gnd.n3212 gnd.n3211 585
R2535 gnd.n2824 gnd.n2823 585
R2536 gnd.n2831 gnd.n2823 585
R2537 gnd.n3206 gnd.n3205 585
R2538 gnd.n3205 gnd.n3204 585
R2539 gnd.n2827 gnd.n2826 585
R2540 gnd.n3194 gnd.n2827 585
R2541 gnd.n3181 gnd.n2851 585
R2542 gnd.n2851 gnd.n2850 585
R2543 gnd.n3183 gnd.n3182 585
R2544 gnd.n3184 gnd.n3183 585
R2545 gnd.n2852 gnd.n2849 585
R2546 gnd.n2859 gnd.n2849 585
R2547 gnd.n3176 gnd.n3175 585
R2548 gnd.n3175 gnd.n3174 585
R2549 gnd.n2855 gnd.n2854 585
R2550 gnd.n3163 gnd.n2855 585
R2551 gnd.n3150 gnd.n2876 585
R2552 gnd.n2876 gnd.n2875 585
R2553 gnd.n3152 gnd.n3151 585
R2554 gnd.n3153 gnd.n3152 585
R2555 gnd.n3146 gnd.n2874 585
R2556 gnd.n3145 gnd.n3144 585
R2557 gnd.n2879 gnd.n2878 585
R2558 gnd.n3142 gnd.n2879 585
R2559 gnd.n2901 gnd.n2900 585
R2560 gnd.n2904 gnd.n2903 585
R2561 gnd.n2902 gnd.n2897 585
R2562 gnd.n2909 gnd.n2908 585
R2563 gnd.n2911 gnd.n2910 585
R2564 gnd.n2914 gnd.n2913 585
R2565 gnd.n2912 gnd.n2895 585
R2566 gnd.n2919 gnd.n2918 585
R2567 gnd.n2921 gnd.n2920 585
R2568 gnd.n2924 gnd.n2923 585
R2569 gnd.n2922 gnd.n2893 585
R2570 gnd.n2929 gnd.n2928 585
R2571 gnd.n2933 gnd.n2930 585
R2572 gnd.n2934 gnd.n2871 585
R2573 gnd.n3812 gnd.n2488 585
R2574 gnd.n3879 gnd.n3878 585
R2575 gnd.n3881 gnd.n3880 585
R2576 gnd.n3883 gnd.n3882 585
R2577 gnd.n3885 gnd.n3884 585
R2578 gnd.n3887 gnd.n3886 585
R2579 gnd.n3889 gnd.n3888 585
R2580 gnd.n3891 gnd.n3890 585
R2581 gnd.n3893 gnd.n3892 585
R2582 gnd.n3895 gnd.n3894 585
R2583 gnd.n3897 gnd.n3896 585
R2584 gnd.n3899 gnd.n3898 585
R2585 gnd.n3901 gnd.n3900 585
R2586 gnd.n3904 gnd.n3903 585
R2587 gnd.n3902 gnd.n2476 585
R2588 gnd.n3908 gnd.n2474 585
R2589 gnd.n3910 gnd.n3909 585
R2590 gnd.n3911 gnd.n3910 585
R2591 gnd.n3813 gnd.n2529 585
R2592 gnd.n3813 gnd.n2450 585
R2593 gnd.n3815 gnd.n3814 585
R2594 gnd.n3814 gnd.n2524 585
R2595 gnd.n3811 gnd.n2528 585
R2596 gnd.n3811 gnd.n3810 585
R2597 gnd.n3790 gnd.n2530 585
R2598 gnd.n2542 gnd.n2530 585
R2599 gnd.n3789 gnd.n2540 585
R2600 gnd.n3798 gnd.n2540 585
R2601 gnd.n3524 gnd.n2547 585
R2602 gnd.n3525 gnd.n3524 585
R2603 gnd.n3523 gnd.n3522 585
R2604 gnd.n3523 gnd.n2551 585
R2605 gnd.n3521 gnd.n2553 585
R2606 gnd.n3514 gnd.n2553 585
R2607 gnd.n2566 gnd.n2554 585
R2608 gnd.n2566 gnd.n2558 585
R2609 gnd.n3470 gnd.n2567 585
R2610 gnd.n3504 gnd.n2567 585
R2611 gnd.n3469 gnd.n3468 585
R2612 gnd.n3468 gnd.n2574 585
R2613 gnd.n3467 gnd.n2582 585
R2614 gnd.n3467 gnd.n2573 585
R2615 gnd.n3466 gnd.n2584 585
R2616 gnd.n3466 gnd.n3465 585
R2617 gnd.n3445 gnd.n2583 585
R2618 gnd.n2596 gnd.n2583 585
R2619 gnd.n3444 gnd.n2594 585
R2620 gnd.n3455 gnd.n2594 585
R2621 gnd.n3435 gnd.n2601 585
R2622 gnd.n3436 gnd.n3435 585
R2623 gnd.n3434 gnd.n3433 585
R2624 gnd.n3434 gnd.n2605 585
R2625 gnd.n3432 gnd.n2607 585
R2626 gnd.n3425 gnd.n2607 585
R2627 gnd.n2622 gnd.n2608 585
R2628 gnd.n2622 gnd.n2612 585
R2629 gnd.n3385 gnd.n2623 585
R2630 gnd.n3415 gnd.n2623 585
R2631 gnd.n3384 gnd.n3383 585
R2632 gnd.n3383 gnd.n2630 585
R2633 gnd.n3382 gnd.n2637 585
R2634 gnd.n3382 gnd.n2629 585
R2635 gnd.n3381 gnd.n2639 585
R2636 gnd.n3381 gnd.n3380 585
R2637 gnd.n3360 gnd.n2638 585
R2638 gnd.n2651 gnd.n2638 585
R2639 gnd.n3359 gnd.n2649 585
R2640 gnd.n3370 gnd.n2649 585
R2641 gnd.n3350 gnd.n2656 585
R2642 gnd.n3351 gnd.n3350 585
R2643 gnd.n3349 gnd.n3348 585
R2644 gnd.n3349 gnd.n2660 585
R2645 gnd.n3347 gnd.n2662 585
R2646 gnd.n3340 gnd.n2662 585
R2647 gnd.n3327 gnd.n2663 585
R2648 gnd.n3328 gnd.n3327 585
R2649 gnd.n3280 gnd.n2676 585
R2650 gnd.n3330 gnd.n2676 585
R2651 gnd.n3282 gnd.n3281 585
R2652 gnd.n3283 gnd.n3282 585
R2653 gnd.n3275 gnd.n2778 585
R2654 gnd.n2778 gnd.n2777 585
R2655 gnd.n3273 gnd.n3272 585
R2656 gnd.n3272 gnd.n2759 585
R2657 gnd.n3270 gnd.n2757 585
R2658 gnd.n3291 gnd.n2757 585
R2659 gnd.n2788 gnd.n2787 585
R2660 gnd.n2787 gnd.n2786 585
R2661 gnd.n3264 gnd.n2747 585
R2662 gnd.n3297 gnd.n2747 585
R2663 gnd.n3263 gnd.n3262 585
R2664 gnd.n3262 gnd.n3261 585
R2665 gnd.n3259 gnd.n2790 585
R2666 gnd.n3259 gnd.n2737 585
R2667 gnd.n3258 gnd.n3257 585
R2668 gnd.n3258 gnd.n2736 585
R2669 gnd.n2793 gnd.n2792 585
R2670 gnd.n3249 gnd.n2792 585
R2671 gnd.n3217 gnd.n3216 585
R2672 gnd.n3216 gnd.n2797 585
R2673 gnd.n3218 gnd.n2806 585
R2674 gnd.n3235 gnd.n2806 585
R2675 gnd.n3215 gnd.n3214 585
R2676 gnd.n3214 gnd.n2812 585
R2677 gnd.n3213 gnd.n2820 585
R2678 gnd.n3213 gnd.n3212 585
R2679 gnd.n3198 gnd.n2821 585
R2680 gnd.n2831 gnd.n2821 585
R2681 gnd.n3197 gnd.n2829 585
R2682 gnd.n3204 gnd.n2829 585
R2683 gnd.n3196 gnd.n3195 585
R2684 gnd.n3195 gnd.n3194 585
R2685 gnd.n2840 gnd.n2837 585
R2686 gnd.n2850 gnd.n2840 585
R2687 gnd.n3186 gnd.n3185 585
R2688 gnd.n3185 gnd.n3184 585
R2689 gnd.n2846 gnd.n2845 585
R2690 gnd.n2859 gnd.n2846 585
R2691 gnd.n3166 gnd.n2857 585
R2692 gnd.n3174 gnd.n2857 585
R2693 gnd.n3165 gnd.n3164 585
R2694 gnd.n3164 gnd.n3163 585
R2695 gnd.n2866 gnd.n2864 585
R2696 gnd.n2875 gnd.n2866 585
R2697 gnd.n3155 gnd.n3154 585
R2698 gnd.n3154 gnd.n3153 585
R2699 gnd.n5413 gnd.n5412 585
R2700 gnd.n5414 gnd.n5413 585
R2701 gnd.n5327 gnd.n1829 585
R2702 gnd.n1836 gnd.n1829 585
R2703 gnd.n5326 gnd.n5325 585
R2704 gnd.n5325 gnd.n5324 585
R2705 gnd.n1832 gnd.n1831 585
R2706 gnd.n5095 gnd.n1832 585
R2707 gnd.n5084 gnd.n1879 585
R2708 gnd.n1879 gnd.n1873 585
R2709 gnd.n5086 gnd.n5085 585
R2710 gnd.n5087 gnd.n5086 585
R2711 gnd.n5083 gnd.n1878 585
R2712 gnd.n5077 gnd.n1878 585
R2713 gnd.n5082 gnd.n5081 585
R2714 gnd.n5081 gnd.n5080 585
R2715 gnd.n1881 gnd.n1880 585
R2716 gnd.n5064 gnd.n1881 585
R2717 gnd.n5039 gnd.n5038 585
R2718 gnd.n5038 gnd.n1892 585
R2719 gnd.n5040 gnd.n1901 585
R2720 gnd.n5053 gnd.n1901 585
R2721 gnd.n5041 gnd.n1911 585
R2722 gnd.n1911 gnd.n1900 585
R2723 gnd.n5043 gnd.n5042 585
R2724 gnd.n5044 gnd.n5043 585
R2725 gnd.n5037 gnd.n1910 585
R2726 gnd.n5032 gnd.n1910 585
R2727 gnd.n5036 gnd.n5035 585
R2728 gnd.n5035 gnd.n5034 585
R2729 gnd.n1913 gnd.n1912 585
R2730 gnd.n5019 gnd.n1913 585
R2731 gnd.n5008 gnd.n1928 585
R2732 gnd.n1928 gnd.n1922 585
R2733 gnd.n5010 gnd.n5009 585
R2734 gnd.n5011 gnd.n5010 585
R2735 gnd.n5007 gnd.n1927 585
R2736 gnd.n1934 gnd.n1927 585
R2737 gnd.n5006 gnd.n5005 585
R2738 gnd.n5005 gnd.n5004 585
R2739 gnd.n1930 gnd.n1929 585
R2740 gnd.n4885 gnd.n1930 585
R2741 gnd.n4992 gnd.n4991 585
R2742 gnd.n4993 gnd.n4992 585
R2743 gnd.n4990 gnd.n1946 585
R2744 gnd.n1946 gnd.n1942 585
R2745 gnd.n4989 gnd.n4988 585
R2746 gnd.n4988 gnd.n4987 585
R2747 gnd.n1948 gnd.n1947 585
R2748 gnd.n4895 gnd.n1948 585
R2749 gnd.n4961 gnd.n4960 585
R2750 gnd.n4962 gnd.n4961 585
R2751 gnd.n4959 gnd.n1959 585
R2752 gnd.n1959 gnd.n1956 585
R2753 gnd.n4958 gnd.n4957 585
R2754 gnd.n4957 gnd.n4956 585
R2755 gnd.n1961 gnd.n1960 585
R2756 gnd.n4902 gnd.n1961 585
R2757 gnd.n4942 gnd.n4941 585
R2758 gnd.n4943 gnd.n4942 585
R2759 gnd.n4940 gnd.n1972 585
R2760 gnd.n4935 gnd.n1972 585
R2761 gnd.n4939 gnd.n4938 585
R2762 gnd.n4938 gnd.n4937 585
R2763 gnd.n1974 gnd.n1973 585
R2764 gnd.n1986 gnd.n1974 585
R2765 gnd.n4871 gnd.n4870 585
R2766 gnd.n4871 gnd.n1985 585
R2767 gnd.n4875 gnd.n4874 585
R2768 gnd.n4874 gnd.n4873 585
R2769 gnd.n4876 gnd.n1992 585
R2770 gnd.n4915 gnd.n1992 585
R2771 gnd.n4877 gnd.n2001 585
R2772 gnd.n4801 gnd.n2001 585
R2773 gnd.n4879 gnd.n4878 585
R2774 gnd.n4880 gnd.n4879 585
R2775 gnd.n4869 gnd.n2000 585
R2776 gnd.n4864 gnd.n2000 585
R2777 gnd.n4868 gnd.n4867 585
R2778 gnd.n4867 gnd.n4866 585
R2779 gnd.n2003 gnd.n2002 585
R2780 gnd.n4853 gnd.n2003 585
R2781 gnd.n4843 gnd.n2021 585
R2782 gnd.n2021 gnd.n2012 585
R2783 gnd.n4845 gnd.n4844 585
R2784 gnd.n4846 gnd.n4845 585
R2785 gnd.n4842 gnd.n2020 585
R2786 gnd.n2025 gnd.n2020 585
R2787 gnd.n4841 gnd.n4840 585
R2788 gnd.n4840 gnd.n4839 585
R2789 gnd.n2023 gnd.n2022 585
R2790 gnd.n4793 gnd.n2023 585
R2791 gnd.n4827 gnd.n4826 585
R2792 gnd.n4828 gnd.n4827 585
R2793 gnd.n4825 gnd.n2036 585
R2794 gnd.n2036 gnd.n2032 585
R2795 gnd.n4824 gnd.n4823 585
R2796 gnd.n4823 gnd.n4822 585
R2797 gnd.n2038 gnd.n2037 585
R2798 gnd.n4783 gnd.n2038 585
R2799 gnd.n4768 gnd.n4767 585
R2800 gnd.n4767 gnd.n2048 585
R2801 gnd.n4769 gnd.n2058 585
R2802 gnd.n4752 gnd.n2058 585
R2803 gnd.n4771 gnd.n4770 585
R2804 gnd.n4772 gnd.n4771 585
R2805 gnd.n4766 gnd.n2057 585
R2806 gnd.n2057 gnd.n2054 585
R2807 gnd.n4765 gnd.n4764 585
R2808 gnd.n4764 gnd.n4763 585
R2809 gnd.n2060 gnd.n2059 585
R2810 gnd.n4743 gnd.n2060 585
R2811 gnd.n4728 gnd.n4727 585
R2812 gnd.n4727 gnd.n2071 585
R2813 gnd.n4729 gnd.n2081 585
R2814 gnd.n4716 gnd.n2081 585
R2815 gnd.n4731 gnd.n4730 585
R2816 gnd.n4732 gnd.n4731 585
R2817 gnd.n4726 gnd.n2080 585
R2818 gnd.n2080 gnd.n2077 585
R2819 gnd.n4725 gnd.n4724 585
R2820 gnd.n4724 gnd.n4723 585
R2821 gnd.n2083 gnd.n2082 585
R2822 gnd.n2096 gnd.n2083 585
R2823 gnd.n4701 gnd.n4700 585
R2824 gnd.n4702 gnd.n4701 585
R2825 gnd.n4699 gnd.n2098 585
R2826 gnd.n4694 gnd.n2098 585
R2827 gnd.n4698 gnd.n4697 585
R2828 gnd.n4697 gnd.n4696 585
R2829 gnd.n2100 gnd.n2099 585
R2830 gnd.n4680 gnd.n2100 585
R2831 gnd.n4668 gnd.n2118 585
R2832 gnd.n2118 gnd.n2110 585
R2833 gnd.n4670 gnd.n4669 585
R2834 gnd.n4671 gnd.n4670 585
R2835 gnd.n4667 gnd.n2117 585
R2836 gnd.n4612 gnd.n2117 585
R2837 gnd.n4666 gnd.n4665 585
R2838 gnd.n4665 gnd.n4664 585
R2839 gnd.n2120 gnd.n2119 585
R2840 gnd.n4638 gnd.n2120 585
R2841 gnd.n4651 gnd.n4650 585
R2842 gnd.n4652 gnd.n4651 585
R2843 gnd.n4649 gnd.n2131 585
R2844 gnd.n4644 gnd.n2131 585
R2845 gnd.n4648 gnd.n4647 585
R2846 gnd.n4647 gnd.n4646 585
R2847 gnd.n2133 gnd.n2132 585
R2848 gnd.n4633 gnd.n2133 585
R2849 gnd.n4585 gnd.n4582 585
R2850 gnd.n4585 gnd.n4584 585
R2851 gnd.n4586 gnd.n4581 585
R2852 gnd.n4586 gnd.n2147 585
R2853 gnd.n4588 gnd.n4587 585
R2854 gnd.n4587 gnd.n2146 585
R2855 gnd.n4589 gnd.n2158 585
R2856 gnd.n4569 gnd.n2158 585
R2857 gnd.n4591 gnd.n4590 585
R2858 gnd.n4592 gnd.n4591 585
R2859 gnd.n4580 gnd.n2157 585
R2860 gnd.n4575 gnd.n2157 585
R2861 gnd.n4579 gnd.n4578 585
R2862 gnd.n4578 gnd.n4577 585
R2863 gnd.n2160 gnd.n2159 585
R2864 gnd.n4560 gnd.n2160 585
R2865 gnd.n2183 gnd.n2182 585
R2866 gnd.n4535 gnd.n2183 585
R2867 gnd.n4539 gnd.n4538 585
R2868 gnd.n4538 gnd.n4537 585
R2869 gnd.n4540 gnd.n2172 585
R2870 gnd.n4551 gnd.n2172 585
R2871 gnd.n4541 gnd.n2180 585
R2872 gnd.n2184 gnd.n2180 585
R2873 gnd.n4543 gnd.n4542 585
R2874 gnd.n4544 gnd.n4543 585
R2875 gnd.n2181 gnd.n2179 585
R2876 gnd.n4517 gnd.n2179 585
R2877 gnd.n4510 gnd.n4509 585
R2878 gnd.n4511 gnd.n4510 585
R2879 gnd.n4508 gnd.n2194 585
R2880 gnd.n2194 gnd.n1492 585
R2881 gnd.n4507 gnd.n4506 585
R2882 gnd.n4506 gnd.n1490 585
R2883 gnd.n4505 gnd.n2195 585
R2884 gnd.n4505 gnd.n4504 585
R2885 gnd.n1478 gnd.n1477 585
R2886 gnd.n2275 gnd.n1478 585
R2887 gnd.n5994 gnd.n5993 585
R2888 gnd.n5993 gnd.n5992 585
R2889 gnd.n5995 gnd.n1456 585
R2890 gnd.n2281 gnd.n1456 585
R2891 gnd.n6060 gnd.n6059 585
R2892 gnd.n6058 gnd.n1455 585
R2893 gnd.n6057 gnd.n1454 585
R2894 gnd.n6062 gnd.n1454 585
R2895 gnd.n6056 gnd.n6055 585
R2896 gnd.n6054 gnd.n6053 585
R2897 gnd.n6052 gnd.n6051 585
R2898 gnd.n6050 gnd.n6049 585
R2899 gnd.n6048 gnd.n6047 585
R2900 gnd.n6046 gnd.n6045 585
R2901 gnd.n6044 gnd.n6043 585
R2902 gnd.n6042 gnd.n6041 585
R2903 gnd.n6040 gnd.n6039 585
R2904 gnd.n6038 gnd.n6037 585
R2905 gnd.n6036 gnd.n6035 585
R2906 gnd.n6034 gnd.n6033 585
R2907 gnd.n6032 gnd.n6031 585
R2908 gnd.n6030 gnd.n6029 585
R2909 gnd.n6028 gnd.n6027 585
R2910 gnd.n6026 gnd.n6025 585
R2911 gnd.n6024 gnd.n6023 585
R2912 gnd.n6022 gnd.n6021 585
R2913 gnd.n6020 gnd.n6019 585
R2914 gnd.n6018 gnd.n6017 585
R2915 gnd.n6016 gnd.n6015 585
R2916 gnd.n6014 gnd.n6013 585
R2917 gnd.n6012 gnd.n6011 585
R2918 gnd.n6010 gnd.n6009 585
R2919 gnd.n6008 gnd.n6007 585
R2920 gnd.n6006 gnd.n6005 585
R2921 gnd.n6004 gnd.n6003 585
R2922 gnd.n6002 gnd.n6001 585
R2923 gnd.n6000 gnd.n1418 585
R2924 gnd.n6065 gnd.n6064 585
R2925 gnd.n1420 gnd.n1417 585
R2926 gnd.n2208 gnd.n2207 585
R2927 gnd.n2210 gnd.n2209 585
R2928 gnd.n2213 gnd.n2212 585
R2929 gnd.n2215 gnd.n2214 585
R2930 gnd.n2217 gnd.n2216 585
R2931 gnd.n2219 gnd.n2218 585
R2932 gnd.n2221 gnd.n2220 585
R2933 gnd.n2223 gnd.n2222 585
R2934 gnd.n2225 gnd.n2224 585
R2935 gnd.n2227 gnd.n2226 585
R2936 gnd.n2229 gnd.n2228 585
R2937 gnd.n2231 gnd.n2230 585
R2938 gnd.n2233 gnd.n2232 585
R2939 gnd.n2235 gnd.n2234 585
R2940 gnd.n2237 gnd.n2236 585
R2941 gnd.n2239 gnd.n2238 585
R2942 gnd.n2241 gnd.n2240 585
R2943 gnd.n2243 gnd.n2242 585
R2944 gnd.n2245 gnd.n2244 585
R2945 gnd.n2247 gnd.n2246 585
R2946 gnd.n2249 gnd.n2248 585
R2947 gnd.n2251 gnd.n2250 585
R2948 gnd.n2253 gnd.n2252 585
R2949 gnd.n2255 gnd.n2254 585
R2950 gnd.n2257 gnd.n2256 585
R2951 gnd.n2259 gnd.n2258 585
R2952 gnd.n2261 gnd.n2260 585
R2953 gnd.n2263 gnd.n2262 585
R2954 gnd.n2265 gnd.n2264 585
R2955 gnd.n2267 gnd.n2266 585
R2956 gnd.n2268 gnd.n2204 585
R2957 gnd.n5417 gnd.n5416 585
R2958 gnd.n5419 gnd.n5418 585
R2959 gnd.n5421 gnd.n5420 585
R2960 gnd.n5423 gnd.n5422 585
R2961 gnd.n5425 gnd.n5424 585
R2962 gnd.n5427 gnd.n5426 585
R2963 gnd.n5429 gnd.n5428 585
R2964 gnd.n5431 gnd.n5430 585
R2965 gnd.n5433 gnd.n5432 585
R2966 gnd.n5435 gnd.n5434 585
R2967 gnd.n5437 gnd.n5436 585
R2968 gnd.n5439 gnd.n5438 585
R2969 gnd.n5441 gnd.n5440 585
R2970 gnd.n5443 gnd.n5442 585
R2971 gnd.n5445 gnd.n5444 585
R2972 gnd.n5447 gnd.n5446 585
R2973 gnd.n5449 gnd.n5448 585
R2974 gnd.n5451 gnd.n5450 585
R2975 gnd.n5453 gnd.n5452 585
R2976 gnd.n5455 gnd.n5454 585
R2977 gnd.n5457 gnd.n5456 585
R2978 gnd.n5459 gnd.n5458 585
R2979 gnd.n5461 gnd.n5460 585
R2980 gnd.n5463 gnd.n5462 585
R2981 gnd.n5465 gnd.n5464 585
R2982 gnd.n5467 gnd.n5466 585
R2983 gnd.n5469 gnd.n5468 585
R2984 gnd.n5471 gnd.n5470 585
R2985 gnd.n5473 gnd.n5472 585
R2986 gnd.n5475 gnd.n1823 585
R2987 gnd.n5477 gnd.n5476 585
R2988 gnd.n5479 gnd.n1787 585
R2989 gnd.n5481 gnd.n5480 585
R2990 gnd.n5484 gnd.n5483 585
R2991 gnd.n1790 gnd.n1788 585
R2992 gnd.n5350 gnd.n5349 585
R2993 gnd.n5352 gnd.n5351 585
R2994 gnd.n5355 gnd.n5354 585
R2995 gnd.n5357 gnd.n5356 585
R2996 gnd.n5359 gnd.n5358 585
R2997 gnd.n5361 gnd.n5360 585
R2998 gnd.n5363 gnd.n5362 585
R2999 gnd.n5365 gnd.n5364 585
R3000 gnd.n5367 gnd.n5366 585
R3001 gnd.n5369 gnd.n5368 585
R3002 gnd.n5371 gnd.n5370 585
R3003 gnd.n5373 gnd.n5372 585
R3004 gnd.n5375 gnd.n5374 585
R3005 gnd.n5377 gnd.n5376 585
R3006 gnd.n5379 gnd.n5378 585
R3007 gnd.n5381 gnd.n5380 585
R3008 gnd.n5383 gnd.n5382 585
R3009 gnd.n5385 gnd.n5384 585
R3010 gnd.n5387 gnd.n5386 585
R3011 gnd.n5389 gnd.n5388 585
R3012 gnd.n5391 gnd.n5390 585
R3013 gnd.n5393 gnd.n5392 585
R3014 gnd.n5395 gnd.n5394 585
R3015 gnd.n5397 gnd.n5396 585
R3016 gnd.n5399 gnd.n5398 585
R3017 gnd.n5401 gnd.n5400 585
R3018 gnd.n5403 gnd.n5402 585
R3019 gnd.n5405 gnd.n5404 585
R3020 gnd.n5407 gnd.n5406 585
R3021 gnd.n5409 gnd.n5408 585
R3022 gnd.n5410 gnd.n1830 585
R3023 gnd.n5415 gnd.n1826 585
R3024 gnd.n5415 gnd.n5414 585
R3025 gnd.n5091 gnd.n1827 585
R3026 gnd.n1836 gnd.n1827 585
R3027 gnd.n5092 gnd.n1834 585
R3028 gnd.n5324 gnd.n1834 585
R3029 gnd.n5094 gnd.n5093 585
R3030 gnd.n5095 gnd.n5094 585
R3031 gnd.n5090 gnd.n1874 585
R3032 gnd.n1874 gnd.n1873 585
R3033 gnd.n5089 gnd.n5088 585
R3034 gnd.n5088 gnd.n5087 585
R3035 gnd.n1876 gnd.n1875 585
R3036 gnd.n5077 gnd.n1876 585
R3037 gnd.n5048 gnd.n1883 585
R3038 gnd.n5080 gnd.n1883 585
R3039 gnd.n5049 gnd.n1893 585
R3040 gnd.n5064 gnd.n1893 585
R3041 gnd.n5050 gnd.n1904 585
R3042 gnd.n1904 gnd.n1892 585
R3043 gnd.n5052 gnd.n5051 585
R3044 gnd.n5053 gnd.n5052 585
R3045 gnd.n5047 gnd.n1903 585
R3046 gnd.n1903 gnd.n1900 585
R3047 gnd.n5046 gnd.n5045 585
R3048 gnd.n5045 gnd.n5044 585
R3049 gnd.n1906 gnd.n1905 585
R3050 gnd.n5032 gnd.n1906 585
R3051 gnd.n5015 gnd.n1914 585
R3052 gnd.n5034 gnd.n1914 585
R3053 gnd.n5017 gnd.n5016 585
R3054 gnd.n5019 gnd.n5017 585
R3055 gnd.n5014 gnd.n1924 585
R3056 gnd.n1924 gnd.n1922 585
R3057 gnd.n5013 gnd.n5012 585
R3058 gnd.n5012 gnd.n5011 585
R3059 gnd.n1926 gnd.n1925 585
R3060 gnd.n1934 gnd.n1926 585
R3061 gnd.n4884 gnd.n1932 585
R3062 gnd.n5004 gnd.n1932 585
R3063 gnd.n4887 gnd.n4886 585
R3064 gnd.n4886 gnd.n4885 585
R3065 gnd.n4888 gnd.n1944 585
R3066 gnd.n4993 gnd.n1944 585
R3067 gnd.n4890 gnd.n4889 585
R3068 gnd.n4889 gnd.n1942 585
R3069 gnd.n4891 gnd.n1949 585
R3070 gnd.n4987 gnd.n1949 585
R3071 gnd.n4897 gnd.n4896 585
R3072 gnd.n4896 gnd.n4895 585
R3073 gnd.n4898 gnd.n1957 585
R3074 gnd.n4962 gnd.n1957 585
R3075 gnd.n4900 gnd.n4899 585
R3076 gnd.n4899 gnd.n1956 585
R3077 gnd.n4901 gnd.n1963 585
R3078 gnd.n4956 gnd.n1963 585
R3079 gnd.n4904 gnd.n4903 585
R3080 gnd.n4903 gnd.n4902 585
R3081 gnd.n4905 gnd.n1970 585
R3082 gnd.n4943 gnd.n1970 585
R3083 gnd.n4906 gnd.n1977 585
R3084 gnd.n4935 gnd.n1977 585
R3085 gnd.n4907 gnd.n1976 585
R3086 gnd.n4937 gnd.n1976 585
R3087 gnd.n4909 gnd.n4908 585
R3088 gnd.n4909 gnd.n1986 585
R3089 gnd.n4911 gnd.n4910 585
R3090 gnd.n4910 gnd.n1985 585
R3091 gnd.n4912 gnd.n1995 585
R3092 gnd.n4873 gnd.n1995 585
R3093 gnd.n4914 gnd.n4913 585
R3094 gnd.n4915 gnd.n4914 585
R3095 gnd.n4883 gnd.n1994 585
R3096 gnd.n4801 gnd.n1994 585
R3097 gnd.n4882 gnd.n4881 585
R3098 gnd.n4881 gnd.n4880 585
R3099 gnd.n1997 gnd.n1996 585
R3100 gnd.n4864 gnd.n1997 585
R3101 gnd.n4850 gnd.n2005 585
R3102 gnd.n4866 gnd.n2005 585
R3103 gnd.n4852 gnd.n4851 585
R3104 gnd.n4853 gnd.n4852 585
R3105 gnd.n4849 gnd.n2014 585
R3106 gnd.n2014 gnd.n2012 585
R3107 gnd.n4848 gnd.n4847 585
R3108 gnd.n4847 gnd.n4846 585
R3109 gnd.n2016 gnd.n2015 585
R3110 gnd.n2025 gnd.n2016 585
R3111 gnd.n4790 gnd.n2024 585
R3112 gnd.n4839 gnd.n2024 585
R3113 gnd.n4792 gnd.n4791 585
R3114 gnd.n4793 gnd.n4792 585
R3115 gnd.n4789 gnd.n2034 585
R3116 gnd.n4828 gnd.n2034 585
R3117 gnd.n4788 gnd.n4787 585
R3118 gnd.n4787 gnd.n2032 585
R3119 gnd.n4786 gnd.n2040 585
R3120 gnd.n4822 gnd.n2040 585
R3121 gnd.n4785 gnd.n4784 585
R3122 gnd.n4784 gnd.n4783 585
R3123 gnd.n2047 gnd.n2046 585
R3124 gnd.n2048 gnd.n2047 585
R3125 gnd.n4751 gnd.n4750 585
R3126 gnd.n4752 gnd.n4751 585
R3127 gnd.n4749 gnd.n2055 585
R3128 gnd.n4772 gnd.n2055 585
R3129 gnd.n4748 gnd.n4747 585
R3130 gnd.n4747 gnd.n2054 585
R3131 gnd.n4746 gnd.n2062 585
R3132 gnd.n4763 gnd.n2062 585
R3133 gnd.n4745 gnd.n4744 585
R3134 gnd.n4744 gnd.n4743 585
R3135 gnd.n2070 gnd.n2069 585
R3136 gnd.n2071 gnd.n2070 585
R3137 gnd.n4718 gnd.n4717 585
R3138 gnd.n4717 gnd.n4716 585
R3139 gnd.n4719 gnd.n2078 585
R3140 gnd.n4732 gnd.n2078 585
R3141 gnd.n4720 gnd.n2086 585
R3142 gnd.n2086 gnd.n2077 585
R3143 gnd.n4722 gnd.n4721 585
R3144 gnd.n4723 gnd.n4722 585
R3145 gnd.n2087 gnd.n2085 585
R3146 gnd.n2096 gnd.n2085 585
R3147 gnd.n4675 gnd.n2095 585
R3148 gnd.n4702 gnd.n2095 585
R3149 gnd.n4676 gnd.n2103 585
R3150 gnd.n4694 gnd.n2103 585
R3151 gnd.n4677 gnd.n2102 585
R3152 gnd.n4696 gnd.n2102 585
R3153 gnd.n4679 gnd.n4678 585
R3154 gnd.n4680 gnd.n4679 585
R3155 gnd.n4674 gnd.n2112 585
R3156 gnd.n2112 gnd.n2110 585
R3157 gnd.n4673 gnd.n4672 585
R3158 gnd.n4672 gnd.n4671 585
R3159 gnd.n2114 gnd.n2113 585
R3160 gnd.n4612 gnd.n2114 585
R3161 gnd.n4637 gnd.n2122 585
R3162 gnd.n4664 gnd.n2122 585
R3163 gnd.n4640 gnd.n4639 585
R3164 gnd.n4639 gnd.n4638 585
R3165 gnd.n4641 gnd.n2129 585
R3166 gnd.n4652 gnd.n2129 585
R3167 gnd.n4643 gnd.n4642 585
R3168 gnd.n4644 gnd.n4643 585
R3169 gnd.n4636 gnd.n2135 585
R3170 gnd.n4646 gnd.n2135 585
R3171 gnd.n4635 gnd.n4634 585
R3172 gnd.n4634 gnd.n4633 585
R3173 gnd.n2138 gnd.n2137 585
R3174 gnd.n4584 gnd.n2138 585
R3175 gnd.n4566 gnd.n4565 585
R3176 gnd.n4566 gnd.n2147 585
R3177 gnd.n4567 gnd.n4564 585
R3178 gnd.n4567 gnd.n2146 585
R3179 gnd.n4571 gnd.n4570 585
R3180 gnd.n4570 gnd.n4569 585
R3181 gnd.n4572 gnd.n2155 585
R3182 gnd.n4592 gnd.n2155 585
R3183 gnd.n4574 gnd.n4573 585
R3184 gnd.n4575 gnd.n4574 585
R3185 gnd.n4563 gnd.n2162 585
R3186 gnd.n4577 gnd.n2162 585
R3187 gnd.n4562 gnd.n4561 585
R3188 gnd.n4561 gnd.n4560 585
R3189 gnd.n2164 gnd.n2163 585
R3190 gnd.n4535 gnd.n2164 585
R3191 gnd.n4548 gnd.n2174 585
R3192 gnd.n4537 gnd.n2174 585
R3193 gnd.n4550 gnd.n4549 585
R3194 gnd.n4551 gnd.n4550 585
R3195 gnd.n4547 gnd.n2173 585
R3196 gnd.n2184 gnd.n2173 585
R3197 gnd.n4546 gnd.n4545 585
R3198 gnd.n4545 gnd.n4544 585
R3199 gnd.n2176 gnd.n2175 585
R3200 gnd.n4517 gnd.n2176 585
R3201 gnd.n2269 gnd.n2193 585
R3202 gnd.n4511 gnd.n2193 585
R3203 gnd.n2271 gnd.n2270 585
R3204 gnd.n2271 gnd.n1492 585
R3205 gnd.n2273 gnd.n2272 585
R3206 gnd.n2272 gnd.n1490 585
R3207 gnd.n2274 gnd.n2197 585
R3208 gnd.n4504 gnd.n2197 585
R3209 gnd.n2277 gnd.n2276 585
R3210 gnd.n2276 gnd.n2275 585
R3211 gnd.n2278 gnd.n1480 585
R3212 gnd.n5992 gnd.n1480 585
R3213 gnd.n2280 gnd.n2279 585
R3214 gnd.n2281 gnd.n2280 585
R3215 gnd.n6201 gnd.n6200 585
R3216 gnd.n6200 gnd.n6199 585
R3217 gnd.n6202 gnd.n1132 585
R3218 gnd.n6192 gnd.n1132 585
R3219 gnd.n6204 gnd.n6203 585
R3220 gnd.n6205 gnd.n6204 585
R3221 gnd.n1117 gnd.n1116 585
R3222 gnd.n4398 gnd.n1117 585
R3223 gnd.n6213 gnd.n6212 585
R3224 gnd.n6212 gnd.n6211 585
R3225 gnd.n6214 gnd.n1111 585
R3226 gnd.n4392 gnd.n1111 585
R3227 gnd.n6216 gnd.n6215 585
R3228 gnd.n6217 gnd.n6216 585
R3229 gnd.n1097 gnd.n1096 585
R3230 gnd.n4409 gnd.n1097 585
R3231 gnd.n6225 gnd.n6224 585
R3232 gnd.n6224 gnd.n6223 585
R3233 gnd.n6226 gnd.n1091 585
R3234 gnd.n4385 gnd.n1091 585
R3235 gnd.n6228 gnd.n6227 585
R3236 gnd.n6229 gnd.n6228 585
R3237 gnd.n1077 gnd.n1076 585
R3238 gnd.n4377 gnd.n1077 585
R3239 gnd.n6237 gnd.n6236 585
R3240 gnd.n6236 gnd.n6235 585
R3241 gnd.n6238 gnd.n1071 585
R3242 gnd.n4371 gnd.n1071 585
R3243 gnd.n6240 gnd.n6239 585
R3244 gnd.n6241 gnd.n6240 585
R3245 gnd.n1057 gnd.n1056 585
R3246 gnd.n4363 gnd.n1057 585
R3247 gnd.n6249 gnd.n6248 585
R3248 gnd.n6248 gnd.n6247 585
R3249 gnd.n6250 gnd.n1054 585
R3250 gnd.n4307 gnd.n1054 585
R3251 gnd.n6253 gnd.n6252 585
R3252 gnd.n6254 gnd.n6253 585
R3253 gnd.n1055 gnd.n1040 585
R3254 gnd.n4315 gnd.n1040 585
R3255 gnd.n6262 gnd.n6261 585
R3256 gnd.n6261 gnd.n6260 585
R3257 gnd.n6263 gnd.n1037 585
R3258 gnd.n4296 gnd.n1037 585
R3259 gnd.n6266 gnd.n6265 585
R3260 gnd.n6267 gnd.n6266 585
R3261 gnd.n1038 gnd.n1021 585
R3262 gnd.n4326 gnd.n1021 585
R3263 gnd.n6275 gnd.n6274 585
R3264 gnd.n6274 gnd.n6273 585
R3265 gnd.n6276 gnd.n1019 585
R3266 gnd.n4332 gnd.n1019 585
R3267 gnd.n6278 gnd.n1015 585
R3268 gnd.n2370 gnd.n1015 585
R3269 gnd.n6280 gnd.n6279 585
R3270 gnd.n6281 gnd.n6280 585
R3271 gnd.n1001 gnd.n1000 585
R3272 gnd.n4279 gnd.n1001 585
R3273 gnd.n6289 gnd.n6288 585
R3274 gnd.n6288 gnd.n6287 585
R3275 gnd.n6290 gnd.n995 585
R3276 gnd.n4267 gnd.n995 585
R3277 gnd.n6292 gnd.n6291 585
R3278 gnd.n6293 gnd.n6292 585
R3279 gnd.n979 gnd.n978 585
R3280 gnd.n4260 gnd.n979 585
R3281 gnd.n6301 gnd.n6300 585
R3282 gnd.n6300 gnd.n6299 585
R3283 gnd.n6302 gnd.n973 585
R3284 gnd.n4252 gnd.n973 585
R3285 gnd.n6304 gnd.n6303 585
R3286 gnd.n6305 gnd.n6304 585
R3287 gnd.n974 gnd.n972 585
R3288 gnd.n972 gnd.n967 585
R3289 gnd.n4242 gnd.n4241 585
R3290 gnd.n4243 gnd.n4242 585
R3291 gnd.n2427 gnd.n2426 585
R3292 gnd.n2434 gnd.n2426 585
R3293 gnd.n4236 gnd.n4235 585
R3294 gnd.n4235 gnd.n4234 585
R3295 gnd.n2430 gnd.n2429 585
R3296 gnd.n2431 gnd.n2430 585
R3297 gnd.n4219 gnd.n4218 585
R3298 gnd.n4220 gnd.n4219 585
R3299 gnd.n2446 gnd.n2445 585
R3300 gnd.n2445 gnd.n2442 585
R3301 gnd.n4214 gnd.n4213 585
R3302 gnd.n2449 gnd.n2448 585
R3303 gnd.n4210 gnd.n4209 585
R3304 gnd.n4211 gnd.n4210 585
R3305 gnd.n4208 gnd.n3950 585
R3306 gnd.n4207 gnd.n4206 585
R3307 gnd.n4205 gnd.n4204 585
R3308 gnd.n4203 gnd.n4202 585
R3309 gnd.n4201 gnd.n4200 585
R3310 gnd.n4199 gnd.n4198 585
R3311 gnd.n4197 gnd.n4196 585
R3312 gnd.n4195 gnd.n4194 585
R3313 gnd.n4193 gnd.n4192 585
R3314 gnd.n4191 gnd.n4190 585
R3315 gnd.n4189 gnd.n4188 585
R3316 gnd.n4187 gnd.n4186 585
R3317 gnd.n4185 gnd.n4184 585
R3318 gnd.n4183 gnd.n4182 585
R3319 gnd.n4181 gnd.n4180 585
R3320 gnd.n4178 gnd.n4177 585
R3321 gnd.n4176 gnd.n4175 585
R3322 gnd.n4174 gnd.n4173 585
R3323 gnd.n4172 gnd.n4171 585
R3324 gnd.n4170 gnd.n4169 585
R3325 gnd.n4168 gnd.n4167 585
R3326 gnd.n4166 gnd.n4165 585
R3327 gnd.n4164 gnd.n4163 585
R3328 gnd.n4162 gnd.n4161 585
R3329 gnd.n4160 gnd.n4159 585
R3330 gnd.n4158 gnd.n4157 585
R3331 gnd.n4156 gnd.n4155 585
R3332 gnd.n4154 gnd.n4153 585
R3333 gnd.n4152 gnd.n4151 585
R3334 gnd.n4150 gnd.n4149 585
R3335 gnd.n4148 gnd.n4147 585
R3336 gnd.n4146 gnd.n4145 585
R3337 gnd.n4144 gnd.n4143 585
R3338 gnd.n4142 gnd.n4141 585
R3339 gnd.n4140 gnd.n4139 585
R3340 gnd.n4138 gnd.n4137 585
R3341 gnd.n4136 gnd.n4135 585
R3342 gnd.n4134 gnd.n4133 585
R3343 gnd.n4132 gnd.n4131 585
R3344 gnd.n4130 gnd.n4129 585
R3345 gnd.n4128 gnd.n4127 585
R3346 gnd.n4126 gnd.n4125 585
R3347 gnd.n4124 gnd.n4123 585
R3348 gnd.n4122 gnd.n4121 585
R3349 gnd.n4120 gnd.n4119 585
R3350 gnd.n4118 gnd.n4117 585
R3351 gnd.n4116 gnd.n4115 585
R3352 gnd.n4114 gnd.n4113 585
R3353 gnd.n4112 gnd.n4111 585
R3354 gnd.n4110 gnd.n4109 585
R3355 gnd.n4108 gnd.n4107 585
R3356 gnd.n4106 gnd.n4105 585
R3357 gnd.n4104 gnd.n4103 585
R3358 gnd.n4102 gnd.n4101 585
R3359 gnd.n4100 gnd.n4099 585
R3360 gnd.n4011 gnd.n4010 585
R3361 gnd.n1348 gnd.n1347 585
R3362 gnd.n1354 gnd.n1353 585
R3363 gnd.n1356 gnd.n1355 585
R3364 gnd.n1358 gnd.n1357 585
R3365 gnd.n1360 gnd.n1359 585
R3366 gnd.n1362 gnd.n1361 585
R3367 gnd.n1364 gnd.n1363 585
R3368 gnd.n1366 gnd.n1365 585
R3369 gnd.n1368 gnd.n1367 585
R3370 gnd.n1370 gnd.n1369 585
R3371 gnd.n1372 gnd.n1371 585
R3372 gnd.n1374 gnd.n1373 585
R3373 gnd.n1376 gnd.n1375 585
R3374 gnd.n1378 gnd.n1377 585
R3375 gnd.n1380 gnd.n1379 585
R3376 gnd.n1382 gnd.n1381 585
R3377 gnd.n1384 gnd.n1383 585
R3378 gnd.n1386 gnd.n1385 585
R3379 gnd.n1388 gnd.n1387 585
R3380 gnd.n1391 gnd.n1390 585
R3381 gnd.n1389 gnd.n1327 585
R3382 gnd.n1396 gnd.n1395 585
R3383 gnd.n1398 gnd.n1397 585
R3384 gnd.n1400 gnd.n1399 585
R3385 gnd.n1402 gnd.n1401 585
R3386 gnd.n1404 gnd.n1403 585
R3387 gnd.n1406 gnd.n1405 585
R3388 gnd.n1408 gnd.n1407 585
R3389 gnd.n1410 gnd.n1409 585
R3390 gnd.n1413 gnd.n1412 585
R3391 gnd.n1411 gnd.n1318 585
R3392 gnd.n6068 gnd.n6067 585
R3393 gnd.n6070 gnd.n6069 585
R3394 gnd.n6072 gnd.n6071 585
R3395 gnd.n6074 gnd.n6073 585
R3396 gnd.n6076 gnd.n6075 585
R3397 gnd.n6078 gnd.n6077 585
R3398 gnd.n6080 gnd.n6079 585
R3399 gnd.n6082 gnd.n6081 585
R3400 gnd.n6085 gnd.n6084 585
R3401 gnd.n6087 gnd.n6086 585
R3402 gnd.n6089 gnd.n6088 585
R3403 gnd.n6091 gnd.n6090 585
R3404 gnd.n6093 gnd.n6092 585
R3405 gnd.n6095 gnd.n6094 585
R3406 gnd.n6097 gnd.n6096 585
R3407 gnd.n6099 gnd.n6098 585
R3408 gnd.n6101 gnd.n6100 585
R3409 gnd.n6103 gnd.n6102 585
R3410 gnd.n6105 gnd.n6104 585
R3411 gnd.n6107 gnd.n6106 585
R3412 gnd.n6109 gnd.n6108 585
R3413 gnd.n6111 gnd.n6110 585
R3414 gnd.n6112 gnd.n1287 585
R3415 gnd.n6114 gnd.n6113 585
R3416 gnd.n1288 gnd.n1286 585
R3417 gnd.n1289 gnd.n1137 585
R3418 gnd.n6116 gnd.n1137 585
R3419 gnd.n6195 gnd.n1139 585
R3420 gnd.n6199 gnd.n1139 585
R3421 gnd.n6194 gnd.n6193 585
R3422 gnd.n6193 gnd.n6192 585
R3423 gnd.n1145 gnd.n1129 585
R3424 gnd.n6205 gnd.n1129 585
R3425 gnd.n4397 gnd.n4396 585
R3426 gnd.n4398 gnd.n4397 585
R3427 gnd.n4395 gnd.n1119 585
R3428 gnd.n6211 gnd.n1119 585
R3429 gnd.n4394 gnd.n4393 585
R3430 gnd.n4393 gnd.n4392 585
R3431 gnd.n4390 gnd.n1108 585
R3432 gnd.n6217 gnd.n1108 585
R3433 gnd.n4389 gnd.n2339 585
R3434 gnd.n4409 gnd.n2339 585
R3435 gnd.n4388 gnd.n1099 585
R3436 gnd.n6223 gnd.n1099 585
R3437 gnd.n4387 gnd.n4386 585
R3438 gnd.n4386 gnd.n4385 585
R3439 gnd.n2345 gnd.n1088 585
R3440 gnd.n6229 gnd.n1088 585
R3441 gnd.n4376 gnd.n4375 585
R3442 gnd.n4377 gnd.n4376 585
R3443 gnd.n4374 gnd.n1079 585
R3444 gnd.n6235 gnd.n1079 585
R3445 gnd.n4373 gnd.n4372 585
R3446 gnd.n4372 gnd.n4371 585
R3447 gnd.n2351 gnd.n1068 585
R3448 gnd.n6241 gnd.n1068 585
R3449 gnd.n4303 gnd.n2356 585
R3450 gnd.n4363 gnd.n2356 585
R3451 gnd.n4304 gnd.n1059 585
R3452 gnd.n6247 gnd.n1059 585
R3453 gnd.n4306 gnd.n4305 585
R3454 gnd.n4307 gnd.n4306 585
R3455 gnd.n4301 gnd.n1051 585
R3456 gnd.n6254 gnd.n1051 585
R3457 gnd.n4300 gnd.n2388 585
R3458 gnd.n4315 gnd.n2388 585
R3459 gnd.n4299 gnd.n1042 585
R3460 gnd.n6260 gnd.n1042 585
R3461 gnd.n4298 gnd.n4297 585
R3462 gnd.n4297 gnd.n4296 585
R3463 gnd.n4290 gnd.n1034 585
R3464 gnd.n6267 gnd.n1034 585
R3465 gnd.n4289 gnd.n2378 585
R3466 gnd.n4326 gnd.n2378 585
R3467 gnd.n4288 gnd.n1023 585
R3468 gnd.n6273 gnd.n1023 585
R3469 gnd.n4287 gnd.n2371 585
R3470 gnd.n4332 gnd.n2371 585
R3471 gnd.n4284 gnd.n4283 585
R3472 gnd.n4283 gnd.n2370 585
R3473 gnd.n4282 gnd.n1012 585
R3474 gnd.n6281 gnd.n1012 585
R3475 gnd.n4281 gnd.n4280 585
R3476 gnd.n4280 gnd.n4279 585
R3477 gnd.n2392 gnd.n1003 585
R3478 gnd.n6287 gnd.n1003 585
R3479 gnd.n4266 gnd.n4265 585
R3480 gnd.n4267 gnd.n4266 585
R3481 gnd.n4263 gnd.n992 585
R3482 gnd.n6293 gnd.n992 585
R3483 gnd.n4262 gnd.n4261 585
R3484 gnd.n4261 gnd.n4260 585
R3485 gnd.n2396 gnd.n981 585
R3486 gnd.n6299 gnd.n981 585
R3487 gnd.n4251 gnd.n4250 585
R3488 gnd.n4252 gnd.n4251 585
R3489 gnd.n2419 gnd.n968 585
R3490 gnd.n6305 gnd.n968 585
R3491 gnd.n4226 gnd.n4225 585
R3492 gnd.n4225 gnd.n967 585
R3493 gnd.n4227 gnd.n2424 585
R3494 gnd.n4243 gnd.n2424 585
R3495 gnd.n4229 gnd.n4228 585
R3496 gnd.n4228 gnd.n2434 585
R3497 gnd.n4224 gnd.n2432 585
R3498 gnd.n4234 gnd.n2432 585
R3499 gnd.n4223 gnd.n4222 585
R3500 gnd.n4222 gnd.n2431 585
R3501 gnd.n4221 gnd.n2439 585
R3502 gnd.n4221 gnd.n4220 585
R3503 gnd.n4094 gnd.n2441 585
R3504 gnd.n2442 gnd.n2441 585
R3505 gnd.n7285 gnd.n7284 585
R3506 gnd.n7284 gnd.n7283 585
R3507 gnd.n7286 gnd.n161 585
R3508 gnd.n167 gnd.n161 585
R3509 gnd.n7288 gnd.n7287 585
R3510 gnd.n7289 gnd.n7288 585
R3511 gnd.n148 gnd.n147 585
R3512 gnd.n152 gnd.n148 585
R3513 gnd.n7297 gnd.n7296 585
R3514 gnd.n7296 gnd.n7295 585
R3515 gnd.n7298 gnd.n142 585
R3516 gnd.n142 gnd.n141 585
R3517 gnd.n7300 gnd.n7299 585
R3518 gnd.n7301 gnd.n7300 585
R3519 gnd.n127 gnd.n126 585
R3520 gnd.n7266 gnd.n127 585
R3521 gnd.n7309 gnd.n7308 585
R3522 gnd.n7308 gnd.n7307 585
R3523 gnd.n7310 gnd.n121 585
R3524 gnd.n7174 gnd.n121 585
R3525 gnd.n7312 gnd.n7311 585
R3526 gnd.n7313 gnd.n7312 585
R3527 gnd.n107 gnd.n106 585
R3528 gnd.n7167 gnd.n107 585
R3529 gnd.n7321 gnd.n7320 585
R3530 gnd.n7320 gnd.n7319 585
R3531 gnd.n7322 gnd.n102 585
R3532 gnd.n7159 gnd.n102 585
R3533 gnd.n7324 gnd.n7323 585
R3534 gnd.n7325 gnd.n7324 585
R3535 gnd.n85 gnd.n83 585
R3536 gnd.n7152 gnd.n85 585
R3537 gnd.n7333 gnd.n7332 585
R3538 gnd.n7332 gnd.n7331 585
R3539 gnd.n84 gnd.n76 585
R3540 gnd.n7144 gnd.n84 585
R3541 gnd.n7336 gnd.n74 585
R3542 gnd.n7137 gnd.n74 585
R3543 gnd.n7338 gnd.n7337 585
R3544 gnd.n7339 gnd.n7338 585
R3545 gnd.n1712 gnd.n73 585
R3546 gnd.n5785 gnd.n73 585
R3547 gnd.n5793 gnd.n1713 585
R3548 gnd.n5793 gnd.n5792 585
R3549 gnd.n5796 gnd.n5795 585
R3550 gnd.n5797 gnd.n5796 585
R3551 gnd.n5794 gnd.n1711 585
R3552 gnd.n1711 gnd.n1706 585
R3553 gnd.n1695 gnd.n1694 585
R3554 gnd.n1699 gnd.n1694 585
R3555 gnd.n5807 gnd.n1696 585
R3556 gnd.n5807 gnd.n5806 585
R3557 gnd.n5809 gnd.n5808 585
R3558 gnd.n5810 gnd.n5809 585
R3559 gnd.n1680 gnd.n1679 585
R3560 gnd.n5767 gnd.n1680 585
R3561 gnd.n5818 gnd.n5817 585
R3562 gnd.n5817 gnd.n5816 585
R3563 gnd.n5819 gnd.n1674 585
R3564 gnd.n5749 gnd.n1674 585
R3565 gnd.n5821 gnd.n5820 585
R3566 gnd.n5822 gnd.n5821 585
R3567 gnd.n1660 gnd.n1659 585
R3568 gnd.n5742 gnd.n1660 585
R3569 gnd.n5830 gnd.n5829 585
R3570 gnd.n5829 gnd.n5828 585
R3571 gnd.n5831 gnd.n1654 585
R3572 gnd.n5686 gnd.n1654 585
R3573 gnd.n5833 gnd.n5832 585
R3574 gnd.n5834 gnd.n5833 585
R3575 gnd.n1640 gnd.n1639 585
R3576 gnd.n5697 gnd.n1640 585
R3577 gnd.n5842 gnd.n5841 585
R3578 gnd.n5841 gnd.n5840 585
R3579 gnd.n5843 gnd.n1634 585
R3580 gnd.n5677 gnd.n1634 585
R3581 gnd.n5845 gnd.n5844 585
R3582 gnd.n5846 gnd.n5845 585
R3583 gnd.n1617 gnd.n1616 585
R3584 gnd.n5669 gnd.n1617 585
R3585 gnd.n5854 gnd.n5853 585
R3586 gnd.n5853 gnd.n5852 585
R3587 gnd.n5855 gnd.n1612 585
R3588 gnd.n5121 gnd.n1612 585
R3589 gnd.n5857 gnd.n5856 585
R3590 gnd.n5858 gnd.n5857 585
R3591 gnd.n5510 gnd.n1611 585
R3592 gnd.n5515 gnd.n5513 585
R3593 gnd.n5516 gnd.n5509 585
R3594 gnd.n5516 gnd.n1598 585
R3595 gnd.n5519 gnd.n5518 585
R3596 gnd.n5507 gnd.n5506 585
R3597 gnd.n5524 gnd.n5523 585
R3598 gnd.n5526 gnd.n5505 585
R3599 gnd.n5529 gnd.n5528 585
R3600 gnd.n5503 gnd.n5502 585
R3601 gnd.n5534 gnd.n5533 585
R3602 gnd.n5536 gnd.n5501 585
R3603 gnd.n5539 gnd.n5538 585
R3604 gnd.n5499 gnd.n5498 585
R3605 gnd.n5544 gnd.n5543 585
R3606 gnd.n5546 gnd.n5497 585
R3607 gnd.n5549 gnd.n5548 585
R3608 gnd.n5495 gnd.n5494 585
R3609 gnd.n5557 gnd.n5556 585
R3610 gnd.n5559 gnd.n5493 585
R3611 gnd.n5562 gnd.n5561 585
R3612 gnd.n5491 gnd.n5490 585
R3613 gnd.n5567 gnd.n5566 585
R3614 gnd.n5569 gnd.n5489 585
R3615 gnd.n5572 gnd.n5571 585
R3616 gnd.n5487 gnd.n5486 585
R3617 gnd.n5578 gnd.n5577 585
R3618 gnd.n5582 gnd.n1786 585
R3619 gnd.n5585 gnd.n5584 585
R3620 gnd.n1784 gnd.n1783 585
R3621 gnd.n5590 gnd.n5589 585
R3622 gnd.n5592 gnd.n1782 585
R3623 gnd.n5595 gnd.n5594 585
R3624 gnd.n1780 gnd.n1779 585
R3625 gnd.n5600 gnd.n5599 585
R3626 gnd.n5602 gnd.n1778 585
R3627 gnd.n5607 gnd.n5604 585
R3628 gnd.n1776 gnd.n1775 585
R3629 gnd.n5612 gnd.n5611 585
R3630 gnd.n5614 gnd.n1774 585
R3631 gnd.n5617 gnd.n5616 585
R3632 gnd.n1772 gnd.n1771 585
R3633 gnd.n5622 gnd.n5621 585
R3634 gnd.n5624 gnd.n1770 585
R3635 gnd.n5627 gnd.n5626 585
R3636 gnd.n1768 gnd.n1767 585
R3637 gnd.n5632 gnd.n5631 585
R3638 gnd.n5634 gnd.n1766 585
R3639 gnd.n5637 gnd.n5636 585
R3640 gnd.n1764 gnd.n1763 585
R3641 gnd.n5642 gnd.n5641 585
R3642 gnd.n5644 gnd.n1762 585
R3643 gnd.n5647 gnd.n5646 585
R3644 gnd.n1760 gnd.n1759 585
R3645 gnd.n5653 gnd.n5652 585
R3646 gnd.n5655 gnd.n1758 585
R3647 gnd.n5656 gnd.n1757 585
R3648 gnd.n5659 gnd.n5658 585
R3649 gnd.n383 gnd.n382 585
R3650 gnd.n380 gnd.n176 585
R3651 gnd.n379 gnd.n378 585
R3652 gnd.n372 gnd.n178 585
R3653 gnd.n374 gnd.n373 585
R3654 gnd.n370 gnd.n180 585
R3655 gnd.n369 gnd.n368 585
R3656 gnd.n362 gnd.n182 585
R3657 gnd.n364 gnd.n363 585
R3658 gnd.n360 gnd.n184 585
R3659 gnd.n359 gnd.n358 585
R3660 gnd.n352 gnd.n186 585
R3661 gnd.n354 gnd.n353 585
R3662 gnd.n350 gnd.n188 585
R3663 gnd.n349 gnd.n348 585
R3664 gnd.n342 gnd.n190 585
R3665 gnd.n344 gnd.n343 585
R3666 gnd.n340 gnd.n192 585
R3667 gnd.n339 gnd.n338 585
R3668 gnd.n332 gnd.n194 585
R3669 gnd.n334 gnd.n333 585
R3670 gnd.n330 gnd.n198 585
R3671 gnd.n329 gnd.n328 585
R3672 gnd.n322 gnd.n200 585
R3673 gnd.n324 gnd.n323 585
R3674 gnd.n320 gnd.n202 585
R3675 gnd.n319 gnd.n318 585
R3676 gnd.n312 gnd.n204 585
R3677 gnd.n314 gnd.n313 585
R3678 gnd.n310 gnd.n206 585
R3679 gnd.n309 gnd.n308 585
R3680 gnd.n302 gnd.n208 585
R3681 gnd.n304 gnd.n303 585
R3682 gnd.n300 gnd.n210 585
R3683 gnd.n299 gnd.n298 585
R3684 gnd.n292 gnd.n212 585
R3685 gnd.n294 gnd.n293 585
R3686 gnd.n290 gnd.n214 585
R3687 gnd.n289 gnd.n288 585
R3688 gnd.n282 gnd.n216 585
R3689 gnd.n284 gnd.n283 585
R3690 gnd.n280 gnd.n279 585
R3691 gnd.n278 gnd.n221 585
R3692 gnd.n272 gnd.n222 585
R3693 gnd.n274 gnd.n273 585
R3694 gnd.n269 gnd.n224 585
R3695 gnd.n268 gnd.n267 585
R3696 gnd.n261 gnd.n226 585
R3697 gnd.n263 gnd.n262 585
R3698 gnd.n259 gnd.n228 585
R3699 gnd.n258 gnd.n257 585
R3700 gnd.n251 gnd.n230 585
R3701 gnd.n253 gnd.n252 585
R3702 gnd.n249 gnd.n232 585
R3703 gnd.n248 gnd.n247 585
R3704 gnd.n241 gnd.n234 585
R3705 gnd.n243 gnd.n242 585
R3706 gnd.n239 gnd.n238 585
R3707 gnd.n237 gnd.n166 585
R3708 gnd.n170 gnd.n166 585
R3709 gnd.n7279 gnd.n168 585
R3710 gnd.n7283 gnd.n168 585
R3711 gnd.n7278 gnd.n7277 585
R3712 gnd.n7277 gnd.n167 585
R3713 gnd.n7276 gnd.n159 585
R3714 gnd.n7289 gnd.n159 585
R3715 gnd.n7275 gnd.n7274 585
R3716 gnd.n7274 gnd.n152 585
R3717 gnd.n7273 gnd.n150 585
R3718 gnd.n7295 gnd.n150 585
R3719 gnd.n7272 gnd.n7271 585
R3720 gnd.n7271 gnd.n141 585
R3721 gnd.n7269 gnd.n139 585
R3722 gnd.n7301 gnd.n139 585
R3723 gnd.n7268 gnd.n7267 585
R3724 gnd.n7267 gnd.n7266 585
R3725 gnd.n386 gnd.n129 585
R3726 gnd.n7307 gnd.n129 585
R3727 gnd.n7173 gnd.n7172 585
R3728 gnd.n7174 gnd.n7173 585
R3729 gnd.n7170 gnd.n118 585
R3730 gnd.n7313 gnd.n118 585
R3731 gnd.n7169 gnd.n7168 585
R3732 gnd.n7168 gnd.n7167 585
R3733 gnd.n390 gnd.n109 585
R3734 gnd.n7319 gnd.n109 585
R3735 gnd.n7158 gnd.n7157 585
R3736 gnd.n7159 gnd.n7158 585
R3737 gnd.n7155 gnd.n99 585
R3738 gnd.n7325 gnd.n99 585
R3739 gnd.n7154 gnd.n7153 585
R3740 gnd.n7153 gnd.n7152 585
R3741 gnd.n395 gnd.n87 585
R3742 gnd.n7331 gnd.n87 585
R3743 gnd.n7143 gnd.n7142 585
R3744 gnd.n7144 gnd.n7143 585
R3745 gnd.n399 gnd.n398 585
R3746 gnd.n7137 gnd.n398 585
R3747 gnd.n5784 gnd.n70 585
R3748 gnd.n7339 gnd.n70 585
R3749 gnd.n5787 gnd.n5786 585
R3750 gnd.n5786 gnd.n5785 585
R3751 gnd.n5783 gnd.n1714 585
R3752 gnd.n5792 gnd.n1714 585
R3753 gnd.n5782 gnd.n1707 585
R3754 gnd.n5797 gnd.n1707 585
R3755 gnd.n5772 gnd.n1726 585
R3756 gnd.n5772 gnd.n1706 585
R3757 gnd.n5774 gnd.n5773 585
R3758 gnd.n5773 gnd.n1699 585
R3759 gnd.n5771 gnd.n1697 585
R3760 gnd.n5806 gnd.n1697 585
R3761 gnd.n5770 gnd.n1691 585
R3762 gnd.n5810 gnd.n1691 585
R3763 gnd.n5769 gnd.n5768 585
R3764 gnd.n5768 gnd.n5767 585
R3765 gnd.n1728 gnd.n1682 585
R3766 gnd.n5816 gnd.n1682 585
R3767 gnd.n5748 gnd.n5747 585
R3768 gnd.n5749 gnd.n5748 585
R3769 gnd.n5745 gnd.n1671 585
R3770 gnd.n5822 gnd.n1671 585
R3771 gnd.n5744 gnd.n5743 585
R3772 gnd.n5743 gnd.n5742 585
R3773 gnd.n1734 gnd.n1662 585
R3774 gnd.n5828 gnd.n1662 585
R3775 gnd.n5685 gnd.n5684 585
R3776 gnd.n5686 gnd.n5685 585
R3777 gnd.n5682 gnd.n1651 585
R3778 gnd.n5834 gnd.n1651 585
R3779 gnd.n5681 gnd.n1741 585
R3780 gnd.n5697 gnd.n1741 585
R3781 gnd.n5680 gnd.n1642 585
R3782 gnd.n5840 gnd.n1642 585
R3783 gnd.n5679 gnd.n5678 585
R3784 gnd.n5678 gnd.n5677 585
R3785 gnd.n1746 gnd.n1631 585
R3786 gnd.n5846 gnd.n1631 585
R3787 gnd.n5668 gnd.n5667 585
R3788 gnd.n5669 gnd.n5668 585
R3789 gnd.n5666 gnd.n1619 585
R3790 gnd.n5852 gnd.n1619 585
R3791 gnd.n5665 gnd.n1752 585
R3792 gnd.n5121 gnd.n1752 585
R3793 gnd.n1751 gnd.n1607 585
R3794 gnd.n5858 gnd.n1607 585
R3795 gnd.n6311 gnd.n961 585
R3796 gnd.n2423 gnd.n961 585
R3797 gnd.n7116 gnd.n7115 585
R3798 gnd.n7116 gnd.n149 585
R3799 gnd.n7117 gnd.n418 585
R3800 gnd.n7117 gnd.n138 585
R3801 gnd.n7119 gnd.n7118 585
R3802 gnd.n7118 gnd.n131 585
R3803 gnd.n7120 gnd.n413 585
R3804 gnd.n413 gnd.n128 585
R3805 gnd.n7122 gnd.n7121 585
R3806 gnd.n7122 gnd.n120 585
R3807 gnd.n7123 gnd.n412 585
R3808 gnd.n7123 gnd.n117 585
R3809 gnd.n7125 gnd.n7124 585
R3810 gnd.n7124 gnd.n391 585
R3811 gnd.n7126 gnd.n407 585
R3812 gnd.n407 gnd.n108 585
R3813 gnd.n7128 gnd.n7127 585
R3814 gnd.n7128 gnd.n101 585
R3815 gnd.n7129 gnd.n406 585
R3816 gnd.n7129 gnd.n98 585
R3817 gnd.n7131 gnd.n7130 585
R3818 gnd.n7130 gnd.n89 585
R3819 gnd.n7132 gnd.n403 585
R3820 gnd.n403 gnd.n86 585
R3821 gnd.n7135 gnd.n7134 585
R3822 gnd.n7136 gnd.n7135 585
R3823 gnd.n404 gnd.n402 585
R3824 gnd.n402 gnd.n71 585
R3825 gnd.n1719 gnd.n1716 585
R3826 gnd.n1716 gnd.n69 585
R3827 gnd.n1721 gnd.n1720 585
R3828 gnd.n1722 gnd.n1721 585
R3829 gnd.n1704 gnd.n1703 585
R3830 gnd.n1709 gnd.n1704 585
R3831 gnd.n5800 gnd.n5799 585
R3832 gnd.n5799 gnd.n5798 585
R3833 gnd.n5802 gnd.n1701 585
R3834 gnd.n1705 gnd.n1701 585
R3835 gnd.n5804 gnd.n5803 585
R3836 gnd.n5805 gnd.n5804 585
R3837 gnd.n5732 gnd.n1700 585
R3838 gnd.n1700 gnd.n1693 585
R3839 gnd.n5734 gnd.n5733 585
R3840 gnd.n5734 gnd.n1690 585
R3841 gnd.n5735 gnd.n5729 585
R3842 gnd.n5735 gnd.n1729 585
R3843 gnd.n5737 gnd.n5736 585
R3844 gnd.n5736 gnd.n1681 585
R3845 gnd.n5738 gnd.n1737 585
R3846 gnd.n1737 gnd.n1673 585
R3847 gnd.n5740 gnd.n5739 585
R3848 gnd.n5741 gnd.n5740 585
R3849 gnd.n1738 gnd.n1736 585
R3850 gnd.n1736 gnd.n1664 585
R3851 gnd.n5723 gnd.n5722 585
R3852 gnd.n5722 gnd.n1661 585
R3853 gnd.n5721 gnd.n1740 585
R3854 gnd.n5721 gnd.n1653 585
R3855 gnd.n5720 gnd.n5719 585
R3856 gnd.n5720 gnd.n1650 585
R3857 gnd.n5700 gnd.n5699 585
R3858 gnd.n5699 gnd.n5698 585
R3859 gnd.n5715 gnd.n5714 585
R3860 gnd.n5714 gnd.n1641 585
R3861 gnd.n5713 gnd.n5702 585
R3862 gnd.n5713 gnd.n1633 585
R3863 gnd.n5712 gnd.n5711 585
R3864 gnd.n5712 gnd.n1630 585
R3865 gnd.n5704 gnd.n5703 585
R3866 gnd.n5703 gnd.n1621 585
R3867 gnd.n5707 gnd.n5706 585
R3868 gnd.n5706 gnd.n1618 585
R3869 gnd.n1605 gnd.n1604 585
R3870 gnd.n1609 gnd.n1605 585
R3871 gnd.n5861 gnd.n5860 585
R3872 gnd.n5860 gnd.n5859 585
R3873 gnd.n5862 gnd.n1599 585
R3874 gnd.n1606 gnd.n1599 585
R3875 gnd.n5864 gnd.n5863 585
R3876 gnd.n5865 gnd.n5864 585
R3877 gnd.n1596 gnd.n1595 585
R3878 gnd.n5866 gnd.n1596 585
R3879 gnd.n5869 gnd.n5868 585
R3880 gnd.n5868 gnd.n5867 585
R3881 gnd.n5870 gnd.n1590 585
R3882 gnd.n1590 gnd.n1588 585
R3883 gnd.n5872 gnd.n5871 585
R3884 gnd.n5873 gnd.n5872 585
R3885 gnd.n1591 gnd.n1589 585
R3886 gnd.n1589 gnd.n1586 585
R3887 gnd.n1859 gnd.n1858 585
R3888 gnd.n5302 gnd.n1859 585
R3889 gnd.n5306 gnd.n5305 585
R3890 gnd.n5305 gnd.n5304 585
R3891 gnd.n5307 gnd.n1849 585
R3892 gnd.n1860 gnd.n1849 585
R3893 gnd.n5309 gnd.n5308 585
R3894 gnd.n5310 gnd.n5309 585
R3895 gnd.n1850 gnd.n1844 585
R3896 gnd.n5313 gnd.n1844 585
R3897 gnd.n5316 gnd.n1843 585
R3898 gnd.n5316 gnd.n5315 585
R3899 gnd.n5318 gnd.n5317 585
R3900 gnd.n5317 gnd.n1791 585
R3901 gnd.n5319 gnd.n1838 585
R3902 gnd.n1838 gnd.n1828 585
R3903 gnd.n5321 gnd.n5320 585
R3904 gnd.n5322 gnd.n5321 585
R3905 gnd.n1839 gnd.n1837 585
R3906 gnd.n1837 gnd.n1833 585
R3907 gnd.n5073 gnd.n1887 585
R3908 gnd.n1887 gnd.n1886 585
R3909 gnd.n5075 gnd.n5074 585
R3910 gnd.n5076 gnd.n5075 585
R3911 gnd.n1888 gnd.n1885 585
R3912 gnd.n1885 gnd.n1882 585
R3913 gnd.n5067 gnd.n5066 585
R3914 gnd.n5066 gnd.n5065 585
R3915 gnd.n1891 gnd.n1890 585
R3916 gnd.n5053 gnd.n1891 585
R3917 gnd.n5028 gnd.n1917 585
R3918 gnd.n1917 gnd.n1909 585
R3919 gnd.n5030 gnd.n5029 585
R3920 gnd.n5031 gnd.n5030 585
R3921 gnd.n1918 gnd.n1916 585
R3922 gnd.n5018 gnd.n1916 585
R3923 gnd.n5023 gnd.n5022 585
R3924 gnd.n5022 gnd.n5021 585
R3925 gnd.n1921 gnd.n1920 585
R3926 gnd.n1933 gnd.n1921 585
R3927 gnd.n5002 gnd.n5001 585
R3928 gnd.n5003 gnd.n5002 585
R3929 gnd.n1938 gnd.n1937 585
R3930 gnd.n1945 gnd.n1937 585
R3931 gnd.n4997 gnd.n4996 585
R3932 gnd.n4996 gnd.n4995 585
R3933 gnd.n1941 gnd.n1940 585
R3934 gnd.n4892 gnd.n1941 585
R3935 gnd.n4951 gnd.n1965 585
R3936 gnd.n1965 gnd.n1958 585
R3937 gnd.n4953 gnd.n4952 585
R3938 gnd.n4954 gnd.n4953 585
R3939 gnd.n1966 gnd.n1964 585
R3940 gnd.n1964 gnd.n1962 585
R3941 gnd.n4946 gnd.n4945 585
R3942 gnd.n4945 gnd.n4944 585
R3943 gnd.n1969 gnd.n1968 585
R3944 gnd.n4936 gnd.n1969 585
R3945 gnd.n4922 gnd.n4921 585
R3946 gnd.n4923 gnd.n4922 585
R3947 gnd.n1988 gnd.n1987 585
R3948 gnd.n4872 gnd.n1987 585
R3949 gnd.n4917 gnd.n4916 585
R3950 gnd.n4916 gnd.n4915 585
R3951 gnd.n1991 gnd.n1990 585
R3952 gnd.n1999 gnd.n1991 585
R3953 gnd.n4862 gnd.n4861 585
R3954 gnd.n4863 gnd.n4862 585
R3955 gnd.n2008 gnd.n2007 585
R3956 gnd.n2007 gnd.n2004 585
R3957 gnd.n4857 gnd.n4856 585
R3958 gnd.n4856 gnd.n4855 585
R3959 gnd.n2011 gnd.n2010 585
R3960 gnd.n2017 gnd.n2011 585
R3961 gnd.n4837 gnd.n4836 585
R3962 gnd.n4838 gnd.n4837 585
R3963 gnd.n2028 gnd.n2027 585
R3964 gnd.n2035 gnd.n2027 585
R3965 gnd.n4832 gnd.n4831 585
R3966 gnd.n4831 gnd.n4830 585
R3967 gnd.n2031 gnd.n2030 585
R3968 gnd.n2039 gnd.n2031 585
R3969 gnd.n4780 gnd.n4779 585
R3970 gnd.n4781 gnd.n4780 585
R3971 gnd.n2050 gnd.n2049 585
R3972 gnd.n2068 gnd.n2049 585
R3973 gnd.n4775 gnd.n4774 585
R3974 gnd.n4774 gnd.n4773 585
R3975 gnd.n2053 gnd.n2052 585
R3976 gnd.n2061 gnd.n2053 585
R3977 gnd.n4740 gnd.n4739 585
R3978 gnd.n4741 gnd.n4740 585
R3979 gnd.n2073 gnd.n2072 585
R3980 gnd.n2088 gnd.n2072 585
R3981 gnd.n4735 gnd.n4734 585
R3982 gnd.n4734 gnd.n4733 585
R3983 gnd.n2076 gnd.n2075 585
R3984 gnd.n4723 gnd.n2076 585
R3985 gnd.n4690 gnd.n2105 585
R3986 gnd.n2105 gnd.n2097 585
R3987 gnd.n4692 gnd.n4691 585
R3988 gnd.n4693 gnd.n4692 585
R3989 gnd.n2106 gnd.n2104 585
R3990 gnd.n2104 gnd.n2101 585
R3991 gnd.n4685 gnd.n4684 585
R3992 gnd.n4684 gnd.n4683 585
R3993 gnd.n2109 gnd.n2108 585
R3994 gnd.n2115 gnd.n2109 585
R3995 gnd.n4662 gnd.n4661 585
R3996 gnd.n4663 gnd.n4662 585
R3997 gnd.n2124 gnd.n2123 585
R3998 gnd.n2130 gnd.n2123 585
R3999 gnd.n4657 gnd.n4656 585
R4000 gnd.n4656 gnd.n4655 585
R4001 gnd.n2127 gnd.n2126 585
R4002 gnd.n2134 gnd.n2127 585
R4003 gnd.n4600 gnd.n2149 585
R4004 gnd.n2149 gnd.n2139 585
R4005 gnd.n4602 gnd.n4601 585
R4006 gnd.n4603 gnd.n4602 585
R4007 gnd.n2150 gnd.n2148 585
R4008 gnd.n4568 gnd.n2148 585
R4009 gnd.n4595 gnd.n4594 585
R4010 gnd.n4594 gnd.n4593 585
R4011 gnd.n2153 gnd.n2152 585
R4012 gnd.n4576 gnd.n2153 585
R4013 gnd.n4558 gnd.n4557 585
R4014 gnd.n4559 gnd.n4558 585
R4015 gnd.n2168 gnd.n2167 585
R4016 gnd.n4536 gnd.n2167 585
R4017 gnd.n4553 gnd.n4552 585
R4018 gnd.n4552 gnd.n4551 585
R4019 gnd.n2171 gnd.n2170 585
R4020 gnd.n2178 gnd.n2171 585
R4021 gnd.n4515 gnd.n4514 585
R4022 gnd.n4516 gnd.n4515 585
R4023 gnd.n1489 gnd.n1488 585
R4024 gnd.n2192 gnd.n1489 585
R4025 gnd.n5987 gnd.n5986 585
R4026 gnd.n5986 gnd.n5985 585
R4027 gnd.n5988 gnd.n1483 585
R4028 gnd.n2196 gnd.n1483 585
R4029 gnd.n5990 gnd.n5989 585
R4030 gnd.n5991 gnd.n5990 585
R4031 gnd.n1484 gnd.n1482 585
R4032 gnd.n2282 gnd.n1482 585
R4033 gnd.n4477 gnd.n2293 585
R4034 gnd.n2293 gnd.n1453 585
R4035 gnd.n4479 gnd.n4478 585
R4036 gnd.n4480 gnd.n4479 585
R4037 gnd.n2294 gnd.n2292 585
R4038 gnd.n2292 gnd.n2290 585
R4039 gnd.n4471 gnd.n4470 585
R4040 gnd.n4470 gnd.n4469 585
R4041 gnd.n2297 gnd.n2296 585
R4042 gnd.n2306 gnd.n2297 585
R4043 gnd.n4444 gnd.n2321 585
R4044 gnd.n2321 gnd.n2305 585
R4045 gnd.n4446 gnd.n4445 585
R4046 gnd.n4447 gnd.n4446 585
R4047 gnd.n2322 gnd.n2320 585
R4048 gnd.n2320 gnd.n2313 585
R4049 gnd.n4439 gnd.n4438 585
R4050 gnd.n4438 gnd.n4437 585
R4051 gnd.n4435 gnd.n2324 585
R4052 gnd.n4435 gnd.n1168 585
R4053 gnd.n4434 gnd.n4433 585
R4054 gnd.n4434 gnd.n1154 585
R4055 gnd.n2327 gnd.n2326 585
R4056 gnd.n2326 gnd.n2325 585
R4057 gnd.n4429 gnd.n4428 585
R4058 gnd.n4428 gnd.n1257 585
R4059 gnd.n4427 gnd.n2329 585
R4060 gnd.n4427 gnd.n1243 585
R4061 gnd.n4426 gnd.n4425 585
R4062 gnd.n4426 gnd.n1141 585
R4063 gnd.n2331 gnd.n2330 585
R4064 gnd.n2330 gnd.n1138 585
R4065 gnd.n4421 gnd.n4420 585
R4066 gnd.n4420 gnd.n1131 585
R4067 gnd.n4419 gnd.n2333 585
R4068 gnd.n4419 gnd.n1128 585
R4069 gnd.n4418 gnd.n4417 585
R4070 gnd.n4418 gnd.n1121 585
R4071 gnd.n2335 gnd.n2334 585
R4072 gnd.n2334 gnd.n1118 585
R4073 gnd.n4413 gnd.n4412 585
R4074 gnd.n4412 gnd.n1110 585
R4075 gnd.n4411 gnd.n2337 585
R4076 gnd.n4411 gnd.n4410 585
R4077 gnd.n4350 gnd.n2338 585
R4078 gnd.n2338 gnd.n1101 585
R4079 gnd.n4352 gnd.n4351 585
R4080 gnd.n4351 gnd.n1098 585
R4081 gnd.n4353 gnd.n4344 585
R4082 gnd.n4344 gnd.n1090 585
R4083 gnd.n4355 gnd.n4354 585
R4084 gnd.n4355 gnd.n1087 585
R4085 gnd.n4356 gnd.n4343 585
R4086 gnd.n4356 gnd.n2350 585
R4087 gnd.n4358 gnd.n4357 585
R4088 gnd.n4357 gnd.n1078 585
R4089 gnd.n4359 gnd.n2358 585
R4090 gnd.n2358 gnd.n1070 585
R4091 gnd.n4361 gnd.n4360 585
R4092 gnd.n4362 gnd.n4361 585
R4093 gnd.n2359 gnd.n2357 585
R4094 gnd.n2357 gnd.n1061 585
R4095 gnd.n2383 gnd.n2382 585
R4096 gnd.n2383 gnd.n1058 585
R4097 gnd.n2385 gnd.n2384 585
R4098 gnd.n2384 gnd.n1053 585
R4099 gnd.n2387 gnd.n2386 585
R4100 gnd.n2387 gnd.n1050 585
R4101 gnd.n4318 gnd.n4317 585
R4102 gnd.n4317 gnd.n4316 585
R4103 gnd.n4320 gnd.n4319 585
R4104 gnd.n4320 gnd.n1041 585
R4105 gnd.n4322 gnd.n4321 585
R4106 gnd.n4321 gnd.n1036 585
R4107 gnd.n4324 gnd.n4323 585
R4108 gnd.n4325 gnd.n4324 585
R4109 gnd.n2381 gnd.n2380 585
R4110 gnd.n2381 gnd.n1025 585
R4111 gnd.n2379 gnd.n2369 585
R4112 gnd.n2369 gnd.n1022 585
R4113 gnd.n4334 gnd.n2367 585
R4114 gnd.n4334 gnd.n4333 585
R4115 gnd.n4336 gnd.n4335 585
R4116 gnd.n4335 gnd.n1014 585
R4117 gnd.n2368 gnd.n2366 585
R4118 gnd.n4278 gnd.n2368 585
R4119 gnd.n2408 gnd.n2407 585
R4120 gnd.n2408 gnd.n1005 585
R4121 gnd.n2409 gnd.n2404 585
R4122 gnd.n2409 gnd.n1002 585
R4123 gnd.n2411 gnd.n2410 585
R4124 gnd.n2410 gnd.n994 585
R4125 gnd.n2412 gnd.n2398 585
R4126 gnd.n2398 gnd.n991 585
R4127 gnd.n2414 gnd.n2413 585
R4128 gnd.n2415 gnd.n2414 585
R4129 gnd.n2399 gnd.n2397 585
R4130 gnd.n2397 gnd.n980 585
R4131 gnd.n966 gnd.n965 585
R4132 gnd.n970 gnd.n966 585
R4133 gnd.n6308 gnd.n6307 585
R4134 gnd.n6307 gnd.n6306 585
R4135 gnd.n5876 gnd.n5875 585
R4136 gnd.n5875 gnd.n5874 585
R4137 gnd.n1584 gnd.n1582 585
R4138 gnd.n5301 gnd.n1584 585
R4139 gnd.n5880 gnd.n1581 585
R4140 gnd.n5303 gnd.n1581 585
R4141 gnd.n5881 gnd.n1580 585
R4142 gnd.n1861 gnd.n1580 585
R4143 gnd.n5882 gnd.n1579 585
R4144 gnd.n1848 gnd.n1579 585
R4145 gnd.n5311 gnd.n1577 585
R4146 gnd.n5312 gnd.n5311 585
R4147 gnd.n5886 gnd.n1576 585
R4148 gnd.n5314 gnd.n1576 585
R4149 gnd.n5887 gnd.n1575 585
R4150 gnd.n1845 gnd.n1575 585
R4151 gnd.n5888 gnd.n1574 585
R4152 gnd.n5106 gnd.n1574 585
R4153 gnd.n5103 gnd.n1572 585
R4154 gnd.n5104 gnd.n5103 585
R4155 gnd.n5892 gnd.n1571 585
R4156 gnd.n5323 gnd.n1571 585
R4157 gnd.n5893 gnd.n1570 585
R4158 gnd.n5096 gnd.n1570 585
R4159 gnd.n5894 gnd.n1569 585
R4160 gnd.n1877 gnd.n1569 585
R4161 gnd.n5078 gnd.n1567 585
R4162 gnd.n5079 gnd.n5078 585
R4163 gnd.n5898 gnd.n1566 585
R4164 gnd.n5063 gnd.n1566 585
R4165 gnd.n5899 gnd.n1565 585
R4166 gnd.n1902 gnd.n1565 585
R4167 gnd.n5900 gnd.n1564 585
R4168 gnd.n5054 gnd.n1564 585
R4169 gnd.n1907 gnd.n1562 585
R4170 gnd.n1908 gnd.n1907 585
R4171 gnd.n5904 gnd.n1561 585
R4172 gnd.n5033 gnd.n1561 585
R4173 gnd.n5905 gnd.n1560 585
R4174 gnd.n5020 gnd.n1560 585
R4175 gnd.n5906 gnd.n1559 585
R4176 gnd.n4971 gnd.n1559 585
R4177 gnd.n1935 gnd.n1557 585
R4178 gnd.n1936 gnd.n1935 585
R4179 gnd.n5910 gnd.n1556 585
R4180 gnd.n1931 gnd.n1556 585
R4181 gnd.n5911 gnd.n1555 585
R4182 gnd.n4994 gnd.n1555 585
R4183 gnd.n5912 gnd.n1554 585
R4184 gnd.n4986 gnd.n1554 585
R4185 gnd.n4893 gnd.n1552 585
R4186 gnd.n4894 gnd.n4893 585
R4187 gnd.n5916 gnd.n1551 585
R4188 gnd.n4963 gnd.n1551 585
R4189 gnd.n5917 gnd.n1550 585
R4190 gnd.n4955 gnd.n1550 585
R4191 gnd.n5918 gnd.n1549 585
R4192 gnd.n1971 gnd.n1549 585
R4193 gnd.n4933 gnd.n1547 585
R4194 gnd.n4934 gnd.n4933 585
R4195 gnd.n5922 gnd.n1546 585
R4196 gnd.n1975 gnd.n1546 585
R4197 gnd.n5923 gnd.n1545 585
R4198 gnd.n4924 gnd.n1545 585
R4199 gnd.n5924 gnd.n1544 585
R4200 gnd.n1993 gnd.n1544 585
R4201 gnd.n4802 gnd.n1542 585
R4202 gnd.n4803 gnd.n4802 585
R4203 gnd.n5928 gnd.n1541 585
R4204 gnd.n1998 gnd.n1541 585
R4205 gnd.n5929 gnd.n1540 585
R4206 gnd.n4865 gnd.n1540 585
R4207 gnd.n5930 gnd.n1539 585
R4208 gnd.n4854 gnd.n1539 585
R4209 gnd.n2018 gnd.n1537 585
R4210 gnd.n2019 gnd.n2018 585
R4211 gnd.n5934 gnd.n1536 585
R4212 gnd.n2026 gnd.n1536 585
R4213 gnd.n5935 gnd.n1535 585
R4214 gnd.n4794 gnd.n1535 585
R4215 gnd.n5936 gnd.n1534 585
R4216 gnd.n4829 gnd.n1534 585
R4217 gnd.n4820 gnd.n1532 585
R4218 gnd.n4821 gnd.n4820 585
R4219 gnd.n5940 gnd.n1531 585
R4220 gnd.n4782 gnd.n1531 585
R4221 gnd.n5941 gnd.n1530 585
R4222 gnd.n4753 gnd.n1530 585
R4223 gnd.n5942 gnd.n1529 585
R4224 gnd.n2056 gnd.n1529 585
R4225 gnd.n4761 gnd.n1527 585
R4226 gnd.n4762 gnd.n4761 585
R4227 gnd.n5946 gnd.n1526 585
R4228 gnd.n4742 gnd.n1526 585
R4229 gnd.n5947 gnd.n1525 585
R4230 gnd.n4715 gnd.n1525 585
R4231 gnd.n5948 gnd.n1524 585
R4232 gnd.n2079 gnd.n1524 585
R4233 gnd.n4706 gnd.n1522 585
R4234 gnd.n4707 gnd.n4706 585
R4235 gnd.n5952 gnd.n1521 585
R4236 gnd.n2084 gnd.n1521 585
R4237 gnd.n5953 gnd.n1520 585
R4238 gnd.n4703 gnd.n1520 585
R4239 gnd.n5954 gnd.n1519 585
R4240 gnd.n4695 gnd.n1519 585
R4241 gnd.n4681 gnd.n1517 585
R4242 gnd.n4682 gnd.n4681 585
R4243 gnd.n5958 gnd.n1516 585
R4244 gnd.n2116 gnd.n1516 585
R4245 gnd.n5959 gnd.n1515 585
R4246 gnd.n4613 gnd.n1515 585
R4247 gnd.n5960 gnd.n1514 585
R4248 gnd.n2121 gnd.n1514 585
R4249 gnd.n4653 gnd.n1512 585
R4250 gnd.n4654 gnd.n4653 585
R4251 gnd.n5964 gnd.n1511 585
R4252 gnd.n4645 gnd.n1511 585
R4253 gnd.n5965 gnd.n1510 585
R4254 gnd.n4632 gnd.n1510 585
R4255 gnd.n5966 gnd.n1509 585
R4256 gnd.n4583 gnd.n1509 585
R4257 gnd.n4604 gnd.n1507 585
R4258 gnd.n4605 gnd.n4604 585
R4259 gnd.n5970 gnd.n1506 585
R4260 gnd.n2156 gnd.n1506 585
R4261 gnd.n5971 gnd.n1505 585
R4262 gnd.n2154 gnd.n1505 585
R4263 gnd.n5972 gnd.n1504 585
R4264 gnd.n2161 gnd.n1504 585
R4265 gnd.n2165 gnd.n1502 585
R4266 gnd.n2166 gnd.n2165 585
R4267 gnd.n5976 gnd.n1501 585
R4268 gnd.n4534 gnd.n1501 585
R4269 gnd.n5977 gnd.n1500 585
R4270 gnd.n2185 gnd.n1500 585
R4271 gnd.n5978 gnd.n1499 585
R4272 gnd.n2177 gnd.n1499 585
R4273 gnd.n1496 gnd.n1494 585
R4274 gnd.n4518 gnd.n1494 585
R4275 gnd.n5983 gnd.n5982 585
R4276 gnd.n5984 gnd.n5983 585
R4277 gnd.n1495 gnd.n1493 585
R4278 gnd.n4503 gnd.n1493 585
R4279 gnd.n4487 gnd.n4486 585
R4280 gnd.n4486 gnd.n1481 585
R4281 gnd.n2286 gnd.n2284 585
R4282 gnd.n2284 gnd.n1479 585
R4283 gnd.n4492 gnd.n4491 585
R4284 gnd.n4493 gnd.n4492 585
R4285 gnd.n2285 gnd.n2283 585
R4286 gnd.n2283 gnd.n1421 585
R4287 gnd.n4483 gnd.n4482 585
R4288 gnd.n4482 gnd.n4481 585
R4289 gnd.n2289 gnd.n2288 585
R4290 gnd.n4468 gnd.n2289 585
R4291 gnd.n2310 gnd.n2308 585
R4292 gnd.n2308 gnd.n2298 585
R4293 gnd.n4456 gnd.n4455 585
R4294 gnd.n4457 gnd.n4456 585
R4295 gnd.n2309 gnd.n2307 585
R4296 gnd.n2319 gnd.n2307 585
R4297 gnd.n4450 gnd.n4449 585
R4298 gnd.n4449 gnd.n4448 585
R4299 gnd.n2312 gnd.n1171 585
R4300 gnd.n4436 gnd.n1171 585
R4301 gnd.n6179 gnd.n6178 585
R4302 gnd.n6177 gnd.n1170 585
R4303 gnd.n1173 gnd.n1169 585
R4304 gnd.n6181 gnd.n1169 585
R4305 gnd.n6173 gnd.n1175 585
R4306 gnd.n6172 gnd.n1176 585
R4307 gnd.n6171 gnd.n1177 585
R4308 gnd.n1180 gnd.n1178 585
R4309 gnd.n6166 gnd.n1181 585
R4310 gnd.n6165 gnd.n1182 585
R4311 gnd.n6164 gnd.n1183 585
R4312 gnd.n1192 gnd.n1184 585
R4313 gnd.n6157 gnd.n1193 585
R4314 gnd.n6156 gnd.n1194 585
R4315 gnd.n1196 gnd.n1195 585
R4316 gnd.n6149 gnd.n1202 585
R4317 gnd.n6148 gnd.n1203 585
R4318 gnd.n1210 gnd.n1204 585
R4319 gnd.n6141 gnd.n1211 585
R4320 gnd.n6140 gnd.n1212 585
R4321 gnd.n1214 gnd.n1213 585
R4322 gnd.n6133 gnd.n1220 585
R4323 gnd.n6132 gnd.n1221 585
R4324 gnd.n1228 gnd.n1222 585
R4325 gnd.n6125 gnd.n1229 585
R4326 gnd.n6124 gnd.n1230 585
R4327 gnd.n1235 gnd.n1234 585
R4328 gnd.n1166 gnd.n1151 585
R4329 gnd.n6185 gnd.n1152 585
R4330 gnd.n6184 gnd.n6183 585
R4331 gnd.n1864 gnd.n1587 585
R4332 gnd.n5874 gnd.n1587 585
R4333 gnd.n5300 gnd.n5299 585
R4334 gnd.n5301 gnd.n5300 585
R4335 gnd.n1863 gnd.n1862 585
R4336 gnd.n5303 gnd.n1862 585
R4337 gnd.n5117 gnd.n5116 585
R4338 gnd.n5116 gnd.n1861 585
R4339 gnd.n5115 gnd.n5114 585
R4340 gnd.n5115 gnd.n1848 585
R4341 gnd.n5113 gnd.n1847 585
R4342 gnd.n5312 gnd.n1847 585
R4343 gnd.n1866 gnd.n1846 585
R4344 gnd.n5314 gnd.n1846 585
R4345 gnd.n5109 gnd.n5108 585
R4346 gnd.n5108 gnd.n1845 585
R4347 gnd.n5107 gnd.n1868 585
R4348 gnd.n5107 gnd.n5106 585
R4349 gnd.n5105 gnd.n5102 585
R4350 gnd.n5105 gnd.n5104 585
R4351 gnd.n1869 gnd.n1835 585
R4352 gnd.n5323 gnd.n1835 585
R4353 gnd.n5098 gnd.n5097 585
R4354 gnd.n5097 gnd.n5096 585
R4355 gnd.n1872 gnd.n1871 585
R4356 gnd.n1877 gnd.n1872 585
R4357 gnd.n1896 gnd.n1884 585
R4358 gnd.n5079 gnd.n1884 585
R4359 gnd.n5062 gnd.n5061 585
R4360 gnd.n5063 gnd.n5062 585
R4361 gnd.n1895 gnd.n1894 585
R4362 gnd.n1902 gnd.n1894 585
R4363 gnd.n5056 gnd.n5055 585
R4364 gnd.n5055 gnd.n5054 585
R4365 gnd.n1899 gnd.n1898 585
R4366 gnd.n1908 gnd.n1899 585
R4367 gnd.n4974 gnd.n1915 585
R4368 gnd.n5033 gnd.n1915 585
R4369 gnd.n4973 gnd.n1923 585
R4370 gnd.n5020 gnd.n1923 585
R4371 gnd.n4978 gnd.n4972 585
R4372 gnd.n4972 gnd.n4971 585
R4373 gnd.n4979 gnd.n4970 585
R4374 gnd.n4970 gnd.n1936 585
R4375 gnd.n4980 gnd.n4969 585
R4376 gnd.n4969 gnd.n1931 585
R4377 gnd.n1952 gnd.n1943 585
R4378 gnd.n4994 gnd.n1943 585
R4379 gnd.n4985 gnd.n4984 585
R4380 gnd.n4986 gnd.n4985 585
R4381 gnd.n1951 gnd.n1950 585
R4382 gnd.n4894 gnd.n1950 585
R4383 gnd.n4965 gnd.n4964 585
R4384 gnd.n4964 gnd.n4963 585
R4385 gnd.n1955 gnd.n1954 585
R4386 gnd.n4955 gnd.n1955 585
R4387 gnd.n1981 gnd.n1979 585
R4388 gnd.n1979 gnd.n1971 585
R4389 gnd.n4932 gnd.n4931 585
R4390 gnd.n4934 gnd.n4932 585
R4391 gnd.n1980 gnd.n1978 585
R4392 gnd.n1978 gnd.n1975 585
R4393 gnd.n4926 gnd.n4925 585
R4394 gnd.n4925 gnd.n4924 585
R4395 gnd.n1984 gnd.n1983 585
R4396 gnd.n1993 gnd.n1984 585
R4397 gnd.n4806 gnd.n4804 585
R4398 gnd.n4804 gnd.n4803 585
R4399 gnd.n4807 gnd.n4800 585
R4400 gnd.n4800 gnd.n1998 585
R4401 gnd.n4808 gnd.n2006 585
R4402 gnd.n4865 gnd.n2006 585
R4403 gnd.n4798 gnd.n2013 585
R4404 gnd.n4854 gnd.n2013 585
R4405 gnd.n4812 gnd.n4797 585
R4406 gnd.n4797 gnd.n2019 585
R4407 gnd.n4813 gnd.n4796 585
R4408 gnd.n4796 gnd.n2026 585
R4409 gnd.n4814 gnd.n4795 585
R4410 gnd.n4795 gnd.n4794 585
R4411 gnd.n2043 gnd.n2033 585
R4412 gnd.n4829 gnd.n2033 585
R4413 gnd.n4819 gnd.n4818 585
R4414 gnd.n4821 gnd.n4819 585
R4415 gnd.n2042 gnd.n2041 585
R4416 gnd.n4782 gnd.n2041 585
R4417 gnd.n4755 gnd.n4754 585
R4418 gnd.n4754 gnd.n4753 585
R4419 gnd.n2066 gnd.n2064 585
R4420 gnd.n2064 gnd.n2056 585
R4421 gnd.n4760 gnd.n4759 585
R4422 gnd.n4762 gnd.n4760 585
R4423 gnd.n2065 gnd.n2063 585
R4424 gnd.n4742 gnd.n2063 585
R4425 gnd.n4714 gnd.n4713 585
R4426 gnd.n4715 gnd.n4714 585
R4427 gnd.n2090 gnd.n2089 585
R4428 gnd.n2089 gnd.n2079 585
R4429 gnd.n4709 gnd.n4708 585
R4430 gnd.n4708 gnd.n4707 585
R4431 gnd.n4705 gnd.n2092 585
R4432 gnd.n4705 gnd.n2084 585
R4433 gnd.n4704 gnd.n2094 585
R4434 gnd.n4704 gnd.n4703 585
R4435 gnd.n4619 gnd.n2093 585
R4436 gnd.n4695 gnd.n2093 585
R4437 gnd.n4620 gnd.n2111 585
R4438 gnd.n4682 gnd.n2111 585
R4439 gnd.n4616 gnd.n4615 585
R4440 gnd.n4615 gnd.n2116 585
R4441 gnd.n4624 gnd.n4614 585
R4442 gnd.n4614 gnd.n4613 585
R4443 gnd.n4625 gnd.n4611 585
R4444 gnd.n4611 gnd.n2121 585
R4445 gnd.n4626 gnd.n2128 585
R4446 gnd.n4654 gnd.n2128 585
R4447 gnd.n2142 gnd.n2136 585
R4448 gnd.n4645 gnd.n2136 585
R4449 gnd.n4631 gnd.n4630 585
R4450 gnd.n4632 gnd.n4631 585
R4451 gnd.n2141 gnd.n2140 585
R4452 gnd.n4583 gnd.n2140 585
R4453 gnd.n4607 gnd.n4606 585
R4454 gnd.n4606 gnd.n4605 585
R4455 gnd.n2145 gnd.n2144 585
R4456 gnd.n2156 gnd.n2145 585
R4457 gnd.n4527 gnd.n4526 585
R4458 gnd.n4526 gnd.n2154 585
R4459 gnd.n4528 gnd.n4525 585
R4460 gnd.n4525 gnd.n2161 585
R4461 gnd.n2189 gnd.n2187 585
R4462 gnd.n2187 gnd.n2166 585
R4463 gnd.n4533 gnd.n4532 585
R4464 gnd.n4534 gnd.n4533 585
R4465 gnd.n2188 gnd.n2186 585
R4466 gnd.n2186 gnd.n2185 585
R4467 gnd.n4521 gnd.n4520 585
R4468 gnd.n4520 gnd.n2177 585
R4469 gnd.n4519 gnd.n2191 585
R4470 gnd.n4519 gnd.n4518 585
R4471 gnd.n2200 gnd.n1491 585
R4472 gnd.n5984 gnd.n1491 585
R4473 gnd.n4502 gnd.n4501 585
R4474 gnd.n4503 gnd.n4502 585
R4475 gnd.n2199 gnd.n2198 585
R4476 gnd.n2198 gnd.n1481 585
R4477 gnd.n4496 gnd.n4495 585
R4478 gnd.n4495 gnd.n1479 585
R4479 gnd.n4494 gnd.n2202 585
R4480 gnd.n4494 gnd.n4493 585
R4481 gnd.n4462 gnd.n2203 585
R4482 gnd.n2203 gnd.n1421 585
R4483 gnd.n2301 gnd.n2291 585
R4484 gnd.n4481 gnd.n2291 585
R4485 gnd.n4467 gnd.n4466 585
R4486 gnd.n4468 gnd.n4467 585
R4487 gnd.n2300 gnd.n2299 585
R4488 gnd.n2299 gnd.n2298 585
R4489 gnd.n4459 gnd.n4458 585
R4490 gnd.n4458 gnd.n4457 585
R4491 gnd.n2304 gnd.n2303 585
R4492 gnd.n2319 gnd.n2304 585
R4493 gnd.n2318 gnd.n2317 585
R4494 gnd.n4448 gnd.n2318 585
R4495 gnd.n2314 gnd.n1153 585
R4496 gnd.n4436 gnd.n1153 585
R4497 gnd.n5274 gnd.n5129 585
R4498 gnd.n5129 gnd.n1597 585
R4499 gnd.n5275 gnd.n5272 585
R4500 gnd.n5270 gnd.n5147 585
R4501 gnd.n5269 gnd.n5268 585
R4502 gnd.n5253 gnd.n5149 585
R4503 gnd.n5255 gnd.n5254 585
R4504 gnd.n5251 gnd.n5156 585
R4505 gnd.n5250 gnd.n5249 585
R4506 gnd.n5234 gnd.n5158 585
R4507 gnd.n5236 gnd.n5235 585
R4508 gnd.n5232 gnd.n5165 585
R4509 gnd.n5231 gnd.n5230 585
R4510 gnd.n5215 gnd.n5167 585
R4511 gnd.n5217 gnd.n5216 585
R4512 gnd.n5213 gnd.n5174 585
R4513 gnd.n5212 gnd.n5211 585
R4514 gnd.n5200 gnd.n5176 585
R4515 gnd.n5202 gnd.n5201 585
R4516 gnd.n5198 gnd.n5177 585
R4517 gnd.n5197 gnd.n5196 585
R4518 gnd.n5189 gnd.n5179 585
R4519 gnd.n5191 gnd.n5190 585
R4520 gnd.n5187 gnd.n5181 585
R4521 gnd.n5186 gnd.n5185 585
R4522 gnd.n5183 gnd.n1585 585
R4523 gnd.n5295 gnd.n5294 585
R4524 gnd.n5292 gnd.n5127 585
R4525 gnd.n5291 gnd.n5128 585
R4526 gnd.n5289 gnd.n5288 585
R4527 gnd.n6484 gnd.n795 530.795
R4528 gnd.n5413 gnd.n1830 482.89
R4529 gnd.n5416 gnd.n5415 482.89
R4530 gnd.n2280 gnd.n2204 482.89
R4531 gnd.n6060 gnd.n1456 482.89
R4532 gnd.n2205 gnd.t79 443.966
R4533 gnd.n1824 gnd.t105 443.966
R4534 gnd.n5997 gnd.t131 443.966
R4535 gnd.n5347 gnd.t32 443.966
R4536 gnd.n1231 gnd.t72 371.625
R4537 gnd.n5140 gnd.t99 371.625
R4538 gnd.n1238 gnd.t121 371.625
R4539 gnd.n5553 gnd.t96 371.625
R4540 gnd.n5605 gnd.t86 371.625
R4541 gnd.n1755 gnd.t25 371.625
R4542 gnd.n174 gnd.t36 371.625
R4543 gnd.n196 gnd.t21 371.625
R4544 gnd.n218 gnd.t89 371.625
R4545 gnd.n7187 gnd.t114 371.625
R4546 gnd.n3967 gnd.t56 371.625
R4547 gnd.n3989 gnd.t42 371.625
R4548 gnd.n4012 gnd.t66 371.625
R4549 gnd.n4031 gnd.t17 371.625
R4550 gnd.n1308 gnd.t111 371.625
R4551 gnd.n1349 gnd.t45 371.625
R4552 gnd.n1328 gnd.t69 371.625
R4553 gnd.n5130 gnd.t49 371.625
R4554 gnd.n2931 gnd.t59 323.425
R4555 gnd.n2489 gnd.t92 323.425
R4556 gnd.n3779 gnd.n3753 289.615
R4557 gnd.n3747 gnd.n3721 289.615
R4558 gnd.n3715 gnd.n3689 289.615
R4559 gnd.n3684 gnd.n3658 289.615
R4560 gnd.n3652 gnd.n3626 289.615
R4561 gnd.n3620 gnd.n3594 289.615
R4562 gnd.n3588 gnd.n3562 289.615
R4563 gnd.n3557 gnd.n3531 289.615
R4564 gnd.n3005 gnd.t124 279.217
R4565 gnd.n2515 gnd.t117 279.217
R4566 gnd.n1463 gnd.t110 260.649
R4567 gnd.n5339 gnd.t31 260.649
R4568 gnd.n6062 gnd.n6061 256.663
R4569 gnd.n6062 gnd.n1422 256.663
R4570 gnd.n6062 gnd.n1423 256.663
R4571 gnd.n6062 gnd.n1424 256.663
R4572 gnd.n6062 gnd.n1425 256.663
R4573 gnd.n6062 gnd.n1426 256.663
R4574 gnd.n6062 gnd.n1427 256.663
R4575 gnd.n6062 gnd.n1428 256.663
R4576 gnd.n6062 gnd.n1429 256.663
R4577 gnd.n6062 gnd.n1430 256.663
R4578 gnd.n6062 gnd.n1431 256.663
R4579 gnd.n6062 gnd.n1432 256.663
R4580 gnd.n6062 gnd.n1433 256.663
R4581 gnd.n6062 gnd.n1434 256.663
R4582 gnd.n6062 gnd.n1435 256.663
R4583 gnd.n6062 gnd.n1436 256.663
R4584 gnd.n6065 gnd.n1419 256.663
R4585 gnd.n6063 gnd.n6062 256.663
R4586 gnd.n6062 gnd.n1437 256.663
R4587 gnd.n6062 gnd.n1438 256.663
R4588 gnd.n6062 gnd.n1439 256.663
R4589 gnd.n6062 gnd.n1440 256.663
R4590 gnd.n6062 gnd.n1441 256.663
R4591 gnd.n6062 gnd.n1442 256.663
R4592 gnd.n6062 gnd.n1443 256.663
R4593 gnd.n6062 gnd.n1444 256.663
R4594 gnd.n6062 gnd.n1445 256.663
R4595 gnd.n6062 gnd.n1446 256.663
R4596 gnd.n6062 gnd.n1447 256.663
R4597 gnd.n6062 gnd.n1448 256.663
R4598 gnd.n6062 gnd.n1449 256.663
R4599 gnd.n6062 gnd.n1450 256.663
R4600 gnd.n6062 gnd.n1451 256.663
R4601 gnd.n6062 gnd.n1452 256.663
R4602 gnd.n5481 gnd.n1808 256.663
R4603 gnd.n5481 gnd.n1809 256.663
R4604 gnd.n5481 gnd.n1810 256.663
R4605 gnd.n5481 gnd.n1811 256.663
R4606 gnd.n5481 gnd.n1812 256.663
R4607 gnd.n5481 gnd.n1813 256.663
R4608 gnd.n5481 gnd.n1814 256.663
R4609 gnd.n5481 gnd.n1815 256.663
R4610 gnd.n5481 gnd.n1816 256.663
R4611 gnd.n5481 gnd.n1817 256.663
R4612 gnd.n5481 gnd.n1818 256.663
R4613 gnd.n5481 gnd.n1819 256.663
R4614 gnd.n5481 gnd.n1820 256.663
R4615 gnd.n5481 gnd.n1821 256.663
R4616 gnd.n5481 gnd.n1822 256.663
R4617 gnd.n5481 gnd.n5478 256.663
R4618 gnd.n5484 gnd.n1789 256.663
R4619 gnd.n5482 gnd.n5481 256.663
R4620 gnd.n5481 gnd.n1807 256.663
R4621 gnd.n5481 gnd.n1806 256.663
R4622 gnd.n5481 gnd.n1805 256.663
R4623 gnd.n5481 gnd.n1804 256.663
R4624 gnd.n5481 gnd.n1803 256.663
R4625 gnd.n5481 gnd.n1802 256.663
R4626 gnd.n5481 gnd.n1801 256.663
R4627 gnd.n5481 gnd.n1800 256.663
R4628 gnd.n5481 gnd.n1799 256.663
R4629 gnd.n5481 gnd.n1798 256.663
R4630 gnd.n5481 gnd.n1797 256.663
R4631 gnd.n5481 gnd.n1796 256.663
R4632 gnd.n5481 gnd.n1795 256.663
R4633 gnd.n5481 gnd.n1794 256.663
R4634 gnd.n5481 gnd.n1793 256.663
R4635 gnd.n5481 gnd.n1792 256.663
R4636 gnd.n4211 gnd.n3940 242.672
R4637 gnd.n4211 gnd.n3941 242.672
R4638 gnd.n4211 gnd.n3942 242.672
R4639 gnd.n4211 gnd.n3943 242.672
R4640 gnd.n4211 gnd.n3944 242.672
R4641 gnd.n4211 gnd.n3945 242.672
R4642 gnd.n4211 gnd.n3946 242.672
R4643 gnd.n4211 gnd.n3947 242.672
R4644 gnd.n4211 gnd.n3948 242.672
R4645 gnd.n6117 gnd.n6116 242.672
R4646 gnd.n6116 gnd.n1256 242.672
R4647 gnd.n6116 gnd.n1254 242.672
R4648 gnd.n6116 gnd.n1253 242.672
R4649 gnd.n6116 gnd.n1251 242.672
R4650 gnd.n6116 gnd.n1249 242.672
R4651 gnd.n6116 gnd.n1248 242.672
R4652 gnd.n6116 gnd.n1246 242.672
R4653 gnd.n6116 gnd.n1244 242.672
R4654 gnd.n3059 gnd.n3058 242.672
R4655 gnd.n3059 gnd.n2969 242.672
R4656 gnd.n3059 gnd.n2970 242.672
R4657 gnd.n3059 gnd.n2971 242.672
R4658 gnd.n3059 gnd.n2972 242.672
R4659 gnd.n3059 gnd.n2973 242.672
R4660 gnd.n3059 gnd.n2974 242.672
R4661 gnd.n3059 gnd.n2975 242.672
R4662 gnd.n3059 gnd.n2976 242.672
R4663 gnd.n3059 gnd.n2977 242.672
R4664 gnd.n3059 gnd.n2978 242.672
R4665 gnd.n3059 gnd.n2979 242.672
R4666 gnd.n3060 gnd.n3059 242.672
R4667 gnd.n3911 gnd.n2464 242.672
R4668 gnd.n3911 gnd.n2463 242.672
R4669 gnd.n3911 gnd.n2462 242.672
R4670 gnd.n3911 gnd.n2461 242.672
R4671 gnd.n3911 gnd.n2460 242.672
R4672 gnd.n3911 gnd.n2459 242.672
R4673 gnd.n3911 gnd.n2458 242.672
R4674 gnd.n3911 gnd.n2457 242.672
R4675 gnd.n3911 gnd.n2456 242.672
R4676 gnd.n3911 gnd.n2455 242.672
R4677 gnd.n3911 gnd.n2454 242.672
R4678 gnd.n3911 gnd.n2453 242.672
R4679 gnd.n3911 gnd.n2452 242.672
R4680 gnd.n5205 gnd.n1598 242.672
R4681 gnd.n5222 gnd.n1598 242.672
R4682 gnd.n5224 gnd.n1598 242.672
R4683 gnd.n5241 gnd.n1598 242.672
R4684 gnd.n5243 gnd.n1598 242.672
R4685 gnd.n5260 gnd.n1598 242.672
R4686 gnd.n5262 gnd.n1598 242.672
R4687 gnd.n5280 gnd.n1598 242.672
R4688 gnd.n5282 gnd.n1598 242.672
R4689 gnd.n7249 gnd.n170 242.672
R4690 gnd.n7190 gnd.n170 242.672
R4691 gnd.n7239 gnd.n170 242.672
R4692 gnd.n7194 gnd.n170 242.672
R4693 gnd.n7229 gnd.n170 242.672
R4694 gnd.n7198 gnd.n170 242.672
R4695 gnd.n7219 gnd.n170 242.672
R4696 gnd.n7202 gnd.n170 242.672
R4697 gnd.n7209 gnd.n170 242.672
R4698 gnd.n3143 gnd.n3142 242.672
R4699 gnd.n3142 gnd.n2881 242.672
R4700 gnd.n3142 gnd.n2882 242.672
R4701 gnd.n3142 gnd.n2883 242.672
R4702 gnd.n3142 gnd.n2884 242.672
R4703 gnd.n3142 gnd.n2885 242.672
R4704 gnd.n3142 gnd.n2886 242.672
R4705 gnd.n3142 gnd.n2887 242.672
R4706 gnd.n3911 gnd.n2465 242.672
R4707 gnd.n3911 gnd.n2466 242.672
R4708 gnd.n3911 gnd.n2467 242.672
R4709 gnd.n3911 gnd.n2468 242.672
R4710 gnd.n3911 gnd.n2469 242.672
R4711 gnd.n3911 gnd.n2470 242.672
R4712 gnd.n3911 gnd.n2471 242.672
R4713 gnd.n3911 gnd.n2472 242.672
R4714 gnd.n4212 gnd.n4211 242.672
R4715 gnd.n4211 gnd.n3912 242.672
R4716 gnd.n4211 gnd.n3913 242.672
R4717 gnd.n4211 gnd.n3914 242.672
R4718 gnd.n4211 gnd.n3915 242.672
R4719 gnd.n4211 gnd.n3916 242.672
R4720 gnd.n4211 gnd.n3917 242.672
R4721 gnd.n4211 gnd.n3918 242.672
R4722 gnd.n4211 gnd.n3919 242.672
R4723 gnd.n4211 gnd.n3920 242.672
R4724 gnd.n4211 gnd.n3921 242.672
R4725 gnd.n4211 gnd.n3922 242.672
R4726 gnd.n4211 gnd.n3923 242.672
R4727 gnd.n4211 gnd.n3924 242.672
R4728 gnd.n4211 gnd.n3925 242.672
R4729 gnd.n4211 gnd.n3926 242.672
R4730 gnd.n4211 gnd.n3927 242.672
R4731 gnd.n4211 gnd.n3928 242.672
R4732 gnd.n4211 gnd.n3929 242.672
R4733 gnd.n4211 gnd.n3930 242.672
R4734 gnd.n4211 gnd.n3931 242.672
R4735 gnd.n4211 gnd.n3932 242.672
R4736 gnd.n4211 gnd.n3933 242.672
R4737 gnd.n4211 gnd.n3934 242.672
R4738 gnd.n4211 gnd.n3935 242.672
R4739 gnd.n4211 gnd.n3936 242.672
R4740 gnd.n4211 gnd.n3937 242.672
R4741 gnd.n4211 gnd.n3938 242.672
R4742 gnd.n4211 gnd.n3939 242.672
R4743 gnd.n6116 gnd.n1258 242.672
R4744 gnd.n6116 gnd.n1259 242.672
R4745 gnd.n6116 gnd.n1260 242.672
R4746 gnd.n6116 gnd.n1261 242.672
R4747 gnd.n6116 gnd.n1262 242.672
R4748 gnd.n6116 gnd.n1263 242.672
R4749 gnd.n6116 gnd.n1264 242.672
R4750 gnd.n6116 gnd.n1265 242.672
R4751 gnd.n6116 gnd.n1266 242.672
R4752 gnd.n6116 gnd.n1267 242.672
R4753 gnd.n6116 gnd.n1268 242.672
R4754 gnd.n6116 gnd.n1269 242.672
R4755 gnd.n6116 gnd.n1270 242.672
R4756 gnd.n6116 gnd.n1271 242.672
R4757 gnd.n6116 gnd.n1272 242.672
R4758 gnd.n6116 gnd.n1273 242.672
R4759 gnd.n6066 gnd.n1319 242.672
R4760 gnd.n6116 gnd.n1274 242.672
R4761 gnd.n6116 gnd.n1275 242.672
R4762 gnd.n6116 gnd.n1276 242.672
R4763 gnd.n6116 gnd.n1277 242.672
R4764 gnd.n6116 gnd.n1278 242.672
R4765 gnd.n6116 gnd.n1279 242.672
R4766 gnd.n6116 gnd.n1280 242.672
R4767 gnd.n6116 gnd.n1281 242.672
R4768 gnd.n6116 gnd.n1282 242.672
R4769 gnd.n6116 gnd.n1283 242.672
R4770 gnd.n6116 gnd.n1284 242.672
R4771 gnd.n6116 gnd.n1285 242.672
R4772 gnd.n6116 gnd.n6115 242.672
R4773 gnd.n5514 gnd.n1598 242.672
R4774 gnd.n5517 gnd.n1598 242.672
R4775 gnd.n5525 gnd.n1598 242.672
R4776 gnd.n5527 gnd.n1598 242.672
R4777 gnd.n5535 gnd.n1598 242.672
R4778 gnd.n5537 gnd.n1598 242.672
R4779 gnd.n5545 gnd.n1598 242.672
R4780 gnd.n5547 gnd.n1598 242.672
R4781 gnd.n5558 gnd.n1598 242.672
R4782 gnd.n5560 gnd.n1598 242.672
R4783 gnd.n5568 gnd.n1598 242.672
R4784 gnd.n5570 gnd.n1598 242.672
R4785 gnd.n5579 gnd.n1598 242.672
R4786 gnd.n5580 gnd.n5485 242.672
R4787 gnd.n5581 gnd.n1598 242.672
R4788 gnd.n5583 gnd.n1598 242.672
R4789 gnd.n5591 gnd.n1598 242.672
R4790 gnd.n5593 gnd.n1598 242.672
R4791 gnd.n5601 gnd.n1598 242.672
R4792 gnd.n5603 gnd.n1598 242.672
R4793 gnd.n5613 gnd.n1598 242.672
R4794 gnd.n5615 gnd.n1598 242.672
R4795 gnd.n5623 gnd.n1598 242.672
R4796 gnd.n5625 gnd.n1598 242.672
R4797 gnd.n5633 gnd.n1598 242.672
R4798 gnd.n5635 gnd.n1598 242.672
R4799 gnd.n5643 gnd.n1598 242.672
R4800 gnd.n5645 gnd.n1598 242.672
R4801 gnd.n5654 gnd.n1598 242.672
R4802 gnd.n5657 gnd.n1598 242.672
R4803 gnd.n381 gnd.n170 242.672
R4804 gnd.n177 gnd.n170 242.672
R4805 gnd.n371 gnd.n170 242.672
R4806 gnd.n181 gnd.n170 242.672
R4807 gnd.n361 gnd.n170 242.672
R4808 gnd.n185 gnd.n170 242.672
R4809 gnd.n351 gnd.n170 242.672
R4810 gnd.n189 gnd.n170 242.672
R4811 gnd.n341 gnd.n170 242.672
R4812 gnd.n193 gnd.n170 242.672
R4813 gnd.n331 gnd.n170 242.672
R4814 gnd.n199 gnd.n170 242.672
R4815 gnd.n321 gnd.n170 242.672
R4816 gnd.n203 gnd.n170 242.672
R4817 gnd.n311 gnd.n170 242.672
R4818 gnd.n207 gnd.n170 242.672
R4819 gnd.n301 gnd.n170 242.672
R4820 gnd.n211 gnd.n170 242.672
R4821 gnd.n291 gnd.n170 242.672
R4822 gnd.n215 gnd.n170 242.672
R4823 gnd.n281 gnd.n170 242.672
R4824 gnd.n271 gnd.n170 242.672
R4825 gnd.n270 gnd.n170 242.672
R4826 gnd.n225 gnd.n170 242.672
R4827 gnd.n260 gnd.n170 242.672
R4828 gnd.n229 gnd.n170 242.672
R4829 gnd.n250 gnd.n170 242.672
R4830 gnd.n233 gnd.n170 242.672
R4831 gnd.n240 gnd.n170 242.672
R4832 gnd.n6181 gnd.n6180 242.672
R4833 gnd.n6181 gnd.n1155 242.672
R4834 gnd.n6181 gnd.n1156 242.672
R4835 gnd.n6181 gnd.n1157 242.672
R4836 gnd.n6181 gnd.n1158 242.672
R4837 gnd.n6181 gnd.n1159 242.672
R4838 gnd.n6181 gnd.n1160 242.672
R4839 gnd.n6181 gnd.n1161 242.672
R4840 gnd.n6181 gnd.n1162 242.672
R4841 gnd.n6181 gnd.n1163 242.672
R4842 gnd.n6181 gnd.n1164 242.672
R4843 gnd.n6181 gnd.n1165 242.672
R4844 gnd.n6181 gnd.n1167 242.672
R4845 gnd.n6182 gnd.n6181 242.672
R4846 gnd.n5271 gnd.n1597 242.672
R4847 gnd.n5148 gnd.n1597 242.672
R4848 gnd.n5252 gnd.n1597 242.672
R4849 gnd.n5157 gnd.n1597 242.672
R4850 gnd.n5233 gnd.n1597 242.672
R4851 gnd.n5166 gnd.n1597 242.672
R4852 gnd.n5214 gnd.n1597 242.672
R4853 gnd.n5175 gnd.n1597 242.672
R4854 gnd.n5199 gnd.n1597 242.672
R4855 gnd.n5178 gnd.n1597 242.672
R4856 gnd.n5188 gnd.n1597 242.672
R4857 gnd.n5182 gnd.n1597 242.672
R4858 gnd.n5293 gnd.n1597 242.672
R4859 gnd.n5290 gnd.n1597 242.672
R4860 gnd.n239 gnd.n166 240.244
R4861 gnd.n242 gnd.n241 240.244
R4862 gnd.n249 gnd.n248 240.244
R4863 gnd.n252 gnd.n251 240.244
R4864 gnd.n259 gnd.n258 240.244
R4865 gnd.n262 gnd.n261 240.244
R4866 gnd.n269 gnd.n268 240.244
R4867 gnd.n273 gnd.n272 240.244
R4868 gnd.n280 gnd.n221 240.244
R4869 gnd.n283 gnd.n282 240.244
R4870 gnd.n290 gnd.n289 240.244
R4871 gnd.n293 gnd.n292 240.244
R4872 gnd.n300 gnd.n299 240.244
R4873 gnd.n303 gnd.n302 240.244
R4874 gnd.n310 gnd.n309 240.244
R4875 gnd.n313 gnd.n312 240.244
R4876 gnd.n320 gnd.n319 240.244
R4877 gnd.n323 gnd.n322 240.244
R4878 gnd.n330 gnd.n329 240.244
R4879 gnd.n333 gnd.n332 240.244
R4880 gnd.n340 gnd.n339 240.244
R4881 gnd.n343 gnd.n342 240.244
R4882 gnd.n350 gnd.n349 240.244
R4883 gnd.n353 gnd.n352 240.244
R4884 gnd.n360 gnd.n359 240.244
R4885 gnd.n363 gnd.n362 240.244
R4886 gnd.n370 gnd.n369 240.244
R4887 gnd.n373 gnd.n372 240.244
R4888 gnd.n380 gnd.n379 240.244
R4889 gnd.n1752 gnd.n1607 240.244
R4890 gnd.n1752 gnd.n1619 240.244
R4891 gnd.n5668 gnd.n1619 240.244
R4892 gnd.n5668 gnd.n1631 240.244
R4893 gnd.n5678 gnd.n1631 240.244
R4894 gnd.n5678 gnd.n1642 240.244
R4895 gnd.n1741 gnd.n1642 240.244
R4896 gnd.n1741 gnd.n1651 240.244
R4897 gnd.n5685 gnd.n1651 240.244
R4898 gnd.n5685 gnd.n1662 240.244
R4899 gnd.n5743 gnd.n1662 240.244
R4900 gnd.n5743 gnd.n1671 240.244
R4901 gnd.n5748 gnd.n1671 240.244
R4902 gnd.n5748 gnd.n1682 240.244
R4903 gnd.n5768 gnd.n1682 240.244
R4904 gnd.n5768 gnd.n1691 240.244
R4905 gnd.n1697 gnd.n1691 240.244
R4906 gnd.n5773 gnd.n1697 240.244
R4907 gnd.n5773 gnd.n5772 240.244
R4908 gnd.n5772 gnd.n1707 240.244
R4909 gnd.n1714 gnd.n1707 240.244
R4910 gnd.n5786 gnd.n1714 240.244
R4911 gnd.n5786 gnd.n70 240.244
R4912 gnd.n398 gnd.n70 240.244
R4913 gnd.n7143 gnd.n398 240.244
R4914 gnd.n7143 gnd.n87 240.244
R4915 gnd.n7153 gnd.n87 240.244
R4916 gnd.n7153 gnd.n99 240.244
R4917 gnd.n7158 gnd.n99 240.244
R4918 gnd.n7158 gnd.n109 240.244
R4919 gnd.n7168 gnd.n109 240.244
R4920 gnd.n7168 gnd.n118 240.244
R4921 gnd.n7173 gnd.n118 240.244
R4922 gnd.n7173 gnd.n129 240.244
R4923 gnd.n7267 gnd.n129 240.244
R4924 gnd.n7267 gnd.n139 240.244
R4925 gnd.n7271 gnd.n139 240.244
R4926 gnd.n7271 gnd.n150 240.244
R4927 gnd.n7274 gnd.n150 240.244
R4928 gnd.n7274 gnd.n159 240.244
R4929 gnd.n7277 gnd.n159 240.244
R4930 gnd.n7277 gnd.n168 240.244
R4931 gnd.n5516 gnd.n5515 240.244
R4932 gnd.n5518 gnd.n5516 240.244
R4933 gnd.n5524 gnd.n5506 240.244
R4934 gnd.n5528 gnd.n5526 240.244
R4935 gnd.n5534 gnd.n5502 240.244
R4936 gnd.n5538 gnd.n5536 240.244
R4937 gnd.n5544 gnd.n5498 240.244
R4938 gnd.n5548 gnd.n5546 240.244
R4939 gnd.n5557 gnd.n5494 240.244
R4940 gnd.n5561 gnd.n5559 240.244
R4941 gnd.n5567 gnd.n5490 240.244
R4942 gnd.n5571 gnd.n5569 240.244
R4943 gnd.n5578 gnd.n5486 240.244
R4944 gnd.n5584 gnd.n5582 240.244
R4945 gnd.n5590 gnd.n1783 240.244
R4946 gnd.n5594 gnd.n5592 240.244
R4947 gnd.n5600 gnd.n1779 240.244
R4948 gnd.n5604 gnd.n5602 240.244
R4949 gnd.n5612 gnd.n1775 240.244
R4950 gnd.n5616 gnd.n5614 240.244
R4951 gnd.n5622 gnd.n1771 240.244
R4952 gnd.n5626 gnd.n5624 240.244
R4953 gnd.n5632 gnd.n1767 240.244
R4954 gnd.n5636 gnd.n5634 240.244
R4955 gnd.n5642 gnd.n1763 240.244
R4956 gnd.n5646 gnd.n5644 240.244
R4957 gnd.n5653 gnd.n1759 240.244
R4958 gnd.n5656 gnd.n5655 240.244
R4959 gnd.n5857 gnd.n1612 240.244
R4960 gnd.n5853 gnd.n1612 240.244
R4961 gnd.n5853 gnd.n1617 240.244
R4962 gnd.n5845 gnd.n1617 240.244
R4963 gnd.n5845 gnd.n1634 240.244
R4964 gnd.n5841 gnd.n1634 240.244
R4965 gnd.n5841 gnd.n1640 240.244
R4966 gnd.n5833 gnd.n1640 240.244
R4967 gnd.n5833 gnd.n1654 240.244
R4968 gnd.n5829 gnd.n1654 240.244
R4969 gnd.n5829 gnd.n1660 240.244
R4970 gnd.n5821 gnd.n1660 240.244
R4971 gnd.n5821 gnd.n1674 240.244
R4972 gnd.n5817 gnd.n1674 240.244
R4973 gnd.n5817 gnd.n1680 240.244
R4974 gnd.n5809 gnd.n1680 240.244
R4975 gnd.n5809 gnd.n5807 240.244
R4976 gnd.n5807 gnd.n1694 240.244
R4977 gnd.n1711 gnd.n1694 240.244
R4978 gnd.n5796 gnd.n1711 240.244
R4979 gnd.n5796 gnd.n5793 240.244
R4980 gnd.n5793 gnd.n73 240.244
R4981 gnd.n7338 gnd.n73 240.244
R4982 gnd.n7338 gnd.n74 240.244
R4983 gnd.n84 gnd.n74 240.244
R4984 gnd.n7332 gnd.n84 240.244
R4985 gnd.n7332 gnd.n85 240.244
R4986 gnd.n7324 gnd.n85 240.244
R4987 gnd.n7324 gnd.n102 240.244
R4988 gnd.n7320 gnd.n102 240.244
R4989 gnd.n7320 gnd.n107 240.244
R4990 gnd.n7312 gnd.n107 240.244
R4991 gnd.n7312 gnd.n121 240.244
R4992 gnd.n7308 gnd.n121 240.244
R4993 gnd.n7308 gnd.n127 240.244
R4994 gnd.n7300 gnd.n127 240.244
R4995 gnd.n7300 gnd.n142 240.244
R4996 gnd.n7296 gnd.n142 240.244
R4997 gnd.n7296 gnd.n148 240.244
R4998 gnd.n7288 gnd.n148 240.244
R4999 gnd.n7288 gnd.n161 240.244
R5000 gnd.n7284 gnd.n161 240.244
R5001 gnd.n1286 gnd.n1137 240.244
R5002 gnd.n6114 gnd.n1287 240.244
R5003 gnd.n6110 gnd.n6109 240.244
R5004 gnd.n6106 gnd.n6105 240.244
R5005 gnd.n6102 gnd.n6101 240.244
R5006 gnd.n6098 gnd.n6097 240.244
R5007 gnd.n6094 gnd.n6093 240.244
R5008 gnd.n6090 gnd.n6089 240.244
R5009 gnd.n6086 gnd.n6085 240.244
R5010 gnd.n6081 gnd.n6080 240.244
R5011 gnd.n6077 gnd.n6076 240.244
R5012 gnd.n6073 gnd.n6072 240.244
R5013 gnd.n6069 gnd.n6068 240.244
R5014 gnd.n1412 gnd.n1411 240.244
R5015 gnd.n1409 gnd.n1408 240.244
R5016 gnd.n1405 gnd.n1404 240.244
R5017 gnd.n1401 gnd.n1400 240.244
R5018 gnd.n1397 gnd.n1396 240.244
R5019 gnd.n1390 gnd.n1389 240.244
R5020 gnd.n1387 gnd.n1386 240.244
R5021 gnd.n1383 gnd.n1382 240.244
R5022 gnd.n1379 gnd.n1378 240.244
R5023 gnd.n1375 gnd.n1374 240.244
R5024 gnd.n1371 gnd.n1370 240.244
R5025 gnd.n1367 gnd.n1366 240.244
R5026 gnd.n1363 gnd.n1362 240.244
R5027 gnd.n1359 gnd.n1358 240.244
R5028 gnd.n1355 gnd.n1354 240.244
R5029 gnd.n4221 gnd.n2441 240.244
R5030 gnd.n4222 gnd.n4221 240.244
R5031 gnd.n4222 gnd.n2432 240.244
R5032 gnd.n4228 gnd.n2432 240.244
R5033 gnd.n4228 gnd.n2424 240.244
R5034 gnd.n4225 gnd.n2424 240.244
R5035 gnd.n4225 gnd.n968 240.244
R5036 gnd.n4251 gnd.n968 240.244
R5037 gnd.n4251 gnd.n981 240.244
R5038 gnd.n4261 gnd.n981 240.244
R5039 gnd.n4261 gnd.n992 240.244
R5040 gnd.n4266 gnd.n992 240.244
R5041 gnd.n4266 gnd.n1003 240.244
R5042 gnd.n4280 gnd.n1003 240.244
R5043 gnd.n4280 gnd.n1012 240.244
R5044 gnd.n4283 gnd.n1012 240.244
R5045 gnd.n4283 gnd.n2371 240.244
R5046 gnd.n2371 gnd.n1023 240.244
R5047 gnd.n2378 gnd.n1023 240.244
R5048 gnd.n2378 gnd.n1034 240.244
R5049 gnd.n4297 gnd.n1034 240.244
R5050 gnd.n4297 gnd.n1042 240.244
R5051 gnd.n2388 gnd.n1042 240.244
R5052 gnd.n2388 gnd.n1051 240.244
R5053 gnd.n4306 gnd.n1051 240.244
R5054 gnd.n4306 gnd.n1059 240.244
R5055 gnd.n2356 gnd.n1059 240.244
R5056 gnd.n2356 gnd.n1068 240.244
R5057 gnd.n4372 gnd.n1068 240.244
R5058 gnd.n4372 gnd.n1079 240.244
R5059 gnd.n4376 gnd.n1079 240.244
R5060 gnd.n4376 gnd.n1088 240.244
R5061 gnd.n4386 gnd.n1088 240.244
R5062 gnd.n4386 gnd.n1099 240.244
R5063 gnd.n2339 gnd.n1099 240.244
R5064 gnd.n2339 gnd.n1108 240.244
R5065 gnd.n4393 gnd.n1108 240.244
R5066 gnd.n4393 gnd.n1119 240.244
R5067 gnd.n4397 gnd.n1119 240.244
R5068 gnd.n4397 gnd.n1129 240.244
R5069 gnd.n6193 gnd.n1129 240.244
R5070 gnd.n6193 gnd.n1139 240.244
R5071 gnd.n4210 gnd.n2449 240.244
R5072 gnd.n4210 gnd.n3950 240.244
R5073 gnd.n4206 gnd.n4205 240.244
R5074 gnd.n4202 gnd.n4201 240.244
R5075 gnd.n4198 gnd.n4197 240.244
R5076 gnd.n4194 gnd.n4193 240.244
R5077 gnd.n4190 gnd.n4189 240.244
R5078 gnd.n4186 gnd.n4185 240.244
R5079 gnd.n4182 gnd.n4181 240.244
R5080 gnd.n4177 gnd.n4176 240.244
R5081 gnd.n4173 gnd.n4172 240.244
R5082 gnd.n4169 gnd.n4168 240.244
R5083 gnd.n4165 gnd.n4164 240.244
R5084 gnd.n4161 gnd.n4160 240.244
R5085 gnd.n4157 gnd.n4156 240.244
R5086 gnd.n4153 gnd.n4152 240.244
R5087 gnd.n4149 gnd.n4148 240.244
R5088 gnd.n4145 gnd.n4144 240.244
R5089 gnd.n4141 gnd.n4140 240.244
R5090 gnd.n4137 gnd.n4136 240.244
R5091 gnd.n4133 gnd.n4132 240.244
R5092 gnd.n4129 gnd.n4128 240.244
R5093 gnd.n4125 gnd.n4124 240.244
R5094 gnd.n4121 gnd.n4120 240.244
R5095 gnd.n4117 gnd.n4116 240.244
R5096 gnd.n4113 gnd.n4112 240.244
R5097 gnd.n4109 gnd.n4108 240.244
R5098 gnd.n4105 gnd.n4104 240.244
R5099 gnd.n4101 gnd.n4100 240.244
R5100 gnd.n4219 gnd.n2445 240.244
R5101 gnd.n4219 gnd.n2430 240.244
R5102 gnd.n4235 gnd.n2430 240.244
R5103 gnd.n4235 gnd.n2426 240.244
R5104 gnd.n4242 gnd.n2426 240.244
R5105 gnd.n4242 gnd.n972 240.244
R5106 gnd.n6304 gnd.n972 240.244
R5107 gnd.n6304 gnd.n973 240.244
R5108 gnd.n6300 gnd.n973 240.244
R5109 gnd.n6300 gnd.n979 240.244
R5110 gnd.n6292 gnd.n979 240.244
R5111 gnd.n6292 gnd.n995 240.244
R5112 gnd.n6288 gnd.n995 240.244
R5113 gnd.n6288 gnd.n1001 240.244
R5114 gnd.n6280 gnd.n1001 240.244
R5115 gnd.n6280 gnd.n1015 240.244
R5116 gnd.n1019 gnd.n1015 240.244
R5117 gnd.n6274 gnd.n1019 240.244
R5118 gnd.n6274 gnd.n1021 240.244
R5119 gnd.n6266 gnd.n1021 240.244
R5120 gnd.n6266 gnd.n1037 240.244
R5121 gnd.n6261 gnd.n1037 240.244
R5122 gnd.n6261 gnd.n1040 240.244
R5123 gnd.n6253 gnd.n1040 240.244
R5124 gnd.n6253 gnd.n1054 240.244
R5125 gnd.n6248 gnd.n1054 240.244
R5126 gnd.n6248 gnd.n1057 240.244
R5127 gnd.n6240 gnd.n1057 240.244
R5128 gnd.n6240 gnd.n1071 240.244
R5129 gnd.n6236 gnd.n1071 240.244
R5130 gnd.n6236 gnd.n1077 240.244
R5131 gnd.n6228 gnd.n1077 240.244
R5132 gnd.n6228 gnd.n1091 240.244
R5133 gnd.n6224 gnd.n1091 240.244
R5134 gnd.n6224 gnd.n1097 240.244
R5135 gnd.n6216 gnd.n1097 240.244
R5136 gnd.n6216 gnd.n1111 240.244
R5137 gnd.n6212 gnd.n1111 240.244
R5138 gnd.n6212 gnd.n1117 240.244
R5139 gnd.n6204 gnd.n1117 240.244
R5140 gnd.n6204 gnd.n1132 240.244
R5141 gnd.n6200 gnd.n1132 240.244
R5142 gnd.n3910 gnd.n2474 240.244
R5143 gnd.n3903 gnd.n3902 240.244
R5144 gnd.n3900 gnd.n3899 240.244
R5145 gnd.n3896 gnd.n3895 240.244
R5146 gnd.n3892 gnd.n3891 240.244
R5147 gnd.n3888 gnd.n3887 240.244
R5148 gnd.n3884 gnd.n3883 240.244
R5149 gnd.n3880 gnd.n3879 240.244
R5150 gnd.n3154 gnd.n2866 240.244
R5151 gnd.n3164 gnd.n2866 240.244
R5152 gnd.n3164 gnd.n2857 240.244
R5153 gnd.n2857 gnd.n2846 240.244
R5154 gnd.n3185 gnd.n2846 240.244
R5155 gnd.n3185 gnd.n2840 240.244
R5156 gnd.n3195 gnd.n2840 240.244
R5157 gnd.n3195 gnd.n2829 240.244
R5158 gnd.n2829 gnd.n2821 240.244
R5159 gnd.n3213 gnd.n2821 240.244
R5160 gnd.n3214 gnd.n3213 240.244
R5161 gnd.n3214 gnd.n2806 240.244
R5162 gnd.n3216 gnd.n2806 240.244
R5163 gnd.n3216 gnd.n2792 240.244
R5164 gnd.n3258 gnd.n2792 240.244
R5165 gnd.n3259 gnd.n3258 240.244
R5166 gnd.n3262 gnd.n3259 240.244
R5167 gnd.n3262 gnd.n2747 240.244
R5168 gnd.n2787 gnd.n2747 240.244
R5169 gnd.n2787 gnd.n2757 240.244
R5170 gnd.n3272 gnd.n2757 240.244
R5171 gnd.n3272 gnd.n2778 240.244
R5172 gnd.n3282 gnd.n2778 240.244
R5173 gnd.n3282 gnd.n2676 240.244
R5174 gnd.n3327 gnd.n2676 240.244
R5175 gnd.n3327 gnd.n2662 240.244
R5176 gnd.n3349 gnd.n2662 240.244
R5177 gnd.n3350 gnd.n3349 240.244
R5178 gnd.n3350 gnd.n2649 240.244
R5179 gnd.n2649 gnd.n2638 240.244
R5180 gnd.n3381 gnd.n2638 240.244
R5181 gnd.n3382 gnd.n3381 240.244
R5182 gnd.n3383 gnd.n3382 240.244
R5183 gnd.n3383 gnd.n2623 240.244
R5184 gnd.n2623 gnd.n2622 240.244
R5185 gnd.n2622 gnd.n2607 240.244
R5186 gnd.n3434 gnd.n2607 240.244
R5187 gnd.n3435 gnd.n3434 240.244
R5188 gnd.n3435 gnd.n2594 240.244
R5189 gnd.n2594 gnd.n2583 240.244
R5190 gnd.n3466 gnd.n2583 240.244
R5191 gnd.n3467 gnd.n3466 240.244
R5192 gnd.n3468 gnd.n3467 240.244
R5193 gnd.n3468 gnd.n2567 240.244
R5194 gnd.n2567 gnd.n2566 240.244
R5195 gnd.n2566 gnd.n2553 240.244
R5196 gnd.n3523 gnd.n2553 240.244
R5197 gnd.n3524 gnd.n3523 240.244
R5198 gnd.n3524 gnd.n2540 240.244
R5199 gnd.n2540 gnd.n2530 240.244
R5200 gnd.n3811 gnd.n2530 240.244
R5201 gnd.n3814 gnd.n3811 240.244
R5202 gnd.n3814 gnd.n3813 240.244
R5203 gnd.n3144 gnd.n2879 240.244
R5204 gnd.n2900 gnd.n2879 240.244
R5205 gnd.n2903 gnd.n2902 240.244
R5206 gnd.n2910 gnd.n2909 240.244
R5207 gnd.n2913 gnd.n2912 240.244
R5208 gnd.n2920 gnd.n2919 240.244
R5209 gnd.n2923 gnd.n2922 240.244
R5210 gnd.n2930 gnd.n2929 240.244
R5211 gnd.n3152 gnd.n2876 240.244
R5212 gnd.n2876 gnd.n2855 240.244
R5213 gnd.n3175 gnd.n2855 240.244
R5214 gnd.n3175 gnd.n2849 240.244
R5215 gnd.n3183 gnd.n2849 240.244
R5216 gnd.n3183 gnd.n2851 240.244
R5217 gnd.n2851 gnd.n2827 240.244
R5218 gnd.n3205 gnd.n2827 240.244
R5219 gnd.n3205 gnd.n2823 240.244
R5220 gnd.n3211 gnd.n2823 240.244
R5221 gnd.n3211 gnd.n2805 240.244
R5222 gnd.n3236 gnd.n2805 240.244
R5223 gnd.n3236 gnd.n2800 240.244
R5224 gnd.n3248 gnd.n2800 240.244
R5225 gnd.n3248 gnd.n2801 240.244
R5226 gnd.n3244 gnd.n2801 240.244
R5227 gnd.n3244 gnd.n2749 240.244
R5228 gnd.n3296 gnd.n2749 240.244
R5229 gnd.n3296 gnd.n2750 240.244
R5230 gnd.n3292 gnd.n2750 240.244
R5231 gnd.n3292 gnd.n2756 240.244
R5232 gnd.n2776 gnd.n2756 240.244
R5233 gnd.n2776 gnd.n2674 240.244
R5234 gnd.n3331 gnd.n2674 240.244
R5235 gnd.n3331 gnd.n2669 240.244
R5236 gnd.n3339 gnd.n2669 240.244
R5237 gnd.n3339 gnd.n2670 240.244
R5238 gnd.n2670 gnd.n2647 240.244
R5239 gnd.n3371 gnd.n2647 240.244
R5240 gnd.n3371 gnd.n2642 240.244
R5241 gnd.n3379 gnd.n2642 240.244
R5242 gnd.n3379 gnd.n2643 240.244
R5243 gnd.n2643 gnd.n2620 240.244
R5244 gnd.n3416 gnd.n2620 240.244
R5245 gnd.n3416 gnd.n2615 240.244
R5246 gnd.n3424 gnd.n2615 240.244
R5247 gnd.n3424 gnd.n2616 240.244
R5248 gnd.n2616 gnd.n2592 240.244
R5249 gnd.n3456 gnd.n2592 240.244
R5250 gnd.n3456 gnd.n2587 240.244
R5251 gnd.n3464 gnd.n2587 240.244
R5252 gnd.n3464 gnd.n2588 240.244
R5253 gnd.n2588 gnd.n2565 240.244
R5254 gnd.n3505 gnd.n2565 240.244
R5255 gnd.n3505 gnd.n2560 240.244
R5256 gnd.n3513 gnd.n2560 240.244
R5257 gnd.n3513 gnd.n2561 240.244
R5258 gnd.n2561 gnd.n2538 240.244
R5259 gnd.n3799 gnd.n2538 240.244
R5260 gnd.n3799 gnd.n2533 240.244
R5261 gnd.n3809 gnd.n2533 240.244
R5262 gnd.n3809 gnd.n2534 240.244
R5263 gnd.n2534 gnd.n2473 240.244
R5264 gnd.n7208 gnd.n171 240.244
R5265 gnd.n7211 gnd.n7210 240.244
R5266 gnd.n7218 gnd.n7217 240.244
R5267 gnd.n7221 gnd.n7220 240.244
R5268 gnd.n7228 gnd.n7227 240.244
R5269 gnd.n7231 gnd.n7230 240.244
R5270 gnd.n7238 gnd.n7237 240.244
R5271 gnd.n7241 gnd.n7240 240.244
R5272 gnd.n7248 gnd.n7247 240.244
R5273 gnd.n5122 gnd.n1608 240.244
R5274 gnd.n5122 gnd.n1620 240.244
R5275 gnd.n5670 gnd.n1620 240.244
R5276 gnd.n5670 gnd.n1632 240.244
R5277 gnd.n5676 gnd.n1632 240.244
R5278 gnd.n5676 gnd.n1643 240.244
R5279 gnd.n5696 gnd.n1643 240.244
R5280 gnd.n5696 gnd.n1652 240.244
R5281 gnd.n5687 gnd.n1652 240.244
R5282 gnd.n5687 gnd.n1663 240.244
R5283 gnd.n1735 gnd.n1663 240.244
R5284 gnd.n1735 gnd.n1672 240.244
R5285 gnd.n5750 gnd.n1672 240.244
R5286 gnd.n5750 gnd.n1683 240.244
R5287 gnd.n5766 gnd.n1683 240.244
R5288 gnd.n5766 gnd.n1692 240.244
R5289 gnd.n1698 gnd.n1692 240.244
R5290 gnd.n5755 gnd.n1698 240.244
R5291 gnd.n5756 gnd.n5755 240.244
R5292 gnd.n5756 gnd.n1708 240.244
R5293 gnd.n1715 gnd.n1708 240.244
R5294 gnd.n1715 gnd.n66 240.244
R5295 gnd.n7340 gnd.n66 240.244
R5296 gnd.n7340 gnd.n68 240.244
R5297 gnd.n7145 gnd.n68 240.244
R5298 gnd.n7145 gnd.n88 240.244
R5299 gnd.n7151 gnd.n88 240.244
R5300 gnd.n7151 gnd.n100 240.244
R5301 gnd.n7160 gnd.n100 240.244
R5302 gnd.n7160 gnd.n110 240.244
R5303 gnd.n7166 gnd.n110 240.244
R5304 gnd.n7166 gnd.n119 240.244
R5305 gnd.n7175 gnd.n119 240.244
R5306 gnd.n7175 gnd.n130 240.244
R5307 gnd.n7265 gnd.n130 240.244
R5308 gnd.n7265 gnd.n140 240.244
R5309 gnd.n7261 gnd.n140 240.244
R5310 gnd.n7261 gnd.n151 240.244
R5311 gnd.n7258 gnd.n151 240.244
R5312 gnd.n7258 gnd.n160 240.244
R5313 gnd.n7255 gnd.n160 240.244
R5314 gnd.n7255 gnd.n169 240.244
R5315 gnd.n5221 gnd.n5170 240.244
R5316 gnd.n5225 gnd.n5223 240.244
R5317 gnd.n5240 gnd.n5161 240.244
R5318 gnd.n5244 gnd.n5242 240.244
R5319 gnd.n5259 gnd.n5152 240.244
R5320 gnd.n5263 gnd.n5261 240.244
R5321 gnd.n5279 gnd.n5143 240.244
R5322 gnd.n5283 gnd.n5281 240.244
R5323 gnd.n5139 gnd.n5138 240.244
R5324 gnd.n1622 gnd.n1610 240.244
R5325 gnd.n5851 gnd.n1622 240.244
R5326 gnd.n5851 gnd.n1623 240.244
R5327 gnd.n5847 gnd.n1623 240.244
R5328 gnd.n5847 gnd.n1629 240.244
R5329 gnd.n5839 gnd.n1629 240.244
R5330 gnd.n5839 gnd.n1644 240.244
R5331 gnd.n5835 gnd.n1644 240.244
R5332 gnd.n5835 gnd.n1649 240.244
R5333 gnd.n5827 gnd.n1649 240.244
R5334 gnd.n5827 gnd.n1665 240.244
R5335 gnd.n5823 gnd.n1665 240.244
R5336 gnd.n5823 gnd.n1670 240.244
R5337 gnd.n5815 gnd.n1670 240.244
R5338 gnd.n5815 gnd.n1684 240.244
R5339 gnd.n5811 gnd.n1684 240.244
R5340 gnd.n5811 gnd.n1689 240.244
R5341 gnd.n5777 gnd.n1689 240.244
R5342 gnd.n5778 gnd.n5777 240.244
R5343 gnd.n5778 gnd.n1710 240.244
R5344 gnd.n5791 gnd.n1710 240.244
R5345 gnd.n5791 gnd.n1723 240.244
R5346 gnd.n1723 gnd.n72 240.244
R5347 gnd.n7138 gnd.n72 240.244
R5348 gnd.n7138 gnd.n90 240.244
R5349 gnd.n7330 gnd.n90 240.244
R5350 gnd.n7330 gnd.n91 240.244
R5351 gnd.n7326 gnd.n91 240.244
R5352 gnd.n7326 gnd.n97 240.244
R5353 gnd.n7318 gnd.n97 240.244
R5354 gnd.n7318 gnd.n111 240.244
R5355 gnd.n7314 gnd.n111 240.244
R5356 gnd.n7314 gnd.n116 240.244
R5357 gnd.n7306 gnd.n116 240.244
R5358 gnd.n7306 gnd.n132 240.244
R5359 gnd.n7302 gnd.n132 240.244
R5360 gnd.n7302 gnd.n137 240.244
R5361 gnd.n7294 gnd.n137 240.244
R5362 gnd.n7294 gnd.n153 240.244
R5363 gnd.n7290 gnd.n153 240.244
R5364 gnd.n7290 gnd.n158 240.244
R5365 gnd.n7282 gnd.n158 240.244
R5366 gnd.n2493 gnd.n2451 240.244
R5367 gnd.n3870 gnd.n3869 240.244
R5368 gnd.n3866 gnd.n3865 240.244
R5369 gnd.n3862 gnd.n3861 240.244
R5370 gnd.n3858 gnd.n3857 240.244
R5371 gnd.n3854 gnd.n3853 240.244
R5372 gnd.n3850 gnd.n3849 240.244
R5373 gnd.n3846 gnd.n3845 240.244
R5374 gnd.n3842 gnd.n3841 240.244
R5375 gnd.n3838 gnd.n3837 240.244
R5376 gnd.n3834 gnd.n3833 240.244
R5377 gnd.n3830 gnd.n3829 240.244
R5378 gnd.n3826 gnd.n3825 240.244
R5379 gnd.n3067 gnd.n2964 240.244
R5380 gnd.n3067 gnd.n2957 240.244
R5381 gnd.n3078 gnd.n2957 240.244
R5382 gnd.n3078 gnd.n2953 240.244
R5383 gnd.n3084 gnd.n2953 240.244
R5384 gnd.n3084 gnd.n2945 240.244
R5385 gnd.n3094 gnd.n2945 240.244
R5386 gnd.n3094 gnd.n2940 240.244
R5387 gnd.n3130 gnd.n2940 240.244
R5388 gnd.n3130 gnd.n2941 240.244
R5389 gnd.n2941 gnd.n2888 240.244
R5390 gnd.n3125 gnd.n2888 240.244
R5391 gnd.n3125 gnd.n3124 240.244
R5392 gnd.n3124 gnd.n2867 240.244
R5393 gnd.n3120 gnd.n2867 240.244
R5394 gnd.n3120 gnd.n2858 240.244
R5395 gnd.n3117 gnd.n2858 240.244
R5396 gnd.n3117 gnd.n3116 240.244
R5397 gnd.n3116 gnd.n2841 240.244
R5398 gnd.n3112 gnd.n2841 240.244
R5399 gnd.n3112 gnd.n2830 240.244
R5400 gnd.n2830 gnd.n2811 240.244
R5401 gnd.n3225 gnd.n2811 240.244
R5402 gnd.n3225 gnd.n2807 240.244
R5403 gnd.n3233 gnd.n2807 240.244
R5404 gnd.n3233 gnd.n2798 240.244
R5405 gnd.n2798 gnd.n2734 240.244
R5406 gnd.n3305 gnd.n2734 240.244
R5407 gnd.n3305 gnd.n2735 240.244
R5408 gnd.n2746 gnd.n2735 240.244
R5409 gnd.n2781 gnd.n2746 240.244
R5410 gnd.n2784 gnd.n2781 240.244
R5411 gnd.n2784 gnd.n2758 240.244
R5412 gnd.n2771 gnd.n2758 240.244
R5413 gnd.n2771 gnd.n2768 240.244
R5414 gnd.n2768 gnd.n2677 240.244
R5415 gnd.n3326 gnd.n2677 240.244
R5416 gnd.n3326 gnd.n2667 240.244
R5417 gnd.n3322 gnd.n2667 240.244
R5418 gnd.n3322 gnd.n2661 240.244
R5419 gnd.n3319 gnd.n2661 240.244
R5420 gnd.n3319 gnd.n2650 240.244
R5421 gnd.n3316 gnd.n2650 240.244
R5422 gnd.n3316 gnd.n2628 240.244
R5423 gnd.n3392 gnd.n2628 240.244
R5424 gnd.n3392 gnd.n2624 240.244
R5425 gnd.n3413 gnd.n2624 240.244
R5426 gnd.n3413 gnd.n2613 240.244
R5427 gnd.n3409 gnd.n2613 240.244
R5428 gnd.n3409 gnd.n2606 240.244
R5429 gnd.n3406 gnd.n2606 240.244
R5430 gnd.n3406 gnd.n2595 240.244
R5431 gnd.n3403 gnd.n2595 240.244
R5432 gnd.n3403 gnd.n2572 240.244
R5433 gnd.n3477 gnd.n2572 240.244
R5434 gnd.n3477 gnd.n2568 240.244
R5435 gnd.n3502 gnd.n2568 240.244
R5436 gnd.n3502 gnd.n2559 240.244
R5437 gnd.n3498 gnd.n2559 240.244
R5438 gnd.n3498 gnd.n2552 240.244
R5439 gnd.n3494 gnd.n2552 240.244
R5440 gnd.n3494 gnd.n2541 240.244
R5441 gnd.n3491 gnd.n2541 240.244
R5442 gnd.n3491 gnd.n2522 240.244
R5443 gnd.n3821 gnd.n2522 240.244
R5444 gnd.n2981 gnd.n2980 240.244
R5445 gnd.n3052 gnd.n2980 240.244
R5446 gnd.n3050 gnd.n3049 240.244
R5447 gnd.n3046 gnd.n3045 240.244
R5448 gnd.n3042 gnd.n3041 240.244
R5449 gnd.n3038 gnd.n3037 240.244
R5450 gnd.n3034 gnd.n3033 240.244
R5451 gnd.n3030 gnd.n3029 240.244
R5452 gnd.n3026 gnd.n3025 240.244
R5453 gnd.n3022 gnd.n3021 240.244
R5454 gnd.n3018 gnd.n3017 240.244
R5455 gnd.n3014 gnd.n3013 240.244
R5456 gnd.n3010 gnd.n2968 240.244
R5457 gnd.n3070 gnd.n2962 240.244
R5458 gnd.n3070 gnd.n2958 240.244
R5459 gnd.n3076 gnd.n2958 240.244
R5460 gnd.n3076 gnd.n2951 240.244
R5461 gnd.n3086 gnd.n2951 240.244
R5462 gnd.n3086 gnd.n2947 240.244
R5463 gnd.n3092 gnd.n2947 240.244
R5464 gnd.n3092 gnd.n2938 240.244
R5465 gnd.n3132 gnd.n2938 240.244
R5466 gnd.n3132 gnd.n2889 240.244
R5467 gnd.n3140 gnd.n2889 240.244
R5468 gnd.n3140 gnd.n2890 240.244
R5469 gnd.n2890 gnd.n2868 240.244
R5470 gnd.n3161 gnd.n2868 240.244
R5471 gnd.n3161 gnd.n2860 240.244
R5472 gnd.n3172 gnd.n2860 240.244
R5473 gnd.n3172 gnd.n2861 240.244
R5474 gnd.n2861 gnd.n2842 240.244
R5475 gnd.n3192 gnd.n2842 240.244
R5476 gnd.n3192 gnd.n2832 240.244
R5477 gnd.n3202 gnd.n2832 240.244
R5478 gnd.n3202 gnd.n2813 240.244
R5479 gnd.n3223 gnd.n2813 240.244
R5480 gnd.n3223 gnd.n2815 240.244
R5481 gnd.n2815 gnd.n2796 240.244
R5482 gnd.n3251 gnd.n2796 240.244
R5483 gnd.n3251 gnd.n2738 240.244
R5484 gnd.n3303 gnd.n2738 240.244
R5485 gnd.n3303 gnd.n2739 240.244
R5486 gnd.n3299 gnd.n2739 240.244
R5487 gnd.n3299 gnd.n2745 240.244
R5488 gnd.n2760 gnd.n2745 240.244
R5489 gnd.n3289 gnd.n2760 240.244
R5490 gnd.n3289 gnd.n2761 240.244
R5491 gnd.n3285 gnd.n2761 240.244
R5492 gnd.n3285 gnd.n2767 240.244
R5493 gnd.n2767 gnd.n2666 240.244
R5494 gnd.n3342 gnd.n2666 240.244
R5495 gnd.n3342 gnd.n2659 240.244
R5496 gnd.n3353 gnd.n2659 240.244
R5497 gnd.n3353 gnd.n2652 240.244
R5498 gnd.n3368 gnd.n2652 240.244
R5499 gnd.n3368 gnd.n2653 240.244
R5500 gnd.n2653 gnd.n2631 240.244
R5501 gnd.n3390 gnd.n2631 240.244
R5502 gnd.n3390 gnd.n2632 240.244
R5503 gnd.n2632 gnd.n2611 240.244
R5504 gnd.n3427 gnd.n2611 240.244
R5505 gnd.n3427 gnd.n2604 240.244
R5506 gnd.n3438 gnd.n2604 240.244
R5507 gnd.n3438 gnd.n2597 240.244
R5508 gnd.n3453 gnd.n2597 240.244
R5509 gnd.n3453 gnd.n2598 240.244
R5510 gnd.n2598 gnd.n2575 240.244
R5511 gnd.n3475 gnd.n2575 240.244
R5512 gnd.n3475 gnd.n2577 240.244
R5513 gnd.n2577 gnd.n2557 240.244
R5514 gnd.n3516 gnd.n2557 240.244
R5515 gnd.n3516 gnd.n2550 240.244
R5516 gnd.n3527 gnd.n2550 240.244
R5517 gnd.n3527 gnd.n2543 240.244
R5518 gnd.n3796 gnd.n2543 240.244
R5519 gnd.n3796 gnd.n2544 240.244
R5520 gnd.n2544 gnd.n2525 240.244
R5521 gnd.n3819 gnd.n2525 240.244
R5522 gnd.n1188 gnd.n1142 240.244
R5523 gnd.n1245 gnd.n1189 240.244
R5524 gnd.n1199 gnd.n1198 240.244
R5525 gnd.n1247 gnd.n1206 240.244
R5526 gnd.n1250 gnd.n1207 240.244
R5527 gnd.n1217 gnd.n1216 240.244
R5528 gnd.n1252 gnd.n1224 240.244
R5529 gnd.n1255 gnd.n1225 240.244
R5530 gnd.n1242 gnd.n1237 240.244
R5531 gnd.n4049 gnd.n2443 240.244
R5532 gnd.n4046 gnd.n2443 240.244
R5533 gnd.n4046 gnd.n2433 240.244
R5534 gnd.n4043 gnd.n2433 240.244
R5535 gnd.n4043 gnd.n2425 240.244
R5536 gnd.n4040 gnd.n2425 240.244
R5537 gnd.n4040 gnd.n969 240.244
R5538 gnd.n4253 gnd.n969 240.244
R5539 gnd.n4253 gnd.n982 240.244
R5540 gnd.n4259 gnd.n982 240.244
R5541 gnd.n4259 gnd.n993 240.244
R5542 gnd.n4268 gnd.n993 240.244
R5543 gnd.n4268 gnd.n1004 240.244
R5544 gnd.n4277 gnd.n1004 240.244
R5545 gnd.n4277 gnd.n1013 240.244
R5546 gnd.n2372 gnd.n1013 240.244
R5547 gnd.n4331 gnd.n2372 240.244
R5548 gnd.n4331 gnd.n1024 240.244
R5549 gnd.n4327 gnd.n1024 240.244
R5550 gnd.n4327 gnd.n1035 240.244
R5551 gnd.n4295 gnd.n1035 240.244
R5552 gnd.n4295 gnd.n1043 240.244
R5553 gnd.n4314 gnd.n1043 240.244
R5554 gnd.n4314 gnd.n1052 240.244
R5555 gnd.n4308 gnd.n1052 240.244
R5556 gnd.n4308 gnd.n1060 240.244
R5557 gnd.n4364 gnd.n1060 240.244
R5558 gnd.n4364 gnd.n1069 240.244
R5559 gnd.n4370 gnd.n1069 240.244
R5560 gnd.n4370 gnd.n1080 240.244
R5561 gnd.n4378 gnd.n1080 240.244
R5562 gnd.n4378 gnd.n1089 240.244
R5563 gnd.n4384 gnd.n1089 240.244
R5564 gnd.n4384 gnd.n1100 240.244
R5565 gnd.n4408 gnd.n1100 240.244
R5566 gnd.n4408 gnd.n1109 240.244
R5567 gnd.n2344 gnd.n1109 240.244
R5568 gnd.n2344 gnd.n1120 240.244
R5569 gnd.n4399 gnd.n1120 240.244
R5570 gnd.n4399 gnd.n1130 240.244
R5571 gnd.n6191 gnd.n1130 240.244
R5572 gnd.n6191 gnd.n1140 240.244
R5573 gnd.n4086 gnd.n4085 240.244
R5574 gnd.n4082 gnd.n4081 240.244
R5575 gnd.n4078 gnd.n4077 240.244
R5576 gnd.n4074 gnd.n4073 240.244
R5577 gnd.n4070 gnd.n4069 240.244
R5578 gnd.n4066 gnd.n4065 240.244
R5579 gnd.n4062 gnd.n4061 240.244
R5580 gnd.n4058 gnd.n4057 240.244
R5581 gnd.n4030 gnd.n3949 240.244
R5582 gnd.n4090 gnd.n2444 240.244
R5583 gnd.n2444 gnd.n2435 240.244
R5584 gnd.n4233 gnd.n2435 240.244
R5585 gnd.n4233 gnd.n2422 240.244
R5586 gnd.n4244 gnd.n2422 240.244
R5587 gnd.n4245 gnd.n4244 240.244
R5588 gnd.n4245 gnd.n971 240.244
R5589 gnd.n983 gnd.n971 240.244
R5590 gnd.n6298 gnd.n983 240.244
R5591 gnd.n6298 gnd.n984 240.244
R5592 gnd.n6294 gnd.n984 240.244
R5593 gnd.n6294 gnd.n990 240.244
R5594 gnd.n6286 gnd.n990 240.244
R5595 gnd.n6286 gnd.n1006 240.244
R5596 gnd.n6282 gnd.n1006 240.244
R5597 gnd.n6282 gnd.n1011 240.244
R5598 gnd.n1026 gnd.n1011 240.244
R5599 gnd.n6272 gnd.n1026 240.244
R5600 gnd.n6272 gnd.n1027 240.244
R5601 gnd.n6268 gnd.n1027 240.244
R5602 gnd.n6268 gnd.n1033 240.244
R5603 gnd.n6259 gnd.n1033 240.244
R5604 gnd.n6259 gnd.n1044 240.244
R5605 gnd.n6255 gnd.n1044 240.244
R5606 gnd.n6255 gnd.n1049 240.244
R5607 gnd.n6246 gnd.n1049 240.244
R5608 gnd.n6246 gnd.n1062 240.244
R5609 gnd.n6242 gnd.n1062 240.244
R5610 gnd.n6242 gnd.n1067 240.244
R5611 gnd.n6234 gnd.n1067 240.244
R5612 gnd.n6234 gnd.n1081 240.244
R5613 gnd.n6230 gnd.n1081 240.244
R5614 gnd.n6230 gnd.n1086 240.244
R5615 gnd.n6222 gnd.n1086 240.244
R5616 gnd.n6222 gnd.n1102 240.244
R5617 gnd.n6218 gnd.n1102 240.244
R5618 gnd.n6218 gnd.n1107 240.244
R5619 gnd.n6210 gnd.n1107 240.244
R5620 gnd.n6210 gnd.n1122 240.244
R5621 gnd.n6206 gnd.n1122 240.244
R5622 gnd.n6206 gnd.n1127 240.244
R5623 gnd.n6198 gnd.n1127 240.244
R5624 gnd.n6483 gnd.n794 240.244
R5625 gnd.n6487 gnd.n794 240.244
R5626 gnd.n6487 gnd.n790 240.244
R5627 gnd.n6493 gnd.n790 240.244
R5628 gnd.n6493 gnd.n788 240.244
R5629 gnd.n6497 gnd.n788 240.244
R5630 gnd.n6497 gnd.n784 240.244
R5631 gnd.n6503 gnd.n784 240.244
R5632 gnd.n6503 gnd.n782 240.244
R5633 gnd.n6507 gnd.n782 240.244
R5634 gnd.n6507 gnd.n778 240.244
R5635 gnd.n6513 gnd.n778 240.244
R5636 gnd.n6513 gnd.n776 240.244
R5637 gnd.n6517 gnd.n776 240.244
R5638 gnd.n6517 gnd.n772 240.244
R5639 gnd.n6523 gnd.n772 240.244
R5640 gnd.n6523 gnd.n770 240.244
R5641 gnd.n6527 gnd.n770 240.244
R5642 gnd.n6527 gnd.n766 240.244
R5643 gnd.n6533 gnd.n766 240.244
R5644 gnd.n6533 gnd.n764 240.244
R5645 gnd.n6537 gnd.n764 240.244
R5646 gnd.n6537 gnd.n760 240.244
R5647 gnd.n6543 gnd.n760 240.244
R5648 gnd.n6543 gnd.n758 240.244
R5649 gnd.n6547 gnd.n758 240.244
R5650 gnd.n6547 gnd.n754 240.244
R5651 gnd.n6553 gnd.n754 240.244
R5652 gnd.n6553 gnd.n752 240.244
R5653 gnd.n6557 gnd.n752 240.244
R5654 gnd.n6557 gnd.n748 240.244
R5655 gnd.n6563 gnd.n748 240.244
R5656 gnd.n6563 gnd.n746 240.244
R5657 gnd.n6567 gnd.n746 240.244
R5658 gnd.n6567 gnd.n742 240.244
R5659 gnd.n6573 gnd.n742 240.244
R5660 gnd.n6573 gnd.n740 240.244
R5661 gnd.n6577 gnd.n740 240.244
R5662 gnd.n6577 gnd.n736 240.244
R5663 gnd.n6583 gnd.n736 240.244
R5664 gnd.n6583 gnd.n734 240.244
R5665 gnd.n6587 gnd.n734 240.244
R5666 gnd.n6587 gnd.n730 240.244
R5667 gnd.n6593 gnd.n730 240.244
R5668 gnd.n6593 gnd.n728 240.244
R5669 gnd.n6597 gnd.n728 240.244
R5670 gnd.n6597 gnd.n724 240.244
R5671 gnd.n6603 gnd.n724 240.244
R5672 gnd.n6603 gnd.n722 240.244
R5673 gnd.n6607 gnd.n722 240.244
R5674 gnd.n6607 gnd.n718 240.244
R5675 gnd.n6613 gnd.n718 240.244
R5676 gnd.n6613 gnd.n716 240.244
R5677 gnd.n6617 gnd.n716 240.244
R5678 gnd.n6617 gnd.n712 240.244
R5679 gnd.n6623 gnd.n712 240.244
R5680 gnd.n6623 gnd.n710 240.244
R5681 gnd.n6627 gnd.n710 240.244
R5682 gnd.n6627 gnd.n706 240.244
R5683 gnd.n6633 gnd.n706 240.244
R5684 gnd.n6633 gnd.n704 240.244
R5685 gnd.n6637 gnd.n704 240.244
R5686 gnd.n6637 gnd.n700 240.244
R5687 gnd.n6643 gnd.n700 240.244
R5688 gnd.n6643 gnd.n698 240.244
R5689 gnd.n6647 gnd.n698 240.244
R5690 gnd.n6647 gnd.n694 240.244
R5691 gnd.n6653 gnd.n694 240.244
R5692 gnd.n6653 gnd.n692 240.244
R5693 gnd.n6657 gnd.n692 240.244
R5694 gnd.n6657 gnd.n688 240.244
R5695 gnd.n6663 gnd.n688 240.244
R5696 gnd.n6663 gnd.n686 240.244
R5697 gnd.n6667 gnd.n686 240.244
R5698 gnd.n6667 gnd.n682 240.244
R5699 gnd.n6673 gnd.n682 240.244
R5700 gnd.n6673 gnd.n680 240.244
R5701 gnd.n6677 gnd.n680 240.244
R5702 gnd.n6677 gnd.n676 240.244
R5703 gnd.n6683 gnd.n676 240.244
R5704 gnd.n6683 gnd.n674 240.244
R5705 gnd.n6687 gnd.n674 240.244
R5706 gnd.n6687 gnd.n670 240.244
R5707 gnd.n6693 gnd.n670 240.244
R5708 gnd.n6693 gnd.n668 240.244
R5709 gnd.n6697 gnd.n668 240.244
R5710 gnd.n6697 gnd.n664 240.244
R5711 gnd.n6703 gnd.n664 240.244
R5712 gnd.n6703 gnd.n662 240.244
R5713 gnd.n6707 gnd.n662 240.244
R5714 gnd.n6707 gnd.n658 240.244
R5715 gnd.n6713 gnd.n658 240.244
R5716 gnd.n6713 gnd.n656 240.244
R5717 gnd.n6717 gnd.n656 240.244
R5718 gnd.n6717 gnd.n652 240.244
R5719 gnd.n6723 gnd.n652 240.244
R5720 gnd.n6723 gnd.n650 240.244
R5721 gnd.n6727 gnd.n650 240.244
R5722 gnd.n6727 gnd.n646 240.244
R5723 gnd.n6733 gnd.n646 240.244
R5724 gnd.n6733 gnd.n644 240.244
R5725 gnd.n6737 gnd.n644 240.244
R5726 gnd.n6737 gnd.n640 240.244
R5727 gnd.n6743 gnd.n640 240.244
R5728 gnd.n6743 gnd.n638 240.244
R5729 gnd.n6747 gnd.n638 240.244
R5730 gnd.n6747 gnd.n634 240.244
R5731 gnd.n6753 gnd.n634 240.244
R5732 gnd.n6753 gnd.n632 240.244
R5733 gnd.n6757 gnd.n632 240.244
R5734 gnd.n6757 gnd.n628 240.244
R5735 gnd.n6763 gnd.n628 240.244
R5736 gnd.n6763 gnd.n626 240.244
R5737 gnd.n6767 gnd.n626 240.244
R5738 gnd.n6767 gnd.n622 240.244
R5739 gnd.n6773 gnd.n622 240.244
R5740 gnd.n6773 gnd.n620 240.244
R5741 gnd.n6777 gnd.n620 240.244
R5742 gnd.n6777 gnd.n616 240.244
R5743 gnd.n6783 gnd.n616 240.244
R5744 gnd.n6783 gnd.n614 240.244
R5745 gnd.n6787 gnd.n614 240.244
R5746 gnd.n6787 gnd.n610 240.244
R5747 gnd.n6793 gnd.n610 240.244
R5748 gnd.n6793 gnd.n608 240.244
R5749 gnd.n6797 gnd.n608 240.244
R5750 gnd.n6797 gnd.n604 240.244
R5751 gnd.n6803 gnd.n604 240.244
R5752 gnd.n6803 gnd.n602 240.244
R5753 gnd.n6807 gnd.n602 240.244
R5754 gnd.n6807 gnd.n598 240.244
R5755 gnd.n6813 gnd.n598 240.244
R5756 gnd.n6813 gnd.n596 240.244
R5757 gnd.n6817 gnd.n596 240.244
R5758 gnd.n6817 gnd.n592 240.244
R5759 gnd.n6823 gnd.n592 240.244
R5760 gnd.n6823 gnd.n590 240.244
R5761 gnd.n6827 gnd.n590 240.244
R5762 gnd.n6827 gnd.n586 240.244
R5763 gnd.n6833 gnd.n586 240.244
R5764 gnd.n6833 gnd.n584 240.244
R5765 gnd.n6837 gnd.n584 240.244
R5766 gnd.n6837 gnd.n580 240.244
R5767 gnd.n6843 gnd.n580 240.244
R5768 gnd.n6843 gnd.n578 240.244
R5769 gnd.n6847 gnd.n578 240.244
R5770 gnd.n6847 gnd.n574 240.244
R5771 gnd.n6853 gnd.n574 240.244
R5772 gnd.n6853 gnd.n572 240.244
R5773 gnd.n6857 gnd.n572 240.244
R5774 gnd.n6857 gnd.n568 240.244
R5775 gnd.n6863 gnd.n568 240.244
R5776 gnd.n6863 gnd.n566 240.244
R5777 gnd.n6867 gnd.n566 240.244
R5778 gnd.n6867 gnd.n562 240.244
R5779 gnd.n6873 gnd.n562 240.244
R5780 gnd.n6873 gnd.n560 240.244
R5781 gnd.n6877 gnd.n560 240.244
R5782 gnd.n6877 gnd.n556 240.244
R5783 gnd.n6883 gnd.n556 240.244
R5784 gnd.n6883 gnd.n554 240.244
R5785 gnd.n6887 gnd.n554 240.244
R5786 gnd.n6887 gnd.n550 240.244
R5787 gnd.n6894 gnd.n550 240.244
R5788 gnd.n6894 gnd.n548 240.244
R5789 gnd.n6898 gnd.n548 240.244
R5790 gnd.n6898 gnd.n545 240.244
R5791 gnd.n6904 gnd.n543 240.244
R5792 gnd.n6908 gnd.n543 240.244
R5793 gnd.n6908 gnd.n539 240.244
R5794 gnd.n6914 gnd.n539 240.244
R5795 gnd.n6914 gnd.n537 240.244
R5796 gnd.n6918 gnd.n537 240.244
R5797 gnd.n6918 gnd.n533 240.244
R5798 gnd.n6924 gnd.n533 240.244
R5799 gnd.n6924 gnd.n531 240.244
R5800 gnd.n6928 gnd.n531 240.244
R5801 gnd.n6928 gnd.n527 240.244
R5802 gnd.n6934 gnd.n527 240.244
R5803 gnd.n6934 gnd.n525 240.244
R5804 gnd.n6938 gnd.n525 240.244
R5805 gnd.n6938 gnd.n521 240.244
R5806 gnd.n6944 gnd.n521 240.244
R5807 gnd.n6944 gnd.n519 240.244
R5808 gnd.n6948 gnd.n519 240.244
R5809 gnd.n6948 gnd.n515 240.244
R5810 gnd.n6954 gnd.n515 240.244
R5811 gnd.n6954 gnd.n513 240.244
R5812 gnd.n6958 gnd.n513 240.244
R5813 gnd.n6958 gnd.n509 240.244
R5814 gnd.n6964 gnd.n509 240.244
R5815 gnd.n6964 gnd.n507 240.244
R5816 gnd.n6968 gnd.n507 240.244
R5817 gnd.n6968 gnd.n503 240.244
R5818 gnd.n6974 gnd.n503 240.244
R5819 gnd.n6974 gnd.n501 240.244
R5820 gnd.n6978 gnd.n501 240.244
R5821 gnd.n6978 gnd.n497 240.244
R5822 gnd.n6984 gnd.n497 240.244
R5823 gnd.n6984 gnd.n495 240.244
R5824 gnd.n6988 gnd.n495 240.244
R5825 gnd.n6988 gnd.n491 240.244
R5826 gnd.n6994 gnd.n491 240.244
R5827 gnd.n6994 gnd.n489 240.244
R5828 gnd.n6998 gnd.n489 240.244
R5829 gnd.n6998 gnd.n485 240.244
R5830 gnd.n7004 gnd.n485 240.244
R5831 gnd.n7004 gnd.n483 240.244
R5832 gnd.n7008 gnd.n483 240.244
R5833 gnd.n7008 gnd.n479 240.244
R5834 gnd.n7014 gnd.n479 240.244
R5835 gnd.n7014 gnd.n477 240.244
R5836 gnd.n7018 gnd.n477 240.244
R5837 gnd.n7018 gnd.n473 240.244
R5838 gnd.n7024 gnd.n473 240.244
R5839 gnd.n7024 gnd.n471 240.244
R5840 gnd.n7028 gnd.n471 240.244
R5841 gnd.n7028 gnd.n467 240.244
R5842 gnd.n7034 gnd.n467 240.244
R5843 gnd.n7034 gnd.n465 240.244
R5844 gnd.n7038 gnd.n465 240.244
R5845 gnd.n7038 gnd.n461 240.244
R5846 gnd.n7044 gnd.n461 240.244
R5847 gnd.n7044 gnd.n459 240.244
R5848 gnd.n7048 gnd.n459 240.244
R5849 gnd.n7048 gnd.n455 240.244
R5850 gnd.n7054 gnd.n455 240.244
R5851 gnd.n7054 gnd.n453 240.244
R5852 gnd.n7058 gnd.n453 240.244
R5853 gnd.n7058 gnd.n449 240.244
R5854 gnd.n7064 gnd.n449 240.244
R5855 gnd.n7064 gnd.n447 240.244
R5856 gnd.n7068 gnd.n447 240.244
R5857 gnd.n7068 gnd.n443 240.244
R5858 gnd.n7074 gnd.n443 240.244
R5859 gnd.n7074 gnd.n441 240.244
R5860 gnd.n7078 gnd.n441 240.244
R5861 gnd.n7078 gnd.n437 240.244
R5862 gnd.n7084 gnd.n437 240.244
R5863 gnd.n7084 gnd.n435 240.244
R5864 gnd.n7088 gnd.n435 240.244
R5865 gnd.n7088 gnd.n431 240.244
R5866 gnd.n7094 gnd.n431 240.244
R5867 gnd.n7094 gnd.n429 240.244
R5868 gnd.n7098 gnd.n429 240.244
R5869 gnd.n7098 gnd.n425 240.244
R5870 gnd.n7104 gnd.n425 240.244
R5871 gnd.n7104 gnd.n423 240.244
R5872 gnd.n7109 gnd.n423 240.244
R5873 gnd.n7109 gnd.n419 240.244
R5874 gnd.n7116 gnd.n419 240.244
R5875 gnd.n6307 gnd.n966 240.244
R5876 gnd.n2397 gnd.n966 240.244
R5877 gnd.n2414 gnd.n2397 240.244
R5878 gnd.n2414 gnd.n2398 240.244
R5879 gnd.n2410 gnd.n2398 240.244
R5880 gnd.n2410 gnd.n2409 240.244
R5881 gnd.n2409 gnd.n2408 240.244
R5882 gnd.n2408 gnd.n2368 240.244
R5883 gnd.n4335 gnd.n2368 240.244
R5884 gnd.n4335 gnd.n4334 240.244
R5885 gnd.n4334 gnd.n2369 240.244
R5886 gnd.n2381 gnd.n2369 240.244
R5887 gnd.n4324 gnd.n2381 240.244
R5888 gnd.n4324 gnd.n4321 240.244
R5889 gnd.n4321 gnd.n4320 240.244
R5890 gnd.n4320 gnd.n4317 240.244
R5891 gnd.n4317 gnd.n2387 240.244
R5892 gnd.n2387 gnd.n2384 240.244
R5893 gnd.n2384 gnd.n2383 240.244
R5894 gnd.n2383 gnd.n2357 240.244
R5895 gnd.n4361 gnd.n2357 240.244
R5896 gnd.n4361 gnd.n2358 240.244
R5897 gnd.n4357 gnd.n2358 240.244
R5898 gnd.n4357 gnd.n4356 240.244
R5899 gnd.n4356 gnd.n4355 240.244
R5900 gnd.n4355 gnd.n4344 240.244
R5901 gnd.n4351 gnd.n4344 240.244
R5902 gnd.n4351 gnd.n2338 240.244
R5903 gnd.n4411 gnd.n2338 240.244
R5904 gnd.n4412 gnd.n4411 240.244
R5905 gnd.n4412 gnd.n2334 240.244
R5906 gnd.n4418 gnd.n2334 240.244
R5907 gnd.n4419 gnd.n4418 240.244
R5908 gnd.n4420 gnd.n4419 240.244
R5909 gnd.n4420 gnd.n2330 240.244
R5910 gnd.n4426 gnd.n2330 240.244
R5911 gnd.n4427 gnd.n4426 240.244
R5912 gnd.n4428 gnd.n4427 240.244
R5913 gnd.n4428 gnd.n2326 240.244
R5914 gnd.n4434 gnd.n2326 240.244
R5915 gnd.n4435 gnd.n4434 240.244
R5916 gnd.n4438 gnd.n4435 240.244
R5917 gnd.n4438 gnd.n2320 240.244
R5918 gnd.n4446 gnd.n2320 240.244
R5919 gnd.n4446 gnd.n2321 240.244
R5920 gnd.n2321 gnd.n2297 240.244
R5921 gnd.n4470 gnd.n2297 240.244
R5922 gnd.n4470 gnd.n2292 240.244
R5923 gnd.n4479 gnd.n2292 240.244
R5924 gnd.n4479 gnd.n2293 240.244
R5925 gnd.n2293 gnd.n1482 240.244
R5926 gnd.n5990 gnd.n1482 240.244
R5927 gnd.n5990 gnd.n1483 240.244
R5928 gnd.n5986 gnd.n1483 240.244
R5929 gnd.n5986 gnd.n1489 240.244
R5930 gnd.n4515 gnd.n1489 240.244
R5931 gnd.n4515 gnd.n2171 240.244
R5932 gnd.n4552 gnd.n2171 240.244
R5933 gnd.n4552 gnd.n2167 240.244
R5934 gnd.n4558 gnd.n2167 240.244
R5935 gnd.n4558 gnd.n2153 240.244
R5936 gnd.n4594 gnd.n2153 240.244
R5937 gnd.n4594 gnd.n2148 240.244
R5938 gnd.n4602 gnd.n2148 240.244
R5939 gnd.n4602 gnd.n2149 240.244
R5940 gnd.n2149 gnd.n2127 240.244
R5941 gnd.n4656 gnd.n2127 240.244
R5942 gnd.n4656 gnd.n2123 240.244
R5943 gnd.n4662 gnd.n2123 240.244
R5944 gnd.n4662 gnd.n2109 240.244
R5945 gnd.n4684 gnd.n2109 240.244
R5946 gnd.n4684 gnd.n2104 240.244
R5947 gnd.n4692 gnd.n2104 240.244
R5948 gnd.n4692 gnd.n2105 240.244
R5949 gnd.n2105 gnd.n2076 240.244
R5950 gnd.n4734 gnd.n2076 240.244
R5951 gnd.n4734 gnd.n2072 240.244
R5952 gnd.n4740 gnd.n2072 240.244
R5953 gnd.n4740 gnd.n2053 240.244
R5954 gnd.n4774 gnd.n2053 240.244
R5955 gnd.n4774 gnd.n2049 240.244
R5956 gnd.n4780 gnd.n2049 240.244
R5957 gnd.n4780 gnd.n2031 240.244
R5958 gnd.n4831 gnd.n2031 240.244
R5959 gnd.n4831 gnd.n2027 240.244
R5960 gnd.n4837 gnd.n2027 240.244
R5961 gnd.n4837 gnd.n2011 240.244
R5962 gnd.n4856 gnd.n2011 240.244
R5963 gnd.n4856 gnd.n2007 240.244
R5964 gnd.n4862 gnd.n2007 240.244
R5965 gnd.n4862 gnd.n1991 240.244
R5966 gnd.n4916 gnd.n1991 240.244
R5967 gnd.n4916 gnd.n1987 240.244
R5968 gnd.n4922 gnd.n1987 240.244
R5969 gnd.n4922 gnd.n1969 240.244
R5970 gnd.n4945 gnd.n1969 240.244
R5971 gnd.n4945 gnd.n1964 240.244
R5972 gnd.n4953 gnd.n1964 240.244
R5973 gnd.n4953 gnd.n1965 240.244
R5974 gnd.n1965 gnd.n1941 240.244
R5975 gnd.n4996 gnd.n1941 240.244
R5976 gnd.n4996 gnd.n1937 240.244
R5977 gnd.n5002 gnd.n1937 240.244
R5978 gnd.n5002 gnd.n1921 240.244
R5979 gnd.n5022 gnd.n1921 240.244
R5980 gnd.n5022 gnd.n1916 240.244
R5981 gnd.n5030 gnd.n1916 240.244
R5982 gnd.n5030 gnd.n1917 240.244
R5983 gnd.n1917 gnd.n1891 240.244
R5984 gnd.n5066 gnd.n1891 240.244
R5985 gnd.n5066 gnd.n1885 240.244
R5986 gnd.n5075 gnd.n1885 240.244
R5987 gnd.n5075 gnd.n1887 240.244
R5988 gnd.n1887 gnd.n1837 240.244
R5989 gnd.n5321 gnd.n1837 240.244
R5990 gnd.n5321 gnd.n1838 240.244
R5991 gnd.n5317 gnd.n1838 240.244
R5992 gnd.n5317 gnd.n5316 240.244
R5993 gnd.n5316 gnd.n1844 240.244
R5994 gnd.n5309 gnd.n1844 240.244
R5995 gnd.n5309 gnd.n1849 240.244
R5996 gnd.n5305 gnd.n1849 240.244
R5997 gnd.n5305 gnd.n1859 240.244
R5998 gnd.n1859 gnd.n1589 240.244
R5999 gnd.n5872 gnd.n1589 240.244
R6000 gnd.n5872 gnd.n1590 240.244
R6001 gnd.n5868 gnd.n1590 240.244
R6002 gnd.n5868 gnd.n1596 240.244
R6003 gnd.n5864 gnd.n1596 240.244
R6004 gnd.n5864 gnd.n1599 240.244
R6005 gnd.n5860 gnd.n1599 240.244
R6006 gnd.n5860 gnd.n1605 240.244
R6007 gnd.n5706 gnd.n1605 240.244
R6008 gnd.n5706 gnd.n5703 240.244
R6009 gnd.n5712 gnd.n5703 240.244
R6010 gnd.n5713 gnd.n5712 240.244
R6011 gnd.n5714 gnd.n5713 240.244
R6012 gnd.n5714 gnd.n5699 240.244
R6013 gnd.n5720 gnd.n5699 240.244
R6014 gnd.n5721 gnd.n5720 240.244
R6015 gnd.n5722 gnd.n5721 240.244
R6016 gnd.n5722 gnd.n1736 240.244
R6017 gnd.n5740 gnd.n1736 240.244
R6018 gnd.n5740 gnd.n1737 240.244
R6019 gnd.n5736 gnd.n1737 240.244
R6020 gnd.n5736 gnd.n5735 240.244
R6021 gnd.n5735 gnd.n5734 240.244
R6022 gnd.n5734 gnd.n1700 240.244
R6023 gnd.n5804 gnd.n1700 240.244
R6024 gnd.n5804 gnd.n1701 240.244
R6025 gnd.n5799 gnd.n1701 240.244
R6026 gnd.n5799 gnd.n1704 240.244
R6027 gnd.n1721 gnd.n1704 240.244
R6028 gnd.n1721 gnd.n1716 240.244
R6029 gnd.n1716 gnd.n402 240.244
R6030 gnd.n7135 gnd.n402 240.244
R6031 gnd.n7135 gnd.n403 240.244
R6032 gnd.n7130 gnd.n403 240.244
R6033 gnd.n7130 gnd.n7129 240.244
R6034 gnd.n7129 gnd.n7128 240.244
R6035 gnd.n7128 gnd.n407 240.244
R6036 gnd.n7124 gnd.n407 240.244
R6037 gnd.n7124 gnd.n7123 240.244
R6038 gnd.n7123 gnd.n7122 240.244
R6039 gnd.n7122 gnd.n413 240.244
R6040 gnd.n7118 gnd.n413 240.244
R6041 gnd.n7118 gnd.n7117 240.244
R6042 gnd.n6477 gnd.n796 240.244
R6043 gnd.n6477 gnd.n799 240.244
R6044 gnd.n6473 gnd.n799 240.244
R6045 gnd.n6473 gnd.n801 240.244
R6046 gnd.n6469 gnd.n801 240.244
R6047 gnd.n6469 gnd.n807 240.244
R6048 gnd.n6465 gnd.n807 240.244
R6049 gnd.n6465 gnd.n809 240.244
R6050 gnd.n6461 gnd.n809 240.244
R6051 gnd.n6461 gnd.n815 240.244
R6052 gnd.n6457 gnd.n815 240.244
R6053 gnd.n6457 gnd.n817 240.244
R6054 gnd.n6453 gnd.n817 240.244
R6055 gnd.n6453 gnd.n823 240.244
R6056 gnd.n6449 gnd.n823 240.244
R6057 gnd.n6449 gnd.n825 240.244
R6058 gnd.n6445 gnd.n825 240.244
R6059 gnd.n6445 gnd.n831 240.244
R6060 gnd.n6441 gnd.n831 240.244
R6061 gnd.n6441 gnd.n833 240.244
R6062 gnd.n6437 gnd.n833 240.244
R6063 gnd.n6437 gnd.n839 240.244
R6064 gnd.n6433 gnd.n839 240.244
R6065 gnd.n6433 gnd.n841 240.244
R6066 gnd.n6429 gnd.n841 240.244
R6067 gnd.n6429 gnd.n847 240.244
R6068 gnd.n6425 gnd.n847 240.244
R6069 gnd.n6425 gnd.n849 240.244
R6070 gnd.n6421 gnd.n849 240.244
R6071 gnd.n6421 gnd.n855 240.244
R6072 gnd.n6417 gnd.n855 240.244
R6073 gnd.n6417 gnd.n857 240.244
R6074 gnd.n6413 gnd.n857 240.244
R6075 gnd.n6413 gnd.n863 240.244
R6076 gnd.n6409 gnd.n863 240.244
R6077 gnd.n6409 gnd.n865 240.244
R6078 gnd.n6405 gnd.n865 240.244
R6079 gnd.n6405 gnd.n871 240.244
R6080 gnd.n6401 gnd.n871 240.244
R6081 gnd.n6401 gnd.n873 240.244
R6082 gnd.n6397 gnd.n873 240.244
R6083 gnd.n6397 gnd.n879 240.244
R6084 gnd.n6393 gnd.n879 240.244
R6085 gnd.n6393 gnd.n881 240.244
R6086 gnd.n6389 gnd.n881 240.244
R6087 gnd.n6389 gnd.n887 240.244
R6088 gnd.n6385 gnd.n887 240.244
R6089 gnd.n6385 gnd.n889 240.244
R6090 gnd.n6381 gnd.n889 240.244
R6091 gnd.n6381 gnd.n895 240.244
R6092 gnd.n6377 gnd.n895 240.244
R6093 gnd.n6377 gnd.n897 240.244
R6094 gnd.n6373 gnd.n897 240.244
R6095 gnd.n6373 gnd.n903 240.244
R6096 gnd.n6369 gnd.n903 240.244
R6097 gnd.n6369 gnd.n905 240.244
R6098 gnd.n6365 gnd.n905 240.244
R6099 gnd.n6365 gnd.n911 240.244
R6100 gnd.n6361 gnd.n911 240.244
R6101 gnd.n6361 gnd.n913 240.244
R6102 gnd.n6357 gnd.n913 240.244
R6103 gnd.n6357 gnd.n919 240.244
R6104 gnd.n6353 gnd.n919 240.244
R6105 gnd.n6353 gnd.n921 240.244
R6106 gnd.n6349 gnd.n921 240.244
R6107 gnd.n6349 gnd.n927 240.244
R6108 gnd.n6345 gnd.n927 240.244
R6109 gnd.n6345 gnd.n929 240.244
R6110 gnd.n6341 gnd.n929 240.244
R6111 gnd.n6341 gnd.n935 240.244
R6112 gnd.n6337 gnd.n935 240.244
R6113 gnd.n6337 gnd.n937 240.244
R6114 gnd.n6333 gnd.n937 240.244
R6115 gnd.n6333 gnd.n943 240.244
R6116 gnd.n6329 gnd.n943 240.244
R6117 gnd.n6329 gnd.n945 240.244
R6118 gnd.n6325 gnd.n945 240.244
R6119 gnd.n6325 gnd.n951 240.244
R6120 gnd.n6321 gnd.n951 240.244
R6121 gnd.n6321 gnd.n953 240.244
R6122 gnd.n6317 gnd.n953 240.244
R6123 gnd.n6317 gnd.n959 240.244
R6124 gnd.n6313 gnd.n959 240.244
R6125 gnd.n6313 gnd.n961 240.244
R6126 gnd.n4449 gnd.n1171 240.244
R6127 gnd.n4449 gnd.n2307 240.244
R6128 gnd.n4456 gnd.n2307 240.244
R6129 gnd.n4456 gnd.n2308 240.244
R6130 gnd.n2308 gnd.n2289 240.244
R6131 gnd.n4482 gnd.n2289 240.244
R6132 gnd.n4482 gnd.n2283 240.244
R6133 gnd.n4492 gnd.n2283 240.244
R6134 gnd.n4492 gnd.n2284 240.244
R6135 gnd.n4486 gnd.n2284 240.244
R6136 gnd.n4486 gnd.n1493 240.244
R6137 gnd.n5983 gnd.n1493 240.244
R6138 gnd.n5983 gnd.n1494 240.244
R6139 gnd.n1499 gnd.n1494 240.244
R6140 gnd.n1500 gnd.n1499 240.244
R6141 gnd.n1501 gnd.n1500 240.244
R6142 gnd.n2165 gnd.n1501 240.244
R6143 gnd.n2165 gnd.n1504 240.244
R6144 gnd.n1505 gnd.n1504 240.244
R6145 gnd.n1506 gnd.n1505 240.244
R6146 gnd.n4604 gnd.n1506 240.244
R6147 gnd.n4604 gnd.n1509 240.244
R6148 gnd.n1510 gnd.n1509 240.244
R6149 gnd.n1511 gnd.n1510 240.244
R6150 gnd.n4653 gnd.n1511 240.244
R6151 gnd.n4653 gnd.n1514 240.244
R6152 gnd.n1515 gnd.n1514 240.244
R6153 gnd.n1516 gnd.n1515 240.244
R6154 gnd.n4681 gnd.n1516 240.244
R6155 gnd.n4681 gnd.n1519 240.244
R6156 gnd.n1520 gnd.n1519 240.244
R6157 gnd.n1521 gnd.n1520 240.244
R6158 gnd.n4706 gnd.n1521 240.244
R6159 gnd.n4706 gnd.n1524 240.244
R6160 gnd.n1525 gnd.n1524 240.244
R6161 gnd.n1526 gnd.n1525 240.244
R6162 gnd.n4761 gnd.n1526 240.244
R6163 gnd.n4761 gnd.n1529 240.244
R6164 gnd.n1530 gnd.n1529 240.244
R6165 gnd.n1531 gnd.n1530 240.244
R6166 gnd.n4820 gnd.n1531 240.244
R6167 gnd.n4820 gnd.n1534 240.244
R6168 gnd.n1535 gnd.n1534 240.244
R6169 gnd.n1536 gnd.n1535 240.244
R6170 gnd.n2018 gnd.n1536 240.244
R6171 gnd.n2018 gnd.n1539 240.244
R6172 gnd.n1540 gnd.n1539 240.244
R6173 gnd.n1541 gnd.n1540 240.244
R6174 gnd.n4802 gnd.n1541 240.244
R6175 gnd.n4802 gnd.n1544 240.244
R6176 gnd.n1545 gnd.n1544 240.244
R6177 gnd.n1546 gnd.n1545 240.244
R6178 gnd.n4933 gnd.n1546 240.244
R6179 gnd.n4933 gnd.n1549 240.244
R6180 gnd.n1550 gnd.n1549 240.244
R6181 gnd.n1551 gnd.n1550 240.244
R6182 gnd.n4893 gnd.n1551 240.244
R6183 gnd.n4893 gnd.n1554 240.244
R6184 gnd.n1555 gnd.n1554 240.244
R6185 gnd.n1556 gnd.n1555 240.244
R6186 gnd.n1935 gnd.n1556 240.244
R6187 gnd.n1935 gnd.n1559 240.244
R6188 gnd.n1560 gnd.n1559 240.244
R6189 gnd.n1561 gnd.n1560 240.244
R6190 gnd.n1907 gnd.n1561 240.244
R6191 gnd.n1907 gnd.n1564 240.244
R6192 gnd.n1565 gnd.n1564 240.244
R6193 gnd.n1566 gnd.n1565 240.244
R6194 gnd.n5078 gnd.n1566 240.244
R6195 gnd.n5078 gnd.n1569 240.244
R6196 gnd.n1570 gnd.n1569 240.244
R6197 gnd.n1571 gnd.n1570 240.244
R6198 gnd.n5103 gnd.n1571 240.244
R6199 gnd.n5103 gnd.n1574 240.244
R6200 gnd.n1575 gnd.n1574 240.244
R6201 gnd.n1576 gnd.n1575 240.244
R6202 gnd.n5311 gnd.n1576 240.244
R6203 gnd.n5311 gnd.n1579 240.244
R6204 gnd.n1580 gnd.n1579 240.244
R6205 gnd.n1581 gnd.n1580 240.244
R6206 gnd.n1584 gnd.n1581 240.244
R6207 gnd.n5875 gnd.n1584 240.244
R6208 gnd.n1170 gnd.n1169 240.244
R6209 gnd.n1175 gnd.n1169 240.244
R6210 gnd.n1177 gnd.n1176 240.244
R6211 gnd.n1181 gnd.n1180 240.244
R6212 gnd.n1183 gnd.n1182 240.244
R6213 gnd.n1193 gnd.n1192 240.244
R6214 gnd.n1195 gnd.n1194 240.244
R6215 gnd.n1203 gnd.n1202 240.244
R6216 gnd.n1211 gnd.n1210 240.244
R6217 gnd.n1213 gnd.n1212 240.244
R6218 gnd.n1221 gnd.n1220 240.244
R6219 gnd.n1229 gnd.n1228 240.244
R6220 gnd.n1234 gnd.n1230 240.244
R6221 gnd.n1166 gnd.n1152 240.244
R6222 gnd.n2318 gnd.n1153 240.244
R6223 gnd.n2318 gnd.n2304 240.244
R6224 gnd.n4458 gnd.n2304 240.244
R6225 gnd.n4458 gnd.n2299 240.244
R6226 gnd.n4467 gnd.n2299 240.244
R6227 gnd.n4467 gnd.n2291 240.244
R6228 gnd.n2291 gnd.n2203 240.244
R6229 gnd.n4494 gnd.n2203 240.244
R6230 gnd.n4495 gnd.n4494 240.244
R6231 gnd.n4495 gnd.n2198 240.244
R6232 gnd.n4502 gnd.n2198 240.244
R6233 gnd.n4502 gnd.n1491 240.244
R6234 gnd.n4519 gnd.n1491 240.244
R6235 gnd.n4520 gnd.n4519 240.244
R6236 gnd.n4520 gnd.n2186 240.244
R6237 gnd.n4533 gnd.n2186 240.244
R6238 gnd.n4533 gnd.n2187 240.244
R6239 gnd.n4525 gnd.n2187 240.244
R6240 gnd.n4526 gnd.n4525 240.244
R6241 gnd.n4526 gnd.n2145 240.244
R6242 gnd.n4606 gnd.n2145 240.244
R6243 gnd.n4606 gnd.n2140 240.244
R6244 gnd.n4631 gnd.n2140 240.244
R6245 gnd.n4631 gnd.n2136 240.244
R6246 gnd.n2136 gnd.n2128 240.244
R6247 gnd.n4611 gnd.n2128 240.244
R6248 gnd.n4614 gnd.n4611 240.244
R6249 gnd.n4615 gnd.n4614 240.244
R6250 gnd.n4615 gnd.n2111 240.244
R6251 gnd.n2111 gnd.n2093 240.244
R6252 gnd.n4704 gnd.n2093 240.244
R6253 gnd.n4705 gnd.n4704 240.244
R6254 gnd.n4708 gnd.n4705 240.244
R6255 gnd.n4708 gnd.n2089 240.244
R6256 gnd.n4714 gnd.n2089 240.244
R6257 gnd.n4714 gnd.n2063 240.244
R6258 gnd.n4760 gnd.n2063 240.244
R6259 gnd.n4760 gnd.n2064 240.244
R6260 gnd.n4754 gnd.n2064 240.244
R6261 gnd.n4754 gnd.n2041 240.244
R6262 gnd.n4819 gnd.n2041 240.244
R6263 gnd.n4819 gnd.n2033 240.244
R6264 gnd.n4795 gnd.n2033 240.244
R6265 gnd.n4796 gnd.n4795 240.244
R6266 gnd.n4797 gnd.n4796 240.244
R6267 gnd.n4797 gnd.n2013 240.244
R6268 gnd.n2013 gnd.n2006 240.244
R6269 gnd.n4800 gnd.n2006 240.244
R6270 gnd.n4804 gnd.n4800 240.244
R6271 gnd.n4804 gnd.n1984 240.244
R6272 gnd.n4925 gnd.n1984 240.244
R6273 gnd.n4925 gnd.n1978 240.244
R6274 gnd.n4932 gnd.n1978 240.244
R6275 gnd.n4932 gnd.n1979 240.244
R6276 gnd.n1979 gnd.n1955 240.244
R6277 gnd.n4964 gnd.n1955 240.244
R6278 gnd.n4964 gnd.n1950 240.244
R6279 gnd.n4985 gnd.n1950 240.244
R6280 gnd.n4985 gnd.n1943 240.244
R6281 gnd.n4969 gnd.n1943 240.244
R6282 gnd.n4970 gnd.n4969 240.244
R6283 gnd.n4972 gnd.n4970 240.244
R6284 gnd.n4972 gnd.n1923 240.244
R6285 gnd.n1923 gnd.n1915 240.244
R6286 gnd.n1915 gnd.n1899 240.244
R6287 gnd.n5055 gnd.n1899 240.244
R6288 gnd.n5055 gnd.n1894 240.244
R6289 gnd.n5062 gnd.n1894 240.244
R6290 gnd.n5062 gnd.n1884 240.244
R6291 gnd.n1884 gnd.n1872 240.244
R6292 gnd.n5097 gnd.n1872 240.244
R6293 gnd.n5097 gnd.n1835 240.244
R6294 gnd.n5105 gnd.n1835 240.244
R6295 gnd.n5107 gnd.n5105 240.244
R6296 gnd.n5108 gnd.n5107 240.244
R6297 gnd.n5108 gnd.n1846 240.244
R6298 gnd.n1847 gnd.n1846 240.244
R6299 gnd.n5115 gnd.n1847 240.244
R6300 gnd.n5116 gnd.n5115 240.244
R6301 gnd.n5116 gnd.n1862 240.244
R6302 gnd.n5300 gnd.n1862 240.244
R6303 gnd.n5300 gnd.n1587 240.244
R6304 gnd.n5187 gnd.n5186 240.244
R6305 gnd.n5190 gnd.n5189 240.244
R6306 gnd.n5198 gnd.n5197 240.244
R6307 gnd.n5201 gnd.n5200 240.244
R6308 gnd.n5213 gnd.n5212 240.244
R6309 gnd.n5216 gnd.n5215 240.244
R6310 gnd.n5232 gnd.n5231 240.244
R6311 gnd.n5235 gnd.n5234 240.244
R6312 gnd.n5251 gnd.n5250 240.244
R6313 gnd.n5254 gnd.n5253 240.244
R6314 gnd.n5270 gnd.n5269 240.244
R6315 gnd.n5272 gnd.n5129 240.244
R6316 gnd.n5289 gnd.n5129 240.244
R6317 gnd.n5292 gnd.n5291 240.244
R6318 gnd.n1463 gnd.n1462 240.132
R6319 gnd.n5339 gnd.n5338 240.132
R6320 gnd.n6485 gnd.n6484 225.874
R6321 gnd.n6486 gnd.n6485 225.874
R6322 gnd.n6486 gnd.n789 225.874
R6323 gnd.n6494 gnd.n789 225.874
R6324 gnd.n6495 gnd.n6494 225.874
R6325 gnd.n6496 gnd.n6495 225.874
R6326 gnd.n6496 gnd.n783 225.874
R6327 gnd.n6504 gnd.n783 225.874
R6328 gnd.n6505 gnd.n6504 225.874
R6329 gnd.n6506 gnd.n6505 225.874
R6330 gnd.n6506 gnd.n777 225.874
R6331 gnd.n6514 gnd.n777 225.874
R6332 gnd.n6515 gnd.n6514 225.874
R6333 gnd.n6516 gnd.n6515 225.874
R6334 gnd.n6516 gnd.n771 225.874
R6335 gnd.n6524 gnd.n771 225.874
R6336 gnd.n6525 gnd.n6524 225.874
R6337 gnd.n6526 gnd.n6525 225.874
R6338 gnd.n6526 gnd.n765 225.874
R6339 gnd.n6534 gnd.n765 225.874
R6340 gnd.n6535 gnd.n6534 225.874
R6341 gnd.n6536 gnd.n6535 225.874
R6342 gnd.n6536 gnd.n759 225.874
R6343 gnd.n6544 gnd.n759 225.874
R6344 gnd.n6545 gnd.n6544 225.874
R6345 gnd.n6546 gnd.n6545 225.874
R6346 gnd.n6546 gnd.n753 225.874
R6347 gnd.n6554 gnd.n753 225.874
R6348 gnd.n6555 gnd.n6554 225.874
R6349 gnd.n6556 gnd.n6555 225.874
R6350 gnd.n6556 gnd.n747 225.874
R6351 gnd.n6564 gnd.n747 225.874
R6352 gnd.n6565 gnd.n6564 225.874
R6353 gnd.n6566 gnd.n6565 225.874
R6354 gnd.n6566 gnd.n741 225.874
R6355 gnd.n6574 gnd.n741 225.874
R6356 gnd.n6575 gnd.n6574 225.874
R6357 gnd.n6576 gnd.n6575 225.874
R6358 gnd.n6576 gnd.n735 225.874
R6359 gnd.n6584 gnd.n735 225.874
R6360 gnd.n6585 gnd.n6584 225.874
R6361 gnd.n6586 gnd.n6585 225.874
R6362 gnd.n6586 gnd.n729 225.874
R6363 gnd.n6594 gnd.n729 225.874
R6364 gnd.n6595 gnd.n6594 225.874
R6365 gnd.n6596 gnd.n6595 225.874
R6366 gnd.n6596 gnd.n723 225.874
R6367 gnd.n6604 gnd.n723 225.874
R6368 gnd.n6605 gnd.n6604 225.874
R6369 gnd.n6606 gnd.n6605 225.874
R6370 gnd.n6606 gnd.n717 225.874
R6371 gnd.n6614 gnd.n717 225.874
R6372 gnd.n6615 gnd.n6614 225.874
R6373 gnd.n6616 gnd.n6615 225.874
R6374 gnd.n6616 gnd.n711 225.874
R6375 gnd.n6624 gnd.n711 225.874
R6376 gnd.n6625 gnd.n6624 225.874
R6377 gnd.n6626 gnd.n6625 225.874
R6378 gnd.n6626 gnd.n705 225.874
R6379 gnd.n6634 gnd.n705 225.874
R6380 gnd.n6635 gnd.n6634 225.874
R6381 gnd.n6636 gnd.n6635 225.874
R6382 gnd.n6636 gnd.n699 225.874
R6383 gnd.n6644 gnd.n699 225.874
R6384 gnd.n6645 gnd.n6644 225.874
R6385 gnd.n6646 gnd.n6645 225.874
R6386 gnd.n6646 gnd.n693 225.874
R6387 gnd.n6654 gnd.n693 225.874
R6388 gnd.n6655 gnd.n6654 225.874
R6389 gnd.n6656 gnd.n6655 225.874
R6390 gnd.n6656 gnd.n687 225.874
R6391 gnd.n6664 gnd.n687 225.874
R6392 gnd.n6665 gnd.n6664 225.874
R6393 gnd.n6666 gnd.n6665 225.874
R6394 gnd.n6666 gnd.n681 225.874
R6395 gnd.n6674 gnd.n681 225.874
R6396 gnd.n6675 gnd.n6674 225.874
R6397 gnd.n6676 gnd.n6675 225.874
R6398 gnd.n6676 gnd.n675 225.874
R6399 gnd.n6684 gnd.n675 225.874
R6400 gnd.n6685 gnd.n6684 225.874
R6401 gnd.n6686 gnd.n6685 225.874
R6402 gnd.n6686 gnd.n669 225.874
R6403 gnd.n6694 gnd.n669 225.874
R6404 gnd.n6695 gnd.n6694 225.874
R6405 gnd.n6696 gnd.n6695 225.874
R6406 gnd.n6696 gnd.n663 225.874
R6407 gnd.n6704 gnd.n663 225.874
R6408 gnd.n6705 gnd.n6704 225.874
R6409 gnd.n6706 gnd.n6705 225.874
R6410 gnd.n6706 gnd.n657 225.874
R6411 gnd.n6714 gnd.n657 225.874
R6412 gnd.n6715 gnd.n6714 225.874
R6413 gnd.n6716 gnd.n6715 225.874
R6414 gnd.n6716 gnd.n651 225.874
R6415 gnd.n6724 gnd.n651 225.874
R6416 gnd.n6725 gnd.n6724 225.874
R6417 gnd.n6726 gnd.n6725 225.874
R6418 gnd.n6726 gnd.n645 225.874
R6419 gnd.n6734 gnd.n645 225.874
R6420 gnd.n6735 gnd.n6734 225.874
R6421 gnd.n6736 gnd.n6735 225.874
R6422 gnd.n6736 gnd.n639 225.874
R6423 gnd.n6744 gnd.n639 225.874
R6424 gnd.n6745 gnd.n6744 225.874
R6425 gnd.n6746 gnd.n6745 225.874
R6426 gnd.n6746 gnd.n633 225.874
R6427 gnd.n6754 gnd.n633 225.874
R6428 gnd.n6755 gnd.n6754 225.874
R6429 gnd.n6756 gnd.n6755 225.874
R6430 gnd.n6756 gnd.n627 225.874
R6431 gnd.n6764 gnd.n627 225.874
R6432 gnd.n6765 gnd.n6764 225.874
R6433 gnd.n6766 gnd.n6765 225.874
R6434 gnd.n6766 gnd.n621 225.874
R6435 gnd.n6774 gnd.n621 225.874
R6436 gnd.n6775 gnd.n6774 225.874
R6437 gnd.n6776 gnd.n6775 225.874
R6438 gnd.n6776 gnd.n615 225.874
R6439 gnd.n6784 gnd.n615 225.874
R6440 gnd.n6785 gnd.n6784 225.874
R6441 gnd.n6786 gnd.n6785 225.874
R6442 gnd.n6786 gnd.n609 225.874
R6443 gnd.n6794 gnd.n609 225.874
R6444 gnd.n6795 gnd.n6794 225.874
R6445 gnd.n6796 gnd.n6795 225.874
R6446 gnd.n6796 gnd.n603 225.874
R6447 gnd.n6804 gnd.n603 225.874
R6448 gnd.n6805 gnd.n6804 225.874
R6449 gnd.n6806 gnd.n6805 225.874
R6450 gnd.n6806 gnd.n597 225.874
R6451 gnd.n6814 gnd.n597 225.874
R6452 gnd.n6815 gnd.n6814 225.874
R6453 gnd.n6816 gnd.n6815 225.874
R6454 gnd.n6816 gnd.n591 225.874
R6455 gnd.n6824 gnd.n591 225.874
R6456 gnd.n6825 gnd.n6824 225.874
R6457 gnd.n6826 gnd.n6825 225.874
R6458 gnd.n6826 gnd.n585 225.874
R6459 gnd.n6834 gnd.n585 225.874
R6460 gnd.n6835 gnd.n6834 225.874
R6461 gnd.n6836 gnd.n6835 225.874
R6462 gnd.n6836 gnd.n579 225.874
R6463 gnd.n6844 gnd.n579 225.874
R6464 gnd.n6845 gnd.n6844 225.874
R6465 gnd.n6846 gnd.n6845 225.874
R6466 gnd.n6846 gnd.n573 225.874
R6467 gnd.n6854 gnd.n573 225.874
R6468 gnd.n6855 gnd.n6854 225.874
R6469 gnd.n6856 gnd.n6855 225.874
R6470 gnd.n6856 gnd.n567 225.874
R6471 gnd.n6864 gnd.n567 225.874
R6472 gnd.n6865 gnd.n6864 225.874
R6473 gnd.n6866 gnd.n6865 225.874
R6474 gnd.n6866 gnd.n561 225.874
R6475 gnd.n6874 gnd.n561 225.874
R6476 gnd.n6875 gnd.n6874 225.874
R6477 gnd.n6876 gnd.n6875 225.874
R6478 gnd.n6876 gnd.n555 225.874
R6479 gnd.n6884 gnd.n555 225.874
R6480 gnd.n6885 gnd.n6884 225.874
R6481 gnd.n6886 gnd.n6885 225.874
R6482 gnd.n6886 gnd.n549 225.874
R6483 gnd.n6895 gnd.n549 225.874
R6484 gnd.n6896 gnd.n6895 225.874
R6485 gnd.n6897 gnd.n6896 225.874
R6486 gnd.n6897 gnd.n544 225.874
R6487 gnd.n3005 gnd.t127 224.174
R6488 gnd.n2515 gnd.t119 224.174
R6489 gnd.n7107 gnd.n170 215.659
R6490 gnd.n6906 gnd.n6905 206.476
R6491 gnd.n6907 gnd.n6906 206.476
R6492 gnd.n6907 gnd.n538 206.476
R6493 gnd.n6915 gnd.n538 206.476
R6494 gnd.n6916 gnd.n6915 206.476
R6495 gnd.n6917 gnd.n6916 206.476
R6496 gnd.n6917 gnd.n532 206.476
R6497 gnd.n6925 gnd.n532 206.476
R6498 gnd.n6926 gnd.n6925 206.476
R6499 gnd.n6927 gnd.n6926 206.476
R6500 gnd.n6927 gnd.n526 206.476
R6501 gnd.n6935 gnd.n526 206.476
R6502 gnd.n6936 gnd.n6935 206.476
R6503 gnd.n6937 gnd.n6936 206.476
R6504 gnd.n6937 gnd.n520 206.476
R6505 gnd.n6945 gnd.n520 206.476
R6506 gnd.n6946 gnd.n6945 206.476
R6507 gnd.n6947 gnd.n6946 206.476
R6508 gnd.n6947 gnd.n514 206.476
R6509 gnd.n6955 gnd.n514 206.476
R6510 gnd.n6956 gnd.n6955 206.476
R6511 gnd.n6957 gnd.n6956 206.476
R6512 gnd.n6957 gnd.n508 206.476
R6513 gnd.n6965 gnd.n508 206.476
R6514 gnd.n6966 gnd.n6965 206.476
R6515 gnd.n6967 gnd.n6966 206.476
R6516 gnd.n6967 gnd.n502 206.476
R6517 gnd.n6975 gnd.n502 206.476
R6518 gnd.n6976 gnd.n6975 206.476
R6519 gnd.n6977 gnd.n6976 206.476
R6520 gnd.n6977 gnd.n496 206.476
R6521 gnd.n6985 gnd.n496 206.476
R6522 gnd.n6986 gnd.n6985 206.476
R6523 gnd.n6987 gnd.n6986 206.476
R6524 gnd.n6987 gnd.n490 206.476
R6525 gnd.n6995 gnd.n490 206.476
R6526 gnd.n6996 gnd.n6995 206.476
R6527 gnd.n6997 gnd.n6996 206.476
R6528 gnd.n6997 gnd.n484 206.476
R6529 gnd.n7005 gnd.n484 206.476
R6530 gnd.n7006 gnd.n7005 206.476
R6531 gnd.n7007 gnd.n7006 206.476
R6532 gnd.n7007 gnd.n478 206.476
R6533 gnd.n7015 gnd.n478 206.476
R6534 gnd.n7016 gnd.n7015 206.476
R6535 gnd.n7017 gnd.n7016 206.476
R6536 gnd.n7017 gnd.n472 206.476
R6537 gnd.n7025 gnd.n472 206.476
R6538 gnd.n7026 gnd.n7025 206.476
R6539 gnd.n7027 gnd.n7026 206.476
R6540 gnd.n7027 gnd.n466 206.476
R6541 gnd.n7035 gnd.n466 206.476
R6542 gnd.n7036 gnd.n7035 206.476
R6543 gnd.n7037 gnd.n7036 206.476
R6544 gnd.n7037 gnd.n460 206.476
R6545 gnd.n7045 gnd.n460 206.476
R6546 gnd.n7046 gnd.n7045 206.476
R6547 gnd.n7047 gnd.n7046 206.476
R6548 gnd.n7047 gnd.n454 206.476
R6549 gnd.n7055 gnd.n454 206.476
R6550 gnd.n7056 gnd.n7055 206.476
R6551 gnd.n7057 gnd.n7056 206.476
R6552 gnd.n7057 gnd.n448 206.476
R6553 gnd.n7065 gnd.n448 206.476
R6554 gnd.n7066 gnd.n7065 206.476
R6555 gnd.n7067 gnd.n7066 206.476
R6556 gnd.n7067 gnd.n442 206.476
R6557 gnd.n7075 gnd.n442 206.476
R6558 gnd.n7076 gnd.n7075 206.476
R6559 gnd.n7077 gnd.n7076 206.476
R6560 gnd.n7077 gnd.n436 206.476
R6561 gnd.n7085 gnd.n436 206.476
R6562 gnd.n7086 gnd.n7085 206.476
R6563 gnd.n7087 gnd.n7086 206.476
R6564 gnd.n7087 gnd.n430 206.476
R6565 gnd.n7095 gnd.n430 206.476
R6566 gnd.n7096 gnd.n7095 206.476
R6567 gnd.n7097 gnd.n7096 206.476
R6568 gnd.n7097 gnd.n424 206.476
R6569 gnd.n7105 gnd.n424 206.476
R6570 gnd.n7106 gnd.n7105 206.476
R6571 gnd.n7108 gnd.n7106 206.476
R6572 gnd.n7108 gnd.n7107 206.476
R6573 gnd.n5580 gnd.n5579 199.319
R6574 gnd.n5581 gnd.n5580 199.319
R6575 gnd.n1319 gnd.n1274 199.319
R6576 gnd.n1319 gnd.n1273 199.319
R6577 gnd.n1464 gnd.n1461 186.49
R6578 gnd.n5340 gnd.n5337 186.49
R6579 gnd.n3780 gnd.n3779 185
R6580 gnd.n3778 gnd.n3777 185
R6581 gnd.n3757 gnd.n3756 185
R6582 gnd.n3772 gnd.n3771 185
R6583 gnd.n3770 gnd.n3769 185
R6584 gnd.n3761 gnd.n3760 185
R6585 gnd.n3764 gnd.n3763 185
R6586 gnd.n3748 gnd.n3747 185
R6587 gnd.n3746 gnd.n3745 185
R6588 gnd.n3725 gnd.n3724 185
R6589 gnd.n3740 gnd.n3739 185
R6590 gnd.n3738 gnd.n3737 185
R6591 gnd.n3729 gnd.n3728 185
R6592 gnd.n3732 gnd.n3731 185
R6593 gnd.n3716 gnd.n3715 185
R6594 gnd.n3714 gnd.n3713 185
R6595 gnd.n3693 gnd.n3692 185
R6596 gnd.n3708 gnd.n3707 185
R6597 gnd.n3706 gnd.n3705 185
R6598 gnd.n3697 gnd.n3696 185
R6599 gnd.n3700 gnd.n3699 185
R6600 gnd.n3685 gnd.n3684 185
R6601 gnd.n3683 gnd.n3682 185
R6602 gnd.n3662 gnd.n3661 185
R6603 gnd.n3677 gnd.n3676 185
R6604 gnd.n3675 gnd.n3674 185
R6605 gnd.n3666 gnd.n3665 185
R6606 gnd.n3669 gnd.n3668 185
R6607 gnd.n3653 gnd.n3652 185
R6608 gnd.n3651 gnd.n3650 185
R6609 gnd.n3630 gnd.n3629 185
R6610 gnd.n3645 gnd.n3644 185
R6611 gnd.n3643 gnd.n3642 185
R6612 gnd.n3634 gnd.n3633 185
R6613 gnd.n3637 gnd.n3636 185
R6614 gnd.n3621 gnd.n3620 185
R6615 gnd.n3619 gnd.n3618 185
R6616 gnd.n3598 gnd.n3597 185
R6617 gnd.n3613 gnd.n3612 185
R6618 gnd.n3611 gnd.n3610 185
R6619 gnd.n3602 gnd.n3601 185
R6620 gnd.n3605 gnd.n3604 185
R6621 gnd.n3589 gnd.n3588 185
R6622 gnd.n3587 gnd.n3586 185
R6623 gnd.n3566 gnd.n3565 185
R6624 gnd.n3581 gnd.n3580 185
R6625 gnd.n3579 gnd.n3578 185
R6626 gnd.n3570 gnd.n3569 185
R6627 gnd.n3573 gnd.n3572 185
R6628 gnd.n3558 gnd.n3557 185
R6629 gnd.n3556 gnd.n3555 185
R6630 gnd.n3535 gnd.n3534 185
R6631 gnd.n3550 gnd.n3549 185
R6632 gnd.n3548 gnd.n3547 185
R6633 gnd.n3539 gnd.n3538 185
R6634 gnd.n3542 gnd.n3541 185
R6635 gnd.n3006 gnd.t126 178.987
R6636 gnd.n2516 gnd.t120 178.987
R6637 gnd.n1 gnd.t247 170.774
R6638 gnd.n7 gnd.t202 170.103
R6639 gnd.n6 gnd.t318 170.103
R6640 gnd.n5 gnd.t146 170.103
R6641 gnd.n4 gnd.t228 170.103
R6642 gnd.n3 gnd.t200 170.103
R6643 gnd.n2 gnd.t212 170.103
R6644 gnd.n1 gnd.t276 170.103
R6645 gnd.n5408 gnd.n5407 163.367
R6646 gnd.n5404 gnd.n5403 163.367
R6647 gnd.n5400 gnd.n5399 163.367
R6648 gnd.n5396 gnd.n5395 163.367
R6649 gnd.n5392 gnd.n5391 163.367
R6650 gnd.n5388 gnd.n5387 163.367
R6651 gnd.n5384 gnd.n5383 163.367
R6652 gnd.n5380 gnd.n5379 163.367
R6653 gnd.n5376 gnd.n5375 163.367
R6654 gnd.n5372 gnd.n5371 163.367
R6655 gnd.n5368 gnd.n5367 163.367
R6656 gnd.n5364 gnd.n5363 163.367
R6657 gnd.n5360 gnd.n5359 163.367
R6658 gnd.n5356 gnd.n5355 163.367
R6659 gnd.n5351 gnd.n5350 163.367
R6660 gnd.n5483 gnd.n1790 163.367
R6661 gnd.n5480 gnd.n5479 163.367
R6662 gnd.n5477 gnd.n1823 163.367
R6663 gnd.n5472 gnd.n5471 163.367
R6664 gnd.n5468 gnd.n5467 163.367
R6665 gnd.n5464 gnd.n5463 163.367
R6666 gnd.n5460 gnd.n5459 163.367
R6667 gnd.n5456 gnd.n5455 163.367
R6668 gnd.n5452 gnd.n5451 163.367
R6669 gnd.n5448 gnd.n5447 163.367
R6670 gnd.n5444 gnd.n5443 163.367
R6671 gnd.n5440 gnd.n5439 163.367
R6672 gnd.n5436 gnd.n5435 163.367
R6673 gnd.n5432 gnd.n5431 163.367
R6674 gnd.n5428 gnd.n5427 163.367
R6675 gnd.n5424 gnd.n5423 163.367
R6676 gnd.n5420 gnd.n5419 163.367
R6677 gnd.n2280 gnd.n1480 163.367
R6678 gnd.n2276 gnd.n1480 163.367
R6679 gnd.n2276 gnd.n2197 163.367
R6680 gnd.n2272 gnd.n2197 163.367
R6681 gnd.n2272 gnd.n2271 163.367
R6682 gnd.n2271 gnd.n2193 163.367
R6683 gnd.n2193 gnd.n2176 163.367
R6684 gnd.n4545 gnd.n2176 163.367
R6685 gnd.n4545 gnd.n2173 163.367
R6686 gnd.n4550 gnd.n2173 163.367
R6687 gnd.n4550 gnd.n2174 163.367
R6688 gnd.n2174 gnd.n2164 163.367
R6689 gnd.n4561 gnd.n2164 163.367
R6690 gnd.n4561 gnd.n2162 163.367
R6691 gnd.n4574 gnd.n2162 163.367
R6692 gnd.n4574 gnd.n2155 163.367
R6693 gnd.n4570 gnd.n2155 163.367
R6694 gnd.n4570 gnd.n4567 163.367
R6695 gnd.n4567 gnd.n4566 163.367
R6696 gnd.n4566 gnd.n2138 163.367
R6697 gnd.n4634 gnd.n2138 163.367
R6698 gnd.n4634 gnd.n2135 163.367
R6699 gnd.n4643 gnd.n2135 163.367
R6700 gnd.n4643 gnd.n2129 163.367
R6701 gnd.n4639 gnd.n2129 163.367
R6702 gnd.n4639 gnd.n2122 163.367
R6703 gnd.n2122 gnd.n2114 163.367
R6704 gnd.n4672 gnd.n2114 163.367
R6705 gnd.n4672 gnd.n2112 163.367
R6706 gnd.n4679 gnd.n2112 163.367
R6707 gnd.n4679 gnd.n2102 163.367
R6708 gnd.n2103 gnd.n2102 163.367
R6709 gnd.n2103 gnd.n2095 163.367
R6710 gnd.n2095 gnd.n2085 163.367
R6711 gnd.n4722 gnd.n2085 163.367
R6712 gnd.n4722 gnd.n2086 163.367
R6713 gnd.n2086 gnd.n2078 163.367
R6714 gnd.n4717 gnd.n2078 163.367
R6715 gnd.n4717 gnd.n2070 163.367
R6716 gnd.n4744 gnd.n2070 163.367
R6717 gnd.n4744 gnd.n2062 163.367
R6718 gnd.n4747 gnd.n2062 163.367
R6719 gnd.n4747 gnd.n2055 163.367
R6720 gnd.n4751 gnd.n2055 163.367
R6721 gnd.n4751 gnd.n2047 163.367
R6722 gnd.n4784 gnd.n2047 163.367
R6723 gnd.n4784 gnd.n2040 163.367
R6724 gnd.n4787 gnd.n2040 163.367
R6725 gnd.n4787 gnd.n2034 163.367
R6726 gnd.n4792 gnd.n2034 163.367
R6727 gnd.n4792 gnd.n2024 163.367
R6728 gnd.n2024 gnd.n2016 163.367
R6729 gnd.n4847 gnd.n2016 163.367
R6730 gnd.n4847 gnd.n2014 163.367
R6731 gnd.n4852 gnd.n2014 163.367
R6732 gnd.n4852 gnd.n2005 163.367
R6733 gnd.n2005 gnd.n1997 163.367
R6734 gnd.n4881 gnd.n1997 163.367
R6735 gnd.n4881 gnd.n1994 163.367
R6736 gnd.n4914 gnd.n1994 163.367
R6737 gnd.n4914 gnd.n1995 163.367
R6738 gnd.n4910 gnd.n1995 163.367
R6739 gnd.n4910 gnd.n4909 163.367
R6740 gnd.n4909 gnd.n1976 163.367
R6741 gnd.n1977 gnd.n1976 163.367
R6742 gnd.n1977 gnd.n1970 163.367
R6743 gnd.n4903 gnd.n1970 163.367
R6744 gnd.n4903 gnd.n1963 163.367
R6745 gnd.n4899 gnd.n1963 163.367
R6746 gnd.n4899 gnd.n1957 163.367
R6747 gnd.n4896 gnd.n1957 163.367
R6748 gnd.n4896 gnd.n1949 163.367
R6749 gnd.n4889 gnd.n1949 163.367
R6750 gnd.n4889 gnd.n1944 163.367
R6751 gnd.n4886 gnd.n1944 163.367
R6752 gnd.n4886 gnd.n1932 163.367
R6753 gnd.n1932 gnd.n1926 163.367
R6754 gnd.n5012 gnd.n1926 163.367
R6755 gnd.n5012 gnd.n1924 163.367
R6756 gnd.n5017 gnd.n1924 163.367
R6757 gnd.n5017 gnd.n1914 163.367
R6758 gnd.n1914 gnd.n1906 163.367
R6759 gnd.n5045 gnd.n1906 163.367
R6760 gnd.n5045 gnd.n1903 163.367
R6761 gnd.n5052 gnd.n1903 163.367
R6762 gnd.n5052 gnd.n1904 163.367
R6763 gnd.n1904 gnd.n1893 163.367
R6764 gnd.n1893 gnd.n1883 163.367
R6765 gnd.n1883 gnd.n1876 163.367
R6766 gnd.n5088 gnd.n1876 163.367
R6767 gnd.n5088 gnd.n1874 163.367
R6768 gnd.n5094 gnd.n1874 163.367
R6769 gnd.n5094 gnd.n1834 163.367
R6770 gnd.n1834 gnd.n1827 163.367
R6771 gnd.n5415 gnd.n1827 163.367
R6772 gnd.n1455 gnd.n1454 163.367
R6773 gnd.n6055 gnd.n1454 163.367
R6774 gnd.n6053 gnd.n6052 163.367
R6775 gnd.n6049 gnd.n6048 163.367
R6776 gnd.n6045 gnd.n6044 163.367
R6777 gnd.n6041 gnd.n6040 163.367
R6778 gnd.n6037 gnd.n6036 163.367
R6779 gnd.n6033 gnd.n6032 163.367
R6780 gnd.n6029 gnd.n6028 163.367
R6781 gnd.n6025 gnd.n6024 163.367
R6782 gnd.n6021 gnd.n6020 163.367
R6783 gnd.n6017 gnd.n6016 163.367
R6784 gnd.n6013 gnd.n6012 163.367
R6785 gnd.n6009 gnd.n6008 163.367
R6786 gnd.n6005 gnd.n6004 163.367
R6787 gnd.n6001 gnd.n6000 163.367
R6788 gnd.n6064 gnd.n1420 163.367
R6789 gnd.n2209 gnd.n2208 163.367
R6790 gnd.n2214 gnd.n2213 163.367
R6791 gnd.n2218 gnd.n2217 163.367
R6792 gnd.n2222 gnd.n2221 163.367
R6793 gnd.n2226 gnd.n2225 163.367
R6794 gnd.n2230 gnd.n2229 163.367
R6795 gnd.n2234 gnd.n2233 163.367
R6796 gnd.n2238 gnd.n2237 163.367
R6797 gnd.n2242 gnd.n2241 163.367
R6798 gnd.n2246 gnd.n2245 163.367
R6799 gnd.n2250 gnd.n2249 163.367
R6800 gnd.n2254 gnd.n2253 163.367
R6801 gnd.n2258 gnd.n2257 163.367
R6802 gnd.n2262 gnd.n2261 163.367
R6803 gnd.n2266 gnd.n2265 163.367
R6804 gnd.n5993 gnd.n1456 163.367
R6805 gnd.n5993 gnd.n1478 163.367
R6806 gnd.n4505 gnd.n1478 163.367
R6807 gnd.n4506 gnd.n4505 163.367
R6808 gnd.n4506 gnd.n2194 163.367
R6809 gnd.n4510 gnd.n2194 163.367
R6810 gnd.n4510 gnd.n2179 163.367
R6811 gnd.n4543 gnd.n2179 163.367
R6812 gnd.n4543 gnd.n2180 163.367
R6813 gnd.n2180 gnd.n2172 163.367
R6814 gnd.n4538 gnd.n2172 163.367
R6815 gnd.n4538 gnd.n2183 163.367
R6816 gnd.n2183 gnd.n2160 163.367
R6817 gnd.n4578 gnd.n2160 163.367
R6818 gnd.n4578 gnd.n2157 163.367
R6819 gnd.n4591 gnd.n2157 163.367
R6820 gnd.n4591 gnd.n2158 163.367
R6821 gnd.n4587 gnd.n2158 163.367
R6822 gnd.n4587 gnd.n4586 163.367
R6823 gnd.n4586 gnd.n4585 163.367
R6824 gnd.n4585 gnd.n2133 163.367
R6825 gnd.n4647 gnd.n2133 163.367
R6826 gnd.n4647 gnd.n2131 163.367
R6827 gnd.n4651 gnd.n2131 163.367
R6828 gnd.n4651 gnd.n2120 163.367
R6829 gnd.n4665 gnd.n2120 163.367
R6830 gnd.n4665 gnd.n2117 163.367
R6831 gnd.n4670 gnd.n2117 163.367
R6832 gnd.n4670 gnd.n2118 163.367
R6833 gnd.n2118 gnd.n2100 163.367
R6834 gnd.n4697 gnd.n2100 163.367
R6835 gnd.n4697 gnd.n2098 163.367
R6836 gnd.n4701 gnd.n2098 163.367
R6837 gnd.n4701 gnd.n2083 163.367
R6838 gnd.n4724 gnd.n2083 163.367
R6839 gnd.n4724 gnd.n2080 163.367
R6840 gnd.n4731 gnd.n2080 163.367
R6841 gnd.n4731 gnd.n2081 163.367
R6842 gnd.n4727 gnd.n2081 163.367
R6843 gnd.n4727 gnd.n2060 163.367
R6844 gnd.n4764 gnd.n2060 163.367
R6845 gnd.n4764 gnd.n2057 163.367
R6846 gnd.n4771 gnd.n2057 163.367
R6847 gnd.n4771 gnd.n2058 163.367
R6848 gnd.n4767 gnd.n2058 163.367
R6849 gnd.n4767 gnd.n2038 163.367
R6850 gnd.n4823 gnd.n2038 163.367
R6851 gnd.n4823 gnd.n2036 163.367
R6852 gnd.n4827 gnd.n2036 163.367
R6853 gnd.n4827 gnd.n2023 163.367
R6854 gnd.n4840 gnd.n2023 163.367
R6855 gnd.n4840 gnd.n2020 163.367
R6856 gnd.n4845 gnd.n2020 163.367
R6857 gnd.n4845 gnd.n2021 163.367
R6858 gnd.n2021 gnd.n2003 163.367
R6859 gnd.n4867 gnd.n2003 163.367
R6860 gnd.n4867 gnd.n2000 163.367
R6861 gnd.n4879 gnd.n2000 163.367
R6862 gnd.n4879 gnd.n2001 163.367
R6863 gnd.n2001 gnd.n1992 163.367
R6864 gnd.n4874 gnd.n1992 163.367
R6865 gnd.n4874 gnd.n4871 163.367
R6866 gnd.n4871 gnd.n1974 163.367
R6867 gnd.n4938 gnd.n1974 163.367
R6868 gnd.n4938 gnd.n1972 163.367
R6869 gnd.n4942 gnd.n1972 163.367
R6870 gnd.n4942 gnd.n1961 163.367
R6871 gnd.n4957 gnd.n1961 163.367
R6872 gnd.n4957 gnd.n1959 163.367
R6873 gnd.n4961 gnd.n1959 163.367
R6874 gnd.n4961 gnd.n1948 163.367
R6875 gnd.n4988 gnd.n1948 163.367
R6876 gnd.n4988 gnd.n1946 163.367
R6877 gnd.n4992 gnd.n1946 163.367
R6878 gnd.n4992 gnd.n1930 163.367
R6879 gnd.n5005 gnd.n1930 163.367
R6880 gnd.n5005 gnd.n1927 163.367
R6881 gnd.n5010 gnd.n1927 163.367
R6882 gnd.n5010 gnd.n1928 163.367
R6883 gnd.n1928 gnd.n1913 163.367
R6884 gnd.n5035 gnd.n1913 163.367
R6885 gnd.n5035 gnd.n1910 163.367
R6886 gnd.n5043 gnd.n1910 163.367
R6887 gnd.n5043 gnd.n1911 163.367
R6888 gnd.n1911 gnd.n1901 163.367
R6889 gnd.n5038 gnd.n1901 163.367
R6890 gnd.n5038 gnd.n1881 163.367
R6891 gnd.n5081 gnd.n1881 163.367
R6892 gnd.n5081 gnd.n1878 163.367
R6893 gnd.n5086 gnd.n1878 163.367
R6894 gnd.n5086 gnd.n1879 163.367
R6895 gnd.n1879 gnd.n1832 163.367
R6896 gnd.n5325 gnd.n1832 163.367
R6897 gnd.n5325 gnd.n1829 163.367
R6898 gnd.n5413 gnd.n1829 163.367
R6899 gnd.n5346 gnd.n5345 156.462
R6900 gnd.n3720 gnd.n3688 153.042
R6901 gnd.n3784 gnd.n3783 152.079
R6902 gnd.n3752 gnd.n3751 152.079
R6903 gnd.n3720 gnd.n3719 152.079
R6904 gnd.n1469 gnd.n1468 152
R6905 gnd.n1470 gnd.n1459 152
R6906 gnd.n1472 gnd.n1471 152
R6907 gnd.n1474 gnd.n1457 152
R6908 gnd.n1476 gnd.n1475 152
R6909 gnd.n5344 gnd.n5328 152
R6910 gnd.n5336 gnd.n5329 152
R6911 gnd.n5335 gnd.n5334 152
R6912 gnd.n5333 gnd.n5330 152
R6913 gnd.n5331 gnd.t29 150.546
R6914 gnd.t193 gnd.n3762 147.661
R6915 gnd.t311 gnd.n3730 147.661
R6916 gnd.t221 gnd.n3698 147.661
R6917 gnd.t290 gnd.n3667 147.661
R6918 gnd.t144 gnd.n3635 147.661
R6919 gnd.t323 gnd.n3603 147.661
R6920 gnd.t327 gnd.n3571 147.661
R6921 gnd.t325 gnd.n3540 147.661
R6922 gnd.n5482 gnd.n1789 143.351
R6923 gnd.n1436 gnd.n1419 143.351
R6924 gnd.n6063 gnd.n1419 143.351
R6925 gnd.n1466 gnd.t83 130.484
R6926 gnd.n1475 gnd.t108 126.766
R6927 gnd.n1473 gnd.t39 126.766
R6928 gnd.n1459 gnd.t102 126.766
R6929 gnd.n1467 gnd.t63 126.766
R6930 gnd.n5332 gnd.t14 126.766
R6931 gnd.n5334 gnd.t128 126.766
R6932 gnd.n5343 gnd.t76 126.766
R6933 gnd.n5345 gnd.t53 126.766
R6934 gnd.n3779 gnd.n3778 104.615
R6935 gnd.n3778 gnd.n3756 104.615
R6936 gnd.n3771 gnd.n3756 104.615
R6937 gnd.n3771 gnd.n3770 104.615
R6938 gnd.n3770 gnd.n3760 104.615
R6939 gnd.n3763 gnd.n3760 104.615
R6940 gnd.n3747 gnd.n3746 104.615
R6941 gnd.n3746 gnd.n3724 104.615
R6942 gnd.n3739 gnd.n3724 104.615
R6943 gnd.n3739 gnd.n3738 104.615
R6944 gnd.n3738 gnd.n3728 104.615
R6945 gnd.n3731 gnd.n3728 104.615
R6946 gnd.n3715 gnd.n3714 104.615
R6947 gnd.n3714 gnd.n3692 104.615
R6948 gnd.n3707 gnd.n3692 104.615
R6949 gnd.n3707 gnd.n3706 104.615
R6950 gnd.n3706 gnd.n3696 104.615
R6951 gnd.n3699 gnd.n3696 104.615
R6952 gnd.n3684 gnd.n3683 104.615
R6953 gnd.n3683 gnd.n3661 104.615
R6954 gnd.n3676 gnd.n3661 104.615
R6955 gnd.n3676 gnd.n3675 104.615
R6956 gnd.n3675 gnd.n3665 104.615
R6957 gnd.n3668 gnd.n3665 104.615
R6958 gnd.n3652 gnd.n3651 104.615
R6959 gnd.n3651 gnd.n3629 104.615
R6960 gnd.n3644 gnd.n3629 104.615
R6961 gnd.n3644 gnd.n3643 104.615
R6962 gnd.n3643 gnd.n3633 104.615
R6963 gnd.n3636 gnd.n3633 104.615
R6964 gnd.n3620 gnd.n3619 104.615
R6965 gnd.n3619 gnd.n3597 104.615
R6966 gnd.n3612 gnd.n3597 104.615
R6967 gnd.n3612 gnd.n3611 104.615
R6968 gnd.n3611 gnd.n3601 104.615
R6969 gnd.n3604 gnd.n3601 104.615
R6970 gnd.n3588 gnd.n3587 104.615
R6971 gnd.n3587 gnd.n3565 104.615
R6972 gnd.n3580 gnd.n3565 104.615
R6973 gnd.n3580 gnd.n3579 104.615
R6974 gnd.n3579 gnd.n3569 104.615
R6975 gnd.n3572 gnd.n3569 104.615
R6976 gnd.n3557 gnd.n3556 104.615
R6977 gnd.n3556 gnd.n3534 104.615
R6978 gnd.n3549 gnd.n3534 104.615
R6979 gnd.n3549 gnd.n3548 104.615
R6980 gnd.n3548 gnd.n3538 104.615
R6981 gnd.n3541 gnd.n3538 104.615
R6982 gnd.n2931 gnd.t62 100.632
R6983 gnd.n2489 gnd.t94 100.632
R6984 gnd.n242 gnd.n240 99.6594
R6985 gnd.n248 gnd.n233 99.6594
R6986 gnd.n252 gnd.n250 99.6594
R6987 gnd.n258 gnd.n229 99.6594
R6988 gnd.n262 gnd.n260 99.6594
R6989 gnd.n268 gnd.n225 99.6594
R6990 gnd.n273 gnd.n270 99.6594
R6991 gnd.n271 gnd.n221 99.6594
R6992 gnd.n283 gnd.n281 99.6594
R6993 gnd.n289 gnd.n215 99.6594
R6994 gnd.n293 gnd.n291 99.6594
R6995 gnd.n299 gnd.n211 99.6594
R6996 gnd.n303 gnd.n301 99.6594
R6997 gnd.n309 gnd.n207 99.6594
R6998 gnd.n313 gnd.n311 99.6594
R6999 gnd.n319 gnd.n203 99.6594
R7000 gnd.n323 gnd.n321 99.6594
R7001 gnd.n329 gnd.n199 99.6594
R7002 gnd.n333 gnd.n331 99.6594
R7003 gnd.n339 gnd.n193 99.6594
R7004 gnd.n343 gnd.n341 99.6594
R7005 gnd.n349 gnd.n189 99.6594
R7006 gnd.n353 gnd.n351 99.6594
R7007 gnd.n359 gnd.n185 99.6594
R7008 gnd.n363 gnd.n361 99.6594
R7009 gnd.n369 gnd.n181 99.6594
R7010 gnd.n373 gnd.n371 99.6594
R7011 gnd.n379 gnd.n177 99.6594
R7012 gnd.n382 gnd.n381 99.6594
R7013 gnd.n5514 gnd.n1611 99.6594
R7014 gnd.n5518 gnd.n5517 99.6594
R7015 gnd.n5525 gnd.n5524 99.6594
R7016 gnd.n5528 gnd.n5527 99.6594
R7017 gnd.n5535 gnd.n5534 99.6594
R7018 gnd.n5538 gnd.n5537 99.6594
R7019 gnd.n5545 gnd.n5544 99.6594
R7020 gnd.n5548 gnd.n5547 99.6594
R7021 gnd.n5558 gnd.n5557 99.6594
R7022 gnd.n5561 gnd.n5560 99.6594
R7023 gnd.n5568 gnd.n5567 99.6594
R7024 gnd.n5571 gnd.n5570 99.6594
R7025 gnd.n5579 gnd.n5578 99.6594
R7026 gnd.n5584 gnd.n5583 99.6594
R7027 gnd.n5591 gnd.n5590 99.6594
R7028 gnd.n5594 gnd.n5593 99.6594
R7029 gnd.n5601 gnd.n5600 99.6594
R7030 gnd.n5604 gnd.n5603 99.6594
R7031 gnd.n5613 gnd.n5612 99.6594
R7032 gnd.n5616 gnd.n5615 99.6594
R7033 gnd.n5623 gnd.n5622 99.6594
R7034 gnd.n5626 gnd.n5625 99.6594
R7035 gnd.n5633 gnd.n5632 99.6594
R7036 gnd.n5636 gnd.n5635 99.6594
R7037 gnd.n5643 gnd.n5642 99.6594
R7038 gnd.n5646 gnd.n5645 99.6594
R7039 gnd.n5654 gnd.n5653 99.6594
R7040 gnd.n5657 gnd.n5656 99.6594
R7041 gnd.n6115 gnd.n6114 99.6594
R7042 gnd.n6110 gnd.n1285 99.6594
R7043 gnd.n6106 gnd.n1284 99.6594
R7044 gnd.n6102 gnd.n1283 99.6594
R7045 gnd.n6098 gnd.n1282 99.6594
R7046 gnd.n6094 gnd.n1281 99.6594
R7047 gnd.n6090 gnd.n1280 99.6594
R7048 gnd.n6086 gnd.n1279 99.6594
R7049 gnd.n6081 gnd.n1278 99.6594
R7050 gnd.n6077 gnd.n1277 99.6594
R7051 gnd.n6073 gnd.n1276 99.6594
R7052 gnd.n6069 gnd.n1275 99.6594
R7053 gnd.n1411 gnd.n1273 99.6594
R7054 gnd.n1409 gnd.n1272 99.6594
R7055 gnd.n1405 gnd.n1271 99.6594
R7056 gnd.n1401 gnd.n1270 99.6594
R7057 gnd.n1397 gnd.n1269 99.6594
R7058 gnd.n1389 gnd.n1268 99.6594
R7059 gnd.n1387 gnd.n1267 99.6594
R7060 gnd.n1383 gnd.n1266 99.6594
R7061 gnd.n1379 gnd.n1265 99.6594
R7062 gnd.n1375 gnd.n1264 99.6594
R7063 gnd.n1371 gnd.n1263 99.6594
R7064 gnd.n1367 gnd.n1262 99.6594
R7065 gnd.n1363 gnd.n1261 99.6594
R7066 gnd.n1359 gnd.n1260 99.6594
R7067 gnd.n1355 gnd.n1259 99.6594
R7068 gnd.n1347 gnd.n1258 99.6594
R7069 gnd.n4213 gnd.n4212 99.6594
R7070 gnd.n3950 gnd.n3912 99.6594
R7071 gnd.n4205 gnd.n3913 99.6594
R7072 gnd.n4201 gnd.n3914 99.6594
R7073 gnd.n4197 gnd.n3915 99.6594
R7074 gnd.n4193 gnd.n3916 99.6594
R7075 gnd.n4189 gnd.n3917 99.6594
R7076 gnd.n4185 gnd.n3918 99.6594
R7077 gnd.n4181 gnd.n3919 99.6594
R7078 gnd.n4176 gnd.n3920 99.6594
R7079 gnd.n4172 gnd.n3921 99.6594
R7080 gnd.n4168 gnd.n3922 99.6594
R7081 gnd.n4164 gnd.n3923 99.6594
R7082 gnd.n4160 gnd.n3924 99.6594
R7083 gnd.n4156 gnd.n3925 99.6594
R7084 gnd.n4152 gnd.n3926 99.6594
R7085 gnd.n4148 gnd.n3927 99.6594
R7086 gnd.n4144 gnd.n3928 99.6594
R7087 gnd.n4140 gnd.n3929 99.6594
R7088 gnd.n4136 gnd.n3930 99.6594
R7089 gnd.n4132 gnd.n3931 99.6594
R7090 gnd.n4128 gnd.n3932 99.6594
R7091 gnd.n4124 gnd.n3933 99.6594
R7092 gnd.n4120 gnd.n3934 99.6594
R7093 gnd.n4116 gnd.n3935 99.6594
R7094 gnd.n4112 gnd.n3936 99.6594
R7095 gnd.n4108 gnd.n3937 99.6594
R7096 gnd.n4104 gnd.n3938 99.6594
R7097 gnd.n4100 gnd.n3939 99.6594
R7098 gnd.n3902 gnd.n2472 99.6594
R7099 gnd.n3900 gnd.n2471 99.6594
R7100 gnd.n3896 gnd.n2470 99.6594
R7101 gnd.n3892 gnd.n2469 99.6594
R7102 gnd.n3888 gnd.n2468 99.6594
R7103 gnd.n3884 gnd.n2467 99.6594
R7104 gnd.n3880 gnd.n2466 99.6594
R7105 gnd.n3812 gnd.n2465 99.6594
R7106 gnd.n3143 gnd.n2874 99.6594
R7107 gnd.n2900 gnd.n2881 99.6594
R7108 gnd.n2902 gnd.n2882 99.6594
R7109 gnd.n2910 gnd.n2883 99.6594
R7110 gnd.n2912 gnd.n2884 99.6594
R7111 gnd.n2920 gnd.n2885 99.6594
R7112 gnd.n2922 gnd.n2886 99.6594
R7113 gnd.n2930 gnd.n2887 99.6594
R7114 gnd.n7211 gnd.n7209 99.6594
R7115 gnd.n7217 gnd.n7202 99.6594
R7116 gnd.n7221 gnd.n7219 99.6594
R7117 gnd.n7227 gnd.n7198 99.6594
R7118 gnd.n7231 gnd.n7229 99.6594
R7119 gnd.n7237 gnd.n7194 99.6594
R7120 gnd.n7241 gnd.n7239 99.6594
R7121 gnd.n7247 gnd.n7190 99.6594
R7122 gnd.n7250 gnd.n7249 99.6594
R7123 gnd.n5206 gnd.n5205 99.6594
R7124 gnd.n5222 gnd.n5221 99.6594
R7125 gnd.n5225 gnd.n5224 99.6594
R7126 gnd.n5241 gnd.n5240 99.6594
R7127 gnd.n5244 gnd.n5243 99.6594
R7128 gnd.n5260 gnd.n5259 99.6594
R7129 gnd.n5263 gnd.n5262 99.6594
R7130 gnd.n5280 gnd.n5279 99.6594
R7131 gnd.n5283 gnd.n5282 99.6594
R7132 gnd.n3870 gnd.n2452 99.6594
R7133 gnd.n3866 gnd.n2453 99.6594
R7134 gnd.n3862 gnd.n2454 99.6594
R7135 gnd.n3858 gnd.n2455 99.6594
R7136 gnd.n3854 gnd.n2456 99.6594
R7137 gnd.n3850 gnd.n2457 99.6594
R7138 gnd.n3846 gnd.n2458 99.6594
R7139 gnd.n3842 gnd.n2459 99.6594
R7140 gnd.n3838 gnd.n2460 99.6594
R7141 gnd.n3834 gnd.n2461 99.6594
R7142 gnd.n3830 gnd.n2462 99.6594
R7143 gnd.n3826 gnd.n2463 99.6594
R7144 gnd.n3822 gnd.n2464 99.6594
R7145 gnd.n3058 gnd.n3057 99.6594
R7146 gnd.n3052 gnd.n2969 99.6594
R7147 gnd.n3049 gnd.n2970 99.6594
R7148 gnd.n3045 gnd.n2971 99.6594
R7149 gnd.n3041 gnd.n2972 99.6594
R7150 gnd.n3037 gnd.n2973 99.6594
R7151 gnd.n3033 gnd.n2974 99.6594
R7152 gnd.n3029 gnd.n2975 99.6594
R7153 gnd.n3025 gnd.n2976 99.6594
R7154 gnd.n3021 gnd.n2977 99.6594
R7155 gnd.n3017 gnd.n2978 99.6594
R7156 gnd.n3013 gnd.n2979 99.6594
R7157 gnd.n3060 gnd.n2968 99.6594
R7158 gnd.n1244 gnd.n1189 99.6594
R7159 gnd.n1246 gnd.n1198 99.6594
R7160 gnd.n1248 gnd.n1247 99.6594
R7161 gnd.n1249 gnd.n1207 99.6594
R7162 gnd.n1251 gnd.n1216 99.6594
R7163 gnd.n1253 gnd.n1252 99.6594
R7164 gnd.n1254 gnd.n1225 99.6594
R7165 gnd.n1256 gnd.n1237 99.6594
R7166 gnd.n6118 gnd.n6117 99.6594
R7167 gnd.n4089 gnd.n3940 99.6594
R7168 gnd.n4085 gnd.n3941 99.6594
R7169 gnd.n4081 gnd.n3942 99.6594
R7170 gnd.n4077 gnd.n3943 99.6594
R7171 gnd.n4073 gnd.n3944 99.6594
R7172 gnd.n4069 gnd.n3945 99.6594
R7173 gnd.n4065 gnd.n3946 99.6594
R7174 gnd.n4061 gnd.n3947 99.6594
R7175 gnd.n4057 gnd.n3948 99.6594
R7176 gnd.n4086 gnd.n3940 99.6594
R7177 gnd.n4082 gnd.n3941 99.6594
R7178 gnd.n4078 gnd.n3942 99.6594
R7179 gnd.n4074 gnd.n3943 99.6594
R7180 gnd.n4070 gnd.n3944 99.6594
R7181 gnd.n4066 gnd.n3945 99.6594
R7182 gnd.n4062 gnd.n3946 99.6594
R7183 gnd.n4058 gnd.n3947 99.6594
R7184 gnd.n4030 gnd.n3948 99.6594
R7185 gnd.n6117 gnd.n1242 99.6594
R7186 gnd.n1256 gnd.n1255 99.6594
R7187 gnd.n1254 gnd.n1224 99.6594
R7188 gnd.n1253 gnd.n1217 99.6594
R7189 gnd.n1251 gnd.n1250 99.6594
R7190 gnd.n1249 gnd.n1206 99.6594
R7191 gnd.n1248 gnd.n1199 99.6594
R7192 gnd.n1246 gnd.n1245 99.6594
R7193 gnd.n1244 gnd.n1188 99.6594
R7194 gnd.n3058 gnd.n2981 99.6594
R7195 gnd.n3050 gnd.n2969 99.6594
R7196 gnd.n3046 gnd.n2970 99.6594
R7197 gnd.n3042 gnd.n2971 99.6594
R7198 gnd.n3038 gnd.n2972 99.6594
R7199 gnd.n3034 gnd.n2973 99.6594
R7200 gnd.n3030 gnd.n2974 99.6594
R7201 gnd.n3026 gnd.n2975 99.6594
R7202 gnd.n3022 gnd.n2976 99.6594
R7203 gnd.n3018 gnd.n2977 99.6594
R7204 gnd.n3014 gnd.n2978 99.6594
R7205 gnd.n3010 gnd.n2979 99.6594
R7206 gnd.n3061 gnd.n3060 99.6594
R7207 gnd.n3825 gnd.n2464 99.6594
R7208 gnd.n3829 gnd.n2463 99.6594
R7209 gnd.n3833 gnd.n2462 99.6594
R7210 gnd.n3837 gnd.n2461 99.6594
R7211 gnd.n3841 gnd.n2460 99.6594
R7212 gnd.n3845 gnd.n2459 99.6594
R7213 gnd.n3849 gnd.n2458 99.6594
R7214 gnd.n3853 gnd.n2457 99.6594
R7215 gnd.n3857 gnd.n2456 99.6594
R7216 gnd.n3861 gnd.n2455 99.6594
R7217 gnd.n3865 gnd.n2454 99.6594
R7218 gnd.n3869 gnd.n2453 99.6594
R7219 gnd.n2493 gnd.n2452 99.6594
R7220 gnd.n5205 gnd.n5170 99.6594
R7221 gnd.n5223 gnd.n5222 99.6594
R7222 gnd.n5224 gnd.n5161 99.6594
R7223 gnd.n5242 gnd.n5241 99.6594
R7224 gnd.n5243 gnd.n5152 99.6594
R7225 gnd.n5261 gnd.n5260 99.6594
R7226 gnd.n5262 gnd.n5143 99.6594
R7227 gnd.n5281 gnd.n5280 99.6594
R7228 gnd.n5282 gnd.n5139 99.6594
R7229 gnd.n7249 gnd.n7248 99.6594
R7230 gnd.n7240 gnd.n7190 99.6594
R7231 gnd.n7239 gnd.n7238 99.6594
R7232 gnd.n7230 gnd.n7194 99.6594
R7233 gnd.n7229 gnd.n7228 99.6594
R7234 gnd.n7220 gnd.n7198 99.6594
R7235 gnd.n7219 gnd.n7218 99.6594
R7236 gnd.n7210 gnd.n7202 99.6594
R7237 gnd.n7209 gnd.n7208 99.6594
R7238 gnd.n3144 gnd.n3143 99.6594
R7239 gnd.n2903 gnd.n2881 99.6594
R7240 gnd.n2909 gnd.n2882 99.6594
R7241 gnd.n2913 gnd.n2883 99.6594
R7242 gnd.n2919 gnd.n2884 99.6594
R7243 gnd.n2923 gnd.n2885 99.6594
R7244 gnd.n2929 gnd.n2886 99.6594
R7245 gnd.n2887 gnd.n2871 99.6594
R7246 gnd.n3879 gnd.n2465 99.6594
R7247 gnd.n3883 gnd.n2466 99.6594
R7248 gnd.n3887 gnd.n2467 99.6594
R7249 gnd.n3891 gnd.n2468 99.6594
R7250 gnd.n3895 gnd.n2469 99.6594
R7251 gnd.n3899 gnd.n2470 99.6594
R7252 gnd.n3903 gnd.n2471 99.6594
R7253 gnd.n2474 gnd.n2472 99.6594
R7254 gnd.n4212 gnd.n2449 99.6594
R7255 gnd.n4206 gnd.n3912 99.6594
R7256 gnd.n4202 gnd.n3913 99.6594
R7257 gnd.n4198 gnd.n3914 99.6594
R7258 gnd.n4194 gnd.n3915 99.6594
R7259 gnd.n4190 gnd.n3916 99.6594
R7260 gnd.n4186 gnd.n3917 99.6594
R7261 gnd.n4182 gnd.n3918 99.6594
R7262 gnd.n4177 gnd.n3919 99.6594
R7263 gnd.n4173 gnd.n3920 99.6594
R7264 gnd.n4169 gnd.n3921 99.6594
R7265 gnd.n4165 gnd.n3922 99.6594
R7266 gnd.n4161 gnd.n3923 99.6594
R7267 gnd.n4157 gnd.n3924 99.6594
R7268 gnd.n4153 gnd.n3925 99.6594
R7269 gnd.n4149 gnd.n3926 99.6594
R7270 gnd.n4145 gnd.n3927 99.6594
R7271 gnd.n4141 gnd.n3928 99.6594
R7272 gnd.n4137 gnd.n3929 99.6594
R7273 gnd.n4133 gnd.n3930 99.6594
R7274 gnd.n4129 gnd.n3931 99.6594
R7275 gnd.n4125 gnd.n3932 99.6594
R7276 gnd.n4121 gnd.n3933 99.6594
R7277 gnd.n4117 gnd.n3934 99.6594
R7278 gnd.n4113 gnd.n3935 99.6594
R7279 gnd.n4109 gnd.n3936 99.6594
R7280 gnd.n4105 gnd.n3937 99.6594
R7281 gnd.n4101 gnd.n3938 99.6594
R7282 gnd.n4010 gnd.n3939 99.6594
R7283 gnd.n1354 gnd.n1258 99.6594
R7284 gnd.n1358 gnd.n1259 99.6594
R7285 gnd.n1362 gnd.n1260 99.6594
R7286 gnd.n1366 gnd.n1261 99.6594
R7287 gnd.n1370 gnd.n1262 99.6594
R7288 gnd.n1374 gnd.n1263 99.6594
R7289 gnd.n1378 gnd.n1264 99.6594
R7290 gnd.n1382 gnd.n1265 99.6594
R7291 gnd.n1386 gnd.n1266 99.6594
R7292 gnd.n1390 gnd.n1267 99.6594
R7293 gnd.n1396 gnd.n1268 99.6594
R7294 gnd.n1400 gnd.n1269 99.6594
R7295 gnd.n1404 gnd.n1270 99.6594
R7296 gnd.n1408 gnd.n1271 99.6594
R7297 gnd.n1412 gnd.n1272 99.6594
R7298 gnd.n6068 gnd.n1274 99.6594
R7299 gnd.n6072 gnd.n1275 99.6594
R7300 gnd.n6076 gnd.n1276 99.6594
R7301 gnd.n6080 gnd.n1277 99.6594
R7302 gnd.n6085 gnd.n1278 99.6594
R7303 gnd.n6089 gnd.n1279 99.6594
R7304 gnd.n6093 gnd.n1280 99.6594
R7305 gnd.n6097 gnd.n1281 99.6594
R7306 gnd.n6101 gnd.n1282 99.6594
R7307 gnd.n6105 gnd.n1283 99.6594
R7308 gnd.n6109 gnd.n1284 99.6594
R7309 gnd.n1287 gnd.n1285 99.6594
R7310 gnd.n6115 gnd.n1286 99.6594
R7311 gnd.n5515 gnd.n5514 99.6594
R7312 gnd.n5517 gnd.n5506 99.6594
R7313 gnd.n5526 gnd.n5525 99.6594
R7314 gnd.n5527 gnd.n5502 99.6594
R7315 gnd.n5536 gnd.n5535 99.6594
R7316 gnd.n5537 gnd.n5498 99.6594
R7317 gnd.n5546 gnd.n5545 99.6594
R7318 gnd.n5547 gnd.n5494 99.6594
R7319 gnd.n5559 gnd.n5558 99.6594
R7320 gnd.n5560 gnd.n5490 99.6594
R7321 gnd.n5569 gnd.n5568 99.6594
R7322 gnd.n5570 gnd.n5486 99.6594
R7323 gnd.n5582 gnd.n5581 99.6594
R7324 gnd.n5583 gnd.n1783 99.6594
R7325 gnd.n5592 gnd.n5591 99.6594
R7326 gnd.n5593 gnd.n1779 99.6594
R7327 gnd.n5602 gnd.n5601 99.6594
R7328 gnd.n5603 gnd.n1775 99.6594
R7329 gnd.n5614 gnd.n5613 99.6594
R7330 gnd.n5615 gnd.n1771 99.6594
R7331 gnd.n5624 gnd.n5623 99.6594
R7332 gnd.n5625 gnd.n1767 99.6594
R7333 gnd.n5634 gnd.n5633 99.6594
R7334 gnd.n5635 gnd.n1763 99.6594
R7335 gnd.n5644 gnd.n5643 99.6594
R7336 gnd.n5645 gnd.n1759 99.6594
R7337 gnd.n5655 gnd.n5654 99.6594
R7338 gnd.n5658 gnd.n5657 99.6594
R7339 gnd.n381 gnd.n380 99.6594
R7340 gnd.n372 gnd.n177 99.6594
R7341 gnd.n371 gnd.n370 99.6594
R7342 gnd.n362 gnd.n181 99.6594
R7343 gnd.n361 gnd.n360 99.6594
R7344 gnd.n352 gnd.n185 99.6594
R7345 gnd.n351 gnd.n350 99.6594
R7346 gnd.n342 gnd.n189 99.6594
R7347 gnd.n341 gnd.n340 99.6594
R7348 gnd.n332 gnd.n193 99.6594
R7349 gnd.n331 gnd.n330 99.6594
R7350 gnd.n322 gnd.n199 99.6594
R7351 gnd.n321 gnd.n320 99.6594
R7352 gnd.n312 gnd.n203 99.6594
R7353 gnd.n311 gnd.n310 99.6594
R7354 gnd.n302 gnd.n207 99.6594
R7355 gnd.n301 gnd.n300 99.6594
R7356 gnd.n292 gnd.n211 99.6594
R7357 gnd.n291 gnd.n290 99.6594
R7358 gnd.n282 gnd.n215 99.6594
R7359 gnd.n281 gnd.n280 99.6594
R7360 gnd.n272 gnd.n271 99.6594
R7361 gnd.n270 gnd.n269 99.6594
R7362 gnd.n261 gnd.n225 99.6594
R7363 gnd.n260 gnd.n259 99.6594
R7364 gnd.n251 gnd.n229 99.6594
R7365 gnd.n250 gnd.n249 99.6594
R7366 gnd.n241 gnd.n233 99.6594
R7367 gnd.n240 gnd.n239 99.6594
R7368 gnd.n6180 gnd.n6179 99.6594
R7369 gnd.n1175 gnd.n1155 99.6594
R7370 gnd.n1177 gnd.n1156 99.6594
R7371 gnd.n1181 gnd.n1157 99.6594
R7372 gnd.n1183 gnd.n1158 99.6594
R7373 gnd.n1193 gnd.n1159 99.6594
R7374 gnd.n1195 gnd.n1160 99.6594
R7375 gnd.n1203 gnd.n1161 99.6594
R7376 gnd.n1211 gnd.n1162 99.6594
R7377 gnd.n1213 gnd.n1163 99.6594
R7378 gnd.n1221 gnd.n1164 99.6594
R7379 gnd.n1229 gnd.n1165 99.6594
R7380 gnd.n1234 gnd.n1167 99.6594
R7381 gnd.n6182 gnd.n1152 99.6594
R7382 gnd.n6180 gnd.n1170 99.6594
R7383 gnd.n1176 gnd.n1155 99.6594
R7384 gnd.n1180 gnd.n1156 99.6594
R7385 gnd.n1182 gnd.n1157 99.6594
R7386 gnd.n1192 gnd.n1158 99.6594
R7387 gnd.n1194 gnd.n1159 99.6594
R7388 gnd.n1202 gnd.n1160 99.6594
R7389 gnd.n1210 gnd.n1161 99.6594
R7390 gnd.n1212 gnd.n1162 99.6594
R7391 gnd.n1220 gnd.n1163 99.6594
R7392 gnd.n1228 gnd.n1164 99.6594
R7393 gnd.n1230 gnd.n1165 99.6594
R7394 gnd.n1167 gnd.n1166 99.6594
R7395 gnd.n6183 gnd.n6182 99.6594
R7396 gnd.n5186 gnd.n5182 99.6594
R7397 gnd.n5190 gnd.n5188 99.6594
R7398 gnd.n5197 gnd.n5178 99.6594
R7399 gnd.n5201 gnd.n5199 99.6594
R7400 gnd.n5212 gnd.n5175 99.6594
R7401 gnd.n5216 gnd.n5214 99.6594
R7402 gnd.n5231 gnd.n5166 99.6594
R7403 gnd.n5235 gnd.n5233 99.6594
R7404 gnd.n5250 gnd.n5157 99.6594
R7405 gnd.n5254 gnd.n5252 99.6594
R7406 gnd.n5269 gnd.n5148 99.6594
R7407 gnd.n5272 gnd.n5271 99.6594
R7408 gnd.n5290 gnd.n5289 99.6594
R7409 gnd.n5293 gnd.n5292 99.6594
R7410 gnd.n5271 gnd.n5270 99.6594
R7411 gnd.n5253 gnd.n5148 99.6594
R7412 gnd.n5252 gnd.n5251 99.6594
R7413 gnd.n5234 gnd.n5157 99.6594
R7414 gnd.n5233 gnd.n5232 99.6594
R7415 gnd.n5215 gnd.n5166 99.6594
R7416 gnd.n5214 gnd.n5213 99.6594
R7417 gnd.n5200 gnd.n5175 99.6594
R7418 gnd.n5199 gnd.n5198 99.6594
R7419 gnd.n5189 gnd.n5178 99.6594
R7420 gnd.n5188 gnd.n5187 99.6594
R7421 gnd.n5182 gnd.n1585 99.6594
R7422 gnd.n5294 gnd.n5293 99.6594
R7423 gnd.n5291 gnd.n5290 99.6594
R7424 gnd.n1231 gnd.t75 98.63
R7425 gnd.n5140 gnd.t101 98.63
R7426 gnd.n1238 gnd.t122 98.63
R7427 gnd.n5553 gnd.t98 98.63
R7428 gnd.n5605 gnd.t88 98.63
R7429 gnd.n1755 gnd.t28 98.63
R7430 gnd.n174 gnd.t37 98.63
R7431 gnd.n196 gnd.t23 98.63
R7432 gnd.n218 gnd.t90 98.63
R7433 gnd.n7187 gnd.t115 98.63
R7434 gnd.n3967 gnd.t58 98.63
R7435 gnd.n3989 gnd.t44 98.63
R7436 gnd.n4012 gnd.t68 98.63
R7437 gnd.n4031 gnd.t20 98.63
R7438 gnd.n1308 gnd.t112 98.63
R7439 gnd.n1349 gnd.t47 98.63
R7440 gnd.n1328 gnd.t70 98.63
R7441 gnd.n5130 gnd.t51 98.63
R7442 gnd.n2205 gnd.t82 92.8196
R7443 gnd.n1824 gnd.t106 92.8196
R7444 gnd.n5997 gnd.t133 92.8118
R7445 gnd.n5347 gnd.t34 92.8118
R7446 gnd.n1466 gnd.n1465 81.8399
R7447 gnd.n5485 gnd.n5484 78.9125
R7448 gnd.n6066 gnd.n6065 78.9125
R7449 gnd.n2932 gnd.t61 74.8376
R7450 gnd.n2490 gnd.t95 74.8376
R7451 gnd.n2206 gnd.t81 72.8438
R7452 gnd.n1825 gnd.t107 72.8438
R7453 gnd.n1467 gnd.n1460 72.8411
R7454 gnd.n1473 gnd.n1458 72.8411
R7455 gnd.n5343 gnd.n5342 72.8411
R7456 gnd.n1232 gnd.t74 72.836
R7457 gnd.n5998 gnd.t132 72.836
R7458 gnd.n5348 gnd.t35 72.836
R7459 gnd.n5141 gnd.t100 72.836
R7460 gnd.n1239 gnd.t123 72.836
R7461 gnd.n5554 gnd.t97 72.836
R7462 gnd.n5606 gnd.t87 72.836
R7463 gnd.n1756 gnd.t27 72.836
R7464 gnd.n175 gnd.t38 72.836
R7465 gnd.n197 gnd.t24 72.836
R7466 gnd.n219 gnd.t91 72.836
R7467 gnd.n7188 gnd.t116 72.836
R7468 gnd.n3968 gnd.t57 72.836
R7469 gnd.n3990 gnd.t43 72.836
R7470 gnd.n4013 gnd.t67 72.836
R7471 gnd.n4032 gnd.t19 72.836
R7472 gnd.n1309 gnd.t113 72.836
R7473 gnd.n1350 gnd.t48 72.836
R7474 gnd.n1329 gnd.t71 72.836
R7475 gnd.n5131 gnd.t52 72.836
R7476 gnd.n5408 gnd.n1792 71.676
R7477 gnd.n5404 gnd.n1793 71.676
R7478 gnd.n5400 gnd.n1794 71.676
R7479 gnd.n5396 gnd.n1795 71.676
R7480 gnd.n5392 gnd.n1796 71.676
R7481 gnd.n5388 gnd.n1797 71.676
R7482 gnd.n5384 gnd.n1798 71.676
R7483 gnd.n5380 gnd.n1799 71.676
R7484 gnd.n5376 gnd.n1800 71.676
R7485 gnd.n5372 gnd.n1801 71.676
R7486 gnd.n5368 gnd.n1802 71.676
R7487 gnd.n5364 gnd.n1803 71.676
R7488 gnd.n5360 gnd.n1804 71.676
R7489 gnd.n5356 gnd.n1805 71.676
R7490 gnd.n5351 gnd.n1806 71.676
R7491 gnd.n1807 gnd.n1790 71.676
R7492 gnd.n5480 gnd.n1789 71.676
R7493 gnd.n5478 gnd.n5477 71.676
R7494 gnd.n5472 gnd.n1822 71.676
R7495 gnd.n5468 gnd.n1821 71.676
R7496 gnd.n5464 gnd.n1820 71.676
R7497 gnd.n5460 gnd.n1819 71.676
R7498 gnd.n5456 gnd.n1818 71.676
R7499 gnd.n5452 gnd.n1817 71.676
R7500 gnd.n5448 gnd.n1816 71.676
R7501 gnd.n5444 gnd.n1815 71.676
R7502 gnd.n5440 gnd.n1814 71.676
R7503 gnd.n5436 gnd.n1813 71.676
R7504 gnd.n5432 gnd.n1812 71.676
R7505 gnd.n5428 gnd.n1811 71.676
R7506 gnd.n5424 gnd.n1810 71.676
R7507 gnd.n5420 gnd.n1809 71.676
R7508 gnd.n5416 gnd.n1808 71.676
R7509 gnd.n6061 gnd.n6060 71.676
R7510 gnd.n6055 gnd.n1422 71.676
R7511 gnd.n6052 gnd.n1423 71.676
R7512 gnd.n6048 gnd.n1424 71.676
R7513 gnd.n6044 gnd.n1425 71.676
R7514 gnd.n6040 gnd.n1426 71.676
R7515 gnd.n6036 gnd.n1427 71.676
R7516 gnd.n6032 gnd.n1428 71.676
R7517 gnd.n6028 gnd.n1429 71.676
R7518 gnd.n6024 gnd.n1430 71.676
R7519 gnd.n6020 gnd.n1431 71.676
R7520 gnd.n6016 gnd.n1432 71.676
R7521 gnd.n6012 gnd.n1433 71.676
R7522 gnd.n6008 gnd.n1434 71.676
R7523 gnd.n6004 gnd.n1435 71.676
R7524 gnd.n6000 gnd.n1436 71.676
R7525 gnd.n1437 gnd.n1420 71.676
R7526 gnd.n2209 gnd.n1438 71.676
R7527 gnd.n2214 gnd.n1439 71.676
R7528 gnd.n2218 gnd.n1440 71.676
R7529 gnd.n2222 gnd.n1441 71.676
R7530 gnd.n2226 gnd.n1442 71.676
R7531 gnd.n2230 gnd.n1443 71.676
R7532 gnd.n2234 gnd.n1444 71.676
R7533 gnd.n2238 gnd.n1445 71.676
R7534 gnd.n2242 gnd.n1446 71.676
R7535 gnd.n2246 gnd.n1447 71.676
R7536 gnd.n2250 gnd.n1448 71.676
R7537 gnd.n2254 gnd.n1449 71.676
R7538 gnd.n2258 gnd.n1450 71.676
R7539 gnd.n2262 gnd.n1451 71.676
R7540 gnd.n2266 gnd.n1452 71.676
R7541 gnd.n6061 gnd.n1455 71.676
R7542 gnd.n6053 gnd.n1422 71.676
R7543 gnd.n6049 gnd.n1423 71.676
R7544 gnd.n6045 gnd.n1424 71.676
R7545 gnd.n6041 gnd.n1425 71.676
R7546 gnd.n6037 gnd.n1426 71.676
R7547 gnd.n6033 gnd.n1427 71.676
R7548 gnd.n6029 gnd.n1428 71.676
R7549 gnd.n6025 gnd.n1429 71.676
R7550 gnd.n6021 gnd.n1430 71.676
R7551 gnd.n6017 gnd.n1431 71.676
R7552 gnd.n6013 gnd.n1432 71.676
R7553 gnd.n6009 gnd.n1433 71.676
R7554 gnd.n6005 gnd.n1434 71.676
R7555 gnd.n6001 gnd.n1435 71.676
R7556 gnd.n6064 gnd.n6063 71.676
R7557 gnd.n2208 gnd.n1437 71.676
R7558 gnd.n2213 gnd.n1438 71.676
R7559 gnd.n2217 gnd.n1439 71.676
R7560 gnd.n2221 gnd.n1440 71.676
R7561 gnd.n2225 gnd.n1441 71.676
R7562 gnd.n2229 gnd.n1442 71.676
R7563 gnd.n2233 gnd.n1443 71.676
R7564 gnd.n2237 gnd.n1444 71.676
R7565 gnd.n2241 gnd.n1445 71.676
R7566 gnd.n2245 gnd.n1446 71.676
R7567 gnd.n2249 gnd.n1447 71.676
R7568 gnd.n2253 gnd.n1448 71.676
R7569 gnd.n2257 gnd.n1449 71.676
R7570 gnd.n2261 gnd.n1450 71.676
R7571 gnd.n2265 gnd.n1451 71.676
R7572 gnd.n2204 gnd.n1452 71.676
R7573 gnd.n5419 gnd.n1808 71.676
R7574 gnd.n5423 gnd.n1809 71.676
R7575 gnd.n5427 gnd.n1810 71.676
R7576 gnd.n5431 gnd.n1811 71.676
R7577 gnd.n5435 gnd.n1812 71.676
R7578 gnd.n5439 gnd.n1813 71.676
R7579 gnd.n5443 gnd.n1814 71.676
R7580 gnd.n5447 gnd.n1815 71.676
R7581 gnd.n5451 gnd.n1816 71.676
R7582 gnd.n5455 gnd.n1817 71.676
R7583 gnd.n5459 gnd.n1818 71.676
R7584 gnd.n5463 gnd.n1819 71.676
R7585 gnd.n5467 gnd.n1820 71.676
R7586 gnd.n5471 gnd.n1821 71.676
R7587 gnd.n1823 gnd.n1822 71.676
R7588 gnd.n5479 gnd.n5478 71.676
R7589 gnd.n5483 gnd.n5482 71.676
R7590 gnd.n5350 gnd.n1807 71.676
R7591 gnd.n5355 gnd.n1806 71.676
R7592 gnd.n5359 gnd.n1805 71.676
R7593 gnd.n5363 gnd.n1804 71.676
R7594 gnd.n5367 gnd.n1803 71.676
R7595 gnd.n5371 gnd.n1802 71.676
R7596 gnd.n5375 gnd.n1801 71.676
R7597 gnd.n5379 gnd.n1800 71.676
R7598 gnd.n5383 gnd.n1799 71.676
R7599 gnd.n5387 gnd.n1798 71.676
R7600 gnd.n5391 gnd.n1797 71.676
R7601 gnd.n5395 gnd.n1796 71.676
R7602 gnd.n5399 gnd.n1795 71.676
R7603 gnd.n5403 gnd.n1794 71.676
R7604 gnd.n5407 gnd.n1793 71.676
R7605 gnd.n1830 gnd.n1792 71.676
R7606 gnd.n8 gnd.t223 69.1507
R7607 gnd.n14 gnd.t313 68.4792
R7608 gnd.n13 gnd.t230 68.4792
R7609 gnd.n12 gnd.t300 68.4792
R7610 gnd.n11 gnd.t320 68.4792
R7611 gnd.n10 gnd.t264 68.4792
R7612 gnd.n9 gnd.t148 68.4792
R7613 gnd.n8 gnd.t278 68.4792
R7614 gnd.n3059 gnd.n2963 64.369
R7615 gnd.n4211 gnd.n2442 63.0944
R7616 gnd.n7283 gnd.n170 63.0944
R7617 gnd.n2211 gnd.n2206 59.5399
R7618 gnd.n5474 gnd.n1825 59.5399
R7619 gnd.n5999 gnd.n5998 59.5399
R7620 gnd.n5353 gnd.n5348 59.5399
R7621 gnd.n5996 gnd.n1476 59.1804
R7622 gnd.n3911 gnd.n2450 57.3586
R7623 gnd.n2718 gnd.t244 56.407
R7624 gnd.n2683 gnd.t268 56.407
R7625 gnd.n2694 gnd.t137 56.407
R7626 gnd.n2706 gnd.t161 56.407
R7627 gnd.n52 gnd.t152 56.407
R7628 gnd.n17 gnd.t171 56.407
R7629 gnd.n28 gnd.t195 56.407
R7630 gnd.n40 gnd.t303 56.407
R7631 gnd.n2727 gnd.t209 55.8337
R7632 gnd.n2692 gnd.t170 55.8337
R7633 gnd.n2703 gnd.t274 55.8337
R7634 gnd.n2715 gnd.t205 55.8337
R7635 gnd.n61 gnd.t164 55.8337
R7636 gnd.n26 gnd.t254 55.8337
R7637 gnd.n37 gnd.t7 55.8337
R7638 gnd.n49 gnd.t315 55.8337
R7639 gnd.n1464 gnd.n1463 54.358
R7640 gnd.n5340 gnd.n5339 54.358
R7641 gnd.n2718 gnd.n2717 53.0052
R7642 gnd.n2720 gnd.n2719 53.0052
R7643 gnd.n2722 gnd.n2721 53.0052
R7644 gnd.n2724 gnd.n2723 53.0052
R7645 gnd.n2726 gnd.n2725 53.0052
R7646 gnd.n2683 gnd.n2682 53.0052
R7647 gnd.n2685 gnd.n2684 53.0052
R7648 gnd.n2687 gnd.n2686 53.0052
R7649 gnd.n2689 gnd.n2688 53.0052
R7650 gnd.n2691 gnd.n2690 53.0052
R7651 gnd.n2694 gnd.n2693 53.0052
R7652 gnd.n2696 gnd.n2695 53.0052
R7653 gnd.n2698 gnd.n2697 53.0052
R7654 gnd.n2700 gnd.n2699 53.0052
R7655 gnd.n2702 gnd.n2701 53.0052
R7656 gnd.n2706 gnd.n2705 53.0052
R7657 gnd.n2708 gnd.n2707 53.0052
R7658 gnd.n2710 gnd.n2709 53.0052
R7659 gnd.n2712 gnd.n2711 53.0052
R7660 gnd.n2714 gnd.n2713 53.0052
R7661 gnd.n60 gnd.n59 53.0052
R7662 gnd.n58 gnd.n57 53.0052
R7663 gnd.n56 gnd.n55 53.0052
R7664 gnd.n54 gnd.n53 53.0052
R7665 gnd.n52 gnd.n51 53.0052
R7666 gnd.n25 gnd.n24 53.0052
R7667 gnd.n23 gnd.n22 53.0052
R7668 gnd.n21 gnd.n20 53.0052
R7669 gnd.n19 gnd.n18 53.0052
R7670 gnd.n17 gnd.n16 53.0052
R7671 gnd.n36 gnd.n35 53.0052
R7672 gnd.n34 gnd.n33 53.0052
R7673 gnd.n32 gnd.n31 53.0052
R7674 gnd.n30 gnd.n29 53.0052
R7675 gnd.n28 gnd.n27 53.0052
R7676 gnd.n48 gnd.n47 53.0052
R7677 gnd.n46 gnd.n45 53.0052
R7678 gnd.n44 gnd.n43 53.0052
R7679 gnd.n42 gnd.n41 53.0052
R7680 gnd.n40 gnd.n39 53.0052
R7681 gnd.n5331 gnd.n5330 52.4801
R7682 gnd.n3763 gnd.t193 52.3082
R7683 gnd.n3731 gnd.t311 52.3082
R7684 gnd.n3699 gnd.t221 52.3082
R7685 gnd.n3668 gnd.t290 52.3082
R7686 gnd.n3636 gnd.t144 52.3082
R7687 gnd.n3604 gnd.t323 52.3082
R7688 gnd.n3572 gnd.t327 52.3082
R7689 gnd.n3541 gnd.t325 52.3082
R7690 gnd.n3593 gnd.n3561 51.4173
R7691 gnd.n3657 gnd.n3656 50.455
R7692 gnd.n3625 gnd.n3624 50.455
R7693 gnd.n3593 gnd.n3592 50.455
R7694 gnd.n3006 gnd.n3005 45.1884
R7695 gnd.n2516 gnd.n2515 45.1884
R7696 gnd.n5411 gnd.n5346 44.3322
R7697 gnd.n1467 gnd.n1466 44.3189
R7698 gnd.n1233 gnd.n1232 42.2793
R7699 gnd.n5285 gnd.n5141 42.2793
R7700 gnd.n3007 gnd.n3006 42.2793
R7701 gnd.n2517 gnd.n2516 42.2793
R7702 gnd.n2933 gnd.n2932 42.2793
R7703 gnd.n3878 gnd.n2490 42.2793
R7704 gnd.n6120 gnd.n1239 42.2793
R7705 gnd.n5555 gnd.n5554 42.2793
R7706 gnd.n5607 gnd.n5606 42.2793
R7707 gnd.n1757 gnd.n1756 42.2793
R7708 gnd.n176 gnd.n175 42.2793
R7709 gnd.n198 gnd.n197 42.2793
R7710 gnd.n220 gnd.n219 42.2793
R7711 gnd.n7189 gnd.n7188 42.2793
R7712 gnd.n4179 gnd.n3968 42.2793
R7713 gnd.n4139 gnd.n3990 42.2793
R7714 gnd.n4099 gnd.n4013 42.2793
R7715 gnd.n4033 gnd.n4032 42.2793
R7716 gnd.n6083 gnd.n1309 42.2793
R7717 gnd.n1353 gnd.n1350 42.2793
R7718 gnd.n1395 gnd.n1329 42.2793
R7719 gnd.n5132 gnd.n5131 42.2793
R7720 gnd.n1465 gnd.n1464 41.6274
R7721 gnd.n5341 gnd.n5340 41.6274
R7722 gnd.n6476 gnd.n795 41.1297
R7723 gnd.n6476 gnd.n6475 41.1297
R7724 gnd.n6475 gnd.n6474 41.1297
R7725 gnd.n6474 gnd.n800 41.1297
R7726 gnd.n6468 gnd.n800 41.1297
R7727 gnd.n6468 gnd.n6467 41.1297
R7728 gnd.n6467 gnd.n6466 41.1297
R7729 gnd.n6466 gnd.n808 41.1297
R7730 gnd.n6460 gnd.n808 41.1297
R7731 gnd.n6460 gnd.n6459 41.1297
R7732 gnd.n6459 gnd.n6458 41.1297
R7733 gnd.n6458 gnd.n816 41.1297
R7734 gnd.n6452 gnd.n816 41.1297
R7735 gnd.n6452 gnd.n6451 41.1297
R7736 gnd.n6451 gnd.n6450 41.1297
R7737 gnd.n6450 gnd.n824 41.1297
R7738 gnd.n6444 gnd.n824 41.1297
R7739 gnd.n6444 gnd.n6443 41.1297
R7740 gnd.n6443 gnd.n6442 41.1297
R7741 gnd.n6442 gnd.n832 41.1297
R7742 gnd.n6436 gnd.n832 41.1297
R7743 gnd.n6436 gnd.n6435 41.1297
R7744 gnd.n6435 gnd.n6434 41.1297
R7745 gnd.n6434 gnd.n840 41.1297
R7746 gnd.n6428 gnd.n840 41.1297
R7747 gnd.n6428 gnd.n6427 41.1297
R7748 gnd.n6427 gnd.n6426 41.1297
R7749 gnd.n6426 gnd.n848 41.1297
R7750 gnd.n6420 gnd.n848 41.1297
R7751 gnd.n6420 gnd.n6419 41.1297
R7752 gnd.n6419 gnd.n6418 41.1297
R7753 gnd.n6418 gnd.n856 41.1297
R7754 gnd.n6412 gnd.n856 41.1297
R7755 gnd.n6412 gnd.n6411 41.1297
R7756 gnd.n6411 gnd.n6410 41.1297
R7757 gnd.n6410 gnd.n864 41.1297
R7758 gnd.n6404 gnd.n864 41.1297
R7759 gnd.n6404 gnd.n6403 41.1297
R7760 gnd.n6403 gnd.n6402 41.1297
R7761 gnd.n6402 gnd.n872 41.1297
R7762 gnd.n6396 gnd.n872 41.1297
R7763 gnd.n6396 gnd.n6395 41.1297
R7764 gnd.n6395 gnd.n6394 41.1297
R7765 gnd.n6394 gnd.n880 41.1297
R7766 gnd.n6388 gnd.n880 41.1297
R7767 gnd.n6388 gnd.n6387 41.1297
R7768 gnd.n6387 gnd.n6386 41.1297
R7769 gnd.n6386 gnd.n888 41.1297
R7770 gnd.n6380 gnd.n888 41.1297
R7771 gnd.n6380 gnd.n6379 41.1297
R7772 gnd.n6379 gnd.n6378 41.1297
R7773 gnd.n6378 gnd.n896 41.1297
R7774 gnd.n6372 gnd.n896 41.1297
R7775 gnd.n6372 gnd.n6371 41.1297
R7776 gnd.n6371 gnd.n6370 41.1297
R7777 gnd.n6370 gnd.n904 41.1297
R7778 gnd.n6364 gnd.n904 41.1297
R7779 gnd.n6364 gnd.n6363 41.1297
R7780 gnd.n6363 gnd.n6362 41.1297
R7781 gnd.n6362 gnd.n912 41.1297
R7782 gnd.n6356 gnd.n912 41.1297
R7783 gnd.n6356 gnd.n6355 41.1297
R7784 gnd.n6355 gnd.n6354 41.1297
R7785 gnd.n6354 gnd.n920 41.1297
R7786 gnd.n6348 gnd.n920 41.1297
R7787 gnd.n6348 gnd.n6347 41.1297
R7788 gnd.n6347 gnd.n6346 41.1297
R7789 gnd.n6346 gnd.n928 41.1297
R7790 gnd.n6340 gnd.n928 41.1297
R7791 gnd.n6340 gnd.n6339 41.1297
R7792 gnd.n6339 gnd.n6338 41.1297
R7793 gnd.n6338 gnd.n936 41.1297
R7794 gnd.n6332 gnd.n936 41.1297
R7795 gnd.n6332 gnd.n6331 41.1297
R7796 gnd.n6331 gnd.n6330 41.1297
R7797 gnd.n6330 gnd.n944 41.1297
R7798 gnd.n6324 gnd.n944 41.1297
R7799 gnd.n6324 gnd.n6323 41.1297
R7800 gnd.n6323 gnd.n6322 41.1297
R7801 gnd.n6322 gnd.n952 41.1297
R7802 gnd.n6316 gnd.n952 41.1297
R7803 gnd.n6316 gnd.n6315 41.1297
R7804 gnd.n6315 gnd.n6314 41.1297
R7805 gnd.n1474 gnd.n1473 40.8975
R7806 gnd.n5344 gnd.n5343 40.8975
R7807 gnd.n1473 gnd.n1472 35.055
R7808 gnd.n1468 gnd.n1467 35.055
R7809 gnd.n5333 gnd.n5332 35.055
R7810 gnd.n5343 gnd.n5329 35.055
R7811 gnd.n3069 gnd.n2963 31.8661
R7812 gnd.n3069 gnd.n3068 31.8661
R7813 gnd.n3077 gnd.n2952 31.8661
R7814 gnd.n3085 gnd.n2952 31.8661
R7815 gnd.n3085 gnd.n2946 31.8661
R7816 gnd.n3093 gnd.n2946 31.8661
R7817 gnd.n3093 gnd.n2939 31.8661
R7818 gnd.n3131 gnd.n2939 31.8661
R7819 gnd.n3141 gnd.n2872 31.8661
R7820 gnd.n4220 gnd.n2442 31.8661
R7821 gnd.n4234 gnd.n2431 31.8661
R7822 gnd.n4234 gnd.n2434 31.8661
R7823 gnd.n4243 gnd.n967 31.8661
R7824 gnd.n1243 gnd.n1141 31.8661
R7825 gnd.n2325 gnd.n1257 31.8661
R7826 gnd.n2325 gnd.n1154 31.8661
R7827 gnd.n4437 gnd.n1168 31.8661
R7828 gnd.n5873 gnd.n1588 31.8661
R7829 gnd.n5867 gnd.n5866 31.8661
R7830 gnd.n5866 gnd.n5865 31.8661
R7831 gnd.n5859 gnd.n1606 31.8661
R7832 gnd.n7301 gnd.n141 31.8661
R7833 gnd.n7295 gnd.n152 31.8661
R7834 gnd.n7289 gnd.n152 31.8661
R7835 gnd.n7283 gnd.n167 31.8661
R7836 gnd.n5417 gnd.n1826 31.3761
R7837 gnd.n2279 gnd.n2268 31.3761
R7838 gnd.n1232 gnd.n1231 25.7944
R7839 gnd.n5141 gnd.n5140 25.7944
R7840 gnd.n2932 gnd.n2931 25.7944
R7841 gnd.n2490 gnd.n2489 25.7944
R7842 gnd.n1239 gnd.n1238 25.7944
R7843 gnd.n5554 gnd.n5553 25.7944
R7844 gnd.n5606 gnd.n5605 25.7944
R7845 gnd.n1756 gnd.n1755 25.7944
R7846 gnd.n175 gnd.n174 25.7944
R7847 gnd.n197 gnd.n196 25.7944
R7848 gnd.n219 gnd.n218 25.7944
R7849 gnd.n7188 gnd.n7187 25.7944
R7850 gnd.n3968 gnd.n3967 25.7944
R7851 gnd.n3990 gnd.n3989 25.7944
R7852 gnd.n4013 gnd.n4012 25.7944
R7853 gnd.n4032 gnd.n4031 25.7944
R7854 gnd.n1309 gnd.n1308 25.7944
R7855 gnd.n1350 gnd.n1349 25.7944
R7856 gnd.n1329 gnd.n1328 25.7944
R7857 gnd.n5131 gnd.n5130 25.7944
R7858 gnd.n3153 gnd.n2873 24.8557
R7859 gnd.n3163 gnd.n2856 24.8557
R7860 gnd.n2859 gnd.n2847 24.8557
R7861 gnd.n3184 gnd.n2848 24.8557
R7862 gnd.n3194 gnd.n2828 24.8557
R7863 gnd.n3204 gnd.n3203 24.8557
R7864 gnd.n2814 gnd.n2812 24.8557
R7865 gnd.n3235 gnd.n3234 24.8557
R7866 gnd.n3250 gnd.n2797 24.8557
R7867 gnd.n3304 gnd.n2736 24.8557
R7868 gnd.n3260 gnd.n2737 24.8557
R7869 gnd.n3297 gnd.n2748 24.8557
R7870 gnd.n2786 gnd.n2785 24.8557
R7871 gnd.n3291 gnd.n3290 24.8557
R7872 gnd.n2772 gnd.n2759 24.8557
R7873 gnd.n3330 gnd.n3329 24.8557
R7874 gnd.n3340 gnd.n2668 24.8557
R7875 gnd.n3352 gnd.n2660 24.8557
R7876 gnd.n3351 gnd.n2648 24.8557
R7877 gnd.n3370 gnd.n3369 24.8557
R7878 gnd.n3380 gnd.n2641 24.8557
R7879 gnd.n3391 gnd.n2629 24.8557
R7880 gnd.n3415 gnd.n3414 24.8557
R7881 gnd.n3426 gnd.n2612 24.8557
R7882 gnd.n3425 gnd.n2614 24.8557
R7883 gnd.n3437 gnd.n2605 24.8557
R7884 gnd.n3455 gnd.n3454 24.8557
R7885 gnd.n2596 gnd.n2585 24.8557
R7886 gnd.n3476 gnd.n2573 24.8557
R7887 gnd.n3504 gnd.n3503 24.8557
R7888 gnd.n3515 gnd.n2558 24.8557
R7889 gnd.n3526 gnd.n2551 24.8557
R7890 gnd.n3525 gnd.n2539 24.8557
R7891 gnd.n3798 gnd.n3797 24.8557
R7892 gnd.n3820 gnd.n2524 24.8557
R7893 gnd.n6314 gnd.n960 24.678
R7894 gnd.n3174 gnd.t324 23.2624
R7895 gnd.n2875 gnd.t60 22.6251
R7896 gnd.t289 gnd.n2880 21.3504
R7897 gnd.n4252 gnd.n970 21.0318
R7898 gnd.n6299 gnd.n980 21.0318
R7899 gnd.n4260 gnd.n2415 21.0318
R7900 gnd.n6293 gnd.n991 21.0318
R7901 gnd.n6287 gnd.n1002 21.0318
R7902 gnd.n4279 gnd.n1005 21.0318
R7903 gnd.n2370 gnd.n1014 21.0318
R7904 gnd.n4333 gnd.n4332 21.0318
R7905 gnd.n6273 gnd.n1022 21.0318
R7906 gnd.n4326 gnd.n1025 21.0318
R7907 gnd.n4296 gnd.n1036 21.0318
R7908 gnd.n6260 gnd.n1041 21.0318
R7909 gnd.n4316 gnd.n4315 21.0318
R7910 gnd.n6254 gnd.n1050 21.0318
R7911 gnd.n6247 gnd.n1058 21.0318
R7912 gnd.n4363 gnd.n1061 21.0318
R7913 gnd.n4371 gnd.n1070 21.0318
R7914 gnd.n6235 gnd.n1078 21.0318
R7915 gnd.n4377 gnd.n2350 21.0318
R7916 gnd.n6229 gnd.n1087 21.0318
R7917 gnd.n6223 gnd.n1098 21.0318
R7918 gnd.n4409 gnd.n1101 21.0318
R7919 gnd.n4392 gnd.n1110 21.0318
R7920 gnd.n6211 gnd.n1118 21.0318
R7921 gnd.n4398 gnd.n1121 21.0318
R7922 gnd.n6205 gnd.n1128 21.0318
R7923 gnd.n6199 gnd.n1138 21.0318
R7924 gnd.n5858 gnd.n1609 21.0318
R7925 gnd.n5852 gnd.n1621 21.0318
R7926 gnd.n5669 gnd.n1630 21.0318
R7927 gnd.n5846 gnd.n1633 21.0318
R7928 gnd.n5677 gnd.n1641 21.0318
R7929 gnd.n5697 gnd.n1650 21.0318
R7930 gnd.n5834 gnd.n1653 21.0318
R7931 gnd.n5828 gnd.n1664 21.0318
R7932 gnd.n5742 gnd.n5741 21.0318
R7933 gnd.n5822 gnd.n1673 21.0318
R7934 gnd.n5749 gnd.n1681 21.0318
R7935 gnd.n5767 gnd.n1690 21.0318
R7936 gnd.n5810 gnd.n1693 21.0318
R7937 gnd.n1705 gnd.n1699 21.0318
R7938 gnd.n5798 gnd.n1706 21.0318
R7939 gnd.n5797 gnd.n1709 21.0318
R7940 gnd.n5792 gnd.n1722 21.0318
R7941 gnd.n7339 gnd.n71 21.0318
R7942 gnd.n7137 gnd.n7136 21.0318
R7943 gnd.n7144 gnd.n86 21.0318
R7944 gnd.n7331 gnd.n89 21.0318
R7945 gnd.n7325 gnd.n101 21.0318
R7946 gnd.n7159 gnd.n108 21.0318
R7947 gnd.n7167 gnd.n117 21.0318
R7948 gnd.n7313 gnd.n120 21.0318
R7949 gnd.n7174 gnd.n128 21.0318
R7950 gnd.n7307 gnd.n131 21.0318
R7951 gnd.t292 gnd.n2586 20.7131
R7952 gnd.n6281 gnd.t138 20.7131
R7953 gnd.t185 gnd.n1053 20.7131
R7954 gnd.t153 gnd.n5805 20.7131
R7955 gnd.n7152 gnd.t188 20.7131
R7956 gnd.n6116 gnd.n1243 20.3945
R7957 gnd.n1606 gnd.n1598 20.3945
R7958 gnd.t218 gnd.n2621 20.0758
R7959 gnd.t169 gnd.n6305 20.0758
R7960 gnd.t206 gnd.n1090 20.0758
R7961 gnd.t190 gnd.n1661 20.0758
R7962 gnd.n7266 gnd.t6 20.0758
R7963 gnd.n2206 gnd.n2205 19.9763
R7964 gnd.n1825 gnd.n1824 19.9763
R7965 gnd.n5998 gnd.n5997 19.9763
R7966 gnd.n5348 gnd.n5347 19.9763
R7967 gnd.n1462 gnd.t41 19.8005
R7968 gnd.n1462 gnd.t104 19.8005
R7969 gnd.n1461 gnd.t65 19.8005
R7970 gnd.n1461 gnd.t85 19.8005
R7971 gnd.n5338 gnd.t16 19.8005
R7972 gnd.n5338 gnd.t130 19.8005
R7973 gnd.n5337 gnd.t78 19.8005
R7974 gnd.n5337 gnd.t55 19.8005
R7975 gnd.n1458 gnd.n1457 19.5087
R7976 gnd.n1471 gnd.n1458 19.5087
R7977 gnd.n1469 gnd.n1460 19.5087
R7978 gnd.n5342 gnd.n5336 19.5087
R7979 gnd.n3341 gnd.t11 19.4385
R7980 gnd.n4243 gnd.n2423 19.4385
R7981 gnd.n149 gnd.n141 19.4385
R7982 gnd.n2317 gnd.n2314 19.3944
R7983 gnd.n2317 gnd.n2303 19.3944
R7984 gnd.n4459 gnd.n2303 19.3944
R7985 gnd.n4459 gnd.n2300 19.3944
R7986 gnd.n4466 gnd.n2300 19.3944
R7987 gnd.n4466 gnd.n2301 19.3944
R7988 gnd.n4462 gnd.n2301 19.3944
R7989 gnd.n4462 gnd.n2202 19.3944
R7990 gnd.n4496 gnd.n2202 19.3944
R7991 gnd.n4496 gnd.n2199 19.3944
R7992 gnd.n4501 gnd.n2199 19.3944
R7993 gnd.n4501 gnd.n2200 19.3944
R7994 gnd.n2200 gnd.n2191 19.3944
R7995 gnd.n4521 gnd.n2191 19.3944
R7996 gnd.n4521 gnd.n2188 19.3944
R7997 gnd.n4532 gnd.n2188 19.3944
R7998 gnd.n4532 gnd.n2189 19.3944
R7999 gnd.n4528 gnd.n2189 19.3944
R8000 gnd.n4528 gnd.n4527 19.3944
R8001 gnd.n4527 gnd.n2144 19.3944
R8002 gnd.n4607 gnd.n2144 19.3944
R8003 gnd.n4607 gnd.n2141 19.3944
R8004 gnd.n4630 gnd.n2141 19.3944
R8005 gnd.n4630 gnd.n2142 19.3944
R8006 gnd.n4626 gnd.n2142 19.3944
R8007 gnd.n4626 gnd.n4625 19.3944
R8008 gnd.n4625 gnd.n4624 19.3944
R8009 gnd.n4624 gnd.n4616 19.3944
R8010 gnd.n4620 gnd.n4616 19.3944
R8011 gnd.n4620 gnd.n4619 19.3944
R8012 gnd.n4619 gnd.n2094 19.3944
R8013 gnd.n2094 gnd.n2092 19.3944
R8014 gnd.n4709 gnd.n2092 19.3944
R8015 gnd.n4709 gnd.n2090 19.3944
R8016 gnd.n4713 gnd.n2090 19.3944
R8017 gnd.n4713 gnd.n2065 19.3944
R8018 gnd.n4759 gnd.n2065 19.3944
R8019 gnd.n4759 gnd.n2066 19.3944
R8020 gnd.n4755 gnd.n2066 19.3944
R8021 gnd.n4755 gnd.n2042 19.3944
R8022 gnd.n4818 gnd.n2042 19.3944
R8023 gnd.n4818 gnd.n2043 19.3944
R8024 gnd.n4814 gnd.n2043 19.3944
R8025 gnd.n4814 gnd.n4813 19.3944
R8026 gnd.n4813 gnd.n4812 19.3944
R8027 gnd.n4812 gnd.n4798 19.3944
R8028 gnd.n4808 gnd.n4798 19.3944
R8029 gnd.n4808 gnd.n4807 19.3944
R8030 gnd.n4807 gnd.n4806 19.3944
R8031 gnd.n4806 gnd.n1983 19.3944
R8032 gnd.n4926 gnd.n1983 19.3944
R8033 gnd.n4926 gnd.n1980 19.3944
R8034 gnd.n4931 gnd.n1980 19.3944
R8035 gnd.n4931 gnd.n1981 19.3944
R8036 gnd.n1981 gnd.n1954 19.3944
R8037 gnd.n4965 gnd.n1954 19.3944
R8038 gnd.n4965 gnd.n1951 19.3944
R8039 gnd.n4984 gnd.n1951 19.3944
R8040 gnd.n4984 gnd.n1952 19.3944
R8041 gnd.n4980 gnd.n1952 19.3944
R8042 gnd.n4980 gnd.n4979 19.3944
R8043 gnd.n4979 gnd.n4978 19.3944
R8044 gnd.n4978 gnd.n4973 19.3944
R8045 gnd.n4974 gnd.n4973 19.3944
R8046 gnd.n4974 gnd.n1898 19.3944
R8047 gnd.n5056 gnd.n1898 19.3944
R8048 gnd.n5056 gnd.n1895 19.3944
R8049 gnd.n5061 gnd.n1895 19.3944
R8050 gnd.n5061 gnd.n1896 19.3944
R8051 gnd.n1896 gnd.n1871 19.3944
R8052 gnd.n5098 gnd.n1871 19.3944
R8053 gnd.n5098 gnd.n1869 19.3944
R8054 gnd.n5102 gnd.n1869 19.3944
R8055 gnd.n5102 gnd.n1868 19.3944
R8056 gnd.n5109 gnd.n1868 19.3944
R8057 gnd.n5109 gnd.n1866 19.3944
R8058 gnd.n5113 gnd.n1866 19.3944
R8059 gnd.n5114 gnd.n5113 19.3944
R8060 gnd.n5117 gnd.n5114 19.3944
R8061 gnd.n5117 gnd.n1863 19.3944
R8062 gnd.n5299 gnd.n1863 19.3944
R8063 gnd.n5299 gnd.n1864 19.3944
R8064 gnd.n1235 gnd.n1151 19.3944
R8065 gnd.n6185 gnd.n1151 19.3944
R8066 gnd.n6185 gnd.n6184 19.3944
R8067 gnd.n6178 gnd.n6177 19.3944
R8068 gnd.n6177 gnd.n1173 19.3944
R8069 gnd.n6173 gnd.n1173 19.3944
R8070 gnd.n6173 gnd.n6172 19.3944
R8071 gnd.n6172 gnd.n6171 19.3944
R8072 gnd.n6171 gnd.n1178 19.3944
R8073 gnd.n6166 gnd.n1178 19.3944
R8074 gnd.n6166 gnd.n6165 19.3944
R8075 gnd.n6165 gnd.n6164 19.3944
R8076 gnd.n6164 gnd.n1184 19.3944
R8077 gnd.n6157 gnd.n1184 19.3944
R8078 gnd.n6157 gnd.n6156 19.3944
R8079 gnd.n6156 gnd.n1196 19.3944
R8080 gnd.n6149 gnd.n1196 19.3944
R8081 gnd.n6149 gnd.n6148 19.3944
R8082 gnd.n6148 gnd.n1204 19.3944
R8083 gnd.n6141 gnd.n1204 19.3944
R8084 gnd.n6141 gnd.n6140 19.3944
R8085 gnd.n6140 gnd.n1214 19.3944
R8086 gnd.n6133 gnd.n1214 19.3944
R8087 gnd.n6133 gnd.n6132 19.3944
R8088 gnd.n6132 gnd.n1222 19.3944
R8089 gnd.n6125 gnd.n1222 19.3944
R8090 gnd.n6125 gnd.n6124 19.3944
R8091 gnd.n5207 gnd.n5171 19.3944
R8092 gnd.n5220 gnd.n5171 19.3944
R8093 gnd.n5220 gnd.n5169 19.3944
R8094 gnd.n5226 gnd.n5169 19.3944
R8095 gnd.n5226 gnd.n5162 19.3944
R8096 gnd.n5239 gnd.n5162 19.3944
R8097 gnd.n5239 gnd.n5160 19.3944
R8098 gnd.n5245 gnd.n5160 19.3944
R8099 gnd.n5245 gnd.n5153 19.3944
R8100 gnd.n5258 gnd.n5153 19.3944
R8101 gnd.n5258 gnd.n5151 19.3944
R8102 gnd.n5264 gnd.n5151 19.3944
R8103 gnd.n5264 gnd.n5144 19.3944
R8104 gnd.n5278 gnd.n5144 19.3944
R8105 gnd.n5278 gnd.n5142 19.3944
R8106 gnd.n5284 gnd.n5142 19.3944
R8107 gnd.n3056 gnd.n3055 19.3944
R8108 gnd.n3055 gnd.n3054 19.3944
R8109 gnd.n3054 gnd.n3053 19.3944
R8110 gnd.n3053 gnd.n3051 19.3944
R8111 gnd.n3051 gnd.n3048 19.3944
R8112 gnd.n3048 gnd.n3047 19.3944
R8113 gnd.n3047 gnd.n3044 19.3944
R8114 gnd.n3044 gnd.n3043 19.3944
R8115 gnd.n3043 gnd.n3040 19.3944
R8116 gnd.n3040 gnd.n3039 19.3944
R8117 gnd.n3039 gnd.n3036 19.3944
R8118 gnd.n3036 gnd.n3035 19.3944
R8119 gnd.n3035 gnd.n3032 19.3944
R8120 gnd.n3032 gnd.n3031 19.3944
R8121 gnd.n3031 gnd.n3028 19.3944
R8122 gnd.n3028 gnd.n3027 19.3944
R8123 gnd.n3027 gnd.n3024 19.3944
R8124 gnd.n3024 gnd.n3023 19.3944
R8125 gnd.n3023 gnd.n3020 19.3944
R8126 gnd.n3020 gnd.n3019 19.3944
R8127 gnd.n3019 gnd.n3016 19.3944
R8128 gnd.n3016 gnd.n3015 19.3944
R8129 gnd.n3012 gnd.n3011 19.3944
R8130 gnd.n3011 gnd.n2967 19.3944
R8131 gnd.n3062 gnd.n2967 19.3944
R8132 gnd.n3828 gnd.n3827 19.3944
R8133 gnd.n3827 gnd.n3824 19.3944
R8134 gnd.n3824 gnd.n3823 19.3944
R8135 gnd.n3873 gnd.n3872 19.3944
R8136 gnd.n3872 gnd.n3871 19.3944
R8137 gnd.n3871 gnd.n3868 19.3944
R8138 gnd.n3868 gnd.n3867 19.3944
R8139 gnd.n3867 gnd.n3864 19.3944
R8140 gnd.n3864 gnd.n3863 19.3944
R8141 gnd.n3863 gnd.n3860 19.3944
R8142 gnd.n3860 gnd.n3859 19.3944
R8143 gnd.n3859 gnd.n3856 19.3944
R8144 gnd.n3856 gnd.n3855 19.3944
R8145 gnd.n3855 gnd.n3852 19.3944
R8146 gnd.n3852 gnd.n3851 19.3944
R8147 gnd.n3851 gnd.n3848 19.3944
R8148 gnd.n3848 gnd.n3847 19.3944
R8149 gnd.n3847 gnd.n3844 19.3944
R8150 gnd.n3844 gnd.n3843 19.3944
R8151 gnd.n3843 gnd.n3840 19.3944
R8152 gnd.n3840 gnd.n3839 19.3944
R8153 gnd.n3839 gnd.n3836 19.3944
R8154 gnd.n3836 gnd.n3835 19.3944
R8155 gnd.n3835 gnd.n3832 19.3944
R8156 gnd.n3832 gnd.n3831 19.3944
R8157 gnd.n3155 gnd.n2864 19.3944
R8158 gnd.n3165 gnd.n2864 19.3944
R8159 gnd.n3166 gnd.n3165 19.3944
R8160 gnd.n3166 gnd.n2845 19.3944
R8161 gnd.n3186 gnd.n2845 19.3944
R8162 gnd.n3186 gnd.n2837 19.3944
R8163 gnd.n3196 gnd.n2837 19.3944
R8164 gnd.n3197 gnd.n3196 19.3944
R8165 gnd.n3198 gnd.n3197 19.3944
R8166 gnd.n3198 gnd.n2820 19.3944
R8167 gnd.n3215 gnd.n2820 19.3944
R8168 gnd.n3218 gnd.n3215 19.3944
R8169 gnd.n3218 gnd.n3217 19.3944
R8170 gnd.n3217 gnd.n2793 19.3944
R8171 gnd.n3257 gnd.n2793 19.3944
R8172 gnd.n3257 gnd.n2790 19.3944
R8173 gnd.n3263 gnd.n2790 19.3944
R8174 gnd.n3264 gnd.n3263 19.3944
R8175 gnd.n3264 gnd.n2788 19.3944
R8176 gnd.n3270 gnd.n2788 19.3944
R8177 gnd.n3273 gnd.n3270 19.3944
R8178 gnd.n3275 gnd.n3273 19.3944
R8179 gnd.n3281 gnd.n3275 19.3944
R8180 gnd.n3281 gnd.n3280 19.3944
R8181 gnd.n3280 gnd.n2663 19.3944
R8182 gnd.n3347 gnd.n2663 19.3944
R8183 gnd.n3348 gnd.n3347 19.3944
R8184 gnd.n3348 gnd.n2656 19.3944
R8185 gnd.n3359 gnd.n2656 19.3944
R8186 gnd.n3360 gnd.n3359 19.3944
R8187 gnd.n3360 gnd.n2639 19.3944
R8188 gnd.n2639 gnd.n2637 19.3944
R8189 gnd.n3384 gnd.n2637 19.3944
R8190 gnd.n3385 gnd.n3384 19.3944
R8191 gnd.n3385 gnd.n2608 19.3944
R8192 gnd.n3432 gnd.n2608 19.3944
R8193 gnd.n3433 gnd.n3432 19.3944
R8194 gnd.n3433 gnd.n2601 19.3944
R8195 gnd.n3444 gnd.n2601 19.3944
R8196 gnd.n3445 gnd.n3444 19.3944
R8197 gnd.n3445 gnd.n2584 19.3944
R8198 gnd.n2584 gnd.n2582 19.3944
R8199 gnd.n3469 gnd.n2582 19.3944
R8200 gnd.n3470 gnd.n3469 19.3944
R8201 gnd.n3470 gnd.n2554 19.3944
R8202 gnd.n3521 gnd.n2554 19.3944
R8203 gnd.n3522 gnd.n3521 19.3944
R8204 gnd.n3522 gnd.n2547 19.3944
R8205 gnd.n3789 gnd.n2547 19.3944
R8206 gnd.n3790 gnd.n3789 19.3944
R8207 gnd.n3790 gnd.n2528 19.3944
R8208 gnd.n3815 gnd.n2528 19.3944
R8209 gnd.n3815 gnd.n2529 19.3944
R8210 gnd.n3146 gnd.n3145 19.3944
R8211 gnd.n3145 gnd.n2878 19.3944
R8212 gnd.n2901 gnd.n2878 19.3944
R8213 gnd.n2904 gnd.n2901 19.3944
R8214 gnd.n2904 gnd.n2897 19.3944
R8215 gnd.n2908 gnd.n2897 19.3944
R8216 gnd.n2911 gnd.n2908 19.3944
R8217 gnd.n2914 gnd.n2911 19.3944
R8218 gnd.n2914 gnd.n2895 19.3944
R8219 gnd.n2918 gnd.n2895 19.3944
R8220 gnd.n2921 gnd.n2918 19.3944
R8221 gnd.n2924 gnd.n2921 19.3944
R8222 gnd.n2924 gnd.n2893 19.3944
R8223 gnd.n2928 gnd.n2893 19.3944
R8224 gnd.n3151 gnd.n3150 19.3944
R8225 gnd.n3150 gnd.n2854 19.3944
R8226 gnd.n3176 gnd.n2854 19.3944
R8227 gnd.n3176 gnd.n2852 19.3944
R8228 gnd.n3182 gnd.n2852 19.3944
R8229 gnd.n3182 gnd.n3181 19.3944
R8230 gnd.n3181 gnd.n2826 19.3944
R8231 gnd.n3206 gnd.n2826 19.3944
R8232 gnd.n3206 gnd.n2824 19.3944
R8233 gnd.n3210 gnd.n2824 19.3944
R8234 gnd.n3210 gnd.n2804 19.3944
R8235 gnd.n3237 gnd.n2804 19.3944
R8236 gnd.n3237 gnd.n2802 19.3944
R8237 gnd.n3247 gnd.n2802 19.3944
R8238 gnd.n3247 gnd.n3246 19.3944
R8239 gnd.n3246 gnd.n3245 19.3944
R8240 gnd.n3245 gnd.n2751 19.3944
R8241 gnd.n3295 gnd.n2751 19.3944
R8242 gnd.n3295 gnd.n3294 19.3944
R8243 gnd.n3294 gnd.n3293 19.3944
R8244 gnd.n3293 gnd.n2755 19.3944
R8245 gnd.n2775 gnd.n2755 19.3944
R8246 gnd.n2775 gnd.n2673 19.3944
R8247 gnd.n3332 gnd.n2673 19.3944
R8248 gnd.n3332 gnd.n2671 19.3944
R8249 gnd.n3338 gnd.n2671 19.3944
R8250 gnd.n3338 gnd.n3337 19.3944
R8251 gnd.n3337 gnd.n2646 19.3944
R8252 gnd.n3372 gnd.n2646 19.3944
R8253 gnd.n3372 gnd.n2644 19.3944
R8254 gnd.n3378 gnd.n2644 19.3944
R8255 gnd.n3378 gnd.n3377 19.3944
R8256 gnd.n3377 gnd.n2619 19.3944
R8257 gnd.n3417 gnd.n2619 19.3944
R8258 gnd.n3417 gnd.n2617 19.3944
R8259 gnd.n3423 gnd.n2617 19.3944
R8260 gnd.n3423 gnd.n3422 19.3944
R8261 gnd.n3422 gnd.n2591 19.3944
R8262 gnd.n3457 gnd.n2591 19.3944
R8263 gnd.n3457 gnd.n2589 19.3944
R8264 gnd.n3463 gnd.n2589 19.3944
R8265 gnd.n3463 gnd.n3462 19.3944
R8266 gnd.n3462 gnd.n2564 19.3944
R8267 gnd.n3506 gnd.n2564 19.3944
R8268 gnd.n3506 gnd.n2562 19.3944
R8269 gnd.n3512 gnd.n2562 19.3944
R8270 gnd.n3512 gnd.n3511 19.3944
R8271 gnd.n3511 gnd.n2537 19.3944
R8272 gnd.n3800 gnd.n2537 19.3944
R8273 gnd.n3800 gnd.n2535 19.3944
R8274 gnd.n3808 gnd.n2535 19.3944
R8275 gnd.n3808 gnd.n3807 19.3944
R8276 gnd.n3807 gnd.n3806 19.3944
R8277 gnd.n3909 gnd.n3908 19.3944
R8278 gnd.n3908 gnd.n2476 19.3944
R8279 gnd.n3904 gnd.n2476 19.3944
R8280 gnd.n3904 gnd.n3901 19.3944
R8281 gnd.n3901 gnd.n3898 19.3944
R8282 gnd.n3898 gnd.n3897 19.3944
R8283 gnd.n3897 gnd.n3894 19.3944
R8284 gnd.n3894 gnd.n3893 19.3944
R8285 gnd.n3893 gnd.n3890 19.3944
R8286 gnd.n3890 gnd.n3889 19.3944
R8287 gnd.n3889 gnd.n3886 19.3944
R8288 gnd.n3886 gnd.n3885 19.3944
R8289 gnd.n3885 gnd.n3882 19.3944
R8290 gnd.n3882 gnd.n3881 19.3944
R8291 gnd.n3066 gnd.n2965 19.3944
R8292 gnd.n3066 gnd.n2956 19.3944
R8293 gnd.n3079 gnd.n2956 19.3944
R8294 gnd.n3079 gnd.n2954 19.3944
R8295 gnd.n3083 gnd.n2954 19.3944
R8296 gnd.n3083 gnd.n2944 19.3944
R8297 gnd.n3095 gnd.n2944 19.3944
R8298 gnd.n3095 gnd.n2942 19.3944
R8299 gnd.n3129 gnd.n2942 19.3944
R8300 gnd.n3129 gnd.n3128 19.3944
R8301 gnd.n3128 gnd.n3127 19.3944
R8302 gnd.n3127 gnd.n3126 19.3944
R8303 gnd.n3126 gnd.n3123 19.3944
R8304 gnd.n3123 gnd.n3122 19.3944
R8305 gnd.n3122 gnd.n3121 19.3944
R8306 gnd.n3121 gnd.n3119 19.3944
R8307 gnd.n3119 gnd.n3118 19.3944
R8308 gnd.n3118 gnd.n3115 19.3944
R8309 gnd.n3115 gnd.n3114 19.3944
R8310 gnd.n3114 gnd.n3113 19.3944
R8311 gnd.n3113 gnd.n3111 19.3944
R8312 gnd.n3111 gnd.n2810 19.3944
R8313 gnd.n3226 gnd.n2810 19.3944
R8314 gnd.n3226 gnd.n2808 19.3944
R8315 gnd.n3232 gnd.n2808 19.3944
R8316 gnd.n3232 gnd.n3231 19.3944
R8317 gnd.n3231 gnd.n2732 19.3944
R8318 gnd.n3306 gnd.n2732 19.3944
R8319 gnd.n3306 gnd.n2733 19.3944
R8320 gnd.n2780 gnd.n2779 19.3944
R8321 gnd.n2783 gnd.n2782 19.3944
R8322 gnd.n2770 gnd.n2769 19.3944
R8323 gnd.n3325 gnd.n2678 19.3944
R8324 gnd.n3325 gnd.n3324 19.3944
R8325 gnd.n3324 gnd.n3323 19.3944
R8326 gnd.n3323 gnd.n3321 19.3944
R8327 gnd.n3321 gnd.n3320 19.3944
R8328 gnd.n3320 gnd.n3318 19.3944
R8329 gnd.n3318 gnd.n3317 19.3944
R8330 gnd.n3317 gnd.n2627 19.3944
R8331 gnd.n3393 gnd.n2627 19.3944
R8332 gnd.n3393 gnd.n2625 19.3944
R8333 gnd.n3412 gnd.n2625 19.3944
R8334 gnd.n3412 gnd.n3411 19.3944
R8335 gnd.n3411 gnd.n3410 19.3944
R8336 gnd.n3410 gnd.n3408 19.3944
R8337 gnd.n3408 gnd.n3407 19.3944
R8338 gnd.n3407 gnd.n3405 19.3944
R8339 gnd.n3405 gnd.n3404 19.3944
R8340 gnd.n3404 gnd.n2571 19.3944
R8341 gnd.n3478 gnd.n2571 19.3944
R8342 gnd.n3478 gnd.n2569 19.3944
R8343 gnd.n3501 gnd.n2569 19.3944
R8344 gnd.n3501 gnd.n3500 19.3944
R8345 gnd.n3500 gnd.n3499 19.3944
R8346 gnd.n3499 gnd.n3496 19.3944
R8347 gnd.n3496 gnd.n3495 19.3944
R8348 gnd.n3495 gnd.n3493 19.3944
R8349 gnd.n3493 gnd.n3492 19.3944
R8350 gnd.n3492 gnd.n3490 19.3944
R8351 gnd.n3490 gnd.n2523 19.3944
R8352 gnd.n3071 gnd.n2961 19.3944
R8353 gnd.n3071 gnd.n2959 19.3944
R8354 gnd.n3075 gnd.n2959 19.3944
R8355 gnd.n3075 gnd.n2950 19.3944
R8356 gnd.n3087 gnd.n2950 19.3944
R8357 gnd.n3087 gnd.n2948 19.3944
R8358 gnd.n3091 gnd.n2948 19.3944
R8359 gnd.n3091 gnd.n2937 19.3944
R8360 gnd.n3133 gnd.n2937 19.3944
R8361 gnd.n3133 gnd.n2891 19.3944
R8362 gnd.n3139 gnd.n2891 19.3944
R8363 gnd.n3139 gnd.n3138 19.3944
R8364 gnd.n3138 gnd.n2869 19.3944
R8365 gnd.n3160 gnd.n2869 19.3944
R8366 gnd.n3160 gnd.n2862 19.3944
R8367 gnd.n3171 gnd.n2862 19.3944
R8368 gnd.n3171 gnd.n3170 19.3944
R8369 gnd.n3170 gnd.n2843 19.3944
R8370 gnd.n3191 gnd.n2843 19.3944
R8371 gnd.n3191 gnd.n2833 19.3944
R8372 gnd.n3201 gnd.n2833 19.3944
R8373 gnd.n3201 gnd.n2816 19.3944
R8374 gnd.n3222 gnd.n2816 19.3944
R8375 gnd.n3222 gnd.n3221 19.3944
R8376 gnd.n3221 gnd.n2795 19.3944
R8377 gnd.n3252 gnd.n2795 19.3944
R8378 gnd.n3252 gnd.n2740 19.3944
R8379 gnd.n3302 gnd.n2740 19.3944
R8380 gnd.n3302 gnd.n3301 19.3944
R8381 gnd.n3301 gnd.n3300 19.3944
R8382 gnd.n3300 gnd.n2744 19.3944
R8383 gnd.n2762 gnd.n2744 19.3944
R8384 gnd.n3288 gnd.n2762 19.3944
R8385 gnd.n3288 gnd.n3287 19.3944
R8386 gnd.n3287 gnd.n3286 19.3944
R8387 gnd.n3286 gnd.n2766 19.3944
R8388 gnd.n2766 gnd.n2665 19.3944
R8389 gnd.n3343 gnd.n2665 19.3944
R8390 gnd.n3343 gnd.n2658 19.3944
R8391 gnd.n3354 gnd.n2658 19.3944
R8392 gnd.n3354 gnd.n2654 19.3944
R8393 gnd.n3367 gnd.n2654 19.3944
R8394 gnd.n3367 gnd.n3366 19.3944
R8395 gnd.n3366 gnd.n2633 19.3944
R8396 gnd.n3389 gnd.n2633 19.3944
R8397 gnd.n3389 gnd.n3388 19.3944
R8398 gnd.n3388 gnd.n2610 19.3944
R8399 gnd.n3428 gnd.n2610 19.3944
R8400 gnd.n3428 gnd.n2603 19.3944
R8401 gnd.n3439 gnd.n2603 19.3944
R8402 gnd.n3439 gnd.n2599 19.3944
R8403 gnd.n3452 gnd.n2599 19.3944
R8404 gnd.n3452 gnd.n3451 19.3944
R8405 gnd.n3451 gnd.n2578 19.3944
R8406 gnd.n3474 gnd.n2578 19.3944
R8407 gnd.n3474 gnd.n3473 19.3944
R8408 gnd.n3473 gnd.n2556 19.3944
R8409 gnd.n3517 gnd.n2556 19.3944
R8410 gnd.n3517 gnd.n2549 19.3944
R8411 gnd.n3528 gnd.n2549 19.3944
R8412 gnd.n3528 gnd.n2545 19.3944
R8413 gnd.n3795 gnd.n2545 19.3944
R8414 gnd.n3795 gnd.n3794 19.3944
R8415 gnd.n3794 gnd.n2526 19.3944
R8416 gnd.n3818 gnd.n2526 19.3944
R8417 gnd.n6161 gnd.n1187 19.3944
R8418 gnd.n6161 gnd.n6160 19.3944
R8419 gnd.n6160 gnd.n1190 19.3944
R8420 gnd.n6153 gnd.n1190 19.3944
R8421 gnd.n6153 gnd.n6152 19.3944
R8422 gnd.n6152 gnd.n1200 19.3944
R8423 gnd.n6145 gnd.n1200 19.3944
R8424 gnd.n6145 gnd.n6144 19.3944
R8425 gnd.n6144 gnd.n1208 19.3944
R8426 gnd.n6137 gnd.n1208 19.3944
R8427 gnd.n6137 gnd.n6136 19.3944
R8428 gnd.n6136 gnd.n1218 19.3944
R8429 gnd.n6129 gnd.n1218 19.3944
R8430 gnd.n6129 gnd.n6128 19.3944
R8431 gnd.n6128 gnd.n1226 19.3944
R8432 gnd.n6121 gnd.n1226 19.3944
R8433 gnd.n6903 gnd.n542 19.3944
R8434 gnd.n6909 gnd.n542 19.3944
R8435 gnd.n6909 gnd.n540 19.3944
R8436 gnd.n6913 gnd.n540 19.3944
R8437 gnd.n6913 gnd.n536 19.3944
R8438 gnd.n6919 gnd.n536 19.3944
R8439 gnd.n6919 gnd.n534 19.3944
R8440 gnd.n6923 gnd.n534 19.3944
R8441 gnd.n6923 gnd.n530 19.3944
R8442 gnd.n6929 gnd.n530 19.3944
R8443 gnd.n6929 gnd.n528 19.3944
R8444 gnd.n6933 gnd.n528 19.3944
R8445 gnd.n6933 gnd.n524 19.3944
R8446 gnd.n6939 gnd.n524 19.3944
R8447 gnd.n6939 gnd.n522 19.3944
R8448 gnd.n6943 gnd.n522 19.3944
R8449 gnd.n6943 gnd.n518 19.3944
R8450 gnd.n6949 gnd.n518 19.3944
R8451 gnd.n6949 gnd.n516 19.3944
R8452 gnd.n6953 gnd.n516 19.3944
R8453 gnd.n6953 gnd.n512 19.3944
R8454 gnd.n6959 gnd.n512 19.3944
R8455 gnd.n6959 gnd.n510 19.3944
R8456 gnd.n6963 gnd.n510 19.3944
R8457 gnd.n6963 gnd.n506 19.3944
R8458 gnd.n6969 gnd.n506 19.3944
R8459 gnd.n6969 gnd.n504 19.3944
R8460 gnd.n6973 gnd.n504 19.3944
R8461 gnd.n6973 gnd.n500 19.3944
R8462 gnd.n6979 gnd.n500 19.3944
R8463 gnd.n6979 gnd.n498 19.3944
R8464 gnd.n6983 gnd.n498 19.3944
R8465 gnd.n6983 gnd.n494 19.3944
R8466 gnd.n6989 gnd.n494 19.3944
R8467 gnd.n6989 gnd.n492 19.3944
R8468 gnd.n6993 gnd.n492 19.3944
R8469 gnd.n6993 gnd.n488 19.3944
R8470 gnd.n6999 gnd.n488 19.3944
R8471 gnd.n6999 gnd.n486 19.3944
R8472 gnd.n7003 gnd.n486 19.3944
R8473 gnd.n7003 gnd.n482 19.3944
R8474 gnd.n7009 gnd.n482 19.3944
R8475 gnd.n7009 gnd.n480 19.3944
R8476 gnd.n7013 gnd.n480 19.3944
R8477 gnd.n7013 gnd.n476 19.3944
R8478 gnd.n7019 gnd.n476 19.3944
R8479 gnd.n7019 gnd.n474 19.3944
R8480 gnd.n7023 gnd.n474 19.3944
R8481 gnd.n7023 gnd.n470 19.3944
R8482 gnd.n7029 gnd.n470 19.3944
R8483 gnd.n7029 gnd.n468 19.3944
R8484 gnd.n7033 gnd.n468 19.3944
R8485 gnd.n7033 gnd.n464 19.3944
R8486 gnd.n7039 gnd.n464 19.3944
R8487 gnd.n7039 gnd.n462 19.3944
R8488 gnd.n7043 gnd.n462 19.3944
R8489 gnd.n7043 gnd.n458 19.3944
R8490 gnd.n7049 gnd.n458 19.3944
R8491 gnd.n7049 gnd.n456 19.3944
R8492 gnd.n7053 gnd.n456 19.3944
R8493 gnd.n7053 gnd.n452 19.3944
R8494 gnd.n7059 gnd.n452 19.3944
R8495 gnd.n7059 gnd.n450 19.3944
R8496 gnd.n7063 gnd.n450 19.3944
R8497 gnd.n7063 gnd.n446 19.3944
R8498 gnd.n7069 gnd.n446 19.3944
R8499 gnd.n7069 gnd.n444 19.3944
R8500 gnd.n7073 gnd.n444 19.3944
R8501 gnd.n7073 gnd.n440 19.3944
R8502 gnd.n7079 gnd.n440 19.3944
R8503 gnd.n7079 gnd.n438 19.3944
R8504 gnd.n7083 gnd.n438 19.3944
R8505 gnd.n7083 gnd.n434 19.3944
R8506 gnd.n7089 gnd.n434 19.3944
R8507 gnd.n7089 gnd.n432 19.3944
R8508 gnd.n7093 gnd.n432 19.3944
R8509 gnd.n7093 gnd.n428 19.3944
R8510 gnd.n7099 gnd.n428 19.3944
R8511 gnd.n7099 gnd.n426 19.3944
R8512 gnd.n7103 gnd.n426 19.3944
R8513 gnd.n7103 gnd.n422 19.3944
R8514 gnd.n7110 gnd.n422 19.3944
R8515 gnd.n7110 gnd.n420 19.3944
R8516 gnd.n7115 gnd.n420 19.3944
R8517 gnd.n6482 gnd.n793 19.3944
R8518 gnd.n6488 gnd.n793 19.3944
R8519 gnd.n6488 gnd.n791 19.3944
R8520 gnd.n6492 gnd.n791 19.3944
R8521 gnd.n6492 gnd.n787 19.3944
R8522 gnd.n6498 gnd.n787 19.3944
R8523 gnd.n6498 gnd.n785 19.3944
R8524 gnd.n6502 gnd.n785 19.3944
R8525 gnd.n6502 gnd.n781 19.3944
R8526 gnd.n6508 gnd.n781 19.3944
R8527 gnd.n6508 gnd.n779 19.3944
R8528 gnd.n6512 gnd.n779 19.3944
R8529 gnd.n6512 gnd.n775 19.3944
R8530 gnd.n6518 gnd.n775 19.3944
R8531 gnd.n6518 gnd.n773 19.3944
R8532 gnd.n6522 gnd.n773 19.3944
R8533 gnd.n6522 gnd.n769 19.3944
R8534 gnd.n6528 gnd.n769 19.3944
R8535 gnd.n6528 gnd.n767 19.3944
R8536 gnd.n6532 gnd.n767 19.3944
R8537 gnd.n6532 gnd.n763 19.3944
R8538 gnd.n6538 gnd.n763 19.3944
R8539 gnd.n6538 gnd.n761 19.3944
R8540 gnd.n6542 gnd.n761 19.3944
R8541 gnd.n6542 gnd.n757 19.3944
R8542 gnd.n6548 gnd.n757 19.3944
R8543 gnd.n6548 gnd.n755 19.3944
R8544 gnd.n6552 gnd.n755 19.3944
R8545 gnd.n6552 gnd.n751 19.3944
R8546 gnd.n6558 gnd.n751 19.3944
R8547 gnd.n6558 gnd.n749 19.3944
R8548 gnd.n6562 gnd.n749 19.3944
R8549 gnd.n6562 gnd.n745 19.3944
R8550 gnd.n6568 gnd.n745 19.3944
R8551 gnd.n6568 gnd.n743 19.3944
R8552 gnd.n6572 gnd.n743 19.3944
R8553 gnd.n6572 gnd.n739 19.3944
R8554 gnd.n6578 gnd.n739 19.3944
R8555 gnd.n6578 gnd.n737 19.3944
R8556 gnd.n6582 gnd.n737 19.3944
R8557 gnd.n6582 gnd.n733 19.3944
R8558 gnd.n6588 gnd.n733 19.3944
R8559 gnd.n6588 gnd.n731 19.3944
R8560 gnd.n6592 gnd.n731 19.3944
R8561 gnd.n6592 gnd.n727 19.3944
R8562 gnd.n6598 gnd.n727 19.3944
R8563 gnd.n6598 gnd.n725 19.3944
R8564 gnd.n6602 gnd.n725 19.3944
R8565 gnd.n6602 gnd.n721 19.3944
R8566 gnd.n6608 gnd.n721 19.3944
R8567 gnd.n6608 gnd.n719 19.3944
R8568 gnd.n6612 gnd.n719 19.3944
R8569 gnd.n6612 gnd.n715 19.3944
R8570 gnd.n6618 gnd.n715 19.3944
R8571 gnd.n6618 gnd.n713 19.3944
R8572 gnd.n6622 gnd.n713 19.3944
R8573 gnd.n6622 gnd.n709 19.3944
R8574 gnd.n6628 gnd.n709 19.3944
R8575 gnd.n6628 gnd.n707 19.3944
R8576 gnd.n6632 gnd.n707 19.3944
R8577 gnd.n6632 gnd.n703 19.3944
R8578 gnd.n6638 gnd.n703 19.3944
R8579 gnd.n6638 gnd.n701 19.3944
R8580 gnd.n6642 gnd.n701 19.3944
R8581 gnd.n6642 gnd.n697 19.3944
R8582 gnd.n6648 gnd.n697 19.3944
R8583 gnd.n6648 gnd.n695 19.3944
R8584 gnd.n6652 gnd.n695 19.3944
R8585 gnd.n6652 gnd.n691 19.3944
R8586 gnd.n6658 gnd.n691 19.3944
R8587 gnd.n6658 gnd.n689 19.3944
R8588 gnd.n6662 gnd.n689 19.3944
R8589 gnd.n6662 gnd.n685 19.3944
R8590 gnd.n6668 gnd.n685 19.3944
R8591 gnd.n6668 gnd.n683 19.3944
R8592 gnd.n6672 gnd.n683 19.3944
R8593 gnd.n6672 gnd.n679 19.3944
R8594 gnd.n6678 gnd.n679 19.3944
R8595 gnd.n6678 gnd.n677 19.3944
R8596 gnd.n6682 gnd.n677 19.3944
R8597 gnd.n6682 gnd.n673 19.3944
R8598 gnd.n6688 gnd.n673 19.3944
R8599 gnd.n6688 gnd.n671 19.3944
R8600 gnd.n6692 gnd.n671 19.3944
R8601 gnd.n6692 gnd.n667 19.3944
R8602 gnd.n6698 gnd.n667 19.3944
R8603 gnd.n6698 gnd.n665 19.3944
R8604 gnd.n6702 gnd.n665 19.3944
R8605 gnd.n6702 gnd.n661 19.3944
R8606 gnd.n6708 gnd.n661 19.3944
R8607 gnd.n6708 gnd.n659 19.3944
R8608 gnd.n6712 gnd.n659 19.3944
R8609 gnd.n6712 gnd.n655 19.3944
R8610 gnd.n6718 gnd.n655 19.3944
R8611 gnd.n6718 gnd.n653 19.3944
R8612 gnd.n6722 gnd.n653 19.3944
R8613 gnd.n6722 gnd.n649 19.3944
R8614 gnd.n6728 gnd.n649 19.3944
R8615 gnd.n6728 gnd.n647 19.3944
R8616 gnd.n6732 gnd.n647 19.3944
R8617 gnd.n6732 gnd.n643 19.3944
R8618 gnd.n6738 gnd.n643 19.3944
R8619 gnd.n6738 gnd.n641 19.3944
R8620 gnd.n6742 gnd.n641 19.3944
R8621 gnd.n6742 gnd.n637 19.3944
R8622 gnd.n6748 gnd.n637 19.3944
R8623 gnd.n6748 gnd.n635 19.3944
R8624 gnd.n6752 gnd.n635 19.3944
R8625 gnd.n6752 gnd.n631 19.3944
R8626 gnd.n6758 gnd.n631 19.3944
R8627 gnd.n6758 gnd.n629 19.3944
R8628 gnd.n6762 gnd.n629 19.3944
R8629 gnd.n6762 gnd.n625 19.3944
R8630 gnd.n6768 gnd.n625 19.3944
R8631 gnd.n6768 gnd.n623 19.3944
R8632 gnd.n6772 gnd.n623 19.3944
R8633 gnd.n6772 gnd.n619 19.3944
R8634 gnd.n6778 gnd.n619 19.3944
R8635 gnd.n6778 gnd.n617 19.3944
R8636 gnd.n6782 gnd.n617 19.3944
R8637 gnd.n6782 gnd.n613 19.3944
R8638 gnd.n6788 gnd.n613 19.3944
R8639 gnd.n6788 gnd.n611 19.3944
R8640 gnd.n6792 gnd.n611 19.3944
R8641 gnd.n6792 gnd.n607 19.3944
R8642 gnd.n6798 gnd.n607 19.3944
R8643 gnd.n6798 gnd.n605 19.3944
R8644 gnd.n6802 gnd.n605 19.3944
R8645 gnd.n6802 gnd.n601 19.3944
R8646 gnd.n6808 gnd.n601 19.3944
R8647 gnd.n6808 gnd.n599 19.3944
R8648 gnd.n6812 gnd.n599 19.3944
R8649 gnd.n6812 gnd.n595 19.3944
R8650 gnd.n6818 gnd.n595 19.3944
R8651 gnd.n6818 gnd.n593 19.3944
R8652 gnd.n6822 gnd.n593 19.3944
R8653 gnd.n6822 gnd.n589 19.3944
R8654 gnd.n6828 gnd.n589 19.3944
R8655 gnd.n6828 gnd.n587 19.3944
R8656 gnd.n6832 gnd.n587 19.3944
R8657 gnd.n6832 gnd.n583 19.3944
R8658 gnd.n6838 gnd.n583 19.3944
R8659 gnd.n6838 gnd.n581 19.3944
R8660 gnd.n6842 gnd.n581 19.3944
R8661 gnd.n6842 gnd.n577 19.3944
R8662 gnd.n6848 gnd.n577 19.3944
R8663 gnd.n6848 gnd.n575 19.3944
R8664 gnd.n6852 gnd.n575 19.3944
R8665 gnd.n6852 gnd.n571 19.3944
R8666 gnd.n6858 gnd.n571 19.3944
R8667 gnd.n6858 gnd.n569 19.3944
R8668 gnd.n6862 gnd.n569 19.3944
R8669 gnd.n6862 gnd.n565 19.3944
R8670 gnd.n6868 gnd.n565 19.3944
R8671 gnd.n6868 gnd.n563 19.3944
R8672 gnd.n6872 gnd.n563 19.3944
R8673 gnd.n6872 gnd.n559 19.3944
R8674 gnd.n6878 gnd.n559 19.3944
R8675 gnd.n6878 gnd.n557 19.3944
R8676 gnd.n6882 gnd.n557 19.3944
R8677 gnd.n6882 gnd.n553 19.3944
R8678 gnd.n6888 gnd.n553 19.3944
R8679 gnd.n6888 gnd.n551 19.3944
R8680 gnd.n6893 gnd.n551 19.3944
R8681 gnd.n6893 gnd.n547 19.3944
R8682 gnd.n6899 gnd.n547 19.3944
R8683 gnd.n6900 gnd.n6899 19.3944
R8684 gnd.n5513 gnd.n5510 19.3944
R8685 gnd.n5513 gnd.n5509 19.3944
R8686 gnd.n5519 gnd.n5509 19.3944
R8687 gnd.n5519 gnd.n5507 19.3944
R8688 gnd.n5523 gnd.n5507 19.3944
R8689 gnd.n5523 gnd.n5505 19.3944
R8690 gnd.n5529 gnd.n5505 19.3944
R8691 gnd.n5529 gnd.n5503 19.3944
R8692 gnd.n5533 gnd.n5503 19.3944
R8693 gnd.n5533 gnd.n5501 19.3944
R8694 gnd.n5539 gnd.n5501 19.3944
R8695 gnd.n5539 gnd.n5499 19.3944
R8696 gnd.n5543 gnd.n5499 19.3944
R8697 gnd.n5543 gnd.n5497 19.3944
R8698 gnd.n5549 gnd.n5497 19.3944
R8699 gnd.n5549 gnd.n5495 19.3944
R8700 gnd.n5556 gnd.n5495 19.3944
R8701 gnd.n5562 gnd.n5493 19.3944
R8702 gnd.n5562 gnd.n5491 19.3944
R8703 gnd.n5566 gnd.n5491 19.3944
R8704 gnd.n5566 gnd.n5489 19.3944
R8705 gnd.n5572 gnd.n5489 19.3944
R8706 gnd.n5572 gnd.n5487 19.3944
R8707 gnd.n5577 gnd.n5487 19.3944
R8708 gnd.n5585 gnd.n1786 19.3944
R8709 gnd.n5585 gnd.n1784 19.3944
R8710 gnd.n5589 gnd.n1784 19.3944
R8711 gnd.n5589 gnd.n1782 19.3944
R8712 gnd.n5595 gnd.n1782 19.3944
R8713 gnd.n5595 gnd.n1780 19.3944
R8714 gnd.n5599 gnd.n1780 19.3944
R8715 gnd.n5599 gnd.n1778 19.3944
R8716 gnd.n5611 gnd.n1776 19.3944
R8717 gnd.n5611 gnd.n1774 19.3944
R8718 gnd.n5617 gnd.n1774 19.3944
R8719 gnd.n5617 gnd.n1772 19.3944
R8720 gnd.n5621 gnd.n1772 19.3944
R8721 gnd.n5621 gnd.n1770 19.3944
R8722 gnd.n5627 gnd.n1770 19.3944
R8723 gnd.n5627 gnd.n1768 19.3944
R8724 gnd.n5631 gnd.n1768 19.3944
R8725 gnd.n5631 gnd.n1766 19.3944
R8726 gnd.n5637 gnd.n1766 19.3944
R8727 gnd.n5637 gnd.n1764 19.3944
R8728 gnd.n5641 gnd.n1764 19.3944
R8729 gnd.n5641 gnd.n1762 19.3944
R8730 gnd.n5647 gnd.n1762 19.3944
R8731 gnd.n5647 gnd.n1760 19.3944
R8732 gnd.n5652 gnd.n1760 19.3944
R8733 gnd.n5652 gnd.n1758 19.3944
R8734 gnd.n5665 gnd.n1751 19.3944
R8735 gnd.n5666 gnd.n5665 19.3944
R8736 gnd.n5667 gnd.n5666 19.3944
R8737 gnd.n5667 gnd.n1746 19.3944
R8738 gnd.n5679 gnd.n1746 19.3944
R8739 gnd.n5680 gnd.n5679 19.3944
R8740 gnd.n5681 gnd.n5680 19.3944
R8741 gnd.n5682 gnd.n5681 19.3944
R8742 gnd.n5684 gnd.n5682 19.3944
R8743 gnd.n5684 gnd.n1734 19.3944
R8744 gnd.n5744 gnd.n1734 19.3944
R8745 gnd.n5745 gnd.n5744 19.3944
R8746 gnd.n5747 gnd.n5745 19.3944
R8747 gnd.n5747 gnd.n1728 19.3944
R8748 gnd.n5769 gnd.n1728 19.3944
R8749 gnd.n5770 gnd.n5769 19.3944
R8750 gnd.n5771 gnd.n5770 19.3944
R8751 gnd.n5774 gnd.n5771 19.3944
R8752 gnd.n5774 gnd.n1726 19.3944
R8753 gnd.n5782 gnd.n1726 19.3944
R8754 gnd.n5783 gnd.n5782 19.3944
R8755 gnd.n5787 gnd.n5783 19.3944
R8756 gnd.n5787 gnd.n5784 19.3944
R8757 gnd.n5784 gnd.n399 19.3944
R8758 gnd.n7142 gnd.n399 19.3944
R8759 gnd.n7142 gnd.n395 19.3944
R8760 gnd.n7154 gnd.n395 19.3944
R8761 gnd.n7155 gnd.n7154 19.3944
R8762 gnd.n7157 gnd.n7155 19.3944
R8763 gnd.n7157 gnd.n390 19.3944
R8764 gnd.n7169 gnd.n390 19.3944
R8765 gnd.n7170 gnd.n7169 19.3944
R8766 gnd.n7172 gnd.n7170 19.3944
R8767 gnd.n7172 gnd.n386 19.3944
R8768 gnd.n7268 gnd.n386 19.3944
R8769 gnd.n7269 gnd.n7268 19.3944
R8770 gnd.n7272 gnd.n7269 19.3944
R8771 gnd.n7273 gnd.n7272 19.3944
R8772 gnd.n7275 gnd.n7273 19.3944
R8773 gnd.n7276 gnd.n7275 19.3944
R8774 gnd.n7278 gnd.n7276 19.3944
R8775 gnd.n7279 gnd.n7278 19.3944
R8776 gnd.n5662 gnd.n1624 19.3944
R8777 gnd.n5850 gnd.n1624 19.3944
R8778 gnd.n5850 gnd.n5849 19.3944
R8779 gnd.n5849 gnd.n5848 19.3944
R8780 gnd.n5848 gnd.n1628 19.3944
R8781 gnd.n5838 gnd.n1628 19.3944
R8782 gnd.n5838 gnd.n5837 19.3944
R8783 gnd.n5837 gnd.n5836 19.3944
R8784 gnd.n5836 gnd.n1648 19.3944
R8785 gnd.n5826 gnd.n1648 19.3944
R8786 gnd.n5826 gnd.n5825 19.3944
R8787 gnd.n5825 gnd.n5824 19.3944
R8788 gnd.n5824 gnd.n1669 19.3944
R8789 gnd.n5814 gnd.n1669 19.3944
R8790 gnd.n5814 gnd.n5813 19.3944
R8791 gnd.n5813 gnd.n5812 19.3944
R8792 gnd.n5812 gnd.n1688 19.3944
R8793 gnd.n5776 gnd.n1688 19.3944
R8794 gnd.n5779 gnd.n5776 19.3944
R8795 gnd.n5779 gnd.n1724 19.3944
R8796 gnd.n5790 gnd.n1724 19.3944
R8797 gnd.n5790 gnd.n5789 19.3944
R8798 gnd.n5789 gnd.n401 19.3944
R8799 gnd.n7139 gnd.n401 19.3944
R8800 gnd.n7139 gnd.n92 19.3944
R8801 gnd.n7329 gnd.n92 19.3944
R8802 gnd.n7329 gnd.n7328 19.3944
R8803 gnd.n7328 gnd.n7327 19.3944
R8804 gnd.n7327 gnd.n96 19.3944
R8805 gnd.n7317 gnd.n96 19.3944
R8806 gnd.n7317 gnd.n7316 19.3944
R8807 gnd.n7316 gnd.n7315 19.3944
R8808 gnd.n7315 gnd.n115 19.3944
R8809 gnd.n7305 gnd.n115 19.3944
R8810 gnd.n7305 gnd.n7304 19.3944
R8811 gnd.n7304 gnd.n7303 19.3944
R8812 gnd.n7303 gnd.n136 19.3944
R8813 gnd.n7293 gnd.n136 19.3944
R8814 gnd.n7293 gnd.n7292 19.3944
R8815 gnd.n7292 gnd.n7291 19.3944
R8816 gnd.n7291 gnd.n157 19.3944
R8817 gnd.n7281 gnd.n157 19.3944
R8818 gnd.n334 gnd.n194 19.3944
R8819 gnd.n338 gnd.n194 19.3944
R8820 gnd.n338 gnd.n192 19.3944
R8821 gnd.n344 gnd.n192 19.3944
R8822 gnd.n344 gnd.n190 19.3944
R8823 gnd.n348 gnd.n190 19.3944
R8824 gnd.n348 gnd.n188 19.3944
R8825 gnd.n354 gnd.n188 19.3944
R8826 gnd.n354 gnd.n186 19.3944
R8827 gnd.n358 gnd.n186 19.3944
R8828 gnd.n358 gnd.n184 19.3944
R8829 gnd.n364 gnd.n184 19.3944
R8830 gnd.n364 gnd.n182 19.3944
R8831 gnd.n368 gnd.n182 19.3944
R8832 gnd.n368 gnd.n180 19.3944
R8833 gnd.n374 gnd.n180 19.3944
R8834 gnd.n374 gnd.n178 19.3944
R8835 gnd.n378 gnd.n178 19.3944
R8836 gnd.n284 gnd.n216 19.3944
R8837 gnd.n288 gnd.n216 19.3944
R8838 gnd.n288 gnd.n214 19.3944
R8839 gnd.n294 gnd.n214 19.3944
R8840 gnd.n294 gnd.n212 19.3944
R8841 gnd.n298 gnd.n212 19.3944
R8842 gnd.n298 gnd.n210 19.3944
R8843 gnd.n304 gnd.n210 19.3944
R8844 gnd.n304 gnd.n208 19.3944
R8845 gnd.n308 gnd.n208 19.3944
R8846 gnd.n308 gnd.n206 19.3944
R8847 gnd.n314 gnd.n206 19.3944
R8848 gnd.n314 gnd.n204 19.3944
R8849 gnd.n318 gnd.n204 19.3944
R8850 gnd.n318 gnd.n202 19.3944
R8851 gnd.n324 gnd.n202 19.3944
R8852 gnd.n324 gnd.n200 19.3944
R8853 gnd.n328 gnd.n200 19.3944
R8854 gnd.n238 gnd.n237 19.3944
R8855 gnd.n243 gnd.n238 19.3944
R8856 gnd.n243 gnd.n234 19.3944
R8857 gnd.n247 gnd.n234 19.3944
R8858 gnd.n247 gnd.n232 19.3944
R8859 gnd.n253 gnd.n232 19.3944
R8860 gnd.n253 gnd.n230 19.3944
R8861 gnd.n257 gnd.n230 19.3944
R8862 gnd.n257 gnd.n228 19.3944
R8863 gnd.n263 gnd.n228 19.3944
R8864 gnd.n263 gnd.n226 19.3944
R8865 gnd.n267 gnd.n226 19.3944
R8866 gnd.n267 gnd.n224 19.3944
R8867 gnd.n274 gnd.n224 19.3944
R8868 gnd.n274 gnd.n222 19.3944
R8869 gnd.n278 gnd.n222 19.3944
R8870 gnd.n279 gnd.n278 19.3944
R8871 gnd.n7207 gnd.n7206 19.3944
R8872 gnd.n7212 gnd.n7207 19.3944
R8873 gnd.n7212 gnd.n7203 19.3944
R8874 gnd.n7216 gnd.n7203 19.3944
R8875 gnd.n7216 gnd.n7201 19.3944
R8876 gnd.n7222 gnd.n7201 19.3944
R8877 gnd.n7222 gnd.n7199 19.3944
R8878 gnd.n7226 gnd.n7199 19.3944
R8879 gnd.n7226 gnd.n7197 19.3944
R8880 gnd.n7232 gnd.n7197 19.3944
R8881 gnd.n7232 gnd.n7195 19.3944
R8882 gnd.n7236 gnd.n7195 19.3944
R8883 gnd.n7236 gnd.n7193 19.3944
R8884 gnd.n7242 gnd.n7193 19.3944
R8885 gnd.n7242 gnd.n7191 19.3944
R8886 gnd.n7246 gnd.n7191 19.3944
R8887 gnd.n5124 gnd.n5123 19.3944
R8888 gnd.n5123 gnd.n1750 19.3944
R8889 gnd.n5671 gnd.n1750 19.3944
R8890 gnd.n5671 gnd.n1748 19.3944
R8891 gnd.n5675 gnd.n1748 19.3944
R8892 gnd.n5675 gnd.n1742 19.3944
R8893 gnd.n5695 gnd.n1742 19.3944
R8894 gnd.n5695 gnd.n1743 19.3944
R8895 gnd.n5691 gnd.n1743 19.3944
R8896 gnd.n5691 gnd.n5690 19.3944
R8897 gnd.n5690 gnd.n5689 19.3944
R8898 gnd.n5689 gnd.n1733 19.3944
R8899 gnd.n5751 gnd.n1733 19.3944
R8900 gnd.n5751 gnd.n1730 19.3944
R8901 gnd.n5765 gnd.n1730 19.3944
R8902 gnd.n5765 gnd.n1731 19.3944
R8903 gnd.n5761 gnd.n1731 19.3944
R8904 gnd.n5761 gnd.n5760 19.3944
R8905 gnd.n5760 gnd.n5759 19.3944
R8906 gnd.n5759 gnd.n5757 19.3944
R8907 gnd.n5757 gnd.n64 19.3944
R8908 gnd.n7342 gnd.n64 19.3944
R8909 gnd.n7342 gnd.n7341 19.3944
R8910 gnd.n7341 gnd.n67 19.3944
R8911 gnd.n7146 gnd.n67 19.3944
R8912 gnd.n7146 gnd.n396 19.3944
R8913 gnd.n7150 gnd.n396 19.3944
R8914 gnd.n7150 gnd.n394 19.3944
R8915 gnd.n7161 gnd.n394 19.3944
R8916 gnd.n7161 gnd.n392 19.3944
R8917 gnd.n7165 gnd.n392 19.3944
R8918 gnd.n7165 gnd.n389 19.3944
R8919 gnd.n7176 gnd.n389 19.3944
R8920 gnd.n7176 gnd.n387 19.3944
R8921 gnd.n7264 gnd.n387 19.3944
R8922 gnd.n7264 gnd.n7263 19.3944
R8923 gnd.n7263 gnd.n7262 19.3944
R8924 gnd.n7262 gnd.n7260 19.3944
R8925 gnd.n7260 gnd.n7259 19.3944
R8926 gnd.n7259 gnd.n7257 19.3944
R8927 gnd.n7257 gnd.n7256 19.3944
R8928 gnd.n7256 gnd.n7254 19.3944
R8929 gnd.n5856 gnd.n5855 19.3944
R8930 gnd.n5855 gnd.n5854 19.3944
R8931 gnd.n5854 gnd.n1616 19.3944
R8932 gnd.n5844 gnd.n1616 19.3944
R8933 gnd.n5844 gnd.n5843 19.3944
R8934 gnd.n5843 gnd.n5842 19.3944
R8935 gnd.n5842 gnd.n1639 19.3944
R8936 gnd.n5832 gnd.n1639 19.3944
R8937 gnd.n5832 gnd.n5831 19.3944
R8938 gnd.n5831 gnd.n5830 19.3944
R8939 gnd.n5830 gnd.n1659 19.3944
R8940 gnd.n5820 gnd.n1659 19.3944
R8941 gnd.n5820 gnd.n5819 19.3944
R8942 gnd.n5819 gnd.n5818 19.3944
R8943 gnd.n5818 gnd.n1679 19.3944
R8944 gnd.n5808 gnd.n1679 19.3944
R8945 gnd.n1696 gnd.n1695 19.3944
R8946 gnd.n5795 gnd.n5794 19.3944
R8947 gnd.n1713 gnd.n1712 19.3944
R8948 gnd.n7337 gnd.n7336 19.3944
R8949 gnd.n7333 gnd.n76 19.3944
R8950 gnd.n7333 gnd.n83 19.3944
R8951 gnd.n7323 gnd.n83 19.3944
R8952 gnd.n7323 gnd.n7322 19.3944
R8953 gnd.n7322 gnd.n7321 19.3944
R8954 gnd.n7321 gnd.n106 19.3944
R8955 gnd.n7311 gnd.n106 19.3944
R8956 gnd.n7311 gnd.n7310 19.3944
R8957 gnd.n7310 gnd.n7309 19.3944
R8958 gnd.n7309 gnd.n126 19.3944
R8959 gnd.n7299 gnd.n126 19.3944
R8960 gnd.n7299 gnd.n7298 19.3944
R8961 gnd.n7298 gnd.n7297 19.3944
R8962 gnd.n7297 gnd.n147 19.3944
R8963 gnd.n7287 gnd.n147 19.3944
R8964 gnd.n7287 gnd.n7286 19.3944
R8965 gnd.n7286 gnd.n7285 19.3944
R8966 gnd.n6308 gnd.n965 19.3944
R8967 gnd.n2399 gnd.n965 19.3944
R8968 gnd.n2413 gnd.n2399 19.3944
R8969 gnd.n2413 gnd.n2412 19.3944
R8970 gnd.n2412 gnd.n2411 19.3944
R8971 gnd.n2411 gnd.n2404 19.3944
R8972 gnd.n2407 gnd.n2404 19.3944
R8973 gnd.n2407 gnd.n2366 19.3944
R8974 gnd.n4336 gnd.n2366 19.3944
R8975 gnd.n4336 gnd.n2367 19.3944
R8976 gnd.n2380 gnd.n2379 19.3944
R8977 gnd.n4323 gnd.n4322 19.3944
R8978 gnd.n4319 gnd.n4318 19.3944
R8979 gnd.n2386 gnd.n2385 19.3944
R8980 gnd.n2382 gnd.n2359 19.3944
R8981 gnd.n4360 gnd.n2359 19.3944
R8982 gnd.n4360 gnd.n4359 19.3944
R8983 gnd.n4359 gnd.n4358 19.3944
R8984 gnd.n4358 gnd.n4343 19.3944
R8985 gnd.n4354 gnd.n4343 19.3944
R8986 gnd.n4354 gnd.n4353 19.3944
R8987 gnd.n4353 gnd.n4352 19.3944
R8988 gnd.n4352 gnd.n4350 19.3944
R8989 gnd.n4350 gnd.n2337 19.3944
R8990 gnd.n4413 gnd.n2337 19.3944
R8991 gnd.n4413 gnd.n2335 19.3944
R8992 gnd.n4417 gnd.n2335 19.3944
R8993 gnd.n4417 gnd.n2333 19.3944
R8994 gnd.n4421 gnd.n2333 19.3944
R8995 gnd.n4421 gnd.n2331 19.3944
R8996 gnd.n4425 gnd.n2331 19.3944
R8997 gnd.n4425 gnd.n2329 19.3944
R8998 gnd.n4429 gnd.n2329 19.3944
R8999 gnd.n4429 gnd.n2327 19.3944
R9000 gnd.n4433 gnd.n2327 19.3944
R9001 gnd.n4433 gnd.n2324 19.3944
R9002 gnd.n4439 gnd.n2324 19.3944
R9003 gnd.n4439 gnd.n2322 19.3944
R9004 gnd.n4445 gnd.n2322 19.3944
R9005 gnd.n4445 gnd.n4444 19.3944
R9006 gnd.n4444 gnd.n2296 19.3944
R9007 gnd.n4471 gnd.n2296 19.3944
R9008 gnd.n4471 gnd.n2294 19.3944
R9009 gnd.n4478 gnd.n2294 19.3944
R9010 gnd.n4478 gnd.n4477 19.3944
R9011 gnd.n4477 gnd.n1484 19.3944
R9012 gnd.n5989 gnd.n1484 19.3944
R9013 gnd.n5989 gnd.n5988 19.3944
R9014 gnd.n5988 gnd.n5987 19.3944
R9015 gnd.n5987 gnd.n1488 19.3944
R9016 gnd.n4514 gnd.n1488 19.3944
R9017 gnd.n4514 gnd.n2170 19.3944
R9018 gnd.n4553 gnd.n2170 19.3944
R9019 gnd.n4553 gnd.n2168 19.3944
R9020 gnd.n4557 gnd.n2168 19.3944
R9021 gnd.n4557 gnd.n2152 19.3944
R9022 gnd.n4595 gnd.n2152 19.3944
R9023 gnd.n4595 gnd.n2150 19.3944
R9024 gnd.n4601 gnd.n2150 19.3944
R9025 gnd.n4601 gnd.n4600 19.3944
R9026 gnd.n4600 gnd.n2126 19.3944
R9027 gnd.n4657 gnd.n2126 19.3944
R9028 gnd.n4657 gnd.n2124 19.3944
R9029 gnd.n4661 gnd.n2124 19.3944
R9030 gnd.n4661 gnd.n2108 19.3944
R9031 gnd.n4685 gnd.n2108 19.3944
R9032 gnd.n4685 gnd.n2106 19.3944
R9033 gnd.n4691 gnd.n2106 19.3944
R9034 gnd.n4691 gnd.n4690 19.3944
R9035 gnd.n4690 gnd.n2075 19.3944
R9036 gnd.n4735 gnd.n2075 19.3944
R9037 gnd.n4735 gnd.n2073 19.3944
R9038 gnd.n4739 gnd.n2073 19.3944
R9039 gnd.n4739 gnd.n2052 19.3944
R9040 gnd.n4775 gnd.n2052 19.3944
R9041 gnd.n4775 gnd.n2050 19.3944
R9042 gnd.n4779 gnd.n2050 19.3944
R9043 gnd.n4779 gnd.n2030 19.3944
R9044 gnd.n4832 gnd.n2030 19.3944
R9045 gnd.n4832 gnd.n2028 19.3944
R9046 gnd.n4836 gnd.n2028 19.3944
R9047 gnd.n4836 gnd.n2010 19.3944
R9048 gnd.n4857 gnd.n2010 19.3944
R9049 gnd.n4857 gnd.n2008 19.3944
R9050 gnd.n4861 gnd.n2008 19.3944
R9051 gnd.n4861 gnd.n1990 19.3944
R9052 gnd.n4917 gnd.n1990 19.3944
R9053 gnd.n4917 gnd.n1988 19.3944
R9054 gnd.n4921 gnd.n1988 19.3944
R9055 gnd.n4921 gnd.n1968 19.3944
R9056 gnd.n4946 gnd.n1968 19.3944
R9057 gnd.n4946 gnd.n1966 19.3944
R9058 gnd.n4952 gnd.n1966 19.3944
R9059 gnd.n4952 gnd.n4951 19.3944
R9060 gnd.n4951 gnd.n1940 19.3944
R9061 gnd.n4997 gnd.n1940 19.3944
R9062 gnd.n4997 gnd.n1938 19.3944
R9063 gnd.n5001 gnd.n1938 19.3944
R9064 gnd.n5001 gnd.n1920 19.3944
R9065 gnd.n5023 gnd.n1920 19.3944
R9066 gnd.n5023 gnd.n1918 19.3944
R9067 gnd.n5029 gnd.n1918 19.3944
R9068 gnd.n5029 gnd.n5028 19.3944
R9069 gnd.n5028 gnd.n1890 19.3944
R9070 gnd.n5067 gnd.n1890 19.3944
R9071 gnd.n5067 gnd.n1888 19.3944
R9072 gnd.n5074 gnd.n1888 19.3944
R9073 gnd.n5074 gnd.n5073 19.3944
R9074 gnd.n5073 gnd.n1839 19.3944
R9075 gnd.n5320 gnd.n1839 19.3944
R9076 gnd.n5320 gnd.n5319 19.3944
R9077 gnd.n5319 gnd.n5318 19.3944
R9078 gnd.n5318 gnd.n1843 19.3944
R9079 gnd.n1850 gnd.n1843 19.3944
R9080 gnd.n5308 gnd.n1850 19.3944
R9081 gnd.n5308 gnd.n5307 19.3944
R9082 gnd.n5307 gnd.n5306 19.3944
R9083 gnd.n5306 gnd.n1858 19.3944
R9084 gnd.n1858 gnd.n1591 19.3944
R9085 gnd.n5871 gnd.n1591 19.3944
R9086 gnd.n5871 gnd.n5870 19.3944
R9087 gnd.n5870 gnd.n5869 19.3944
R9088 gnd.n5869 gnd.n1595 19.3944
R9089 gnd.n5863 gnd.n1595 19.3944
R9090 gnd.n5863 gnd.n5862 19.3944
R9091 gnd.n5862 gnd.n5861 19.3944
R9092 gnd.n5861 gnd.n1604 19.3944
R9093 gnd.n5707 gnd.n1604 19.3944
R9094 gnd.n5707 gnd.n5704 19.3944
R9095 gnd.n5711 gnd.n5704 19.3944
R9096 gnd.n5711 gnd.n5702 19.3944
R9097 gnd.n5715 gnd.n5702 19.3944
R9098 gnd.n5715 gnd.n5700 19.3944
R9099 gnd.n5719 gnd.n5700 19.3944
R9100 gnd.n5719 gnd.n1740 19.3944
R9101 gnd.n5723 gnd.n1740 19.3944
R9102 gnd.n5723 gnd.n1738 19.3944
R9103 gnd.n5739 gnd.n1738 19.3944
R9104 gnd.n5739 gnd.n5738 19.3944
R9105 gnd.n5738 gnd.n5737 19.3944
R9106 gnd.n5737 gnd.n5729 19.3944
R9107 gnd.n5733 gnd.n5729 19.3944
R9108 gnd.n5733 gnd.n5732 19.3944
R9109 gnd.n5803 gnd.n5802 19.3944
R9110 gnd.n5800 gnd.n1703 19.3944
R9111 gnd.n1720 gnd.n1719 19.3944
R9112 gnd.n7134 gnd.n404 19.3944
R9113 gnd.n7132 gnd.n7131 19.3944
R9114 gnd.n7131 gnd.n406 19.3944
R9115 gnd.n7127 gnd.n406 19.3944
R9116 gnd.n7127 gnd.n7126 19.3944
R9117 gnd.n7126 gnd.n7125 19.3944
R9118 gnd.n7125 gnd.n412 19.3944
R9119 gnd.n7121 gnd.n412 19.3944
R9120 gnd.n7121 gnd.n7120 19.3944
R9121 gnd.n7120 gnd.n7119 19.3944
R9122 gnd.n7119 gnd.n418 19.3944
R9123 gnd.n4214 gnd.n2448 19.3944
R9124 gnd.n4209 gnd.n2448 19.3944
R9125 gnd.n4209 gnd.n4208 19.3944
R9126 gnd.n4208 gnd.n4207 19.3944
R9127 gnd.n4207 gnd.n4204 19.3944
R9128 gnd.n4204 gnd.n4203 19.3944
R9129 gnd.n4203 gnd.n4200 19.3944
R9130 gnd.n4200 gnd.n4199 19.3944
R9131 gnd.n4199 gnd.n4196 19.3944
R9132 gnd.n4196 gnd.n4195 19.3944
R9133 gnd.n4195 gnd.n4192 19.3944
R9134 gnd.n4192 gnd.n4191 19.3944
R9135 gnd.n4191 gnd.n4188 19.3944
R9136 gnd.n4188 gnd.n4187 19.3944
R9137 gnd.n4187 gnd.n4184 19.3944
R9138 gnd.n4184 gnd.n4183 19.3944
R9139 gnd.n4183 gnd.n4180 19.3944
R9140 gnd.n4178 gnd.n4175 19.3944
R9141 gnd.n4175 gnd.n4174 19.3944
R9142 gnd.n4174 gnd.n4171 19.3944
R9143 gnd.n4171 gnd.n4170 19.3944
R9144 gnd.n4170 gnd.n4167 19.3944
R9145 gnd.n4167 gnd.n4166 19.3944
R9146 gnd.n4166 gnd.n4163 19.3944
R9147 gnd.n4163 gnd.n4162 19.3944
R9148 gnd.n4162 gnd.n4159 19.3944
R9149 gnd.n4159 gnd.n4158 19.3944
R9150 gnd.n4158 gnd.n4155 19.3944
R9151 gnd.n4155 gnd.n4154 19.3944
R9152 gnd.n4154 gnd.n4151 19.3944
R9153 gnd.n4151 gnd.n4150 19.3944
R9154 gnd.n4150 gnd.n4147 19.3944
R9155 gnd.n4147 gnd.n4146 19.3944
R9156 gnd.n4146 gnd.n4143 19.3944
R9157 gnd.n4143 gnd.n4142 19.3944
R9158 gnd.n4138 gnd.n4135 19.3944
R9159 gnd.n4135 gnd.n4134 19.3944
R9160 gnd.n4134 gnd.n4131 19.3944
R9161 gnd.n4131 gnd.n4130 19.3944
R9162 gnd.n4130 gnd.n4127 19.3944
R9163 gnd.n4127 gnd.n4126 19.3944
R9164 gnd.n4126 gnd.n4123 19.3944
R9165 gnd.n4123 gnd.n4122 19.3944
R9166 gnd.n4122 gnd.n4119 19.3944
R9167 gnd.n4119 gnd.n4118 19.3944
R9168 gnd.n4118 gnd.n4115 19.3944
R9169 gnd.n4115 gnd.n4114 19.3944
R9170 gnd.n4114 gnd.n4111 19.3944
R9171 gnd.n4111 gnd.n4110 19.3944
R9172 gnd.n4110 gnd.n4107 19.3944
R9173 gnd.n4107 gnd.n4106 19.3944
R9174 gnd.n4106 gnd.n4103 19.3944
R9175 gnd.n4103 gnd.n4102 19.3944
R9176 gnd.n4088 gnd.n4087 19.3944
R9177 gnd.n4087 gnd.n4084 19.3944
R9178 gnd.n4084 gnd.n4083 19.3944
R9179 gnd.n4083 gnd.n4080 19.3944
R9180 gnd.n4080 gnd.n4079 19.3944
R9181 gnd.n4079 gnd.n4076 19.3944
R9182 gnd.n4076 gnd.n4075 19.3944
R9183 gnd.n4075 gnd.n4072 19.3944
R9184 gnd.n4072 gnd.n4071 19.3944
R9185 gnd.n4071 gnd.n4068 19.3944
R9186 gnd.n4068 gnd.n4067 19.3944
R9187 gnd.n4067 gnd.n4064 19.3944
R9188 gnd.n4064 gnd.n4063 19.3944
R9189 gnd.n4063 gnd.n4060 19.3944
R9190 gnd.n4060 gnd.n4059 19.3944
R9191 gnd.n4059 gnd.n4056 19.3944
R9192 gnd.n4050 gnd.n4048 19.3944
R9193 gnd.n4048 gnd.n4047 19.3944
R9194 gnd.n4047 gnd.n4045 19.3944
R9195 gnd.n4045 gnd.n4044 19.3944
R9196 gnd.n4044 gnd.n4042 19.3944
R9197 gnd.n4042 gnd.n4041 19.3944
R9198 gnd.n4041 gnd.n2418 19.3944
R9199 gnd.n4254 gnd.n2418 19.3944
R9200 gnd.n4254 gnd.n2416 19.3944
R9201 gnd.n4258 gnd.n2416 19.3944
R9202 gnd.n4258 gnd.n2395 19.3944
R9203 gnd.n4269 gnd.n2395 19.3944
R9204 gnd.n4269 gnd.n2393 19.3944
R9205 gnd.n4276 gnd.n2393 19.3944
R9206 gnd.n4276 gnd.n4275 19.3944
R9207 gnd.n4275 gnd.n2373 19.3944
R9208 gnd.n4330 gnd.n2373 19.3944
R9209 gnd.n4330 gnd.n4329 19.3944
R9210 gnd.n4329 gnd.n4328 19.3944
R9211 gnd.n4328 gnd.n2377 19.3944
R9212 gnd.n4294 gnd.n2377 19.3944
R9213 gnd.n4294 gnd.n2389 19.3944
R9214 gnd.n4313 gnd.n2389 19.3944
R9215 gnd.n4313 gnd.n2390 19.3944
R9216 gnd.n4309 gnd.n2390 19.3944
R9217 gnd.n4309 gnd.n2355 19.3944
R9218 gnd.n4365 gnd.n2355 19.3944
R9219 gnd.n4365 gnd.n2353 19.3944
R9220 gnd.n4369 gnd.n2353 19.3944
R9221 gnd.n4369 gnd.n2349 19.3944
R9222 gnd.n4379 gnd.n2349 19.3944
R9223 gnd.n4379 gnd.n2347 19.3944
R9224 gnd.n4383 gnd.n2347 19.3944
R9225 gnd.n4383 gnd.n2340 19.3944
R9226 gnd.n4407 gnd.n2340 19.3944
R9227 gnd.n4407 gnd.n2341 19.3944
R9228 gnd.n4403 gnd.n2341 19.3944
R9229 gnd.n4403 gnd.n4402 19.3944
R9230 gnd.n4402 gnd.n4401 19.3944
R9231 gnd.n4401 gnd.n1146 19.3944
R9232 gnd.n6190 gnd.n1146 19.3944
R9233 gnd.n6190 gnd.n1147 19.3944
R9234 gnd.n4094 gnd.n2439 19.3944
R9235 gnd.n4223 gnd.n2439 19.3944
R9236 gnd.n4224 gnd.n4223 19.3944
R9237 gnd.n4229 gnd.n4224 19.3944
R9238 gnd.n4229 gnd.n4227 19.3944
R9239 gnd.n4227 gnd.n4226 19.3944
R9240 gnd.n4226 gnd.n2419 19.3944
R9241 gnd.n4250 gnd.n2419 19.3944
R9242 gnd.n4250 gnd.n2396 19.3944
R9243 gnd.n4262 gnd.n2396 19.3944
R9244 gnd.n4263 gnd.n4262 19.3944
R9245 gnd.n4265 gnd.n4263 19.3944
R9246 gnd.n4265 gnd.n2392 19.3944
R9247 gnd.n4281 gnd.n2392 19.3944
R9248 gnd.n4282 gnd.n4281 19.3944
R9249 gnd.n4284 gnd.n4282 19.3944
R9250 gnd.n4287 gnd.n4284 19.3944
R9251 gnd.n4288 gnd.n4287 19.3944
R9252 gnd.n4289 gnd.n4288 19.3944
R9253 gnd.n4290 gnd.n4289 19.3944
R9254 gnd.n4298 gnd.n4290 19.3944
R9255 gnd.n4299 gnd.n4298 19.3944
R9256 gnd.n4300 gnd.n4299 19.3944
R9257 gnd.n4301 gnd.n4300 19.3944
R9258 gnd.n4305 gnd.n4301 19.3944
R9259 gnd.n4305 gnd.n4304 19.3944
R9260 gnd.n4304 gnd.n4303 19.3944
R9261 gnd.n4303 gnd.n2351 19.3944
R9262 gnd.n4373 gnd.n2351 19.3944
R9263 gnd.n4374 gnd.n4373 19.3944
R9264 gnd.n4375 gnd.n4374 19.3944
R9265 gnd.n4375 gnd.n2345 19.3944
R9266 gnd.n4387 gnd.n2345 19.3944
R9267 gnd.n4388 gnd.n4387 19.3944
R9268 gnd.n4389 gnd.n4388 19.3944
R9269 gnd.n4390 gnd.n4389 19.3944
R9270 gnd.n4394 gnd.n4390 19.3944
R9271 gnd.n4395 gnd.n4394 19.3944
R9272 gnd.n4396 gnd.n4395 19.3944
R9273 gnd.n4396 gnd.n1145 19.3944
R9274 gnd.n6194 gnd.n1145 19.3944
R9275 gnd.n6195 gnd.n6194 19.3944
R9276 gnd.n4092 gnd.n4091 19.3944
R9277 gnd.n4092 gnd.n2436 19.3944
R9278 gnd.n4232 gnd.n2436 19.3944
R9279 gnd.n4232 gnd.n4231 19.3944
R9280 gnd.n4231 gnd.n2421 19.3944
R9281 gnd.n4246 gnd.n2421 19.3944
R9282 gnd.n4247 gnd.n4246 19.3944
R9283 gnd.n4247 gnd.n985 19.3944
R9284 gnd.n6297 gnd.n985 19.3944
R9285 gnd.n6297 gnd.n6296 19.3944
R9286 gnd.n6296 gnd.n6295 19.3944
R9287 gnd.n6295 gnd.n989 19.3944
R9288 gnd.n6285 gnd.n989 19.3944
R9289 gnd.n6285 gnd.n6284 19.3944
R9290 gnd.n6284 gnd.n6283 19.3944
R9291 gnd.n6283 gnd.n1010 19.3944
R9292 gnd.n1028 gnd.n1010 19.3944
R9293 gnd.n6271 gnd.n1028 19.3944
R9294 gnd.n6271 gnd.n6270 19.3944
R9295 gnd.n6270 gnd.n6269 19.3944
R9296 gnd.n6269 gnd.n1032 19.3944
R9297 gnd.n6258 gnd.n1032 19.3944
R9298 gnd.n6258 gnd.n6257 19.3944
R9299 gnd.n6257 gnd.n6256 19.3944
R9300 gnd.n6256 gnd.n1048 19.3944
R9301 gnd.n6245 gnd.n1048 19.3944
R9302 gnd.n6245 gnd.n6244 19.3944
R9303 gnd.n6244 gnd.n6243 19.3944
R9304 gnd.n6243 gnd.n1066 19.3944
R9305 gnd.n6233 gnd.n1066 19.3944
R9306 gnd.n6233 gnd.n6232 19.3944
R9307 gnd.n6232 gnd.n6231 19.3944
R9308 gnd.n6231 gnd.n1085 19.3944
R9309 gnd.n6221 gnd.n1085 19.3944
R9310 gnd.n6221 gnd.n6220 19.3944
R9311 gnd.n6220 gnd.n6219 19.3944
R9312 gnd.n6219 gnd.n1106 19.3944
R9313 gnd.n6209 gnd.n1106 19.3944
R9314 gnd.n6209 gnd.n6208 19.3944
R9315 gnd.n6208 gnd.n6207 19.3944
R9316 gnd.n6207 gnd.n1126 19.3944
R9317 gnd.n6197 gnd.n1126 19.3944
R9318 gnd.n1289 gnd.n1288 19.3944
R9319 gnd.n6113 gnd.n1288 19.3944
R9320 gnd.n6113 gnd.n6112 19.3944
R9321 gnd.n6112 gnd.n6111 19.3944
R9322 gnd.n6111 gnd.n6108 19.3944
R9323 gnd.n6108 gnd.n6107 19.3944
R9324 gnd.n6107 gnd.n6104 19.3944
R9325 gnd.n6104 gnd.n6103 19.3944
R9326 gnd.n6103 gnd.n6100 19.3944
R9327 gnd.n6100 gnd.n6099 19.3944
R9328 gnd.n6099 gnd.n6096 19.3944
R9329 gnd.n6096 gnd.n6095 19.3944
R9330 gnd.n6095 gnd.n6092 19.3944
R9331 gnd.n6092 gnd.n6091 19.3944
R9332 gnd.n6091 gnd.n6088 19.3944
R9333 gnd.n6088 gnd.n6087 19.3944
R9334 gnd.n6087 gnd.n6084 19.3944
R9335 gnd.n1391 gnd.n1327 19.3944
R9336 gnd.n1391 gnd.n1388 19.3944
R9337 gnd.n1388 gnd.n1385 19.3944
R9338 gnd.n1385 gnd.n1384 19.3944
R9339 gnd.n1384 gnd.n1381 19.3944
R9340 gnd.n1381 gnd.n1380 19.3944
R9341 gnd.n1380 gnd.n1377 19.3944
R9342 gnd.n1377 gnd.n1376 19.3944
R9343 gnd.n1376 gnd.n1373 19.3944
R9344 gnd.n1373 gnd.n1372 19.3944
R9345 gnd.n1372 gnd.n1369 19.3944
R9346 gnd.n1369 gnd.n1368 19.3944
R9347 gnd.n1368 gnd.n1365 19.3944
R9348 gnd.n1365 gnd.n1364 19.3944
R9349 gnd.n1364 gnd.n1361 19.3944
R9350 gnd.n1361 gnd.n1360 19.3944
R9351 gnd.n1360 gnd.n1357 19.3944
R9352 gnd.n1357 gnd.n1356 19.3944
R9353 gnd.n1413 gnd.n1318 19.3944
R9354 gnd.n1413 gnd.n1410 19.3944
R9355 gnd.n1410 gnd.n1407 19.3944
R9356 gnd.n1407 gnd.n1406 19.3944
R9357 gnd.n1406 gnd.n1403 19.3944
R9358 gnd.n1403 gnd.n1402 19.3944
R9359 gnd.n1402 gnd.n1399 19.3944
R9360 gnd.n1399 gnd.n1398 19.3944
R9361 gnd.n6082 gnd.n6079 19.3944
R9362 gnd.n6079 gnd.n6078 19.3944
R9363 gnd.n6078 gnd.n6075 19.3944
R9364 gnd.n6075 gnd.n6074 19.3944
R9365 gnd.n6074 gnd.n6071 19.3944
R9366 gnd.n6071 gnd.n6070 19.3944
R9367 gnd.n6070 gnd.n6067 19.3944
R9368 gnd.n4218 gnd.n2446 19.3944
R9369 gnd.n4218 gnd.n2429 19.3944
R9370 gnd.n4236 gnd.n2429 19.3944
R9371 gnd.n4236 gnd.n2427 19.3944
R9372 gnd.n4241 gnd.n2427 19.3944
R9373 gnd.n4241 gnd.n974 19.3944
R9374 gnd.n6303 gnd.n974 19.3944
R9375 gnd.n6303 gnd.n6302 19.3944
R9376 gnd.n6302 gnd.n6301 19.3944
R9377 gnd.n6301 gnd.n978 19.3944
R9378 gnd.n6291 gnd.n978 19.3944
R9379 gnd.n6291 gnd.n6290 19.3944
R9380 gnd.n6290 gnd.n6289 19.3944
R9381 gnd.n6289 gnd.n1000 19.3944
R9382 gnd.n6279 gnd.n1000 19.3944
R9383 gnd.n6279 gnd.n6278 19.3944
R9384 gnd.n6276 gnd.n6275 19.3944
R9385 gnd.n6265 gnd.n1038 19.3944
R9386 gnd.n6263 gnd.n6262 19.3944
R9387 gnd.n6252 gnd.n1055 19.3944
R9388 gnd.n6250 gnd.n6249 19.3944
R9389 gnd.n6249 gnd.n1056 19.3944
R9390 gnd.n6239 gnd.n1056 19.3944
R9391 gnd.n6239 gnd.n6238 19.3944
R9392 gnd.n6238 gnd.n6237 19.3944
R9393 gnd.n6237 gnd.n1076 19.3944
R9394 gnd.n6227 gnd.n1076 19.3944
R9395 gnd.n6227 gnd.n6226 19.3944
R9396 gnd.n6226 gnd.n6225 19.3944
R9397 gnd.n6225 gnd.n1096 19.3944
R9398 gnd.n6215 gnd.n1096 19.3944
R9399 gnd.n6215 gnd.n6214 19.3944
R9400 gnd.n6214 gnd.n6213 19.3944
R9401 gnd.n6213 gnd.n1116 19.3944
R9402 gnd.n6203 gnd.n1116 19.3944
R9403 gnd.n6203 gnd.n6202 19.3944
R9404 gnd.n6202 gnd.n6201 19.3944
R9405 gnd.n6479 gnd.n6478 19.3944
R9406 gnd.n6478 gnd.n798 19.3944
R9407 gnd.n6472 gnd.n798 19.3944
R9408 gnd.n6472 gnd.n6471 19.3944
R9409 gnd.n6471 gnd.n6470 19.3944
R9410 gnd.n6470 gnd.n806 19.3944
R9411 gnd.n6464 gnd.n806 19.3944
R9412 gnd.n6464 gnd.n6463 19.3944
R9413 gnd.n6463 gnd.n6462 19.3944
R9414 gnd.n6462 gnd.n814 19.3944
R9415 gnd.n6456 gnd.n814 19.3944
R9416 gnd.n6456 gnd.n6455 19.3944
R9417 gnd.n6455 gnd.n6454 19.3944
R9418 gnd.n6454 gnd.n822 19.3944
R9419 gnd.n6448 gnd.n822 19.3944
R9420 gnd.n6448 gnd.n6447 19.3944
R9421 gnd.n6447 gnd.n6446 19.3944
R9422 gnd.n6446 gnd.n830 19.3944
R9423 gnd.n6440 gnd.n830 19.3944
R9424 gnd.n6440 gnd.n6439 19.3944
R9425 gnd.n6439 gnd.n6438 19.3944
R9426 gnd.n6438 gnd.n838 19.3944
R9427 gnd.n6432 gnd.n838 19.3944
R9428 gnd.n6432 gnd.n6431 19.3944
R9429 gnd.n6431 gnd.n6430 19.3944
R9430 gnd.n6430 gnd.n846 19.3944
R9431 gnd.n6424 gnd.n846 19.3944
R9432 gnd.n6424 gnd.n6423 19.3944
R9433 gnd.n6423 gnd.n6422 19.3944
R9434 gnd.n6422 gnd.n854 19.3944
R9435 gnd.n6416 gnd.n854 19.3944
R9436 gnd.n6416 gnd.n6415 19.3944
R9437 gnd.n6415 gnd.n6414 19.3944
R9438 gnd.n6414 gnd.n862 19.3944
R9439 gnd.n6408 gnd.n862 19.3944
R9440 gnd.n6408 gnd.n6407 19.3944
R9441 gnd.n6407 gnd.n6406 19.3944
R9442 gnd.n6406 gnd.n870 19.3944
R9443 gnd.n6400 gnd.n870 19.3944
R9444 gnd.n6400 gnd.n6399 19.3944
R9445 gnd.n6399 gnd.n6398 19.3944
R9446 gnd.n6398 gnd.n878 19.3944
R9447 gnd.n6392 gnd.n878 19.3944
R9448 gnd.n6392 gnd.n6391 19.3944
R9449 gnd.n6391 gnd.n6390 19.3944
R9450 gnd.n6390 gnd.n886 19.3944
R9451 gnd.n6384 gnd.n886 19.3944
R9452 gnd.n6384 gnd.n6383 19.3944
R9453 gnd.n6383 gnd.n6382 19.3944
R9454 gnd.n6382 gnd.n894 19.3944
R9455 gnd.n6376 gnd.n894 19.3944
R9456 gnd.n6376 gnd.n6375 19.3944
R9457 gnd.n6375 gnd.n6374 19.3944
R9458 gnd.n6374 gnd.n902 19.3944
R9459 gnd.n6368 gnd.n902 19.3944
R9460 gnd.n6368 gnd.n6367 19.3944
R9461 gnd.n6367 gnd.n6366 19.3944
R9462 gnd.n6366 gnd.n910 19.3944
R9463 gnd.n6360 gnd.n910 19.3944
R9464 gnd.n6360 gnd.n6359 19.3944
R9465 gnd.n6359 gnd.n6358 19.3944
R9466 gnd.n6358 gnd.n918 19.3944
R9467 gnd.n6352 gnd.n918 19.3944
R9468 gnd.n6352 gnd.n6351 19.3944
R9469 gnd.n6351 gnd.n6350 19.3944
R9470 gnd.n6350 gnd.n926 19.3944
R9471 gnd.n6344 gnd.n926 19.3944
R9472 gnd.n6344 gnd.n6343 19.3944
R9473 gnd.n6343 gnd.n6342 19.3944
R9474 gnd.n6342 gnd.n934 19.3944
R9475 gnd.n6336 gnd.n934 19.3944
R9476 gnd.n6336 gnd.n6335 19.3944
R9477 gnd.n6335 gnd.n6334 19.3944
R9478 gnd.n6334 gnd.n942 19.3944
R9479 gnd.n6328 gnd.n942 19.3944
R9480 gnd.n6328 gnd.n6327 19.3944
R9481 gnd.n6327 gnd.n6326 19.3944
R9482 gnd.n6326 gnd.n950 19.3944
R9483 gnd.n6320 gnd.n950 19.3944
R9484 gnd.n6320 gnd.n6319 19.3944
R9485 gnd.n6319 gnd.n6318 19.3944
R9486 gnd.n6318 gnd.n958 19.3944
R9487 gnd.n6312 gnd.n958 19.3944
R9488 gnd.n6312 gnd.n6311 19.3944
R9489 gnd.n4450 gnd.n2312 19.3944
R9490 gnd.n4450 gnd.n2309 19.3944
R9491 gnd.n4455 gnd.n2309 19.3944
R9492 gnd.n4455 gnd.n2310 19.3944
R9493 gnd.n2310 gnd.n2288 19.3944
R9494 gnd.n4483 gnd.n2288 19.3944
R9495 gnd.n4483 gnd.n2285 19.3944
R9496 gnd.n4491 gnd.n2285 19.3944
R9497 gnd.n4491 gnd.n2286 19.3944
R9498 gnd.n4487 gnd.n2286 19.3944
R9499 gnd.n4487 gnd.n1495 19.3944
R9500 gnd.n5982 gnd.n1495 19.3944
R9501 gnd.n5982 gnd.n1496 19.3944
R9502 gnd.n5978 gnd.n1496 19.3944
R9503 gnd.n5978 gnd.n5977 19.3944
R9504 gnd.n5977 gnd.n5976 19.3944
R9505 gnd.n5976 gnd.n1502 19.3944
R9506 gnd.n5972 gnd.n1502 19.3944
R9507 gnd.n5972 gnd.n5971 19.3944
R9508 gnd.n5971 gnd.n5970 19.3944
R9509 gnd.n5970 gnd.n1507 19.3944
R9510 gnd.n5966 gnd.n1507 19.3944
R9511 gnd.n5966 gnd.n5965 19.3944
R9512 gnd.n5965 gnd.n5964 19.3944
R9513 gnd.n5964 gnd.n1512 19.3944
R9514 gnd.n5960 gnd.n1512 19.3944
R9515 gnd.n5960 gnd.n5959 19.3944
R9516 gnd.n5959 gnd.n5958 19.3944
R9517 gnd.n5958 gnd.n1517 19.3944
R9518 gnd.n5954 gnd.n1517 19.3944
R9519 gnd.n5954 gnd.n5953 19.3944
R9520 gnd.n5953 gnd.n5952 19.3944
R9521 gnd.n5952 gnd.n1522 19.3944
R9522 gnd.n5948 gnd.n1522 19.3944
R9523 gnd.n5948 gnd.n5947 19.3944
R9524 gnd.n5947 gnd.n5946 19.3944
R9525 gnd.n5946 gnd.n1527 19.3944
R9526 gnd.n5942 gnd.n1527 19.3944
R9527 gnd.n5942 gnd.n5941 19.3944
R9528 gnd.n5941 gnd.n5940 19.3944
R9529 gnd.n5940 gnd.n1532 19.3944
R9530 gnd.n5936 gnd.n1532 19.3944
R9531 gnd.n5936 gnd.n5935 19.3944
R9532 gnd.n5935 gnd.n5934 19.3944
R9533 gnd.n5934 gnd.n1537 19.3944
R9534 gnd.n5930 gnd.n1537 19.3944
R9535 gnd.n5930 gnd.n5929 19.3944
R9536 gnd.n5929 gnd.n5928 19.3944
R9537 gnd.n5928 gnd.n1542 19.3944
R9538 gnd.n5924 gnd.n1542 19.3944
R9539 gnd.n5924 gnd.n5923 19.3944
R9540 gnd.n5923 gnd.n5922 19.3944
R9541 gnd.n5922 gnd.n1547 19.3944
R9542 gnd.n5918 gnd.n1547 19.3944
R9543 gnd.n5918 gnd.n5917 19.3944
R9544 gnd.n5917 gnd.n5916 19.3944
R9545 gnd.n5916 gnd.n1552 19.3944
R9546 gnd.n5912 gnd.n1552 19.3944
R9547 gnd.n5912 gnd.n5911 19.3944
R9548 gnd.n5911 gnd.n5910 19.3944
R9549 gnd.n5910 gnd.n1557 19.3944
R9550 gnd.n5906 gnd.n1557 19.3944
R9551 gnd.n5906 gnd.n5905 19.3944
R9552 gnd.n5905 gnd.n5904 19.3944
R9553 gnd.n5904 gnd.n1562 19.3944
R9554 gnd.n5900 gnd.n1562 19.3944
R9555 gnd.n5900 gnd.n5899 19.3944
R9556 gnd.n5899 gnd.n5898 19.3944
R9557 gnd.n5898 gnd.n1567 19.3944
R9558 gnd.n5894 gnd.n1567 19.3944
R9559 gnd.n5894 gnd.n5893 19.3944
R9560 gnd.n5893 gnd.n5892 19.3944
R9561 gnd.n5892 gnd.n1572 19.3944
R9562 gnd.n5888 gnd.n1572 19.3944
R9563 gnd.n5888 gnd.n5887 19.3944
R9564 gnd.n5887 gnd.n5886 19.3944
R9565 gnd.n5886 gnd.n1577 19.3944
R9566 gnd.n5882 gnd.n1577 19.3944
R9567 gnd.n5882 gnd.n5881 19.3944
R9568 gnd.n5881 gnd.n5880 19.3944
R9569 gnd.n5880 gnd.n1582 19.3944
R9570 gnd.n5876 gnd.n1582 19.3944
R9571 gnd.n5185 gnd.n5183 19.3944
R9572 gnd.n5185 gnd.n5181 19.3944
R9573 gnd.n5191 gnd.n5181 19.3944
R9574 gnd.n5191 gnd.n5179 19.3944
R9575 gnd.n5196 gnd.n5179 19.3944
R9576 gnd.n5196 gnd.n5177 19.3944
R9577 gnd.n5202 gnd.n5177 19.3944
R9578 gnd.n5202 gnd.n5176 19.3944
R9579 gnd.n5211 gnd.n5176 19.3944
R9580 gnd.n5211 gnd.n5174 19.3944
R9581 gnd.n5217 gnd.n5174 19.3944
R9582 gnd.n5217 gnd.n5167 19.3944
R9583 gnd.n5230 gnd.n5167 19.3944
R9584 gnd.n5230 gnd.n5165 19.3944
R9585 gnd.n5236 gnd.n5165 19.3944
R9586 gnd.n5236 gnd.n5158 19.3944
R9587 gnd.n5249 gnd.n5158 19.3944
R9588 gnd.n5249 gnd.n5156 19.3944
R9589 gnd.n5255 gnd.n5156 19.3944
R9590 gnd.n5255 gnd.n5149 19.3944
R9591 gnd.n5268 gnd.n5149 19.3944
R9592 gnd.n5268 gnd.n5147 19.3944
R9593 gnd.n5275 gnd.n5147 19.3944
R9594 gnd.n5275 gnd.n5274 19.3944
R9595 gnd.n5288 gnd.n5128 19.3944
R9596 gnd.n5128 gnd.n5127 19.3944
R9597 gnd.n5295 gnd.n5127 19.3944
R9598 gnd.n5996 gnd.n5995 19.2005
R9599 gnd.n5412 gnd.n5411 19.2005
R9600 gnd.n3298 gnd.t167 18.8012
R9601 gnd.n3283 gnd.t310 18.8012
R9602 gnd.n3142 gnd.n3141 18.4825
R9603 gnd.n5577 gnd.n5485 18.4247
R9604 gnd.n6067 gnd.n6066 18.4247
R9605 gnd.n5285 gnd.n5284 18.2308
R9606 gnd.n6121 gnd.n6120 18.2308
R9607 gnd.n7246 gnd.n7189 18.2308
R9608 gnd.n4056 gnd.n4033 18.2308
R9609 gnd.t166 gnd.n2822 18.1639
R9610 gnd.n2850 gnd.t174 17.5266
R9611 gnd.n3249 gnd.t12 16.8893
R9612 gnd.n4220 gnd.t18 16.8893
R9613 gnd.n6192 gnd.t46 16.8893
R9614 gnd.n5121 gnd.t26 16.8893
R9615 gnd.n167 gnd.t22 16.8893
R9616 gnd.n5607 gnd.n1778 16.6793
R9617 gnd.n328 gnd.n198 16.6793
R9618 gnd.n4142 gnd.n4139 16.6793
R9619 gnd.n1398 gnd.n1395 16.6793
R9620 gnd.n3077 gnd.t125 16.2519
R9621 gnd.n2777 gnd.t293 16.2519
R9622 gnd.n6181 gnd.n1154 15.9333
R9623 gnd.n6181 gnd.n1168 15.9333
R9624 gnd.n4437 gnd.n4436 15.9333
R9625 gnd.n4436 gnd.n2313 15.9333
R9626 gnd.n4448 gnd.n2313 15.9333
R9627 gnd.n4448 gnd.n4447 15.9333
R9628 gnd.n2319 gnd.n2305 15.9333
R9629 gnd.n4457 gnd.n2305 15.9333
R9630 gnd.n4457 gnd.n2306 15.9333
R9631 gnd.n2306 gnd.n2298 15.9333
R9632 gnd.n4469 gnd.n2298 15.9333
R9633 gnd.n4469 gnd.n4468 15.9333
R9634 gnd.n4468 gnd.n2290 15.9333
R9635 gnd.n4481 gnd.n2290 15.9333
R9636 gnd.n4480 gnd.n1421 15.9333
R9637 gnd.n4493 gnd.n1453 15.9333
R9638 gnd.n5991 gnd.n1481 15.9333
R9639 gnd.n4516 gnd.n2177 15.9333
R9640 gnd.n4559 gnd.n2166 15.9333
R9641 gnd.n4593 gnd.n2154 15.9333
R9642 gnd.n4605 gnd.n4603 15.9333
R9643 gnd.n4632 gnd.n2134 15.9333
R9644 gnd.n4723 gnd.n2084 15.9333
R9645 gnd.n4742 gnd.n2061 15.9333
R9646 gnd.n2068 gnd.n2056 15.9333
R9647 gnd.n4782 gnd.n2039 15.9333
R9648 gnd.n4830 gnd.n4829 15.9333
R9649 gnd.n4838 gnd.n2026 15.9333
R9650 gnd.n4855 gnd.n4854 15.9333
R9651 gnd.n4915 gnd.n1993 15.9333
R9652 gnd.n4995 gnd.n4994 15.9333
R9653 gnd.n5003 gnd.n1936 15.9333
R9654 gnd.n5021 gnd.n5020 15.9333
R9655 gnd.n5031 gnd.n1908 15.9333
R9656 gnd.n5053 gnd.n1902 15.9333
R9657 gnd.n5323 gnd.n5322 15.9333
R9658 gnd.n5106 gnd.n1828 15.9333
R9659 gnd.n5106 gnd.n1791 15.9333
R9660 gnd.n5315 gnd.n1845 15.9333
R9661 gnd.n5314 gnd.n5313 15.9333
R9662 gnd.n5313 gnd.n5312 15.9333
R9663 gnd.n5312 gnd.n5310 15.9333
R9664 gnd.n5310 gnd.n1848 15.9333
R9665 gnd.n1860 gnd.n1848 15.9333
R9666 gnd.n1861 gnd.n1860 15.9333
R9667 gnd.n5304 gnd.n1861 15.9333
R9668 gnd.n5304 gnd.n5303 15.9333
R9669 gnd.n5302 gnd.n5301 15.9333
R9670 gnd.n5301 gnd.n1586 15.9333
R9671 gnd.n5874 gnd.n1586 15.9333
R9672 gnd.n5874 gnd.n5873 15.9333
R9673 gnd.n1597 gnd.n1588 15.9333
R9674 gnd.n5867 gnd.n1597 15.9333
R9675 gnd.n3764 gnd.n3762 15.6674
R9676 gnd.n3732 gnd.n3730 15.6674
R9677 gnd.n3700 gnd.n3698 15.6674
R9678 gnd.n3669 gnd.n3667 15.6674
R9679 gnd.n3637 gnd.n3635 15.6674
R9680 gnd.n3605 gnd.n3603 15.6674
R9681 gnd.n3573 gnd.n3571 15.6674
R9682 gnd.n3542 gnd.n3540 15.6674
R9683 gnd.n3068 gnd.t125 15.6146
R9684 gnd.t118 gnd.n2531 15.6146
R9685 gnd.t93 gnd.n2532 15.6146
R9686 gnd.t73 gnd.n2319 15.6146
R9687 gnd.n5303 gnd.t50 15.6146
R9688 gnd.n5659 gnd.n1757 15.3217
R9689 gnd.n383 gnd.n176 15.3217
R9690 gnd.n4099 gnd.n4011 15.3217
R9691 gnd.n1353 gnd.n1348 15.3217
R9692 gnd.n4633 gnd.n2139 15.296
R9693 gnd.n4652 gnd.n2130 15.296
R9694 gnd.n4613 gnd.t262 15.296
R9695 gnd.n4783 gnd.n4781 15.296
R9696 gnd.n4828 gnd.n2035 15.296
R9697 gnd.n4955 gnd.t5 15.296
R9698 gnd.n4895 gnd.n1958 15.296
R9699 gnd.n4993 gnd.n1945 15.296
R9700 gnd.n1886 gnd.t33 15.296
R9701 gnd.n5332 gnd.n5331 15.0827
R9702 gnd.n1465 gnd.n1460 15.0481
R9703 gnd.n5342 gnd.n5341 15.0481
R9704 gnd.n3436 gnd.t173 14.9773
R9705 gnd.t18 gnd.n2431 14.9773
R9706 gnd.n6062 gnd.n1421 14.9773
R9707 gnd.n7289 gnd.t22 14.9773
R9708 gnd.n4493 gnd.t109 14.6587
R9709 gnd.n4560 gnd.n2161 14.6587
R9710 gnd.n4695 gnd.n4694 14.6587
R9711 gnd.n1986 gnd.n1975 14.6587
R9712 gnd.n5033 gnd.n5032 14.6587
R9713 gnd.t30 gnd.n1882 14.6587
R9714 gnd.n5080 gnd.n5079 14.6587
R9715 gnd.t143 gnd.n2574 14.34
R9716 gnd.n3514 gnd.t165 14.34
R9717 gnd.n4518 gnd.t64 14.0214
R9718 gnd.n4568 gnd.n2146 14.0214
R9719 gnd.n4612 gnd.n2115 14.0214
R9720 gnd.n4773 gnd.n4772 14.0214
R9721 gnd.n2025 gnd.n2017 14.0214
R9722 gnd.n4956 gnd.n1962 14.0214
R9723 gnd.n1934 gnd.n1933 14.0214
R9724 gnd.n5324 gnd.n1833 14.0214
R9725 gnd.n3224 gnd.t220 13.7027
R9726 gnd.n2088 gnd.t199 13.7027
R9727 gnd.n4863 gnd.t319 13.7027
R9728 gnd.n2934 gnd.n2933 13.5763
R9729 gnd.n3878 gnd.n2488 13.5763
R9730 gnd.n3142 gnd.n2880 13.384
R9731 gnd.n4503 gnd.n1490 13.384
R9732 gnd.n4592 gnd.n2156 13.384
R9733 gnd.n2116 gnd.n2110 13.384
R9734 gnd.t248 gnd.n4682 13.384
R9735 gnd.n4934 gnd.t1 13.384
R9736 gnd.n4943 gnd.n1971 13.384
R9737 gnd.n4971 gnd.n1922 13.384
R9738 gnd.n5096 gnd.n1873 13.384
R9739 gnd.n1476 gnd.n1457 13.1884
R9740 gnd.n1471 gnd.n1470 13.1884
R9741 gnd.n1470 gnd.n1469 13.1884
R9742 gnd.n5335 gnd.n5330 13.1884
R9743 gnd.n5336 gnd.n5335 13.1884
R9744 gnd.n1472 gnd.n1459 13.146
R9745 gnd.n1468 gnd.n1459 13.146
R9746 gnd.n5334 gnd.n5333 13.146
R9747 gnd.n5334 gnd.n5329 13.146
R9748 gnd.n4534 gnd.t275 13.0654
R9749 gnd.n5054 gnd.t229 13.0654
R9750 gnd.n3765 gnd.n3761 12.8005
R9751 gnd.n3733 gnd.n3729 12.8005
R9752 gnd.n3701 gnd.n3697 12.8005
R9753 gnd.n3670 gnd.n3666 12.8005
R9754 gnd.n3638 gnd.n3634 12.8005
R9755 gnd.n3606 gnd.n3602 12.8005
R9756 gnd.n3574 gnd.n3570 12.8005
R9757 gnd.n3543 gnd.n3539 12.8005
R9758 gnd.n2192 gnd.n1492 12.7467
R9759 gnd.n4551 gnd.t84 12.7467
R9760 gnd.n4576 gnd.n4575 12.7467
R9761 gnd.n4743 gnd.n4741 12.7467
R9762 gnd.n4853 gnd.n2004 12.7467
R9763 gnd.n5019 gnd.n5018 12.7467
R9764 gnd.n2434 gnd.n2423 12.4281
R9765 gnd.n7295 gnd.n149 12.4281
R9766 gnd.n2933 gnd.n2928 12.4126
R9767 gnd.n3881 gnd.n3878 12.4126
R9768 gnd.n6059 gnd.n5996 12.1761
R9769 gnd.n5411 gnd.n5410 12.1761
R9770 gnd.n5992 gnd.n1479 12.1094
R9771 gnd.t40 gnd.n2196 12.1094
R9772 gnd.n4583 gnd.n2147 12.1094
R9773 gnd.n4664 gnd.n2121 12.1094
R9774 gnd.n4963 gnd.n1956 12.1094
R9775 gnd.n5004 gnd.n1931 12.1094
R9776 gnd.n5104 gnd.n1836 12.1094
R9777 gnd.n3769 gnd.n3768 12.0247
R9778 gnd.n3737 gnd.n3736 12.0247
R9779 gnd.n3705 gnd.n3704 12.0247
R9780 gnd.n3674 gnd.n3673 12.0247
R9781 gnd.n3642 gnd.n3641 12.0247
R9782 gnd.n3610 gnd.n3609 12.0247
R9783 gnd.n3578 gnd.n3577 12.0247
R9784 gnd.n3547 gnd.n3546 12.0247
R9785 gnd.n6217 gnd.t136 11.7908
R9786 gnd.n5840 gnd.t151 11.7908
R9787 gnd.n6116 gnd.n1257 11.4721
R9788 gnd.n4544 gnd.n2178 11.4721
R9789 gnd.n4536 gnd.n4535 11.4721
R9790 gnd.n4703 gnd.t213 11.4721
R9791 gnd.n4702 gnd.n2097 11.4721
R9792 gnd.n4733 gnd.n4732 11.4721
R9793 gnd.n4880 gnd.n1999 11.4721
R9794 gnd.n4872 gnd.n1985 11.4721
R9795 gnd.n4924 gnd.t2 11.4721
R9796 gnd.n5044 gnd.n1909 11.4721
R9797 gnd.n5065 gnd.n5064 11.4721
R9798 gnd.n5865 gnd.n1598 11.4721
R9799 gnd.n3772 gnd.n3759 11.249
R9800 gnd.n3740 gnd.n3727 11.249
R9801 gnd.n3708 gnd.n3695 11.249
R9802 gnd.n3677 gnd.n3664 11.249
R9803 gnd.n3645 gnd.n3632 11.249
R9804 gnd.n3613 gnd.n3600 11.249
R9805 gnd.n3581 gnd.n3568 11.249
R9806 gnd.n3550 gnd.n3537 11.249
R9807 gnd.n3212 gnd.t220 11.1535
R9808 gnd.t266 gnd.n994 11.1535
R9809 gnd.n6241 gnd.t203 11.1535
R9810 gnd.n4481 gnd.t246 11.1535
R9811 gnd.n4680 gnd.t147 11.1535
R9812 gnd.t145 gnd.n4935 11.1535
R9813 gnd.t312 gnd.n5314 11.1535
R9814 gnd.n5816 gnd.t179 11.1535
R9815 gnd.n391 gnd.t162 11.1535
R9816 gnd.n6306 gnd.n967 10.8348
R9817 gnd.n6305 gnd.n970 10.8348
R9818 gnd.n4252 gnd.n980 10.8348
R9819 gnd.n4260 gnd.n991 10.8348
R9820 gnd.n6293 gnd.n994 10.8348
R9821 gnd.n4267 gnd.n1002 10.8348
R9822 gnd.n6287 gnd.n1005 10.8348
R9823 gnd.n4279 gnd.n4278 10.8348
R9824 gnd.n6281 gnd.n1014 10.8348
R9825 gnd.n4333 gnd.n2370 10.8348
R9826 gnd.n6273 gnd.n1025 10.8348
R9827 gnd.n4326 gnd.n4325 10.8348
R9828 gnd.n6267 gnd.n1036 10.8348
R9829 gnd.n4296 gnd.n1041 10.8348
R9830 gnd.n4315 gnd.n1050 10.8348
R9831 gnd.n6254 gnd.n1053 10.8348
R9832 gnd.n4307 gnd.n1058 10.8348
R9833 gnd.n6247 gnd.n1061 10.8348
R9834 gnd.n4363 gnd.n4362 10.8348
R9835 gnd.n6241 gnd.n1070 10.8348
R9836 gnd.n4371 gnd.n1078 10.8348
R9837 gnd.n4377 gnd.n1087 10.8348
R9838 gnd.n6229 gnd.n1090 10.8348
R9839 gnd.n4385 gnd.n1098 10.8348
R9840 gnd.n6223 gnd.n1101 10.8348
R9841 gnd.n4410 gnd.n4409 10.8348
R9842 gnd.n6217 gnd.n1110 10.8348
R9843 gnd.n4392 gnd.n1118 10.8348
R9844 gnd.n6211 gnd.n1121 10.8348
R9845 gnd.n4398 gnd.n1128 10.8348
R9846 gnd.n6205 gnd.n1131 10.8348
R9847 gnd.n6192 gnd.n1138 10.8348
R9848 gnd.n6199 gnd.n1141 10.8348
R9849 gnd.n4646 gnd.n4645 10.8348
R9850 gnd.n4645 gnd.n4644 10.8348
R9851 gnd.n4822 gnd.n4821 10.8348
R9852 gnd.n4821 gnd.n2032 10.8348
R9853 gnd.n4987 gnd.n4986 10.8348
R9854 gnd.n4986 gnd.n1942 10.8348
R9855 gnd.n5859 gnd.n5858 10.8348
R9856 gnd.n5121 gnd.n1609 10.8348
R9857 gnd.n5852 gnd.n1618 10.8348
R9858 gnd.n5669 gnd.n1621 10.8348
R9859 gnd.n5846 gnd.n1630 10.8348
R9860 gnd.n5677 gnd.n1633 10.8348
R9861 gnd.n5840 gnd.n1641 10.8348
R9862 gnd.n5698 gnd.n5697 10.8348
R9863 gnd.n5834 gnd.n1650 10.8348
R9864 gnd.n5686 gnd.n1653 10.8348
R9865 gnd.n5828 gnd.n1661 10.8348
R9866 gnd.n5742 gnd.n1664 10.8348
R9867 gnd.n5749 gnd.n1673 10.8348
R9868 gnd.n5816 gnd.n1681 10.8348
R9869 gnd.n5767 gnd.n1729 10.8348
R9870 gnd.n5810 gnd.n1690 10.8348
R9871 gnd.n5806 gnd.n1693 10.8348
R9872 gnd.n5805 gnd.n1699 10.8348
R9873 gnd.n1706 gnd.n1705 10.8348
R9874 gnd.n5792 gnd.n1709 10.8348
R9875 gnd.n5785 gnd.n1722 10.8348
R9876 gnd.n7339 gnd.n69 10.8348
R9877 gnd.n7137 gnd.n71 10.8348
R9878 gnd.n7331 gnd.n86 10.8348
R9879 gnd.n7152 gnd.n89 10.8348
R9880 gnd.n7325 gnd.n98 10.8348
R9881 gnd.n7159 gnd.n101 10.8348
R9882 gnd.n7319 gnd.n108 10.8348
R9883 gnd.n7167 gnd.n391 10.8348
R9884 gnd.n7313 gnd.n117 10.8348
R9885 gnd.n7307 gnd.n128 10.8348
R9886 gnd.n7266 gnd.n131 10.8348
R9887 gnd.n7301 gnd.n138 10.8348
R9888 gnd.n1758 gnd.n1757 10.6672
R9889 gnd.n378 gnd.n176 10.6672
R9890 gnd.n4102 gnd.n4099 10.6672
R9891 gnd.n1356 gnd.n1353 10.6672
R9892 gnd.n5476 gnd.n1787 10.6151
R9893 gnd.n5476 gnd.n5475 10.6151
R9894 gnd.n5473 gnd.n5470 10.6151
R9895 gnd.n5470 gnd.n5469 10.6151
R9896 gnd.n5469 gnd.n5466 10.6151
R9897 gnd.n5466 gnd.n5465 10.6151
R9898 gnd.n5465 gnd.n5462 10.6151
R9899 gnd.n5462 gnd.n5461 10.6151
R9900 gnd.n5461 gnd.n5458 10.6151
R9901 gnd.n5458 gnd.n5457 10.6151
R9902 gnd.n5457 gnd.n5454 10.6151
R9903 gnd.n5454 gnd.n5453 10.6151
R9904 gnd.n5453 gnd.n5450 10.6151
R9905 gnd.n5450 gnd.n5449 10.6151
R9906 gnd.n5449 gnd.n5446 10.6151
R9907 gnd.n5446 gnd.n5445 10.6151
R9908 gnd.n5445 gnd.n5442 10.6151
R9909 gnd.n5442 gnd.n5441 10.6151
R9910 gnd.n5441 gnd.n5438 10.6151
R9911 gnd.n5438 gnd.n5437 10.6151
R9912 gnd.n5437 gnd.n5434 10.6151
R9913 gnd.n5434 gnd.n5433 10.6151
R9914 gnd.n5433 gnd.n5430 10.6151
R9915 gnd.n5430 gnd.n5429 10.6151
R9916 gnd.n5429 gnd.n5426 10.6151
R9917 gnd.n5426 gnd.n5425 10.6151
R9918 gnd.n5425 gnd.n5422 10.6151
R9919 gnd.n5422 gnd.n5421 10.6151
R9920 gnd.n5421 gnd.n5418 10.6151
R9921 gnd.n5418 gnd.n5417 10.6151
R9922 gnd.n2279 gnd.n2278 10.6151
R9923 gnd.n2278 gnd.n2277 10.6151
R9924 gnd.n2277 gnd.n2274 10.6151
R9925 gnd.n2274 gnd.n2273 10.6151
R9926 gnd.n2273 gnd.n2270 10.6151
R9927 gnd.n2270 gnd.n2269 10.6151
R9928 gnd.n2269 gnd.n2175 10.6151
R9929 gnd.n4546 gnd.n2175 10.6151
R9930 gnd.n4547 gnd.n4546 10.6151
R9931 gnd.n4549 gnd.n4547 10.6151
R9932 gnd.n4549 gnd.n4548 10.6151
R9933 gnd.n4548 gnd.n2163 10.6151
R9934 gnd.n4562 gnd.n2163 10.6151
R9935 gnd.n4563 gnd.n4562 10.6151
R9936 gnd.n4573 gnd.n4563 10.6151
R9937 gnd.n4573 gnd.n4572 10.6151
R9938 gnd.n4572 gnd.n4571 10.6151
R9939 gnd.n4571 gnd.n4564 10.6151
R9940 gnd.n4565 gnd.n4564 10.6151
R9941 gnd.n4565 gnd.n2137 10.6151
R9942 gnd.n4635 gnd.n2137 10.6151
R9943 gnd.n4636 gnd.n4635 10.6151
R9944 gnd.n4642 gnd.n4636 10.6151
R9945 gnd.n4642 gnd.n4641 10.6151
R9946 gnd.n4641 gnd.n4640 10.6151
R9947 gnd.n4640 gnd.n4637 10.6151
R9948 gnd.n4637 gnd.n2113 10.6151
R9949 gnd.n4673 gnd.n2113 10.6151
R9950 gnd.n4674 gnd.n4673 10.6151
R9951 gnd.n4678 gnd.n4674 10.6151
R9952 gnd.n4678 gnd.n4677 10.6151
R9953 gnd.n4677 gnd.n4676 10.6151
R9954 gnd.n4676 gnd.n4675 10.6151
R9955 gnd.n4675 gnd.n2087 10.6151
R9956 gnd.n4721 gnd.n2087 10.6151
R9957 gnd.n4721 gnd.n4720 10.6151
R9958 gnd.n4720 gnd.n4719 10.6151
R9959 gnd.n4719 gnd.n4718 10.6151
R9960 gnd.n4718 gnd.n2069 10.6151
R9961 gnd.n4745 gnd.n2069 10.6151
R9962 gnd.n4746 gnd.n4745 10.6151
R9963 gnd.n4748 gnd.n4746 10.6151
R9964 gnd.n4749 gnd.n4748 10.6151
R9965 gnd.n4750 gnd.n4749 10.6151
R9966 gnd.n4750 gnd.n2046 10.6151
R9967 gnd.n4785 gnd.n2046 10.6151
R9968 gnd.n4786 gnd.n4785 10.6151
R9969 gnd.n4788 gnd.n4786 10.6151
R9970 gnd.n4789 gnd.n4788 10.6151
R9971 gnd.n4791 gnd.n4789 10.6151
R9972 gnd.n4791 gnd.n4790 10.6151
R9973 gnd.n4790 gnd.n2015 10.6151
R9974 gnd.n4848 gnd.n2015 10.6151
R9975 gnd.n4849 gnd.n4848 10.6151
R9976 gnd.n4851 gnd.n4849 10.6151
R9977 gnd.n4851 gnd.n4850 10.6151
R9978 gnd.n4850 gnd.n1996 10.6151
R9979 gnd.n4882 gnd.n1996 10.6151
R9980 gnd.n4883 gnd.n4882 10.6151
R9981 gnd.n4913 gnd.n4883 10.6151
R9982 gnd.n4913 gnd.n4912 10.6151
R9983 gnd.n4912 gnd.n4911 10.6151
R9984 gnd.n4911 gnd.n4908 10.6151
R9985 gnd.n4908 gnd.n4907 10.6151
R9986 gnd.n4907 gnd.n4906 10.6151
R9987 gnd.n4906 gnd.n4905 10.6151
R9988 gnd.n4905 gnd.n4904 10.6151
R9989 gnd.n4904 gnd.n4901 10.6151
R9990 gnd.n4901 gnd.n4900 10.6151
R9991 gnd.n4900 gnd.n4898 10.6151
R9992 gnd.n4898 gnd.n4897 10.6151
R9993 gnd.n4897 gnd.n4891 10.6151
R9994 gnd.n4891 gnd.n4890 10.6151
R9995 gnd.n4890 gnd.n4888 10.6151
R9996 gnd.n4888 gnd.n4887 10.6151
R9997 gnd.n4887 gnd.n4884 10.6151
R9998 gnd.n4884 gnd.n1925 10.6151
R9999 gnd.n5013 gnd.n1925 10.6151
R10000 gnd.n5014 gnd.n5013 10.6151
R10001 gnd.n5016 gnd.n5014 10.6151
R10002 gnd.n5016 gnd.n5015 10.6151
R10003 gnd.n5015 gnd.n1905 10.6151
R10004 gnd.n5046 gnd.n1905 10.6151
R10005 gnd.n5047 gnd.n5046 10.6151
R10006 gnd.n5051 gnd.n5047 10.6151
R10007 gnd.n5051 gnd.n5050 10.6151
R10008 gnd.n5050 gnd.n5049 10.6151
R10009 gnd.n5049 gnd.n5048 10.6151
R10010 gnd.n5048 gnd.n1875 10.6151
R10011 gnd.n5089 gnd.n1875 10.6151
R10012 gnd.n5090 gnd.n5089 10.6151
R10013 gnd.n5093 gnd.n5090 10.6151
R10014 gnd.n5093 gnd.n5092 10.6151
R10015 gnd.n5092 gnd.n5091 10.6151
R10016 gnd.n5091 gnd.n1826 10.6151
R10017 gnd.n2207 gnd.n1417 10.6151
R10018 gnd.n2210 gnd.n2207 10.6151
R10019 gnd.n2215 gnd.n2212 10.6151
R10020 gnd.n2216 gnd.n2215 10.6151
R10021 gnd.n2219 gnd.n2216 10.6151
R10022 gnd.n2220 gnd.n2219 10.6151
R10023 gnd.n2223 gnd.n2220 10.6151
R10024 gnd.n2224 gnd.n2223 10.6151
R10025 gnd.n2227 gnd.n2224 10.6151
R10026 gnd.n2228 gnd.n2227 10.6151
R10027 gnd.n2231 gnd.n2228 10.6151
R10028 gnd.n2232 gnd.n2231 10.6151
R10029 gnd.n2235 gnd.n2232 10.6151
R10030 gnd.n2236 gnd.n2235 10.6151
R10031 gnd.n2239 gnd.n2236 10.6151
R10032 gnd.n2240 gnd.n2239 10.6151
R10033 gnd.n2243 gnd.n2240 10.6151
R10034 gnd.n2244 gnd.n2243 10.6151
R10035 gnd.n2247 gnd.n2244 10.6151
R10036 gnd.n2248 gnd.n2247 10.6151
R10037 gnd.n2251 gnd.n2248 10.6151
R10038 gnd.n2252 gnd.n2251 10.6151
R10039 gnd.n2255 gnd.n2252 10.6151
R10040 gnd.n2256 gnd.n2255 10.6151
R10041 gnd.n2259 gnd.n2256 10.6151
R10042 gnd.n2260 gnd.n2259 10.6151
R10043 gnd.n2263 gnd.n2260 10.6151
R10044 gnd.n2264 gnd.n2263 10.6151
R10045 gnd.n2267 gnd.n2264 10.6151
R10046 gnd.n2268 gnd.n2267 10.6151
R10047 gnd.n6059 gnd.n6058 10.6151
R10048 gnd.n6058 gnd.n6057 10.6151
R10049 gnd.n6057 gnd.n6056 10.6151
R10050 gnd.n6056 gnd.n6054 10.6151
R10051 gnd.n6054 gnd.n6051 10.6151
R10052 gnd.n6051 gnd.n6050 10.6151
R10053 gnd.n6050 gnd.n6047 10.6151
R10054 gnd.n6047 gnd.n6046 10.6151
R10055 gnd.n6046 gnd.n6043 10.6151
R10056 gnd.n6043 gnd.n6042 10.6151
R10057 gnd.n6042 gnd.n6039 10.6151
R10058 gnd.n6039 gnd.n6038 10.6151
R10059 gnd.n6038 gnd.n6035 10.6151
R10060 gnd.n6035 gnd.n6034 10.6151
R10061 gnd.n6034 gnd.n6031 10.6151
R10062 gnd.n6031 gnd.n6030 10.6151
R10063 gnd.n6030 gnd.n6027 10.6151
R10064 gnd.n6027 gnd.n6026 10.6151
R10065 gnd.n6026 gnd.n6023 10.6151
R10066 gnd.n6023 gnd.n6022 10.6151
R10067 gnd.n6022 gnd.n6019 10.6151
R10068 gnd.n6019 gnd.n6018 10.6151
R10069 gnd.n6018 gnd.n6015 10.6151
R10070 gnd.n6015 gnd.n6014 10.6151
R10071 gnd.n6014 gnd.n6011 10.6151
R10072 gnd.n6011 gnd.n6010 10.6151
R10073 gnd.n6010 gnd.n6007 10.6151
R10074 gnd.n6007 gnd.n6006 10.6151
R10075 gnd.n6003 gnd.n6002 10.6151
R10076 gnd.n6002 gnd.n1418 10.6151
R10077 gnd.n5410 gnd.n5409 10.6151
R10078 gnd.n5409 gnd.n5406 10.6151
R10079 gnd.n5406 gnd.n5405 10.6151
R10080 gnd.n5405 gnd.n5402 10.6151
R10081 gnd.n5402 gnd.n5401 10.6151
R10082 gnd.n5401 gnd.n5398 10.6151
R10083 gnd.n5398 gnd.n5397 10.6151
R10084 gnd.n5397 gnd.n5394 10.6151
R10085 gnd.n5394 gnd.n5393 10.6151
R10086 gnd.n5393 gnd.n5390 10.6151
R10087 gnd.n5390 gnd.n5389 10.6151
R10088 gnd.n5389 gnd.n5386 10.6151
R10089 gnd.n5386 gnd.n5385 10.6151
R10090 gnd.n5385 gnd.n5382 10.6151
R10091 gnd.n5382 gnd.n5381 10.6151
R10092 gnd.n5381 gnd.n5378 10.6151
R10093 gnd.n5378 gnd.n5377 10.6151
R10094 gnd.n5377 gnd.n5374 10.6151
R10095 gnd.n5374 gnd.n5373 10.6151
R10096 gnd.n5373 gnd.n5370 10.6151
R10097 gnd.n5370 gnd.n5369 10.6151
R10098 gnd.n5369 gnd.n5366 10.6151
R10099 gnd.n5366 gnd.n5365 10.6151
R10100 gnd.n5365 gnd.n5362 10.6151
R10101 gnd.n5362 gnd.n5361 10.6151
R10102 gnd.n5361 gnd.n5358 10.6151
R10103 gnd.n5358 gnd.n5357 10.6151
R10104 gnd.n5357 gnd.n5354 10.6151
R10105 gnd.n5352 gnd.n5349 10.6151
R10106 gnd.n5349 gnd.n1788 10.6151
R10107 gnd.n5995 gnd.n5994 10.6151
R10108 gnd.n5994 gnd.n1477 10.6151
R10109 gnd.n2195 gnd.n1477 10.6151
R10110 gnd.n4507 gnd.n2195 10.6151
R10111 gnd.n4508 gnd.n4507 10.6151
R10112 gnd.n4509 gnd.n4508 10.6151
R10113 gnd.n4509 gnd.n2181 10.6151
R10114 gnd.n4542 gnd.n2181 10.6151
R10115 gnd.n4542 gnd.n4541 10.6151
R10116 gnd.n4541 gnd.n4540 10.6151
R10117 gnd.n4540 gnd.n4539 10.6151
R10118 gnd.n4539 gnd.n2182 10.6151
R10119 gnd.n2182 gnd.n2159 10.6151
R10120 gnd.n4579 gnd.n2159 10.6151
R10121 gnd.n4580 gnd.n4579 10.6151
R10122 gnd.n4590 gnd.n4580 10.6151
R10123 gnd.n4590 gnd.n4589 10.6151
R10124 gnd.n4589 gnd.n4588 10.6151
R10125 gnd.n4588 gnd.n4581 10.6151
R10126 gnd.n4582 gnd.n4581 10.6151
R10127 gnd.n4582 gnd.n2132 10.6151
R10128 gnd.n4648 gnd.n2132 10.6151
R10129 gnd.n4649 gnd.n4648 10.6151
R10130 gnd.n4650 gnd.n4649 10.6151
R10131 gnd.n4650 gnd.n2119 10.6151
R10132 gnd.n4666 gnd.n2119 10.6151
R10133 gnd.n4667 gnd.n4666 10.6151
R10134 gnd.n4669 gnd.n4667 10.6151
R10135 gnd.n4669 gnd.n4668 10.6151
R10136 gnd.n4668 gnd.n2099 10.6151
R10137 gnd.n4698 gnd.n2099 10.6151
R10138 gnd.n4699 gnd.n4698 10.6151
R10139 gnd.n4700 gnd.n4699 10.6151
R10140 gnd.n4700 gnd.n2082 10.6151
R10141 gnd.n4725 gnd.n2082 10.6151
R10142 gnd.n4726 gnd.n4725 10.6151
R10143 gnd.n4730 gnd.n4726 10.6151
R10144 gnd.n4730 gnd.n4729 10.6151
R10145 gnd.n4729 gnd.n4728 10.6151
R10146 gnd.n4728 gnd.n2059 10.6151
R10147 gnd.n4765 gnd.n2059 10.6151
R10148 gnd.n4766 gnd.n4765 10.6151
R10149 gnd.n4770 gnd.n4766 10.6151
R10150 gnd.n4770 gnd.n4769 10.6151
R10151 gnd.n4769 gnd.n4768 10.6151
R10152 gnd.n4768 gnd.n2037 10.6151
R10153 gnd.n4824 gnd.n2037 10.6151
R10154 gnd.n4825 gnd.n4824 10.6151
R10155 gnd.n4826 gnd.n4825 10.6151
R10156 gnd.n4826 gnd.n2022 10.6151
R10157 gnd.n4841 gnd.n2022 10.6151
R10158 gnd.n4842 gnd.n4841 10.6151
R10159 gnd.n4844 gnd.n4842 10.6151
R10160 gnd.n4844 gnd.n4843 10.6151
R10161 gnd.n4843 gnd.n2002 10.6151
R10162 gnd.n4868 gnd.n2002 10.6151
R10163 gnd.n4869 gnd.n4868 10.6151
R10164 gnd.n4878 gnd.n4869 10.6151
R10165 gnd.n4878 gnd.n4877 10.6151
R10166 gnd.n4877 gnd.n4876 10.6151
R10167 gnd.n4876 gnd.n4875 10.6151
R10168 gnd.n4875 gnd.n4870 10.6151
R10169 gnd.n4870 gnd.n1973 10.6151
R10170 gnd.n4939 gnd.n1973 10.6151
R10171 gnd.n4940 gnd.n4939 10.6151
R10172 gnd.n4941 gnd.n4940 10.6151
R10173 gnd.n4941 gnd.n1960 10.6151
R10174 gnd.n4958 gnd.n1960 10.6151
R10175 gnd.n4959 gnd.n4958 10.6151
R10176 gnd.n4960 gnd.n4959 10.6151
R10177 gnd.n4960 gnd.n1947 10.6151
R10178 gnd.n4989 gnd.n1947 10.6151
R10179 gnd.n4990 gnd.n4989 10.6151
R10180 gnd.n4991 gnd.n4990 10.6151
R10181 gnd.n4991 gnd.n1929 10.6151
R10182 gnd.n5006 gnd.n1929 10.6151
R10183 gnd.n5007 gnd.n5006 10.6151
R10184 gnd.n5009 gnd.n5007 10.6151
R10185 gnd.n5009 gnd.n5008 10.6151
R10186 gnd.n5008 gnd.n1912 10.6151
R10187 gnd.n5036 gnd.n1912 10.6151
R10188 gnd.n5037 gnd.n5036 10.6151
R10189 gnd.n5042 gnd.n5037 10.6151
R10190 gnd.n5042 gnd.n5041 10.6151
R10191 gnd.n5041 gnd.n5040 10.6151
R10192 gnd.n5040 gnd.n5039 10.6151
R10193 gnd.n5039 gnd.n1880 10.6151
R10194 gnd.n5082 gnd.n1880 10.6151
R10195 gnd.n5083 gnd.n5082 10.6151
R10196 gnd.n5085 gnd.n5083 10.6151
R10197 gnd.n5085 gnd.n5084 10.6151
R10198 gnd.n5084 gnd.n1831 10.6151
R10199 gnd.n5326 gnd.n1831 10.6151
R10200 gnd.n5327 gnd.n5326 10.6151
R10201 gnd.n5412 gnd.n5327 10.6151
R10202 gnd.n3131 gnd.t289 10.5161
R10203 gnd.n2576 gnd.t143 10.5161
R10204 gnd.n3497 gnd.t165 10.5161
R10205 gnd.t157 gnd.n1022 10.5161
R10206 gnd.n4325 gnd.t155 10.5161
R10207 gnd.n6267 gnd.t155 10.5161
R10208 gnd.n6260 gnd.t197 10.5161
R10209 gnd.n4655 gnd.t211 10.5161
R10210 gnd.t299 gnd.n4892 10.5161
R10211 gnd.t149 gnd.n5797 10.5161
R10212 gnd.n5785 gnd.t8 10.5161
R10213 gnd.t8 gnd.n69 10.5161
R10214 gnd.n7136 gnd.t134 10.5161
R10215 gnd.n3773 gnd.n3757 10.4732
R10216 gnd.n3741 gnd.n3725 10.4732
R10217 gnd.n3709 gnd.n3693 10.4732
R10218 gnd.n3678 gnd.n3662 10.4732
R10219 gnd.n3646 gnd.n3630 10.4732
R10220 gnd.n3614 gnd.n3598 10.4732
R10221 gnd.n3582 gnd.n3566 10.4732
R10222 gnd.n3551 gnd.n3535 10.4732
R10223 gnd.n2184 gnd.n2178 10.1975
R10224 gnd.n2097 gnd.n2096 10.1975
R10225 gnd.n4733 gnd.n2077 10.1975
R10226 gnd.n4801 gnd.n1999 10.1975
R10227 gnd.n4873 gnd.n4872 10.1975
R10228 gnd.n5065 gnd.n1892 10.1975
R10229 gnd.n1845 gnd.t54 10.1975
R10230 gnd.n2415 gnd.t175 9.87883
R10231 gnd.n4267 gnd.t266 9.87883
R10232 gnd.n4362 gnd.t203 9.87883
R10233 gnd.n6235 gnd.t287 9.87883
R10234 gnd.n5822 gnd.t177 9.87883
R10235 gnd.n1729 gnd.t179 9.87883
R10236 gnd.n7319 gnd.t162 9.87883
R10237 gnd.t159 gnd.n120 9.87883
R10238 gnd.n3777 gnd.n3776 9.69747
R10239 gnd.n3745 gnd.n3744 9.69747
R10240 gnd.n3713 gnd.n3712 9.69747
R10241 gnd.n3682 gnd.n3681 9.69747
R10242 gnd.n3650 gnd.n3649 9.69747
R10243 gnd.n3618 gnd.n3617 9.69747
R10244 gnd.n3586 gnd.n3585 9.69747
R10245 gnd.n3555 gnd.n3554 9.69747
R10246 gnd.n2281 gnd.n1479 9.56018
R10247 gnd.n4584 gnd.n4583 9.56018
R10248 gnd.n4638 gnd.n2121 9.56018
R10249 gnd.n4707 gnd.t257 9.56018
R10250 gnd.n4753 gnd.n2048 9.56018
R10251 gnd.n4794 gnd.n4793 9.56018
R10252 gnd.n4803 gnd.t142 9.56018
R10253 gnd.n4963 gnd.n4962 9.56018
R10254 gnd.n4885 gnd.n1931 9.56018
R10255 gnd.n3783 gnd.n3782 9.45567
R10256 gnd.n3751 gnd.n3750 9.45567
R10257 gnd.n3719 gnd.n3718 9.45567
R10258 gnd.n3688 gnd.n3687 9.45567
R10259 gnd.n3656 gnd.n3655 9.45567
R10260 gnd.n3624 gnd.n3623 9.45567
R10261 gnd.n3592 gnd.n3591 9.45567
R10262 gnd.n3561 gnd.n3560 9.45567
R10263 gnd.n5607 gnd.n1776 9.30959
R10264 gnd.n334 gnd.n198 9.30959
R10265 gnd.n4139 gnd.n4138 9.30959
R10266 gnd.n1395 gnd.n1327 9.30959
R10267 gnd.n3782 gnd.n3781 9.3005
R10268 gnd.n3755 gnd.n3754 9.3005
R10269 gnd.n3776 gnd.n3775 9.3005
R10270 gnd.n3774 gnd.n3773 9.3005
R10271 gnd.n3759 gnd.n3758 9.3005
R10272 gnd.n3768 gnd.n3767 9.3005
R10273 gnd.n3766 gnd.n3765 9.3005
R10274 gnd.n3750 gnd.n3749 9.3005
R10275 gnd.n3723 gnd.n3722 9.3005
R10276 gnd.n3744 gnd.n3743 9.3005
R10277 gnd.n3742 gnd.n3741 9.3005
R10278 gnd.n3727 gnd.n3726 9.3005
R10279 gnd.n3736 gnd.n3735 9.3005
R10280 gnd.n3734 gnd.n3733 9.3005
R10281 gnd.n3718 gnd.n3717 9.3005
R10282 gnd.n3691 gnd.n3690 9.3005
R10283 gnd.n3712 gnd.n3711 9.3005
R10284 gnd.n3710 gnd.n3709 9.3005
R10285 gnd.n3695 gnd.n3694 9.3005
R10286 gnd.n3704 gnd.n3703 9.3005
R10287 gnd.n3702 gnd.n3701 9.3005
R10288 gnd.n3687 gnd.n3686 9.3005
R10289 gnd.n3660 gnd.n3659 9.3005
R10290 gnd.n3681 gnd.n3680 9.3005
R10291 gnd.n3679 gnd.n3678 9.3005
R10292 gnd.n3664 gnd.n3663 9.3005
R10293 gnd.n3673 gnd.n3672 9.3005
R10294 gnd.n3671 gnd.n3670 9.3005
R10295 gnd.n3655 gnd.n3654 9.3005
R10296 gnd.n3628 gnd.n3627 9.3005
R10297 gnd.n3649 gnd.n3648 9.3005
R10298 gnd.n3647 gnd.n3646 9.3005
R10299 gnd.n3632 gnd.n3631 9.3005
R10300 gnd.n3641 gnd.n3640 9.3005
R10301 gnd.n3639 gnd.n3638 9.3005
R10302 gnd.n3623 gnd.n3622 9.3005
R10303 gnd.n3596 gnd.n3595 9.3005
R10304 gnd.n3617 gnd.n3616 9.3005
R10305 gnd.n3615 gnd.n3614 9.3005
R10306 gnd.n3600 gnd.n3599 9.3005
R10307 gnd.n3609 gnd.n3608 9.3005
R10308 gnd.n3607 gnd.n3606 9.3005
R10309 gnd.n3591 gnd.n3590 9.3005
R10310 gnd.n3564 gnd.n3563 9.3005
R10311 gnd.n3585 gnd.n3584 9.3005
R10312 gnd.n3583 gnd.n3582 9.3005
R10313 gnd.n3568 gnd.n3567 9.3005
R10314 gnd.n3577 gnd.n3576 9.3005
R10315 gnd.n3575 gnd.n3574 9.3005
R10316 gnd.n3560 gnd.n3559 9.3005
R10317 gnd.n3533 gnd.n3532 9.3005
R10318 gnd.n3554 gnd.n3553 9.3005
R10319 gnd.n3552 gnd.n3551 9.3005
R10320 gnd.n3537 gnd.n3536 9.3005
R10321 gnd.n3546 gnd.n3545 9.3005
R10322 gnd.n3544 gnd.n3543 9.3005
R10323 gnd.n3908 gnd.n3907 9.3005
R10324 gnd.n3906 gnd.n2476 9.3005
R10325 gnd.n3905 gnd.n3904 9.3005
R10326 gnd.n3901 gnd.n2477 9.3005
R10327 gnd.n3898 gnd.n2478 9.3005
R10328 gnd.n3897 gnd.n2479 9.3005
R10329 gnd.n3894 gnd.n2480 9.3005
R10330 gnd.n3893 gnd.n2481 9.3005
R10331 gnd.n3890 gnd.n2482 9.3005
R10332 gnd.n3889 gnd.n2483 9.3005
R10333 gnd.n3886 gnd.n2484 9.3005
R10334 gnd.n3885 gnd.n2485 9.3005
R10335 gnd.n3882 gnd.n2486 9.3005
R10336 gnd.n3881 gnd.n2487 9.3005
R10337 gnd.n3878 gnd.n3877 9.3005
R10338 gnd.n3876 gnd.n2488 9.3005
R10339 gnd.n3909 gnd.n2475 9.3005
R10340 gnd.n3150 gnd.n3149 9.3005
R10341 gnd.n2854 gnd.n2853 9.3005
R10342 gnd.n3177 gnd.n3176 9.3005
R10343 gnd.n3178 gnd.n2852 9.3005
R10344 gnd.n3182 gnd.n3179 9.3005
R10345 gnd.n3181 gnd.n3180 9.3005
R10346 gnd.n2826 gnd.n2825 9.3005
R10347 gnd.n3207 gnd.n3206 9.3005
R10348 gnd.n3208 gnd.n2824 9.3005
R10349 gnd.n3210 gnd.n3209 9.3005
R10350 gnd.n2804 gnd.n2803 9.3005
R10351 gnd.n3238 gnd.n3237 9.3005
R10352 gnd.n3239 gnd.n2802 9.3005
R10353 gnd.n3247 gnd.n3240 9.3005
R10354 gnd.n3246 gnd.n3241 9.3005
R10355 gnd.n3245 gnd.n3243 9.3005
R10356 gnd.n3242 gnd.n2751 9.3005
R10357 gnd.n3295 gnd.n2752 9.3005
R10358 gnd.n3294 gnd.n2753 9.3005
R10359 gnd.n3293 gnd.n2754 9.3005
R10360 gnd.n2773 gnd.n2755 9.3005
R10361 gnd.n2775 gnd.n2774 9.3005
R10362 gnd.n2673 gnd.n2672 9.3005
R10363 gnd.n3333 gnd.n3332 9.3005
R10364 gnd.n3334 gnd.n2671 9.3005
R10365 gnd.n3338 gnd.n3335 9.3005
R10366 gnd.n3337 gnd.n3336 9.3005
R10367 gnd.n2646 gnd.n2645 9.3005
R10368 gnd.n3373 gnd.n3372 9.3005
R10369 gnd.n3374 gnd.n2644 9.3005
R10370 gnd.n3378 gnd.n3375 9.3005
R10371 gnd.n3377 gnd.n3376 9.3005
R10372 gnd.n2619 gnd.n2618 9.3005
R10373 gnd.n3418 gnd.n3417 9.3005
R10374 gnd.n3419 gnd.n2617 9.3005
R10375 gnd.n3423 gnd.n3420 9.3005
R10376 gnd.n3422 gnd.n3421 9.3005
R10377 gnd.n2591 gnd.n2590 9.3005
R10378 gnd.n3458 gnd.n3457 9.3005
R10379 gnd.n3459 gnd.n2589 9.3005
R10380 gnd.n3463 gnd.n3460 9.3005
R10381 gnd.n3462 gnd.n3461 9.3005
R10382 gnd.n2564 gnd.n2563 9.3005
R10383 gnd.n3507 gnd.n3506 9.3005
R10384 gnd.n3508 gnd.n2562 9.3005
R10385 gnd.n3512 gnd.n3509 9.3005
R10386 gnd.n3511 gnd.n3510 9.3005
R10387 gnd.n2537 gnd.n2536 9.3005
R10388 gnd.n3801 gnd.n3800 9.3005
R10389 gnd.n3802 gnd.n2535 9.3005
R10390 gnd.n3808 gnd.n3803 9.3005
R10391 gnd.n3807 gnd.n3804 9.3005
R10392 gnd.n3806 gnd.n3805 9.3005
R10393 gnd.n3151 gnd.n3148 9.3005
R10394 gnd.n2933 gnd.n2892 9.3005
R10395 gnd.n2928 gnd.n2927 9.3005
R10396 gnd.n2926 gnd.n2893 9.3005
R10397 gnd.n2925 gnd.n2924 9.3005
R10398 gnd.n2921 gnd.n2894 9.3005
R10399 gnd.n2918 gnd.n2917 9.3005
R10400 gnd.n2916 gnd.n2895 9.3005
R10401 gnd.n2915 gnd.n2914 9.3005
R10402 gnd.n2911 gnd.n2896 9.3005
R10403 gnd.n2908 gnd.n2907 9.3005
R10404 gnd.n2906 gnd.n2897 9.3005
R10405 gnd.n2905 gnd.n2904 9.3005
R10406 gnd.n2901 gnd.n2899 9.3005
R10407 gnd.n2898 gnd.n2878 9.3005
R10408 gnd.n3145 gnd.n2877 9.3005
R10409 gnd.n3147 gnd.n3146 9.3005
R10410 gnd.n2935 gnd.n2934 9.3005
R10411 gnd.n3158 gnd.n2864 9.3005
R10412 gnd.n3165 gnd.n2865 9.3005
R10413 gnd.n3167 gnd.n3166 9.3005
R10414 gnd.n3168 gnd.n2845 9.3005
R10415 gnd.n3187 gnd.n3186 9.3005
R10416 gnd.n3189 gnd.n2837 9.3005
R10417 gnd.n3196 gnd.n2839 9.3005
R10418 gnd.n3197 gnd.n2834 9.3005
R10419 gnd.n3199 gnd.n3198 9.3005
R10420 gnd.n2835 gnd.n2820 9.3005
R10421 gnd.n3215 gnd.n2818 9.3005
R10422 gnd.n3219 gnd.n3218 9.3005
R10423 gnd.n3217 gnd.n2794 9.3005
R10424 gnd.n3254 gnd.n2793 9.3005
R10425 gnd.n3257 gnd.n3256 9.3005
R10426 gnd.n2790 gnd.n2789 9.3005
R10427 gnd.n3263 gnd.n2791 9.3005
R10428 gnd.n3265 gnd.n3264 9.3005
R10429 gnd.n3267 gnd.n2788 9.3005
R10430 gnd.n3270 gnd.n3269 9.3005
R10431 gnd.n3273 gnd.n3271 9.3005
R10432 gnd.n3275 gnd.n3274 9.3005
R10433 gnd.n3281 gnd.n3276 9.3005
R10434 gnd.n3280 gnd.n3279 9.3005
R10435 gnd.n2664 gnd.n2663 9.3005
R10436 gnd.n3347 gnd.n3346 9.3005
R10437 gnd.n3348 gnd.n2657 9.3005
R10438 gnd.n3356 gnd.n2656 9.3005
R10439 gnd.n3359 gnd.n3358 9.3005
R10440 gnd.n3361 gnd.n3360 9.3005
R10441 gnd.n3364 gnd.n2639 9.3005
R10442 gnd.n3362 gnd.n2637 9.3005
R10443 gnd.n3384 gnd.n2635 9.3005
R10444 gnd.n3386 gnd.n3385 9.3005
R10445 gnd.n2609 gnd.n2608 9.3005
R10446 gnd.n3432 gnd.n3431 9.3005
R10447 gnd.n3433 gnd.n2602 9.3005
R10448 gnd.n3441 gnd.n2601 9.3005
R10449 gnd.n3444 gnd.n3443 9.3005
R10450 gnd.n3446 gnd.n3445 9.3005
R10451 gnd.n3449 gnd.n2584 9.3005
R10452 gnd.n3447 gnd.n2582 9.3005
R10453 gnd.n3469 gnd.n2580 9.3005
R10454 gnd.n3471 gnd.n3470 9.3005
R10455 gnd.n2555 gnd.n2554 9.3005
R10456 gnd.n3521 gnd.n3520 9.3005
R10457 gnd.n3522 gnd.n2548 9.3005
R10458 gnd.n3530 gnd.n2547 9.3005
R10459 gnd.n3789 gnd.n3788 9.3005
R10460 gnd.n3791 gnd.n3790 9.3005
R10461 gnd.n3792 gnd.n2528 9.3005
R10462 gnd.n3816 gnd.n3815 9.3005
R10463 gnd.n2529 gnd.n2491 9.3005
R10464 gnd.n3156 gnd.n3155 9.3005
R10465 gnd.n3872 gnd.n2492 9.3005
R10466 gnd.n3871 gnd.n2494 9.3005
R10467 gnd.n3868 gnd.n2495 9.3005
R10468 gnd.n3867 gnd.n2496 9.3005
R10469 gnd.n3864 gnd.n2497 9.3005
R10470 gnd.n3863 gnd.n2498 9.3005
R10471 gnd.n3860 gnd.n2499 9.3005
R10472 gnd.n3859 gnd.n2500 9.3005
R10473 gnd.n3856 gnd.n2501 9.3005
R10474 gnd.n3855 gnd.n2502 9.3005
R10475 gnd.n3852 gnd.n2503 9.3005
R10476 gnd.n3851 gnd.n2504 9.3005
R10477 gnd.n3848 gnd.n2505 9.3005
R10478 gnd.n3847 gnd.n2506 9.3005
R10479 gnd.n3844 gnd.n2507 9.3005
R10480 gnd.n3843 gnd.n2508 9.3005
R10481 gnd.n3840 gnd.n2509 9.3005
R10482 gnd.n3839 gnd.n2510 9.3005
R10483 gnd.n3836 gnd.n2511 9.3005
R10484 gnd.n3835 gnd.n2512 9.3005
R10485 gnd.n3832 gnd.n2513 9.3005
R10486 gnd.n3831 gnd.n2514 9.3005
R10487 gnd.n3828 gnd.n2518 9.3005
R10488 gnd.n3827 gnd.n2519 9.3005
R10489 gnd.n3824 gnd.n2520 9.3005
R10490 gnd.n3823 gnd.n2521 9.3005
R10491 gnd.n3874 gnd.n3873 9.3005
R10492 gnd.n3325 gnd.n3309 9.3005
R10493 gnd.n3324 gnd.n3310 9.3005
R10494 gnd.n3323 gnd.n3311 9.3005
R10495 gnd.n3321 gnd.n3312 9.3005
R10496 gnd.n3320 gnd.n3313 9.3005
R10497 gnd.n3318 gnd.n3314 9.3005
R10498 gnd.n3317 gnd.n3315 9.3005
R10499 gnd.n2627 gnd.n2626 9.3005
R10500 gnd.n3394 gnd.n3393 9.3005
R10501 gnd.n3395 gnd.n2625 9.3005
R10502 gnd.n3412 gnd.n3396 9.3005
R10503 gnd.n3411 gnd.n3397 9.3005
R10504 gnd.n3410 gnd.n3398 9.3005
R10505 gnd.n3408 gnd.n3399 9.3005
R10506 gnd.n3407 gnd.n3400 9.3005
R10507 gnd.n3405 gnd.n3401 9.3005
R10508 gnd.n3404 gnd.n3402 9.3005
R10509 gnd.n2571 gnd.n2570 9.3005
R10510 gnd.n3479 gnd.n3478 9.3005
R10511 gnd.n3480 gnd.n2569 9.3005
R10512 gnd.n3501 gnd.n3481 9.3005
R10513 gnd.n3500 gnd.n3482 9.3005
R10514 gnd.n3499 gnd.n3483 9.3005
R10515 gnd.n3496 gnd.n3484 9.3005
R10516 gnd.n3495 gnd.n3485 9.3005
R10517 gnd.n3493 gnd.n3486 9.3005
R10518 gnd.n3492 gnd.n3487 9.3005
R10519 gnd.n3490 gnd.n3489 9.3005
R10520 gnd.n3488 gnd.n2523 9.3005
R10521 gnd.n3066 gnd.n3065 9.3005
R10522 gnd.n2956 gnd.n2955 9.3005
R10523 gnd.n3080 gnd.n3079 9.3005
R10524 gnd.n3081 gnd.n2954 9.3005
R10525 gnd.n3083 gnd.n3082 9.3005
R10526 gnd.n2944 gnd.n2943 9.3005
R10527 gnd.n3096 gnd.n3095 9.3005
R10528 gnd.n3097 gnd.n2942 9.3005
R10529 gnd.n3129 gnd.n3098 9.3005
R10530 gnd.n3128 gnd.n3099 9.3005
R10531 gnd.n3127 gnd.n3100 9.3005
R10532 gnd.n3126 gnd.n3101 9.3005
R10533 gnd.n3123 gnd.n3102 9.3005
R10534 gnd.n3122 gnd.n3103 9.3005
R10535 gnd.n3121 gnd.n3104 9.3005
R10536 gnd.n3119 gnd.n3105 9.3005
R10537 gnd.n3118 gnd.n3106 9.3005
R10538 gnd.n3115 gnd.n3107 9.3005
R10539 gnd.n3114 gnd.n3108 9.3005
R10540 gnd.n3113 gnd.n3109 9.3005
R10541 gnd.n3111 gnd.n3110 9.3005
R10542 gnd.n2810 gnd.n2809 9.3005
R10543 gnd.n3227 gnd.n3226 9.3005
R10544 gnd.n3228 gnd.n2808 9.3005
R10545 gnd.n3232 gnd.n3229 9.3005
R10546 gnd.n3231 gnd.n3230 9.3005
R10547 gnd.n2732 gnd.n2731 9.3005
R10548 gnd.n3307 gnd.n3306 9.3005
R10549 gnd.n3064 gnd.n2965 9.3005
R10550 gnd.n2967 gnd.n2966 9.3005
R10551 gnd.n3011 gnd.n3009 9.3005
R10552 gnd.n3012 gnd.n3008 9.3005
R10553 gnd.n3015 gnd.n3004 9.3005
R10554 gnd.n3016 gnd.n3003 9.3005
R10555 gnd.n3019 gnd.n3002 9.3005
R10556 gnd.n3020 gnd.n3001 9.3005
R10557 gnd.n3023 gnd.n3000 9.3005
R10558 gnd.n3024 gnd.n2999 9.3005
R10559 gnd.n3027 gnd.n2998 9.3005
R10560 gnd.n3028 gnd.n2997 9.3005
R10561 gnd.n3031 gnd.n2996 9.3005
R10562 gnd.n3032 gnd.n2995 9.3005
R10563 gnd.n3035 gnd.n2994 9.3005
R10564 gnd.n3036 gnd.n2993 9.3005
R10565 gnd.n3039 gnd.n2992 9.3005
R10566 gnd.n3040 gnd.n2991 9.3005
R10567 gnd.n3043 gnd.n2990 9.3005
R10568 gnd.n3044 gnd.n2989 9.3005
R10569 gnd.n3047 gnd.n2988 9.3005
R10570 gnd.n3048 gnd.n2987 9.3005
R10571 gnd.n3051 gnd.n2986 9.3005
R10572 gnd.n3053 gnd.n2985 9.3005
R10573 gnd.n3054 gnd.n2984 9.3005
R10574 gnd.n3055 gnd.n2983 9.3005
R10575 gnd.n3056 gnd.n2982 9.3005
R10576 gnd.n3063 gnd.n3062 9.3005
R10577 gnd.n3072 gnd.n3071 9.3005
R10578 gnd.n3073 gnd.n2959 9.3005
R10579 gnd.n3075 gnd.n3074 9.3005
R10580 gnd.n2950 gnd.n2949 9.3005
R10581 gnd.n3088 gnd.n3087 9.3005
R10582 gnd.n3089 gnd.n2948 9.3005
R10583 gnd.n3091 gnd.n3090 9.3005
R10584 gnd.n2937 gnd.n2936 9.3005
R10585 gnd.n3134 gnd.n3133 9.3005
R10586 gnd.n3135 gnd.n2891 9.3005
R10587 gnd.n3139 gnd.n3137 9.3005
R10588 gnd.n3138 gnd.n2870 9.3005
R10589 gnd.n3157 gnd.n2869 9.3005
R10590 gnd.n3160 gnd.n3159 9.3005
R10591 gnd.n2863 gnd.n2862 9.3005
R10592 gnd.n3171 gnd.n3169 9.3005
R10593 gnd.n3170 gnd.n2844 9.3005
R10594 gnd.n3188 gnd.n2843 9.3005
R10595 gnd.n3191 gnd.n3190 9.3005
R10596 gnd.n2838 gnd.n2833 9.3005
R10597 gnd.n3201 gnd.n3200 9.3005
R10598 gnd.n2836 gnd.n2816 9.3005
R10599 gnd.n3222 gnd.n2817 9.3005
R10600 gnd.n3221 gnd.n3220 9.3005
R10601 gnd.n2819 gnd.n2795 9.3005
R10602 gnd.n3253 gnd.n3252 9.3005
R10603 gnd.n3255 gnd.n2740 9.3005
R10604 gnd.n3302 gnd.n2741 9.3005
R10605 gnd.n3301 gnd.n2742 9.3005
R10606 gnd.n3300 gnd.n2743 9.3005
R10607 gnd.n3266 gnd.n2744 9.3005
R10608 gnd.n3268 gnd.n2762 9.3005
R10609 gnd.n3288 gnd.n2763 9.3005
R10610 gnd.n3287 gnd.n2764 9.3005
R10611 gnd.n3286 gnd.n2765 9.3005
R10612 gnd.n3277 gnd.n2766 9.3005
R10613 gnd.n3278 gnd.n2665 9.3005
R10614 gnd.n3344 gnd.n3343 9.3005
R10615 gnd.n3345 gnd.n2658 9.3005
R10616 gnd.n3355 gnd.n3354 9.3005
R10617 gnd.n3357 gnd.n2654 9.3005
R10618 gnd.n3367 gnd.n2655 9.3005
R10619 gnd.n3366 gnd.n3365 9.3005
R10620 gnd.n3363 gnd.n2633 9.3005
R10621 gnd.n3389 gnd.n2634 9.3005
R10622 gnd.n3388 gnd.n3387 9.3005
R10623 gnd.n2636 gnd.n2610 9.3005
R10624 gnd.n3429 gnd.n3428 9.3005
R10625 gnd.n3430 gnd.n2603 9.3005
R10626 gnd.n3440 gnd.n3439 9.3005
R10627 gnd.n3442 gnd.n2599 9.3005
R10628 gnd.n3452 gnd.n2600 9.3005
R10629 gnd.n3451 gnd.n3450 9.3005
R10630 gnd.n3448 gnd.n2578 9.3005
R10631 gnd.n3474 gnd.n2579 9.3005
R10632 gnd.n3473 gnd.n3472 9.3005
R10633 gnd.n2581 gnd.n2556 9.3005
R10634 gnd.n3518 gnd.n3517 9.3005
R10635 gnd.n3519 gnd.n2549 9.3005
R10636 gnd.n3529 gnd.n3528 9.3005
R10637 gnd.n3787 gnd.n2545 9.3005
R10638 gnd.n3795 gnd.n2546 9.3005
R10639 gnd.n3794 gnd.n3793 9.3005
R10640 gnd.n2527 gnd.n2526 9.3005
R10641 gnd.n3818 gnd.n3817 9.3005
R10642 gnd.n2961 gnd.n2960 9.3005
R10643 gnd.n6482 gnd.n6481 9.3005
R10644 gnd.n793 gnd.n792 9.3005
R10645 gnd.n6489 gnd.n6488 9.3005
R10646 gnd.n6490 gnd.n791 9.3005
R10647 gnd.n6492 gnd.n6491 9.3005
R10648 gnd.n787 gnd.n786 9.3005
R10649 gnd.n6499 gnd.n6498 9.3005
R10650 gnd.n6500 gnd.n785 9.3005
R10651 gnd.n6502 gnd.n6501 9.3005
R10652 gnd.n781 gnd.n780 9.3005
R10653 gnd.n6509 gnd.n6508 9.3005
R10654 gnd.n6510 gnd.n779 9.3005
R10655 gnd.n6512 gnd.n6511 9.3005
R10656 gnd.n775 gnd.n774 9.3005
R10657 gnd.n6519 gnd.n6518 9.3005
R10658 gnd.n6520 gnd.n773 9.3005
R10659 gnd.n6522 gnd.n6521 9.3005
R10660 gnd.n769 gnd.n768 9.3005
R10661 gnd.n6529 gnd.n6528 9.3005
R10662 gnd.n6530 gnd.n767 9.3005
R10663 gnd.n6532 gnd.n6531 9.3005
R10664 gnd.n763 gnd.n762 9.3005
R10665 gnd.n6539 gnd.n6538 9.3005
R10666 gnd.n6540 gnd.n761 9.3005
R10667 gnd.n6542 gnd.n6541 9.3005
R10668 gnd.n757 gnd.n756 9.3005
R10669 gnd.n6549 gnd.n6548 9.3005
R10670 gnd.n6550 gnd.n755 9.3005
R10671 gnd.n6552 gnd.n6551 9.3005
R10672 gnd.n751 gnd.n750 9.3005
R10673 gnd.n6559 gnd.n6558 9.3005
R10674 gnd.n6560 gnd.n749 9.3005
R10675 gnd.n6562 gnd.n6561 9.3005
R10676 gnd.n745 gnd.n744 9.3005
R10677 gnd.n6569 gnd.n6568 9.3005
R10678 gnd.n6570 gnd.n743 9.3005
R10679 gnd.n6572 gnd.n6571 9.3005
R10680 gnd.n739 gnd.n738 9.3005
R10681 gnd.n6579 gnd.n6578 9.3005
R10682 gnd.n6580 gnd.n737 9.3005
R10683 gnd.n6582 gnd.n6581 9.3005
R10684 gnd.n733 gnd.n732 9.3005
R10685 gnd.n6589 gnd.n6588 9.3005
R10686 gnd.n6590 gnd.n731 9.3005
R10687 gnd.n6592 gnd.n6591 9.3005
R10688 gnd.n727 gnd.n726 9.3005
R10689 gnd.n6599 gnd.n6598 9.3005
R10690 gnd.n6600 gnd.n725 9.3005
R10691 gnd.n6602 gnd.n6601 9.3005
R10692 gnd.n721 gnd.n720 9.3005
R10693 gnd.n6609 gnd.n6608 9.3005
R10694 gnd.n6610 gnd.n719 9.3005
R10695 gnd.n6612 gnd.n6611 9.3005
R10696 gnd.n715 gnd.n714 9.3005
R10697 gnd.n6619 gnd.n6618 9.3005
R10698 gnd.n6620 gnd.n713 9.3005
R10699 gnd.n6622 gnd.n6621 9.3005
R10700 gnd.n709 gnd.n708 9.3005
R10701 gnd.n6629 gnd.n6628 9.3005
R10702 gnd.n6630 gnd.n707 9.3005
R10703 gnd.n6632 gnd.n6631 9.3005
R10704 gnd.n703 gnd.n702 9.3005
R10705 gnd.n6639 gnd.n6638 9.3005
R10706 gnd.n6640 gnd.n701 9.3005
R10707 gnd.n6642 gnd.n6641 9.3005
R10708 gnd.n697 gnd.n696 9.3005
R10709 gnd.n6649 gnd.n6648 9.3005
R10710 gnd.n6650 gnd.n695 9.3005
R10711 gnd.n6652 gnd.n6651 9.3005
R10712 gnd.n691 gnd.n690 9.3005
R10713 gnd.n6659 gnd.n6658 9.3005
R10714 gnd.n6660 gnd.n689 9.3005
R10715 gnd.n6662 gnd.n6661 9.3005
R10716 gnd.n685 gnd.n684 9.3005
R10717 gnd.n6669 gnd.n6668 9.3005
R10718 gnd.n6670 gnd.n683 9.3005
R10719 gnd.n6672 gnd.n6671 9.3005
R10720 gnd.n679 gnd.n678 9.3005
R10721 gnd.n6679 gnd.n6678 9.3005
R10722 gnd.n6680 gnd.n677 9.3005
R10723 gnd.n6682 gnd.n6681 9.3005
R10724 gnd.n673 gnd.n672 9.3005
R10725 gnd.n6689 gnd.n6688 9.3005
R10726 gnd.n6690 gnd.n671 9.3005
R10727 gnd.n6692 gnd.n6691 9.3005
R10728 gnd.n667 gnd.n666 9.3005
R10729 gnd.n6699 gnd.n6698 9.3005
R10730 gnd.n6700 gnd.n665 9.3005
R10731 gnd.n6702 gnd.n6701 9.3005
R10732 gnd.n661 gnd.n660 9.3005
R10733 gnd.n6709 gnd.n6708 9.3005
R10734 gnd.n6710 gnd.n659 9.3005
R10735 gnd.n6712 gnd.n6711 9.3005
R10736 gnd.n655 gnd.n654 9.3005
R10737 gnd.n6719 gnd.n6718 9.3005
R10738 gnd.n6720 gnd.n653 9.3005
R10739 gnd.n6722 gnd.n6721 9.3005
R10740 gnd.n649 gnd.n648 9.3005
R10741 gnd.n6729 gnd.n6728 9.3005
R10742 gnd.n6730 gnd.n647 9.3005
R10743 gnd.n6732 gnd.n6731 9.3005
R10744 gnd.n643 gnd.n642 9.3005
R10745 gnd.n6739 gnd.n6738 9.3005
R10746 gnd.n6740 gnd.n641 9.3005
R10747 gnd.n6742 gnd.n6741 9.3005
R10748 gnd.n637 gnd.n636 9.3005
R10749 gnd.n6749 gnd.n6748 9.3005
R10750 gnd.n6750 gnd.n635 9.3005
R10751 gnd.n6752 gnd.n6751 9.3005
R10752 gnd.n631 gnd.n630 9.3005
R10753 gnd.n6759 gnd.n6758 9.3005
R10754 gnd.n6760 gnd.n629 9.3005
R10755 gnd.n6762 gnd.n6761 9.3005
R10756 gnd.n625 gnd.n624 9.3005
R10757 gnd.n6769 gnd.n6768 9.3005
R10758 gnd.n6770 gnd.n623 9.3005
R10759 gnd.n6772 gnd.n6771 9.3005
R10760 gnd.n619 gnd.n618 9.3005
R10761 gnd.n6779 gnd.n6778 9.3005
R10762 gnd.n6780 gnd.n617 9.3005
R10763 gnd.n6782 gnd.n6781 9.3005
R10764 gnd.n613 gnd.n612 9.3005
R10765 gnd.n6789 gnd.n6788 9.3005
R10766 gnd.n6790 gnd.n611 9.3005
R10767 gnd.n6792 gnd.n6791 9.3005
R10768 gnd.n607 gnd.n606 9.3005
R10769 gnd.n6799 gnd.n6798 9.3005
R10770 gnd.n6800 gnd.n605 9.3005
R10771 gnd.n6802 gnd.n6801 9.3005
R10772 gnd.n601 gnd.n600 9.3005
R10773 gnd.n6809 gnd.n6808 9.3005
R10774 gnd.n6810 gnd.n599 9.3005
R10775 gnd.n6812 gnd.n6811 9.3005
R10776 gnd.n595 gnd.n594 9.3005
R10777 gnd.n6819 gnd.n6818 9.3005
R10778 gnd.n6820 gnd.n593 9.3005
R10779 gnd.n6822 gnd.n6821 9.3005
R10780 gnd.n589 gnd.n588 9.3005
R10781 gnd.n6829 gnd.n6828 9.3005
R10782 gnd.n6830 gnd.n587 9.3005
R10783 gnd.n6832 gnd.n6831 9.3005
R10784 gnd.n583 gnd.n582 9.3005
R10785 gnd.n6839 gnd.n6838 9.3005
R10786 gnd.n6840 gnd.n581 9.3005
R10787 gnd.n6842 gnd.n6841 9.3005
R10788 gnd.n577 gnd.n576 9.3005
R10789 gnd.n6849 gnd.n6848 9.3005
R10790 gnd.n6850 gnd.n575 9.3005
R10791 gnd.n6852 gnd.n6851 9.3005
R10792 gnd.n571 gnd.n570 9.3005
R10793 gnd.n6859 gnd.n6858 9.3005
R10794 gnd.n6860 gnd.n569 9.3005
R10795 gnd.n6862 gnd.n6861 9.3005
R10796 gnd.n565 gnd.n564 9.3005
R10797 gnd.n6869 gnd.n6868 9.3005
R10798 gnd.n6870 gnd.n563 9.3005
R10799 gnd.n6872 gnd.n6871 9.3005
R10800 gnd.n559 gnd.n558 9.3005
R10801 gnd.n6879 gnd.n6878 9.3005
R10802 gnd.n6880 gnd.n557 9.3005
R10803 gnd.n6882 gnd.n6881 9.3005
R10804 gnd.n553 gnd.n552 9.3005
R10805 gnd.n6889 gnd.n6888 9.3005
R10806 gnd.n6890 gnd.n551 9.3005
R10807 gnd.n6893 gnd.n6892 9.3005
R10808 gnd.n6891 gnd.n547 9.3005
R10809 gnd.n6899 gnd.n546 9.3005
R10810 gnd.n6901 gnd.n6900 9.3005
R10811 gnd.n542 gnd.n541 9.3005
R10812 gnd.n6910 gnd.n6909 9.3005
R10813 gnd.n6911 gnd.n540 9.3005
R10814 gnd.n6913 gnd.n6912 9.3005
R10815 gnd.n536 gnd.n535 9.3005
R10816 gnd.n6920 gnd.n6919 9.3005
R10817 gnd.n6921 gnd.n534 9.3005
R10818 gnd.n6923 gnd.n6922 9.3005
R10819 gnd.n530 gnd.n529 9.3005
R10820 gnd.n6930 gnd.n6929 9.3005
R10821 gnd.n6931 gnd.n528 9.3005
R10822 gnd.n6933 gnd.n6932 9.3005
R10823 gnd.n524 gnd.n523 9.3005
R10824 gnd.n6940 gnd.n6939 9.3005
R10825 gnd.n6941 gnd.n522 9.3005
R10826 gnd.n6943 gnd.n6942 9.3005
R10827 gnd.n518 gnd.n517 9.3005
R10828 gnd.n6950 gnd.n6949 9.3005
R10829 gnd.n6951 gnd.n516 9.3005
R10830 gnd.n6953 gnd.n6952 9.3005
R10831 gnd.n512 gnd.n511 9.3005
R10832 gnd.n6960 gnd.n6959 9.3005
R10833 gnd.n6961 gnd.n510 9.3005
R10834 gnd.n6963 gnd.n6962 9.3005
R10835 gnd.n506 gnd.n505 9.3005
R10836 gnd.n6970 gnd.n6969 9.3005
R10837 gnd.n6971 gnd.n504 9.3005
R10838 gnd.n6973 gnd.n6972 9.3005
R10839 gnd.n500 gnd.n499 9.3005
R10840 gnd.n6980 gnd.n6979 9.3005
R10841 gnd.n6981 gnd.n498 9.3005
R10842 gnd.n6983 gnd.n6982 9.3005
R10843 gnd.n494 gnd.n493 9.3005
R10844 gnd.n6990 gnd.n6989 9.3005
R10845 gnd.n6991 gnd.n492 9.3005
R10846 gnd.n6993 gnd.n6992 9.3005
R10847 gnd.n488 gnd.n487 9.3005
R10848 gnd.n7000 gnd.n6999 9.3005
R10849 gnd.n7001 gnd.n486 9.3005
R10850 gnd.n7003 gnd.n7002 9.3005
R10851 gnd.n482 gnd.n481 9.3005
R10852 gnd.n7010 gnd.n7009 9.3005
R10853 gnd.n7011 gnd.n480 9.3005
R10854 gnd.n7013 gnd.n7012 9.3005
R10855 gnd.n476 gnd.n475 9.3005
R10856 gnd.n7020 gnd.n7019 9.3005
R10857 gnd.n7021 gnd.n474 9.3005
R10858 gnd.n7023 gnd.n7022 9.3005
R10859 gnd.n470 gnd.n469 9.3005
R10860 gnd.n7030 gnd.n7029 9.3005
R10861 gnd.n7031 gnd.n468 9.3005
R10862 gnd.n7033 gnd.n7032 9.3005
R10863 gnd.n464 gnd.n463 9.3005
R10864 gnd.n7040 gnd.n7039 9.3005
R10865 gnd.n7041 gnd.n462 9.3005
R10866 gnd.n7043 gnd.n7042 9.3005
R10867 gnd.n458 gnd.n457 9.3005
R10868 gnd.n7050 gnd.n7049 9.3005
R10869 gnd.n7051 gnd.n456 9.3005
R10870 gnd.n7053 gnd.n7052 9.3005
R10871 gnd.n452 gnd.n451 9.3005
R10872 gnd.n7060 gnd.n7059 9.3005
R10873 gnd.n7061 gnd.n450 9.3005
R10874 gnd.n7063 gnd.n7062 9.3005
R10875 gnd.n446 gnd.n445 9.3005
R10876 gnd.n7070 gnd.n7069 9.3005
R10877 gnd.n7071 gnd.n444 9.3005
R10878 gnd.n7073 gnd.n7072 9.3005
R10879 gnd.n440 gnd.n439 9.3005
R10880 gnd.n7080 gnd.n7079 9.3005
R10881 gnd.n7081 gnd.n438 9.3005
R10882 gnd.n7083 gnd.n7082 9.3005
R10883 gnd.n434 gnd.n433 9.3005
R10884 gnd.n7090 gnd.n7089 9.3005
R10885 gnd.n7091 gnd.n432 9.3005
R10886 gnd.n7093 gnd.n7092 9.3005
R10887 gnd.n428 gnd.n427 9.3005
R10888 gnd.n7100 gnd.n7099 9.3005
R10889 gnd.n7101 gnd.n426 9.3005
R10890 gnd.n7103 gnd.n7102 9.3005
R10891 gnd.n422 gnd.n421 9.3005
R10892 gnd.n7111 gnd.n7110 9.3005
R10893 gnd.n7112 gnd.n420 9.3005
R10894 gnd.n7115 gnd.n7114 9.3005
R10895 gnd.n6903 gnd.n6902 9.3005
R10896 gnd.n7343 gnd.n7342 9.3005
R10897 gnd.n7341 gnd.n65 9.3005
R10898 gnd.n397 gnd.n67 9.3005
R10899 gnd.n7147 gnd.n7146 9.3005
R10900 gnd.n7148 gnd.n396 9.3005
R10901 gnd.n7150 gnd.n7149 9.3005
R10902 gnd.n394 gnd.n393 9.3005
R10903 gnd.n7162 gnd.n7161 9.3005
R10904 gnd.n7163 gnd.n392 9.3005
R10905 gnd.n7165 gnd.n7164 9.3005
R10906 gnd.n389 gnd.n388 9.3005
R10907 gnd.n7177 gnd.n7176 9.3005
R10908 gnd.n7178 gnd.n387 9.3005
R10909 gnd.n7264 gnd.n7179 9.3005
R10910 gnd.n7263 gnd.n7180 9.3005
R10911 gnd.n7262 gnd.n7181 9.3005
R10912 gnd.n7260 gnd.n7182 9.3005
R10913 gnd.n7259 gnd.n7183 9.3005
R10914 gnd.n7257 gnd.n7184 9.3005
R10915 gnd.n7256 gnd.n7185 9.3005
R10916 gnd.n7254 gnd.n7253 9.3005
R10917 gnd.n7207 gnd.n7204 9.3005
R10918 gnd.n7213 gnd.n7212 9.3005
R10919 gnd.n7214 gnd.n7203 9.3005
R10920 gnd.n7216 gnd.n7215 9.3005
R10921 gnd.n7201 gnd.n7200 9.3005
R10922 gnd.n7223 gnd.n7222 9.3005
R10923 gnd.n7224 gnd.n7199 9.3005
R10924 gnd.n7226 gnd.n7225 9.3005
R10925 gnd.n7197 gnd.n7196 9.3005
R10926 gnd.n7233 gnd.n7232 9.3005
R10927 gnd.n7234 gnd.n7195 9.3005
R10928 gnd.n7236 gnd.n7235 9.3005
R10929 gnd.n7193 gnd.n7192 9.3005
R10930 gnd.n7243 gnd.n7242 9.3005
R10931 gnd.n7244 gnd.n7191 9.3005
R10932 gnd.n7246 gnd.n7245 9.3005
R10933 gnd.n7189 gnd.n7186 9.3005
R10934 gnd.n7252 gnd.n7251 9.3005
R10935 gnd.n7206 gnd.n7205 9.3005
R10936 gnd.n238 gnd.n235 9.3005
R10937 gnd.n244 gnd.n243 9.3005
R10938 gnd.n245 gnd.n234 9.3005
R10939 gnd.n247 gnd.n246 9.3005
R10940 gnd.n232 gnd.n231 9.3005
R10941 gnd.n254 gnd.n253 9.3005
R10942 gnd.n255 gnd.n230 9.3005
R10943 gnd.n257 gnd.n256 9.3005
R10944 gnd.n228 gnd.n227 9.3005
R10945 gnd.n264 gnd.n263 9.3005
R10946 gnd.n265 gnd.n226 9.3005
R10947 gnd.n267 gnd.n266 9.3005
R10948 gnd.n224 gnd.n223 9.3005
R10949 gnd.n275 gnd.n274 9.3005
R10950 gnd.n276 gnd.n222 9.3005
R10951 gnd.n278 gnd.n277 9.3005
R10952 gnd.n279 gnd.n217 9.3005
R10953 gnd.n285 gnd.n284 9.3005
R10954 gnd.n286 gnd.n216 9.3005
R10955 gnd.n288 gnd.n287 9.3005
R10956 gnd.n214 gnd.n213 9.3005
R10957 gnd.n295 gnd.n294 9.3005
R10958 gnd.n296 gnd.n212 9.3005
R10959 gnd.n298 gnd.n297 9.3005
R10960 gnd.n210 gnd.n209 9.3005
R10961 gnd.n305 gnd.n304 9.3005
R10962 gnd.n306 gnd.n208 9.3005
R10963 gnd.n308 gnd.n307 9.3005
R10964 gnd.n206 gnd.n205 9.3005
R10965 gnd.n315 gnd.n314 9.3005
R10966 gnd.n316 gnd.n204 9.3005
R10967 gnd.n318 gnd.n317 9.3005
R10968 gnd.n202 gnd.n201 9.3005
R10969 gnd.n325 gnd.n324 9.3005
R10970 gnd.n326 gnd.n200 9.3005
R10971 gnd.n328 gnd.n327 9.3005
R10972 gnd.n198 gnd.n195 9.3005
R10973 gnd.n335 gnd.n334 9.3005
R10974 gnd.n336 gnd.n194 9.3005
R10975 gnd.n338 gnd.n337 9.3005
R10976 gnd.n192 gnd.n191 9.3005
R10977 gnd.n345 gnd.n344 9.3005
R10978 gnd.n346 gnd.n190 9.3005
R10979 gnd.n348 gnd.n347 9.3005
R10980 gnd.n188 gnd.n187 9.3005
R10981 gnd.n355 gnd.n354 9.3005
R10982 gnd.n356 gnd.n186 9.3005
R10983 gnd.n358 gnd.n357 9.3005
R10984 gnd.n184 gnd.n183 9.3005
R10985 gnd.n365 gnd.n364 9.3005
R10986 gnd.n366 gnd.n182 9.3005
R10987 gnd.n368 gnd.n367 9.3005
R10988 gnd.n180 gnd.n179 9.3005
R10989 gnd.n375 gnd.n374 9.3005
R10990 gnd.n376 gnd.n178 9.3005
R10991 gnd.n378 gnd.n377 9.3005
R10992 gnd.n176 gnd.n173 9.3005
R10993 gnd.n384 gnd.n383 9.3005
R10994 gnd.n237 gnd.n236 9.3005
R10995 gnd.n5664 gnd.n1624 9.3005
R10996 gnd.n5850 gnd.n1625 9.3005
R10997 gnd.n5849 gnd.n1626 9.3005
R10998 gnd.n5848 gnd.n1627 9.3005
R10999 gnd.n1747 gnd.n1628 9.3005
R11000 gnd.n5838 gnd.n1645 9.3005
R11001 gnd.n5837 gnd.n1646 9.3005
R11002 gnd.n5836 gnd.n1647 9.3005
R11003 gnd.n5683 gnd.n1648 9.3005
R11004 gnd.n5826 gnd.n1666 9.3005
R11005 gnd.n5825 gnd.n1667 9.3005
R11006 gnd.n5824 gnd.n1668 9.3005
R11007 gnd.n5746 gnd.n1669 9.3005
R11008 gnd.n5814 gnd.n1685 9.3005
R11009 gnd.n5813 gnd.n1686 9.3005
R11010 gnd.n5812 gnd.n1687 9.3005
R11011 gnd.n1727 gnd.n1688 9.3005
R11012 gnd.n5776 gnd.n5775 9.3005
R11013 gnd.n5780 gnd.n5779 9.3005
R11014 gnd.n5781 gnd.n1724 9.3005
R11015 gnd.n5790 gnd.n1725 9.3005
R11016 gnd.n5789 gnd.n5788 9.3005
R11017 gnd.n401 gnd.n400 9.3005
R11018 gnd.n7140 gnd.n7139 9.3005
R11019 gnd.n7141 gnd.n92 9.3005
R11020 gnd.n7329 gnd.n93 9.3005
R11021 gnd.n7328 gnd.n94 9.3005
R11022 gnd.n7327 gnd.n95 9.3005
R11023 gnd.n7156 gnd.n96 9.3005
R11024 gnd.n7317 gnd.n112 9.3005
R11025 gnd.n7316 gnd.n113 9.3005
R11026 gnd.n7315 gnd.n114 9.3005
R11027 gnd.n7171 gnd.n115 9.3005
R11028 gnd.n7305 gnd.n133 9.3005
R11029 gnd.n7304 gnd.n134 9.3005
R11030 gnd.n7303 gnd.n135 9.3005
R11031 gnd.n7270 gnd.n136 9.3005
R11032 gnd.n7293 gnd.n154 9.3005
R11033 gnd.n7292 gnd.n155 9.3005
R11034 gnd.n7291 gnd.n156 9.3005
R11035 gnd.n172 gnd.n157 9.3005
R11036 gnd.n7281 gnd.n7280 9.3005
R11037 gnd.n5663 gnd.n5662 9.3005
R11038 gnd.n5665 gnd.n5664 9.3005
R11039 gnd.n5666 gnd.n1625 9.3005
R11040 gnd.n5667 gnd.n1626 9.3005
R11041 gnd.n1746 gnd.n1627 9.3005
R11042 gnd.n5679 gnd.n1747 9.3005
R11043 gnd.n5680 gnd.n1645 9.3005
R11044 gnd.n5681 gnd.n1646 9.3005
R11045 gnd.n5682 gnd.n1647 9.3005
R11046 gnd.n5684 gnd.n5683 9.3005
R11047 gnd.n1734 gnd.n1666 9.3005
R11048 gnd.n5744 gnd.n1667 9.3005
R11049 gnd.n5745 gnd.n1668 9.3005
R11050 gnd.n5747 gnd.n5746 9.3005
R11051 gnd.n1728 gnd.n1685 9.3005
R11052 gnd.n5769 gnd.n1686 9.3005
R11053 gnd.n5770 gnd.n1687 9.3005
R11054 gnd.n5771 gnd.n1727 9.3005
R11055 gnd.n5775 gnd.n5774 9.3005
R11056 gnd.n5780 gnd.n1726 9.3005
R11057 gnd.n5782 gnd.n5781 9.3005
R11058 gnd.n5783 gnd.n1725 9.3005
R11059 gnd.n5788 gnd.n5787 9.3005
R11060 gnd.n5784 gnd.n400 9.3005
R11061 gnd.n7140 gnd.n399 9.3005
R11062 gnd.n7142 gnd.n7141 9.3005
R11063 gnd.n395 gnd.n93 9.3005
R11064 gnd.n7154 gnd.n94 9.3005
R11065 gnd.n7155 gnd.n95 9.3005
R11066 gnd.n7157 gnd.n7156 9.3005
R11067 gnd.n390 gnd.n112 9.3005
R11068 gnd.n7169 gnd.n113 9.3005
R11069 gnd.n7170 gnd.n114 9.3005
R11070 gnd.n7172 gnd.n7171 9.3005
R11071 gnd.n386 gnd.n133 9.3005
R11072 gnd.n7268 gnd.n134 9.3005
R11073 gnd.n7269 gnd.n135 9.3005
R11074 gnd.n7272 gnd.n7270 9.3005
R11075 gnd.n7273 gnd.n154 9.3005
R11076 gnd.n7275 gnd.n155 9.3005
R11077 gnd.n7276 gnd.n156 9.3005
R11078 gnd.n7278 gnd.n172 9.3005
R11079 gnd.n7280 gnd.n7279 9.3005
R11080 gnd.n5663 gnd.n1751 9.3005
R11081 gnd.n1757 gnd.n1754 9.3005
R11082 gnd.n5650 gnd.n1758 9.3005
R11083 gnd.n5652 gnd.n5651 9.3005
R11084 gnd.n5649 gnd.n1760 9.3005
R11085 gnd.n5648 gnd.n5647 9.3005
R11086 gnd.n1762 gnd.n1761 9.3005
R11087 gnd.n5641 gnd.n5640 9.3005
R11088 gnd.n5639 gnd.n1764 9.3005
R11089 gnd.n5638 gnd.n5637 9.3005
R11090 gnd.n1766 gnd.n1765 9.3005
R11091 gnd.n5631 gnd.n5630 9.3005
R11092 gnd.n5629 gnd.n1768 9.3005
R11093 gnd.n5628 gnd.n5627 9.3005
R11094 gnd.n1770 gnd.n1769 9.3005
R11095 gnd.n5621 gnd.n5620 9.3005
R11096 gnd.n5619 gnd.n1772 9.3005
R11097 gnd.n5618 gnd.n5617 9.3005
R11098 gnd.n1774 gnd.n1773 9.3005
R11099 gnd.n5611 gnd.n5610 9.3005
R11100 gnd.n5609 gnd.n1776 9.3005
R11101 gnd.n1778 gnd.n1777 9.3005
R11102 gnd.n5599 gnd.n5598 9.3005
R11103 gnd.n5597 gnd.n1780 9.3005
R11104 gnd.n5596 gnd.n5595 9.3005
R11105 gnd.n1782 gnd.n1781 9.3005
R11106 gnd.n5589 gnd.n5588 9.3005
R11107 gnd.n5587 gnd.n1784 9.3005
R11108 gnd.n5586 gnd.n5585 9.3005
R11109 gnd.n1786 gnd.n1785 9.3005
R11110 gnd.n5577 gnd.n5576 9.3005
R11111 gnd.n5574 gnd.n5487 9.3005
R11112 gnd.n5573 gnd.n5572 9.3005
R11113 gnd.n5489 gnd.n5488 9.3005
R11114 gnd.n5566 gnd.n5565 9.3005
R11115 gnd.n5564 gnd.n5491 9.3005
R11116 gnd.n5563 gnd.n5562 9.3005
R11117 gnd.n5493 gnd.n5492 9.3005
R11118 gnd.n5556 gnd.n5552 9.3005
R11119 gnd.n5551 gnd.n5495 9.3005
R11120 gnd.n5550 gnd.n5549 9.3005
R11121 gnd.n5497 gnd.n5496 9.3005
R11122 gnd.n5543 gnd.n5542 9.3005
R11123 gnd.n5541 gnd.n5499 9.3005
R11124 gnd.n5540 gnd.n5539 9.3005
R11125 gnd.n5501 gnd.n5500 9.3005
R11126 gnd.n5533 gnd.n5532 9.3005
R11127 gnd.n5531 gnd.n5503 9.3005
R11128 gnd.n5530 gnd.n5529 9.3005
R11129 gnd.n5505 gnd.n5504 9.3005
R11130 gnd.n5523 gnd.n5522 9.3005
R11131 gnd.n5521 gnd.n5507 9.3005
R11132 gnd.n5520 gnd.n5519 9.3005
R11133 gnd.n5509 gnd.n5508 9.3005
R11134 gnd.n5513 gnd.n5512 9.3005
R11135 gnd.n5511 gnd.n5510 9.3005
R11136 gnd.n5608 gnd.n5607 9.3005
R11137 gnd.n5660 gnd.n5659 9.3005
R11138 gnd.n5855 gnd.n1614 9.3005
R11139 gnd.n5854 gnd.n1615 9.3005
R11140 gnd.n1635 gnd.n1616 9.3005
R11141 gnd.n5844 gnd.n1636 9.3005
R11142 gnd.n5843 gnd.n1637 9.3005
R11143 gnd.n5842 gnd.n1638 9.3005
R11144 gnd.n1655 gnd.n1639 9.3005
R11145 gnd.n5832 gnd.n1656 9.3005
R11146 gnd.n5831 gnd.n1657 9.3005
R11147 gnd.n5830 gnd.n1658 9.3005
R11148 gnd.n1675 gnd.n1659 9.3005
R11149 gnd.n5820 gnd.n1676 9.3005
R11150 gnd.n5819 gnd.n1677 9.3005
R11151 gnd.n5818 gnd.n1678 9.3005
R11152 gnd.n1679 gnd.n78 9.3005
R11153 gnd.n83 gnd.n77 9.3005
R11154 gnd.n7323 gnd.n103 9.3005
R11155 gnd.n7322 gnd.n104 9.3005
R11156 gnd.n7321 gnd.n105 9.3005
R11157 gnd.n122 gnd.n106 9.3005
R11158 gnd.n7311 gnd.n123 9.3005
R11159 gnd.n7310 gnd.n124 9.3005
R11160 gnd.n7309 gnd.n125 9.3005
R11161 gnd.n143 gnd.n126 9.3005
R11162 gnd.n7299 gnd.n144 9.3005
R11163 gnd.n7298 gnd.n145 9.3005
R11164 gnd.n7297 gnd.n146 9.3005
R11165 gnd.n162 gnd.n147 9.3005
R11166 gnd.n7287 gnd.n163 9.3005
R11167 gnd.n7286 gnd.n164 9.3005
R11168 gnd.n7285 gnd.n165 9.3005
R11169 gnd.n5856 gnd.n1613 9.3005
R11170 gnd.n7334 gnd.n7333 9.3005
R11171 gnd.n4339 gnd.n2359 9.3005
R11172 gnd.n4360 gnd.n4340 9.3005
R11173 gnd.n4359 gnd.n4341 9.3005
R11174 gnd.n4358 gnd.n4342 9.3005
R11175 gnd.n4345 gnd.n4343 9.3005
R11176 gnd.n4354 gnd.n4346 9.3005
R11177 gnd.n4353 gnd.n4347 9.3005
R11178 gnd.n4352 gnd.n4348 9.3005
R11179 gnd.n4350 gnd.n4349 9.3005
R11180 gnd.n2337 gnd.n2336 9.3005
R11181 gnd.n4414 gnd.n4413 9.3005
R11182 gnd.n4415 gnd.n2335 9.3005
R11183 gnd.n4417 gnd.n4416 9.3005
R11184 gnd.n2333 gnd.n2332 9.3005
R11185 gnd.n4422 gnd.n4421 9.3005
R11186 gnd.n4423 gnd.n2331 9.3005
R11187 gnd.n4425 gnd.n4424 9.3005
R11188 gnd.n2329 gnd.n2328 9.3005
R11189 gnd.n4430 gnd.n4429 9.3005
R11190 gnd.n4431 gnd.n2327 9.3005
R11191 gnd.n4433 gnd.n4432 9.3005
R11192 gnd.n2324 gnd.n2323 9.3005
R11193 gnd.n4440 gnd.n4439 9.3005
R11194 gnd.n4441 gnd.n2322 9.3005
R11195 gnd.n4445 gnd.n4442 9.3005
R11196 gnd.n4444 gnd.n4443 9.3005
R11197 gnd.n2296 gnd.n2295 9.3005
R11198 gnd.n4472 gnd.n4471 9.3005
R11199 gnd.n4473 gnd.n2294 9.3005
R11200 gnd.n4478 gnd.n4474 9.3005
R11201 gnd.n4477 gnd.n4476 9.3005
R11202 gnd.n4475 gnd.n1484 9.3005
R11203 gnd.n5989 gnd.n1485 9.3005
R11204 gnd.n5988 gnd.n1486 9.3005
R11205 gnd.n5987 gnd.n1487 9.3005
R11206 gnd.n4512 gnd.n1488 9.3005
R11207 gnd.n4514 gnd.n4513 9.3005
R11208 gnd.n2170 gnd.n2169 9.3005
R11209 gnd.n4554 gnd.n4553 9.3005
R11210 gnd.n4555 gnd.n2168 9.3005
R11211 gnd.n4557 gnd.n4556 9.3005
R11212 gnd.n2152 gnd.n2151 9.3005
R11213 gnd.n4596 gnd.n4595 9.3005
R11214 gnd.n4597 gnd.n2150 9.3005
R11215 gnd.n4601 gnd.n4598 9.3005
R11216 gnd.n4600 gnd.n4599 9.3005
R11217 gnd.n2126 gnd.n2125 9.3005
R11218 gnd.n4658 gnd.n4657 9.3005
R11219 gnd.n4659 gnd.n2124 9.3005
R11220 gnd.n4661 gnd.n4660 9.3005
R11221 gnd.n2108 gnd.n2107 9.3005
R11222 gnd.n4686 gnd.n4685 9.3005
R11223 gnd.n4687 gnd.n2106 9.3005
R11224 gnd.n4691 gnd.n4688 9.3005
R11225 gnd.n4690 gnd.n4689 9.3005
R11226 gnd.n2075 gnd.n2074 9.3005
R11227 gnd.n4736 gnd.n4735 9.3005
R11228 gnd.n4737 gnd.n2073 9.3005
R11229 gnd.n4739 gnd.n4738 9.3005
R11230 gnd.n2052 gnd.n2051 9.3005
R11231 gnd.n4776 gnd.n4775 9.3005
R11232 gnd.n4777 gnd.n2050 9.3005
R11233 gnd.n4779 gnd.n4778 9.3005
R11234 gnd.n2030 gnd.n2029 9.3005
R11235 gnd.n4833 gnd.n4832 9.3005
R11236 gnd.n4834 gnd.n2028 9.3005
R11237 gnd.n4836 gnd.n4835 9.3005
R11238 gnd.n2010 gnd.n2009 9.3005
R11239 gnd.n4858 gnd.n4857 9.3005
R11240 gnd.n4859 gnd.n2008 9.3005
R11241 gnd.n4861 gnd.n4860 9.3005
R11242 gnd.n1990 gnd.n1989 9.3005
R11243 gnd.n4918 gnd.n4917 9.3005
R11244 gnd.n4919 gnd.n1988 9.3005
R11245 gnd.n4921 gnd.n4920 9.3005
R11246 gnd.n1968 gnd.n1967 9.3005
R11247 gnd.n4947 gnd.n4946 9.3005
R11248 gnd.n4948 gnd.n1966 9.3005
R11249 gnd.n4952 gnd.n4949 9.3005
R11250 gnd.n4951 gnd.n4950 9.3005
R11251 gnd.n1940 gnd.n1939 9.3005
R11252 gnd.n4998 gnd.n4997 9.3005
R11253 gnd.n4999 gnd.n1938 9.3005
R11254 gnd.n5001 gnd.n5000 9.3005
R11255 gnd.n1920 gnd.n1919 9.3005
R11256 gnd.n5024 gnd.n5023 9.3005
R11257 gnd.n5025 gnd.n1918 9.3005
R11258 gnd.n5029 gnd.n5026 9.3005
R11259 gnd.n5028 gnd.n5027 9.3005
R11260 gnd.n1890 gnd.n1889 9.3005
R11261 gnd.n5068 gnd.n5067 9.3005
R11262 gnd.n5069 gnd.n1888 9.3005
R11263 gnd.n5074 gnd.n5070 9.3005
R11264 gnd.n5073 gnd.n5072 9.3005
R11265 gnd.n5071 gnd.n1839 9.3005
R11266 gnd.n5320 gnd.n1840 9.3005
R11267 gnd.n5319 gnd.n1841 9.3005
R11268 gnd.n5318 gnd.n1842 9.3005
R11269 gnd.n1851 gnd.n1843 9.3005
R11270 gnd.n1852 gnd.n1850 9.3005
R11271 gnd.n5308 gnd.n1853 9.3005
R11272 gnd.n5307 gnd.n1854 9.3005
R11273 gnd.n5306 gnd.n1855 9.3005
R11274 gnd.n1858 gnd.n1857 9.3005
R11275 gnd.n1856 gnd.n1591 9.3005
R11276 gnd.n5871 gnd.n1592 9.3005
R11277 gnd.n5870 gnd.n1593 9.3005
R11278 gnd.n5869 gnd.n1594 9.3005
R11279 gnd.n1600 gnd.n1595 9.3005
R11280 gnd.n5863 gnd.n1601 9.3005
R11281 gnd.n5862 gnd.n1602 9.3005
R11282 gnd.n5861 gnd.n1603 9.3005
R11283 gnd.n5705 gnd.n1604 9.3005
R11284 gnd.n5708 gnd.n5707 9.3005
R11285 gnd.n5709 gnd.n5704 9.3005
R11286 gnd.n5711 gnd.n5710 9.3005
R11287 gnd.n5702 gnd.n5701 9.3005
R11288 gnd.n5716 gnd.n5715 9.3005
R11289 gnd.n5717 gnd.n5700 9.3005
R11290 gnd.n5719 gnd.n5718 9.3005
R11291 gnd.n1740 gnd.n1739 9.3005
R11292 gnd.n5724 gnd.n5723 9.3005
R11293 gnd.n5725 gnd.n1738 9.3005
R11294 gnd.n5739 gnd.n5726 9.3005
R11295 gnd.n5738 gnd.n5727 9.3005
R11296 gnd.n5737 gnd.n5728 9.3005
R11297 gnd.n5730 gnd.n5729 9.3005
R11298 gnd.n5733 gnd.n5731 9.3005
R11299 gnd.n7131 gnd.n405 9.3005
R11300 gnd.n408 gnd.n406 9.3005
R11301 gnd.n7127 gnd.n409 9.3005
R11302 gnd.n7126 gnd.n410 9.3005
R11303 gnd.n7125 gnd.n411 9.3005
R11304 gnd.n414 gnd.n412 9.3005
R11305 gnd.n7121 gnd.n415 9.3005
R11306 gnd.n7120 gnd.n416 9.3005
R11307 gnd.n7119 gnd.n417 9.3005
R11308 gnd.n7113 gnd.n418 9.3005
R11309 gnd.n4294 gnd.n4293 9.3005
R11310 gnd.n4048 gnd.n4034 9.3005
R11311 gnd.n4047 gnd.n4035 9.3005
R11312 gnd.n4045 gnd.n4036 9.3005
R11313 gnd.n4044 gnd.n4037 9.3005
R11314 gnd.n4042 gnd.n4038 9.3005
R11315 gnd.n4041 gnd.n4039 9.3005
R11316 gnd.n2418 gnd.n2417 9.3005
R11317 gnd.n4255 gnd.n4254 9.3005
R11318 gnd.n4256 gnd.n2416 9.3005
R11319 gnd.n4258 gnd.n4257 9.3005
R11320 gnd.n2395 gnd.n2394 9.3005
R11321 gnd.n4270 gnd.n4269 9.3005
R11322 gnd.n4271 gnd.n2393 9.3005
R11323 gnd.n4276 gnd.n4272 9.3005
R11324 gnd.n4275 gnd.n4274 9.3005
R11325 gnd.n4273 gnd.n2373 9.3005
R11326 gnd.n4330 gnd.n2374 9.3005
R11327 gnd.n4329 gnd.n2375 9.3005
R11328 gnd.n4328 gnd.n2376 9.3005
R11329 gnd.n4292 gnd.n2377 9.3005
R11330 gnd.n4051 gnd.n4050 9.3005
R11331 gnd.n4056 gnd.n4055 9.3005
R11332 gnd.n4059 gnd.n4029 9.3005
R11333 gnd.n4060 gnd.n4028 9.3005
R11334 gnd.n4063 gnd.n4027 9.3005
R11335 gnd.n4064 gnd.n4026 9.3005
R11336 gnd.n4067 gnd.n4025 9.3005
R11337 gnd.n4068 gnd.n4024 9.3005
R11338 gnd.n4071 gnd.n4023 9.3005
R11339 gnd.n4072 gnd.n4022 9.3005
R11340 gnd.n4075 gnd.n4021 9.3005
R11341 gnd.n4076 gnd.n4020 9.3005
R11342 gnd.n4079 gnd.n4019 9.3005
R11343 gnd.n4080 gnd.n4018 9.3005
R11344 gnd.n4083 gnd.n4017 9.3005
R11345 gnd.n4084 gnd.n4016 9.3005
R11346 gnd.n4087 gnd.n4015 9.3005
R11347 gnd.n4088 gnd.n4014 9.3005
R11348 gnd.n4054 gnd.n4033 9.3005
R11349 gnd.n4053 gnd.n4052 9.3005
R11350 gnd.n6067 gnd.n1317 9.3005
R11351 gnd.n6070 gnd.n1316 9.3005
R11352 gnd.n6071 gnd.n1315 9.3005
R11353 gnd.n6074 gnd.n1314 9.3005
R11354 gnd.n6075 gnd.n1313 9.3005
R11355 gnd.n6078 gnd.n1312 9.3005
R11356 gnd.n6079 gnd.n1311 9.3005
R11357 gnd.n6082 gnd.n1310 9.3005
R11358 gnd.n6084 gnd.n1307 9.3005
R11359 gnd.n6087 gnd.n1306 9.3005
R11360 gnd.n6088 gnd.n1305 9.3005
R11361 gnd.n6091 gnd.n1304 9.3005
R11362 gnd.n6092 gnd.n1303 9.3005
R11363 gnd.n6095 gnd.n1302 9.3005
R11364 gnd.n6096 gnd.n1301 9.3005
R11365 gnd.n6099 gnd.n1300 9.3005
R11366 gnd.n6100 gnd.n1299 9.3005
R11367 gnd.n6103 gnd.n1298 9.3005
R11368 gnd.n6104 gnd.n1297 9.3005
R11369 gnd.n6107 gnd.n1296 9.3005
R11370 gnd.n6108 gnd.n1295 9.3005
R11371 gnd.n6111 gnd.n1294 9.3005
R11372 gnd.n6112 gnd.n1293 9.3005
R11373 gnd.n6113 gnd.n1292 9.3005
R11374 gnd.n1291 gnd.n1288 9.3005
R11375 gnd.n1290 gnd.n1289 9.3005
R11376 gnd.n1414 gnd.n1413 9.3005
R11377 gnd.n1410 gnd.n1320 9.3005
R11378 gnd.n1407 gnd.n1321 9.3005
R11379 gnd.n1406 gnd.n1322 9.3005
R11380 gnd.n1403 gnd.n1323 9.3005
R11381 gnd.n1402 gnd.n1324 9.3005
R11382 gnd.n1399 gnd.n1325 9.3005
R11383 gnd.n1398 gnd.n1326 9.3005
R11384 gnd.n1395 gnd.n1394 9.3005
R11385 gnd.n1393 gnd.n1327 9.3005
R11386 gnd.n1392 gnd.n1391 9.3005
R11387 gnd.n1388 gnd.n1330 9.3005
R11388 gnd.n1385 gnd.n1331 9.3005
R11389 gnd.n1384 gnd.n1332 9.3005
R11390 gnd.n1381 gnd.n1333 9.3005
R11391 gnd.n1380 gnd.n1334 9.3005
R11392 gnd.n1377 gnd.n1335 9.3005
R11393 gnd.n1376 gnd.n1336 9.3005
R11394 gnd.n1373 gnd.n1337 9.3005
R11395 gnd.n1372 gnd.n1338 9.3005
R11396 gnd.n1369 gnd.n1339 9.3005
R11397 gnd.n1368 gnd.n1340 9.3005
R11398 gnd.n1365 gnd.n1341 9.3005
R11399 gnd.n1364 gnd.n1342 9.3005
R11400 gnd.n1361 gnd.n1343 9.3005
R11401 gnd.n1360 gnd.n1344 9.3005
R11402 gnd.n1357 gnd.n1345 9.3005
R11403 gnd.n1356 gnd.n1346 9.3005
R11404 gnd.n1353 gnd.n1352 9.3005
R11405 gnd.n1351 gnd.n1348 9.3005
R11406 gnd.n1415 gnd.n1318 9.3005
R11407 gnd.n4093 gnd.n4092 9.3005
R11408 gnd.n2440 gnd.n2436 9.3005
R11409 gnd.n4232 gnd.n2437 9.3005
R11410 gnd.n4231 gnd.n4230 9.3005
R11411 gnd.n2438 gnd.n2421 9.3005
R11412 gnd.n4246 gnd.n2420 9.3005
R11413 gnd.n4248 gnd.n4247 9.3005
R11414 gnd.n4249 gnd.n985 9.3005
R11415 gnd.n6297 gnd.n986 9.3005
R11416 gnd.n6296 gnd.n987 9.3005
R11417 gnd.n6295 gnd.n988 9.3005
R11418 gnd.n4264 gnd.n989 9.3005
R11419 gnd.n6285 gnd.n1007 9.3005
R11420 gnd.n6284 gnd.n1008 9.3005
R11421 gnd.n6283 gnd.n1009 9.3005
R11422 gnd.n4285 gnd.n1010 9.3005
R11423 gnd.n4286 gnd.n1028 9.3005
R11424 gnd.n6271 gnd.n1029 9.3005
R11425 gnd.n6270 gnd.n1030 9.3005
R11426 gnd.n6269 gnd.n1031 9.3005
R11427 gnd.n4291 gnd.n1032 9.3005
R11428 gnd.n6258 gnd.n1045 9.3005
R11429 gnd.n6257 gnd.n1046 9.3005
R11430 gnd.n6256 gnd.n1047 9.3005
R11431 gnd.n4302 gnd.n1048 9.3005
R11432 gnd.n6245 gnd.n1063 9.3005
R11433 gnd.n6244 gnd.n1064 9.3005
R11434 gnd.n6243 gnd.n1065 9.3005
R11435 gnd.n2352 gnd.n1066 9.3005
R11436 gnd.n6233 gnd.n1082 9.3005
R11437 gnd.n6232 gnd.n1083 9.3005
R11438 gnd.n6231 gnd.n1084 9.3005
R11439 gnd.n2346 gnd.n1085 9.3005
R11440 gnd.n6221 gnd.n1103 9.3005
R11441 gnd.n6220 gnd.n1104 9.3005
R11442 gnd.n6219 gnd.n1105 9.3005
R11443 gnd.n4391 gnd.n1106 9.3005
R11444 gnd.n6209 gnd.n1123 9.3005
R11445 gnd.n6208 gnd.n1124 9.3005
R11446 gnd.n6207 gnd.n1125 9.3005
R11447 gnd.n1143 gnd.n1126 9.3005
R11448 gnd.n6197 gnd.n6196 9.3005
R11449 gnd.n4095 gnd.n4091 9.3005
R11450 gnd.n4093 gnd.n2439 9.3005
R11451 gnd.n4223 gnd.n2440 9.3005
R11452 gnd.n4224 gnd.n2437 9.3005
R11453 gnd.n4230 gnd.n4229 9.3005
R11454 gnd.n4227 gnd.n2438 9.3005
R11455 gnd.n4226 gnd.n2420 9.3005
R11456 gnd.n4248 gnd.n2419 9.3005
R11457 gnd.n4250 gnd.n4249 9.3005
R11458 gnd.n2396 gnd.n986 9.3005
R11459 gnd.n4262 gnd.n987 9.3005
R11460 gnd.n4263 gnd.n988 9.3005
R11461 gnd.n4265 gnd.n4264 9.3005
R11462 gnd.n2392 gnd.n1007 9.3005
R11463 gnd.n4281 gnd.n1008 9.3005
R11464 gnd.n4282 gnd.n1009 9.3005
R11465 gnd.n4285 gnd.n4284 9.3005
R11466 gnd.n4287 gnd.n4286 9.3005
R11467 gnd.n4288 gnd.n1029 9.3005
R11468 gnd.n4289 gnd.n1030 9.3005
R11469 gnd.n4290 gnd.n1031 9.3005
R11470 gnd.n4298 gnd.n4291 9.3005
R11471 gnd.n4299 gnd.n1045 9.3005
R11472 gnd.n4300 gnd.n1046 9.3005
R11473 gnd.n4301 gnd.n1047 9.3005
R11474 gnd.n4305 gnd.n4302 9.3005
R11475 gnd.n4304 gnd.n1063 9.3005
R11476 gnd.n4303 gnd.n1064 9.3005
R11477 gnd.n2351 gnd.n1065 9.3005
R11478 gnd.n4373 gnd.n2352 9.3005
R11479 gnd.n4374 gnd.n1082 9.3005
R11480 gnd.n4375 gnd.n1083 9.3005
R11481 gnd.n2345 gnd.n1084 9.3005
R11482 gnd.n4387 gnd.n2346 9.3005
R11483 gnd.n4388 gnd.n1103 9.3005
R11484 gnd.n4389 gnd.n1104 9.3005
R11485 gnd.n4390 gnd.n1105 9.3005
R11486 gnd.n4394 gnd.n4391 9.3005
R11487 gnd.n4395 gnd.n1123 9.3005
R11488 gnd.n4396 gnd.n1124 9.3005
R11489 gnd.n1145 gnd.n1125 9.3005
R11490 gnd.n6194 gnd.n1143 9.3005
R11491 gnd.n6196 gnd.n6195 9.3005
R11492 gnd.n4095 gnd.n4094 9.3005
R11493 gnd.n4099 gnd.n4098 9.3005
R11494 gnd.n4102 gnd.n4009 9.3005
R11495 gnd.n4103 gnd.n4008 9.3005
R11496 gnd.n4106 gnd.n4007 9.3005
R11497 gnd.n4107 gnd.n4006 9.3005
R11498 gnd.n4110 gnd.n4005 9.3005
R11499 gnd.n4111 gnd.n4004 9.3005
R11500 gnd.n4114 gnd.n4003 9.3005
R11501 gnd.n4115 gnd.n4002 9.3005
R11502 gnd.n4118 gnd.n4001 9.3005
R11503 gnd.n4119 gnd.n4000 9.3005
R11504 gnd.n4122 gnd.n3999 9.3005
R11505 gnd.n4123 gnd.n3998 9.3005
R11506 gnd.n4126 gnd.n3997 9.3005
R11507 gnd.n4127 gnd.n3996 9.3005
R11508 gnd.n4130 gnd.n3995 9.3005
R11509 gnd.n4131 gnd.n3994 9.3005
R11510 gnd.n4134 gnd.n3993 9.3005
R11511 gnd.n4135 gnd.n3992 9.3005
R11512 gnd.n4138 gnd.n3991 9.3005
R11513 gnd.n4142 gnd.n3987 9.3005
R11514 gnd.n4143 gnd.n3986 9.3005
R11515 gnd.n4146 gnd.n3985 9.3005
R11516 gnd.n4147 gnd.n3984 9.3005
R11517 gnd.n4150 gnd.n3983 9.3005
R11518 gnd.n4151 gnd.n3982 9.3005
R11519 gnd.n4154 gnd.n3981 9.3005
R11520 gnd.n4155 gnd.n3980 9.3005
R11521 gnd.n4158 gnd.n3979 9.3005
R11522 gnd.n4159 gnd.n3978 9.3005
R11523 gnd.n4162 gnd.n3977 9.3005
R11524 gnd.n4163 gnd.n3976 9.3005
R11525 gnd.n4166 gnd.n3975 9.3005
R11526 gnd.n4167 gnd.n3974 9.3005
R11527 gnd.n4170 gnd.n3973 9.3005
R11528 gnd.n4171 gnd.n3972 9.3005
R11529 gnd.n4174 gnd.n3971 9.3005
R11530 gnd.n4175 gnd.n3970 9.3005
R11531 gnd.n4178 gnd.n3969 9.3005
R11532 gnd.n4180 gnd.n3966 9.3005
R11533 gnd.n4183 gnd.n3965 9.3005
R11534 gnd.n4184 gnd.n3964 9.3005
R11535 gnd.n4187 gnd.n3963 9.3005
R11536 gnd.n4188 gnd.n3962 9.3005
R11537 gnd.n4191 gnd.n3961 9.3005
R11538 gnd.n4192 gnd.n3960 9.3005
R11539 gnd.n4195 gnd.n3959 9.3005
R11540 gnd.n4196 gnd.n3958 9.3005
R11541 gnd.n4199 gnd.n3957 9.3005
R11542 gnd.n4200 gnd.n3956 9.3005
R11543 gnd.n4203 gnd.n3955 9.3005
R11544 gnd.n4204 gnd.n3954 9.3005
R11545 gnd.n4207 gnd.n3953 9.3005
R11546 gnd.n4208 gnd.n3952 9.3005
R11547 gnd.n4209 gnd.n3951 9.3005
R11548 gnd.n2448 gnd.n2447 9.3005
R11549 gnd.n4215 gnd.n4214 9.3005
R11550 gnd.n4139 gnd.n3988 9.3005
R11551 gnd.n4097 gnd.n4011 9.3005
R11552 gnd.n4218 gnd.n4217 9.3005
R11553 gnd.n2429 gnd.n2428 9.3005
R11554 gnd.n4237 gnd.n4236 9.3005
R11555 gnd.n4238 gnd.n2427 9.3005
R11556 gnd.n4241 gnd.n4240 9.3005
R11557 gnd.n4239 gnd.n974 9.3005
R11558 gnd.n6303 gnd.n975 9.3005
R11559 gnd.n6302 gnd.n976 9.3005
R11560 gnd.n6301 gnd.n977 9.3005
R11561 gnd.n996 gnd.n978 9.3005
R11562 gnd.n6291 gnd.n997 9.3005
R11563 gnd.n6290 gnd.n998 9.3005
R11564 gnd.n6289 gnd.n999 9.3005
R11565 gnd.n1016 gnd.n1000 9.3005
R11566 gnd.n6279 gnd.n1017 9.3005
R11567 gnd.n1072 gnd.n1056 9.3005
R11568 gnd.n6239 gnd.n1073 9.3005
R11569 gnd.n6238 gnd.n1074 9.3005
R11570 gnd.n6237 gnd.n1075 9.3005
R11571 gnd.n1092 gnd.n1076 9.3005
R11572 gnd.n6227 gnd.n1093 9.3005
R11573 gnd.n6226 gnd.n1094 9.3005
R11574 gnd.n6225 gnd.n1095 9.3005
R11575 gnd.n1112 gnd.n1096 9.3005
R11576 gnd.n6215 gnd.n1113 9.3005
R11577 gnd.n6214 gnd.n1114 9.3005
R11578 gnd.n6213 gnd.n1115 9.3005
R11579 gnd.n1133 gnd.n1116 9.3005
R11580 gnd.n6203 gnd.n1134 9.3005
R11581 gnd.n6202 gnd.n1135 9.3005
R11582 gnd.n6201 gnd.n1136 9.3005
R11583 gnd.n4216 gnd.n2446 9.3005
R11584 gnd.n6249 gnd.n1018 9.3005
R11585 gnd.n965 gnd.n964 9.3005
R11586 gnd.n2400 gnd.n2399 9.3005
R11587 gnd.n2413 gnd.n2401 9.3005
R11588 gnd.n2412 gnd.n2402 9.3005
R11589 gnd.n2411 gnd.n2403 9.3005
R11590 gnd.n2405 gnd.n2404 9.3005
R11591 gnd.n2407 gnd.n2406 9.3005
R11592 gnd.n2366 gnd.n2365 9.3005
R11593 gnd.n4337 gnd.n4336 9.3005
R11594 gnd.n6309 gnd.n6308 9.3005
R11595 gnd.n6312 gnd.n963 9.3005
R11596 gnd.n962 gnd.n958 9.3005
R11597 gnd.n6318 gnd.n957 9.3005
R11598 gnd.n6319 gnd.n956 9.3005
R11599 gnd.n6320 gnd.n955 9.3005
R11600 gnd.n954 gnd.n950 9.3005
R11601 gnd.n6326 gnd.n949 9.3005
R11602 gnd.n6327 gnd.n948 9.3005
R11603 gnd.n6328 gnd.n947 9.3005
R11604 gnd.n946 gnd.n942 9.3005
R11605 gnd.n6334 gnd.n941 9.3005
R11606 gnd.n6335 gnd.n940 9.3005
R11607 gnd.n6336 gnd.n939 9.3005
R11608 gnd.n938 gnd.n934 9.3005
R11609 gnd.n6342 gnd.n933 9.3005
R11610 gnd.n6343 gnd.n932 9.3005
R11611 gnd.n6344 gnd.n931 9.3005
R11612 gnd.n930 gnd.n926 9.3005
R11613 gnd.n6350 gnd.n925 9.3005
R11614 gnd.n6351 gnd.n924 9.3005
R11615 gnd.n6352 gnd.n923 9.3005
R11616 gnd.n922 gnd.n918 9.3005
R11617 gnd.n6358 gnd.n917 9.3005
R11618 gnd.n6359 gnd.n916 9.3005
R11619 gnd.n6360 gnd.n915 9.3005
R11620 gnd.n914 gnd.n910 9.3005
R11621 gnd.n6366 gnd.n909 9.3005
R11622 gnd.n6367 gnd.n908 9.3005
R11623 gnd.n6368 gnd.n907 9.3005
R11624 gnd.n906 gnd.n902 9.3005
R11625 gnd.n6374 gnd.n901 9.3005
R11626 gnd.n6375 gnd.n900 9.3005
R11627 gnd.n6376 gnd.n899 9.3005
R11628 gnd.n898 gnd.n894 9.3005
R11629 gnd.n6382 gnd.n893 9.3005
R11630 gnd.n6383 gnd.n892 9.3005
R11631 gnd.n6384 gnd.n891 9.3005
R11632 gnd.n890 gnd.n886 9.3005
R11633 gnd.n6390 gnd.n885 9.3005
R11634 gnd.n6391 gnd.n884 9.3005
R11635 gnd.n6392 gnd.n883 9.3005
R11636 gnd.n882 gnd.n878 9.3005
R11637 gnd.n6398 gnd.n877 9.3005
R11638 gnd.n6399 gnd.n876 9.3005
R11639 gnd.n6400 gnd.n875 9.3005
R11640 gnd.n874 gnd.n870 9.3005
R11641 gnd.n6406 gnd.n869 9.3005
R11642 gnd.n6407 gnd.n868 9.3005
R11643 gnd.n6408 gnd.n867 9.3005
R11644 gnd.n866 gnd.n862 9.3005
R11645 gnd.n6414 gnd.n861 9.3005
R11646 gnd.n6415 gnd.n860 9.3005
R11647 gnd.n6416 gnd.n859 9.3005
R11648 gnd.n858 gnd.n854 9.3005
R11649 gnd.n6422 gnd.n853 9.3005
R11650 gnd.n6423 gnd.n852 9.3005
R11651 gnd.n6424 gnd.n851 9.3005
R11652 gnd.n850 gnd.n846 9.3005
R11653 gnd.n6430 gnd.n845 9.3005
R11654 gnd.n6431 gnd.n844 9.3005
R11655 gnd.n6432 gnd.n843 9.3005
R11656 gnd.n842 gnd.n838 9.3005
R11657 gnd.n6438 gnd.n837 9.3005
R11658 gnd.n6439 gnd.n836 9.3005
R11659 gnd.n6440 gnd.n835 9.3005
R11660 gnd.n834 gnd.n830 9.3005
R11661 gnd.n6446 gnd.n829 9.3005
R11662 gnd.n6447 gnd.n828 9.3005
R11663 gnd.n6448 gnd.n827 9.3005
R11664 gnd.n826 gnd.n822 9.3005
R11665 gnd.n6454 gnd.n821 9.3005
R11666 gnd.n6455 gnd.n820 9.3005
R11667 gnd.n6456 gnd.n819 9.3005
R11668 gnd.n818 gnd.n814 9.3005
R11669 gnd.n6462 gnd.n813 9.3005
R11670 gnd.n6463 gnd.n812 9.3005
R11671 gnd.n6464 gnd.n811 9.3005
R11672 gnd.n810 gnd.n806 9.3005
R11673 gnd.n6470 gnd.n805 9.3005
R11674 gnd.n6471 gnd.n804 9.3005
R11675 gnd.n6472 gnd.n803 9.3005
R11676 gnd.n802 gnd.n798 9.3005
R11677 gnd.n6478 gnd.n797 9.3005
R11678 gnd.n6480 gnd.n6479 9.3005
R11679 gnd.n6311 gnd.n6310 9.3005
R11680 gnd.n5296 gnd.n5295 9.3005
R11681 gnd.n2317 gnd.n2316 9.3005
R11682 gnd.n2303 gnd.n2302 9.3005
R11683 gnd.n4460 gnd.n4459 9.3005
R11684 gnd.n4461 gnd.n2300 9.3005
R11685 gnd.n4466 gnd.n4465 9.3005
R11686 gnd.n4464 gnd.n2301 9.3005
R11687 gnd.n4463 gnd.n4462 9.3005
R11688 gnd.n2202 gnd.n2201 9.3005
R11689 gnd.n4497 gnd.n4496 9.3005
R11690 gnd.n4498 gnd.n2199 9.3005
R11691 gnd.n4501 gnd.n4500 9.3005
R11692 gnd.n4499 gnd.n2200 9.3005
R11693 gnd.n2191 gnd.n2190 9.3005
R11694 gnd.n4522 gnd.n4521 9.3005
R11695 gnd.n4523 gnd.n2188 9.3005
R11696 gnd.n4532 gnd.n4531 9.3005
R11697 gnd.n4530 gnd.n2189 9.3005
R11698 gnd.n4529 gnd.n4528 9.3005
R11699 gnd.n4527 gnd.n4524 9.3005
R11700 gnd.n2144 gnd.n2143 9.3005
R11701 gnd.n4608 gnd.n4607 9.3005
R11702 gnd.n4609 gnd.n2141 9.3005
R11703 gnd.n4630 gnd.n4629 9.3005
R11704 gnd.n4628 gnd.n2142 9.3005
R11705 gnd.n4627 gnd.n4626 9.3005
R11706 gnd.n4625 gnd.n4610 9.3005
R11707 gnd.n4624 gnd.n4623 9.3005
R11708 gnd.n4622 gnd.n4616 9.3005
R11709 gnd.n4621 gnd.n4620 9.3005
R11710 gnd.n4619 gnd.n4618 9.3005
R11711 gnd.n4617 gnd.n2094 9.3005
R11712 gnd.n2092 gnd.n2091 9.3005
R11713 gnd.n4710 gnd.n4709 9.3005
R11714 gnd.n4711 gnd.n2090 9.3005
R11715 gnd.n4713 gnd.n4712 9.3005
R11716 gnd.n2067 gnd.n2065 9.3005
R11717 gnd.n4759 gnd.n4758 9.3005
R11718 gnd.n4757 gnd.n2066 9.3005
R11719 gnd.n4756 gnd.n4755 9.3005
R11720 gnd.n2044 gnd.n2042 9.3005
R11721 gnd.n4818 gnd.n4817 9.3005
R11722 gnd.n4816 gnd.n2043 9.3005
R11723 gnd.n4815 gnd.n4814 9.3005
R11724 gnd.n4813 gnd.n2045 9.3005
R11725 gnd.n4812 gnd.n4811 9.3005
R11726 gnd.n4810 gnd.n4798 9.3005
R11727 gnd.n4809 gnd.n4808 9.3005
R11728 gnd.n4807 gnd.n4799 9.3005
R11729 gnd.n4806 gnd.n4805 9.3005
R11730 gnd.n1983 gnd.n1982 9.3005
R11731 gnd.n4927 gnd.n4926 9.3005
R11732 gnd.n4928 gnd.n1980 9.3005
R11733 gnd.n4931 gnd.n4930 9.3005
R11734 gnd.n4929 gnd.n1981 9.3005
R11735 gnd.n1954 gnd.n1953 9.3005
R11736 gnd.n4966 gnd.n4965 9.3005
R11737 gnd.n4967 gnd.n1951 9.3005
R11738 gnd.n4984 gnd.n4983 9.3005
R11739 gnd.n4982 gnd.n1952 9.3005
R11740 gnd.n4981 gnd.n4980 9.3005
R11741 gnd.n4979 gnd.n4968 9.3005
R11742 gnd.n4978 gnd.n4977 9.3005
R11743 gnd.n4976 gnd.n4973 9.3005
R11744 gnd.n4975 gnd.n4974 9.3005
R11745 gnd.n1898 gnd.n1897 9.3005
R11746 gnd.n5057 gnd.n5056 9.3005
R11747 gnd.n5058 gnd.n1895 9.3005
R11748 gnd.n5061 gnd.n5060 9.3005
R11749 gnd.n5059 gnd.n1896 9.3005
R11750 gnd.n1871 gnd.n1870 9.3005
R11751 gnd.n5099 gnd.n5098 9.3005
R11752 gnd.n5100 gnd.n1869 9.3005
R11753 gnd.n5102 gnd.n5101 9.3005
R11754 gnd.n1868 gnd.n1867 9.3005
R11755 gnd.n5110 gnd.n5109 9.3005
R11756 gnd.n5111 gnd.n1866 9.3005
R11757 gnd.n5113 gnd.n5112 9.3005
R11758 gnd.n5114 gnd.n1865 9.3005
R11759 gnd.n5118 gnd.n5117 9.3005
R11760 gnd.n5119 gnd.n1863 9.3005
R11761 gnd.n5299 gnd.n5298 9.3005
R11762 gnd.n5297 gnd.n1864 9.3005
R11763 gnd.n2315 gnd.n2314 9.3005
R11764 gnd.n6184 gnd.n1149 9.3005
R11765 gnd.n2391 gnd.n2389 9.3005
R11766 gnd.n4313 gnd.n4312 9.3005
R11767 gnd.n4311 gnd.n2390 9.3005
R11768 gnd.n4310 gnd.n4309 9.3005
R11769 gnd.n2355 gnd.n2354 9.3005
R11770 gnd.n4366 gnd.n4365 9.3005
R11771 gnd.n4367 gnd.n2353 9.3005
R11772 gnd.n4369 gnd.n4368 9.3005
R11773 gnd.n2349 gnd.n2348 9.3005
R11774 gnd.n4380 gnd.n4379 9.3005
R11775 gnd.n4381 gnd.n2347 9.3005
R11776 gnd.n4383 gnd.n4382 9.3005
R11777 gnd.n2342 gnd.n2340 9.3005
R11778 gnd.n4407 gnd.n4406 9.3005
R11779 gnd.n4405 gnd.n2341 9.3005
R11780 gnd.n4404 gnd.n4403 9.3005
R11781 gnd.n4402 gnd.n2343 9.3005
R11782 gnd.n4401 gnd.n4400 9.3005
R11783 gnd.n1148 gnd.n1146 9.3005
R11784 gnd.n6190 gnd.n6189 9.3005
R11785 gnd.n6188 gnd.n1147 9.3005
R11786 gnd.n6162 gnd.n6161 9.3005
R11787 gnd.n6160 gnd.n6159 9.3005
R11788 gnd.n1191 gnd.n1190 9.3005
R11789 gnd.n6154 gnd.n6153 9.3005
R11790 gnd.n6152 gnd.n6151 9.3005
R11791 gnd.n1201 gnd.n1200 9.3005
R11792 gnd.n6146 gnd.n6145 9.3005
R11793 gnd.n6144 gnd.n6143 9.3005
R11794 gnd.n1209 gnd.n1208 9.3005
R11795 gnd.n6138 gnd.n6137 9.3005
R11796 gnd.n6136 gnd.n6135 9.3005
R11797 gnd.n1219 gnd.n1218 9.3005
R11798 gnd.n6130 gnd.n6129 9.3005
R11799 gnd.n6128 gnd.n6127 9.3005
R11800 gnd.n1227 gnd.n1226 9.3005
R11801 gnd.n6122 gnd.n6121 9.3005
R11802 gnd.n6120 gnd.n1241 9.3005
R11803 gnd.n6119 gnd.n1150 9.3005
R11804 gnd.n1187 gnd.n1185 9.3005
R11805 gnd.n6186 gnd.n6185 9.3005
R11806 gnd.n1240 gnd.n1151 9.3005
R11807 gnd.n1236 gnd.n1235 9.3005
R11808 gnd.n6124 gnd.n6123 9.3005
R11809 gnd.n6126 gnd.n6125 9.3005
R11810 gnd.n1223 gnd.n1222 9.3005
R11811 gnd.n6132 gnd.n6131 9.3005
R11812 gnd.n6134 gnd.n6133 9.3005
R11813 gnd.n1215 gnd.n1214 9.3005
R11814 gnd.n6140 gnd.n6139 9.3005
R11815 gnd.n6142 gnd.n6141 9.3005
R11816 gnd.n1205 gnd.n1204 9.3005
R11817 gnd.n6148 gnd.n6147 9.3005
R11818 gnd.n6150 gnd.n6149 9.3005
R11819 gnd.n1197 gnd.n1196 9.3005
R11820 gnd.n6156 gnd.n6155 9.3005
R11821 gnd.n6158 gnd.n6157 9.3005
R11822 gnd.n1186 gnd.n1184 9.3005
R11823 gnd.n6164 gnd.n6163 9.3005
R11824 gnd.n6165 gnd.n1179 9.3005
R11825 gnd.n6167 gnd.n6166 9.3005
R11826 gnd.n6169 gnd.n1178 9.3005
R11827 gnd.n6171 gnd.n6170 9.3005
R11828 gnd.n6172 gnd.n1174 9.3005
R11829 gnd.n6174 gnd.n6173 9.3005
R11830 gnd.n6175 gnd.n1173 9.3005
R11831 gnd.n6177 gnd.n6176 9.3005
R11832 gnd.n6178 gnd.n1172 9.3005
R11833 gnd.n4451 gnd.n4450 9.3005
R11834 gnd.n4452 gnd.n2309 9.3005
R11835 gnd.n4455 gnd.n4454 9.3005
R11836 gnd.n4453 gnd.n2310 9.3005
R11837 gnd.n2288 gnd.n2287 9.3005
R11838 gnd.n4484 gnd.n4483 9.3005
R11839 gnd.n4485 gnd.n2285 9.3005
R11840 gnd.n4491 gnd.n4490 9.3005
R11841 gnd.n4489 gnd.n2286 9.3005
R11842 gnd.n4488 gnd.n4487 9.3005
R11843 gnd.n1497 gnd.n1495 9.3005
R11844 gnd.n5982 gnd.n5981 9.3005
R11845 gnd.n5980 gnd.n1496 9.3005
R11846 gnd.n5979 gnd.n5978 9.3005
R11847 gnd.n5977 gnd.n1498 9.3005
R11848 gnd.n5976 gnd.n5975 9.3005
R11849 gnd.n5974 gnd.n1502 9.3005
R11850 gnd.n5973 gnd.n5972 9.3005
R11851 gnd.n5971 gnd.n1503 9.3005
R11852 gnd.n5970 gnd.n5969 9.3005
R11853 gnd.n5968 gnd.n1507 9.3005
R11854 gnd.n5967 gnd.n5966 9.3005
R11855 gnd.n5965 gnd.n1508 9.3005
R11856 gnd.n5964 gnd.n5963 9.3005
R11857 gnd.n5962 gnd.n1512 9.3005
R11858 gnd.n5961 gnd.n5960 9.3005
R11859 gnd.n5959 gnd.n1513 9.3005
R11860 gnd.n5958 gnd.n5957 9.3005
R11861 gnd.n5956 gnd.n1517 9.3005
R11862 gnd.n5955 gnd.n5954 9.3005
R11863 gnd.n5953 gnd.n1518 9.3005
R11864 gnd.n5952 gnd.n5951 9.3005
R11865 gnd.n5950 gnd.n1522 9.3005
R11866 gnd.n5949 gnd.n5948 9.3005
R11867 gnd.n5947 gnd.n1523 9.3005
R11868 gnd.n5946 gnd.n5945 9.3005
R11869 gnd.n5944 gnd.n1527 9.3005
R11870 gnd.n5943 gnd.n5942 9.3005
R11871 gnd.n5941 gnd.n1528 9.3005
R11872 gnd.n5940 gnd.n5939 9.3005
R11873 gnd.n5938 gnd.n1532 9.3005
R11874 gnd.n5937 gnd.n5936 9.3005
R11875 gnd.n5935 gnd.n1533 9.3005
R11876 gnd.n5934 gnd.n5933 9.3005
R11877 gnd.n5932 gnd.n1537 9.3005
R11878 gnd.n5931 gnd.n5930 9.3005
R11879 gnd.n5929 gnd.n1538 9.3005
R11880 gnd.n5928 gnd.n5927 9.3005
R11881 gnd.n5926 gnd.n1542 9.3005
R11882 gnd.n5925 gnd.n5924 9.3005
R11883 gnd.n5923 gnd.n1543 9.3005
R11884 gnd.n5922 gnd.n5921 9.3005
R11885 gnd.n5920 gnd.n1547 9.3005
R11886 gnd.n5919 gnd.n5918 9.3005
R11887 gnd.n5917 gnd.n1548 9.3005
R11888 gnd.n5916 gnd.n5915 9.3005
R11889 gnd.n5914 gnd.n1552 9.3005
R11890 gnd.n5913 gnd.n5912 9.3005
R11891 gnd.n5911 gnd.n1553 9.3005
R11892 gnd.n5910 gnd.n5909 9.3005
R11893 gnd.n5908 gnd.n1557 9.3005
R11894 gnd.n5907 gnd.n5906 9.3005
R11895 gnd.n5905 gnd.n1558 9.3005
R11896 gnd.n5904 gnd.n5903 9.3005
R11897 gnd.n5902 gnd.n1562 9.3005
R11898 gnd.n5901 gnd.n5900 9.3005
R11899 gnd.n5899 gnd.n1563 9.3005
R11900 gnd.n5898 gnd.n5897 9.3005
R11901 gnd.n5896 gnd.n1567 9.3005
R11902 gnd.n5895 gnd.n5894 9.3005
R11903 gnd.n5893 gnd.n1568 9.3005
R11904 gnd.n5892 gnd.n5891 9.3005
R11905 gnd.n5890 gnd.n1572 9.3005
R11906 gnd.n5889 gnd.n5888 9.3005
R11907 gnd.n5887 gnd.n1573 9.3005
R11908 gnd.n5886 gnd.n5885 9.3005
R11909 gnd.n5884 gnd.n1577 9.3005
R11910 gnd.n5883 gnd.n5882 9.3005
R11911 gnd.n5881 gnd.n1578 9.3005
R11912 gnd.n5880 gnd.n5879 9.3005
R11913 gnd.n5878 gnd.n1582 9.3005
R11914 gnd.n5877 gnd.n5876 9.3005
R11915 gnd.n2312 gnd.n2311 9.3005
R11916 gnd.n5185 gnd.n5184 9.3005
R11917 gnd.n5181 gnd.n5180 9.3005
R11918 gnd.n5192 gnd.n5191 9.3005
R11919 gnd.n5193 gnd.n5179 9.3005
R11920 gnd.n5196 gnd.n5195 9.3005
R11921 gnd.n5194 gnd.n5177 9.3005
R11922 gnd.n5183 gnd.n1583 9.3005
R11923 gnd.n5284 gnd.n5133 9.3005
R11924 gnd.n5146 gnd.n5142 9.3005
R11925 gnd.n5278 gnd.n5277 9.3005
R11926 gnd.n5266 gnd.n5144 9.3005
R11927 gnd.n5265 gnd.n5264 9.3005
R11928 gnd.n5155 gnd.n5151 9.3005
R11929 gnd.n5258 gnd.n5257 9.3005
R11930 gnd.n5247 gnd.n5153 9.3005
R11931 gnd.n5246 gnd.n5245 9.3005
R11932 gnd.n5164 gnd.n5160 9.3005
R11933 gnd.n5239 gnd.n5238 9.3005
R11934 gnd.n5228 gnd.n5162 9.3005
R11935 gnd.n5227 gnd.n5226 9.3005
R11936 gnd.n5173 gnd.n5169 9.3005
R11937 gnd.n5220 gnd.n5219 9.3005
R11938 gnd.n5209 gnd.n5171 9.3005
R11939 gnd.n5208 gnd.n5207 9.3005
R11940 gnd.n5286 gnd.n5285 9.3005
R11941 gnd.n5137 gnd.n5136 9.3005
R11942 gnd.n5203 gnd.n5202 9.3005
R11943 gnd.n5204 gnd.n5176 9.3005
R11944 gnd.n5211 gnd.n5210 9.3005
R11945 gnd.n5174 gnd.n5172 9.3005
R11946 gnd.n5218 gnd.n5217 9.3005
R11947 gnd.n5168 gnd.n5167 9.3005
R11948 gnd.n5230 gnd.n5229 9.3005
R11949 gnd.n5165 gnd.n5163 9.3005
R11950 gnd.n5237 gnd.n5236 9.3005
R11951 gnd.n5159 gnd.n5158 9.3005
R11952 gnd.n5249 gnd.n5248 9.3005
R11953 gnd.n5156 gnd.n5154 9.3005
R11954 gnd.n5256 gnd.n5255 9.3005
R11955 gnd.n5150 gnd.n5149 9.3005
R11956 gnd.n5268 gnd.n5267 9.3005
R11957 gnd.n5147 gnd.n5145 9.3005
R11958 gnd.n5276 gnd.n5275 9.3005
R11959 gnd.n5274 gnd.n5273 9.3005
R11960 gnd.n5288 gnd.n5287 9.3005
R11961 gnd.n5134 gnd.n5128 9.3005
R11962 gnd.n5135 gnd.n5127 9.3005
R11963 gnd.n5123 gnd.n5120 9.3005
R11964 gnd.n1750 gnd.n1749 9.3005
R11965 gnd.n5672 gnd.n5671 9.3005
R11966 gnd.n5673 gnd.n1748 9.3005
R11967 gnd.n5675 gnd.n5674 9.3005
R11968 gnd.n1744 gnd.n1742 9.3005
R11969 gnd.n5695 gnd.n5694 9.3005
R11970 gnd.n5693 gnd.n1743 9.3005
R11971 gnd.n5692 gnd.n5691 9.3005
R11972 gnd.n5690 gnd.n1745 9.3005
R11973 gnd.n5689 gnd.n5688 9.3005
R11974 gnd.n1733 gnd.n1732 9.3005
R11975 gnd.n5752 gnd.n5751 9.3005
R11976 gnd.n5753 gnd.n1730 9.3005
R11977 gnd.n5765 gnd.n5764 9.3005
R11978 gnd.n5763 gnd.n1731 9.3005
R11979 gnd.n5762 gnd.n5761 9.3005
R11980 gnd.n5760 gnd.n5754 9.3005
R11981 gnd.n5759 gnd.n5758 9.3005
R11982 gnd.n5757 gnd.n63 9.3005
R11983 gnd.n5125 gnd.n5124 9.3005
R11984 gnd.n7344 gnd.n64 9.3005
R11985 gnd.t172 gnd.n2640 9.24152
R11986 gnd.n2542 gnd.t118 9.24152
R11987 gnd.n3810 gnd.t93 9.24152
R11988 gnd.n4410 gnd.t136 9.24152
R11989 gnd.n5698 gnd.t151 9.24152
R11990 gnd.t322 gnd.t172 8.92286
R11991 gnd.n5985 gnd.t103 8.92286
R11992 gnd.n4511 gnd.n2192 8.92286
R11993 gnd.t258 gnd.n4536 8.92286
R11994 gnd.n4696 gnd.n2101 8.92286
R11995 gnd.n4741 gnd.n2071 8.92286
R11996 gnd.n4866 gnd.n2004 8.92286
R11997 gnd.n4937 gnd.n4936 8.92286
R11998 gnd.n1909 gnd.t141 8.92286
R11999 gnd.n5077 gnd.n5076 8.92286
R12000 gnd.n5414 gnd.t77 8.92286
R12001 gnd.n3780 gnd.n3755 8.92171
R12002 gnd.n3748 gnd.n3723 8.92171
R12003 gnd.n3716 gnd.n3691 8.92171
R12004 gnd.n3685 gnd.n3660 8.92171
R12005 gnd.n3653 gnd.n3628 8.92171
R12006 gnd.n3621 gnd.n3596 8.92171
R12007 gnd.n3589 gnd.n3564 8.92171
R12008 gnd.n3558 gnd.n3533 8.92171
R12009 gnd.n5346 gnd.n5328 8.72777
R12010 gnd.n3284 gnd.t293 8.60421
R12011 gnd.n2704 gnd.n2692 8.43656
R12012 gnd.n38 gnd.n26 8.43656
R12013 gnd.n4671 gnd.n2116 8.28555
R12014 gnd.n4762 gnd.n2054 8.28555
R12015 gnd.n4846 gnd.n2019 8.28555
R12016 gnd.n4902 gnd.n1971 8.28555
R12017 gnd.n3781 gnd.n3753 8.14595
R12018 gnd.n3749 gnd.n3721 8.14595
R12019 gnd.n3717 gnd.n3689 8.14595
R12020 gnd.n3686 gnd.n3658 8.14595
R12021 gnd.n3654 gnd.n3626 8.14595
R12022 gnd.n3622 gnd.n3594 8.14595
R12023 gnd.n3590 gnd.n3562 8.14595
R12024 gnd.n3559 gnd.n3531 8.14595
R12025 gnd.n4293 gnd.n0 8.10675
R12026 gnd.n7345 gnd.n7344 8.10675
R12027 gnd.n3786 gnd.n3785 7.97301
R12028 gnd.t12 gnd.n2799 7.9669
R12029 gnd.n7345 gnd.n62 7.78567
R12030 gnd.n5285 gnd.n5137 7.75808
R12031 gnd.n6120 gnd.n6119 7.75808
R12032 gnd.n7251 gnd.n7189 7.75808
R12033 gnd.n4052 gnd.n4033 7.75808
R12034 gnd.n4504 gnd.n2196 7.64824
R12035 gnd.n4671 gnd.n2115 7.64824
R12036 gnd.t259 gnd.n4715 7.64824
R12037 gnd.n4763 gnd.t0 7.64824
R12038 gnd.n4773 gnd.n2054 7.64824
R12039 gnd.n4846 gnd.n2017 7.64824
R12040 gnd.t224 gnd.n2012 7.64824
R12041 gnd.n4865 gnd.t256 7.64824
R12042 gnd.n4902 gnd.n1962 7.64824
R12043 gnd.n2729 gnd.n2728 7.53171
R12044 gnd.n3193 gnd.t174 7.32958
R12045 gnd.n4504 gnd.t222 7.32958
R12046 gnd.t201 gnd.n5095 7.32958
R12047 gnd.n1475 gnd.n1474 7.30353
R12048 gnd.n5345 gnd.n5344 7.30353
R12049 gnd.n3153 gnd.n2872 7.01093
R12050 gnd.n2875 gnd.n2873 7.01093
R12051 gnd.n3163 gnd.n3162 7.01093
R12052 gnd.n3174 gnd.n2856 7.01093
R12053 gnd.n3173 gnd.n2859 7.01093
R12054 gnd.n3184 gnd.n2847 7.01093
R12055 gnd.n2850 gnd.n2848 7.01093
R12056 gnd.n3194 gnd.n3193 7.01093
R12057 gnd.n3204 gnd.n2828 7.01093
R12058 gnd.n3203 gnd.n2831 7.01093
R12059 gnd.n3212 gnd.n2822 7.01093
R12060 gnd.n3224 gnd.n2812 7.01093
R12061 gnd.n3234 gnd.n2797 7.01093
R12062 gnd.n3250 gnd.n3249 7.01093
R12063 gnd.n2799 gnd.n2736 7.01093
R12064 gnd.n3304 gnd.n2737 7.01093
R12065 gnd.n3298 gnd.n3297 7.01093
R12066 gnd.n2786 gnd.n2748 7.01093
R12067 gnd.n3290 gnd.n2759 7.01093
R12068 gnd.n2777 gnd.n2772 7.01093
R12069 gnd.n3284 gnd.n3283 7.01093
R12070 gnd.n3330 gnd.n2675 7.01093
R12071 gnd.n3329 gnd.n3328 7.01093
R12072 gnd.n3341 gnd.n3340 7.01093
R12073 gnd.n2668 gnd.n2660 7.01093
R12074 gnd.n3370 gnd.n2648 7.01093
R12075 gnd.n3369 gnd.n2651 7.01093
R12076 gnd.n3380 gnd.n2640 7.01093
R12077 gnd.n2641 gnd.n2629 7.01093
R12078 gnd.n3391 gnd.n2630 7.01093
R12079 gnd.n3415 gnd.n2621 7.01093
R12080 gnd.n3414 gnd.n2612 7.01093
R12081 gnd.n3437 gnd.n3436 7.01093
R12082 gnd.n3455 gnd.n2593 7.01093
R12083 gnd.n3454 gnd.n2596 7.01093
R12084 gnd.n3465 gnd.n2585 7.01093
R12085 gnd.n2586 gnd.n2573 7.01093
R12086 gnd.n3476 gnd.n2574 7.01093
R12087 gnd.n3503 gnd.n2558 7.01093
R12088 gnd.n3515 gnd.n3514 7.01093
R12089 gnd.n3497 gnd.n2551 7.01093
R12090 gnd.n3526 gnd.n3525 7.01093
R12091 gnd.n3798 gnd.n2539 7.01093
R12092 gnd.n3797 gnd.n2542 7.01093
R12093 gnd.n3810 gnd.n2531 7.01093
R12094 gnd.n2532 gnd.n2524 7.01093
R12095 gnd.n3820 gnd.n2450 7.01093
R12096 gnd.n4518 gnd.n4511 7.01093
R12097 gnd.n4577 gnd.n2161 7.01093
R12098 gnd.t3 gnd.n4576 7.01093
R12099 gnd.n4696 gnd.n4695 7.01093
R12100 gnd.n4716 gnd.t259 7.01093
R12101 gnd.n4715 gnd.n2071 7.01093
R12102 gnd.n4866 gnd.n4865 7.01093
R12103 gnd.t256 gnd.n4864 7.01093
R12104 gnd.n4937 gnd.n1975 7.01093
R12105 gnd.n5018 gnd.t261 7.01093
R12106 gnd.n5034 gnd.n5033 7.01093
R12107 gnd.n5079 gnd.n5077 7.01093
R12108 gnd.n2831 gnd.t166 6.69227
R12109 gnd.n2651 gnd.t322 6.69227
R12110 gnd.n3504 gnd.t13 6.69227
R12111 gnd.t277 gnd.n2156 6.69227
R12112 gnd.n4971 gnd.t317 6.69227
R12113 gnd.n5475 gnd.n5474 6.5566
R12114 gnd.n2211 gnd.n2210 6.5566
R12115 gnd.n6003 gnd.n5999 6.5566
R12116 gnd.n5353 gnd.n5352 6.5566
R12117 gnd.n2593 gnd.n960 6.37362
R12118 gnd.n2282 gnd.n2281 6.37362
R12119 gnd.t103 gnd.t80 6.37362
R12120 gnd.n4638 gnd.n2130 6.37362
R12121 gnd.n4723 gnd.t257 6.37362
R12122 gnd.n4781 gnd.n2048 6.37362
R12123 gnd.n4793 gnd.n2035 6.37362
R12124 gnd.n4915 gnd.t142 6.37362
R12125 gnd.n4962 gnd.n1958 6.37362
R12126 gnd.n5076 gnd.t15 6.37362
R12127 gnd.n5087 gnd.t15 6.37362
R12128 gnd.n5414 gnd.n1828 6.37362
R12129 gnd.n1235 gnd.n1233 6.20656
R12130 gnd.n5288 gnd.n5132 6.20656
R12131 gnd.t326 gnd.n3260 6.05496
R12132 gnd.n3261 gnd.t167 6.05496
R12133 gnd.t310 gnd.n2675 6.05496
R12134 gnd.t10 gnd.n3425 6.05496
R12135 gnd.t225 gnd.t263 6.05496
R12136 gnd.t232 gnd.t227 6.05496
R12137 gnd.n3783 gnd.n3753 5.81868
R12138 gnd.n3751 gnd.n3721 5.81868
R12139 gnd.n3719 gnd.n3689 5.81868
R12140 gnd.n3688 gnd.n3658 5.81868
R12141 gnd.n3656 gnd.n3626 5.81868
R12142 gnd.n3624 gnd.n3594 5.81868
R12143 gnd.n3592 gnd.n3562 5.81868
R12144 gnd.n3561 gnd.n3531 5.81868
R12145 gnd.n2185 gnd.n2184 5.73631
R12146 gnd.n4537 gnd.n4534 5.73631
R12147 gnd.n2096 gnd.n2084 5.73631
R12148 gnd.n4707 gnd.n2077 5.73631
R12149 gnd.t0 gnd.n4762 5.73631
R12150 gnd.n2019 gnd.t224 5.73631
R12151 gnd.n4803 gnd.n4801 5.73631
R12152 gnd.n4873 gnd.n1993 5.73631
R12153 gnd.n5054 gnd.n1900 5.73631
R12154 gnd.n1902 gnd.n1892 5.73631
R12155 gnd.n5484 gnd.n1787 5.62001
R12156 gnd.n6065 gnd.n1417 5.62001
R12157 gnd.n6065 gnd.n1418 5.62001
R12158 gnd.n5484 gnd.n1788 5.62001
R12159 gnd.n3012 gnd.n3007 5.4308
R12160 gnd.n3828 gnd.n2517 5.4308
R12161 gnd.n3328 gnd.t11 5.41765
R12162 gnd.t294 gnd.n3351 5.41765
R12163 gnd.t192 gnd.n2605 5.41765
R12164 gnd.t211 gnd.n4654 5.41765
R12165 gnd.n4894 gnd.t299 5.41765
R12166 gnd.t214 gnd.n4568 5.09899
R12167 gnd.n4646 gnd.n2134 5.09899
R12168 gnd.n4822 gnd.n2039 5.09899
R12169 gnd.n4830 gnd.n2032 5.09899
R12170 gnd.n4995 gnd.n1942 5.09899
R12171 gnd.n1933 gnd.t231 5.09899
R12172 gnd.n3781 gnd.n3780 5.04292
R12173 gnd.n3749 gnd.n3748 5.04292
R12174 gnd.n3717 gnd.n3716 5.04292
R12175 gnd.n3686 gnd.n3685 5.04292
R12176 gnd.n3654 gnd.n3653 5.04292
R12177 gnd.n3622 gnd.n3621 5.04292
R12178 gnd.n3590 gnd.n3589 5.04292
R12179 gnd.n3559 gnd.n3558 5.04292
R12180 gnd.n3291 gnd.t219 4.78034
R12181 gnd.n2630 gnd.t218 4.78034
R12182 gnd.t246 gnd.n4480 4.78034
R12183 gnd.n5481 gnd.t54 4.78034
R12184 gnd.n5315 gnd.t312 4.78034
R12185 gnd.n2733 gnd.n2730 4.74817
R12186 gnd.n2783 gnd.n2681 4.74817
R12187 gnd.n2770 gnd.n2680 4.74817
R12188 gnd.n2679 gnd.n2678 4.74817
R12189 gnd.n2779 gnd.n2730 4.74817
R12190 gnd.n2780 gnd.n2681 4.74817
R12191 gnd.n2782 gnd.n2680 4.74817
R12192 gnd.n2769 gnd.n2679 4.74817
R12193 gnd.n1696 gnd.n82 4.74817
R12194 gnd.n5794 gnd.n81 4.74817
R12195 gnd.n1713 gnd.n80 4.74817
R12196 gnd.n7337 gnd.n75 4.74817
R12197 gnd.n7335 gnd.n76 4.74817
R12198 gnd.n5808 gnd.n82 4.74817
R12199 gnd.n1695 gnd.n81 4.74817
R12200 gnd.n5795 gnd.n80 4.74817
R12201 gnd.n1712 gnd.n75 4.74817
R12202 gnd.n7336 gnd.n7335 4.74817
R12203 gnd.n2367 gnd.n2364 4.74817
R12204 gnd.n4323 gnd.n2363 4.74817
R12205 gnd.n4319 gnd.n2362 4.74817
R12206 gnd.n2386 gnd.n2361 4.74817
R12207 gnd.n2382 gnd.n2360 4.74817
R12208 gnd.n5803 gnd.n1702 4.74817
R12209 gnd.n5801 gnd.n5800 4.74817
R12210 gnd.n1720 gnd.n1717 4.74817
R12211 gnd.n1718 gnd.n404 4.74817
R12212 gnd.n7133 gnd.n7132 4.74817
R12213 gnd.n5732 gnd.n1702 4.74817
R12214 gnd.n5802 gnd.n5801 4.74817
R12215 gnd.n1717 gnd.n1703 4.74817
R12216 gnd.n1719 gnd.n1718 4.74817
R12217 gnd.n7134 gnd.n7133 4.74817
R12218 gnd.n6277 gnd.n6276 4.74817
R12219 gnd.n1038 gnd.n1020 4.74817
R12220 gnd.n6264 gnd.n6263 4.74817
R12221 gnd.n1055 gnd.n1039 4.74817
R12222 gnd.n6251 gnd.n6250 4.74817
R12223 gnd.n6278 gnd.n6277 4.74817
R12224 gnd.n6275 gnd.n1020 4.74817
R12225 gnd.n6265 gnd.n6264 4.74817
R12226 gnd.n6262 gnd.n1039 4.74817
R12227 gnd.n6252 gnd.n6251 4.74817
R12228 gnd.n2379 gnd.n2364 4.74817
R12229 gnd.n2380 gnd.n2363 4.74817
R12230 gnd.n4322 gnd.n2362 4.74817
R12231 gnd.n4318 gnd.n2361 4.74817
R12232 gnd.n2385 gnd.n2360 4.74817
R12233 gnd.n2728 gnd.n2727 4.74296
R12234 gnd.n62 gnd.n61 4.74296
R12235 gnd.n2704 gnd.n2703 4.7074
R12236 gnd.n2716 gnd.n2715 4.7074
R12237 gnd.n38 gnd.n37 4.7074
R12238 gnd.n50 gnd.n49 4.7074
R12239 gnd.n2728 gnd.n2716 4.65959
R12240 gnd.n62 gnd.n50 4.65959
R12241 gnd.n5575 gnd.n5485 4.6132
R12242 gnd.n6066 gnd.n1416 4.6132
R12243 gnd.n4544 gnd.n2177 4.46168
R12244 gnd.n4535 gnd.n2166 4.46168
R12245 gnd.n4693 gnd.t213 4.46168
R12246 gnd.n4703 gnd.n4702 4.46168
R12247 gnd.n4732 gnd.n2079 4.46168
R12248 gnd.n4880 gnd.n1998 4.46168
R12249 gnd.n4924 gnd.n1985 4.46168
R12250 gnd.t2 gnd.n4923 4.46168
R12251 gnd.n5044 gnd.n1908 4.46168
R12252 gnd.n5064 gnd.n5063 4.46168
R12253 gnd.t129 gnd.n1833 4.46168
R12254 gnd.n5341 gnd.n5328 4.46111
R12255 gnd.n3766 gnd.n3762 4.38594
R12256 gnd.n3734 gnd.n3730 4.38594
R12257 gnd.n3702 gnd.n3698 4.38594
R12258 gnd.n3671 gnd.n3667 4.38594
R12259 gnd.n3639 gnd.n3635 4.38594
R12260 gnd.n3607 gnd.n3603 4.38594
R12261 gnd.n3575 gnd.n3571 4.38594
R12262 gnd.n3544 gnd.n3540 4.38594
R12263 gnd.n3777 gnd.n3755 4.26717
R12264 gnd.n3745 gnd.n3723 4.26717
R12265 gnd.n3713 gnd.n3691 4.26717
R12266 gnd.n3682 gnd.n3660 4.26717
R12267 gnd.n3650 gnd.n3628 4.26717
R12268 gnd.n3618 gnd.n3596 4.26717
R12269 gnd.n3586 gnd.n3564 4.26717
R12270 gnd.n3555 gnd.n3533 4.26717
R12271 gnd.n3235 gnd.t217 4.14303
R12272 gnd.n3465 gnd.t292 4.14303
R12273 gnd.t46 gnd.n1131 4.14303
R12274 gnd.t26 gnd.n1618 4.14303
R12275 gnd.n3785 gnd.n3784 4.08274
R12276 gnd.n5474 gnd.n5473 4.05904
R12277 gnd.n2212 gnd.n2211 4.05904
R12278 gnd.n6006 gnd.n5999 4.05904
R12279 gnd.n5354 gnd.n5353 4.05904
R12280 gnd.n15 gnd.n7 3.99943
R12281 gnd.n5992 gnd.n5991 3.82437
R12282 gnd.n4603 gnd.n2147 3.82437
R12283 gnd.n4644 gnd.t226 3.82437
R12284 gnd.n4664 gnd.n4663 3.82437
R12285 gnd.n4752 gnd.n2068 3.82437
R12286 gnd.n4753 gnd.t225 3.82437
R12287 gnd.n4794 gnd.t232 3.82437
R12288 gnd.n4839 gnd.n4838 3.82437
R12289 gnd.n4954 gnd.n1956 3.82437
R12290 gnd.n4987 gnd.t4 3.82437
R12291 gnd.n5004 gnd.n5003 3.82437
R12292 gnd.n5322 gnd.n1836 3.82437
R12293 gnd.n3308 gnd.n2729 3.81325
R12294 gnd.n2716 gnd.n2704 3.72967
R12295 gnd.n50 gnd.n38 3.72967
R12296 gnd.n3785 gnd.n3657 3.70378
R12297 gnd.n15 gnd.n14 3.60163
R12298 gnd.t173 gnd.n960 3.50571
R12299 gnd.n3776 gnd.n3757 3.49141
R12300 gnd.n3744 gnd.n3725 3.49141
R12301 gnd.n3712 gnd.n3693 3.49141
R12302 gnd.n3681 gnd.n3662 3.49141
R12303 gnd.n3649 gnd.n3630 3.49141
R12304 gnd.n3617 gnd.n3598 3.49141
R12305 gnd.n3585 gnd.n3566 3.49141
R12306 gnd.n3554 gnd.n3535 3.49141
R12307 gnd.n5556 gnd.n5555 3.29747
R12308 gnd.n5555 gnd.n5493 3.29747
R12309 gnd.n284 gnd.n220 3.29747
R12310 gnd.n279 gnd.n220 3.29747
R12311 gnd.n4180 gnd.n4179 3.29747
R12312 gnd.n4179 gnd.n4178 3.29747
R12313 gnd.n6084 gnd.n6083 3.29747
R12314 gnd.n6083 gnd.n6082 3.29747
R12315 gnd.n5984 gnd.n1492 3.18706
R12316 gnd.n2185 gnd.t84 3.18706
R12317 gnd.n4575 gnd.n2154 3.18706
R12318 gnd.n4584 gnd.t260 3.18706
R12319 gnd.t260 gnd.n2139 3.18706
R12320 gnd.n4682 gnd.n4680 3.18706
R12321 gnd.n4743 gnd.n4742 3.18706
R12322 gnd.n4854 gnd.n4853 3.18706
R12323 gnd.n4935 gnd.n4934 3.18706
R12324 gnd.t140 gnd.n1945 3.18706
R12325 gnd.n4885 gnd.t140 3.18706
R12326 gnd.n5020 gnd.n5019 3.18706
R12327 gnd.n5087 gnd.n1877 3.18706
R12328 gnd.n5095 gnd.t129 3.18706
R12329 gnd.n2814 gnd.t217 2.8684
R12330 gnd.n4551 gnd.t275 2.8684
R12331 gnd.t229 gnd.n5053 2.8684
R12332 gnd.n2717 gnd.t298 2.82907
R12333 gnd.n2717 gnd.t207 2.82907
R12334 gnd.n2719 gnd.t309 2.82907
R12335 gnd.n2719 gnd.t245 2.82907
R12336 gnd.n2721 gnd.t241 2.82907
R12337 gnd.n2721 gnd.t243 2.82907
R12338 gnd.n2723 gnd.t281 2.82907
R12339 gnd.n2723 gnd.t251 2.82907
R12340 gnd.n2725 gnd.t210 2.82907
R12341 gnd.n2725 gnd.t279 2.82907
R12342 gnd.n2682 gnd.t302 2.82907
R12343 gnd.n2682 gnd.t237 2.82907
R12344 gnd.n2684 gnd.t215 2.82907
R12345 gnd.n2684 gnd.t249 2.82907
R12346 gnd.n2686 gnd.t236 2.82907
R12347 gnd.n2686 gnd.t306 2.82907
R12348 gnd.n2688 gnd.t286 2.82907
R12349 gnd.n2688 gnd.t158 2.82907
R12350 gnd.n2690 gnd.t176 2.82907
R12351 gnd.n2690 gnd.t270 2.82907
R12352 gnd.n2693 gnd.t288 2.82907
R12353 gnd.n2693 gnd.t250 2.82907
R12354 gnd.n2695 gnd.t265 2.82907
R12355 gnd.n2695 gnd.t204 2.82907
R12356 gnd.n2697 gnd.t156 2.82907
R12357 gnd.n2697 gnd.t198 2.82907
R12358 gnd.n2699 gnd.t273 2.82907
R12359 gnd.n2699 gnd.t321 2.82907
R12360 gnd.n2701 gnd.t316 2.82907
R12361 gnd.n2701 gnd.t267 2.82907
R12362 gnd.n2705 gnd.t307 2.82907
R12363 gnd.n2705 gnd.t255 2.82907
R12364 gnd.n2707 gnd.t186 2.82907
R12365 gnd.n2707 gnd.t240 2.82907
R12366 gnd.n2709 gnd.t285 2.82907
R12367 gnd.n2709 gnd.t272 2.82907
R12368 gnd.n2711 gnd.t139 2.82907
R12369 gnd.n2711 gnd.t269 2.82907
R12370 gnd.n2713 gnd.t216 2.82907
R12371 gnd.n2713 gnd.t314 2.82907
R12372 gnd.n59 gnd.t242 2.82907
R12373 gnd.n59 gnd.t160 2.82907
R12374 gnd.n57 gnd.t194 2.82907
R12375 gnd.n57 gnd.t189 2.82907
R12376 gnd.n55 gnd.t150 2.82907
R12377 gnd.n55 gnd.t252 2.82907
R12378 gnd.n53 gnd.t295 2.82907
R12379 gnd.n53 gnd.t208 2.82907
R12380 gnd.n51 gnd.t280 2.82907
R12381 gnd.n51 gnd.t297 2.82907
R12382 gnd.n24 gnd.t181 2.82907
R12383 gnd.n24 gnd.t283 2.82907
R12384 gnd.n22 gnd.t234 2.82907
R12385 gnd.n22 gnd.t282 2.82907
R12386 gnd.n20 gnd.t271 2.82907
R12387 gnd.n20 gnd.t304 2.82907
R12388 gnd.n18 gnd.t180 2.82907
R12389 gnd.n18 gnd.t154 2.82907
R12390 gnd.n16 gnd.t308 2.82907
R12391 gnd.n16 gnd.t183 2.82907
R12392 gnd.n35 gnd.t235 2.82907
R12393 gnd.n35 gnd.t182 2.82907
R12394 gnd.n33 gnd.t135 2.82907
R12395 gnd.n33 gnd.t291 2.82907
R12396 gnd.n31 gnd.t296 2.82907
R12397 gnd.n31 gnd.t9 2.82907
R12398 gnd.n29 gnd.t187 2.82907
R12399 gnd.n29 gnd.t168 2.82907
R12400 gnd.n27 gnd.t191 2.82907
R12401 gnd.n27 gnd.t233 2.82907
R12402 gnd.n47 gnd.t163 2.82907
R12403 gnd.n47 gnd.t238 2.82907
R12404 gnd.n45 gnd.t184 2.82907
R12405 gnd.n45 gnd.t301 2.82907
R12406 gnd.n43 gnd.t305 2.82907
R12407 gnd.n43 gnd.t239 2.82907
R12408 gnd.n41 gnd.t253 2.82907
R12409 gnd.n41 gnd.t284 2.82907
R12410 gnd.n39 gnd.t196 2.82907
R12411 gnd.n39 gnd.t178 2.82907
R12412 gnd.n3773 gnd.n3772 2.71565
R12413 gnd.n3741 gnd.n3740 2.71565
R12414 gnd.n3709 gnd.n3708 2.71565
R12415 gnd.n3678 gnd.n3677 2.71565
R12416 gnd.n3646 gnd.n3645 2.71565
R12417 gnd.n3614 gnd.n3613 2.71565
R12418 gnd.n3582 gnd.n3581 2.71565
R12419 gnd.n3551 gnd.n3550 2.71565
R12420 gnd.n5985 gnd.n1490 2.54975
R12421 gnd.n4593 gnd.n4592 2.54975
R12422 gnd.n4569 gnd.t214 2.54975
R12423 gnd.n4683 gnd.n2110 2.54975
R12424 gnd.n4683 gnd.t248 2.54975
R12425 gnd.n4763 gnd.n2061 2.54975
R12426 gnd.n4855 gnd.n2012 2.54975
R12427 gnd.n4944 gnd.t1 2.54975
R12428 gnd.n4944 gnd.n4943 2.54975
R12429 gnd.n5011 gnd.t231 2.54975
R12430 gnd.n5021 gnd.n1922 2.54975
R12431 gnd.n1886 gnd.n1873 2.54975
R12432 gnd.n3308 gnd.n2730 2.27742
R12433 gnd.n3308 gnd.n2681 2.27742
R12434 gnd.n3308 gnd.n2680 2.27742
R12435 gnd.n3308 gnd.n2679 2.27742
R12436 gnd.n7334 gnd.n82 2.27742
R12437 gnd.n7334 gnd.n81 2.27742
R12438 gnd.n7334 gnd.n80 2.27742
R12439 gnd.n7334 gnd.n75 2.27742
R12440 gnd.n7335 gnd.n7334 2.27742
R12441 gnd.n1702 gnd.n79 2.27742
R12442 gnd.n5801 gnd.n79 2.27742
R12443 gnd.n1717 gnd.n79 2.27742
R12444 gnd.n1718 gnd.n79 2.27742
R12445 gnd.n7133 gnd.n79 2.27742
R12446 gnd.n6277 gnd.n1018 2.27742
R12447 gnd.n1020 gnd.n1018 2.27742
R12448 gnd.n6264 gnd.n1018 2.27742
R12449 gnd.n1039 gnd.n1018 2.27742
R12450 gnd.n6251 gnd.n1018 2.27742
R12451 gnd.n4338 gnd.n2364 2.27742
R12452 gnd.n4338 gnd.n2363 2.27742
R12453 gnd.n4338 gnd.n2362 2.27742
R12454 gnd.n4338 gnd.n2361 2.27742
R12455 gnd.n4338 gnd.n2360 2.27742
R12456 gnd.n3162 gnd.t60 2.23109
R12457 gnd.n2785 gnd.t219 2.23109
R12458 gnd.t199 gnd.n2079 2.23109
R12459 gnd.t263 gnd.n4752 2.23109
R12460 gnd.n4839 gnd.t227 2.23109
R12461 gnd.t319 gnd.n1998 2.23109
R12462 gnd.n3769 gnd.n3759 1.93989
R12463 gnd.n3737 gnd.n3727 1.93989
R12464 gnd.n3705 gnd.n3695 1.93989
R12465 gnd.n3674 gnd.n3664 1.93989
R12466 gnd.n3642 gnd.n3632 1.93989
R12467 gnd.n3610 gnd.n3600 1.93989
R12468 gnd.n3578 gnd.n3568 1.93989
R12469 gnd.n3547 gnd.n3537 1.93989
R12470 gnd.n2275 gnd.n1481 1.91244
R12471 gnd.n2275 gnd.t40 1.91244
R12472 gnd.n4577 gnd.t3 1.91244
R12473 gnd.n4605 gnd.n2146 1.91244
R12474 gnd.n4613 gnd.n4612 1.91244
R12475 gnd.n4772 gnd.n2056 1.91244
R12476 gnd.n2026 gnd.n2025 1.91244
R12477 gnd.n4956 gnd.n4955 1.91244
R12478 gnd.n1936 gnd.n1934 1.91244
R12479 gnd.n5034 gnd.t261 1.91244
R12480 gnd.n5324 gnd.n5323 1.91244
R12481 gnd.t324 gnd.n3173 1.59378
R12482 gnd.n3352 gnd.t294 1.59378
R12483 gnd.n2614 gnd.t192 1.59378
R12484 gnd.n4569 gnd.t277 1.59378
R12485 gnd.t147 gnd.n2101 1.59378
R12486 gnd.n4936 gnd.t145 1.59378
R12487 gnd.n5011 gnd.t317 1.59378
R12488 gnd.t109 gnd.n2282 1.27512
R12489 gnd.n4517 gnd.n4516 1.27512
R12490 gnd.n4537 gnd.t258 1.27512
R12491 gnd.n4560 gnd.n4559 1.27512
R12492 gnd.n4655 gnd.t226 1.27512
R12493 gnd.n4694 gnd.n4693 1.27512
R12494 gnd.n4716 gnd.n2088 1.27512
R12495 gnd.n4864 gnd.n4863 1.27512
R12496 gnd.n4923 gnd.n1986 1.27512
R12497 gnd.n4892 gnd.t4 1.27512
R12498 gnd.n5032 gnd.n5031 1.27512
R12499 gnd.t141 gnd.n1900 1.27512
R12500 gnd.n5063 gnd.t30 1.27512
R12501 gnd.n5080 gnd.n1882 1.27512
R12502 gnd.n3015 gnd.n3007 1.16414
R12503 gnd.n3831 gnd.n2517 1.16414
R12504 gnd.n3768 gnd.n3761 1.16414
R12505 gnd.n3736 gnd.n3729 1.16414
R12506 gnd.n3704 gnd.n3697 1.16414
R12507 gnd.n3673 gnd.n3666 1.16414
R12508 gnd.n3641 gnd.n3634 1.16414
R12509 gnd.n3609 gnd.n3602 1.16414
R12510 gnd.n3577 gnd.n3570 1.16414
R12511 gnd.n3546 gnd.n3539 1.16414
R12512 gnd.n5485 gnd.n1786 0.970197
R12513 gnd.n6066 gnd.n1318 0.970197
R12514 gnd.n3752 gnd.n3720 0.962709
R12515 gnd.n3784 gnd.n3752 0.962709
R12516 gnd.n3625 gnd.n3593 0.962709
R12517 gnd.n3657 gnd.n3625 0.962709
R12518 gnd.n3261 gnd.t326 0.956468
R12519 gnd.n3426 gnd.t10 0.956468
R12520 gnd.n6306 gnd.t169 0.956468
R12521 gnd.n6299 gnd.t175 0.956468
R12522 gnd.n2350 gnd.t287 0.956468
R12523 gnd.n4385 gnd.t206 0.956468
R12524 gnd.n6062 gnd.n1453 0.956468
R12525 gnd.t222 gnd.n4503 0.956468
R12526 gnd.n5096 gnd.t201 0.956468
R12527 gnd.n5481 gnd.n1791 0.956468
R12528 gnd.n5686 gnd.t190 0.956468
R12529 gnd.n5741 gnd.t177 0.956468
R12530 gnd.n7174 gnd.t159 0.956468
R12531 gnd.t6 gnd.n138 0.956468
R12532 gnd.n2 gnd.n1 0.672012
R12533 gnd.n3 gnd.n2 0.672012
R12534 gnd.n4 gnd.n3 0.672012
R12535 gnd.n5 gnd.n4 0.672012
R12536 gnd.n6 gnd.n5 0.672012
R12537 gnd.n7 gnd.n6 0.672012
R12538 gnd.n9 gnd.n8 0.672012
R12539 gnd.n10 gnd.n9 0.672012
R12540 gnd.n11 gnd.n10 0.672012
R12541 gnd.n12 gnd.n11 0.672012
R12542 gnd.n13 gnd.n12 0.672012
R12543 gnd.n14 gnd.n13 0.672012
R12544 gnd.t80 gnd.n5984 0.637812
R12545 gnd.t64 gnd.n4517 0.637812
R12546 gnd.n4633 gnd.n4632 0.637812
R12547 gnd.n4654 gnd.n4652 0.637812
R12548 gnd.n4663 gnd.t262 0.637812
R12549 gnd.n4783 gnd.n4782 0.637812
R12550 gnd.n4829 gnd.n4828 0.637812
R12551 gnd.t5 gnd.n4954 0.637812
R12552 gnd.n4895 gnd.n4894 0.637812
R12553 gnd.n4994 gnd.n4993 0.637812
R12554 gnd.t33 gnd.n1877 0.637812
R12555 gnd.n5104 gnd.t77 0.637812
R12556 gnd.n2727 gnd.n2726 0.573776
R12557 gnd.n2726 gnd.n2724 0.573776
R12558 gnd.n2724 gnd.n2722 0.573776
R12559 gnd.n2722 gnd.n2720 0.573776
R12560 gnd.n2720 gnd.n2718 0.573776
R12561 gnd.n2692 gnd.n2691 0.573776
R12562 gnd.n2691 gnd.n2689 0.573776
R12563 gnd.n2689 gnd.n2687 0.573776
R12564 gnd.n2687 gnd.n2685 0.573776
R12565 gnd.n2685 gnd.n2683 0.573776
R12566 gnd.n2703 gnd.n2702 0.573776
R12567 gnd.n2702 gnd.n2700 0.573776
R12568 gnd.n2700 gnd.n2698 0.573776
R12569 gnd.n2698 gnd.n2696 0.573776
R12570 gnd.n2696 gnd.n2694 0.573776
R12571 gnd.n2715 gnd.n2714 0.573776
R12572 gnd.n2714 gnd.n2712 0.573776
R12573 gnd.n2712 gnd.n2710 0.573776
R12574 gnd.n2710 gnd.n2708 0.573776
R12575 gnd.n2708 gnd.n2706 0.573776
R12576 gnd.n54 gnd.n52 0.573776
R12577 gnd.n56 gnd.n54 0.573776
R12578 gnd.n58 gnd.n56 0.573776
R12579 gnd.n60 gnd.n58 0.573776
R12580 gnd.n61 gnd.n60 0.573776
R12581 gnd.n19 gnd.n17 0.573776
R12582 gnd.n21 gnd.n19 0.573776
R12583 gnd.n23 gnd.n21 0.573776
R12584 gnd.n25 gnd.n23 0.573776
R12585 gnd.n26 gnd.n25 0.573776
R12586 gnd.n30 gnd.n28 0.573776
R12587 gnd.n32 gnd.n30 0.573776
R12588 gnd.n34 gnd.n32 0.573776
R12589 gnd.n36 gnd.n34 0.573776
R12590 gnd.n37 gnd.n36 0.573776
R12591 gnd.n42 gnd.n40 0.573776
R12592 gnd.n44 gnd.n42 0.573776
R12593 gnd.n46 gnd.n44 0.573776
R12594 gnd.n48 gnd.n46 0.573776
R12595 gnd.n49 gnd.n48 0.573776
R12596 gnd gnd.n0 0.551497
R12597 gnd.n7253 gnd.n7252 0.532512
R12598 gnd.n4053 gnd.n4051 0.532512
R12599 gnd.n236 gnd.n165 0.497451
R12600 gnd.n1290 gnd.n1136 0.497451
R12601 gnd.n5511 gnd.n1613 0.497451
R12602 gnd.n4216 gnd.n4215 0.497451
R12603 gnd.n5297 gnd.n5296 0.489829
R12604 gnd.n2315 gnd.n1149 0.489829
R12605 gnd.n2311 gnd.n1172 0.489829
R12606 gnd.n5877 gnd.n1583 0.489829
R12607 gnd.n3488 gnd.n2521 0.486781
R12608 gnd.n3064 gnd.n3063 0.48678
R12609 gnd.n3805 gnd.n2475 0.480683
R12610 gnd.n3148 gnd.n3147 0.480683
R12611 gnd.n6481 gnd.n6480 0.480683
R12612 gnd.n6902 gnd.n6901 0.480683
R12613 gnd.n7114 gnd.n7113 0.480683
R12614 gnd.n6310 gnd.n6309 0.480683
R12615 gnd.n7346 gnd.n7345 0.470187
R12616 gnd.n7334 gnd.n79 0.4255
R12617 gnd.n4338 gnd.n1018 0.4255
R12618 gnd.n6124 gnd.n1233 0.388379
R12619 gnd.n3765 gnd.n3764 0.388379
R12620 gnd.n3733 gnd.n3732 0.388379
R12621 gnd.n3701 gnd.n3700 0.388379
R12622 gnd.n3670 gnd.n3669 0.388379
R12623 gnd.n3638 gnd.n3637 0.388379
R12624 gnd.n3606 gnd.n3605 0.388379
R12625 gnd.n3574 gnd.n3573 0.388379
R12626 gnd.n3543 gnd.n3542 0.388379
R12627 gnd.n5274 gnd.n5132 0.388379
R12628 gnd.n7346 gnd.n15 0.374463
R12629 gnd.n2576 gnd.t13 0.319156
R12630 gnd.n4278 gnd.t138 0.319156
R12631 gnd.n4332 gnd.t157 0.319156
R12632 gnd.n4316 gnd.t197 0.319156
R12633 gnd.n4307 gnd.t185 0.319156
R12634 gnd.n4447 gnd.t73 0.319156
R12635 gnd.t50 gnd.n5302 0.319156
R12636 gnd.n5806 gnd.t153 0.319156
R12637 gnd.n5798 gnd.t149 0.319156
R12638 gnd.n7144 gnd.t134 0.319156
R12639 gnd.t188 gnd.n98 0.319156
R12640 gnd.n2982 gnd.n2960 0.311721
R12641 gnd.n6188 gnd.n6187 0.302329
R12642 gnd.n5126 gnd.n5125 0.302329
R12643 gnd gnd.n7346 0.295112
R12644 gnd.n7205 gnd.n385 0.293183
R12645 gnd.n4096 gnd.n4014 0.293183
R12646 gnd.n3876 gnd.n3875 0.268793
R12647 gnd.n385 gnd.n384 0.258122
R12648 gnd.n5661 gnd.n5660 0.258122
R12649 gnd.n1351 gnd.n1144 0.258122
R12650 gnd.n4097 gnd.n4096 0.258122
R12651 gnd.n3875 gnd.n3874 0.241354
R12652 gnd.n5576 gnd.n5575 0.229039
R12653 gnd.n5575 gnd.n1785 0.229039
R12654 gnd.n1416 gnd.n1317 0.229039
R12655 gnd.n1416 gnd.n1415 0.229039
R12656 gnd.n3136 gnd.n2935 0.206293
R12657 gnd.n3782 gnd.n3754 0.155672
R12658 gnd.n3775 gnd.n3754 0.155672
R12659 gnd.n3775 gnd.n3774 0.155672
R12660 gnd.n3774 gnd.n3758 0.155672
R12661 gnd.n3767 gnd.n3758 0.155672
R12662 gnd.n3767 gnd.n3766 0.155672
R12663 gnd.n3750 gnd.n3722 0.155672
R12664 gnd.n3743 gnd.n3722 0.155672
R12665 gnd.n3743 gnd.n3742 0.155672
R12666 gnd.n3742 gnd.n3726 0.155672
R12667 gnd.n3735 gnd.n3726 0.155672
R12668 gnd.n3735 gnd.n3734 0.155672
R12669 gnd.n3718 gnd.n3690 0.155672
R12670 gnd.n3711 gnd.n3690 0.155672
R12671 gnd.n3711 gnd.n3710 0.155672
R12672 gnd.n3710 gnd.n3694 0.155672
R12673 gnd.n3703 gnd.n3694 0.155672
R12674 gnd.n3703 gnd.n3702 0.155672
R12675 gnd.n3687 gnd.n3659 0.155672
R12676 gnd.n3680 gnd.n3659 0.155672
R12677 gnd.n3680 gnd.n3679 0.155672
R12678 gnd.n3679 gnd.n3663 0.155672
R12679 gnd.n3672 gnd.n3663 0.155672
R12680 gnd.n3672 gnd.n3671 0.155672
R12681 gnd.n3655 gnd.n3627 0.155672
R12682 gnd.n3648 gnd.n3627 0.155672
R12683 gnd.n3648 gnd.n3647 0.155672
R12684 gnd.n3647 gnd.n3631 0.155672
R12685 gnd.n3640 gnd.n3631 0.155672
R12686 gnd.n3640 gnd.n3639 0.155672
R12687 gnd.n3623 gnd.n3595 0.155672
R12688 gnd.n3616 gnd.n3595 0.155672
R12689 gnd.n3616 gnd.n3615 0.155672
R12690 gnd.n3615 gnd.n3599 0.155672
R12691 gnd.n3608 gnd.n3599 0.155672
R12692 gnd.n3608 gnd.n3607 0.155672
R12693 gnd.n3591 gnd.n3563 0.155672
R12694 gnd.n3584 gnd.n3563 0.155672
R12695 gnd.n3584 gnd.n3583 0.155672
R12696 gnd.n3583 gnd.n3567 0.155672
R12697 gnd.n3576 gnd.n3567 0.155672
R12698 gnd.n3576 gnd.n3575 0.155672
R12699 gnd.n3560 gnd.n3532 0.155672
R12700 gnd.n3553 gnd.n3532 0.155672
R12701 gnd.n3553 gnd.n3552 0.155672
R12702 gnd.n3552 gnd.n3536 0.155672
R12703 gnd.n3545 gnd.n3536 0.155672
R12704 gnd.n3545 gnd.n3544 0.155672
R12705 gnd.n3907 gnd.n2475 0.152939
R12706 gnd.n3907 gnd.n3906 0.152939
R12707 gnd.n3906 gnd.n3905 0.152939
R12708 gnd.n3905 gnd.n2477 0.152939
R12709 gnd.n2478 gnd.n2477 0.152939
R12710 gnd.n2479 gnd.n2478 0.152939
R12711 gnd.n2480 gnd.n2479 0.152939
R12712 gnd.n2481 gnd.n2480 0.152939
R12713 gnd.n2482 gnd.n2481 0.152939
R12714 gnd.n2483 gnd.n2482 0.152939
R12715 gnd.n2484 gnd.n2483 0.152939
R12716 gnd.n2485 gnd.n2484 0.152939
R12717 gnd.n2486 gnd.n2485 0.152939
R12718 gnd.n2487 gnd.n2486 0.152939
R12719 gnd.n3877 gnd.n2487 0.152939
R12720 gnd.n3877 gnd.n3876 0.152939
R12721 gnd.n3149 gnd.n3148 0.152939
R12722 gnd.n3149 gnd.n2853 0.152939
R12723 gnd.n3177 gnd.n2853 0.152939
R12724 gnd.n3178 gnd.n3177 0.152939
R12725 gnd.n3179 gnd.n3178 0.152939
R12726 gnd.n3180 gnd.n3179 0.152939
R12727 gnd.n3180 gnd.n2825 0.152939
R12728 gnd.n3207 gnd.n2825 0.152939
R12729 gnd.n3208 gnd.n3207 0.152939
R12730 gnd.n3209 gnd.n3208 0.152939
R12731 gnd.n3209 gnd.n2803 0.152939
R12732 gnd.n3238 gnd.n2803 0.152939
R12733 gnd.n3239 gnd.n3238 0.152939
R12734 gnd.n3240 gnd.n3239 0.152939
R12735 gnd.n3241 gnd.n3240 0.152939
R12736 gnd.n3243 gnd.n3241 0.152939
R12737 gnd.n3243 gnd.n3242 0.152939
R12738 gnd.n3242 gnd.n2752 0.152939
R12739 gnd.n2753 gnd.n2752 0.152939
R12740 gnd.n2754 gnd.n2753 0.152939
R12741 gnd.n2773 gnd.n2754 0.152939
R12742 gnd.n2774 gnd.n2773 0.152939
R12743 gnd.n2774 gnd.n2672 0.152939
R12744 gnd.n3333 gnd.n2672 0.152939
R12745 gnd.n3334 gnd.n3333 0.152939
R12746 gnd.n3335 gnd.n3334 0.152939
R12747 gnd.n3336 gnd.n3335 0.152939
R12748 gnd.n3336 gnd.n2645 0.152939
R12749 gnd.n3373 gnd.n2645 0.152939
R12750 gnd.n3374 gnd.n3373 0.152939
R12751 gnd.n3375 gnd.n3374 0.152939
R12752 gnd.n3376 gnd.n3375 0.152939
R12753 gnd.n3376 gnd.n2618 0.152939
R12754 gnd.n3418 gnd.n2618 0.152939
R12755 gnd.n3419 gnd.n3418 0.152939
R12756 gnd.n3420 gnd.n3419 0.152939
R12757 gnd.n3421 gnd.n3420 0.152939
R12758 gnd.n3421 gnd.n2590 0.152939
R12759 gnd.n3458 gnd.n2590 0.152939
R12760 gnd.n3459 gnd.n3458 0.152939
R12761 gnd.n3460 gnd.n3459 0.152939
R12762 gnd.n3461 gnd.n3460 0.152939
R12763 gnd.n3461 gnd.n2563 0.152939
R12764 gnd.n3507 gnd.n2563 0.152939
R12765 gnd.n3508 gnd.n3507 0.152939
R12766 gnd.n3509 gnd.n3508 0.152939
R12767 gnd.n3510 gnd.n3509 0.152939
R12768 gnd.n3510 gnd.n2536 0.152939
R12769 gnd.n3801 gnd.n2536 0.152939
R12770 gnd.n3802 gnd.n3801 0.152939
R12771 gnd.n3803 gnd.n3802 0.152939
R12772 gnd.n3804 gnd.n3803 0.152939
R12773 gnd.n3805 gnd.n3804 0.152939
R12774 gnd.n3147 gnd.n2877 0.152939
R12775 gnd.n2898 gnd.n2877 0.152939
R12776 gnd.n2899 gnd.n2898 0.152939
R12777 gnd.n2905 gnd.n2899 0.152939
R12778 gnd.n2906 gnd.n2905 0.152939
R12779 gnd.n2907 gnd.n2906 0.152939
R12780 gnd.n2907 gnd.n2896 0.152939
R12781 gnd.n2915 gnd.n2896 0.152939
R12782 gnd.n2916 gnd.n2915 0.152939
R12783 gnd.n2917 gnd.n2916 0.152939
R12784 gnd.n2917 gnd.n2894 0.152939
R12785 gnd.n2925 gnd.n2894 0.152939
R12786 gnd.n2926 gnd.n2925 0.152939
R12787 gnd.n2927 gnd.n2926 0.152939
R12788 gnd.n2927 gnd.n2892 0.152939
R12789 gnd.n2935 gnd.n2892 0.152939
R12790 gnd.n3874 gnd.n2492 0.152939
R12791 gnd.n2494 gnd.n2492 0.152939
R12792 gnd.n2495 gnd.n2494 0.152939
R12793 gnd.n2496 gnd.n2495 0.152939
R12794 gnd.n2497 gnd.n2496 0.152939
R12795 gnd.n2498 gnd.n2497 0.152939
R12796 gnd.n2499 gnd.n2498 0.152939
R12797 gnd.n2500 gnd.n2499 0.152939
R12798 gnd.n2501 gnd.n2500 0.152939
R12799 gnd.n2502 gnd.n2501 0.152939
R12800 gnd.n2503 gnd.n2502 0.152939
R12801 gnd.n2504 gnd.n2503 0.152939
R12802 gnd.n2505 gnd.n2504 0.152939
R12803 gnd.n2506 gnd.n2505 0.152939
R12804 gnd.n2507 gnd.n2506 0.152939
R12805 gnd.n2508 gnd.n2507 0.152939
R12806 gnd.n2509 gnd.n2508 0.152939
R12807 gnd.n2510 gnd.n2509 0.152939
R12808 gnd.n2511 gnd.n2510 0.152939
R12809 gnd.n2512 gnd.n2511 0.152939
R12810 gnd.n2513 gnd.n2512 0.152939
R12811 gnd.n2514 gnd.n2513 0.152939
R12812 gnd.n2518 gnd.n2514 0.152939
R12813 gnd.n2519 gnd.n2518 0.152939
R12814 gnd.n2520 gnd.n2519 0.152939
R12815 gnd.n2521 gnd.n2520 0.152939
R12816 gnd.n3310 gnd.n3309 0.152939
R12817 gnd.n3311 gnd.n3310 0.152939
R12818 gnd.n3312 gnd.n3311 0.152939
R12819 gnd.n3313 gnd.n3312 0.152939
R12820 gnd.n3314 gnd.n3313 0.152939
R12821 gnd.n3315 gnd.n3314 0.152939
R12822 gnd.n3315 gnd.n2626 0.152939
R12823 gnd.n3394 gnd.n2626 0.152939
R12824 gnd.n3395 gnd.n3394 0.152939
R12825 gnd.n3396 gnd.n3395 0.152939
R12826 gnd.n3397 gnd.n3396 0.152939
R12827 gnd.n3398 gnd.n3397 0.152939
R12828 gnd.n3399 gnd.n3398 0.152939
R12829 gnd.n3400 gnd.n3399 0.152939
R12830 gnd.n3401 gnd.n3400 0.152939
R12831 gnd.n3402 gnd.n3401 0.152939
R12832 gnd.n3402 gnd.n2570 0.152939
R12833 gnd.n3479 gnd.n2570 0.152939
R12834 gnd.n3480 gnd.n3479 0.152939
R12835 gnd.n3481 gnd.n3480 0.152939
R12836 gnd.n3482 gnd.n3481 0.152939
R12837 gnd.n3483 gnd.n3482 0.152939
R12838 gnd.n3484 gnd.n3483 0.152939
R12839 gnd.n3485 gnd.n3484 0.152939
R12840 gnd.n3486 gnd.n3485 0.152939
R12841 gnd.n3487 gnd.n3486 0.152939
R12842 gnd.n3489 gnd.n3487 0.152939
R12843 gnd.n3489 gnd.n3488 0.152939
R12844 gnd.n3065 gnd.n3064 0.152939
R12845 gnd.n3065 gnd.n2955 0.152939
R12846 gnd.n3080 gnd.n2955 0.152939
R12847 gnd.n3081 gnd.n3080 0.152939
R12848 gnd.n3082 gnd.n3081 0.152939
R12849 gnd.n3082 gnd.n2943 0.152939
R12850 gnd.n3096 gnd.n2943 0.152939
R12851 gnd.n3097 gnd.n3096 0.152939
R12852 gnd.n3098 gnd.n3097 0.152939
R12853 gnd.n3099 gnd.n3098 0.152939
R12854 gnd.n3100 gnd.n3099 0.152939
R12855 gnd.n3101 gnd.n3100 0.152939
R12856 gnd.n3102 gnd.n3101 0.152939
R12857 gnd.n3103 gnd.n3102 0.152939
R12858 gnd.n3104 gnd.n3103 0.152939
R12859 gnd.n3105 gnd.n3104 0.152939
R12860 gnd.n3106 gnd.n3105 0.152939
R12861 gnd.n3107 gnd.n3106 0.152939
R12862 gnd.n3108 gnd.n3107 0.152939
R12863 gnd.n3109 gnd.n3108 0.152939
R12864 gnd.n3110 gnd.n3109 0.152939
R12865 gnd.n3110 gnd.n2809 0.152939
R12866 gnd.n3227 gnd.n2809 0.152939
R12867 gnd.n3228 gnd.n3227 0.152939
R12868 gnd.n3229 gnd.n3228 0.152939
R12869 gnd.n3230 gnd.n3229 0.152939
R12870 gnd.n3230 gnd.n2731 0.152939
R12871 gnd.n3307 gnd.n2731 0.152939
R12872 gnd.n2983 gnd.n2982 0.152939
R12873 gnd.n2984 gnd.n2983 0.152939
R12874 gnd.n2985 gnd.n2984 0.152939
R12875 gnd.n2986 gnd.n2985 0.152939
R12876 gnd.n2987 gnd.n2986 0.152939
R12877 gnd.n2988 gnd.n2987 0.152939
R12878 gnd.n2989 gnd.n2988 0.152939
R12879 gnd.n2990 gnd.n2989 0.152939
R12880 gnd.n2991 gnd.n2990 0.152939
R12881 gnd.n2992 gnd.n2991 0.152939
R12882 gnd.n2993 gnd.n2992 0.152939
R12883 gnd.n2994 gnd.n2993 0.152939
R12884 gnd.n2995 gnd.n2994 0.152939
R12885 gnd.n2996 gnd.n2995 0.152939
R12886 gnd.n2997 gnd.n2996 0.152939
R12887 gnd.n2998 gnd.n2997 0.152939
R12888 gnd.n2999 gnd.n2998 0.152939
R12889 gnd.n3000 gnd.n2999 0.152939
R12890 gnd.n3001 gnd.n3000 0.152939
R12891 gnd.n3002 gnd.n3001 0.152939
R12892 gnd.n3003 gnd.n3002 0.152939
R12893 gnd.n3004 gnd.n3003 0.152939
R12894 gnd.n3008 gnd.n3004 0.152939
R12895 gnd.n3009 gnd.n3008 0.152939
R12896 gnd.n3009 gnd.n2966 0.152939
R12897 gnd.n3063 gnd.n2966 0.152939
R12898 gnd.n6481 gnd.n792 0.152939
R12899 gnd.n6489 gnd.n792 0.152939
R12900 gnd.n6490 gnd.n6489 0.152939
R12901 gnd.n6491 gnd.n6490 0.152939
R12902 gnd.n6491 gnd.n786 0.152939
R12903 gnd.n6499 gnd.n786 0.152939
R12904 gnd.n6500 gnd.n6499 0.152939
R12905 gnd.n6501 gnd.n6500 0.152939
R12906 gnd.n6501 gnd.n780 0.152939
R12907 gnd.n6509 gnd.n780 0.152939
R12908 gnd.n6510 gnd.n6509 0.152939
R12909 gnd.n6511 gnd.n6510 0.152939
R12910 gnd.n6511 gnd.n774 0.152939
R12911 gnd.n6519 gnd.n774 0.152939
R12912 gnd.n6520 gnd.n6519 0.152939
R12913 gnd.n6521 gnd.n6520 0.152939
R12914 gnd.n6521 gnd.n768 0.152939
R12915 gnd.n6529 gnd.n768 0.152939
R12916 gnd.n6530 gnd.n6529 0.152939
R12917 gnd.n6531 gnd.n6530 0.152939
R12918 gnd.n6531 gnd.n762 0.152939
R12919 gnd.n6539 gnd.n762 0.152939
R12920 gnd.n6540 gnd.n6539 0.152939
R12921 gnd.n6541 gnd.n6540 0.152939
R12922 gnd.n6541 gnd.n756 0.152939
R12923 gnd.n6549 gnd.n756 0.152939
R12924 gnd.n6550 gnd.n6549 0.152939
R12925 gnd.n6551 gnd.n6550 0.152939
R12926 gnd.n6551 gnd.n750 0.152939
R12927 gnd.n6559 gnd.n750 0.152939
R12928 gnd.n6560 gnd.n6559 0.152939
R12929 gnd.n6561 gnd.n6560 0.152939
R12930 gnd.n6561 gnd.n744 0.152939
R12931 gnd.n6569 gnd.n744 0.152939
R12932 gnd.n6570 gnd.n6569 0.152939
R12933 gnd.n6571 gnd.n6570 0.152939
R12934 gnd.n6571 gnd.n738 0.152939
R12935 gnd.n6579 gnd.n738 0.152939
R12936 gnd.n6580 gnd.n6579 0.152939
R12937 gnd.n6581 gnd.n6580 0.152939
R12938 gnd.n6581 gnd.n732 0.152939
R12939 gnd.n6589 gnd.n732 0.152939
R12940 gnd.n6590 gnd.n6589 0.152939
R12941 gnd.n6591 gnd.n6590 0.152939
R12942 gnd.n6591 gnd.n726 0.152939
R12943 gnd.n6599 gnd.n726 0.152939
R12944 gnd.n6600 gnd.n6599 0.152939
R12945 gnd.n6601 gnd.n6600 0.152939
R12946 gnd.n6601 gnd.n720 0.152939
R12947 gnd.n6609 gnd.n720 0.152939
R12948 gnd.n6610 gnd.n6609 0.152939
R12949 gnd.n6611 gnd.n6610 0.152939
R12950 gnd.n6611 gnd.n714 0.152939
R12951 gnd.n6619 gnd.n714 0.152939
R12952 gnd.n6620 gnd.n6619 0.152939
R12953 gnd.n6621 gnd.n6620 0.152939
R12954 gnd.n6621 gnd.n708 0.152939
R12955 gnd.n6629 gnd.n708 0.152939
R12956 gnd.n6630 gnd.n6629 0.152939
R12957 gnd.n6631 gnd.n6630 0.152939
R12958 gnd.n6631 gnd.n702 0.152939
R12959 gnd.n6639 gnd.n702 0.152939
R12960 gnd.n6640 gnd.n6639 0.152939
R12961 gnd.n6641 gnd.n6640 0.152939
R12962 gnd.n6641 gnd.n696 0.152939
R12963 gnd.n6649 gnd.n696 0.152939
R12964 gnd.n6650 gnd.n6649 0.152939
R12965 gnd.n6651 gnd.n6650 0.152939
R12966 gnd.n6651 gnd.n690 0.152939
R12967 gnd.n6659 gnd.n690 0.152939
R12968 gnd.n6660 gnd.n6659 0.152939
R12969 gnd.n6661 gnd.n6660 0.152939
R12970 gnd.n6661 gnd.n684 0.152939
R12971 gnd.n6669 gnd.n684 0.152939
R12972 gnd.n6670 gnd.n6669 0.152939
R12973 gnd.n6671 gnd.n6670 0.152939
R12974 gnd.n6671 gnd.n678 0.152939
R12975 gnd.n6679 gnd.n678 0.152939
R12976 gnd.n6680 gnd.n6679 0.152939
R12977 gnd.n6681 gnd.n6680 0.152939
R12978 gnd.n6681 gnd.n672 0.152939
R12979 gnd.n6689 gnd.n672 0.152939
R12980 gnd.n6690 gnd.n6689 0.152939
R12981 gnd.n6691 gnd.n6690 0.152939
R12982 gnd.n6691 gnd.n666 0.152939
R12983 gnd.n6699 gnd.n666 0.152939
R12984 gnd.n6700 gnd.n6699 0.152939
R12985 gnd.n6701 gnd.n6700 0.152939
R12986 gnd.n6701 gnd.n660 0.152939
R12987 gnd.n6709 gnd.n660 0.152939
R12988 gnd.n6710 gnd.n6709 0.152939
R12989 gnd.n6711 gnd.n6710 0.152939
R12990 gnd.n6711 gnd.n654 0.152939
R12991 gnd.n6719 gnd.n654 0.152939
R12992 gnd.n6720 gnd.n6719 0.152939
R12993 gnd.n6721 gnd.n6720 0.152939
R12994 gnd.n6721 gnd.n648 0.152939
R12995 gnd.n6729 gnd.n648 0.152939
R12996 gnd.n6730 gnd.n6729 0.152939
R12997 gnd.n6731 gnd.n6730 0.152939
R12998 gnd.n6731 gnd.n642 0.152939
R12999 gnd.n6739 gnd.n642 0.152939
R13000 gnd.n6740 gnd.n6739 0.152939
R13001 gnd.n6741 gnd.n6740 0.152939
R13002 gnd.n6741 gnd.n636 0.152939
R13003 gnd.n6749 gnd.n636 0.152939
R13004 gnd.n6750 gnd.n6749 0.152939
R13005 gnd.n6751 gnd.n6750 0.152939
R13006 gnd.n6751 gnd.n630 0.152939
R13007 gnd.n6759 gnd.n630 0.152939
R13008 gnd.n6760 gnd.n6759 0.152939
R13009 gnd.n6761 gnd.n6760 0.152939
R13010 gnd.n6761 gnd.n624 0.152939
R13011 gnd.n6769 gnd.n624 0.152939
R13012 gnd.n6770 gnd.n6769 0.152939
R13013 gnd.n6771 gnd.n6770 0.152939
R13014 gnd.n6771 gnd.n618 0.152939
R13015 gnd.n6779 gnd.n618 0.152939
R13016 gnd.n6780 gnd.n6779 0.152939
R13017 gnd.n6781 gnd.n6780 0.152939
R13018 gnd.n6781 gnd.n612 0.152939
R13019 gnd.n6789 gnd.n612 0.152939
R13020 gnd.n6790 gnd.n6789 0.152939
R13021 gnd.n6791 gnd.n6790 0.152939
R13022 gnd.n6791 gnd.n606 0.152939
R13023 gnd.n6799 gnd.n606 0.152939
R13024 gnd.n6800 gnd.n6799 0.152939
R13025 gnd.n6801 gnd.n6800 0.152939
R13026 gnd.n6801 gnd.n600 0.152939
R13027 gnd.n6809 gnd.n600 0.152939
R13028 gnd.n6810 gnd.n6809 0.152939
R13029 gnd.n6811 gnd.n6810 0.152939
R13030 gnd.n6811 gnd.n594 0.152939
R13031 gnd.n6819 gnd.n594 0.152939
R13032 gnd.n6820 gnd.n6819 0.152939
R13033 gnd.n6821 gnd.n6820 0.152939
R13034 gnd.n6821 gnd.n588 0.152939
R13035 gnd.n6829 gnd.n588 0.152939
R13036 gnd.n6830 gnd.n6829 0.152939
R13037 gnd.n6831 gnd.n6830 0.152939
R13038 gnd.n6831 gnd.n582 0.152939
R13039 gnd.n6839 gnd.n582 0.152939
R13040 gnd.n6840 gnd.n6839 0.152939
R13041 gnd.n6841 gnd.n6840 0.152939
R13042 gnd.n6841 gnd.n576 0.152939
R13043 gnd.n6849 gnd.n576 0.152939
R13044 gnd.n6850 gnd.n6849 0.152939
R13045 gnd.n6851 gnd.n6850 0.152939
R13046 gnd.n6851 gnd.n570 0.152939
R13047 gnd.n6859 gnd.n570 0.152939
R13048 gnd.n6860 gnd.n6859 0.152939
R13049 gnd.n6861 gnd.n6860 0.152939
R13050 gnd.n6861 gnd.n564 0.152939
R13051 gnd.n6869 gnd.n564 0.152939
R13052 gnd.n6870 gnd.n6869 0.152939
R13053 gnd.n6871 gnd.n6870 0.152939
R13054 gnd.n6871 gnd.n558 0.152939
R13055 gnd.n6879 gnd.n558 0.152939
R13056 gnd.n6880 gnd.n6879 0.152939
R13057 gnd.n6881 gnd.n6880 0.152939
R13058 gnd.n6881 gnd.n552 0.152939
R13059 gnd.n6889 gnd.n552 0.152939
R13060 gnd.n6890 gnd.n6889 0.152939
R13061 gnd.n6892 gnd.n6890 0.152939
R13062 gnd.n6892 gnd.n6891 0.152939
R13063 gnd.n6891 gnd.n546 0.152939
R13064 gnd.n6901 gnd.n546 0.152939
R13065 gnd.n6902 gnd.n541 0.152939
R13066 gnd.n6910 gnd.n541 0.152939
R13067 gnd.n6911 gnd.n6910 0.152939
R13068 gnd.n6912 gnd.n6911 0.152939
R13069 gnd.n6912 gnd.n535 0.152939
R13070 gnd.n6920 gnd.n535 0.152939
R13071 gnd.n6921 gnd.n6920 0.152939
R13072 gnd.n6922 gnd.n6921 0.152939
R13073 gnd.n6922 gnd.n529 0.152939
R13074 gnd.n6930 gnd.n529 0.152939
R13075 gnd.n6931 gnd.n6930 0.152939
R13076 gnd.n6932 gnd.n6931 0.152939
R13077 gnd.n6932 gnd.n523 0.152939
R13078 gnd.n6940 gnd.n523 0.152939
R13079 gnd.n6941 gnd.n6940 0.152939
R13080 gnd.n6942 gnd.n6941 0.152939
R13081 gnd.n6942 gnd.n517 0.152939
R13082 gnd.n6950 gnd.n517 0.152939
R13083 gnd.n6951 gnd.n6950 0.152939
R13084 gnd.n6952 gnd.n6951 0.152939
R13085 gnd.n6952 gnd.n511 0.152939
R13086 gnd.n6960 gnd.n511 0.152939
R13087 gnd.n6961 gnd.n6960 0.152939
R13088 gnd.n6962 gnd.n6961 0.152939
R13089 gnd.n6962 gnd.n505 0.152939
R13090 gnd.n6970 gnd.n505 0.152939
R13091 gnd.n6971 gnd.n6970 0.152939
R13092 gnd.n6972 gnd.n6971 0.152939
R13093 gnd.n6972 gnd.n499 0.152939
R13094 gnd.n6980 gnd.n499 0.152939
R13095 gnd.n6981 gnd.n6980 0.152939
R13096 gnd.n6982 gnd.n6981 0.152939
R13097 gnd.n6982 gnd.n493 0.152939
R13098 gnd.n6990 gnd.n493 0.152939
R13099 gnd.n6991 gnd.n6990 0.152939
R13100 gnd.n6992 gnd.n6991 0.152939
R13101 gnd.n6992 gnd.n487 0.152939
R13102 gnd.n7000 gnd.n487 0.152939
R13103 gnd.n7001 gnd.n7000 0.152939
R13104 gnd.n7002 gnd.n7001 0.152939
R13105 gnd.n7002 gnd.n481 0.152939
R13106 gnd.n7010 gnd.n481 0.152939
R13107 gnd.n7011 gnd.n7010 0.152939
R13108 gnd.n7012 gnd.n7011 0.152939
R13109 gnd.n7012 gnd.n475 0.152939
R13110 gnd.n7020 gnd.n475 0.152939
R13111 gnd.n7021 gnd.n7020 0.152939
R13112 gnd.n7022 gnd.n7021 0.152939
R13113 gnd.n7022 gnd.n469 0.152939
R13114 gnd.n7030 gnd.n469 0.152939
R13115 gnd.n7031 gnd.n7030 0.152939
R13116 gnd.n7032 gnd.n7031 0.152939
R13117 gnd.n7032 gnd.n463 0.152939
R13118 gnd.n7040 gnd.n463 0.152939
R13119 gnd.n7041 gnd.n7040 0.152939
R13120 gnd.n7042 gnd.n7041 0.152939
R13121 gnd.n7042 gnd.n457 0.152939
R13122 gnd.n7050 gnd.n457 0.152939
R13123 gnd.n7051 gnd.n7050 0.152939
R13124 gnd.n7052 gnd.n7051 0.152939
R13125 gnd.n7052 gnd.n451 0.152939
R13126 gnd.n7060 gnd.n451 0.152939
R13127 gnd.n7061 gnd.n7060 0.152939
R13128 gnd.n7062 gnd.n7061 0.152939
R13129 gnd.n7062 gnd.n445 0.152939
R13130 gnd.n7070 gnd.n445 0.152939
R13131 gnd.n7071 gnd.n7070 0.152939
R13132 gnd.n7072 gnd.n7071 0.152939
R13133 gnd.n7072 gnd.n439 0.152939
R13134 gnd.n7080 gnd.n439 0.152939
R13135 gnd.n7081 gnd.n7080 0.152939
R13136 gnd.n7082 gnd.n7081 0.152939
R13137 gnd.n7082 gnd.n433 0.152939
R13138 gnd.n7090 gnd.n433 0.152939
R13139 gnd.n7091 gnd.n7090 0.152939
R13140 gnd.n7092 gnd.n7091 0.152939
R13141 gnd.n7092 gnd.n427 0.152939
R13142 gnd.n7100 gnd.n427 0.152939
R13143 gnd.n7101 gnd.n7100 0.152939
R13144 gnd.n7102 gnd.n7101 0.152939
R13145 gnd.n7102 gnd.n421 0.152939
R13146 gnd.n7111 gnd.n421 0.152939
R13147 gnd.n7112 gnd.n7111 0.152939
R13148 gnd.n7114 gnd.n7112 0.152939
R13149 gnd.n408 gnd.n405 0.152939
R13150 gnd.n409 gnd.n408 0.152939
R13151 gnd.n410 gnd.n409 0.152939
R13152 gnd.n411 gnd.n410 0.152939
R13153 gnd.n414 gnd.n411 0.152939
R13154 gnd.n415 gnd.n414 0.152939
R13155 gnd.n416 gnd.n415 0.152939
R13156 gnd.n417 gnd.n416 0.152939
R13157 gnd.n7113 gnd.n417 0.152939
R13158 gnd.n7334 gnd.n77 0.152939
R13159 gnd.n103 gnd.n77 0.152939
R13160 gnd.n104 gnd.n103 0.152939
R13161 gnd.n105 gnd.n104 0.152939
R13162 gnd.n122 gnd.n105 0.152939
R13163 gnd.n123 gnd.n122 0.152939
R13164 gnd.n124 gnd.n123 0.152939
R13165 gnd.n125 gnd.n124 0.152939
R13166 gnd.n143 gnd.n125 0.152939
R13167 gnd.n144 gnd.n143 0.152939
R13168 gnd.n145 gnd.n144 0.152939
R13169 gnd.n146 gnd.n145 0.152939
R13170 gnd.n162 gnd.n146 0.152939
R13171 gnd.n163 gnd.n162 0.152939
R13172 gnd.n164 gnd.n163 0.152939
R13173 gnd.n165 gnd.n164 0.152939
R13174 gnd.n7343 gnd.n65 0.152939
R13175 gnd.n397 gnd.n65 0.152939
R13176 gnd.n7147 gnd.n397 0.152939
R13177 gnd.n7148 gnd.n7147 0.152939
R13178 gnd.n7149 gnd.n7148 0.152939
R13179 gnd.n7149 gnd.n393 0.152939
R13180 gnd.n7162 gnd.n393 0.152939
R13181 gnd.n7163 gnd.n7162 0.152939
R13182 gnd.n7164 gnd.n7163 0.152939
R13183 gnd.n7164 gnd.n388 0.152939
R13184 gnd.n7177 gnd.n388 0.152939
R13185 gnd.n7178 gnd.n7177 0.152939
R13186 gnd.n7179 gnd.n7178 0.152939
R13187 gnd.n7180 gnd.n7179 0.152939
R13188 gnd.n7181 gnd.n7180 0.152939
R13189 gnd.n7182 gnd.n7181 0.152939
R13190 gnd.n7183 gnd.n7182 0.152939
R13191 gnd.n7184 gnd.n7183 0.152939
R13192 gnd.n7185 gnd.n7184 0.152939
R13193 gnd.n7253 gnd.n7185 0.152939
R13194 gnd.n7205 gnd.n7204 0.152939
R13195 gnd.n7213 gnd.n7204 0.152939
R13196 gnd.n7214 gnd.n7213 0.152939
R13197 gnd.n7215 gnd.n7214 0.152939
R13198 gnd.n7215 gnd.n7200 0.152939
R13199 gnd.n7223 gnd.n7200 0.152939
R13200 gnd.n7224 gnd.n7223 0.152939
R13201 gnd.n7225 gnd.n7224 0.152939
R13202 gnd.n7225 gnd.n7196 0.152939
R13203 gnd.n7233 gnd.n7196 0.152939
R13204 gnd.n7234 gnd.n7233 0.152939
R13205 gnd.n7235 gnd.n7234 0.152939
R13206 gnd.n7235 gnd.n7192 0.152939
R13207 gnd.n7243 gnd.n7192 0.152939
R13208 gnd.n7244 gnd.n7243 0.152939
R13209 gnd.n7245 gnd.n7244 0.152939
R13210 gnd.n7245 gnd.n7186 0.152939
R13211 gnd.n7252 gnd.n7186 0.152939
R13212 gnd.n236 gnd.n235 0.152939
R13213 gnd.n244 gnd.n235 0.152939
R13214 gnd.n245 gnd.n244 0.152939
R13215 gnd.n246 gnd.n245 0.152939
R13216 gnd.n246 gnd.n231 0.152939
R13217 gnd.n254 gnd.n231 0.152939
R13218 gnd.n255 gnd.n254 0.152939
R13219 gnd.n256 gnd.n255 0.152939
R13220 gnd.n256 gnd.n227 0.152939
R13221 gnd.n264 gnd.n227 0.152939
R13222 gnd.n265 gnd.n264 0.152939
R13223 gnd.n266 gnd.n265 0.152939
R13224 gnd.n266 gnd.n223 0.152939
R13225 gnd.n275 gnd.n223 0.152939
R13226 gnd.n276 gnd.n275 0.152939
R13227 gnd.n277 gnd.n276 0.152939
R13228 gnd.n277 gnd.n217 0.152939
R13229 gnd.n285 gnd.n217 0.152939
R13230 gnd.n286 gnd.n285 0.152939
R13231 gnd.n287 gnd.n286 0.152939
R13232 gnd.n287 gnd.n213 0.152939
R13233 gnd.n295 gnd.n213 0.152939
R13234 gnd.n296 gnd.n295 0.152939
R13235 gnd.n297 gnd.n296 0.152939
R13236 gnd.n297 gnd.n209 0.152939
R13237 gnd.n305 gnd.n209 0.152939
R13238 gnd.n306 gnd.n305 0.152939
R13239 gnd.n307 gnd.n306 0.152939
R13240 gnd.n307 gnd.n205 0.152939
R13241 gnd.n315 gnd.n205 0.152939
R13242 gnd.n316 gnd.n315 0.152939
R13243 gnd.n317 gnd.n316 0.152939
R13244 gnd.n317 gnd.n201 0.152939
R13245 gnd.n325 gnd.n201 0.152939
R13246 gnd.n326 gnd.n325 0.152939
R13247 gnd.n327 gnd.n326 0.152939
R13248 gnd.n327 gnd.n195 0.152939
R13249 gnd.n335 gnd.n195 0.152939
R13250 gnd.n336 gnd.n335 0.152939
R13251 gnd.n337 gnd.n336 0.152939
R13252 gnd.n337 gnd.n191 0.152939
R13253 gnd.n345 gnd.n191 0.152939
R13254 gnd.n346 gnd.n345 0.152939
R13255 gnd.n347 gnd.n346 0.152939
R13256 gnd.n347 gnd.n187 0.152939
R13257 gnd.n355 gnd.n187 0.152939
R13258 gnd.n356 gnd.n355 0.152939
R13259 gnd.n357 gnd.n356 0.152939
R13260 gnd.n357 gnd.n183 0.152939
R13261 gnd.n365 gnd.n183 0.152939
R13262 gnd.n366 gnd.n365 0.152939
R13263 gnd.n367 gnd.n366 0.152939
R13264 gnd.n367 gnd.n179 0.152939
R13265 gnd.n375 gnd.n179 0.152939
R13266 gnd.n376 gnd.n375 0.152939
R13267 gnd.n377 gnd.n376 0.152939
R13268 gnd.n377 gnd.n173 0.152939
R13269 gnd.n384 gnd.n173 0.152939
R13270 gnd.n5512 gnd.n5511 0.152939
R13271 gnd.n5512 gnd.n5508 0.152939
R13272 gnd.n5520 gnd.n5508 0.152939
R13273 gnd.n5521 gnd.n5520 0.152939
R13274 gnd.n5522 gnd.n5521 0.152939
R13275 gnd.n5522 gnd.n5504 0.152939
R13276 gnd.n5530 gnd.n5504 0.152939
R13277 gnd.n5531 gnd.n5530 0.152939
R13278 gnd.n5532 gnd.n5531 0.152939
R13279 gnd.n5532 gnd.n5500 0.152939
R13280 gnd.n5540 gnd.n5500 0.152939
R13281 gnd.n5541 gnd.n5540 0.152939
R13282 gnd.n5542 gnd.n5541 0.152939
R13283 gnd.n5542 gnd.n5496 0.152939
R13284 gnd.n5550 gnd.n5496 0.152939
R13285 gnd.n5551 gnd.n5550 0.152939
R13286 gnd.n5552 gnd.n5551 0.152939
R13287 gnd.n5552 gnd.n5492 0.152939
R13288 gnd.n5563 gnd.n5492 0.152939
R13289 gnd.n5564 gnd.n5563 0.152939
R13290 gnd.n5565 gnd.n5564 0.152939
R13291 gnd.n5565 gnd.n5488 0.152939
R13292 gnd.n5573 gnd.n5488 0.152939
R13293 gnd.n5574 gnd.n5573 0.152939
R13294 gnd.n5576 gnd.n5574 0.152939
R13295 gnd.n5586 gnd.n1785 0.152939
R13296 gnd.n5587 gnd.n5586 0.152939
R13297 gnd.n5588 gnd.n5587 0.152939
R13298 gnd.n5588 gnd.n1781 0.152939
R13299 gnd.n5596 gnd.n1781 0.152939
R13300 gnd.n5597 gnd.n5596 0.152939
R13301 gnd.n5598 gnd.n5597 0.152939
R13302 gnd.n5598 gnd.n1777 0.152939
R13303 gnd.n5608 gnd.n1777 0.152939
R13304 gnd.n5609 gnd.n5608 0.152939
R13305 gnd.n5610 gnd.n5609 0.152939
R13306 gnd.n5610 gnd.n1773 0.152939
R13307 gnd.n5618 gnd.n1773 0.152939
R13308 gnd.n5619 gnd.n5618 0.152939
R13309 gnd.n5620 gnd.n5619 0.152939
R13310 gnd.n5620 gnd.n1769 0.152939
R13311 gnd.n5628 gnd.n1769 0.152939
R13312 gnd.n5629 gnd.n5628 0.152939
R13313 gnd.n5630 gnd.n5629 0.152939
R13314 gnd.n5630 gnd.n1765 0.152939
R13315 gnd.n5638 gnd.n1765 0.152939
R13316 gnd.n5639 gnd.n5638 0.152939
R13317 gnd.n5640 gnd.n5639 0.152939
R13318 gnd.n5640 gnd.n1761 0.152939
R13319 gnd.n5648 gnd.n1761 0.152939
R13320 gnd.n5649 gnd.n5648 0.152939
R13321 gnd.n5651 gnd.n5649 0.152939
R13322 gnd.n5651 gnd.n5650 0.152939
R13323 gnd.n5650 gnd.n1754 0.152939
R13324 gnd.n5660 gnd.n1754 0.152939
R13325 gnd.n1614 gnd.n1613 0.152939
R13326 gnd.n1615 gnd.n1614 0.152939
R13327 gnd.n1635 gnd.n1615 0.152939
R13328 gnd.n1636 gnd.n1635 0.152939
R13329 gnd.n1637 gnd.n1636 0.152939
R13330 gnd.n1638 gnd.n1637 0.152939
R13331 gnd.n1655 gnd.n1638 0.152939
R13332 gnd.n1656 gnd.n1655 0.152939
R13333 gnd.n1657 gnd.n1656 0.152939
R13334 gnd.n1658 gnd.n1657 0.152939
R13335 gnd.n1675 gnd.n1658 0.152939
R13336 gnd.n1676 gnd.n1675 0.152939
R13337 gnd.n1677 gnd.n1676 0.152939
R13338 gnd.n1678 gnd.n1677 0.152939
R13339 gnd.n1678 gnd.n78 0.152939
R13340 gnd.n7334 gnd.n78 0.152939
R13341 gnd.n4340 gnd.n4339 0.152939
R13342 gnd.n4341 gnd.n4340 0.152939
R13343 gnd.n4342 gnd.n4341 0.152939
R13344 gnd.n4345 gnd.n4342 0.152939
R13345 gnd.n4346 gnd.n4345 0.152939
R13346 gnd.n4347 gnd.n4346 0.152939
R13347 gnd.n4348 gnd.n4347 0.152939
R13348 gnd.n4349 gnd.n4348 0.152939
R13349 gnd.n4349 gnd.n2336 0.152939
R13350 gnd.n4414 gnd.n2336 0.152939
R13351 gnd.n4415 gnd.n4414 0.152939
R13352 gnd.n4416 gnd.n4415 0.152939
R13353 gnd.n4416 gnd.n2332 0.152939
R13354 gnd.n4422 gnd.n2332 0.152939
R13355 gnd.n4423 gnd.n4422 0.152939
R13356 gnd.n4424 gnd.n4423 0.152939
R13357 gnd.n4424 gnd.n2328 0.152939
R13358 gnd.n4430 gnd.n2328 0.152939
R13359 gnd.n4431 gnd.n4430 0.152939
R13360 gnd.n4432 gnd.n4431 0.152939
R13361 gnd.n4432 gnd.n2323 0.152939
R13362 gnd.n4440 gnd.n2323 0.152939
R13363 gnd.n4441 gnd.n4440 0.152939
R13364 gnd.n4442 gnd.n4441 0.152939
R13365 gnd.n4443 gnd.n4442 0.152939
R13366 gnd.n4443 gnd.n2295 0.152939
R13367 gnd.n4472 gnd.n2295 0.152939
R13368 gnd.n4473 gnd.n4472 0.152939
R13369 gnd.n4474 gnd.n4473 0.152939
R13370 gnd.n4476 gnd.n4474 0.152939
R13371 gnd.n4476 gnd.n4475 0.152939
R13372 gnd.n4475 gnd.n1485 0.152939
R13373 gnd.n1486 gnd.n1485 0.152939
R13374 gnd.n1487 gnd.n1486 0.152939
R13375 gnd.n4512 gnd.n1487 0.152939
R13376 gnd.n4513 gnd.n4512 0.152939
R13377 gnd.n4513 gnd.n2169 0.152939
R13378 gnd.n4554 gnd.n2169 0.152939
R13379 gnd.n4555 gnd.n4554 0.152939
R13380 gnd.n4556 gnd.n4555 0.152939
R13381 gnd.n4556 gnd.n2151 0.152939
R13382 gnd.n4596 gnd.n2151 0.152939
R13383 gnd.n4597 gnd.n4596 0.152939
R13384 gnd.n4598 gnd.n4597 0.152939
R13385 gnd.n4599 gnd.n4598 0.152939
R13386 gnd.n4599 gnd.n2125 0.152939
R13387 gnd.n4658 gnd.n2125 0.152939
R13388 gnd.n4659 gnd.n4658 0.152939
R13389 gnd.n4660 gnd.n4659 0.152939
R13390 gnd.n4660 gnd.n2107 0.152939
R13391 gnd.n4686 gnd.n2107 0.152939
R13392 gnd.n4687 gnd.n4686 0.152939
R13393 gnd.n4688 gnd.n4687 0.152939
R13394 gnd.n4689 gnd.n4688 0.152939
R13395 gnd.n4689 gnd.n2074 0.152939
R13396 gnd.n4736 gnd.n2074 0.152939
R13397 gnd.n4737 gnd.n4736 0.152939
R13398 gnd.n4738 gnd.n4737 0.152939
R13399 gnd.n4738 gnd.n2051 0.152939
R13400 gnd.n4776 gnd.n2051 0.152939
R13401 gnd.n4777 gnd.n4776 0.152939
R13402 gnd.n4778 gnd.n4777 0.152939
R13403 gnd.n4778 gnd.n2029 0.152939
R13404 gnd.n4833 gnd.n2029 0.152939
R13405 gnd.n4834 gnd.n4833 0.152939
R13406 gnd.n4835 gnd.n4834 0.152939
R13407 gnd.n4835 gnd.n2009 0.152939
R13408 gnd.n4858 gnd.n2009 0.152939
R13409 gnd.n4859 gnd.n4858 0.152939
R13410 gnd.n4860 gnd.n4859 0.152939
R13411 gnd.n4860 gnd.n1989 0.152939
R13412 gnd.n4918 gnd.n1989 0.152939
R13413 gnd.n4919 gnd.n4918 0.152939
R13414 gnd.n4920 gnd.n4919 0.152939
R13415 gnd.n4920 gnd.n1967 0.152939
R13416 gnd.n4947 gnd.n1967 0.152939
R13417 gnd.n4948 gnd.n4947 0.152939
R13418 gnd.n4949 gnd.n4948 0.152939
R13419 gnd.n4950 gnd.n4949 0.152939
R13420 gnd.n4950 gnd.n1939 0.152939
R13421 gnd.n4998 gnd.n1939 0.152939
R13422 gnd.n4999 gnd.n4998 0.152939
R13423 gnd.n5000 gnd.n4999 0.152939
R13424 gnd.n5000 gnd.n1919 0.152939
R13425 gnd.n5024 gnd.n1919 0.152939
R13426 gnd.n5025 gnd.n5024 0.152939
R13427 gnd.n5026 gnd.n5025 0.152939
R13428 gnd.n5027 gnd.n5026 0.152939
R13429 gnd.n5027 gnd.n1889 0.152939
R13430 gnd.n5068 gnd.n1889 0.152939
R13431 gnd.n5069 gnd.n5068 0.152939
R13432 gnd.n5070 gnd.n5069 0.152939
R13433 gnd.n5072 gnd.n5070 0.152939
R13434 gnd.n5072 gnd.n5071 0.152939
R13435 gnd.n5071 gnd.n1840 0.152939
R13436 gnd.n1841 gnd.n1840 0.152939
R13437 gnd.n1842 gnd.n1841 0.152939
R13438 gnd.n1851 gnd.n1842 0.152939
R13439 gnd.n1852 gnd.n1851 0.152939
R13440 gnd.n1853 gnd.n1852 0.152939
R13441 gnd.n1854 gnd.n1853 0.152939
R13442 gnd.n1855 gnd.n1854 0.152939
R13443 gnd.n1857 gnd.n1855 0.152939
R13444 gnd.n1857 gnd.n1856 0.152939
R13445 gnd.n1856 gnd.n1592 0.152939
R13446 gnd.n1593 gnd.n1592 0.152939
R13447 gnd.n1594 gnd.n1593 0.152939
R13448 gnd.n1600 gnd.n1594 0.152939
R13449 gnd.n1601 gnd.n1600 0.152939
R13450 gnd.n1602 gnd.n1601 0.152939
R13451 gnd.n1603 gnd.n1602 0.152939
R13452 gnd.n5705 gnd.n1603 0.152939
R13453 gnd.n5708 gnd.n5705 0.152939
R13454 gnd.n5709 gnd.n5708 0.152939
R13455 gnd.n5710 gnd.n5709 0.152939
R13456 gnd.n5710 gnd.n5701 0.152939
R13457 gnd.n5716 gnd.n5701 0.152939
R13458 gnd.n5717 gnd.n5716 0.152939
R13459 gnd.n5718 gnd.n5717 0.152939
R13460 gnd.n5718 gnd.n1739 0.152939
R13461 gnd.n5724 gnd.n1739 0.152939
R13462 gnd.n5725 gnd.n5724 0.152939
R13463 gnd.n5726 gnd.n5725 0.152939
R13464 gnd.n5727 gnd.n5726 0.152939
R13465 gnd.n5728 gnd.n5727 0.152939
R13466 gnd.n5730 gnd.n5728 0.152939
R13467 gnd.n5731 gnd.n5730 0.152939
R13468 gnd.n4051 gnd.n4034 0.152939
R13469 gnd.n4035 gnd.n4034 0.152939
R13470 gnd.n4036 gnd.n4035 0.152939
R13471 gnd.n4037 gnd.n4036 0.152939
R13472 gnd.n4038 gnd.n4037 0.152939
R13473 gnd.n4039 gnd.n4038 0.152939
R13474 gnd.n4039 gnd.n2417 0.152939
R13475 gnd.n4255 gnd.n2417 0.152939
R13476 gnd.n4256 gnd.n4255 0.152939
R13477 gnd.n4257 gnd.n4256 0.152939
R13478 gnd.n4257 gnd.n2394 0.152939
R13479 gnd.n4270 gnd.n2394 0.152939
R13480 gnd.n4271 gnd.n4270 0.152939
R13481 gnd.n4272 gnd.n4271 0.152939
R13482 gnd.n4274 gnd.n4272 0.152939
R13483 gnd.n4274 gnd.n4273 0.152939
R13484 gnd.n4273 gnd.n2374 0.152939
R13485 gnd.n2375 gnd.n2374 0.152939
R13486 gnd.n2376 gnd.n2375 0.152939
R13487 gnd.n4292 gnd.n2376 0.152939
R13488 gnd.n4015 gnd.n4014 0.152939
R13489 gnd.n4016 gnd.n4015 0.152939
R13490 gnd.n4017 gnd.n4016 0.152939
R13491 gnd.n4018 gnd.n4017 0.152939
R13492 gnd.n4019 gnd.n4018 0.152939
R13493 gnd.n4020 gnd.n4019 0.152939
R13494 gnd.n4021 gnd.n4020 0.152939
R13495 gnd.n4022 gnd.n4021 0.152939
R13496 gnd.n4023 gnd.n4022 0.152939
R13497 gnd.n4024 gnd.n4023 0.152939
R13498 gnd.n4025 gnd.n4024 0.152939
R13499 gnd.n4026 gnd.n4025 0.152939
R13500 gnd.n4027 gnd.n4026 0.152939
R13501 gnd.n4028 gnd.n4027 0.152939
R13502 gnd.n4029 gnd.n4028 0.152939
R13503 gnd.n4055 gnd.n4029 0.152939
R13504 gnd.n4055 gnd.n4054 0.152939
R13505 gnd.n4054 gnd.n4053 0.152939
R13506 gnd.n1072 gnd.n1018 0.152939
R13507 gnd.n1073 gnd.n1072 0.152939
R13508 gnd.n1074 gnd.n1073 0.152939
R13509 gnd.n1075 gnd.n1074 0.152939
R13510 gnd.n1092 gnd.n1075 0.152939
R13511 gnd.n1093 gnd.n1092 0.152939
R13512 gnd.n1094 gnd.n1093 0.152939
R13513 gnd.n1095 gnd.n1094 0.152939
R13514 gnd.n1112 gnd.n1095 0.152939
R13515 gnd.n1113 gnd.n1112 0.152939
R13516 gnd.n1114 gnd.n1113 0.152939
R13517 gnd.n1115 gnd.n1114 0.152939
R13518 gnd.n1133 gnd.n1115 0.152939
R13519 gnd.n1134 gnd.n1133 0.152939
R13520 gnd.n1135 gnd.n1134 0.152939
R13521 gnd.n1136 gnd.n1135 0.152939
R13522 gnd.n1291 gnd.n1290 0.152939
R13523 gnd.n1292 gnd.n1291 0.152939
R13524 gnd.n1293 gnd.n1292 0.152939
R13525 gnd.n1294 gnd.n1293 0.152939
R13526 gnd.n1295 gnd.n1294 0.152939
R13527 gnd.n1296 gnd.n1295 0.152939
R13528 gnd.n1297 gnd.n1296 0.152939
R13529 gnd.n1298 gnd.n1297 0.152939
R13530 gnd.n1299 gnd.n1298 0.152939
R13531 gnd.n1300 gnd.n1299 0.152939
R13532 gnd.n1301 gnd.n1300 0.152939
R13533 gnd.n1302 gnd.n1301 0.152939
R13534 gnd.n1303 gnd.n1302 0.152939
R13535 gnd.n1304 gnd.n1303 0.152939
R13536 gnd.n1305 gnd.n1304 0.152939
R13537 gnd.n1306 gnd.n1305 0.152939
R13538 gnd.n1307 gnd.n1306 0.152939
R13539 gnd.n1310 gnd.n1307 0.152939
R13540 gnd.n1311 gnd.n1310 0.152939
R13541 gnd.n1312 gnd.n1311 0.152939
R13542 gnd.n1313 gnd.n1312 0.152939
R13543 gnd.n1314 gnd.n1313 0.152939
R13544 gnd.n1315 gnd.n1314 0.152939
R13545 gnd.n1316 gnd.n1315 0.152939
R13546 gnd.n1317 gnd.n1316 0.152939
R13547 gnd.n1415 gnd.n1414 0.152939
R13548 gnd.n1414 gnd.n1320 0.152939
R13549 gnd.n1321 gnd.n1320 0.152939
R13550 gnd.n1322 gnd.n1321 0.152939
R13551 gnd.n1323 gnd.n1322 0.152939
R13552 gnd.n1324 gnd.n1323 0.152939
R13553 gnd.n1325 gnd.n1324 0.152939
R13554 gnd.n1326 gnd.n1325 0.152939
R13555 gnd.n1394 gnd.n1326 0.152939
R13556 gnd.n1394 gnd.n1393 0.152939
R13557 gnd.n1393 gnd.n1392 0.152939
R13558 gnd.n1392 gnd.n1330 0.152939
R13559 gnd.n1331 gnd.n1330 0.152939
R13560 gnd.n1332 gnd.n1331 0.152939
R13561 gnd.n1333 gnd.n1332 0.152939
R13562 gnd.n1334 gnd.n1333 0.152939
R13563 gnd.n1335 gnd.n1334 0.152939
R13564 gnd.n1336 gnd.n1335 0.152939
R13565 gnd.n1337 gnd.n1336 0.152939
R13566 gnd.n1338 gnd.n1337 0.152939
R13567 gnd.n1339 gnd.n1338 0.152939
R13568 gnd.n1340 gnd.n1339 0.152939
R13569 gnd.n1341 gnd.n1340 0.152939
R13570 gnd.n1342 gnd.n1341 0.152939
R13571 gnd.n1343 gnd.n1342 0.152939
R13572 gnd.n1344 gnd.n1343 0.152939
R13573 gnd.n1345 gnd.n1344 0.152939
R13574 gnd.n1346 gnd.n1345 0.152939
R13575 gnd.n1352 gnd.n1346 0.152939
R13576 gnd.n1352 gnd.n1351 0.152939
R13577 gnd.n4215 gnd.n2447 0.152939
R13578 gnd.n3951 gnd.n2447 0.152939
R13579 gnd.n3952 gnd.n3951 0.152939
R13580 gnd.n3953 gnd.n3952 0.152939
R13581 gnd.n3954 gnd.n3953 0.152939
R13582 gnd.n3955 gnd.n3954 0.152939
R13583 gnd.n3956 gnd.n3955 0.152939
R13584 gnd.n3957 gnd.n3956 0.152939
R13585 gnd.n3958 gnd.n3957 0.152939
R13586 gnd.n3959 gnd.n3958 0.152939
R13587 gnd.n3960 gnd.n3959 0.152939
R13588 gnd.n3961 gnd.n3960 0.152939
R13589 gnd.n3962 gnd.n3961 0.152939
R13590 gnd.n3963 gnd.n3962 0.152939
R13591 gnd.n3964 gnd.n3963 0.152939
R13592 gnd.n3965 gnd.n3964 0.152939
R13593 gnd.n3966 gnd.n3965 0.152939
R13594 gnd.n3969 gnd.n3966 0.152939
R13595 gnd.n3970 gnd.n3969 0.152939
R13596 gnd.n3971 gnd.n3970 0.152939
R13597 gnd.n3972 gnd.n3971 0.152939
R13598 gnd.n3973 gnd.n3972 0.152939
R13599 gnd.n3974 gnd.n3973 0.152939
R13600 gnd.n3975 gnd.n3974 0.152939
R13601 gnd.n3976 gnd.n3975 0.152939
R13602 gnd.n3977 gnd.n3976 0.152939
R13603 gnd.n3978 gnd.n3977 0.152939
R13604 gnd.n3979 gnd.n3978 0.152939
R13605 gnd.n3980 gnd.n3979 0.152939
R13606 gnd.n3981 gnd.n3980 0.152939
R13607 gnd.n3982 gnd.n3981 0.152939
R13608 gnd.n3983 gnd.n3982 0.152939
R13609 gnd.n3984 gnd.n3983 0.152939
R13610 gnd.n3985 gnd.n3984 0.152939
R13611 gnd.n3986 gnd.n3985 0.152939
R13612 gnd.n3987 gnd.n3986 0.152939
R13613 gnd.n3988 gnd.n3987 0.152939
R13614 gnd.n3991 gnd.n3988 0.152939
R13615 gnd.n3992 gnd.n3991 0.152939
R13616 gnd.n3993 gnd.n3992 0.152939
R13617 gnd.n3994 gnd.n3993 0.152939
R13618 gnd.n3995 gnd.n3994 0.152939
R13619 gnd.n3996 gnd.n3995 0.152939
R13620 gnd.n3997 gnd.n3996 0.152939
R13621 gnd.n3998 gnd.n3997 0.152939
R13622 gnd.n3999 gnd.n3998 0.152939
R13623 gnd.n4000 gnd.n3999 0.152939
R13624 gnd.n4001 gnd.n4000 0.152939
R13625 gnd.n4002 gnd.n4001 0.152939
R13626 gnd.n4003 gnd.n4002 0.152939
R13627 gnd.n4004 gnd.n4003 0.152939
R13628 gnd.n4005 gnd.n4004 0.152939
R13629 gnd.n4006 gnd.n4005 0.152939
R13630 gnd.n4007 gnd.n4006 0.152939
R13631 gnd.n4008 gnd.n4007 0.152939
R13632 gnd.n4009 gnd.n4008 0.152939
R13633 gnd.n4098 gnd.n4009 0.152939
R13634 gnd.n4098 gnd.n4097 0.152939
R13635 gnd.n4217 gnd.n4216 0.152939
R13636 gnd.n4217 gnd.n2428 0.152939
R13637 gnd.n4237 gnd.n2428 0.152939
R13638 gnd.n4238 gnd.n4237 0.152939
R13639 gnd.n4240 gnd.n4238 0.152939
R13640 gnd.n4240 gnd.n4239 0.152939
R13641 gnd.n4239 gnd.n975 0.152939
R13642 gnd.n976 gnd.n975 0.152939
R13643 gnd.n977 gnd.n976 0.152939
R13644 gnd.n996 gnd.n977 0.152939
R13645 gnd.n997 gnd.n996 0.152939
R13646 gnd.n998 gnd.n997 0.152939
R13647 gnd.n999 gnd.n998 0.152939
R13648 gnd.n1016 gnd.n999 0.152939
R13649 gnd.n1017 gnd.n1016 0.152939
R13650 gnd.n1018 gnd.n1017 0.152939
R13651 gnd.n6309 gnd.n964 0.152939
R13652 gnd.n2400 gnd.n964 0.152939
R13653 gnd.n2401 gnd.n2400 0.152939
R13654 gnd.n2402 gnd.n2401 0.152939
R13655 gnd.n2403 gnd.n2402 0.152939
R13656 gnd.n2405 gnd.n2403 0.152939
R13657 gnd.n2406 gnd.n2405 0.152939
R13658 gnd.n2406 gnd.n2365 0.152939
R13659 gnd.n4337 gnd.n2365 0.152939
R13660 gnd.n6480 gnd.n797 0.152939
R13661 gnd.n802 gnd.n797 0.152939
R13662 gnd.n803 gnd.n802 0.152939
R13663 gnd.n804 gnd.n803 0.152939
R13664 gnd.n805 gnd.n804 0.152939
R13665 gnd.n810 gnd.n805 0.152939
R13666 gnd.n811 gnd.n810 0.152939
R13667 gnd.n812 gnd.n811 0.152939
R13668 gnd.n813 gnd.n812 0.152939
R13669 gnd.n818 gnd.n813 0.152939
R13670 gnd.n819 gnd.n818 0.152939
R13671 gnd.n820 gnd.n819 0.152939
R13672 gnd.n821 gnd.n820 0.152939
R13673 gnd.n826 gnd.n821 0.152939
R13674 gnd.n827 gnd.n826 0.152939
R13675 gnd.n828 gnd.n827 0.152939
R13676 gnd.n829 gnd.n828 0.152939
R13677 gnd.n834 gnd.n829 0.152939
R13678 gnd.n835 gnd.n834 0.152939
R13679 gnd.n836 gnd.n835 0.152939
R13680 gnd.n837 gnd.n836 0.152939
R13681 gnd.n842 gnd.n837 0.152939
R13682 gnd.n843 gnd.n842 0.152939
R13683 gnd.n844 gnd.n843 0.152939
R13684 gnd.n845 gnd.n844 0.152939
R13685 gnd.n850 gnd.n845 0.152939
R13686 gnd.n851 gnd.n850 0.152939
R13687 gnd.n852 gnd.n851 0.152939
R13688 gnd.n853 gnd.n852 0.152939
R13689 gnd.n858 gnd.n853 0.152939
R13690 gnd.n859 gnd.n858 0.152939
R13691 gnd.n860 gnd.n859 0.152939
R13692 gnd.n861 gnd.n860 0.152939
R13693 gnd.n866 gnd.n861 0.152939
R13694 gnd.n867 gnd.n866 0.152939
R13695 gnd.n868 gnd.n867 0.152939
R13696 gnd.n869 gnd.n868 0.152939
R13697 gnd.n874 gnd.n869 0.152939
R13698 gnd.n875 gnd.n874 0.152939
R13699 gnd.n876 gnd.n875 0.152939
R13700 gnd.n877 gnd.n876 0.152939
R13701 gnd.n882 gnd.n877 0.152939
R13702 gnd.n883 gnd.n882 0.152939
R13703 gnd.n884 gnd.n883 0.152939
R13704 gnd.n885 gnd.n884 0.152939
R13705 gnd.n890 gnd.n885 0.152939
R13706 gnd.n891 gnd.n890 0.152939
R13707 gnd.n892 gnd.n891 0.152939
R13708 gnd.n893 gnd.n892 0.152939
R13709 gnd.n898 gnd.n893 0.152939
R13710 gnd.n899 gnd.n898 0.152939
R13711 gnd.n900 gnd.n899 0.152939
R13712 gnd.n901 gnd.n900 0.152939
R13713 gnd.n906 gnd.n901 0.152939
R13714 gnd.n907 gnd.n906 0.152939
R13715 gnd.n908 gnd.n907 0.152939
R13716 gnd.n909 gnd.n908 0.152939
R13717 gnd.n914 gnd.n909 0.152939
R13718 gnd.n915 gnd.n914 0.152939
R13719 gnd.n916 gnd.n915 0.152939
R13720 gnd.n917 gnd.n916 0.152939
R13721 gnd.n922 gnd.n917 0.152939
R13722 gnd.n923 gnd.n922 0.152939
R13723 gnd.n924 gnd.n923 0.152939
R13724 gnd.n925 gnd.n924 0.152939
R13725 gnd.n930 gnd.n925 0.152939
R13726 gnd.n931 gnd.n930 0.152939
R13727 gnd.n932 gnd.n931 0.152939
R13728 gnd.n933 gnd.n932 0.152939
R13729 gnd.n938 gnd.n933 0.152939
R13730 gnd.n939 gnd.n938 0.152939
R13731 gnd.n940 gnd.n939 0.152939
R13732 gnd.n941 gnd.n940 0.152939
R13733 gnd.n946 gnd.n941 0.152939
R13734 gnd.n947 gnd.n946 0.152939
R13735 gnd.n948 gnd.n947 0.152939
R13736 gnd.n949 gnd.n948 0.152939
R13737 gnd.n954 gnd.n949 0.152939
R13738 gnd.n955 gnd.n954 0.152939
R13739 gnd.n956 gnd.n955 0.152939
R13740 gnd.n957 gnd.n956 0.152939
R13741 gnd.n962 gnd.n957 0.152939
R13742 gnd.n963 gnd.n962 0.152939
R13743 gnd.n6310 gnd.n963 0.152939
R13744 gnd.n2316 gnd.n2315 0.152939
R13745 gnd.n2316 gnd.n2302 0.152939
R13746 gnd.n4460 gnd.n2302 0.152939
R13747 gnd.n4461 gnd.n4460 0.152939
R13748 gnd.n4465 gnd.n4461 0.152939
R13749 gnd.n4465 gnd.n4464 0.152939
R13750 gnd.n4464 gnd.n4463 0.152939
R13751 gnd.n4463 gnd.n2201 0.152939
R13752 gnd.n4497 gnd.n2201 0.152939
R13753 gnd.n4498 gnd.n4497 0.152939
R13754 gnd.n4500 gnd.n4498 0.152939
R13755 gnd.n4500 gnd.n4499 0.152939
R13756 gnd.n4499 gnd.n2190 0.152939
R13757 gnd.n4522 gnd.n2190 0.152939
R13758 gnd.n4523 gnd.n4522 0.152939
R13759 gnd.n4531 gnd.n4523 0.152939
R13760 gnd.n4531 gnd.n4530 0.152939
R13761 gnd.n4530 gnd.n4529 0.152939
R13762 gnd.n4529 gnd.n4524 0.152939
R13763 gnd.n4524 gnd.n2143 0.152939
R13764 gnd.n4608 gnd.n2143 0.152939
R13765 gnd.n4609 gnd.n4608 0.152939
R13766 gnd.n4629 gnd.n4609 0.152939
R13767 gnd.n4629 gnd.n4628 0.152939
R13768 gnd.n4628 gnd.n4627 0.152939
R13769 gnd.n4627 gnd.n4610 0.152939
R13770 gnd.n4623 gnd.n4610 0.152939
R13771 gnd.n4623 gnd.n4622 0.152939
R13772 gnd.n4622 gnd.n4621 0.152939
R13773 gnd.n4621 gnd.n4618 0.152939
R13774 gnd.n4618 gnd.n4617 0.152939
R13775 gnd.n4617 gnd.n2091 0.152939
R13776 gnd.n4710 gnd.n2091 0.152939
R13777 gnd.n4711 gnd.n4710 0.152939
R13778 gnd.n4712 gnd.n4711 0.152939
R13779 gnd.n4712 gnd.n2067 0.152939
R13780 gnd.n4758 gnd.n2067 0.152939
R13781 gnd.n4758 gnd.n4757 0.152939
R13782 gnd.n4757 gnd.n4756 0.152939
R13783 gnd.n4756 gnd.n2044 0.152939
R13784 gnd.n4817 gnd.n2044 0.152939
R13785 gnd.n4817 gnd.n4816 0.152939
R13786 gnd.n4816 gnd.n4815 0.152939
R13787 gnd.n4815 gnd.n2045 0.152939
R13788 gnd.n4811 gnd.n2045 0.152939
R13789 gnd.n4811 gnd.n4810 0.152939
R13790 gnd.n4810 gnd.n4809 0.152939
R13791 gnd.n4809 gnd.n4799 0.152939
R13792 gnd.n4805 gnd.n4799 0.152939
R13793 gnd.n4805 gnd.n1982 0.152939
R13794 gnd.n4927 gnd.n1982 0.152939
R13795 gnd.n4928 gnd.n4927 0.152939
R13796 gnd.n4930 gnd.n4928 0.152939
R13797 gnd.n4930 gnd.n4929 0.152939
R13798 gnd.n4929 gnd.n1953 0.152939
R13799 gnd.n4966 gnd.n1953 0.152939
R13800 gnd.n4967 gnd.n4966 0.152939
R13801 gnd.n4983 gnd.n4967 0.152939
R13802 gnd.n4983 gnd.n4982 0.152939
R13803 gnd.n4982 gnd.n4981 0.152939
R13804 gnd.n4981 gnd.n4968 0.152939
R13805 gnd.n4977 gnd.n4968 0.152939
R13806 gnd.n4977 gnd.n4976 0.152939
R13807 gnd.n4976 gnd.n4975 0.152939
R13808 gnd.n4975 gnd.n1897 0.152939
R13809 gnd.n5057 gnd.n1897 0.152939
R13810 gnd.n5058 gnd.n5057 0.152939
R13811 gnd.n5060 gnd.n5058 0.152939
R13812 gnd.n5060 gnd.n5059 0.152939
R13813 gnd.n5059 gnd.n1870 0.152939
R13814 gnd.n5099 gnd.n1870 0.152939
R13815 gnd.n5100 gnd.n5099 0.152939
R13816 gnd.n5101 gnd.n5100 0.152939
R13817 gnd.n5101 gnd.n1867 0.152939
R13818 gnd.n5110 gnd.n1867 0.152939
R13819 gnd.n5111 gnd.n5110 0.152939
R13820 gnd.n5112 gnd.n5111 0.152939
R13821 gnd.n5112 gnd.n1865 0.152939
R13822 gnd.n5118 gnd.n1865 0.152939
R13823 gnd.n5119 gnd.n5118 0.152939
R13824 gnd.n5298 gnd.n5119 0.152939
R13825 gnd.n5298 gnd.n5297 0.152939
R13826 gnd.n4312 gnd.n2391 0.152939
R13827 gnd.n4312 gnd.n4311 0.152939
R13828 gnd.n4311 gnd.n4310 0.152939
R13829 gnd.n4310 gnd.n2354 0.152939
R13830 gnd.n4366 gnd.n2354 0.152939
R13831 gnd.n4367 gnd.n4366 0.152939
R13832 gnd.n4368 gnd.n4367 0.152939
R13833 gnd.n4368 gnd.n2348 0.152939
R13834 gnd.n4380 gnd.n2348 0.152939
R13835 gnd.n4381 gnd.n4380 0.152939
R13836 gnd.n4382 gnd.n4381 0.152939
R13837 gnd.n4382 gnd.n2342 0.152939
R13838 gnd.n4406 gnd.n2342 0.152939
R13839 gnd.n4406 gnd.n4405 0.152939
R13840 gnd.n4405 gnd.n4404 0.152939
R13841 gnd.n4404 gnd.n2343 0.152939
R13842 gnd.n4400 gnd.n2343 0.152939
R13843 gnd.n4400 gnd.n1148 0.152939
R13844 gnd.n6189 gnd.n1148 0.152939
R13845 gnd.n6189 gnd.n6188 0.152939
R13846 gnd.n6176 gnd.n1172 0.152939
R13847 gnd.n6176 gnd.n6175 0.152939
R13848 gnd.n6175 gnd.n6174 0.152939
R13849 gnd.n6174 gnd.n1174 0.152939
R13850 gnd.n6170 gnd.n1174 0.152939
R13851 gnd.n6170 gnd.n6169 0.152939
R13852 gnd.n4451 gnd.n2311 0.152939
R13853 gnd.n4452 gnd.n4451 0.152939
R13854 gnd.n4454 gnd.n4452 0.152939
R13855 gnd.n4454 gnd.n4453 0.152939
R13856 gnd.n4453 gnd.n2287 0.152939
R13857 gnd.n4484 gnd.n2287 0.152939
R13858 gnd.n4485 gnd.n4484 0.152939
R13859 gnd.n4490 gnd.n4485 0.152939
R13860 gnd.n4490 gnd.n4489 0.152939
R13861 gnd.n4489 gnd.n4488 0.152939
R13862 gnd.n4488 gnd.n1497 0.152939
R13863 gnd.n5981 gnd.n1497 0.152939
R13864 gnd.n5981 gnd.n5980 0.152939
R13865 gnd.n5980 gnd.n5979 0.152939
R13866 gnd.n5979 gnd.n1498 0.152939
R13867 gnd.n5975 gnd.n1498 0.152939
R13868 gnd.n5975 gnd.n5974 0.152939
R13869 gnd.n5974 gnd.n5973 0.152939
R13870 gnd.n5973 gnd.n1503 0.152939
R13871 gnd.n5969 gnd.n1503 0.152939
R13872 gnd.n5969 gnd.n5968 0.152939
R13873 gnd.n5968 gnd.n5967 0.152939
R13874 gnd.n5967 gnd.n1508 0.152939
R13875 gnd.n5963 gnd.n1508 0.152939
R13876 gnd.n5963 gnd.n5962 0.152939
R13877 gnd.n5962 gnd.n5961 0.152939
R13878 gnd.n5961 gnd.n1513 0.152939
R13879 gnd.n5957 gnd.n1513 0.152939
R13880 gnd.n5957 gnd.n5956 0.152939
R13881 gnd.n5956 gnd.n5955 0.152939
R13882 gnd.n5955 gnd.n1518 0.152939
R13883 gnd.n5951 gnd.n1518 0.152939
R13884 gnd.n5951 gnd.n5950 0.152939
R13885 gnd.n5950 gnd.n5949 0.152939
R13886 gnd.n5949 gnd.n1523 0.152939
R13887 gnd.n5945 gnd.n1523 0.152939
R13888 gnd.n5945 gnd.n5944 0.152939
R13889 gnd.n5944 gnd.n5943 0.152939
R13890 gnd.n5943 gnd.n1528 0.152939
R13891 gnd.n5939 gnd.n1528 0.152939
R13892 gnd.n5939 gnd.n5938 0.152939
R13893 gnd.n5938 gnd.n5937 0.152939
R13894 gnd.n5937 gnd.n1533 0.152939
R13895 gnd.n5933 gnd.n1533 0.152939
R13896 gnd.n5933 gnd.n5932 0.152939
R13897 gnd.n5932 gnd.n5931 0.152939
R13898 gnd.n5931 gnd.n1538 0.152939
R13899 gnd.n5927 gnd.n1538 0.152939
R13900 gnd.n5927 gnd.n5926 0.152939
R13901 gnd.n5926 gnd.n5925 0.152939
R13902 gnd.n5925 gnd.n1543 0.152939
R13903 gnd.n5921 gnd.n1543 0.152939
R13904 gnd.n5921 gnd.n5920 0.152939
R13905 gnd.n5920 gnd.n5919 0.152939
R13906 gnd.n5919 gnd.n1548 0.152939
R13907 gnd.n5915 gnd.n1548 0.152939
R13908 gnd.n5915 gnd.n5914 0.152939
R13909 gnd.n5914 gnd.n5913 0.152939
R13910 gnd.n5913 gnd.n1553 0.152939
R13911 gnd.n5909 gnd.n1553 0.152939
R13912 gnd.n5909 gnd.n5908 0.152939
R13913 gnd.n5908 gnd.n5907 0.152939
R13914 gnd.n5907 gnd.n1558 0.152939
R13915 gnd.n5903 gnd.n1558 0.152939
R13916 gnd.n5903 gnd.n5902 0.152939
R13917 gnd.n5902 gnd.n5901 0.152939
R13918 gnd.n5901 gnd.n1563 0.152939
R13919 gnd.n5897 gnd.n1563 0.152939
R13920 gnd.n5897 gnd.n5896 0.152939
R13921 gnd.n5896 gnd.n5895 0.152939
R13922 gnd.n5895 gnd.n1568 0.152939
R13923 gnd.n5891 gnd.n1568 0.152939
R13924 gnd.n5891 gnd.n5890 0.152939
R13925 gnd.n5890 gnd.n5889 0.152939
R13926 gnd.n5889 gnd.n1573 0.152939
R13927 gnd.n5885 gnd.n1573 0.152939
R13928 gnd.n5885 gnd.n5884 0.152939
R13929 gnd.n5884 gnd.n5883 0.152939
R13930 gnd.n5883 gnd.n1578 0.152939
R13931 gnd.n5879 gnd.n1578 0.152939
R13932 gnd.n5879 gnd.n5878 0.152939
R13933 gnd.n5878 gnd.n5877 0.152939
R13934 gnd.n5184 gnd.n1583 0.152939
R13935 gnd.n5184 gnd.n5180 0.152939
R13936 gnd.n5192 gnd.n5180 0.152939
R13937 gnd.n5193 gnd.n5192 0.152939
R13938 gnd.n5195 gnd.n5193 0.152939
R13939 gnd.n5195 gnd.n5194 0.152939
R13940 gnd.n5125 gnd.n5120 0.152939
R13941 gnd.n5120 gnd.n1749 0.152939
R13942 gnd.n5672 gnd.n1749 0.152939
R13943 gnd.n5673 gnd.n5672 0.152939
R13944 gnd.n5674 gnd.n5673 0.152939
R13945 gnd.n5674 gnd.n1744 0.152939
R13946 gnd.n5694 gnd.n1744 0.152939
R13947 gnd.n5694 gnd.n5693 0.152939
R13948 gnd.n5693 gnd.n5692 0.152939
R13949 gnd.n5692 gnd.n1745 0.152939
R13950 gnd.n5688 gnd.n1745 0.152939
R13951 gnd.n5688 gnd.n1732 0.152939
R13952 gnd.n5752 gnd.n1732 0.152939
R13953 gnd.n5753 gnd.n5752 0.152939
R13954 gnd.n5764 gnd.n5753 0.152939
R13955 gnd.n5764 gnd.n5763 0.152939
R13956 gnd.n5763 gnd.n5762 0.152939
R13957 gnd.n5762 gnd.n5754 0.152939
R13958 gnd.n5758 gnd.n5754 0.152939
R13959 gnd.n5758 gnd.n63 0.152939
R13960 gnd.n7344 gnd.n7343 0.145814
R13961 gnd.n4293 gnd.n4292 0.145814
R13962 gnd.n4293 gnd.n2391 0.145814
R13963 gnd.n7344 gnd.n63 0.145814
R13964 gnd.n6169 gnd.n6168 0.128549
R13965 gnd.n5194 gnd.n1753 0.128549
R13966 gnd.n2729 gnd.n0 0.127478
R13967 gnd.n405 gnd.n79 0.10111
R13968 gnd.n4338 gnd.n4337 0.10111
R13969 gnd.n3309 gnd.n3308 0.0767195
R13970 gnd.n3308 gnd.n3307 0.0767195
R13971 gnd.n6168 gnd.n1144 0.063
R13972 gnd.n5661 gnd.n1753 0.063
R13973 gnd.n5663 gnd.n5661 0.0538288
R13974 gnd.n7280 gnd.n385 0.0538288
R13975 gnd.n4096 gnd.n4095 0.0538288
R13976 gnd.n6196 gnd.n1144 0.0538288
R13977 gnd.n4339 gnd.n4338 0.0523293
R13978 gnd.n5731 gnd.n79 0.0523293
R13979 gnd.n3875 gnd.n2491 0.0477147
R13980 gnd.n3072 gnd.n2960 0.0442063
R13981 gnd.n3073 gnd.n3072 0.0442063
R13982 gnd.n3074 gnd.n3073 0.0442063
R13983 gnd.n3074 gnd.n2949 0.0442063
R13984 gnd.n3088 gnd.n2949 0.0442063
R13985 gnd.n3089 gnd.n3088 0.0442063
R13986 gnd.n3090 gnd.n3089 0.0442063
R13987 gnd.n3090 gnd.n2936 0.0442063
R13988 gnd.n3134 gnd.n2936 0.0442063
R13989 gnd.n3135 gnd.n3134 0.0442063
R13990 gnd.n3137 gnd.n2870 0.0344674
R13991 gnd.n5664 gnd.n5663 0.0344674
R13992 gnd.n5664 gnd.n1625 0.0344674
R13993 gnd.n1626 gnd.n1625 0.0344674
R13994 gnd.n1627 gnd.n1626 0.0344674
R13995 gnd.n1747 gnd.n1627 0.0344674
R13996 gnd.n1747 gnd.n1645 0.0344674
R13997 gnd.n1646 gnd.n1645 0.0344674
R13998 gnd.n1647 gnd.n1646 0.0344674
R13999 gnd.n5683 gnd.n1647 0.0344674
R14000 gnd.n5683 gnd.n1666 0.0344674
R14001 gnd.n1667 gnd.n1666 0.0344674
R14002 gnd.n1668 gnd.n1667 0.0344674
R14003 gnd.n5746 gnd.n1668 0.0344674
R14004 gnd.n5746 gnd.n1685 0.0344674
R14005 gnd.n1686 gnd.n1685 0.0344674
R14006 gnd.n1687 gnd.n1686 0.0344674
R14007 gnd.n1727 gnd.n1687 0.0344674
R14008 gnd.n5775 gnd.n1727 0.0344674
R14009 gnd.n5780 gnd.n5775 0.0344674
R14010 gnd.n5781 gnd.n5780 0.0344674
R14011 gnd.n5781 gnd.n1725 0.0344674
R14012 gnd.n5788 gnd.n1725 0.0344674
R14013 gnd.n5788 gnd.n400 0.0344674
R14014 gnd.n7140 gnd.n400 0.0344674
R14015 gnd.n7141 gnd.n7140 0.0344674
R14016 gnd.n7141 gnd.n93 0.0344674
R14017 gnd.n94 gnd.n93 0.0344674
R14018 gnd.n95 gnd.n94 0.0344674
R14019 gnd.n7156 gnd.n95 0.0344674
R14020 gnd.n7156 gnd.n112 0.0344674
R14021 gnd.n113 gnd.n112 0.0344674
R14022 gnd.n114 gnd.n113 0.0344674
R14023 gnd.n7171 gnd.n114 0.0344674
R14024 gnd.n7171 gnd.n133 0.0344674
R14025 gnd.n134 gnd.n133 0.0344674
R14026 gnd.n135 gnd.n134 0.0344674
R14027 gnd.n7270 gnd.n135 0.0344674
R14028 gnd.n7270 gnd.n154 0.0344674
R14029 gnd.n155 gnd.n154 0.0344674
R14030 gnd.n156 gnd.n155 0.0344674
R14031 gnd.n172 gnd.n156 0.0344674
R14032 gnd.n7280 gnd.n172 0.0344674
R14033 gnd.n4095 gnd.n4093 0.0344674
R14034 gnd.n4093 gnd.n2440 0.0344674
R14035 gnd.n2440 gnd.n2437 0.0344674
R14036 gnd.n4230 gnd.n2437 0.0344674
R14037 gnd.n4230 gnd.n2438 0.0344674
R14038 gnd.n2438 gnd.n2420 0.0344674
R14039 gnd.n4248 gnd.n2420 0.0344674
R14040 gnd.n4249 gnd.n4248 0.0344674
R14041 gnd.n4249 gnd.n986 0.0344674
R14042 gnd.n987 gnd.n986 0.0344674
R14043 gnd.n988 gnd.n987 0.0344674
R14044 gnd.n4264 gnd.n988 0.0344674
R14045 gnd.n4264 gnd.n1007 0.0344674
R14046 gnd.n1008 gnd.n1007 0.0344674
R14047 gnd.n1009 gnd.n1008 0.0344674
R14048 gnd.n4285 gnd.n1009 0.0344674
R14049 gnd.n4286 gnd.n4285 0.0344674
R14050 gnd.n4286 gnd.n1029 0.0344674
R14051 gnd.n1030 gnd.n1029 0.0344674
R14052 gnd.n1031 gnd.n1030 0.0344674
R14053 gnd.n4291 gnd.n1031 0.0344674
R14054 gnd.n4291 gnd.n1045 0.0344674
R14055 gnd.n1046 gnd.n1045 0.0344674
R14056 gnd.n1047 gnd.n1046 0.0344674
R14057 gnd.n4302 gnd.n1047 0.0344674
R14058 gnd.n4302 gnd.n1063 0.0344674
R14059 gnd.n1064 gnd.n1063 0.0344674
R14060 gnd.n1065 gnd.n1064 0.0344674
R14061 gnd.n2352 gnd.n1065 0.0344674
R14062 gnd.n2352 gnd.n1082 0.0344674
R14063 gnd.n1083 gnd.n1082 0.0344674
R14064 gnd.n1084 gnd.n1083 0.0344674
R14065 gnd.n2346 gnd.n1084 0.0344674
R14066 gnd.n2346 gnd.n1103 0.0344674
R14067 gnd.n1104 gnd.n1103 0.0344674
R14068 gnd.n1105 gnd.n1104 0.0344674
R14069 gnd.n4391 gnd.n1105 0.0344674
R14070 gnd.n4391 gnd.n1123 0.0344674
R14071 gnd.n1124 gnd.n1123 0.0344674
R14072 gnd.n1125 gnd.n1124 0.0344674
R14073 gnd.n1143 gnd.n1125 0.0344674
R14074 gnd.n6196 gnd.n1143 0.0344674
R14075 gnd.n6167 gnd.n1179 0.0344674
R14076 gnd.n5204 gnd.n5203 0.0344674
R14077 gnd.n6187 gnd.n6186 0.029712
R14078 gnd.n5135 gnd.n5126 0.029712
R14079 gnd.n3157 gnd.n3156 0.0269946
R14080 gnd.n3159 gnd.n3158 0.0269946
R14081 gnd.n2865 gnd.n2863 0.0269946
R14082 gnd.n3169 gnd.n3167 0.0269946
R14083 gnd.n3168 gnd.n2844 0.0269946
R14084 gnd.n3188 gnd.n3187 0.0269946
R14085 gnd.n3190 gnd.n3189 0.0269946
R14086 gnd.n2839 gnd.n2838 0.0269946
R14087 gnd.n3200 gnd.n2834 0.0269946
R14088 gnd.n3199 gnd.n2836 0.0269946
R14089 gnd.n2835 gnd.n2817 0.0269946
R14090 gnd.n3220 gnd.n2818 0.0269946
R14091 gnd.n3219 gnd.n2819 0.0269946
R14092 gnd.n3253 gnd.n2794 0.0269946
R14093 gnd.n3255 gnd.n3254 0.0269946
R14094 gnd.n3256 gnd.n2741 0.0269946
R14095 gnd.n2789 gnd.n2742 0.0269946
R14096 gnd.n2791 gnd.n2743 0.0269946
R14097 gnd.n3266 gnd.n3265 0.0269946
R14098 gnd.n3268 gnd.n3267 0.0269946
R14099 gnd.n3269 gnd.n2763 0.0269946
R14100 gnd.n3271 gnd.n2764 0.0269946
R14101 gnd.n3274 gnd.n2765 0.0269946
R14102 gnd.n3277 gnd.n3276 0.0269946
R14103 gnd.n3279 gnd.n3278 0.0269946
R14104 gnd.n3344 gnd.n2664 0.0269946
R14105 gnd.n3346 gnd.n3345 0.0269946
R14106 gnd.n3355 gnd.n2657 0.0269946
R14107 gnd.n3357 gnd.n3356 0.0269946
R14108 gnd.n3358 gnd.n2655 0.0269946
R14109 gnd.n3365 gnd.n3361 0.0269946
R14110 gnd.n3364 gnd.n3363 0.0269946
R14111 gnd.n3362 gnd.n2634 0.0269946
R14112 gnd.n3387 gnd.n2635 0.0269946
R14113 gnd.n3386 gnd.n2636 0.0269946
R14114 gnd.n3429 gnd.n2609 0.0269946
R14115 gnd.n3431 gnd.n3430 0.0269946
R14116 gnd.n3440 gnd.n2602 0.0269946
R14117 gnd.n3442 gnd.n3441 0.0269946
R14118 gnd.n3443 gnd.n2600 0.0269946
R14119 gnd.n3450 gnd.n3446 0.0269946
R14120 gnd.n3449 gnd.n3448 0.0269946
R14121 gnd.n3447 gnd.n2579 0.0269946
R14122 gnd.n3472 gnd.n2580 0.0269946
R14123 gnd.n3471 gnd.n2581 0.0269946
R14124 gnd.n3518 gnd.n2555 0.0269946
R14125 gnd.n3520 gnd.n3519 0.0269946
R14126 gnd.n3529 gnd.n2548 0.0269946
R14127 gnd.n3788 gnd.n2546 0.0269946
R14128 gnd.n3793 gnd.n3791 0.0269946
R14129 gnd.n3792 gnd.n2527 0.0269946
R14130 gnd.n3817 gnd.n3816 0.0269946
R14131 gnd.n6163 gnd.n1185 0.0225788
R14132 gnd.n6162 gnd.n1186 0.0225788
R14133 gnd.n6159 gnd.n6158 0.0225788
R14134 gnd.n6155 gnd.n1191 0.0225788
R14135 gnd.n6154 gnd.n1197 0.0225788
R14136 gnd.n6151 gnd.n6150 0.0225788
R14137 gnd.n6147 gnd.n1201 0.0225788
R14138 gnd.n6146 gnd.n1205 0.0225788
R14139 gnd.n6143 gnd.n6142 0.0225788
R14140 gnd.n6139 gnd.n1209 0.0225788
R14141 gnd.n6138 gnd.n1215 0.0225788
R14142 gnd.n6135 gnd.n6134 0.0225788
R14143 gnd.n6131 gnd.n1219 0.0225788
R14144 gnd.n6130 gnd.n1223 0.0225788
R14145 gnd.n6127 gnd.n6126 0.0225788
R14146 gnd.n6123 gnd.n1227 0.0225788
R14147 gnd.n6122 gnd.n1236 0.0225788
R14148 gnd.n1241 gnd.n1240 0.0225788
R14149 gnd.n6186 gnd.n1150 0.0225788
R14150 gnd.n5210 gnd.n5208 0.0225788
R14151 gnd.n5209 gnd.n5172 0.0225788
R14152 gnd.n5219 gnd.n5218 0.0225788
R14153 gnd.n5173 gnd.n5168 0.0225788
R14154 gnd.n5229 gnd.n5227 0.0225788
R14155 gnd.n5228 gnd.n5163 0.0225788
R14156 gnd.n5238 gnd.n5237 0.0225788
R14157 gnd.n5164 gnd.n5159 0.0225788
R14158 gnd.n5248 gnd.n5246 0.0225788
R14159 gnd.n5247 gnd.n5154 0.0225788
R14160 gnd.n5257 gnd.n5256 0.0225788
R14161 gnd.n5155 gnd.n5150 0.0225788
R14162 gnd.n5267 gnd.n5265 0.0225788
R14163 gnd.n5266 gnd.n5145 0.0225788
R14164 gnd.n5277 gnd.n5276 0.0225788
R14165 gnd.n5273 gnd.n5146 0.0225788
R14166 gnd.n5287 gnd.n5133 0.0225788
R14167 gnd.n5286 gnd.n5134 0.0225788
R14168 gnd.n5136 gnd.n5135 0.0225788
R14169 gnd.n5296 gnd.n5126 0.0218415
R14170 gnd.n6187 gnd.n1149 0.0218415
R14171 gnd.n3137 gnd.n3136 0.0202011
R14172 gnd.n3136 gnd.n3135 0.0148637
R14173 gnd.n3786 gnd.n3530 0.0144266
R14174 gnd.n3787 gnd.n3786 0.0130679
R14175 gnd.n1185 gnd.n1179 0.0123886
R14176 gnd.n6163 gnd.n6162 0.0123886
R14177 gnd.n6159 gnd.n1186 0.0123886
R14178 gnd.n6158 gnd.n1191 0.0123886
R14179 gnd.n6155 gnd.n6154 0.0123886
R14180 gnd.n6151 gnd.n1197 0.0123886
R14181 gnd.n6150 gnd.n1201 0.0123886
R14182 gnd.n6147 gnd.n6146 0.0123886
R14183 gnd.n6143 gnd.n1205 0.0123886
R14184 gnd.n6142 gnd.n1209 0.0123886
R14185 gnd.n6139 gnd.n6138 0.0123886
R14186 gnd.n6135 gnd.n1215 0.0123886
R14187 gnd.n6134 gnd.n1219 0.0123886
R14188 gnd.n6131 gnd.n6130 0.0123886
R14189 gnd.n6127 gnd.n1223 0.0123886
R14190 gnd.n6126 gnd.n1227 0.0123886
R14191 gnd.n6123 gnd.n6122 0.0123886
R14192 gnd.n1241 gnd.n1236 0.0123886
R14193 gnd.n1240 gnd.n1150 0.0123886
R14194 gnd.n5208 gnd.n5204 0.0123886
R14195 gnd.n5210 gnd.n5209 0.0123886
R14196 gnd.n5219 gnd.n5172 0.0123886
R14197 gnd.n5218 gnd.n5173 0.0123886
R14198 gnd.n5227 gnd.n5168 0.0123886
R14199 gnd.n5229 gnd.n5228 0.0123886
R14200 gnd.n5238 gnd.n5163 0.0123886
R14201 gnd.n5237 gnd.n5164 0.0123886
R14202 gnd.n5246 gnd.n5159 0.0123886
R14203 gnd.n5248 gnd.n5247 0.0123886
R14204 gnd.n5257 gnd.n5154 0.0123886
R14205 gnd.n5256 gnd.n5155 0.0123886
R14206 gnd.n5265 gnd.n5150 0.0123886
R14207 gnd.n5267 gnd.n5266 0.0123886
R14208 gnd.n5277 gnd.n5145 0.0123886
R14209 gnd.n5276 gnd.n5146 0.0123886
R14210 gnd.n5273 gnd.n5133 0.0123886
R14211 gnd.n5287 gnd.n5286 0.0123886
R14212 gnd.n5136 gnd.n5134 0.0123886
R14213 gnd.n3156 gnd.n2870 0.00797283
R14214 gnd.n3158 gnd.n3157 0.00797283
R14215 gnd.n3159 gnd.n2865 0.00797283
R14216 gnd.n3167 gnd.n2863 0.00797283
R14217 gnd.n3169 gnd.n3168 0.00797283
R14218 gnd.n3187 gnd.n2844 0.00797283
R14219 gnd.n3189 gnd.n3188 0.00797283
R14220 gnd.n3190 gnd.n2839 0.00797283
R14221 gnd.n2838 gnd.n2834 0.00797283
R14222 gnd.n3200 gnd.n3199 0.00797283
R14223 gnd.n2836 gnd.n2835 0.00797283
R14224 gnd.n2818 gnd.n2817 0.00797283
R14225 gnd.n3220 gnd.n3219 0.00797283
R14226 gnd.n2819 gnd.n2794 0.00797283
R14227 gnd.n3254 gnd.n3253 0.00797283
R14228 gnd.n3256 gnd.n3255 0.00797283
R14229 gnd.n2789 gnd.n2741 0.00797283
R14230 gnd.n2791 gnd.n2742 0.00797283
R14231 gnd.n3265 gnd.n2743 0.00797283
R14232 gnd.n3267 gnd.n3266 0.00797283
R14233 gnd.n3269 gnd.n3268 0.00797283
R14234 gnd.n3271 gnd.n2763 0.00797283
R14235 gnd.n3274 gnd.n2764 0.00797283
R14236 gnd.n3276 gnd.n2765 0.00797283
R14237 gnd.n3279 gnd.n3277 0.00797283
R14238 gnd.n3278 gnd.n2664 0.00797283
R14239 gnd.n3346 gnd.n3344 0.00797283
R14240 gnd.n3345 gnd.n2657 0.00797283
R14241 gnd.n3356 gnd.n3355 0.00797283
R14242 gnd.n3358 gnd.n3357 0.00797283
R14243 gnd.n3361 gnd.n2655 0.00797283
R14244 gnd.n3365 gnd.n3364 0.00797283
R14245 gnd.n3363 gnd.n3362 0.00797283
R14246 gnd.n2635 gnd.n2634 0.00797283
R14247 gnd.n3387 gnd.n3386 0.00797283
R14248 gnd.n2636 gnd.n2609 0.00797283
R14249 gnd.n3431 gnd.n3429 0.00797283
R14250 gnd.n3430 gnd.n2602 0.00797283
R14251 gnd.n3441 gnd.n3440 0.00797283
R14252 gnd.n3443 gnd.n3442 0.00797283
R14253 gnd.n3446 gnd.n2600 0.00797283
R14254 gnd.n3450 gnd.n3449 0.00797283
R14255 gnd.n3448 gnd.n3447 0.00797283
R14256 gnd.n2580 gnd.n2579 0.00797283
R14257 gnd.n3472 gnd.n3471 0.00797283
R14258 gnd.n2581 gnd.n2555 0.00797283
R14259 gnd.n3520 gnd.n3518 0.00797283
R14260 gnd.n3519 gnd.n2548 0.00797283
R14261 gnd.n3530 gnd.n3529 0.00797283
R14262 gnd.n3788 gnd.n3787 0.00797283
R14263 gnd.n3791 gnd.n2546 0.00797283
R14264 gnd.n3793 gnd.n3792 0.00797283
R14265 gnd.n3816 gnd.n2527 0.00797283
R14266 gnd.n3817 gnd.n2491 0.00797283
R14267 gnd.n6168 gnd.n6167 0.00593478
R14268 gnd.n5203 gnd.n1753 0.00593478
R14269 vdd.n327 vdd.n291 756.745
R14270 vdd.n268 vdd.n232 756.745
R14271 vdd.n225 vdd.n189 756.745
R14272 vdd.n166 vdd.n130 756.745
R14273 vdd.n124 vdd.n88 756.745
R14274 vdd.n65 vdd.n29 756.745
R14275 vdd.n1746 vdd.n1710 756.745
R14276 vdd.n1805 vdd.n1769 756.745
R14277 vdd.n1644 vdd.n1608 756.745
R14278 vdd.n1703 vdd.n1667 756.745
R14279 vdd.n1543 vdd.n1507 756.745
R14280 vdd.n1602 vdd.n1566 756.745
R14281 vdd.n2177 vdd.t108 640.208
R14282 vdd.n965 vdd.t93 640.208
R14283 vdd.n2151 vdd.t54 640.208
R14284 vdd.n957 vdd.t118 640.208
R14285 vdd.n2922 vdd.t69 640.208
R14286 vdd.n2642 vdd.t115 640.208
R14287 vdd.n832 vdd.t97 640.208
R14288 vdd.n2639 vdd.t101 640.208
R14289 vdd.n799 vdd.t105 640.208
R14290 vdd.n1027 vdd.t111 640.208
R14291 vdd.n1317 vdd.t84 592.009
R14292 vdd.n1355 vdd.t73 592.009
R14293 vdd.n1251 vdd.t87 592.009
R14294 vdd.n2333 vdd.t65 592.009
R14295 vdd.n1970 vdd.t77 592.009
R14296 vdd.n1930 vdd.t90 592.009
R14297 vdd.n426 vdd.t80 592.009
R14298 vdd.n440 vdd.t121 592.009
R14299 vdd.n452 vdd.t127 592.009
R14300 vdd.n768 vdd.t58 592.009
R14301 vdd.n3184 vdd.t62 592.009
R14302 vdd.n688 vdd.t124 592.009
R14303 vdd.n328 vdd.n327 585
R14304 vdd.n326 vdd.n293 585
R14305 vdd.n325 vdd.n324 585
R14306 vdd.n296 vdd.n294 585
R14307 vdd.n319 vdd.n318 585
R14308 vdd.n317 vdd.n316 585
R14309 vdd.n300 vdd.n299 585
R14310 vdd.n311 vdd.n310 585
R14311 vdd.n309 vdd.n308 585
R14312 vdd.n304 vdd.n303 585
R14313 vdd.n269 vdd.n268 585
R14314 vdd.n267 vdd.n234 585
R14315 vdd.n266 vdd.n265 585
R14316 vdd.n237 vdd.n235 585
R14317 vdd.n260 vdd.n259 585
R14318 vdd.n258 vdd.n257 585
R14319 vdd.n241 vdd.n240 585
R14320 vdd.n252 vdd.n251 585
R14321 vdd.n250 vdd.n249 585
R14322 vdd.n245 vdd.n244 585
R14323 vdd.n226 vdd.n225 585
R14324 vdd.n224 vdd.n191 585
R14325 vdd.n223 vdd.n222 585
R14326 vdd.n194 vdd.n192 585
R14327 vdd.n217 vdd.n216 585
R14328 vdd.n215 vdd.n214 585
R14329 vdd.n198 vdd.n197 585
R14330 vdd.n209 vdd.n208 585
R14331 vdd.n207 vdd.n206 585
R14332 vdd.n202 vdd.n201 585
R14333 vdd.n167 vdd.n166 585
R14334 vdd.n165 vdd.n132 585
R14335 vdd.n164 vdd.n163 585
R14336 vdd.n135 vdd.n133 585
R14337 vdd.n158 vdd.n157 585
R14338 vdd.n156 vdd.n155 585
R14339 vdd.n139 vdd.n138 585
R14340 vdd.n150 vdd.n149 585
R14341 vdd.n148 vdd.n147 585
R14342 vdd.n143 vdd.n142 585
R14343 vdd.n125 vdd.n124 585
R14344 vdd.n123 vdd.n90 585
R14345 vdd.n122 vdd.n121 585
R14346 vdd.n93 vdd.n91 585
R14347 vdd.n116 vdd.n115 585
R14348 vdd.n114 vdd.n113 585
R14349 vdd.n97 vdd.n96 585
R14350 vdd.n108 vdd.n107 585
R14351 vdd.n106 vdd.n105 585
R14352 vdd.n101 vdd.n100 585
R14353 vdd.n66 vdd.n65 585
R14354 vdd.n64 vdd.n31 585
R14355 vdd.n63 vdd.n62 585
R14356 vdd.n34 vdd.n32 585
R14357 vdd.n57 vdd.n56 585
R14358 vdd.n55 vdd.n54 585
R14359 vdd.n38 vdd.n37 585
R14360 vdd.n49 vdd.n48 585
R14361 vdd.n47 vdd.n46 585
R14362 vdd.n42 vdd.n41 585
R14363 vdd.n1747 vdd.n1746 585
R14364 vdd.n1745 vdd.n1712 585
R14365 vdd.n1744 vdd.n1743 585
R14366 vdd.n1715 vdd.n1713 585
R14367 vdd.n1738 vdd.n1737 585
R14368 vdd.n1736 vdd.n1735 585
R14369 vdd.n1719 vdd.n1718 585
R14370 vdd.n1730 vdd.n1729 585
R14371 vdd.n1728 vdd.n1727 585
R14372 vdd.n1723 vdd.n1722 585
R14373 vdd.n1806 vdd.n1805 585
R14374 vdd.n1804 vdd.n1771 585
R14375 vdd.n1803 vdd.n1802 585
R14376 vdd.n1774 vdd.n1772 585
R14377 vdd.n1797 vdd.n1796 585
R14378 vdd.n1795 vdd.n1794 585
R14379 vdd.n1778 vdd.n1777 585
R14380 vdd.n1789 vdd.n1788 585
R14381 vdd.n1787 vdd.n1786 585
R14382 vdd.n1782 vdd.n1781 585
R14383 vdd.n1645 vdd.n1644 585
R14384 vdd.n1643 vdd.n1610 585
R14385 vdd.n1642 vdd.n1641 585
R14386 vdd.n1613 vdd.n1611 585
R14387 vdd.n1636 vdd.n1635 585
R14388 vdd.n1634 vdd.n1633 585
R14389 vdd.n1617 vdd.n1616 585
R14390 vdd.n1628 vdd.n1627 585
R14391 vdd.n1626 vdd.n1625 585
R14392 vdd.n1621 vdd.n1620 585
R14393 vdd.n1704 vdd.n1703 585
R14394 vdd.n1702 vdd.n1669 585
R14395 vdd.n1701 vdd.n1700 585
R14396 vdd.n1672 vdd.n1670 585
R14397 vdd.n1695 vdd.n1694 585
R14398 vdd.n1693 vdd.n1692 585
R14399 vdd.n1676 vdd.n1675 585
R14400 vdd.n1687 vdd.n1686 585
R14401 vdd.n1685 vdd.n1684 585
R14402 vdd.n1680 vdd.n1679 585
R14403 vdd.n1544 vdd.n1543 585
R14404 vdd.n1542 vdd.n1509 585
R14405 vdd.n1541 vdd.n1540 585
R14406 vdd.n1512 vdd.n1510 585
R14407 vdd.n1535 vdd.n1534 585
R14408 vdd.n1533 vdd.n1532 585
R14409 vdd.n1516 vdd.n1515 585
R14410 vdd.n1527 vdd.n1526 585
R14411 vdd.n1525 vdd.n1524 585
R14412 vdd.n1520 vdd.n1519 585
R14413 vdd.n1603 vdd.n1602 585
R14414 vdd.n1601 vdd.n1568 585
R14415 vdd.n1600 vdd.n1599 585
R14416 vdd.n1571 vdd.n1569 585
R14417 vdd.n1594 vdd.n1593 585
R14418 vdd.n1592 vdd.n1591 585
R14419 vdd.n1575 vdd.n1574 585
R14420 vdd.n1586 vdd.n1585 585
R14421 vdd.n1584 vdd.n1583 585
R14422 vdd.n1579 vdd.n1578 585
R14423 vdd.n3356 vdd.n392 509.269
R14424 vdd.n3352 vdd.n393 509.269
R14425 vdd.n3224 vdd.n685 509.269
R14426 vdd.n3221 vdd.n684 509.269
R14427 vdd.n2328 vdd.n1075 509.269
R14428 vdd.n2331 vdd.n2330 509.269
R14429 vdd.n1224 vdd.n1188 509.269
R14430 vdd.n1420 vdd.n1189 509.269
R14431 vdd.n305 vdd.t263 329.043
R14432 vdd.n246 vdd.t240 329.043
R14433 vdd.n203 vdd.t252 329.043
R14434 vdd.n144 vdd.t224 329.043
R14435 vdd.n102 vdd.t203 329.043
R14436 vdd.n43 vdd.t141 329.043
R14437 vdd.n1724 vdd.t283 329.043
R14438 vdd.n1783 vdd.t172 329.043
R14439 vdd.n1622 vdd.t269 329.043
R14440 vdd.n1681 vdd.t149 329.043
R14441 vdd.n1521 vdd.t145 329.043
R14442 vdd.n1580 vdd.t204 329.043
R14443 vdd.n1317 vdd.t86 319.788
R14444 vdd.n1355 vdd.t76 319.788
R14445 vdd.n1251 vdd.t89 319.788
R14446 vdd.n2333 vdd.t67 319.788
R14447 vdd.n1970 vdd.t78 319.788
R14448 vdd.n1930 vdd.t91 319.788
R14449 vdd.n426 vdd.t82 319.788
R14450 vdd.n440 vdd.t122 319.788
R14451 vdd.n452 vdd.t128 319.788
R14452 vdd.n768 vdd.t61 319.788
R14453 vdd.n3184 vdd.t64 319.788
R14454 vdd.n688 vdd.t126 319.788
R14455 vdd.n1318 vdd.t85 303.69
R14456 vdd.n1356 vdd.t75 303.69
R14457 vdd.n1252 vdd.t88 303.69
R14458 vdd.n2334 vdd.t68 303.69
R14459 vdd.n1971 vdd.t79 303.69
R14460 vdd.n1931 vdd.t92 303.69
R14461 vdd.n427 vdd.t83 303.69
R14462 vdd.n441 vdd.t123 303.69
R14463 vdd.n453 vdd.t129 303.69
R14464 vdd.n769 vdd.t60 303.69
R14465 vdd.n3185 vdd.t63 303.69
R14466 vdd.n689 vdd.t125 303.69
R14467 vdd.n2865 vdd.n913 297.074
R14468 vdd.n3058 vdd.n809 297.074
R14469 vdd.n2995 vdd.n806 297.074
R14470 vdd.n2788 vdd.n914 297.074
R14471 vdd.n2603 vdd.n954 297.074
R14472 vdd.n2534 vdd.n2533 297.074
R14473 vdd.n2280 vdd.n1050 297.074
R14474 vdd.n2376 vdd.n1048 297.074
R14475 vdd.n2974 vdd.n807 297.074
R14476 vdd.n3061 vdd.n3060 297.074
R14477 vdd.n2637 vdd.n915 297.074
R14478 vdd.n2863 vdd.n916 297.074
R14479 vdd.n2531 vdd.n963 297.074
R14480 vdd.n961 vdd.n936 297.074
R14481 vdd.n2217 vdd.n1051 297.074
R14482 vdd.n2374 vdd.n1052 297.074
R14483 vdd.n2976 vdd.n807 185
R14484 vdd.n3059 vdd.n807 185
R14485 vdd.n2978 vdd.n2977 185
R14486 vdd.n2977 vdd.n805 185
R14487 vdd.n2979 vdd.n839 185
R14488 vdd.n2989 vdd.n839 185
R14489 vdd.n2980 vdd.n848 185
R14490 vdd.n848 vdd.n846 185
R14491 vdd.n2982 vdd.n2981 185
R14492 vdd.n2983 vdd.n2982 185
R14493 vdd.n2935 vdd.n847 185
R14494 vdd.n847 vdd.n843 185
R14495 vdd.n2934 vdd.n2933 185
R14496 vdd.n2933 vdd.n2932 185
R14497 vdd.n850 vdd.n849 185
R14498 vdd.n851 vdd.n850 185
R14499 vdd.n2925 vdd.n2924 185
R14500 vdd.n2926 vdd.n2925 185
R14501 vdd.n2921 vdd.n860 185
R14502 vdd.n860 vdd.n857 185
R14503 vdd.n2920 vdd.n2919 185
R14504 vdd.n2919 vdd.n2918 185
R14505 vdd.n862 vdd.n861 185
R14506 vdd.n870 vdd.n862 185
R14507 vdd.n2911 vdd.n2910 185
R14508 vdd.n2912 vdd.n2911 185
R14509 vdd.n2909 vdd.n871 185
R14510 vdd.n2760 vdd.n871 185
R14511 vdd.n2908 vdd.n2907 185
R14512 vdd.n2907 vdd.n2906 185
R14513 vdd.n873 vdd.n872 185
R14514 vdd.n874 vdd.n873 185
R14515 vdd.n2899 vdd.n2898 185
R14516 vdd.n2900 vdd.n2899 185
R14517 vdd.n2897 vdd.n883 185
R14518 vdd.n883 vdd.n880 185
R14519 vdd.n2896 vdd.n2895 185
R14520 vdd.n2895 vdd.n2894 185
R14521 vdd.n885 vdd.n884 185
R14522 vdd.n893 vdd.n885 185
R14523 vdd.n2887 vdd.n2886 185
R14524 vdd.n2888 vdd.n2887 185
R14525 vdd.n2885 vdd.n894 185
R14526 vdd.n900 vdd.n894 185
R14527 vdd.n2884 vdd.n2883 185
R14528 vdd.n2883 vdd.n2882 185
R14529 vdd.n896 vdd.n895 185
R14530 vdd.n897 vdd.n896 185
R14531 vdd.n2875 vdd.n2874 185
R14532 vdd.n2876 vdd.n2875 185
R14533 vdd.n2873 vdd.n906 185
R14534 vdd.n2781 vdd.n906 185
R14535 vdd.n2872 vdd.n2871 185
R14536 vdd.n2871 vdd.n2870 185
R14537 vdd.n908 vdd.n907 185
R14538 vdd.t132 vdd.n908 185
R14539 vdd.n2863 vdd.n2862 185
R14540 vdd.n2864 vdd.n2863 185
R14541 vdd.n2861 vdd.n916 185
R14542 vdd.n2860 vdd.n2859 185
R14543 vdd.n918 vdd.n917 185
R14544 vdd.n2646 vdd.n2645 185
R14545 vdd.n2648 vdd.n2647 185
R14546 vdd.n2650 vdd.n2649 185
R14547 vdd.n2652 vdd.n2651 185
R14548 vdd.n2654 vdd.n2653 185
R14549 vdd.n2656 vdd.n2655 185
R14550 vdd.n2658 vdd.n2657 185
R14551 vdd.n2660 vdd.n2659 185
R14552 vdd.n2662 vdd.n2661 185
R14553 vdd.n2664 vdd.n2663 185
R14554 vdd.n2666 vdd.n2665 185
R14555 vdd.n2668 vdd.n2667 185
R14556 vdd.n2670 vdd.n2669 185
R14557 vdd.n2672 vdd.n2671 185
R14558 vdd.n2674 vdd.n2673 185
R14559 vdd.n2676 vdd.n2675 185
R14560 vdd.n2678 vdd.n2677 185
R14561 vdd.n2680 vdd.n2679 185
R14562 vdd.n2682 vdd.n2681 185
R14563 vdd.n2684 vdd.n2683 185
R14564 vdd.n2686 vdd.n2685 185
R14565 vdd.n2688 vdd.n2687 185
R14566 vdd.n2690 vdd.n2689 185
R14567 vdd.n2692 vdd.n2691 185
R14568 vdd.n2694 vdd.n2693 185
R14569 vdd.n2696 vdd.n2695 185
R14570 vdd.n2698 vdd.n2697 185
R14571 vdd.n2700 vdd.n2699 185
R14572 vdd.n2702 vdd.n2701 185
R14573 vdd.n2704 vdd.n2703 185
R14574 vdd.n2706 vdd.n2705 185
R14575 vdd.n2707 vdd.n2637 185
R14576 vdd.n2857 vdd.n2637 185
R14577 vdd.n3062 vdd.n3061 185
R14578 vdd.n3063 vdd.n798 185
R14579 vdd.n3065 vdd.n3064 185
R14580 vdd.n3067 vdd.n796 185
R14581 vdd.n3069 vdd.n3068 185
R14582 vdd.n3070 vdd.n795 185
R14583 vdd.n3072 vdd.n3071 185
R14584 vdd.n3074 vdd.n793 185
R14585 vdd.n3076 vdd.n3075 185
R14586 vdd.n3077 vdd.n792 185
R14587 vdd.n3079 vdd.n3078 185
R14588 vdd.n3081 vdd.n790 185
R14589 vdd.n3083 vdd.n3082 185
R14590 vdd.n3084 vdd.n789 185
R14591 vdd.n3086 vdd.n3085 185
R14592 vdd.n3088 vdd.n788 185
R14593 vdd.n3089 vdd.n786 185
R14594 vdd.n3092 vdd.n3091 185
R14595 vdd.n787 vdd.n785 185
R14596 vdd.n2948 vdd.n2947 185
R14597 vdd.n2950 vdd.n2949 185
R14598 vdd.n2952 vdd.n2944 185
R14599 vdd.n2954 vdd.n2953 185
R14600 vdd.n2955 vdd.n2943 185
R14601 vdd.n2957 vdd.n2956 185
R14602 vdd.n2959 vdd.n2941 185
R14603 vdd.n2961 vdd.n2960 185
R14604 vdd.n2962 vdd.n2940 185
R14605 vdd.n2964 vdd.n2963 185
R14606 vdd.n2966 vdd.n2938 185
R14607 vdd.n2968 vdd.n2967 185
R14608 vdd.n2969 vdd.n2937 185
R14609 vdd.n2971 vdd.n2970 185
R14610 vdd.n2973 vdd.n2936 185
R14611 vdd.n2975 vdd.n2974 185
R14612 vdd.n2974 vdd.n692 185
R14613 vdd.n3060 vdd.n802 185
R14614 vdd.n3060 vdd.n3059 185
R14615 vdd.n2712 vdd.n804 185
R14616 vdd.n805 vdd.n804 185
R14617 vdd.n2713 vdd.n838 185
R14618 vdd.n2989 vdd.n838 185
R14619 vdd.n2715 vdd.n2714 185
R14620 vdd.n2714 vdd.n846 185
R14621 vdd.n2716 vdd.n845 185
R14622 vdd.n2983 vdd.n845 185
R14623 vdd.n2718 vdd.n2717 185
R14624 vdd.n2717 vdd.n843 185
R14625 vdd.n2719 vdd.n853 185
R14626 vdd.n2932 vdd.n853 185
R14627 vdd.n2721 vdd.n2720 185
R14628 vdd.n2720 vdd.n851 185
R14629 vdd.n2722 vdd.n859 185
R14630 vdd.n2926 vdd.n859 185
R14631 vdd.n2724 vdd.n2723 185
R14632 vdd.n2723 vdd.n857 185
R14633 vdd.n2725 vdd.n864 185
R14634 vdd.n2918 vdd.n864 185
R14635 vdd.n2727 vdd.n2726 185
R14636 vdd.n2726 vdd.n870 185
R14637 vdd.n2728 vdd.n869 185
R14638 vdd.n2912 vdd.n869 185
R14639 vdd.n2762 vdd.n2761 185
R14640 vdd.n2761 vdd.n2760 185
R14641 vdd.n2763 vdd.n876 185
R14642 vdd.n2906 vdd.n876 185
R14643 vdd.n2765 vdd.n2764 185
R14644 vdd.n2764 vdd.n874 185
R14645 vdd.n2766 vdd.n882 185
R14646 vdd.n2900 vdd.n882 185
R14647 vdd.n2768 vdd.n2767 185
R14648 vdd.n2767 vdd.n880 185
R14649 vdd.n2769 vdd.n887 185
R14650 vdd.n2894 vdd.n887 185
R14651 vdd.n2771 vdd.n2770 185
R14652 vdd.n2770 vdd.n893 185
R14653 vdd.n2772 vdd.n892 185
R14654 vdd.n2888 vdd.n892 185
R14655 vdd.n2774 vdd.n2773 185
R14656 vdd.n2773 vdd.n900 185
R14657 vdd.n2775 vdd.n899 185
R14658 vdd.n2882 vdd.n899 185
R14659 vdd.n2777 vdd.n2776 185
R14660 vdd.n2776 vdd.n897 185
R14661 vdd.n2778 vdd.n905 185
R14662 vdd.n2876 vdd.n905 185
R14663 vdd.n2780 vdd.n2779 185
R14664 vdd.n2781 vdd.n2780 185
R14665 vdd.n2711 vdd.n910 185
R14666 vdd.n2870 vdd.n910 185
R14667 vdd.n2710 vdd.n2709 185
R14668 vdd.n2709 vdd.t132 185
R14669 vdd.n2708 vdd.n915 185
R14670 vdd.n2864 vdd.n915 185
R14671 vdd.n2328 vdd.n2327 185
R14672 vdd.n2329 vdd.n2328 185
R14673 vdd.n1076 vdd.n1074 185
R14674 vdd.n1894 vdd.n1074 185
R14675 vdd.n1897 vdd.n1896 185
R14676 vdd.n1896 vdd.n1895 185
R14677 vdd.n1079 vdd.n1078 185
R14678 vdd.n1080 vdd.n1079 185
R14679 vdd.n1883 vdd.n1882 185
R14680 vdd.n1884 vdd.n1883 185
R14681 vdd.n1088 vdd.n1087 185
R14682 vdd.n1875 vdd.n1087 185
R14683 vdd.n1878 vdd.n1877 185
R14684 vdd.n1877 vdd.n1876 185
R14685 vdd.n1091 vdd.n1090 185
R14686 vdd.n1098 vdd.n1091 185
R14687 vdd.n1866 vdd.n1865 185
R14688 vdd.n1867 vdd.n1866 185
R14689 vdd.n1100 vdd.n1099 185
R14690 vdd.n1099 vdd.n1097 185
R14691 vdd.n1861 vdd.n1860 185
R14692 vdd.n1860 vdd.n1859 185
R14693 vdd.n1103 vdd.n1102 185
R14694 vdd.n1104 vdd.n1103 185
R14695 vdd.n1850 vdd.n1849 185
R14696 vdd.n1851 vdd.n1850 185
R14697 vdd.n1111 vdd.n1110 185
R14698 vdd.n1842 vdd.n1110 185
R14699 vdd.n1845 vdd.n1844 185
R14700 vdd.n1844 vdd.n1843 185
R14701 vdd.n1114 vdd.n1113 185
R14702 vdd.n1120 vdd.n1114 185
R14703 vdd.n1833 vdd.n1832 185
R14704 vdd.n1834 vdd.n1833 185
R14705 vdd.n1122 vdd.n1121 185
R14706 vdd.n1825 vdd.n1121 185
R14707 vdd.n1828 vdd.n1827 185
R14708 vdd.n1827 vdd.n1826 185
R14709 vdd.n1125 vdd.n1124 185
R14710 vdd.n1126 vdd.n1125 185
R14711 vdd.n1816 vdd.n1815 185
R14712 vdd.n1817 vdd.n1816 185
R14713 vdd.n1134 vdd.n1133 185
R14714 vdd.n1133 vdd.n1132 185
R14715 vdd.n1504 vdd.n1503 185
R14716 vdd.n1503 vdd.n1502 185
R14717 vdd.n1137 vdd.n1136 185
R14718 vdd.n1143 vdd.n1137 185
R14719 vdd.n1493 vdd.n1492 185
R14720 vdd.n1494 vdd.n1493 185
R14721 vdd.n1145 vdd.n1144 185
R14722 vdd.n1485 vdd.n1144 185
R14723 vdd.n1488 vdd.n1487 185
R14724 vdd.n1487 vdd.n1486 185
R14725 vdd.n1148 vdd.n1147 185
R14726 vdd.n1155 vdd.n1148 185
R14727 vdd.n1476 vdd.n1475 185
R14728 vdd.n1477 vdd.n1476 185
R14729 vdd.n1157 vdd.n1156 185
R14730 vdd.n1156 vdd.n1154 185
R14731 vdd.n1471 vdd.n1470 185
R14732 vdd.n1470 vdd.n1469 185
R14733 vdd.n1160 vdd.n1159 185
R14734 vdd.n1161 vdd.n1160 185
R14735 vdd.n1460 vdd.n1459 185
R14736 vdd.n1461 vdd.n1460 185
R14737 vdd.n1168 vdd.n1167 185
R14738 vdd.n1452 vdd.n1167 185
R14739 vdd.n1455 vdd.n1454 185
R14740 vdd.n1454 vdd.n1453 185
R14741 vdd.n1171 vdd.n1170 185
R14742 vdd.n1177 vdd.n1171 185
R14743 vdd.n1443 vdd.n1442 185
R14744 vdd.n1444 vdd.n1443 185
R14745 vdd.n1179 vdd.n1178 185
R14746 vdd.n1435 vdd.n1178 185
R14747 vdd.n1438 vdd.n1437 185
R14748 vdd.n1437 vdd.n1436 185
R14749 vdd.n1182 vdd.n1181 185
R14750 vdd.n1183 vdd.n1182 185
R14751 vdd.n1426 vdd.n1425 185
R14752 vdd.n1427 vdd.n1426 185
R14753 vdd.n1190 vdd.n1189 185
R14754 vdd.n1225 vdd.n1189 185
R14755 vdd.n1421 vdd.n1420 185
R14756 vdd.n1193 vdd.n1192 185
R14757 vdd.n1417 vdd.n1416 185
R14758 vdd.n1418 vdd.n1417 185
R14759 vdd.n1227 vdd.n1226 185
R14760 vdd.n1412 vdd.n1229 185
R14761 vdd.n1411 vdd.n1230 185
R14762 vdd.n1410 vdd.n1231 185
R14763 vdd.n1233 vdd.n1232 185
R14764 vdd.n1406 vdd.n1235 185
R14765 vdd.n1405 vdd.n1236 185
R14766 vdd.n1404 vdd.n1237 185
R14767 vdd.n1239 vdd.n1238 185
R14768 vdd.n1400 vdd.n1241 185
R14769 vdd.n1399 vdd.n1242 185
R14770 vdd.n1398 vdd.n1243 185
R14771 vdd.n1245 vdd.n1244 185
R14772 vdd.n1394 vdd.n1247 185
R14773 vdd.n1393 vdd.n1248 185
R14774 vdd.n1392 vdd.n1249 185
R14775 vdd.n1253 vdd.n1250 185
R14776 vdd.n1388 vdd.n1255 185
R14777 vdd.n1387 vdd.n1256 185
R14778 vdd.n1386 vdd.n1257 185
R14779 vdd.n1259 vdd.n1258 185
R14780 vdd.n1382 vdd.n1261 185
R14781 vdd.n1381 vdd.n1262 185
R14782 vdd.n1380 vdd.n1263 185
R14783 vdd.n1265 vdd.n1264 185
R14784 vdd.n1376 vdd.n1267 185
R14785 vdd.n1375 vdd.n1268 185
R14786 vdd.n1374 vdd.n1269 185
R14787 vdd.n1271 vdd.n1270 185
R14788 vdd.n1370 vdd.n1273 185
R14789 vdd.n1369 vdd.n1274 185
R14790 vdd.n1368 vdd.n1275 185
R14791 vdd.n1277 vdd.n1276 185
R14792 vdd.n1364 vdd.n1279 185
R14793 vdd.n1363 vdd.n1280 185
R14794 vdd.n1362 vdd.n1281 185
R14795 vdd.n1283 vdd.n1282 185
R14796 vdd.n1358 vdd.n1285 185
R14797 vdd.n1357 vdd.n1354 185
R14798 vdd.n1353 vdd.n1286 185
R14799 vdd.n1288 vdd.n1287 185
R14800 vdd.n1349 vdd.n1290 185
R14801 vdd.n1348 vdd.n1291 185
R14802 vdd.n1347 vdd.n1292 185
R14803 vdd.n1294 vdd.n1293 185
R14804 vdd.n1343 vdd.n1296 185
R14805 vdd.n1342 vdd.n1297 185
R14806 vdd.n1341 vdd.n1298 185
R14807 vdd.n1300 vdd.n1299 185
R14808 vdd.n1337 vdd.n1302 185
R14809 vdd.n1336 vdd.n1303 185
R14810 vdd.n1335 vdd.n1304 185
R14811 vdd.n1306 vdd.n1305 185
R14812 vdd.n1331 vdd.n1308 185
R14813 vdd.n1330 vdd.n1309 185
R14814 vdd.n1329 vdd.n1310 185
R14815 vdd.n1312 vdd.n1311 185
R14816 vdd.n1325 vdd.n1314 185
R14817 vdd.n1324 vdd.n1315 185
R14818 vdd.n1323 vdd.n1316 185
R14819 vdd.n1320 vdd.n1224 185
R14820 vdd.n1418 vdd.n1224 185
R14821 vdd.n2332 vdd.n2331 185
R14822 vdd.n2336 vdd.n1069 185
R14823 vdd.n1999 vdd.n1068 185
R14824 vdd.n2002 vdd.n2001 185
R14825 vdd.n2004 vdd.n2003 185
R14826 vdd.n2007 vdd.n2006 185
R14827 vdd.n2009 vdd.n2008 185
R14828 vdd.n2011 vdd.n1997 185
R14829 vdd.n2013 vdd.n2012 185
R14830 vdd.n2014 vdd.n1991 185
R14831 vdd.n2016 vdd.n2015 185
R14832 vdd.n2018 vdd.n1989 185
R14833 vdd.n2020 vdd.n2019 185
R14834 vdd.n2021 vdd.n1984 185
R14835 vdd.n2023 vdd.n2022 185
R14836 vdd.n2025 vdd.n1982 185
R14837 vdd.n2027 vdd.n2026 185
R14838 vdd.n2028 vdd.n1978 185
R14839 vdd.n2030 vdd.n2029 185
R14840 vdd.n2032 vdd.n1975 185
R14841 vdd.n2034 vdd.n2033 185
R14842 vdd.n1976 vdd.n1969 185
R14843 vdd.n2038 vdd.n1973 185
R14844 vdd.n2039 vdd.n1965 185
R14845 vdd.n2041 vdd.n2040 185
R14846 vdd.n2043 vdd.n1963 185
R14847 vdd.n2045 vdd.n2044 185
R14848 vdd.n2046 vdd.n1958 185
R14849 vdd.n2048 vdd.n2047 185
R14850 vdd.n2050 vdd.n1956 185
R14851 vdd.n2052 vdd.n2051 185
R14852 vdd.n2053 vdd.n1951 185
R14853 vdd.n2055 vdd.n2054 185
R14854 vdd.n2057 vdd.n1949 185
R14855 vdd.n2059 vdd.n2058 185
R14856 vdd.n2060 vdd.n1944 185
R14857 vdd.n2062 vdd.n2061 185
R14858 vdd.n2064 vdd.n1942 185
R14859 vdd.n2066 vdd.n2065 185
R14860 vdd.n2067 vdd.n1938 185
R14861 vdd.n2069 vdd.n2068 185
R14862 vdd.n2071 vdd.n1935 185
R14863 vdd.n2073 vdd.n2072 185
R14864 vdd.n1936 vdd.n1929 185
R14865 vdd.n2077 vdd.n1933 185
R14866 vdd.n2078 vdd.n1925 185
R14867 vdd.n2080 vdd.n2079 185
R14868 vdd.n2082 vdd.n1923 185
R14869 vdd.n2084 vdd.n2083 185
R14870 vdd.n2085 vdd.n1918 185
R14871 vdd.n2087 vdd.n2086 185
R14872 vdd.n2089 vdd.n1916 185
R14873 vdd.n2091 vdd.n2090 185
R14874 vdd.n2092 vdd.n1911 185
R14875 vdd.n2094 vdd.n2093 185
R14876 vdd.n2096 vdd.n1910 185
R14877 vdd.n2097 vdd.n1907 185
R14878 vdd.n2100 vdd.n2099 185
R14879 vdd.n1909 vdd.n1905 185
R14880 vdd.n2317 vdd.n1903 185
R14881 vdd.n2319 vdd.n2318 185
R14882 vdd.n2321 vdd.n1901 185
R14883 vdd.n2323 vdd.n2322 185
R14884 vdd.n2324 vdd.n1075 185
R14885 vdd.n2330 vdd.n1072 185
R14886 vdd.n2330 vdd.n2329 185
R14887 vdd.n1083 vdd.n1071 185
R14888 vdd.n1894 vdd.n1071 185
R14889 vdd.n1893 vdd.n1892 185
R14890 vdd.n1895 vdd.n1893 185
R14891 vdd.n1082 vdd.n1081 185
R14892 vdd.n1081 vdd.n1080 185
R14893 vdd.n1886 vdd.n1885 185
R14894 vdd.n1885 vdd.n1884 185
R14895 vdd.n1086 vdd.n1085 185
R14896 vdd.n1875 vdd.n1086 185
R14897 vdd.n1874 vdd.n1873 185
R14898 vdd.n1876 vdd.n1874 185
R14899 vdd.n1093 vdd.n1092 185
R14900 vdd.n1098 vdd.n1092 185
R14901 vdd.n1869 vdd.n1868 185
R14902 vdd.n1868 vdd.n1867 185
R14903 vdd.n1096 vdd.n1095 185
R14904 vdd.n1097 vdd.n1096 185
R14905 vdd.n1858 vdd.n1857 185
R14906 vdd.n1859 vdd.n1858 185
R14907 vdd.n1106 vdd.n1105 185
R14908 vdd.n1105 vdd.n1104 185
R14909 vdd.n1853 vdd.n1852 185
R14910 vdd.n1852 vdd.n1851 185
R14911 vdd.n1109 vdd.n1108 185
R14912 vdd.n1842 vdd.n1109 185
R14913 vdd.n1841 vdd.n1840 185
R14914 vdd.n1843 vdd.n1841 185
R14915 vdd.n1116 vdd.n1115 185
R14916 vdd.n1120 vdd.n1115 185
R14917 vdd.n1836 vdd.n1835 185
R14918 vdd.n1835 vdd.n1834 185
R14919 vdd.n1119 vdd.n1118 185
R14920 vdd.n1825 vdd.n1119 185
R14921 vdd.n1824 vdd.n1823 185
R14922 vdd.n1826 vdd.n1824 185
R14923 vdd.n1128 vdd.n1127 185
R14924 vdd.n1127 vdd.n1126 185
R14925 vdd.n1819 vdd.n1818 185
R14926 vdd.n1818 vdd.n1817 185
R14927 vdd.n1131 vdd.n1130 185
R14928 vdd.n1132 vdd.n1131 185
R14929 vdd.n1501 vdd.n1500 185
R14930 vdd.n1502 vdd.n1501 185
R14931 vdd.n1139 vdd.n1138 185
R14932 vdd.n1143 vdd.n1138 185
R14933 vdd.n1496 vdd.n1495 185
R14934 vdd.n1495 vdd.n1494 185
R14935 vdd.n1142 vdd.n1141 185
R14936 vdd.n1485 vdd.n1142 185
R14937 vdd.n1484 vdd.n1483 185
R14938 vdd.n1486 vdd.n1484 185
R14939 vdd.n1150 vdd.n1149 185
R14940 vdd.n1155 vdd.n1149 185
R14941 vdd.n1479 vdd.n1478 185
R14942 vdd.n1478 vdd.n1477 185
R14943 vdd.n1153 vdd.n1152 185
R14944 vdd.n1154 vdd.n1153 185
R14945 vdd.n1468 vdd.n1467 185
R14946 vdd.n1469 vdd.n1468 185
R14947 vdd.n1163 vdd.n1162 185
R14948 vdd.n1162 vdd.n1161 185
R14949 vdd.n1463 vdd.n1462 185
R14950 vdd.n1462 vdd.n1461 185
R14951 vdd.n1166 vdd.n1165 185
R14952 vdd.n1452 vdd.n1166 185
R14953 vdd.n1451 vdd.n1450 185
R14954 vdd.n1453 vdd.n1451 185
R14955 vdd.n1173 vdd.n1172 185
R14956 vdd.n1177 vdd.n1172 185
R14957 vdd.n1446 vdd.n1445 185
R14958 vdd.n1445 vdd.n1444 185
R14959 vdd.n1176 vdd.n1175 185
R14960 vdd.n1435 vdd.n1176 185
R14961 vdd.n1434 vdd.n1433 185
R14962 vdd.n1436 vdd.n1434 185
R14963 vdd.n1185 vdd.n1184 185
R14964 vdd.n1184 vdd.n1183 185
R14965 vdd.n1429 vdd.n1428 185
R14966 vdd.n1428 vdd.n1427 185
R14967 vdd.n1188 vdd.n1187 185
R14968 vdd.n1225 vdd.n1188 185
R14969 vdd.n956 vdd.n954 185
R14970 vdd.n2532 vdd.n954 185
R14971 vdd.n2454 vdd.n973 185
R14972 vdd.n973 vdd.t35 185
R14973 vdd.n2456 vdd.n2455 185
R14974 vdd.n2457 vdd.n2456 185
R14975 vdd.n2453 vdd.n972 185
R14976 vdd.n2156 vdd.n972 185
R14977 vdd.n2452 vdd.n2451 185
R14978 vdd.n2451 vdd.n2450 185
R14979 vdd.n975 vdd.n974 185
R14980 vdd.n976 vdd.n975 185
R14981 vdd.n2441 vdd.n2440 185
R14982 vdd.n2442 vdd.n2441 185
R14983 vdd.n2439 vdd.n986 185
R14984 vdd.n986 vdd.n983 185
R14985 vdd.n2438 vdd.n2437 185
R14986 vdd.n2437 vdd.n2436 185
R14987 vdd.n988 vdd.n987 185
R14988 vdd.n989 vdd.n988 185
R14989 vdd.n2429 vdd.n2428 185
R14990 vdd.n2430 vdd.n2429 185
R14991 vdd.n2427 vdd.n997 185
R14992 vdd.n1002 vdd.n997 185
R14993 vdd.n2426 vdd.n2425 185
R14994 vdd.n2425 vdd.n2424 185
R14995 vdd.n999 vdd.n998 185
R14996 vdd.n1008 vdd.n999 185
R14997 vdd.n2417 vdd.n2416 185
R14998 vdd.n2418 vdd.n2417 185
R14999 vdd.n2415 vdd.n1009 185
R15000 vdd.n2257 vdd.n1009 185
R15001 vdd.n2414 vdd.n2413 185
R15002 vdd.n2413 vdd.n2412 185
R15003 vdd.n1011 vdd.n1010 185
R15004 vdd.n1012 vdd.n1011 185
R15005 vdd.n2405 vdd.n2404 185
R15006 vdd.n2406 vdd.n2405 185
R15007 vdd.n2403 vdd.n1021 185
R15008 vdd.n1021 vdd.n1018 185
R15009 vdd.n2402 vdd.n2401 185
R15010 vdd.n2401 vdd.n2400 185
R15011 vdd.n1023 vdd.n1022 185
R15012 vdd.n1033 vdd.n1023 185
R15013 vdd.n2392 vdd.n2391 185
R15014 vdd.n2393 vdd.n2392 185
R15015 vdd.n2390 vdd.n1034 185
R15016 vdd.n1034 vdd.n1030 185
R15017 vdd.n2389 vdd.n2388 185
R15018 vdd.n2388 vdd.n2387 185
R15019 vdd.n1036 vdd.n1035 185
R15020 vdd.n1037 vdd.n1036 185
R15021 vdd.n2380 vdd.n2379 185
R15022 vdd.n2381 vdd.n2380 185
R15023 vdd.n2378 vdd.n1046 185
R15024 vdd.n1046 vdd.n1043 185
R15025 vdd.n2377 vdd.n2376 185
R15026 vdd.n2376 vdd.n2375 185
R15027 vdd.n1048 vdd.n1047 185
R15028 vdd.n2112 vdd.n2111 185
R15029 vdd.n2113 vdd.n2109 185
R15030 vdd.n2109 vdd.n1049 185
R15031 vdd.n2115 vdd.n2114 185
R15032 vdd.n2117 vdd.n2108 185
R15033 vdd.n2120 vdd.n2119 185
R15034 vdd.n2121 vdd.n2107 185
R15035 vdd.n2123 vdd.n2122 185
R15036 vdd.n2125 vdd.n2106 185
R15037 vdd.n2128 vdd.n2127 185
R15038 vdd.n2129 vdd.n2105 185
R15039 vdd.n2131 vdd.n2130 185
R15040 vdd.n2133 vdd.n2104 185
R15041 vdd.n2136 vdd.n2135 185
R15042 vdd.n2137 vdd.n2103 185
R15043 vdd.n2139 vdd.n2138 185
R15044 vdd.n2141 vdd.n2102 185
R15045 vdd.n2314 vdd.n2142 185
R15046 vdd.n2313 vdd.n2312 185
R15047 vdd.n2310 vdd.n2143 185
R15048 vdd.n2308 vdd.n2307 185
R15049 vdd.n2306 vdd.n2144 185
R15050 vdd.n2305 vdd.n2304 185
R15051 vdd.n2302 vdd.n2145 185
R15052 vdd.n2300 vdd.n2299 185
R15053 vdd.n2298 vdd.n2146 185
R15054 vdd.n2297 vdd.n2296 185
R15055 vdd.n2294 vdd.n2147 185
R15056 vdd.n2292 vdd.n2291 185
R15057 vdd.n2290 vdd.n2148 185
R15058 vdd.n2289 vdd.n2288 185
R15059 vdd.n2286 vdd.n2149 185
R15060 vdd.n2284 vdd.n2283 185
R15061 vdd.n2282 vdd.n2150 185
R15062 vdd.n2281 vdd.n2280 185
R15063 vdd.n2535 vdd.n2534 185
R15064 vdd.n2537 vdd.n2536 185
R15065 vdd.n2539 vdd.n2538 185
R15066 vdd.n2542 vdd.n2541 185
R15067 vdd.n2544 vdd.n2543 185
R15068 vdd.n2546 vdd.n2545 185
R15069 vdd.n2548 vdd.n2547 185
R15070 vdd.n2550 vdd.n2549 185
R15071 vdd.n2552 vdd.n2551 185
R15072 vdd.n2554 vdd.n2553 185
R15073 vdd.n2556 vdd.n2555 185
R15074 vdd.n2558 vdd.n2557 185
R15075 vdd.n2560 vdd.n2559 185
R15076 vdd.n2562 vdd.n2561 185
R15077 vdd.n2564 vdd.n2563 185
R15078 vdd.n2566 vdd.n2565 185
R15079 vdd.n2568 vdd.n2567 185
R15080 vdd.n2570 vdd.n2569 185
R15081 vdd.n2572 vdd.n2571 185
R15082 vdd.n2574 vdd.n2573 185
R15083 vdd.n2576 vdd.n2575 185
R15084 vdd.n2578 vdd.n2577 185
R15085 vdd.n2580 vdd.n2579 185
R15086 vdd.n2582 vdd.n2581 185
R15087 vdd.n2584 vdd.n2583 185
R15088 vdd.n2586 vdd.n2585 185
R15089 vdd.n2588 vdd.n2587 185
R15090 vdd.n2590 vdd.n2589 185
R15091 vdd.n2592 vdd.n2591 185
R15092 vdd.n2594 vdd.n2593 185
R15093 vdd.n2596 vdd.n2595 185
R15094 vdd.n2598 vdd.n2597 185
R15095 vdd.n2600 vdd.n2599 185
R15096 vdd.n2601 vdd.n955 185
R15097 vdd.n2603 vdd.n2602 185
R15098 vdd.n2604 vdd.n2603 185
R15099 vdd.n2533 vdd.n959 185
R15100 vdd.n2533 vdd.n2532 185
R15101 vdd.n2154 vdd.n960 185
R15102 vdd.t35 vdd.n960 185
R15103 vdd.n2155 vdd.n970 185
R15104 vdd.n2457 vdd.n970 185
R15105 vdd.n2158 vdd.n2157 185
R15106 vdd.n2157 vdd.n2156 185
R15107 vdd.n2159 vdd.n977 185
R15108 vdd.n2450 vdd.n977 185
R15109 vdd.n2161 vdd.n2160 185
R15110 vdd.n2160 vdd.n976 185
R15111 vdd.n2162 vdd.n984 185
R15112 vdd.n2442 vdd.n984 185
R15113 vdd.n2164 vdd.n2163 185
R15114 vdd.n2163 vdd.n983 185
R15115 vdd.n2165 vdd.n990 185
R15116 vdd.n2436 vdd.n990 185
R15117 vdd.n2167 vdd.n2166 185
R15118 vdd.n2166 vdd.n989 185
R15119 vdd.n2168 vdd.n995 185
R15120 vdd.n2430 vdd.n995 185
R15121 vdd.n2170 vdd.n2169 185
R15122 vdd.n2169 vdd.n1002 185
R15123 vdd.n2171 vdd.n1000 185
R15124 vdd.n2424 vdd.n1000 185
R15125 vdd.n2173 vdd.n2172 185
R15126 vdd.n2172 vdd.n1008 185
R15127 vdd.n2174 vdd.n1006 185
R15128 vdd.n2418 vdd.n1006 185
R15129 vdd.n2259 vdd.n2258 185
R15130 vdd.n2258 vdd.n2257 185
R15131 vdd.n2260 vdd.n1013 185
R15132 vdd.n2412 vdd.n1013 185
R15133 vdd.n2262 vdd.n2261 185
R15134 vdd.n2261 vdd.n1012 185
R15135 vdd.n2263 vdd.n1019 185
R15136 vdd.n2406 vdd.n1019 185
R15137 vdd.n2265 vdd.n2264 185
R15138 vdd.n2264 vdd.n1018 185
R15139 vdd.n2266 vdd.n1024 185
R15140 vdd.n2400 vdd.n1024 185
R15141 vdd.n2268 vdd.n2267 185
R15142 vdd.n2267 vdd.n1033 185
R15143 vdd.n2269 vdd.n1031 185
R15144 vdd.n2393 vdd.n1031 185
R15145 vdd.n2271 vdd.n2270 185
R15146 vdd.n2270 vdd.n1030 185
R15147 vdd.n2272 vdd.n1038 185
R15148 vdd.n2387 vdd.n1038 185
R15149 vdd.n2274 vdd.n2273 185
R15150 vdd.n2273 vdd.n1037 185
R15151 vdd.n2275 vdd.n1044 185
R15152 vdd.n2381 vdd.n1044 185
R15153 vdd.n2277 vdd.n2276 185
R15154 vdd.n2276 vdd.n1043 185
R15155 vdd.n2278 vdd.n1050 185
R15156 vdd.n2375 vdd.n1050 185
R15157 vdd.n3357 vdd.n3356 185
R15158 vdd.n3356 vdd.n3355 185
R15159 vdd.n3358 vdd.n387 185
R15160 vdd.n387 vdd.n386 185
R15161 vdd.n3360 vdd.n3359 185
R15162 vdd.n3361 vdd.n3360 185
R15163 vdd.n382 vdd.n381 185
R15164 vdd.n3362 vdd.n382 185
R15165 vdd.n3365 vdd.n3364 185
R15166 vdd.n3364 vdd.n3363 185
R15167 vdd.n3366 vdd.n376 185
R15168 vdd.n376 vdd.n375 185
R15169 vdd.n3368 vdd.n3367 185
R15170 vdd.n3369 vdd.n3368 185
R15171 vdd.n371 vdd.n370 185
R15172 vdd.n3370 vdd.n371 185
R15173 vdd.n3373 vdd.n3372 185
R15174 vdd.n3372 vdd.n3371 185
R15175 vdd.n3374 vdd.n365 185
R15176 vdd.n3331 vdd.n365 185
R15177 vdd.n3376 vdd.n3375 185
R15178 vdd.n3377 vdd.n3376 185
R15179 vdd.n360 vdd.n359 185
R15180 vdd.n3378 vdd.n360 185
R15181 vdd.n3381 vdd.n3380 185
R15182 vdd.n3380 vdd.n3379 185
R15183 vdd.n3382 vdd.n354 185
R15184 vdd.n361 vdd.n354 185
R15185 vdd.n3384 vdd.n3383 185
R15186 vdd.n3385 vdd.n3384 185
R15187 vdd.n350 vdd.n349 185
R15188 vdd.n3386 vdd.n350 185
R15189 vdd.n3389 vdd.n3388 185
R15190 vdd.n3388 vdd.n3387 185
R15191 vdd.n3390 vdd.n345 185
R15192 vdd.n345 vdd.n344 185
R15193 vdd.n3392 vdd.n3391 185
R15194 vdd.n3393 vdd.n3392 185
R15195 vdd.n339 vdd.n337 185
R15196 vdd.n3394 vdd.n339 185
R15197 vdd.n3397 vdd.n3396 185
R15198 vdd.n3396 vdd.n3395 185
R15199 vdd.n338 vdd.n336 185
R15200 vdd.n340 vdd.n338 185
R15201 vdd.n3307 vdd.n3306 185
R15202 vdd.n3308 vdd.n3307 185
R15203 vdd.n635 vdd.n634 185
R15204 vdd.n634 vdd.n633 185
R15205 vdd.n3302 vdd.n3301 185
R15206 vdd.n3301 vdd.n3300 185
R15207 vdd.n638 vdd.n637 185
R15208 vdd.n644 vdd.n638 185
R15209 vdd.n3288 vdd.n3287 185
R15210 vdd.n3289 vdd.n3288 185
R15211 vdd.n646 vdd.n645 185
R15212 vdd.n3280 vdd.n645 185
R15213 vdd.n3283 vdd.n3282 185
R15214 vdd.n3282 vdd.n3281 185
R15215 vdd.n649 vdd.n648 185
R15216 vdd.n656 vdd.n649 185
R15217 vdd.n3271 vdd.n3270 185
R15218 vdd.n3272 vdd.n3271 185
R15219 vdd.n658 vdd.n657 185
R15220 vdd.n657 vdd.n655 185
R15221 vdd.n3266 vdd.n3265 185
R15222 vdd.n3265 vdd.n3264 185
R15223 vdd.n661 vdd.n660 185
R15224 vdd.n662 vdd.n661 185
R15225 vdd.n3255 vdd.n3254 185
R15226 vdd.n3256 vdd.n3255 185
R15227 vdd.n669 vdd.n668 185
R15228 vdd.n3247 vdd.n668 185
R15229 vdd.n3250 vdd.n3249 185
R15230 vdd.n3249 vdd.n3248 185
R15231 vdd.n672 vdd.n671 185
R15232 vdd.n679 vdd.n672 185
R15233 vdd.n3238 vdd.n3237 185
R15234 vdd.n3239 vdd.n3238 185
R15235 vdd.n681 vdd.n680 185
R15236 vdd.n680 vdd.n678 185
R15237 vdd.n3233 vdd.n3232 185
R15238 vdd.n3232 vdd.n3231 185
R15239 vdd.n684 vdd.n683 185
R15240 vdd.n723 vdd.n684 185
R15241 vdd.n3221 vdd.n3220 185
R15242 vdd.n3219 vdd.n725 185
R15243 vdd.n3218 vdd.n724 185
R15244 vdd.n3223 vdd.n724 185
R15245 vdd.n729 vdd.n728 185
R15246 vdd.n733 vdd.n732 185
R15247 vdd.n3214 vdd.n734 185
R15248 vdd.n3213 vdd.n3212 185
R15249 vdd.n3211 vdd.n3210 185
R15250 vdd.n3209 vdd.n3208 185
R15251 vdd.n3207 vdd.n3206 185
R15252 vdd.n3205 vdd.n3204 185
R15253 vdd.n3203 vdd.n3202 185
R15254 vdd.n3201 vdd.n3200 185
R15255 vdd.n3199 vdd.n3198 185
R15256 vdd.n3197 vdd.n3196 185
R15257 vdd.n3195 vdd.n3194 185
R15258 vdd.n3193 vdd.n3192 185
R15259 vdd.n3191 vdd.n3190 185
R15260 vdd.n3189 vdd.n3188 185
R15261 vdd.n3187 vdd.n3186 185
R15262 vdd.n3178 vdd.n747 185
R15263 vdd.n3180 vdd.n3179 185
R15264 vdd.n3177 vdd.n3176 185
R15265 vdd.n3175 vdd.n3174 185
R15266 vdd.n3173 vdd.n3172 185
R15267 vdd.n3171 vdd.n3170 185
R15268 vdd.n3169 vdd.n3168 185
R15269 vdd.n3167 vdd.n3166 185
R15270 vdd.n3165 vdd.n3164 185
R15271 vdd.n3163 vdd.n3162 185
R15272 vdd.n3161 vdd.n3160 185
R15273 vdd.n3159 vdd.n3158 185
R15274 vdd.n3157 vdd.n3156 185
R15275 vdd.n3155 vdd.n3154 185
R15276 vdd.n3153 vdd.n3152 185
R15277 vdd.n3151 vdd.n3150 185
R15278 vdd.n3149 vdd.n3148 185
R15279 vdd.n3147 vdd.n3146 185
R15280 vdd.n3145 vdd.n3144 185
R15281 vdd.n3143 vdd.n3142 185
R15282 vdd.n3141 vdd.n3140 185
R15283 vdd.n3139 vdd.n3138 185
R15284 vdd.n3132 vdd.n767 185
R15285 vdd.n3134 vdd.n3133 185
R15286 vdd.n3131 vdd.n3130 185
R15287 vdd.n3129 vdd.n3128 185
R15288 vdd.n3127 vdd.n3126 185
R15289 vdd.n3125 vdd.n3124 185
R15290 vdd.n3123 vdd.n3122 185
R15291 vdd.n3121 vdd.n3120 185
R15292 vdd.n3119 vdd.n3118 185
R15293 vdd.n3117 vdd.n3116 185
R15294 vdd.n3115 vdd.n3114 185
R15295 vdd.n3113 vdd.n3112 185
R15296 vdd.n3111 vdd.n3110 185
R15297 vdd.n3109 vdd.n3108 185
R15298 vdd.n3107 vdd.n3106 185
R15299 vdd.n3105 vdd.n3104 185
R15300 vdd.n3103 vdd.n3102 185
R15301 vdd.n3101 vdd.n3100 185
R15302 vdd.n3099 vdd.n3098 185
R15303 vdd.n3097 vdd.n3096 185
R15304 vdd.n3095 vdd.n691 185
R15305 vdd.n3225 vdd.n3224 185
R15306 vdd.n3224 vdd.n3223 185
R15307 vdd.n3352 vdd.n3351 185
R15308 vdd.n618 vdd.n425 185
R15309 vdd.n617 vdd.n616 185
R15310 vdd.n615 vdd.n614 185
R15311 vdd.n613 vdd.n430 185
R15312 vdd.n609 vdd.n608 185
R15313 vdd.n607 vdd.n606 185
R15314 vdd.n605 vdd.n604 185
R15315 vdd.n603 vdd.n432 185
R15316 vdd.n599 vdd.n598 185
R15317 vdd.n597 vdd.n596 185
R15318 vdd.n595 vdd.n594 185
R15319 vdd.n593 vdd.n434 185
R15320 vdd.n589 vdd.n588 185
R15321 vdd.n587 vdd.n586 185
R15322 vdd.n585 vdd.n584 185
R15323 vdd.n583 vdd.n436 185
R15324 vdd.n579 vdd.n578 185
R15325 vdd.n577 vdd.n576 185
R15326 vdd.n575 vdd.n574 185
R15327 vdd.n573 vdd.n438 185
R15328 vdd.n569 vdd.n568 185
R15329 vdd.n567 vdd.n566 185
R15330 vdd.n565 vdd.n564 185
R15331 vdd.n563 vdd.n442 185
R15332 vdd.n559 vdd.n558 185
R15333 vdd.n557 vdd.n556 185
R15334 vdd.n555 vdd.n554 185
R15335 vdd.n553 vdd.n444 185
R15336 vdd.n549 vdd.n548 185
R15337 vdd.n547 vdd.n546 185
R15338 vdd.n545 vdd.n544 185
R15339 vdd.n543 vdd.n446 185
R15340 vdd.n539 vdd.n538 185
R15341 vdd.n537 vdd.n536 185
R15342 vdd.n535 vdd.n534 185
R15343 vdd.n533 vdd.n448 185
R15344 vdd.n529 vdd.n528 185
R15345 vdd.n527 vdd.n526 185
R15346 vdd.n525 vdd.n524 185
R15347 vdd.n523 vdd.n450 185
R15348 vdd.n519 vdd.n518 185
R15349 vdd.n517 vdd.n516 185
R15350 vdd.n515 vdd.n514 185
R15351 vdd.n513 vdd.n454 185
R15352 vdd.n509 vdd.n508 185
R15353 vdd.n507 vdd.n506 185
R15354 vdd.n505 vdd.n504 185
R15355 vdd.n503 vdd.n456 185
R15356 vdd.n499 vdd.n498 185
R15357 vdd.n497 vdd.n496 185
R15358 vdd.n495 vdd.n494 185
R15359 vdd.n493 vdd.n458 185
R15360 vdd.n489 vdd.n488 185
R15361 vdd.n487 vdd.n486 185
R15362 vdd.n485 vdd.n484 185
R15363 vdd.n483 vdd.n460 185
R15364 vdd.n479 vdd.n478 185
R15365 vdd.n477 vdd.n476 185
R15366 vdd.n475 vdd.n474 185
R15367 vdd.n473 vdd.n462 185
R15368 vdd.n469 vdd.n468 185
R15369 vdd.n467 vdd.n466 185
R15370 vdd.n465 vdd.n392 185
R15371 vdd.n3348 vdd.n393 185
R15372 vdd.n3355 vdd.n393 185
R15373 vdd.n3347 vdd.n3346 185
R15374 vdd.n3346 vdd.n386 185
R15375 vdd.n3345 vdd.n385 185
R15376 vdd.n3361 vdd.n385 185
R15377 vdd.n621 vdd.n384 185
R15378 vdd.n3362 vdd.n384 185
R15379 vdd.n3341 vdd.n383 185
R15380 vdd.n3363 vdd.n383 185
R15381 vdd.n3340 vdd.n3339 185
R15382 vdd.n3339 vdd.n375 185
R15383 vdd.n3338 vdd.n374 185
R15384 vdd.n3369 vdd.n374 185
R15385 vdd.n623 vdd.n373 185
R15386 vdd.n3370 vdd.n373 185
R15387 vdd.n3334 vdd.n372 185
R15388 vdd.n3371 vdd.n372 185
R15389 vdd.n3333 vdd.n3332 185
R15390 vdd.n3332 vdd.n3331 185
R15391 vdd.n3330 vdd.n364 185
R15392 vdd.n3377 vdd.n364 185
R15393 vdd.n625 vdd.n363 185
R15394 vdd.n3378 vdd.n363 185
R15395 vdd.n3326 vdd.n362 185
R15396 vdd.n3379 vdd.n362 185
R15397 vdd.n3325 vdd.n3324 185
R15398 vdd.n3324 vdd.n361 185
R15399 vdd.n3323 vdd.n353 185
R15400 vdd.n3385 vdd.n353 185
R15401 vdd.n627 vdd.n352 185
R15402 vdd.n3386 vdd.n352 185
R15403 vdd.n3319 vdd.n351 185
R15404 vdd.n3387 vdd.n351 185
R15405 vdd.n3318 vdd.n3317 185
R15406 vdd.n3317 vdd.n344 185
R15407 vdd.n3316 vdd.n343 185
R15408 vdd.n3393 vdd.n343 185
R15409 vdd.n629 vdd.n342 185
R15410 vdd.n3394 vdd.n342 185
R15411 vdd.n3312 vdd.n341 185
R15412 vdd.n3395 vdd.n341 185
R15413 vdd.n3311 vdd.n3310 185
R15414 vdd.n3310 vdd.n340 185
R15415 vdd.n3309 vdd.n631 185
R15416 vdd.n3309 vdd.n3308 185
R15417 vdd.n3297 vdd.n632 185
R15418 vdd.n633 vdd.n632 185
R15419 vdd.n3299 vdd.n3298 185
R15420 vdd.n3300 vdd.n3299 185
R15421 vdd.n640 vdd.n639 185
R15422 vdd.n644 vdd.n639 185
R15423 vdd.n3291 vdd.n3290 185
R15424 vdd.n3290 vdd.n3289 185
R15425 vdd.n643 vdd.n642 185
R15426 vdd.n3280 vdd.n643 185
R15427 vdd.n3279 vdd.n3278 185
R15428 vdd.n3281 vdd.n3279 185
R15429 vdd.n651 vdd.n650 185
R15430 vdd.n656 vdd.n650 185
R15431 vdd.n3274 vdd.n3273 185
R15432 vdd.n3273 vdd.n3272 185
R15433 vdd.n654 vdd.n653 185
R15434 vdd.n655 vdd.n654 185
R15435 vdd.n3263 vdd.n3262 185
R15436 vdd.n3264 vdd.n3263 185
R15437 vdd.n664 vdd.n663 185
R15438 vdd.n663 vdd.n662 185
R15439 vdd.n3258 vdd.n3257 185
R15440 vdd.n3257 vdd.n3256 185
R15441 vdd.n667 vdd.n666 185
R15442 vdd.n3247 vdd.n667 185
R15443 vdd.n3246 vdd.n3245 185
R15444 vdd.n3248 vdd.n3246 185
R15445 vdd.n674 vdd.n673 185
R15446 vdd.n679 vdd.n673 185
R15447 vdd.n3241 vdd.n3240 185
R15448 vdd.n3240 vdd.n3239 185
R15449 vdd.n677 vdd.n676 185
R15450 vdd.n678 vdd.n677 185
R15451 vdd.n3230 vdd.n3229 185
R15452 vdd.n3231 vdd.n3230 185
R15453 vdd.n686 vdd.n685 185
R15454 vdd.n723 vdd.n685 185
R15455 vdd.n913 vdd.n912 185
R15456 vdd.n2855 vdd.n2854 185
R15457 vdd.n2853 vdd.n2638 185
R15458 vdd.n2857 vdd.n2638 185
R15459 vdd.n2852 vdd.n2851 185
R15460 vdd.n2850 vdd.n2849 185
R15461 vdd.n2848 vdd.n2847 185
R15462 vdd.n2846 vdd.n2845 185
R15463 vdd.n2844 vdd.n2843 185
R15464 vdd.n2842 vdd.n2841 185
R15465 vdd.n2840 vdd.n2839 185
R15466 vdd.n2838 vdd.n2837 185
R15467 vdd.n2836 vdd.n2835 185
R15468 vdd.n2834 vdd.n2833 185
R15469 vdd.n2832 vdd.n2831 185
R15470 vdd.n2830 vdd.n2829 185
R15471 vdd.n2828 vdd.n2827 185
R15472 vdd.n2826 vdd.n2825 185
R15473 vdd.n2824 vdd.n2823 185
R15474 vdd.n2822 vdd.n2821 185
R15475 vdd.n2820 vdd.n2819 185
R15476 vdd.n2818 vdd.n2817 185
R15477 vdd.n2816 vdd.n2815 185
R15478 vdd.n2814 vdd.n2813 185
R15479 vdd.n2812 vdd.n2811 185
R15480 vdd.n2810 vdd.n2809 185
R15481 vdd.n2808 vdd.n2807 185
R15482 vdd.n2806 vdd.n2805 185
R15483 vdd.n2804 vdd.n2803 185
R15484 vdd.n2802 vdd.n2801 185
R15485 vdd.n2800 vdd.n2799 185
R15486 vdd.n2798 vdd.n2797 185
R15487 vdd.n2796 vdd.n2795 185
R15488 vdd.n2793 vdd.n2792 185
R15489 vdd.n2791 vdd.n2790 185
R15490 vdd.n2789 vdd.n2788 185
R15491 vdd.n2995 vdd.n2994 185
R15492 vdd.n2997 vdd.n834 185
R15493 vdd.n2999 vdd.n2998 185
R15494 vdd.n3001 vdd.n831 185
R15495 vdd.n3003 vdd.n3002 185
R15496 vdd.n3005 vdd.n829 185
R15497 vdd.n3007 vdd.n3006 185
R15498 vdd.n3008 vdd.n828 185
R15499 vdd.n3010 vdd.n3009 185
R15500 vdd.n3012 vdd.n826 185
R15501 vdd.n3014 vdd.n3013 185
R15502 vdd.n3015 vdd.n825 185
R15503 vdd.n3017 vdd.n3016 185
R15504 vdd.n3019 vdd.n823 185
R15505 vdd.n3021 vdd.n3020 185
R15506 vdd.n3022 vdd.n822 185
R15507 vdd.n3024 vdd.n3023 185
R15508 vdd.n3026 vdd.n731 185
R15509 vdd.n3028 vdd.n3027 185
R15510 vdd.n3030 vdd.n820 185
R15511 vdd.n3032 vdd.n3031 185
R15512 vdd.n3033 vdd.n819 185
R15513 vdd.n3035 vdd.n3034 185
R15514 vdd.n3037 vdd.n817 185
R15515 vdd.n3039 vdd.n3038 185
R15516 vdd.n3040 vdd.n816 185
R15517 vdd.n3042 vdd.n3041 185
R15518 vdd.n3044 vdd.n814 185
R15519 vdd.n3046 vdd.n3045 185
R15520 vdd.n3047 vdd.n813 185
R15521 vdd.n3049 vdd.n3048 185
R15522 vdd.n3051 vdd.n812 185
R15523 vdd.n3052 vdd.n811 185
R15524 vdd.n3055 vdd.n3054 185
R15525 vdd.n3056 vdd.n809 185
R15526 vdd.n809 vdd.n692 185
R15527 vdd.n2993 vdd.n806 185
R15528 vdd.n3059 vdd.n806 185
R15529 vdd.n2992 vdd.n2991 185
R15530 vdd.n2991 vdd.n805 185
R15531 vdd.n2990 vdd.n836 185
R15532 vdd.n2990 vdd.n2989 185
R15533 vdd.n2744 vdd.n837 185
R15534 vdd.n846 vdd.n837 185
R15535 vdd.n2745 vdd.n844 185
R15536 vdd.n2983 vdd.n844 185
R15537 vdd.n2747 vdd.n2746 185
R15538 vdd.n2746 vdd.n843 185
R15539 vdd.n2748 vdd.n852 185
R15540 vdd.n2932 vdd.n852 185
R15541 vdd.n2750 vdd.n2749 185
R15542 vdd.n2749 vdd.n851 185
R15543 vdd.n2751 vdd.n858 185
R15544 vdd.n2926 vdd.n858 185
R15545 vdd.n2753 vdd.n2752 185
R15546 vdd.n2752 vdd.n857 185
R15547 vdd.n2754 vdd.n863 185
R15548 vdd.n2918 vdd.n863 185
R15549 vdd.n2756 vdd.n2755 185
R15550 vdd.n2755 vdd.n870 185
R15551 vdd.n2757 vdd.n868 185
R15552 vdd.n2912 vdd.n868 185
R15553 vdd.n2759 vdd.n2758 185
R15554 vdd.n2760 vdd.n2759 185
R15555 vdd.n2743 vdd.n875 185
R15556 vdd.n2906 vdd.n875 185
R15557 vdd.n2742 vdd.n2741 185
R15558 vdd.n2741 vdd.n874 185
R15559 vdd.n2740 vdd.n881 185
R15560 vdd.n2900 vdd.n881 185
R15561 vdd.n2739 vdd.n2738 185
R15562 vdd.n2738 vdd.n880 185
R15563 vdd.n2737 vdd.n886 185
R15564 vdd.n2894 vdd.n886 185
R15565 vdd.n2736 vdd.n2735 185
R15566 vdd.n2735 vdd.n893 185
R15567 vdd.n2734 vdd.n891 185
R15568 vdd.n2888 vdd.n891 185
R15569 vdd.n2733 vdd.n2732 185
R15570 vdd.n2732 vdd.n900 185
R15571 vdd.n2731 vdd.n898 185
R15572 vdd.n2882 vdd.n898 185
R15573 vdd.n2730 vdd.n2729 185
R15574 vdd.n2729 vdd.n897 185
R15575 vdd.n2641 vdd.n904 185
R15576 vdd.n2876 vdd.n904 185
R15577 vdd.n2783 vdd.n2782 185
R15578 vdd.n2782 vdd.n2781 185
R15579 vdd.n2784 vdd.n909 185
R15580 vdd.n2870 vdd.n909 185
R15581 vdd.n2786 vdd.n2785 185
R15582 vdd.n2785 vdd.t132 185
R15583 vdd.n2787 vdd.n914 185
R15584 vdd.n2864 vdd.n914 185
R15585 vdd.n2866 vdd.n2865 185
R15586 vdd.n2865 vdd.n2864 185
R15587 vdd.n2867 vdd.n911 185
R15588 vdd.n911 vdd.t132 185
R15589 vdd.n2869 vdd.n2868 185
R15590 vdd.n2870 vdd.n2869 185
R15591 vdd.n903 vdd.n902 185
R15592 vdd.n2781 vdd.n903 185
R15593 vdd.n2878 vdd.n2877 185
R15594 vdd.n2877 vdd.n2876 185
R15595 vdd.n2879 vdd.n901 185
R15596 vdd.n901 vdd.n897 185
R15597 vdd.n2881 vdd.n2880 185
R15598 vdd.n2882 vdd.n2881 185
R15599 vdd.n890 vdd.n889 185
R15600 vdd.n900 vdd.n890 185
R15601 vdd.n2890 vdd.n2889 185
R15602 vdd.n2889 vdd.n2888 185
R15603 vdd.n2891 vdd.n888 185
R15604 vdd.n893 vdd.n888 185
R15605 vdd.n2893 vdd.n2892 185
R15606 vdd.n2894 vdd.n2893 185
R15607 vdd.n879 vdd.n878 185
R15608 vdd.n880 vdd.n879 185
R15609 vdd.n2902 vdd.n2901 185
R15610 vdd.n2901 vdd.n2900 185
R15611 vdd.n2903 vdd.n877 185
R15612 vdd.n877 vdd.n874 185
R15613 vdd.n2905 vdd.n2904 185
R15614 vdd.n2906 vdd.n2905 185
R15615 vdd.n867 vdd.n866 185
R15616 vdd.n2760 vdd.n867 185
R15617 vdd.n2914 vdd.n2913 185
R15618 vdd.n2913 vdd.n2912 185
R15619 vdd.n2915 vdd.n865 185
R15620 vdd.n870 vdd.n865 185
R15621 vdd.n2917 vdd.n2916 185
R15622 vdd.n2918 vdd.n2917 185
R15623 vdd.n856 vdd.n855 185
R15624 vdd.n857 vdd.n856 185
R15625 vdd.n2928 vdd.n2927 185
R15626 vdd.n2927 vdd.n2926 185
R15627 vdd.n2929 vdd.n854 185
R15628 vdd.n854 vdd.n851 185
R15629 vdd.n2931 vdd.n2930 185
R15630 vdd.n2932 vdd.n2931 185
R15631 vdd.n842 vdd.n841 185
R15632 vdd.n843 vdd.n842 185
R15633 vdd.n2985 vdd.n2984 185
R15634 vdd.n2984 vdd.n2983 185
R15635 vdd.n2986 vdd.n840 185
R15636 vdd.n846 vdd.n840 185
R15637 vdd.n2988 vdd.n2987 185
R15638 vdd.n2989 vdd.n2988 185
R15639 vdd.n810 vdd.n808 185
R15640 vdd.n808 vdd.n805 185
R15641 vdd.n3058 vdd.n3057 185
R15642 vdd.n3059 vdd.n3058 185
R15643 vdd.n2531 vdd.n2530 185
R15644 vdd.n2532 vdd.n2531 185
R15645 vdd.n964 vdd.n962 185
R15646 vdd.n962 vdd.t35 185
R15647 vdd.n2446 vdd.n971 185
R15648 vdd.n2457 vdd.n971 185
R15649 vdd.n2447 vdd.n980 185
R15650 vdd.n2156 vdd.n980 185
R15651 vdd.n2449 vdd.n2448 185
R15652 vdd.n2450 vdd.n2449 185
R15653 vdd.n2445 vdd.n979 185
R15654 vdd.n979 vdd.n976 185
R15655 vdd.n2444 vdd.n2443 185
R15656 vdd.n2443 vdd.n2442 185
R15657 vdd.n982 vdd.n981 185
R15658 vdd.n983 vdd.n982 185
R15659 vdd.n2435 vdd.n2434 185
R15660 vdd.n2436 vdd.n2435 185
R15661 vdd.n2433 vdd.n992 185
R15662 vdd.n992 vdd.n989 185
R15663 vdd.n2432 vdd.n2431 185
R15664 vdd.n2431 vdd.n2430 185
R15665 vdd.n994 vdd.n993 185
R15666 vdd.n1002 vdd.n994 185
R15667 vdd.n2423 vdd.n2422 185
R15668 vdd.n2424 vdd.n2423 185
R15669 vdd.n2421 vdd.n1003 185
R15670 vdd.n1008 vdd.n1003 185
R15671 vdd.n2420 vdd.n2419 185
R15672 vdd.n2419 vdd.n2418 185
R15673 vdd.n1005 vdd.n1004 185
R15674 vdd.n2257 vdd.n1005 185
R15675 vdd.n2411 vdd.n2410 185
R15676 vdd.n2412 vdd.n2411 185
R15677 vdd.n2409 vdd.n1015 185
R15678 vdd.n1015 vdd.n1012 185
R15679 vdd.n2408 vdd.n2407 185
R15680 vdd.n2407 vdd.n2406 185
R15681 vdd.n1017 vdd.n1016 185
R15682 vdd.n1018 vdd.n1017 185
R15683 vdd.n2399 vdd.n2398 185
R15684 vdd.n2400 vdd.n2399 185
R15685 vdd.n2396 vdd.n1026 185
R15686 vdd.n1033 vdd.n1026 185
R15687 vdd.n2395 vdd.n2394 185
R15688 vdd.n2394 vdd.n2393 185
R15689 vdd.n1029 vdd.n1028 185
R15690 vdd.n1030 vdd.n1029 185
R15691 vdd.n2386 vdd.n2385 185
R15692 vdd.n2387 vdd.n2386 185
R15693 vdd.n2384 vdd.n1040 185
R15694 vdd.n1040 vdd.n1037 185
R15695 vdd.n2383 vdd.n2382 185
R15696 vdd.n2382 vdd.n2381 185
R15697 vdd.n1042 vdd.n1041 185
R15698 vdd.n1043 vdd.n1042 185
R15699 vdd.n2374 vdd.n2373 185
R15700 vdd.n2375 vdd.n2374 185
R15701 vdd.n2462 vdd.n936 185
R15702 vdd.n2604 vdd.n936 185
R15703 vdd.n2464 vdd.n2463 185
R15704 vdd.n2466 vdd.n2465 185
R15705 vdd.n2468 vdd.n2467 185
R15706 vdd.n2470 vdd.n2469 185
R15707 vdd.n2472 vdd.n2471 185
R15708 vdd.n2474 vdd.n2473 185
R15709 vdd.n2476 vdd.n2475 185
R15710 vdd.n2478 vdd.n2477 185
R15711 vdd.n2480 vdd.n2479 185
R15712 vdd.n2482 vdd.n2481 185
R15713 vdd.n2484 vdd.n2483 185
R15714 vdd.n2486 vdd.n2485 185
R15715 vdd.n2488 vdd.n2487 185
R15716 vdd.n2490 vdd.n2489 185
R15717 vdd.n2492 vdd.n2491 185
R15718 vdd.n2494 vdd.n2493 185
R15719 vdd.n2496 vdd.n2495 185
R15720 vdd.n2498 vdd.n2497 185
R15721 vdd.n2500 vdd.n2499 185
R15722 vdd.n2502 vdd.n2501 185
R15723 vdd.n2504 vdd.n2503 185
R15724 vdd.n2506 vdd.n2505 185
R15725 vdd.n2508 vdd.n2507 185
R15726 vdd.n2510 vdd.n2509 185
R15727 vdd.n2512 vdd.n2511 185
R15728 vdd.n2514 vdd.n2513 185
R15729 vdd.n2516 vdd.n2515 185
R15730 vdd.n2518 vdd.n2517 185
R15731 vdd.n2520 vdd.n2519 185
R15732 vdd.n2522 vdd.n2521 185
R15733 vdd.n2524 vdd.n2523 185
R15734 vdd.n2526 vdd.n2525 185
R15735 vdd.n2528 vdd.n2527 185
R15736 vdd.n2529 vdd.n963 185
R15737 vdd.n2461 vdd.n961 185
R15738 vdd.n2532 vdd.n961 185
R15739 vdd.n2460 vdd.n2459 185
R15740 vdd.n2459 vdd.t35 185
R15741 vdd.n2458 vdd.n968 185
R15742 vdd.n2458 vdd.n2457 185
R15743 vdd.n2238 vdd.n969 185
R15744 vdd.n2156 vdd.n969 185
R15745 vdd.n2239 vdd.n978 185
R15746 vdd.n2450 vdd.n978 185
R15747 vdd.n2241 vdd.n2240 185
R15748 vdd.n2240 vdd.n976 185
R15749 vdd.n2242 vdd.n985 185
R15750 vdd.n2442 vdd.n985 185
R15751 vdd.n2244 vdd.n2243 185
R15752 vdd.n2243 vdd.n983 185
R15753 vdd.n2245 vdd.n991 185
R15754 vdd.n2436 vdd.n991 185
R15755 vdd.n2247 vdd.n2246 185
R15756 vdd.n2246 vdd.n989 185
R15757 vdd.n2248 vdd.n996 185
R15758 vdd.n2430 vdd.n996 185
R15759 vdd.n2250 vdd.n2249 185
R15760 vdd.n2249 vdd.n1002 185
R15761 vdd.n2251 vdd.n1001 185
R15762 vdd.n2424 vdd.n1001 185
R15763 vdd.n2253 vdd.n2252 185
R15764 vdd.n2252 vdd.n1008 185
R15765 vdd.n2254 vdd.n1007 185
R15766 vdd.n2418 vdd.n1007 185
R15767 vdd.n2256 vdd.n2255 185
R15768 vdd.n2257 vdd.n2256 185
R15769 vdd.n2237 vdd.n1014 185
R15770 vdd.n2412 vdd.n1014 185
R15771 vdd.n2236 vdd.n2235 185
R15772 vdd.n2235 vdd.n1012 185
R15773 vdd.n2234 vdd.n1020 185
R15774 vdd.n2406 vdd.n1020 185
R15775 vdd.n2233 vdd.n2232 185
R15776 vdd.n2232 vdd.n1018 185
R15777 vdd.n2231 vdd.n1025 185
R15778 vdd.n2400 vdd.n1025 185
R15779 vdd.n2230 vdd.n2229 185
R15780 vdd.n2229 vdd.n1033 185
R15781 vdd.n2228 vdd.n1032 185
R15782 vdd.n2393 vdd.n1032 185
R15783 vdd.n2227 vdd.n2226 185
R15784 vdd.n2226 vdd.n1030 185
R15785 vdd.n2225 vdd.n1039 185
R15786 vdd.n2387 vdd.n1039 185
R15787 vdd.n2224 vdd.n2223 185
R15788 vdd.n2223 vdd.n1037 185
R15789 vdd.n2222 vdd.n1045 185
R15790 vdd.n2381 vdd.n1045 185
R15791 vdd.n2221 vdd.n2220 185
R15792 vdd.n2220 vdd.n1043 185
R15793 vdd.n2219 vdd.n1051 185
R15794 vdd.n2375 vdd.n1051 185
R15795 vdd.n2372 vdd.n1052 185
R15796 vdd.n2371 vdd.n2370 185
R15797 vdd.n2368 vdd.n1053 185
R15798 vdd.n2366 vdd.n2365 185
R15799 vdd.n2364 vdd.n1054 185
R15800 vdd.n2363 vdd.n2362 185
R15801 vdd.n2360 vdd.n1055 185
R15802 vdd.n2358 vdd.n2357 185
R15803 vdd.n2356 vdd.n1056 185
R15804 vdd.n2355 vdd.n2354 185
R15805 vdd.n2352 vdd.n1057 185
R15806 vdd.n2350 vdd.n2349 185
R15807 vdd.n2348 vdd.n1058 185
R15808 vdd.n2347 vdd.n2346 185
R15809 vdd.n2344 vdd.n1059 185
R15810 vdd.n2342 vdd.n2341 185
R15811 vdd.n2340 vdd.n1060 185
R15812 vdd.n2339 vdd.n1062 185
R15813 vdd.n2184 vdd.n1063 185
R15814 vdd.n2187 vdd.n2186 185
R15815 vdd.n2189 vdd.n2188 185
R15816 vdd.n2191 vdd.n2183 185
R15817 vdd.n2194 vdd.n2193 185
R15818 vdd.n2195 vdd.n2182 185
R15819 vdd.n2197 vdd.n2196 185
R15820 vdd.n2199 vdd.n2181 185
R15821 vdd.n2202 vdd.n2201 185
R15822 vdd.n2203 vdd.n2180 185
R15823 vdd.n2205 vdd.n2204 185
R15824 vdd.n2207 vdd.n2179 185
R15825 vdd.n2210 vdd.n2209 185
R15826 vdd.n2211 vdd.n2176 185
R15827 vdd.n2214 vdd.n2213 185
R15828 vdd.n2216 vdd.n2175 185
R15829 vdd.n2218 vdd.n2217 185
R15830 vdd.n2217 vdd.n1049 185
R15831 vdd.n327 vdd.n326 171.744
R15832 vdd.n326 vdd.n325 171.744
R15833 vdd.n325 vdd.n294 171.744
R15834 vdd.n318 vdd.n294 171.744
R15835 vdd.n318 vdd.n317 171.744
R15836 vdd.n317 vdd.n299 171.744
R15837 vdd.n310 vdd.n299 171.744
R15838 vdd.n310 vdd.n309 171.744
R15839 vdd.n309 vdd.n303 171.744
R15840 vdd.n268 vdd.n267 171.744
R15841 vdd.n267 vdd.n266 171.744
R15842 vdd.n266 vdd.n235 171.744
R15843 vdd.n259 vdd.n235 171.744
R15844 vdd.n259 vdd.n258 171.744
R15845 vdd.n258 vdd.n240 171.744
R15846 vdd.n251 vdd.n240 171.744
R15847 vdd.n251 vdd.n250 171.744
R15848 vdd.n250 vdd.n244 171.744
R15849 vdd.n225 vdd.n224 171.744
R15850 vdd.n224 vdd.n223 171.744
R15851 vdd.n223 vdd.n192 171.744
R15852 vdd.n216 vdd.n192 171.744
R15853 vdd.n216 vdd.n215 171.744
R15854 vdd.n215 vdd.n197 171.744
R15855 vdd.n208 vdd.n197 171.744
R15856 vdd.n208 vdd.n207 171.744
R15857 vdd.n207 vdd.n201 171.744
R15858 vdd.n166 vdd.n165 171.744
R15859 vdd.n165 vdd.n164 171.744
R15860 vdd.n164 vdd.n133 171.744
R15861 vdd.n157 vdd.n133 171.744
R15862 vdd.n157 vdd.n156 171.744
R15863 vdd.n156 vdd.n138 171.744
R15864 vdd.n149 vdd.n138 171.744
R15865 vdd.n149 vdd.n148 171.744
R15866 vdd.n148 vdd.n142 171.744
R15867 vdd.n124 vdd.n123 171.744
R15868 vdd.n123 vdd.n122 171.744
R15869 vdd.n122 vdd.n91 171.744
R15870 vdd.n115 vdd.n91 171.744
R15871 vdd.n115 vdd.n114 171.744
R15872 vdd.n114 vdd.n96 171.744
R15873 vdd.n107 vdd.n96 171.744
R15874 vdd.n107 vdd.n106 171.744
R15875 vdd.n106 vdd.n100 171.744
R15876 vdd.n65 vdd.n64 171.744
R15877 vdd.n64 vdd.n63 171.744
R15878 vdd.n63 vdd.n32 171.744
R15879 vdd.n56 vdd.n32 171.744
R15880 vdd.n56 vdd.n55 171.744
R15881 vdd.n55 vdd.n37 171.744
R15882 vdd.n48 vdd.n37 171.744
R15883 vdd.n48 vdd.n47 171.744
R15884 vdd.n47 vdd.n41 171.744
R15885 vdd.n1746 vdd.n1745 171.744
R15886 vdd.n1745 vdd.n1744 171.744
R15887 vdd.n1744 vdd.n1713 171.744
R15888 vdd.n1737 vdd.n1713 171.744
R15889 vdd.n1737 vdd.n1736 171.744
R15890 vdd.n1736 vdd.n1718 171.744
R15891 vdd.n1729 vdd.n1718 171.744
R15892 vdd.n1729 vdd.n1728 171.744
R15893 vdd.n1728 vdd.n1722 171.744
R15894 vdd.n1805 vdd.n1804 171.744
R15895 vdd.n1804 vdd.n1803 171.744
R15896 vdd.n1803 vdd.n1772 171.744
R15897 vdd.n1796 vdd.n1772 171.744
R15898 vdd.n1796 vdd.n1795 171.744
R15899 vdd.n1795 vdd.n1777 171.744
R15900 vdd.n1788 vdd.n1777 171.744
R15901 vdd.n1788 vdd.n1787 171.744
R15902 vdd.n1787 vdd.n1781 171.744
R15903 vdd.n1644 vdd.n1643 171.744
R15904 vdd.n1643 vdd.n1642 171.744
R15905 vdd.n1642 vdd.n1611 171.744
R15906 vdd.n1635 vdd.n1611 171.744
R15907 vdd.n1635 vdd.n1634 171.744
R15908 vdd.n1634 vdd.n1616 171.744
R15909 vdd.n1627 vdd.n1616 171.744
R15910 vdd.n1627 vdd.n1626 171.744
R15911 vdd.n1626 vdd.n1620 171.744
R15912 vdd.n1703 vdd.n1702 171.744
R15913 vdd.n1702 vdd.n1701 171.744
R15914 vdd.n1701 vdd.n1670 171.744
R15915 vdd.n1694 vdd.n1670 171.744
R15916 vdd.n1694 vdd.n1693 171.744
R15917 vdd.n1693 vdd.n1675 171.744
R15918 vdd.n1686 vdd.n1675 171.744
R15919 vdd.n1686 vdd.n1685 171.744
R15920 vdd.n1685 vdd.n1679 171.744
R15921 vdd.n1543 vdd.n1542 171.744
R15922 vdd.n1542 vdd.n1541 171.744
R15923 vdd.n1541 vdd.n1510 171.744
R15924 vdd.n1534 vdd.n1510 171.744
R15925 vdd.n1534 vdd.n1533 171.744
R15926 vdd.n1533 vdd.n1515 171.744
R15927 vdd.n1526 vdd.n1515 171.744
R15928 vdd.n1526 vdd.n1525 171.744
R15929 vdd.n1525 vdd.n1519 171.744
R15930 vdd.n1602 vdd.n1601 171.744
R15931 vdd.n1601 vdd.n1600 171.744
R15932 vdd.n1600 vdd.n1569 171.744
R15933 vdd.n1593 vdd.n1569 171.744
R15934 vdd.n1593 vdd.n1592 171.744
R15935 vdd.n1592 vdd.n1574 171.744
R15936 vdd.n1585 vdd.n1574 171.744
R15937 vdd.n1585 vdd.n1584 171.744
R15938 vdd.n1584 vdd.n1578 171.744
R15939 vdd.n468 vdd.n467 146.341
R15940 vdd.n474 vdd.n473 146.341
R15941 vdd.n478 vdd.n477 146.341
R15942 vdd.n484 vdd.n483 146.341
R15943 vdd.n488 vdd.n487 146.341
R15944 vdd.n494 vdd.n493 146.341
R15945 vdd.n498 vdd.n497 146.341
R15946 vdd.n504 vdd.n503 146.341
R15947 vdd.n508 vdd.n507 146.341
R15948 vdd.n514 vdd.n513 146.341
R15949 vdd.n518 vdd.n517 146.341
R15950 vdd.n524 vdd.n523 146.341
R15951 vdd.n528 vdd.n527 146.341
R15952 vdd.n534 vdd.n533 146.341
R15953 vdd.n538 vdd.n537 146.341
R15954 vdd.n544 vdd.n543 146.341
R15955 vdd.n548 vdd.n547 146.341
R15956 vdd.n554 vdd.n553 146.341
R15957 vdd.n558 vdd.n557 146.341
R15958 vdd.n564 vdd.n563 146.341
R15959 vdd.n568 vdd.n567 146.341
R15960 vdd.n574 vdd.n573 146.341
R15961 vdd.n578 vdd.n577 146.341
R15962 vdd.n584 vdd.n583 146.341
R15963 vdd.n588 vdd.n587 146.341
R15964 vdd.n594 vdd.n593 146.341
R15965 vdd.n598 vdd.n597 146.341
R15966 vdd.n604 vdd.n603 146.341
R15967 vdd.n608 vdd.n607 146.341
R15968 vdd.n614 vdd.n613 146.341
R15969 vdd.n616 vdd.n425 146.341
R15970 vdd.n3230 vdd.n685 146.341
R15971 vdd.n3230 vdd.n677 146.341
R15972 vdd.n3240 vdd.n677 146.341
R15973 vdd.n3240 vdd.n673 146.341
R15974 vdd.n3246 vdd.n673 146.341
R15975 vdd.n3246 vdd.n667 146.341
R15976 vdd.n3257 vdd.n667 146.341
R15977 vdd.n3257 vdd.n663 146.341
R15978 vdd.n3263 vdd.n663 146.341
R15979 vdd.n3263 vdd.n654 146.341
R15980 vdd.n3273 vdd.n654 146.341
R15981 vdd.n3273 vdd.n650 146.341
R15982 vdd.n3279 vdd.n650 146.341
R15983 vdd.n3279 vdd.n643 146.341
R15984 vdd.n3290 vdd.n643 146.341
R15985 vdd.n3290 vdd.n639 146.341
R15986 vdd.n3299 vdd.n639 146.341
R15987 vdd.n3299 vdd.n632 146.341
R15988 vdd.n3309 vdd.n632 146.341
R15989 vdd.n3310 vdd.n3309 146.341
R15990 vdd.n3310 vdd.n341 146.341
R15991 vdd.n342 vdd.n341 146.341
R15992 vdd.n343 vdd.n342 146.341
R15993 vdd.n3317 vdd.n343 146.341
R15994 vdd.n3317 vdd.n351 146.341
R15995 vdd.n352 vdd.n351 146.341
R15996 vdd.n353 vdd.n352 146.341
R15997 vdd.n3324 vdd.n353 146.341
R15998 vdd.n3324 vdd.n362 146.341
R15999 vdd.n363 vdd.n362 146.341
R16000 vdd.n364 vdd.n363 146.341
R16001 vdd.n3332 vdd.n364 146.341
R16002 vdd.n3332 vdd.n372 146.341
R16003 vdd.n373 vdd.n372 146.341
R16004 vdd.n374 vdd.n373 146.341
R16005 vdd.n3339 vdd.n374 146.341
R16006 vdd.n3339 vdd.n383 146.341
R16007 vdd.n384 vdd.n383 146.341
R16008 vdd.n385 vdd.n384 146.341
R16009 vdd.n3346 vdd.n385 146.341
R16010 vdd.n3346 vdd.n393 146.341
R16011 vdd.n725 vdd.n724 146.341
R16012 vdd.n728 vdd.n724 146.341
R16013 vdd.n734 vdd.n733 146.341
R16014 vdd.n3212 vdd.n3211 146.341
R16015 vdd.n3208 vdd.n3207 146.341
R16016 vdd.n3204 vdd.n3203 146.341
R16017 vdd.n3200 vdd.n3199 146.341
R16018 vdd.n3196 vdd.n3195 146.341
R16019 vdd.n3192 vdd.n3191 146.341
R16020 vdd.n3188 vdd.n3187 146.341
R16021 vdd.n3179 vdd.n3178 146.341
R16022 vdd.n3176 vdd.n3175 146.341
R16023 vdd.n3172 vdd.n3171 146.341
R16024 vdd.n3168 vdd.n3167 146.341
R16025 vdd.n3164 vdd.n3163 146.341
R16026 vdd.n3160 vdd.n3159 146.341
R16027 vdd.n3156 vdd.n3155 146.341
R16028 vdd.n3152 vdd.n3151 146.341
R16029 vdd.n3148 vdd.n3147 146.341
R16030 vdd.n3144 vdd.n3143 146.341
R16031 vdd.n3140 vdd.n3139 146.341
R16032 vdd.n3133 vdd.n3132 146.341
R16033 vdd.n3130 vdd.n3129 146.341
R16034 vdd.n3126 vdd.n3125 146.341
R16035 vdd.n3122 vdd.n3121 146.341
R16036 vdd.n3118 vdd.n3117 146.341
R16037 vdd.n3114 vdd.n3113 146.341
R16038 vdd.n3110 vdd.n3109 146.341
R16039 vdd.n3106 vdd.n3105 146.341
R16040 vdd.n3102 vdd.n3101 146.341
R16041 vdd.n3098 vdd.n3097 146.341
R16042 vdd.n3224 vdd.n691 146.341
R16043 vdd.n3232 vdd.n684 146.341
R16044 vdd.n3232 vdd.n680 146.341
R16045 vdd.n3238 vdd.n680 146.341
R16046 vdd.n3238 vdd.n672 146.341
R16047 vdd.n3249 vdd.n672 146.341
R16048 vdd.n3249 vdd.n668 146.341
R16049 vdd.n3255 vdd.n668 146.341
R16050 vdd.n3255 vdd.n661 146.341
R16051 vdd.n3265 vdd.n661 146.341
R16052 vdd.n3265 vdd.n657 146.341
R16053 vdd.n3271 vdd.n657 146.341
R16054 vdd.n3271 vdd.n649 146.341
R16055 vdd.n3282 vdd.n649 146.341
R16056 vdd.n3282 vdd.n645 146.341
R16057 vdd.n3288 vdd.n645 146.341
R16058 vdd.n3288 vdd.n638 146.341
R16059 vdd.n3301 vdd.n638 146.341
R16060 vdd.n3301 vdd.n634 146.341
R16061 vdd.n3307 vdd.n634 146.341
R16062 vdd.n3307 vdd.n338 146.341
R16063 vdd.n3396 vdd.n338 146.341
R16064 vdd.n3396 vdd.n339 146.341
R16065 vdd.n3392 vdd.n339 146.341
R16066 vdd.n3392 vdd.n345 146.341
R16067 vdd.n3388 vdd.n345 146.341
R16068 vdd.n3388 vdd.n350 146.341
R16069 vdd.n3384 vdd.n350 146.341
R16070 vdd.n3384 vdd.n354 146.341
R16071 vdd.n3380 vdd.n354 146.341
R16072 vdd.n3380 vdd.n360 146.341
R16073 vdd.n3376 vdd.n360 146.341
R16074 vdd.n3376 vdd.n365 146.341
R16075 vdd.n3372 vdd.n365 146.341
R16076 vdd.n3372 vdd.n371 146.341
R16077 vdd.n3368 vdd.n371 146.341
R16078 vdd.n3368 vdd.n376 146.341
R16079 vdd.n3364 vdd.n376 146.341
R16080 vdd.n3364 vdd.n382 146.341
R16081 vdd.n3360 vdd.n382 146.341
R16082 vdd.n3360 vdd.n387 146.341
R16083 vdd.n3356 vdd.n387 146.341
R16084 vdd.n2322 vdd.n2321 146.341
R16085 vdd.n2319 vdd.n1903 146.341
R16086 vdd.n2099 vdd.n1909 146.341
R16087 vdd.n2097 vdd.n2096 146.341
R16088 vdd.n2094 vdd.n1911 146.341
R16089 vdd.n2090 vdd.n2089 146.341
R16090 vdd.n2087 vdd.n1918 146.341
R16091 vdd.n2083 vdd.n2082 146.341
R16092 vdd.n2080 vdd.n1925 146.341
R16093 vdd.n1936 vdd.n1933 146.341
R16094 vdd.n2072 vdd.n2071 146.341
R16095 vdd.n2069 vdd.n1938 146.341
R16096 vdd.n2065 vdd.n2064 146.341
R16097 vdd.n2062 vdd.n1944 146.341
R16098 vdd.n2058 vdd.n2057 146.341
R16099 vdd.n2055 vdd.n1951 146.341
R16100 vdd.n2051 vdd.n2050 146.341
R16101 vdd.n2048 vdd.n1958 146.341
R16102 vdd.n2044 vdd.n2043 146.341
R16103 vdd.n2041 vdd.n1965 146.341
R16104 vdd.n1976 vdd.n1973 146.341
R16105 vdd.n2033 vdd.n2032 146.341
R16106 vdd.n2030 vdd.n1978 146.341
R16107 vdd.n2026 vdd.n2025 146.341
R16108 vdd.n2023 vdd.n1984 146.341
R16109 vdd.n2019 vdd.n2018 146.341
R16110 vdd.n2016 vdd.n1991 146.341
R16111 vdd.n2012 vdd.n2011 146.341
R16112 vdd.n2009 vdd.n2006 146.341
R16113 vdd.n2004 vdd.n2001 146.341
R16114 vdd.n1999 vdd.n1069 146.341
R16115 vdd.n1428 vdd.n1188 146.341
R16116 vdd.n1428 vdd.n1184 146.341
R16117 vdd.n1434 vdd.n1184 146.341
R16118 vdd.n1434 vdd.n1176 146.341
R16119 vdd.n1445 vdd.n1176 146.341
R16120 vdd.n1445 vdd.n1172 146.341
R16121 vdd.n1451 vdd.n1172 146.341
R16122 vdd.n1451 vdd.n1166 146.341
R16123 vdd.n1462 vdd.n1166 146.341
R16124 vdd.n1462 vdd.n1162 146.341
R16125 vdd.n1468 vdd.n1162 146.341
R16126 vdd.n1468 vdd.n1153 146.341
R16127 vdd.n1478 vdd.n1153 146.341
R16128 vdd.n1478 vdd.n1149 146.341
R16129 vdd.n1484 vdd.n1149 146.341
R16130 vdd.n1484 vdd.n1142 146.341
R16131 vdd.n1495 vdd.n1142 146.341
R16132 vdd.n1495 vdd.n1138 146.341
R16133 vdd.n1501 vdd.n1138 146.341
R16134 vdd.n1501 vdd.n1131 146.341
R16135 vdd.n1818 vdd.n1131 146.341
R16136 vdd.n1818 vdd.n1127 146.341
R16137 vdd.n1824 vdd.n1127 146.341
R16138 vdd.n1824 vdd.n1119 146.341
R16139 vdd.n1835 vdd.n1119 146.341
R16140 vdd.n1835 vdd.n1115 146.341
R16141 vdd.n1841 vdd.n1115 146.341
R16142 vdd.n1841 vdd.n1109 146.341
R16143 vdd.n1852 vdd.n1109 146.341
R16144 vdd.n1852 vdd.n1105 146.341
R16145 vdd.n1858 vdd.n1105 146.341
R16146 vdd.n1858 vdd.n1096 146.341
R16147 vdd.n1868 vdd.n1096 146.341
R16148 vdd.n1868 vdd.n1092 146.341
R16149 vdd.n1874 vdd.n1092 146.341
R16150 vdd.n1874 vdd.n1086 146.341
R16151 vdd.n1885 vdd.n1086 146.341
R16152 vdd.n1885 vdd.n1081 146.341
R16153 vdd.n1893 vdd.n1081 146.341
R16154 vdd.n1893 vdd.n1071 146.341
R16155 vdd.n2330 vdd.n1071 146.341
R16156 vdd.n1417 vdd.n1193 146.341
R16157 vdd.n1417 vdd.n1226 146.341
R16158 vdd.n1230 vdd.n1229 146.341
R16159 vdd.n1232 vdd.n1231 146.341
R16160 vdd.n1236 vdd.n1235 146.341
R16161 vdd.n1238 vdd.n1237 146.341
R16162 vdd.n1242 vdd.n1241 146.341
R16163 vdd.n1244 vdd.n1243 146.341
R16164 vdd.n1248 vdd.n1247 146.341
R16165 vdd.n1250 vdd.n1249 146.341
R16166 vdd.n1256 vdd.n1255 146.341
R16167 vdd.n1258 vdd.n1257 146.341
R16168 vdd.n1262 vdd.n1261 146.341
R16169 vdd.n1264 vdd.n1263 146.341
R16170 vdd.n1268 vdd.n1267 146.341
R16171 vdd.n1270 vdd.n1269 146.341
R16172 vdd.n1274 vdd.n1273 146.341
R16173 vdd.n1276 vdd.n1275 146.341
R16174 vdd.n1280 vdd.n1279 146.341
R16175 vdd.n1282 vdd.n1281 146.341
R16176 vdd.n1354 vdd.n1285 146.341
R16177 vdd.n1287 vdd.n1286 146.341
R16178 vdd.n1291 vdd.n1290 146.341
R16179 vdd.n1293 vdd.n1292 146.341
R16180 vdd.n1297 vdd.n1296 146.341
R16181 vdd.n1299 vdd.n1298 146.341
R16182 vdd.n1303 vdd.n1302 146.341
R16183 vdd.n1305 vdd.n1304 146.341
R16184 vdd.n1309 vdd.n1308 146.341
R16185 vdd.n1311 vdd.n1310 146.341
R16186 vdd.n1315 vdd.n1314 146.341
R16187 vdd.n1316 vdd.n1224 146.341
R16188 vdd.n1426 vdd.n1189 146.341
R16189 vdd.n1426 vdd.n1182 146.341
R16190 vdd.n1437 vdd.n1182 146.341
R16191 vdd.n1437 vdd.n1178 146.341
R16192 vdd.n1443 vdd.n1178 146.341
R16193 vdd.n1443 vdd.n1171 146.341
R16194 vdd.n1454 vdd.n1171 146.341
R16195 vdd.n1454 vdd.n1167 146.341
R16196 vdd.n1460 vdd.n1167 146.341
R16197 vdd.n1460 vdd.n1160 146.341
R16198 vdd.n1470 vdd.n1160 146.341
R16199 vdd.n1470 vdd.n1156 146.341
R16200 vdd.n1476 vdd.n1156 146.341
R16201 vdd.n1476 vdd.n1148 146.341
R16202 vdd.n1487 vdd.n1148 146.341
R16203 vdd.n1487 vdd.n1144 146.341
R16204 vdd.n1493 vdd.n1144 146.341
R16205 vdd.n1493 vdd.n1137 146.341
R16206 vdd.n1503 vdd.n1137 146.341
R16207 vdd.n1503 vdd.n1133 146.341
R16208 vdd.n1816 vdd.n1133 146.341
R16209 vdd.n1816 vdd.n1125 146.341
R16210 vdd.n1827 vdd.n1125 146.341
R16211 vdd.n1827 vdd.n1121 146.341
R16212 vdd.n1833 vdd.n1121 146.341
R16213 vdd.n1833 vdd.n1114 146.341
R16214 vdd.n1844 vdd.n1114 146.341
R16215 vdd.n1844 vdd.n1110 146.341
R16216 vdd.n1850 vdd.n1110 146.341
R16217 vdd.n1850 vdd.n1103 146.341
R16218 vdd.n1860 vdd.n1103 146.341
R16219 vdd.n1860 vdd.n1099 146.341
R16220 vdd.n1866 vdd.n1099 146.341
R16221 vdd.n1866 vdd.n1091 146.341
R16222 vdd.n1877 vdd.n1091 146.341
R16223 vdd.n1877 vdd.n1087 146.341
R16224 vdd.n1883 vdd.n1087 146.341
R16225 vdd.n1883 vdd.n1079 146.341
R16226 vdd.n1896 vdd.n1079 146.341
R16227 vdd.n1896 vdd.n1074 146.341
R16228 vdd.n2328 vdd.n1074 146.341
R16229 vdd.n1073 vdd.n1049 141.707
R16230 vdd.n3223 vdd.n692 141.707
R16231 vdd.n2177 vdd.t110 127.284
R16232 vdd.n965 vdd.t95 127.284
R16233 vdd.n2151 vdd.t57 127.284
R16234 vdd.n957 vdd.t119 127.284
R16235 vdd.n2922 vdd.t71 127.284
R16236 vdd.n2922 vdd.t72 127.284
R16237 vdd.n2642 vdd.t117 127.284
R16238 vdd.n832 vdd.t99 127.284
R16239 vdd.n2639 vdd.t104 127.284
R16240 vdd.n799 vdd.t106 127.284
R16241 vdd.n1027 vdd.t113 127.284
R16242 vdd.n1027 vdd.t114 127.284
R16243 vdd.n22 vdd.n20 117.314
R16244 vdd.n17 vdd.n15 117.314
R16245 vdd.n27 vdd.n26 116.927
R16246 vdd.n24 vdd.n23 116.927
R16247 vdd.n22 vdd.n21 116.927
R16248 vdd.n17 vdd.n16 116.927
R16249 vdd.n19 vdd.n18 116.927
R16250 vdd.n27 vdd.n25 116.927
R16251 vdd.n2178 vdd.t109 111.188
R16252 vdd.n966 vdd.t96 111.188
R16253 vdd.n2152 vdd.t56 111.188
R16254 vdd.n958 vdd.t120 111.188
R16255 vdd.n2643 vdd.t116 111.188
R16256 vdd.n833 vdd.t100 111.188
R16257 vdd.n2640 vdd.t103 111.188
R16258 vdd.n800 vdd.t107 111.188
R16259 vdd.n2865 vdd.n911 99.5127
R16260 vdd.n2869 vdd.n911 99.5127
R16261 vdd.n2869 vdd.n903 99.5127
R16262 vdd.n2877 vdd.n903 99.5127
R16263 vdd.n2877 vdd.n901 99.5127
R16264 vdd.n2881 vdd.n901 99.5127
R16265 vdd.n2881 vdd.n890 99.5127
R16266 vdd.n2889 vdd.n890 99.5127
R16267 vdd.n2889 vdd.n888 99.5127
R16268 vdd.n2893 vdd.n888 99.5127
R16269 vdd.n2893 vdd.n879 99.5127
R16270 vdd.n2901 vdd.n879 99.5127
R16271 vdd.n2901 vdd.n877 99.5127
R16272 vdd.n2905 vdd.n877 99.5127
R16273 vdd.n2905 vdd.n867 99.5127
R16274 vdd.n2913 vdd.n867 99.5127
R16275 vdd.n2913 vdd.n865 99.5127
R16276 vdd.n2917 vdd.n865 99.5127
R16277 vdd.n2917 vdd.n856 99.5127
R16278 vdd.n2927 vdd.n856 99.5127
R16279 vdd.n2927 vdd.n854 99.5127
R16280 vdd.n2931 vdd.n854 99.5127
R16281 vdd.n2931 vdd.n842 99.5127
R16282 vdd.n2984 vdd.n842 99.5127
R16283 vdd.n2984 vdd.n840 99.5127
R16284 vdd.n2988 vdd.n840 99.5127
R16285 vdd.n2988 vdd.n808 99.5127
R16286 vdd.n3058 vdd.n808 99.5127
R16287 vdd.n3054 vdd.n809 99.5127
R16288 vdd.n3052 vdd.n3051 99.5127
R16289 vdd.n3049 vdd.n813 99.5127
R16290 vdd.n3045 vdd.n3044 99.5127
R16291 vdd.n3042 vdd.n816 99.5127
R16292 vdd.n3038 vdd.n3037 99.5127
R16293 vdd.n3035 vdd.n819 99.5127
R16294 vdd.n3031 vdd.n3030 99.5127
R16295 vdd.n3028 vdd.n3026 99.5127
R16296 vdd.n3024 vdd.n822 99.5127
R16297 vdd.n3020 vdd.n3019 99.5127
R16298 vdd.n3017 vdd.n825 99.5127
R16299 vdd.n3013 vdd.n3012 99.5127
R16300 vdd.n3010 vdd.n828 99.5127
R16301 vdd.n3006 vdd.n3005 99.5127
R16302 vdd.n3003 vdd.n831 99.5127
R16303 vdd.n2998 vdd.n2997 99.5127
R16304 vdd.n2785 vdd.n914 99.5127
R16305 vdd.n2785 vdd.n909 99.5127
R16306 vdd.n2782 vdd.n909 99.5127
R16307 vdd.n2782 vdd.n904 99.5127
R16308 vdd.n2729 vdd.n904 99.5127
R16309 vdd.n2729 vdd.n898 99.5127
R16310 vdd.n2732 vdd.n898 99.5127
R16311 vdd.n2732 vdd.n891 99.5127
R16312 vdd.n2735 vdd.n891 99.5127
R16313 vdd.n2735 vdd.n886 99.5127
R16314 vdd.n2738 vdd.n886 99.5127
R16315 vdd.n2738 vdd.n881 99.5127
R16316 vdd.n2741 vdd.n881 99.5127
R16317 vdd.n2741 vdd.n875 99.5127
R16318 vdd.n2759 vdd.n875 99.5127
R16319 vdd.n2759 vdd.n868 99.5127
R16320 vdd.n2755 vdd.n868 99.5127
R16321 vdd.n2755 vdd.n863 99.5127
R16322 vdd.n2752 vdd.n863 99.5127
R16323 vdd.n2752 vdd.n858 99.5127
R16324 vdd.n2749 vdd.n858 99.5127
R16325 vdd.n2749 vdd.n852 99.5127
R16326 vdd.n2746 vdd.n852 99.5127
R16327 vdd.n2746 vdd.n844 99.5127
R16328 vdd.n844 vdd.n837 99.5127
R16329 vdd.n2990 vdd.n837 99.5127
R16330 vdd.n2991 vdd.n2990 99.5127
R16331 vdd.n2991 vdd.n806 99.5127
R16332 vdd.n2855 vdd.n2638 99.5127
R16333 vdd.n2851 vdd.n2638 99.5127
R16334 vdd.n2849 vdd.n2848 99.5127
R16335 vdd.n2845 vdd.n2844 99.5127
R16336 vdd.n2841 vdd.n2840 99.5127
R16337 vdd.n2837 vdd.n2836 99.5127
R16338 vdd.n2833 vdd.n2832 99.5127
R16339 vdd.n2829 vdd.n2828 99.5127
R16340 vdd.n2825 vdd.n2824 99.5127
R16341 vdd.n2821 vdd.n2820 99.5127
R16342 vdd.n2817 vdd.n2816 99.5127
R16343 vdd.n2813 vdd.n2812 99.5127
R16344 vdd.n2809 vdd.n2808 99.5127
R16345 vdd.n2805 vdd.n2804 99.5127
R16346 vdd.n2801 vdd.n2800 99.5127
R16347 vdd.n2797 vdd.n2796 99.5127
R16348 vdd.n2792 vdd.n2791 99.5127
R16349 vdd.n2603 vdd.n955 99.5127
R16350 vdd.n2599 vdd.n2598 99.5127
R16351 vdd.n2595 vdd.n2594 99.5127
R16352 vdd.n2591 vdd.n2590 99.5127
R16353 vdd.n2587 vdd.n2586 99.5127
R16354 vdd.n2583 vdd.n2582 99.5127
R16355 vdd.n2579 vdd.n2578 99.5127
R16356 vdd.n2575 vdd.n2574 99.5127
R16357 vdd.n2571 vdd.n2570 99.5127
R16358 vdd.n2567 vdd.n2566 99.5127
R16359 vdd.n2563 vdd.n2562 99.5127
R16360 vdd.n2559 vdd.n2558 99.5127
R16361 vdd.n2555 vdd.n2554 99.5127
R16362 vdd.n2551 vdd.n2550 99.5127
R16363 vdd.n2547 vdd.n2546 99.5127
R16364 vdd.n2543 vdd.n2542 99.5127
R16365 vdd.n2538 vdd.n2537 99.5127
R16366 vdd.n2276 vdd.n1050 99.5127
R16367 vdd.n2276 vdd.n1044 99.5127
R16368 vdd.n2273 vdd.n1044 99.5127
R16369 vdd.n2273 vdd.n1038 99.5127
R16370 vdd.n2270 vdd.n1038 99.5127
R16371 vdd.n2270 vdd.n1031 99.5127
R16372 vdd.n2267 vdd.n1031 99.5127
R16373 vdd.n2267 vdd.n1024 99.5127
R16374 vdd.n2264 vdd.n1024 99.5127
R16375 vdd.n2264 vdd.n1019 99.5127
R16376 vdd.n2261 vdd.n1019 99.5127
R16377 vdd.n2261 vdd.n1013 99.5127
R16378 vdd.n2258 vdd.n1013 99.5127
R16379 vdd.n2258 vdd.n1006 99.5127
R16380 vdd.n2172 vdd.n1006 99.5127
R16381 vdd.n2172 vdd.n1000 99.5127
R16382 vdd.n2169 vdd.n1000 99.5127
R16383 vdd.n2169 vdd.n995 99.5127
R16384 vdd.n2166 vdd.n995 99.5127
R16385 vdd.n2166 vdd.n990 99.5127
R16386 vdd.n2163 vdd.n990 99.5127
R16387 vdd.n2163 vdd.n984 99.5127
R16388 vdd.n2160 vdd.n984 99.5127
R16389 vdd.n2160 vdd.n977 99.5127
R16390 vdd.n2157 vdd.n977 99.5127
R16391 vdd.n2157 vdd.n970 99.5127
R16392 vdd.n970 vdd.n960 99.5127
R16393 vdd.n2533 vdd.n960 99.5127
R16394 vdd.n2111 vdd.n2109 99.5127
R16395 vdd.n2115 vdd.n2109 99.5127
R16396 vdd.n2119 vdd.n2117 99.5127
R16397 vdd.n2123 vdd.n2107 99.5127
R16398 vdd.n2127 vdd.n2125 99.5127
R16399 vdd.n2131 vdd.n2105 99.5127
R16400 vdd.n2135 vdd.n2133 99.5127
R16401 vdd.n2139 vdd.n2103 99.5127
R16402 vdd.n2142 vdd.n2141 99.5127
R16403 vdd.n2312 vdd.n2310 99.5127
R16404 vdd.n2308 vdd.n2144 99.5127
R16405 vdd.n2304 vdd.n2302 99.5127
R16406 vdd.n2300 vdd.n2146 99.5127
R16407 vdd.n2296 vdd.n2294 99.5127
R16408 vdd.n2292 vdd.n2148 99.5127
R16409 vdd.n2288 vdd.n2286 99.5127
R16410 vdd.n2284 vdd.n2150 99.5127
R16411 vdd.n2376 vdd.n1046 99.5127
R16412 vdd.n2380 vdd.n1046 99.5127
R16413 vdd.n2380 vdd.n1036 99.5127
R16414 vdd.n2388 vdd.n1036 99.5127
R16415 vdd.n2388 vdd.n1034 99.5127
R16416 vdd.n2392 vdd.n1034 99.5127
R16417 vdd.n2392 vdd.n1023 99.5127
R16418 vdd.n2401 vdd.n1023 99.5127
R16419 vdd.n2401 vdd.n1021 99.5127
R16420 vdd.n2405 vdd.n1021 99.5127
R16421 vdd.n2405 vdd.n1011 99.5127
R16422 vdd.n2413 vdd.n1011 99.5127
R16423 vdd.n2413 vdd.n1009 99.5127
R16424 vdd.n2417 vdd.n1009 99.5127
R16425 vdd.n2417 vdd.n999 99.5127
R16426 vdd.n2425 vdd.n999 99.5127
R16427 vdd.n2425 vdd.n997 99.5127
R16428 vdd.n2429 vdd.n997 99.5127
R16429 vdd.n2429 vdd.n988 99.5127
R16430 vdd.n2437 vdd.n988 99.5127
R16431 vdd.n2437 vdd.n986 99.5127
R16432 vdd.n2441 vdd.n986 99.5127
R16433 vdd.n2441 vdd.n975 99.5127
R16434 vdd.n2451 vdd.n975 99.5127
R16435 vdd.n2451 vdd.n972 99.5127
R16436 vdd.n2456 vdd.n972 99.5127
R16437 vdd.n2456 vdd.n973 99.5127
R16438 vdd.n973 vdd.n954 99.5127
R16439 vdd.n2974 vdd.n2973 99.5127
R16440 vdd.n2971 vdd.n2937 99.5127
R16441 vdd.n2967 vdd.n2966 99.5127
R16442 vdd.n2964 vdd.n2940 99.5127
R16443 vdd.n2960 vdd.n2959 99.5127
R16444 vdd.n2957 vdd.n2943 99.5127
R16445 vdd.n2953 vdd.n2952 99.5127
R16446 vdd.n2950 vdd.n2947 99.5127
R16447 vdd.n3091 vdd.n787 99.5127
R16448 vdd.n3089 vdd.n3088 99.5127
R16449 vdd.n3086 vdd.n789 99.5127
R16450 vdd.n3082 vdd.n3081 99.5127
R16451 vdd.n3079 vdd.n792 99.5127
R16452 vdd.n3075 vdd.n3074 99.5127
R16453 vdd.n3072 vdd.n795 99.5127
R16454 vdd.n3068 vdd.n3067 99.5127
R16455 vdd.n3065 vdd.n798 99.5127
R16456 vdd.n2709 vdd.n915 99.5127
R16457 vdd.n2709 vdd.n910 99.5127
R16458 vdd.n2780 vdd.n910 99.5127
R16459 vdd.n2780 vdd.n905 99.5127
R16460 vdd.n2776 vdd.n905 99.5127
R16461 vdd.n2776 vdd.n899 99.5127
R16462 vdd.n2773 vdd.n899 99.5127
R16463 vdd.n2773 vdd.n892 99.5127
R16464 vdd.n2770 vdd.n892 99.5127
R16465 vdd.n2770 vdd.n887 99.5127
R16466 vdd.n2767 vdd.n887 99.5127
R16467 vdd.n2767 vdd.n882 99.5127
R16468 vdd.n2764 vdd.n882 99.5127
R16469 vdd.n2764 vdd.n876 99.5127
R16470 vdd.n2761 vdd.n876 99.5127
R16471 vdd.n2761 vdd.n869 99.5127
R16472 vdd.n2726 vdd.n869 99.5127
R16473 vdd.n2726 vdd.n864 99.5127
R16474 vdd.n2723 vdd.n864 99.5127
R16475 vdd.n2723 vdd.n859 99.5127
R16476 vdd.n2720 vdd.n859 99.5127
R16477 vdd.n2720 vdd.n853 99.5127
R16478 vdd.n2717 vdd.n853 99.5127
R16479 vdd.n2717 vdd.n845 99.5127
R16480 vdd.n2714 vdd.n845 99.5127
R16481 vdd.n2714 vdd.n838 99.5127
R16482 vdd.n838 vdd.n804 99.5127
R16483 vdd.n3060 vdd.n804 99.5127
R16484 vdd.n2859 vdd.n918 99.5127
R16485 vdd.n2647 vdd.n2646 99.5127
R16486 vdd.n2651 vdd.n2650 99.5127
R16487 vdd.n2655 vdd.n2654 99.5127
R16488 vdd.n2659 vdd.n2658 99.5127
R16489 vdd.n2663 vdd.n2662 99.5127
R16490 vdd.n2667 vdd.n2666 99.5127
R16491 vdd.n2671 vdd.n2670 99.5127
R16492 vdd.n2675 vdd.n2674 99.5127
R16493 vdd.n2679 vdd.n2678 99.5127
R16494 vdd.n2683 vdd.n2682 99.5127
R16495 vdd.n2687 vdd.n2686 99.5127
R16496 vdd.n2691 vdd.n2690 99.5127
R16497 vdd.n2695 vdd.n2694 99.5127
R16498 vdd.n2699 vdd.n2698 99.5127
R16499 vdd.n2703 vdd.n2702 99.5127
R16500 vdd.n2705 vdd.n2637 99.5127
R16501 vdd.n2863 vdd.n908 99.5127
R16502 vdd.n2871 vdd.n908 99.5127
R16503 vdd.n2871 vdd.n906 99.5127
R16504 vdd.n2875 vdd.n906 99.5127
R16505 vdd.n2875 vdd.n896 99.5127
R16506 vdd.n2883 vdd.n896 99.5127
R16507 vdd.n2883 vdd.n894 99.5127
R16508 vdd.n2887 vdd.n894 99.5127
R16509 vdd.n2887 vdd.n885 99.5127
R16510 vdd.n2895 vdd.n885 99.5127
R16511 vdd.n2895 vdd.n883 99.5127
R16512 vdd.n2899 vdd.n883 99.5127
R16513 vdd.n2899 vdd.n873 99.5127
R16514 vdd.n2907 vdd.n873 99.5127
R16515 vdd.n2907 vdd.n871 99.5127
R16516 vdd.n2911 vdd.n871 99.5127
R16517 vdd.n2911 vdd.n862 99.5127
R16518 vdd.n2919 vdd.n862 99.5127
R16519 vdd.n2919 vdd.n860 99.5127
R16520 vdd.n2925 vdd.n860 99.5127
R16521 vdd.n2925 vdd.n850 99.5127
R16522 vdd.n2933 vdd.n850 99.5127
R16523 vdd.n2933 vdd.n847 99.5127
R16524 vdd.n2982 vdd.n847 99.5127
R16525 vdd.n2982 vdd.n848 99.5127
R16526 vdd.n848 vdd.n839 99.5127
R16527 vdd.n2977 vdd.n839 99.5127
R16528 vdd.n2977 vdd.n807 99.5127
R16529 vdd.n2527 vdd.n2526 99.5127
R16530 vdd.n2523 vdd.n2522 99.5127
R16531 vdd.n2519 vdd.n2518 99.5127
R16532 vdd.n2515 vdd.n2514 99.5127
R16533 vdd.n2511 vdd.n2510 99.5127
R16534 vdd.n2507 vdd.n2506 99.5127
R16535 vdd.n2503 vdd.n2502 99.5127
R16536 vdd.n2499 vdd.n2498 99.5127
R16537 vdd.n2495 vdd.n2494 99.5127
R16538 vdd.n2491 vdd.n2490 99.5127
R16539 vdd.n2487 vdd.n2486 99.5127
R16540 vdd.n2483 vdd.n2482 99.5127
R16541 vdd.n2479 vdd.n2478 99.5127
R16542 vdd.n2475 vdd.n2474 99.5127
R16543 vdd.n2471 vdd.n2470 99.5127
R16544 vdd.n2467 vdd.n2466 99.5127
R16545 vdd.n2463 vdd.n936 99.5127
R16546 vdd.n2220 vdd.n1051 99.5127
R16547 vdd.n2220 vdd.n1045 99.5127
R16548 vdd.n2223 vdd.n1045 99.5127
R16549 vdd.n2223 vdd.n1039 99.5127
R16550 vdd.n2226 vdd.n1039 99.5127
R16551 vdd.n2226 vdd.n1032 99.5127
R16552 vdd.n2229 vdd.n1032 99.5127
R16553 vdd.n2229 vdd.n1025 99.5127
R16554 vdd.n2232 vdd.n1025 99.5127
R16555 vdd.n2232 vdd.n1020 99.5127
R16556 vdd.n2235 vdd.n1020 99.5127
R16557 vdd.n2235 vdd.n1014 99.5127
R16558 vdd.n2256 vdd.n1014 99.5127
R16559 vdd.n2256 vdd.n1007 99.5127
R16560 vdd.n2252 vdd.n1007 99.5127
R16561 vdd.n2252 vdd.n1001 99.5127
R16562 vdd.n2249 vdd.n1001 99.5127
R16563 vdd.n2249 vdd.n996 99.5127
R16564 vdd.n2246 vdd.n996 99.5127
R16565 vdd.n2246 vdd.n991 99.5127
R16566 vdd.n2243 vdd.n991 99.5127
R16567 vdd.n2243 vdd.n985 99.5127
R16568 vdd.n2240 vdd.n985 99.5127
R16569 vdd.n2240 vdd.n978 99.5127
R16570 vdd.n978 vdd.n969 99.5127
R16571 vdd.n2458 vdd.n969 99.5127
R16572 vdd.n2459 vdd.n2458 99.5127
R16573 vdd.n2459 vdd.n961 99.5127
R16574 vdd.n2370 vdd.n2368 99.5127
R16575 vdd.n2366 vdd.n1054 99.5127
R16576 vdd.n2362 vdd.n2360 99.5127
R16577 vdd.n2358 vdd.n1056 99.5127
R16578 vdd.n2354 vdd.n2352 99.5127
R16579 vdd.n2350 vdd.n1058 99.5127
R16580 vdd.n2346 vdd.n2344 99.5127
R16581 vdd.n2342 vdd.n1060 99.5127
R16582 vdd.n2184 vdd.n1062 99.5127
R16583 vdd.n2189 vdd.n2186 99.5127
R16584 vdd.n2193 vdd.n2191 99.5127
R16585 vdd.n2197 vdd.n2182 99.5127
R16586 vdd.n2201 vdd.n2199 99.5127
R16587 vdd.n2205 vdd.n2180 99.5127
R16588 vdd.n2209 vdd.n2207 99.5127
R16589 vdd.n2214 vdd.n2176 99.5127
R16590 vdd.n2217 vdd.n2216 99.5127
R16591 vdd.n2374 vdd.n1042 99.5127
R16592 vdd.n2382 vdd.n1042 99.5127
R16593 vdd.n2382 vdd.n1040 99.5127
R16594 vdd.n2386 vdd.n1040 99.5127
R16595 vdd.n2386 vdd.n1029 99.5127
R16596 vdd.n2394 vdd.n1029 99.5127
R16597 vdd.n2394 vdd.n1026 99.5127
R16598 vdd.n2399 vdd.n1026 99.5127
R16599 vdd.n2399 vdd.n1017 99.5127
R16600 vdd.n2407 vdd.n1017 99.5127
R16601 vdd.n2407 vdd.n1015 99.5127
R16602 vdd.n2411 vdd.n1015 99.5127
R16603 vdd.n2411 vdd.n1005 99.5127
R16604 vdd.n2419 vdd.n1005 99.5127
R16605 vdd.n2419 vdd.n1003 99.5127
R16606 vdd.n2423 vdd.n1003 99.5127
R16607 vdd.n2423 vdd.n994 99.5127
R16608 vdd.n2431 vdd.n994 99.5127
R16609 vdd.n2431 vdd.n992 99.5127
R16610 vdd.n2435 vdd.n992 99.5127
R16611 vdd.n2435 vdd.n982 99.5127
R16612 vdd.n2443 vdd.n982 99.5127
R16613 vdd.n2443 vdd.n979 99.5127
R16614 vdd.n2449 vdd.n979 99.5127
R16615 vdd.n2449 vdd.n980 99.5127
R16616 vdd.n980 vdd.n971 99.5127
R16617 vdd.n971 vdd.n962 99.5127
R16618 vdd.n2531 vdd.n962 99.5127
R16619 vdd.n9 vdd.n7 98.9633
R16620 vdd.n2 vdd.n0 98.9633
R16621 vdd.n9 vdd.n8 98.6055
R16622 vdd.n11 vdd.n10 98.6055
R16623 vdd.n13 vdd.n12 98.6055
R16624 vdd.n6 vdd.n5 98.6055
R16625 vdd.n4 vdd.n3 98.6055
R16626 vdd.n2 vdd.n1 98.6055
R16627 vdd.t263 vdd.n303 85.8723
R16628 vdd.t240 vdd.n244 85.8723
R16629 vdd.t252 vdd.n201 85.8723
R16630 vdd.t224 vdd.n142 85.8723
R16631 vdd.t203 vdd.n100 85.8723
R16632 vdd.t141 vdd.n41 85.8723
R16633 vdd.t283 vdd.n1722 85.8723
R16634 vdd.t172 vdd.n1781 85.8723
R16635 vdd.t269 vdd.n1620 85.8723
R16636 vdd.t149 vdd.n1679 85.8723
R16637 vdd.t145 vdd.n1519 85.8723
R16638 vdd.t204 vdd.n1578 85.8723
R16639 vdd.n2923 vdd.n2922 78.546
R16640 vdd.n2397 vdd.n1027 78.546
R16641 vdd.n290 vdd.n289 75.1835
R16642 vdd.n288 vdd.n287 75.1835
R16643 vdd.n286 vdd.n285 75.1835
R16644 vdd.n284 vdd.n283 75.1835
R16645 vdd.n282 vdd.n281 75.1835
R16646 vdd.n280 vdd.n279 75.1835
R16647 vdd.n278 vdd.n277 75.1835
R16648 vdd.n276 vdd.n275 75.1835
R16649 vdd.n274 vdd.n273 75.1835
R16650 vdd.n188 vdd.n187 75.1835
R16651 vdd.n186 vdd.n185 75.1835
R16652 vdd.n184 vdd.n183 75.1835
R16653 vdd.n182 vdd.n181 75.1835
R16654 vdd.n180 vdd.n179 75.1835
R16655 vdd.n178 vdd.n177 75.1835
R16656 vdd.n176 vdd.n175 75.1835
R16657 vdd.n174 vdd.n173 75.1835
R16658 vdd.n172 vdd.n171 75.1835
R16659 vdd.n87 vdd.n86 75.1835
R16660 vdd.n85 vdd.n84 75.1835
R16661 vdd.n83 vdd.n82 75.1835
R16662 vdd.n81 vdd.n80 75.1835
R16663 vdd.n79 vdd.n78 75.1835
R16664 vdd.n77 vdd.n76 75.1835
R16665 vdd.n75 vdd.n74 75.1835
R16666 vdd.n73 vdd.n72 75.1835
R16667 vdd.n71 vdd.n70 75.1835
R16668 vdd.n1752 vdd.n1751 75.1835
R16669 vdd.n1754 vdd.n1753 75.1835
R16670 vdd.n1756 vdd.n1755 75.1835
R16671 vdd.n1758 vdd.n1757 75.1835
R16672 vdd.n1760 vdd.n1759 75.1835
R16673 vdd.n1762 vdd.n1761 75.1835
R16674 vdd.n1764 vdd.n1763 75.1835
R16675 vdd.n1766 vdd.n1765 75.1835
R16676 vdd.n1768 vdd.n1767 75.1835
R16677 vdd.n1650 vdd.n1649 75.1835
R16678 vdd.n1652 vdd.n1651 75.1835
R16679 vdd.n1654 vdd.n1653 75.1835
R16680 vdd.n1656 vdd.n1655 75.1835
R16681 vdd.n1658 vdd.n1657 75.1835
R16682 vdd.n1660 vdd.n1659 75.1835
R16683 vdd.n1662 vdd.n1661 75.1835
R16684 vdd.n1664 vdd.n1663 75.1835
R16685 vdd.n1666 vdd.n1665 75.1835
R16686 vdd.n1549 vdd.n1548 75.1835
R16687 vdd.n1551 vdd.n1550 75.1835
R16688 vdd.n1553 vdd.n1552 75.1835
R16689 vdd.n1555 vdd.n1554 75.1835
R16690 vdd.n1557 vdd.n1556 75.1835
R16691 vdd.n1559 vdd.n1558 75.1835
R16692 vdd.n1561 vdd.n1560 75.1835
R16693 vdd.n1563 vdd.n1562 75.1835
R16694 vdd.n1565 vdd.n1564 75.1835
R16695 vdd.n2858 vdd.n2857 72.8958
R16696 vdd.n2857 vdd.n2621 72.8958
R16697 vdd.n2857 vdd.n2622 72.8958
R16698 vdd.n2857 vdd.n2623 72.8958
R16699 vdd.n2857 vdd.n2624 72.8958
R16700 vdd.n2857 vdd.n2625 72.8958
R16701 vdd.n2857 vdd.n2626 72.8958
R16702 vdd.n2857 vdd.n2627 72.8958
R16703 vdd.n2857 vdd.n2628 72.8958
R16704 vdd.n2857 vdd.n2629 72.8958
R16705 vdd.n2857 vdd.n2630 72.8958
R16706 vdd.n2857 vdd.n2631 72.8958
R16707 vdd.n2857 vdd.n2632 72.8958
R16708 vdd.n2857 vdd.n2633 72.8958
R16709 vdd.n2857 vdd.n2634 72.8958
R16710 vdd.n2857 vdd.n2635 72.8958
R16711 vdd.n2857 vdd.n2636 72.8958
R16712 vdd.n803 vdd.n692 72.8958
R16713 vdd.n3066 vdd.n692 72.8958
R16714 vdd.n797 vdd.n692 72.8958
R16715 vdd.n3073 vdd.n692 72.8958
R16716 vdd.n794 vdd.n692 72.8958
R16717 vdd.n3080 vdd.n692 72.8958
R16718 vdd.n791 vdd.n692 72.8958
R16719 vdd.n3087 vdd.n692 72.8958
R16720 vdd.n3090 vdd.n692 72.8958
R16721 vdd.n2946 vdd.n692 72.8958
R16722 vdd.n2951 vdd.n692 72.8958
R16723 vdd.n2945 vdd.n692 72.8958
R16724 vdd.n2958 vdd.n692 72.8958
R16725 vdd.n2942 vdd.n692 72.8958
R16726 vdd.n2965 vdd.n692 72.8958
R16727 vdd.n2939 vdd.n692 72.8958
R16728 vdd.n2972 vdd.n692 72.8958
R16729 vdd.n2110 vdd.n1049 72.8958
R16730 vdd.n2116 vdd.n1049 72.8958
R16731 vdd.n2118 vdd.n1049 72.8958
R16732 vdd.n2124 vdd.n1049 72.8958
R16733 vdd.n2126 vdd.n1049 72.8958
R16734 vdd.n2132 vdd.n1049 72.8958
R16735 vdd.n2134 vdd.n1049 72.8958
R16736 vdd.n2140 vdd.n1049 72.8958
R16737 vdd.n2311 vdd.n1049 72.8958
R16738 vdd.n2309 vdd.n1049 72.8958
R16739 vdd.n2303 vdd.n1049 72.8958
R16740 vdd.n2301 vdd.n1049 72.8958
R16741 vdd.n2295 vdd.n1049 72.8958
R16742 vdd.n2293 vdd.n1049 72.8958
R16743 vdd.n2287 vdd.n1049 72.8958
R16744 vdd.n2285 vdd.n1049 72.8958
R16745 vdd.n2279 vdd.n1049 72.8958
R16746 vdd.n2604 vdd.n937 72.8958
R16747 vdd.n2604 vdd.n938 72.8958
R16748 vdd.n2604 vdd.n939 72.8958
R16749 vdd.n2604 vdd.n940 72.8958
R16750 vdd.n2604 vdd.n941 72.8958
R16751 vdd.n2604 vdd.n942 72.8958
R16752 vdd.n2604 vdd.n943 72.8958
R16753 vdd.n2604 vdd.n944 72.8958
R16754 vdd.n2604 vdd.n945 72.8958
R16755 vdd.n2604 vdd.n946 72.8958
R16756 vdd.n2604 vdd.n947 72.8958
R16757 vdd.n2604 vdd.n948 72.8958
R16758 vdd.n2604 vdd.n949 72.8958
R16759 vdd.n2604 vdd.n950 72.8958
R16760 vdd.n2604 vdd.n951 72.8958
R16761 vdd.n2604 vdd.n952 72.8958
R16762 vdd.n2604 vdd.n953 72.8958
R16763 vdd.n2857 vdd.n2856 72.8958
R16764 vdd.n2857 vdd.n2605 72.8958
R16765 vdd.n2857 vdd.n2606 72.8958
R16766 vdd.n2857 vdd.n2607 72.8958
R16767 vdd.n2857 vdd.n2608 72.8958
R16768 vdd.n2857 vdd.n2609 72.8958
R16769 vdd.n2857 vdd.n2610 72.8958
R16770 vdd.n2857 vdd.n2611 72.8958
R16771 vdd.n2857 vdd.n2612 72.8958
R16772 vdd.n2857 vdd.n2613 72.8958
R16773 vdd.n2857 vdd.n2614 72.8958
R16774 vdd.n2857 vdd.n2615 72.8958
R16775 vdd.n2857 vdd.n2616 72.8958
R16776 vdd.n2857 vdd.n2617 72.8958
R16777 vdd.n2857 vdd.n2618 72.8958
R16778 vdd.n2857 vdd.n2619 72.8958
R16779 vdd.n2857 vdd.n2620 72.8958
R16780 vdd.n2996 vdd.n692 72.8958
R16781 vdd.n835 vdd.n692 72.8958
R16782 vdd.n3004 vdd.n692 72.8958
R16783 vdd.n830 vdd.n692 72.8958
R16784 vdd.n3011 vdd.n692 72.8958
R16785 vdd.n827 vdd.n692 72.8958
R16786 vdd.n3018 vdd.n692 72.8958
R16787 vdd.n824 vdd.n692 72.8958
R16788 vdd.n3025 vdd.n692 72.8958
R16789 vdd.n3029 vdd.n692 72.8958
R16790 vdd.n821 vdd.n692 72.8958
R16791 vdd.n3036 vdd.n692 72.8958
R16792 vdd.n818 vdd.n692 72.8958
R16793 vdd.n3043 vdd.n692 72.8958
R16794 vdd.n815 vdd.n692 72.8958
R16795 vdd.n3050 vdd.n692 72.8958
R16796 vdd.n3053 vdd.n692 72.8958
R16797 vdd.n2604 vdd.n935 72.8958
R16798 vdd.n2604 vdd.n934 72.8958
R16799 vdd.n2604 vdd.n933 72.8958
R16800 vdd.n2604 vdd.n932 72.8958
R16801 vdd.n2604 vdd.n931 72.8958
R16802 vdd.n2604 vdd.n930 72.8958
R16803 vdd.n2604 vdd.n929 72.8958
R16804 vdd.n2604 vdd.n928 72.8958
R16805 vdd.n2604 vdd.n927 72.8958
R16806 vdd.n2604 vdd.n926 72.8958
R16807 vdd.n2604 vdd.n925 72.8958
R16808 vdd.n2604 vdd.n924 72.8958
R16809 vdd.n2604 vdd.n923 72.8958
R16810 vdd.n2604 vdd.n922 72.8958
R16811 vdd.n2604 vdd.n921 72.8958
R16812 vdd.n2604 vdd.n920 72.8958
R16813 vdd.n2604 vdd.n919 72.8958
R16814 vdd.n2369 vdd.n1049 72.8958
R16815 vdd.n2367 vdd.n1049 72.8958
R16816 vdd.n2361 vdd.n1049 72.8958
R16817 vdd.n2359 vdd.n1049 72.8958
R16818 vdd.n2353 vdd.n1049 72.8958
R16819 vdd.n2351 vdd.n1049 72.8958
R16820 vdd.n2345 vdd.n1049 72.8958
R16821 vdd.n2343 vdd.n1049 72.8958
R16822 vdd.n1061 vdd.n1049 72.8958
R16823 vdd.n2185 vdd.n1049 72.8958
R16824 vdd.n2190 vdd.n1049 72.8958
R16825 vdd.n2192 vdd.n1049 72.8958
R16826 vdd.n2198 vdd.n1049 72.8958
R16827 vdd.n2200 vdd.n1049 72.8958
R16828 vdd.n2206 vdd.n1049 72.8958
R16829 vdd.n2208 vdd.n1049 72.8958
R16830 vdd.n2215 vdd.n1049 72.8958
R16831 vdd.n1419 vdd.n1418 66.2847
R16832 vdd.n1418 vdd.n1194 66.2847
R16833 vdd.n1418 vdd.n1195 66.2847
R16834 vdd.n1418 vdd.n1196 66.2847
R16835 vdd.n1418 vdd.n1197 66.2847
R16836 vdd.n1418 vdd.n1198 66.2847
R16837 vdd.n1418 vdd.n1199 66.2847
R16838 vdd.n1418 vdd.n1200 66.2847
R16839 vdd.n1418 vdd.n1201 66.2847
R16840 vdd.n1418 vdd.n1202 66.2847
R16841 vdd.n1418 vdd.n1203 66.2847
R16842 vdd.n1418 vdd.n1204 66.2847
R16843 vdd.n1418 vdd.n1205 66.2847
R16844 vdd.n1418 vdd.n1206 66.2847
R16845 vdd.n1418 vdd.n1207 66.2847
R16846 vdd.n1418 vdd.n1208 66.2847
R16847 vdd.n1418 vdd.n1209 66.2847
R16848 vdd.n1418 vdd.n1210 66.2847
R16849 vdd.n1418 vdd.n1211 66.2847
R16850 vdd.n1418 vdd.n1212 66.2847
R16851 vdd.n1418 vdd.n1213 66.2847
R16852 vdd.n1418 vdd.n1214 66.2847
R16853 vdd.n1418 vdd.n1215 66.2847
R16854 vdd.n1418 vdd.n1216 66.2847
R16855 vdd.n1418 vdd.n1217 66.2847
R16856 vdd.n1418 vdd.n1218 66.2847
R16857 vdd.n1418 vdd.n1219 66.2847
R16858 vdd.n1418 vdd.n1220 66.2847
R16859 vdd.n1418 vdd.n1221 66.2847
R16860 vdd.n1418 vdd.n1222 66.2847
R16861 vdd.n1418 vdd.n1223 66.2847
R16862 vdd.n1073 vdd.n1070 66.2847
R16863 vdd.n2000 vdd.n1073 66.2847
R16864 vdd.n2005 vdd.n1073 66.2847
R16865 vdd.n2010 vdd.n1073 66.2847
R16866 vdd.n1998 vdd.n1073 66.2847
R16867 vdd.n2017 vdd.n1073 66.2847
R16868 vdd.n1990 vdd.n1073 66.2847
R16869 vdd.n2024 vdd.n1073 66.2847
R16870 vdd.n1983 vdd.n1073 66.2847
R16871 vdd.n2031 vdd.n1073 66.2847
R16872 vdd.n1977 vdd.n1073 66.2847
R16873 vdd.n1972 vdd.n1073 66.2847
R16874 vdd.n2042 vdd.n1073 66.2847
R16875 vdd.n1964 vdd.n1073 66.2847
R16876 vdd.n2049 vdd.n1073 66.2847
R16877 vdd.n1957 vdd.n1073 66.2847
R16878 vdd.n2056 vdd.n1073 66.2847
R16879 vdd.n1950 vdd.n1073 66.2847
R16880 vdd.n2063 vdd.n1073 66.2847
R16881 vdd.n1943 vdd.n1073 66.2847
R16882 vdd.n2070 vdd.n1073 66.2847
R16883 vdd.n1937 vdd.n1073 66.2847
R16884 vdd.n1932 vdd.n1073 66.2847
R16885 vdd.n2081 vdd.n1073 66.2847
R16886 vdd.n1924 vdd.n1073 66.2847
R16887 vdd.n2088 vdd.n1073 66.2847
R16888 vdd.n1917 vdd.n1073 66.2847
R16889 vdd.n2095 vdd.n1073 66.2847
R16890 vdd.n2098 vdd.n1073 66.2847
R16891 vdd.n1908 vdd.n1073 66.2847
R16892 vdd.n2320 vdd.n1073 66.2847
R16893 vdd.n1902 vdd.n1073 66.2847
R16894 vdd.n3223 vdd.n3222 66.2847
R16895 vdd.n3223 vdd.n693 66.2847
R16896 vdd.n3223 vdd.n694 66.2847
R16897 vdd.n3223 vdd.n695 66.2847
R16898 vdd.n3223 vdd.n696 66.2847
R16899 vdd.n3223 vdd.n697 66.2847
R16900 vdd.n3223 vdd.n698 66.2847
R16901 vdd.n3223 vdd.n699 66.2847
R16902 vdd.n3223 vdd.n700 66.2847
R16903 vdd.n3223 vdd.n701 66.2847
R16904 vdd.n3223 vdd.n702 66.2847
R16905 vdd.n3223 vdd.n703 66.2847
R16906 vdd.n3223 vdd.n704 66.2847
R16907 vdd.n3223 vdd.n705 66.2847
R16908 vdd.n3223 vdd.n706 66.2847
R16909 vdd.n3223 vdd.n707 66.2847
R16910 vdd.n3223 vdd.n708 66.2847
R16911 vdd.n3223 vdd.n709 66.2847
R16912 vdd.n3223 vdd.n710 66.2847
R16913 vdd.n3223 vdd.n711 66.2847
R16914 vdd.n3223 vdd.n712 66.2847
R16915 vdd.n3223 vdd.n713 66.2847
R16916 vdd.n3223 vdd.n714 66.2847
R16917 vdd.n3223 vdd.n715 66.2847
R16918 vdd.n3223 vdd.n716 66.2847
R16919 vdd.n3223 vdd.n717 66.2847
R16920 vdd.n3223 vdd.n718 66.2847
R16921 vdd.n3223 vdd.n719 66.2847
R16922 vdd.n3223 vdd.n720 66.2847
R16923 vdd.n3223 vdd.n721 66.2847
R16924 vdd.n3223 vdd.n722 66.2847
R16925 vdd.n3354 vdd.n3353 66.2847
R16926 vdd.n3354 vdd.n424 66.2847
R16927 vdd.n3354 vdd.n423 66.2847
R16928 vdd.n3354 vdd.n422 66.2847
R16929 vdd.n3354 vdd.n421 66.2847
R16930 vdd.n3354 vdd.n420 66.2847
R16931 vdd.n3354 vdd.n419 66.2847
R16932 vdd.n3354 vdd.n418 66.2847
R16933 vdd.n3354 vdd.n417 66.2847
R16934 vdd.n3354 vdd.n416 66.2847
R16935 vdd.n3354 vdd.n415 66.2847
R16936 vdd.n3354 vdd.n414 66.2847
R16937 vdd.n3354 vdd.n413 66.2847
R16938 vdd.n3354 vdd.n412 66.2847
R16939 vdd.n3354 vdd.n411 66.2847
R16940 vdd.n3354 vdd.n410 66.2847
R16941 vdd.n3354 vdd.n409 66.2847
R16942 vdd.n3354 vdd.n408 66.2847
R16943 vdd.n3354 vdd.n407 66.2847
R16944 vdd.n3354 vdd.n406 66.2847
R16945 vdd.n3354 vdd.n405 66.2847
R16946 vdd.n3354 vdd.n404 66.2847
R16947 vdd.n3354 vdd.n403 66.2847
R16948 vdd.n3354 vdd.n402 66.2847
R16949 vdd.n3354 vdd.n401 66.2847
R16950 vdd.n3354 vdd.n400 66.2847
R16951 vdd.n3354 vdd.n399 66.2847
R16952 vdd.n3354 vdd.n398 66.2847
R16953 vdd.n3354 vdd.n397 66.2847
R16954 vdd.n3354 vdd.n396 66.2847
R16955 vdd.n3354 vdd.n395 66.2847
R16956 vdd.n3354 vdd.n394 66.2847
R16957 vdd.n467 vdd.n394 52.4337
R16958 vdd.n473 vdd.n395 52.4337
R16959 vdd.n477 vdd.n396 52.4337
R16960 vdd.n483 vdd.n397 52.4337
R16961 vdd.n487 vdd.n398 52.4337
R16962 vdd.n493 vdd.n399 52.4337
R16963 vdd.n497 vdd.n400 52.4337
R16964 vdd.n503 vdd.n401 52.4337
R16965 vdd.n507 vdd.n402 52.4337
R16966 vdd.n513 vdd.n403 52.4337
R16967 vdd.n517 vdd.n404 52.4337
R16968 vdd.n523 vdd.n405 52.4337
R16969 vdd.n527 vdd.n406 52.4337
R16970 vdd.n533 vdd.n407 52.4337
R16971 vdd.n537 vdd.n408 52.4337
R16972 vdd.n543 vdd.n409 52.4337
R16973 vdd.n547 vdd.n410 52.4337
R16974 vdd.n553 vdd.n411 52.4337
R16975 vdd.n557 vdd.n412 52.4337
R16976 vdd.n563 vdd.n413 52.4337
R16977 vdd.n567 vdd.n414 52.4337
R16978 vdd.n573 vdd.n415 52.4337
R16979 vdd.n577 vdd.n416 52.4337
R16980 vdd.n583 vdd.n417 52.4337
R16981 vdd.n587 vdd.n418 52.4337
R16982 vdd.n593 vdd.n419 52.4337
R16983 vdd.n597 vdd.n420 52.4337
R16984 vdd.n603 vdd.n421 52.4337
R16985 vdd.n607 vdd.n422 52.4337
R16986 vdd.n613 vdd.n423 52.4337
R16987 vdd.n616 vdd.n424 52.4337
R16988 vdd.n3353 vdd.n3352 52.4337
R16989 vdd.n3222 vdd.n3221 52.4337
R16990 vdd.n728 vdd.n693 52.4337
R16991 vdd.n734 vdd.n694 52.4337
R16992 vdd.n3211 vdd.n695 52.4337
R16993 vdd.n3207 vdd.n696 52.4337
R16994 vdd.n3203 vdd.n697 52.4337
R16995 vdd.n3199 vdd.n698 52.4337
R16996 vdd.n3195 vdd.n699 52.4337
R16997 vdd.n3191 vdd.n700 52.4337
R16998 vdd.n3187 vdd.n701 52.4337
R16999 vdd.n3179 vdd.n702 52.4337
R17000 vdd.n3175 vdd.n703 52.4337
R17001 vdd.n3171 vdd.n704 52.4337
R17002 vdd.n3167 vdd.n705 52.4337
R17003 vdd.n3163 vdd.n706 52.4337
R17004 vdd.n3159 vdd.n707 52.4337
R17005 vdd.n3155 vdd.n708 52.4337
R17006 vdd.n3151 vdd.n709 52.4337
R17007 vdd.n3147 vdd.n710 52.4337
R17008 vdd.n3143 vdd.n711 52.4337
R17009 vdd.n3139 vdd.n712 52.4337
R17010 vdd.n3133 vdd.n713 52.4337
R17011 vdd.n3129 vdd.n714 52.4337
R17012 vdd.n3125 vdd.n715 52.4337
R17013 vdd.n3121 vdd.n716 52.4337
R17014 vdd.n3117 vdd.n717 52.4337
R17015 vdd.n3113 vdd.n718 52.4337
R17016 vdd.n3109 vdd.n719 52.4337
R17017 vdd.n3105 vdd.n720 52.4337
R17018 vdd.n3101 vdd.n721 52.4337
R17019 vdd.n3097 vdd.n722 52.4337
R17020 vdd.n2322 vdd.n1902 52.4337
R17021 vdd.n2320 vdd.n2319 52.4337
R17022 vdd.n1909 vdd.n1908 52.4337
R17023 vdd.n2098 vdd.n2097 52.4337
R17024 vdd.n2095 vdd.n2094 52.4337
R17025 vdd.n2090 vdd.n1917 52.4337
R17026 vdd.n2088 vdd.n2087 52.4337
R17027 vdd.n2083 vdd.n1924 52.4337
R17028 vdd.n2081 vdd.n2080 52.4337
R17029 vdd.n1933 vdd.n1932 52.4337
R17030 vdd.n2072 vdd.n1937 52.4337
R17031 vdd.n2070 vdd.n2069 52.4337
R17032 vdd.n2065 vdd.n1943 52.4337
R17033 vdd.n2063 vdd.n2062 52.4337
R17034 vdd.n2058 vdd.n1950 52.4337
R17035 vdd.n2056 vdd.n2055 52.4337
R17036 vdd.n2051 vdd.n1957 52.4337
R17037 vdd.n2049 vdd.n2048 52.4337
R17038 vdd.n2044 vdd.n1964 52.4337
R17039 vdd.n2042 vdd.n2041 52.4337
R17040 vdd.n1973 vdd.n1972 52.4337
R17041 vdd.n2033 vdd.n1977 52.4337
R17042 vdd.n2031 vdd.n2030 52.4337
R17043 vdd.n2026 vdd.n1983 52.4337
R17044 vdd.n2024 vdd.n2023 52.4337
R17045 vdd.n2019 vdd.n1990 52.4337
R17046 vdd.n2017 vdd.n2016 52.4337
R17047 vdd.n2012 vdd.n1998 52.4337
R17048 vdd.n2010 vdd.n2009 52.4337
R17049 vdd.n2005 vdd.n2004 52.4337
R17050 vdd.n2000 vdd.n1999 52.4337
R17051 vdd.n2331 vdd.n1070 52.4337
R17052 vdd.n1420 vdd.n1419 52.4337
R17053 vdd.n1226 vdd.n1194 52.4337
R17054 vdd.n1230 vdd.n1195 52.4337
R17055 vdd.n1232 vdd.n1196 52.4337
R17056 vdd.n1236 vdd.n1197 52.4337
R17057 vdd.n1238 vdd.n1198 52.4337
R17058 vdd.n1242 vdd.n1199 52.4337
R17059 vdd.n1244 vdd.n1200 52.4337
R17060 vdd.n1248 vdd.n1201 52.4337
R17061 vdd.n1250 vdd.n1202 52.4337
R17062 vdd.n1256 vdd.n1203 52.4337
R17063 vdd.n1258 vdd.n1204 52.4337
R17064 vdd.n1262 vdd.n1205 52.4337
R17065 vdd.n1264 vdd.n1206 52.4337
R17066 vdd.n1268 vdd.n1207 52.4337
R17067 vdd.n1270 vdd.n1208 52.4337
R17068 vdd.n1274 vdd.n1209 52.4337
R17069 vdd.n1276 vdd.n1210 52.4337
R17070 vdd.n1280 vdd.n1211 52.4337
R17071 vdd.n1282 vdd.n1212 52.4337
R17072 vdd.n1354 vdd.n1213 52.4337
R17073 vdd.n1287 vdd.n1214 52.4337
R17074 vdd.n1291 vdd.n1215 52.4337
R17075 vdd.n1293 vdd.n1216 52.4337
R17076 vdd.n1297 vdd.n1217 52.4337
R17077 vdd.n1299 vdd.n1218 52.4337
R17078 vdd.n1303 vdd.n1219 52.4337
R17079 vdd.n1305 vdd.n1220 52.4337
R17080 vdd.n1309 vdd.n1221 52.4337
R17081 vdd.n1311 vdd.n1222 52.4337
R17082 vdd.n1315 vdd.n1223 52.4337
R17083 vdd.n1419 vdd.n1193 52.4337
R17084 vdd.n1229 vdd.n1194 52.4337
R17085 vdd.n1231 vdd.n1195 52.4337
R17086 vdd.n1235 vdd.n1196 52.4337
R17087 vdd.n1237 vdd.n1197 52.4337
R17088 vdd.n1241 vdd.n1198 52.4337
R17089 vdd.n1243 vdd.n1199 52.4337
R17090 vdd.n1247 vdd.n1200 52.4337
R17091 vdd.n1249 vdd.n1201 52.4337
R17092 vdd.n1255 vdd.n1202 52.4337
R17093 vdd.n1257 vdd.n1203 52.4337
R17094 vdd.n1261 vdd.n1204 52.4337
R17095 vdd.n1263 vdd.n1205 52.4337
R17096 vdd.n1267 vdd.n1206 52.4337
R17097 vdd.n1269 vdd.n1207 52.4337
R17098 vdd.n1273 vdd.n1208 52.4337
R17099 vdd.n1275 vdd.n1209 52.4337
R17100 vdd.n1279 vdd.n1210 52.4337
R17101 vdd.n1281 vdd.n1211 52.4337
R17102 vdd.n1285 vdd.n1212 52.4337
R17103 vdd.n1286 vdd.n1213 52.4337
R17104 vdd.n1290 vdd.n1214 52.4337
R17105 vdd.n1292 vdd.n1215 52.4337
R17106 vdd.n1296 vdd.n1216 52.4337
R17107 vdd.n1298 vdd.n1217 52.4337
R17108 vdd.n1302 vdd.n1218 52.4337
R17109 vdd.n1304 vdd.n1219 52.4337
R17110 vdd.n1308 vdd.n1220 52.4337
R17111 vdd.n1310 vdd.n1221 52.4337
R17112 vdd.n1314 vdd.n1222 52.4337
R17113 vdd.n1316 vdd.n1223 52.4337
R17114 vdd.n1070 vdd.n1069 52.4337
R17115 vdd.n2001 vdd.n2000 52.4337
R17116 vdd.n2006 vdd.n2005 52.4337
R17117 vdd.n2011 vdd.n2010 52.4337
R17118 vdd.n1998 vdd.n1991 52.4337
R17119 vdd.n2018 vdd.n2017 52.4337
R17120 vdd.n1990 vdd.n1984 52.4337
R17121 vdd.n2025 vdd.n2024 52.4337
R17122 vdd.n1983 vdd.n1978 52.4337
R17123 vdd.n2032 vdd.n2031 52.4337
R17124 vdd.n1977 vdd.n1976 52.4337
R17125 vdd.n1972 vdd.n1965 52.4337
R17126 vdd.n2043 vdd.n2042 52.4337
R17127 vdd.n1964 vdd.n1958 52.4337
R17128 vdd.n2050 vdd.n2049 52.4337
R17129 vdd.n1957 vdd.n1951 52.4337
R17130 vdd.n2057 vdd.n2056 52.4337
R17131 vdd.n1950 vdd.n1944 52.4337
R17132 vdd.n2064 vdd.n2063 52.4337
R17133 vdd.n1943 vdd.n1938 52.4337
R17134 vdd.n2071 vdd.n2070 52.4337
R17135 vdd.n1937 vdd.n1936 52.4337
R17136 vdd.n1932 vdd.n1925 52.4337
R17137 vdd.n2082 vdd.n2081 52.4337
R17138 vdd.n1924 vdd.n1918 52.4337
R17139 vdd.n2089 vdd.n2088 52.4337
R17140 vdd.n1917 vdd.n1911 52.4337
R17141 vdd.n2096 vdd.n2095 52.4337
R17142 vdd.n2099 vdd.n2098 52.4337
R17143 vdd.n1908 vdd.n1903 52.4337
R17144 vdd.n2321 vdd.n2320 52.4337
R17145 vdd.n1902 vdd.n1075 52.4337
R17146 vdd.n3222 vdd.n725 52.4337
R17147 vdd.n733 vdd.n693 52.4337
R17148 vdd.n3212 vdd.n694 52.4337
R17149 vdd.n3208 vdd.n695 52.4337
R17150 vdd.n3204 vdd.n696 52.4337
R17151 vdd.n3200 vdd.n697 52.4337
R17152 vdd.n3196 vdd.n698 52.4337
R17153 vdd.n3192 vdd.n699 52.4337
R17154 vdd.n3188 vdd.n700 52.4337
R17155 vdd.n3178 vdd.n701 52.4337
R17156 vdd.n3176 vdd.n702 52.4337
R17157 vdd.n3172 vdd.n703 52.4337
R17158 vdd.n3168 vdd.n704 52.4337
R17159 vdd.n3164 vdd.n705 52.4337
R17160 vdd.n3160 vdd.n706 52.4337
R17161 vdd.n3156 vdd.n707 52.4337
R17162 vdd.n3152 vdd.n708 52.4337
R17163 vdd.n3148 vdd.n709 52.4337
R17164 vdd.n3144 vdd.n710 52.4337
R17165 vdd.n3140 vdd.n711 52.4337
R17166 vdd.n3132 vdd.n712 52.4337
R17167 vdd.n3130 vdd.n713 52.4337
R17168 vdd.n3126 vdd.n714 52.4337
R17169 vdd.n3122 vdd.n715 52.4337
R17170 vdd.n3118 vdd.n716 52.4337
R17171 vdd.n3114 vdd.n717 52.4337
R17172 vdd.n3110 vdd.n718 52.4337
R17173 vdd.n3106 vdd.n719 52.4337
R17174 vdd.n3102 vdd.n720 52.4337
R17175 vdd.n3098 vdd.n721 52.4337
R17176 vdd.n722 vdd.n691 52.4337
R17177 vdd.n3353 vdd.n425 52.4337
R17178 vdd.n614 vdd.n424 52.4337
R17179 vdd.n608 vdd.n423 52.4337
R17180 vdd.n604 vdd.n422 52.4337
R17181 vdd.n598 vdd.n421 52.4337
R17182 vdd.n594 vdd.n420 52.4337
R17183 vdd.n588 vdd.n419 52.4337
R17184 vdd.n584 vdd.n418 52.4337
R17185 vdd.n578 vdd.n417 52.4337
R17186 vdd.n574 vdd.n416 52.4337
R17187 vdd.n568 vdd.n415 52.4337
R17188 vdd.n564 vdd.n414 52.4337
R17189 vdd.n558 vdd.n413 52.4337
R17190 vdd.n554 vdd.n412 52.4337
R17191 vdd.n548 vdd.n411 52.4337
R17192 vdd.n544 vdd.n410 52.4337
R17193 vdd.n538 vdd.n409 52.4337
R17194 vdd.n534 vdd.n408 52.4337
R17195 vdd.n528 vdd.n407 52.4337
R17196 vdd.n524 vdd.n406 52.4337
R17197 vdd.n518 vdd.n405 52.4337
R17198 vdd.n514 vdd.n404 52.4337
R17199 vdd.n508 vdd.n403 52.4337
R17200 vdd.n504 vdd.n402 52.4337
R17201 vdd.n498 vdd.n401 52.4337
R17202 vdd.n494 vdd.n400 52.4337
R17203 vdd.n488 vdd.n399 52.4337
R17204 vdd.n484 vdd.n398 52.4337
R17205 vdd.n478 vdd.n397 52.4337
R17206 vdd.n474 vdd.n396 52.4337
R17207 vdd.n468 vdd.n395 52.4337
R17208 vdd.n394 vdd.n392 52.4337
R17209 vdd.t48 vdd.t26 51.4683
R17210 vdd.n274 vdd.n272 42.0461
R17211 vdd.n172 vdd.n170 42.0461
R17212 vdd.n71 vdd.n69 42.0461
R17213 vdd.n1752 vdd.n1750 42.0461
R17214 vdd.n1650 vdd.n1648 42.0461
R17215 vdd.n1549 vdd.n1547 42.0461
R17216 vdd.n332 vdd.n331 41.6884
R17217 vdd.n230 vdd.n229 41.6884
R17218 vdd.n129 vdd.n128 41.6884
R17219 vdd.n1810 vdd.n1809 41.6884
R17220 vdd.n1708 vdd.n1707 41.6884
R17221 vdd.n1607 vdd.n1606 41.6884
R17222 vdd.n1319 vdd.n1318 41.1157
R17223 vdd.n1357 vdd.n1356 41.1157
R17224 vdd.n1253 vdd.n1252 41.1157
R17225 vdd.n428 vdd.n427 41.1157
R17226 vdd.n566 vdd.n441 41.1157
R17227 vdd.n454 vdd.n453 41.1157
R17228 vdd.n3053 vdd.n3052 39.2114
R17229 vdd.n3050 vdd.n3049 39.2114
R17230 vdd.n3045 vdd.n815 39.2114
R17231 vdd.n3043 vdd.n3042 39.2114
R17232 vdd.n3038 vdd.n818 39.2114
R17233 vdd.n3036 vdd.n3035 39.2114
R17234 vdd.n3031 vdd.n821 39.2114
R17235 vdd.n3029 vdd.n3028 39.2114
R17236 vdd.n3025 vdd.n3024 39.2114
R17237 vdd.n3020 vdd.n824 39.2114
R17238 vdd.n3018 vdd.n3017 39.2114
R17239 vdd.n3013 vdd.n827 39.2114
R17240 vdd.n3011 vdd.n3010 39.2114
R17241 vdd.n3006 vdd.n830 39.2114
R17242 vdd.n3004 vdd.n3003 39.2114
R17243 vdd.n2998 vdd.n835 39.2114
R17244 vdd.n2996 vdd.n2995 39.2114
R17245 vdd.n2856 vdd.n913 39.2114
R17246 vdd.n2851 vdd.n2605 39.2114
R17247 vdd.n2848 vdd.n2606 39.2114
R17248 vdd.n2844 vdd.n2607 39.2114
R17249 vdd.n2840 vdd.n2608 39.2114
R17250 vdd.n2836 vdd.n2609 39.2114
R17251 vdd.n2832 vdd.n2610 39.2114
R17252 vdd.n2828 vdd.n2611 39.2114
R17253 vdd.n2824 vdd.n2612 39.2114
R17254 vdd.n2820 vdd.n2613 39.2114
R17255 vdd.n2816 vdd.n2614 39.2114
R17256 vdd.n2812 vdd.n2615 39.2114
R17257 vdd.n2808 vdd.n2616 39.2114
R17258 vdd.n2804 vdd.n2617 39.2114
R17259 vdd.n2800 vdd.n2618 39.2114
R17260 vdd.n2796 vdd.n2619 39.2114
R17261 vdd.n2791 vdd.n2620 39.2114
R17262 vdd.n2599 vdd.n953 39.2114
R17263 vdd.n2595 vdd.n952 39.2114
R17264 vdd.n2591 vdd.n951 39.2114
R17265 vdd.n2587 vdd.n950 39.2114
R17266 vdd.n2583 vdd.n949 39.2114
R17267 vdd.n2579 vdd.n948 39.2114
R17268 vdd.n2575 vdd.n947 39.2114
R17269 vdd.n2571 vdd.n946 39.2114
R17270 vdd.n2567 vdd.n945 39.2114
R17271 vdd.n2563 vdd.n944 39.2114
R17272 vdd.n2559 vdd.n943 39.2114
R17273 vdd.n2555 vdd.n942 39.2114
R17274 vdd.n2551 vdd.n941 39.2114
R17275 vdd.n2547 vdd.n940 39.2114
R17276 vdd.n2543 vdd.n939 39.2114
R17277 vdd.n2538 vdd.n938 39.2114
R17278 vdd.n2534 vdd.n937 39.2114
R17279 vdd.n2110 vdd.n1048 39.2114
R17280 vdd.n2116 vdd.n2115 39.2114
R17281 vdd.n2119 vdd.n2118 39.2114
R17282 vdd.n2124 vdd.n2123 39.2114
R17283 vdd.n2127 vdd.n2126 39.2114
R17284 vdd.n2132 vdd.n2131 39.2114
R17285 vdd.n2135 vdd.n2134 39.2114
R17286 vdd.n2140 vdd.n2139 39.2114
R17287 vdd.n2311 vdd.n2142 39.2114
R17288 vdd.n2310 vdd.n2309 39.2114
R17289 vdd.n2303 vdd.n2144 39.2114
R17290 vdd.n2302 vdd.n2301 39.2114
R17291 vdd.n2295 vdd.n2146 39.2114
R17292 vdd.n2294 vdd.n2293 39.2114
R17293 vdd.n2287 vdd.n2148 39.2114
R17294 vdd.n2286 vdd.n2285 39.2114
R17295 vdd.n2279 vdd.n2150 39.2114
R17296 vdd.n2972 vdd.n2971 39.2114
R17297 vdd.n2967 vdd.n2939 39.2114
R17298 vdd.n2965 vdd.n2964 39.2114
R17299 vdd.n2960 vdd.n2942 39.2114
R17300 vdd.n2958 vdd.n2957 39.2114
R17301 vdd.n2953 vdd.n2945 39.2114
R17302 vdd.n2951 vdd.n2950 39.2114
R17303 vdd.n2946 vdd.n787 39.2114
R17304 vdd.n3090 vdd.n3089 39.2114
R17305 vdd.n3087 vdd.n3086 39.2114
R17306 vdd.n3082 vdd.n791 39.2114
R17307 vdd.n3080 vdd.n3079 39.2114
R17308 vdd.n3075 vdd.n794 39.2114
R17309 vdd.n3073 vdd.n3072 39.2114
R17310 vdd.n3068 vdd.n797 39.2114
R17311 vdd.n3066 vdd.n3065 39.2114
R17312 vdd.n3061 vdd.n803 39.2114
R17313 vdd.n2858 vdd.n916 39.2114
R17314 vdd.n2621 vdd.n918 39.2114
R17315 vdd.n2647 vdd.n2622 39.2114
R17316 vdd.n2651 vdd.n2623 39.2114
R17317 vdd.n2655 vdd.n2624 39.2114
R17318 vdd.n2659 vdd.n2625 39.2114
R17319 vdd.n2663 vdd.n2626 39.2114
R17320 vdd.n2667 vdd.n2627 39.2114
R17321 vdd.n2671 vdd.n2628 39.2114
R17322 vdd.n2675 vdd.n2629 39.2114
R17323 vdd.n2679 vdd.n2630 39.2114
R17324 vdd.n2683 vdd.n2631 39.2114
R17325 vdd.n2687 vdd.n2632 39.2114
R17326 vdd.n2691 vdd.n2633 39.2114
R17327 vdd.n2695 vdd.n2634 39.2114
R17328 vdd.n2699 vdd.n2635 39.2114
R17329 vdd.n2703 vdd.n2636 39.2114
R17330 vdd.n2859 vdd.n2858 39.2114
R17331 vdd.n2646 vdd.n2621 39.2114
R17332 vdd.n2650 vdd.n2622 39.2114
R17333 vdd.n2654 vdd.n2623 39.2114
R17334 vdd.n2658 vdd.n2624 39.2114
R17335 vdd.n2662 vdd.n2625 39.2114
R17336 vdd.n2666 vdd.n2626 39.2114
R17337 vdd.n2670 vdd.n2627 39.2114
R17338 vdd.n2674 vdd.n2628 39.2114
R17339 vdd.n2678 vdd.n2629 39.2114
R17340 vdd.n2682 vdd.n2630 39.2114
R17341 vdd.n2686 vdd.n2631 39.2114
R17342 vdd.n2690 vdd.n2632 39.2114
R17343 vdd.n2694 vdd.n2633 39.2114
R17344 vdd.n2698 vdd.n2634 39.2114
R17345 vdd.n2702 vdd.n2635 39.2114
R17346 vdd.n2705 vdd.n2636 39.2114
R17347 vdd.n803 vdd.n798 39.2114
R17348 vdd.n3067 vdd.n3066 39.2114
R17349 vdd.n797 vdd.n795 39.2114
R17350 vdd.n3074 vdd.n3073 39.2114
R17351 vdd.n794 vdd.n792 39.2114
R17352 vdd.n3081 vdd.n3080 39.2114
R17353 vdd.n791 vdd.n789 39.2114
R17354 vdd.n3088 vdd.n3087 39.2114
R17355 vdd.n3091 vdd.n3090 39.2114
R17356 vdd.n2947 vdd.n2946 39.2114
R17357 vdd.n2952 vdd.n2951 39.2114
R17358 vdd.n2945 vdd.n2943 39.2114
R17359 vdd.n2959 vdd.n2958 39.2114
R17360 vdd.n2942 vdd.n2940 39.2114
R17361 vdd.n2966 vdd.n2965 39.2114
R17362 vdd.n2939 vdd.n2937 39.2114
R17363 vdd.n2973 vdd.n2972 39.2114
R17364 vdd.n2111 vdd.n2110 39.2114
R17365 vdd.n2117 vdd.n2116 39.2114
R17366 vdd.n2118 vdd.n2107 39.2114
R17367 vdd.n2125 vdd.n2124 39.2114
R17368 vdd.n2126 vdd.n2105 39.2114
R17369 vdd.n2133 vdd.n2132 39.2114
R17370 vdd.n2134 vdd.n2103 39.2114
R17371 vdd.n2141 vdd.n2140 39.2114
R17372 vdd.n2312 vdd.n2311 39.2114
R17373 vdd.n2309 vdd.n2308 39.2114
R17374 vdd.n2304 vdd.n2303 39.2114
R17375 vdd.n2301 vdd.n2300 39.2114
R17376 vdd.n2296 vdd.n2295 39.2114
R17377 vdd.n2293 vdd.n2292 39.2114
R17378 vdd.n2288 vdd.n2287 39.2114
R17379 vdd.n2285 vdd.n2284 39.2114
R17380 vdd.n2280 vdd.n2279 39.2114
R17381 vdd.n2537 vdd.n937 39.2114
R17382 vdd.n2542 vdd.n938 39.2114
R17383 vdd.n2546 vdd.n939 39.2114
R17384 vdd.n2550 vdd.n940 39.2114
R17385 vdd.n2554 vdd.n941 39.2114
R17386 vdd.n2558 vdd.n942 39.2114
R17387 vdd.n2562 vdd.n943 39.2114
R17388 vdd.n2566 vdd.n944 39.2114
R17389 vdd.n2570 vdd.n945 39.2114
R17390 vdd.n2574 vdd.n946 39.2114
R17391 vdd.n2578 vdd.n947 39.2114
R17392 vdd.n2582 vdd.n948 39.2114
R17393 vdd.n2586 vdd.n949 39.2114
R17394 vdd.n2590 vdd.n950 39.2114
R17395 vdd.n2594 vdd.n951 39.2114
R17396 vdd.n2598 vdd.n952 39.2114
R17397 vdd.n955 vdd.n953 39.2114
R17398 vdd.n2856 vdd.n2855 39.2114
R17399 vdd.n2849 vdd.n2605 39.2114
R17400 vdd.n2845 vdd.n2606 39.2114
R17401 vdd.n2841 vdd.n2607 39.2114
R17402 vdd.n2837 vdd.n2608 39.2114
R17403 vdd.n2833 vdd.n2609 39.2114
R17404 vdd.n2829 vdd.n2610 39.2114
R17405 vdd.n2825 vdd.n2611 39.2114
R17406 vdd.n2821 vdd.n2612 39.2114
R17407 vdd.n2817 vdd.n2613 39.2114
R17408 vdd.n2813 vdd.n2614 39.2114
R17409 vdd.n2809 vdd.n2615 39.2114
R17410 vdd.n2805 vdd.n2616 39.2114
R17411 vdd.n2801 vdd.n2617 39.2114
R17412 vdd.n2797 vdd.n2618 39.2114
R17413 vdd.n2792 vdd.n2619 39.2114
R17414 vdd.n2788 vdd.n2620 39.2114
R17415 vdd.n2997 vdd.n2996 39.2114
R17416 vdd.n835 vdd.n831 39.2114
R17417 vdd.n3005 vdd.n3004 39.2114
R17418 vdd.n830 vdd.n828 39.2114
R17419 vdd.n3012 vdd.n3011 39.2114
R17420 vdd.n827 vdd.n825 39.2114
R17421 vdd.n3019 vdd.n3018 39.2114
R17422 vdd.n824 vdd.n822 39.2114
R17423 vdd.n3026 vdd.n3025 39.2114
R17424 vdd.n3030 vdd.n3029 39.2114
R17425 vdd.n821 vdd.n819 39.2114
R17426 vdd.n3037 vdd.n3036 39.2114
R17427 vdd.n818 vdd.n816 39.2114
R17428 vdd.n3044 vdd.n3043 39.2114
R17429 vdd.n815 vdd.n813 39.2114
R17430 vdd.n3051 vdd.n3050 39.2114
R17431 vdd.n3054 vdd.n3053 39.2114
R17432 vdd.n963 vdd.n919 39.2114
R17433 vdd.n2526 vdd.n920 39.2114
R17434 vdd.n2522 vdd.n921 39.2114
R17435 vdd.n2518 vdd.n922 39.2114
R17436 vdd.n2514 vdd.n923 39.2114
R17437 vdd.n2510 vdd.n924 39.2114
R17438 vdd.n2506 vdd.n925 39.2114
R17439 vdd.n2502 vdd.n926 39.2114
R17440 vdd.n2498 vdd.n927 39.2114
R17441 vdd.n2494 vdd.n928 39.2114
R17442 vdd.n2490 vdd.n929 39.2114
R17443 vdd.n2486 vdd.n930 39.2114
R17444 vdd.n2482 vdd.n931 39.2114
R17445 vdd.n2478 vdd.n932 39.2114
R17446 vdd.n2474 vdd.n933 39.2114
R17447 vdd.n2470 vdd.n934 39.2114
R17448 vdd.n2466 vdd.n935 39.2114
R17449 vdd.n2369 vdd.n1052 39.2114
R17450 vdd.n2368 vdd.n2367 39.2114
R17451 vdd.n2361 vdd.n1054 39.2114
R17452 vdd.n2360 vdd.n2359 39.2114
R17453 vdd.n2353 vdd.n1056 39.2114
R17454 vdd.n2352 vdd.n2351 39.2114
R17455 vdd.n2345 vdd.n1058 39.2114
R17456 vdd.n2344 vdd.n2343 39.2114
R17457 vdd.n1061 vdd.n1060 39.2114
R17458 vdd.n2185 vdd.n2184 39.2114
R17459 vdd.n2190 vdd.n2189 39.2114
R17460 vdd.n2193 vdd.n2192 39.2114
R17461 vdd.n2198 vdd.n2197 39.2114
R17462 vdd.n2201 vdd.n2200 39.2114
R17463 vdd.n2206 vdd.n2205 39.2114
R17464 vdd.n2209 vdd.n2208 39.2114
R17465 vdd.n2215 vdd.n2214 39.2114
R17466 vdd.n2463 vdd.n935 39.2114
R17467 vdd.n2467 vdd.n934 39.2114
R17468 vdd.n2471 vdd.n933 39.2114
R17469 vdd.n2475 vdd.n932 39.2114
R17470 vdd.n2479 vdd.n931 39.2114
R17471 vdd.n2483 vdd.n930 39.2114
R17472 vdd.n2487 vdd.n929 39.2114
R17473 vdd.n2491 vdd.n928 39.2114
R17474 vdd.n2495 vdd.n927 39.2114
R17475 vdd.n2499 vdd.n926 39.2114
R17476 vdd.n2503 vdd.n925 39.2114
R17477 vdd.n2507 vdd.n924 39.2114
R17478 vdd.n2511 vdd.n923 39.2114
R17479 vdd.n2515 vdd.n922 39.2114
R17480 vdd.n2519 vdd.n921 39.2114
R17481 vdd.n2523 vdd.n920 39.2114
R17482 vdd.n2527 vdd.n919 39.2114
R17483 vdd.n2370 vdd.n2369 39.2114
R17484 vdd.n2367 vdd.n2366 39.2114
R17485 vdd.n2362 vdd.n2361 39.2114
R17486 vdd.n2359 vdd.n2358 39.2114
R17487 vdd.n2354 vdd.n2353 39.2114
R17488 vdd.n2351 vdd.n2350 39.2114
R17489 vdd.n2346 vdd.n2345 39.2114
R17490 vdd.n2343 vdd.n2342 39.2114
R17491 vdd.n1062 vdd.n1061 39.2114
R17492 vdd.n2186 vdd.n2185 39.2114
R17493 vdd.n2191 vdd.n2190 39.2114
R17494 vdd.n2192 vdd.n2182 39.2114
R17495 vdd.n2199 vdd.n2198 39.2114
R17496 vdd.n2200 vdd.n2180 39.2114
R17497 vdd.n2207 vdd.n2206 39.2114
R17498 vdd.n2208 vdd.n2176 39.2114
R17499 vdd.n2216 vdd.n2215 39.2114
R17500 vdd.n2335 vdd.n2334 37.2369
R17501 vdd.n2038 vdd.n1971 37.2369
R17502 vdd.n2077 vdd.n1931 37.2369
R17503 vdd.n3138 vdd.n769 37.2369
R17504 vdd.n3186 vdd.n3185 37.2369
R17505 vdd.n690 vdd.n689 37.2369
R17506 vdd.n2377 vdd.n1047 31.6883
R17507 vdd.n2602 vdd.n956 31.6883
R17508 vdd.n2535 vdd.n959 31.6883
R17509 vdd.n2281 vdd.n2278 31.6883
R17510 vdd.n2789 vdd.n2787 31.6883
R17511 vdd.n2994 vdd.n2993 31.6883
R17512 vdd.n2866 vdd.n912 31.6883
R17513 vdd.n3057 vdd.n3056 31.6883
R17514 vdd.n2976 vdd.n2975 31.6883
R17515 vdd.n3062 vdd.n802 31.6883
R17516 vdd.n2708 vdd.n2707 31.6883
R17517 vdd.n2862 vdd.n2861 31.6883
R17518 vdd.n2373 vdd.n2372 31.6883
R17519 vdd.n2530 vdd.n2529 31.6883
R17520 vdd.n2462 vdd.n2461 31.6883
R17521 vdd.n2219 vdd.n2218 31.6883
R17522 vdd.n2212 vdd.n2178 30.449
R17523 vdd.n967 vdd.n966 30.449
R17524 vdd.n2153 vdd.n2152 30.449
R17525 vdd.n2540 vdd.n958 30.449
R17526 vdd.n2644 vdd.n2643 30.449
R17527 vdd.n3000 vdd.n833 30.449
R17528 vdd.n2794 vdd.n2640 30.449
R17529 vdd.n801 vdd.n800 30.449
R17530 vdd.n1418 vdd.n1225 22.2201
R17531 vdd.n2329 vdd.n1073 22.2201
R17532 vdd.n3223 vdd.n723 22.2201
R17533 vdd.n3355 vdd.n3354 22.2201
R17534 vdd.n1429 vdd.n1187 19.3944
R17535 vdd.n1429 vdd.n1185 19.3944
R17536 vdd.n1433 vdd.n1185 19.3944
R17537 vdd.n1433 vdd.n1175 19.3944
R17538 vdd.n1446 vdd.n1175 19.3944
R17539 vdd.n1446 vdd.n1173 19.3944
R17540 vdd.n1450 vdd.n1173 19.3944
R17541 vdd.n1450 vdd.n1165 19.3944
R17542 vdd.n1463 vdd.n1165 19.3944
R17543 vdd.n1463 vdd.n1163 19.3944
R17544 vdd.n1467 vdd.n1163 19.3944
R17545 vdd.n1467 vdd.n1152 19.3944
R17546 vdd.n1479 vdd.n1152 19.3944
R17547 vdd.n1479 vdd.n1150 19.3944
R17548 vdd.n1483 vdd.n1150 19.3944
R17549 vdd.n1483 vdd.n1141 19.3944
R17550 vdd.n1496 vdd.n1141 19.3944
R17551 vdd.n1496 vdd.n1139 19.3944
R17552 vdd.n1500 vdd.n1139 19.3944
R17553 vdd.n1500 vdd.n1130 19.3944
R17554 vdd.n1819 vdd.n1130 19.3944
R17555 vdd.n1819 vdd.n1128 19.3944
R17556 vdd.n1823 vdd.n1128 19.3944
R17557 vdd.n1823 vdd.n1118 19.3944
R17558 vdd.n1836 vdd.n1118 19.3944
R17559 vdd.n1836 vdd.n1116 19.3944
R17560 vdd.n1840 vdd.n1116 19.3944
R17561 vdd.n1840 vdd.n1108 19.3944
R17562 vdd.n1853 vdd.n1108 19.3944
R17563 vdd.n1853 vdd.n1106 19.3944
R17564 vdd.n1857 vdd.n1106 19.3944
R17565 vdd.n1857 vdd.n1095 19.3944
R17566 vdd.n1869 vdd.n1095 19.3944
R17567 vdd.n1869 vdd.n1093 19.3944
R17568 vdd.n1873 vdd.n1093 19.3944
R17569 vdd.n1873 vdd.n1085 19.3944
R17570 vdd.n1886 vdd.n1085 19.3944
R17571 vdd.n1886 vdd.n1082 19.3944
R17572 vdd.n1892 vdd.n1082 19.3944
R17573 vdd.n1892 vdd.n1083 19.3944
R17574 vdd.n1083 vdd.n1072 19.3944
R17575 vdd.n1353 vdd.n1288 19.3944
R17576 vdd.n1349 vdd.n1288 19.3944
R17577 vdd.n1349 vdd.n1348 19.3944
R17578 vdd.n1348 vdd.n1347 19.3944
R17579 vdd.n1347 vdd.n1294 19.3944
R17580 vdd.n1343 vdd.n1294 19.3944
R17581 vdd.n1343 vdd.n1342 19.3944
R17582 vdd.n1342 vdd.n1341 19.3944
R17583 vdd.n1341 vdd.n1300 19.3944
R17584 vdd.n1337 vdd.n1300 19.3944
R17585 vdd.n1337 vdd.n1336 19.3944
R17586 vdd.n1336 vdd.n1335 19.3944
R17587 vdd.n1335 vdd.n1306 19.3944
R17588 vdd.n1331 vdd.n1306 19.3944
R17589 vdd.n1331 vdd.n1330 19.3944
R17590 vdd.n1330 vdd.n1329 19.3944
R17591 vdd.n1329 vdd.n1312 19.3944
R17592 vdd.n1325 vdd.n1312 19.3944
R17593 vdd.n1325 vdd.n1324 19.3944
R17594 vdd.n1324 vdd.n1323 19.3944
R17595 vdd.n1388 vdd.n1387 19.3944
R17596 vdd.n1387 vdd.n1386 19.3944
R17597 vdd.n1386 vdd.n1259 19.3944
R17598 vdd.n1382 vdd.n1259 19.3944
R17599 vdd.n1382 vdd.n1381 19.3944
R17600 vdd.n1381 vdd.n1380 19.3944
R17601 vdd.n1380 vdd.n1265 19.3944
R17602 vdd.n1376 vdd.n1265 19.3944
R17603 vdd.n1376 vdd.n1375 19.3944
R17604 vdd.n1375 vdd.n1374 19.3944
R17605 vdd.n1374 vdd.n1271 19.3944
R17606 vdd.n1370 vdd.n1271 19.3944
R17607 vdd.n1370 vdd.n1369 19.3944
R17608 vdd.n1369 vdd.n1368 19.3944
R17609 vdd.n1368 vdd.n1277 19.3944
R17610 vdd.n1364 vdd.n1277 19.3944
R17611 vdd.n1364 vdd.n1363 19.3944
R17612 vdd.n1363 vdd.n1362 19.3944
R17613 vdd.n1362 vdd.n1283 19.3944
R17614 vdd.n1358 vdd.n1283 19.3944
R17615 vdd.n1421 vdd.n1192 19.3944
R17616 vdd.n1416 vdd.n1192 19.3944
R17617 vdd.n1416 vdd.n1227 19.3944
R17618 vdd.n1412 vdd.n1227 19.3944
R17619 vdd.n1412 vdd.n1411 19.3944
R17620 vdd.n1411 vdd.n1410 19.3944
R17621 vdd.n1410 vdd.n1233 19.3944
R17622 vdd.n1406 vdd.n1233 19.3944
R17623 vdd.n1406 vdd.n1405 19.3944
R17624 vdd.n1405 vdd.n1404 19.3944
R17625 vdd.n1404 vdd.n1239 19.3944
R17626 vdd.n1400 vdd.n1239 19.3944
R17627 vdd.n1400 vdd.n1399 19.3944
R17628 vdd.n1399 vdd.n1398 19.3944
R17629 vdd.n1398 vdd.n1245 19.3944
R17630 vdd.n1394 vdd.n1245 19.3944
R17631 vdd.n1394 vdd.n1393 19.3944
R17632 vdd.n1393 vdd.n1392 19.3944
R17633 vdd.n2034 vdd.n1969 19.3944
R17634 vdd.n2034 vdd.n1975 19.3944
R17635 vdd.n2029 vdd.n1975 19.3944
R17636 vdd.n2029 vdd.n2028 19.3944
R17637 vdd.n2028 vdd.n2027 19.3944
R17638 vdd.n2027 vdd.n1982 19.3944
R17639 vdd.n2022 vdd.n1982 19.3944
R17640 vdd.n2022 vdd.n2021 19.3944
R17641 vdd.n2021 vdd.n2020 19.3944
R17642 vdd.n2020 vdd.n1989 19.3944
R17643 vdd.n2015 vdd.n1989 19.3944
R17644 vdd.n2015 vdd.n2014 19.3944
R17645 vdd.n2014 vdd.n2013 19.3944
R17646 vdd.n2013 vdd.n1997 19.3944
R17647 vdd.n2008 vdd.n1997 19.3944
R17648 vdd.n2008 vdd.n2007 19.3944
R17649 vdd.n2003 vdd.n2002 19.3944
R17650 vdd.n2336 vdd.n1068 19.3944
R17651 vdd.n2073 vdd.n1929 19.3944
R17652 vdd.n2073 vdd.n1935 19.3944
R17653 vdd.n2068 vdd.n1935 19.3944
R17654 vdd.n2068 vdd.n2067 19.3944
R17655 vdd.n2067 vdd.n2066 19.3944
R17656 vdd.n2066 vdd.n1942 19.3944
R17657 vdd.n2061 vdd.n1942 19.3944
R17658 vdd.n2061 vdd.n2060 19.3944
R17659 vdd.n2060 vdd.n2059 19.3944
R17660 vdd.n2059 vdd.n1949 19.3944
R17661 vdd.n2054 vdd.n1949 19.3944
R17662 vdd.n2054 vdd.n2053 19.3944
R17663 vdd.n2053 vdd.n2052 19.3944
R17664 vdd.n2052 vdd.n1956 19.3944
R17665 vdd.n2047 vdd.n1956 19.3944
R17666 vdd.n2047 vdd.n2046 19.3944
R17667 vdd.n2046 vdd.n2045 19.3944
R17668 vdd.n2045 vdd.n1963 19.3944
R17669 vdd.n2040 vdd.n1963 19.3944
R17670 vdd.n2040 vdd.n2039 19.3944
R17671 vdd.n2324 vdd.n2323 19.3944
R17672 vdd.n2323 vdd.n1901 19.3944
R17673 vdd.n2318 vdd.n2317 19.3944
R17674 vdd.n2100 vdd.n1905 19.3944
R17675 vdd.n2100 vdd.n1907 19.3944
R17676 vdd.n1910 vdd.n1907 19.3944
R17677 vdd.n2093 vdd.n1910 19.3944
R17678 vdd.n2093 vdd.n2092 19.3944
R17679 vdd.n2092 vdd.n2091 19.3944
R17680 vdd.n2091 vdd.n1916 19.3944
R17681 vdd.n2086 vdd.n1916 19.3944
R17682 vdd.n2086 vdd.n2085 19.3944
R17683 vdd.n2085 vdd.n2084 19.3944
R17684 vdd.n2084 vdd.n1923 19.3944
R17685 vdd.n2079 vdd.n1923 19.3944
R17686 vdd.n2079 vdd.n2078 19.3944
R17687 vdd.n1425 vdd.n1190 19.3944
R17688 vdd.n1425 vdd.n1181 19.3944
R17689 vdd.n1438 vdd.n1181 19.3944
R17690 vdd.n1438 vdd.n1179 19.3944
R17691 vdd.n1442 vdd.n1179 19.3944
R17692 vdd.n1442 vdd.n1170 19.3944
R17693 vdd.n1455 vdd.n1170 19.3944
R17694 vdd.n1455 vdd.n1168 19.3944
R17695 vdd.n1459 vdd.n1168 19.3944
R17696 vdd.n1459 vdd.n1159 19.3944
R17697 vdd.n1471 vdd.n1159 19.3944
R17698 vdd.n1471 vdd.n1157 19.3944
R17699 vdd.n1475 vdd.n1157 19.3944
R17700 vdd.n1475 vdd.n1147 19.3944
R17701 vdd.n1488 vdd.n1147 19.3944
R17702 vdd.n1488 vdd.n1145 19.3944
R17703 vdd.n1492 vdd.n1145 19.3944
R17704 vdd.n1492 vdd.n1136 19.3944
R17705 vdd.n1504 vdd.n1136 19.3944
R17706 vdd.n1504 vdd.n1134 19.3944
R17707 vdd.n1815 vdd.n1134 19.3944
R17708 vdd.n1815 vdd.n1124 19.3944
R17709 vdd.n1828 vdd.n1124 19.3944
R17710 vdd.n1828 vdd.n1122 19.3944
R17711 vdd.n1832 vdd.n1122 19.3944
R17712 vdd.n1832 vdd.n1113 19.3944
R17713 vdd.n1845 vdd.n1113 19.3944
R17714 vdd.n1845 vdd.n1111 19.3944
R17715 vdd.n1849 vdd.n1111 19.3944
R17716 vdd.n1849 vdd.n1102 19.3944
R17717 vdd.n1861 vdd.n1102 19.3944
R17718 vdd.n1861 vdd.n1100 19.3944
R17719 vdd.n1865 vdd.n1100 19.3944
R17720 vdd.n1865 vdd.n1090 19.3944
R17721 vdd.n1878 vdd.n1090 19.3944
R17722 vdd.n1878 vdd.n1088 19.3944
R17723 vdd.n1882 vdd.n1088 19.3944
R17724 vdd.n1882 vdd.n1078 19.3944
R17725 vdd.n1897 vdd.n1078 19.3944
R17726 vdd.n1897 vdd.n1076 19.3944
R17727 vdd.n2327 vdd.n1076 19.3944
R17728 vdd.n3229 vdd.n686 19.3944
R17729 vdd.n3229 vdd.n676 19.3944
R17730 vdd.n3241 vdd.n676 19.3944
R17731 vdd.n3241 vdd.n674 19.3944
R17732 vdd.n3245 vdd.n674 19.3944
R17733 vdd.n3245 vdd.n666 19.3944
R17734 vdd.n3258 vdd.n666 19.3944
R17735 vdd.n3258 vdd.n664 19.3944
R17736 vdd.n3262 vdd.n664 19.3944
R17737 vdd.n3262 vdd.n653 19.3944
R17738 vdd.n3274 vdd.n653 19.3944
R17739 vdd.n3274 vdd.n651 19.3944
R17740 vdd.n3278 vdd.n651 19.3944
R17741 vdd.n3278 vdd.n642 19.3944
R17742 vdd.n3291 vdd.n642 19.3944
R17743 vdd.n3291 vdd.n640 19.3944
R17744 vdd.n3298 vdd.n640 19.3944
R17745 vdd.n3298 vdd.n3297 19.3944
R17746 vdd.n3297 vdd.n631 19.3944
R17747 vdd.n3311 vdd.n631 19.3944
R17748 vdd.n3312 vdd.n3311 19.3944
R17749 vdd.n3312 vdd.n629 19.3944
R17750 vdd.n3316 vdd.n629 19.3944
R17751 vdd.n3318 vdd.n3316 19.3944
R17752 vdd.n3319 vdd.n3318 19.3944
R17753 vdd.n3319 vdd.n627 19.3944
R17754 vdd.n3323 vdd.n627 19.3944
R17755 vdd.n3325 vdd.n3323 19.3944
R17756 vdd.n3326 vdd.n3325 19.3944
R17757 vdd.n3326 vdd.n625 19.3944
R17758 vdd.n3330 vdd.n625 19.3944
R17759 vdd.n3333 vdd.n3330 19.3944
R17760 vdd.n3334 vdd.n3333 19.3944
R17761 vdd.n3334 vdd.n623 19.3944
R17762 vdd.n3338 vdd.n623 19.3944
R17763 vdd.n3340 vdd.n3338 19.3944
R17764 vdd.n3341 vdd.n3340 19.3944
R17765 vdd.n3341 vdd.n621 19.3944
R17766 vdd.n3345 vdd.n621 19.3944
R17767 vdd.n3347 vdd.n3345 19.3944
R17768 vdd.n3348 vdd.n3347 19.3944
R17769 vdd.n569 vdd.n438 19.3944
R17770 vdd.n575 vdd.n438 19.3944
R17771 vdd.n576 vdd.n575 19.3944
R17772 vdd.n579 vdd.n576 19.3944
R17773 vdd.n579 vdd.n436 19.3944
R17774 vdd.n585 vdd.n436 19.3944
R17775 vdd.n586 vdd.n585 19.3944
R17776 vdd.n589 vdd.n586 19.3944
R17777 vdd.n589 vdd.n434 19.3944
R17778 vdd.n595 vdd.n434 19.3944
R17779 vdd.n596 vdd.n595 19.3944
R17780 vdd.n599 vdd.n596 19.3944
R17781 vdd.n599 vdd.n432 19.3944
R17782 vdd.n605 vdd.n432 19.3944
R17783 vdd.n606 vdd.n605 19.3944
R17784 vdd.n609 vdd.n606 19.3944
R17785 vdd.n609 vdd.n430 19.3944
R17786 vdd.n615 vdd.n430 19.3944
R17787 vdd.n617 vdd.n615 19.3944
R17788 vdd.n618 vdd.n617 19.3944
R17789 vdd.n516 vdd.n515 19.3944
R17790 vdd.n519 vdd.n516 19.3944
R17791 vdd.n519 vdd.n450 19.3944
R17792 vdd.n525 vdd.n450 19.3944
R17793 vdd.n526 vdd.n525 19.3944
R17794 vdd.n529 vdd.n526 19.3944
R17795 vdd.n529 vdd.n448 19.3944
R17796 vdd.n535 vdd.n448 19.3944
R17797 vdd.n536 vdd.n535 19.3944
R17798 vdd.n539 vdd.n536 19.3944
R17799 vdd.n539 vdd.n446 19.3944
R17800 vdd.n545 vdd.n446 19.3944
R17801 vdd.n546 vdd.n545 19.3944
R17802 vdd.n549 vdd.n546 19.3944
R17803 vdd.n549 vdd.n444 19.3944
R17804 vdd.n555 vdd.n444 19.3944
R17805 vdd.n556 vdd.n555 19.3944
R17806 vdd.n559 vdd.n556 19.3944
R17807 vdd.n559 vdd.n442 19.3944
R17808 vdd.n565 vdd.n442 19.3944
R17809 vdd.n466 vdd.n465 19.3944
R17810 vdd.n469 vdd.n466 19.3944
R17811 vdd.n469 vdd.n462 19.3944
R17812 vdd.n475 vdd.n462 19.3944
R17813 vdd.n476 vdd.n475 19.3944
R17814 vdd.n479 vdd.n476 19.3944
R17815 vdd.n479 vdd.n460 19.3944
R17816 vdd.n485 vdd.n460 19.3944
R17817 vdd.n486 vdd.n485 19.3944
R17818 vdd.n489 vdd.n486 19.3944
R17819 vdd.n489 vdd.n458 19.3944
R17820 vdd.n495 vdd.n458 19.3944
R17821 vdd.n496 vdd.n495 19.3944
R17822 vdd.n499 vdd.n496 19.3944
R17823 vdd.n499 vdd.n456 19.3944
R17824 vdd.n505 vdd.n456 19.3944
R17825 vdd.n506 vdd.n505 19.3944
R17826 vdd.n509 vdd.n506 19.3944
R17827 vdd.n3233 vdd.n683 19.3944
R17828 vdd.n3233 vdd.n681 19.3944
R17829 vdd.n3237 vdd.n681 19.3944
R17830 vdd.n3237 vdd.n671 19.3944
R17831 vdd.n3250 vdd.n671 19.3944
R17832 vdd.n3250 vdd.n669 19.3944
R17833 vdd.n3254 vdd.n669 19.3944
R17834 vdd.n3254 vdd.n660 19.3944
R17835 vdd.n3266 vdd.n660 19.3944
R17836 vdd.n3266 vdd.n658 19.3944
R17837 vdd.n3270 vdd.n658 19.3944
R17838 vdd.n3270 vdd.n648 19.3944
R17839 vdd.n3283 vdd.n648 19.3944
R17840 vdd.n3283 vdd.n646 19.3944
R17841 vdd.n3287 vdd.n646 19.3944
R17842 vdd.n3287 vdd.n637 19.3944
R17843 vdd.n3302 vdd.n637 19.3944
R17844 vdd.n3302 vdd.n635 19.3944
R17845 vdd.n3306 vdd.n635 19.3944
R17846 vdd.n3306 vdd.n336 19.3944
R17847 vdd.n3397 vdd.n336 19.3944
R17848 vdd.n3397 vdd.n337 19.3944
R17849 vdd.n3391 vdd.n337 19.3944
R17850 vdd.n3391 vdd.n3390 19.3944
R17851 vdd.n3390 vdd.n3389 19.3944
R17852 vdd.n3389 vdd.n349 19.3944
R17853 vdd.n3383 vdd.n349 19.3944
R17854 vdd.n3383 vdd.n3382 19.3944
R17855 vdd.n3382 vdd.n3381 19.3944
R17856 vdd.n3381 vdd.n359 19.3944
R17857 vdd.n3375 vdd.n359 19.3944
R17858 vdd.n3375 vdd.n3374 19.3944
R17859 vdd.n3374 vdd.n3373 19.3944
R17860 vdd.n3373 vdd.n370 19.3944
R17861 vdd.n3367 vdd.n370 19.3944
R17862 vdd.n3367 vdd.n3366 19.3944
R17863 vdd.n3366 vdd.n3365 19.3944
R17864 vdd.n3365 vdd.n381 19.3944
R17865 vdd.n3359 vdd.n381 19.3944
R17866 vdd.n3359 vdd.n3358 19.3944
R17867 vdd.n3358 vdd.n3357 19.3944
R17868 vdd.n3180 vdd.n747 19.3944
R17869 vdd.n3180 vdd.n3177 19.3944
R17870 vdd.n3177 vdd.n3174 19.3944
R17871 vdd.n3174 vdd.n3173 19.3944
R17872 vdd.n3173 vdd.n3170 19.3944
R17873 vdd.n3170 vdd.n3169 19.3944
R17874 vdd.n3169 vdd.n3166 19.3944
R17875 vdd.n3166 vdd.n3165 19.3944
R17876 vdd.n3165 vdd.n3162 19.3944
R17877 vdd.n3162 vdd.n3161 19.3944
R17878 vdd.n3161 vdd.n3158 19.3944
R17879 vdd.n3158 vdd.n3157 19.3944
R17880 vdd.n3157 vdd.n3154 19.3944
R17881 vdd.n3154 vdd.n3153 19.3944
R17882 vdd.n3153 vdd.n3150 19.3944
R17883 vdd.n3150 vdd.n3149 19.3944
R17884 vdd.n3149 vdd.n3146 19.3944
R17885 vdd.n3146 vdd.n3145 19.3944
R17886 vdd.n3145 vdd.n3142 19.3944
R17887 vdd.n3142 vdd.n3141 19.3944
R17888 vdd.n3220 vdd.n3219 19.3944
R17889 vdd.n3219 vdd.n3218 19.3944
R17890 vdd.n732 vdd.n729 19.3944
R17891 vdd.n3214 vdd.n3213 19.3944
R17892 vdd.n3213 vdd.n3210 19.3944
R17893 vdd.n3210 vdd.n3209 19.3944
R17894 vdd.n3209 vdd.n3206 19.3944
R17895 vdd.n3206 vdd.n3205 19.3944
R17896 vdd.n3205 vdd.n3202 19.3944
R17897 vdd.n3202 vdd.n3201 19.3944
R17898 vdd.n3201 vdd.n3198 19.3944
R17899 vdd.n3198 vdd.n3197 19.3944
R17900 vdd.n3197 vdd.n3194 19.3944
R17901 vdd.n3194 vdd.n3193 19.3944
R17902 vdd.n3193 vdd.n3190 19.3944
R17903 vdd.n3190 vdd.n3189 19.3944
R17904 vdd.n3134 vdd.n767 19.3944
R17905 vdd.n3134 vdd.n3131 19.3944
R17906 vdd.n3131 vdd.n3128 19.3944
R17907 vdd.n3128 vdd.n3127 19.3944
R17908 vdd.n3127 vdd.n3124 19.3944
R17909 vdd.n3124 vdd.n3123 19.3944
R17910 vdd.n3123 vdd.n3120 19.3944
R17911 vdd.n3120 vdd.n3119 19.3944
R17912 vdd.n3119 vdd.n3116 19.3944
R17913 vdd.n3116 vdd.n3115 19.3944
R17914 vdd.n3115 vdd.n3112 19.3944
R17915 vdd.n3112 vdd.n3111 19.3944
R17916 vdd.n3111 vdd.n3108 19.3944
R17917 vdd.n3108 vdd.n3107 19.3944
R17918 vdd.n3107 vdd.n3104 19.3944
R17919 vdd.n3104 vdd.n3103 19.3944
R17920 vdd.n3100 vdd.n3099 19.3944
R17921 vdd.n3096 vdd.n3095 19.3944
R17922 vdd.n1357 vdd.n1353 19.0066
R17923 vdd.n2038 vdd.n1969 19.0066
R17924 vdd.n569 vdd.n566 19.0066
R17925 vdd.n3138 vdd.n767 19.0066
R17926 vdd.n2178 vdd.n2177 16.0975
R17927 vdd.n966 vdd.n965 16.0975
R17928 vdd.n1318 vdd.n1317 16.0975
R17929 vdd.n1356 vdd.n1355 16.0975
R17930 vdd.n1252 vdd.n1251 16.0975
R17931 vdd.n2334 vdd.n2333 16.0975
R17932 vdd.n1971 vdd.n1970 16.0975
R17933 vdd.n1931 vdd.n1930 16.0975
R17934 vdd.n2152 vdd.n2151 16.0975
R17935 vdd.n958 vdd.n957 16.0975
R17936 vdd.n2643 vdd.n2642 16.0975
R17937 vdd.n427 vdd.n426 16.0975
R17938 vdd.n441 vdd.n440 16.0975
R17939 vdd.n453 vdd.n452 16.0975
R17940 vdd.n769 vdd.n768 16.0975
R17941 vdd.n3185 vdd.n3184 16.0975
R17942 vdd.n833 vdd.n832 16.0975
R17943 vdd.n2640 vdd.n2639 16.0975
R17944 vdd.n689 vdd.n688 16.0975
R17945 vdd.n800 vdd.n799 16.0975
R17946 vdd.t26 vdd.n2604 15.4182
R17947 vdd.n2857 vdd.t48 15.4182
R17948 vdd.n2375 vdd.n1049 14.5112
R17949 vdd.n3059 vdd.n692 14.5112
R17950 vdd.n28 vdd.n27 14.4007
R17951 vdd.n328 vdd.n293 13.1884
R17952 vdd.n269 vdd.n234 13.1884
R17953 vdd.n226 vdd.n191 13.1884
R17954 vdd.n167 vdd.n132 13.1884
R17955 vdd.n125 vdd.n90 13.1884
R17956 vdd.n66 vdd.n31 13.1884
R17957 vdd.n1747 vdd.n1712 13.1884
R17958 vdd.n1806 vdd.n1771 13.1884
R17959 vdd.n1645 vdd.n1610 13.1884
R17960 vdd.n1704 vdd.n1669 13.1884
R17961 vdd.n1544 vdd.n1509 13.1884
R17962 vdd.n1603 vdd.n1568 13.1884
R17963 vdd.n1388 vdd.n1253 12.9944
R17964 vdd.n1392 vdd.n1253 12.9944
R17965 vdd.n2077 vdd.n1929 12.9944
R17966 vdd.n2078 vdd.n2077 12.9944
R17967 vdd.n515 vdd.n454 12.9944
R17968 vdd.n509 vdd.n454 12.9944
R17969 vdd.n3186 vdd.n747 12.9944
R17970 vdd.n3189 vdd.n3186 12.9944
R17971 vdd.n329 vdd.n291 12.8005
R17972 vdd.n324 vdd.n295 12.8005
R17973 vdd.n270 vdd.n232 12.8005
R17974 vdd.n265 vdd.n236 12.8005
R17975 vdd.n227 vdd.n189 12.8005
R17976 vdd.n222 vdd.n193 12.8005
R17977 vdd.n168 vdd.n130 12.8005
R17978 vdd.n163 vdd.n134 12.8005
R17979 vdd.n126 vdd.n88 12.8005
R17980 vdd.n121 vdd.n92 12.8005
R17981 vdd.n67 vdd.n29 12.8005
R17982 vdd.n62 vdd.n33 12.8005
R17983 vdd.n1748 vdd.n1710 12.8005
R17984 vdd.n1743 vdd.n1714 12.8005
R17985 vdd.n1807 vdd.n1769 12.8005
R17986 vdd.n1802 vdd.n1773 12.8005
R17987 vdd.n1646 vdd.n1608 12.8005
R17988 vdd.n1641 vdd.n1612 12.8005
R17989 vdd.n1705 vdd.n1667 12.8005
R17990 vdd.n1700 vdd.n1671 12.8005
R17991 vdd.n1545 vdd.n1507 12.8005
R17992 vdd.n1540 vdd.n1511 12.8005
R17993 vdd.n1604 vdd.n1566 12.8005
R17994 vdd.n1599 vdd.n1570 12.8005
R17995 vdd.n323 vdd.n296 12.0247
R17996 vdd.n264 vdd.n237 12.0247
R17997 vdd.n221 vdd.n194 12.0247
R17998 vdd.n162 vdd.n135 12.0247
R17999 vdd.n120 vdd.n93 12.0247
R18000 vdd.n61 vdd.n34 12.0247
R18001 vdd.n1742 vdd.n1715 12.0247
R18002 vdd.n1801 vdd.n1774 12.0247
R18003 vdd.n1640 vdd.n1613 12.0247
R18004 vdd.n1699 vdd.n1672 12.0247
R18005 vdd.n1539 vdd.n1512 12.0247
R18006 vdd.n1598 vdd.n1571 12.0247
R18007 vdd.n1427 vdd.n1183 11.337
R18008 vdd.n1436 vdd.n1183 11.337
R18009 vdd.n1436 vdd.n1435 11.337
R18010 vdd.n1444 vdd.n1177 11.337
R18011 vdd.n1453 vdd.n1452 11.337
R18012 vdd.n1469 vdd.n1161 11.337
R18013 vdd.n1477 vdd.n1154 11.337
R18014 vdd.n1486 vdd.n1485 11.337
R18015 vdd.n1494 vdd.n1143 11.337
R18016 vdd.n1817 vdd.n1132 11.337
R18017 vdd.n1826 vdd.n1126 11.337
R18018 vdd.n1834 vdd.n1120 11.337
R18019 vdd.n1843 vdd.n1842 11.337
R18020 vdd.n1859 vdd.n1104 11.337
R18021 vdd.n1867 vdd.n1097 11.337
R18022 vdd.n1876 vdd.n1875 11.337
R18023 vdd.n1884 vdd.n1080 11.337
R18024 vdd.n1895 vdd.n1080 11.337
R18025 vdd.n1895 vdd.n1894 11.337
R18026 vdd.n3231 vdd.n678 11.337
R18027 vdd.n3239 vdd.n678 11.337
R18028 vdd.n3239 vdd.n679 11.337
R18029 vdd.n3248 vdd.n3247 11.337
R18030 vdd.n3264 vdd.n662 11.337
R18031 vdd.n3272 vdd.n655 11.337
R18032 vdd.n3281 vdd.n3280 11.337
R18033 vdd.n3289 vdd.n644 11.337
R18034 vdd.n3308 vdd.n633 11.337
R18035 vdd.n3395 vdd.n340 11.337
R18036 vdd.n3393 vdd.n344 11.337
R18037 vdd.n3387 vdd.n3386 11.337
R18038 vdd.n3379 vdd.n361 11.337
R18039 vdd.n3378 vdd.n3377 11.337
R18040 vdd.n3371 vdd.n3370 11.337
R18041 vdd.n3369 vdd.n375 11.337
R18042 vdd.n3363 vdd.n3362 11.337
R18043 vdd.n3362 vdd.n3361 11.337
R18044 vdd.n3361 vdd.n386 11.337
R18045 vdd.n320 vdd.n319 11.249
R18046 vdd.n261 vdd.n260 11.249
R18047 vdd.n218 vdd.n217 11.249
R18048 vdd.n159 vdd.n158 11.249
R18049 vdd.n117 vdd.n116 11.249
R18050 vdd.n58 vdd.n57 11.249
R18051 vdd.n1739 vdd.n1738 11.249
R18052 vdd.n1798 vdd.n1797 11.249
R18053 vdd.n1637 vdd.n1636 11.249
R18054 vdd.n1696 vdd.n1695 11.249
R18055 vdd.n1536 vdd.n1535 11.249
R18056 vdd.n1595 vdd.n1594 11.249
R18057 vdd.n1225 vdd.t74 11.2237
R18058 vdd.n3355 vdd.t81 11.2237
R18059 vdd.n2532 vdd.t37 11.1103
R18060 vdd.n2864 vdd.t44 11.1103
R18061 vdd.t157 vdd.n1098 10.7702
R18062 vdd.n3256 vdd.t217 10.7702
R18063 vdd.n305 vdd.n304 10.7238
R18064 vdd.n246 vdd.n245 10.7238
R18065 vdd.n203 vdd.n202 10.7238
R18066 vdd.n144 vdd.n143 10.7238
R18067 vdd.n102 vdd.n101 10.7238
R18068 vdd.n43 vdd.n42 10.7238
R18069 vdd.n1724 vdd.n1723 10.7238
R18070 vdd.n1783 vdd.n1782 10.7238
R18071 vdd.n1622 vdd.n1621 10.7238
R18072 vdd.n1681 vdd.n1680 10.7238
R18073 vdd.n1521 vdd.n1520 10.7238
R18074 vdd.n1580 vdd.n1579 10.7238
R18075 vdd.n2378 vdd.n2377 10.6151
R18076 vdd.n2379 vdd.n2378 10.6151
R18077 vdd.n2379 vdd.n1035 10.6151
R18078 vdd.n2389 vdd.n1035 10.6151
R18079 vdd.n2390 vdd.n2389 10.6151
R18080 vdd.n2391 vdd.n2390 10.6151
R18081 vdd.n2391 vdd.n1022 10.6151
R18082 vdd.n2402 vdd.n1022 10.6151
R18083 vdd.n2403 vdd.n2402 10.6151
R18084 vdd.n2404 vdd.n2403 10.6151
R18085 vdd.n2404 vdd.n1010 10.6151
R18086 vdd.n2414 vdd.n1010 10.6151
R18087 vdd.n2415 vdd.n2414 10.6151
R18088 vdd.n2416 vdd.n2415 10.6151
R18089 vdd.n2416 vdd.n998 10.6151
R18090 vdd.n2426 vdd.n998 10.6151
R18091 vdd.n2427 vdd.n2426 10.6151
R18092 vdd.n2428 vdd.n2427 10.6151
R18093 vdd.n2428 vdd.n987 10.6151
R18094 vdd.n2438 vdd.n987 10.6151
R18095 vdd.n2439 vdd.n2438 10.6151
R18096 vdd.n2440 vdd.n2439 10.6151
R18097 vdd.n2440 vdd.n974 10.6151
R18098 vdd.n2452 vdd.n974 10.6151
R18099 vdd.n2453 vdd.n2452 10.6151
R18100 vdd.n2455 vdd.n2453 10.6151
R18101 vdd.n2455 vdd.n2454 10.6151
R18102 vdd.n2454 vdd.n956 10.6151
R18103 vdd.n2602 vdd.n2601 10.6151
R18104 vdd.n2601 vdd.n2600 10.6151
R18105 vdd.n2600 vdd.n2597 10.6151
R18106 vdd.n2597 vdd.n2596 10.6151
R18107 vdd.n2596 vdd.n2593 10.6151
R18108 vdd.n2593 vdd.n2592 10.6151
R18109 vdd.n2592 vdd.n2589 10.6151
R18110 vdd.n2589 vdd.n2588 10.6151
R18111 vdd.n2588 vdd.n2585 10.6151
R18112 vdd.n2585 vdd.n2584 10.6151
R18113 vdd.n2584 vdd.n2581 10.6151
R18114 vdd.n2581 vdd.n2580 10.6151
R18115 vdd.n2580 vdd.n2577 10.6151
R18116 vdd.n2577 vdd.n2576 10.6151
R18117 vdd.n2576 vdd.n2573 10.6151
R18118 vdd.n2573 vdd.n2572 10.6151
R18119 vdd.n2572 vdd.n2569 10.6151
R18120 vdd.n2569 vdd.n2568 10.6151
R18121 vdd.n2568 vdd.n2565 10.6151
R18122 vdd.n2565 vdd.n2564 10.6151
R18123 vdd.n2564 vdd.n2561 10.6151
R18124 vdd.n2561 vdd.n2560 10.6151
R18125 vdd.n2560 vdd.n2557 10.6151
R18126 vdd.n2557 vdd.n2556 10.6151
R18127 vdd.n2556 vdd.n2553 10.6151
R18128 vdd.n2553 vdd.n2552 10.6151
R18129 vdd.n2552 vdd.n2549 10.6151
R18130 vdd.n2549 vdd.n2548 10.6151
R18131 vdd.n2548 vdd.n2545 10.6151
R18132 vdd.n2545 vdd.n2544 10.6151
R18133 vdd.n2544 vdd.n2541 10.6151
R18134 vdd.n2539 vdd.n2536 10.6151
R18135 vdd.n2536 vdd.n2535 10.6151
R18136 vdd.n2278 vdd.n2277 10.6151
R18137 vdd.n2277 vdd.n2275 10.6151
R18138 vdd.n2275 vdd.n2274 10.6151
R18139 vdd.n2274 vdd.n2272 10.6151
R18140 vdd.n2272 vdd.n2271 10.6151
R18141 vdd.n2271 vdd.n2269 10.6151
R18142 vdd.n2269 vdd.n2268 10.6151
R18143 vdd.n2268 vdd.n2266 10.6151
R18144 vdd.n2266 vdd.n2265 10.6151
R18145 vdd.n2265 vdd.n2263 10.6151
R18146 vdd.n2263 vdd.n2262 10.6151
R18147 vdd.n2262 vdd.n2260 10.6151
R18148 vdd.n2260 vdd.n2259 10.6151
R18149 vdd.n2259 vdd.n2174 10.6151
R18150 vdd.n2174 vdd.n2173 10.6151
R18151 vdd.n2173 vdd.n2171 10.6151
R18152 vdd.n2171 vdd.n2170 10.6151
R18153 vdd.n2170 vdd.n2168 10.6151
R18154 vdd.n2168 vdd.n2167 10.6151
R18155 vdd.n2167 vdd.n2165 10.6151
R18156 vdd.n2165 vdd.n2164 10.6151
R18157 vdd.n2164 vdd.n2162 10.6151
R18158 vdd.n2162 vdd.n2161 10.6151
R18159 vdd.n2161 vdd.n2159 10.6151
R18160 vdd.n2159 vdd.n2158 10.6151
R18161 vdd.n2158 vdd.n2155 10.6151
R18162 vdd.n2155 vdd.n2154 10.6151
R18163 vdd.n2154 vdd.n959 10.6151
R18164 vdd.n2112 vdd.n1047 10.6151
R18165 vdd.n2113 vdd.n2112 10.6151
R18166 vdd.n2114 vdd.n2113 10.6151
R18167 vdd.n2114 vdd.n2108 10.6151
R18168 vdd.n2120 vdd.n2108 10.6151
R18169 vdd.n2121 vdd.n2120 10.6151
R18170 vdd.n2122 vdd.n2121 10.6151
R18171 vdd.n2122 vdd.n2106 10.6151
R18172 vdd.n2128 vdd.n2106 10.6151
R18173 vdd.n2129 vdd.n2128 10.6151
R18174 vdd.n2130 vdd.n2129 10.6151
R18175 vdd.n2130 vdd.n2104 10.6151
R18176 vdd.n2136 vdd.n2104 10.6151
R18177 vdd.n2137 vdd.n2136 10.6151
R18178 vdd.n2138 vdd.n2137 10.6151
R18179 vdd.n2138 vdd.n2102 10.6151
R18180 vdd.n2314 vdd.n2102 10.6151
R18181 vdd.n2314 vdd.n2313 10.6151
R18182 vdd.n2313 vdd.n2143 10.6151
R18183 vdd.n2307 vdd.n2143 10.6151
R18184 vdd.n2307 vdd.n2306 10.6151
R18185 vdd.n2306 vdd.n2305 10.6151
R18186 vdd.n2305 vdd.n2145 10.6151
R18187 vdd.n2299 vdd.n2145 10.6151
R18188 vdd.n2299 vdd.n2298 10.6151
R18189 vdd.n2298 vdd.n2297 10.6151
R18190 vdd.n2297 vdd.n2147 10.6151
R18191 vdd.n2291 vdd.n2147 10.6151
R18192 vdd.n2291 vdd.n2290 10.6151
R18193 vdd.n2290 vdd.n2289 10.6151
R18194 vdd.n2289 vdd.n2149 10.6151
R18195 vdd.n2283 vdd.n2282 10.6151
R18196 vdd.n2282 vdd.n2281 10.6151
R18197 vdd.n2787 vdd.n2786 10.6151
R18198 vdd.n2786 vdd.n2784 10.6151
R18199 vdd.n2784 vdd.n2783 10.6151
R18200 vdd.n2783 vdd.n2641 10.6151
R18201 vdd.n2730 vdd.n2641 10.6151
R18202 vdd.n2731 vdd.n2730 10.6151
R18203 vdd.n2733 vdd.n2731 10.6151
R18204 vdd.n2734 vdd.n2733 10.6151
R18205 vdd.n2736 vdd.n2734 10.6151
R18206 vdd.n2737 vdd.n2736 10.6151
R18207 vdd.n2739 vdd.n2737 10.6151
R18208 vdd.n2740 vdd.n2739 10.6151
R18209 vdd.n2742 vdd.n2740 10.6151
R18210 vdd.n2743 vdd.n2742 10.6151
R18211 vdd.n2758 vdd.n2743 10.6151
R18212 vdd.n2758 vdd.n2757 10.6151
R18213 vdd.n2757 vdd.n2756 10.6151
R18214 vdd.n2756 vdd.n2754 10.6151
R18215 vdd.n2754 vdd.n2753 10.6151
R18216 vdd.n2753 vdd.n2751 10.6151
R18217 vdd.n2751 vdd.n2750 10.6151
R18218 vdd.n2750 vdd.n2748 10.6151
R18219 vdd.n2748 vdd.n2747 10.6151
R18220 vdd.n2747 vdd.n2745 10.6151
R18221 vdd.n2745 vdd.n2744 10.6151
R18222 vdd.n2744 vdd.n836 10.6151
R18223 vdd.n2992 vdd.n836 10.6151
R18224 vdd.n2993 vdd.n2992 10.6151
R18225 vdd.n2854 vdd.n912 10.6151
R18226 vdd.n2854 vdd.n2853 10.6151
R18227 vdd.n2853 vdd.n2852 10.6151
R18228 vdd.n2852 vdd.n2850 10.6151
R18229 vdd.n2850 vdd.n2847 10.6151
R18230 vdd.n2847 vdd.n2846 10.6151
R18231 vdd.n2846 vdd.n2843 10.6151
R18232 vdd.n2843 vdd.n2842 10.6151
R18233 vdd.n2842 vdd.n2839 10.6151
R18234 vdd.n2839 vdd.n2838 10.6151
R18235 vdd.n2838 vdd.n2835 10.6151
R18236 vdd.n2835 vdd.n2834 10.6151
R18237 vdd.n2834 vdd.n2831 10.6151
R18238 vdd.n2831 vdd.n2830 10.6151
R18239 vdd.n2830 vdd.n2827 10.6151
R18240 vdd.n2827 vdd.n2826 10.6151
R18241 vdd.n2826 vdd.n2823 10.6151
R18242 vdd.n2823 vdd.n2822 10.6151
R18243 vdd.n2822 vdd.n2819 10.6151
R18244 vdd.n2819 vdd.n2818 10.6151
R18245 vdd.n2818 vdd.n2815 10.6151
R18246 vdd.n2815 vdd.n2814 10.6151
R18247 vdd.n2814 vdd.n2811 10.6151
R18248 vdd.n2811 vdd.n2810 10.6151
R18249 vdd.n2810 vdd.n2807 10.6151
R18250 vdd.n2807 vdd.n2806 10.6151
R18251 vdd.n2806 vdd.n2803 10.6151
R18252 vdd.n2803 vdd.n2802 10.6151
R18253 vdd.n2802 vdd.n2799 10.6151
R18254 vdd.n2799 vdd.n2798 10.6151
R18255 vdd.n2798 vdd.n2795 10.6151
R18256 vdd.n2793 vdd.n2790 10.6151
R18257 vdd.n2790 vdd.n2789 10.6151
R18258 vdd.n2867 vdd.n2866 10.6151
R18259 vdd.n2868 vdd.n2867 10.6151
R18260 vdd.n2868 vdd.n902 10.6151
R18261 vdd.n2878 vdd.n902 10.6151
R18262 vdd.n2879 vdd.n2878 10.6151
R18263 vdd.n2880 vdd.n2879 10.6151
R18264 vdd.n2880 vdd.n889 10.6151
R18265 vdd.n2890 vdd.n889 10.6151
R18266 vdd.n2891 vdd.n2890 10.6151
R18267 vdd.n2892 vdd.n2891 10.6151
R18268 vdd.n2892 vdd.n878 10.6151
R18269 vdd.n2902 vdd.n878 10.6151
R18270 vdd.n2903 vdd.n2902 10.6151
R18271 vdd.n2904 vdd.n2903 10.6151
R18272 vdd.n2904 vdd.n866 10.6151
R18273 vdd.n2914 vdd.n866 10.6151
R18274 vdd.n2915 vdd.n2914 10.6151
R18275 vdd.n2916 vdd.n2915 10.6151
R18276 vdd.n2916 vdd.n855 10.6151
R18277 vdd.n2928 vdd.n855 10.6151
R18278 vdd.n2929 vdd.n2928 10.6151
R18279 vdd.n2930 vdd.n2929 10.6151
R18280 vdd.n2930 vdd.n841 10.6151
R18281 vdd.n2985 vdd.n841 10.6151
R18282 vdd.n2986 vdd.n2985 10.6151
R18283 vdd.n2987 vdd.n2986 10.6151
R18284 vdd.n2987 vdd.n810 10.6151
R18285 vdd.n3057 vdd.n810 10.6151
R18286 vdd.n3056 vdd.n3055 10.6151
R18287 vdd.n3055 vdd.n811 10.6151
R18288 vdd.n812 vdd.n811 10.6151
R18289 vdd.n3048 vdd.n812 10.6151
R18290 vdd.n3048 vdd.n3047 10.6151
R18291 vdd.n3047 vdd.n3046 10.6151
R18292 vdd.n3046 vdd.n814 10.6151
R18293 vdd.n3041 vdd.n814 10.6151
R18294 vdd.n3041 vdd.n3040 10.6151
R18295 vdd.n3040 vdd.n3039 10.6151
R18296 vdd.n3039 vdd.n817 10.6151
R18297 vdd.n3034 vdd.n817 10.6151
R18298 vdd.n3034 vdd.n3033 10.6151
R18299 vdd.n3033 vdd.n3032 10.6151
R18300 vdd.n3032 vdd.n820 10.6151
R18301 vdd.n3027 vdd.n820 10.6151
R18302 vdd.n3027 vdd.n731 10.6151
R18303 vdd.n3023 vdd.n731 10.6151
R18304 vdd.n3023 vdd.n3022 10.6151
R18305 vdd.n3022 vdd.n3021 10.6151
R18306 vdd.n3021 vdd.n823 10.6151
R18307 vdd.n3016 vdd.n823 10.6151
R18308 vdd.n3016 vdd.n3015 10.6151
R18309 vdd.n3015 vdd.n3014 10.6151
R18310 vdd.n3014 vdd.n826 10.6151
R18311 vdd.n3009 vdd.n826 10.6151
R18312 vdd.n3009 vdd.n3008 10.6151
R18313 vdd.n3008 vdd.n3007 10.6151
R18314 vdd.n3007 vdd.n829 10.6151
R18315 vdd.n3002 vdd.n829 10.6151
R18316 vdd.n3002 vdd.n3001 10.6151
R18317 vdd.n2999 vdd.n834 10.6151
R18318 vdd.n2994 vdd.n834 10.6151
R18319 vdd.n2975 vdd.n2936 10.6151
R18320 vdd.n2970 vdd.n2936 10.6151
R18321 vdd.n2970 vdd.n2969 10.6151
R18322 vdd.n2969 vdd.n2968 10.6151
R18323 vdd.n2968 vdd.n2938 10.6151
R18324 vdd.n2963 vdd.n2938 10.6151
R18325 vdd.n2963 vdd.n2962 10.6151
R18326 vdd.n2962 vdd.n2961 10.6151
R18327 vdd.n2961 vdd.n2941 10.6151
R18328 vdd.n2956 vdd.n2941 10.6151
R18329 vdd.n2956 vdd.n2955 10.6151
R18330 vdd.n2955 vdd.n2954 10.6151
R18331 vdd.n2954 vdd.n2944 10.6151
R18332 vdd.n2949 vdd.n2944 10.6151
R18333 vdd.n2949 vdd.n2948 10.6151
R18334 vdd.n2948 vdd.n785 10.6151
R18335 vdd.n3092 vdd.n785 10.6151
R18336 vdd.n3092 vdd.n786 10.6151
R18337 vdd.n788 vdd.n786 10.6151
R18338 vdd.n3085 vdd.n788 10.6151
R18339 vdd.n3085 vdd.n3084 10.6151
R18340 vdd.n3084 vdd.n3083 10.6151
R18341 vdd.n3083 vdd.n790 10.6151
R18342 vdd.n3078 vdd.n790 10.6151
R18343 vdd.n3078 vdd.n3077 10.6151
R18344 vdd.n3077 vdd.n3076 10.6151
R18345 vdd.n3076 vdd.n793 10.6151
R18346 vdd.n3071 vdd.n793 10.6151
R18347 vdd.n3071 vdd.n3070 10.6151
R18348 vdd.n3070 vdd.n3069 10.6151
R18349 vdd.n3069 vdd.n796 10.6151
R18350 vdd.n3064 vdd.n3063 10.6151
R18351 vdd.n3063 vdd.n3062 10.6151
R18352 vdd.n2710 vdd.n2708 10.6151
R18353 vdd.n2711 vdd.n2710 10.6151
R18354 vdd.n2779 vdd.n2711 10.6151
R18355 vdd.n2779 vdd.n2778 10.6151
R18356 vdd.n2778 vdd.n2777 10.6151
R18357 vdd.n2777 vdd.n2775 10.6151
R18358 vdd.n2775 vdd.n2774 10.6151
R18359 vdd.n2774 vdd.n2772 10.6151
R18360 vdd.n2772 vdd.n2771 10.6151
R18361 vdd.n2771 vdd.n2769 10.6151
R18362 vdd.n2769 vdd.n2768 10.6151
R18363 vdd.n2768 vdd.n2766 10.6151
R18364 vdd.n2766 vdd.n2765 10.6151
R18365 vdd.n2765 vdd.n2763 10.6151
R18366 vdd.n2763 vdd.n2762 10.6151
R18367 vdd.n2762 vdd.n2728 10.6151
R18368 vdd.n2728 vdd.n2727 10.6151
R18369 vdd.n2727 vdd.n2725 10.6151
R18370 vdd.n2725 vdd.n2724 10.6151
R18371 vdd.n2724 vdd.n2722 10.6151
R18372 vdd.n2722 vdd.n2721 10.6151
R18373 vdd.n2721 vdd.n2719 10.6151
R18374 vdd.n2719 vdd.n2718 10.6151
R18375 vdd.n2718 vdd.n2716 10.6151
R18376 vdd.n2716 vdd.n2715 10.6151
R18377 vdd.n2715 vdd.n2713 10.6151
R18378 vdd.n2713 vdd.n2712 10.6151
R18379 vdd.n2712 vdd.n802 10.6151
R18380 vdd.n2861 vdd.n2860 10.6151
R18381 vdd.n2860 vdd.n917 10.6151
R18382 vdd.n2645 vdd.n917 10.6151
R18383 vdd.n2648 vdd.n2645 10.6151
R18384 vdd.n2649 vdd.n2648 10.6151
R18385 vdd.n2652 vdd.n2649 10.6151
R18386 vdd.n2653 vdd.n2652 10.6151
R18387 vdd.n2656 vdd.n2653 10.6151
R18388 vdd.n2657 vdd.n2656 10.6151
R18389 vdd.n2660 vdd.n2657 10.6151
R18390 vdd.n2661 vdd.n2660 10.6151
R18391 vdd.n2664 vdd.n2661 10.6151
R18392 vdd.n2665 vdd.n2664 10.6151
R18393 vdd.n2668 vdd.n2665 10.6151
R18394 vdd.n2669 vdd.n2668 10.6151
R18395 vdd.n2672 vdd.n2669 10.6151
R18396 vdd.n2673 vdd.n2672 10.6151
R18397 vdd.n2676 vdd.n2673 10.6151
R18398 vdd.n2677 vdd.n2676 10.6151
R18399 vdd.n2680 vdd.n2677 10.6151
R18400 vdd.n2681 vdd.n2680 10.6151
R18401 vdd.n2684 vdd.n2681 10.6151
R18402 vdd.n2685 vdd.n2684 10.6151
R18403 vdd.n2688 vdd.n2685 10.6151
R18404 vdd.n2689 vdd.n2688 10.6151
R18405 vdd.n2692 vdd.n2689 10.6151
R18406 vdd.n2693 vdd.n2692 10.6151
R18407 vdd.n2696 vdd.n2693 10.6151
R18408 vdd.n2697 vdd.n2696 10.6151
R18409 vdd.n2700 vdd.n2697 10.6151
R18410 vdd.n2701 vdd.n2700 10.6151
R18411 vdd.n2706 vdd.n2704 10.6151
R18412 vdd.n2707 vdd.n2706 10.6151
R18413 vdd.n2862 vdd.n907 10.6151
R18414 vdd.n2872 vdd.n907 10.6151
R18415 vdd.n2873 vdd.n2872 10.6151
R18416 vdd.n2874 vdd.n2873 10.6151
R18417 vdd.n2874 vdd.n895 10.6151
R18418 vdd.n2884 vdd.n895 10.6151
R18419 vdd.n2885 vdd.n2884 10.6151
R18420 vdd.n2886 vdd.n2885 10.6151
R18421 vdd.n2886 vdd.n884 10.6151
R18422 vdd.n2896 vdd.n884 10.6151
R18423 vdd.n2897 vdd.n2896 10.6151
R18424 vdd.n2898 vdd.n2897 10.6151
R18425 vdd.n2898 vdd.n872 10.6151
R18426 vdd.n2908 vdd.n872 10.6151
R18427 vdd.n2909 vdd.n2908 10.6151
R18428 vdd.n2910 vdd.n2909 10.6151
R18429 vdd.n2910 vdd.n861 10.6151
R18430 vdd.n2920 vdd.n861 10.6151
R18431 vdd.n2921 vdd.n2920 10.6151
R18432 vdd.n2924 vdd.n2921 10.6151
R18433 vdd.n2934 vdd.n849 10.6151
R18434 vdd.n2935 vdd.n2934 10.6151
R18435 vdd.n2981 vdd.n2935 10.6151
R18436 vdd.n2981 vdd.n2980 10.6151
R18437 vdd.n2980 vdd.n2979 10.6151
R18438 vdd.n2979 vdd.n2978 10.6151
R18439 vdd.n2978 vdd.n2976 10.6151
R18440 vdd.n2373 vdd.n1041 10.6151
R18441 vdd.n2383 vdd.n1041 10.6151
R18442 vdd.n2384 vdd.n2383 10.6151
R18443 vdd.n2385 vdd.n2384 10.6151
R18444 vdd.n2385 vdd.n1028 10.6151
R18445 vdd.n2395 vdd.n1028 10.6151
R18446 vdd.n2396 vdd.n2395 10.6151
R18447 vdd.n2398 vdd.n1016 10.6151
R18448 vdd.n2408 vdd.n1016 10.6151
R18449 vdd.n2409 vdd.n2408 10.6151
R18450 vdd.n2410 vdd.n2409 10.6151
R18451 vdd.n2410 vdd.n1004 10.6151
R18452 vdd.n2420 vdd.n1004 10.6151
R18453 vdd.n2421 vdd.n2420 10.6151
R18454 vdd.n2422 vdd.n2421 10.6151
R18455 vdd.n2422 vdd.n993 10.6151
R18456 vdd.n2432 vdd.n993 10.6151
R18457 vdd.n2433 vdd.n2432 10.6151
R18458 vdd.n2434 vdd.n2433 10.6151
R18459 vdd.n2434 vdd.n981 10.6151
R18460 vdd.n2444 vdd.n981 10.6151
R18461 vdd.n2445 vdd.n2444 10.6151
R18462 vdd.n2448 vdd.n2445 10.6151
R18463 vdd.n2448 vdd.n2447 10.6151
R18464 vdd.n2447 vdd.n2446 10.6151
R18465 vdd.n2446 vdd.n964 10.6151
R18466 vdd.n2530 vdd.n964 10.6151
R18467 vdd.n2529 vdd.n2528 10.6151
R18468 vdd.n2528 vdd.n2525 10.6151
R18469 vdd.n2525 vdd.n2524 10.6151
R18470 vdd.n2524 vdd.n2521 10.6151
R18471 vdd.n2521 vdd.n2520 10.6151
R18472 vdd.n2520 vdd.n2517 10.6151
R18473 vdd.n2517 vdd.n2516 10.6151
R18474 vdd.n2516 vdd.n2513 10.6151
R18475 vdd.n2513 vdd.n2512 10.6151
R18476 vdd.n2512 vdd.n2509 10.6151
R18477 vdd.n2509 vdd.n2508 10.6151
R18478 vdd.n2508 vdd.n2505 10.6151
R18479 vdd.n2505 vdd.n2504 10.6151
R18480 vdd.n2504 vdd.n2501 10.6151
R18481 vdd.n2501 vdd.n2500 10.6151
R18482 vdd.n2500 vdd.n2497 10.6151
R18483 vdd.n2497 vdd.n2496 10.6151
R18484 vdd.n2496 vdd.n2493 10.6151
R18485 vdd.n2493 vdd.n2492 10.6151
R18486 vdd.n2492 vdd.n2489 10.6151
R18487 vdd.n2489 vdd.n2488 10.6151
R18488 vdd.n2488 vdd.n2485 10.6151
R18489 vdd.n2485 vdd.n2484 10.6151
R18490 vdd.n2484 vdd.n2481 10.6151
R18491 vdd.n2481 vdd.n2480 10.6151
R18492 vdd.n2480 vdd.n2477 10.6151
R18493 vdd.n2477 vdd.n2476 10.6151
R18494 vdd.n2476 vdd.n2473 10.6151
R18495 vdd.n2473 vdd.n2472 10.6151
R18496 vdd.n2472 vdd.n2469 10.6151
R18497 vdd.n2469 vdd.n2468 10.6151
R18498 vdd.n2465 vdd.n2464 10.6151
R18499 vdd.n2464 vdd.n2462 10.6151
R18500 vdd.n2221 vdd.n2219 10.6151
R18501 vdd.n2222 vdd.n2221 10.6151
R18502 vdd.n2224 vdd.n2222 10.6151
R18503 vdd.n2225 vdd.n2224 10.6151
R18504 vdd.n2227 vdd.n2225 10.6151
R18505 vdd.n2228 vdd.n2227 10.6151
R18506 vdd.n2230 vdd.n2228 10.6151
R18507 vdd.n2231 vdd.n2230 10.6151
R18508 vdd.n2233 vdd.n2231 10.6151
R18509 vdd.n2234 vdd.n2233 10.6151
R18510 vdd.n2236 vdd.n2234 10.6151
R18511 vdd.n2237 vdd.n2236 10.6151
R18512 vdd.n2255 vdd.n2237 10.6151
R18513 vdd.n2255 vdd.n2254 10.6151
R18514 vdd.n2254 vdd.n2253 10.6151
R18515 vdd.n2253 vdd.n2251 10.6151
R18516 vdd.n2251 vdd.n2250 10.6151
R18517 vdd.n2250 vdd.n2248 10.6151
R18518 vdd.n2248 vdd.n2247 10.6151
R18519 vdd.n2247 vdd.n2245 10.6151
R18520 vdd.n2245 vdd.n2244 10.6151
R18521 vdd.n2244 vdd.n2242 10.6151
R18522 vdd.n2242 vdd.n2241 10.6151
R18523 vdd.n2241 vdd.n2239 10.6151
R18524 vdd.n2239 vdd.n2238 10.6151
R18525 vdd.n2238 vdd.n968 10.6151
R18526 vdd.n2460 vdd.n968 10.6151
R18527 vdd.n2461 vdd.n2460 10.6151
R18528 vdd.n2372 vdd.n2371 10.6151
R18529 vdd.n2371 vdd.n1053 10.6151
R18530 vdd.n2365 vdd.n1053 10.6151
R18531 vdd.n2365 vdd.n2364 10.6151
R18532 vdd.n2364 vdd.n2363 10.6151
R18533 vdd.n2363 vdd.n1055 10.6151
R18534 vdd.n2357 vdd.n1055 10.6151
R18535 vdd.n2357 vdd.n2356 10.6151
R18536 vdd.n2356 vdd.n2355 10.6151
R18537 vdd.n2355 vdd.n1057 10.6151
R18538 vdd.n2349 vdd.n1057 10.6151
R18539 vdd.n2349 vdd.n2348 10.6151
R18540 vdd.n2348 vdd.n2347 10.6151
R18541 vdd.n2347 vdd.n1059 10.6151
R18542 vdd.n2341 vdd.n1059 10.6151
R18543 vdd.n2341 vdd.n2340 10.6151
R18544 vdd.n2340 vdd.n2339 10.6151
R18545 vdd.n2339 vdd.n1063 10.6151
R18546 vdd.n2187 vdd.n1063 10.6151
R18547 vdd.n2188 vdd.n2187 10.6151
R18548 vdd.n2188 vdd.n2183 10.6151
R18549 vdd.n2194 vdd.n2183 10.6151
R18550 vdd.n2195 vdd.n2194 10.6151
R18551 vdd.n2196 vdd.n2195 10.6151
R18552 vdd.n2196 vdd.n2181 10.6151
R18553 vdd.n2202 vdd.n2181 10.6151
R18554 vdd.n2203 vdd.n2202 10.6151
R18555 vdd.n2204 vdd.n2203 10.6151
R18556 vdd.n2204 vdd.n2179 10.6151
R18557 vdd.n2210 vdd.n2179 10.6151
R18558 vdd.n2211 vdd.n2210 10.6151
R18559 vdd.n2213 vdd.n2175 10.6151
R18560 vdd.n2218 vdd.n2175 10.6151
R18561 vdd.n1851 vdd.t146 10.5435
R18562 vdd.n656 vdd.t253 10.5435
R18563 vdd.n316 vdd.n298 10.4732
R18564 vdd.n257 vdd.n239 10.4732
R18565 vdd.n214 vdd.n196 10.4732
R18566 vdd.n155 vdd.n137 10.4732
R18567 vdd.n113 vdd.n95 10.4732
R18568 vdd.n54 vdd.n36 10.4732
R18569 vdd.n1735 vdd.n1717 10.4732
R18570 vdd.n1794 vdd.n1776 10.4732
R18571 vdd.n1633 vdd.n1615 10.4732
R18572 vdd.n1692 vdd.n1674 10.4732
R18573 vdd.n1532 vdd.n1514 10.4732
R18574 vdd.n1591 vdd.n1573 10.4732
R18575 vdd.t234 vdd.n1825 10.3167
R18576 vdd.n3300 vdd.t195 10.3167
R18577 vdd.n1502 vdd.t165 10.09
R18578 vdd.n3394 vdd.t163 10.09
R18579 vdd.t229 vdd.n1155 9.86327
R18580 vdd.n3385 vdd.t161 9.86327
R18581 vdd.n315 vdd.n300 9.69747
R18582 vdd.n256 vdd.n241 9.69747
R18583 vdd.n213 vdd.n198 9.69747
R18584 vdd.n154 vdd.n139 9.69747
R18585 vdd.n112 vdd.n97 9.69747
R18586 vdd.n53 vdd.n38 9.69747
R18587 vdd.n1734 vdd.n1719 9.69747
R18588 vdd.n1793 vdd.n1778 9.69747
R18589 vdd.n1632 vdd.n1617 9.69747
R18590 vdd.n1691 vdd.n1676 9.69747
R18591 vdd.n1531 vdd.n1516 9.69747
R18592 vdd.n1590 vdd.n1575 9.69747
R18593 vdd.n2315 vdd.n2314 9.67831
R18594 vdd.n3216 vdd.n731 9.67831
R18595 vdd.n3093 vdd.n3092 9.67831
R18596 vdd.n2339 vdd.n2338 9.67831
R18597 vdd.n1461 vdd.t180 9.63654
R18598 vdd.n3331 vdd.t159 9.63654
R18599 vdd.n331 vdd.n330 9.45567
R18600 vdd.n272 vdd.n271 9.45567
R18601 vdd.n229 vdd.n228 9.45567
R18602 vdd.n170 vdd.n169 9.45567
R18603 vdd.n128 vdd.n127 9.45567
R18604 vdd.n69 vdd.n68 9.45567
R18605 vdd.n1750 vdd.n1749 9.45567
R18606 vdd.n1809 vdd.n1808 9.45567
R18607 vdd.n1648 vdd.n1647 9.45567
R18608 vdd.n1707 vdd.n1706 9.45567
R18609 vdd.n1547 vdd.n1546 9.45567
R18610 vdd.n1606 vdd.n1605 9.45567
R18611 vdd.n1435 vdd.t148 9.40981
R18612 vdd.n3363 vdd.t202 9.40981
R18613 vdd.n2075 vdd.n1929 9.3005
R18614 vdd.n2074 vdd.n2073 9.3005
R18615 vdd.n1935 vdd.n1934 9.3005
R18616 vdd.n2068 vdd.n1939 9.3005
R18617 vdd.n2067 vdd.n1940 9.3005
R18618 vdd.n2066 vdd.n1941 9.3005
R18619 vdd.n1945 vdd.n1942 9.3005
R18620 vdd.n2061 vdd.n1946 9.3005
R18621 vdd.n2060 vdd.n1947 9.3005
R18622 vdd.n2059 vdd.n1948 9.3005
R18623 vdd.n1952 vdd.n1949 9.3005
R18624 vdd.n2054 vdd.n1953 9.3005
R18625 vdd.n2053 vdd.n1954 9.3005
R18626 vdd.n2052 vdd.n1955 9.3005
R18627 vdd.n1959 vdd.n1956 9.3005
R18628 vdd.n2047 vdd.n1960 9.3005
R18629 vdd.n2046 vdd.n1961 9.3005
R18630 vdd.n2045 vdd.n1962 9.3005
R18631 vdd.n1966 vdd.n1963 9.3005
R18632 vdd.n2040 vdd.n1967 9.3005
R18633 vdd.n2039 vdd.n1968 9.3005
R18634 vdd.n2038 vdd.n2037 9.3005
R18635 vdd.n2036 vdd.n1969 9.3005
R18636 vdd.n2035 vdd.n2034 9.3005
R18637 vdd.n1975 vdd.n1974 9.3005
R18638 vdd.n2029 vdd.n1979 9.3005
R18639 vdd.n2028 vdd.n1980 9.3005
R18640 vdd.n2027 vdd.n1981 9.3005
R18641 vdd.n1985 vdd.n1982 9.3005
R18642 vdd.n2022 vdd.n1986 9.3005
R18643 vdd.n2021 vdd.n1987 9.3005
R18644 vdd.n2020 vdd.n1988 9.3005
R18645 vdd.n1992 vdd.n1989 9.3005
R18646 vdd.n2015 vdd.n1993 9.3005
R18647 vdd.n2014 vdd.n1994 9.3005
R18648 vdd.n2013 vdd.n1995 9.3005
R18649 vdd.n1997 vdd.n1996 9.3005
R18650 vdd.n2008 vdd.n1064 9.3005
R18651 vdd.n2077 vdd.n2076 9.3005
R18652 vdd.n2101 vdd.n2100 9.3005
R18653 vdd.n1907 vdd.n1906 9.3005
R18654 vdd.n1912 vdd.n1910 9.3005
R18655 vdd.n2093 vdd.n1913 9.3005
R18656 vdd.n2092 vdd.n1914 9.3005
R18657 vdd.n2091 vdd.n1915 9.3005
R18658 vdd.n1919 vdd.n1916 9.3005
R18659 vdd.n2086 vdd.n1920 9.3005
R18660 vdd.n2085 vdd.n1921 9.3005
R18661 vdd.n2084 vdd.n1922 9.3005
R18662 vdd.n1926 vdd.n1923 9.3005
R18663 vdd.n2079 vdd.n1927 9.3005
R18664 vdd.n2078 vdd.n1928 9.3005
R18665 vdd.n2323 vdd.n1900 9.3005
R18666 vdd.n2325 vdd.n2324 9.3005
R18667 vdd.n1815 vdd.n1814 9.3005
R18668 vdd.n1124 vdd.n1123 9.3005
R18669 vdd.n1829 vdd.n1828 9.3005
R18670 vdd.n1830 vdd.n1122 9.3005
R18671 vdd.n1832 vdd.n1831 9.3005
R18672 vdd.n1113 vdd.n1112 9.3005
R18673 vdd.n1846 vdd.n1845 9.3005
R18674 vdd.n1847 vdd.n1111 9.3005
R18675 vdd.n1849 vdd.n1848 9.3005
R18676 vdd.n1102 vdd.n1101 9.3005
R18677 vdd.n1862 vdd.n1861 9.3005
R18678 vdd.n1863 vdd.n1100 9.3005
R18679 vdd.n1865 vdd.n1864 9.3005
R18680 vdd.n1090 vdd.n1089 9.3005
R18681 vdd.n1879 vdd.n1878 9.3005
R18682 vdd.n1880 vdd.n1088 9.3005
R18683 vdd.n1882 vdd.n1881 9.3005
R18684 vdd.n1078 vdd.n1077 9.3005
R18685 vdd.n1898 vdd.n1897 9.3005
R18686 vdd.n1899 vdd.n1076 9.3005
R18687 vdd.n2327 vdd.n2326 9.3005
R18688 vdd.n307 vdd.n306 9.3005
R18689 vdd.n302 vdd.n301 9.3005
R18690 vdd.n313 vdd.n312 9.3005
R18691 vdd.n315 vdd.n314 9.3005
R18692 vdd.n298 vdd.n297 9.3005
R18693 vdd.n321 vdd.n320 9.3005
R18694 vdd.n323 vdd.n322 9.3005
R18695 vdd.n295 vdd.n292 9.3005
R18696 vdd.n330 vdd.n329 9.3005
R18697 vdd.n248 vdd.n247 9.3005
R18698 vdd.n243 vdd.n242 9.3005
R18699 vdd.n254 vdd.n253 9.3005
R18700 vdd.n256 vdd.n255 9.3005
R18701 vdd.n239 vdd.n238 9.3005
R18702 vdd.n262 vdd.n261 9.3005
R18703 vdd.n264 vdd.n263 9.3005
R18704 vdd.n236 vdd.n233 9.3005
R18705 vdd.n271 vdd.n270 9.3005
R18706 vdd.n205 vdd.n204 9.3005
R18707 vdd.n200 vdd.n199 9.3005
R18708 vdd.n211 vdd.n210 9.3005
R18709 vdd.n213 vdd.n212 9.3005
R18710 vdd.n196 vdd.n195 9.3005
R18711 vdd.n219 vdd.n218 9.3005
R18712 vdd.n221 vdd.n220 9.3005
R18713 vdd.n193 vdd.n190 9.3005
R18714 vdd.n228 vdd.n227 9.3005
R18715 vdd.n146 vdd.n145 9.3005
R18716 vdd.n141 vdd.n140 9.3005
R18717 vdd.n152 vdd.n151 9.3005
R18718 vdd.n154 vdd.n153 9.3005
R18719 vdd.n137 vdd.n136 9.3005
R18720 vdd.n160 vdd.n159 9.3005
R18721 vdd.n162 vdd.n161 9.3005
R18722 vdd.n134 vdd.n131 9.3005
R18723 vdd.n169 vdd.n168 9.3005
R18724 vdd.n104 vdd.n103 9.3005
R18725 vdd.n99 vdd.n98 9.3005
R18726 vdd.n110 vdd.n109 9.3005
R18727 vdd.n112 vdd.n111 9.3005
R18728 vdd.n95 vdd.n94 9.3005
R18729 vdd.n118 vdd.n117 9.3005
R18730 vdd.n120 vdd.n119 9.3005
R18731 vdd.n92 vdd.n89 9.3005
R18732 vdd.n127 vdd.n126 9.3005
R18733 vdd.n45 vdd.n44 9.3005
R18734 vdd.n40 vdd.n39 9.3005
R18735 vdd.n51 vdd.n50 9.3005
R18736 vdd.n53 vdd.n52 9.3005
R18737 vdd.n36 vdd.n35 9.3005
R18738 vdd.n59 vdd.n58 9.3005
R18739 vdd.n61 vdd.n60 9.3005
R18740 vdd.n33 vdd.n30 9.3005
R18741 vdd.n68 vdd.n67 9.3005
R18742 vdd.n3138 vdd.n3137 9.3005
R18743 vdd.n3141 vdd.n766 9.3005
R18744 vdd.n3142 vdd.n765 9.3005
R18745 vdd.n3145 vdd.n764 9.3005
R18746 vdd.n3146 vdd.n763 9.3005
R18747 vdd.n3149 vdd.n762 9.3005
R18748 vdd.n3150 vdd.n761 9.3005
R18749 vdd.n3153 vdd.n760 9.3005
R18750 vdd.n3154 vdd.n759 9.3005
R18751 vdd.n3157 vdd.n758 9.3005
R18752 vdd.n3158 vdd.n757 9.3005
R18753 vdd.n3161 vdd.n756 9.3005
R18754 vdd.n3162 vdd.n755 9.3005
R18755 vdd.n3165 vdd.n754 9.3005
R18756 vdd.n3166 vdd.n753 9.3005
R18757 vdd.n3169 vdd.n752 9.3005
R18758 vdd.n3170 vdd.n751 9.3005
R18759 vdd.n3173 vdd.n750 9.3005
R18760 vdd.n3174 vdd.n749 9.3005
R18761 vdd.n3177 vdd.n748 9.3005
R18762 vdd.n3181 vdd.n3180 9.3005
R18763 vdd.n3182 vdd.n747 9.3005
R18764 vdd.n3186 vdd.n3183 9.3005
R18765 vdd.n3189 vdd.n746 9.3005
R18766 vdd.n3190 vdd.n745 9.3005
R18767 vdd.n3193 vdd.n744 9.3005
R18768 vdd.n3194 vdd.n743 9.3005
R18769 vdd.n3197 vdd.n742 9.3005
R18770 vdd.n3198 vdd.n741 9.3005
R18771 vdd.n3201 vdd.n740 9.3005
R18772 vdd.n3202 vdd.n739 9.3005
R18773 vdd.n3205 vdd.n738 9.3005
R18774 vdd.n3206 vdd.n737 9.3005
R18775 vdd.n3209 vdd.n736 9.3005
R18776 vdd.n3210 vdd.n735 9.3005
R18777 vdd.n3213 vdd.n730 9.3005
R18778 vdd.n3219 vdd.n727 9.3005
R18779 vdd.n3220 vdd.n726 9.3005
R18780 vdd.n3234 vdd.n3233 9.3005
R18781 vdd.n3235 vdd.n681 9.3005
R18782 vdd.n3237 vdd.n3236 9.3005
R18783 vdd.n671 vdd.n670 9.3005
R18784 vdd.n3251 vdd.n3250 9.3005
R18785 vdd.n3252 vdd.n669 9.3005
R18786 vdd.n3254 vdd.n3253 9.3005
R18787 vdd.n660 vdd.n659 9.3005
R18788 vdd.n3267 vdd.n3266 9.3005
R18789 vdd.n3268 vdd.n658 9.3005
R18790 vdd.n3270 vdd.n3269 9.3005
R18791 vdd.n648 vdd.n647 9.3005
R18792 vdd.n3284 vdd.n3283 9.3005
R18793 vdd.n3285 vdd.n646 9.3005
R18794 vdd.n3287 vdd.n3286 9.3005
R18795 vdd.n637 vdd.n636 9.3005
R18796 vdd.n3303 vdd.n3302 9.3005
R18797 vdd.n3304 vdd.n635 9.3005
R18798 vdd.n3306 vdd.n3305 9.3005
R18799 vdd.n336 vdd.n334 9.3005
R18800 vdd.n683 vdd.n682 9.3005
R18801 vdd.n3398 vdd.n3397 9.3005
R18802 vdd.n337 vdd.n335 9.3005
R18803 vdd.n3391 vdd.n346 9.3005
R18804 vdd.n3390 vdd.n347 9.3005
R18805 vdd.n3389 vdd.n348 9.3005
R18806 vdd.n355 vdd.n349 9.3005
R18807 vdd.n3383 vdd.n356 9.3005
R18808 vdd.n3382 vdd.n357 9.3005
R18809 vdd.n3381 vdd.n358 9.3005
R18810 vdd.n366 vdd.n359 9.3005
R18811 vdd.n3375 vdd.n367 9.3005
R18812 vdd.n3374 vdd.n368 9.3005
R18813 vdd.n3373 vdd.n369 9.3005
R18814 vdd.n377 vdd.n370 9.3005
R18815 vdd.n3367 vdd.n378 9.3005
R18816 vdd.n3366 vdd.n379 9.3005
R18817 vdd.n3365 vdd.n380 9.3005
R18818 vdd.n388 vdd.n381 9.3005
R18819 vdd.n3359 vdd.n389 9.3005
R18820 vdd.n3358 vdd.n390 9.3005
R18821 vdd.n3357 vdd.n391 9.3005
R18822 vdd.n466 vdd.n463 9.3005
R18823 vdd.n470 vdd.n469 9.3005
R18824 vdd.n471 vdd.n462 9.3005
R18825 vdd.n475 vdd.n472 9.3005
R18826 vdd.n476 vdd.n461 9.3005
R18827 vdd.n480 vdd.n479 9.3005
R18828 vdd.n481 vdd.n460 9.3005
R18829 vdd.n485 vdd.n482 9.3005
R18830 vdd.n486 vdd.n459 9.3005
R18831 vdd.n490 vdd.n489 9.3005
R18832 vdd.n491 vdd.n458 9.3005
R18833 vdd.n495 vdd.n492 9.3005
R18834 vdd.n496 vdd.n457 9.3005
R18835 vdd.n500 vdd.n499 9.3005
R18836 vdd.n501 vdd.n456 9.3005
R18837 vdd.n505 vdd.n502 9.3005
R18838 vdd.n506 vdd.n455 9.3005
R18839 vdd.n510 vdd.n509 9.3005
R18840 vdd.n511 vdd.n454 9.3005
R18841 vdd.n515 vdd.n512 9.3005
R18842 vdd.n516 vdd.n451 9.3005
R18843 vdd.n520 vdd.n519 9.3005
R18844 vdd.n521 vdd.n450 9.3005
R18845 vdd.n525 vdd.n522 9.3005
R18846 vdd.n526 vdd.n449 9.3005
R18847 vdd.n530 vdd.n529 9.3005
R18848 vdd.n531 vdd.n448 9.3005
R18849 vdd.n535 vdd.n532 9.3005
R18850 vdd.n536 vdd.n447 9.3005
R18851 vdd.n540 vdd.n539 9.3005
R18852 vdd.n541 vdd.n446 9.3005
R18853 vdd.n545 vdd.n542 9.3005
R18854 vdd.n546 vdd.n445 9.3005
R18855 vdd.n550 vdd.n549 9.3005
R18856 vdd.n551 vdd.n444 9.3005
R18857 vdd.n555 vdd.n552 9.3005
R18858 vdd.n556 vdd.n443 9.3005
R18859 vdd.n560 vdd.n559 9.3005
R18860 vdd.n561 vdd.n442 9.3005
R18861 vdd.n565 vdd.n562 9.3005
R18862 vdd.n566 vdd.n439 9.3005
R18863 vdd.n570 vdd.n569 9.3005
R18864 vdd.n571 vdd.n438 9.3005
R18865 vdd.n575 vdd.n572 9.3005
R18866 vdd.n576 vdd.n437 9.3005
R18867 vdd.n580 vdd.n579 9.3005
R18868 vdd.n581 vdd.n436 9.3005
R18869 vdd.n585 vdd.n582 9.3005
R18870 vdd.n586 vdd.n435 9.3005
R18871 vdd.n590 vdd.n589 9.3005
R18872 vdd.n591 vdd.n434 9.3005
R18873 vdd.n595 vdd.n592 9.3005
R18874 vdd.n596 vdd.n433 9.3005
R18875 vdd.n600 vdd.n599 9.3005
R18876 vdd.n601 vdd.n432 9.3005
R18877 vdd.n605 vdd.n602 9.3005
R18878 vdd.n606 vdd.n431 9.3005
R18879 vdd.n610 vdd.n609 9.3005
R18880 vdd.n611 vdd.n430 9.3005
R18881 vdd.n615 vdd.n612 9.3005
R18882 vdd.n617 vdd.n429 9.3005
R18883 vdd.n619 vdd.n618 9.3005
R18884 vdd.n3351 vdd.n3350 9.3005
R18885 vdd.n465 vdd.n464 9.3005
R18886 vdd.n3229 vdd.n3228 9.3005
R18887 vdd.n676 vdd.n675 9.3005
R18888 vdd.n3242 vdd.n3241 9.3005
R18889 vdd.n3243 vdd.n674 9.3005
R18890 vdd.n3245 vdd.n3244 9.3005
R18891 vdd.n666 vdd.n665 9.3005
R18892 vdd.n3259 vdd.n3258 9.3005
R18893 vdd.n3260 vdd.n664 9.3005
R18894 vdd.n3262 vdd.n3261 9.3005
R18895 vdd.n653 vdd.n652 9.3005
R18896 vdd.n3275 vdd.n3274 9.3005
R18897 vdd.n3276 vdd.n651 9.3005
R18898 vdd.n3278 vdd.n3277 9.3005
R18899 vdd.n642 vdd.n641 9.3005
R18900 vdd.n3292 vdd.n3291 9.3005
R18901 vdd.n3293 vdd.n640 9.3005
R18902 vdd.n3298 vdd.n3294 9.3005
R18903 vdd.n3297 vdd.n3296 9.3005
R18904 vdd.n3295 vdd.n631 9.3005
R18905 vdd.n3311 vdd.n630 9.3005
R18906 vdd.n3313 vdd.n3312 9.3005
R18907 vdd.n3314 vdd.n629 9.3005
R18908 vdd.n3316 vdd.n3315 9.3005
R18909 vdd.n3318 vdd.n628 9.3005
R18910 vdd.n3320 vdd.n3319 9.3005
R18911 vdd.n3321 vdd.n627 9.3005
R18912 vdd.n3323 vdd.n3322 9.3005
R18913 vdd.n3325 vdd.n626 9.3005
R18914 vdd.n3327 vdd.n3326 9.3005
R18915 vdd.n3328 vdd.n625 9.3005
R18916 vdd.n3330 vdd.n3329 9.3005
R18917 vdd.n3333 vdd.n624 9.3005
R18918 vdd.n3335 vdd.n3334 9.3005
R18919 vdd.n3336 vdd.n623 9.3005
R18920 vdd.n3338 vdd.n3337 9.3005
R18921 vdd.n3340 vdd.n622 9.3005
R18922 vdd.n3342 vdd.n3341 9.3005
R18923 vdd.n3343 vdd.n621 9.3005
R18924 vdd.n3345 vdd.n3344 9.3005
R18925 vdd.n3347 vdd.n620 9.3005
R18926 vdd.n3349 vdd.n3348 9.3005
R18927 vdd.n3227 vdd.n686 9.3005
R18928 vdd.n3226 vdd.n3225 9.3005
R18929 vdd.n3095 vdd.n687 9.3005
R18930 vdd.n3104 vdd.n783 9.3005
R18931 vdd.n3107 vdd.n782 9.3005
R18932 vdd.n3108 vdd.n781 9.3005
R18933 vdd.n3111 vdd.n780 9.3005
R18934 vdd.n3112 vdd.n779 9.3005
R18935 vdd.n3115 vdd.n778 9.3005
R18936 vdd.n3116 vdd.n777 9.3005
R18937 vdd.n3119 vdd.n776 9.3005
R18938 vdd.n3120 vdd.n775 9.3005
R18939 vdd.n3123 vdd.n774 9.3005
R18940 vdd.n3124 vdd.n773 9.3005
R18941 vdd.n3127 vdd.n772 9.3005
R18942 vdd.n3128 vdd.n771 9.3005
R18943 vdd.n3131 vdd.n770 9.3005
R18944 vdd.n3135 vdd.n3134 9.3005
R18945 vdd.n3136 vdd.n767 9.3005
R18946 vdd.n2337 vdd.n2336 9.3005
R18947 vdd.n2332 vdd.n1067 9.3005
R18948 vdd.n1430 vdd.n1429 9.3005
R18949 vdd.n1431 vdd.n1185 9.3005
R18950 vdd.n1433 vdd.n1432 9.3005
R18951 vdd.n1175 vdd.n1174 9.3005
R18952 vdd.n1447 vdd.n1446 9.3005
R18953 vdd.n1448 vdd.n1173 9.3005
R18954 vdd.n1450 vdd.n1449 9.3005
R18955 vdd.n1165 vdd.n1164 9.3005
R18956 vdd.n1464 vdd.n1463 9.3005
R18957 vdd.n1465 vdd.n1163 9.3005
R18958 vdd.n1467 vdd.n1466 9.3005
R18959 vdd.n1152 vdd.n1151 9.3005
R18960 vdd.n1480 vdd.n1479 9.3005
R18961 vdd.n1481 vdd.n1150 9.3005
R18962 vdd.n1483 vdd.n1482 9.3005
R18963 vdd.n1141 vdd.n1140 9.3005
R18964 vdd.n1497 vdd.n1496 9.3005
R18965 vdd.n1498 vdd.n1139 9.3005
R18966 vdd.n1500 vdd.n1499 9.3005
R18967 vdd.n1130 vdd.n1129 9.3005
R18968 vdd.n1820 vdd.n1819 9.3005
R18969 vdd.n1821 vdd.n1128 9.3005
R18970 vdd.n1823 vdd.n1822 9.3005
R18971 vdd.n1118 vdd.n1117 9.3005
R18972 vdd.n1837 vdd.n1836 9.3005
R18973 vdd.n1838 vdd.n1116 9.3005
R18974 vdd.n1840 vdd.n1839 9.3005
R18975 vdd.n1108 vdd.n1107 9.3005
R18976 vdd.n1854 vdd.n1853 9.3005
R18977 vdd.n1855 vdd.n1106 9.3005
R18978 vdd.n1857 vdd.n1856 9.3005
R18979 vdd.n1095 vdd.n1094 9.3005
R18980 vdd.n1870 vdd.n1869 9.3005
R18981 vdd.n1871 vdd.n1093 9.3005
R18982 vdd.n1873 vdd.n1872 9.3005
R18983 vdd.n1085 vdd.n1084 9.3005
R18984 vdd.n1887 vdd.n1886 9.3005
R18985 vdd.n1888 vdd.n1082 9.3005
R18986 vdd.n1892 vdd.n1891 9.3005
R18987 vdd.n1890 vdd.n1083 9.3005
R18988 vdd.n1889 vdd.n1072 9.3005
R18989 vdd.n1187 vdd.n1186 9.3005
R18990 vdd.n1323 vdd.n1322 9.3005
R18991 vdd.n1324 vdd.n1313 9.3005
R18992 vdd.n1326 vdd.n1325 9.3005
R18993 vdd.n1327 vdd.n1312 9.3005
R18994 vdd.n1329 vdd.n1328 9.3005
R18995 vdd.n1330 vdd.n1307 9.3005
R18996 vdd.n1332 vdd.n1331 9.3005
R18997 vdd.n1333 vdd.n1306 9.3005
R18998 vdd.n1335 vdd.n1334 9.3005
R18999 vdd.n1336 vdd.n1301 9.3005
R19000 vdd.n1338 vdd.n1337 9.3005
R19001 vdd.n1339 vdd.n1300 9.3005
R19002 vdd.n1341 vdd.n1340 9.3005
R19003 vdd.n1342 vdd.n1295 9.3005
R19004 vdd.n1344 vdd.n1343 9.3005
R19005 vdd.n1345 vdd.n1294 9.3005
R19006 vdd.n1347 vdd.n1346 9.3005
R19007 vdd.n1348 vdd.n1289 9.3005
R19008 vdd.n1350 vdd.n1349 9.3005
R19009 vdd.n1351 vdd.n1288 9.3005
R19010 vdd.n1353 vdd.n1352 9.3005
R19011 vdd.n1357 vdd.n1284 9.3005
R19012 vdd.n1359 vdd.n1358 9.3005
R19013 vdd.n1360 vdd.n1283 9.3005
R19014 vdd.n1362 vdd.n1361 9.3005
R19015 vdd.n1363 vdd.n1278 9.3005
R19016 vdd.n1365 vdd.n1364 9.3005
R19017 vdd.n1366 vdd.n1277 9.3005
R19018 vdd.n1368 vdd.n1367 9.3005
R19019 vdd.n1369 vdd.n1272 9.3005
R19020 vdd.n1371 vdd.n1370 9.3005
R19021 vdd.n1372 vdd.n1271 9.3005
R19022 vdd.n1374 vdd.n1373 9.3005
R19023 vdd.n1375 vdd.n1266 9.3005
R19024 vdd.n1377 vdd.n1376 9.3005
R19025 vdd.n1378 vdd.n1265 9.3005
R19026 vdd.n1380 vdd.n1379 9.3005
R19027 vdd.n1381 vdd.n1260 9.3005
R19028 vdd.n1383 vdd.n1382 9.3005
R19029 vdd.n1384 vdd.n1259 9.3005
R19030 vdd.n1386 vdd.n1385 9.3005
R19031 vdd.n1387 vdd.n1254 9.3005
R19032 vdd.n1389 vdd.n1388 9.3005
R19033 vdd.n1390 vdd.n1253 9.3005
R19034 vdd.n1392 vdd.n1391 9.3005
R19035 vdd.n1393 vdd.n1246 9.3005
R19036 vdd.n1395 vdd.n1394 9.3005
R19037 vdd.n1396 vdd.n1245 9.3005
R19038 vdd.n1398 vdd.n1397 9.3005
R19039 vdd.n1399 vdd.n1240 9.3005
R19040 vdd.n1401 vdd.n1400 9.3005
R19041 vdd.n1402 vdd.n1239 9.3005
R19042 vdd.n1404 vdd.n1403 9.3005
R19043 vdd.n1405 vdd.n1234 9.3005
R19044 vdd.n1407 vdd.n1406 9.3005
R19045 vdd.n1408 vdd.n1233 9.3005
R19046 vdd.n1410 vdd.n1409 9.3005
R19047 vdd.n1411 vdd.n1228 9.3005
R19048 vdd.n1413 vdd.n1412 9.3005
R19049 vdd.n1414 vdd.n1227 9.3005
R19050 vdd.n1416 vdd.n1415 9.3005
R19051 vdd.n1192 vdd.n1191 9.3005
R19052 vdd.n1422 vdd.n1421 9.3005
R19053 vdd.n1321 vdd.n1320 9.3005
R19054 vdd.n1425 vdd.n1424 9.3005
R19055 vdd.n1181 vdd.n1180 9.3005
R19056 vdd.n1439 vdd.n1438 9.3005
R19057 vdd.n1440 vdd.n1179 9.3005
R19058 vdd.n1442 vdd.n1441 9.3005
R19059 vdd.n1170 vdd.n1169 9.3005
R19060 vdd.n1456 vdd.n1455 9.3005
R19061 vdd.n1457 vdd.n1168 9.3005
R19062 vdd.n1459 vdd.n1458 9.3005
R19063 vdd.n1159 vdd.n1158 9.3005
R19064 vdd.n1472 vdd.n1471 9.3005
R19065 vdd.n1473 vdd.n1157 9.3005
R19066 vdd.n1475 vdd.n1474 9.3005
R19067 vdd.n1147 vdd.n1146 9.3005
R19068 vdd.n1489 vdd.n1488 9.3005
R19069 vdd.n1490 vdd.n1145 9.3005
R19070 vdd.n1492 vdd.n1491 9.3005
R19071 vdd.n1136 vdd.n1135 9.3005
R19072 vdd.n1505 vdd.n1504 9.3005
R19073 vdd.n1506 vdd.n1134 9.3005
R19074 vdd.n1423 vdd.n1190 9.3005
R19075 vdd.n1726 vdd.n1725 9.3005
R19076 vdd.n1721 vdd.n1720 9.3005
R19077 vdd.n1732 vdd.n1731 9.3005
R19078 vdd.n1734 vdd.n1733 9.3005
R19079 vdd.n1717 vdd.n1716 9.3005
R19080 vdd.n1740 vdd.n1739 9.3005
R19081 vdd.n1742 vdd.n1741 9.3005
R19082 vdd.n1714 vdd.n1711 9.3005
R19083 vdd.n1749 vdd.n1748 9.3005
R19084 vdd.n1785 vdd.n1784 9.3005
R19085 vdd.n1780 vdd.n1779 9.3005
R19086 vdd.n1791 vdd.n1790 9.3005
R19087 vdd.n1793 vdd.n1792 9.3005
R19088 vdd.n1776 vdd.n1775 9.3005
R19089 vdd.n1799 vdd.n1798 9.3005
R19090 vdd.n1801 vdd.n1800 9.3005
R19091 vdd.n1773 vdd.n1770 9.3005
R19092 vdd.n1808 vdd.n1807 9.3005
R19093 vdd.n1624 vdd.n1623 9.3005
R19094 vdd.n1619 vdd.n1618 9.3005
R19095 vdd.n1630 vdd.n1629 9.3005
R19096 vdd.n1632 vdd.n1631 9.3005
R19097 vdd.n1615 vdd.n1614 9.3005
R19098 vdd.n1638 vdd.n1637 9.3005
R19099 vdd.n1640 vdd.n1639 9.3005
R19100 vdd.n1612 vdd.n1609 9.3005
R19101 vdd.n1647 vdd.n1646 9.3005
R19102 vdd.n1683 vdd.n1682 9.3005
R19103 vdd.n1678 vdd.n1677 9.3005
R19104 vdd.n1689 vdd.n1688 9.3005
R19105 vdd.n1691 vdd.n1690 9.3005
R19106 vdd.n1674 vdd.n1673 9.3005
R19107 vdd.n1697 vdd.n1696 9.3005
R19108 vdd.n1699 vdd.n1698 9.3005
R19109 vdd.n1671 vdd.n1668 9.3005
R19110 vdd.n1706 vdd.n1705 9.3005
R19111 vdd.n1523 vdd.n1522 9.3005
R19112 vdd.n1518 vdd.n1517 9.3005
R19113 vdd.n1529 vdd.n1528 9.3005
R19114 vdd.n1531 vdd.n1530 9.3005
R19115 vdd.n1514 vdd.n1513 9.3005
R19116 vdd.n1537 vdd.n1536 9.3005
R19117 vdd.n1539 vdd.n1538 9.3005
R19118 vdd.n1511 vdd.n1508 9.3005
R19119 vdd.n1546 vdd.n1545 9.3005
R19120 vdd.n1582 vdd.n1581 9.3005
R19121 vdd.n1577 vdd.n1576 9.3005
R19122 vdd.n1588 vdd.n1587 9.3005
R19123 vdd.n1590 vdd.n1589 9.3005
R19124 vdd.n1573 vdd.n1572 9.3005
R19125 vdd.n1596 vdd.n1595 9.3005
R19126 vdd.n1598 vdd.n1597 9.3005
R19127 vdd.n1570 vdd.n1567 9.3005
R19128 vdd.n1605 vdd.n1604 9.3005
R19129 vdd.n1461 vdd.t178 9.18308
R19130 vdd.n3331 vdd.t245 9.18308
R19131 vdd.n1155 vdd.t227 8.95635
R19132 vdd.n2329 vdd.t66 8.95635
R19133 vdd.n723 vdd.t59 8.95635
R19134 vdd.t191 vdd.n3385 8.95635
R19135 vdd.n312 vdd.n311 8.92171
R19136 vdd.n253 vdd.n252 8.92171
R19137 vdd.n210 vdd.n209 8.92171
R19138 vdd.n151 vdd.n150 8.92171
R19139 vdd.n109 vdd.n108 8.92171
R19140 vdd.n50 vdd.n49 8.92171
R19141 vdd.n1731 vdd.n1730 8.92171
R19142 vdd.n1790 vdd.n1789 8.92171
R19143 vdd.n1629 vdd.n1628 8.92171
R19144 vdd.n1688 vdd.n1687 8.92171
R19145 vdd.n1528 vdd.n1527 8.92171
R19146 vdd.n1587 vdd.n1586 8.92171
R19147 vdd.n231 vdd.n129 8.81535
R19148 vdd.n1709 vdd.n1607 8.81535
R19149 vdd.n1502 vdd.t199 8.72962
R19150 vdd.t136 vdd.n3394 8.72962
R19151 vdd.n1825 vdd.t248 8.50289
R19152 vdd.n3300 vdd.t193 8.50289
R19153 vdd.n28 vdd.n14 8.42249
R19154 vdd.n1851 vdd.t187 8.27616
R19155 vdd.t185 vdd.n656 8.27616
R19156 vdd.n3400 vdd.n3399 8.16225
R19157 vdd.n1813 vdd.n1812 8.16225
R19158 vdd.n308 vdd.n302 8.14595
R19159 vdd.n249 vdd.n243 8.14595
R19160 vdd.n206 vdd.n200 8.14595
R19161 vdd.n147 vdd.n141 8.14595
R19162 vdd.n105 vdd.n99 8.14595
R19163 vdd.n46 vdd.n40 8.14595
R19164 vdd.n1727 vdd.n1721 8.14595
R19165 vdd.n1786 vdd.n1780 8.14595
R19166 vdd.n1625 vdd.n1619 8.14595
R19167 vdd.n1684 vdd.n1678 8.14595
R19168 vdd.n1524 vdd.n1518 8.14595
R19169 vdd.n1583 vdd.n1577 8.14595
R19170 vdd.n2923 vdd.n849 8.11757
R19171 vdd.n2397 vdd.n2396 8.11757
R19172 vdd.n1098 vdd.t271 8.04943
R19173 vdd.n3256 vdd.t225 8.04943
R19174 vdd.n2375 vdd.n1043 7.70933
R19175 vdd.n2381 vdd.n1043 7.70933
R19176 vdd.n2387 vdd.n1037 7.70933
R19177 vdd.n2387 vdd.n1030 7.70933
R19178 vdd.n2393 vdd.n1030 7.70933
R19179 vdd.n2393 vdd.n1033 7.70933
R19180 vdd.n2400 vdd.n1018 7.70933
R19181 vdd.n2406 vdd.n1018 7.70933
R19182 vdd.n2412 vdd.n1012 7.70933
R19183 vdd.n2418 vdd.n1008 7.70933
R19184 vdd.n2424 vdd.n1002 7.70933
R19185 vdd.n2436 vdd.n989 7.70933
R19186 vdd.n2442 vdd.n983 7.70933
R19187 vdd.n2442 vdd.n976 7.70933
R19188 vdd.n2450 vdd.n976 7.70933
R19189 vdd.n2457 vdd.t35 7.70933
R19190 vdd.n2532 vdd.t35 7.70933
R19191 vdd.n2864 vdd.t132 7.70933
R19192 vdd.n2870 vdd.t132 7.70933
R19193 vdd.n2876 vdd.n897 7.70933
R19194 vdd.n2882 vdd.n897 7.70933
R19195 vdd.n2882 vdd.n900 7.70933
R19196 vdd.n2888 vdd.n893 7.70933
R19197 vdd.n2900 vdd.n880 7.70933
R19198 vdd.n2906 vdd.n874 7.70933
R19199 vdd.n2912 vdd.n870 7.70933
R19200 vdd.n2918 vdd.n857 7.70933
R19201 vdd.n2926 vdd.n857 7.70933
R19202 vdd.n2932 vdd.n851 7.70933
R19203 vdd.n2932 vdd.n843 7.70933
R19204 vdd.n2983 vdd.n843 7.70933
R19205 vdd.n2983 vdd.n846 7.70933
R19206 vdd.n2989 vdd.n805 7.70933
R19207 vdd.n3059 vdd.n805 7.70933
R19208 vdd.n307 vdd.n304 7.3702
R19209 vdd.n248 vdd.n245 7.3702
R19210 vdd.n205 vdd.n202 7.3702
R19211 vdd.n146 vdd.n143 7.3702
R19212 vdd.n104 vdd.n101 7.3702
R19213 vdd.n45 vdd.n42 7.3702
R19214 vdd.n1726 vdd.n1723 7.3702
R19215 vdd.n1785 vdd.n1782 7.3702
R19216 vdd.n1624 vdd.n1621 7.3702
R19217 vdd.n1683 vdd.n1680 7.3702
R19218 vdd.n1523 vdd.n1520 7.3702
R19219 vdd.n1582 vdd.n1579 7.3702
R19220 vdd.n1884 vdd.t144 7.1425
R19221 vdd.n679 vdd.t140 7.1425
R19222 vdd.n1358 vdd.n1357 6.98232
R19223 vdd.n2039 vdd.n2038 6.98232
R19224 vdd.n566 vdd.n565 6.98232
R19225 vdd.n3141 vdd.n3138 6.98232
R19226 vdd.t250 vdd.n1097 6.91577
R19227 vdd.n3264 vdd.t150 6.91577
R19228 vdd.n1843 vdd.t209 6.68904
R19229 vdd.n3280 vdd.t134 6.68904
R19230 vdd.t155 vdd.n1126 6.46231
R19231 vdd.n3308 vdd.t152 6.46231
R19232 vdd.n3400 vdd.n333 6.38151
R19233 vdd.n1812 vdd.n1811 6.38151
R19234 vdd.n1494 vdd.t182 6.23558
R19235 vdd.t220 vdd.n344 6.23558
R19236 vdd.t138 vdd.n1154 6.00885
R19237 vdd.n2412 vdd.t24 6.00885
R19238 vdd.n2912 vdd.t22 6.00885
R19239 vdd.n3379 vdd.t168 6.00885
R19240 vdd.n1033 vdd.t112 5.89549
R19241 vdd.t70 vdd.n851 5.89549
R19242 vdd.n308 vdd.n307 5.81868
R19243 vdd.n249 vdd.n248 5.81868
R19244 vdd.n206 vdd.n205 5.81868
R19245 vdd.n147 vdd.n146 5.81868
R19246 vdd.n105 vdd.n104 5.81868
R19247 vdd.n46 vdd.n45 5.81868
R19248 vdd.n1727 vdd.n1726 5.81868
R19249 vdd.n1786 vdd.n1785 5.81868
R19250 vdd.n1625 vdd.n1624 5.81868
R19251 vdd.n1684 vdd.n1683 5.81868
R19252 vdd.n1524 vdd.n1523 5.81868
R19253 vdd.n1583 vdd.n1582 5.81868
R19254 vdd.n1453 vdd.t142 5.78212
R19255 vdd.t55 vdd.n1037 5.78212
R19256 vdd.n2156 vdd.t94 5.78212
R19257 vdd.n2781 vdd.t102 5.78212
R19258 vdd.n846 vdd.t98 5.78212
R19259 vdd.n3370 vdd.t214 5.78212
R19260 vdd.n2540 vdd.n2539 5.77611
R19261 vdd.n2283 vdd.n2153 5.77611
R19262 vdd.n2794 vdd.n2793 5.77611
R19263 vdd.n3000 vdd.n2999 5.77611
R19264 vdd.n3064 vdd.n801 5.77611
R19265 vdd.n2704 vdd.n2644 5.77611
R19266 vdd.n2465 vdd.n967 5.77611
R19267 vdd.n2213 vdd.n2212 5.77611
R19268 vdd.n1320 vdd.n1319 5.62474
R19269 vdd.n2335 vdd.n2332 5.62474
R19270 vdd.n3351 vdd.n428 5.62474
R19271 vdd.n3225 vdd.n690 5.62474
R19272 vdd.n1177 vdd.t142 5.55539
R19273 vdd.t214 vdd.n3369 5.55539
R19274 vdd.t11 vdd.n989 5.44203
R19275 vdd.n893 vdd.t31 5.44203
R19276 vdd.n1469 vdd.t138 5.32866
R19277 vdd.t168 vdd.n3378 5.32866
R19278 vdd.n1485 vdd.t182 5.10193
R19279 vdd.t47 vdd.n1012 5.10193
R19280 vdd.n1002 vdd.t25 5.10193
R19281 vdd.t30 vdd.n880 5.10193
R19282 vdd.n870 vdd.t19 5.10193
R19283 vdd.n3387 vdd.t220 5.10193
R19284 vdd.n311 vdd.n302 5.04292
R19285 vdd.n252 vdd.n243 5.04292
R19286 vdd.n209 vdd.n200 5.04292
R19287 vdd.n150 vdd.n141 5.04292
R19288 vdd.n108 vdd.n99 5.04292
R19289 vdd.n49 vdd.n40 5.04292
R19290 vdd.n1730 vdd.n1721 5.04292
R19291 vdd.n1789 vdd.n1780 5.04292
R19292 vdd.n1628 vdd.n1619 5.04292
R19293 vdd.n1687 vdd.n1678 5.04292
R19294 vdd.n1527 vdd.n1518 5.04292
R19295 vdd.n1586 vdd.n1577 5.04292
R19296 vdd.n1817 vdd.t155 4.8752
R19297 vdd.t23 vdd.t39 4.8752
R19298 vdd.t50 vdd.t130 4.8752
R19299 vdd.t28 vdd.t10 4.8752
R19300 vdd.t294 vdd.t46 4.8752
R19301 vdd.t152 vdd.n340 4.8752
R19302 vdd.n2541 vdd.n2540 4.83952
R19303 vdd.n2153 vdd.n2149 4.83952
R19304 vdd.n2795 vdd.n2794 4.83952
R19305 vdd.n3001 vdd.n3000 4.83952
R19306 vdd.n801 vdd.n796 4.83952
R19307 vdd.n2701 vdd.n2644 4.83952
R19308 vdd.n2468 vdd.n967 4.83952
R19309 vdd.n2212 vdd.n2211 4.83952
R19310 vdd.n2007 vdd.n1065 4.74817
R19311 vdd.n2002 vdd.n1066 4.74817
R19312 vdd.n1904 vdd.n1901 4.74817
R19313 vdd.n2316 vdd.n1905 4.74817
R19314 vdd.n2318 vdd.n1904 4.74817
R19315 vdd.n2317 vdd.n2316 4.74817
R19316 vdd.n3218 vdd.n3217 4.74817
R19317 vdd.n3215 vdd.n3214 4.74817
R19318 vdd.n3215 vdd.n732 4.74817
R19319 vdd.n3217 vdd.n729 4.74817
R19320 vdd.n3100 vdd.n784 4.74817
R19321 vdd.n3096 vdd.n3094 4.74817
R19322 vdd.n3099 vdd.n3094 4.74817
R19323 vdd.n3103 vdd.n784 4.74817
R19324 vdd.n2003 vdd.n1065 4.74817
R19325 vdd.n1068 vdd.n1066 4.74817
R19326 vdd.n333 vdd.n332 4.7074
R19327 vdd.n231 vdd.n230 4.7074
R19328 vdd.n1811 vdd.n1810 4.7074
R19329 vdd.n1709 vdd.n1708 4.7074
R19330 vdd.n1120 vdd.t209 4.64847
R19331 vdd.n3289 vdd.t134 4.64847
R19332 vdd.n2418 vdd.t33 4.53511
R19333 vdd.n2906 vdd.t41 4.53511
R19334 vdd.n1859 vdd.t250 4.42174
R19335 vdd.t150 vdd.n655 4.42174
R19336 vdd.n2450 vdd.t20 4.30838
R19337 vdd.n2876 vdd.t14 4.30838
R19338 vdd.n312 vdd.n300 4.26717
R19339 vdd.n253 vdd.n241 4.26717
R19340 vdd.n210 vdd.n198 4.26717
R19341 vdd.n151 vdd.n139 4.26717
R19342 vdd.n109 vdd.n97 4.26717
R19343 vdd.n50 vdd.n38 4.26717
R19344 vdd.n1731 vdd.n1719 4.26717
R19345 vdd.n1790 vdd.n1778 4.26717
R19346 vdd.n1629 vdd.n1617 4.26717
R19347 vdd.n1688 vdd.n1676 4.26717
R19348 vdd.n1528 vdd.n1516 4.26717
R19349 vdd.n1587 vdd.n1575 4.26717
R19350 vdd.n1875 vdd.t144 4.19501
R19351 vdd.n3248 vdd.t140 4.19501
R19352 vdd.n333 vdd.n231 4.10845
R19353 vdd.n1811 vdd.n1709 4.10845
R19354 vdd.n289 vdd.t177 4.06363
R19355 vdd.n289 vdd.t238 4.06363
R19356 vdd.n287 vdd.t268 4.06363
R19357 vdd.n287 vdd.t285 4.06363
R19358 vdd.n285 vdd.t289 4.06363
R19359 vdd.n285 vdd.t184 4.06363
R19360 vdd.n283 vdd.t207 4.06363
R19361 vdd.n283 vdd.t288 4.06363
R19362 vdd.n281 vdd.t290 4.06363
R19363 vdd.n281 vdd.t206 4.06363
R19364 vdd.n279 vdd.t211 4.06363
R19365 vdd.n279 vdd.t213 4.06363
R19366 vdd.n277 vdd.t264 4.06363
R19367 vdd.n277 vdd.t167 4.06363
R19368 vdd.n275 vdd.t173 4.06363
R19369 vdd.n275 vdd.t237 4.06363
R19370 vdd.n273 vdd.t241 4.06363
R19371 vdd.n273 vdd.t270 4.06363
R19372 vdd.n187 vdd.t160 4.06363
R19373 vdd.n187 vdd.t215 4.06363
R19374 vdd.n185 vdd.t255 4.06363
R19375 vdd.n185 vdd.t273 4.06363
R19376 vdd.n183 vdd.t277 4.06363
R19377 vdd.n183 vdd.t162 4.06363
R19378 vdd.n181 vdd.t190 4.06363
R19379 vdd.n181 vdd.t276 4.06363
R19380 vdd.n179 vdd.t280 4.06363
R19381 vdd.n179 vdd.t137 4.06363
R19382 vdd.n177 vdd.t194 4.06363
R19383 vdd.n177 vdd.t196 4.06363
R19384 vdd.n175 vdd.t254 4.06363
R19385 vdd.n175 vdd.t135 4.06363
R19386 vdd.n173 vdd.t151 4.06363
R19387 vdd.n173 vdd.t216 4.06363
R19388 vdd.n171 vdd.t226 4.06363
R19389 vdd.n171 vdd.t256 4.06363
R19390 vdd.n86 vdd.t176 4.06363
R19391 vdd.n86 vdd.t261 4.06363
R19392 vdd.n84 vdd.t169 4.06363
R19393 vdd.n84 vdd.t246 4.06363
R19394 vdd.n82 vdd.t192 4.06363
R19395 vdd.n82 vdd.t274 4.06363
R19396 vdd.n80 vdd.t164 4.06363
R19397 vdd.n80 vdd.t221 4.06363
R19398 vdd.n78 vdd.t153 4.06363
R19399 vdd.n78 vdd.t197 4.06363
R19400 vdd.n76 vdd.t286 4.06363
R19401 vdd.n76 vdd.t260 4.06363
R19402 vdd.n74 vdd.t266 4.06363
R19403 vdd.n74 vdd.t208 4.06363
R19404 vdd.n72 vdd.t291 4.06363
R19405 vdd.n72 vdd.t186 4.06363
R19406 vdd.n70 vdd.t278 4.06363
R19407 vdd.n70 vdd.t218 4.06363
R19408 vdd.n1751 vdd.t175 4.06363
R19409 vdd.n1751 vdd.t284 4.06363
R19410 vdd.n1753 vdd.t281 4.06363
R19411 vdd.n1753 vdd.t262 4.06363
R19412 vdd.n1755 vdd.t231 4.06363
R19413 vdd.n1755 vdd.t171 4.06363
R19414 vdd.n1757 vdd.t293 4.06363
R19415 vdd.n1757 vdd.t259 4.06363
R19416 vdd.n1759 vdd.t257 4.06363
R19417 vdd.n1759 vdd.t205 4.06363
R19418 vdd.n1761 vdd.t201 4.06363
R19419 vdd.n1761 vdd.t232 4.06363
R19420 vdd.n1763 vdd.t233 4.06363
R19421 vdd.n1763 vdd.t242 4.06363
R19422 vdd.n1765 vdd.t198 4.06363
R19423 vdd.n1765 vdd.t174 4.06363
R19424 vdd.n1767 vdd.t170 4.06363
R19425 vdd.n1767 vdd.t239 4.06363
R19426 vdd.n1649 vdd.t158 4.06363
R19427 vdd.n1649 vdd.t272 4.06363
R19428 vdd.n1651 vdd.t265 4.06363
R19429 vdd.n1651 vdd.t251 4.06363
R19430 vdd.n1653 vdd.t212 4.06363
R19431 vdd.n1653 vdd.t147 4.06363
R19432 vdd.n1655 vdd.t282 4.06363
R19433 vdd.n1655 vdd.t249 4.06363
R19434 vdd.n1657 vdd.t243 4.06363
R19435 vdd.n1657 vdd.t189 4.06363
R19436 vdd.n1659 vdd.t183 4.06363
R19437 vdd.n1659 vdd.t244 4.06363
R19438 vdd.n1661 vdd.t230 4.06363
R19439 vdd.n1661 vdd.t228 4.06363
R19440 vdd.n1663 vdd.t179 4.06363
R19441 vdd.n1663 vdd.t154 4.06363
R19442 vdd.n1665 vdd.t143 4.06363
R19443 vdd.n1665 vdd.t223 4.06363
R19444 vdd.n1548 vdd.t219 4.06363
R19445 vdd.n1548 vdd.t279 4.06363
R19446 vdd.n1550 vdd.t188 4.06363
R19447 vdd.n1550 vdd.t258 4.06363
R19448 vdd.n1552 vdd.t210 4.06363
R19449 vdd.n1552 vdd.t267 4.06363
R19450 vdd.n1554 vdd.t235 4.06363
R19451 vdd.n1554 vdd.t287 4.06363
R19452 vdd.n1556 vdd.t200 4.06363
R19453 vdd.n1556 vdd.t156 4.06363
R19454 vdd.n1558 vdd.t222 4.06363
R19455 vdd.n1558 vdd.t166 4.06363
R19456 vdd.n1560 vdd.t275 4.06363
R19457 vdd.n1560 vdd.t292 4.06363
R19458 vdd.n1562 vdd.t247 4.06363
R19459 vdd.n1562 vdd.t139 4.06363
R19460 vdd.n1564 vdd.t236 4.06363
R19461 vdd.n1564 vdd.t181 4.06363
R19462 vdd.n26 vdd.t53 3.9605
R19463 vdd.n26 vdd.t7 3.9605
R19464 vdd.n23 vdd.t6 3.9605
R19465 vdd.n23 vdd.t18 3.9605
R19466 vdd.n21 vdd.t16 3.9605
R19467 vdd.n21 vdd.t2 3.9605
R19468 vdd.n20 vdd.t9 3.9605
R19469 vdd.n20 vdd.t5 3.9605
R19470 vdd.n15 vdd.t3 3.9605
R19471 vdd.n15 vdd.t4 3.9605
R19472 vdd.n16 vdd.t8 3.9605
R19473 vdd.n16 vdd.t51 3.9605
R19474 vdd.n18 vdd.t17 3.9605
R19475 vdd.n18 vdd.t0 3.9605
R19476 vdd.n25 vdd.t52 3.9605
R19477 vdd.n25 vdd.t1 3.9605
R19478 vdd.n7 vdd.t295 3.61217
R19479 vdd.n7 vdd.t42 3.61217
R19480 vdd.n8 vdd.t29 3.61217
R19481 vdd.n8 vdd.t32 3.61217
R19482 vdd.n10 vdd.t133 3.61217
R19483 vdd.n10 vdd.t15 3.61217
R19484 vdd.n12 vdd.t49 3.61217
R19485 vdd.n12 vdd.t45 3.61217
R19486 vdd.n5 vdd.t38 3.61217
R19487 vdd.n5 vdd.t27 3.61217
R19488 vdd.n3 vdd.t21 3.61217
R19489 vdd.n3 vdd.t36 3.61217
R19490 vdd.n1 vdd.t12 3.61217
R19491 vdd.n1 vdd.t131 3.61217
R19492 vdd.n0 vdd.t34 3.61217
R19493 vdd.n0 vdd.t40 3.61217
R19494 vdd.n316 vdd.n315 3.49141
R19495 vdd.n257 vdd.n256 3.49141
R19496 vdd.n214 vdd.n213 3.49141
R19497 vdd.n155 vdd.n154 3.49141
R19498 vdd.n113 vdd.n112 3.49141
R19499 vdd.n54 vdd.n53 3.49141
R19500 vdd.n1735 vdd.n1734 3.49141
R19501 vdd.n1794 vdd.n1793 3.49141
R19502 vdd.n1633 vdd.n1632 3.49141
R19503 vdd.n1692 vdd.n1691 3.49141
R19504 vdd.n1532 vdd.n1531 3.49141
R19505 vdd.n1591 vdd.n1590 3.49141
R19506 vdd.n2156 vdd.t20 3.40145
R19507 vdd.n2604 vdd.t37 3.40145
R19508 vdd.n2857 vdd.t44 3.40145
R19509 vdd.n2781 vdd.t14 3.40145
R19510 vdd.n1876 vdd.t271 3.28809
R19511 vdd.n3247 vdd.t225 3.28809
R19512 vdd.n2257 vdd.t33 3.17472
R19513 vdd.n2760 vdd.t41 3.17472
R19514 vdd.t187 vdd.n1104 3.06136
R19515 vdd.n3272 vdd.t185 3.06136
R19516 vdd.n1834 vdd.t248 2.83463
R19517 vdd.n644 vdd.t193 2.83463
R19518 vdd.n319 vdd.n298 2.71565
R19519 vdd.n260 vdd.n239 2.71565
R19520 vdd.n217 vdd.n196 2.71565
R19521 vdd.n158 vdd.n137 2.71565
R19522 vdd.n116 vdd.n95 2.71565
R19523 vdd.n57 vdd.n36 2.71565
R19524 vdd.n1738 vdd.n1717 2.71565
R19525 vdd.n1797 vdd.n1776 2.71565
R19526 vdd.n1636 vdd.n1615 2.71565
R19527 vdd.n1695 vdd.n1674 2.71565
R19528 vdd.n1535 vdd.n1514 2.71565
R19529 vdd.n1594 vdd.n1573 2.71565
R19530 vdd.t199 vdd.n1132 2.6079
R19531 vdd.n2406 vdd.t47 2.6079
R19532 vdd.n2430 vdd.t25 2.6079
R19533 vdd.n2894 vdd.t30 2.6079
R19534 vdd.n2918 vdd.t19 2.6079
R19535 vdd.n3395 vdd.t136 2.6079
R19536 vdd.n2924 vdd.n2923 2.49806
R19537 vdd.n2398 vdd.n2397 2.49806
R19538 vdd.n306 vdd.n305 2.4129
R19539 vdd.n247 vdd.n246 2.4129
R19540 vdd.n204 vdd.n203 2.4129
R19541 vdd.n145 vdd.n144 2.4129
R19542 vdd.n103 vdd.n102 2.4129
R19543 vdd.n44 vdd.n43 2.4129
R19544 vdd.n1725 vdd.n1724 2.4129
R19545 vdd.n1784 vdd.n1783 2.4129
R19546 vdd.n1623 vdd.n1622 2.4129
R19547 vdd.n1682 vdd.n1681 2.4129
R19548 vdd.n1522 vdd.n1521 2.4129
R19549 vdd.n1581 vdd.n1580 2.4129
R19550 vdd.n1486 vdd.t227 2.38117
R19551 vdd.n1894 vdd.t66 2.38117
R19552 vdd.n3231 vdd.t59 2.38117
R19553 vdd.n3386 vdd.t191 2.38117
R19554 vdd.n2315 vdd.n1904 2.27742
R19555 vdd.n2316 vdd.n2315 2.27742
R19556 vdd.n3216 vdd.n3215 2.27742
R19557 vdd.n3217 vdd.n3216 2.27742
R19558 vdd.n3094 vdd.n3093 2.27742
R19559 vdd.n3093 vdd.n784 2.27742
R19560 vdd.n2338 vdd.n1065 2.27742
R19561 vdd.n2338 vdd.n1066 2.27742
R19562 vdd.n2430 vdd.t11 2.2678
R19563 vdd.n2894 vdd.t31 2.2678
R19564 vdd.t178 vdd.n1161 2.15444
R19565 vdd.n3377 vdd.t245 2.15444
R19566 vdd.t130 vdd.n983 2.04107
R19567 vdd.n900 vdd.t28 2.04107
R19568 vdd.n320 vdd.n296 1.93989
R19569 vdd.n261 vdd.n237 1.93989
R19570 vdd.n218 vdd.n194 1.93989
R19571 vdd.n159 vdd.n135 1.93989
R19572 vdd.n117 vdd.n93 1.93989
R19573 vdd.n58 vdd.n34 1.93989
R19574 vdd.n1739 vdd.n1715 1.93989
R19575 vdd.n1798 vdd.n1774 1.93989
R19576 vdd.n1637 vdd.n1613 1.93989
R19577 vdd.n1696 vdd.n1672 1.93989
R19578 vdd.n1536 vdd.n1512 1.93989
R19579 vdd.n1595 vdd.n1571 1.93989
R19580 vdd.n1444 vdd.t148 1.92771
R19581 vdd.n2381 vdd.t55 1.92771
R19582 vdd.n2457 vdd.t94 1.92771
R19583 vdd.n2870 vdd.t102 1.92771
R19584 vdd.n2989 vdd.t98 1.92771
R19585 vdd.t202 vdd.n375 1.92771
R19586 vdd.n1452 vdd.t180 1.70098
R19587 vdd.n2257 vdd.t24 1.70098
R19588 vdd.n1008 vdd.t23 1.70098
R19589 vdd.t46 vdd.n874 1.70098
R19590 vdd.n2760 vdd.t22 1.70098
R19591 vdd.n3371 vdd.t159 1.70098
R19592 vdd.n1477 vdd.t229 1.47425
R19593 vdd.n361 vdd.t161 1.47425
R19594 vdd.n1143 vdd.t165 1.24752
R19595 vdd.t163 vdd.n3393 1.24752
R19596 vdd.n331 vdd.n291 1.16414
R19597 vdd.n324 vdd.n323 1.16414
R19598 vdd.n272 vdd.n232 1.16414
R19599 vdd.n265 vdd.n264 1.16414
R19600 vdd.n229 vdd.n189 1.16414
R19601 vdd.n222 vdd.n221 1.16414
R19602 vdd.n170 vdd.n130 1.16414
R19603 vdd.n163 vdd.n162 1.16414
R19604 vdd.n128 vdd.n88 1.16414
R19605 vdd.n121 vdd.n120 1.16414
R19606 vdd.n69 vdd.n29 1.16414
R19607 vdd.n62 vdd.n61 1.16414
R19608 vdd.n1750 vdd.n1710 1.16414
R19609 vdd.n1743 vdd.n1742 1.16414
R19610 vdd.n1809 vdd.n1769 1.16414
R19611 vdd.n1802 vdd.n1801 1.16414
R19612 vdd.n1648 vdd.n1608 1.16414
R19613 vdd.n1641 vdd.n1640 1.16414
R19614 vdd.n1707 vdd.n1667 1.16414
R19615 vdd.n1700 vdd.n1699 1.16414
R19616 vdd.n1547 vdd.n1507 1.16414
R19617 vdd.n1540 vdd.n1539 1.16414
R19618 vdd.n1606 vdd.n1566 1.16414
R19619 vdd.n1599 vdd.n1598 1.16414
R19620 vdd.n2424 vdd.t39 1.13415
R19621 vdd.n2900 vdd.t294 1.13415
R19622 vdd.n1826 vdd.t234 1.02079
R19623 vdd.t112 vdd.t43 1.02079
R19624 vdd.t13 vdd.t70 1.02079
R19625 vdd.t195 vdd.n633 1.02079
R19626 vdd.n1323 vdd.n1319 0.970197
R19627 vdd.n2336 vdd.n2335 0.970197
R19628 vdd.n618 vdd.n428 0.970197
R19629 vdd.n3095 vdd.n690 0.970197
R19630 vdd.n1812 vdd.n28 0.90431
R19631 vdd vdd.n3400 0.896477
R19632 vdd.n1842 vdd.t146 0.794056
R19633 vdd.n2400 vdd.t43 0.794056
R19634 vdd.n2436 vdd.t50 0.794056
R19635 vdd.n2888 vdd.t10 0.794056
R19636 vdd.n2926 vdd.t13 0.794056
R19637 vdd.n3281 vdd.t253 0.794056
R19638 vdd.n1867 vdd.t157 0.567326
R19639 vdd.t217 vdd.n662 0.567326
R19640 vdd.n2326 vdd.n2325 0.530988
R19641 vdd.n726 vdd.n682 0.530988
R19642 vdd.n464 vdd.n391 0.530988
R19643 vdd.n3350 vdd.n3349 0.530988
R19644 vdd.n3227 vdd.n3226 0.530988
R19645 vdd.n1889 vdd.n1067 0.530988
R19646 vdd.n1321 vdd.n1186 0.530988
R19647 vdd.n1423 vdd.n1422 0.530988
R19648 vdd.n4 vdd.n2 0.459552
R19649 vdd.n11 vdd.n9 0.459552
R19650 vdd.n329 vdd.n328 0.388379
R19651 vdd.n295 vdd.n293 0.388379
R19652 vdd.n270 vdd.n269 0.388379
R19653 vdd.n236 vdd.n234 0.388379
R19654 vdd.n227 vdd.n226 0.388379
R19655 vdd.n193 vdd.n191 0.388379
R19656 vdd.n168 vdd.n167 0.388379
R19657 vdd.n134 vdd.n132 0.388379
R19658 vdd.n126 vdd.n125 0.388379
R19659 vdd.n92 vdd.n90 0.388379
R19660 vdd.n67 vdd.n66 0.388379
R19661 vdd.n33 vdd.n31 0.388379
R19662 vdd.n1748 vdd.n1747 0.388379
R19663 vdd.n1714 vdd.n1712 0.388379
R19664 vdd.n1807 vdd.n1806 0.388379
R19665 vdd.n1773 vdd.n1771 0.388379
R19666 vdd.n1646 vdd.n1645 0.388379
R19667 vdd.n1612 vdd.n1610 0.388379
R19668 vdd.n1705 vdd.n1704 0.388379
R19669 vdd.n1671 vdd.n1669 0.388379
R19670 vdd.n1545 vdd.n1544 0.388379
R19671 vdd.n1511 vdd.n1509 0.388379
R19672 vdd.n1604 vdd.n1603 0.388379
R19673 vdd.n1570 vdd.n1568 0.388379
R19674 vdd.n19 vdd.n17 0.387128
R19675 vdd.n24 vdd.n22 0.387128
R19676 vdd.n6 vdd.n4 0.358259
R19677 vdd.n13 vdd.n11 0.358259
R19678 vdd.n276 vdd.n274 0.358259
R19679 vdd.n278 vdd.n276 0.358259
R19680 vdd.n280 vdd.n278 0.358259
R19681 vdd.n282 vdd.n280 0.358259
R19682 vdd.n284 vdd.n282 0.358259
R19683 vdd.n286 vdd.n284 0.358259
R19684 vdd.n288 vdd.n286 0.358259
R19685 vdd.n290 vdd.n288 0.358259
R19686 vdd.n332 vdd.n290 0.358259
R19687 vdd.n174 vdd.n172 0.358259
R19688 vdd.n176 vdd.n174 0.358259
R19689 vdd.n178 vdd.n176 0.358259
R19690 vdd.n180 vdd.n178 0.358259
R19691 vdd.n182 vdd.n180 0.358259
R19692 vdd.n184 vdd.n182 0.358259
R19693 vdd.n186 vdd.n184 0.358259
R19694 vdd.n188 vdd.n186 0.358259
R19695 vdd.n230 vdd.n188 0.358259
R19696 vdd.n73 vdd.n71 0.358259
R19697 vdd.n75 vdd.n73 0.358259
R19698 vdd.n77 vdd.n75 0.358259
R19699 vdd.n79 vdd.n77 0.358259
R19700 vdd.n81 vdd.n79 0.358259
R19701 vdd.n83 vdd.n81 0.358259
R19702 vdd.n85 vdd.n83 0.358259
R19703 vdd.n87 vdd.n85 0.358259
R19704 vdd.n129 vdd.n87 0.358259
R19705 vdd.n1810 vdd.n1768 0.358259
R19706 vdd.n1768 vdd.n1766 0.358259
R19707 vdd.n1766 vdd.n1764 0.358259
R19708 vdd.n1764 vdd.n1762 0.358259
R19709 vdd.n1762 vdd.n1760 0.358259
R19710 vdd.n1760 vdd.n1758 0.358259
R19711 vdd.n1758 vdd.n1756 0.358259
R19712 vdd.n1756 vdd.n1754 0.358259
R19713 vdd.n1754 vdd.n1752 0.358259
R19714 vdd.n1708 vdd.n1666 0.358259
R19715 vdd.n1666 vdd.n1664 0.358259
R19716 vdd.n1664 vdd.n1662 0.358259
R19717 vdd.n1662 vdd.n1660 0.358259
R19718 vdd.n1660 vdd.n1658 0.358259
R19719 vdd.n1658 vdd.n1656 0.358259
R19720 vdd.n1656 vdd.n1654 0.358259
R19721 vdd.n1654 vdd.n1652 0.358259
R19722 vdd.n1652 vdd.n1650 0.358259
R19723 vdd.n1607 vdd.n1565 0.358259
R19724 vdd.n1565 vdd.n1563 0.358259
R19725 vdd.n1563 vdd.n1561 0.358259
R19726 vdd.n1561 vdd.n1559 0.358259
R19727 vdd.n1559 vdd.n1557 0.358259
R19728 vdd.n1557 vdd.n1555 0.358259
R19729 vdd.n1555 vdd.n1553 0.358259
R19730 vdd.n1553 vdd.n1551 0.358259
R19731 vdd.n1551 vdd.n1549 0.358259
R19732 vdd.n14 vdd.n6 0.334552
R19733 vdd.n14 vdd.n13 0.334552
R19734 vdd.n27 vdd.n19 0.21707
R19735 vdd.n27 vdd.n24 0.21707
R19736 vdd.n330 vdd.n292 0.155672
R19737 vdd.n322 vdd.n292 0.155672
R19738 vdd.n322 vdd.n321 0.155672
R19739 vdd.n321 vdd.n297 0.155672
R19740 vdd.n314 vdd.n297 0.155672
R19741 vdd.n314 vdd.n313 0.155672
R19742 vdd.n313 vdd.n301 0.155672
R19743 vdd.n306 vdd.n301 0.155672
R19744 vdd.n271 vdd.n233 0.155672
R19745 vdd.n263 vdd.n233 0.155672
R19746 vdd.n263 vdd.n262 0.155672
R19747 vdd.n262 vdd.n238 0.155672
R19748 vdd.n255 vdd.n238 0.155672
R19749 vdd.n255 vdd.n254 0.155672
R19750 vdd.n254 vdd.n242 0.155672
R19751 vdd.n247 vdd.n242 0.155672
R19752 vdd.n228 vdd.n190 0.155672
R19753 vdd.n220 vdd.n190 0.155672
R19754 vdd.n220 vdd.n219 0.155672
R19755 vdd.n219 vdd.n195 0.155672
R19756 vdd.n212 vdd.n195 0.155672
R19757 vdd.n212 vdd.n211 0.155672
R19758 vdd.n211 vdd.n199 0.155672
R19759 vdd.n204 vdd.n199 0.155672
R19760 vdd.n169 vdd.n131 0.155672
R19761 vdd.n161 vdd.n131 0.155672
R19762 vdd.n161 vdd.n160 0.155672
R19763 vdd.n160 vdd.n136 0.155672
R19764 vdd.n153 vdd.n136 0.155672
R19765 vdd.n153 vdd.n152 0.155672
R19766 vdd.n152 vdd.n140 0.155672
R19767 vdd.n145 vdd.n140 0.155672
R19768 vdd.n127 vdd.n89 0.155672
R19769 vdd.n119 vdd.n89 0.155672
R19770 vdd.n119 vdd.n118 0.155672
R19771 vdd.n118 vdd.n94 0.155672
R19772 vdd.n111 vdd.n94 0.155672
R19773 vdd.n111 vdd.n110 0.155672
R19774 vdd.n110 vdd.n98 0.155672
R19775 vdd.n103 vdd.n98 0.155672
R19776 vdd.n68 vdd.n30 0.155672
R19777 vdd.n60 vdd.n30 0.155672
R19778 vdd.n60 vdd.n59 0.155672
R19779 vdd.n59 vdd.n35 0.155672
R19780 vdd.n52 vdd.n35 0.155672
R19781 vdd.n52 vdd.n51 0.155672
R19782 vdd.n51 vdd.n39 0.155672
R19783 vdd.n44 vdd.n39 0.155672
R19784 vdd.n1749 vdd.n1711 0.155672
R19785 vdd.n1741 vdd.n1711 0.155672
R19786 vdd.n1741 vdd.n1740 0.155672
R19787 vdd.n1740 vdd.n1716 0.155672
R19788 vdd.n1733 vdd.n1716 0.155672
R19789 vdd.n1733 vdd.n1732 0.155672
R19790 vdd.n1732 vdd.n1720 0.155672
R19791 vdd.n1725 vdd.n1720 0.155672
R19792 vdd.n1808 vdd.n1770 0.155672
R19793 vdd.n1800 vdd.n1770 0.155672
R19794 vdd.n1800 vdd.n1799 0.155672
R19795 vdd.n1799 vdd.n1775 0.155672
R19796 vdd.n1792 vdd.n1775 0.155672
R19797 vdd.n1792 vdd.n1791 0.155672
R19798 vdd.n1791 vdd.n1779 0.155672
R19799 vdd.n1784 vdd.n1779 0.155672
R19800 vdd.n1647 vdd.n1609 0.155672
R19801 vdd.n1639 vdd.n1609 0.155672
R19802 vdd.n1639 vdd.n1638 0.155672
R19803 vdd.n1638 vdd.n1614 0.155672
R19804 vdd.n1631 vdd.n1614 0.155672
R19805 vdd.n1631 vdd.n1630 0.155672
R19806 vdd.n1630 vdd.n1618 0.155672
R19807 vdd.n1623 vdd.n1618 0.155672
R19808 vdd.n1706 vdd.n1668 0.155672
R19809 vdd.n1698 vdd.n1668 0.155672
R19810 vdd.n1698 vdd.n1697 0.155672
R19811 vdd.n1697 vdd.n1673 0.155672
R19812 vdd.n1690 vdd.n1673 0.155672
R19813 vdd.n1690 vdd.n1689 0.155672
R19814 vdd.n1689 vdd.n1677 0.155672
R19815 vdd.n1682 vdd.n1677 0.155672
R19816 vdd.n1546 vdd.n1508 0.155672
R19817 vdd.n1538 vdd.n1508 0.155672
R19818 vdd.n1538 vdd.n1537 0.155672
R19819 vdd.n1537 vdd.n1513 0.155672
R19820 vdd.n1530 vdd.n1513 0.155672
R19821 vdd.n1530 vdd.n1529 0.155672
R19822 vdd.n1529 vdd.n1517 0.155672
R19823 vdd.n1522 vdd.n1517 0.155672
R19824 vdd.n1605 vdd.n1567 0.155672
R19825 vdd.n1597 vdd.n1567 0.155672
R19826 vdd.n1597 vdd.n1596 0.155672
R19827 vdd.n1596 vdd.n1572 0.155672
R19828 vdd.n1589 vdd.n1572 0.155672
R19829 vdd.n1589 vdd.n1588 0.155672
R19830 vdd.n1588 vdd.n1576 0.155672
R19831 vdd.n1581 vdd.n1576 0.155672
R19832 vdd.n2101 vdd.n1906 0.152939
R19833 vdd.n1912 vdd.n1906 0.152939
R19834 vdd.n1913 vdd.n1912 0.152939
R19835 vdd.n1914 vdd.n1913 0.152939
R19836 vdd.n1915 vdd.n1914 0.152939
R19837 vdd.n1919 vdd.n1915 0.152939
R19838 vdd.n1920 vdd.n1919 0.152939
R19839 vdd.n1921 vdd.n1920 0.152939
R19840 vdd.n1922 vdd.n1921 0.152939
R19841 vdd.n1926 vdd.n1922 0.152939
R19842 vdd.n1927 vdd.n1926 0.152939
R19843 vdd.n1928 vdd.n1927 0.152939
R19844 vdd.n2076 vdd.n1928 0.152939
R19845 vdd.n2076 vdd.n2075 0.152939
R19846 vdd.n2075 vdd.n2074 0.152939
R19847 vdd.n2074 vdd.n1934 0.152939
R19848 vdd.n1939 vdd.n1934 0.152939
R19849 vdd.n1940 vdd.n1939 0.152939
R19850 vdd.n1941 vdd.n1940 0.152939
R19851 vdd.n1945 vdd.n1941 0.152939
R19852 vdd.n1946 vdd.n1945 0.152939
R19853 vdd.n1947 vdd.n1946 0.152939
R19854 vdd.n1948 vdd.n1947 0.152939
R19855 vdd.n1952 vdd.n1948 0.152939
R19856 vdd.n1953 vdd.n1952 0.152939
R19857 vdd.n1954 vdd.n1953 0.152939
R19858 vdd.n1955 vdd.n1954 0.152939
R19859 vdd.n1959 vdd.n1955 0.152939
R19860 vdd.n1960 vdd.n1959 0.152939
R19861 vdd.n1961 vdd.n1960 0.152939
R19862 vdd.n1962 vdd.n1961 0.152939
R19863 vdd.n1966 vdd.n1962 0.152939
R19864 vdd.n1967 vdd.n1966 0.152939
R19865 vdd.n1968 vdd.n1967 0.152939
R19866 vdd.n2037 vdd.n1968 0.152939
R19867 vdd.n2037 vdd.n2036 0.152939
R19868 vdd.n2036 vdd.n2035 0.152939
R19869 vdd.n2035 vdd.n1974 0.152939
R19870 vdd.n1979 vdd.n1974 0.152939
R19871 vdd.n1980 vdd.n1979 0.152939
R19872 vdd.n1981 vdd.n1980 0.152939
R19873 vdd.n1985 vdd.n1981 0.152939
R19874 vdd.n1986 vdd.n1985 0.152939
R19875 vdd.n1987 vdd.n1986 0.152939
R19876 vdd.n1988 vdd.n1987 0.152939
R19877 vdd.n1992 vdd.n1988 0.152939
R19878 vdd.n1993 vdd.n1992 0.152939
R19879 vdd.n1994 vdd.n1993 0.152939
R19880 vdd.n1995 vdd.n1994 0.152939
R19881 vdd.n1996 vdd.n1995 0.152939
R19882 vdd.n1996 vdd.n1064 0.152939
R19883 vdd.n2325 vdd.n1900 0.152939
R19884 vdd.n1814 vdd.n1123 0.152939
R19885 vdd.n1829 vdd.n1123 0.152939
R19886 vdd.n1830 vdd.n1829 0.152939
R19887 vdd.n1831 vdd.n1830 0.152939
R19888 vdd.n1831 vdd.n1112 0.152939
R19889 vdd.n1846 vdd.n1112 0.152939
R19890 vdd.n1847 vdd.n1846 0.152939
R19891 vdd.n1848 vdd.n1847 0.152939
R19892 vdd.n1848 vdd.n1101 0.152939
R19893 vdd.n1862 vdd.n1101 0.152939
R19894 vdd.n1863 vdd.n1862 0.152939
R19895 vdd.n1864 vdd.n1863 0.152939
R19896 vdd.n1864 vdd.n1089 0.152939
R19897 vdd.n1879 vdd.n1089 0.152939
R19898 vdd.n1880 vdd.n1879 0.152939
R19899 vdd.n1881 vdd.n1880 0.152939
R19900 vdd.n1881 vdd.n1077 0.152939
R19901 vdd.n1898 vdd.n1077 0.152939
R19902 vdd.n1899 vdd.n1898 0.152939
R19903 vdd.n2326 vdd.n1899 0.152939
R19904 vdd.n735 vdd.n730 0.152939
R19905 vdd.n736 vdd.n735 0.152939
R19906 vdd.n737 vdd.n736 0.152939
R19907 vdd.n738 vdd.n737 0.152939
R19908 vdd.n739 vdd.n738 0.152939
R19909 vdd.n740 vdd.n739 0.152939
R19910 vdd.n741 vdd.n740 0.152939
R19911 vdd.n742 vdd.n741 0.152939
R19912 vdd.n743 vdd.n742 0.152939
R19913 vdd.n744 vdd.n743 0.152939
R19914 vdd.n745 vdd.n744 0.152939
R19915 vdd.n746 vdd.n745 0.152939
R19916 vdd.n3183 vdd.n746 0.152939
R19917 vdd.n3183 vdd.n3182 0.152939
R19918 vdd.n3182 vdd.n3181 0.152939
R19919 vdd.n3181 vdd.n748 0.152939
R19920 vdd.n749 vdd.n748 0.152939
R19921 vdd.n750 vdd.n749 0.152939
R19922 vdd.n751 vdd.n750 0.152939
R19923 vdd.n752 vdd.n751 0.152939
R19924 vdd.n753 vdd.n752 0.152939
R19925 vdd.n754 vdd.n753 0.152939
R19926 vdd.n755 vdd.n754 0.152939
R19927 vdd.n756 vdd.n755 0.152939
R19928 vdd.n757 vdd.n756 0.152939
R19929 vdd.n758 vdd.n757 0.152939
R19930 vdd.n759 vdd.n758 0.152939
R19931 vdd.n760 vdd.n759 0.152939
R19932 vdd.n761 vdd.n760 0.152939
R19933 vdd.n762 vdd.n761 0.152939
R19934 vdd.n763 vdd.n762 0.152939
R19935 vdd.n764 vdd.n763 0.152939
R19936 vdd.n765 vdd.n764 0.152939
R19937 vdd.n766 vdd.n765 0.152939
R19938 vdd.n3137 vdd.n766 0.152939
R19939 vdd.n3137 vdd.n3136 0.152939
R19940 vdd.n3136 vdd.n3135 0.152939
R19941 vdd.n3135 vdd.n770 0.152939
R19942 vdd.n771 vdd.n770 0.152939
R19943 vdd.n772 vdd.n771 0.152939
R19944 vdd.n773 vdd.n772 0.152939
R19945 vdd.n774 vdd.n773 0.152939
R19946 vdd.n775 vdd.n774 0.152939
R19947 vdd.n776 vdd.n775 0.152939
R19948 vdd.n777 vdd.n776 0.152939
R19949 vdd.n778 vdd.n777 0.152939
R19950 vdd.n779 vdd.n778 0.152939
R19951 vdd.n780 vdd.n779 0.152939
R19952 vdd.n781 vdd.n780 0.152939
R19953 vdd.n782 vdd.n781 0.152939
R19954 vdd.n783 vdd.n782 0.152939
R19955 vdd.n727 vdd.n726 0.152939
R19956 vdd.n3234 vdd.n682 0.152939
R19957 vdd.n3235 vdd.n3234 0.152939
R19958 vdd.n3236 vdd.n3235 0.152939
R19959 vdd.n3236 vdd.n670 0.152939
R19960 vdd.n3251 vdd.n670 0.152939
R19961 vdd.n3252 vdd.n3251 0.152939
R19962 vdd.n3253 vdd.n3252 0.152939
R19963 vdd.n3253 vdd.n659 0.152939
R19964 vdd.n3267 vdd.n659 0.152939
R19965 vdd.n3268 vdd.n3267 0.152939
R19966 vdd.n3269 vdd.n3268 0.152939
R19967 vdd.n3269 vdd.n647 0.152939
R19968 vdd.n3284 vdd.n647 0.152939
R19969 vdd.n3285 vdd.n3284 0.152939
R19970 vdd.n3286 vdd.n3285 0.152939
R19971 vdd.n3286 vdd.n636 0.152939
R19972 vdd.n3303 vdd.n636 0.152939
R19973 vdd.n3304 vdd.n3303 0.152939
R19974 vdd.n3305 vdd.n3304 0.152939
R19975 vdd.n3305 vdd.n334 0.152939
R19976 vdd.n3398 vdd.n335 0.152939
R19977 vdd.n346 vdd.n335 0.152939
R19978 vdd.n347 vdd.n346 0.152939
R19979 vdd.n348 vdd.n347 0.152939
R19980 vdd.n355 vdd.n348 0.152939
R19981 vdd.n356 vdd.n355 0.152939
R19982 vdd.n357 vdd.n356 0.152939
R19983 vdd.n358 vdd.n357 0.152939
R19984 vdd.n366 vdd.n358 0.152939
R19985 vdd.n367 vdd.n366 0.152939
R19986 vdd.n368 vdd.n367 0.152939
R19987 vdd.n369 vdd.n368 0.152939
R19988 vdd.n377 vdd.n369 0.152939
R19989 vdd.n378 vdd.n377 0.152939
R19990 vdd.n379 vdd.n378 0.152939
R19991 vdd.n380 vdd.n379 0.152939
R19992 vdd.n388 vdd.n380 0.152939
R19993 vdd.n389 vdd.n388 0.152939
R19994 vdd.n390 vdd.n389 0.152939
R19995 vdd.n391 vdd.n390 0.152939
R19996 vdd.n464 vdd.n463 0.152939
R19997 vdd.n470 vdd.n463 0.152939
R19998 vdd.n471 vdd.n470 0.152939
R19999 vdd.n472 vdd.n471 0.152939
R20000 vdd.n472 vdd.n461 0.152939
R20001 vdd.n480 vdd.n461 0.152939
R20002 vdd.n481 vdd.n480 0.152939
R20003 vdd.n482 vdd.n481 0.152939
R20004 vdd.n482 vdd.n459 0.152939
R20005 vdd.n490 vdd.n459 0.152939
R20006 vdd.n491 vdd.n490 0.152939
R20007 vdd.n492 vdd.n491 0.152939
R20008 vdd.n492 vdd.n457 0.152939
R20009 vdd.n500 vdd.n457 0.152939
R20010 vdd.n501 vdd.n500 0.152939
R20011 vdd.n502 vdd.n501 0.152939
R20012 vdd.n502 vdd.n455 0.152939
R20013 vdd.n510 vdd.n455 0.152939
R20014 vdd.n511 vdd.n510 0.152939
R20015 vdd.n512 vdd.n511 0.152939
R20016 vdd.n512 vdd.n451 0.152939
R20017 vdd.n520 vdd.n451 0.152939
R20018 vdd.n521 vdd.n520 0.152939
R20019 vdd.n522 vdd.n521 0.152939
R20020 vdd.n522 vdd.n449 0.152939
R20021 vdd.n530 vdd.n449 0.152939
R20022 vdd.n531 vdd.n530 0.152939
R20023 vdd.n532 vdd.n531 0.152939
R20024 vdd.n532 vdd.n447 0.152939
R20025 vdd.n540 vdd.n447 0.152939
R20026 vdd.n541 vdd.n540 0.152939
R20027 vdd.n542 vdd.n541 0.152939
R20028 vdd.n542 vdd.n445 0.152939
R20029 vdd.n550 vdd.n445 0.152939
R20030 vdd.n551 vdd.n550 0.152939
R20031 vdd.n552 vdd.n551 0.152939
R20032 vdd.n552 vdd.n443 0.152939
R20033 vdd.n560 vdd.n443 0.152939
R20034 vdd.n561 vdd.n560 0.152939
R20035 vdd.n562 vdd.n561 0.152939
R20036 vdd.n562 vdd.n439 0.152939
R20037 vdd.n570 vdd.n439 0.152939
R20038 vdd.n571 vdd.n570 0.152939
R20039 vdd.n572 vdd.n571 0.152939
R20040 vdd.n572 vdd.n437 0.152939
R20041 vdd.n580 vdd.n437 0.152939
R20042 vdd.n581 vdd.n580 0.152939
R20043 vdd.n582 vdd.n581 0.152939
R20044 vdd.n582 vdd.n435 0.152939
R20045 vdd.n590 vdd.n435 0.152939
R20046 vdd.n591 vdd.n590 0.152939
R20047 vdd.n592 vdd.n591 0.152939
R20048 vdd.n592 vdd.n433 0.152939
R20049 vdd.n600 vdd.n433 0.152939
R20050 vdd.n601 vdd.n600 0.152939
R20051 vdd.n602 vdd.n601 0.152939
R20052 vdd.n602 vdd.n431 0.152939
R20053 vdd.n610 vdd.n431 0.152939
R20054 vdd.n611 vdd.n610 0.152939
R20055 vdd.n612 vdd.n611 0.152939
R20056 vdd.n612 vdd.n429 0.152939
R20057 vdd.n619 vdd.n429 0.152939
R20058 vdd.n3350 vdd.n619 0.152939
R20059 vdd.n3228 vdd.n3227 0.152939
R20060 vdd.n3228 vdd.n675 0.152939
R20061 vdd.n3242 vdd.n675 0.152939
R20062 vdd.n3243 vdd.n3242 0.152939
R20063 vdd.n3244 vdd.n3243 0.152939
R20064 vdd.n3244 vdd.n665 0.152939
R20065 vdd.n3259 vdd.n665 0.152939
R20066 vdd.n3260 vdd.n3259 0.152939
R20067 vdd.n3261 vdd.n3260 0.152939
R20068 vdd.n3261 vdd.n652 0.152939
R20069 vdd.n3275 vdd.n652 0.152939
R20070 vdd.n3276 vdd.n3275 0.152939
R20071 vdd.n3277 vdd.n3276 0.152939
R20072 vdd.n3277 vdd.n641 0.152939
R20073 vdd.n3292 vdd.n641 0.152939
R20074 vdd.n3293 vdd.n3292 0.152939
R20075 vdd.n3294 vdd.n3293 0.152939
R20076 vdd.n3296 vdd.n3294 0.152939
R20077 vdd.n3296 vdd.n3295 0.152939
R20078 vdd.n3295 vdd.n630 0.152939
R20079 vdd.n3313 vdd.n630 0.152939
R20080 vdd.n3314 vdd.n3313 0.152939
R20081 vdd.n3315 vdd.n3314 0.152939
R20082 vdd.n3315 vdd.n628 0.152939
R20083 vdd.n3320 vdd.n628 0.152939
R20084 vdd.n3321 vdd.n3320 0.152939
R20085 vdd.n3322 vdd.n3321 0.152939
R20086 vdd.n3322 vdd.n626 0.152939
R20087 vdd.n3327 vdd.n626 0.152939
R20088 vdd.n3328 vdd.n3327 0.152939
R20089 vdd.n3329 vdd.n3328 0.152939
R20090 vdd.n3329 vdd.n624 0.152939
R20091 vdd.n3335 vdd.n624 0.152939
R20092 vdd.n3336 vdd.n3335 0.152939
R20093 vdd.n3337 vdd.n3336 0.152939
R20094 vdd.n3337 vdd.n622 0.152939
R20095 vdd.n3342 vdd.n622 0.152939
R20096 vdd.n3343 vdd.n3342 0.152939
R20097 vdd.n3344 vdd.n3343 0.152939
R20098 vdd.n3344 vdd.n620 0.152939
R20099 vdd.n3349 vdd.n620 0.152939
R20100 vdd.n3226 vdd.n687 0.152939
R20101 vdd.n2337 vdd.n1067 0.152939
R20102 vdd.n1430 vdd.n1186 0.152939
R20103 vdd.n1431 vdd.n1430 0.152939
R20104 vdd.n1432 vdd.n1431 0.152939
R20105 vdd.n1432 vdd.n1174 0.152939
R20106 vdd.n1447 vdd.n1174 0.152939
R20107 vdd.n1448 vdd.n1447 0.152939
R20108 vdd.n1449 vdd.n1448 0.152939
R20109 vdd.n1449 vdd.n1164 0.152939
R20110 vdd.n1464 vdd.n1164 0.152939
R20111 vdd.n1465 vdd.n1464 0.152939
R20112 vdd.n1466 vdd.n1465 0.152939
R20113 vdd.n1466 vdd.n1151 0.152939
R20114 vdd.n1480 vdd.n1151 0.152939
R20115 vdd.n1481 vdd.n1480 0.152939
R20116 vdd.n1482 vdd.n1481 0.152939
R20117 vdd.n1482 vdd.n1140 0.152939
R20118 vdd.n1497 vdd.n1140 0.152939
R20119 vdd.n1498 vdd.n1497 0.152939
R20120 vdd.n1499 vdd.n1498 0.152939
R20121 vdd.n1499 vdd.n1129 0.152939
R20122 vdd.n1820 vdd.n1129 0.152939
R20123 vdd.n1821 vdd.n1820 0.152939
R20124 vdd.n1822 vdd.n1821 0.152939
R20125 vdd.n1822 vdd.n1117 0.152939
R20126 vdd.n1837 vdd.n1117 0.152939
R20127 vdd.n1838 vdd.n1837 0.152939
R20128 vdd.n1839 vdd.n1838 0.152939
R20129 vdd.n1839 vdd.n1107 0.152939
R20130 vdd.n1854 vdd.n1107 0.152939
R20131 vdd.n1855 vdd.n1854 0.152939
R20132 vdd.n1856 vdd.n1855 0.152939
R20133 vdd.n1856 vdd.n1094 0.152939
R20134 vdd.n1870 vdd.n1094 0.152939
R20135 vdd.n1871 vdd.n1870 0.152939
R20136 vdd.n1872 vdd.n1871 0.152939
R20137 vdd.n1872 vdd.n1084 0.152939
R20138 vdd.n1887 vdd.n1084 0.152939
R20139 vdd.n1888 vdd.n1887 0.152939
R20140 vdd.n1891 vdd.n1888 0.152939
R20141 vdd.n1891 vdd.n1890 0.152939
R20142 vdd.n1890 vdd.n1889 0.152939
R20143 vdd.n1422 vdd.n1191 0.152939
R20144 vdd.n1415 vdd.n1191 0.152939
R20145 vdd.n1415 vdd.n1414 0.152939
R20146 vdd.n1414 vdd.n1413 0.152939
R20147 vdd.n1413 vdd.n1228 0.152939
R20148 vdd.n1409 vdd.n1228 0.152939
R20149 vdd.n1409 vdd.n1408 0.152939
R20150 vdd.n1408 vdd.n1407 0.152939
R20151 vdd.n1407 vdd.n1234 0.152939
R20152 vdd.n1403 vdd.n1234 0.152939
R20153 vdd.n1403 vdd.n1402 0.152939
R20154 vdd.n1402 vdd.n1401 0.152939
R20155 vdd.n1401 vdd.n1240 0.152939
R20156 vdd.n1397 vdd.n1240 0.152939
R20157 vdd.n1397 vdd.n1396 0.152939
R20158 vdd.n1396 vdd.n1395 0.152939
R20159 vdd.n1395 vdd.n1246 0.152939
R20160 vdd.n1391 vdd.n1246 0.152939
R20161 vdd.n1391 vdd.n1390 0.152939
R20162 vdd.n1390 vdd.n1389 0.152939
R20163 vdd.n1389 vdd.n1254 0.152939
R20164 vdd.n1385 vdd.n1254 0.152939
R20165 vdd.n1385 vdd.n1384 0.152939
R20166 vdd.n1384 vdd.n1383 0.152939
R20167 vdd.n1383 vdd.n1260 0.152939
R20168 vdd.n1379 vdd.n1260 0.152939
R20169 vdd.n1379 vdd.n1378 0.152939
R20170 vdd.n1378 vdd.n1377 0.152939
R20171 vdd.n1377 vdd.n1266 0.152939
R20172 vdd.n1373 vdd.n1266 0.152939
R20173 vdd.n1373 vdd.n1372 0.152939
R20174 vdd.n1372 vdd.n1371 0.152939
R20175 vdd.n1371 vdd.n1272 0.152939
R20176 vdd.n1367 vdd.n1272 0.152939
R20177 vdd.n1367 vdd.n1366 0.152939
R20178 vdd.n1366 vdd.n1365 0.152939
R20179 vdd.n1365 vdd.n1278 0.152939
R20180 vdd.n1361 vdd.n1278 0.152939
R20181 vdd.n1361 vdd.n1360 0.152939
R20182 vdd.n1360 vdd.n1359 0.152939
R20183 vdd.n1359 vdd.n1284 0.152939
R20184 vdd.n1352 vdd.n1284 0.152939
R20185 vdd.n1352 vdd.n1351 0.152939
R20186 vdd.n1351 vdd.n1350 0.152939
R20187 vdd.n1350 vdd.n1289 0.152939
R20188 vdd.n1346 vdd.n1289 0.152939
R20189 vdd.n1346 vdd.n1345 0.152939
R20190 vdd.n1345 vdd.n1344 0.152939
R20191 vdd.n1344 vdd.n1295 0.152939
R20192 vdd.n1340 vdd.n1295 0.152939
R20193 vdd.n1340 vdd.n1339 0.152939
R20194 vdd.n1339 vdd.n1338 0.152939
R20195 vdd.n1338 vdd.n1301 0.152939
R20196 vdd.n1334 vdd.n1301 0.152939
R20197 vdd.n1334 vdd.n1333 0.152939
R20198 vdd.n1333 vdd.n1332 0.152939
R20199 vdd.n1332 vdd.n1307 0.152939
R20200 vdd.n1328 vdd.n1307 0.152939
R20201 vdd.n1328 vdd.n1327 0.152939
R20202 vdd.n1327 vdd.n1326 0.152939
R20203 vdd.n1326 vdd.n1313 0.152939
R20204 vdd.n1322 vdd.n1313 0.152939
R20205 vdd.n1322 vdd.n1321 0.152939
R20206 vdd.n1424 vdd.n1423 0.152939
R20207 vdd.n1424 vdd.n1180 0.152939
R20208 vdd.n1439 vdd.n1180 0.152939
R20209 vdd.n1440 vdd.n1439 0.152939
R20210 vdd.n1441 vdd.n1440 0.152939
R20211 vdd.n1441 vdd.n1169 0.152939
R20212 vdd.n1456 vdd.n1169 0.152939
R20213 vdd.n1457 vdd.n1456 0.152939
R20214 vdd.n1458 vdd.n1457 0.152939
R20215 vdd.n1458 vdd.n1158 0.152939
R20216 vdd.n1472 vdd.n1158 0.152939
R20217 vdd.n1473 vdd.n1472 0.152939
R20218 vdd.n1474 vdd.n1473 0.152939
R20219 vdd.n1474 vdd.n1146 0.152939
R20220 vdd.n1489 vdd.n1146 0.152939
R20221 vdd.n1490 vdd.n1489 0.152939
R20222 vdd.n1491 vdd.n1490 0.152939
R20223 vdd.n1491 vdd.n1135 0.152939
R20224 vdd.n1505 vdd.n1135 0.152939
R20225 vdd.n1506 vdd.n1505 0.152939
R20226 vdd.n1427 vdd.t74 0.113865
R20227 vdd.t81 vdd.n386 0.113865
R20228 vdd.n2315 vdd.n1900 0.110256
R20229 vdd.n3216 vdd.n727 0.110256
R20230 vdd.n3093 vdd.n687 0.110256
R20231 vdd.n2338 vdd.n2337 0.110256
R20232 vdd.n1814 vdd.n1813 0.0695946
R20233 vdd.n3399 vdd.n334 0.0695946
R20234 vdd.n3399 vdd.n3398 0.0695946
R20235 vdd.n1813 vdd.n1506 0.0695946
R20236 vdd.n2315 vdd.n2101 0.0431829
R20237 vdd.n2338 vdd.n1064 0.0431829
R20238 vdd.n3216 vdd.n730 0.0431829
R20239 vdd.n3093 vdd.n783 0.0431829
R20240 vdd vdd.n28 0.00833333
R20241 CSoutput.n19 CSoutput.t206 184.661
R20242 CSoutput.n78 CSoutput.n77 165.8
R20243 CSoutput.n76 CSoutput.n0 165.8
R20244 CSoutput.n75 CSoutput.n74 165.8
R20245 CSoutput.n73 CSoutput.n72 165.8
R20246 CSoutput.n71 CSoutput.n2 165.8
R20247 CSoutput.n69 CSoutput.n68 165.8
R20248 CSoutput.n67 CSoutput.n3 165.8
R20249 CSoutput.n66 CSoutput.n65 165.8
R20250 CSoutput.n63 CSoutput.n4 165.8
R20251 CSoutput.n61 CSoutput.n60 165.8
R20252 CSoutput.n59 CSoutput.n5 165.8
R20253 CSoutput.n58 CSoutput.n57 165.8
R20254 CSoutput.n55 CSoutput.n6 165.8
R20255 CSoutput.n54 CSoutput.n53 165.8
R20256 CSoutput.n52 CSoutput.n51 165.8
R20257 CSoutput.n50 CSoutput.n8 165.8
R20258 CSoutput.n48 CSoutput.n47 165.8
R20259 CSoutput.n46 CSoutput.n9 165.8
R20260 CSoutput.n45 CSoutput.n44 165.8
R20261 CSoutput.n42 CSoutput.n10 165.8
R20262 CSoutput.n41 CSoutput.n40 165.8
R20263 CSoutput.n39 CSoutput.n38 165.8
R20264 CSoutput.n37 CSoutput.n12 165.8
R20265 CSoutput.n35 CSoutput.n34 165.8
R20266 CSoutput.n33 CSoutput.n13 165.8
R20267 CSoutput.n32 CSoutput.n31 165.8
R20268 CSoutput.n29 CSoutput.n14 165.8
R20269 CSoutput.n28 CSoutput.n27 165.8
R20270 CSoutput.n26 CSoutput.n25 165.8
R20271 CSoutput.n24 CSoutput.n16 165.8
R20272 CSoutput.n22 CSoutput.n21 165.8
R20273 CSoutput.n20 CSoutput.n17 165.8
R20274 CSoutput.n77 CSoutput.t208 162.194
R20275 CSoutput.n18 CSoutput.t209 120.501
R20276 CSoutput.n23 CSoutput.t195 120.501
R20277 CSoutput.n15 CSoutput.t192 120.501
R20278 CSoutput.n30 CSoutput.t210 120.501
R20279 CSoutput.n36 CSoutput.t198 120.501
R20280 CSoutput.n11 CSoutput.t200 120.501
R20281 CSoutput.n43 CSoutput.t212 120.501
R20282 CSoutput.n49 CSoutput.t202 120.501
R20283 CSoutput.n7 CSoutput.t204 120.501
R20284 CSoutput.n56 CSoutput.t196 120.501
R20285 CSoutput.n62 CSoutput.t211 120.501
R20286 CSoutput.n64 CSoutput.t205 120.501
R20287 CSoutput.n70 CSoutput.t199 120.501
R20288 CSoutput.n1 CSoutput.t194 120.501
R20289 CSoutput.n330 CSoutput.n328 103.469
R20290 CSoutput.n310 CSoutput.n308 103.469
R20291 CSoutput.n291 CSoutput.n289 103.469
R20292 CSoutput.n120 CSoutput.n118 103.469
R20293 CSoutput.n100 CSoutput.n98 103.469
R20294 CSoutput.n81 CSoutput.n79 103.469
R20295 CSoutput.n344 CSoutput.n343 103.111
R20296 CSoutput.n342 CSoutput.n341 103.111
R20297 CSoutput.n340 CSoutput.n339 103.111
R20298 CSoutput.n338 CSoutput.n337 103.111
R20299 CSoutput.n336 CSoutput.n335 103.111
R20300 CSoutput.n334 CSoutput.n333 103.111
R20301 CSoutput.n332 CSoutput.n331 103.111
R20302 CSoutput.n330 CSoutput.n329 103.111
R20303 CSoutput.n326 CSoutput.n325 103.111
R20304 CSoutput.n324 CSoutput.n323 103.111
R20305 CSoutput.n322 CSoutput.n321 103.111
R20306 CSoutput.n320 CSoutput.n319 103.111
R20307 CSoutput.n318 CSoutput.n317 103.111
R20308 CSoutput.n316 CSoutput.n315 103.111
R20309 CSoutput.n314 CSoutput.n313 103.111
R20310 CSoutput.n312 CSoutput.n311 103.111
R20311 CSoutput.n310 CSoutput.n309 103.111
R20312 CSoutput.n307 CSoutput.n306 103.111
R20313 CSoutput.n305 CSoutput.n304 103.111
R20314 CSoutput.n303 CSoutput.n302 103.111
R20315 CSoutput.n301 CSoutput.n300 103.111
R20316 CSoutput.n299 CSoutput.n298 103.111
R20317 CSoutput.n297 CSoutput.n296 103.111
R20318 CSoutput.n295 CSoutput.n294 103.111
R20319 CSoutput.n293 CSoutput.n292 103.111
R20320 CSoutput.n291 CSoutput.n290 103.111
R20321 CSoutput.n120 CSoutput.n119 103.111
R20322 CSoutput.n122 CSoutput.n121 103.111
R20323 CSoutput.n124 CSoutput.n123 103.111
R20324 CSoutput.n126 CSoutput.n125 103.111
R20325 CSoutput.n128 CSoutput.n127 103.111
R20326 CSoutput.n130 CSoutput.n129 103.111
R20327 CSoutput.n132 CSoutput.n131 103.111
R20328 CSoutput.n134 CSoutput.n133 103.111
R20329 CSoutput.n136 CSoutput.n135 103.111
R20330 CSoutput.n100 CSoutput.n99 103.111
R20331 CSoutput.n102 CSoutput.n101 103.111
R20332 CSoutput.n104 CSoutput.n103 103.111
R20333 CSoutput.n106 CSoutput.n105 103.111
R20334 CSoutput.n108 CSoutput.n107 103.111
R20335 CSoutput.n110 CSoutput.n109 103.111
R20336 CSoutput.n112 CSoutput.n111 103.111
R20337 CSoutput.n114 CSoutput.n113 103.111
R20338 CSoutput.n116 CSoutput.n115 103.111
R20339 CSoutput.n81 CSoutput.n80 103.111
R20340 CSoutput.n83 CSoutput.n82 103.111
R20341 CSoutput.n85 CSoutput.n84 103.111
R20342 CSoutput.n87 CSoutput.n86 103.111
R20343 CSoutput.n89 CSoutput.n88 103.111
R20344 CSoutput.n91 CSoutput.n90 103.111
R20345 CSoutput.n93 CSoutput.n92 103.111
R20346 CSoutput.n95 CSoutput.n94 103.111
R20347 CSoutput.n97 CSoutput.n96 103.111
R20348 CSoutput.n346 CSoutput.n345 103.111
R20349 CSoutput.n374 CSoutput.n372 81.5057
R20350 CSoutput.n362 CSoutput.n360 81.5057
R20351 CSoutput.n351 CSoutput.n349 81.5057
R20352 CSoutput.n410 CSoutput.n408 81.5057
R20353 CSoutput.n398 CSoutput.n396 81.5057
R20354 CSoutput.n387 CSoutput.n385 81.5057
R20355 CSoutput.n382 CSoutput.n381 80.9324
R20356 CSoutput.n380 CSoutput.n379 80.9324
R20357 CSoutput.n378 CSoutput.n377 80.9324
R20358 CSoutput.n376 CSoutput.n375 80.9324
R20359 CSoutput.n374 CSoutput.n373 80.9324
R20360 CSoutput.n370 CSoutput.n369 80.9324
R20361 CSoutput.n368 CSoutput.n367 80.9324
R20362 CSoutput.n366 CSoutput.n365 80.9324
R20363 CSoutput.n364 CSoutput.n363 80.9324
R20364 CSoutput.n362 CSoutput.n361 80.9324
R20365 CSoutput.n359 CSoutput.n358 80.9324
R20366 CSoutput.n357 CSoutput.n356 80.9324
R20367 CSoutput.n355 CSoutput.n354 80.9324
R20368 CSoutput.n353 CSoutput.n352 80.9324
R20369 CSoutput.n351 CSoutput.n350 80.9324
R20370 CSoutput.n410 CSoutput.n409 80.9324
R20371 CSoutput.n412 CSoutput.n411 80.9324
R20372 CSoutput.n414 CSoutput.n413 80.9324
R20373 CSoutput.n416 CSoutput.n415 80.9324
R20374 CSoutput.n418 CSoutput.n417 80.9324
R20375 CSoutput.n398 CSoutput.n397 80.9324
R20376 CSoutput.n400 CSoutput.n399 80.9324
R20377 CSoutput.n402 CSoutput.n401 80.9324
R20378 CSoutput.n404 CSoutput.n403 80.9324
R20379 CSoutput.n406 CSoutput.n405 80.9324
R20380 CSoutput.n387 CSoutput.n386 80.9324
R20381 CSoutput.n389 CSoutput.n388 80.9324
R20382 CSoutput.n391 CSoutput.n390 80.9324
R20383 CSoutput.n393 CSoutput.n392 80.9324
R20384 CSoutput.n395 CSoutput.n394 80.9324
R20385 CSoutput.n25 CSoutput.n24 48.1486
R20386 CSoutput.n69 CSoutput.n3 48.1486
R20387 CSoutput.n38 CSoutput.n37 48.1486
R20388 CSoutput.n42 CSoutput.n41 48.1486
R20389 CSoutput.n51 CSoutput.n50 48.1486
R20390 CSoutput.n55 CSoutput.n54 48.1486
R20391 CSoutput.n22 CSoutput.n17 46.462
R20392 CSoutput.n72 CSoutput.n71 46.462
R20393 CSoutput.n20 CSoutput.n19 44.9055
R20394 CSoutput.n29 CSoutput.n28 43.7635
R20395 CSoutput.n65 CSoutput.n63 43.7635
R20396 CSoutput.n35 CSoutput.n13 41.7396
R20397 CSoutput.n57 CSoutput.n5 41.7396
R20398 CSoutput.n44 CSoutput.n9 37.0171
R20399 CSoutput.n48 CSoutput.n9 37.0171
R20400 CSoutput.n76 CSoutput.n75 34.9932
R20401 CSoutput.n31 CSoutput.n13 32.2947
R20402 CSoutput.n61 CSoutput.n5 32.2947
R20403 CSoutput.n30 CSoutput.n29 29.6014
R20404 CSoutput.n63 CSoutput.n62 29.6014
R20405 CSoutput.n19 CSoutput.n18 28.4085
R20406 CSoutput.n18 CSoutput.n17 25.1176
R20407 CSoutput.n72 CSoutput.n1 25.1176
R20408 CSoutput.n43 CSoutput.n42 22.0922
R20409 CSoutput.n50 CSoutput.n49 22.0922
R20410 CSoutput.n77 CSoutput.n76 21.8586
R20411 CSoutput.n37 CSoutput.n36 18.9681
R20412 CSoutput.n56 CSoutput.n55 18.9681
R20413 CSoutput.n25 CSoutput.n15 17.6292
R20414 CSoutput.n64 CSoutput.n3 17.6292
R20415 CSoutput.n24 CSoutput.n23 15.844
R20416 CSoutput.n70 CSoutput.n69 15.844
R20417 CSoutput.n38 CSoutput.n11 14.5051
R20418 CSoutput.n54 CSoutput.n7 14.5051
R20419 CSoutput.n421 CSoutput.n78 11.4982
R20420 CSoutput.n41 CSoutput.n11 11.3811
R20421 CSoutput.n51 CSoutput.n7 11.3811
R20422 CSoutput.n23 CSoutput.n22 10.0422
R20423 CSoutput.n71 CSoutput.n70 10.0422
R20424 CSoutput.n327 CSoutput.n307 9.25285
R20425 CSoutput.n117 CSoutput.n97 9.25285
R20426 CSoutput.n371 CSoutput.n359 8.98182
R20427 CSoutput.n407 CSoutput.n395 8.98182
R20428 CSoutput.n384 CSoutput.n348 8.61621
R20429 CSoutput.n28 CSoutput.n15 8.25698
R20430 CSoutput.n65 CSoutput.n64 8.25698
R20431 CSoutput.n348 CSoutput.n347 7.12641
R20432 CSoutput.n138 CSoutput.n137 7.12641
R20433 CSoutput.n36 CSoutput.n35 6.91809
R20434 CSoutput.n57 CSoutput.n56 6.91809
R20435 CSoutput.n384 CSoutput.n383 6.02792
R20436 CSoutput.n420 CSoutput.n419 6.02792
R20437 CSoutput.n383 CSoutput.n382 5.25266
R20438 CSoutput.n371 CSoutput.n370 5.25266
R20439 CSoutput.n419 CSoutput.n418 5.25266
R20440 CSoutput.n407 CSoutput.n406 5.25266
R20441 CSoutput.n347 CSoutput.n346 5.1449
R20442 CSoutput.n327 CSoutput.n326 5.1449
R20443 CSoutput.n137 CSoutput.n136 5.1449
R20444 CSoutput.n117 CSoutput.n116 5.1449
R20445 CSoutput.n421 CSoutput.n138 5.02377
R20446 CSoutput.n229 CSoutput.n182 4.5005
R20447 CSoutput.n198 CSoutput.n182 4.5005
R20448 CSoutput.n193 CSoutput.n177 4.5005
R20449 CSoutput.n193 CSoutput.n179 4.5005
R20450 CSoutput.n193 CSoutput.n176 4.5005
R20451 CSoutput.n193 CSoutput.n180 4.5005
R20452 CSoutput.n193 CSoutput.n175 4.5005
R20453 CSoutput.n193 CSoutput.t197 4.5005
R20454 CSoutput.n193 CSoutput.n174 4.5005
R20455 CSoutput.n193 CSoutput.n181 4.5005
R20456 CSoutput.n193 CSoutput.n182 4.5005
R20457 CSoutput.n191 CSoutput.n177 4.5005
R20458 CSoutput.n191 CSoutput.n179 4.5005
R20459 CSoutput.n191 CSoutput.n176 4.5005
R20460 CSoutput.n191 CSoutput.n180 4.5005
R20461 CSoutput.n191 CSoutput.n175 4.5005
R20462 CSoutput.n191 CSoutput.t197 4.5005
R20463 CSoutput.n191 CSoutput.n174 4.5005
R20464 CSoutput.n191 CSoutput.n181 4.5005
R20465 CSoutput.n191 CSoutput.n182 4.5005
R20466 CSoutput.n190 CSoutput.n177 4.5005
R20467 CSoutput.n190 CSoutput.n179 4.5005
R20468 CSoutput.n190 CSoutput.n176 4.5005
R20469 CSoutput.n190 CSoutput.n180 4.5005
R20470 CSoutput.n190 CSoutput.n175 4.5005
R20471 CSoutput.n190 CSoutput.t197 4.5005
R20472 CSoutput.n190 CSoutput.n174 4.5005
R20473 CSoutput.n190 CSoutput.n181 4.5005
R20474 CSoutput.n190 CSoutput.n182 4.5005
R20475 CSoutput.n275 CSoutput.n177 4.5005
R20476 CSoutput.n275 CSoutput.n179 4.5005
R20477 CSoutput.n275 CSoutput.n176 4.5005
R20478 CSoutput.n275 CSoutput.n180 4.5005
R20479 CSoutput.n275 CSoutput.n175 4.5005
R20480 CSoutput.n275 CSoutput.t197 4.5005
R20481 CSoutput.n275 CSoutput.n174 4.5005
R20482 CSoutput.n275 CSoutput.n181 4.5005
R20483 CSoutput.n275 CSoutput.n182 4.5005
R20484 CSoutput.n273 CSoutput.n177 4.5005
R20485 CSoutput.n273 CSoutput.n179 4.5005
R20486 CSoutput.n273 CSoutput.n176 4.5005
R20487 CSoutput.n273 CSoutput.n180 4.5005
R20488 CSoutput.n273 CSoutput.n175 4.5005
R20489 CSoutput.n273 CSoutput.t197 4.5005
R20490 CSoutput.n273 CSoutput.n174 4.5005
R20491 CSoutput.n273 CSoutput.n181 4.5005
R20492 CSoutput.n271 CSoutput.n177 4.5005
R20493 CSoutput.n271 CSoutput.n179 4.5005
R20494 CSoutput.n271 CSoutput.n176 4.5005
R20495 CSoutput.n271 CSoutput.n180 4.5005
R20496 CSoutput.n271 CSoutput.n175 4.5005
R20497 CSoutput.n271 CSoutput.t197 4.5005
R20498 CSoutput.n271 CSoutput.n174 4.5005
R20499 CSoutput.n271 CSoutput.n181 4.5005
R20500 CSoutput.n201 CSoutput.n177 4.5005
R20501 CSoutput.n201 CSoutput.n179 4.5005
R20502 CSoutput.n201 CSoutput.n176 4.5005
R20503 CSoutput.n201 CSoutput.n180 4.5005
R20504 CSoutput.n201 CSoutput.n175 4.5005
R20505 CSoutput.n201 CSoutput.t197 4.5005
R20506 CSoutput.n201 CSoutput.n174 4.5005
R20507 CSoutput.n201 CSoutput.n181 4.5005
R20508 CSoutput.n201 CSoutput.n182 4.5005
R20509 CSoutput.n200 CSoutput.n177 4.5005
R20510 CSoutput.n200 CSoutput.n179 4.5005
R20511 CSoutput.n200 CSoutput.n176 4.5005
R20512 CSoutput.n200 CSoutput.n180 4.5005
R20513 CSoutput.n200 CSoutput.n175 4.5005
R20514 CSoutput.n200 CSoutput.t197 4.5005
R20515 CSoutput.n200 CSoutput.n174 4.5005
R20516 CSoutput.n200 CSoutput.n181 4.5005
R20517 CSoutput.n200 CSoutput.n182 4.5005
R20518 CSoutput.n204 CSoutput.n177 4.5005
R20519 CSoutput.n204 CSoutput.n179 4.5005
R20520 CSoutput.n204 CSoutput.n176 4.5005
R20521 CSoutput.n204 CSoutput.n180 4.5005
R20522 CSoutput.n204 CSoutput.n175 4.5005
R20523 CSoutput.n204 CSoutput.t197 4.5005
R20524 CSoutput.n204 CSoutput.n174 4.5005
R20525 CSoutput.n204 CSoutput.n181 4.5005
R20526 CSoutput.n204 CSoutput.n182 4.5005
R20527 CSoutput.n203 CSoutput.n177 4.5005
R20528 CSoutput.n203 CSoutput.n179 4.5005
R20529 CSoutput.n203 CSoutput.n176 4.5005
R20530 CSoutput.n203 CSoutput.n180 4.5005
R20531 CSoutput.n203 CSoutput.n175 4.5005
R20532 CSoutput.n203 CSoutput.t197 4.5005
R20533 CSoutput.n203 CSoutput.n174 4.5005
R20534 CSoutput.n203 CSoutput.n181 4.5005
R20535 CSoutput.n203 CSoutput.n182 4.5005
R20536 CSoutput.n186 CSoutput.n177 4.5005
R20537 CSoutput.n186 CSoutput.n179 4.5005
R20538 CSoutput.n186 CSoutput.n176 4.5005
R20539 CSoutput.n186 CSoutput.n180 4.5005
R20540 CSoutput.n186 CSoutput.n175 4.5005
R20541 CSoutput.n186 CSoutput.t197 4.5005
R20542 CSoutput.n186 CSoutput.n174 4.5005
R20543 CSoutput.n186 CSoutput.n181 4.5005
R20544 CSoutput.n186 CSoutput.n182 4.5005
R20545 CSoutput.n278 CSoutput.n177 4.5005
R20546 CSoutput.n278 CSoutput.n179 4.5005
R20547 CSoutput.n278 CSoutput.n176 4.5005
R20548 CSoutput.n278 CSoutput.n180 4.5005
R20549 CSoutput.n278 CSoutput.n175 4.5005
R20550 CSoutput.n278 CSoutput.t197 4.5005
R20551 CSoutput.n278 CSoutput.n174 4.5005
R20552 CSoutput.n278 CSoutput.n181 4.5005
R20553 CSoutput.n278 CSoutput.n182 4.5005
R20554 CSoutput.n265 CSoutput.n236 4.5005
R20555 CSoutput.n265 CSoutput.n242 4.5005
R20556 CSoutput.n223 CSoutput.n212 4.5005
R20557 CSoutput.n223 CSoutput.n214 4.5005
R20558 CSoutput.n223 CSoutput.n211 4.5005
R20559 CSoutput.n223 CSoutput.n215 4.5005
R20560 CSoutput.n223 CSoutput.n210 4.5005
R20561 CSoutput.n223 CSoutput.t193 4.5005
R20562 CSoutput.n223 CSoutput.n209 4.5005
R20563 CSoutput.n223 CSoutput.n216 4.5005
R20564 CSoutput.n265 CSoutput.n223 4.5005
R20565 CSoutput.n244 CSoutput.n212 4.5005
R20566 CSoutput.n244 CSoutput.n214 4.5005
R20567 CSoutput.n244 CSoutput.n211 4.5005
R20568 CSoutput.n244 CSoutput.n215 4.5005
R20569 CSoutput.n244 CSoutput.n210 4.5005
R20570 CSoutput.n244 CSoutput.t193 4.5005
R20571 CSoutput.n244 CSoutput.n209 4.5005
R20572 CSoutput.n244 CSoutput.n216 4.5005
R20573 CSoutput.n265 CSoutput.n244 4.5005
R20574 CSoutput.n222 CSoutput.n212 4.5005
R20575 CSoutput.n222 CSoutput.n214 4.5005
R20576 CSoutput.n222 CSoutput.n211 4.5005
R20577 CSoutput.n222 CSoutput.n215 4.5005
R20578 CSoutput.n222 CSoutput.n210 4.5005
R20579 CSoutput.n222 CSoutput.t193 4.5005
R20580 CSoutput.n222 CSoutput.n209 4.5005
R20581 CSoutput.n222 CSoutput.n216 4.5005
R20582 CSoutput.n265 CSoutput.n222 4.5005
R20583 CSoutput.n246 CSoutput.n212 4.5005
R20584 CSoutput.n246 CSoutput.n214 4.5005
R20585 CSoutput.n246 CSoutput.n211 4.5005
R20586 CSoutput.n246 CSoutput.n215 4.5005
R20587 CSoutput.n246 CSoutput.n210 4.5005
R20588 CSoutput.n246 CSoutput.t193 4.5005
R20589 CSoutput.n246 CSoutput.n209 4.5005
R20590 CSoutput.n246 CSoutput.n216 4.5005
R20591 CSoutput.n265 CSoutput.n246 4.5005
R20592 CSoutput.n212 CSoutput.n207 4.5005
R20593 CSoutput.n214 CSoutput.n207 4.5005
R20594 CSoutput.n211 CSoutput.n207 4.5005
R20595 CSoutput.n215 CSoutput.n207 4.5005
R20596 CSoutput.n210 CSoutput.n207 4.5005
R20597 CSoutput.t193 CSoutput.n207 4.5005
R20598 CSoutput.n209 CSoutput.n207 4.5005
R20599 CSoutput.n216 CSoutput.n207 4.5005
R20600 CSoutput.n268 CSoutput.n212 4.5005
R20601 CSoutput.n268 CSoutput.n214 4.5005
R20602 CSoutput.n268 CSoutput.n211 4.5005
R20603 CSoutput.n268 CSoutput.n215 4.5005
R20604 CSoutput.n268 CSoutput.n210 4.5005
R20605 CSoutput.n268 CSoutput.t193 4.5005
R20606 CSoutput.n268 CSoutput.n209 4.5005
R20607 CSoutput.n268 CSoutput.n216 4.5005
R20608 CSoutput.n266 CSoutput.n212 4.5005
R20609 CSoutput.n266 CSoutput.n214 4.5005
R20610 CSoutput.n266 CSoutput.n211 4.5005
R20611 CSoutput.n266 CSoutput.n215 4.5005
R20612 CSoutput.n266 CSoutput.n210 4.5005
R20613 CSoutput.n266 CSoutput.t193 4.5005
R20614 CSoutput.n266 CSoutput.n209 4.5005
R20615 CSoutput.n266 CSoutput.n216 4.5005
R20616 CSoutput.n266 CSoutput.n265 4.5005
R20617 CSoutput.n248 CSoutput.n212 4.5005
R20618 CSoutput.n248 CSoutput.n214 4.5005
R20619 CSoutput.n248 CSoutput.n211 4.5005
R20620 CSoutput.n248 CSoutput.n215 4.5005
R20621 CSoutput.n248 CSoutput.n210 4.5005
R20622 CSoutput.n248 CSoutput.t193 4.5005
R20623 CSoutput.n248 CSoutput.n209 4.5005
R20624 CSoutput.n248 CSoutput.n216 4.5005
R20625 CSoutput.n265 CSoutput.n248 4.5005
R20626 CSoutput.n220 CSoutput.n212 4.5005
R20627 CSoutput.n220 CSoutput.n214 4.5005
R20628 CSoutput.n220 CSoutput.n211 4.5005
R20629 CSoutput.n220 CSoutput.n215 4.5005
R20630 CSoutput.n220 CSoutput.n210 4.5005
R20631 CSoutput.n220 CSoutput.t193 4.5005
R20632 CSoutput.n220 CSoutput.n209 4.5005
R20633 CSoutput.n220 CSoutput.n216 4.5005
R20634 CSoutput.n265 CSoutput.n220 4.5005
R20635 CSoutput.n250 CSoutput.n212 4.5005
R20636 CSoutput.n250 CSoutput.n214 4.5005
R20637 CSoutput.n250 CSoutput.n211 4.5005
R20638 CSoutput.n250 CSoutput.n215 4.5005
R20639 CSoutput.n250 CSoutput.n210 4.5005
R20640 CSoutput.n250 CSoutput.t193 4.5005
R20641 CSoutput.n250 CSoutput.n209 4.5005
R20642 CSoutput.n250 CSoutput.n216 4.5005
R20643 CSoutput.n265 CSoutput.n250 4.5005
R20644 CSoutput.n219 CSoutput.n212 4.5005
R20645 CSoutput.n219 CSoutput.n214 4.5005
R20646 CSoutput.n219 CSoutput.n211 4.5005
R20647 CSoutput.n219 CSoutput.n215 4.5005
R20648 CSoutput.n219 CSoutput.n210 4.5005
R20649 CSoutput.n219 CSoutput.t193 4.5005
R20650 CSoutput.n219 CSoutput.n209 4.5005
R20651 CSoutput.n219 CSoutput.n216 4.5005
R20652 CSoutput.n265 CSoutput.n219 4.5005
R20653 CSoutput.n264 CSoutput.n212 4.5005
R20654 CSoutput.n264 CSoutput.n214 4.5005
R20655 CSoutput.n264 CSoutput.n211 4.5005
R20656 CSoutput.n264 CSoutput.n215 4.5005
R20657 CSoutput.n264 CSoutput.n210 4.5005
R20658 CSoutput.n264 CSoutput.t193 4.5005
R20659 CSoutput.n264 CSoutput.n209 4.5005
R20660 CSoutput.n264 CSoutput.n216 4.5005
R20661 CSoutput.n265 CSoutput.n264 4.5005
R20662 CSoutput.n263 CSoutput.n148 4.5005
R20663 CSoutput.n164 CSoutput.n148 4.5005
R20664 CSoutput.n159 CSoutput.n143 4.5005
R20665 CSoutput.n159 CSoutput.n145 4.5005
R20666 CSoutput.n159 CSoutput.n142 4.5005
R20667 CSoutput.n159 CSoutput.n146 4.5005
R20668 CSoutput.n159 CSoutput.n141 4.5005
R20669 CSoutput.n159 CSoutput.t213 4.5005
R20670 CSoutput.n159 CSoutput.n140 4.5005
R20671 CSoutput.n159 CSoutput.n147 4.5005
R20672 CSoutput.n159 CSoutput.n148 4.5005
R20673 CSoutput.n157 CSoutput.n143 4.5005
R20674 CSoutput.n157 CSoutput.n145 4.5005
R20675 CSoutput.n157 CSoutput.n142 4.5005
R20676 CSoutput.n157 CSoutput.n146 4.5005
R20677 CSoutput.n157 CSoutput.n141 4.5005
R20678 CSoutput.n157 CSoutput.t213 4.5005
R20679 CSoutput.n157 CSoutput.n140 4.5005
R20680 CSoutput.n157 CSoutput.n147 4.5005
R20681 CSoutput.n157 CSoutput.n148 4.5005
R20682 CSoutput.n156 CSoutput.n143 4.5005
R20683 CSoutput.n156 CSoutput.n145 4.5005
R20684 CSoutput.n156 CSoutput.n142 4.5005
R20685 CSoutput.n156 CSoutput.n146 4.5005
R20686 CSoutput.n156 CSoutput.n141 4.5005
R20687 CSoutput.n156 CSoutput.t213 4.5005
R20688 CSoutput.n156 CSoutput.n140 4.5005
R20689 CSoutput.n156 CSoutput.n147 4.5005
R20690 CSoutput.n156 CSoutput.n148 4.5005
R20691 CSoutput.n285 CSoutput.n143 4.5005
R20692 CSoutput.n285 CSoutput.n145 4.5005
R20693 CSoutput.n285 CSoutput.n142 4.5005
R20694 CSoutput.n285 CSoutput.n146 4.5005
R20695 CSoutput.n285 CSoutput.n141 4.5005
R20696 CSoutput.n285 CSoutput.t213 4.5005
R20697 CSoutput.n285 CSoutput.n140 4.5005
R20698 CSoutput.n285 CSoutput.n147 4.5005
R20699 CSoutput.n285 CSoutput.n148 4.5005
R20700 CSoutput.n283 CSoutput.n143 4.5005
R20701 CSoutput.n283 CSoutput.n145 4.5005
R20702 CSoutput.n283 CSoutput.n142 4.5005
R20703 CSoutput.n283 CSoutput.n146 4.5005
R20704 CSoutput.n283 CSoutput.n141 4.5005
R20705 CSoutput.n283 CSoutput.t213 4.5005
R20706 CSoutput.n283 CSoutput.n140 4.5005
R20707 CSoutput.n283 CSoutput.n147 4.5005
R20708 CSoutput.n281 CSoutput.n143 4.5005
R20709 CSoutput.n281 CSoutput.n145 4.5005
R20710 CSoutput.n281 CSoutput.n142 4.5005
R20711 CSoutput.n281 CSoutput.n146 4.5005
R20712 CSoutput.n281 CSoutput.n141 4.5005
R20713 CSoutput.n281 CSoutput.t213 4.5005
R20714 CSoutput.n281 CSoutput.n140 4.5005
R20715 CSoutput.n281 CSoutput.n147 4.5005
R20716 CSoutput.n167 CSoutput.n143 4.5005
R20717 CSoutput.n167 CSoutput.n145 4.5005
R20718 CSoutput.n167 CSoutput.n142 4.5005
R20719 CSoutput.n167 CSoutput.n146 4.5005
R20720 CSoutput.n167 CSoutput.n141 4.5005
R20721 CSoutput.n167 CSoutput.t213 4.5005
R20722 CSoutput.n167 CSoutput.n140 4.5005
R20723 CSoutput.n167 CSoutput.n147 4.5005
R20724 CSoutput.n167 CSoutput.n148 4.5005
R20725 CSoutput.n166 CSoutput.n143 4.5005
R20726 CSoutput.n166 CSoutput.n145 4.5005
R20727 CSoutput.n166 CSoutput.n142 4.5005
R20728 CSoutput.n166 CSoutput.n146 4.5005
R20729 CSoutput.n166 CSoutput.n141 4.5005
R20730 CSoutput.n166 CSoutput.t213 4.5005
R20731 CSoutput.n166 CSoutput.n140 4.5005
R20732 CSoutput.n166 CSoutput.n147 4.5005
R20733 CSoutput.n166 CSoutput.n148 4.5005
R20734 CSoutput.n170 CSoutput.n143 4.5005
R20735 CSoutput.n170 CSoutput.n145 4.5005
R20736 CSoutput.n170 CSoutput.n142 4.5005
R20737 CSoutput.n170 CSoutput.n146 4.5005
R20738 CSoutput.n170 CSoutput.n141 4.5005
R20739 CSoutput.n170 CSoutput.t213 4.5005
R20740 CSoutput.n170 CSoutput.n140 4.5005
R20741 CSoutput.n170 CSoutput.n147 4.5005
R20742 CSoutput.n170 CSoutput.n148 4.5005
R20743 CSoutput.n169 CSoutput.n143 4.5005
R20744 CSoutput.n169 CSoutput.n145 4.5005
R20745 CSoutput.n169 CSoutput.n142 4.5005
R20746 CSoutput.n169 CSoutput.n146 4.5005
R20747 CSoutput.n169 CSoutput.n141 4.5005
R20748 CSoutput.n169 CSoutput.t213 4.5005
R20749 CSoutput.n169 CSoutput.n140 4.5005
R20750 CSoutput.n169 CSoutput.n147 4.5005
R20751 CSoutput.n169 CSoutput.n148 4.5005
R20752 CSoutput.n152 CSoutput.n143 4.5005
R20753 CSoutput.n152 CSoutput.n145 4.5005
R20754 CSoutput.n152 CSoutput.n142 4.5005
R20755 CSoutput.n152 CSoutput.n146 4.5005
R20756 CSoutput.n152 CSoutput.n141 4.5005
R20757 CSoutput.n152 CSoutput.t213 4.5005
R20758 CSoutput.n152 CSoutput.n140 4.5005
R20759 CSoutput.n152 CSoutput.n147 4.5005
R20760 CSoutput.n152 CSoutput.n148 4.5005
R20761 CSoutput.n288 CSoutput.n143 4.5005
R20762 CSoutput.n288 CSoutput.n145 4.5005
R20763 CSoutput.n288 CSoutput.n142 4.5005
R20764 CSoutput.n288 CSoutput.n146 4.5005
R20765 CSoutput.n288 CSoutput.n141 4.5005
R20766 CSoutput.n288 CSoutput.t213 4.5005
R20767 CSoutput.n288 CSoutput.n140 4.5005
R20768 CSoutput.n288 CSoutput.n147 4.5005
R20769 CSoutput.n288 CSoutput.n148 4.5005
R20770 CSoutput.n347 CSoutput.n327 4.10845
R20771 CSoutput.n137 CSoutput.n117 4.10845
R20772 CSoutput.n345 CSoutput.t127 4.06363
R20773 CSoutput.n345 CSoutput.t151 4.06363
R20774 CSoutput.n343 CSoutput.t171 4.06363
R20775 CSoutput.n343 CSoutput.t85 4.06363
R20776 CSoutput.n341 CSoutput.t89 4.06363
R20777 CSoutput.n341 CSoutput.t155 4.06363
R20778 CSoutput.n339 CSoutput.t174 4.06363
R20779 CSoutput.n339 CSoutput.t175 4.06363
R20780 CSoutput.n337 CSoutput.t105 4.06363
R20781 CSoutput.n337 CSoutput.t106 4.06363
R20782 CSoutput.n335 CSoutput.t111 4.06363
R20783 CSoutput.n335 CSoutput.t176 4.06363
R20784 CSoutput.n333 CSoutput.t75 4.06363
R20785 CSoutput.n333 CSoutput.t109 4.06363
R20786 CSoutput.n331 CSoutput.t126 4.06363
R20787 CSoutput.n331 CSoutput.t150 4.06363
R20788 CSoutput.n329 CSoutput.t157 4.06363
R20789 CSoutput.n329 CSoutput.t81 4.06363
R20790 CSoutput.n328 CSoutput.t129 4.06363
R20791 CSoutput.n328 CSoutput.t130 4.06363
R20792 CSoutput.n325 CSoutput.t112 4.06363
R20793 CSoutput.n325 CSoutput.t139 4.06363
R20794 CSoutput.n323 CSoutput.t159 4.06363
R20795 CSoutput.n323 CSoutput.t71 4.06363
R20796 CSoutput.n321 CSoutput.t72 4.06363
R20797 CSoutput.n321 CSoutput.t141 4.06363
R20798 CSoutput.n319 CSoutput.t162 4.06363
R20799 CSoutput.n319 CSoutput.t163 4.06363
R20800 CSoutput.n317 CSoutput.t93 4.06363
R20801 CSoutput.n317 CSoutput.t94 4.06363
R20802 CSoutput.n315 CSoutput.t97 4.06363
R20803 CSoutput.n315 CSoutput.t166 4.06363
R20804 CSoutput.n313 CSoutput.t60 4.06363
R20805 CSoutput.n313 CSoutput.t96 4.06363
R20806 CSoutput.n311 CSoutput.t113 4.06363
R20807 CSoutput.n311 CSoutput.t140 4.06363
R20808 CSoutput.n309 CSoutput.t142 4.06363
R20809 CSoutput.n309 CSoutput.t66 4.06363
R20810 CSoutput.n308 CSoutput.t119 4.06363
R20811 CSoutput.n308 CSoutput.t120 4.06363
R20812 CSoutput.n306 CSoutput.t148 4.06363
R20813 CSoutput.n306 CSoutput.t102 4.06363
R20814 CSoutput.n304 CSoutput.t135 4.06363
R20815 CSoutput.n304 CSoutput.t84 4.06363
R20816 CSoutput.n302 CSoutput.t160 4.06363
R20817 CSoutput.n302 CSoutput.t76 4.06363
R20818 CSoutput.n300 CSoutput.t116 4.06363
R20819 CSoutput.n300 CSoutput.t95 4.06363
R20820 CSoutput.n298 CSoutput.t98 4.06363
R20821 CSoutput.n298 CSoutput.t73 4.06363
R20822 CSoutput.n296 CSoutput.t147 4.06363
R20823 CSoutput.n296 CSoutput.t67 4.06363
R20824 CSoutput.n294 CSoutput.t107 4.06363
R20825 CSoutput.n294 CSoutput.t172 4.06363
R20826 CSoutput.n292 CSoutput.t90 4.06363
R20827 CSoutput.n292 CSoutput.t153 4.06363
R20828 CSoutput.n290 CSoutput.t114 4.06363
R20829 CSoutput.n290 CSoutput.t177 4.06363
R20830 CSoutput.n289 CSoutput.t61 4.06363
R20831 CSoutput.n289 CSoutput.t164 4.06363
R20832 CSoutput.n118 CSoutput.t170 4.06363
R20833 CSoutput.n118 CSoutput.t169 4.06363
R20834 CSoutput.n119 CSoutput.t149 4.06363
R20835 CSoutput.n119 CSoutput.t83 4.06363
R20836 CSoutput.n121 CSoutput.t79 4.06363
R20837 CSoutput.n121 CSoutput.t167 4.06363
R20838 CSoutput.n123 CSoutput.t146 4.06363
R20839 CSoutput.n123 CSoutput.t123 4.06363
R20840 CSoutput.n125 CSoutput.t104 4.06363
R20841 CSoutput.n125 CSoutput.t179 4.06363
R20842 CSoutput.n127 CSoutput.t144 4.06363
R20843 CSoutput.n127 CSoutput.t143 4.06363
R20844 CSoutput.n129 CSoutput.t131 4.06363
R20845 CSoutput.n129 CSoutput.t101 4.06363
R20846 CSoutput.n131 CSoutput.t82 4.06363
R20847 CSoutput.n131 CSoutput.t132 4.06363
R20848 CSoutput.n133 CSoutput.t128 4.06363
R20849 CSoutput.n133 CSoutput.t99 4.06363
R20850 CSoutput.n135 CSoutput.t80 4.06363
R20851 CSoutput.n135 CSoutput.t78 4.06363
R20852 CSoutput.n98 CSoutput.t158 4.06363
R20853 CSoutput.n98 CSoutput.t156 4.06363
R20854 CSoutput.n99 CSoutput.t138 4.06363
R20855 CSoutput.n99 CSoutput.t70 4.06363
R20856 CSoutput.n101 CSoutput.t64 4.06363
R20857 CSoutput.n101 CSoutput.t152 4.06363
R20858 CSoutput.n103 CSoutput.t137 4.06363
R20859 CSoutput.n103 CSoutput.t110 4.06363
R20860 CSoutput.n105 CSoutput.t92 4.06363
R20861 CSoutput.n105 CSoutput.t168 4.06363
R20862 CSoutput.n107 CSoutput.t134 4.06363
R20863 CSoutput.n107 CSoutput.t133 4.06363
R20864 CSoutput.n109 CSoutput.t121 4.06363
R20865 CSoutput.n109 CSoutput.t88 4.06363
R20866 CSoutput.n111 CSoutput.t68 4.06363
R20867 CSoutput.n111 CSoutput.t122 4.06363
R20868 CSoutput.n113 CSoutput.t118 4.06363
R20869 CSoutput.n113 CSoutput.t86 4.06363
R20870 CSoutput.n115 CSoutput.t65 4.06363
R20871 CSoutput.n115 CSoutput.t62 4.06363
R20872 CSoutput.n79 CSoutput.t165 4.06363
R20873 CSoutput.n79 CSoutput.t63 4.06363
R20874 CSoutput.n80 CSoutput.t145 4.06363
R20875 CSoutput.n80 CSoutput.t115 4.06363
R20876 CSoutput.n82 CSoutput.t154 4.06363
R20877 CSoutput.n82 CSoutput.t91 4.06363
R20878 CSoutput.n84 CSoutput.t173 4.06363
R20879 CSoutput.n84 CSoutput.t108 4.06363
R20880 CSoutput.n86 CSoutput.t69 4.06363
R20881 CSoutput.n86 CSoutput.t124 4.06363
R20882 CSoutput.n88 CSoutput.t74 4.06363
R20883 CSoutput.n88 CSoutput.t100 4.06363
R20884 CSoutput.n90 CSoutput.t178 4.06363
R20885 CSoutput.n90 CSoutput.t117 4.06363
R20886 CSoutput.n92 CSoutput.t77 4.06363
R20887 CSoutput.n92 CSoutput.t161 4.06363
R20888 CSoutput.n94 CSoutput.t87 4.06363
R20889 CSoutput.n94 CSoutput.t136 4.06363
R20890 CSoutput.n96 CSoutput.t103 4.06363
R20891 CSoutput.n96 CSoutput.t125 4.06363
R20892 CSoutput.n44 CSoutput.n43 3.79402
R20893 CSoutput.n49 CSoutput.n48 3.79402
R20894 CSoutput.n383 CSoutput.n371 3.72967
R20895 CSoutput.n419 CSoutput.n407 3.72967
R20896 CSoutput.n421 CSoutput.n420 3.57343
R20897 CSoutput.n381 CSoutput.t53 2.82907
R20898 CSoutput.n381 CSoutput.t41 2.82907
R20899 CSoutput.n379 CSoutput.t52 2.82907
R20900 CSoutput.n379 CSoutput.t16 2.82907
R20901 CSoutput.n377 CSoutput.t183 2.82907
R20902 CSoutput.n377 CSoutput.t31 2.82907
R20903 CSoutput.n375 CSoutput.t5 2.82907
R20904 CSoutput.n375 CSoutput.t48 2.82907
R20905 CSoutput.n373 CSoutput.t18 2.82907
R20906 CSoutput.n373 CSoutput.t15 2.82907
R20907 CSoutput.n372 CSoutput.t12 2.82907
R20908 CSoutput.n372 CSoutput.t187 2.82907
R20909 CSoutput.n369 CSoutput.t17 2.82907
R20910 CSoutput.n369 CSoutput.t0 2.82907
R20911 CSoutput.n367 CSoutput.t58 2.82907
R20912 CSoutput.n367 CSoutput.t32 2.82907
R20913 CSoutput.n365 CSoutput.t1 2.82907
R20914 CSoutput.n365 CSoutput.t2 2.82907
R20915 CSoutput.n363 CSoutput.t10 2.82907
R20916 CSoutput.n363 CSoutput.t59 2.82907
R20917 CSoutput.n361 CSoutput.t30 2.82907
R20918 CSoutput.n361 CSoutput.t21 2.82907
R20919 CSoutput.n360 CSoutput.t23 2.82907
R20920 CSoutput.n360 CSoutput.t22 2.82907
R20921 CSoutput.n358 CSoutput.t35 2.82907
R20922 CSoutput.n358 CSoutput.t189 2.82907
R20923 CSoutput.n356 CSoutput.t180 2.82907
R20924 CSoutput.n356 CSoutput.t9 2.82907
R20925 CSoutput.n354 CSoutput.t36 2.82907
R20926 CSoutput.n354 CSoutput.t19 2.82907
R20927 CSoutput.n352 CSoutput.t54 2.82907
R20928 CSoutput.n352 CSoutput.t184 2.82907
R20929 CSoutput.n350 CSoutput.t14 2.82907
R20930 CSoutput.n350 CSoutput.t40 2.82907
R20931 CSoutput.n349 CSoutput.t182 2.82907
R20932 CSoutput.n349 CSoutput.t24 2.82907
R20933 CSoutput.n408 CSoutput.t34 2.82907
R20934 CSoutput.n408 CSoutput.t45 2.82907
R20935 CSoutput.n409 CSoutput.t38 2.82907
R20936 CSoutput.n409 CSoutput.t181 2.82907
R20937 CSoutput.n411 CSoutput.t185 2.82907
R20938 CSoutput.n411 CSoutput.t28 2.82907
R20939 CSoutput.n413 CSoutput.t7 2.82907
R20940 CSoutput.n413 CSoutput.t33 2.82907
R20941 CSoutput.n415 CSoutput.t47 2.82907
R20942 CSoutput.n415 CSoutput.t56 2.82907
R20943 CSoutput.n417 CSoutput.t11 2.82907
R20944 CSoutput.n417 CSoutput.t13 2.82907
R20945 CSoutput.n396 CSoutput.t39 2.82907
R20946 CSoutput.n396 CSoutput.t3 2.82907
R20947 CSoutput.n397 CSoutput.t26 2.82907
R20948 CSoutput.n397 CSoutput.t57 2.82907
R20949 CSoutput.n399 CSoutput.t25 2.82907
R20950 CSoutput.n399 CSoutput.t43 2.82907
R20951 CSoutput.n401 CSoutput.t191 2.82907
R20952 CSoutput.n401 CSoutput.t6 2.82907
R20953 CSoutput.n403 CSoutput.t44 2.82907
R20954 CSoutput.n403 CSoutput.t50 2.82907
R20955 CSoutput.n405 CSoutput.t51 2.82907
R20956 CSoutput.n405 CSoutput.t190 2.82907
R20957 CSoutput.n385 CSoutput.t42 2.82907
R20958 CSoutput.n385 CSoutput.t8 2.82907
R20959 CSoutput.n386 CSoutput.t37 2.82907
R20960 CSoutput.n386 CSoutput.t186 2.82907
R20961 CSoutput.n388 CSoutput.t49 2.82907
R20962 CSoutput.n388 CSoutput.t20 2.82907
R20963 CSoutput.n390 CSoutput.t46 2.82907
R20964 CSoutput.n390 CSoutput.t55 2.82907
R20965 CSoutput.n392 CSoutput.t188 2.82907
R20966 CSoutput.n392 CSoutput.t4 2.82907
R20967 CSoutput.n394 CSoutput.t27 2.82907
R20968 CSoutput.n394 CSoutput.t29 2.82907
R20969 CSoutput.n420 CSoutput.n384 2.75627
R20970 CSoutput.n348 CSoutput.n138 2.57547
R20971 CSoutput.n75 CSoutput.n1 2.45513
R20972 CSoutput.n229 CSoutput.n227 2.251
R20973 CSoutput.n229 CSoutput.n226 2.251
R20974 CSoutput.n229 CSoutput.n225 2.251
R20975 CSoutput.n229 CSoutput.n224 2.251
R20976 CSoutput.n198 CSoutput.n197 2.251
R20977 CSoutput.n198 CSoutput.n196 2.251
R20978 CSoutput.n198 CSoutput.n195 2.251
R20979 CSoutput.n198 CSoutput.n194 2.251
R20980 CSoutput.n271 CSoutput.n270 2.251
R20981 CSoutput.n236 CSoutput.n234 2.251
R20982 CSoutput.n236 CSoutput.n233 2.251
R20983 CSoutput.n236 CSoutput.n232 2.251
R20984 CSoutput.n254 CSoutput.n236 2.251
R20985 CSoutput.n242 CSoutput.n241 2.251
R20986 CSoutput.n242 CSoutput.n240 2.251
R20987 CSoutput.n242 CSoutput.n239 2.251
R20988 CSoutput.n242 CSoutput.n238 2.251
R20989 CSoutput.n268 CSoutput.n208 2.251
R20990 CSoutput.n263 CSoutput.n261 2.251
R20991 CSoutput.n263 CSoutput.n260 2.251
R20992 CSoutput.n263 CSoutput.n259 2.251
R20993 CSoutput.n263 CSoutput.n258 2.251
R20994 CSoutput.n164 CSoutput.n163 2.251
R20995 CSoutput.n164 CSoutput.n162 2.251
R20996 CSoutput.n164 CSoutput.n161 2.251
R20997 CSoutput.n164 CSoutput.n160 2.251
R20998 CSoutput.n281 CSoutput.n280 2.251
R20999 CSoutput.n198 CSoutput.n178 2.2505
R21000 CSoutput.n193 CSoutput.n178 2.2505
R21001 CSoutput.n191 CSoutput.n178 2.2505
R21002 CSoutput.n190 CSoutput.n178 2.2505
R21003 CSoutput.n275 CSoutput.n178 2.2505
R21004 CSoutput.n273 CSoutput.n178 2.2505
R21005 CSoutput.n271 CSoutput.n178 2.2505
R21006 CSoutput.n201 CSoutput.n178 2.2505
R21007 CSoutput.n200 CSoutput.n178 2.2505
R21008 CSoutput.n204 CSoutput.n178 2.2505
R21009 CSoutput.n203 CSoutput.n178 2.2505
R21010 CSoutput.n186 CSoutput.n178 2.2505
R21011 CSoutput.n278 CSoutput.n178 2.2505
R21012 CSoutput.n278 CSoutput.n277 2.2505
R21013 CSoutput.n242 CSoutput.n213 2.2505
R21014 CSoutput.n223 CSoutput.n213 2.2505
R21015 CSoutput.n244 CSoutput.n213 2.2505
R21016 CSoutput.n222 CSoutput.n213 2.2505
R21017 CSoutput.n246 CSoutput.n213 2.2505
R21018 CSoutput.n213 CSoutput.n207 2.2505
R21019 CSoutput.n268 CSoutput.n213 2.2505
R21020 CSoutput.n266 CSoutput.n213 2.2505
R21021 CSoutput.n248 CSoutput.n213 2.2505
R21022 CSoutput.n220 CSoutput.n213 2.2505
R21023 CSoutput.n250 CSoutput.n213 2.2505
R21024 CSoutput.n219 CSoutput.n213 2.2505
R21025 CSoutput.n264 CSoutput.n213 2.2505
R21026 CSoutput.n264 CSoutput.n217 2.2505
R21027 CSoutput.n164 CSoutput.n144 2.2505
R21028 CSoutput.n159 CSoutput.n144 2.2505
R21029 CSoutput.n157 CSoutput.n144 2.2505
R21030 CSoutput.n156 CSoutput.n144 2.2505
R21031 CSoutput.n285 CSoutput.n144 2.2505
R21032 CSoutput.n283 CSoutput.n144 2.2505
R21033 CSoutput.n281 CSoutput.n144 2.2505
R21034 CSoutput.n167 CSoutput.n144 2.2505
R21035 CSoutput.n166 CSoutput.n144 2.2505
R21036 CSoutput.n170 CSoutput.n144 2.2505
R21037 CSoutput.n169 CSoutput.n144 2.2505
R21038 CSoutput.n152 CSoutput.n144 2.2505
R21039 CSoutput.n288 CSoutput.n144 2.2505
R21040 CSoutput.n288 CSoutput.n287 2.2505
R21041 CSoutput.n206 CSoutput.n199 2.25024
R21042 CSoutput.n206 CSoutput.n192 2.25024
R21043 CSoutput.n274 CSoutput.n206 2.25024
R21044 CSoutput.n206 CSoutput.n202 2.25024
R21045 CSoutput.n206 CSoutput.n205 2.25024
R21046 CSoutput.n206 CSoutput.n173 2.25024
R21047 CSoutput.n256 CSoutput.n253 2.25024
R21048 CSoutput.n256 CSoutput.n252 2.25024
R21049 CSoutput.n256 CSoutput.n251 2.25024
R21050 CSoutput.n256 CSoutput.n218 2.25024
R21051 CSoutput.n256 CSoutput.n255 2.25024
R21052 CSoutput.n257 CSoutput.n256 2.25024
R21053 CSoutput.n172 CSoutput.n165 2.25024
R21054 CSoutput.n172 CSoutput.n158 2.25024
R21055 CSoutput.n284 CSoutput.n172 2.25024
R21056 CSoutput.n172 CSoutput.n168 2.25024
R21057 CSoutput.n172 CSoutput.n171 2.25024
R21058 CSoutput.n172 CSoutput.n139 2.25024
R21059 CSoutput.n273 CSoutput.n183 1.50111
R21060 CSoutput.n221 CSoutput.n207 1.50111
R21061 CSoutput.n283 CSoutput.n149 1.50111
R21062 CSoutput.n229 CSoutput.n228 1.501
R21063 CSoutput.n236 CSoutput.n235 1.501
R21064 CSoutput.n263 CSoutput.n262 1.501
R21065 CSoutput.n277 CSoutput.n188 1.12536
R21066 CSoutput.n277 CSoutput.n189 1.12536
R21067 CSoutput.n277 CSoutput.n276 1.12536
R21068 CSoutput.n237 CSoutput.n217 1.12536
R21069 CSoutput.n243 CSoutput.n217 1.12536
R21070 CSoutput.n245 CSoutput.n217 1.12536
R21071 CSoutput.n287 CSoutput.n154 1.12536
R21072 CSoutput.n287 CSoutput.n155 1.12536
R21073 CSoutput.n287 CSoutput.n286 1.12536
R21074 CSoutput.n277 CSoutput.n184 1.12536
R21075 CSoutput.n277 CSoutput.n185 1.12536
R21076 CSoutput.n277 CSoutput.n187 1.12536
R21077 CSoutput.n267 CSoutput.n217 1.12536
R21078 CSoutput.n247 CSoutput.n217 1.12536
R21079 CSoutput.n249 CSoutput.n217 1.12536
R21080 CSoutput.n287 CSoutput.n150 1.12536
R21081 CSoutput.n287 CSoutput.n151 1.12536
R21082 CSoutput.n287 CSoutput.n153 1.12536
R21083 CSoutput.n31 CSoutput.n30 0.669944
R21084 CSoutput.n62 CSoutput.n61 0.669944
R21085 CSoutput.n376 CSoutput.n374 0.573776
R21086 CSoutput.n378 CSoutput.n376 0.573776
R21087 CSoutput.n380 CSoutput.n378 0.573776
R21088 CSoutput.n382 CSoutput.n380 0.573776
R21089 CSoutput.n364 CSoutput.n362 0.573776
R21090 CSoutput.n366 CSoutput.n364 0.573776
R21091 CSoutput.n368 CSoutput.n366 0.573776
R21092 CSoutput.n370 CSoutput.n368 0.573776
R21093 CSoutput.n353 CSoutput.n351 0.573776
R21094 CSoutput.n355 CSoutput.n353 0.573776
R21095 CSoutput.n357 CSoutput.n355 0.573776
R21096 CSoutput.n359 CSoutput.n357 0.573776
R21097 CSoutput.n418 CSoutput.n416 0.573776
R21098 CSoutput.n416 CSoutput.n414 0.573776
R21099 CSoutput.n414 CSoutput.n412 0.573776
R21100 CSoutput.n412 CSoutput.n410 0.573776
R21101 CSoutput.n406 CSoutput.n404 0.573776
R21102 CSoutput.n404 CSoutput.n402 0.573776
R21103 CSoutput.n402 CSoutput.n400 0.573776
R21104 CSoutput.n400 CSoutput.n398 0.573776
R21105 CSoutput.n395 CSoutput.n393 0.573776
R21106 CSoutput.n393 CSoutput.n391 0.573776
R21107 CSoutput.n391 CSoutput.n389 0.573776
R21108 CSoutput.n389 CSoutput.n387 0.573776
R21109 CSoutput.n421 CSoutput.n288 0.53442
R21110 CSoutput.n332 CSoutput.n330 0.358259
R21111 CSoutput.n334 CSoutput.n332 0.358259
R21112 CSoutput.n336 CSoutput.n334 0.358259
R21113 CSoutput.n338 CSoutput.n336 0.358259
R21114 CSoutput.n340 CSoutput.n338 0.358259
R21115 CSoutput.n342 CSoutput.n340 0.358259
R21116 CSoutput.n344 CSoutput.n342 0.358259
R21117 CSoutput.n346 CSoutput.n344 0.358259
R21118 CSoutput.n312 CSoutput.n310 0.358259
R21119 CSoutput.n314 CSoutput.n312 0.358259
R21120 CSoutput.n316 CSoutput.n314 0.358259
R21121 CSoutput.n318 CSoutput.n316 0.358259
R21122 CSoutput.n320 CSoutput.n318 0.358259
R21123 CSoutput.n322 CSoutput.n320 0.358259
R21124 CSoutput.n324 CSoutput.n322 0.358259
R21125 CSoutput.n326 CSoutput.n324 0.358259
R21126 CSoutput.n293 CSoutput.n291 0.358259
R21127 CSoutput.n295 CSoutput.n293 0.358259
R21128 CSoutput.n297 CSoutput.n295 0.358259
R21129 CSoutput.n299 CSoutput.n297 0.358259
R21130 CSoutput.n301 CSoutput.n299 0.358259
R21131 CSoutput.n303 CSoutput.n301 0.358259
R21132 CSoutput.n305 CSoutput.n303 0.358259
R21133 CSoutput.n307 CSoutput.n305 0.358259
R21134 CSoutput.n136 CSoutput.n134 0.358259
R21135 CSoutput.n134 CSoutput.n132 0.358259
R21136 CSoutput.n132 CSoutput.n130 0.358259
R21137 CSoutput.n130 CSoutput.n128 0.358259
R21138 CSoutput.n128 CSoutput.n126 0.358259
R21139 CSoutput.n126 CSoutput.n124 0.358259
R21140 CSoutput.n124 CSoutput.n122 0.358259
R21141 CSoutput.n122 CSoutput.n120 0.358259
R21142 CSoutput.n116 CSoutput.n114 0.358259
R21143 CSoutput.n114 CSoutput.n112 0.358259
R21144 CSoutput.n112 CSoutput.n110 0.358259
R21145 CSoutput.n110 CSoutput.n108 0.358259
R21146 CSoutput.n108 CSoutput.n106 0.358259
R21147 CSoutput.n106 CSoutput.n104 0.358259
R21148 CSoutput.n104 CSoutput.n102 0.358259
R21149 CSoutput.n102 CSoutput.n100 0.358259
R21150 CSoutput.n97 CSoutput.n95 0.358259
R21151 CSoutput.n95 CSoutput.n93 0.358259
R21152 CSoutput.n93 CSoutput.n91 0.358259
R21153 CSoutput.n91 CSoutput.n89 0.358259
R21154 CSoutput.n89 CSoutput.n87 0.358259
R21155 CSoutput.n87 CSoutput.n85 0.358259
R21156 CSoutput.n85 CSoutput.n83 0.358259
R21157 CSoutput.n83 CSoutput.n81 0.358259
R21158 CSoutput.n21 CSoutput.n20 0.169105
R21159 CSoutput.n21 CSoutput.n16 0.169105
R21160 CSoutput.n26 CSoutput.n16 0.169105
R21161 CSoutput.n27 CSoutput.n26 0.169105
R21162 CSoutput.n27 CSoutput.n14 0.169105
R21163 CSoutput.n32 CSoutput.n14 0.169105
R21164 CSoutput.n33 CSoutput.n32 0.169105
R21165 CSoutput.n34 CSoutput.n33 0.169105
R21166 CSoutput.n34 CSoutput.n12 0.169105
R21167 CSoutput.n39 CSoutput.n12 0.169105
R21168 CSoutput.n40 CSoutput.n39 0.169105
R21169 CSoutput.n40 CSoutput.n10 0.169105
R21170 CSoutput.n45 CSoutput.n10 0.169105
R21171 CSoutput.n46 CSoutput.n45 0.169105
R21172 CSoutput.n47 CSoutput.n46 0.169105
R21173 CSoutput.n47 CSoutput.n8 0.169105
R21174 CSoutput.n52 CSoutput.n8 0.169105
R21175 CSoutput.n53 CSoutput.n52 0.169105
R21176 CSoutput.n53 CSoutput.n6 0.169105
R21177 CSoutput.n58 CSoutput.n6 0.169105
R21178 CSoutput.n59 CSoutput.n58 0.169105
R21179 CSoutput.n60 CSoutput.n59 0.169105
R21180 CSoutput.n60 CSoutput.n4 0.169105
R21181 CSoutput.n66 CSoutput.n4 0.169105
R21182 CSoutput.n67 CSoutput.n66 0.169105
R21183 CSoutput.n68 CSoutput.n67 0.169105
R21184 CSoutput.n68 CSoutput.n2 0.169105
R21185 CSoutput.n73 CSoutput.n2 0.169105
R21186 CSoutput.n74 CSoutput.n73 0.169105
R21187 CSoutput.n74 CSoutput.n0 0.169105
R21188 CSoutput.n78 CSoutput.n0 0.169105
R21189 CSoutput.n231 CSoutput.n230 0.0910737
R21190 CSoutput.n282 CSoutput.n279 0.0723685
R21191 CSoutput.n236 CSoutput.n231 0.0522944
R21192 CSoutput.n279 CSoutput.n278 0.0499135
R21193 CSoutput.n230 CSoutput.n229 0.0499135
R21194 CSoutput.n264 CSoutput.n263 0.0464294
R21195 CSoutput.n272 CSoutput.n269 0.0391444
R21196 CSoutput.n231 CSoutput.t203 0.023435
R21197 CSoutput.n279 CSoutput.t201 0.02262
R21198 CSoutput.n230 CSoutput.t207 0.02262
R21199 CSoutput CSoutput.n421 0.0052
R21200 CSoutput.n201 CSoutput.n184 0.00365111
R21201 CSoutput.n204 CSoutput.n185 0.00365111
R21202 CSoutput.n187 CSoutput.n186 0.00365111
R21203 CSoutput.n229 CSoutput.n188 0.00365111
R21204 CSoutput.n193 CSoutput.n189 0.00365111
R21205 CSoutput.n276 CSoutput.n190 0.00365111
R21206 CSoutput.n267 CSoutput.n266 0.00365111
R21207 CSoutput.n247 CSoutput.n220 0.00365111
R21208 CSoutput.n249 CSoutput.n219 0.00365111
R21209 CSoutput.n237 CSoutput.n236 0.00365111
R21210 CSoutput.n243 CSoutput.n223 0.00365111
R21211 CSoutput.n245 CSoutput.n222 0.00365111
R21212 CSoutput.n167 CSoutput.n150 0.00365111
R21213 CSoutput.n170 CSoutput.n151 0.00365111
R21214 CSoutput.n153 CSoutput.n152 0.00365111
R21215 CSoutput.n263 CSoutput.n154 0.00365111
R21216 CSoutput.n159 CSoutput.n155 0.00365111
R21217 CSoutput.n286 CSoutput.n156 0.00365111
R21218 CSoutput.n198 CSoutput.n188 0.00340054
R21219 CSoutput.n191 CSoutput.n189 0.00340054
R21220 CSoutput.n276 CSoutput.n275 0.00340054
R21221 CSoutput.n271 CSoutput.n184 0.00340054
R21222 CSoutput.n200 CSoutput.n185 0.00340054
R21223 CSoutput.n203 CSoutput.n187 0.00340054
R21224 CSoutput.n242 CSoutput.n237 0.00340054
R21225 CSoutput.n244 CSoutput.n243 0.00340054
R21226 CSoutput.n246 CSoutput.n245 0.00340054
R21227 CSoutput.n268 CSoutput.n267 0.00340054
R21228 CSoutput.n248 CSoutput.n247 0.00340054
R21229 CSoutput.n250 CSoutput.n249 0.00340054
R21230 CSoutput.n164 CSoutput.n154 0.00340054
R21231 CSoutput.n157 CSoutput.n155 0.00340054
R21232 CSoutput.n286 CSoutput.n285 0.00340054
R21233 CSoutput.n281 CSoutput.n150 0.00340054
R21234 CSoutput.n166 CSoutput.n151 0.00340054
R21235 CSoutput.n169 CSoutput.n153 0.00340054
R21236 CSoutput.n199 CSoutput.n193 0.00252698
R21237 CSoutput.n192 CSoutput.n190 0.00252698
R21238 CSoutput.n274 CSoutput.n273 0.00252698
R21239 CSoutput.n202 CSoutput.n200 0.00252698
R21240 CSoutput.n205 CSoutput.n203 0.00252698
R21241 CSoutput.n278 CSoutput.n173 0.00252698
R21242 CSoutput.n199 CSoutput.n198 0.00252698
R21243 CSoutput.n192 CSoutput.n191 0.00252698
R21244 CSoutput.n275 CSoutput.n274 0.00252698
R21245 CSoutput.n202 CSoutput.n201 0.00252698
R21246 CSoutput.n205 CSoutput.n204 0.00252698
R21247 CSoutput.n186 CSoutput.n173 0.00252698
R21248 CSoutput.n253 CSoutput.n223 0.00252698
R21249 CSoutput.n252 CSoutput.n222 0.00252698
R21250 CSoutput.n251 CSoutput.n207 0.00252698
R21251 CSoutput.n248 CSoutput.n218 0.00252698
R21252 CSoutput.n255 CSoutput.n250 0.00252698
R21253 CSoutput.n264 CSoutput.n257 0.00252698
R21254 CSoutput.n253 CSoutput.n242 0.00252698
R21255 CSoutput.n252 CSoutput.n244 0.00252698
R21256 CSoutput.n251 CSoutput.n246 0.00252698
R21257 CSoutput.n266 CSoutput.n218 0.00252698
R21258 CSoutput.n255 CSoutput.n220 0.00252698
R21259 CSoutput.n257 CSoutput.n219 0.00252698
R21260 CSoutput.n165 CSoutput.n159 0.00252698
R21261 CSoutput.n158 CSoutput.n156 0.00252698
R21262 CSoutput.n284 CSoutput.n283 0.00252698
R21263 CSoutput.n168 CSoutput.n166 0.00252698
R21264 CSoutput.n171 CSoutput.n169 0.00252698
R21265 CSoutput.n288 CSoutput.n139 0.00252698
R21266 CSoutput.n165 CSoutput.n164 0.00252698
R21267 CSoutput.n158 CSoutput.n157 0.00252698
R21268 CSoutput.n285 CSoutput.n284 0.00252698
R21269 CSoutput.n168 CSoutput.n167 0.00252698
R21270 CSoutput.n171 CSoutput.n170 0.00252698
R21271 CSoutput.n152 CSoutput.n139 0.00252698
R21272 CSoutput.n273 CSoutput.n272 0.0020275
R21273 CSoutput.n272 CSoutput.n271 0.0020275
R21274 CSoutput.n269 CSoutput.n207 0.0020275
R21275 CSoutput.n269 CSoutput.n268 0.0020275
R21276 CSoutput.n283 CSoutput.n282 0.0020275
R21277 CSoutput.n282 CSoutput.n281 0.0020275
R21278 CSoutput.n183 CSoutput.n182 0.00166668
R21279 CSoutput.n265 CSoutput.n221 0.00166668
R21280 CSoutput.n149 CSoutput.n148 0.00166668
R21281 CSoutput.n287 CSoutput.n149 0.00133328
R21282 CSoutput.n221 CSoutput.n217 0.00133328
R21283 CSoutput.n277 CSoutput.n183 0.00133328
R21284 CSoutput.n280 CSoutput.n172 0.001
R21285 CSoutput.n258 CSoutput.n172 0.001
R21286 CSoutput.n160 CSoutput.n140 0.001
R21287 CSoutput.n259 CSoutput.n140 0.001
R21288 CSoutput.n161 CSoutput.n141 0.001
R21289 CSoutput.n260 CSoutput.n141 0.001
R21290 CSoutput.n162 CSoutput.n142 0.001
R21291 CSoutput.n261 CSoutput.n142 0.001
R21292 CSoutput.n163 CSoutput.n143 0.001
R21293 CSoutput.n262 CSoutput.n143 0.001
R21294 CSoutput.n256 CSoutput.n208 0.001
R21295 CSoutput.n256 CSoutput.n254 0.001
R21296 CSoutput.n238 CSoutput.n209 0.001
R21297 CSoutput.n232 CSoutput.n209 0.001
R21298 CSoutput.n239 CSoutput.n210 0.001
R21299 CSoutput.n233 CSoutput.n210 0.001
R21300 CSoutput.n240 CSoutput.n211 0.001
R21301 CSoutput.n234 CSoutput.n211 0.001
R21302 CSoutput.n241 CSoutput.n212 0.001
R21303 CSoutput.n235 CSoutput.n212 0.001
R21304 CSoutput.n270 CSoutput.n206 0.001
R21305 CSoutput.n224 CSoutput.n206 0.001
R21306 CSoutput.n194 CSoutput.n174 0.001
R21307 CSoutput.n225 CSoutput.n174 0.001
R21308 CSoutput.n195 CSoutput.n175 0.001
R21309 CSoutput.n226 CSoutput.n175 0.001
R21310 CSoutput.n196 CSoutput.n176 0.001
R21311 CSoutput.n227 CSoutput.n176 0.001
R21312 CSoutput.n197 CSoutput.n177 0.001
R21313 CSoutput.n228 CSoutput.n177 0.001
R21314 CSoutput.n228 CSoutput.n178 0.001
R21315 CSoutput.n227 CSoutput.n179 0.001
R21316 CSoutput.n226 CSoutput.n180 0.001
R21317 CSoutput.n225 CSoutput.t197 0.001
R21318 CSoutput.n224 CSoutput.n181 0.001
R21319 CSoutput.n197 CSoutput.n179 0.001
R21320 CSoutput.n196 CSoutput.n180 0.001
R21321 CSoutput.n195 CSoutput.t197 0.001
R21322 CSoutput.n194 CSoutput.n181 0.001
R21323 CSoutput.n270 CSoutput.n182 0.001
R21324 CSoutput.n235 CSoutput.n213 0.001
R21325 CSoutput.n234 CSoutput.n214 0.001
R21326 CSoutput.n233 CSoutput.n215 0.001
R21327 CSoutput.n232 CSoutput.t193 0.001
R21328 CSoutput.n254 CSoutput.n216 0.001
R21329 CSoutput.n241 CSoutput.n214 0.001
R21330 CSoutput.n240 CSoutput.n215 0.001
R21331 CSoutput.n239 CSoutput.t193 0.001
R21332 CSoutput.n238 CSoutput.n216 0.001
R21333 CSoutput.n265 CSoutput.n208 0.001
R21334 CSoutput.n262 CSoutput.n144 0.001
R21335 CSoutput.n261 CSoutput.n145 0.001
R21336 CSoutput.n260 CSoutput.n146 0.001
R21337 CSoutput.n259 CSoutput.t213 0.001
R21338 CSoutput.n258 CSoutput.n147 0.001
R21339 CSoutput.n163 CSoutput.n145 0.001
R21340 CSoutput.n162 CSoutput.n146 0.001
R21341 CSoutput.n161 CSoutput.t213 0.001
R21342 CSoutput.n160 CSoutput.n147 0.001
R21343 CSoutput.n280 CSoutput.n148 0.001
R21344 commonsourceibias.n25 commonsourceibias.t22 230.006
R21345 commonsourceibias.n91 commonsourceibias.t73 230.006
R21346 commonsourceibias.n218 commonsourceibias.t98 230.006
R21347 commonsourceibias.n154 commonsourceibias.t70 230.006
R21348 commonsourceibias.n322 commonsourceibias.t40 230.006
R21349 commonsourceibias.n281 commonsourceibias.t111 230.006
R21350 commonsourceibias.n483 commonsourceibias.t113 230.006
R21351 commonsourceibias.n419 commonsourceibias.t52 230.006
R21352 commonsourceibias.n70 commonsourceibias.t8 207.983
R21353 commonsourceibias.n136 commonsourceibias.t89 207.983
R21354 commonsourceibias.n263 commonsourceibias.t109 207.983
R21355 commonsourceibias.n199 commonsourceibias.t54 207.983
R21356 commonsourceibias.n368 commonsourceibias.t26 207.983
R21357 commonsourceibias.n402 commonsourceibias.t69 207.983
R21358 commonsourceibias.n529 commonsourceibias.t63 207.983
R21359 commonsourceibias.n465 commonsourceibias.t112 207.983
R21360 commonsourceibias.n10 commonsourceibias.t38 168.701
R21361 commonsourceibias.n63 commonsourceibias.t0 168.701
R21362 commonsourceibias.n57 commonsourceibias.t6 168.701
R21363 commonsourceibias.n16 commonsourceibias.t44 168.701
R21364 commonsourceibias.n49 commonsourceibias.t12 168.701
R21365 commonsourceibias.n43 commonsourceibias.t20 168.701
R21366 commonsourceibias.n19 commonsourceibias.t2 168.701
R21367 commonsourceibias.n21 commonsourceibias.t10 168.701
R21368 commonsourceibias.n23 commonsourceibias.t34 168.701
R21369 commonsourceibias.n26 commonsourceibias.t16 168.701
R21370 commonsourceibias.n1 commonsourceibias.t51 168.701
R21371 commonsourceibias.n129 commonsourceibias.t95 168.701
R21372 commonsourceibias.n123 commonsourceibias.t90 168.701
R21373 commonsourceibias.n7 commonsourceibias.t101 168.701
R21374 commonsourceibias.n115 commonsourceibias.t86 168.701
R21375 commonsourceibias.n109 commonsourceibias.t77 168.701
R21376 commonsourceibias.n85 commonsourceibias.t94 168.701
R21377 commonsourceibias.n87 commonsourceibias.t87 168.701
R21378 commonsourceibias.n89 commonsourceibias.t58 168.701
R21379 commonsourceibias.n92 commonsourceibias.t80 168.701
R21380 commonsourceibias.n219 commonsourceibias.t102 168.701
R21381 commonsourceibias.n216 commonsourceibias.t48 168.701
R21382 commonsourceibias.n214 commonsourceibias.t103 168.701
R21383 commonsourceibias.n212 commonsourceibias.t108 168.701
R21384 commonsourceibias.n236 commonsourceibias.t88 168.701
R21385 commonsourceibias.n242 commonsourceibias.t68 168.701
R21386 commonsourceibias.n209 commonsourceibias.t115 168.701
R21387 commonsourceibias.n250 commonsourceibias.t93 168.701
R21388 commonsourceibias.n256 commonsourceibias.t96 168.701
R21389 commonsourceibias.n203 commonsourceibias.t57 168.701
R21390 commonsourceibias.n139 commonsourceibias.t119 168.701
R21391 commonsourceibias.n192 commonsourceibias.t110 168.701
R21392 commonsourceibias.n186 commonsourceibias.t60 168.701
R21393 commonsourceibias.n145 commonsourceibias.t117 168.701
R21394 commonsourceibias.n178 commonsourceibias.t65 168.701
R21395 commonsourceibias.n172 commonsourceibias.t59 168.701
R21396 commonsourceibias.n148 commonsourceibias.t118 168.701
R21397 commonsourceibias.n150 commonsourceibias.t71 168.701
R21398 commonsourceibias.n152 commonsourceibias.t83 168.701
R21399 commonsourceibias.n155 commonsourceibias.t116 168.701
R21400 commonsourceibias.n323 commonsourceibias.t32 168.701
R21401 commonsourceibias.n320 commonsourceibias.t42 168.701
R21402 commonsourceibias.n318 commonsourceibias.t28 168.701
R21403 commonsourceibias.n316 commonsourceibias.t18 168.701
R21404 commonsourceibias.n340 commonsourceibias.t36 168.701
R21405 commonsourceibias.n346 commonsourceibias.t30 168.701
R21406 commonsourceibias.n348 commonsourceibias.t4 168.701
R21407 commonsourceibias.n355 commonsourceibias.t24 168.701
R21408 commonsourceibias.n361 commonsourceibias.t14 168.701
R21409 commonsourceibias.n308 commonsourceibias.t46 168.701
R21410 commonsourceibias.n267 commonsourceibias.t99 168.701
R21411 commonsourceibias.n395 commonsourceibias.t84 168.701
R21412 commonsourceibias.n389 commonsourceibias.t72 168.701
R21413 commonsourceibias.n382 commonsourceibias.t92 168.701
R21414 commonsourceibias.n380 commonsourceibias.t66 168.701
R21415 commonsourceibias.n282 commonsourceibias.t64 168.701
R21416 commonsourceibias.n279 commonsourceibias.t104 168.701
R21417 commonsourceibias.n277 commonsourceibias.t67 168.701
R21418 commonsourceibias.n275 commonsourceibias.t79 168.701
R21419 commonsourceibias.n299 commonsourceibias.t56 168.701
R21420 commonsourceibias.n484 commonsourceibias.t97 168.701
R21421 commonsourceibias.n481 commonsourceibias.t78 168.701
R21422 commonsourceibias.n479 commonsourceibias.t53 168.701
R21423 commonsourceibias.n477 commonsourceibias.t62 168.701
R21424 commonsourceibias.n501 commonsourceibias.t82 168.701
R21425 commonsourceibias.n507 commonsourceibias.t85 168.701
R21426 commonsourceibias.n509 commonsourceibias.t76 168.701
R21427 commonsourceibias.n516 commonsourceibias.t100 168.701
R21428 commonsourceibias.n522 commonsourceibias.t91 168.701
R21429 commonsourceibias.n469 commonsourceibias.t81 168.701
R21430 commonsourceibias.n420 commonsourceibias.t61 168.701
R21431 commonsourceibias.n417 commonsourceibias.t75 168.701
R21432 commonsourceibias.n415 commonsourceibias.t55 168.701
R21433 commonsourceibias.n413 commonsourceibias.t105 168.701
R21434 commonsourceibias.n437 commonsourceibias.t74 168.701
R21435 commonsourceibias.n443 commonsourceibias.t49 168.701
R21436 commonsourceibias.n445 commonsourceibias.t106 168.701
R21437 commonsourceibias.n452 commonsourceibias.t114 168.701
R21438 commonsourceibias.n458 commonsourceibias.t50 168.701
R21439 commonsourceibias.n405 commonsourceibias.t107 168.701
R21440 commonsourceibias.n27 commonsourceibias.n24 161.3
R21441 commonsourceibias.n29 commonsourceibias.n28 161.3
R21442 commonsourceibias.n31 commonsourceibias.n30 161.3
R21443 commonsourceibias.n32 commonsourceibias.n22 161.3
R21444 commonsourceibias.n34 commonsourceibias.n33 161.3
R21445 commonsourceibias.n36 commonsourceibias.n35 161.3
R21446 commonsourceibias.n37 commonsourceibias.n20 161.3
R21447 commonsourceibias.n39 commonsourceibias.n38 161.3
R21448 commonsourceibias.n41 commonsourceibias.n40 161.3
R21449 commonsourceibias.n42 commonsourceibias.n18 161.3
R21450 commonsourceibias.n45 commonsourceibias.n44 161.3
R21451 commonsourceibias.n46 commonsourceibias.n17 161.3
R21452 commonsourceibias.n48 commonsourceibias.n47 161.3
R21453 commonsourceibias.n50 commonsourceibias.n15 161.3
R21454 commonsourceibias.n52 commonsourceibias.n51 161.3
R21455 commonsourceibias.n53 commonsourceibias.n14 161.3
R21456 commonsourceibias.n55 commonsourceibias.n54 161.3
R21457 commonsourceibias.n56 commonsourceibias.n13 161.3
R21458 commonsourceibias.n59 commonsourceibias.n58 161.3
R21459 commonsourceibias.n60 commonsourceibias.n12 161.3
R21460 commonsourceibias.n62 commonsourceibias.n61 161.3
R21461 commonsourceibias.n64 commonsourceibias.n11 161.3
R21462 commonsourceibias.n66 commonsourceibias.n65 161.3
R21463 commonsourceibias.n68 commonsourceibias.n67 161.3
R21464 commonsourceibias.n69 commonsourceibias.n9 161.3
R21465 commonsourceibias.n93 commonsourceibias.n90 161.3
R21466 commonsourceibias.n95 commonsourceibias.n94 161.3
R21467 commonsourceibias.n97 commonsourceibias.n96 161.3
R21468 commonsourceibias.n98 commonsourceibias.n88 161.3
R21469 commonsourceibias.n100 commonsourceibias.n99 161.3
R21470 commonsourceibias.n102 commonsourceibias.n101 161.3
R21471 commonsourceibias.n103 commonsourceibias.n86 161.3
R21472 commonsourceibias.n105 commonsourceibias.n104 161.3
R21473 commonsourceibias.n107 commonsourceibias.n106 161.3
R21474 commonsourceibias.n108 commonsourceibias.n84 161.3
R21475 commonsourceibias.n111 commonsourceibias.n110 161.3
R21476 commonsourceibias.n112 commonsourceibias.n8 161.3
R21477 commonsourceibias.n114 commonsourceibias.n113 161.3
R21478 commonsourceibias.n116 commonsourceibias.n6 161.3
R21479 commonsourceibias.n118 commonsourceibias.n117 161.3
R21480 commonsourceibias.n119 commonsourceibias.n5 161.3
R21481 commonsourceibias.n121 commonsourceibias.n120 161.3
R21482 commonsourceibias.n122 commonsourceibias.n4 161.3
R21483 commonsourceibias.n125 commonsourceibias.n124 161.3
R21484 commonsourceibias.n126 commonsourceibias.n3 161.3
R21485 commonsourceibias.n128 commonsourceibias.n127 161.3
R21486 commonsourceibias.n130 commonsourceibias.n2 161.3
R21487 commonsourceibias.n132 commonsourceibias.n131 161.3
R21488 commonsourceibias.n134 commonsourceibias.n133 161.3
R21489 commonsourceibias.n135 commonsourceibias.n0 161.3
R21490 commonsourceibias.n262 commonsourceibias.n202 161.3
R21491 commonsourceibias.n261 commonsourceibias.n260 161.3
R21492 commonsourceibias.n259 commonsourceibias.n258 161.3
R21493 commonsourceibias.n257 commonsourceibias.n204 161.3
R21494 commonsourceibias.n255 commonsourceibias.n254 161.3
R21495 commonsourceibias.n253 commonsourceibias.n205 161.3
R21496 commonsourceibias.n252 commonsourceibias.n251 161.3
R21497 commonsourceibias.n249 commonsourceibias.n206 161.3
R21498 commonsourceibias.n248 commonsourceibias.n247 161.3
R21499 commonsourceibias.n246 commonsourceibias.n207 161.3
R21500 commonsourceibias.n245 commonsourceibias.n244 161.3
R21501 commonsourceibias.n243 commonsourceibias.n208 161.3
R21502 commonsourceibias.n241 commonsourceibias.n240 161.3
R21503 commonsourceibias.n239 commonsourceibias.n210 161.3
R21504 commonsourceibias.n238 commonsourceibias.n237 161.3
R21505 commonsourceibias.n235 commonsourceibias.n211 161.3
R21506 commonsourceibias.n234 commonsourceibias.n233 161.3
R21507 commonsourceibias.n232 commonsourceibias.n231 161.3
R21508 commonsourceibias.n230 commonsourceibias.n213 161.3
R21509 commonsourceibias.n229 commonsourceibias.n228 161.3
R21510 commonsourceibias.n227 commonsourceibias.n226 161.3
R21511 commonsourceibias.n225 commonsourceibias.n215 161.3
R21512 commonsourceibias.n224 commonsourceibias.n223 161.3
R21513 commonsourceibias.n222 commonsourceibias.n221 161.3
R21514 commonsourceibias.n220 commonsourceibias.n217 161.3
R21515 commonsourceibias.n156 commonsourceibias.n153 161.3
R21516 commonsourceibias.n158 commonsourceibias.n157 161.3
R21517 commonsourceibias.n160 commonsourceibias.n159 161.3
R21518 commonsourceibias.n161 commonsourceibias.n151 161.3
R21519 commonsourceibias.n163 commonsourceibias.n162 161.3
R21520 commonsourceibias.n165 commonsourceibias.n164 161.3
R21521 commonsourceibias.n166 commonsourceibias.n149 161.3
R21522 commonsourceibias.n168 commonsourceibias.n167 161.3
R21523 commonsourceibias.n170 commonsourceibias.n169 161.3
R21524 commonsourceibias.n171 commonsourceibias.n147 161.3
R21525 commonsourceibias.n174 commonsourceibias.n173 161.3
R21526 commonsourceibias.n175 commonsourceibias.n146 161.3
R21527 commonsourceibias.n177 commonsourceibias.n176 161.3
R21528 commonsourceibias.n179 commonsourceibias.n144 161.3
R21529 commonsourceibias.n181 commonsourceibias.n180 161.3
R21530 commonsourceibias.n182 commonsourceibias.n143 161.3
R21531 commonsourceibias.n184 commonsourceibias.n183 161.3
R21532 commonsourceibias.n185 commonsourceibias.n142 161.3
R21533 commonsourceibias.n188 commonsourceibias.n187 161.3
R21534 commonsourceibias.n189 commonsourceibias.n141 161.3
R21535 commonsourceibias.n191 commonsourceibias.n190 161.3
R21536 commonsourceibias.n193 commonsourceibias.n140 161.3
R21537 commonsourceibias.n195 commonsourceibias.n194 161.3
R21538 commonsourceibias.n197 commonsourceibias.n196 161.3
R21539 commonsourceibias.n198 commonsourceibias.n138 161.3
R21540 commonsourceibias.n367 commonsourceibias.n307 161.3
R21541 commonsourceibias.n366 commonsourceibias.n365 161.3
R21542 commonsourceibias.n364 commonsourceibias.n363 161.3
R21543 commonsourceibias.n362 commonsourceibias.n309 161.3
R21544 commonsourceibias.n360 commonsourceibias.n359 161.3
R21545 commonsourceibias.n358 commonsourceibias.n310 161.3
R21546 commonsourceibias.n357 commonsourceibias.n356 161.3
R21547 commonsourceibias.n354 commonsourceibias.n311 161.3
R21548 commonsourceibias.n353 commonsourceibias.n352 161.3
R21549 commonsourceibias.n351 commonsourceibias.n312 161.3
R21550 commonsourceibias.n350 commonsourceibias.n349 161.3
R21551 commonsourceibias.n347 commonsourceibias.n313 161.3
R21552 commonsourceibias.n345 commonsourceibias.n344 161.3
R21553 commonsourceibias.n343 commonsourceibias.n314 161.3
R21554 commonsourceibias.n342 commonsourceibias.n341 161.3
R21555 commonsourceibias.n339 commonsourceibias.n315 161.3
R21556 commonsourceibias.n338 commonsourceibias.n337 161.3
R21557 commonsourceibias.n336 commonsourceibias.n335 161.3
R21558 commonsourceibias.n334 commonsourceibias.n317 161.3
R21559 commonsourceibias.n333 commonsourceibias.n332 161.3
R21560 commonsourceibias.n331 commonsourceibias.n330 161.3
R21561 commonsourceibias.n329 commonsourceibias.n319 161.3
R21562 commonsourceibias.n328 commonsourceibias.n327 161.3
R21563 commonsourceibias.n326 commonsourceibias.n325 161.3
R21564 commonsourceibias.n324 commonsourceibias.n321 161.3
R21565 commonsourceibias.n301 commonsourceibias.n300 161.3
R21566 commonsourceibias.n298 commonsourceibias.n274 161.3
R21567 commonsourceibias.n297 commonsourceibias.n296 161.3
R21568 commonsourceibias.n295 commonsourceibias.n294 161.3
R21569 commonsourceibias.n293 commonsourceibias.n276 161.3
R21570 commonsourceibias.n292 commonsourceibias.n291 161.3
R21571 commonsourceibias.n290 commonsourceibias.n289 161.3
R21572 commonsourceibias.n288 commonsourceibias.n278 161.3
R21573 commonsourceibias.n287 commonsourceibias.n286 161.3
R21574 commonsourceibias.n285 commonsourceibias.n284 161.3
R21575 commonsourceibias.n283 commonsourceibias.n280 161.3
R21576 commonsourceibias.n377 commonsourceibias.n273 161.3
R21577 commonsourceibias.n401 commonsourceibias.n266 161.3
R21578 commonsourceibias.n400 commonsourceibias.n399 161.3
R21579 commonsourceibias.n398 commonsourceibias.n397 161.3
R21580 commonsourceibias.n396 commonsourceibias.n268 161.3
R21581 commonsourceibias.n394 commonsourceibias.n393 161.3
R21582 commonsourceibias.n392 commonsourceibias.n269 161.3
R21583 commonsourceibias.n391 commonsourceibias.n390 161.3
R21584 commonsourceibias.n388 commonsourceibias.n270 161.3
R21585 commonsourceibias.n387 commonsourceibias.n386 161.3
R21586 commonsourceibias.n385 commonsourceibias.n271 161.3
R21587 commonsourceibias.n384 commonsourceibias.n383 161.3
R21588 commonsourceibias.n381 commonsourceibias.n272 161.3
R21589 commonsourceibias.n379 commonsourceibias.n378 161.3
R21590 commonsourceibias.n528 commonsourceibias.n468 161.3
R21591 commonsourceibias.n527 commonsourceibias.n526 161.3
R21592 commonsourceibias.n525 commonsourceibias.n524 161.3
R21593 commonsourceibias.n523 commonsourceibias.n470 161.3
R21594 commonsourceibias.n521 commonsourceibias.n520 161.3
R21595 commonsourceibias.n519 commonsourceibias.n471 161.3
R21596 commonsourceibias.n518 commonsourceibias.n517 161.3
R21597 commonsourceibias.n515 commonsourceibias.n472 161.3
R21598 commonsourceibias.n514 commonsourceibias.n513 161.3
R21599 commonsourceibias.n512 commonsourceibias.n473 161.3
R21600 commonsourceibias.n511 commonsourceibias.n510 161.3
R21601 commonsourceibias.n508 commonsourceibias.n474 161.3
R21602 commonsourceibias.n506 commonsourceibias.n505 161.3
R21603 commonsourceibias.n504 commonsourceibias.n475 161.3
R21604 commonsourceibias.n503 commonsourceibias.n502 161.3
R21605 commonsourceibias.n500 commonsourceibias.n476 161.3
R21606 commonsourceibias.n499 commonsourceibias.n498 161.3
R21607 commonsourceibias.n497 commonsourceibias.n496 161.3
R21608 commonsourceibias.n495 commonsourceibias.n478 161.3
R21609 commonsourceibias.n494 commonsourceibias.n493 161.3
R21610 commonsourceibias.n492 commonsourceibias.n491 161.3
R21611 commonsourceibias.n490 commonsourceibias.n480 161.3
R21612 commonsourceibias.n489 commonsourceibias.n488 161.3
R21613 commonsourceibias.n487 commonsourceibias.n486 161.3
R21614 commonsourceibias.n485 commonsourceibias.n482 161.3
R21615 commonsourceibias.n464 commonsourceibias.n404 161.3
R21616 commonsourceibias.n463 commonsourceibias.n462 161.3
R21617 commonsourceibias.n461 commonsourceibias.n460 161.3
R21618 commonsourceibias.n459 commonsourceibias.n406 161.3
R21619 commonsourceibias.n457 commonsourceibias.n456 161.3
R21620 commonsourceibias.n455 commonsourceibias.n407 161.3
R21621 commonsourceibias.n454 commonsourceibias.n453 161.3
R21622 commonsourceibias.n451 commonsourceibias.n408 161.3
R21623 commonsourceibias.n450 commonsourceibias.n449 161.3
R21624 commonsourceibias.n448 commonsourceibias.n409 161.3
R21625 commonsourceibias.n447 commonsourceibias.n446 161.3
R21626 commonsourceibias.n444 commonsourceibias.n410 161.3
R21627 commonsourceibias.n442 commonsourceibias.n441 161.3
R21628 commonsourceibias.n440 commonsourceibias.n411 161.3
R21629 commonsourceibias.n439 commonsourceibias.n438 161.3
R21630 commonsourceibias.n436 commonsourceibias.n412 161.3
R21631 commonsourceibias.n435 commonsourceibias.n434 161.3
R21632 commonsourceibias.n433 commonsourceibias.n432 161.3
R21633 commonsourceibias.n431 commonsourceibias.n414 161.3
R21634 commonsourceibias.n430 commonsourceibias.n429 161.3
R21635 commonsourceibias.n428 commonsourceibias.n427 161.3
R21636 commonsourceibias.n426 commonsourceibias.n416 161.3
R21637 commonsourceibias.n425 commonsourceibias.n424 161.3
R21638 commonsourceibias.n423 commonsourceibias.n422 161.3
R21639 commonsourceibias.n421 commonsourceibias.n418 161.3
R21640 commonsourceibias.n80 commonsourceibias.n78 81.5057
R21641 commonsourceibias.n304 commonsourceibias.n302 81.5057
R21642 commonsourceibias.n80 commonsourceibias.n79 80.9324
R21643 commonsourceibias.n82 commonsourceibias.n81 80.9324
R21644 commonsourceibias.n77 commonsourceibias.n76 80.9324
R21645 commonsourceibias.n75 commonsourceibias.n74 80.9324
R21646 commonsourceibias.n73 commonsourceibias.n72 80.9324
R21647 commonsourceibias.n371 commonsourceibias.n370 80.9324
R21648 commonsourceibias.n373 commonsourceibias.n372 80.9324
R21649 commonsourceibias.n375 commonsourceibias.n374 80.9324
R21650 commonsourceibias.n306 commonsourceibias.n305 80.9324
R21651 commonsourceibias.n304 commonsourceibias.n303 80.9324
R21652 commonsourceibias.n71 commonsourceibias.n70 80.6037
R21653 commonsourceibias.n137 commonsourceibias.n136 80.6037
R21654 commonsourceibias.n264 commonsourceibias.n263 80.6037
R21655 commonsourceibias.n200 commonsourceibias.n199 80.6037
R21656 commonsourceibias.n369 commonsourceibias.n368 80.6037
R21657 commonsourceibias.n403 commonsourceibias.n402 80.6037
R21658 commonsourceibias.n530 commonsourceibias.n529 80.6037
R21659 commonsourceibias.n466 commonsourceibias.n465 80.6037
R21660 commonsourceibias.n65 commonsourceibias.n64 56.5617
R21661 commonsourceibias.n51 commonsourceibias.n50 56.5617
R21662 commonsourceibias.n42 commonsourceibias.n41 56.5617
R21663 commonsourceibias.n28 commonsourceibias.n27 56.5617
R21664 commonsourceibias.n131 commonsourceibias.n130 56.5617
R21665 commonsourceibias.n117 commonsourceibias.n116 56.5617
R21666 commonsourceibias.n108 commonsourceibias.n107 56.5617
R21667 commonsourceibias.n94 commonsourceibias.n93 56.5617
R21668 commonsourceibias.n221 commonsourceibias.n220 56.5617
R21669 commonsourceibias.n235 commonsourceibias.n234 56.5617
R21670 commonsourceibias.n244 commonsourceibias.n243 56.5617
R21671 commonsourceibias.n258 commonsourceibias.n257 56.5617
R21672 commonsourceibias.n194 commonsourceibias.n193 56.5617
R21673 commonsourceibias.n180 commonsourceibias.n179 56.5617
R21674 commonsourceibias.n171 commonsourceibias.n170 56.5617
R21675 commonsourceibias.n157 commonsourceibias.n156 56.5617
R21676 commonsourceibias.n325 commonsourceibias.n324 56.5617
R21677 commonsourceibias.n339 commonsourceibias.n338 56.5617
R21678 commonsourceibias.n349 commonsourceibias.n347 56.5617
R21679 commonsourceibias.n363 commonsourceibias.n362 56.5617
R21680 commonsourceibias.n397 commonsourceibias.n396 56.5617
R21681 commonsourceibias.n383 commonsourceibias.n381 56.5617
R21682 commonsourceibias.n284 commonsourceibias.n283 56.5617
R21683 commonsourceibias.n298 commonsourceibias.n297 56.5617
R21684 commonsourceibias.n486 commonsourceibias.n485 56.5617
R21685 commonsourceibias.n500 commonsourceibias.n499 56.5617
R21686 commonsourceibias.n510 commonsourceibias.n508 56.5617
R21687 commonsourceibias.n524 commonsourceibias.n523 56.5617
R21688 commonsourceibias.n422 commonsourceibias.n421 56.5617
R21689 commonsourceibias.n436 commonsourceibias.n435 56.5617
R21690 commonsourceibias.n446 commonsourceibias.n444 56.5617
R21691 commonsourceibias.n460 commonsourceibias.n459 56.5617
R21692 commonsourceibias.n56 commonsourceibias.n55 56.0773
R21693 commonsourceibias.n37 commonsourceibias.n36 56.0773
R21694 commonsourceibias.n122 commonsourceibias.n121 56.0773
R21695 commonsourceibias.n103 commonsourceibias.n102 56.0773
R21696 commonsourceibias.n230 commonsourceibias.n229 56.0773
R21697 commonsourceibias.n249 commonsourceibias.n248 56.0773
R21698 commonsourceibias.n185 commonsourceibias.n184 56.0773
R21699 commonsourceibias.n166 commonsourceibias.n165 56.0773
R21700 commonsourceibias.n334 commonsourceibias.n333 56.0773
R21701 commonsourceibias.n354 commonsourceibias.n353 56.0773
R21702 commonsourceibias.n388 commonsourceibias.n387 56.0773
R21703 commonsourceibias.n293 commonsourceibias.n292 56.0773
R21704 commonsourceibias.n495 commonsourceibias.n494 56.0773
R21705 commonsourceibias.n515 commonsourceibias.n514 56.0773
R21706 commonsourceibias.n431 commonsourceibias.n430 56.0773
R21707 commonsourceibias.n451 commonsourceibias.n450 56.0773
R21708 commonsourceibias.n70 commonsourceibias.n69 46.0096
R21709 commonsourceibias.n136 commonsourceibias.n135 46.0096
R21710 commonsourceibias.n263 commonsourceibias.n262 46.0096
R21711 commonsourceibias.n199 commonsourceibias.n198 46.0096
R21712 commonsourceibias.n368 commonsourceibias.n367 46.0096
R21713 commonsourceibias.n402 commonsourceibias.n401 46.0096
R21714 commonsourceibias.n529 commonsourceibias.n528 46.0096
R21715 commonsourceibias.n465 commonsourceibias.n464 46.0096
R21716 commonsourceibias.n58 commonsourceibias.n12 41.5458
R21717 commonsourceibias.n33 commonsourceibias.n32 41.5458
R21718 commonsourceibias.n124 commonsourceibias.n3 41.5458
R21719 commonsourceibias.n99 commonsourceibias.n98 41.5458
R21720 commonsourceibias.n226 commonsourceibias.n225 41.5458
R21721 commonsourceibias.n251 commonsourceibias.n205 41.5458
R21722 commonsourceibias.n187 commonsourceibias.n141 41.5458
R21723 commonsourceibias.n162 commonsourceibias.n161 41.5458
R21724 commonsourceibias.n330 commonsourceibias.n329 41.5458
R21725 commonsourceibias.n356 commonsourceibias.n310 41.5458
R21726 commonsourceibias.n390 commonsourceibias.n269 41.5458
R21727 commonsourceibias.n289 commonsourceibias.n288 41.5458
R21728 commonsourceibias.n491 commonsourceibias.n490 41.5458
R21729 commonsourceibias.n517 commonsourceibias.n471 41.5458
R21730 commonsourceibias.n427 commonsourceibias.n426 41.5458
R21731 commonsourceibias.n453 commonsourceibias.n407 41.5458
R21732 commonsourceibias.n48 commonsourceibias.n17 40.577
R21733 commonsourceibias.n44 commonsourceibias.n17 40.577
R21734 commonsourceibias.n114 commonsourceibias.n8 40.577
R21735 commonsourceibias.n110 commonsourceibias.n8 40.577
R21736 commonsourceibias.n237 commonsourceibias.n210 40.577
R21737 commonsourceibias.n241 commonsourceibias.n210 40.577
R21738 commonsourceibias.n177 commonsourceibias.n146 40.577
R21739 commonsourceibias.n173 commonsourceibias.n146 40.577
R21740 commonsourceibias.n341 commonsourceibias.n314 40.577
R21741 commonsourceibias.n345 commonsourceibias.n314 40.577
R21742 commonsourceibias.n379 commonsourceibias.n273 40.577
R21743 commonsourceibias.n300 commonsourceibias.n273 40.577
R21744 commonsourceibias.n502 commonsourceibias.n475 40.577
R21745 commonsourceibias.n506 commonsourceibias.n475 40.577
R21746 commonsourceibias.n438 commonsourceibias.n411 40.577
R21747 commonsourceibias.n442 commonsourceibias.n411 40.577
R21748 commonsourceibias.n62 commonsourceibias.n12 39.6083
R21749 commonsourceibias.n32 commonsourceibias.n31 39.6083
R21750 commonsourceibias.n128 commonsourceibias.n3 39.6083
R21751 commonsourceibias.n98 commonsourceibias.n97 39.6083
R21752 commonsourceibias.n225 commonsourceibias.n224 39.6083
R21753 commonsourceibias.n255 commonsourceibias.n205 39.6083
R21754 commonsourceibias.n191 commonsourceibias.n141 39.6083
R21755 commonsourceibias.n161 commonsourceibias.n160 39.6083
R21756 commonsourceibias.n329 commonsourceibias.n328 39.6083
R21757 commonsourceibias.n360 commonsourceibias.n310 39.6083
R21758 commonsourceibias.n394 commonsourceibias.n269 39.6083
R21759 commonsourceibias.n288 commonsourceibias.n287 39.6083
R21760 commonsourceibias.n490 commonsourceibias.n489 39.6083
R21761 commonsourceibias.n521 commonsourceibias.n471 39.6083
R21762 commonsourceibias.n426 commonsourceibias.n425 39.6083
R21763 commonsourceibias.n457 commonsourceibias.n407 39.6083
R21764 commonsourceibias.n26 commonsourceibias.n25 33.0515
R21765 commonsourceibias.n92 commonsourceibias.n91 33.0515
R21766 commonsourceibias.n155 commonsourceibias.n154 33.0515
R21767 commonsourceibias.n219 commonsourceibias.n218 33.0515
R21768 commonsourceibias.n323 commonsourceibias.n322 33.0515
R21769 commonsourceibias.n282 commonsourceibias.n281 33.0515
R21770 commonsourceibias.n484 commonsourceibias.n483 33.0515
R21771 commonsourceibias.n420 commonsourceibias.n419 33.0515
R21772 commonsourceibias.n25 commonsourceibias.n24 28.5514
R21773 commonsourceibias.n91 commonsourceibias.n90 28.5514
R21774 commonsourceibias.n218 commonsourceibias.n217 28.5514
R21775 commonsourceibias.n154 commonsourceibias.n153 28.5514
R21776 commonsourceibias.n322 commonsourceibias.n321 28.5514
R21777 commonsourceibias.n281 commonsourceibias.n280 28.5514
R21778 commonsourceibias.n483 commonsourceibias.n482 28.5514
R21779 commonsourceibias.n419 commonsourceibias.n418 28.5514
R21780 commonsourceibias.n69 commonsourceibias.n68 26.0455
R21781 commonsourceibias.n135 commonsourceibias.n134 26.0455
R21782 commonsourceibias.n262 commonsourceibias.n261 26.0455
R21783 commonsourceibias.n198 commonsourceibias.n197 26.0455
R21784 commonsourceibias.n367 commonsourceibias.n366 26.0455
R21785 commonsourceibias.n401 commonsourceibias.n400 26.0455
R21786 commonsourceibias.n528 commonsourceibias.n527 26.0455
R21787 commonsourceibias.n464 commonsourceibias.n463 26.0455
R21788 commonsourceibias.n55 commonsourceibias.n14 25.0767
R21789 commonsourceibias.n38 commonsourceibias.n37 25.0767
R21790 commonsourceibias.n121 commonsourceibias.n5 25.0767
R21791 commonsourceibias.n104 commonsourceibias.n103 25.0767
R21792 commonsourceibias.n231 commonsourceibias.n230 25.0767
R21793 commonsourceibias.n248 commonsourceibias.n207 25.0767
R21794 commonsourceibias.n184 commonsourceibias.n143 25.0767
R21795 commonsourceibias.n167 commonsourceibias.n166 25.0767
R21796 commonsourceibias.n335 commonsourceibias.n334 25.0767
R21797 commonsourceibias.n353 commonsourceibias.n312 25.0767
R21798 commonsourceibias.n387 commonsourceibias.n271 25.0767
R21799 commonsourceibias.n294 commonsourceibias.n293 25.0767
R21800 commonsourceibias.n496 commonsourceibias.n495 25.0767
R21801 commonsourceibias.n514 commonsourceibias.n473 25.0767
R21802 commonsourceibias.n432 commonsourceibias.n431 25.0767
R21803 commonsourceibias.n450 commonsourceibias.n409 25.0767
R21804 commonsourceibias.n51 commonsourceibias.n16 24.3464
R21805 commonsourceibias.n41 commonsourceibias.n19 24.3464
R21806 commonsourceibias.n117 commonsourceibias.n7 24.3464
R21807 commonsourceibias.n107 commonsourceibias.n85 24.3464
R21808 commonsourceibias.n234 commonsourceibias.n212 24.3464
R21809 commonsourceibias.n244 commonsourceibias.n209 24.3464
R21810 commonsourceibias.n180 commonsourceibias.n145 24.3464
R21811 commonsourceibias.n170 commonsourceibias.n148 24.3464
R21812 commonsourceibias.n338 commonsourceibias.n316 24.3464
R21813 commonsourceibias.n349 commonsourceibias.n348 24.3464
R21814 commonsourceibias.n383 commonsourceibias.n382 24.3464
R21815 commonsourceibias.n297 commonsourceibias.n275 24.3464
R21816 commonsourceibias.n499 commonsourceibias.n477 24.3464
R21817 commonsourceibias.n510 commonsourceibias.n509 24.3464
R21818 commonsourceibias.n435 commonsourceibias.n413 24.3464
R21819 commonsourceibias.n446 commonsourceibias.n445 24.3464
R21820 commonsourceibias.n65 commonsourceibias.n10 23.8546
R21821 commonsourceibias.n27 commonsourceibias.n26 23.8546
R21822 commonsourceibias.n131 commonsourceibias.n1 23.8546
R21823 commonsourceibias.n93 commonsourceibias.n92 23.8546
R21824 commonsourceibias.n220 commonsourceibias.n219 23.8546
R21825 commonsourceibias.n258 commonsourceibias.n203 23.8546
R21826 commonsourceibias.n194 commonsourceibias.n139 23.8546
R21827 commonsourceibias.n156 commonsourceibias.n155 23.8546
R21828 commonsourceibias.n324 commonsourceibias.n323 23.8546
R21829 commonsourceibias.n363 commonsourceibias.n308 23.8546
R21830 commonsourceibias.n397 commonsourceibias.n267 23.8546
R21831 commonsourceibias.n283 commonsourceibias.n282 23.8546
R21832 commonsourceibias.n485 commonsourceibias.n484 23.8546
R21833 commonsourceibias.n524 commonsourceibias.n469 23.8546
R21834 commonsourceibias.n421 commonsourceibias.n420 23.8546
R21835 commonsourceibias.n460 commonsourceibias.n405 23.8546
R21836 commonsourceibias.n64 commonsourceibias.n63 16.9689
R21837 commonsourceibias.n28 commonsourceibias.n23 16.9689
R21838 commonsourceibias.n130 commonsourceibias.n129 16.9689
R21839 commonsourceibias.n94 commonsourceibias.n89 16.9689
R21840 commonsourceibias.n221 commonsourceibias.n216 16.9689
R21841 commonsourceibias.n257 commonsourceibias.n256 16.9689
R21842 commonsourceibias.n193 commonsourceibias.n192 16.9689
R21843 commonsourceibias.n157 commonsourceibias.n152 16.9689
R21844 commonsourceibias.n325 commonsourceibias.n320 16.9689
R21845 commonsourceibias.n362 commonsourceibias.n361 16.9689
R21846 commonsourceibias.n396 commonsourceibias.n395 16.9689
R21847 commonsourceibias.n284 commonsourceibias.n279 16.9689
R21848 commonsourceibias.n486 commonsourceibias.n481 16.9689
R21849 commonsourceibias.n523 commonsourceibias.n522 16.9689
R21850 commonsourceibias.n422 commonsourceibias.n417 16.9689
R21851 commonsourceibias.n459 commonsourceibias.n458 16.9689
R21852 commonsourceibias.n50 commonsourceibias.n49 16.477
R21853 commonsourceibias.n43 commonsourceibias.n42 16.477
R21854 commonsourceibias.n116 commonsourceibias.n115 16.477
R21855 commonsourceibias.n109 commonsourceibias.n108 16.477
R21856 commonsourceibias.n236 commonsourceibias.n235 16.477
R21857 commonsourceibias.n243 commonsourceibias.n242 16.477
R21858 commonsourceibias.n179 commonsourceibias.n178 16.477
R21859 commonsourceibias.n172 commonsourceibias.n171 16.477
R21860 commonsourceibias.n340 commonsourceibias.n339 16.477
R21861 commonsourceibias.n347 commonsourceibias.n346 16.477
R21862 commonsourceibias.n381 commonsourceibias.n380 16.477
R21863 commonsourceibias.n299 commonsourceibias.n298 16.477
R21864 commonsourceibias.n501 commonsourceibias.n500 16.477
R21865 commonsourceibias.n508 commonsourceibias.n507 16.477
R21866 commonsourceibias.n437 commonsourceibias.n436 16.477
R21867 commonsourceibias.n444 commonsourceibias.n443 16.477
R21868 commonsourceibias.n57 commonsourceibias.n56 15.9852
R21869 commonsourceibias.n36 commonsourceibias.n21 15.9852
R21870 commonsourceibias.n123 commonsourceibias.n122 15.9852
R21871 commonsourceibias.n102 commonsourceibias.n87 15.9852
R21872 commonsourceibias.n229 commonsourceibias.n214 15.9852
R21873 commonsourceibias.n250 commonsourceibias.n249 15.9852
R21874 commonsourceibias.n186 commonsourceibias.n185 15.9852
R21875 commonsourceibias.n165 commonsourceibias.n150 15.9852
R21876 commonsourceibias.n333 commonsourceibias.n318 15.9852
R21877 commonsourceibias.n355 commonsourceibias.n354 15.9852
R21878 commonsourceibias.n389 commonsourceibias.n388 15.9852
R21879 commonsourceibias.n292 commonsourceibias.n277 15.9852
R21880 commonsourceibias.n494 commonsourceibias.n479 15.9852
R21881 commonsourceibias.n516 commonsourceibias.n515 15.9852
R21882 commonsourceibias.n430 commonsourceibias.n415 15.9852
R21883 commonsourceibias.n452 commonsourceibias.n451 15.9852
R21884 commonsourceibias.n73 commonsourceibias.n71 13.2057
R21885 commonsourceibias.n371 commonsourceibias.n369 13.2057
R21886 commonsourceibias.n532 commonsourceibias.n265 10.122
R21887 commonsourceibias.n112 commonsourceibias.n83 9.50363
R21888 commonsourceibias.n377 commonsourceibias.n376 9.50363
R21889 commonsourceibias.n201 commonsourceibias.n137 8.7339
R21890 commonsourceibias.n467 commonsourceibias.n403 8.7339
R21891 commonsourceibias.n58 commonsourceibias.n57 8.60764
R21892 commonsourceibias.n33 commonsourceibias.n21 8.60764
R21893 commonsourceibias.n124 commonsourceibias.n123 8.60764
R21894 commonsourceibias.n99 commonsourceibias.n87 8.60764
R21895 commonsourceibias.n226 commonsourceibias.n214 8.60764
R21896 commonsourceibias.n251 commonsourceibias.n250 8.60764
R21897 commonsourceibias.n187 commonsourceibias.n186 8.60764
R21898 commonsourceibias.n162 commonsourceibias.n150 8.60764
R21899 commonsourceibias.n330 commonsourceibias.n318 8.60764
R21900 commonsourceibias.n356 commonsourceibias.n355 8.60764
R21901 commonsourceibias.n390 commonsourceibias.n389 8.60764
R21902 commonsourceibias.n289 commonsourceibias.n277 8.60764
R21903 commonsourceibias.n491 commonsourceibias.n479 8.60764
R21904 commonsourceibias.n517 commonsourceibias.n516 8.60764
R21905 commonsourceibias.n427 commonsourceibias.n415 8.60764
R21906 commonsourceibias.n453 commonsourceibias.n452 8.60764
R21907 commonsourceibias.n532 commonsourceibias.n531 8.46921
R21908 commonsourceibias.n49 commonsourceibias.n48 8.11581
R21909 commonsourceibias.n44 commonsourceibias.n43 8.11581
R21910 commonsourceibias.n115 commonsourceibias.n114 8.11581
R21911 commonsourceibias.n110 commonsourceibias.n109 8.11581
R21912 commonsourceibias.n237 commonsourceibias.n236 8.11581
R21913 commonsourceibias.n242 commonsourceibias.n241 8.11581
R21914 commonsourceibias.n178 commonsourceibias.n177 8.11581
R21915 commonsourceibias.n173 commonsourceibias.n172 8.11581
R21916 commonsourceibias.n341 commonsourceibias.n340 8.11581
R21917 commonsourceibias.n346 commonsourceibias.n345 8.11581
R21918 commonsourceibias.n380 commonsourceibias.n379 8.11581
R21919 commonsourceibias.n300 commonsourceibias.n299 8.11581
R21920 commonsourceibias.n502 commonsourceibias.n501 8.11581
R21921 commonsourceibias.n507 commonsourceibias.n506 8.11581
R21922 commonsourceibias.n438 commonsourceibias.n437 8.11581
R21923 commonsourceibias.n443 commonsourceibias.n442 8.11581
R21924 commonsourceibias.n63 commonsourceibias.n62 7.62397
R21925 commonsourceibias.n31 commonsourceibias.n23 7.62397
R21926 commonsourceibias.n129 commonsourceibias.n128 7.62397
R21927 commonsourceibias.n97 commonsourceibias.n89 7.62397
R21928 commonsourceibias.n224 commonsourceibias.n216 7.62397
R21929 commonsourceibias.n256 commonsourceibias.n255 7.62397
R21930 commonsourceibias.n192 commonsourceibias.n191 7.62397
R21931 commonsourceibias.n160 commonsourceibias.n152 7.62397
R21932 commonsourceibias.n328 commonsourceibias.n320 7.62397
R21933 commonsourceibias.n361 commonsourceibias.n360 7.62397
R21934 commonsourceibias.n395 commonsourceibias.n394 7.62397
R21935 commonsourceibias.n287 commonsourceibias.n279 7.62397
R21936 commonsourceibias.n489 commonsourceibias.n481 7.62397
R21937 commonsourceibias.n522 commonsourceibias.n521 7.62397
R21938 commonsourceibias.n425 commonsourceibias.n417 7.62397
R21939 commonsourceibias.n458 commonsourceibias.n457 7.62397
R21940 commonsourceibias.n265 commonsourceibias.n264 5.00473
R21941 commonsourceibias.n201 commonsourceibias.n200 5.00473
R21942 commonsourceibias.n531 commonsourceibias.n530 5.00473
R21943 commonsourceibias.n467 commonsourceibias.n466 5.00473
R21944 commonsourceibias commonsourceibias.n532 3.87639
R21945 commonsourceibias.n265 commonsourceibias.n201 3.72967
R21946 commonsourceibias.n531 commonsourceibias.n467 3.72967
R21947 commonsourceibias.n78 commonsourceibias.t17 2.82907
R21948 commonsourceibias.n78 commonsourceibias.t23 2.82907
R21949 commonsourceibias.n79 commonsourceibias.t11 2.82907
R21950 commonsourceibias.n79 commonsourceibias.t35 2.82907
R21951 commonsourceibias.n81 commonsourceibias.t21 2.82907
R21952 commonsourceibias.n81 commonsourceibias.t3 2.82907
R21953 commonsourceibias.n76 commonsourceibias.t45 2.82907
R21954 commonsourceibias.n76 commonsourceibias.t13 2.82907
R21955 commonsourceibias.n74 commonsourceibias.t1 2.82907
R21956 commonsourceibias.n74 commonsourceibias.t7 2.82907
R21957 commonsourceibias.n72 commonsourceibias.t9 2.82907
R21958 commonsourceibias.n72 commonsourceibias.t39 2.82907
R21959 commonsourceibias.n370 commonsourceibias.t47 2.82907
R21960 commonsourceibias.n370 commonsourceibias.t27 2.82907
R21961 commonsourceibias.n372 commonsourceibias.t25 2.82907
R21962 commonsourceibias.n372 commonsourceibias.t15 2.82907
R21963 commonsourceibias.n374 commonsourceibias.t31 2.82907
R21964 commonsourceibias.n374 commonsourceibias.t5 2.82907
R21965 commonsourceibias.n305 commonsourceibias.t19 2.82907
R21966 commonsourceibias.n305 commonsourceibias.t37 2.82907
R21967 commonsourceibias.n303 commonsourceibias.t43 2.82907
R21968 commonsourceibias.n303 commonsourceibias.t29 2.82907
R21969 commonsourceibias.n302 commonsourceibias.t41 2.82907
R21970 commonsourceibias.n302 commonsourceibias.t33 2.82907
R21971 commonsourceibias.n68 commonsourceibias.n10 0.738255
R21972 commonsourceibias.n134 commonsourceibias.n1 0.738255
R21973 commonsourceibias.n261 commonsourceibias.n203 0.738255
R21974 commonsourceibias.n197 commonsourceibias.n139 0.738255
R21975 commonsourceibias.n366 commonsourceibias.n308 0.738255
R21976 commonsourceibias.n400 commonsourceibias.n267 0.738255
R21977 commonsourceibias.n527 commonsourceibias.n469 0.738255
R21978 commonsourceibias.n463 commonsourceibias.n405 0.738255
R21979 commonsourceibias.n75 commonsourceibias.n73 0.573776
R21980 commonsourceibias.n77 commonsourceibias.n75 0.573776
R21981 commonsourceibias.n82 commonsourceibias.n80 0.573776
R21982 commonsourceibias.n306 commonsourceibias.n304 0.573776
R21983 commonsourceibias.n375 commonsourceibias.n373 0.573776
R21984 commonsourceibias.n373 commonsourceibias.n371 0.573776
R21985 commonsourceibias.n83 commonsourceibias.n77 0.287138
R21986 commonsourceibias.n83 commonsourceibias.n82 0.287138
R21987 commonsourceibias.n376 commonsourceibias.n306 0.287138
R21988 commonsourceibias.n376 commonsourceibias.n375 0.287138
R21989 commonsourceibias.n71 commonsourceibias.n9 0.285035
R21990 commonsourceibias.n137 commonsourceibias.n0 0.285035
R21991 commonsourceibias.n264 commonsourceibias.n202 0.285035
R21992 commonsourceibias.n200 commonsourceibias.n138 0.285035
R21993 commonsourceibias.n369 commonsourceibias.n307 0.285035
R21994 commonsourceibias.n403 commonsourceibias.n266 0.285035
R21995 commonsourceibias.n530 commonsourceibias.n468 0.285035
R21996 commonsourceibias.n466 commonsourceibias.n404 0.285035
R21997 commonsourceibias.n16 commonsourceibias.n14 0.246418
R21998 commonsourceibias.n38 commonsourceibias.n19 0.246418
R21999 commonsourceibias.n7 commonsourceibias.n5 0.246418
R22000 commonsourceibias.n104 commonsourceibias.n85 0.246418
R22001 commonsourceibias.n231 commonsourceibias.n212 0.246418
R22002 commonsourceibias.n209 commonsourceibias.n207 0.246418
R22003 commonsourceibias.n145 commonsourceibias.n143 0.246418
R22004 commonsourceibias.n167 commonsourceibias.n148 0.246418
R22005 commonsourceibias.n335 commonsourceibias.n316 0.246418
R22006 commonsourceibias.n348 commonsourceibias.n312 0.246418
R22007 commonsourceibias.n382 commonsourceibias.n271 0.246418
R22008 commonsourceibias.n294 commonsourceibias.n275 0.246418
R22009 commonsourceibias.n496 commonsourceibias.n477 0.246418
R22010 commonsourceibias.n509 commonsourceibias.n473 0.246418
R22011 commonsourceibias.n432 commonsourceibias.n413 0.246418
R22012 commonsourceibias.n445 commonsourceibias.n409 0.246418
R22013 commonsourceibias.n67 commonsourceibias.n9 0.189894
R22014 commonsourceibias.n67 commonsourceibias.n66 0.189894
R22015 commonsourceibias.n66 commonsourceibias.n11 0.189894
R22016 commonsourceibias.n61 commonsourceibias.n11 0.189894
R22017 commonsourceibias.n61 commonsourceibias.n60 0.189894
R22018 commonsourceibias.n60 commonsourceibias.n59 0.189894
R22019 commonsourceibias.n59 commonsourceibias.n13 0.189894
R22020 commonsourceibias.n54 commonsourceibias.n13 0.189894
R22021 commonsourceibias.n54 commonsourceibias.n53 0.189894
R22022 commonsourceibias.n53 commonsourceibias.n52 0.189894
R22023 commonsourceibias.n52 commonsourceibias.n15 0.189894
R22024 commonsourceibias.n47 commonsourceibias.n15 0.189894
R22025 commonsourceibias.n47 commonsourceibias.n46 0.189894
R22026 commonsourceibias.n46 commonsourceibias.n45 0.189894
R22027 commonsourceibias.n45 commonsourceibias.n18 0.189894
R22028 commonsourceibias.n40 commonsourceibias.n18 0.189894
R22029 commonsourceibias.n40 commonsourceibias.n39 0.189894
R22030 commonsourceibias.n39 commonsourceibias.n20 0.189894
R22031 commonsourceibias.n35 commonsourceibias.n20 0.189894
R22032 commonsourceibias.n35 commonsourceibias.n34 0.189894
R22033 commonsourceibias.n34 commonsourceibias.n22 0.189894
R22034 commonsourceibias.n30 commonsourceibias.n22 0.189894
R22035 commonsourceibias.n30 commonsourceibias.n29 0.189894
R22036 commonsourceibias.n29 commonsourceibias.n24 0.189894
R22037 commonsourceibias.n111 commonsourceibias.n84 0.189894
R22038 commonsourceibias.n106 commonsourceibias.n84 0.189894
R22039 commonsourceibias.n106 commonsourceibias.n105 0.189894
R22040 commonsourceibias.n105 commonsourceibias.n86 0.189894
R22041 commonsourceibias.n101 commonsourceibias.n86 0.189894
R22042 commonsourceibias.n101 commonsourceibias.n100 0.189894
R22043 commonsourceibias.n100 commonsourceibias.n88 0.189894
R22044 commonsourceibias.n96 commonsourceibias.n88 0.189894
R22045 commonsourceibias.n96 commonsourceibias.n95 0.189894
R22046 commonsourceibias.n95 commonsourceibias.n90 0.189894
R22047 commonsourceibias.n133 commonsourceibias.n0 0.189894
R22048 commonsourceibias.n133 commonsourceibias.n132 0.189894
R22049 commonsourceibias.n132 commonsourceibias.n2 0.189894
R22050 commonsourceibias.n127 commonsourceibias.n2 0.189894
R22051 commonsourceibias.n127 commonsourceibias.n126 0.189894
R22052 commonsourceibias.n126 commonsourceibias.n125 0.189894
R22053 commonsourceibias.n125 commonsourceibias.n4 0.189894
R22054 commonsourceibias.n120 commonsourceibias.n4 0.189894
R22055 commonsourceibias.n120 commonsourceibias.n119 0.189894
R22056 commonsourceibias.n119 commonsourceibias.n118 0.189894
R22057 commonsourceibias.n118 commonsourceibias.n6 0.189894
R22058 commonsourceibias.n113 commonsourceibias.n6 0.189894
R22059 commonsourceibias.n260 commonsourceibias.n202 0.189894
R22060 commonsourceibias.n260 commonsourceibias.n259 0.189894
R22061 commonsourceibias.n259 commonsourceibias.n204 0.189894
R22062 commonsourceibias.n254 commonsourceibias.n204 0.189894
R22063 commonsourceibias.n254 commonsourceibias.n253 0.189894
R22064 commonsourceibias.n253 commonsourceibias.n252 0.189894
R22065 commonsourceibias.n252 commonsourceibias.n206 0.189894
R22066 commonsourceibias.n247 commonsourceibias.n206 0.189894
R22067 commonsourceibias.n247 commonsourceibias.n246 0.189894
R22068 commonsourceibias.n246 commonsourceibias.n245 0.189894
R22069 commonsourceibias.n245 commonsourceibias.n208 0.189894
R22070 commonsourceibias.n240 commonsourceibias.n208 0.189894
R22071 commonsourceibias.n240 commonsourceibias.n239 0.189894
R22072 commonsourceibias.n239 commonsourceibias.n238 0.189894
R22073 commonsourceibias.n238 commonsourceibias.n211 0.189894
R22074 commonsourceibias.n233 commonsourceibias.n211 0.189894
R22075 commonsourceibias.n233 commonsourceibias.n232 0.189894
R22076 commonsourceibias.n232 commonsourceibias.n213 0.189894
R22077 commonsourceibias.n228 commonsourceibias.n213 0.189894
R22078 commonsourceibias.n228 commonsourceibias.n227 0.189894
R22079 commonsourceibias.n227 commonsourceibias.n215 0.189894
R22080 commonsourceibias.n223 commonsourceibias.n215 0.189894
R22081 commonsourceibias.n223 commonsourceibias.n222 0.189894
R22082 commonsourceibias.n222 commonsourceibias.n217 0.189894
R22083 commonsourceibias.n196 commonsourceibias.n138 0.189894
R22084 commonsourceibias.n196 commonsourceibias.n195 0.189894
R22085 commonsourceibias.n195 commonsourceibias.n140 0.189894
R22086 commonsourceibias.n190 commonsourceibias.n140 0.189894
R22087 commonsourceibias.n190 commonsourceibias.n189 0.189894
R22088 commonsourceibias.n189 commonsourceibias.n188 0.189894
R22089 commonsourceibias.n188 commonsourceibias.n142 0.189894
R22090 commonsourceibias.n183 commonsourceibias.n142 0.189894
R22091 commonsourceibias.n183 commonsourceibias.n182 0.189894
R22092 commonsourceibias.n182 commonsourceibias.n181 0.189894
R22093 commonsourceibias.n181 commonsourceibias.n144 0.189894
R22094 commonsourceibias.n176 commonsourceibias.n144 0.189894
R22095 commonsourceibias.n176 commonsourceibias.n175 0.189894
R22096 commonsourceibias.n175 commonsourceibias.n174 0.189894
R22097 commonsourceibias.n174 commonsourceibias.n147 0.189894
R22098 commonsourceibias.n169 commonsourceibias.n147 0.189894
R22099 commonsourceibias.n169 commonsourceibias.n168 0.189894
R22100 commonsourceibias.n168 commonsourceibias.n149 0.189894
R22101 commonsourceibias.n164 commonsourceibias.n149 0.189894
R22102 commonsourceibias.n164 commonsourceibias.n163 0.189894
R22103 commonsourceibias.n163 commonsourceibias.n151 0.189894
R22104 commonsourceibias.n159 commonsourceibias.n151 0.189894
R22105 commonsourceibias.n159 commonsourceibias.n158 0.189894
R22106 commonsourceibias.n158 commonsourceibias.n153 0.189894
R22107 commonsourceibias.n326 commonsourceibias.n321 0.189894
R22108 commonsourceibias.n327 commonsourceibias.n326 0.189894
R22109 commonsourceibias.n327 commonsourceibias.n319 0.189894
R22110 commonsourceibias.n331 commonsourceibias.n319 0.189894
R22111 commonsourceibias.n332 commonsourceibias.n331 0.189894
R22112 commonsourceibias.n332 commonsourceibias.n317 0.189894
R22113 commonsourceibias.n336 commonsourceibias.n317 0.189894
R22114 commonsourceibias.n337 commonsourceibias.n336 0.189894
R22115 commonsourceibias.n337 commonsourceibias.n315 0.189894
R22116 commonsourceibias.n342 commonsourceibias.n315 0.189894
R22117 commonsourceibias.n343 commonsourceibias.n342 0.189894
R22118 commonsourceibias.n344 commonsourceibias.n343 0.189894
R22119 commonsourceibias.n344 commonsourceibias.n313 0.189894
R22120 commonsourceibias.n350 commonsourceibias.n313 0.189894
R22121 commonsourceibias.n351 commonsourceibias.n350 0.189894
R22122 commonsourceibias.n352 commonsourceibias.n351 0.189894
R22123 commonsourceibias.n352 commonsourceibias.n311 0.189894
R22124 commonsourceibias.n357 commonsourceibias.n311 0.189894
R22125 commonsourceibias.n358 commonsourceibias.n357 0.189894
R22126 commonsourceibias.n359 commonsourceibias.n358 0.189894
R22127 commonsourceibias.n359 commonsourceibias.n309 0.189894
R22128 commonsourceibias.n364 commonsourceibias.n309 0.189894
R22129 commonsourceibias.n365 commonsourceibias.n364 0.189894
R22130 commonsourceibias.n365 commonsourceibias.n307 0.189894
R22131 commonsourceibias.n285 commonsourceibias.n280 0.189894
R22132 commonsourceibias.n286 commonsourceibias.n285 0.189894
R22133 commonsourceibias.n286 commonsourceibias.n278 0.189894
R22134 commonsourceibias.n290 commonsourceibias.n278 0.189894
R22135 commonsourceibias.n291 commonsourceibias.n290 0.189894
R22136 commonsourceibias.n291 commonsourceibias.n276 0.189894
R22137 commonsourceibias.n295 commonsourceibias.n276 0.189894
R22138 commonsourceibias.n296 commonsourceibias.n295 0.189894
R22139 commonsourceibias.n296 commonsourceibias.n274 0.189894
R22140 commonsourceibias.n301 commonsourceibias.n274 0.189894
R22141 commonsourceibias.n378 commonsourceibias.n272 0.189894
R22142 commonsourceibias.n384 commonsourceibias.n272 0.189894
R22143 commonsourceibias.n385 commonsourceibias.n384 0.189894
R22144 commonsourceibias.n386 commonsourceibias.n385 0.189894
R22145 commonsourceibias.n386 commonsourceibias.n270 0.189894
R22146 commonsourceibias.n391 commonsourceibias.n270 0.189894
R22147 commonsourceibias.n392 commonsourceibias.n391 0.189894
R22148 commonsourceibias.n393 commonsourceibias.n392 0.189894
R22149 commonsourceibias.n393 commonsourceibias.n268 0.189894
R22150 commonsourceibias.n398 commonsourceibias.n268 0.189894
R22151 commonsourceibias.n399 commonsourceibias.n398 0.189894
R22152 commonsourceibias.n399 commonsourceibias.n266 0.189894
R22153 commonsourceibias.n487 commonsourceibias.n482 0.189894
R22154 commonsourceibias.n488 commonsourceibias.n487 0.189894
R22155 commonsourceibias.n488 commonsourceibias.n480 0.189894
R22156 commonsourceibias.n492 commonsourceibias.n480 0.189894
R22157 commonsourceibias.n493 commonsourceibias.n492 0.189894
R22158 commonsourceibias.n493 commonsourceibias.n478 0.189894
R22159 commonsourceibias.n497 commonsourceibias.n478 0.189894
R22160 commonsourceibias.n498 commonsourceibias.n497 0.189894
R22161 commonsourceibias.n498 commonsourceibias.n476 0.189894
R22162 commonsourceibias.n503 commonsourceibias.n476 0.189894
R22163 commonsourceibias.n504 commonsourceibias.n503 0.189894
R22164 commonsourceibias.n505 commonsourceibias.n504 0.189894
R22165 commonsourceibias.n505 commonsourceibias.n474 0.189894
R22166 commonsourceibias.n511 commonsourceibias.n474 0.189894
R22167 commonsourceibias.n512 commonsourceibias.n511 0.189894
R22168 commonsourceibias.n513 commonsourceibias.n512 0.189894
R22169 commonsourceibias.n513 commonsourceibias.n472 0.189894
R22170 commonsourceibias.n518 commonsourceibias.n472 0.189894
R22171 commonsourceibias.n519 commonsourceibias.n518 0.189894
R22172 commonsourceibias.n520 commonsourceibias.n519 0.189894
R22173 commonsourceibias.n520 commonsourceibias.n470 0.189894
R22174 commonsourceibias.n525 commonsourceibias.n470 0.189894
R22175 commonsourceibias.n526 commonsourceibias.n525 0.189894
R22176 commonsourceibias.n526 commonsourceibias.n468 0.189894
R22177 commonsourceibias.n423 commonsourceibias.n418 0.189894
R22178 commonsourceibias.n424 commonsourceibias.n423 0.189894
R22179 commonsourceibias.n424 commonsourceibias.n416 0.189894
R22180 commonsourceibias.n428 commonsourceibias.n416 0.189894
R22181 commonsourceibias.n429 commonsourceibias.n428 0.189894
R22182 commonsourceibias.n429 commonsourceibias.n414 0.189894
R22183 commonsourceibias.n433 commonsourceibias.n414 0.189894
R22184 commonsourceibias.n434 commonsourceibias.n433 0.189894
R22185 commonsourceibias.n434 commonsourceibias.n412 0.189894
R22186 commonsourceibias.n439 commonsourceibias.n412 0.189894
R22187 commonsourceibias.n440 commonsourceibias.n439 0.189894
R22188 commonsourceibias.n441 commonsourceibias.n440 0.189894
R22189 commonsourceibias.n441 commonsourceibias.n410 0.189894
R22190 commonsourceibias.n447 commonsourceibias.n410 0.189894
R22191 commonsourceibias.n448 commonsourceibias.n447 0.189894
R22192 commonsourceibias.n449 commonsourceibias.n448 0.189894
R22193 commonsourceibias.n449 commonsourceibias.n408 0.189894
R22194 commonsourceibias.n454 commonsourceibias.n408 0.189894
R22195 commonsourceibias.n455 commonsourceibias.n454 0.189894
R22196 commonsourceibias.n456 commonsourceibias.n455 0.189894
R22197 commonsourceibias.n456 commonsourceibias.n406 0.189894
R22198 commonsourceibias.n461 commonsourceibias.n406 0.189894
R22199 commonsourceibias.n462 commonsourceibias.n461 0.189894
R22200 commonsourceibias.n462 commonsourceibias.n404 0.189894
R22201 commonsourceibias.n112 commonsourceibias.n111 0.170955
R22202 commonsourceibias.n113 commonsourceibias.n112 0.170955
R22203 commonsourceibias.n377 commonsourceibias.n301 0.170955
R22204 commonsourceibias.n378 commonsourceibias.n377 0.170955
R22205 a_n2408_n452.n75 a_n2408_n452.t63 512.366
R22206 a_n2408_n452.n65 a_n2408_n452.t54 512.366
R22207 a_n2408_n452.n76 a_n2408_n452.t48 512.366
R22208 a_n2408_n452.n73 a_n2408_n452.t71 512.366
R22209 a_n2408_n452.n66 a_n2408_n452.t60 512.366
R22210 a_n2408_n452.n74 a_n2408_n452.t59 512.366
R22211 a_n2408_n452.n71 a_n2408_n452.t67 512.366
R22212 a_n2408_n452.n67 a_n2408_n452.t52 512.366
R22213 a_n2408_n452.n72 a_n2408_n452.t53 512.366
R22214 a_n2408_n452.n69 a_n2408_n452.t55 512.366
R22215 a_n2408_n452.n68 a_n2408_n452.t64 512.366
R22216 a_n2408_n452.n70 a_n2408_n452.t75 512.366
R22217 a_n2408_n452.n25 a_n2408_n452.t74 539.01
R22218 a_n2408_n452.n80 a_n2408_n452.t57 512.366
R22219 a_n2408_n452.n79 a_n2408_n452.t61 512.366
R22220 a_n2408_n452.n53 a_n2408_n452.t51 512.366
R22221 a_n2408_n452.n78 a_n2408_n452.t66 512.366
R22222 a_n2408_n452.n27 a_n2408_n452.t17 539.01
R22223 a_n2408_n452.n81 a_n2408_n452.t9 512.366
R22224 a_n2408_n452.n52 a_n2408_n452.t11 512.366
R22225 a_n2408_n452.n29 a_n2408_n452.t21 539.01
R22226 a_n2408_n452.n95 a_n2408_n452.t19 512.366
R22227 a_n2408_n452.n94 a_n2408_n452.t25 512.366
R22228 a_n2408_n452.n17 a_n2408_n452.t29 539.01
R22229 a_n2408_n452.n61 a_n2408_n452.t31 512.366
R22230 a_n2408_n452.n62 a_n2408_n452.t15 512.366
R22231 a_n2408_n452.n56 a_n2408_n452.t27 512.366
R22232 a_n2408_n452.n63 a_n2408_n452.t23 512.366
R22233 a_n2408_n452.n21 a_n2408_n452.t69 539.01
R22234 a_n2408_n452.n58 a_n2408_n452.t70 512.366
R22235 a_n2408_n452.n59 a_n2408_n452.t49 512.366
R22236 a_n2408_n452.n57 a_n2408_n452.t56 512.366
R22237 a_n2408_n452.n60 a_n2408_n452.t65 512.366
R22238 a_n2408_n452.n5 a_n2408_n452.n51 70.1674
R22239 a_n2408_n452.n7 a_n2408_n452.n49 70.1674
R22240 a_n2408_n452.n9 a_n2408_n452.n47 70.1674
R22241 a_n2408_n452.n12 a_n2408_n452.n45 70.1674
R22242 a_n2408_n452.n37 a_n2408_n452.n23 70.3058
R22243 a_n2408_n452.n34 a_n2408_n452.n26 44.5595
R22244 a_n2408_n452.n94 a_n2408_n452.n34 20.9685
R22245 a_n2408_n452.n28 a_n2408_n452.n29 44.8194
R22246 a_n2408_n452.n27 a_n2408_n452.n26 44.8194
R22247 a_n2408_n452.n27 a_n2408_n452.n81 13.6566
R22248 a_n2408_n452.n24 a_n2408_n452.n36 70.1674
R22249 a_n2408_n452.n36 a_n2408_n452.n53 20.9683
R22250 a_n2408_n452.n35 a_n2408_n452.n24 75.0448
R22251 a_n2408_n452.n79 a_n2408_n452.n35 11.2134
R22252 a_n2408_n452.n22 a_n2408_n452.n25 44.8194
R22253 a_n2408_n452.n14 a_n2408_n452.n43 70.3058
R22254 a_n2408_n452.n18 a_n2408_n452.n40 70.3058
R22255 a_n2408_n452.n39 a_n2408_n452.n19 70.1674
R22256 a_n2408_n452.n39 a_n2408_n452.n57 20.9683
R22257 a_n2408_n452.n19 a_n2408_n452.n38 75.0448
R22258 a_n2408_n452.n59 a_n2408_n452.n38 11.2134
R22259 a_n2408_n452.n20 a_n2408_n452.n21 44.8194
R22260 a_n2408_n452.n42 a_n2408_n452.n15 70.1674
R22261 a_n2408_n452.n42 a_n2408_n452.n56 20.9683
R22262 a_n2408_n452.n15 a_n2408_n452.n41 75.0448
R22263 a_n2408_n452.n62 a_n2408_n452.n41 11.2134
R22264 a_n2408_n452.n16 a_n2408_n452.n17 44.8194
R22265 a_n2408_n452.n70 a_n2408_n452.n45 20.9683
R22266 a_n2408_n452.n44 a_n2408_n452.n13 75.0448
R22267 a_n2408_n452.n44 a_n2408_n452.n68 11.2134
R22268 a_n2408_n452.n13 a_n2408_n452.n69 161.3
R22269 a_n2408_n452.n72 a_n2408_n452.n47 20.9683
R22270 a_n2408_n452.n46 a_n2408_n452.n10 75.0448
R22271 a_n2408_n452.n46 a_n2408_n452.n67 11.2134
R22272 a_n2408_n452.n10 a_n2408_n452.n71 161.3
R22273 a_n2408_n452.n74 a_n2408_n452.n49 20.9683
R22274 a_n2408_n452.n48 a_n2408_n452.n8 75.0448
R22275 a_n2408_n452.n48 a_n2408_n452.n66 11.2134
R22276 a_n2408_n452.n8 a_n2408_n452.n73 161.3
R22277 a_n2408_n452.n76 a_n2408_n452.n51 20.9683
R22278 a_n2408_n452.n50 a_n2408_n452.n6 75.0448
R22279 a_n2408_n452.n50 a_n2408_n452.n65 11.2134
R22280 a_n2408_n452.n6 a_n2408_n452.n75 161.3
R22281 a_n2408_n452.n3 a_n2408_n452.n91 81.3764
R22282 a_n2408_n452.n4 a_n2408_n452.n85 81.3764
R22283 a_n2408_n452.n0 a_n2408_n452.n82 81.3764
R22284 a_n2408_n452.n3 a_n2408_n452.n92 80.9324
R22285 a_n2408_n452.n2 a_n2408_n452.n93 80.9324
R22286 a_n2408_n452.n2 a_n2408_n452.n90 80.9324
R22287 a_n2408_n452.n2 a_n2408_n452.n89 80.9324
R22288 a_n2408_n452.n1 a_n2408_n452.n88 80.9324
R22289 a_n2408_n452.n4 a_n2408_n452.n86 80.9324
R22290 a_n2408_n452.n0 a_n2408_n452.n87 80.9324
R22291 a_n2408_n452.n0 a_n2408_n452.n84 80.9324
R22292 a_n2408_n452.n0 a_n2408_n452.n83 80.9324
R22293 a_n2408_n452.n33 a_n2408_n452.t18 74.6477
R22294 a_n2408_n452.n30 a_n2408_n452.t30 74.6477
R22295 a_n2408_n452.n32 a_n2408_n452.t22 74.2899
R22296 a_n2408_n452.n31 a_n2408_n452.t14 74.2897
R22297 a_n2408_n452.n33 a_n2408_n452.n97 70.6783
R22298 a_n2408_n452.n31 a_n2408_n452.n55 70.6783
R22299 a_n2408_n452.n30 a_n2408_n452.n54 70.6783
R22300 a_n2408_n452.n98 a_n2408_n452.n33 70.6782
R22301 a_n2408_n452.n75 a_n2408_n452.n65 48.2005
R22302 a_n2408_n452.t68 a_n2408_n452.n51 533.335
R22303 a_n2408_n452.n73 a_n2408_n452.n66 48.2005
R22304 a_n2408_n452.t73 a_n2408_n452.n49 533.335
R22305 a_n2408_n452.n71 a_n2408_n452.n67 48.2005
R22306 a_n2408_n452.t62 a_n2408_n452.n47 533.335
R22307 a_n2408_n452.n69 a_n2408_n452.n68 48.2005
R22308 a_n2408_n452.t58 a_n2408_n452.n45 533.335
R22309 a_n2408_n452.n80 a_n2408_n452.n79 48.2005
R22310 a_n2408_n452.n78 a_n2408_n452.n36 20.9683
R22311 a_n2408_n452.n81 a_n2408_n452.n52 48.2005
R22312 a_n2408_n452.n95 a_n2408_n452.n94 48.2005
R22313 a_n2408_n452.n62 a_n2408_n452.n61 48.2005
R22314 a_n2408_n452.n63 a_n2408_n452.n42 20.9683
R22315 a_n2408_n452.n59 a_n2408_n452.n58 48.2005
R22316 a_n2408_n452.n60 a_n2408_n452.n39 20.9683
R22317 a_n2408_n452.n37 a_n2408_n452.t72 533.058
R22318 a_n2408_n452.t13 a_n2408_n452.n43 533.058
R22319 a_n2408_n452.t50 a_n2408_n452.n40 533.058
R22320 a_n2408_n452.n1 a_n2408_n452.n0 32.6799
R22321 a_n2408_n452.n76 a_n2408_n452.n50 35.3134
R22322 a_n2408_n452.n74 a_n2408_n452.n48 35.3134
R22323 a_n2408_n452.n72 a_n2408_n452.n46 35.3134
R22324 a_n2408_n452.n70 a_n2408_n452.n44 35.3134
R22325 a_n2408_n452.n35 a_n2408_n452.n53 35.3134
R22326 a_n2408_n452.n34 a_n2408_n452.n52 20.9689
R22327 a_n2408_n452.n56 a_n2408_n452.n41 35.3134
R22328 a_n2408_n452.n57 a_n2408_n452.n38 35.3134
R22329 a_n2408_n452.n26 a_n2408_n452.n2 23.891
R22330 a_n2408_n452.n20 a_n2408_n452.n11 12.046
R22331 a_n2408_n452.n23 a_n2408_n452.n77 11.8414
R22332 a_n2408_n452.n96 a_n2408_n452.n28 10.5365
R22333 a_n2408_n452.n64 a_n2408_n452.n31 9.50122
R22334 a_n2408_n452.n77 a_n2408_n452.n5 7.47588
R22335 a_n2408_n452.n13 a_n2408_n452.n11 7.47588
R22336 a_n2408_n452.n64 a_n2408_n452.n14 6.70126
R22337 a_n2408_n452.n32 a_n2408_n452.n96 5.65783
R22338 a_n2408_n452.n77 a_n2408_n452.n64 5.3452
R22339 a_n2408_n452.n26 a_n2408_n452.n22 3.95126
R22340 a_n2408_n452.n16 a_n2408_n452.n18 3.95126
R22341 a_n2408_n452.n97 a_n2408_n452.t20 3.61217
R22342 a_n2408_n452.n97 a_n2408_n452.t26 3.61217
R22343 a_n2408_n452.n55 a_n2408_n452.t28 3.61217
R22344 a_n2408_n452.n55 a_n2408_n452.t24 3.61217
R22345 a_n2408_n452.n54 a_n2408_n452.t32 3.61217
R22346 a_n2408_n452.n54 a_n2408_n452.t16 3.61217
R22347 a_n2408_n452.n98 a_n2408_n452.t12 3.61217
R22348 a_n2408_n452.t10 a_n2408_n452.n98 3.61217
R22349 a_n2408_n452.n91 a_n2408_n452.t0 2.82907
R22350 a_n2408_n452.n91 a_n2408_n452.t36 2.82907
R22351 a_n2408_n452.n92 a_n2408_n452.t44 2.82907
R22352 a_n2408_n452.n92 a_n2408_n452.t47 2.82907
R22353 a_n2408_n452.n93 a_n2408_n452.t40 2.82907
R22354 a_n2408_n452.n93 a_n2408_n452.t33 2.82907
R22355 a_n2408_n452.n90 a_n2408_n452.t37 2.82907
R22356 a_n2408_n452.n90 a_n2408_n452.t43 2.82907
R22357 a_n2408_n452.n89 a_n2408_n452.t34 2.82907
R22358 a_n2408_n452.n89 a_n2408_n452.t42 2.82907
R22359 a_n2408_n452.n88 a_n2408_n452.t45 2.82907
R22360 a_n2408_n452.n88 a_n2408_n452.t3 2.82907
R22361 a_n2408_n452.n85 a_n2408_n452.t46 2.82907
R22362 a_n2408_n452.n85 a_n2408_n452.t7 2.82907
R22363 a_n2408_n452.n86 a_n2408_n452.t6 2.82907
R22364 a_n2408_n452.n86 a_n2408_n452.t38 2.82907
R22365 a_n2408_n452.n87 a_n2408_n452.t5 2.82907
R22366 a_n2408_n452.n87 a_n2408_n452.t4 2.82907
R22367 a_n2408_n452.n84 a_n2408_n452.t2 2.82907
R22368 a_n2408_n452.n84 a_n2408_n452.t1 2.82907
R22369 a_n2408_n452.n83 a_n2408_n452.t41 2.82907
R22370 a_n2408_n452.n83 a_n2408_n452.t8 2.82907
R22371 a_n2408_n452.n82 a_n2408_n452.t39 2.82907
R22372 a_n2408_n452.n82 a_n2408_n452.t35 2.82907
R22373 a_n2408_n452.n96 a_n2408_n452.n11 1.30542
R22374 a_n2408_n452.n8 a_n2408_n452.n9 1.04595
R22375 a_n2408_n452.n25 a_n2408_n452.n80 13.657
R22376 a_n2408_n452.n78 a_n2408_n452.n37 21.4216
R22377 a_n2408_n452.n29 a_n2408_n452.n95 13.657
R22378 a_n2408_n452.n61 a_n2408_n452.n17 13.657
R22379 a_n2408_n452.n43 a_n2408_n452.n63 21.4216
R22380 a_n2408_n452.n58 a_n2408_n452.n21 13.657
R22381 a_n2408_n452.n40 a_n2408_n452.n60 21.4216
R22382 a_n2408_n452.n26 a_n2408_n452.n28 1.47777
R22383 a_n2408_n452.n0 a_n2408_n452.n4 1.3324
R22384 a_n2408_n452.n2 a_n2408_n452.n3 0.888431
R22385 a_n2408_n452.n2 a_n2408_n452.n1 0.888431
R22386 a_n2408_n452.n24 a_n2408_n452.n22 0.758076
R22387 a_n2408_n452.n24 a_n2408_n452.n23 0.758076
R22388 a_n2408_n452.n20 a_n2408_n452.n19 0.758076
R22389 a_n2408_n452.n19 a_n2408_n452.n18 0.758076
R22390 a_n2408_n452.n16 a_n2408_n452.n15 0.758076
R22391 a_n2408_n452.n15 a_n2408_n452.n14 0.758076
R22392 a_n2408_n452.n13 a_n2408_n452.n12 0.758076
R22393 a_n2408_n452.n10 a_n2408_n452.n9 0.758076
R22394 a_n2408_n452.n8 a_n2408_n452.n7 0.758076
R22395 a_n2408_n452.n6 a_n2408_n452.n5 0.758076
R22396 a_n2408_n452.n33 a_n2408_n452.n32 0.716017
R22397 a_n2408_n452.n31 a_n2408_n452.n30 0.716017
R22398 a_n2408_n452.n10 a_n2408_n452.n12 0.67853
R22399 a_n2408_n452.n6 a_n2408_n452.n7 0.67853
R22400 a_n1808_13878.n17 a_n1808_13878.n16 98.9632
R22401 a_n1808_13878.n2 a_n1808_13878.n0 98.7517
R22402 a_n1808_13878.n16 a_n1808_13878.n15 98.6055
R22403 a_n1808_13878.n4 a_n1808_13878.n3 98.6055
R22404 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R22405 a_n1808_13878.n14 a_n1808_13878.n13 98.6054
R22406 a_n1808_13878.n6 a_n1808_13878.t13 74.6477
R22407 a_n1808_13878.n11 a_n1808_13878.t14 74.2899
R22408 a_n1808_13878.n8 a_n1808_13878.t15 74.2899
R22409 a_n1808_13878.n7 a_n1808_13878.t12 74.2899
R22410 a_n1808_13878.n10 a_n1808_13878.n9 70.6783
R22411 a_n1808_13878.n6 a_n1808_13878.n5 70.6783
R22412 a_n1808_13878.n12 a_n1808_13878.n4 13.5694
R22413 a_n1808_13878.n14 a_n1808_13878.n12 11.5762
R22414 a_n1808_13878.n12 a_n1808_13878.n11 6.2408
R22415 a_n1808_13878.n13 a_n1808_13878.t9 3.61217
R22416 a_n1808_13878.n13 a_n1808_13878.t10 3.61217
R22417 a_n1808_13878.n15 a_n1808_13878.t0 3.61217
R22418 a_n1808_13878.n15 a_n1808_13878.t5 3.61217
R22419 a_n1808_13878.n9 a_n1808_13878.t18 3.61217
R22420 a_n1808_13878.n9 a_n1808_13878.t19 3.61217
R22421 a_n1808_13878.n5 a_n1808_13878.t16 3.61217
R22422 a_n1808_13878.n5 a_n1808_13878.t17 3.61217
R22423 a_n1808_13878.n3 a_n1808_13878.t6 3.61217
R22424 a_n1808_13878.n3 a_n1808_13878.t1 3.61217
R22425 a_n1808_13878.n1 a_n1808_13878.t8 3.61217
R22426 a_n1808_13878.n1 a_n1808_13878.t3 3.61217
R22427 a_n1808_13878.n0 a_n1808_13878.t2 3.61217
R22428 a_n1808_13878.n0 a_n1808_13878.t4 3.61217
R22429 a_n1808_13878.n17 a_n1808_13878.t7 3.61217
R22430 a_n1808_13878.t11 a_n1808_13878.n17 3.61217
R22431 a_n1808_13878.n7 a_n1808_13878.n6 0.358259
R22432 a_n1808_13878.n10 a_n1808_13878.n8 0.358259
R22433 a_n1808_13878.n11 a_n1808_13878.n10 0.358259
R22434 a_n1808_13878.n16 a_n1808_13878.n14 0.358259
R22435 a_n1808_13878.n4 a_n1808_13878.n2 0.146627
R22436 a_n1808_13878.n8 a_n1808_13878.n7 0.101793
R22437 minus.n53 minus.t28 323.478
R22438 minus.n11 minus.t8 323.478
R22439 minus.n82 minus.t13 297.12
R22440 minus.n80 minus.t15 297.12
R22441 minus.n44 minus.t5 297.12
R22442 minus.n74 minus.t6 297.12
R22443 minus.n46 minus.t26 297.12
R22444 minus.n68 minus.t21 297.12
R22445 minus.n48 minus.t23 297.12
R22446 minus.n62 minus.t16 297.12
R22447 minus.n50 minus.t17 297.12
R22448 minus.n56 minus.t9 297.12
R22449 minus.n52 minus.t27 297.12
R22450 minus.n10 minus.t7 297.12
R22451 minus.n14 minus.t11 297.12
R22452 minus.n16 minus.t10 297.12
R22453 minus.n20 minus.t12 297.12
R22454 minus.n22 minus.t20 297.12
R22455 minus.n26 minus.t18 297.12
R22456 minus.n28 minus.t25 297.12
R22457 minus.n32 minus.t24 297.12
R22458 minus.n34 minus.t14 297.12
R22459 minus.n38 minus.t22 297.12
R22460 minus.n40 minus.t19 297.12
R22461 minus.n88 minus.t2 243.255
R22462 minus.n87 minus.n85 224.169
R22463 minus.n87 minus.n86 223.454
R22464 minus.n55 minus.n54 161.3
R22465 minus.n56 minus.n51 161.3
R22466 minus.n58 minus.n57 161.3
R22467 minus.n59 minus.n50 161.3
R22468 minus.n61 minus.n60 161.3
R22469 minus.n62 minus.n49 161.3
R22470 minus.n64 minus.n63 161.3
R22471 minus.n65 minus.n48 161.3
R22472 minus.n67 minus.n66 161.3
R22473 minus.n68 minus.n47 161.3
R22474 minus.n70 minus.n69 161.3
R22475 minus.n71 minus.n46 161.3
R22476 minus.n73 minus.n72 161.3
R22477 minus.n74 minus.n45 161.3
R22478 minus.n76 minus.n75 161.3
R22479 minus.n77 minus.n44 161.3
R22480 minus.n79 minus.n78 161.3
R22481 minus.n80 minus.n43 161.3
R22482 minus.n81 minus.n42 161.3
R22483 minus.n83 minus.n82 161.3
R22484 minus.n41 minus.n40 161.3
R22485 minus.n39 minus.n0 161.3
R22486 minus.n38 minus.n37 161.3
R22487 minus.n36 minus.n1 161.3
R22488 minus.n35 minus.n34 161.3
R22489 minus.n33 minus.n2 161.3
R22490 minus.n32 minus.n31 161.3
R22491 minus.n30 minus.n3 161.3
R22492 minus.n29 minus.n28 161.3
R22493 minus.n27 minus.n4 161.3
R22494 minus.n26 minus.n25 161.3
R22495 minus.n24 minus.n5 161.3
R22496 minus.n23 minus.n22 161.3
R22497 minus.n21 minus.n6 161.3
R22498 minus.n20 minus.n19 161.3
R22499 minus.n18 minus.n7 161.3
R22500 minus.n17 minus.n16 161.3
R22501 minus.n15 minus.n8 161.3
R22502 minus.n14 minus.n13 161.3
R22503 minus.n12 minus.n9 161.3
R22504 minus.n82 minus.n81 46.0096
R22505 minus.n40 minus.n39 46.0096
R22506 minus.n12 minus.n11 45.0871
R22507 minus.n54 minus.n53 45.0871
R22508 minus.n80 minus.n79 41.6278
R22509 minus.n55 minus.n52 41.6278
R22510 minus.n10 minus.n9 41.6278
R22511 minus.n38 minus.n1 41.6278
R22512 minus.n75 minus.n44 37.246
R22513 minus.n57 minus.n56 37.246
R22514 minus.n15 minus.n14 37.246
R22515 minus.n34 minus.n33 37.246
R22516 minus.n84 minus.n83 33.3925
R22517 minus.n74 minus.n73 32.8641
R22518 minus.n61 minus.n50 32.8641
R22519 minus.n16 minus.n7 32.8641
R22520 minus.n32 minus.n3 32.8641
R22521 minus.n69 minus.n46 28.4823
R22522 minus.n63 minus.n62 28.4823
R22523 minus.n21 minus.n20 28.4823
R22524 minus.n28 minus.n27 28.4823
R22525 minus.n68 minus.n67 24.1005
R22526 minus.n67 minus.n48 24.1005
R22527 minus.n22 minus.n5 24.1005
R22528 minus.n26 minus.n5 24.1005
R22529 minus.n86 minus.t4 19.8005
R22530 minus.n86 minus.t3 19.8005
R22531 minus.n85 minus.t1 19.8005
R22532 minus.n85 minus.t0 19.8005
R22533 minus.n69 minus.n68 19.7187
R22534 minus.n63 minus.n48 19.7187
R22535 minus.n22 minus.n21 19.7187
R22536 minus.n27 minus.n26 19.7187
R22537 minus.n73 minus.n46 15.3369
R22538 minus.n62 minus.n61 15.3369
R22539 minus.n20 minus.n7 15.3369
R22540 minus.n28 minus.n3 15.3369
R22541 minus.n53 minus.n52 14.1472
R22542 minus.n11 minus.n10 14.1472
R22543 minus.n84 minus.n41 12.0933
R22544 minus minus.n89 11.0787
R22545 minus.n75 minus.n74 10.955
R22546 minus.n57 minus.n50 10.955
R22547 minus.n16 minus.n15 10.955
R22548 minus.n33 minus.n32 10.955
R22549 minus.n79 minus.n44 6.57323
R22550 minus.n56 minus.n55 6.57323
R22551 minus.n14 minus.n9 6.57323
R22552 minus.n34 minus.n1 6.57323
R22553 minus.n89 minus.n88 4.80222
R22554 minus.n81 minus.n80 2.19141
R22555 minus.n39 minus.n38 2.19141
R22556 minus.n89 minus.n84 0.972091
R22557 minus.n88 minus.n87 0.716017
R22558 minus.n83 minus.n42 0.189894
R22559 minus.n43 minus.n42 0.189894
R22560 minus.n78 minus.n43 0.189894
R22561 minus.n78 minus.n77 0.189894
R22562 minus.n77 minus.n76 0.189894
R22563 minus.n76 minus.n45 0.189894
R22564 minus.n72 minus.n45 0.189894
R22565 minus.n72 minus.n71 0.189894
R22566 minus.n71 minus.n70 0.189894
R22567 minus.n70 minus.n47 0.189894
R22568 minus.n66 minus.n47 0.189894
R22569 minus.n66 minus.n65 0.189894
R22570 minus.n65 minus.n64 0.189894
R22571 minus.n64 minus.n49 0.189894
R22572 minus.n60 minus.n49 0.189894
R22573 minus.n60 minus.n59 0.189894
R22574 minus.n59 minus.n58 0.189894
R22575 minus.n58 minus.n51 0.189894
R22576 minus.n54 minus.n51 0.189894
R22577 minus.n13 minus.n12 0.189894
R22578 minus.n13 minus.n8 0.189894
R22579 minus.n17 minus.n8 0.189894
R22580 minus.n18 minus.n17 0.189894
R22581 minus.n19 minus.n18 0.189894
R22582 minus.n19 minus.n6 0.189894
R22583 minus.n23 minus.n6 0.189894
R22584 minus.n24 minus.n23 0.189894
R22585 minus.n25 minus.n24 0.189894
R22586 minus.n25 minus.n4 0.189894
R22587 minus.n29 minus.n4 0.189894
R22588 minus.n30 minus.n29 0.189894
R22589 minus.n31 minus.n30 0.189894
R22590 minus.n31 minus.n2 0.189894
R22591 minus.n35 minus.n2 0.189894
R22592 minus.n36 minus.n35 0.189894
R22593 minus.n37 minus.n36 0.189894
R22594 minus.n37 minus.n0 0.189894
R22595 minus.n41 minus.n0 0.189894
R22596 outputibias.n27 outputibias.n1 289.615
R22597 outputibias.n58 outputibias.n32 289.615
R22598 outputibias.n90 outputibias.n64 289.615
R22599 outputibias.n122 outputibias.n96 289.615
R22600 outputibias.n28 outputibias.n27 185
R22601 outputibias.n26 outputibias.n25 185
R22602 outputibias.n5 outputibias.n4 185
R22603 outputibias.n20 outputibias.n19 185
R22604 outputibias.n18 outputibias.n17 185
R22605 outputibias.n9 outputibias.n8 185
R22606 outputibias.n12 outputibias.n11 185
R22607 outputibias.n59 outputibias.n58 185
R22608 outputibias.n57 outputibias.n56 185
R22609 outputibias.n36 outputibias.n35 185
R22610 outputibias.n51 outputibias.n50 185
R22611 outputibias.n49 outputibias.n48 185
R22612 outputibias.n40 outputibias.n39 185
R22613 outputibias.n43 outputibias.n42 185
R22614 outputibias.n91 outputibias.n90 185
R22615 outputibias.n89 outputibias.n88 185
R22616 outputibias.n68 outputibias.n67 185
R22617 outputibias.n83 outputibias.n82 185
R22618 outputibias.n81 outputibias.n80 185
R22619 outputibias.n72 outputibias.n71 185
R22620 outputibias.n75 outputibias.n74 185
R22621 outputibias.n123 outputibias.n122 185
R22622 outputibias.n121 outputibias.n120 185
R22623 outputibias.n100 outputibias.n99 185
R22624 outputibias.n115 outputibias.n114 185
R22625 outputibias.n113 outputibias.n112 185
R22626 outputibias.n104 outputibias.n103 185
R22627 outputibias.n107 outputibias.n106 185
R22628 outputibias.n0 outputibias.t9 178.945
R22629 outputibias.n133 outputibias.t8 177.018
R22630 outputibias.n132 outputibias.t11 177.018
R22631 outputibias.n0 outputibias.t10 177.018
R22632 outputibias.t5 outputibias.n10 147.661
R22633 outputibias.t7 outputibias.n41 147.661
R22634 outputibias.t1 outputibias.n73 147.661
R22635 outputibias.t3 outputibias.n105 147.661
R22636 outputibias.n128 outputibias.t4 132.363
R22637 outputibias.n128 outputibias.t6 130.436
R22638 outputibias.n129 outputibias.t0 130.436
R22639 outputibias.n130 outputibias.t2 130.436
R22640 outputibias.n27 outputibias.n26 104.615
R22641 outputibias.n26 outputibias.n4 104.615
R22642 outputibias.n19 outputibias.n4 104.615
R22643 outputibias.n19 outputibias.n18 104.615
R22644 outputibias.n18 outputibias.n8 104.615
R22645 outputibias.n11 outputibias.n8 104.615
R22646 outputibias.n58 outputibias.n57 104.615
R22647 outputibias.n57 outputibias.n35 104.615
R22648 outputibias.n50 outputibias.n35 104.615
R22649 outputibias.n50 outputibias.n49 104.615
R22650 outputibias.n49 outputibias.n39 104.615
R22651 outputibias.n42 outputibias.n39 104.615
R22652 outputibias.n90 outputibias.n89 104.615
R22653 outputibias.n89 outputibias.n67 104.615
R22654 outputibias.n82 outputibias.n67 104.615
R22655 outputibias.n82 outputibias.n81 104.615
R22656 outputibias.n81 outputibias.n71 104.615
R22657 outputibias.n74 outputibias.n71 104.615
R22658 outputibias.n122 outputibias.n121 104.615
R22659 outputibias.n121 outputibias.n99 104.615
R22660 outputibias.n114 outputibias.n99 104.615
R22661 outputibias.n114 outputibias.n113 104.615
R22662 outputibias.n113 outputibias.n103 104.615
R22663 outputibias.n106 outputibias.n103 104.615
R22664 outputibias.n63 outputibias.n31 95.6354
R22665 outputibias.n63 outputibias.n62 94.6732
R22666 outputibias.n95 outputibias.n94 94.6732
R22667 outputibias.n127 outputibias.n126 94.6732
R22668 outputibias.n11 outputibias.t5 52.3082
R22669 outputibias.n42 outputibias.t7 52.3082
R22670 outputibias.n74 outputibias.t1 52.3082
R22671 outputibias.n106 outputibias.t3 52.3082
R22672 outputibias.n12 outputibias.n10 15.6674
R22673 outputibias.n43 outputibias.n41 15.6674
R22674 outputibias.n75 outputibias.n73 15.6674
R22675 outputibias.n107 outputibias.n105 15.6674
R22676 outputibias.n13 outputibias.n9 12.8005
R22677 outputibias.n44 outputibias.n40 12.8005
R22678 outputibias.n76 outputibias.n72 12.8005
R22679 outputibias.n108 outputibias.n104 12.8005
R22680 outputibias.n17 outputibias.n16 12.0247
R22681 outputibias.n48 outputibias.n47 12.0247
R22682 outputibias.n80 outputibias.n79 12.0247
R22683 outputibias.n112 outputibias.n111 12.0247
R22684 outputibias.n20 outputibias.n7 11.249
R22685 outputibias.n51 outputibias.n38 11.249
R22686 outputibias.n83 outputibias.n70 11.249
R22687 outputibias.n115 outputibias.n102 11.249
R22688 outputibias.n21 outputibias.n5 10.4732
R22689 outputibias.n52 outputibias.n36 10.4732
R22690 outputibias.n84 outputibias.n68 10.4732
R22691 outputibias.n116 outputibias.n100 10.4732
R22692 outputibias.n25 outputibias.n24 9.69747
R22693 outputibias.n56 outputibias.n55 9.69747
R22694 outputibias.n88 outputibias.n87 9.69747
R22695 outputibias.n120 outputibias.n119 9.69747
R22696 outputibias.n31 outputibias.n30 9.45567
R22697 outputibias.n62 outputibias.n61 9.45567
R22698 outputibias.n94 outputibias.n93 9.45567
R22699 outputibias.n126 outputibias.n125 9.45567
R22700 outputibias.n30 outputibias.n29 9.3005
R22701 outputibias.n3 outputibias.n2 9.3005
R22702 outputibias.n24 outputibias.n23 9.3005
R22703 outputibias.n22 outputibias.n21 9.3005
R22704 outputibias.n7 outputibias.n6 9.3005
R22705 outputibias.n16 outputibias.n15 9.3005
R22706 outputibias.n14 outputibias.n13 9.3005
R22707 outputibias.n61 outputibias.n60 9.3005
R22708 outputibias.n34 outputibias.n33 9.3005
R22709 outputibias.n55 outputibias.n54 9.3005
R22710 outputibias.n53 outputibias.n52 9.3005
R22711 outputibias.n38 outputibias.n37 9.3005
R22712 outputibias.n47 outputibias.n46 9.3005
R22713 outputibias.n45 outputibias.n44 9.3005
R22714 outputibias.n93 outputibias.n92 9.3005
R22715 outputibias.n66 outputibias.n65 9.3005
R22716 outputibias.n87 outputibias.n86 9.3005
R22717 outputibias.n85 outputibias.n84 9.3005
R22718 outputibias.n70 outputibias.n69 9.3005
R22719 outputibias.n79 outputibias.n78 9.3005
R22720 outputibias.n77 outputibias.n76 9.3005
R22721 outputibias.n125 outputibias.n124 9.3005
R22722 outputibias.n98 outputibias.n97 9.3005
R22723 outputibias.n119 outputibias.n118 9.3005
R22724 outputibias.n117 outputibias.n116 9.3005
R22725 outputibias.n102 outputibias.n101 9.3005
R22726 outputibias.n111 outputibias.n110 9.3005
R22727 outputibias.n109 outputibias.n108 9.3005
R22728 outputibias.n28 outputibias.n3 8.92171
R22729 outputibias.n59 outputibias.n34 8.92171
R22730 outputibias.n91 outputibias.n66 8.92171
R22731 outputibias.n123 outputibias.n98 8.92171
R22732 outputibias.n29 outputibias.n1 8.14595
R22733 outputibias.n60 outputibias.n32 8.14595
R22734 outputibias.n92 outputibias.n64 8.14595
R22735 outputibias.n124 outputibias.n96 8.14595
R22736 outputibias.n31 outputibias.n1 5.81868
R22737 outputibias.n62 outputibias.n32 5.81868
R22738 outputibias.n94 outputibias.n64 5.81868
R22739 outputibias.n126 outputibias.n96 5.81868
R22740 outputibias.n131 outputibias.n130 5.20947
R22741 outputibias.n29 outputibias.n28 5.04292
R22742 outputibias.n60 outputibias.n59 5.04292
R22743 outputibias.n92 outputibias.n91 5.04292
R22744 outputibias.n124 outputibias.n123 5.04292
R22745 outputibias.n131 outputibias.n127 4.42209
R22746 outputibias.n14 outputibias.n10 4.38594
R22747 outputibias.n45 outputibias.n41 4.38594
R22748 outputibias.n77 outputibias.n73 4.38594
R22749 outputibias.n109 outputibias.n105 4.38594
R22750 outputibias.n132 outputibias.n131 4.28454
R22751 outputibias.n25 outputibias.n3 4.26717
R22752 outputibias.n56 outputibias.n34 4.26717
R22753 outputibias.n88 outputibias.n66 4.26717
R22754 outputibias.n120 outputibias.n98 4.26717
R22755 outputibias.n24 outputibias.n5 3.49141
R22756 outputibias.n55 outputibias.n36 3.49141
R22757 outputibias.n87 outputibias.n68 3.49141
R22758 outputibias.n119 outputibias.n100 3.49141
R22759 outputibias.n21 outputibias.n20 2.71565
R22760 outputibias.n52 outputibias.n51 2.71565
R22761 outputibias.n84 outputibias.n83 2.71565
R22762 outputibias.n116 outputibias.n115 2.71565
R22763 outputibias.n17 outputibias.n7 1.93989
R22764 outputibias.n48 outputibias.n38 1.93989
R22765 outputibias.n80 outputibias.n70 1.93989
R22766 outputibias.n112 outputibias.n102 1.93989
R22767 outputibias.n130 outputibias.n129 1.9266
R22768 outputibias.n129 outputibias.n128 1.9266
R22769 outputibias.n133 outputibias.n132 1.92658
R22770 outputibias.n134 outputibias.n133 1.29913
R22771 outputibias.n16 outputibias.n9 1.16414
R22772 outputibias.n47 outputibias.n40 1.16414
R22773 outputibias.n79 outputibias.n72 1.16414
R22774 outputibias.n111 outputibias.n104 1.16414
R22775 outputibias.n127 outputibias.n95 0.962709
R22776 outputibias.n95 outputibias.n63 0.962709
R22777 outputibias.n13 outputibias.n12 0.388379
R22778 outputibias.n44 outputibias.n43 0.388379
R22779 outputibias.n76 outputibias.n75 0.388379
R22780 outputibias.n108 outputibias.n107 0.388379
R22781 outputibias.n134 outputibias.n0 0.337251
R22782 outputibias outputibias.n134 0.302375
R22783 outputibias.n30 outputibias.n2 0.155672
R22784 outputibias.n23 outputibias.n2 0.155672
R22785 outputibias.n23 outputibias.n22 0.155672
R22786 outputibias.n22 outputibias.n6 0.155672
R22787 outputibias.n15 outputibias.n6 0.155672
R22788 outputibias.n15 outputibias.n14 0.155672
R22789 outputibias.n61 outputibias.n33 0.155672
R22790 outputibias.n54 outputibias.n33 0.155672
R22791 outputibias.n54 outputibias.n53 0.155672
R22792 outputibias.n53 outputibias.n37 0.155672
R22793 outputibias.n46 outputibias.n37 0.155672
R22794 outputibias.n46 outputibias.n45 0.155672
R22795 outputibias.n93 outputibias.n65 0.155672
R22796 outputibias.n86 outputibias.n65 0.155672
R22797 outputibias.n86 outputibias.n85 0.155672
R22798 outputibias.n85 outputibias.n69 0.155672
R22799 outputibias.n78 outputibias.n69 0.155672
R22800 outputibias.n78 outputibias.n77 0.155672
R22801 outputibias.n125 outputibias.n97 0.155672
R22802 outputibias.n118 outputibias.n97 0.155672
R22803 outputibias.n118 outputibias.n117 0.155672
R22804 outputibias.n117 outputibias.n101 0.155672
R22805 outputibias.n110 outputibias.n101 0.155672
R22806 outputibias.n110 outputibias.n109 0.155672
R22807 output.n41 output.n15 289.615
R22808 output.n72 output.n46 289.615
R22809 output.n104 output.n78 289.615
R22810 output.n136 output.n110 289.615
R22811 output.n77 output.n45 197.26
R22812 output.n77 output.n76 196.298
R22813 output.n109 output.n108 196.298
R22814 output.n141 output.n140 196.298
R22815 output.n42 output.n41 185
R22816 output.n40 output.n39 185
R22817 output.n19 output.n18 185
R22818 output.n34 output.n33 185
R22819 output.n32 output.n31 185
R22820 output.n23 output.n22 185
R22821 output.n26 output.n25 185
R22822 output.n73 output.n72 185
R22823 output.n71 output.n70 185
R22824 output.n50 output.n49 185
R22825 output.n65 output.n64 185
R22826 output.n63 output.n62 185
R22827 output.n54 output.n53 185
R22828 output.n57 output.n56 185
R22829 output.n105 output.n104 185
R22830 output.n103 output.n102 185
R22831 output.n82 output.n81 185
R22832 output.n97 output.n96 185
R22833 output.n95 output.n94 185
R22834 output.n86 output.n85 185
R22835 output.n89 output.n88 185
R22836 output.n137 output.n136 185
R22837 output.n135 output.n134 185
R22838 output.n114 output.n113 185
R22839 output.n129 output.n128 185
R22840 output.n127 output.n126 185
R22841 output.n118 output.n117 185
R22842 output.n121 output.n120 185
R22843 output.t18 output.n24 147.661
R22844 output.t17 output.n55 147.661
R22845 output.t19 output.n87 147.661
R22846 output.t16 output.n119 147.661
R22847 output.n41 output.n40 104.615
R22848 output.n40 output.n18 104.615
R22849 output.n33 output.n18 104.615
R22850 output.n33 output.n32 104.615
R22851 output.n32 output.n22 104.615
R22852 output.n25 output.n22 104.615
R22853 output.n72 output.n71 104.615
R22854 output.n71 output.n49 104.615
R22855 output.n64 output.n49 104.615
R22856 output.n64 output.n63 104.615
R22857 output.n63 output.n53 104.615
R22858 output.n56 output.n53 104.615
R22859 output.n104 output.n103 104.615
R22860 output.n103 output.n81 104.615
R22861 output.n96 output.n81 104.615
R22862 output.n96 output.n95 104.615
R22863 output.n95 output.n85 104.615
R22864 output.n88 output.n85 104.615
R22865 output.n136 output.n135 104.615
R22866 output.n135 output.n113 104.615
R22867 output.n128 output.n113 104.615
R22868 output.n128 output.n127 104.615
R22869 output.n127 output.n117 104.615
R22870 output.n120 output.n117 104.615
R22871 output.n1 output.t4 77.056
R22872 output.n14 output.t5 76.6694
R22873 output.n1 output.n0 72.7095
R22874 output.n3 output.n2 72.7095
R22875 output.n5 output.n4 72.7095
R22876 output.n7 output.n6 72.7095
R22877 output.n9 output.n8 72.7095
R22878 output.n11 output.n10 72.7095
R22879 output.n13 output.n12 72.7095
R22880 output.n25 output.t18 52.3082
R22881 output.n56 output.t17 52.3082
R22882 output.n88 output.t19 52.3082
R22883 output.n120 output.t16 52.3082
R22884 output.n26 output.n24 15.6674
R22885 output.n57 output.n55 15.6674
R22886 output.n89 output.n87 15.6674
R22887 output.n121 output.n119 15.6674
R22888 output.n27 output.n23 12.8005
R22889 output.n58 output.n54 12.8005
R22890 output.n90 output.n86 12.8005
R22891 output.n122 output.n118 12.8005
R22892 output.n31 output.n30 12.0247
R22893 output.n62 output.n61 12.0247
R22894 output.n94 output.n93 12.0247
R22895 output.n126 output.n125 12.0247
R22896 output.n34 output.n21 11.249
R22897 output.n65 output.n52 11.249
R22898 output.n97 output.n84 11.249
R22899 output.n129 output.n116 11.249
R22900 output.n35 output.n19 10.4732
R22901 output.n66 output.n50 10.4732
R22902 output.n98 output.n82 10.4732
R22903 output.n130 output.n114 10.4732
R22904 output.n39 output.n38 9.69747
R22905 output.n70 output.n69 9.69747
R22906 output.n102 output.n101 9.69747
R22907 output.n134 output.n133 9.69747
R22908 output.n45 output.n44 9.45567
R22909 output.n76 output.n75 9.45567
R22910 output.n108 output.n107 9.45567
R22911 output.n140 output.n139 9.45567
R22912 output.n44 output.n43 9.3005
R22913 output.n17 output.n16 9.3005
R22914 output.n38 output.n37 9.3005
R22915 output.n36 output.n35 9.3005
R22916 output.n21 output.n20 9.3005
R22917 output.n30 output.n29 9.3005
R22918 output.n28 output.n27 9.3005
R22919 output.n75 output.n74 9.3005
R22920 output.n48 output.n47 9.3005
R22921 output.n69 output.n68 9.3005
R22922 output.n67 output.n66 9.3005
R22923 output.n52 output.n51 9.3005
R22924 output.n61 output.n60 9.3005
R22925 output.n59 output.n58 9.3005
R22926 output.n107 output.n106 9.3005
R22927 output.n80 output.n79 9.3005
R22928 output.n101 output.n100 9.3005
R22929 output.n99 output.n98 9.3005
R22930 output.n84 output.n83 9.3005
R22931 output.n93 output.n92 9.3005
R22932 output.n91 output.n90 9.3005
R22933 output.n139 output.n138 9.3005
R22934 output.n112 output.n111 9.3005
R22935 output.n133 output.n132 9.3005
R22936 output.n131 output.n130 9.3005
R22937 output.n116 output.n115 9.3005
R22938 output.n125 output.n124 9.3005
R22939 output.n123 output.n122 9.3005
R22940 output.n42 output.n17 8.92171
R22941 output.n73 output.n48 8.92171
R22942 output.n105 output.n80 8.92171
R22943 output.n137 output.n112 8.92171
R22944 output output.n141 8.15037
R22945 output.n43 output.n15 8.14595
R22946 output.n74 output.n46 8.14595
R22947 output.n106 output.n78 8.14595
R22948 output.n138 output.n110 8.14595
R22949 output.n45 output.n15 5.81868
R22950 output.n76 output.n46 5.81868
R22951 output.n108 output.n78 5.81868
R22952 output.n140 output.n110 5.81868
R22953 output.n43 output.n42 5.04292
R22954 output.n74 output.n73 5.04292
R22955 output.n106 output.n105 5.04292
R22956 output.n138 output.n137 5.04292
R22957 output.n28 output.n24 4.38594
R22958 output.n59 output.n55 4.38594
R22959 output.n91 output.n87 4.38594
R22960 output.n123 output.n119 4.38594
R22961 output.n39 output.n17 4.26717
R22962 output.n70 output.n48 4.26717
R22963 output.n102 output.n80 4.26717
R22964 output.n134 output.n112 4.26717
R22965 output.n0 output.t10 3.9605
R22966 output.n0 output.t14 3.9605
R22967 output.n2 output.t1 3.9605
R22968 output.n2 output.t6 3.9605
R22969 output.n4 output.t7 3.9605
R22970 output.n4 output.t12 3.9605
R22971 output.n6 output.t0 3.9605
R22972 output.n6 output.t8 3.9605
R22973 output.n8 output.t11 3.9605
R22974 output.n8 output.t9 3.9605
R22975 output.n10 output.t15 3.9605
R22976 output.n10 output.t2 3.9605
R22977 output.n12 output.t3 3.9605
R22978 output.n12 output.t13 3.9605
R22979 output.n38 output.n19 3.49141
R22980 output.n69 output.n50 3.49141
R22981 output.n101 output.n82 3.49141
R22982 output.n133 output.n114 3.49141
R22983 output.n35 output.n34 2.71565
R22984 output.n66 output.n65 2.71565
R22985 output.n98 output.n97 2.71565
R22986 output.n130 output.n129 2.71565
R22987 output.n31 output.n21 1.93989
R22988 output.n62 output.n52 1.93989
R22989 output.n94 output.n84 1.93989
R22990 output.n126 output.n116 1.93989
R22991 output.n30 output.n23 1.16414
R22992 output.n61 output.n54 1.16414
R22993 output.n93 output.n86 1.16414
R22994 output.n125 output.n118 1.16414
R22995 output.n141 output.n109 0.962709
R22996 output.n109 output.n77 0.962709
R22997 output.n27 output.n26 0.388379
R22998 output.n58 output.n57 0.388379
R22999 output.n90 output.n89 0.388379
R23000 output.n122 output.n121 0.388379
R23001 output.n14 output.n13 0.387128
R23002 output.n13 output.n11 0.387128
R23003 output.n11 output.n9 0.387128
R23004 output.n9 output.n7 0.387128
R23005 output.n7 output.n5 0.387128
R23006 output.n5 output.n3 0.387128
R23007 output.n3 output.n1 0.387128
R23008 output.n44 output.n16 0.155672
R23009 output.n37 output.n16 0.155672
R23010 output.n37 output.n36 0.155672
R23011 output.n36 output.n20 0.155672
R23012 output.n29 output.n20 0.155672
R23013 output.n29 output.n28 0.155672
R23014 output.n75 output.n47 0.155672
R23015 output.n68 output.n47 0.155672
R23016 output.n68 output.n67 0.155672
R23017 output.n67 output.n51 0.155672
R23018 output.n60 output.n51 0.155672
R23019 output.n60 output.n59 0.155672
R23020 output.n107 output.n79 0.155672
R23021 output.n100 output.n79 0.155672
R23022 output.n100 output.n99 0.155672
R23023 output.n99 output.n83 0.155672
R23024 output.n92 output.n83 0.155672
R23025 output.n92 output.n91 0.155672
R23026 output.n139 output.n111 0.155672
R23027 output.n132 output.n111 0.155672
R23028 output.n132 output.n131 0.155672
R23029 output.n131 output.n115 0.155672
R23030 output.n124 output.n115 0.155672
R23031 output.n124 output.n123 0.155672
R23032 output output.n14 0.126227
R23033 a_n1986_8322.n6 a_n1986_8322.t3 74.6477
R23034 a_n1986_8322.n1 a_n1986_8322.t9 74.6477
R23035 a_n1986_8322.n16 a_n1986_8322.t18 74.6474
R23036 a_n1986_8322.n14 a_n1986_8322.t11 74.2899
R23037 a_n1986_8322.n7 a_n1986_8322.t1 74.2899
R23038 a_n1986_8322.n8 a_n1986_8322.t4 74.2899
R23039 a_n1986_8322.n11 a_n1986_8322.t5 74.2899
R23040 a_n1986_8322.n4 a_n1986_8322.t8 74.2899
R23041 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R23042 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R23043 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R23044 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R23045 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R23046 a_n1986_8322.n18 a_n1986_8322.n17 70.6782
R23047 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R23048 a_n1986_8322.n13 a_n1986_8322.t20 9.7972
R23049 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R23050 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R23051 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R23052 a_n1986_8322.n15 a_n1986_8322.t16 3.61217
R23053 a_n1986_8322.n15 a_n1986_8322.t13 3.61217
R23054 a_n1986_8322.n5 a_n1986_8322.t7 3.61217
R23055 a_n1986_8322.n5 a_n1986_8322.t6 3.61217
R23056 a_n1986_8322.n9 a_n1986_8322.t2 3.61217
R23057 a_n1986_8322.n9 a_n1986_8322.t0 3.61217
R23058 a_n1986_8322.n0 a_n1986_8322.t17 3.61217
R23059 a_n1986_8322.n0 a_n1986_8322.t12 3.61217
R23060 a_n1986_8322.n2 a_n1986_8322.t15 3.61217
R23061 a_n1986_8322.n2 a_n1986_8322.t14 3.61217
R23062 a_n1986_8322.n18 a_n1986_8322.t10 3.61217
R23063 a_n1986_8322.t19 a_n1986_8322.n18 3.61217
R23064 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R23065 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R23066 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R23067 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R23068 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R23069 a_n1986_8322.n17 a_n1986_8322.n14 0.358259
R23070 a_n1986_8322.n17 a_n1986_8322.n16 0.358259
R23071 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R23072 a_n1986_8322.t20 a_n1986_8322.t21 0.057021
R23073 diffpairibias.n0 diffpairibias.t18 436.822
R23074 diffpairibias.n21 diffpairibias.t19 435.479
R23075 diffpairibias.n20 diffpairibias.t16 435.479
R23076 diffpairibias.n19 diffpairibias.t17 435.479
R23077 diffpairibias.n18 diffpairibias.t21 435.479
R23078 diffpairibias.n0 diffpairibias.t22 435.479
R23079 diffpairibias.n1 diffpairibias.t20 435.479
R23080 diffpairibias.n2 diffpairibias.t23 435.479
R23081 diffpairibias.n10 diffpairibias.t0 377.536
R23082 diffpairibias.n10 diffpairibias.t8 376.193
R23083 diffpairibias.n11 diffpairibias.t10 376.193
R23084 diffpairibias.n12 diffpairibias.t6 376.193
R23085 diffpairibias.n13 diffpairibias.t2 376.193
R23086 diffpairibias.n14 diffpairibias.t12 376.193
R23087 diffpairibias.n15 diffpairibias.t4 376.193
R23088 diffpairibias.n16 diffpairibias.t14 376.193
R23089 diffpairibias.n3 diffpairibias.t1 113.368
R23090 diffpairibias.n3 diffpairibias.t9 112.698
R23091 diffpairibias.n4 diffpairibias.t11 112.698
R23092 diffpairibias.n5 diffpairibias.t7 112.698
R23093 diffpairibias.n6 diffpairibias.t3 112.698
R23094 diffpairibias.n7 diffpairibias.t13 112.698
R23095 diffpairibias.n8 diffpairibias.t5 112.698
R23096 diffpairibias.n9 diffpairibias.t15 112.698
R23097 diffpairibias.n17 diffpairibias.n16 4.77242
R23098 diffpairibias.n17 diffpairibias.n9 4.30807
R23099 diffpairibias.n18 diffpairibias.n17 4.13945
R23100 diffpairibias.n16 diffpairibias.n15 1.34352
R23101 diffpairibias.n15 diffpairibias.n14 1.34352
R23102 diffpairibias.n14 diffpairibias.n13 1.34352
R23103 diffpairibias.n13 diffpairibias.n12 1.34352
R23104 diffpairibias.n12 diffpairibias.n11 1.34352
R23105 diffpairibias.n11 diffpairibias.n10 1.34352
R23106 diffpairibias.n2 diffpairibias.n1 1.34352
R23107 diffpairibias.n1 diffpairibias.n0 1.34352
R23108 diffpairibias.n19 diffpairibias.n18 1.34352
R23109 diffpairibias.n20 diffpairibias.n19 1.34352
R23110 diffpairibias.n21 diffpairibias.n20 1.34352
R23111 diffpairibias.n22 diffpairibias.n21 0.862419
R23112 diffpairibias diffpairibias.n22 0.684875
R23113 diffpairibias.n9 diffpairibias.n8 0.672012
R23114 diffpairibias.n8 diffpairibias.n7 0.672012
R23115 diffpairibias.n7 diffpairibias.n6 0.672012
R23116 diffpairibias.n6 diffpairibias.n5 0.672012
R23117 diffpairibias.n5 diffpairibias.n4 0.672012
R23118 diffpairibias.n4 diffpairibias.n3 0.672012
R23119 diffpairibias.n22 diffpairibias.n2 0.190907
C0 CSoutput outputibias 0.032386f
C1 vdd CSoutput 0.140836p
C2 minus diffpairibias 4.33e-19
C3 commonsourceibias output 0.006808f
C4 vdd plus 0.093192f
C5 CSoutput minus 2.38478f
C6 plus diffpairibias 4.56e-19
C7 commonsourceibias outputibias 0.003832f
C8 vdd commonsourceibias 0.004218f
C9 CSoutput plus 0.854911f
C10 commonsourceibias diffpairibias 0.06482f
C11 CSoutput commonsourceibias 41.846302f
C12 minus plus 9.21292f
C13 minus commonsourceibias 0.460231f
C14 plus commonsourceibias 0.415048f
C15 output outputibias 2.34152f
C16 vdd output 7.23429f
C17 CSoutput output 6.13881f
C18 diffpairibias gnd 48.980137f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.144047p
C22 plus gnd 34.995f
C23 minus gnd 27.488161f
C24 CSoutput gnd 0.106364p
C25 vdd gnd 0.438396p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 a_n1986_8322.t21 gnd 49.3579f
C74 a_n1986_8322.t20 gnd 74.7673f
C75 a_n1986_8322.t10 gnd 0.093533f
C76 a_n1986_8322.t9 gnd 0.875792f
C77 a_n1986_8322.t17 gnd 0.093533f
C78 a_n1986_8322.t12 gnd 0.093533f
C79 a_n1986_8322.n0 gnd 0.658844f
C80 a_n1986_8322.n1 gnd 0.736161f
C81 a_n1986_8322.t15 gnd 0.093533f
C82 a_n1986_8322.t14 gnd 0.093533f
C83 a_n1986_8322.n2 gnd 0.658844f
C84 a_n1986_8322.n3 gnd 0.374034f
C85 a_n1986_8322.t8 gnd 0.874048f
C86 a_n1986_8322.n4 gnd 1.39896f
C87 a_n1986_8322.t3 gnd 0.875792f
C88 a_n1986_8322.t7 gnd 0.093533f
C89 a_n1986_8322.t6 gnd 0.093533f
C90 a_n1986_8322.n5 gnd 0.658844f
C91 a_n1986_8322.n6 gnd 0.736161f
C92 a_n1986_8322.t1 gnd 0.874048f
C93 a_n1986_8322.n7 gnd 0.370446f
C94 a_n1986_8322.t4 gnd 0.874048f
C95 a_n1986_8322.n8 gnd 0.370446f
C96 a_n1986_8322.t2 gnd 0.093533f
C97 a_n1986_8322.t0 gnd 0.093533f
C98 a_n1986_8322.n9 gnd 0.658844f
C99 a_n1986_8322.n10 gnd 0.374034f
C100 a_n1986_8322.t5 gnd 0.874048f
C101 a_n1986_8322.n11 gnd 0.872317f
C102 a_n1986_8322.n12 gnd 1.59071f
C103 a_n1986_8322.n13 gnd 3.20172f
C104 a_n1986_8322.t11 gnd 0.874048f
C105 a_n1986_8322.n14 gnd 0.76652f
C106 a_n1986_8322.t18 gnd 0.875789f
C107 a_n1986_8322.t16 gnd 0.093533f
C108 a_n1986_8322.t13 gnd 0.093533f
C109 a_n1986_8322.n15 gnd 0.658844f
C110 a_n1986_8322.n16 gnd 0.736163f
C111 a_n1986_8322.n17 gnd 0.374032f
C112 a_n1986_8322.n18 gnd 0.658845f
C113 a_n1986_8322.t19 gnd 0.093533f
C114 output.t4 gnd 0.464308f
C115 output.t10 gnd 0.044422f
C116 output.t14 gnd 0.044422f
C117 output.n0 gnd 0.364624f
C118 output.n1 gnd 0.614102f
C119 output.t1 gnd 0.044422f
C120 output.t6 gnd 0.044422f
C121 output.n2 gnd 0.364624f
C122 output.n3 gnd 0.350265f
C123 output.t7 gnd 0.044422f
C124 output.t12 gnd 0.044422f
C125 output.n4 gnd 0.364624f
C126 output.n5 gnd 0.350265f
C127 output.t0 gnd 0.044422f
C128 output.t8 gnd 0.044422f
C129 output.n6 gnd 0.364624f
C130 output.n7 gnd 0.350265f
C131 output.t11 gnd 0.044422f
C132 output.t9 gnd 0.044422f
C133 output.n8 gnd 0.364624f
C134 output.n9 gnd 0.350265f
C135 output.t15 gnd 0.044422f
C136 output.t2 gnd 0.044422f
C137 output.n10 gnd 0.364624f
C138 output.n11 gnd 0.350265f
C139 output.t3 gnd 0.044422f
C140 output.t13 gnd 0.044422f
C141 output.n12 gnd 0.364624f
C142 output.n13 gnd 0.350265f
C143 output.t5 gnd 0.462979f
C144 output.n14 gnd 0.28994f
C145 output.n15 gnd 0.015803f
C146 output.n16 gnd 0.011243f
C147 output.n17 gnd 0.006041f
C148 output.n18 gnd 0.01428f
C149 output.n19 gnd 0.006397f
C150 output.n20 gnd 0.011243f
C151 output.n21 gnd 0.006041f
C152 output.n22 gnd 0.01428f
C153 output.n23 gnd 0.006397f
C154 output.n24 gnd 0.048111f
C155 output.t18 gnd 0.023274f
C156 output.n25 gnd 0.01071f
C157 output.n26 gnd 0.008435f
C158 output.n27 gnd 0.006041f
C159 output.n28 gnd 0.267512f
C160 output.n29 gnd 0.011243f
C161 output.n30 gnd 0.006041f
C162 output.n31 gnd 0.006397f
C163 output.n32 gnd 0.01428f
C164 output.n33 gnd 0.01428f
C165 output.n34 gnd 0.006397f
C166 output.n35 gnd 0.006041f
C167 output.n36 gnd 0.011243f
C168 output.n37 gnd 0.011243f
C169 output.n38 gnd 0.006041f
C170 output.n39 gnd 0.006397f
C171 output.n40 gnd 0.01428f
C172 output.n41 gnd 0.030913f
C173 output.n42 gnd 0.006397f
C174 output.n43 gnd 0.006041f
C175 output.n44 gnd 0.025987f
C176 output.n45 gnd 0.097665f
C177 output.n46 gnd 0.015803f
C178 output.n47 gnd 0.011243f
C179 output.n48 gnd 0.006041f
C180 output.n49 gnd 0.01428f
C181 output.n50 gnd 0.006397f
C182 output.n51 gnd 0.011243f
C183 output.n52 gnd 0.006041f
C184 output.n53 gnd 0.01428f
C185 output.n54 gnd 0.006397f
C186 output.n55 gnd 0.048111f
C187 output.t17 gnd 0.023274f
C188 output.n56 gnd 0.01071f
C189 output.n57 gnd 0.008435f
C190 output.n58 gnd 0.006041f
C191 output.n59 gnd 0.267512f
C192 output.n60 gnd 0.011243f
C193 output.n61 gnd 0.006041f
C194 output.n62 gnd 0.006397f
C195 output.n63 gnd 0.01428f
C196 output.n64 gnd 0.01428f
C197 output.n65 gnd 0.006397f
C198 output.n66 gnd 0.006041f
C199 output.n67 gnd 0.011243f
C200 output.n68 gnd 0.011243f
C201 output.n69 gnd 0.006041f
C202 output.n70 gnd 0.006397f
C203 output.n71 gnd 0.01428f
C204 output.n72 gnd 0.030913f
C205 output.n73 gnd 0.006397f
C206 output.n74 gnd 0.006041f
C207 output.n75 gnd 0.025987f
C208 output.n76 gnd 0.09306f
C209 output.n77 gnd 1.65264f
C210 output.n78 gnd 0.015803f
C211 output.n79 gnd 0.011243f
C212 output.n80 gnd 0.006041f
C213 output.n81 gnd 0.01428f
C214 output.n82 gnd 0.006397f
C215 output.n83 gnd 0.011243f
C216 output.n84 gnd 0.006041f
C217 output.n85 gnd 0.01428f
C218 output.n86 gnd 0.006397f
C219 output.n87 gnd 0.048111f
C220 output.t19 gnd 0.023274f
C221 output.n88 gnd 0.01071f
C222 output.n89 gnd 0.008435f
C223 output.n90 gnd 0.006041f
C224 output.n91 gnd 0.267512f
C225 output.n92 gnd 0.011243f
C226 output.n93 gnd 0.006041f
C227 output.n94 gnd 0.006397f
C228 output.n95 gnd 0.01428f
C229 output.n96 gnd 0.01428f
C230 output.n97 gnd 0.006397f
C231 output.n98 gnd 0.006041f
C232 output.n99 gnd 0.011243f
C233 output.n100 gnd 0.011243f
C234 output.n101 gnd 0.006041f
C235 output.n102 gnd 0.006397f
C236 output.n103 gnd 0.01428f
C237 output.n104 gnd 0.030913f
C238 output.n105 gnd 0.006397f
C239 output.n106 gnd 0.006041f
C240 output.n107 gnd 0.025987f
C241 output.n108 gnd 0.09306f
C242 output.n109 gnd 0.713089f
C243 output.n110 gnd 0.015803f
C244 output.n111 gnd 0.011243f
C245 output.n112 gnd 0.006041f
C246 output.n113 gnd 0.01428f
C247 output.n114 gnd 0.006397f
C248 output.n115 gnd 0.011243f
C249 output.n116 gnd 0.006041f
C250 output.n117 gnd 0.01428f
C251 output.n118 gnd 0.006397f
C252 output.n119 gnd 0.048111f
C253 output.t16 gnd 0.023274f
C254 output.n120 gnd 0.01071f
C255 output.n121 gnd 0.008435f
C256 output.n122 gnd 0.006041f
C257 output.n123 gnd 0.267512f
C258 output.n124 gnd 0.011243f
C259 output.n125 gnd 0.006041f
C260 output.n126 gnd 0.006397f
C261 output.n127 gnd 0.01428f
C262 output.n128 gnd 0.01428f
C263 output.n129 gnd 0.006397f
C264 output.n130 gnd 0.006041f
C265 output.n131 gnd 0.011243f
C266 output.n132 gnd 0.011243f
C267 output.n133 gnd 0.006041f
C268 output.n134 gnd 0.006397f
C269 output.n135 gnd 0.01428f
C270 output.n136 gnd 0.030913f
C271 output.n137 gnd 0.006397f
C272 output.n138 gnd 0.006041f
C273 output.n139 gnd 0.025987f
C274 output.n140 gnd 0.09306f
C275 output.n141 gnd 1.67353f
C276 outputibias.t10 gnd 0.11477f
C277 outputibias.t9 gnd 0.115567f
C278 outputibias.n0 gnd 0.130108f
C279 outputibias.n1 gnd 0.001372f
C280 outputibias.n2 gnd 9.76e-19
C281 outputibias.n3 gnd 5.24e-19
C282 outputibias.n4 gnd 0.001239f
C283 outputibias.n5 gnd 5.55e-19
C284 outputibias.n6 gnd 9.76e-19
C285 outputibias.n7 gnd 5.24e-19
C286 outputibias.n8 gnd 0.001239f
C287 outputibias.n9 gnd 5.55e-19
C288 outputibias.n10 gnd 0.004176f
C289 outputibias.t5 gnd 0.00202f
C290 outputibias.n11 gnd 9.3e-19
C291 outputibias.n12 gnd 7.32e-19
C292 outputibias.n13 gnd 5.24e-19
C293 outputibias.n14 gnd 0.02322f
C294 outputibias.n15 gnd 9.76e-19
C295 outputibias.n16 gnd 5.24e-19
C296 outputibias.n17 gnd 5.55e-19
C297 outputibias.n18 gnd 0.001239f
C298 outputibias.n19 gnd 0.001239f
C299 outputibias.n20 gnd 5.55e-19
C300 outputibias.n21 gnd 5.24e-19
C301 outputibias.n22 gnd 9.76e-19
C302 outputibias.n23 gnd 9.76e-19
C303 outputibias.n24 gnd 5.24e-19
C304 outputibias.n25 gnd 5.55e-19
C305 outputibias.n26 gnd 0.001239f
C306 outputibias.n27 gnd 0.002683f
C307 outputibias.n28 gnd 5.55e-19
C308 outputibias.n29 gnd 5.24e-19
C309 outputibias.n30 gnd 0.002256f
C310 outputibias.n31 gnd 0.005781f
C311 outputibias.n32 gnd 0.001372f
C312 outputibias.n33 gnd 9.76e-19
C313 outputibias.n34 gnd 5.24e-19
C314 outputibias.n35 gnd 0.001239f
C315 outputibias.n36 gnd 5.55e-19
C316 outputibias.n37 gnd 9.76e-19
C317 outputibias.n38 gnd 5.24e-19
C318 outputibias.n39 gnd 0.001239f
C319 outputibias.n40 gnd 5.55e-19
C320 outputibias.n41 gnd 0.004176f
C321 outputibias.t7 gnd 0.00202f
C322 outputibias.n42 gnd 9.3e-19
C323 outputibias.n43 gnd 7.32e-19
C324 outputibias.n44 gnd 5.24e-19
C325 outputibias.n45 gnd 0.02322f
C326 outputibias.n46 gnd 9.76e-19
C327 outputibias.n47 gnd 5.24e-19
C328 outputibias.n48 gnd 5.55e-19
C329 outputibias.n49 gnd 0.001239f
C330 outputibias.n50 gnd 0.001239f
C331 outputibias.n51 gnd 5.55e-19
C332 outputibias.n52 gnd 5.24e-19
C333 outputibias.n53 gnd 9.76e-19
C334 outputibias.n54 gnd 9.76e-19
C335 outputibias.n55 gnd 5.24e-19
C336 outputibias.n56 gnd 5.55e-19
C337 outputibias.n57 gnd 0.001239f
C338 outputibias.n58 gnd 0.002683f
C339 outputibias.n59 gnd 5.55e-19
C340 outputibias.n60 gnd 5.24e-19
C341 outputibias.n61 gnd 0.002256f
C342 outputibias.n62 gnd 0.005197f
C343 outputibias.n63 gnd 0.121892f
C344 outputibias.n64 gnd 0.001372f
C345 outputibias.n65 gnd 9.76e-19
C346 outputibias.n66 gnd 5.24e-19
C347 outputibias.n67 gnd 0.001239f
C348 outputibias.n68 gnd 5.55e-19
C349 outputibias.n69 gnd 9.76e-19
C350 outputibias.n70 gnd 5.24e-19
C351 outputibias.n71 gnd 0.001239f
C352 outputibias.n72 gnd 5.55e-19
C353 outputibias.n73 gnd 0.004176f
C354 outputibias.t1 gnd 0.00202f
C355 outputibias.n74 gnd 9.3e-19
C356 outputibias.n75 gnd 7.32e-19
C357 outputibias.n76 gnd 5.24e-19
C358 outputibias.n77 gnd 0.02322f
C359 outputibias.n78 gnd 9.76e-19
C360 outputibias.n79 gnd 5.24e-19
C361 outputibias.n80 gnd 5.55e-19
C362 outputibias.n81 gnd 0.001239f
C363 outputibias.n82 gnd 0.001239f
C364 outputibias.n83 gnd 5.55e-19
C365 outputibias.n84 gnd 5.24e-19
C366 outputibias.n85 gnd 9.76e-19
C367 outputibias.n86 gnd 9.76e-19
C368 outputibias.n87 gnd 5.24e-19
C369 outputibias.n88 gnd 5.55e-19
C370 outputibias.n89 gnd 0.001239f
C371 outputibias.n90 gnd 0.002683f
C372 outputibias.n91 gnd 5.55e-19
C373 outputibias.n92 gnd 5.24e-19
C374 outputibias.n93 gnd 0.002256f
C375 outputibias.n94 gnd 0.005197f
C376 outputibias.n95 gnd 0.064513f
C377 outputibias.n96 gnd 0.001372f
C378 outputibias.n97 gnd 9.76e-19
C379 outputibias.n98 gnd 5.24e-19
C380 outputibias.n99 gnd 0.001239f
C381 outputibias.n100 gnd 5.55e-19
C382 outputibias.n101 gnd 9.76e-19
C383 outputibias.n102 gnd 5.24e-19
C384 outputibias.n103 gnd 0.001239f
C385 outputibias.n104 gnd 5.55e-19
C386 outputibias.n105 gnd 0.004176f
C387 outputibias.t3 gnd 0.00202f
C388 outputibias.n106 gnd 9.3e-19
C389 outputibias.n107 gnd 7.32e-19
C390 outputibias.n108 gnd 5.24e-19
C391 outputibias.n109 gnd 0.02322f
C392 outputibias.n110 gnd 9.76e-19
C393 outputibias.n111 gnd 5.24e-19
C394 outputibias.n112 gnd 5.55e-19
C395 outputibias.n113 gnd 0.001239f
C396 outputibias.n114 gnd 0.001239f
C397 outputibias.n115 gnd 5.55e-19
C398 outputibias.n116 gnd 5.24e-19
C399 outputibias.n117 gnd 9.76e-19
C400 outputibias.n118 gnd 9.76e-19
C401 outputibias.n119 gnd 5.24e-19
C402 outputibias.n120 gnd 5.55e-19
C403 outputibias.n121 gnd 0.001239f
C404 outputibias.n122 gnd 0.002683f
C405 outputibias.n123 gnd 5.55e-19
C406 outputibias.n124 gnd 5.24e-19
C407 outputibias.n125 gnd 0.002256f
C408 outputibias.n126 gnd 0.005197f
C409 outputibias.n127 gnd 0.084814f
C410 outputibias.t2 gnd 0.108319f
C411 outputibias.t0 gnd 0.108319f
C412 outputibias.t6 gnd 0.108319f
C413 outputibias.t4 gnd 0.109238f
C414 outputibias.n128 gnd 0.134674f
C415 outputibias.n129 gnd 0.07244f
C416 outputibias.n130 gnd 0.079818f
C417 outputibias.n131 gnd 0.164901f
C418 outputibias.t11 gnd 0.11477f
C419 outputibias.n132 gnd 0.067481f
C420 outputibias.t8 gnd 0.11477f
C421 outputibias.n133 gnd 0.065115f
C422 outputibias.n134 gnd 0.029159f
C423 minus.n0 gnd 0.033059f
C424 minus.n1 gnd 0.007502f
C425 minus.n2 gnd 0.033059f
C426 minus.n3 gnd 0.007502f
C427 minus.n4 gnd 0.033059f
C428 minus.n5 gnd 0.007502f
C429 minus.n6 gnd 0.033059f
C430 minus.n7 gnd 0.007502f
C431 minus.n8 gnd 0.033059f
C432 minus.n9 gnd 0.007502f
C433 minus.t8 gnd 0.484567f
C434 minus.t7 gnd 0.467594f
C435 minus.n10 gnd 0.214486f
C436 minus.n11 gnd 0.192507f
C437 minus.n12 gnd 0.142322f
C438 minus.n13 gnd 0.033059f
C439 minus.t11 gnd 0.467594f
C440 minus.n14 gnd 0.20772f
C441 minus.n15 gnd 0.007502f
C442 minus.t10 gnd 0.467594f
C443 minus.n16 gnd 0.20772f
C444 minus.n17 gnd 0.033059f
C445 minus.n18 gnd 0.033059f
C446 minus.n19 gnd 0.033059f
C447 minus.t12 gnd 0.467594f
C448 minus.n20 gnd 0.20772f
C449 minus.n21 gnd 0.007502f
C450 minus.t20 gnd 0.467594f
C451 minus.n22 gnd 0.20772f
C452 minus.n23 gnd 0.033059f
C453 minus.n24 gnd 0.033059f
C454 minus.n25 gnd 0.033059f
C455 minus.t18 gnd 0.467594f
C456 minus.n26 gnd 0.20772f
C457 minus.n27 gnd 0.007502f
C458 minus.t25 gnd 0.467594f
C459 minus.n28 gnd 0.20772f
C460 minus.n29 gnd 0.033059f
C461 minus.n30 gnd 0.033059f
C462 minus.n31 gnd 0.033059f
C463 minus.t24 gnd 0.467594f
C464 minus.n32 gnd 0.20772f
C465 minus.n33 gnd 0.007502f
C466 minus.t14 gnd 0.467594f
C467 minus.n34 gnd 0.20772f
C468 minus.n35 gnd 0.033059f
C469 minus.n36 gnd 0.033059f
C470 minus.n37 gnd 0.033059f
C471 minus.t22 gnd 0.467594f
C472 minus.n38 gnd 0.20772f
C473 minus.n39 gnd 0.007502f
C474 minus.t19 gnd 0.467594f
C475 minus.n40 gnd 0.208026f
C476 minus.n41 gnd 0.38286f
C477 minus.n42 gnd 0.033059f
C478 minus.t13 gnd 0.467594f
C479 minus.t15 gnd 0.467594f
C480 minus.n43 gnd 0.033059f
C481 minus.t5 gnd 0.467594f
C482 minus.n44 gnd 0.20772f
C483 minus.n45 gnd 0.033059f
C484 minus.t6 gnd 0.467594f
C485 minus.t26 gnd 0.467594f
C486 minus.n46 gnd 0.20772f
C487 minus.n47 gnd 0.033059f
C488 minus.t21 gnd 0.467594f
C489 minus.t23 gnd 0.467594f
C490 minus.n48 gnd 0.20772f
C491 minus.n49 gnd 0.033059f
C492 minus.t16 gnd 0.467594f
C493 minus.t17 gnd 0.467594f
C494 minus.n50 gnd 0.20772f
C495 minus.n51 gnd 0.033059f
C496 minus.t9 gnd 0.467594f
C497 minus.t27 gnd 0.467594f
C498 minus.n52 gnd 0.214486f
C499 minus.t28 gnd 0.484567f
C500 minus.n53 gnd 0.192507f
C501 minus.n54 gnd 0.142322f
C502 minus.n55 gnd 0.007502f
C503 minus.n56 gnd 0.20772f
C504 minus.n57 gnd 0.007502f
C505 minus.n58 gnd 0.033059f
C506 minus.n59 gnd 0.033059f
C507 minus.n60 gnd 0.033059f
C508 minus.n61 gnd 0.007502f
C509 minus.n62 gnd 0.20772f
C510 minus.n63 gnd 0.007502f
C511 minus.n64 gnd 0.033059f
C512 minus.n65 gnd 0.033059f
C513 minus.n66 gnd 0.033059f
C514 minus.n67 gnd 0.007502f
C515 minus.n68 gnd 0.20772f
C516 minus.n69 gnd 0.007502f
C517 minus.n70 gnd 0.033059f
C518 minus.n71 gnd 0.033059f
C519 minus.n72 gnd 0.033059f
C520 minus.n73 gnd 0.007502f
C521 minus.n74 gnd 0.20772f
C522 minus.n75 gnd 0.007502f
C523 minus.n76 gnd 0.033059f
C524 minus.n77 gnd 0.033059f
C525 minus.n78 gnd 0.033059f
C526 minus.n79 gnd 0.007502f
C527 minus.n80 gnd 0.20772f
C528 minus.n81 gnd 0.007502f
C529 minus.n82 gnd 0.208026f
C530 minus.n83 gnd 1.10752f
C531 minus.n84 gnd 1.65019f
C532 minus.t1 gnd 0.010191f
C533 minus.t0 gnd 0.010191f
C534 minus.n85 gnd 0.033511f
C535 minus.t4 gnd 0.010191f
C536 minus.t3 gnd 0.010191f
C537 minus.n86 gnd 0.033052f
C538 minus.n87 gnd 0.282084f
C539 minus.t2 gnd 0.056723f
C540 minus.n88 gnd 0.15393f
C541 minus.n89 gnd 1.77478f
C542 a_n1808_13878.t7 gnd 0.185195f
C543 a_n1808_13878.t2 gnd 0.185195f
C544 a_n1808_13878.t4 gnd 0.185195f
C545 a_n1808_13878.n0 gnd 1.4598f
C546 a_n1808_13878.t8 gnd 0.185195f
C547 a_n1808_13878.t3 gnd 0.185195f
C548 a_n1808_13878.n1 gnd 1.45825f
C549 a_n1808_13878.n2 gnd 2.03762f
C550 a_n1808_13878.t6 gnd 0.185195f
C551 a_n1808_13878.t1 gnd 0.185195f
C552 a_n1808_13878.n3 gnd 1.45825f
C553 a_n1808_13878.n4 gnd 3.69301f
C554 a_n1808_13878.t13 gnd 1.73408f
C555 a_n1808_13878.t16 gnd 0.185195f
C556 a_n1808_13878.t17 gnd 0.185195f
C557 a_n1808_13878.n5 gnd 1.30452f
C558 a_n1808_13878.n6 gnd 1.4576f
C559 a_n1808_13878.t12 gnd 1.73062f
C560 a_n1808_13878.n7 gnd 0.733487f
C561 a_n1808_13878.t15 gnd 1.73062f
C562 a_n1808_13878.n8 gnd 0.733487f
C563 a_n1808_13878.t18 gnd 0.185195f
C564 a_n1808_13878.t19 gnd 0.185195f
C565 a_n1808_13878.n9 gnd 1.30452f
C566 a_n1808_13878.n10 gnd 0.74059f
C567 a_n1808_13878.t14 gnd 1.73062f
C568 a_n1808_13878.n11 gnd 1.7272f
C569 a_n1808_13878.n12 gnd 2.51438f
C570 a_n1808_13878.t9 gnd 0.185195f
C571 a_n1808_13878.t10 gnd 0.185195f
C572 a_n1808_13878.n13 gnd 1.45825f
C573 a_n1808_13878.n14 gnd 1.80025f
C574 a_n1808_13878.t0 gnd 0.185195f
C575 a_n1808_13878.t5 gnd 0.185195f
C576 a_n1808_13878.n15 gnd 1.45825f
C577 a_n1808_13878.n16 gnd 1.31079f
C578 a_n1808_13878.n17 gnd 1.46067f
C579 a_n1808_13878.t11 gnd 0.185195f
C580 a_n2408_n452.n0 gnd 3.99939f
C581 a_n2408_n452.n1 gnd 2.94086f
C582 a_n2408_n452.n2 gnd 3.93642f
C583 a_n2408_n452.n3 gnd 0.830148f
C584 a_n2408_n452.n4 gnd 0.83015f
C585 a_n2408_n452.n5 gnd 0.532573f
C586 a_n2408_n452.n6 gnd 0.207439f
C587 a_n2408_n452.n7 gnd 0.152783f
C588 a_n2408_n452.n8 gnd 0.240126f
C589 a_n2408_n452.n9 gnd 0.18547f
C590 a_n2408_n452.n10 gnd 0.207439f
C591 a_n2408_n452.n11 gnd 1.0188f
C592 a_n2408_n452.n12 gnd 0.152783f
C593 a_n2408_n452.n13 gnd 0.587229f
C594 a_n2408_n452.n14 gnd 0.43766f
C595 a_n2408_n452.n15 gnd 0.218625f
C596 a_n2408_n452.n16 gnd 0.49859f
C597 a_n2408_n452.n17 gnd 0.286021f
C598 a_n2408_n452.n18 gnd 0.443934f
C599 a_n2408_n452.n19 gnd 0.218625f
C600 a_n2408_n452.n20 gnd 0.740623f
C601 a_n2408_n452.n21 gnd 0.286021f
C602 a_n2408_n452.n22 gnd 0.49859f
C603 a_n2408_n452.n23 gnd 0.67269f
C604 a_n2408_n452.n24 gnd 0.218625f
C605 a_n2408_n452.n25 gnd 0.286021f
C606 a_n2408_n452.n26 gnd 3.36354f
C607 a_n2408_n452.n27 gnd 0.286021f
C608 a_n2408_n452.n28 gnd 0.647141f
C609 a_n2408_n452.n29 gnd 0.286021f
C610 a_n2408_n452.n30 gnd 1.19351f
C611 a_n2408_n452.n31 gnd 1.93948f
C612 a_n2408_n452.n32 gnd 1.1588f
C613 a_n2408_n452.n33 gnd 1.79991f
C614 a_n2408_n452.n34 gnd 0.004526f
C615 a_n2408_n452.n35 gnd 0.008464f
C616 a_n2408_n452.n37 gnd 0.289215f
C617 a_n2408_n452.n38 gnd 0.008464f
C618 a_n2408_n452.n40 gnd 0.289215f
C619 a_n2408_n452.n41 gnd 0.008464f
C620 a_n2408_n452.n43 gnd 0.289215f
C621 a_n2408_n452.n44 gnd 0.008464f
C622 a_n2408_n452.n45 gnd 0.288804f
C623 a_n2408_n452.n46 gnd 0.008464f
C624 a_n2408_n452.n47 gnd 0.288804f
C625 a_n2408_n452.n48 gnd 0.008464f
C626 a_n2408_n452.n49 gnd 0.288804f
C627 a_n2408_n452.n50 gnd 0.008464f
C628 a_n2408_n452.n51 gnd 0.288804f
C629 a_n2408_n452.n52 gnd 0.310121f
C630 a_n2408_n452.t12 gnd 0.151641f
C631 a_n2408_n452.t21 gnd 0.720216f
C632 a_n2408_n452.t19 gnd 0.70536f
C633 a_n2408_n452.t25 gnd 0.70536f
C634 a_n2408_n452.t11 gnd 0.70536f
C635 a_n2408_n452.t17 gnd 0.720216f
C636 a_n2408_n452.t74 gnd 0.720216f
C637 a_n2408_n452.t57 gnd 0.70536f
C638 a_n2408_n452.t61 gnd 0.70536f
C639 a_n2408_n452.t51 gnd 0.70536f
C640 a_n2408_n452.n53 gnd 0.310121f
C641 a_n2408_n452.t66 gnd 0.70536f
C642 a_n2408_n452.t72 gnd 0.717022f
C643 a_n2408_n452.t30 gnd 1.41989f
C644 a_n2408_n452.t32 gnd 0.151641f
C645 a_n2408_n452.t16 gnd 0.151641f
C646 a_n2408_n452.n54 gnd 1.06816f
C647 a_n2408_n452.t28 gnd 0.151641f
C648 a_n2408_n452.t24 gnd 0.151641f
C649 a_n2408_n452.n55 gnd 1.06816f
C650 a_n2408_n452.t14 gnd 1.41706f
C651 a_n2408_n452.t27 gnd 0.70536f
C652 a_n2408_n452.n56 gnd 0.310121f
C653 a_n2408_n452.t23 gnd 0.70536f
C654 a_n2408_n452.t31 gnd 0.70536f
C655 a_n2408_n452.t56 gnd 0.70536f
C656 a_n2408_n452.n57 gnd 0.310121f
C657 a_n2408_n452.t65 gnd 0.70536f
C658 a_n2408_n452.t70 gnd 0.70536f
C659 a_n2408_n452.t69 gnd 0.720216f
C660 a_n2408_n452.n58 gnd 0.31277f
C661 a_n2408_n452.t49 gnd 0.70536f
C662 a_n2408_n452.n59 gnd 0.306183f
C663 a_n2408_n452.n60 gnd 0.312771f
C664 a_n2408_n452.t50 gnd 0.717022f
C665 a_n2408_n452.t29 gnd 0.720216f
C666 a_n2408_n452.n61 gnd 0.31277f
C667 a_n2408_n452.t15 gnd 0.70536f
C668 a_n2408_n452.n62 gnd 0.306183f
C669 a_n2408_n452.n63 gnd 0.312771f
C670 a_n2408_n452.t13 gnd 0.717022f
C671 a_n2408_n452.n64 gnd 1.1461f
C672 a_n2408_n452.t54 gnd 0.70536f
C673 a_n2408_n452.n65 gnd 0.306183f
C674 a_n2408_n452.t60 gnd 0.70536f
C675 a_n2408_n452.n66 gnd 0.306183f
C676 a_n2408_n452.t52 gnd 0.70536f
C677 a_n2408_n452.n67 gnd 0.306183f
C678 a_n2408_n452.t64 gnd 0.70536f
C679 a_n2408_n452.n68 gnd 0.306183f
C680 a_n2408_n452.t55 gnd 0.70536f
C681 a_n2408_n452.n69 gnd 0.300622f
C682 a_n2408_n452.t75 gnd 0.70536f
C683 a_n2408_n452.n70 gnd 0.310121f
C684 a_n2408_n452.t58 gnd 0.717179f
C685 a_n2408_n452.t67 gnd 0.70536f
C686 a_n2408_n452.n71 gnd 0.300622f
C687 a_n2408_n452.t53 gnd 0.70536f
C688 a_n2408_n452.n72 gnd 0.310121f
C689 a_n2408_n452.t62 gnd 0.717179f
C690 a_n2408_n452.t71 gnd 0.70536f
C691 a_n2408_n452.n73 gnd 0.300622f
C692 a_n2408_n452.t59 gnd 0.70536f
C693 a_n2408_n452.n74 gnd 0.310121f
C694 a_n2408_n452.t73 gnd 0.717179f
C695 a_n2408_n452.t63 gnd 0.70536f
C696 a_n2408_n452.n75 gnd 0.300622f
C697 a_n2408_n452.t48 gnd 0.70536f
C698 a_n2408_n452.n76 gnd 0.310121f
C699 a_n2408_n452.t68 gnd 0.717179f
C700 a_n2408_n452.n77 gnd 1.35508f
C701 a_n2408_n452.n78 gnd 0.312771f
C702 a_n2408_n452.n79 gnd 0.306183f
C703 a_n2408_n452.n80 gnd 0.31277f
C704 a_n2408_n452.t9 gnd 0.70536f
C705 a_n2408_n452.n81 gnd 0.312771f
C706 a_n2408_n452.t39 gnd 0.117943f
C707 a_n2408_n452.t35 gnd 0.117943f
C708 a_n2408_n452.n82 gnd 1.0445f
C709 a_n2408_n452.t41 gnd 0.117943f
C710 a_n2408_n452.t8 gnd 0.117943f
C711 a_n2408_n452.n83 gnd 1.04218f
C712 a_n2408_n452.t2 gnd 0.117943f
C713 a_n2408_n452.t1 gnd 0.117943f
C714 a_n2408_n452.n84 gnd 1.04218f
C715 a_n2408_n452.t46 gnd 0.117943f
C716 a_n2408_n452.t7 gnd 0.117943f
C717 a_n2408_n452.n85 gnd 1.0445f
C718 a_n2408_n452.t6 gnd 0.117943f
C719 a_n2408_n452.t38 gnd 0.117943f
C720 a_n2408_n452.n86 gnd 1.04218f
C721 a_n2408_n452.t5 gnd 0.117943f
C722 a_n2408_n452.t4 gnd 0.117943f
C723 a_n2408_n452.n87 gnd 1.04218f
C724 a_n2408_n452.t45 gnd 0.117943f
C725 a_n2408_n452.t3 gnd 0.117943f
C726 a_n2408_n452.n88 gnd 1.04218f
C727 a_n2408_n452.t34 gnd 0.117943f
C728 a_n2408_n452.t42 gnd 0.117943f
C729 a_n2408_n452.n89 gnd 1.04218f
C730 a_n2408_n452.t37 gnd 0.117943f
C731 a_n2408_n452.t43 gnd 0.117943f
C732 a_n2408_n452.n90 gnd 1.04218f
C733 a_n2408_n452.t0 gnd 0.117943f
C734 a_n2408_n452.t36 gnd 0.117943f
C735 a_n2408_n452.n91 gnd 1.0445f
C736 a_n2408_n452.t44 gnd 0.117943f
C737 a_n2408_n452.t47 gnd 0.117943f
C738 a_n2408_n452.n92 gnd 1.04218f
C739 a_n2408_n452.t40 gnd 0.117943f
C740 a_n2408_n452.t33 gnd 0.117943f
C741 a_n2408_n452.n93 gnd 1.04218f
C742 a_n2408_n452.n94 gnd 0.310121f
C743 a_n2408_n452.n95 gnd 0.31277f
C744 a_n2408_n452.n96 gnd 0.796711f
C745 a_n2408_n452.t22 gnd 1.41706f
C746 a_n2408_n452.t20 gnd 0.151641f
C747 a_n2408_n452.t26 gnd 0.151641f
C748 a_n2408_n452.n97 gnd 1.06816f
C749 a_n2408_n452.t18 gnd 1.41989f
C750 a_n2408_n452.n98 gnd 1.06816f
C751 a_n2408_n452.t10 gnd 0.151641f
C752 commonsourceibias.n0 gnd 0.012292f
C753 commonsourceibias.t89 gnd 0.186134f
C754 commonsourceibias.t51 gnd 0.172107f
C755 commonsourceibias.n1 gnd 0.068671f
C756 commonsourceibias.n2 gnd 0.009212f
C757 commonsourceibias.t95 gnd 0.172107f
C758 commonsourceibias.n3 gnd 0.007452f
C759 commonsourceibias.n4 gnd 0.009212f
C760 commonsourceibias.t90 gnd 0.172107f
C761 commonsourceibias.n5 gnd 0.008893f
C762 commonsourceibias.n6 gnd 0.009212f
C763 commonsourceibias.t101 gnd 0.172107f
C764 commonsourceibias.n7 gnd 0.068671f
C765 commonsourceibias.t86 gnd 0.172107f
C766 commonsourceibias.n8 gnd 0.00744f
C767 commonsourceibias.n9 gnd 0.012292f
C768 commonsourceibias.t8 gnd 0.186134f
C769 commonsourceibias.t38 gnd 0.172107f
C770 commonsourceibias.n10 gnd 0.068671f
C771 commonsourceibias.n11 gnd 0.009212f
C772 commonsourceibias.t0 gnd 0.172107f
C773 commonsourceibias.n12 gnd 0.007452f
C774 commonsourceibias.n13 gnd 0.009212f
C775 commonsourceibias.t6 gnd 0.172107f
C776 commonsourceibias.n14 gnd 0.008893f
C777 commonsourceibias.n15 gnd 0.009212f
C778 commonsourceibias.t44 gnd 0.172107f
C779 commonsourceibias.n16 gnd 0.068671f
C780 commonsourceibias.t12 gnd 0.172107f
C781 commonsourceibias.n17 gnd 0.00744f
C782 commonsourceibias.n18 gnd 0.009212f
C783 commonsourceibias.t20 gnd 0.172107f
C784 commonsourceibias.t2 gnd 0.172107f
C785 commonsourceibias.n19 gnd 0.068671f
C786 commonsourceibias.n20 gnd 0.009212f
C787 commonsourceibias.t10 gnd 0.172107f
C788 commonsourceibias.n21 gnd 0.068671f
C789 commonsourceibias.n22 gnd 0.009212f
C790 commonsourceibias.t34 gnd 0.172107f
C791 commonsourceibias.n23 gnd 0.068671f
C792 commonsourceibias.n24 gnd 0.046375f
C793 commonsourceibias.t16 gnd 0.172107f
C794 commonsourceibias.t22 gnd 0.194203f
C795 commonsourceibias.n25 gnd 0.079692f
C796 commonsourceibias.n26 gnd 0.082502f
C797 commonsourceibias.n27 gnd 0.011354f
C798 commonsourceibias.n28 gnd 0.012561f
C799 commonsourceibias.n29 gnd 0.009212f
C800 commonsourceibias.n30 gnd 0.009212f
C801 commonsourceibias.n31 gnd 0.012479f
C802 commonsourceibias.n32 gnd 0.007452f
C803 commonsourceibias.n33 gnd 0.012633f
C804 commonsourceibias.n34 gnd 0.009212f
C805 commonsourceibias.n35 gnd 0.009212f
C806 commonsourceibias.n36 gnd 0.01271f
C807 commonsourceibias.n37 gnd 0.01096f
C808 commonsourceibias.n38 gnd 0.008893f
C809 commonsourceibias.n39 gnd 0.009212f
C810 commonsourceibias.n40 gnd 0.009212f
C811 commonsourceibias.n41 gnd 0.011268f
C812 commonsourceibias.n42 gnd 0.012647f
C813 commonsourceibias.n43 gnd 0.068671f
C814 commonsourceibias.n44 gnd 0.012562f
C815 commonsourceibias.n45 gnd 0.009212f
C816 commonsourceibias.n46 gnd 0.009212f
C817 commonsourceibias.n47 gnd 0.009212f
C818 commonsourceibias.n48 gnd 0.012562f
C819 commonsourceibias.n49 gnd 0.068671f
C820 commonsourceibias.n50 gnd 0.012647f
C821 commonsourceibias.n51 gnd 0.011268f
C822 commonsourceibias.n52 gnd 0.009212f
C823 commonsourceibias.n53 gnd 0.009212f
C824 commonsourceibias.n54 gnd 0.009212f
C825 commonsourceibias.n55 gnd 0.01096f
C826 commonsourceibias.n56 gnd 0.01271f
C827 commonsourceibias.n57 gnd 0.068671f
C828 commonsourceibias.n58 gnd 0.012633f
C829 commonsourceibias.n59 gnd 0.009212f
C830 commonsourceibias.n60 gnd 0.009212f
C831 commonsourceibias.n61 gnd 0.009212f
C832 commonsourceibias.n62 gnd 0.012479f
C833 commonsourceibias.n63 gnd 0.068671f
C834 commonsourceibias.n64 gnd 0.012561f
C835 commonsourceibias.n65 gnd 0.011354f
C836 commonsourceibias.n66 gnd 0.009212f
C837 commonsourceibias.n67 gnd 0.009212f
C838 commonsourceibias.n68 gnd 0.009345f
C839 commonsourceibias.n69 gnd 0.009661f
C840 commonsourceibias.n70 gnd 0.082165f
C841 commonsourceibias.n71 gnd 0.09115f
C842 commonsourceibias.t9 gnd 0.019878f
C843 commonsourceibias.t39 gnd 0.019878f
C844 commonsourceibias.n72 gnd 0.175652f
C845 commonsourceibias.n73 gnd 0.151777f
C846 commonsourceibias.t1 gnd 0.019878f
C847 commonsourceibias.t7 gnd 0.019878f
C848 commonsourceibias.n74 gnd 0.175652f
C849 commonsourceibias.n75 gnd 0.080684f
C850 commonsourceibias.t45 gnd 0.019878f
C851 commonsourceibias.t13 gnd 0.019878f
C852 commonsourceibias.n76 gnd 0.175652f
C853 commonsourceibias.n77 gnd 0.067408f
C854 commonsourceibias.t17 gnd 0.019878f
C855 commonsourceibias.t23 gnd 0.019878f
C856 commonsourceibias.n78 gnd 0.17624f
C857 commonsourceibias.t11 gnd 0.019878f
C858 commonsourceibias.t35 gnd 0.019878f
C859 commonsourceibias.n79 gnd 0.175652f
C860 commonsourceibias.n80 gnd 0.163675f
C861 commonsourceibias.t21 gnd 0.019878f
C862 commonsourceibias.t3 gnd 0.019878f
C863 commonsourceibias.n81 gnd 0.175652f
C864 commonsourceibias.n82 gnd 0.067408f
C865 commonsourceibias.n83 gnd 0.081623f
C866 commonsourceibias.n84 gnd 0.009212f
C867 commonsourceibias.t77 gnd 0.172107f
C868 commonsourceibias.t94 gnd 0.172107f
C869 commonsourceibias.n85 gnd 0.068671f
C870 commonsourceibias.n86 gnd 0.009212f
C871 commonsourceibias.t87 gnd 0.172107f
C872 commonsourceibias.n87 gnd 0.068671f
C873 commonsourceibias.n88 gnd 0.009212f
C874 commonsourceibias.t58 gnd 0.172107f
C875 commonsourceibias.n89 gnd 0.068671f
C876 commonsourceibias.n90 gnd 0.046375f
C877 commonsourceibias.t80 gnd 0.172107f
C878 commonsourceibias.t73 gnd 0.194203f
C879 commonsourceibias.n91 gnd 0.079692f
C880 commonsourceibias.n92 gnd 0.082502f
C881 commonsourceibias.n93 gnd 0.011354f
C882 commonsourceibias.n94 gnd 0.012561f
C883 commonsourceibias.n95 gnd 0.009212f
C884 commonsourceibias.n96 gnd 0.009212f
C885 commonsourceibias.n97 gnd 0.012479f
C886 commonsourceibias.n98 gnd 0.007452f
C887 commonsourceibias.n99 gnd 0.012633f
C888 commonsourceibias.n100 gnd 0.009212f
C889 commonsourceibias.n101 gnd 0.009212f
C890 commonsourceibias.n102 gnd 0.01271f
C891 commonsourceibias.n103 gnd 0.01096f
C892 commonsourceibias.n104 gnd 0.008893f
C893 commonsourceibias.n105 gnd 0.009212f
C894 commonsourceibias.n106 gnd 0.009212f
C895 commonsourceibias.n107 gnd 0.011268f
C896 commonsourceibias.n108 gnd 0.012647f
C897 commonsourceibias.n109 gnd 0.068671f
C898 commonsourceibias.n110 gnd 0.012562f
C899 commonsourceibias.n111 gnd 0.009168f
C900 commonsourceibias.n112 gnd 0.066591f
C901 commonsourceibias.n113 gnd 0.009168f
C902 commonsourceibias.n114 gnd 0.012562f
C903 commonsourceibias.n115 gnd 0.068671f
C904 commonsourceibias.n116 gnd 0.012647f
C905 commonsourceibias.n117 gnd 0.011268f
C906 commonsourceibias.n118 gnd 0.009212f
C907 commonsourceibias.n119 gnd 0.009212f
C908 commonsourceibias.n120 gnd 0.009212f
C909 commonsourceibias.n121 gnd 0.01096f
C910 commonsourceibias.n122 gnd 0.01271f
C911 commonsourceibias.n123 gnd 0.068671f
C912 commonsourceibias.n124 gnd 0.012633f
C913 commonsourceibias.n125 gnd 0.009212f
C914 commonsourceibias.n126 gnd 0.009212f
C915 commonsourceibias.n127 gnd 0.009212f
C916 commonsourceibias.n128 gnd 0.012479f
C917 commonsourceibias.n129 gnd 0.068671f
C918 commonsourceibias.n130 gnd 0.012561f
C919 commonsourceibias.n131 gnd 0.011354f
C920 commonsourceibias.n132 gnd 0.009212f
C921 commonsourceibias.n133 gnd 0.009212f
C922 commonsourceibias.n134 gnd 0.009345f
C923 commonsourceibias.n135 gnd 0.009661f
C924 commonsourceibias.n136 gnd 0.082165f
C925 commonsourceibias.n137 gnd 0.053193f
C926 commonsourceibias.n138 gnd 0.012292f
C927 commonsourceibias.t54 gnd 0.186134f
C928 commonsourceibias.t119 gnd 0.172107f
C929 commonsourceibias.n139 gnd 0.068671f
C930 commonsourceibias.n140 gnd 0.009212f
C931 commonsourceibias.t110 gnd 0.172107f
C932 commonsourceibias.n141 gnd 0.007452f
C933 commonsourceibias.n142 gnd 0.009212f
C934 commonsourceibias.t60 gnd 0.172107f
C935 commonsourceibias.n143 gnd 0.008893f
C936 commonsourceibias.n144 gnd 0.009212f
C937 commonsourceibias.t117 gnd 0.172107f
C938 commonsourceibias.n145 gnd 0.068671f
C939 commonsourceibias.t65 gnd 0.172107f
C940 commonsourceibias.n146 gnd 0.00744f
C941 commonsourceibias.n147 gnd 0.009212f
C942 commonsourceibias.t59 gnd 0.172107f
C943 commonsourceibias.t118 gnd 0.172107f
C944 commonsourceibias.n148 gnd 0.068671f
C945 commonsourceibias.n149 gnd 0.009212f
C946 commonsourceibias.t71 gnd 0.172107f
C947 commonsourceibias.n150 gnd 0.068671f
C948 commonsourceibias.n151 gnd 0.009212f
C949 commonsourceibias.t83 gnd 0.172107f
C950 commonsourceibias.n152 gnd 0.068671f
C951 commonsourceibias.n153 gnd 0.046375f
C952 commonsourceibias.t116 gnd 0.172107f
C953 commonsourceibias.t70 gnd 0.194203f
C954 commonsourceibias.n154 gnd 0.079692f
C955 commonsourceibias.n155 gnd 0.082502f
C956 commonsourceibias.n156 gnd 0.011354f
C957 commonsourceibias.n157 gnd 0.012561f
C958 commonsourceibias.n158 gnd 0.009212f
C959 commonsourceibias.n159 gnd 0.009212f
C960 commonsourceibias.n160 gnd 0.012479f
C961 commonsourceibias.n161 gnd 0.007452f
C962 commonsourceibias.n162 gnd 0.012633f
C963 commonsourceibias.n163 gnd 0.009212f
C964 commonsourceibias.n164 gnd 0.009212f
C965 commonsourceibias.n165 gnd 0.01271f
C966 commonsourceibias.n166 gnd 0.01096f
C967 commonsourceibias.n167 gnd 0.008893f
C968 commonsourceibias.n168 gnd 0.009212f
C969 commonsourceibias.n169 gnd 0.009212f
C970 commonsourceibias.n170 gnd 0.011268f
C971 commonsourceibias.n171 gnd 0.012647f
C972 commonsourceibias.n172 gnd 0.068671f
C973 commonsourceibias.n173 gnd 0.012562f
C974 commonsourceibias.n174 gnd 0.009212f
C975 commonsourceibias.n175 gnd 0.009212f
C976 commonsourceibias.n176 gnd 0.009212f
C977 commonsourceibias.n177 gnd 0.012562f
C978 commonsourceibias.n178 gnd 0.068671f
C979 commonsourceibias.n179 gnd 0.012647f
C980 commonsourceibias.n180 gnd 0.011268f
C981 commonsourceibias.n181 gnd 0.009212f
C982 commonsourceibias.n182 gnd 0.009212f
C983 commonsourceibias.n183 gnd 0.009212f
C984 commonsourceibias.n184 gnd 0.01096f
C985 commonsourceibias.n185 gnd 0.01271f
C986 commonsourceibias.n186 gnd 0.068671f
C987 commonsourceibias.n187 gnd 0.012633f
C988 commonsourceibias.n188 gnd 0.009212f
C989 commonsourceibias.n189 gnd 0.009212f
C990 commonsourceibias.n190 gnd 0.009212f
C991 commonsourceibias.n191 gnd 0.012479f
C992 commonsourceibias.n192 gnd 0.068671f
C993 commonsourceibias.n193 gnd 0.012561f
C994 commonsourceibias.n194 gnd 0.011354f
C995 commonsourceibias.n195 gnd 0.009212f
C996 commonsourceibias.n196 gnd 0.009212f
C997 commonsourceibias.n197 gnd 0.009345f
C998 commonsourceibias.n198 gnd 0.009661f
C999 commonsourceibias.n199 gnd 0.082165f
C1000 commonsourceibias.n200 gnd 0.027962f
C1001 commonsourceibias.n201 gnd 0.146988f
C1002 commonsourceibias.n202 gnd 0.012292f
C1003 commonsourceibias.t57 gnd 0.172107f
C1004 commonsourceibias.n203 gnd 0.068671f
C1005 commonsourceibias.n204 gnd 0.009212f
C1006 commonsourceibias.t96 gnd 0.172107f
C1007 commonsourceibias.n205 gnd 0.007452f
C1008 commonsourceibias.n206 gnd 0.009212f
C1009 commonsourceibias.t93 gnd 0.172107f
C1010 commonsourceibias.n207 gnd 0.008893f
C1011 commonsourceibias.n208 gnd 0.009212f
C1012 commonsourceibias.t115 gnd 0.172107f
C1013 commonsourceibias.n209 gnd 0.068671f
C1014 commonsourceibias.t68 gnd 0.172107f
C1015 commonsourceibias.n210 gnd 0.00744f
C1016 commonsourceibias.n211 gnd 0.009212f
C1017 commonsourceibias.t88 gnd 0.172107f
C1018 commonsourceibias.t108 gnd 0.172107f
C1019 commonsourceibias.n212 gnd 0.068671f
C1020 commonsourceibias.n213 gnd 0.009212f
C1021 commonsourceibias.t103 gnd 0.172107f
C1022 commonsourceibias.n214 gnd 0.068671f
C1023 commonsourceibias.n215 gnd 0.009212f
C1024 commonsourceibias.t48 gnd 0.172107f
C1025 commonsourceibias.n216 gnd 0.068671f
C1026 commonsourceibias.n217 gnd 0.046375f
C1027 commonsourceibias.t102 gnd 0.172107f
C1028 commonsourceibias.t98 gnd 0.194203f
C1029 commonsourceibias.n218 gnd 0.079692f
C1030 commonsourceibias.n219 gnd 0.082502f
C1031 commonsourceibias.n220 gnd 0.011354f
C1032 commonsourceibias.n221 gnd 0.012561f
C1033 commonsourceibias.n222 gnd 0.009212f
C1034 commonsourceibias.n223 gnd 0.009212f
C1035 commonsourceibias.n224 gnd 0.012479f
C1036 commonsourceibias.n225 gnd 0.007452f
C1037 commonsourceibias.n226 gnd 0.012633f
C1038 commonsourceibias.n227 gnd 0.009212f
C1039 commonsourceibias.n228 gnd 0.009212f
C1040 commonsourceibias.n229 gnd 0.01271f
C1041 commonsourceibias.n230 gnd 0.01096f
C1042 commonsourceibias.n231 gnd 0.008893f
C1043 commonsourceibias.n232 gnd 0.009212f
C1044 commonsourceibias.n233 gnd 0.009212f
C1045 commonsourceibias.n234 gnd 0.011268f
C1046 commonsourceibias.n235 gnd 0.012647f
C1047 commonsourceibias.n236 gnd 0.068671f
C1048 commonsourceibias.n237 gnd 0.012562f
C1049 commonsourceibias.n238 gnd 0.009212f
C1050 commonsourceibias.n239 gnd 0.009212f
C1051 commonsourceibias.n240 gnd 0.009212f
C1052 commonsourceibias.n241 gnd 0.012562f
C1053 commonsourceibias.n242 gnd 0.068671f
C1054 commonsourceibias.n243 gnd 0.012647f
C1055 commonsourceibias.n244 gnd 0.011268f
C1056 commonsourceibias.n245 gnd 0.009212f
C1057 commonsourceibias.n246 gnd 0.009212f
C1058 commonsourceibias.n247 gnd 0.009212f
C1059 commonsourceibias.n248 gnd 0.01096f
C1060 commonsourceibias.n249 gnd 0.01271f
C1061 commonsourceibias.n250 gnd 0.068671f
C1062 commonsourceibias.n251 gnd 0.012633f
C1063 commonsourceibias.n252 gnd 0.009212f
C1064 commonsourceibias.n253 gnd 0.009212f
C1065 commonsourceibias.n254 gnd 0.009212f
C1066 commonsourceibias.n255 gnd 0.012479f
C1067 commonsourceibias.n256 gnd 0.068671f
C1068 commonsourceibias.n257 gnd 0.012561f
C1069 commonsourceibias.n258 gnd 0.011354f
C1070 commonsourceibias.n259 gnd 0.009212f
C1071 commonsourceibias.n260 gnd 0.009212f
C1072 commonsourceibias.n261 gnd 0.009345f
C1073 commonsourceibias.n262 gnd 0.009661f
C1074 commonsourceibias.t109 gnd 0.186134f
C1075 commonsourceibias.n263 gnd 0.082165f
C1076 commonsourceibias.n264 gnd 0.027962f
C1077 commonsourceibias.n265 gnd 0.437625f
C1078 commonsourceibias.n266 gnd 0.012292f
C1079 commonsourceibias.t69 gnd 0.186134f
C1080 commonsourceibias.t99 gnd 0.172107f
C1081 commonsourceibias.n267 gnd 0.068671f
C1082 commonsourceibias.n268 gnd 0.009212f
C1083 commonsourceibias.t84 gnd 0.172107f
C1084 commonsourceibias.n269 gnd 0.007452f
C1085 commonsourceibias.n270 gnd 0.009212f
C1086 commonsourceibias.t72 gnd 0.172107f
C1087 commonsourceibias.n271 gnd 0.008893f
C1088 commonsourceibias.n272 gnd 0.009212f
C1089 commonsourceibias.t66 gnd 0.172107f
C1090 commonsourceibias.n273 gnd 0.00744f
C1091 commonsourceibias.n274 gnd 0.009212f
C1092 commonsourceibias.t56 gnd 0.172107f
C1093 commonsourceibias.t79 gnd 0.172107f
C1094 commonsourceibias.n275 gnd 0.068671f
C1095 commonsourceibias.n276 gnd 0.009212f
C1096 commonsourceibias.t67 gnd 0.172107f
C1097 commonsourceibias.n277 gnd 0.068671f
C1098 commonsourceibias.n278 gnd 0.009212f
C1099 commonsourceibias.t104 gnd 0.172107f
C1100 commonsourceibias.n279 gnd 0.068671f
C1101 commonsourceibias.n280 gnd 0.046375f
C1102 commonsourceibias.t64 gnd 0.172107f
C1103 commonsourceibias.t111 gnd 0.194203f
C1104 commonsourceibias.n281 gnd 0.079692f
C1105 commonsourceibias.n282 gnd 0.082502f
C1106 commonsourceibias.n283 gnd 0.011354f
C1107 commonsourceibias.n284 gnd 0.012561f
C1108 commonsourceibias.n285 gnd 0.009212f
C1109 commonsourceibias.n286 gnd 0.009212f
C1110 commonsourceibias.n287 gnd 0.012479f
C1111 commonsourceibias.n288 gnd 0.007452f
C1112 commonsourceibias.n289 gnd 0.012633f
C1113 commonsourceibias.n290 gnd 0.009212f
C1114 commonsourceibias.n291 gnd 0.009212f
C1115 commonsourceibias.n292 gnd 0.01271f
C1116 commonsourceibias.n293 gnd 0.01096f
C1117 commonsourceibias.n294 gnd 0.008893f
C1118 commonsourceibias.n295 gnd 0.009212f
C1119 commonsourceibias.n296 gnd 0.009212f
C1120 commonsourceibias.n297 gnd 0.011268f
C1121 commonsourceibias.n298 gnd 0.012647f
C1122 commonsourceibias.n299 gnd 0.068671f
C1123 commonsourceibias.n300 gnd 0.012562f
C1124 commonsourceibias.n301 gnd 0.009168f
C1125 commonsourceibias.t41 gnd 0.019878f
C1126 commonsourceibias.t33 gnd 0.019878f
C1127 commonsourceibias.n302 gnd 0.17624f
C1128 commonsourceibias.t43 gnd 0.019878f
C1129 commonsourceibias.t29 gnd 0.019878f
C1130 commonsourceibias.n303 gnd 0.175652f
C1131 commonsourceibias.n304 gnd 0.163675f
C1132 commonsourceibias.t19 gnd 0.019878f
C1133 commonsourceibias.t37 gnd 0.019878f
C1134 commonsourceibias.n305 gnd 0.175652f
C1135 commonsourceibias.n306 gnd 0.067408f
C1136 commonsourceibias.n307 gnd 0.012292f
C1137 commonsourceibias.t46 gnd 0.172107f
C1138 commonsourceibias.n308 gnd 0.068671f
C1139 commonsourceibias.n309 gnd 0.009212f
C1140 commonsourceibias.t14 gnd 0.172107f
C1141 commonsourceibias.n310 gnd 0.007452f
C1142 commonsourceibias.n311 gnd 0.009212f
C1143 commonsourceibias.t24 gnd 0.172107f
C1144 commonsourceibias.n312 gnd 0.008893f
C1145 commonsourceibias.n313 gnd 0.009212f
C1146 commonsourceibias.t30 gnd 0.172107f
C1147 commonsourceibias.n314 gnd 0.00744f
C1148 commonsourceibias.n315 gnd 0.009212f
C1149 commonsourceibias.t36 gnd 0.172107f
C1150 commonsourceibias.t18 gnd 0.172107f
C1151 commonsourceibias.n316 gnd 0.068671f
C1152 commonsourceibias.n317 gnd 0.009212f
C1153 commonsourceibias.t28 gnd 0.172107f
C1154 commonsourceibias.n318 gnd 0.068671f
C1155 commonsourceibias.n319 gnd 0.009212f
C1156 commonsourceibias.t42 gnd 0.172107f
C1157 commonsourceibias.n320 gnd 0.068671f
C1158 commonsourceibias.n321 gnd 0.046375f
C1159 commonsourceibias.t32 gnd 0.172107f
C1160 commonsourceibias.t40 gnd 0.194203f
C1161 commonsourceibias.n322 gnd 0.079692f
C1162 commonsourceibias.n323 gnd 0.082502f
C1163 commonsourceibias.n324 gnd 0.011354f
C1164 commonsourceibias.n325 gnd 0.012561f
C1165 commonsourceibias.n326 gnd 0.009212f
C1166 commonsourceibias.n327 gnd 0.009212f
C1167 commonsourceibias.n328 gnd 0.012479f
C1168 commonsourceibias.n329 gnd 0.007452f
C1169 commonsourceibias.n330 gnd 0.012633f
C1170 commonsourceibias.n331 gnd 0.009212f
C1171 commonsourceibias.n332 gnd 0.009212f
C1172 commonsourceibias.n333 gnd 0.01271f
C1173 commonsourceibias.n334 gnd 0.01096f
C1174 commonsourceibias.n335 gnd 0.008893f
C1175 commonsourceibias.n336 gnd 0.009212f
C1176 commonsourceibias.n337 gnd 0.009212f
C1177 commonsourceibias.n338 gnd 0.011268f
C1178 commonsourceibias.n339 gnd 0.012647f
C1179 commonsourceibias.n340 gnd 0.068671f
C1180 commonsourceibias.n341 gnd 0.012562f
C1181 commonsourceibias.n342 gnd 0.009212f
C1182 commonsourceibias.n343 gnd 0.009212f
C1183 commonsourceibias.n344 gnd 0.009212f
C1184 commonsourceibias.n345 gnd 0.012562f
C1185 commonsourceibias.n346 gnd 0.068671f
C1186 commonsourceibias.n347 gnd 0.012647f
C1187 commonsourceibias.t4 gnd 0.172107f
C1188 commonsourceibias.n348 gnd 0.068671f
C1189 commonsourceibias.n349 gnd 0.011268f
C1190 commonsourceibias.n350 gnd 0.009212f
C1191 commonsourceibias.n351 gnd 0.009212f
C1192 commonsourceibias.n352 gnd 0.009212f
C1193 commonsourceibias.n353 gnd 0.01096f
C1194 commonsourceibias.n354 gnd 0.01271f
C1195 commonsourceibias.n355 gnd 0.068671f
C1196 commonsourceibias.n356 gnd 0.012633f
C1197 commonsourceibias.n357 gnd 0.009212f
C1198 commonsourceibias.n358 gnd 0.009212f
C1199 commonsourceibias.n359 gnd 0.009212f
C1200 commonsourceibias.n360 gnd 0.012479f
C1201 commonsourceibias.n361 gnd 0.068671f
C1202 commonsourceibias.n362 gnd 0.012561f
C1203 commonsourceibias.n363 gnd 0.011354f
C1204 commonsourceibias.n364 gnd 0.009212f
C1205 commonsourceibias.n365 gnd 0.009212f
C1206 commonsourceibias.n366 gnd 0.009345f
C1207 commonsourceibias.n367 gnd 0.009661f
C1208 commonsourceibias.t26 gnd 0.186134f
C1209 commonsourceibias.n368 gnd 0.082165f
C1210 commonsourceibias.n369 gnd 0.09115f
C1211 commonsourceibias.t47 gnd 0.019878f
C1212 commonsourceibias.t27 gnd 0.019878f
C1213 commonsourceibias.n370 gnd 0.175652f
C1214 commonsourceibias.n371 gnd 0.151777f
C1215 commonsourceibias.t25 gnd 0.019878f
C1216 commonsourceibias.t15 gnd 0.019878f
C1217 commonsourceibias.n372 gnd 0.175652f
C1218 commonsourceibias.n373 gnd 0.080684f
C1219 commonsourceibias.t31 gnd 0.019878f
C1220 commonsourceibias.t5 gnd 0.019878f
C1221 commonsourceibias.n374 gnd 0.175652f
C1222 commonsourceibias.n375 gnd 0.067408f
C1223 commonsourceibias.n376 gnd 0.081623f
C1224 commonsourceibias.n377 gnd 0.066591f
C1225 commonsourceibias.n378 gnd 0.009168f
C1226 commonsourceibias.n379 gnd 0.012562f
C1227 commonsourceibias.n380 gnd 0.068671f
C1228 commonsourceibias.n381 gnd 0.012647f
C1229 commonsourceibias.t92 gnd 0.172107f
C1230 commonsourceibias.n382 gnd 0.068671f
C1231 commonsourceibias.n383 gnd 0.011268f
C1232 commonsourceibias.n384 gnd 0.009212f
C1233 commonsourceibias.n385 gnd 0.009212f
C1234 commonsourceibias.n386 gnd 0.009212f
C1235 commonsourceibias.n387 gnd 0.01096f
C1236 commonsourceibias.n388 gnd 0.01271f
C1237 commonsourceibias.n389 gnd 0.068671f
C1238 commonsourceibias.n390 gnd 0.012633f
C1239 commonsourceibias.n391 gnd 0.009212f
C1240 commonsourceibias.n392 gnd 0.009212f
C1241 commonsourceibias.n393 gnd 0.009212f
C1242 commonsourceibias.n394 gnd 0.012479f
C1243 commonsourceibias.n395 gnd 0.068671f
C1244 commonsourceibias.n396 gnd 0.012561f
C1245 commonsourceibias.n397 gnd 0.011354f
C1246 commonsourceibias.n398 gnd 0.009212f
C1247 commonsourceibias.n399 gnd 0.009212f
C1248 commonsourceibias.n400 gnd 0.009345f
C1249 commonsourceibias.n401 gnd 0.009661f
C1250 commonsourceibias.n402 gnd 0.082165f
C1251 commonsourceibias.n403 gnd 0.053193f
C1252 commonsourceibias.n404 gnd 0.012292f
C1253 commonsourceibias.t107 gnd 0.172107f
C1254 commonsourceibias.n405 gnd 0.068671f
C1255 commonsourceibias.n406 gnd 0.009212f
C1256 commonsourceibias.t50 gnd 0.172107f
C1257 commonsourceibias.n407 gnd 0.007452f
C1258 commonsourceibias.n408 gnd 0.009212f
C1259 commonsourceibias.t114 gnd 0.172107f
C1260 commonsourceibias.n409 gnd 0.008893f
C1261 commonsourceibias.n410 gnd 0.009212f
C1262 commonsourceibias.t49 gnd 0.172107f
C1263 commonsourceibias.n411 gnd 0.00744f
C1264 commonsourceibias.n412 gnd 0.009212f
C1265 commonsourceibias.t74 gnd 0.172107f
C1266 commonsourceibias.t105 gnd 0.172107f
C1267 commonsourceibias.n413 gnd 0.068671f
C1268 commonsourceibias.n414 gnd 0.009212f
C1269 commonsourceibias.t55 gnd 0.172107f
C1270 commonsourceibias.n415 gnd 0.068671f
C1271 commonsourceibias.n416 gnd 0.009212f
C1272 commonsourceibias.t75 gnd 0.172107f
C1273 commonsourceibias.n417 gnd 0.068671f
C1274 commonsourceibias.n418 gnd 0.046375f
C1275 commonsourceibias.t61 gnd 0.172107f
C1276 commonsourceibias.t52 gnd 0.194203f
C1277 commonsourceibias.n419 gnd 0.079692f
C1278 commonsourceibias.n420 gnd 0.082502f
C1279 commonsourceibias.n421 gnd 0.011354f
C1280 commonsourceibias.n422 gnd 0.012561f
C1281 commonsourceibias.n423 gnd 0.009212f
C1282 commonsourceibias.n424 gnd 0.009212f
C1283 commonsourceibias.n425 gnd 0.012479f
C1284 commonsourceibias.n426 gnd 0.007452f
C1285 commonsourceibias.n427 gnd 0.012633f
C1286 commonsourceibias.n428 gnd 0.009212f
C1287 commonsourceibias.n429 gnd 0.009212f
C1288 commonsourceibias.n430 gnd 0.01271f
C1289 commonsourceibias.n431 gnd 0.01096f
C1290 commonsourceibias.n432 gnd 0.008893f
C1291 commonsourceibias.n433 gnd 0.009212f
C1292 commonsourceibias.n434 gnd 0.009212f
C1293 commonsourceibias.n435 gnd 0.011268f
C1294 commonsourceibias.n436 gnd 0.012647f
C1295 commonsourceibias.n437 gnd 0.068671f
C1296 commonsourceibias.n438 gnd 0.012562f
C1297 commonsourceibias.n439 gnd 0.009212f
C1298 commonsourceibias.n440 gnd 0.009212f
C1299 commonsourceibias.n441 gnd 0.009212f
C1300 commonsourceibias.n442 gnd 0.012562f
C1301 commonsourceibias.n443 gnd 0.068671f
C1302 commonsourceibias.n444 gnd 0.012647f
C1303 commonsourceibias.t106 gnd 0.172107f
C1304 commonsourceibias.n445 gnd 0.068671f
C1305 commonsourceibias.n446 gnd 0.011268f
C1306 commonsourceibias.n447 gnd 0.009212f
C1307 commonsourceibias.n448 gnd 0.009212f
C1308 commonsourceibias.n449 gnd 0.009212f
C1309 commonsourceibias.n450 gnd 0.01096f
C1310 commonsourceibias.n451 gnd 0.01271f
C1311 commonsourceibias.n452 gnd 0.068671f
C1312 commonsourceibias.n453 gnd 0.012633f
C1313 commonsourceibias.n454 gnd 0.009212f
C1314 commonsourceibias.n455 gnd 0.009212f
C1315 commonsourceibias.n456 gnd 0.009212f
C1316 commonsourceibias.n457 gnd 0.012479f
C1317 commonsourceibias.n458 gnd 0.068671f
C1318 commonsourceibias.n459 gnd 0.012561f
C1319 commonsourceibias.n460 gnd 0.011354f
C1320 commonsourceibias.n461 gnd 0.009212f
C1321 commonsourceibias.n462 gnd 0.009212f
C1322 commonsourceibias.n463 gnd 0.009345f
C1323 commonsourceibias.n464 gnd 0.009661f
C1324 commonsourceibias.t112 gnd 0.186134f
C1325 commonsourceibias.n465 gnd 0.082165f
C1326 commonsourceibias.n466 gnd 0.027962f
C1327 commonsourceibias.n467 gnd 0.146988f
C1328 commonsourceibias.n468 gnd 0.012292f
C1329 commonsourceibias.t81 gnd 0.172107f
C1330 commonsourceibias.n469 gnd 0.068671f
C1331 commonsourceibias.n470 gnd 0.009212f
C1332 commonsourceibias.t91 gnd 0.172107f
C1333 commonsourceibias.n471 gnd 0.007452f
C1334 commonsourceibias.n472 gnd 0.009212f
C1335 commonsourceibias.t100 gnd 0.172107f
C1336 commonsourceibias.n473 gnd 0.008893f
C1337 commonsourceibias.n474 gnd 0.009212f
C1338 commonsourceibias.t85 gnd 0.172107f
C1339 commonsourceibias.n475 gnd 0.00744f
C1340 commonsourceibias.n476 gnd 0.009212f
C1341 commonsourceibias.t82 gnd 0.172107f
C1342 commonsourceibias.t62 gnd 0.172107f
C1343 commonsourceibias.n477 gnd 0.068671f
C1344 commonsourceibias.n478 gnd 0.009212f
C1345 commonsourceibias.t53 gnd 0.172107f
C1346 commonsourceibias.n479 gnd 0.068671f
C1347 commonsourceibias.n480 gnd 0.009212f
C1348 commonsourceibias.t78 gnd 0.172107f
C1349 commonsourceibias.n481 gnd 0.068671f
C1350 commonsourceibias.n482 gnd 0.046375f
C1351 commonsourceibias.t97 gnd 0.172107f
C1352 commonsourceibias.t113 gnd 0.194203f
C1353 commonsourceibias.n483 gnd 0.079692f
C1354 commonsourceibias.n484 gnd 0.082502f
C1355 commonsourceibias.n485 gnd 0.011354f
C1356 commonsourceibias.n486 gnd 0.012561f
C1357 commonsourceibias.n487 gnd 0.009212f
C1358 commonsourceibias.n488 gnd 0.009212f
C1359 commonsourceibias.n489 gnd 0.012479f
C1360 commonsourceibias.n490 gnd 0.007452f
C1361 commonsourceibias.n491 gnd 0.012633f
C1362 commonsourceibias.n492 gnd 0.009212f
C1363 commonsourceibias.n493 gnd 0.009212f
C1364 commonsourceibias.n494 gnd 0.01271f
C1365 commonsourceibias.n495 gnd 0.01096f
C1366 commonsourceibias.n496 gnd 0.008893f
C1367 commonsourceibias.n497 gnd 0.009212f
C1368 commonsourceibias.n498 gnd 0.009212f
C1369 commonsourceibias.n499 gnd 0.011268f
C1370 commonsourceibias.n500 gnd 0.012647f
C1371 commonsourceibias.n501 gnd 0.068671f
C1372 commonsourceibias.n502 gnd 0.012562f
C1373 commonsourceibias.n503 gnd 0.009212f
C1374 commonsourceibias.n504 gnd 0.009212f
C1375 commonsourceibias.n505 gnd 0.009212f
C1376 commonsourceibias.n506 gnd 0.012562f
C1377 commonsourceibias.n507 gnd 0.068671f
C1378 commonsourceibias.n508 gnd 0.012647f
C1379 commonsourceibias.t76 gnd 0.172107f
C1380 commonsourceibias.n509 gnd 0.068671f
C1381 commonsourceibias.n510 gnd 0.011268f
C1382 commonsourceibias.n511 gnd 0.009212f
C1383 commonsourceibias.n512 gnd 0.009212f
C1384 commonsourceibias.n513 gnd 0.009212f
C1385 commonsourceibias.n514 gnd 0.01096f
C1386 commonsourceibias.n515 gnd 0.01271f
C1387 commonsourceibias.n516 gnd 0.068671f
C1388 commonsourceibias.n517 gnd 0.012633f
C1389 commonsourceibias.n518 gnd 0.009212f
C1390 commonsourceibias.n519 gnd 0.009212f
C1391 commonsourceibias.n520 gnd 0.009212f
C1392 commonsourceibias.n521 gnd 0.012479f
C1393 commonsourceibias.n522 gnd 0.068671f
C1394 commonsourceibias.n523 gnd 0.012561f
C1395 commonsourceibias.n524 gnd 0.011354f
C1396 commonsourceibias.n525 gnd 0.009212f
C1397 commonsourceibias.n526 gnd 0.009212f
C1398 commonsourceibias.n527 gnd 0.009345f
C1399 commonsourceibias.n528 gnd 0.009661f
C1400 commonsourceibias.t63 gnd 0.186134f
C1401 commonsourceibias.n529 gnd 0.082165f
C1402 commonsourceibias.n530 gnd 0.027962f
C1403 commonsourceibias.n531 gnd 0.194173f
C1404 commonsourceibias.n532 gnd 4.69557f
C1405 CSoutput.n0 gnd 0.049151f
C1406 CSoutput.t194 gnd 0.325123f
C1407 CSoutput.n1 gnd 0.146809f
C1408 CSoutput.n2 gnd 0.049151f
C1409 CSoutput.t199 gnd 0.325123f
C1410 CSoutput.n3 gnd 0.038956f
C1411 CSoutput.n4 gnd 0.049151f
C1412 CSoutput.t211 gnd 0.325123f
C1413 CSoutput.n5 gnd 0.033592f
C1414 CSoutput.n6 gnd 0.049151f
C1415 CSoutput.t196 gnd 0.325123f
C1416 CSoutput.t204 gnd 0.325123f
C1417 CSoutput.n7 gnd 0.145209f
C1418 CSoutput.n8 gnd 0.049151f
C1419 CSoutput.t202 gnd 0.325123f
C1420 CSoutput.n9 gnd 0.032028f
C1421 CSoutput.n10 gnd 0.049151f
C1422 CSoutput.t212 gnd 0.325123f
C1423 CSoutput.t200 gnd 0.325123f
C1424 CSoutput.n11 gnd 0.145209f
C1425 CSoutput.n12 gnd 0.049151f
C1426 CSoutput.t198 gnd 0.325123f
C1427 CSoutput.n13 gnd 0.033592f
C1428 CSoutput.n14 gnd 0.049151f
C1429 CSoutput.t210 gnd 0.325123f
C1430 CSoutput.t192 gnd 0.325123f
C1431 CSoutput.n15 gnd 0.145209f
C1432 CSoutput.n16 gnd 0.049151f
C1433 CSoutput.t195 gnd 0.325123f
C1434 CSoutput.n17 gnd 0.035878f
C1435 CSoutput.t206 gnd 0.388531f
C1436 CSoutput.t209 gnd 0.325123f
C1437 CSoutput.n18 gnd 0.185376f
C1438 CSoutput.n19 gnd 0.179879f
C1439 CSoutput.n20 gnd 0.208681f
C1440 CSoutput.n21 gnd 0.049151f
C1441 CSoutput.n22 gnd 0.041022f
C1442 CSoutput.n23 gnd 0.145209f
C1443 CSoutput.n24 gnd 0.039544f
C1444 CSoutput.n25 gnd 0.038956f
C1445 CSoutput.n26 gnd 0.049151f
C1446 CSoutput.n27 gnd 0.049151f
C1447 CSoutput.n28 gnd 0.040707f
C1448 CSoutput.n29 gnd 0.034561f
C1449 CSoutput.n30 gnd 0.148442f
C1450 CSoutput.n31 gnd 0.035037f
C1451 CSoutput.n32 gnd 0.049151f
C1452 CSoutput.n33 gnd 0.049151f
C1453 CSoutput.n34 gnd 0.049151f
C1454 CSoutput.n35 gnd 0.040273f
C1455 CSoutput.n36 gnd 0.145209f
C1456 CSoutput.n37 gnd 0.038515f
C1457 CSoutput.n38 gnd 0.039985f
C1458 CSoutput.n39 gnd 0.049151f
C1459 CSoutput.n40 gnd 0.049151f
C1460 CSoutput.n41 gnd 0.041014f
C1461 CSoutput.n42 gnd 0.037486f
C1462 CSoutput.n43 gnd 0.145209f
C1463 CSoutput.n44 gnd 0.038437f
C1464 CSoutput.n45 gnd 0.049151f
C1465 CSoutput.n46 gnd 0.049151f
C1466 CSoutput.n47 gnd 0.049151f
C1467 CSoutput.n48 gnd 0.038437f
C1468 CSoutput.n49 gnd 0.145209f
C1469 CSoutput.n50 gnd 0.037486f
C1470 CSoutput.n51 gnd 0.041014f
C1471 CSoutput.n52 gnd 0.049151f
C1472 CSoutput.n53 gnd 0.049151f
C1473 CSoutput.n54 gnd 0.039985f
C1474 CSoutput.n55 gnd 0.038515f
C1475 CSoutput.n56 gnd 0.145209f
C1476 CSoutput.n57 gnd 0.040273f
C1477 CSoutput.n58 gnd 0.049151f
C1478 CSoutput.n59 gnd 0.049151f
C1479 CSoutput.n60 gnd 0.049151f
C1480 CSoutput.n61 gnd 0.035037f
C1481 CSoutput.n62 gnd 0.148442f
C1482 CSoutput.n63 gnd 0.034561f
C1483 CSoutput.t205 gnd 0.325123f
C1484 CSoutput.n64 gnd 0.145209f
C1485 CSoutput.n65 gnd 0.040707f
C1486 CSoutput.n66 gnd 0.049151f
C1487 CSoutput.n67 gnd 0.049151f
C1488 CSoutput.n68 gnd 0.049151f
C1489 CSoutput.n69 gnd 0.039544f
C1490 CSoutput.n70 gnd 0.145209f
C1491 CSoutput.n71 gnd 0.041022f
C1492 CSoutput.n72 gnd 0.035878f
C1493 CSoutput.n73 gnd 0.049151f
C1494 CSoutput.n74 gnd 0.049151f
C1495 CSoutput.n75 gnd 0.037208f
C1496 CSoutput.n76 gnd 0.022098f
C1497 CSoutput.t208 gnd 0.365299f
C1498 CSoutput.n77 gnd 0.181466f
C1499 CSoutput.n78 gnd 0.742368f
C1500 CSoutput.t165 gnd 0.061309f
C1501 CSoutput.t63 gnd 0.061309f
C1502 CSoutput.n79 gnd 0.474674f
C1503 CSoutput.t145 gnd 0.061309f
C1504 CSoutput.t115 gnd 0.061309f
C1505 CSoutput.n80 gnd 0.473828f
C1506 CSoutput.n81 gnd 0.480935f
C1507 CSoutput.t154 gnd 0.061309f
C1508 CSoutput.t91 gnd 0.061309f
C1509 CSoutput.n82 gnd 0.473828f
C1510 CSoutput.n83 gnd 0.236984f
C1511 CSoutput.t173 gnd 0.061309f
C1512 CSoutput.t108 gnd 0.061309f
C1513 CSoutput.n84 gnd 0.473828f
C1514 CSoutput.n85 gnd 0.236984f
C1515 CSoutput.t69 gnd 0.061309f
C1516 CSoutput.t124 gnd 0.061309f
C1517 CSoutput.n86 gnd 0.473828f
C1518 CSoutput.n87 gnd 0.236984f
C1519 CSoutput.t74 gnd 0.061309f
C1520 CSoutput.t100 gnd 0.061309f
C1521 CSoutput.n88 gnd 0.473828f
C1522 CSoutput.n89 gnd 0.236984f
C1523 CSoutput.t178 gnd 0.061309f
C1524 CSoutput.t117 gnd 0.061309f
C1525 CSoutput.n90 gnd 0.473828f
C1526 CSoutput.n91 gnd 0.236984f
C1527 CSoutput.t77 gnd 0.061309f
C1528 CSoutput.t161 gnd 0.061309f
C1529 CSoutput.n92 gnd 0.473828f
C1530 CSoutput.n93 gnd 0.236984f
C1531 CSoutput.t87 gnd 0.061309f
C1532 CSoutput.t136 gnd 0.061309f
C1533 CSoutput.n94 gnd 0.473828f
C1534 CSoutput.n95 gnd 0.236984f
C1535 CSoutput.t103 gnd 0.061309f
C1536 CSoutput.t125 gnd 0.061309f
C1537 CSoutput.n96 gnd 0.473828f
C1538 CSoutput.n97 gnd 0.434574f
C1539 CSoutput.t158 gnd 0.061309f
C1540 CSoutput.t156 gnd 0.061309f
C1541 CSoutput.n98 gnd 0.474674f
C1542 CSoutput.t138 gnd 0.061309f
C1543 CSoutput.t70 gnd 0.061309f
C1544 CSoutput.n99 gnd 0.473828f
C1545 CSoutput.n100 gnd 0.480935f
C1546 CSoutput.t64 gnd 0.061309f
C1547 CSoutput.t152 gnd 0.061309f
C1548 CSoutput.n101 gnd 0.473828f
C1549 CSoutput.n102 gnd 0.236984f
C1550 CSoutput.t137 gnd 0.061309f
C1551 CSoutput.t110 gnd 0.061309f
C1552 CSoutput.n103 gnd 0.473828f
C1553 CSoutput.n104 gnd 0.236984f
C1554 CSoutput.t92 gnd 0.061309f
C1555 CSoutput.t168 gnd 0.061309f
C1556 CSoutput.n105 gnd 0.473828f
C1557 CSoutput.n106 gnd 0.236984f
C1558 CSoutput.t134 gnd 0.061309f
C1559 CSoutput.t133 gnd 0.061309f
C1560 CSoutput.n107 gnd 0.473828f
C1561 CSoutput.n108 gnd 0.236984f
C1562 CSoutput.t121 gnd 0.061309f
C1563 CSoutput.t88 gnd 0.061309f
C1564 CSoutput.n109 gnd 0.473828f
C1565 CSoutput.n110 gnd 0.236984f
C1566 CSoutput.t68 gnd 0.061309f
C1567 CSoutput.t122 gnd 0.061309f
C1568 CSoutput.n111 gnd 0.473828f
C1569 CSoutput.n112 gnd 0.236984f
C1570 CSoutput.t118 gnd 0.061309f
C1571 CSoutput.t86 gnd 0.061309f
C1572 CSoutput.n113 gnd 0.473828f
C1573 CSoutput.n114 gnd 0.236984f
C1574 CSoutput.t65 gnd 0.061309f
C1575 CSoutput.t62 gnd 0.061309f
C1576 CSoutput.n115 gnd 0.473828f
C1577 CSoutput.n116 gnd 0.353403f
C1578 CSoutput.n117 gnd 0.445639f
C1579 CSoutput.t170 gnd 0.061309f
C1580 CSoutput.t169 gnd 0.061309f
C1581 CSoutput.n118 gnd 0.474674f
C1582 CSoutput.t149 gnd 0.061309f
C1583 CSoutput.t83 gnd 0.061309f
C1584 CSoutput.n119 gnd 0.473828f
C1585 CSoutput.n120 gnd 0.480935f
C1586 CSoutput.t79 gnd 0.061309f
C1587 CSoutput.t167 gnd 0.061309f
C1588 CSoutput.n121 gnd 0.473828f
C1589 CSoutput.n122 gnd 0.236984f
C1590 CSoutput.t146 gnd 0.061309f
C1591 CSoutput.t123 gnd 0.061309f
C1592 CSoutput.n123 gnd 0.473828f
C1593 CSoutput.n124 gnd 0.236984f
C1594 CSoutput.t104 gnd 0.061309f
C1595 CSoutput.t179 gnd 0.061309f
C1596 CSoutput.n125 gnd 0.473828f
C1597 CSoutput.n126 gnd 0.236984f
C1598 CSoutput.t144 gnd 0.061309f
C1599 CSoutput.t143 gnd 0.061309f
C1600 CSoutput.n127 gnd 0.473828f
C1601 CSoutput.n128 gnd 0.236984f
C1602 CSoutput.t131 gnd 0.061309f
C1603 CSoutput.t101 gnd 0.061309f
C1604 CSoutput.n129 gnd 0.473828f
C1605 CSoutput.n130 gnd 0.236984f
C1606 CSoutput.t82 gnd 0.061309f
C1607 CSoutput.t132 gnd 0.061309f
C1608 CSoutput.n131 gnd 0.473828f
C1609 CSoutput.n132 gnd 0.236984f
C1610 CSoutput.t128 gnd 0.061309f
C1611 CSoutput.t99 gnd 0.061309f
C1612 CSoutput.n133 gnd 0.473828f
C1613 CSoutput.n134 gnd 0.236984f
C1614 CSoutput.t80 gnd 0.061309f
C1615 CSoutput.t78 gnd 0.061309f
C1616 CSoutput.n135 gnd 0.473828f
C1617 CSoutput.n136 gnd 0.353403f
C1618 CSoutput.n137 gnd 0.49811f
C1619 CSoutput.n138 gnd 8.57102f
C1620 CSoutput.n140 gnd 0.869472f
C1621 CSoutput.n141 gnd 0.652104f
C1622 CSoutput.n142 gnd 0.869472f
C1623 CSoutput.n143 gnd 0.869472f
C1624 CSoutput.n144 gnd 2.34089f
C1625 CSoutput.n145 gnd 0.869472f
C1626 CSoutput.n146 gnd 0.869472f
C1627 CSoutput.t213 gnd 1.08684f
C1628 CSoutput.n147 gnd 0.869472f
C1629 CSoutput.n148 gnd 0.869472f
C1630 CSoutput.n152 gnd 0.869472f
C1631 CSoutput.n156 gnd 0.869472f
C1632 CSoutput.n157 gnd 0.869472f
C1633 CSoutput.n159 gnd 0.869472f
C1634 CSoutput.n164 gnd 0.869472f
C1635 CSoutput.n166 gnd 0.869472f
C1636 CSoutput.n167 gnd 0.869472f
C1637 CSoutput.n169 gnd 0.869472f
C1638 CSoutput.n170 gnd 0.869472f
C1639 CSoutput.n172 gnd 0.869472f
C1640 CSoutput.t201 gnd 14.5288f
C1641 CSoutput.n174 gnd 0.869472f
C1642 CSoutput.n175 gnd 0.652104f
C1643 CSoutput.n176 gnd 0.869472f
C1644 CSoutput.n177 gnd 0.869472f
C1645 CSoutput.n178 gnd 2.34089f
C1646 CSoutput.n179 gnd 0.869472f
C1647 CSoutput.n180 gnd 0.869472f
C1648 CSoutput.t197 gnd 1.08684f
C1649 CSoutput.n181 gnd 0.869472f
C1650 CSoutput.n182 gnd 0.869472f
C1651 CSoutput.n186 gnd 0.869472f
C1652 CSoutput.n190 gnd 0.869472f
C1653 CSoutput.n191 gnd 0.869472f
C1654 CSoutput.n193 gnd 0.869472f
C1655 CSoutput.n198 gnd 0.869472f
C1656 CSoutput.n200 gnd 0.869472f
C1657 CSoutput.n201 gnd 0.869472f
C1658 CSoutput.n203 gnd 0.869472f
C1659 CSoutput.n204 gnd 0.869472f
C1660 CSoutput.n206 gnd 0.869472f
C1661 CSoutput.n207 gnd 0.652104f
C1662 CSoutput.n209 gnd 0.869472f
C1663 CSoutput.n210 gnd 0.652104f
C1664 CSoutput.n211 gnd 0.869472f
C1665 CSoutput.n212 gnd 0.869472f
C1666 CSoutput.n213 gnd 2.34089f
C1667 CSoutput.n214 gnd 0.869472f
C1668 CSoutput.n215 gnd 0.869472f
C1669 CSoutput.t193 gnd 1.08684f
C1670 CSoutput.n216 gnd 0.869472f
C1671 CSoutput.n217 gnd 2.34089f
C1672 CSoutput.n219 gnd 0.869472f
C1673 CSoutput.n220 gnd 0.869472f
C1674 CSoutput.n222 gnd 0.869472f
C1675 CSoutput.n223 gnd 0.869472f
C1676 CSoutput.t203 gnd 14.292001f
C1677 CSoutput.t207 gnd 14.5288f
C1678 CSoutput.n229 gnd 2.72766f
C1679 CSoutput.n230 gnd 11.1115f
C1680 CSoutput.n231 gnd 11.5765f
C1681 CSoutput.n236 gnd 2.95479f
C1682 CSoutput.n242 gnd 0.869472f
C1683 CSoutput.n244 gnd 0.869472f
C1684 CSoutput.n246 gnd 0.869472f
C1685 CSoutput.n248 gnd 0.869472f
C1686 CSoutput.n250 gnd 0.869472f
C1687 CSoutput.n256 gnd 0.869472f
C1688 CSoutput.n263 gnd 1.59515f
C1689 CSoutput.n264 gnd 1.59515f
C1690 CSoutput.n265 gnd 0.869472f
C1691 CSoutput.n266 gnd 0.869472f
C1692 CSoutput.n268 gnd 0.652104f
C1693 CSoutput.n269 gnd 0.558469f
C1694 CSoutput.n271 gnd 0.652104f
C1695 CSoutput.n272 gnd 0.558469f
C1696 CSoutput.n273 gnd 0.652104f
C1697 CSoutput.n275 gnd 0.869472f
C1698 CSoutput.n277 gnd 2.34089f
C1699 CSoutput.n278 gnd 2.72766f
C1700 CSoutput.n279 gnd 10.2197f
C1701 CSoutput.n281 gnd 0.652104f
C1702 CSoutput.n282 gnd 1.6779f
C1703 CSoutput.n283 gnd 0.652104f
C1704 CSoutput.n285 gnd 0.869472f
C1705 CSoutput.n287 gnd 2.34089f
C1706 CSoutput.n288 gnd 5.09883f
C1707 CSoutput.t61 gnd 0.061309f
C1708 CSoutput.t164 gnd 0.061309f
C1709 CSoutput.n289 gnd 0.474674f
C1710 CSoutput.t114 gnd 0.061309f
C1711 CSoutput.t177 gnd 0.061309f
C1712 CSoutput.n290 gnd 0.473828f
C1713 CSoutput.n291 gnd 0.480934f
C1714 CSoutput.t90 gnd 0.061309f
C1715 CSoutput.t153 gnd 0.061309f
C1716 CSoutput.n292 gnd 0.473828f
C1717 CSoutput.n293 gnd 0.236984f
C1718 CSoutput.t107 gnd 0.061309f
C1719 CSoutput.t172 gnd 0.061309f
C1720 CSoutput.n294 gnd 0.473828f
C1721 CSoutput.n295 gnd 0.236984f
C1722 CSoutput.t147 gnd 0.061309f
C1723 CSoutput.t67 gnd 0.061309f
C1724 CSoutput.n296 gnd 0.473828f
C1725 CSoutput.n297 gnd 0.236984f
C1726 CSoutput.t98 gnd 0.061309f
C1727 CSoutput.t73 gnd 0.061309f
C1728 CSoutput.n298 gnd 0.473828f
C1729 CSoutput.n299 gnd 0.236984f
C1730 CSoutput.t116 gnd 0.061309f
C1731 CSoutput.t95 gnd 0.061309f
C1732 CSoutput.n300 gnd 0.473828f
C1733 CSoutput.n301 gnd 0.236984f
C1734 CSoutput.t160 gnd 0.061309f
C1735 CSoutput.t76 gnd 0.061309f
C1736 CSoutput.n302 gnd 0.473828f
C1737 CSoutput.n303 gnd 0.236984f
C1738 CSoutput.t135 gnd 0.061309f
C1739 CSoutput.t84 gnd 0.061309f
C1740 CSoutput.n304 gnd 0.473828f
C1741 CSoutput.n305 gnd 0.236984f
C1742 CSoutput.t148 gnd 0.061309f
C1743 CSoutput.t102 gnd 0.061309f
C1744 CSoutput.n306 gnd 0.473828f
C1745 CSoutput.n307 gnd 0.434574f
C1746 CSoutput.t119 gnd 0.061309f
C1747 CSoutput.t120 gnd 0.061309f
C1748 CSoutput.n308 gnd 0.474674f
C1749 CSoutput.t142 gnd 0.061309f
C1750 CSoutput.t66 gnd 0.061309f
C1751 CSoutput.n309 gnd 0.473828f
C1752 CSoutput.n310 gnd 0.480934f
C1753 CSoutput.t113 gnd 0.061309f
C1754 CSoutput.t140 gnd 0.061309f
C1755 CSoutput.n311 gnd 0.473828f
C1756 CSoutput.n312 gnd 0.236984f
C1757 CSoutput.t60 gnd 0.061309f
C1758 CSoutput.t96 gnd 0.061309f
C1759 CSoutput.n313 gnd 0.473828f
C1760 CSoutput.n314 gnd 0.236984f
C1761 CSoutput.t97 gnd 0.061309f
C1762 CSoutput.t166 gnd 0.061309f
C1763 CSoutput.n315 gnd 0.473828f
C1764 CSoutput.n316 gnd 0.236984f
C1765 CSoutput.t93 gnd 0.061309f
C1766 CSoutput.t94 gnd 0.061309f
C1767 CSoutput.n317 gnd 0.473828f
C1768 CSoutput.n318 gnd 0.236984f
C1769 CSoutput.t162 gnd 0.061309f
C1770 CSoutput.t163 gnd 0.061309f
C1771 CSoutput.n319 gnd 0.473828f
C1772 CSoutput.n320 gnd 0.236984f
C1773 CSoutput.t72 gnd 0.061309f
C1774 CSoutput.t141 gnd 0.061309f
C1775 CSoutput.n321 gnd 0.473828f
C1776 CSoutput.n322 gnd 0.236984f
C1777 CSoutput.t159 gnd 0.061309f
C1778 CSoutput.t71 gnd 0.061309f
C1779 CSoutput.n323 gnd 0.473828f
C1780 CSoutput.n324 gnd 0.236984f
C1781 CSoutput.t112 gnd 0.061309f
C1782 CSoutput.t139 gnd 0.061309f
C1783 CSoutput.n325 gnd 0.473828f
C1784 CSoutput.n326 gnd 0.353403f
C1785 CSoutput.n327 gnd 0.445639f
C1786 CSoutput.t129 gnd 0.061309f
C1787 CSoutput.t130 gnd 0.061309f
C1788 CSoutput.n328 gnd 0.474674f
C1789 CSoutput.t157 gnd 0.061309f
C1790 CSoutput.t81 gnd 0.061309f
C1791 CSoutput.n329 gnd 0.473828f
C1792 CSoutput.n330 gnd 0.480934f
C1793 CSoutput.t126 gnd 0.061309f
C1794 CSoutput.t150 gnd 0.061309f
C1795 CSoutput.n331 gnd 0.473828f
C1796 CSoutput.n332 gnd 0.236984f
C1797 CSoutput.t75 gnd 0.061309f
C1798 CSoutput.t109 gnd 0.061309f
C1799 CSoutput.n333 gnd 0.473828f
C1800 CSoutput.n334 gnd 0.236984f
C1801 CSoutput.t111 gnd 0.061309f
C1802 CSoutput.t176 gnd 0.061309f
C1803 CSoutput.n335 gnd 0.473828f
C1804 CSoutput.n336 gnd 0.236984f
C1805 CSoutput.t105 gnd 0.061309f
C1806 CSoutput.t106 gnd 0.061309f
C1807 CSoutput.n337 gnd 0.473828f
C1808 CSoutput.n338 gnd 0.236984f
C1809 CSoutput.t174 gnd 0.061309f
C1810 CSoutput.t175 gnd 0.061309f
C1811 CSoutput.n339 gnd 0.473828f
C1812 CSoutput.n340 gnd 0.236984f
C1813 CSoutput.t89 gnd 0.061309f
C1814 CSoutput.t155 gnd 0.061309f
C1815 CSoutput.n341 gnd 0.473828f
C1816 CSoutput.n342 gnd 0.236984f
C1817 CSoutput.t171 gnd 0.061309f
C1818 CSoutput.t85 gnd 0.061309f
C1819 CSoutput.n343 gnd 0.473828f
C1820 CSoutput.n344 gnd 0.236984f
C1821 CSoutput.t127 gnd 0.061309f
C1822 CSoutput.t151 gnd 0.061309f
C1823 CSoutput.n345 gnd 0.473826f
C1824 CSoutput.n346 gnd 0.353405f
C1825 CSoutput.n347 gnd 0.49811f
C1826 CSoutput.n348 gnd 12.5568f
C1827 CSoutput.t182 gnd 0.053645f
C1828 CSoutput.t24 gnd 0.053645f
C1829 CSoutput.n349 gnd 0.475615f
C1830 CSoutput.t14 gnd 0.053645f
C1831 CSoutput.t40 gnd 0.053645f
C1832 CSoutput.n350 gnd 0.474029f
C1833 CSoutput.n351 gnd 0.441706f
C1834 CSoutput.t54 gnd 0.053645f
C1835 CSoutput.t184 gnd 0.053645f
C1836 CSoutput.n352 gnd 0.474029f
C1837 CSoutput.n353 gnd 0.21774f
C1838 CSoutput.t36 gnd 0.053645f
C1839 CSoutput.t19 gnd 0.053645f
C1840 CSoutput.n354 gnd 0.474029f
C1841 CSoutput.n355 gnd 0.21774f
C1842 CSoutput.t180 gnd 0.053645f
C1843 CSoutput.t9 gnd 0.053645f
C1844 CSoutput.n356 gnd 0.474029f
C1845 CSoutput.n357 gnd 0.21774f
C1846 CSoutput.t35 gnd 0.053645f
C1847 CSoutput.t189 gnd 0.053645f
C1848 CSoutput.n358 gnd 0.474029f
C1849 CSoutput.n359 gnd 0.40161f
C1850 CSoutput.t23 gnd 0.053645f
C1851 CSoutput.t22 gnd 0.053645f
C1852 CSoutput.n360 gnd 0.475615f
C1853 CSoutput.t30 gnd 0.053645f
C1854 CSoutput.t21 gnd 0.053645f
C1855 CSoutput.n361 gnd 0.474029f
C1856 CSoutput.n362 gnd 0.441706f
C1857 CSoutput.t10 gnd 0.053645f
C1858 CSoutput.t59 gnd 0.053645f
C1859 CSoutput.n363 gnd 0.474029f
C1860 CSoutput.n364 gnd 0.21774f
C1861 CSoutput.t1 gnd 0.053645f
C1862 CSoutput.t2 gnd 0.053645f
C1863 CSoutput.n365 gnd 0.474029f
C1864 CSoutput.n366 gnd 0.21774f
C1865 CSoutput.t58 gnd 0.053645f
C1866 CSoutput.t32 gnd 0.053645f
C1867 CSoutput.n367 gnd 0.474029f
C1868 CSoutput.n368 gnd 0.21774f
C1869 CSoutput.t17 gnd 0.053645f
C1870 CSoutput.t0 gnd 0.053645f
C1871 CSoutput.n369 gnd 0.474029f
C1872 CSoutput.n370 gnd 0.330577f
C1873 CSoutput.n371 gnd 0.41696f
C1874 CSoutput.t12 gnd 0.053645f
C1875 CSoutput.t187 gnd 0.053645f
C1876 CSoutput.n372 gnd 0.475615f
C1877 CSoutput.t18 gnd 0.053645f
C1878 CSoutput.t15 gnd 0.053645f
C1879 CSoutput.n373 gnd 0.474029f
C1880 CSoutput.n374 gnd 0.441706f
C1881 CSoutput.t5 gnd 0.053645f
C1882 CSoutput.t48 gnd 0.053645f
C1883 CSoutput.n375 gnd 0.474029f
C1884 CSoutput.n376 gnd 0.21774f
C1885 CSoutput.t183 gnd 0.053645f
C1886 CSoutput.t31 gnd 0.053645f
C1887 CSoutput.n377 gnd 0.474029f
C1888 CSoutput.n378 gnd 0.21774f
C1889 CSoutput.t52 gnd 0.053645f
C1890 CSoutput.t16 gnd 0.053645f
C1891 CSoutput.n379 gnd 0.474029f
C1892 CSoutput.n380 gnd 0.21774f
C1893 CSoutput.t53 gnd 0.053645f
C1894 CSoutput.t41 gnd 0.053645f
C1895 CSoutput.n381 gnd 0.474029f
C1896 CSoutput.n382 gnd 0.330577f
C1897 CSoutput.n383 gnd 0.447749f
C1898 CSoutput.n384 gnd 12.6432f
C1899 CSoutput.t42 gnd 0.053645f
C1900 CSoutput.t8 gnd 0.053645f
C1901 CSoutput.n385 gnd 0.475615f
C1902 CSoutput.t37 gnd 0.053645f
C1903 CSoutput.t186 gnd 0.053645f
C1904 CSoutput.n386 gnd 0.474029f
C1905 CSoutput.n387 gnd 0.441706f
C1906 CSoutput.t49 gnd 0.053645f
C1907 CSoutput.t20 gnd 0.053645f
C1908 CSoutput.n388 gnd 0.474029f
C1909 CSoutput.n389 gnd 0.21774f
C1910 CSoutput.t46 gnd 0.053645f
C1911 CSoutput.t55 gnd 0.053645f
C1912 CSoutput.n390 gnd 0.474029f
C1913 CSoutput.n391 gnd 0.21774f
C1914 CSoutput.t188 gnd 0.053645f
C1915 CSoutput.t4 gnd 0.053645f
C1916 CSoutput.n392 gnd 0.474029f
C1917 CSoutput.n393 gnd 0.21774f
C1918 CSoutput.t27 gnd 0.053645f
C1919 CSoutput.t29 gnd 0.053645f
C1920 CSoutput.n394 gnd 0.474029f
C1921 CSoutput.n395 gnd 0.40161f
C1922 CSoutput.t39 gnd 0.053645f
C1923 CSoutput.t3 gnd 0.053645f
C1924 CSoutput.n396 gnd 0.475615f
C1925 CSoutput.t26 gnd 0.053645f
C1926 CSoutput.t57 gnd 0.053645f
C1927 CSoutput.n397 gnd 0.474029f
C1928 CSoutput.n398 gnd 0.441706f
C1929 CSoutput.t25 gnd 0.053645f
C1930 CSoutput.t43 gnd 0.053645f
C1931 CSoutput.n399 gnd 0.474029f
C1932 CSoutput.n400 gnd 0.21774f
C1933 CSoutput.t191 gnd 0.053645f
C1934 CSoutput.t6 gnd 0.053645f
C1935 CSoutput.n401 gnd 0.474029f
C1936 CSoutput.n402 gnd 0.21774f
C1937 CSoutput.t44 gnd 0.053645f
C1938 CSoutput.t50 gnd 0.053645f
C1939 CSoutput.n403 gnd 0.474029f
C1940 CSoutput.n404 gnd 0.21774f
C1941 CSoutput.t51 gnd 0.053645f
C1942 CSoutput.t190 gnd 0.053645f
C1943 CSoutput.n405 gnd 0.474029f
C1944 CSoutput.n406 gnd 0.330577f
C1945 CSoutput.n407 gnd 0.41696f
C1946 CSoutput.t34 gnd 0.053645f
C1947 CSoutput.t45 gnd 0.053645f
C1948 CSoutput.n408 gnd 0.475615f
C1949 CSoutput.t38 gnd 0.053645f
C1950 CSoutput.t181 gnd 0.053645f
C1951 CSoutput.n409 gnd 0.474029f
C1952 CSoutput.n410 gnd 0.441706f
C1953 CSoutput.t185 gnd 0.053645f
C1954 CSoutput.t28 gnd 0.053645f
C1955 CSoutput.n411 gnd 0.474029f
C1956 CSoutput.n412 gnd 0.21774f
C1957 CSoutput.t7 gnd 0.053645f
C1958 CSoutput.t33 gnd 0.053645f
C1959 CSoutput.n413 gnd 0.474029f
C1960 CSoutput.n414 gnd 0.21774f
C1961 CSoutput.t47 gnd 0.053645f
C1962 CSoutput.t56 gnd 0.053645f
C1963 CSoutput.n415 gnd 0.474029f
C1964 CSoutput.n416 gnd 0.21774f
C1965 CSoutput.t11 gnd 0.053645f
C1966 CSoutput.t13 gnd 0.053645f
C1967 CSoutput.n417 gnd 0.474029f
C1968 CSoutput.n418 gnd 0.330577f
C1969 CSoutput.n419 gnd 0.447749f
C1970 CSoutput.n420 gnd 7.06923f
C1971 CSoutput.n421 gnd 14.8174f
C1972 vdd.t34 gnd 0.040766f
C1973 vdd.t40 gnd 0.040766f
C1974 vdd.n0 gnd 0.321531f
C1975 vdd.t12 gnd 0.040766f
C1976 vdd.t131 gnd 0.040766f
C1977 vdd.n1 gnd 0.321f
C1978 vdd.n2 gnd 0.296023f
C1979 vdd.t21 gnd 0.040766f
C1980 vdd.t36 gnd 0.040766f
C1981 vdd.n3 gnd 0.321f
C1982 vdd.n4 gnd 0.14971f
C1983 vdd.t38 gnd 0.040766f
C1984 vdd.t27 gnd 0.040766f
C1985 vdd.n5 gnd 0.321f
C1986 vdd.n6 gnd 0.140475f
C1987 vdd.t295 gnd 0.040766f
C1988 vdd.t42 gnd 0.040766f
C1989 vdd.n7 gnd 0.321531f
C1990 vdd.t29 gnd 0.040766f
C1991 vdd.t32 gnd 0.040766f
C1992 vdd.n8 gnd 0.321f
C1993 vdd.n9 gnd 0.296023f
C1994 vdd.t133 gnd 0.040766f
C1995 vdd.t15 gnd 0.040766f
C1996 vdd.n10 gnd 0.321f
C1997 vdd.n11 gnd 0.14971f
C1998 vdd.t49 gnd 0.040766f
C1999 vdd.t45 gnd 0.040766f
C2000 vdd.n12 gnd 0.321f
C2001 vdd.n13 gnd 0.140475f
C2002 vdd.n14 gnd 0.099313f
C2003 vdd.t3 gnd 0.022648f
C2004 vdd.t4 gnd 0.022648f
C2005 vdd.n15 gnd 0.208465f
C2006 vdd.t8 gnd 0.022648f
C2007 vdd.t51 gnd 0.022648f
C2008 vdd.n16 gnd 0.207855f
C2009 vdd.n17 gnd 0.361732f
C2010 vdd.t17 gnd 0.022648f
C2011 vdd.t0 gnd 0.022648f
C2012 vdd.n18 gnd 0.207855f
C2013 vdd.n19 gnd 0.149653f
C2014 vdd.t9 gnd 0.022648f
C2015 vdd.t5 gnd 0.022648f
C2016 vdd.n20 gnd 0.208465f
C2017 vdd.t16 gnd 0.022648f
C2018 vdd.t2 gnd 0.022648f
C2019 vdd.n21 gnd 0.207855f
C2020 vdd.n22 gnd 0.361732f
C2021 vdd.t6 gnd 0.022648f
C2022 vdd.t18 gnd 0.022648f
C2023 vdd.n23 gnd 0.207855f
C2024 vdd.n24 gnd 0.149653f
C2025 vdd.t52 gnd 0.022648f
C2026 vdd.t1 gnd 0.022648f
C2027 vdd.n25 gnd 0.207855f
C2028 vdd.t53 gnd 0.022648f
C2029 vdd.t7 gnd 0.022648f
C2030 vdd.n26 gnd 0.207855f
C2031 vdd.n27 gnd 22.5395f
C2032 vdd.n28 gnd 8.528549f
C2033 vdd.n29 gnd 0.006177f
C2034 vdd.n30 gnd 0.005732f
C2035 vdd.n31 gnd 0.003171f
C2036 vdd.n32 gnd 0.00728f
C2037 vdd.n33 gnd 0.00308f
C2038 vdd.n34 gnd 0.003261f
C2039 vdd.n35 gnd 0.005732f
C2040 vdd.n36 gnd 0.00308f
C2041 vdd.n37 gnd 0.00728f
C2042 vdd.n38 gnd 0.003261f
C2043 vdd.n39 gnd 0.005732f
C2044 vdd.n40 gnd 0.00308f
C2045 vdd.n41 gnd 0.00546f
C2046 vdd.n42 gnd 0.005477f
C2047 vdd.t141 gnd 0.015641f
C2048 vdd.n43 gnd 0.034801f
C2049 vdd.n44 gnd 0.181113f
C2050 vdd.n45 gnd 0.00308f
C2051 vdd.n46 gnd 0.003261f
C2052 vdd.n47 gnd 0.00728f
C2053 vdd.n48 gnd 0.00728f
C2054 vdd.n49 gnd 0.003261f
C2055 vdd.n50 gnd 0.00308f
C2056 vdd.n51 gnd 0.005732f
C2057 vdd.n52 gnd 0.005732f
C2058 vdd.n53 gnd 0.00308f
C2059 vdd.n54 gnd 0.003261f
C2060 vdd.n55 gnd 0.00728f
C2061 vdd.n56 gnd 0.00728f
C2062 vdd.n57 gnd 0.003261f
C2063 vdd.n58 gnd 0.00308f
C2064 vdd.n59 gnd 0.005732f
C2065 vdd.n60 gnd 0.005732f
C2066 vdd.n61 gnd 0.00308f
C2067 vdd.n62 gnd 0.003261f
C2068 vdd.n63 gnd 0.00728f
C2069 vdd.n64 gnd 0.00728f
C2070 vdd.n65 gnd 0.017212f
C2071 vdd.n66 gnd 0.003171f
C2072 vdd.n67 gnd 0.00308f
C2073 vdd.n68 gnd 0.014815f
C2074 vdd.n69 gnd 0.010343f
C2075 vdd.t278 gnd 0.036237f
C2076 vdd.t218 gnd 0.036237f
C2077 vdd.n70 gnd 0.249044f
C2078 vdd.n71 gnd 0.195835f
C2079 vdd.t291 gnd 0.036237f
C2080 vdd.t186 gnd 0.036237f
C2081 vdd.n72 gnd 0.249044f
C2082 vdd.n73 gnd 0.158038f
C2083 vdd.t266 gnd 0.036237f
C2084 vdd.t208 gnd 0.036237f
C2085 vdd.n74 gnd 0.249044f
C2086 vdd.n75 gnd 0.158038f
C2087 vdd.t286 gnd 0.036237f
C2088 vdd.t260 gnd 0.036237f
C2089 vdd.n76 gnd 0.249044f
C2090 vdd.n77 gnd 0.158038f
C2091 vdd.t153 gnd 0.036237f
C2092 vdd.t197 gnd 0.036237f
C2093 vdd.n78 gnd 0.249044f
C2094 vdd.n79 gnd 0.158038f
C2095 vdd.t164 gnd 0.036237f
C2096 vdd.t221 gnd 0.036237f
C2097 vdd.n80 gnd 0.249044f
C2098 vdd.n81 gnd 0.158038f
C2099 vdd.t192 gnd 0.036237f
C2100 vdd.t274 gnd 0.036237f
C2101 vdd.n82 gnd 0.249044f
C2102 vdd.n83 gnd 0.158038f
C2103 vdd.t169 gnd 0.036237f
C2104 vdd.t246 gnd 0.036237f
C2105 vdd.n84 gnd 0.249044f
C2106 vdd.n85 gnd 0.158038f
C2107 vdd.t176 gnd 0.036237f
C2108 vdd.t261 gnd 0.036237f
C2109 vdd.n86 gnd 0.249044f
C2110 vdd.n87 gnd 0.158038f
C2111 vdd.n88 gnd 0.006177f
C2112 vdd.n89 gnd 0.005732f
C2113 vdd.n90 gnd 0.003171f
C2114 vdd.n91 gnd 0.00728f
C2115 vdd.n92 gnd 0.00308f
C2116 vdd.n93 gnd 0.003261f
C2117 vdd.n94 gnd 0.005732f
C2118 vdd.n95 gnd 0.00308f
C2119 vdd.n96 gnd 0.00728f
C2120 vdd.n97 gnd 0.003261f
C2121 vdd.n98 gnd 0.005732f
C2122 vdd.n99 gnd 0.00308f
C2123 vdd.n100 gnd 0.00546f
C2124 vdd.n101 gnd 0.005477f
C2125 vdd.t203 gnd 0.015641f
C2126 vdd.n102 gnd 0.034801f
C2127 vdd.n103 gnd 0.181113f
C2128 vdd.n104 gnd 0.00308f
C2129 vdd.n105 gnd 0.003261f
C2130 vdd.n106 gnd 0.00728f
C2131 vdd.n107 gnd 0.00728f
C2132 vdd.n108 gnd 0.003261f
C2133 vdd.n109 gnd 0.00308f
C2134 vdd.n110 gnd 0.005732f
C2135 vdd.n111 gnd 0.005732f
C2136 vdd.n112 gnd 0.00308f
C2137 vdd.n113 gnd 0.003261f
C2138 vdd.n114 gnd 0.00728f
C2139 vdd.n115 gnd 0.00728f
C2140 vdd.n116 gnd 0.003261f
C2141 vdd.n117 gnd 0.00308f
C2142 vdd.n118 gnd 0.005732f
C2143 vdd.n119 gnd 0.005732f
C2144 vdd.n120 gnd 0.00308f
C2145 vdd.n121 gnd 0.003261f
C2146 vdd.n122 gnd 0.00728f
C2147 vdd.n123 gnd 0.00728f
C2148 vdd.n124 gnd 0.017212f
C2149 vdd.n125 gnd 0.003171f
C2150 vdd.n126 gnd 0.00308f
C2151 vdd.n127 gnd 0.014815f
C2152 vdd.n128 gnd 0.010019f
C2153 vdd.n129 gnd 0.117581f
C2154 vdd.n130 gnd 0.006177f
C2155 vdd.n131 gnd 0.005732f
C2156 vdd.n132 gnd 0.003171f
C2157 vdd.n133 gnd 0.00728f
C2158 vdd.n134 gnd 0.00308f
C2159 vdd.n135 gnd 0.003261f
C2160 vdd.n136 gnd 0.005732f
C2161 vdd.n137 gnd 0.00308f
C2162 vdd.n138 gnd 0.00728f
C2163 vdd.n139 gnd 0.003261f
C2164 vdd.n140 gnd 0.005732f
C2165 vdd.n141 gnd 0.00308f
C2166 vdd.n142 gnd 0.00546f
C2167 vdd.n143 gnd 0.005477f
C2168 vdd.t224 gnd 0.015641f
C2169 vdd.n144 gnd 0.034801f
C2170 vdd.n145 gnd 0.181113f
C2171 vdd.n146 gnd 0.00308f
C2172 vdd.n147 gnd 0.003261f
C2173 vdd.n148 gnd 0.00728f
C2174 vdd.n149 gnd 0.00728f
C2175 vdd.n150 gnd 0.003261f
C2176 vdd.n151 gnd 0.00308f
C2177 vdd.n152 gnd 0.005732f
C2178 vdd.n153 gnd 0.005732f
C2179 vdd.n154 gnd 0.00308f
C2180 vdd.n155 gnd 0.003261f
C2181 vdd.n156 gnd 0.00728f
C2182 vdd.n157 gnd 0.00728f
C2183 vdd.n158 gnd 0.003261f
C2184 vdd.n159 gnd 0.00308f
C2185 vdd.n160 gnd 0.005732f
C2186 vdd.n161 gnd 0.005732f
C2187 vdd.n162 gnd 0.00308f
C2188 vdd.n163 gnd 0.003261f
C2189 vdd.n164 gnd 0.00728f
C2190 vdd.n165 gnd 0.00728f
C2191 vdd.n166 gnd 0.017212f
C2192 vdd.n167 gnd 0.003171f
C2193 vdd.n168 gnd 0.00308f
C2194 vdd.n169 gnd 0.014815f
C2195 vdd.n170 gnd 0.010343f
C2196 vdd.t226 gnd 0.036237f
C2197 vdd.t256 gnd 0.036237f
C2198 vdd.n171 gnd 0.249044f
C2199 vdd.n172 gnd 0.195835f
C2200 vdd.t151 gnd 0.036237f
C2201 vdd.t216 gnd 0.036237f
C2202 vdd.n173 gnd 0.249044f
C2203 vdd.n174 gnd 0.158038f
C2204 vdd.t254 gnd 0.036237f
C2205 vdd.t135 gnd 0.036237f
C2206 vdd.n175 gnd 0.249044f
C2207 vdd.n176 gnd 0.158038f
C2208 vdd.t194 gnd 0.036237f
C2209 vdd.t196 gnd 0.036237f
C2210 vdd.n177 gnd 0.249044f
C2211 vdd.n178 gnd 0.158038f
C2212 vdd.t280 gnd 0.036237f
C2213 vdd.t137 gnd 0.036237f
C2214 vdd.n179 gnd 0.249044f
C2215 vdd.n180 gnd 0.158038f
C2216 vdd.t190 gnd 0.036237f
C2217 vdd.t276 gnd 0.036237f
C2218 vdd.n181 gnd 0.249044f
C2219 vdd.n182 gnd 0.158038f
C2220 vdd.t277 gnd 0.036237f
C2221 vdd.t162 gnd 0.036237f
C2222 vdd.n183 gnd 0.249044f
C2223 vdd.n184 gnd 0.158038f
C2224 vdd.t255 gnd 0.036237f
C2225 vdd.t273 gnd 0.036237f
C2226 vdd.n185 gnd 0.249044f
C2227 vdd.n186 gnd 0.158038f
C2228 vdd.t160 gnd 0.036237f
C2229 vdd.t215 gnd 0.036237f
C2230 vdd.n187 gnd 0.249044f
C2231 vdd.n188 gnd 0.158038f
C2232 vdd.n189 gnd 0.006177f
C2233 vdd.n190 gnd 0.005732f
C2234 vdd.n191 gnd 0.003171f
C2235 vdd.n192 gnd 0.00728f
C2236 vdd.n193 gnd 0.00308f
C2237 vdd.n194 gnd 0.003261f
C2238 vdd.n195 gnd 0.005732f
C2239 vdd.n196 gnd 0.00308f
C2240 vdd.n197 gnd 0.00728f
C2241 vdd.n198 gnd 0.003261f
C2242 vdd.n199 gnd 0.005732f
C2243 vdd.n200 gnd 0.00308f
C2244 vdd.n201 gnd 0.00546f
C2245 vdd.n202 gnd 0.005477f
C2246 vdd.t252 gnd 0.015641f
C2247 vdd.n203 gnd 0.034801f
C2248 vdd.n204 gnd 0.181113f
C2249 vdd.n205 gnd 0.00308f
C2250 vdd.n206 gnd 0.003261f
C2251 vdd.n207 gnd 0.00728f
C2252 vdd.n208 gnd 0.00728f
C2253 vdd.n209 gnd 0.003261f
C2254 vdd.n210 gnd 0.00308f
C2255 vdd.n211 gnd 0.005732f
C2256 vdd.n212 gnd 0.005732f
C2257 vdd.n213 gnd 0.00308f
C2258 vdd.n214 gnd 0.003261f
C2259 vdd.n215 gnd 0.00728f
C2260 vdd.n216 gnd 0.00728f
C2261 vdd.n217 gnd 0.003261f
C2262 vdd.n218 gnd 0.00308f
C2263 vdd.n219 gnd 0.005732f
C2264 vdd.n220 gnd 0.005732f
C2265 vdd.n221 gnd 0.00308f
C2266 vdd.n222 gnd 0.003261f
C2267 vdd.n223 gnd 0.00728f
C2268 vdd.n224 gnd 0.00728f
C2269 vdd.n225 gnd 0.017212f
C2270 vdd.n226 gnd 0.003171f
C2271 vdd.n227 gnd 0.00308f
C2272 vdd.n228 gnd 0.014815f
C2273 vdd.n229 gnd 0.010019f
C2274 vdd.n230 gnd 0.069949f
C2275 vdd.n231 gnd 0.252044f
C2276 vdd.n232 gnd 0.006177f
C2277 vdd.n233 gnd 0.005732f
C2278 vdd.n234 gnd 0.003171f
C2279 vdd.n235 gnd 0.00728f
C2280 vdd.n236 gnd 0.00308f
C2281 vdd.n237 gnd 0.003261f
C2282 vdd.n238 gnd 0.005732f
C2283 vdd.n239 gnd 0.00308f
C2284 vdd.n240 gnd 0.00728f
C2285 vdd.n241 gnd 0.003261f
C2286 vdd.n242 gnd 0.005732f
C2287 vdd.n243 gnd 0.00308f
C2288 vdd.n244 gnd 0.00546f
C2289 vdd.n245 gnd 0.005477f
C2290 vdd.t240 gnd 0.015641f
C2291 vdd.n246 gnd 0.034801f
C2292 vdd.n247 gnd 0.181113f
C2293 vdd.n248 gnd 0.00308f
C2294 vdd.n249 gnd 0.003261f
C2295 vdd.n250 gnd 0.00728f
C2296 vdd.n251 gnd 0.00728f
C2297 vdd.n252 gnd 0.003261f
C2298 vdd.n253 gnd 0.00308f
C2299 vdd.n254 gnd 0.005732f
C2300 vdd.n255 gnd 0.005732f
C2301 vdd.n256 gnd 0.00308f
C2302 vdd.n257 gnd 0.003261f
C2303 vdd.n258 gnd 0.00728f
C2304 vdd.n259 gnd 0.00728f
C2305 vdd.n260 gnd 0.003261f
C2306 vdd.n261 gnd 0.00308f
C2307 vdd.n262 gnd 0.005732f
C2308 vdd.n263 gnd 0.005732f
C2309 vdd.n264 gnd 0.00308f
C2310 vdd.n265 gnd 0.003261f
C2311 vdd.n266 gnd 0.00728f
C2312 vdd.n267 gnd 0.00728f
C2313 vdd.n268 gnd 0.017212f
C2314 vdd.n269 gnd 0.003171f
C2315 vdd.n270 gnd 0.00308f
C2316 vdd.n271 gnd 0.014815f
C2317 vdd.n272 gnd 0.010343f
C2318 vdd.t241 gnd 0.036237f
C2319 vdd.t270 gnd 0.036237f
C2320 vdd.n273 gnd 0.249044f
C2321 vdd.n274 gnd 0.195835f
C2322 vdd.t173 gnd 0.036237f
C2323 vdd.t237 gnd 0.036237f
C2324 vdd.n275 gnd 0.249044f
C2325 vdd.n276 gnd 0.158038f
C2326 vdd.t264 gnd 0.036237f
C2327 vdd.t167 gnd 0.036237f
C2328 vdd.n277 gnd 0.249044f
C2329 vdd.n278 gnd 0.158038f
C2330 vdd.t211 gnd 0.036237f
C2331 vdd.t213 gnd 0.036237f
C2332 vdd.n279 gnd 0.249044f
C2333 vdd.n280 gnd 0.158038f
C2334 vdd.t290 gnd 0.036237f
C2335 vdd.t206 gnd 0.036237f
C2336 vdd.n281 gnd 0.249044f
C2337 vdd.n282 gnd 0.158038f
C2338 vdd.t207 gnd 0.036237f
C2339 vdd.t288 gnd 0.036237f
C2340 vdd.n283 gnd 0.249044f
C2341 vdd.n284 gnd 0.158038f
C2342 vdd.t289 gnd 0.036237f
C2343 vdd.t184 gnd 0.036237f
C2344 vdd.n285 gnd 0.249044f
C2345 vdd.n286 gnd 0.158038f
C2346 vdd.t268 gnd 0.036237f
C2347 vdd.t285 gnd 0.036237f
C2348 vdd.n287 gnd 0.249044f
C2349 vdd.n288 gnd 0.158038f
C2350 vdd.t177 gnd 0.036237f
C2351 vdd.t238 gnd 0.036237f
C2352 vdd.n289 gnd 0.249044f
C2353 vdd.n290 gnd 0.158038f
C2354 vdd.n291 gnd 0.006177f
C2355 vdd.n292 gnd 0.005732f
C2356 vdd.n293 gnd 0.003171f
C2357 vdd.n294 gnd 0.00728f
C2358 vdd.n295 gnd 0.00308f
C2359 vdd.n296 gnd 0.003261f
C2360 vdd.n297 gnd 0.005732f
C2361 vdd.n298 gnd 0.00308f
C2362 vdd.n299 gnd 0.00728f
C2363 vdd.n300 gnd 0.003261f
C2364 vdd.n301 gnd 0.005732f
C2365 vdd.n302 gnd 0.00308f
C2366 vdd.n303 gnd 0.00546f
C2367 vdd.n304 gnd 0.005477f
C2368 vdd.t263 gnd 0.015641f
C2369 vdd.n305 gnd 0.034801f
C2370 vdd.n306 gnd 0.181113f
C2371 vdd.n307 gnd 0.00308f
C2372 vdd.n308 gnd 0.003261f
C2373 vdd.n309 gnd 0.00728f
C2374 vdd.n310 gnd 0.00728f
C2375 vdd.n311 gnd 0.003261f
C2376 vdd.n312 gnd 0.00308f
C2377 vdd.n313 gnd 0.005732f
C2378 vdd.n314 gnd 0.005732f
C2379 vdd.n315 gnd 0.00308f
C2380 vdd.n316 gnd 0.003261f
C2381 vdd.n317 gnd 0.00728f
C2382 vdd.n318 gnd 0.00728f
C2383 vdd.n319 gnd 0.003261f
C2384 vdd.n320 gnd 0.00308f
C2385 vdd.n321 gnd 0.005732f
C2386 vdd.n322 gnd 0.005732f
C2387 vdd.n323 gnd 0.00308f
C2388 vdd.n324 gnd 0.003261f
C2389 vdd.n325 gnd 0.00728f
C2390 vdd.n326 gnd 0.00728f
C2391 vdd.n327 gnd 0.017212f
C2392 vdd.n328 gnd 0.003171f
C2393 vdd.n329 gnd 0.00308f
C2394 vdd.n330 gnd 0.014815f
C2395 vdd.n331 gnd 0.010019f
C2396 vdd.n332 gnd 0.069949f
C2397 vdd.n333 gnd 0.288535f
C2398 vdd.n334 gnd 0.00865f
C2399 vdd.n335 gnd 0.011255f
C2400 vdd.n336 gnd 0.009059f
C2401 vdd.n337 gnd 0.009059f
C2402 vdd.n338 gnd 0.011255f
C2403 vdd.n339 gnd 0.011255f
C2404 vdd.n340 gnd 0.822423f
C2405 vdd.n341 gnd 0.011255f
C2406 vdd.n342 gnd 0.011255f
C2407 vdd.n343 gnd 0.011255f
C2408 vdd.n344 gnd 0.891437f
C2409 vdd.n345 gnd 0.011255f
C2410 vdd.n346 gnd 0.011255f
C2411 vdd.n347 gnd 0.011255f
C2412 vdd.n348 gnd 0.011255f
C2413 vdd.n349 gnd 0.009059f
C2414 vdd.n350 gnd 0.011255f
C2415 vdd.t220 gnd 0.575121f
C2416 vdd.n351 gnd 0.011255f
C2417 vdd.n352 gnd 0.011255f
C2418 vdd.n353 gnd 0.011255f
C2419 vdd.t161 gnd 0.575121f
C2420 vdd.n354 gnd 0.011255f
C2421 vdd.n355 gnd 0.011255f
C2422 vdd.n356 gnd 0.011255f
C2423 vdd.n357 gnd 0.011255f
C2424 vdd.n358 gnd 0.011255f
C2425 vdd.n359 gnd 0.009059f
C2426 vdd.n360 gnd 0.011255f
C2427 vdd.n361 gnd 0.649887f
C2428 vdd.n362 gnd 0.011255f
C2429 vdd.n363 gnd 0.011255f
C2430 vdd.n364 gnd 0.011255f
C2431 vdd.t245 gnd 0.575121f
C2432 vdd.n365 gnd 0.011255f
C2433 vdd.n366 gnd 0.011255f
C2434 vdd.n367 gnd 0.011255f
C2435 vdd.n368 gnd 0.011255f
C2436 vdd.n369 gnd 0.011255f
C2437 vdd.n370 gnd 0.009059f
C2438 vdd.n371 gnd 0.011255f
C2439 vdd.t159 gnd 0.575121f
C2440 vdd.n372 gnd 0.011255f
C2441 vdd.n373 gnd 0.011255f
C2442 vdd.n374 gnd 0.011255f
C2443 vdd.n375 gnd 0.672891f
C2444 vdd.n376 gnd 0.011255f
C2445 vdd.n377 gnd 0.011255f
C2446 vdd.n378 gnd 0.011255f
C2447 vdd.n379 gnd 0.011255f
C2448 vdd.n380 gnd 0.011255f
C2449 vdd.n381 gnd 0.009059f
C2450 vdd.n382 gnd 0.011255f
C2451 vdd.t202 gnd 0.575121f
C2452 vdd.n383 gnd 0.011255f
C2453 vdd.n384 gnd 0.011255f
C2454 vdd.n385 gnd 0.011255f
C2455 vdd.n386 gnd 0.580872f
C2456 vdd.n387 gnd 0.011255f
C2457 vdd.n388 gnd 0.011255f
C2458 vdd.n389 gnd 0.011255f
C2459 vdd.n390 gnd 0.011255f
C2460 vdd.n391 gnd 0.027228f
C2461 vdd.n392 gnd 0.027811f
C2462 vdd.t81 gnd 0.575121f
C2463 vdd.n393 gnd 0.027228f
C2464 vdd.n425 gnd 0.011255f
C2465 vdd.t83 gnd 0.13847f
C2466 vdd.t82 gnd 0.147986f
C2467 vdd.t80 gnd 0.18084f
C2468 vdd.n426 gnd 0.231812f
C2469 vdd.n427 gnd 0.19567f
C2470 vdd.n428 gnd 0.014857f
C2471 vdd.n429 gnd 0.011255f
C2472 vdd.n430 gnd 0.009059f
C2473 vdd.n431 gnd 0.011255f
C2474 vdd.n432 gnd 0.009059f
C2475 vdd.n433 gnd 0.011255f
C2476 vdd.n434 gnd 0.009059f
C2477 vdd.n435 gnd 0.011255f
C2478 vdd.n436 gnd 0.009059f
C2479 vdd.n437 gnd 0.011255f
C2480 vdd.n438 gnd 0.009059f
C2481 vdd.n439 gnd 0.011255f
C2482 vdd.t123 gnd 0.13847f
C2483 vdd.t122 gnd 0.147986f
C2484 vdd.t121 gnd 0.18084f
C2485 vdd.n440 gnd 0.231812f
C2486 vdd.n441 gnd 0.19567f
C2487 vdd.n442 gnd 0.009059f
C2488 vdd.n443 gnd 0.011255f
C2489 vdd.n444 gnd 0.009059f
C2490 vdd.n445 gnd 0.011255f
C2491 vdd.n446 gnd 0.009059f
C2492 vdd.n447 gnd 0.011255f
C2493 vdd.n448 gnd 0.009059f
C2494 vdd.n449 gnd 0.011255f
C2495 vdd.n450 gnd 0.009059f
C2496 vdd.n451 gnd 0.011255f
C2497 vdd.t129 gnd 0.13847f
C2498 vdd.t128 gnd 0.147986f
C2499 vdd.t127 gnd 0.18084f
C2500 vdd.n452 gnd 0.231812f
C2501 vdd.n453 gnd 0.19567f
C2502 vdd.n454 gnd 0.019387f
C2503 vdd.n455 gnd 0.011255f
C2504 vdd.n456 gnd 0.009059f
C2505 vdd.n457 gnd 0.011255f
C2506 vdd.n458 gnd 0.009059f
C2507 vdd.n459 gnd 0.011255f
C2508 vdd.n460 gnd 0.009059f
C2509 vdd.n461 gnd 0.011255f
C2510 vdd.n462 gnd 0.009059f
C2511 vdd.n463 gnd 0.011255f
C2512 vdd.n464 gnd 0.027811f
C2513 vdd.n465 gnd 0.007519f
C2514 vdd.n466 gnd 0.009059f
C2515 vdd.n467 gnd 0.011255f
C2516 vdd.n468 gnd 0.011255f
C2517 vdd.n469 gnd 0.009059f
C2518 vdd.n470 gnd 0.011255f
C2519 vdd.n471 gnd 0.011255f
C2520 vdd.n472 gnd 0.011255f
C2521 vdd.n473 gnd 0.011255f
C2522 vdd.n474 gnd 0.011255f
C2523 vdd.n475 gnd 0.009059f
C2524 vdd.n476 gnd 0.009059f
C2525 vdd.n477 gnd 0.011255f
C2526 vdd.n478 gnd 0.011255f
C2527 vdd.n479 gnd 0.009059f
C2528 vdd.n480 gnd 0.011255f
C2529 vdd.n481 gnd 0.011255f
C2530 vdd.n482 gnd 0.011255f
C2531 vdd.n483 gnd 0.011255f
C2532 vdd.n484 gnd 0.011255f
C2533 vdd.n485 gnd 0.009059f
C2534 vdd.n486 gnd 0.009059f
C2535 vdd.n487 gnd 0.011255f
C2536 vdd.n488 gnd 0.011255f
C2537 vdd.n489 gnd 0.009059f
C2538 vdd.n490 gnd 0.011255f
C2539 vdd.n491 gnd 0.011255f
C2540 vdd.n492 gnd 0.011255f
C2541 vdd.n493 gnd 0.011255f
C2542 vdd.n494 gnd 0.011255f
C2543 vdd.n495 gnd 0.009059f
C2544 vdd.n496 gnd 0.009059f
C2545 vdd.n497 gnd 0.011255f
C2546 vdd.n498 gnd 0.011255f
C2547 vdd.n499 gnd 0.009059f
C2548 vdd.n500 gnd 0.011255f
C2549 vdd.n501 gnd 0.011255f
C2550 vdd.n502 gnd 0.011255f
C2551 vdd.n503 gnd 0.011255f
C2552 vdd.n504 gnd 0.011255f
C2553 vdd.n505 gnd 0.009059f
C2554 vdd.n506 gnd 0.009059f
C2555 vdd.n507 gnd 0.011255f
C2556 vdd.n508 gnd 0.011255f
C2557 vdd.n509 gnd 0.007564f
C2558 vdd.n510 gnd 0.011255f
C2559 vdd.n511 gnd 0.011255f
C2560 vdd.n512 gnd 0.011255f
C2561 vdd.n513 gnd 0.011255f
C2562 vdd.n514 gnd 0.011255f
C2563 vdd.n515 gnd 0.007564f
C2564 vdd.n516 gnd 0.009059f
C2565 vdd.n517 gnd 0.011255f
C2566 vdd.n518 gnd 0.011255f
C2567 vdd.n519 gnd 0.009059f
C2568 vdd.n520 gnd 0.011255f
C2569 vdd.n521 gnd 0.011255f
C2570 vdd.n522 gnd 0.011255f
C2571 vdd.n523 gnd 0.011255f
C2572 vdd.n524 gnd 0.011255f
C2573 vdd.n525 gnd 0.009059f
C2574 vdd.n526 gnd 0.009059f
C2575 vdd.n527 gnd 0.011255f
C2576 vdd.n528 gnd 0.011255f
C2577 vdd.n529 gnd 0.009059f
C2578 vdd.n530 gnd 0.011255f
C2579 vdd.n531 gnd 0.011255f
C2580 vdd.n532 gnd 0.011255f
C2581 vdd.n533 gnd 0.011255f
C2582 vdd.n534 gnd 0.011255f
C2583 vdd.n535 gnd 0.009059f
C2584 vdd.n536 gnd 0.009059f
C2585 vdd.n537 gnd 0.011255f
C2586 vdd.n538 gnd 0.011255f
C2587 vdd.n539 gnd 0.009059f
C2588 vdd.n540 gnd 0.011255f
C2589 vdd.n541 gnd 0.011255f
C2590 vdd.n542 gnd 0.011255f
C2591 vdd.n543 gnd 0.011255f
C2592 vdd.n544 gnd 0.011255f
C2593 vdd.n545 gnd 0.009059f
C2594 vdd.n546 gnd 0.009059f
C2595 vdd.n547 gnd 0.011255f
C2596 vdd.n548 gnd 0.011255f
C2597 vdd.n549 gnd 0.009059f
C2598 vdd.n550 gnd 0.011255f
C2599 vdd.n551 gnd 0.011255f
C2600 vdd.n552 gnd 0.011255f
C2601 vdd.n553 gnd 0.011255f
C2602 vdd.n554 gnd 0.011255f
C2603 vdd.n555 gnd 0.009059f
C2604 vdd.n556 gnd 0.009059f
C2605 vdd.n557 gnd 0.011255f
C2606 vdd.n558 gnd 0.011255f
C2607 vdd.n559 gnd 0.009059f
C2608 vdd.n560 gnd 0.011255f
C2609 vdd.n561 gnd 0.011255f
C2610 vdd.n562 gnd 0.011255f
C2611 vdd.n563 gnd 0.011255f
C2612 vdd.n564 gnd 0.011255f
C2613 vdd.n565 gnd 0.00616f
C2614 vdd.n566 gnd 0.019387f
C2615 vdd.n567 gnd 0.011255f
C2616 vdd.n568 gnd 0.011255f
C2617 vdd.n569 gnd 0.008969f
C2618 vdd.n570 gnd 0.011255f
C2619 vdd.n571 gnd 0.011255f
C2620 vdd.n572 gnd 0.011255f
C2621 vdd.n573 gnd 0.011255f
C2622 vdd.n574 gnd 0.011255f
C2623 vdd.n575 gnd 0.009059f
C2624 vdd.n576 gnd 0.009059f
C2625 vdd.n577 gnd 0.011255f
C2626 vdd.n578 gnd 0.011255f
C2627 vdd.n579 gnd 0.009059f
C2628 vdd.n580 gnd 0.011255f
C2629 vdd.n581 gnd 0.011255f
C2630 vdd.n582 gnd 0.011255f
C2631 vdd.n583 gnd 0.011255f
C2632 vdd.n584 gnd 0.011255f
C2633 vdd.n585 gnd 0.009059f
C2634 vdd.n586 gnd 0.009059f
C2635 vdd.n587 gnd 0.011255f
C2636 vdd.n588 gnd 0.011255f
C2637 vdd.n589 gnd 0.009059f
C2638 vdd.n590 gnd 0.011255f
C2639 vdd.n591 gnd 0.011255f
C2640 vdd.n592 gnd 0.011255f
C2641 vdd.n593 gnd 0.011255f
C2642 vdd.n594 gnd 0.011255f
C2643 vdd.n595 gnd 0.009059f
C2644 vdd.n596 gnd 0.009059f
C2645 vdd.n597 gnd 0.011255f
C2646 vdd.n598 gnd 0.011255f
C2647 vdd.n599 gnd 0.009059f
C2648 vdd.n600 gnd 0.011255f
C2649 vdd.n601 gnd 0.011255f
C2650 vdd.n602 gnd 0.011255f
C2651 vdd.n603 gnd 0.011255f
C2652 vdd.n604 gnd 0.011255f
C2653 vdd.n605 gnd 0.009059f
C2654 vdd.n606 gnd 0.009059f
C2655 vdd.n607 gnd 0.011255f
C2656 vdd.n608 gnd 0.011255f
C2657 vdd.n609 gnd 0.009059f
C2658 vdd.n610 gnd 0.011255f
C2659 vdd.n611 gnd 0.011255f
C2660 vdd.n612 gnd 0.011255f
C2661 vdd.n613 gnd 0.011255f
C2662 vdd.n614 gnd 0.011255f
C2663 vdd.n615 gnd 0.009059f
C2664 vdd.n616 gnd 0.011255f
C2665 vdd.n617 gnd 0.009059f
C2666 vdd.n618 gnd 0.004756f
C2667 vdd.n619 gnd 0.011255f
C2668 vdd.n620 gnd 0.011255f
C2669 vdd.n621 gnd 0.009059f
C2670 vdd.n622 gnd 0.011255f
C2671 vdd.n623 gnd 0.009059f
C2672 vdd.n624 gnd 0.011255f
C2673 vdd.n625 gnd 0.009059f
C2674 vdd.n626 gnd 0.011255f
C2675 vdd.n627 gnd 0.009059f
C2676 vdd.n628 gnd 0.011255f
C2677 vdd.n629 gnd 0.009059f
C2678 vdd.n630 gnd 0.011255f
C2679 vdd.n631 gnd 0.009059f
C2680 vdd.n632 gnd 0.011255f
C2681 vdd.n633 gnd 0.626882f
C2682 vdd.t152 gnd 0.575121f
C2683 vdd.n634 gnd 0.011255f
C2684 vdd.n635 gnd 0.009059f
C2685 vdd.n636 gnd 0.011255f
C2686 vdd.n637 gnd 0.009059f
C2687 vdd.n638 gnd 0.011255f
C2688 vdd.t193 gnd 0.575121f
C2689 vdd.n639 gnd 0.011255f
C2690 vdd.n640 gnd 0.009059f
C2691 vdd.n641 gnd 0.011255f
C2692 vdd.n642 gnd 0.009059f
C2693 vdd.n643 gnd 0.011255f
C2694 vdd.t134 gnd 0.575121f
C2695 vdd.n644 gnd 0.718901f
C2696 vdd.n645 gnd 0.011255f
C2697 vdd.n646 gnd 0.009059f
C2698 vdd.n647 gnd 0.011255f
C2699 vdd.n648 gnd 0.009059f
C2700 vdd.n649 gnd 0.011255f
C2701 vdd.t253 gnd 0.575121f
C2702 vdd.n650 gnd 0.011255f
C2703 vdd.n651 gnd 0.009059f
C2704 vdd.n652 gnd 0.011255f
C2705 vdd.n653 gnd 0.009059f
C2706 vdd.n654 gnd 0.011255f
C2707 vdd.n655 gnd 0.799418f
C2708 vdd.n656 gnd 0.954701f
C2709 vdd.t185 gnd 0.575121f
C2710 vdd.n657 gnd 0.011255f
C2711 vdd.n658 gnd 0.009059f
C2712 vdd.n659 gnd 0.011255f
C2713 vdd.n660 gnd 0.009059f
C2714 vdd.n661 gnd 0.011255f
C2715 vdd.n662 gnd 0.603877f
C2716 vdd.n663 gnd 0.011255f
C2717 vdd.n664 gnd 0.009059f
C2718 vdd.n665 gnd 0.011255f
C2719 vdd.n666 gnd 0.009059f
C2720 vdd.n667 gnd 0.011255f
C2721 vdd.t225 gnd 0.575121f
C2722 vdd.t217 gnd 0.575121f
C2723 vdd.n668 gnd 0.011255f
C2724 vdd.n669 gnd 0.009059f
C2725 vdd.n670 gnd 0.011255f
C2726 vdd.n671 gnd 0.009059f
C2727 vdd.n672 gnd 0.011255f
C2728 vdd.t140 gnd 0.575121f
C2729 vdd.n673 gnd 0.011255f
C2730 vdd.n674 gnd 0.009059f
C2731 vdd.n675 gnd 0.011255f
C2732 vdd.n676 gnd 0.009059f
C2733 vdd.n677 gnd 0.011255f
C2734 vdd.n678 gnd 1.15024f
C2735 vdd.n679 gnd 0.937447f
C2736 vdd.n680 gnd 0.011255f
C2737 vdd.n681 gnd 0.009059f
C2738 vdd.n682 gnd 0.027228f
C2739 vdd.n683 gnd 0.007519f
C2740 vdd.n684 gnd 0.027228f
C2741 vdd.t59 gnd 0.575121f
C2742 vdd.n685 gnd 0.027228f
C2743 vdd.n686 gnd 0.007519f
C2744 vdd.n687 gnd 0.00968f
C2745 vdd.t125 gnd 0.13847f
C2746 vdd.t126 gnd 0.147986f
C2747 vdd.t124 gnd 0.18084f
C2748 vdd.n688 gnd 0.231812f
C2749 vdd.n689 gnd 0.194764f
C2750 vdd.n690 gnd 0.013951f
C2751 vdd.n691 gnd 0.011255f
C2752 vdd.n692 gnd 7.92517f
C2753 vdd.n723 gnd 1.58158f
C2754 vdd.n724 gnd 0.011255f
C2755 vdd.n725 gnd 0.011255f
C2756 vdd.n726 gnd 0.027811f
C2757 vdd.n727 gnd 0.00968f
C2758 vdd.n728 gnd 0.011255f
C2759 vdd.n729 gnd 0.009059f
C2760 vdd.n730 gnd 0.007203f
C2761 vdd.n731 gnd 0.018392f
C2762 vdd.n732 gnd 0.009059f
C2763 vdd.n733 gnd 0.011255f
C2764 vdd.n734 gnd 0.011255f
C2765 vdd.n735 gnd 0.011255f
C2766 vdd.n736 gnd 0.011255f
C2767 vdd.n737 gnd 0.011255f
C2768 vdd.n738 gnd 0.011255f
C2769 vdd.n739 gnd 0.011255f
C2770 vdd.n740 gnd 0.011255f
C2771 vdd.n741 gnd 0.011255f
C2772 vdd.n742 gnd 0.011255f
C2773 vdd.n743 gnd 0.011255f
C2774 vdd.n744 gnd 0.011255f
C2775 vdd.n745 gnd 0.011255f
C2776 vdd.n746 gnd 0.011255f
C2777 vdd.n747 gnd 0.007564f
C2778 vdd.n748 gnd 0.011255f
C2779 vdd.n749 gnd 0.011255f
C2780 vdd.n750 gnd 0.011255f
C2781 vdd.n751 gnd 0.011255f
C2782 vdd.n752 gnd 0.011255f
C2783 vdd.n753 gnd 0.011255f
C2784 vdd.n754 gnd 0.011255f
C2785 vdd.n755 gnd 0.011255f
C2786 vdd.n756 gnd 0.011255f
C2787 vdd.n757 gnd 0.011255f
C2788 vdd.n758 gnd 0.011255f
C2789 vdd.n759 gnd 0.011255f
C2790 vdd.n760 gnd 0.011255f
C2791 vdd.n761 gnd 0.011255f
C2792 vdd.n762 gnd 0.011255f
C2793 vdd.n763 gnd 0.011255f
C2794 vdd.n764 gnd 0.011255f
C2795 vdd.n765 gnd 0.011255f
C2796 vdd.n766 gnd 0.011255f
C2797 vdd.n767 gnd 0.008969f
C2798 vdd.t60 gnd 0.13847f
C2799 vdd.t61 gnd 0.147986f
C2800 vdd.t58 gnd 0.18084f
C2801 vdd.n768 gnd 0.231812f
C2802 vdd.n769 gnd 0.194764f
C2803 vdd.n770 gnd 0.011255f
C2804 vdd.n771 gnd 0.011255f
C2805 vdd.n772 gnd 0.011255f
C2806 vdd.n773 gnd 0.011255f
C2807 vdd.n774 gnd 0.011255f
C2808 vdd.n775 gnd 0.011255f
C2809 vdd.n776 gnd 0.011255f
C2810 vdd.n777 gnd 0.011255f
C2811 vdd.n778 gnd 0.011255f
C2812 vdd.n779 gnd 0.011255f
C2813 vdd.n780 gnd 0.011255f
C2814 vdd.n781 gnd 0.011255f
C2815 vdd.n782 gnd 0.011255f
C2816 vdd.n783 gnd 0.007203f
C2817 vdd.n785 gnd 0.007654f
C2818 vdd.n786 gnd 0.007654f
C2819 vdd.n787 gnd 0.007654f
C2820 vdd.n788 gnd 0.007654f
C2821 vdd.n789 gnd 0.007654f
C2822 vdd.n790 gnd 0.007654f
C2823 vdd.n792 gnd 0.007654f
C2824 vdd.n793 gnd 0.007654f
C2825 vdd.n795 gnd 0.007654f
C2826 vdd.n796 gnd 0.005571f
C2827 vdd.n798 gnd 0.007654f
C2828 vdd.t107 gnd 0.309282f
C2829 vdd.t106 gnd 0.316589f
C2830 vdd.t105 gnd 0.201911f
C2831 vdd.n799 gnd 0.109122f
C2832 vdd.n800 gnd 0.061898f
C2833 vdd.n801 gnd 0.010938f
C2834 vdd.n802 gnd 0.017888f
C2835 vdd.n804 gnd 0.007654f
C2836 vdd.n805 gnd 0.782164f
C2837 vdd.n806 gnd 0.016956f
C2838 vdd.n807 gnd 0.016956f
C2839 vdd.n808 gnd 0.007654f
C2840 vdd.n809 gnd 0.018161f
C2841 vdd.n810 gnd 0.007654f
C2842 vdd.n811 gnd 0.007654f
C2843 vdd.n812 gnd 0.007654f
C2844 vdd.n813 gnd 0.007654f
C2845 vdd.n814 gnd 0.007654f
C2846 vdd.n816 gnd 0.007654f
C2847 vdd.n817 gnd 0.007654f
C2848 vdd.n819 gnd 0.007654f
C2849 vdd.n820 gnd 0.007654f
C2850 vdd.n822 gnd 0.007654f
C2851 vdd.n823 gnd 0.007654f
C2852 vdd.n825 gnd 0.007654f
C2853 vdd.n826 gnd 0.007654f
C2854 vdd.n828 gnd 0.007654f
C2855 vdd.n829 gnd 0.007654f
C2856 vdd.n831 gnd 0.007654f
C2857 vdd.t100 gnd 0.309282f
C2858 vdd.t99 gnd 0.316589f
C2859 vdd.t97 gnd 0.201911f
C2860 vdd.n832 gnd 0.109122f
C2861 vdd.n833 gnd 0.061898f
C2862 vdd.n834 gnd 0.007654f
C2863 vdd.n836 gnd 0.007654f
C2864 vdd.n837 gnd 0.007654f
C2865 vdd.t98 gnd 0.391082f
C2866 vdd.n838 gnd 0.007654f
C2867 vdd.n839 gnd 0.007654f
C2868 vdd.n840 gnd 0.007654f
C2869 vdd.n841 gnd 0.007654f
C2870 vdd.n842 gnd 0.007654f
C2871 vdd.n843 gnd 0.782164f
C2872 vdd.n844 gnd 0.007654f
C2873 vdd.n845 gnd 0.007654f
C2874 vdd.n846 gnd 0.684394f
C2875 vdd.n847 gnd 0.007654f
C2876 vdd.n848 gnd 0.007654f
C2877 vdd.n849 gnd 0.006753f
C2878 vdd.n850 gnd 0.007654f
C2879 vdd.n851 gnd 0.690145f
C2880 vdd.n852 gnd 0.007654f
C2881 vdd.n853 gnd 0.007654f
C2882 vdd.n854 gnd 0.007654f
C2883 vdd.n855 gnd 0.007654f
C2884 vdd.n856 gnd 0.007654f
C2885 vdd.n857 gnd 0.782164f
C2886 vdd.n858 gnd 0.007654f
C2887 vdd.n859 gnd 0.007654f
C2888 vdd.t70 gnd 0.350824f
C2889 vdd.t13 gnd 0.092019f
C2890 vdd.n860 gnd 0.007654f
C2891 vdd.n861 gnd 0.007654f
C2892 vdd.n862 gnd 0.007654f
C2893 vdd.t19 gnd 0.391082f
C2894 vdd.n863 gnd 0.007654f
C2895 vdd.n864 gnd 0.007654f
C2896 vdd.n865 gnd 0.007654f
C2897 vdd.n866 gnd 0.007654f
C2898 vdd.n867 gnd 0.007654f
C2899 vdd.t22 gnd 0.391082f
C2900 vdd.n868 gnd 0.007654f
C2901 vdd.n869 gnd 0.007654f
C2902 vdd.n870 gnd 0.649887f
C2903 vdd.n871 gnd 0.007654f
C2904 vdd.n872 gnd 0.007654f
C2905 vdd.n873 gnd 0.007654f
C2906 vdd.n874 gnd 0.47735f
C2907 vdd.n875 gnd 0.007654f
C2908 vdd.n876 gnd 0.007654f
C2909 vdd.t41 gnd 0.391082f
C2910 vdd.n877 gnd 0.007654f
C2911 vdd.n878 gnd 0.007654f
C2912 vdd.n879 gnd 0.007654f
C2913 vdd.n880 gnd 0.649887f
C2914 vdd.n881 gnd 0.007654f
C2915 vdd.n882 gnd 0.007654f
C2916 vdd.t46 gnd 0.33357f
C2917 vdd.t294 gnd 0.304814f
C2918 vdd.n883 gnd 0.007654f
C2919 vdd.n884 gnd 0.007654f
C2920 vdd.n885 gnd 0.007654f
C2921 vdd.t31 gnd 0.391082f
C2922 vdd.n886 gnd 0.007654f
C2923 vdd.n887 gnd 0.007654f
C2924 vdd.t30 gnd 0.391082f
C2925 vdd.n888 gnd 0.007654f
C2926 vdd.n889 gnd 0.007654f
C2927 vdd.n890 gnd 0.007654f
C2928 vdd.t10 gnd 0.28756f
C2929 vdd.n891 gnd 0.007654f
C2930 vdd.n892 gnd 0.007654f
C2931 vdd.n893 gnd 0.66714f
C2932 vdd.n894 gnd 0.007654f
C2933 vdd.n895 gnd 0.007654f
C2934 vdd.n896 gnd 0.007654f
C2935 vdd.n897 gnd 0.782164f
C2936 vdd.n898 gnd 0.007654f
C2937 vdd.n899 gnd 0.007654f
C2938 vdd.t28 gnd 0.350824f
C2939 vdd.n900 gnd 0.494604f
C2940 vdd.n901 gnd 0.007654f
C2941 vdd.n902 gnd 0.007654f
C2942 vdd.n903 gnd 0.007654f
C2943 vdd.t14 gnd 0.391082f
C2944 vdd.n904 gnd 0.007654f
C2945 vdd.n905 gnd 0.007654f
C2946 vdd.n906 gnd 0.007654f
C2947 vdd.n907 gnd 0.007654f
C2948 vdd.n908 gnd 0.007654f
C2949 vdd.t132 gnd 0.782164f
C2950 vdd.n909 gnd 0.007654f
C2951 vdd.n910 gnd 0.007654f
C2952 vdd.t102 gnd 0.391082f
C2953 vdd.n911 gnd 0.007654f
C2954 vdd.n912 gnd 0.018161f
C2955 vdd.n913 gnd 0.018161f
C2956 vdd.t44 gnd 0.736155f
C2957 vdd.n914 gnd 0.016956f
C2958 vdd.n915 gnd 0.016956f
C2959 vdd.n916 gnd 0.018161f
C2960 vdd.n917 gnd 0.007654f
C2961 vdd.n918 gnd 0.007654f
C2962 vdd.t37 gnd 0.736155f
C2963 vdd.n936 gnd 0.018161f
C2964 vdd.n954 gnd 0.016956f
C2965 vdd.n955 gnd 0.007654f
C2966 vdd.n956 gnd 0.016956f
C2967 vdd.t120 gnd 0.309282f
C2968 vdd.t119 gnd 0.316589f
C2969 vdd.t118 gnd 0.201911f
C2970 vdd.n957 gnd 0.109122f
C2971 vdd.n958 gnd 0.061898f
C2972 vdd.n959 gnd 0.017888f
C2973 vdd.n960 gnd 0.007654f
C2974 vdd.t35 gnd 0.782164f
C2975 vdd.n961 gnd 0.016956f
C2976 vdd.n962 gnd 0.007654f
C2977 vdd.n963 gnd 0.018161f
C2978 vdd.n964 gnd 0.007654f
C2979 vdd.t96 gnd 0.309282f
C2980 vdd.t95 gnd 0.316589f
C2981 vdd.t93 gnd 0.201911f
C2982 vdd.n965 gnd 0.109122f
C2983 vdd.n966 gnd 0.061898f
C2984 vdd.n967 gnd 0.010938f
C2985 vdd.n968 gnd 0.007654f
C2986 vdd.n969 gnd 0.007654f
C2987 vdd.t94 gnd 0.391082f
C2988 vdd.n970 gnd 0.007654f
C2989 vdd.n971 gnd 0.007654f
C2990 vdd.n972 gnd 0.007654f
C2991 vdd.n973 gnd 0.007654f
C2992 vdd.n974 gnd 0.007654f
C2993 vdd.n975 gnd 0.007654f
C2994 vdd.n976 gnd 0.782164f
C2995 vdd.n977 gnd 0.007654f
C2996 vdd.n978 gnd 0.007654f
C2997 vdd.t20 gnd 0.391082f
C2998 vdd.n979 gnd 0.007654f
C2999 vdd.n980 gnd 0.007654f
C3000 vdd.n981 gnd 0.007654f
C3001 vdd.n982 gnd 0.007654f
C3002 vdd.n983 gnd 0.494604f
C3003 vdd.n984 gnd 0.007654f
C3004 vdd.n985 gnd 0.007654f
C3005 vdd.n986 gnd 0.007654f
C3006 vdd.n987 gnd 0.007654f
C3007 vdd.n988 gnd 0.007654f
C3008 vdd.n989 gnd 0.66714f
C3009 vdd.n990 gnd 0.007654f
C3010 vdd.n991 gnd 0.007654f
C3011 vdd.t130 gnd 0.350824f
C3012 vdd.t50 gnd 0.28756f
C3013 vdd.n992 gnd 0.007654f
C3014 vdd.n993 gnd 0.007654f
C3015 vdd.n994 gnd 0.007654f
C3016 vdd.t25 gnd 0.391082f
C3017 vdd.n995 gnd 0.007654f
C3018 vdd.n996 gnd 0.007654f
C3019 vdd.t11 gnd 0.391082f
C3020 vdd.n997 gnd 0.007654f
C3021 vdd.n998 gnd 0.007654f
C3022 vdd.n999 gnd 0.007654f
C3023 vdd.t39 gnd 0.304814f
C3024 vdd.n1000 gnd 0.007654f
C3025 vdd.n1001 gnd 0.007654f
C3026 vdd.n1002 gnd 0.649887f
C3027 vdd.n1003 gnd 0.007654f
C3028 vdd.n1004 gnd 0.007654f
C3029 vdd.n1005 gnd 0.007654f
C3030 vdd.t33 gnd 0.391082f
C3031 vdd.n1006 gnd 0.007654f
C3032 vdd.n1007 gnd 0.007654f
C3033 vdd.t23 gnd 0.33357f
C3034 vdd.n1008 gnd 0.47735f
C3035 vdd.n1009 gnd 0.007654f
C3036 vdd.n1010 gnd 0.007654f
C3037 vdd.n1011 gnd 0.007654f
C3038 vdd.n1012 gnd 0.649887f
C3039 vdd.n1013 gnd 0.007654f
C3040 vdd.n1014 gnd 0.007654f
C3041 vdd.t24 gnd 0.391082f
C3042 vdd.n1015 gnd 0.007654f
C3043 vdd.n1016 gnd 0.007654f
C3044 vdd.n1017 gnd 0.007654f
C3045 vdd.n1018 gnd 0.782164f
C3046 vdd.n1019 gnd 0.007654f
C3047 vdd.n1020 gnd 0.007654f
C3048 vdd.t47 gnd 0.391082f
C3049 vdd.n1021 gnd 0.007654f
C3050 vdd.n1022 gnd 0.007654f
C3051 vdd.n1023 gnd 0.007654f
C3052 vdd.t43 gnd 0.092019f
C3053 vdd.n1024 gnd 0.007654f
C3054 vdd.n1025 gnd 0.007654f
C3055 vdd.n1026 gnd 0.007654f
C3056 vdd.t113 gnd 0.316589f
C3057 vdd.t111 gnd 0.201911f
C3058 vdd.t114 gnd 0.316589f
C3059 vdd.n1027 gnd 0.177936f
C3060 vdd.n1028 gnd 0.007654f
C3061 vdd.n1029 gnd 0.007654f
C3062 vdd.n1030 gnd 0.782164f
C3063 vdd.n1031 gnd 0.007654f
C3064 vdd.n1032 gnd 0.007654f
C3065 vdd.t112 gnd 0.350824f
C3066 vdd.n1033 gnd 0.690145f
C3067 vdd.n1034 gnd 0.007654f
C3068 vdd.n1035 gnd 0.007654f
C3069 vdd.n1036 gnd 0.007654f
C3070 vdd.n1037 gnd 0.684394f
C3071 vdd.n1038 gnd 0.007654f
C3072 vdd.n1039 gnd 0.007654f
C3073 vdd.n1040 gnd 0.007654f
C3074 vdd.n1041 gnd 0.007654f
C3075 vdd.n1042 gnd 0.007654f
C3076 vdd.n1043 gnd 0.782164f
C3077 vdd.n1044 gnd 0.007654f
C3078 vdd.n1045 gnd 0.007654f
C3079 vdd.t55 gnd 0.391082f
C3080 vdd.n1046 gnd 0.007654f
C3081 vdd.n1047 gnd 0.018161f
C3082 vdd.n1048 gnd 0.018161f
C3083 vdd.n1049 gnd 7.92517f
C3084 vdd.n1050 gnd 0.016956f
C3085 vdd.n1051 gnd 0.016956f
C3086 vdd.n1052 gnd 0.018161f
C3087 vdd.n1053 gnd 0.007654f
C3088 vdd.n1054 gnd 0.007654f
C3089 vdd.n1055 gnd 0.007654f
C3090 vdd.n1056 gnd 0.007654f
C3091 vdd.n1057 gnd 0.007654f
C3092 vdd.n1058 gnd 0.007654f
C3093 vdd.n1059 gnd 0.007654f
C3094 vdd.n1060 gnd 0.007654f
C3095 vdd.n1062 gnd 0.007654f
C3096 vdd.n1063 gnd 0.007654f
C3097 vdd.n1064 gnd 0.007203f
C3098 vdd.n1067 gnd 0.027811f
C3099 vdd.n1068 gnd 0.009059f
C3100 vdd.n1069 gnd 0.011255f
C3101 vdd.n1071 gnd 0.011255f
C3102 vdd.n1072 gnd 0.007519f
C3103 vdd.t66 gnd 0.575121f
C3104 vdd.n1073 gnd 8.31625f
C3105 vdd.n1074 gnd 0.011255f
C3106 vdd.n1075 gnd 0.027811f
C3107 vdd.n1076 gnd 0.009059f
C3108 vdd.n1077 gnd 0.011255f
C3109 vdd.n1078 gnd 0.009059f
C3110 vdd.n1079 gnd 0.011255f
C3111 vdd.n1080 gnd 1.15024f
C3112 vdd.n1081 gnd 0.011255f
C3113 vdd.n1082 gnd 0.009059f
C3114 vdd.n1083 gnd 0.009059f
C3115 vdd.n1084 gnd 0.011255f
C3116 vdd.n1085 gnd 0.009059f
C3117 vdd.n1086 gnd 0.011255f
C3118 vdd.t144 gnd 0.575121f
C3119 vdd.n1087 gnd 0.011255f
C3120 vdd.n1088 gnd 0.009059f
C3121 vdd.n1089 gnd 0.011255f
C3122 vdd.n1090 gnd 0.009059f
C3123 vdd.n1091 gnd 0.011255f
C3124 vdd.t271 gnd 0.575121f
C3125 vdd.n1092 gnd 0.011255f
C3126 vdd.n1093 gnd 0.009059f
C3127 vdd.n1094 gnd 0.011255f
C3128 vdd.n1095 gnd 0.009059f
C3129 vdd.n1096 gnd 0.011255f
C3130 vdd.n1097 gnd 0.925945f
C3131 vdd.n1098 gnd 0.954701f
C3132 vdd.t157 gnd 0.575121f
C3133 vdd.n1099 gnd 0.011255f
C3134 vdd.n1100 gnd 0.009059f
C3135 vdd.n1101 gnd 0.011255f
C3136 vdd.n1102 gnd 0.009059f
C3137 vdd.n1103 gnd 0.011255f
C3138 vdd.n1104 gnd 0.730404f
C3139 vdd.n1105 gnd 0.011255f
C3140 vdd.n1106 gnd 0.009059f
C3141 vdd.n1107 gnd 0.011255f
C3142 vdd.n1108 gnd 0.009059f
C3143 vdd.n1109 gnd 0.011255f
C3144 vdd.t146 gnd 0.575121f
C3145 vdd.t187 gnd 0.575121f
C3146 vdd.n1110 gnd 0.011255f
C3147 vdd.n1111 gnd 0.009059f
C3148 vdd.n1112 gnd 0.011255f
C3149 vdd.n1113 gnd 0.009059f
C3150 vdd.n1114 gnd 0.011255f
C3151 vdd.t209 gnd 0.575121f
C3152 vdd.n1115 gnd 0.011255f
C3153 vdd.n1116 gnd 0.009059f
C3154 vdd.n1117 gnd 0.011255f
C3155 vdd.n1118 gnd 0.009059f
C3156 vdd.n1119 gnd 0.011255f
C3157 vdd.t248 gnd 0.575121f
C3158 vdd.n1120 gnd 0.81092f
C3159 vdd.n1121 gnd 0.011255f
C3160 vdd.n1122 gnd 0.009059f
C3161 vdd.n1123 gnd 0.011255f
C3162 vdd.n1124 gnd 0.009059f
C3163 vdd.n1125 gnd 0.011255f
C3164 vdd.n1126 gnd 0.90294f
C3165 vdd.n1127 gnd 0.011255f
C3166 vdd.n1128 gnd 0.009059f
C3167 vdd.n1129 gnd 0.011255f
C3168 vdd.n1130 gnd 0.009059f
C3169 vdd.n1131 gnd 0.011255f
C3170 vdd.n1132 gnd 0.707399f
C3171 vdd.t155 gnd 0.575121f
C3172 vdd.n1133 gnd 0.011255f
C3173 vdd.n1134 gnd 0.009059f
C3174 vdd.n1135 gnd 0.011255f
C3175 vdd.n1136 gnd 0.009059f
C3176 vdd.n1137 gnd 0.011255f
C3177 vdd.t165 gnd 0.575121f
C3178 vdd.n1138 gnd 0.011255f
C3179 vdd.n1139 gnd 0.009059f
C3180 vdd.n1140 gnd 0.011255f
C3181 vdd.n1141 gnd 0.009059f
C3182 vdd.n1142 gnd 0.011255f
C3183 vdd.t182 gnd 0.575121f
C3184 vdd.n1143 gnd 0.638384f
C3185 vdd.n1144 gnd 0.011255f
C3186 vdd.n1145 gnd 0.009059f
C3187 vdd.n1146 gnd 0.011255f
C3188 vdd.n1147 gnd 0.009059f
C3189 vdd.n1148 gnd 0.011255f
C3190 vdd.t227 gnd 0.575121f
C3191 vdd.n1149 gnd 0.011255f
C3192 vdd.n1150 gnd 0.009059f
C3193 vdd.n1151 gnd 0.011255f
C3194 vdd.n1152 gnd 0.009059f
C3195 vdd.n1153 gnd 0.011255f
C3196 vdd.n1154 gnd 0.879935f
C3197 vdd.n1155 gnd 0.954701f
C3198 vdd.t229 gnd 0.575121f
C3199 vdd.n1156 gnd 0.011255f
C3200 vdd.n1157 gnd 0.009059f
C3201 vdd.n1158 gnd 0.011255f
C3202 vdd.n1159 gnd 0.009059f
C3203 vdd.n1160 gnd 0.011255f
C3204 vdd.n1161 gnd 0.684394f
C3205 vdd.n1162 gnd 0.011255f
C3206 vdd.n1163 gnd 0.009059f
C3207 vdd.n1164 gnd 0.011255f
C3208 vdd.n1165 gnd 0.009059f
C3209 vdd.n1166 gnd 0.011255f
C3210 vdd.t180 gnd 0.575121f
C3211 vdd.t178 gnd 0.575121f
C3212 vdd.n1167 gnd 0.011255f
C3213 vdd.n1168 gnd 0.009059f
C3214 vdd.n1169 gnd 0.011255f
C3215 vdd.n1170 gnd 0.009059f
C3216 vdd.n1171 gnd 0.011255f
C3217 vdd.t142 gnd 0.575121f
C3218 vdd.n1172 gnd 0.011255f
C3219 vdd.n1173 gnd 0.009059f
C3220 vdd.n1174 gnd 0.011255f
C3221 vdd.n1175 gnd 0.009059f
C3222 vdd.n1176 gnd 0.011255f
C3223 vdd.t148 gnd 0.575121f
C3224 vdd.n1177 gnd 0.85693f
C3225 vdd.n1178 gnd 0.011255f
C3226 vdd.n1179 gnd 0.009059f
C3227 vdd.n1180 gnd 0.011255f
C3228 vdd.n1181 gnd 0.009059f
C3229 vdd.n1182 gnd 0.011255f
C3230 vdd.n1183 gnd 1.15024f
C3231 vdd.n1184 gnd 0.011255f
C3232 vdd.n1185 gnd 0.009059f
C3233 vdd.n1186 gnd 0.027228f
C3234 vdd.n1187 gnd 0.007519f
C3235 vdd.n1188 gnd 0.027228f
C3236 vdd.t74 gnd 0.575121f
C3237 vdd.n1189 gnd 0.027228f
C3238 vdd.n1190 gnd 0.007519f
C3239 vdd.n1191 gnd 0.011255f
C3240 vdd.n1192 gnd 0.009059f
C3241 vdd.n1193 gnd 0.011255f
C3242 vdd.n1224 gnd 0.027811f
C3243 vdd.n1225 gnd 1.69661f
C3244 vdd.n1226 gnd 0.011255f
C3245 vdd.n1227 gnd 0.009059f
C3246 vdd.n1228 gnd 0.011255f
C3247 vdd.n1229 gnd 0.011255f
C3248 vdd.n1230 gnd 0.011255f
C3249 vdd.n1231 gnd 0.011255f
C3250 vdd.n1232 gnd 0.011255f
C3251 vdd.n1233 gnd 0.009059f
C3252 vdd.n1234 gnd 0.011255f
C3253 vdd.n1235 gnd 0.011255f
C3254 vdd.n1236 gnd 0.011255f
C3255 vdd.n1237 gnd 0.011255f
C3256 vdd.n1238 gnd 0.011255f
C3257 vdd.n1239 gnd 0.009059f
C3258 vdd.n1240 gnd 0.011255f
C3259 vdd.n1241 gnd 0.011255f
C3260 vdd.n1242 gnd 0.011255f
C3261 vdd.n1243 gnd 0.011255f
C3262 vdd.n1244 gnd 0.011255f
C3263 vdd.n1245 gnd 0.009059f
C3264 vdd.n1246 gnd 0.011255f
C3265 vdd.n1247 gnd 0.011255f
C3266 vdd.n1248 gnd 0.011255f
C3267 vdd.n1249 gnd 0.011255f
C3268 vdd.n1250 gnd 0.011255f
C3269 vdd.t88 gnd 0.13847f
C3270 vdd.t89 gnd 0.147986f
C3271 vdd.t87 gnd 0.18084f
C3272 vdd.n1251 gnd 0.231812f
C3273 vdd.n1252 gnd 0.19567f
C3274 vdd.n1253 gnd 0.019387f
C3275 vdd.n1254 gnd 0.011255f
C3276 vdd.n1255 gnd 0.011255f
C3277 vdd.n1256 gnd 0.011255f
C3278 vdd.n1257 gnd 0.011255f
C3279 vdd.n1258 gnd 0.011255f
C3280 vdd.n1259 gnd 0.009059f
C3281 vdd.n1260 gnd 0.011255f
C3282 vdd.n1261 gnd 0.011255f
C3283 vdd.n1262 gnd 0.011255f
C3284 vdd.n1263 gnd 0.011255f
C3285 vdd.n1264 gnd 0.011255f
C3286 vdd.n1265 gnd 0.009059f
C3287 vdd.n1266 gnd 0.011255f
C3288 vdd.n1267 gnd 0.011255f
C3289 vdd.n1268 gnd 0.011255f
C3290 vdd.n1269 gnd 0.011255f
C3291 vdd.n1270 gnd 0.011255f
C3292 vdd.n1271 gnd 0.009059f
C3293 vdd.n1272 gnd 0.011255f
C3294 vdd.n1273 gnd 0.011255f
C3295 vdd.n1274 gnd 0.011255f
C3296 vdd.n1275 gnd 0.011255f
C3297 vdd.n1276 gnd 0.011255f
C3298 vdd.n1277 gnd 0.009059f
C3299 vdd.n1278 gnd 0.011255f
C3300 vdd.n1279 gnd 0.011255f
C3301 vdd.n1280 gnd 0.011255f
C3302 vdd.n1281 gnd 0.011255f
C3303 vdd.n1282 gnd 0.011255f
C3304 vdd.n1283 gnd 0.009059f
C3305 vdd.n1284 gnd 0.011255f
C3306 vdd.n1285 gnd 0.011255f
C3307 vdd.n1286 gnd 0.011255f
C3308 vdd.n1287 gnd 0.011255f
C3309 vdd.n1288 gnd 0.009059f
C3310 vdd.n1289 gnd 0.011255f
C3311 vdd.n1290 gnd 0.011255f
C3312 vdd.n1291 gnd 0.011255f
C3313 vdd.n1292 gnd 0.011255f
C3314 vdd.n1293 gnd 0.011255f
C3315 vdd.n1294 gnd 0.009059f
C3316 vdd.n1295 gnd 0.011255f
C3317 vdd.n1296 gnd 0.011255f
C3318 vdd.n1297 gnd 0.011255f
C3319 vdd.n1298 gnd 0.011255f
C3320 vdd.n1299 gnd 0.011255f
C3321 vdd.n1300 gnd 0.009059f
C3322 vdd.n1301 gnd 0.011255f
C3323 vdd.n1302 gnd 0.011255f
C3324 vdd.n1303 gnd 0.011255f
C3325 vdd.n1304 gnd 0.011255f
C3326 vdd.n1305 gnd 0.011255f
C3327 vdd.n1306 gnd 0.009059f
C3328 vdd.n1307 gnd 0.011255f
C3329 vdd.n1308 gnd 0.011255f
C3330 vdd.n1309 gnd 0.011255f
C3331 vdd.n1310 gnd 0.011255f
C3332 vdd.n1311 gnd 0.011255f
C3333 vdd.n1312 gnd 0.009059f
C3334 vdd.n1313 gnd 0.011255f
C3335 vdd.n1314 gnd 0.011255f
C3336 vdd.n1315 gnd 0.011255f
C3337 vdd.n1316 gnd 0.011255f
C3338 vdd.t85 gnd 0.13847f
C3339 vdd.t86 gnd 0.147986f
C3340 vdd.t84 gnd 0.18084f
C3341 vdd.n1317 gnd 0.231812f
C3342 vdd.n1318 gnd 0.19567f
C3343 vdd.n1319 gnd 0.014857f
C3344 vdd.n1320 gnd 0.004303f
C3345 vdd.n1321 gnd 0.027811f
C3346 vdd.n1322 gnd 0.011255f
C3347 vdd.n1323 gnd 0.004756f
C3348 vdd.n1324 gnd 0.009059f
C3349 vdd.n1325 gnd 0.009059f
C3350 vdd.n1326 gnd 0.011255f
C3351 vdd.n1327 gnd 0.011255f
C3352 vdd.n1328 gnd 0.011255f
C3353 vdd.n1329 gnd 0.009059f
C3354 vdd.n1330 gnd 0.009059f
C3355 vdd.n1331 gnd 0.009059f
C3356 vdd.n1332 gnd 0.011255f
C3357 vdd.n1333 gnd 0.011255f
C3358 vdd.n1334 gnd 0.011255f
C3359 vdd.n1335 gnd 0.009059f
C3360 vdd.n1336 gnd 0.009059f
C3361 vdd.n1337 gnd 0.009059f
C3362 vdd.n1338 gnd 0.011255f
C3363 vdd.n1339 gnd 0.011255f
C3364 vdd.n1340 gnd 0.011255f
C3365 vdd.n1341 gnd 0.009059f
C3366 vdd.n1342 gnd 0.009059f
C3367 vdd.n1343 gnd 0.009059f
C3368 vdd.n1344 gnd 0.011255f
C3369 vdd.n1345 gnd 0.011255f
C3370 vdd.n1346 gnd 0.011255f
C3371 vdd.n1347 gnd 0.009059f
C3372 vdd.n1348 gnd 0.009059f
C3373 vdd.n1349 gnd 0.009059f
C3374 vdd.n1350 gnd 0.011255f
C3375 vdd.n1351 gnd 0.011255f
C3376 vdd.n1352 gnd 0.011255f
C3377 vdd.n1353 gnd 0.008969f
C3378 vdd.n1354 gnd 0.011255f
C3379 vdd.t75 gnd 0.13847f
C3380 vdd.t76 gnd 0.147986f
C3381 vdd.t73 gnd 0.18084f
C3382 vdd.n1355 gnd 0.231812f
C3383 vdd.n1356 gnd 0.19567f
C3384 vdd.n1357 gnd 0.019387f
C3385 vdd.n1358 gnd 0.00616f
C3386 vdd.n1359 gnd 0.011255f
C3387 vdd.n1360 gnd 0.011255f
C3388 vdd.n1361 gnd 0.011255f
C3389 vdd.n1362 gnd 0.009059f
C3390 vdd.n1363 gnd 0.009059f
C3391 vdd.n1364 gnd 0.009059f
C3392 vdd.n1365 gnd 0.011255f
C3393 vdd.n1366 gnd 0.011255f
C3394 vdd.n1367 gnd 0.011255f
C3395 vdd.n1368 gnd 0.009059f
C3396 vdd.n1369 gnd 0.009059f
C3397 vdd.n1370 gnd 0.009059f
C3398 vdd.n1371 gnd 0.011255f
C3399 vdd.n1372 gnd 0.011255f
C3400 vdd.n1373 gnd 0.011255f
C3401 vdd.n1374 gnd 0.009059f
C3402 vdd.n1375 gnd 0.009059f
C3403 vdd.n1376 gnd 0.009059f
C3404 vdd.n1377 gnd 0.011255f
C3405 vdd.n1378 gnd 0.011255f
C3406 vdd.n1379 gnd 0.011255f
C3407 vdd.n1380 gnd 0.009059f
C3408 vdd.n1381 gnd 0.009059f
C3409 vdd.n1382 gnd 0.009059f
C3410 vdd.n1383 gnd 0.011255f
C3411 vdd.n1384 gnd 0.011255f
C3412 vdd.n1385 gnd 0.011255f
C3413 vdd.n1386 gnd 0.009059f
C3414 vdd.n1387 gnd 0.009059f
C3415 vdd.n1388 gnd 0.007564f
C3416 vdd.n1389 gnd 0.011255f
C3417 vdd.n1390 gnd 0.011255f
C3418 vdd.n1391 gnd 0.011255f
C3419 vdd.n1392 gnd 0.007564f
C3420 vdd.n1393 gnd 0.009059f
C3421 vdd.n1394 gnd 0.009059f
C3422 vdd.n1395 gnd 0.011255f
C3423 vdd.n1396 gnd 0.011255f
C3424 vdd.n1397 gnd 0.011255f
C3425 vdd.n1398 gnd 0.009059f
C3426 vdd.n1399 gnd 0.009059f
C3427 vdd.n1400 gnd 0.009059f
C3428 vdd.n1401 gnd 0.011255f
C3429 vdd.n1402 gnd 0.011255f
C3430 vdd.n1403 gnd 0.011255f
C3431 vdd.n1404 gnd 0.009059f
C3432 vdd.n1405 gnd 0.009059f
C3433 vdd.n1406 gnd 0.009059f
C3434 vdd.n1407 gnd 0.011255f
C3435 vdd.n1408 gnd 0.011255f
C3436 vdd.n1409 gnd 0.011255f
C3437 vdd.n1410 gnd 0.009059f
C3438 vdd.n1411 gnd 0.009059f
C3439 vdd.n1412 gnd 0.009059f
C3440 vdd.n1413 gnd 0.011255f
C3441 vdd.n1414 gnd 0.011255f
C3442 vdd.n1415 gnd 0.011255f
C3443 vdd.n1416 gnd 0.009059f
C3444 vdd.n1417 gnd 0.011255f
C3445 vdd.n1418 gnd 2.72607f
C3446 vdd.n1420 gnd 0.027811f
C3447 vdd.n1421 gnd 0.007519f
C3448 vdd.n1422 gnd 0.027811f
C3449 vdd.n1423 gnd 0.027228f
C3450 vdd.n1424 gnd 0.011255f
C3451 vdd.n1425 gnd 0.009059f
C3452 vdd.n1426 gnd 0.011255f
C3453 vdd.n1427 gnd 0.580872f
C3454 vdd.n1428 gnd 0.011255f
C3455 vdd.n1429 gnd 0.009059f
C3456 vdd.n1430 gnd 0.011255f
C3457 vdd.n1431 gnd 0.011255f
C3458 vdd.n1432 gnd 0.011255f
C3459 vdd.n1433 gnd 0.009059f
C3460 vdd.n1434 gnd 0.011255f
C3461 vdd.n1435 gnd 1.05247f
C3462 vdd.n1436 gnd 1.15024f
C3463 vdd.n1437 gnd 0.011255f
C3464 vdd.n1438 gnd 0.009059f
C3465 vdd.n1439 gnd 0.011255f
C3466 vdd.n1440 gnd 0.011255f
C3467 vdd.n1441 gnd 0.011255f
C3468 vdd.n1442 gnd 0.009059f
C3469 vdd.n1443 gnd 0.011255f
C3470 vdd.n1444 gnd 0.672891f
C3471 vdd.n1445 gnd 0.011255f
C3472 vdd.n1446 gnd 0.009059f
C3473 vdd.n1447 gnd 0.011255f
C3474 vdd.n1448 gnd 0.011255f
C3475 vdd.n1449 gnd 0.011255f
C3476 vdd.n1450 gnd 0.009059f
C3477 vdd.n1451 gnd 0.011255f
C3478 vdd.n1452 gnd 0.661389f
C3479 vdd.n1453 gnd 0.868433f
C3480 vdd.n1454 gnd 0.011255f
C3481 vdd.n1455 gnd 0.009059f
C3482 vdd.n1456 gnd 0.011255f
C3483 vdd.n1457 gnd 0.011255f
C3484 vdd.n1458 gnd 0.011255f
C3485 vdd.n1459 gnd 0.009059f
C3486 vdd.n1460 gnd 0.011255f
C3487 vdd.n1461 gnd 0.954701f
C3488 vdd.n1462 gnd 0.011255f
C3489 vdd.n1463 gnd 0.009059f
C3490 vdd.n1464 gnd 0.011255f
C3491 vdd.n1465 gnd 0.011255f
C3492 vdd.n1466 gnd 0.011255f
C3493 vdd.n1467 gnd 0.009059f
C3494 vdd.n1468 gnd 0.011255f
C3495 vdd.t138 gnd 0.575121f
C3496 vdd.n1469 gnd 0.845428f
C3497 vdd.n1470 gnd 0.011255f
C3498 vdd.n1471 gnd 0.009059f
C3499 vdd.n1472 gnd 0.011255f
C3500 vdd.n1473 gnd 0.011255f
C3501 vdd.n1474 gnd 0.011255f
C3502 vdd.n1475 gnd 0.009059f
C3503 vdd.n1476 gnd 0.011255f
C3504 vdd.n1477 gnd 0.649887f
C3505 vdd.n1478 gnd 0.011255f
C3506 vdd.n1479 gnd 0.009059f
C3507 vdd.n1480 gnd 0.011255f
C3508 vdd.n1481 gnd 0.011255f
C3509 vdd.n1482 gnd 0.011255f
C3510 vdd.n1483 gnd 0.009059f
C3511 vdd.n1484 gnd 0.011255f
C3512 vdd.n1485 gnd 0.833925f
C3513 vdd.n1486 gnd 0.695896f
C3514 vdd.n1487 gnd 0.011255f
C3515 vdd.n1488 gnd 0.009059f
C3516 vdd.n1489 gnd 0.011255f
C3517 vdd.n1490 gnd 0.011255f
C3518 vdd.n1491 gnd 0.011255f
C3519 vdd.n1492 gnd 0.009059f
C3520 vdd.n1493 gnd 0.011255f
C3521 vdd.n1494 gnd 0.891437f
C3522 vdd.n1495 gnd 0.011255f
C3523 vdd.n1496 gnd 0.009059f
C3524 vdd.n1497 gnd 0.011255f
C3525 vdd.n1498 gnd 0.011255f
C3526 vdd.n1499 gnd 0.011255f
C3527 vdd.n1500 gnd 0.009059f
C3528 vdd.n1501 gnd 0.011255f
C3529 vdd.t199 gnd 0.575121f
C3530 vdd.n1502 gnd 0.954701f
C3531 vdd.n1503 gnd 0.011255f
C3532 vdd.n1504 gnd 0.009059f
C3533 vdd.n1505 gnd 0.011255f
C3534 vdd.n1506 gnd 0.00865f
C3535 vdd.n1507 gnd 0.006177f
C3536 vdd.n1508 gnd 0.005732f
C3537 vdd.n1509 gnd 0.003171f
C3538 vdd.n1510 gnd 0.00728f
C3539 vdd.n1511 gnd 0.00308f
C3540 vdd.n1512 gnd 0.003261f
C3541 vdd.n1513 gnd 0.005732f
C3542 vdd.n1514 gnd 0.00308f
C3543 vdd.n1515 gnd 0.00728f
C3544 vdd.n1516 gnd 0.003261f
C3545 vdd.n1517 gnd 0.005732f
C3546 vdd.n1518 gnd 0.00308f
C3547 vdd.n1519 gnd 0.00546f
C3548 vdd.n1520 gnd 0.005477f
C3549 vdd.t145 gnd 0.015641f
C3550 vdd.n1521 gnd 0.034801f
C3551 vdd.n1522 gnd 0.181113f
C3552 vdd.n1523 gnd 0.00308f
C3553 vdd.n1524 gnd 0.003261f
C3554 vdd.n1525 gnd 0.00728f
C3555 vdd.n1526 gnd 0.00728f
C3556 vdd.n1527 gnd 0.003261f
C3557 vdd.n1528 gnd 0.00308f
C3558 vdd.n1529 gnd 0.005732f
C3559 vdd.n1530 gnd 0.005732f
C3560 vdd.n1531 gnd 0.00308f
C3561 vdd.n1532 gnd 0.003261f
C3562 vdd.n1533 gnd 0.00728f
C3563 vdd.n1534 gnd 0.00728f
C3564 vdd.n1535 gnd 0.003261f
C3565 vdd.n1536 gnd 0.00308f
C3566 vdd.n1537 gnd 0.005732f
C3567 vdd.n1538 gnd 0.005732f
C3568 vdd.n1539 gnd 0.00308f
C3569 vdd.n1540 gnd 0.003261f
C3570 vdd.n1541 gnd 0.00728f
C3571 vdd.n1542 gnd 0.00728f
C3572 vdd.n1543 gnd 0.017212f
C3573 vdd.n1544 gnd 0.003171f
C3574 vdd.n1545 gnd 0.00308f
C3575 vdd.n1546 gnd 0.014815f
C3576 vdd.n1547 gnd 0.010343f
C3577 vdd.t219 gnd 0.036237f
C3578 vdd.t279 gnd 0.036237f
C3579 vdd.n1548 gnd 0.249044f
C3580 vdd.n1549 gnd 0.195835f
C3581 vdd.t188 gnd 0.036237f
C3582 vdd.t258 gnd 0.036237f
C3583 vdd.n1550 gnd 0.249044f
C3584 vdd.n1551 gnd 0.158038f
C3585 vdd.t210 gnd 0.036237f
C3586 vdd.t267 gnd 0.036237f
C3587 vdd.n1552 gnd 0.249044f
C3588 vdd.n1553 gnd 0.158038f
C3589 vdd.t235 gnd 0.036237f
C3590 vdd.t287 gnd 0.036237f
C3591 vdd.n1554 gnd 0.249044f
C3592 vdd.n1555 gnd 0.158038f
C3593 vdd.t200 gnd 0.036237f
C3594 vdd.t156 gnd 0.036237f
C3595 vdd.n1556 gnd 0.249044f
C3596 vdd.n1557 gnd 0.158038f
C3597 vdd.t222 gnd 0.036237f
C3598 vdd.t166 gnd 0.036237f
C3599 vdd.n1558 gnd 0.249044f
C3600 vdd.n1559 gnd 0.158038f
C3601 vdd.t275 gnd 0.036237f
C3602 vdd.t292 gnd 0.036237f
C3603 vdd.n1560 gnd 0.249044f
C3604 vdd.n1561 gnd 0.158038f
C3605 vdd.t247 gnd 0.036237f
C3606 vdd.t139 gnd 0.036237f
C3607 vdd.n1562 gnd 0.249044f
C3608 vdd.n1563 gnd 0.158038f
C3609 vdd.t236 gnd 0.036237f
C3610 vdd.t181 gnd 0.036237f
C3611 vdd.n1564 gnd 0.249044f
C3612 vdd.n1565 gnd 0.158038f
C3613 vdd.n1566 gnd 0.006177f
C3614 vdd.n1567 gnd 0.005732f
C3615 vdd.n1568 gnd 0.003171f
C3616 vdd.n1569 gnd 0.00728f
C3617 vdd.n1570 gnd 0.00308f
C3618 vdd.n1571 gnd 0.003261f
C3619 vdd.n1572 gnd 0.005732f
C3620 vdd.n1573 gnd 0.00308f
C3621 vdd.n1574 gnd 0.00728f
C3622 vdd.n1575 gnd 0.003261f
C3623 vdd.n1576 gnd 0.005732f
C3624 vdd.n1577 gnd 0.00308f
C3625 vdd.n1578 gnd 0.00546f
C3626 vdd.n1579 gnd 0.005477f
C3627 vdd.t204 gnd 0.015641f
C3628 vdd.n1580 gnd 0.034801f
C3629 vdd.n1581 gnd 0.181113f
C3630 vdd.n1582 gnd 0.00308f
C3631 vdd.n1583 gnd 0.003261f
C3632 vdd.n1584 gnd 0.00728f
C3633 vdd.n1585 gnd 0.00728f
C3634 vdd.n1586 gnd 0.003261f
C3635 vdd.n1587 gnd 0.00308f
C3636 vdd.n1588 gnd 0.005732f
C3637 vdd.n1589 gnd 0.005732f
C3638 vdd.n1590 gnd 0.00308f
C3639 vdd.n1591 gnd 0.003261f
C3640 vdd.n1592 gnd 0.00728f
C3641 vdd.n1593 gnd 0.00728f
C3642 vdd.n1594 gnd 0.003261f
C3643 vdd.n1595 gnd 0.00308f
C3644 vdd.n1596 gnd 0.005732f
C3645 vdd.n1597 gnd 0.005732f
C3646 vdd.n1598 gnd 0.00308f
C3647 vdd.n1599 gnd 0.003261f
C3648 vdd.n1600 gnd 0.00728f
C3649 vdd.n1601 gnd 0.00728f
C3650 vdd.n1602 gnd 0.017212f
C3651 vdd.n1603 gnd 0.003171f
C3652 vdd.n1604 gnd 0.00308f
C3653 vdd.n1605 gnd 0.014815f
C3654 vdd.n1606 gnd 0.010019f
C3655 vdd.n1607 gnd 0.117581f
C3656 vdd.n1608 gnd 0.006177f
C3657 vdd.n1609 gnd 0.005732f
C3658 vdd.n1610 gnd 0.003171f
C3659 vdd.n1611 gnd 0.00728f
C3660 vdd.n1612 gnd 0.00308f
C3661 vdd.n1613 gnd 0.003261f
C3662 vdd.n1614 gnd 0.005732f
C3663 vdd.n1615 gnd 0.00308f
C3664 vdd.n1616 gnd 0.00728f
C3665 vdd.n1617 gnd 0.003261f
C3666 vdd.n1618 gnd 0.005732f
C3667 vdd.n1619 gnd 0.00308f
C3668 vdd.n1620 gnd 0.00546f
C3669 vdd.n1621 gnd 0.005477f
C3670 vdd.t269 gnd 0.015641f
C3671 vdd.n1622 gnd 0.034801f
C3672 vdd.n1623 gnd 0.181113f
C3673 vdd.n1624 gnd 0.00308f
C3674 vdd.n1625 gnd 0.003261f
C3675 vdd.n1626 gnd 0.00728f
C3676 vdd.n1627 gnd 0.00728f
C3677 vdd.n1628 gnd 0.003261f
C3678 vdd.n1629 gnd 0.00308f
C3679 vdd.n1630 gnd 0.005732f
C3680 vdd.n1631 gnd 0.005732f
C3681 vdd.n1632 gnd 0.00308f
C3682 vdd.n1633 gnd 0.003261f
C3683 vdd.n1634 gnd 0.00728f
C3684 vdd.n1635 gnd 0.00728f
C3685 vdd.n1636 gnd 0.003261f
C3686 vdd.n1637 gnd 0.00308f
C3687 vdd.n1638 gnd 0.005732f
C3688 vdd.n1639 gnd 0.005732f
C3689 vdd.n1640 gnd 0.00308f
C3690 vdd.n1641 gnd 0.003261f
C3691 vdd.n1642 gnd 0.00728f
C3692 vdd.n1643 gnd 0.00728f
C3693 vdd.n1644 gnd 0.017212f
C3694 vdd.n1645 gnd 0.003171f
C3695 vdd.n1646 gnd 0.00308f
C3696 vdd.n1647 gnd 0.014815f
C3697 vdd.n1648 gnd 0.010343f
C3698 vdd.t158 gnd 0.036237f
C3699 vdd.t272 gnd 0.036237f
C3700 vdd.n1649 gnd 0.249044f
C3701 vdd.n1650 gnd 0.195835f
C3702 vdd.t265 gnd 0.036237f
C3703 vdd.t251 gnd 0.036237f
C3704 vdd.n1651 gnd 0.249044f
C3705 vdd.n1652 gnd 0.158038f
C3706 vdd.t212 gnd 0.036237f
C3707 vdd.t147 gnd 0.036237f
C3708 vdd.n1653 gnd 0.249044f
C3709 vdd.n1654 gnd 0.158038f
C3710 vdd.t282 gnd 0.036237f
C3711 vdd.t249 gnd 0.036237f
C3712 vdd.n1655 gnd 0.249044f
C3713 vdd.n1656 gnd 0.158038f
C3714 vdd.t243 gnd 0.036237f
C3715 vdd.t189 gnd 0.036237f
C3716 vdd.n1657 gnd 0.249044f
C3717 vdd.n1658 gnd 0.158038f
C3718 vdd.t183 gnd 0.036237f
C3719 vdd.t244 gnd 0.036237f
C3720 vdd.n1659 gnd 0.249044f
C3721 vdd.n1660 gnd 0.158038f
C3722 vdd.t230 gnd 0.036237f
C3723 vdd.t228 gnd 0.036237f
C3724 vdd.n1661 gnd 0.249044f
C3725 vdd.n1662 gnd 0.158038f
C3726 vdd.t179 gnd 0.036237f
C3727 vdd.t154 gnd 0.036237f
C3728 vdd.n1663 gnd 0.249044f
C3729 vdd.n1664 gnd 0.158038f
C3730 vdd.t143 gnd 0.036237f
C3731 vdd.t223 gnd 0.036237f
C3732 vdd.n1665 gnd 0.249044f
C3733 vdd.n1666 gnd 0.158038f
C3734 vdd.n1667 gnd 0.006177f
C3735 vdd.n1668 gnd 0.005732f
C3736 vdd.n1669 gnd 0.003171f
C3737 vdd.n1670 gnd 0.00728f
C3738 vdd.n1671 gnd 0.00308f
C3739 vdd.n1672 gnd 0.003261f
C3740 vdd.n1673 gnd 0.005732f
C3741 vdd.n1674 gnd 0.00308f
C3742 vdd.n1675 gnd 0.00728f
C3743 vdd.n1676 gnd 0.003261f
C3744 vdd.n1677 gnd 0.005732f
C3745 vdd.n1678 gnd 0.00308f
C3746 vdd.n1679 gnd 0.00546f
C3747 vdd.n1680 gnd 0.005477f
C3748 vdd.t149 gnd 0.015641f
C3749 vdd.n1681 gnd 0.034801f
C3750 vdd.n1682 gnd 0.181113f
C3751 vdd.n1683 gnd 0.00308f
C3752 vdd.n1684 gnd 0.003261f
C3753 vdd.n1685 gnd 0.00728f
C3754 vdd.n1686 gnd 0.00728f
C3755 vdd.n1687 gnd 0.003261f
C3756 vdd.n1688 gnd 0.00308f
C3757 vdd.n1689 gnd 0.005732f
C3758 vdd.n1690 gnd 0.005732f
C3759 vdd.n1691 gnd 0.00308f
C3760 vdd.n1692 gnd 0.003261f
C3761 vdd.n1693 gnd 0.00728f
C3762 vdd.n1694 gnd 0.00728f
C3763 vdd.n1695 gnd 0.003261f
C3764 vdd.n1696 gnd 0.00308f
C3765 vdd.n1697 gnd 0.005732f
C3766 vdd.n1698 gnd 0.005732f
C3767 vdd.n1699 gnd 0.00308f
C3768 vdd.n1700 gnd 0.003261f
C3769 vdd.n1701 gnd 0.00728f
C3770 vdd.n1702 gnd 0.00728f
C3771 vdd.n1703 gnd 0.017212f
C3772 vdd.n1704 gnd 0.003171f
C3773 vdd.n1705 gnd 0.00308f
C3774 vdd.n1706 gnd 0.014815f
C3775 vdd.n1707 gnd 0.010019f
C3776 vdd.n1708 gnd 0.069949f
C3777 vdd.n1709 gnd 0.252044f
C3778 vdd.n1710 gnd 0.006177f
C3779 vdd.n1711 gnd 0.005732f
C3780 vdd.n1712 gnd 0.003171f
C3781 vdd.n1713 gnd 0.00728f
C3782 vdd.n1714 gnd 0.00308f
C3783 vdd.n1715 gnd 0.003261f
C3784 vdd.n1716 gnd 0.005732f
C3785 vdd.n1717 gnd 0.00308f
C3786 vdd.n1718 gnd 0.00728f
C3787 vdd.n1719 gnd 0.003261f
C3788 vdd.n1720 gnd 0.005732f
C3789 vdd.n1721 gnd 0.00308f
C3790 vdd.n1722 gnd 0.00546f
C3791 vdd.n1723 gnd 0.005477f
C3792 vdd.t283 gnd 0.015641f
C3793 vdd.n1724 gnd 0.034801f
C3794 vdd.n1725 gnd 0.181113f
C3795 vdd.n1726 gnd 0.00308f
C3796 vdd.n1727 gnd 0.003261f
C3797 vdd.n1728 gnd 0.00728f
C3798 vdd.n1729 gnd 0.00728f
C3799 vdd.n1730 gnd 0.003261f
C3800 vdd.n1731 gnd 0.00308f
C3801 vdd.n1732 gnd 0.005732f
C3802 vdd.n1733 gnd 0.005732f
C3803 vdd.n1734 gnd 0.00308f
C3804 vdd.n1735 gnd 0.003261f
C3805 vdd.n1736 gnd 0.00728f
C3806 vdd.n1737 gnd 0.00728f
C3807 vdd.n1738 gnd 0.003261f
C3808 vdd.n1739 gnd 0.00308f
C3809 vdd.n1740 gnd 0.005732f
C3810 vdd.n1741 gnd 0.005732f
C3811 vdd.n1742 gnd 0.00308f
C3812 vdd.n1743 gnd 0.003261f
C3813 vdd.n1744 gnd 0.00728f
C3814 vdd.n1745 gnd 0.00728f
C3815 vdd.n1746 gnd 0.017212f
C3816 vdd.n1747 gnd 0.003171f
C3817 vdd.n1748 gnd 0.00308f
C3818 vdd.n1749 gnd 0.014815f
C3819 vdd.n1750 gnd 0.010343f
C3820 vdd.t175 gnd 0.036237f
C3821 vdd.t284 gnd 0.036237f
C3822 vdd.n1751 gnd 0.249044f
C3823 vdd.n1752 gnd 0.195835f
C3824 vdd.t281 gnd 0.036237f
C3825 vdd.t262 gnd 0.036237f
C3826 vdd.n1753 gnd 0.249044f
C3827 vdd.n1754 gnd 0.158038f
C3828 vdd.t231 gnd 0.036237f
C3829 vdd.t171 gnd 0.036237f
C3830 vdd.n1755 gnd 0.249044f
C3831 vdd.n1756 gnd 0.158038f
C3832 vdd.t293 gnd 0.036237f
C3833 vdd.t259 gnd 0.036237f
C3834 vdd.n1757 gnd 0.249044f
C3835 vdd.n1758 gnd 0.158038f
C3836 vdd.t257 gnd 0.036237f
C3837 vdd.t205 gnd 0.036237f
C3838 vdd.n1759 gnd 0.249044f
C3839 vdd.n1760 gnd 0.158038f
C3840 vdd.t201 gnd 0.036237f
C3841 vdd.t232 gnd 0.036237f
C3842 vdd.n1761 gnd 0.249044f
C3843 vdd.n1762 gnd 0.158038f
C3844 vdd.t233 gnd 0.036237f
C3845 vdd.t242 gnd 0.036237f
C3846 vdd.n1763 gnd 0.249044f
C3847 vdd.n1764 gnd 0.158038f
C3848 vdd.t198 gnd 0.036237f
C3849 vdd.t174 gnd 0.036237f
C3850 vdd.n1765 gnd 0.249044f
C3851 vdd.n1766 gnd 0.158038f
C3852 vdd.t170 gnd 0.036237f
C3853 vdd.t239 gnd 0.036237f
C3854 vdd.n1767 gnd 0.249044f
C3855 vdd.n1768 gnd 0.158038f
C3856 vdd.n1769 gnd 0.006177f
C3857 vdd.n1770 gnd 0.005732f
C3858 vdd.n1771 gnd 0.003171f
C3859 vdd.n1772 gnd 0.00728f
C3860 vdd.n1773 gnd 0.00308f
C3861 vdd.n1774 gnd 0.003261f
C3862 vdd.n1775 gnd 0.005732f
C3863 vdd.n1776 gnd 0.00308f
C3864 vdd.n1777 gnd 0.00728f
C3865 vdd.n1778 gnd 0.003261f
C3866 vdd.n1779 gnd 0.005732f
C3867 vdd.n1780 gnd 0.00308f
C3868 vdd.n1781 gnd 0.00546f
C3869 vdd.n1782 gnd 0.005477f
C3870 vdd.t172 gnd 0.015641f
C3871 vdd.n1783 gnd 0.034801f
C3872 vdd.n1784 gnd 0.181113f
C3873 vdd.n1785 gnd 0.00308f
C3874 vdd.n1786 gnd 0.003261f
C3875 vdd.n1787 gnd 0.00728f
C3876 vdd.n1788 gnd 0.00728f
C3877 vdd.n1789 gnd 0.003261f
C3878 vdd.n1790 gnd 0.00308f
C3879 vdd.n1791 gnd 0.005732f
C3880 vdd.n1792 gnd 0.005732f
C3881 vdd.n1793 gnd 0.00308f
C3882 vdd.n1794 gnd 0.003261f
C3883 vdd.n1795 gnd 0.00728f
C3884 vdd.n1796 gnd 0.00728f
C3885 vdd.n1797 gnd 0.003261f
C3886 vdd.n1798 gnd 0.00308f
C3887 vdd.n1799 gnd 0.005732f
C3888 vdd.n1800 gnd 0.005732f
C3889 vdd.n1801 gnd 0.00308f
C3890 vdd.n1802 gnd 0.003261f
C3891 vdd.n1803 gnd 0.00728f
C3892 vdd.n1804 gnd 0.00728f
C3893 vdd.n1805 gnd 0.017212f
C3894 vdd.n1806 gnd 0.003171f
C3895 vdd.n1807 gnd 0.00308f
C3896 vdd.n1808 gnd 0.014815f
C3897 vdd.n1809 gnd 0.010019f
C3898 vdd.n1810 gnd 0.069949f
C3899 vdd.n1811 gnd 0.288535f
C3900 vdd.n1812 gnd 2.89082f
C3901 vdd.n1813 gnd 0.663882f
C3902 vdd.n1814 gnd 0.00865f
C3903 vdd.n1815 gnd 0.009059f
C3904 vdd.n1816 gnd 0.011255f
C3905 vdd.n1817 gnd 0.822423f
C3906 vdd.n1818 gnd 0.011255f
C3907 vdd.n1819 gnd 0.009059f
C3908 vdd.n1820 gnd 0.011255f
C3909 vdd.n1821 gnd 0.011255f
C3910 vdd.n1822 gnd 0.011255f
C3911 vdd.n1823 gnd 0.009059f
C3912 vdd.n1824 gnd 0.011255f
C3913 vdd.n1825 gnd 0.954701f
C3914 vdd.t234 gnd 0.575121f
C3915 vdd.n1826 gnd 0.626882f
C3916 vdd.n1827 gnd 0.011255f
C3917 vdd.n1828 gnd 0.009059f
C3918 vdd.n1829 gnd 0.011255f
C3919 vdd.n1830 gnd 0.011255f
C3920 vdd.n1831 gnd 0.011255f
C3921 vdd.n1832 gnd 0.009059f
C3922 vdd.n1833 gnd 0.011255f
C3923 vdd.n1834 gnd 0.718901f
C3924 vdd.n1835 gnd 0.011255f
C3925 vdd.n1836 gnd 0.009059f
C3926 vdd.n1837 gnd 0.011255f
C3927 vdd.n1838 gnd 0.011255f
C3928 vdd.n1839 gnd 0.011255f
C3929 vdd.n1840 gnd 0.009059f
C3930 vdd.n1841 gnd 0.011255f
C3931 vdd.n1842 gnd 0.615379f
C3932 vdd.n1843 gnd 0.914442f
C3933 vdd.n1844 gnd 0.011255f
C3934 vdd.n1845 gnd 0.009059f
C3935 vdd.n1846 gnd 0.011255f
C3936 vdd.n1847 gnd 0.011255f
C3937 vdd.n1848 gnd 0.011255f
C3938 vdd.n1849 gnd 0.009059f
C3939 vdd.n1850 gnd 0.011255f
C3940 vdd.n1851 gnd 0.954701f
C3941 vdd.n1852 gnd 0.011255f
C3942 vdd.n1853 gnd 0.009059f
C3943 vdd.n1854 gnd 0.011255f
C3944 vdd.n1855 gnd 0.011255f
C3945 vdd.n1856 gnd 0.011255f
C3946 vdd.n1857 gnd 0.009059f
C3947 vdd.n1858 gnd 0.011255f
C3948 vdd.t250 gnd 0.575121f
C3949 vdd.n1859 gnd 0.799418f
C3950 vdd.n1860 gnd 0.011255f
C3951 vdd.n1861 gnd 0.009059f
C3952 vdd.n1862 gnd 0.011255f
C3953 vdd.n1863 gnd 0.011255f
C3954 vdd.n1864 gnd 0.011255f
C3955 vdd.n1865 gnd 0.009059f
C3956 vdd.n1866 gnd 0.011255f
C3957 vdd.n1867 gnd 0.603877f
C3958 vdd.n1868 gnd 0.011255f
C3959 vdd.n1869 gnd 0.009059f
C3960 vdd.n1870 gnd 0.011255f
C3961 vdd.n1871 gnd 0.011255f
C3962 vdd.n1872 gnd 0.011255f
C3963 vdd.n1873 gnd 0.009059f
C3964 vdd.n1874 gnd 0.011255f
C3965 vdd.n1875 gnd 0.787916f
C3966 vdd.n1876 gnd 0.741906f
C3967 vdd.n1877 gnd 0.011255f
C3968 vdd.n1878 gnd 0.009059f
C3969 vdd.n1879 gnd 0.011255f
C3970 vdd.n1880 gnd 0.011255f
C3971 vdd.n1881 gnd 0.011255f
C3972 vdd.n1882 gnd 0.009059f
C3973 vdd.n1883 gnd 0.011255f
C3974 vdd.n1884 gnd 0.937447f
C3975 vdd.n1885 gnd 0.011255f
C3976 vdd.n1886 gnd 0.009059f
C3977 vdd.n1887 gnd 0.011255f
C3978 vdd.n1888 gnd 0.011255f
C3979 vdd.n1889 gnd 0.027228f
C3980 vdd.n1890 gnd 0.011255f
C3981 vdd.n1891 gnd 0.011255f
C3982 vdd.n1892 gnd 0.009059f
C3983 vdd.n1893 gnd 0.011255f
C3984 vdd.n1894 gnd 0.695896f
C3985 vdd.n1895 gnd 1.15024f
C3986 vdd.n1896 gnd 0.011255f
C3987 vdd.n1897 gnd 0.009059f
C3988 vdd.n1898 gnd 0.011255f
C3989 vdd.n1899 gnd 0.011255f
C3990 vdd.n1900 gnd 0.00968f
C3991 vdd.n1901 gnd 0.009059f
C3992 vdd.n1903 gnd 0.011255f
C3993 vdd.n1905 gnd 0.009059f
C3994 vdd.n1906 gnd 0.011255f
C3995 vdd.n1907 gnd 0.009059f
C3996 vdd.n1909 gnd 0.011255f
C3997 vdd.n1910 gnd 0.009059f
C3998 vdd.n1911 gnd 0.011255f
C3999 vdd.n1912 gnd 0.011255f
C4000 vdd.n1913 gnd 0.011255f
C4001 vdd.n1914 gnd 0.011255f
C4002 vdd.n1915 gnd 0.011255f
C4003 vdd.n1916 gnd 0.009059f
C4004 vdd.n1918 gnd 0.011255f
C4005 vdd.n1919 gnd 0.011255f
C4006 vdd.n1920 gnd 0.011255f
C4007 vdd.n1921 gnd 0.011255f
C4008 vdd.n1922 gnd 0.011255f
C4009 vdd.n1923 gnd 0.009059f
C4010 vdd.n1925 gnd 0.011255f
C4011 vdd.n1926 gnd 0.011255f
C4012 vdd.n1927 gnd 0.011255f
C4013 vdd.n1928 gnd 0.011255f
C4014 vdd.n1929 gnd 0.007564f
C4015 vdd.t92 gnd 0.13847f
C4016 vdd.t91 gnd 0.147986f
C4017 vdd.t90 gnd 0.18084f
C4018 vdd.n1930 gnd 0.231812f
C4019 vdd.n1931 gnd 0.194764f
C4020 vdd.n1933 gnd 0.011255f
C4021 vdd.n1934 gnd 0.011255f
C4022 vdd.n1935 gnd 0.009059f
C4023 vdd.n1936 gnd 0.011255f
C4024 vdd.n1938 gnd 0.011255f
C4025 vdd.n1939 gnd 0.011255f
C4026 vdd.n1940 gnd 0.011255f
C4027 vdd.n1941 gnd 0.011255f
C4028 vdd.n1942 gnd 0.009059f
C4029 vdd.n1944 gnd 0.011255f
C4030 vdd.n1945 gnd 0.011255f
C4031 vdd.n1946 gnd 0.011255f
C4032 vdd.n1947 gnd 0.011255f
C4033 vdd.n1948 gnd 0.011255f
C4034 vdd.n1949 gnd 0.009059f
C4035 vdd.n1951 gnd 0.011255f
C4036 vdd.n1952 gnd 0.011255f
C4037 vdd.n1953 gnd 0.011255f
C4038 vdd.n1954 gnd 0.011255f
C4039 vdd.n1955 gnd 0.011255f
C4040 vdd.n1956 gnd 0.009059f
C4041 vdd.n1958 gnd 0.011255f
C4042 vdd.n1959 gnd 0.011255f
C4043 vdd.n1960 gnd 0.011255f
C4044 vdd.n1961 gnd 0.011255f
C4045 vdd.n1962 gnd 0.011255f
C4046 vdd.n1963 gnd 0.009059f
C4047 vdd.n1965 gnd 0.011255f
C4048 vdd.n1966 gnd 0.011255f
C4049 vdd.n1967 gnd 0.011255f
C4050 vdd.n1968 gnd 0.011255f
C4051 vdd.n1969 gnd 0.008969f
C4052 vdd.t79 gnd 0.13847f
C4053 vdd.t78 gnd 0.147986f
C4054 vdd.t77 gnd 0.18084f
C4055 vdd.n1970 gnd 0.231812f
C4056 vdd.n1971 gnd 0.194764f
C4057 vdd.n1973 gnd 0.011255f
C4058 vdd.n1974 gnd 0.011255f
C4059 vdd.n1975 gnd 0.009059f
C4060 vdd.n1976 gnd 0.011255f
C4061 vdd.n1978 gnd 0.011255f
C4062 vdd.n1979 gnd 0.011255f
C4063 vdd.n1980 gnd 0.011255f
C4064 vdd.n1981 gnd 0.011255f
C4065 vdd.n1982 gnd 0.009059f
C4066 vdd.n1984 gnd 0.011255f
C4067 vdd.n1985 gnd 0.011255f
C4068 vdd.n1986 gnd 0.011255f
C4069 vdd.n1987 gnd 0.011255f
C4070 vdd.n1988 gnd 0.011255f
C4071 vdd.n1989 gnd 0.009059f
C4072 vdd.n1991 gnd 0.011255f
C4073 vdd.n1992 gnd 0.011255f
C4074 vdd.n1993 gnd 0.011255f
C4075 vdd.n1994 gnd 0.011255f
C4076 vdd.n1995 gnd 0.011255f
C4077 vdd.n1996 gnd 0.011255f
C4078 vdd.n1997 gnd 0.009059f
C4079 vdd.n1999 gnd 0.011255f
C4080 vdd.n2001 gnd 0.011255f
C4081 vdd.n2002 gnd 0.009059f
C4082 vdd.n2003 gnd 0.009059f
C4083 vdd.n2004 gnd 0.011255f
C4084 vdd.n2006 gnd 0.011255f
C4085 vdd.n2007 gnd 0.009059f
C4086 vdd.n2008 gnd 0.009059f
C4087 vdd.n2009 gnd 0.011255f
C4088 vdd.n2011 gnd 0.011255f
C4089 vdd.n2012 gnd 0.011255f
C4090 vdd.n2013 gnd 0.009059f
C4091 vdd.n2014 gnd 0.009059f
C4092 vdd.n2015 gnd 0.009059f
C4093 vdd.n2016 gnd 0.011255f
C4094 vdd.n2018 gnd 0.011255f
C4095 vdd.n2019 gnd 0.011255f
C4096 vdd.n2020 gnd 0.009059f
C4097 vdd.n2021 gnd 0.009059f
C4098 vdd.n2022 gnd 0.009059f
C4099 vdd.n2023 gnd 0.011255f
C4100 vdd.n2025 gnd 0.011255f
C4101 vdd.n2026 gnd 0.011255f
C4102 vdd.n2027 gnd 0.009059f
C4103 vdd.n2028 gnd 0.009059f
C4104 vdd.n2029 gnd 0.009059f
C4105 vdd.n2030 gnd 0.011255f
C4106 vdd.n2032 gnd 0.011255f
C4107 vdd.n2033 gnd 0.011255f
C4108 vdd.n2034 gnd 0.009059f
C4109 vdd.n2035 gnd 0.011255f
C4110 vdd.n2036 gnd 0.011255f
C4111 vdd.n2037 gnd 0.011255f
C4112 vdd.n2038 gnd 0.018481f
C4113 vdd.n2039 gnd 0.00616f
C4114 vdd.n2040 gnd 0.009059f
C4115 vdd.n2041 gnd 0.011255f
C4116 vdd.n2043 gnd 0.011255f
C4117 vdd.n2044 gnd 0.011255f
C4118 vdd.n2045 gnd 0.009059f
C4119 vdd.n2046 gnd 0.009059f
C4120 vdd.n2047 gnd 0.009059f
C4121 vdd.n2048 gnd 0.011255f
C4122 vdd.n2050 gnd 0.011255f
C4123 vdd.n2051 gnd 0.011255f
C4124 vdd.n2052 gnd 0.009059f
C4125 vdd.n2053 gnd 0.009059f
C4126 vdd.n2054 gnd 0.009059f
C4127 vdd.n2055 gnd 0.011255f
C4128 vdd.n2057 gnd 0.011255f
C4129 vdd.n2058 gnd 0.011255f
C4130 vdd.n2059 gnd 0.009059f
C4131 vdd.n2060 gnd 0.009059f
C4132 vdd.n2061 gnd 0.009059f
C4133 vdd.n2062 gnd 0.011255f
C4134 vdd.n2064 gnd 0.011255f
C4135 vdd.n2065 gnd 0.011255f
C4136 vdd.n2066 gnd 0.009059f
C4137 vdd.n2067 gnd 0.009059f
C4138 vdd.n2068 gnd 0.009059f
C4139 vdd.n2069 gnd 0.011255f
C4140 vdd.n2071 gnd 0.011255f
C4141 vdd.n2072 gnd 0.011255f
C4142 vdd.n2073 gnd 0.009059f
C4143 vdd.n2074 gnd 0.011255f
C4144 vdd.n2075 gnd 0.011255f
C4145 vdd.n2076 gnd 0.011255f
C4146 vdd.n2077 gnd 0.018481f
C4147 vdd.n2078 gnd 0.007564f
C4148 vdd.n2079 gnd 0.009059f
C4149 vdd.n2080 gnd 0.011255f
C4150 vdd.n2082 gnd 0.011255f
C4151 vdd.n2083 gnd 0.011255f
C4152 vdd.n2084 gnd 0.009059f
C4153 vdd.n2085 gnd 0.009059f
C4154 vdd.n2086 gnd 0.009059f
C4155 vdd.n2087 gnd 0.011255f
C4156 vdd.n2089 gnd 0.011255f
C4157 vdd.n2090 gnd 0.011255f
C4158 vdd.n2091 gnd 0.009059f
C4159 vdd.n2092 gnd 0.009059f
C4160 vdd.n2093 gnd 0.009059f
C4161 vdd.n2094 gnd 0.011255f
C4162 vdd.n2096 gnd 0.011255f
C4163 vdd.n2097 gnd 0.011255f
C4164 vdd.n2099 gnd 0.011255f
C4165 vdd.n2100 gnd 0.009059f
C4166 vdd.n2101 gnd 0.007203f
C4167 vdd.n2102 gnd 0.007654f
C4168 vdd.n2103 gnd 0.007654f
C4169 vdd.n2104 gnd 0.007654f
C4170 vdd.n2105 gnd 0.007654f
C4171 vdd.n2106 gnd 0.007654f
C4172 vdd.n2107 gnd 0.007654f
C4173 vdd.n2108 gnd 0.007654f
C4174 vdd.n2109 gnd 0.007654f
C4175 vdd.n2111 gnd 0.007654f
C4176 vdd.n2112 gnd 0.007654f
C4177 vdd.n2113 gnd 0.007654f
C4178 vdd.n2114 gnd 0.007654f
C4179 vdd.n2115 gnd 0.007654f
C4180 vdd.n2117 gnd 0.007654f
C4181 vdd.n2119 gnd 0.007654f
C4182 vdd.n2120 gnd 0.007654f
C4183 vdd.n2121 gnd 0.007654f
C4184 vdd.n2122 gnd 0.007654f
C4185 vdd.n2123 gnd 0.007654f
C4186 vdd.n2125 gnd 0.007654f
C4187 vdd.n2127 gnd 0.007654f
C4188 vdd.n2128 gnd 0.007654f
C4189 vdd.n2129 gnd 0.007654f
C4190 vdd.n2130 gnd 0.007654f
C4191 vdd.n2131 gnd 0.007654f
C4192 vdd.n2133 gnd 0.007654f
C4193 vdd.n2135 gnd 0.007654f
C4194 vdd.n2136 gnd 0.007654f
C4195 vdd.n2137 gnd 0.007654f
C4196 vdd.n2138 gnd 0.007654f
C4197 vdd.n2139 gnd 0.007654f
C4198 vdd.n2141 gnd 0.007654f
C4199 vdd.n2142 gnd 0.007654f
C4200 vdd.n2143 gnd 0.007654f
C4201 vdd.n2144 gnd 0.007654f
C4202 vdd.n2145 gnd 0.007654f
C4203 vdd.n2146 gnd 0.007654f
C4204 vdd.n2147 gnd 0.007654f
C4205 vdd.n2148 gnd 0.007654f
C4206 vdd.n2149 gnd 0.005571f
C4207 vdd.n2150 gnd 0.007654f
C4208 vdd.t56 gnd 0.309282f
C4209 vdd.t57 gnd 0.316589f
C4210 vdd.t54 gnd 0.201911f
C4211 vdd.n2151 gnd 0.109122f
C4212 vdd.n2152 gnd 0.061898f
C4213 vdd.n2153 gnd 0.010938f
C4214 vdd.n2154 gnd 0.007654f
C4215 vdd.n2155 gnd 0.007654f
C4216 vdd.n2156 gnd 0.465848f
C4217 vdd.n2157 gnd 0.007654f
C4218 vdd.n2158 gnd 0.007654f
C4219 vdd.n2159 gnd 0.007654f
C4220 vdd.n2160 gnd 0.007654f
C4221 vdd.n2161 gnd 0.007654f
C4222 vdd.n2162 gnd 0.007654f
C4223 vdd.n2163 gnd 0.007654f
C4224 vdd.n2164 gnd 0.007654f
C4225 vdd.n2165 gnd 0.007654f
C4226 vdd.n2166 gnd 0.007654f
C4227 vdd.n2167 gnd 0.007654f
C4228 vdd.n2168 gnd 0.007654f
C4229 vdd.n2169 gnd 0.007654f
C4230 vdd.n2170 gnd 0.007654f
C4231 vdd.n2171 gnd 0.007654f
C4232 vdd.n2172 gnd 0.007654f
C4233 vdd.n2173 gnd 0.007654f
C4234 vdd.n2174 gnd 0.007654f
C4235 vdd.n2175 gnd 0.007654f
C4236 vdd.n2176 gnd 0.007654f
C4237 vdd.t109 gnd 0.309282f
C4238 vdd.t110 gnd 0.316589f
C4239 vdd.t108 gnd 0.201911f
C4240 vdd.n2177 gnd 0.109122f
C4241 vdd.n2178 gnd 0.061898f
C4242 vdd.n2179 gnd 0.007654f
C4243 vdd.n2180 gnd 0.007654f
C4244 vdd.n2181 gnd 0.007654f
C4245 vdd.n2182 gnd 0.007654f
C4246 vdd.n2183 gnd 0.007654f
C4247 vdd.n2184 gnd 0.007654f
C4248 vdd.n2186 gnd 0.007654f
C4249 vdd.n2187 gnd 0.007654f
C4250 vdd.n2188 gnd 0.007654f
C4251 vdd.n2189 gnd 0.007654f
C4252 vdd.n2191 gnd 0.007654f
C4253 vdd.n2193 gnd 0.007654f
C4254 vdd.n2194 gnd 0.007654f
C4255 vdd.n2195 gnd 0.007654f
C4256 vdd.n2196 gnd 0.007654f
C4257 vdd.n2197 gnd 0.007654f
C4258 vdd.n2199 gnd 0.007654f
C4259 vdd.n2201 gnd 0.007654f
C4260 vdd.n2202 gnd 0.007654f
C4261 vdd.n2203 gnd 0.007654f
C4262 vdd.n2204 gnd 0.007654f
C4263 vdd.n2205 gnd 0.007654f
C4264 vdd.n2207 gnd 0.007654f
C4265 vdd.n2209 gnd 0.007654f
C4266 vdd.n2210 gnd 0.007654f
C4267 vdd.n2211 gnd 0.005571f
C4268 vdd.n2212 gnd 0.010938f
C4269 vdd.n2213 gnd 0.005909f
C4270 vdd.n2214 gnd 0.007654f
C4271 vdd.n2216 gnd 0.007654f
C4272 vdd.n2217 gnd 0.018161f
C4273 vdd.n2218 gnd 0.018161f
C4274 vdd.n2219 gnd 0.016956f
C4275 vdd.n2220 gnd 0.007654f
C4276 vdd.n2221 gnd 0.007654f
C4277 vdd.n2222 gnd 0.007654f
C4278 vdd.n2223 gnd 0.007654f
C4279 vdd.n2224 gnd 0.007654f
C4280 vdd.n2225 gnd 0.007654f
C4281 vdd.n2226 gnd 0.007654f
C4282 vdd.n2227 gnd 0.007654f
C4283 vdd.n2228 gnd 0.007654f
C4284 vdd.n2229 gnd 0.007654f
C4285 vdd.n2230 gnd 0.007654f
C4286 vdd.n2231 gnd 0.007654f
C4287 vdd.n2232 gnd 0.007654f
C4288 vdd.n2233 gnd 0.007654f
C4289 vdd.n2234 gnd 0.007654f
C4290 vdd.n2235 gnd 0.007654f
C4291 vdd.n2236 gnd 0.007654f
C4292 vdd.n2237 gnd 0.007654f
C4293 vdd.n2238 gnd 0.007654f
C4294 vdd.n2239 gnd 0.007654f
C4295 vdd.n2240 gnd 0.007654f
C4296 vdd.n2241 gnd 0.007654f
C4297 vdd.n2242 gnd 0.007654f
C4298 vdd.n2243 gnd 0.007654f
C4299 vdd.n2244 gnd 0.007654f
C4300 vdd.n2245 gnd 0.007654f
C4301 vdd.n2246 gnd 0.007654f
C4302 vdd.n2247 gnd 0.007654f
C4303 vdd.n2248 gnd 0.007654f
C4304 vdd.n2249 gnd 0.007654f
C4305 vdd.n2250 gnd 0.007654f
C4306 vdd.n2251 gnd 0.007654f
C4307 vdd.n2252 gnd 0.007654f
C4308 vdd.n2253 gnd 0.007654f
C4309 vdd.n2254 gnd 0.007654f
C4310 vdd.n2255 gnd 0.007654f
C4311 vdd.n2256 gnd 0.007654f
C4312 vdd.n2257 gnd 0.247302f
C4313 vdd.n2258 gnd 0.007654f
C4314 vdd.n2259 gnd 0.007654f
C4315 vdd.n2260 gnd 0.007654f
C4316 vdd.n2261 gnd 0.007654f
C4317 vdd.n2262 gnd 0.007654f
C4318 vdd.n2263 gnd 0.007654f
C4319 vdd.n2264 gnd 0.007654f
C4320 vdd.n2265 gnd 0.007654f
C4321 vdd.n2266 gnd 0.007654f
C4322 vdd.n2267 gnd 0.007654f
C4323 vdd.n2268 gnd 0.007654f
C4324 vdd.n2269 gnd 0.007654f
C4325 vdd.n2270 gnd 0.007654f
C4326 vdd.n2271 gnd 0.007654f
C4327 vdd.n2272 gnd 0.007654f
C4328 vdd.n2273 gnd 0.007654f
C4329 vdd.n2274 gnd 0.007654f
C4330 vdd.n2275 gnd 0.007654f
C4331 vdd.n2276 gnd 0.007654f
C4332 vdd.n2277 gnd 0.007654f
C4333 vdd.n2278 gnd 0.016956f
C4334 vdd.n2280 gnd 0.018161f
C4335 vdd.n2281 gnd 0.018161f
C4336 vdd.n2282 gnd 0.007654f
C4337 vdd.n2283 gnd 0.005909f
C4338 vdd.n2284 gnd 0.007654f
C4339 vdd.n2286 gnd 0.007654f
C4340 vdd.n2288 gnd 0.007654f
C4341 vdd.n2289 gnd 0.007654f
C4342 vdd.n2290 gnd 0.007654f
C4343 vdd.n2291 gnd 0.007654f
C4344 vdd.n2292 gnd 0.007654f
C4345 vdd.n2294 gnd 0.007654f
C4346 vdd.n2296 gnd 0.007654f
C4347 vdd.n2297 gnd 0.007654f
C4348 vdd.n2298 gnd 0.007654f
C4349 vdd.n2299 gnd 0.007654f
C4350 vdd.n2300 gnd 0.007654f
C4351 vdd.n2302 gnd 0.007654f
C4352 vdd.n2304 gnd 0.007654f
C4353 vdd.n2305 gnd 0.007654f
C4354 vdd.n2306 gnd 0.007654f
C4355 vdd.n2307 gnd 0.007654f
C4356 vdd.n2308 gnd 0.007654f
C4357 vdd.n2310 gnd 0.007654f
C4358 vdd.n2312 gnd 0.007654f
C4359 vdd.n2313 gnd 0.007654f
C4360 vdd.n2314 gnd 0.022829f
C4361 vdd.n2315 gnd 0.676754f
C4362 vdd.n2317 gnd 0.009059f
C4363 vdd.n2318 gnd 0.009059f
C4364 vdd.n2319 gnd 0.011255f
C4365 vdd.n2321 gnd 0.011255f
C4366 vdd.n2322 gnd 0.011255f
C4367 vdd.n2323 gnd 0.009059f
C4368 vdd.n2324 gnd 0.007519f
C4369 vdd.n2325 gnd 0.027811f
C4370 vdd.n2326 gnd 0.027228f
C4371 vdd.n2327 gnd 0.007519f
C4372 vdd.n2328 gnd 0.027228f
C4373 vdd.n2329 gnd 1.58158f
C4374 vdd.n2330 gnd 0.027228f
C4375 vdd.n2331 gnd 0.027811f
C4376 vdd.n2332 gnd 0.004303f
C4377 vdd.t68 gnd 0.13847f
C4378 vdd.t67 gnd 0.147986f
C4379 vdd.t65 gnd 0.18084f
C4380 vdd.n2333 gnd 0.231812f
C4381 vdd.n2334 gnd 0.194764f
C4382 vdd.n2335 gnd 0.013951f
C4383 vdd.n2336 gnd 0.004756f
C4384 vdd.n2337 gnd 0.00968f
C4385 vdd.n2338 gnd 0.676754f
C4386 vdd.n2339 gnd 0.022829f
C4387 vdd.n2340 gnd 0.007654f
C4388 vdd.n2341 gnd 0.007654f
C4389 vdd.n2342 gnd 0.007654f
C4390 vdd.n2344 gnd 0.007654f
C4391 vdd.n2346 gnd 0.007654f
C4392 vdd.n2347 gnd 0.007654f
C4393 vdd.n2348 gnd 0.007654f
C4394 vdd.n2349 gnd 0.007654f
C4395 vdd.n2350 gnd 0.007654f
C4396 vdd.n2352 gnd 0.007654f
C4397 vdd.n2354 gnd 0.007654f
C4398 vdd.n2355 gnd 0.007654f
C4399 vdd.n2356 gnd 0.007654f
C4400 vdd.n2357 gnd 0.007654f
C4401 vdd.n2358 gnd 0.007654f
C4402 vdd.n2360 gnd 0.007654f
C4403 vdd.n2362 gnd 0.007654f
C4404 vdd.n2363 gnd 0.007654f
C4405 vdd.n2364 gnd 0.007654f
C4406 vdd.n2365 gnd 0.007654f
C4407 vdd.n2366 gnd 0.007654f
C4408 vdd.n2368 gnd 0.007654f
C4409 vdd.n2370 gnd 0.007654f
C4410 vdd.n2371 gnd 0.007654f
C4411 vdd.n2372 gnd 0.018161f
C4412 vdd.n2373 gnd 0.016956f
C4413 vdd.n2374 gnd 0.016956f
C4414 vdd.n2375 gnd 1.12724f
C4415 vdd.n2376 gnd 0.016956f
C4416 vdd.n2377 gnd 0.016956f
C4417 vdd.n2378 gnd 0.007654f
C4418 vdd.n2379 gnd 0.007654f
C4419 vdd.n2380 gnd 0.007654f
C4420 vdd.n2381 gnd 0.488853f
C4421 vdd.n2382 gnd 0.007654f
C4422 vdd.n2383 gnd 0.007654f
C4423 vdd.n2384 gnd 0.007654f
C4424 vdd.n2385 gnd 0.007654f
C4425 vdd.n2386 gnd 0.007654f
C4426 vdd.n2387 gnd 0.782164f
C4427 vdd.n2388 gnd 0.007654f
C4428 vdd.n2389 gnd 0.007654f
C4429 vdd.n2390 gnd 0.007654f
C4430 vdd.n2391 gnd 0.007654f
C4431 vdd.n2392 gnd 0.007654f
C4432 vdd.n2393 gnd 0.782164f
C4433 vdd.n2394 gnd 0.007654f
C4434 vdd.n2395 gnd 0.007654f
C4435 vdd.n2396 gnd 0.006753f
C4436 vdd.n2397 gnd 0.022172f
C4437 vdd.n2398 gnd 0.004727f
C4438 vdd.n2399 gnd 0.007654f
C4439 vdd.n2400 gnd 0.431341f
C4440 vdd.n2401 gnd 0.007654f
C4441 vdd.n2402 gnd 0.007654f
C4442 vdd.n2403 gnd 0.007654f
C4443 vdd.n2404 gnd 0.007654f
C4444 vdd.n2405 gnd 0.007654f
C4445 vdd.n2406 gnd 0.52336f
C4446 vdd.n2407 gnd 0.007654f
C4447 vdd.n2408 gnd 0.007654f
C4448 vdd.n2409 gnd 0.007654f
C4449 vdd.n2410 gnd 0.007654f
C4450 vdd.n2411 gnd 0.007654f
C4451 vdd.n2412 gnd 0.695896f
C4452 vdd.n2413 gnd 0.007654f
C4453 vdd.n2414 gnd 0.007654f
C4454 vdd.n2415 gnd 0.007654f
C4455 vdd.n2416 gnd 0.007654f
C4456 vdd.n2417 gnd 0.007654f
C4457 vdd.n2418 gnd 0.621131f
C4458 vdd.n2419 gnd 0.007654f
C4459 vdd.n2420 gnd 0.007654f
C4460 vdd.n2421 gnd 0.007654f
C4461 vdd.n2422 gnd 0.007654f
C4462 vdd.n2423 gnd 0.007654f
C4463 vdd.n2424 gnd 0.448594f
C4464 vdd.n2425 gnd 0.007654f
C4465 vdd.n2426 gnd 0.007654f
C4466 vdd.n2427 gnd 0.007654f
C4467 vdd.n2428 gnd 0.007654f
C4468 vdd.n2429 gnd 0.007654f
C4469 vdd.n2430 gnd 0.247302f
C4470 vdd.n2431 gnd 0.007654f
C4471 vdd.n2432 gnd 0.007654f
C4472 vdd.n2433 gnd 0.007654f
C4473 vdd.n2434 gnd 0.007654f
C4474 vdd.n2435 gnd 0.007654f
C4475 vdd.n2436 gnd 0.431341f
C4476 vdd.n2437 gnd 0.007654f
C4477 vdd.n2438 gnd 0.007654f
C4478 vdd.n2439 gnd 0.007654f
C4479 vdd.n2440 gnd 0.007654f
C4480 vdd.n2441 gnd 0.007654f
C4481 vdd.n2442 gnd 0.782164f
C4482 vdd.n2443 gnd 0.007654f
C4483 vdd.n2444 gnd 0.007654f
C4484 vdd.n2445 gnd 0.007654f
C4485 vdd.n2446 gnd 0.007654f
C4486 vdd.n2447 gnd 0.007654f
C4487 vdd.n2448 gnd 0.007654f
C4488 vdd.n2449 gnd 0.007654f
C4489 vdd.n2450 gnd 0.609628f
C4490 vdd.n2451 gnd 0.007654f
C4491 vdd.n2452 gnd 0.007654f
C4492 vdd.n2453 gnd 0.007654f
C4493 vdd.n2454 gnd 0.007654f
C4494 vdd.n2455 gnd 0.007654f
C4495 vdd.n2456 gnd 0.007654f
C4496 vdd.n2457 gnd 0.488853f
C4497 vdd.n2458 gnd 0.007654f
C4498 vdd.n2459 gnd 0.007654f
C4499 vdd.n2460 gnd 0.007654f
C4500 vdd.n2461 gnd 0.017888f
C4501 vdd.n2462 gnd 0.017229f
C4502 vdd.n2463 gnd 0.007654f
C4503 vdd.n2464 gnd 0.007654f
C4504 vdd.n2465 gnd 0.005909f
C4505 vdd.n2466 gnd 0.007654f
C4506 vdd.n2467 gnd 0.007654f
C4507 vdd.n2468 gnd 0.005571f
C4508 vdd.n2469 gnd 0.007654f
C4509 vdd.n2470 gnd 0.007654f
C4510 vdd.n2471 gnd 0.007654f
C4511 vdd.n2472 gnd 0.007654f
C4512 vdd.n2473 gnd 0.007654f
C4513 vdd.n2474 gnd 0.007654f
C4514 vdd.n2475 gnd 0.007654f
C4515 vdd.n2476 gnd 0.007654f
C4516 vdd.n2477 gnd 0.007654f
C4517 vdd.n2478 gnd 0.007654f
C4518 vdd.n2479 gnd 0.007654f
C4519 vdd.n2480 gnd 0.007654f
C4520 vdd.n2481 gnd 0.007654f
C4521 vdd.n2482 gnd 0.007654f
C4522 vdd.n2483 gnd 0.007654f
C4523 vdd.n2484 gnd 0.007654f
C4524 vdd.n2485 gnd 0.007654f
C4525 vdd.n2486 gnd 0.007654f
C4526 vdd.n2487 gnd 0.007654f
C4527 vdd.n2488 gnd 0.007654f
C4528 vdd.n2489 gnd 0.007654f
C4529 vdd.n2490 gnd 0.007654f
C4530 vdd.n2491 gnd 0.007654f
C4531 vdd.n2492 gnd 0.007654f
C4532 vdd.n2493 gnd 0.007654f
C4533 vdd.n2494 gnd 0.007654f
C4534 vdd.n2495 gnd 0.007654f
C4535 vdd.n2496 gnd 0.007654f
C4536 vdd.n2497 gnd 0.007654f
C4537 vdd.n2498 gnd 0.007654f
C4538 vdd.n2499 gnd 0.007654f
C4539 vdd.n2500 gnd 0.007654f
C4540 vdd.n2501 gnd 0.007654f
C4541 vdd.n2502 gnd 0.007654f
C4542 vdd.n2503 gnd 0.007654f
C4543 vdd.n2504 gnd 0.007654f
C4544 vdd.n2505 gnd 0.007654f
C4545 vdd.n2506 gnd 0.007654f
C4546 vdd.n2507 gnd 0.007654f
C4547 vdd.n2508 gnd 0.007654f
C4548 vdd.n2509 gnd 0.007654f
C4549 vdd.n2510 gnd 0.007654f
C4550 vdd.n2511 gnd 0.007654f
C4551 vdd.n2512 gnd 0.007654f
C4552 vdd.n2513 gnd 0.007654f
C4553 vdd.n2514 gnd 0.007654f
C4554 vdd.n2515 gnd 0.007654f
C4555 vdd.n2516 gnd 0.007654f
C4556 vdd.n2517 gnd 0.007654f
C4557 vdd.n2518 gnd 0.007654f
C4558 vdd.n2519 gnd 0.007654f
C4559 vdd.n2520 gnd 0.007654f
C4560 vdd.n2521 gnd 0.007654f
C4561 vdd.n2522 gnd 0.007654f
C4562 vdd.n2523 gnd 0.007654f
C4563 vdd.n2524 gnd 0.007654f
C4564 vdd.n2525 gnd 0.007654f
C4565 vdd.n2526 gnd 0.007654f
C4566 vdd.n2527 gnd 0.007654f
C4567 vdd.n2528 gnd 0.007654f
C4568 vdd.n2529 gnd 0.018161f
C4569 vdd.n2530 gnd 0.016956f
C4570 vdd.n2531 gnd 0.016956f
C4571 vdd.n2532 gnd 0.954701f
C4572 vdd.n2533 gnd 0.016956f
C4573 vdd.n2534 gnd 0.018161f
C4574 vdd.n2535 gnd 0.017229f
C4575 vdd.n2536 gnd 0.007654f
C4576 vdd.n2537 gnd 0.007654f
C4577 vdd.n2538 gnd 0.007654f
C4578 vdd.n2539 gnd 0.005909f
C4579 vdd.n2540 gnd 0.010938f
C4580 vdd.n2541 gnd 0.005571f
C4581 vdd.n2542 gnd 0.007654f
C4582 vdd.n2543 gnd 0.007654f
C4583 vdd.n2544 gnd 0.007654f
C4584 vdd.n2545 gnd 0.007654f
C4585 vdd.n2546 gnd 0.007654f
C4586 vdd.n2547 gnd 0.007654f
C4587 vdd.n2548 gnd 0.007654f
C4588 vdd.n2549 gnd 0.007654f
C4589 vdd.n2550 gnd 0.007654f
C4590 vdd.n2551 gnd 0.007654f
C4591 vdd.n2552 gnd 0.007654f
C4592 vdd.n2553 gnd 0.007654f
C4593 vdd.n2554 gnd 0.007654f
C4594 vdd.n2555 gnd 0.007654f
C4595 vdd.n2556 gnd 0.007654f
C4596 vdd.n2557 gnd 0.007654f
C4597 vdd.n2558 gnd 0.007654f
C4598 vdd.n2559 gnd 0.007654f
C4599 vdd.n2560 gnd 0.007654f
C4600 vdd.n2561 gnd 0.007654f
C4601 vdd.n2562 gnd 0.007654f
C4602 vdd.n2563 gnd 0.007654f
C4603 vdd.n2564 gnd 0.007654f
C4604 vdd.n2565 gnd 0.007654f
C4605 vdd.n2566 gnd 0.007654f
C4606 vdd.n2567 gnd 0.007654f
C4607 vdd.n2568 gnd 0.007654f
C4608 vdd.n2569 gnd 0.007654f
C4609 vdd.n2570 gnd 0.007654f
C4610 vdd.n2571 gnd 0.007654f
C4611 vdd.n2572 gnd 0.007654f
C4612 vdd.n2573 gnd 0.007654f
C4613 vdd.n2574 gnd 0.007654f
C4614 vdd.n2575 gnd 0.007654f
C4615 vdd.n2576 gnd 0.007654f
C4616 vdd.n2577 gnd 0.007654f
C4617 vdd.n2578 gnd 0.007654f
C4618 vdd.n2579 gnd 0.007654f
C4619 vdd.n2580 gnd 0.007654f
C4620 vdd.n2581 gnd 0.007654f
C4621 vdd.n2582 gnd 0.007654f
C4622 vdd.n2583 gnd 0.007654f
C4623 vdd.n2584 gnd 0.007654f
C4624 vdd.n2585 gnd 0.007654f
C4625 vdd.n2586 gnd 0.007654f
C4626 vdd.n2587 gnd 0.007654f
C4627 vdd.n2588 gnd 0.007654f
C4628 vdd.n2589 gnd 0.007654f
C4629 vdd.n2590 gnd 0.007654f
C4630 vdd.n2591 gnd 0.007654f
C4631 vdd.n2592 gnd 0.007654f
C4632 vdd.n2593 gnd 0.007654f
C4633 vdd.n2594 gnd 0.007654f
C4634 vdd.n2595 gnd 0.007654f
C4635 vdd.n2596 gnd 0.007654f
C4636 vdd.n2597 gnd 0.007654f
C4637 vdd.n2598 gnd 0.007654f
C4638 vdd.n2599 gnd 0.007654f
C4639 vdd.n2600 gnd 0.007654f
C4640 vdd.n2601 gnd 0.007654f
C4641 vdd.n2602 gnd 0.018161f
C4642 vdd.n2603 gnd 0.018161f
C4643 vdd.n2604 gnd 0.954701f
C4644 vdd.t26 gnd 3.39321f
C4645 vdd.t48 gnd 3.39321f
C4646 vdd.n2637 gnd 0.018161f
C4647 vdd.n2638 gnd 0.007654f
C4648 vdd.t103 gnd 0.309282f
C4649 vdd.t104 gnd 0.316589f
C4650 vdd.t101 gnd 0.201911f
C4651 vdd.n2639 gnd 0.109122f
C4652 vdd.n2640 gnd 0.061898f
C4653 vdd.n2641 gnd 0.007654f
C4654 vdd.t116 gnd 0.309282f
C4655 vdd.t117 gnd 0.316589f
C4656 vdd.t115 gnd 0.201911f
C4657 vdd.n2642 gnd 0.109122f
C4658 vdd.n2643 gnd 0.061898f
C4659 vdd.n2644 gnd 0.010938f
C4660 vdd.n2645 gnd 0.007654f
C4661 vdd.n2646 gnd 0.007654f
C4662 vdd.n2647 gnd 0.007654f
C4663 vdd.n2648 gnd 0.007654f
C4664 vdd.n2649 gnd 0.007654f
C4665 vdd.n2650 gnd 0.007654f
C4666 vdd.n2651 gnd 0.007654f
C4667 vdd.n2652 gnd 0.007654f
C4668 vdd.n2653 gnd 0.007654f
C4669 vdd.n2654 gnd 0.007654f
C4670 vdd.n2655 gnd 0.007654f
C4671 vdd.n2656 gnd 0.007654f
C4672 vdd.n2657 gnd 0.007654f
C4673 vdd.n2658 gnd 0.007654f
C4674 vdd.n2659 gnd 0.007654f
C4675 vdd.n2660 gnd 0.007654f
C4676 vdd.n2661 gnd 0.007654f
C4677 vdd.n2662 gnd 0.007654f
C4678 vdd.n2663 gnd 0.007654f
C4679 vdd.n2664 gnd 0.007654f
C4680 vdd.n2665 gnd 0.007654f
C4681 vdd.n2666 gnd 0.007654f
C4682 vdd.n2667 gnd 0.007654f
C4683 vdd.n2668 gnd 0.007654f
C4684 vdd.n2669 gnd 0.007654f
C4685 vdd.n2670 gnd 0.007654f
C4686 vdd.n2671 gnd 0.007654f
C4687 vdd.n2672 gnd 0.007654f
C4688 vdd.n2673 gnd 0.007654f
C4689 vdd.n2674 gnd 0.007654f
C4690 vdd.n2675 gnd 0.007654f
C4691 vdd.n2676 gnd 0.007654f
C4692 vdd.n2677 gnd 0.007654f
C4693 vdd.n2678 gnd 0.007654f
C4694 vdd.n2679 gnd 0.007654f
C4695 vdd.n2680 gnd 0.007654f
C4696 vdd.n2681 gnd 0.007654f
C4697 vdd.n2682 gnd 0.007654f
C4698 vdd.n2683 gnd 0.007654f
C4699 vdd.n2684 gnd 0.007654f
C4700 vdd.n2685 gnd 0.007654f
C4701 vdd.n2686 gnd 0.007654f
C4702 vdd.n2687 gnd 0.007654f
C4703 vdd.n2688 gnd 0.007654f
C4704 vdd.n2689 gnd 0.007654f
C4705 vdd.n2690 gnd 0.007654f
C4706 vdd.n2691 gnd 0.007654f
C4707 vdd.n2692 gnd 0.007654f
C4708 vdd.n2693 gnd 0.007654f
C4709 vdd.n2694 gnd 0.007654f
C4710 vdd.n2695 gnd 0.007654f
C4711 vdd.n2696 gnd 0.007654f
C4712 vdd.n2697 gnd 0.007654f
C4713 vdd.n2698 gnd 0.007654f
C4714 vdd.n2699 gnd 0.007654f
C4715 vdd.n2700 gnd 0.007654f
C4716 vdd.n2701 gnd 0.005571f
C4717 vdd.n2702 gnd 0.007654f
C4718 vdd.n2703 gnd 0.007654f
C4719 vdd.n2704 gnd 0.005909f
C4720 vdd.n2705 gnd 0.007654f
C4721 vdd.n2706 gnd 0.007654f
C4722 vdd.n2707 gnd 0.018161f
C4723 vdd.n2708 gnd 0.016956f
C4724 vdd.n2709 gnd 0.007654f
C4725 vdd.n2710 gnd 0.007654f
C4726 vdd.n2711 gnd 0.007654f
C4727 vdd.n2712 gnd 0.007654f
C4728 vdd.n2713 gnd 0.007654f
C4729 vdd.n2714 gnd 0.007654f
C4730 vdd.n2715 gnd 0.007654f
C4731 vdd.n2716 gnd 0.007654f
C4732 vdd.n2717 gnd 0.007654f
C4733 vdd.n2718 gnd 0.007654f
C4734 vdd.n2719 gnd 0.007654f
C4735 vdd.n2720 gnd 0.007654f
C4736 vdd.n2721 gnd 0.007654f
C4737 vdd.n2722 gnd 0.007654f
C4738 vdd.n2723 gnd 0.007654f
C4739 vdd.n2724 gnd 0.007654f
C4740 vdd.n2725 gnd 0.007654f
C4741 vdd.n2726 gnd 0.007654f
C4742 vdd.n2727 gnd 0.007654f
C4743 vdd.n2728 gnd 0.007654f
C4744 vdd.n2729 gnd 0.007654f
C4745 vdd.n2730 gnd 0.007654f
C4746 vdd.n2731 gnd 0.007654f
C4747 vdd.n2732 gnd 0.007654f
C4748 vdd.n2733 gnd 0.007654f
C4749 vdd.n2734 gnd 0.007654f
C4750 vdd.n2735 gnd 0.007654f
C4751 vdd.n2736 gnd 0.007654f
C4752 vdd.n2737 gnd 0.007654f
C4753 vdd.n2738 gnd 0.007654f
C4754 vdd.n2739 gnd 0.007654f
C4755 vdd.n2740 gnd 0.007654f
C4756 vdd.n2741 gnd 0.007654f
C4757 vdd.n2742 gnd 0.007654f
C4758 vdd.n2743 gnd 0.007654f
C4759 vdd.n2744 gnd 0.007654f
C4760 vdd.n2745 gnd 0.007654f
C4761 vdd.n2746 gnd 0.007654f
C4762 vdd.n2747 gnd 0.007654f
C4763 vdd.n2748 gnd 0.007654f
C4764 vdd.n2749 gnd 0.007654f
C4765 vdd.n2750 gnd 0.007654f
C4766 vdd.n2751 gnd 0.007654f
C4767 vdd.n2752 gnd 0.007654f
C4768 vdd.n2753 gnd 0.007654f
C4769 vdd.n2754 gnd 0.007654f
C4770 vdd.n2755 gnd 0.007654f
C4771 vdd.n2756 gnd 0.007654f
C4772 vdd.n2757 gnd 0.007654f
C4773 vdd.n2758 gnd 0.007654f
C4774 vdd.n2759 gnd 0.007654f
C4775 vdd.n2760 gnd 0.247302f
C4776 vdd.n2761 gnd 0.007654f
C4777 vdd.n2762 gnd 0.007654f
C4778 vdd.n2763 gnd 0.007654f
C4779 vdd.n2764 gnd 0.007654f
C4780 vdd.n2765 gnd 0.007654f
C4781 vdd.n2766 gnd 0.007654f
C4782 vdd.n2767 gnd 0.007654f
C4783 vdd.n2768 gnd 0.007654f
C4784 vdd.n2769 gnd 0.007654f
C4785 vdd.n2770 gnd 0.007654f
C4786 vdd.n2771 gnd 0.007654f
C4787 vdd.n2772 gnd 0.007654f
C4788 vdd.n2773 gnd 0.007654f
C4789 vdd.n2774 gnd 0.007654f
C4790 vdd.n2775 gnd 0.007654f
C4791 vdd.n2776 gnd 0.007654f
C4792 vdd.n2777 gnd 0.007654f
C4793 vdd.n2778 gnd 0.007654f
C4794 vdd.n2779 gnd 0.007654f
C4795 vdd.n2780 gnd 0.007654f
C4796 vdd.n2781 gnd 0.465848f
C4797 vdd.n2782 gnd 0.007654f
C4798 vdd.n2783 gnd 0.007654f
C4799 vdd.n2784 gnd 0.007654f
C4800 vdd.n2785 gnd 0.007654f
C4801 vdd.n2786 gnd 0.007654f
C4802 vdd.n2787 gnd 0.016956f
C4803 vdd.n2788 gnd 0.018161f
C4804 vdd.n2789 gnd 0.018161f
C4805 vdd.n2790 gnd 0.007654f
C4806 vdd.n2791 gnd 0.007654f
C4807 vdd.n2792 gnd 0.007654f
C4808 vdd.n2793 gnd 0.005909f
C4809 vdd.n2794 gnd 0.010938f
C4810 vdd.n2795 gnd 0.005571f
C4811 vdd.n2796 gnd 0.007654f
C4812 vdd.n2797 gnd 0.007654f
C4813 vdd.n2798 gnd 0.007654f
C4814 vdd.n2799 gnd 0.007654f
C4815 vdd.n2800 gnd 0.007654f
C4816 vdd.n2801 gnd 0.007654f
C4817 vdd.n2802 gnd 0.007654f
C4818 vdd.n2803 gnd 0.007654f
C4819 vdd.n2804 gnd 0.007654f
C4820 vdd.n2805 gnd 0.007654f
C4821 vdd.n2806 gnd 0.007654f
C4822 vdd.n2807 gnd 0.007654f
C4823 vdd.n2808 gnd 0.007654f
C4824 vdd.n2809 gnd 0.007654f
C4825 vdd.n2810 gnd 0.007654f
C4826 vdd.n2811 gnd 0.007654f
C4827 vdd.n2812 gnd 0.007654f
C4828 vdd.n2813 gnd 0.007654f
C4829 vdd.n2814 gnd 0.007654f
C4830 vdd.n2815 gnd 0.007654f
C4831 vdd.n2816 gnd 0.007654f
C4832 vdd.n2817 gnd 0.007654f
C4833 vdd.n2818 gnd 0.007654f
C4834 vdd.n2819 gnd 0.007654f
C4835 vdd.n2820 gnd 0.007654f
C4836 vdd.n2821 gnd 0.007654f
C4837 vdd.n2822 gnd 0.007654f
C4838 vdd.n2823 gnd 0.007654f
C4839 vdd.n2824 gnd 0.007654f
C4840 vdd.n2825 gnd 0.007654f
C4841 vdd.n2826 gnd 0.007654f
C4842 vdd.n2827 gnd 0.007654f
C4843 vdd.n2828 gnd 0.007654f
C4844 vdd.n2829 gnd 0.007654f
C4845 vdd.n2830 gnd 0.007654f
C4846 vdd.n2831 gnd 0.007654f
C4847 vdd.n2832 gnd 0.007654f
C4848 vdd.n2833 gnd 0.007654f
C4849 vdd.n2834 gnd 0.007654f
C4850 vdd.n2835 gnd 0.007654f
C4851 vdd.n2836 gnd 0.007654f
C4852 vdd.n2837 gnd 0.007654f
C4853 vdd.n2838 gnd 0.007654f
C4854 vdd.n2839 gnd 0.007654f
C4855 vdd.n2840 gnd 0.007654f
C4856 vdd.n2841 gnd 0.007654f
C4857 vdd.n2842 gnd 0.007654f
C4858 vdd.n2843 gnd 0.007654f
C4859 vdd.n2844 gnd 0.007654f
C4860 vdd.n2845 gnd 0.007654f
C4861 vdd.n2846 gnd 0.007654f
C4862 vdd.n2847 gnd 0.007654f
C4863 vdd.n2848 gnd 0.007654f
C4864 vdd.n2849 gnd 0.007654f
C4865 vdd.n2850 gnd 0.007654f
C4866 vdd.n2851 gnd 0.007654f
C4867 vdd.n2852 gnd 0.007654f
C4868 vdd.n2853 gnd 0.007654f
C4869 vdd.n2854 gnd 0.007654f
C4870 vdd.n2855 gnd 0.007654f
C4871 vdd.n2857 gnd 0.954701f
C4872 vdd.n2859 gnd 0.007654f
C4873 vdd.n2860 gnd 0.007654f
C4874 vdd.n2861 gnd 0.018161f
C4875 vdd.n2862 gnd 0.016956f
C4876 vdd.n2863 gnd 0.016956f
C4877 vdd.n2864 gnd 0.954701f
C4878 vdd.n2865 gnd 0.016956f
C4879 vdd.n2866 gnd 0.016956f
C4880 vdd.n2867 gnd 0.007654f
C4881 vdd.n2868 gnd 0.007654f
C4882 vdd.n2869 gnd 0.007654f
C4883 vdd.n2870 gnd 0.488853f
C4884 vdd.n2871 gnd 0.007654f
C4885 vdd.n2872 gnd 0.007654f
C4886 vdd.n2873 gnd 0.007654f
C4887 vdd.n2874 gnd 0.007654f
C4888 vdd.n2875 gnd 0.007654f
C4889 vdd.n2876 gnd 0.609628f
C4890 vdd.n2877 gnd 0.007654f
C4891 vdd.n2878 gnd 0.007654f
C4892 vdd.n2879 gnd 0.007654f
C4893 vdd.n2880 gnd 0.007654f
C4894 vdd.n2881 gnd 0.007654f
C4895 vdd.n2882 gnd 0.782164f
C4896 vdd.n2883 gnd 0.007654f
C4897 vdd.n2884 gnd 0.007654f
C4898 vdd.n2885 gnd 0.007654f
C4899 vdd.n2886 gnd 0.007654f
C4900 vdd.n2887 gnd 0.007654f
C4901 vdd.n2888 gnd 0.431341f
C4902 vdd.n2889 gnd 0.007654f
C4903 vdd.n2890 gnd 0.007654f
C4904 vdd.n2891 gnd 0.007654f
C4905 vdd.n2892 gnd 0.007654f
C4906 vdd.n2893 gnd 0.007654f
C4907 vdd.n2894 gnd 0.247302f
C4908 vdd.n2895 gnd 0.007654f
C4909 vdd.n2896 gnd 0.007654f
C4910 vdd.n2897 gnd 0.007654f
C4911 vdd.n2898 gnd 0.007654f
C4912 vdd.n2899 gnd 0.007654f
C4913 vdd.n2900 gnd 0.448594f
C4914 vdd.n2901 gnd 0.007654f
C4915 vdd.n2902 gnd 0.007654f
C4916 vdd.n2903 gnd 0.007654f
C4917 vdd.n2904 gnd 0.007654f
C4918 vdd.n2905 gnd 0.007654f
C4919 vdd.n2906 gnd 0.621131f
C4920 vdd.n2907 gnd 0.007654f
C4921 vdd.n2908 gnd 0.007654f
C4922 vdd.n2909 gnd 0.007654f
C4923 vdd.n2910 gnd 0.007654f
C4924 vdd.n2911 gnd 0.007654f
C4925 vdd.n2912 gnd 0.695896f
C4926 vdd.n2913 gnd 0.007654f
C4927 vdd.n2914 gnd 0.007654f
C4928 vdd.n2915 gnd 0.007654f
C4929 vdd.n2916 gnd 0.007654f
C4930 vdd.n2917 gnd 0.007654f
C4931 vdd.n2918 gnd 0.52336f
C4932 vdd.n2919 gnd 0.007654f
C4933 vdd.n2920 gnd 0.007654f
C4934 vdd.n2921 gnd 0.007654f
C4935 vdd.t71 gnd 0.316589f
C4936 vdd.t69 gnd 0.201911f
C4937 vdd.t72 gnd 0.316589f
C4938 vdd.n2922 gnd 0.177936f
C4939 vdd.n2923 gnd 0.022172f
C4940 vdd.n2924 gnd 0.004727f
C4941 vdd.n2925 gnd 0.007654f
C4942 vdd.n2926 gnd 0.431341f
C4943 vdd.n2927 gnd 0.007654f
C4944 vdd.n2928 gnd 0.007654f
C4945 vdd.n2929 gnd 0.007654f
C4946 vdd.n2930 gnd 0.007654f
C4947 vdd.n2931 gnd 0.007654f
C4948 vdd.n2932 gnd 0.782164f
C4949 vdd.n2933 gnd 0.007654f
C4950 vdd.n2934 gnd 0.007654f
C4951 vdd.n2935 gnd 0.007654f
C4952 vdd.n2936 gnd 0.007654f
C4953 vdd.n2937 gnd 0.007654f
C4954 vdd.n2938 gnd 0.007654f
C4955 vdd.n2940 gnd 0.007654f
C4956 vdd.n2941 gnd 0.007654f
C4957 vdd.n2943 gnd 0.007654f
C4958 vdd.n2944 gnd 0.007654f
C4959 vdd.n2947 gnd 0.007654f
C4960 vdd.n2948 gnd 0.007654f
C4961 vdd.n2949 gnd 0.007654f
C4962 vdd.n2950 gnd 0.007654f
C4963 vdd.n2952 gnd 0.007654f
C4964 vdd.n2953 gnd 0.007654f
C4965 vdd.n2954 gnd 0.007654f
C4966 vdd.n2955 gnd 0.007654f
C4967 vdd.n2956 gnd 0.007654f
C4968 vdd.n2957 gnd 0.007654f
C4969 vdd.n2959 gnd 0.007654f
C4970 vdd.n2960 gnd 0.007654f
C4971 vdd.n2961 gnd 0.007654f
C4972 vdd.n2962 gnd 0.007654f
C4973 vdd.n2963 gnd 0.007654f
C4974 vdd.n2964 gnd 0.007654f
C4975 vdd.n2966 gnd 0.007654f
C4976 vdd.n2967 gnd 0.007654f
C4977 vdd.n2968 gnd 0.007654f
C4978 vdd.n2969 gnd 0.007654f
C4979 vdd.n2970 gnd 0.007654f
C4980 vdd.n2971 gnd 0.007654f
C4981 vdd.n2973 gnd 0.007654f
C4982 vdd.n2974 gnd 0.018161f
C4983 vdd.n2975 gnd 0.018161f
C4984 vdd.n2976 gnd 0.016956f
C4985 vdd.n2977 gnd 0.007654f
C4986 vdd.n2978 gnd 0.007654f
C4987 vdd.n2979 gnd 0.007654f
C4988 vdd.n2980 gnd 0.007654f
C4989 vdd.n2981 gnd 0.007654f
C4990 vdd.n2982 gnd 0.007654f
C4991 vdd.n2983 gnd 0.782164f
C4992 vdd.n2984 gnd 0.007654f
C4993 vdd.n2985 gnd 0.007654f
C4994 vdd.n2986 gnd 0.007654f
C4995 vdd.n2987 gnd 0.007654f
C4996 vdd.n2988 gnd 0.007654f
C4997 vdd.n2989 gnd 0.488853f
C4998 vdd.n2990 gnd 0.007654f
C4999 vdd.n2991 gnd 0.007654f
C5000 vdd.n2992 gnd 0.007654f
C5001 vdd.n2993 gnd 0.017888f
C5002 vdd.n2994 gnd 0.017229f
C5003 vdd.n2995 gnd 0.018161f
C5004 vdd.n2997 gnd 0.007654f
C5005 vdd.n2998 gnd 0.007654f
C5006 vdd.n2999 gnd 0.005909f
C5007 vdd.n3000 gnd 0.010938f
C5008 vdd.n3001 gnd 0.005571f
C5009 vdd.n3002 gnd 0.007654f
C5010 vdd.n3003 gnd 0.007654f
C5011 vdd.n3005 gnd 0.007654f
C5012 vdd.n3006 gnd 0.007654f
C5013 vdd.n3007 gnd 0.007654f
C5014 vdd.n3008 gnd 0.007654f
C5015 vdd.n3009 gnd 0.007654f
C5016 vdd.n3010 gnd 0.007654f
C5017 vdd.n3012 gnd 0.007654f
C5018 vdd.n3013 gnd 0.007654f
C5019 vdd.n3014 gnd 0.007654f
C5020 vdd.n3015 gnd 0.007654f
C5021 vdd.n3016 gnd 0.007654f
C5022 vdd.n3017 gnd 0.007654f
C5023 vdd.n3019 gnd 0.007654f
C5024 vdd.n3020 gnd 0.007654f
C5025 vdd.n3021 gnd 0.007654f
C5026 vdd.n3022 gnd 0.007654f
C5027 vdd.n3023 gnd 0.007654f
C5028 vdd.n3024 gnd 0.007654f
C5029 vdd.n3026 gnd 0.007654f
C5030 vdd.n3027 gnd 0.007654f
C5031 vdd.n3028 gnd 0.007654f
C5032 vdd.n3030 gnd 0.007654f
C5033 vdd.n3031 gnd 0.007654f
C5034 vdd.n3032 gnd 0.007654f
C5035 vdd.n3033 gnd 0.007654f
C5036 vdd.n3034 gnd 0.007654f
C5037 vdd.n3035 gnd 0.007654f
C5038 vdd.n3037 gnd 0.007654f
C5039 vdd.n3038 gnd 0.007654f
C5040 vdd.n3039 gnd 0.007654f
C5041 vdd.n3040 gnd 0.007654f
C5042 vdd.n3041 gnd 0.007654f
C5043 vdd.n3042 gnd 0.007654f
C5044 vdd.n3044 gnd 0.007654f
C5045 vdd.n3045 gnd 0.007654f
C5046 vdd.n3046 gnd 0.007654f
C5047 vdd.n3047 gnd 0.007654f
C5048 vdd.n3048 gnd 0.007654f
C5049 vdd.n3049 gnd 0.007654f
C5050 vdd.n3051 gnd 0.007654f
C5051 vdd.n3052 gnd 0.007654f
C5052 vdd.n3054 gnd 0.007654f
C5053 vdd.n3055 gnd 0.007654f
C5054 vdd.n3056 gnd 0.018161f
C5055 vdd.n3057 gnd 0.016956f
C5056 vdd.n3058 gnd 0.016956f
C5057 vdd.n3059 gnd 1.12724f
C5058 vdd.n3060 gnd 0.016956f
C5059 vdd.n3061 gnd 0.018161f
C5060 vdd.n3062 gnd 0.017229f
C5061 vdd.n3063 gnd 0.007654f
C5062 vdd.n3064 gnd 0.005909f
C5063 vdd.n3065 gnd 0.007654f
C5064 vdd.n3067 gnd 0.007654f
C5065 vdd.n3068 gnd 0.007654f
C5066 vdd.n3069 gnd 0.007654f
C5067 vdd.n3070 gnd 0.007654f
C5068 vdd.n3071 gnd 0.007654f
C5069 vdd.n3072 gnd 0.007654f
C5070 vdd.n3074 gnd 0.007654f
C5071 vdd.n3075 gnd 0.007654f
C5072 vdd.n3076 gnd 0.007654f
C5073 vdd.n3077 gnd 0.007654f
C5074 vdd.n3078 gnd 0.007654f
C5075 vdd.n3079 gnd 0.007654f
C5076 vdd.n3081 gnd 0.007654f
C5077 vdd.n3082 gnd 0.007654f
C5078 vdd.n3083 gnd 0.007654f
C5079 vdd.n3084 gnd 0.007654f
C5080 vdd.n3085 gnd 0.007654f
C5081 vdd.n3086 gnd 0.007654f
C5082 vdd.n3088 gnd 0.007654f
C5083 vdd.n3089 gnd 0.007654f
C5084 vdd.n3091 gnd 0.007654f
C5085 vdd.n3092 gnd 0.018392f
C5086 vdd.n3093 gnd 0.681191f
C5087 vdd.n3095 gnd 0.004756f
C5088 vdd.n3096 gnd 0.009059f
C5089 vdd.n3097 gnd 0.011255f
C5090 vdd.n3098 gnd 0.011255f
C5091 vdd.n3099 gnd 0.009059f
C5092 vdd.n3100 gnd 0.009059f
C5093 vdd.n3101 gnd 0.011255f
C5094 vdd.n3102 gnd 0.011255f
C5095 vdd.n3103 gnd 0.009059f
C5096 vdd.n3104 gnd 0.009059f
C5097 vdd.n3105 gnd 0.011255f
C5098 vdd.n3106 gnd 0.011255f
C5099 vdd.n3107 gnd 0.009059f
C5100 vdd.n3108 gnd 0.009059f
C5101 vdd.n3109 gnd 0.011255f
C5102 vdd.n3110 gnd 0.011255f
C5103 vdd.n3111 gnd 0.009059f
C5104 vdd.n3112 gnd 0.009059f
C5105 vdd.n3113 gnd 0.011255f
C5106 vdd.n3114 gnd 0.011255f
C5107 vdd.n3115 gnd 0.009059f
C5108 vdd.n3116 gnd 0.009059f
C5109 vdd.n3117 gnd 0.011255f
C5110 vdd.n3118 gnd 0.011255f
C5111 vdd.n3119 gnd 0.009059f
C5112 vdd.n3120 gnd 0.009059f
C5113 vdd.n3121 gnd 0.011255f
C5114 vdd.n3122 gnd 0.011255f
C5115 vdd.n3123 gnd 0.009059f
C5116 vdd.n3124 gnd 0.009059f
C5117 vdd.n3125 gnd 0.011255f
C5118 vdd.n3126 gnd 0.011255f
C5119 vdd.n3127 gnd 0.009059f
C5120 vdd.n3128 gnd 0.009059f
C5121 vdd.n3129 gnd 0.011255f
C5122 vdd.n3130 gnd 0.011255f
C5123 vdd.n3131 gnd 0.009059f
C5124 vdd.n3132 gnd 0.011255f
C5125 vdd.n3133 gnd 0.011255f
C5126 vdd.n3134 gnd 0.009059f
C5127 vdd.n3135 gnd 0.011255f
C5128 vdd.n3136 gnd 0.011255f
C5129 vdd.n3137 gnd 0.011255f
C5130 vdd.n3138 gnd 0.018481f
C5131 vdd.n3139 gnd 0.011255f
C5132 vdd.n3140 gnd 0.011255f
C5133 vdd.n3141 gnd 0.00616f
C5134 vdd.n3142 gnd 0.009059f
C5135 vdd.n3143 gnd 0.011255f
C5136 vdd.n3144 gnd 0.011255f
C5137 vdd.n3145 gnd 0.009059f
C5138 vdd.n3146 gnd 0.009059f
C5139 vdd.n3147 gnd 0.011255f
C5140 vdd.n3148 gnd 0.011255f
C5141 vdd.n3149 gnd 0.009059f
C5142 vdd.n3150 gnd 0.009059f
C5143 vdd.n3151 gnd 0.011255f
C5144 vdd.n3152 gnd 0.011255f
C5145 vdd.n3153 gnd 0.009059f
C5146 vdd.n3154 gnd 0.009059f
C5147 vdd.n3155 gnd 0.011255f
C5148 vdd.n3156 gnd 0.011255f
C5149 vdd.n3157 gnd 0.009059f
C5150 vdd.n3158 gnd 0.009059f
C5151 vdd.n3159 gnd 0.011255f
C5152 vdd.n3160 gnd 0.011255f
C5153 vdd.n3161 gnd 0.009059f
C5154 vdd.n3162 gnd 0.009059f
C5155 vdd.n3163 gnd 0.011255f
C5156 vdd.n3164 gnd 0.011255f
C5157 vdd.n3165 gnd 0.009059f
C5158 vdd.n3166 gnd 0.009059f
C5159 vdd.n3167 gnd 0.011255f
C5160 vdd.n3168 gnd 0.011255f
C5161 vdd.n3169 gnd 0.009059f
C5162 vdd.n3170 gnd 0.009059f
C5163 vdd.n3171 gnd 0.011255f
C5164 vdd.n3172 gnd 0.011255f
C5165 vdd.n3173 gnd 0.009059f
C5166 vdd.n3174 gnd 0.009059f
C5167 vdd.n3175 gnd 0.011255f
C5168 vdd.n3176 gnd 0.011255f
C5169 vdd.n3177 gnd 0.009059f
C5170 vdd.n3178 gnd 0.011255f
C5171 vdd.n3179 gnd 0.011255f
C5172 vdd.n3180 gnd 0.009059f
C5173 vdd.n3181 gnd 0.011255f
C5174 vdd.n3182 gnd 0.011255f
C5175 vdd.n3183 gnd 0.011255f
C5176 vdd.t63 gnd 0.13847f
C5177 vdd.t64 gnd 0.147986f
C5178 vdd.t62 gnd 0.18084f
C5179 vdd.n3184 gnd 0.231812f
C5180 vdd.n3185 gnd 0.194764f
C5181 vdd.n3186 gnd 0.018481f
C5182 vdd.n3187 gnd 0.011255f
C5183 vdd.n3188 gnd 0.011255f
C5184 vdd.n3189 gnd 0.007564f
C5185 vdd.n3190 gnd 0.009059f
C5186 vdd.n3191 gnd 0.011255f
C5187 vdd.n3192 gnd 0.011255f
C5188 vdd.n3193 gnd 0.009059f
C5189 vdd.n3194 gnd 0.009059f
C5190 vdd.n3195 gnd 0.011255f
C5191 vdd.n3196 gnd 0.011255f
C5192 vdd.n3197 gnd 0.009059f
C5193 vdd.n3198 gnd 0.009059f
C5194 vdd.n3199 gnd 0.011255f
C5195 vdd.n3200 gnd 0.011255f
C5196 vdd.n3201 gnd 0.009059f
C5197 vdd.n3202 gnd 0.009059f
C5198 vdd.n3203 gnd 0.011255f
C5199 vdd.n3204 gnd 0.011255f
C5200 vdd.n3205 gnd 0.009059f
C5201 vdd.n3206 gnd 0.009059f
C5202 vdd.n3207 gnd 0.011255f
C5203 vdd.n3208 gnd 0.011255f
C5204 vdd.n3209 gnd 0.009059f
C5205 vdd.n3210 gnd 0.009059f
C5206 vdd.n3211 gnd 0.011255f
C5207 vdd.n3212 gnd 0.011255f
C5208 vdd.n3213 gnd 0.009059f
C5209 vdd.n3214 gnd 0.009059f
C5210 vdd.n3216 gnd 0.681191f
C5211 vdd.n3218 gnd 0.009059f
C5212 vdd.n3219 gnd 0.009059f
C5213 vdd.n3220 gnd 0.007519f
C5214 vdd.n3221 gnd 0.027811f
C5215 vdd.n3223 gnd 8.31625f
C5216 vdd.n3224 gnd 0.027811f
C5217 vdd.n3225 gnd 0.004303f
C5218 vdd.n3226 gnd 0.027811f
C5219 vdd.n3227 gnd 0.027228f
C5220 vdd.n3228 gnd 0.011255f
C5221 vdd.n3229 gnd 0.009059f
C5222 vdd.n3230 gnd 0.011255f
C5223 vdd.n3231 gnd 0.695896f
C5224 vdd.n3232 gnd 0.011255f
C5225 vdd.n3233 gnd 0.009059f
C5226 vdd.n3234 gnd 0.011255f
C5227 vdd.n3235 gnd 0.011255f
C5228 vdd.n3236 gnd 0.011255f
C5229 vdd.n3237 gnd 0.009059f
C5230 vdd.n3238 gnd 0.011255f
C5231 vdd.n3239 gnd 1.15024f
C5232 vdd.n3240 gnd 0.011255f
C5233 vdd.n3241 gnd 0.009059f
C5234 vdd.n3242 gnd 0.011255f
C5235 vdd.n3243 gnd 0.011255f
C5236 vdd.n3244 gnd 0.011255f
C5237 vdd.n3245 gnd 0.009059f
C5238 vdd.n3246 gnd 0.011255f
C5239 vdd.n3247 gnd 0.741906f
C5240 vdd.n3248 gnd 0.787916f
C5241 vdd.n3249 gnd 0.011255f
C5242 vdd.n3250 gnd 0.009059f
C5243 vdd.n3251 gnd 0.011255f
C5244 vdd.n3252 gnd 0.011255f
C5245 vdd.n3253 gnd 0.011255f
C5246 vdd.n3254 gnd 0.009059f
C5247 vdd.n3255 gnd 0.011255f
C5248 vdd.n3256 gnd 0.954701f
C5249 vdd.n3257 gnd 0.011255f
C5250 vdd.n3258 gnd 0.009059f
C5251 vdd.n3259 gnd 0.011255f
C5252 vdd.n3260 gnd 0.011255f
C5253 vdd.n3261 gnd 0.011255f
C5254 vdd.n3262 gnd 0.009059f
C5255 vdd.n3263 gnd 0.011255f
C5256 vdd.t150 gnd 0.575121f
C5257 vdd.n3264 gnd 0.925945f
C5258 vdd.n3265 gnd 0.011255f
C5259 vdd.n3266 gnd 0.009059f
C5260 vdd.n3267 gnd 0.011255f
C5261 vdd.n3268 gnd 0.011255f
C5262 vdd.n3269 gnd 0.011255f
C5263 vdd.n3270 gnd 0.009059f
C5264 vdd.n3271 gnd 0.011255f
C5265 vdd.n3272 gnd 0.730404f
C5266 vdd.n3273 gnd 0.011255f
C5267 vdd.n3274 gnd 0.009059f
C5268 vdd.n3275 gnd 0.011255f
C5269 vdd.n3276 gnd 0.011255f
C5270 vdd.n3277 gnd 0.011255f
C5271 vdd.n3278 gnd 0.009059f
C5272 vdd.n3279 gnd 0.011255f
C5273 vdd.n3280 gnd 0.914442f
C5274 vdd.n3281 gnd 0.615379f
C5275 vdd.n3282 gnd 0.011255f
C5276 vdd.n3283 gnd 0.009059f
C5277 vdd.n3284 gnd 0.011255f
C5278 vdd.n3285 gnd 0.011255f
C5279 vdd.n3286 gnd 0.011255f
C5280 vdd.n3287 gnd 0.009059f
C5281 vdd.n3288 gnd 0.011255f
C5282 vdd.n3289 gnd 0.81092f
C5283 vdd.n3290 gnd 0.011255f
C5284 vdd.n3291 gnd 0.009059f
C5285 vdd.n3292 gnd 0.011255f
C5286 vdd.n3293 gnd 0.011255f
C5287 vdd.n3294 gnd 0.011255f
C5288 vdd.n3295 gnd 0.011255f
C5289 vdd.n3296 gnd 0.011255f
C5290 vdd.n3297 gnd 0.009059f
C5291 vdd.n3298 gnd 0.009059f
C5292 vdd.n3299 gnd 0.011255f
C5293 vdd.t195 gnd 0.575121f
C5294 vdd.n3300 gnd 0.954701f
C5295 vdd.n3301 gnd 0.011255f
C5296 vdd.n3302 gnd 0.009059f
C5297 vdd.n3303 gnd 0.011255f
C5298 vdd.n3304 gnd 0.011255f
C5299 vdd.n3305 gnd 0.011255f
C5300 vdd.n3306 gnd 0.009059f
C5301 vdd.n3307 gnd 0.011255f
C5302 vdd.n3308 gnd 0.90294f
C5303 vdd.n3309 gnd 0.011255f
C5304 vdd.n3310 gnd 0.011255f
C5305 vdd.n3311 gnd 0.009059f
C5306 vdd.n3312 gnd 0.009059f
C5307 vdd.n3313 gnd 0.011255f
C5308 vdd.n3314 gnd 0.011255f
C5309 vdd.n3315 gnd 0.011255f
C5310 vdd.n3316 gnd 0.009059f
C5311 vdd.n3317 gnd 0.011255f
C5312 vdd.n3318 gnd 0.009059f
C5313 vdd.n3319 gnd 0.009059f
C5314 vdd.n3320 gnd 0.011255f
C5315 vdd.n3321 gnd 0.011255f
C5316 vdd.n3322 gnd 0.011255f
C5317 vdd.n3323 gnd 0.009059f
C5318 vdd.n3324 gnd 0.011255f
C5319 vdd.n3325 gnd 0.009059f
C5320 vdd.n3326 gnd 0.009059f
C5321 vdd.n3327 gnd 0.011255f
C5322 vdd.n3328 gnd 0.011255f
C5323 vdd.n3329 gnd 0.011255f
C5324 vdd.n3330 gnd 0.009059f
C5325 vdd.n3331 gnd 0.954701f
C5326 vdd.n3332 gnd 0.011255f
C5327 vdd.n3333 gnd 0.009059f
C5328 vdd.n3334 gnd 0.009059f
C5329 vdd.n3335 gnd 0.011255f
C5330 vdd.n3336 gnd 0.011255f
C5331 vdd.n3337 gnd 0.011255f
C5332 vdd.n3338 gnd 0.009059f
C5333 vdd.n3339 gnd 0.011255f
C5334 vdd.n3340 gnd 0.009059f
C5335 vdd.n3341 gnd 0.009059f
C5336 vdd.n3342 gnd 0.011255f
C5337 vdd.n3343 gnd 0.011255f
C5338 vdd.n3344 gnd 0.011255f
C5339 vdd.n3345 gnd 0.009059f
C5340 vdd.n3346 gnd 0.011255f
C5341 vdd.n3347 gnd 0.009059f
C5342 vdd.n3348 gnd 0.007519f
C5343 vdd.n3349 gnd 0.027228f
C5344 vdd.n3350 gnd 0.027811f
C5345 vdd.n3351 gnd 0.004303f
C5346 vdd.n3352 gnd 0.027811f
C5347 vdd.n3354 gnd 2.72607f
C5348 vdd.n3355 gnd 1.69661f
C5349 vdd.n3356 gnd 0.027228f
C5350 vdd.n3357 gnd 0.007519f
C5351 vdd.n3358 gnd 0.009059f
C5352 vdd.n3359 gnd 0.009059f
C5353 vdd.n3360 gnd 0.011255f
C5354 vdd.n3361 gnd 1.15024f
C5355 vdd.n3362 gnd 1.15024f
C5356 vdd.n3363 gnd 1.05247f
C5357 vdd.n3364 gnd 0.011255f
C5358 vdd.n3365 gnd 0.009059f
C5359 vdd.n3366 gnd 0.009059f
C5360 vdd.n3367 gnd 0.009059f
C5361 vdd.n3368 gnd 0.011255f
C5362 vdd.n3369 gnd 0.85693f
C5363 vdd.t214 gnd 0.575121f
C5364 vdd.n3370 gnd 0.868433f
C5365 vdd.n3371 gnd 0.661389f
C5366 vdd.n3372 gnd 0.011255f
C5367 vdd.n3373 gnd 0.009059f
C5368 vdd.n3374 gnd 0.009059f
C5369 vdd.n3375 gnd 0.009059f
C5370 vdd.n3376 gnd 0.011255f
C5371 vdd.n3377 gnd 0.684394f
C5372 vdd.n3378 gnd 0.845428f
C5373 vdd.t168 gnd 0.575121f
C5374 vdd.n3379 gnd 0.879935f
C5375 vdd.n3380 gnd 0.011255f
C5376 vdd.n3381 gnd 0.009059f
C5377 vdd.n3382 gnd 0.009059f
C5378 vdd.n3383 gnd 0.009059f
C5379 vdd.n3384 gnd 0.011255f
C5380 vdd.n3385 gnd 0.954701f
C5381 vdd.t191 gnd 0.575121f
C5382 vdd.n3386 gnd 0.695896f
C5383 vdd.n3387 gnd 0.833925f
C5384 vdd.n3388 gnd 0.011255f
C5385 vdd.n3389 gnd 0.009059f
C5386 vdd.n3390 gnd 0.009059f
C5387 vdd.n3391 gnd 0.009059f
C5388 vdd.n3392 gnd 0.011255f
C5389 vdd.n3393 gnd 0.638384f
C5390 vdd.t163 gnd 0.575121f
C5391 vdd.n3394 gnd 0.954701f
C5392 vdd.t136 gnd 0.575121f
C5393 vdd.n3395 gnd 0.707399f
C5394 vdd.n3396 gnd 0.011255f
C5395 vdd.n3397 gnd 0.009059f
C5396 vdd.n3398 gnd 0.00865f
C5397 vdd.n3399 gnd 0.663882f
C5398 vdd.n3400 gnd 2.87815f
C5399 a_n7636_8799.t22 gnd 0.112804f
C5400 a_n7636_8799.t12 gnd 0.112804f
C5401 a_n7636_8799.t11 gnd 0.112804f
C5402 a_n7636_8799.n0 gnd 0.998992f
C5403 a_n7636_8799.t17 gnd 0.112804f
C5404 a_n7636_8799.t16 gnd 0.112804f
C5405 a_n7636_8799.n1 gnd 0.996775f
C5406 a_n7636_8799.n2 gnd 0.793979f
C5407 a_n7636_8799.t29 gnd 0.145034f
C5408 a_n7636_8799.t33 gnd 0.145034f
C5409 a_n7636_8799.n3 gnd 1.1439f
C5410 a_n7636_8799.t35 gnd 0.145034f
C5411 a_n7636_8799.t3 gnd 0.145034f
C5412 a_n7636_8799.n4 gnd 1.14202f
C5413 a_n7636_8799.n5 gnd 1.02654f
C5414 a_n7636_8799.t30 gnd 0.145034f
C5415 a_n7636_8799.t32 gnd 0.145034f
C5416 a_n7636_8799.n6 gnd 1.14202f
C5417 a_n7636_8799.n7 gnd 2.99722f
C5418 a_n7636_8799.t0 gnd 0.145034f
C5419 a_n7636_8799.t4 gnd 0.145034f
C5420 a_n7636_8799.n8 gnd 1.1439f
C5421 a_n7636_8799.t31 gnd 0.145034f
C5422 a_n7636_8799.t34 gnd 0.145034f
C5423 a_n7636_8799.n9 gnd 1.14202f
C5424 a_n7636_8799.n10 gnd 1.02653f
C5425 a_n7636_8799.t2 gnd 0.145034f
C5426 a_n7636_8799.t1 gnd 0.145034f
C5427 a_n7636_8799.n11 gnd 1.14202f
C5428 a_n7636_8799.n12 gnd 1.80385f
C5429 a_n7636_8799.n13 gnd 5.71928f
C5430 a_n7636_8799.n14 gnd 0.052275f
C5431 a_n7636_8799.t132 gnd 0.601377f
C5432 a_n7636_8799.n15 gnd 0.268587f
C5433 a_n7636_8799.n16 gnd 0.052275f
C5434 a_n7636_8799.n17 gnd 0.011862f
C5435 a_n7636_8799.t48 gnd 0.601377f
C5436 a_n7636_8799.n18 gnd 0.052275f
C5437 a_n7636_8799.t69 gnd 0.601377f
C5438 a_n7636_8799.n19 gnd 0.265525f
C5439 a_n7636_8799.t92 gnd 0.601377f
C5440 a_n7636_8799.n20 gnd 0.052275f
C5441 a_n7636_8799.t111 gnd 0.601377f
C5442 a_n7636_8799.n21 gnd 0.265847f
C5443 a_n7636_8799.n22 gnd 0.052275f
C5444 a_n7636_8799.n23 gnd 0.011862f
C5445 a_n7636_8799.t71 gnd 0.601377f
C5446 a_n7636_8799.n24 gnd 0.052275f
C5447 a_n7636_8799.t83 gnd 0.601377f
C5448 a_n7636_8799.n25 gnd 0.268587f
C5449 a_n7636_8799.n26 gnd 0.052275f
C5450 a_n7636_8799.n27 gnd 0.011862f
C5451 a_n7636_8799.t116 gnd 0.601377f
C5452 a_n7636_8799.n28 gnd 0.165151f
C5453 a_n7636_8799.t137 gnd 0.601377f
C5454 a_n7636_8799.t135 gnd 0.612759f
C5455 a_n7636_8799.n29 gnd 0.252102f
C5456 a_n7636_8799.n30 gnd 0.26488f
C5457 a_n7636_8799.n31 gnd 0.011862f
C5458 a_n7636_8799.t87 gnd 0.601377f
C5459 a_n7636_8799.n32 gnd 0.268587f
C5460 a_n7636_8799.n33 gnd 0.052275f
C5461 a_n7636_8799.n34 gnd 0.052275f
C5462 a_n7636_8799.n35 gnd 0.052275f
C5463 a_n7636_8799.n36 gnd 0.266492f
C5464 a_n7636_8799.t133 gnd 0.601377f
C5465 a_n7636_8799.n37 gnd 0.265202f
C5466 a_n7636_8799.n38 gnd 0.011862f
C5467 a_n7636_8799.n39 gnd 0.052275f
C5468 a_n7636_8799.n40 gnd 0.052275f
C5469 a_n7636_8799.n41 gnd 0.052275f
C5470 a_n7636_8799.n42 gnd 0.011862f
C5471 a_n7636_8799.t84 gnd 0.601377f
C5472 a_n7636_8799.n43 gnd 0.266169f
C5473 a_n7636_8799.t114 gnd 0.601377f
C5474 a_n7636_8799.n44 gnd 0.265525f
C5475 a_n7636_8799.n45 gnd 0.052275f
C5476 a_n7636_8799.n46 gnd 0.052275f
C5477 a_n7636_8799.n47 gnd 0.052275f
C5478 a_n7636_8799.n48 gnd 0.268587f
C5479 a_n7636_8799.n49 gnd 0.011862f
C5480 a_n7636_8799.t72 gnd 0.601377f
C5481 a_n7636_8799.n50 gnd 0.265847f
C5482 a_n7636_8799.n51 gnd 0.052275f
C5483 a_n7636_8799.n52 gnd 0.052275f
C5484 a_n7636_8799.n53 gnd 0.052275f
C5485 a_n7636_8799.n54 gnd 0.011862f
C5486 a_n7636_8799.t36 gnd 0.601377f
C5487 a_n7636_8799.n55 gnd 0.268587f
C5488 a_n7636_8799.n56 gnd 0.011862f
C5489 a_n7636_8799.n57 gnd 0.052275f
C5490 a_n7636_8799.n58 gnd 0.052275f
C5491 a_n7636_8799.n59 gnd 0.052275f
C5492 a_n7636_8799.n60 gnd 0.266169f
C5493 a_n7636_8799.n61 gnd 0.011862f
C5494 a_n7636_8799.t136 gnd 0.601377f
C5495 a_n7636_8799.n62 gnd 0.268587f
C5496 a_n7636_8799.n63 gnd 0.052275f
C5497 a_n7636_8799.n64 gnd 0.052275f
C5498 a_n7636_8799.n65 gnd 0.052275f
C5499 a_n7636_8799.n66 gnd 0.265202f
C5500 a_n7636_8799.t66 gnd 0.601377f
C5501 a_n7636_8799.n67 gnd 0.266492f
C5502 a_n7636_8799.n68 gnd 0.011862f
C5503 a_n7636_8799.n69 gnd 0.052275f
C5504 a_n7636_8799.n70 gnd 0.052275f
C5505 a_n7636_8799.n71 gnd 0.052275f
C5506 a_n7636_8799.n72 gnd 0.011862f
C5507 a_n7636_8799.t45 gnd 0.601377f
C5508 a_n7636_8799.n73 gnd 0.26488f
C5509 a_n7636_8799.t46 gnd 0.601377f
C5510 a_n7636_8799.n74 gnd 0.263108f
C5511 a_n7636_8799.n75 gnd 0.296385f
C5512 a_n7636_8799.n76 gnd 0.052275f
C5513 a_n7636_8799.t145 gnd 0.601377f
C5514 a_n7636_8799.n77 gnd 0.268587f
C5515 a_n7636_8799.n78 gnd 0.052275f
C5516 a_n7636_8799.n79 gnd 0.011862f
C5517 a_n7636_8799.t63 gnd 0.601377f
C5518 a_n7636_8799.n80 gnd 0.052275f
C5519 a_n7636_8799.t78 gnd 0.601377f
C5520 a_n7636_8799.n81 gnd 0.265525f
C5521 a_n7636_8799.t105 gnd 0.601377f
C5522 a_n7636_8799.n82 gnd 0.052275f
C5523 a_n7636_8799.t123 gnd 0.601377f
C5524 a_n7636_8799.n83 gnd 0.265847f
C5525 a_n7636_8799.n84 gnd 0.052275f
C5526 a_n7636_8799.n85 gnd 0.011862f
C5527 a_n7636_8799.t81 gnd 0.601377f
C5528 a_n7636_8799.n86 gnd 0.052275f
C5529 a_n7636_8799.t93 gnd 0.601377f
C5530 a_n7636_8799.n87 gnd 0.268587f
C5531 a_n7636_8799.n88 gnd 0.052275f
C5532 a_n7636_8799.n89 gnd 0.011862f
C5533 a_n7636_8799.t129 gnd 0.601377f
C5534 a_n7636_8799.n90 gnd 0.165151f
C5535 a_n7636_8799.t153 gnd 0.601377f
C5536 a_n7636_8799.t150 gnd 0.612759f
C5537 a_n7636_8799.n91 gnd 0.252102f
C5538 a_n7636_8799.n92 gnd 0.26488f
C5539 a_n7636_8799.n93 gnd 0.011862f
C5540 a_n7636_8799.t97 gnd 0.601377f
C5541 a_n7636_8799.n94 gnd 0.268587f
C5542 a_n7636_8799.n95 gnd 0.052275f
C5543 a_n7636_8799.n96 gnd 0.052275f
C5544 a_n7636_8799.n97 gnd 0.052275f
C5545 a_n7636_8799.n98 gnd 0.266492f
C5546 a_n7636_8799.t147 gnd 0.601377f
C5547 a_n7636_8799.n99 gnd 0.265202f
C5548 a_n7636_8799.n100 gnd 0.011862f
C5549 a_n7636_8799.n101 gnd 0.052275f
C5550 a_n7636_8799.n102 gnd 0.052275f
C5551 a_n7636_8799.n103 gnd 0.052275f
C5552 a_n7636_8799.n104 gnd 0.011862f
C5553 a_n7636_8799.t94 gnd 0.601377f
C5554 a_n7636_8799.n105 gnd 0.266169f
C5555 a_n7636_8799.t127 gnd 0.601377f
C5556 a_n7636_8799.n106 gnd 0.265525f
C5557 a_n7636_8799.n107 gnd 0.052275f
C5558 a_n7636_8799.n108 gnd 0.052275f
C5559 a_n7636_8799.n109 gnd 0.052275f
C5560 a_n7636_8799.n110 gnd 0.268587f
C5561 a_n7636_8799.n111 gnd 0.011862f
C5562 a_n7636_8799.t82 gnd 0.601377f
C5563 a_n7636_8799.n112 gnd 0.265847f
C5564 a_n7636_8799.n113 gnd 0.052275f
C5565 a_n7636_8799.n114 gnd 0.052275f
C5566 a_n7636_8799.n115 gnd 0.052275f
C5567 a_n7636_8799.n116 gnd 0.011862f
C5568 a_n7636_8799.t47 gnd 0.601377f
C5569 a_n7636_8799.n117 gnd 0.268587f
C5570 a_n7636_8799.n118 gnd 0.011862f
C5571 a_n7636_8799.n119 gnd 0.052275f
C5572 a_n7636_8799.n120 gnd 0.052275f
C5573 a_n7636_8799.n121 gnd 0.052275f
C5574 a_n7636_8799.n122 gnd 0.266169f
C5575 a_n7636_8799.n123 gnd 0.011862f
C5576 a_n7636_8799.t151 gnd 0.601377f
C5577 a_n7636_8799.n124 gnd 0.268587f
C5578 a_n7636_8799.n125 gnd 0.052275f
C5579 a_n7636_8799.n126 gnd 0.052275f
C5580 a_n7636_8799.n127 gnd 0.052275f
C5581 a_n7636_8799.n128 gnd 0.265202f
C5582 a_n7636_8799.t77 gnd 0.601377f
C5583 a_n7636_8799.n129 gnd 0.266492f
C5584 a_n7636_8799.n130 gnd 0.011862f
C5585 a_n7636_8799.n131 gnd 0.052275f
C5586 a_n7636_8799.n132 gnd 0.052275f
C5587 a_n7636_8799.n133 gnd 0.052275f
C5588 a_n7636_8799.n134 gnd 0.011862f
C5589 a_n7636_8799.t57 gnd 0.601377f
C5590 a_n7636_8799.n135 gnd 0.26488f
C5591 a_n7636_8799.t59 gnd 0.601377f
C5592 a_n7636_8799.n136 gnd 0.263108f
C5593 a_n7636_8799.n137 gnd 0.130296f
C5594 a_n7636_8799.n138 gnd 0.904087f
C5595 a_n7636_8799.n139 gnd 0.052275f
C5596 a_n7636_8799.t100 gnd 0.601377f
C5597 a_n7636_8799.n140 gnd 0.268587f
C5598 a_n7636_8799.n141 gnd 0.052275f
C5599 a_n7636_8799.n142 gnd 0.011862f
C5600 a_n7636_8799.t124 gnd 0.601377f
C5601 a_n7636_8799.n143 gnd 0.052275f
C5602 a_n7636_8799.t42 gnd 0.601377f
C5603 a_n7636_8799.n144 gnd 0.265525f
C5604 a_n7636_8799.t107 gnd 0.601377f
C5605 a_n7636_8799.n145 gnd 0.052275f
C5606 a_n7636_8799.t146 gnd 0.601377f
C5607 a_n7636_8799.n146 gnd 0.265847f
C5608 a_n7636_8799.n147 gnd 0.052275f
C5609 a_n7636_8799.n148 gnd 0.011862f
C5610 a_n7636_8799.t141 gnd 0.601377f
C5611 a_n7636_8799.n149 gnd 0.052275f
C5612 a_n7636_8799.t54 gnd 0.601377f
C5613 a_n7636_8799.n150 gnd 0.268587f
C5614 a_n7636_8799.n151 gnd 0.052275f
C5615 a_n7636_8799.n152 gnd 0.011862f
C5616 a_n7636_8799.t79 gnd 0.601377f
C5617 a_n7636_8799.n153 gnd 0.165151f
C5618 a_n7636_8799.t90 gnd 0.601377f
C5619 a_n7636_8799.t112 gnd 0.612759f
C5620 a_n7636_8799.n154 gnd 0.252102f
C5621 a_n7636_8799.n155 gnd 0.26488f
C5622 a_n7636_8799.n156 gnd 0.011862f
C5623 a_n7636_8799.t128 gnd 0.601377f
C5624 a_n7636_8799.n157 gnd 0.268587f
C5625 a_n7636_8799.n158 gnd 0.052275f
C5626 a_n7636_8799.n159 gnd 0.052275f
C5627 a_n7636_8799.n160 gnd 0.052275f
C5628 a_n7636_8799.n161 gnd 0.266492f
C5629 a_n7636_8799.t138 gnd 0.601377f
C5630 a_n7636_8799.n162 gnd 0.265202f
C5631 a_n7636_8799.n163 gnd 0.011862f
C5632 a_n7636_8799.n164 gnd 0.052275f
C5633 a_n7636_8799.n165 gnd 0.052275f
C5634 a_n7636_8799.n166 gnd 0.052275f
C5635 a_n7636_8799.n167 gnd 0.011862f
C5636 a_n7636_8799.t37 gnd 0.601377f
C5637 a_n7636_8799.n168 gnd 0.266169f
C5638 a_n7636_8799.t98 gnd 0.601377f
C5639 a_n7636_8799.n169 gnd 0.265525f
C5640 a_n7636_8799.n170 gnd 0.052275f
C5641 a_n7636_8799.n171 gnd 0.052275f
C5642 a_n7636_8799.n172 gnd 0.052275f
C5643 a_n7636_8799.n173 gnd 0.268587f
C5644 a_n7636_8799.n174 gnd 0.011862f
C5645 a_n7636_8799.t115 gnd 0.601377f
C5646 a_n7636_8799.n175 gnd 0.265847f
C5647 a_n7636_8799.n176 gnd 0.052275f
C5648 a_n7636_8799.n177 gnd 0.052275f
C5649 a_n7636_8799.n178 gnd 0.052275f
C5650 a_n7636_8799.n179 gnd 0.011862f
C5651 a_n7636_8799.t91 gnd 0.601377f
C5652 a_n7636_8799.n180 gnd 0.268587f
C5653 a_n7636_8799.n181 gnd 0.011862f
C5654 a_n7636_8799.n182 gnd 0.052275f
C5655 a_n7636_8799.n183 gnd 0.052275f
C5656 a_n7636_8799.n184 gnd 0.052275f
C5657 a_n7636_8799.n185 gnd 0.266169f
C5658 a_n7636_8799.n186 gnd 0.011862f
C5659 a_n7636_8799.t61 gnd 0.601377f
C5660 a_n7636_8799.n187 gnd 0.268587f
C5661 a_n7636_8799.n188 gnd 0.052275f
C5662 a_n7636_8799.n189 gnd 0.052275f
C5663 a_n7636_8799.n190 gnd 0.052275f
C5664 a_n7636_8799.n191 gnd 0.265202f
C5665 a_n7636_8799.t70 gnd 0.601377f
C5666 a_n7636_8799.n192 gnd 0.266492f
C5667 a_n7636_8799.n193 gnd 0.011862f
C5668 a_n7636_8799.n194 gnd 0.052275f
C5669 a_n7636_8799.n195 gnd 0.052275f
C5670 a_n7636_8799.n196 gnd 0.052275f
C5671 a_n7636_8799.n197 gnd 0.011862f
C5672 a_n7636_8799.t50 gnd 0.601377f
C5673 a_n7636_8799.n198 gnd 0.26488f
C5674 a_n7636_8799.t152 gnd 0.601377f
C5675 a_n7636_8799.n199 gnd 0.263108f
C5676 a_n7636_8799.n200 gnd 0.130296f
C5677 a_n7636_8799.n201 gnd 1.50453f
C5678 a_n7636_8799.n202 gnd 0.052275f
C5679 a_n7636_8799.t86 gnd 0.601377f
C5680 a_n7636_8799.t85 gnd 0.601377f
C5681 a_n7636_8799.t58 gnd 0.601377f
C5682 a_n7636_8799.n203 gnd 0.268587f
C5683 a_n7636_8799.n204 gnd 0.052275f
C5684 a_n7636_8799.t134 gnd 0.601377f
C5685 a_n7636_8799.t89 gnd 0.601377f
C5686 a_n7636_8799.n205 gnd 0.052275f
C5687 a_n7636_8799.t65 gnd 0.601377f
C5688 a_n7636_8799.n206 gnd 0.268587f
C5689 a_n7636_8799.n207 gnd 0.052275f
C5690 a_n7636_8799.t140 gnd 0.601377f
C5691 a_n7636_8799.t106 gnd 0.601377f
C5692 a_n7636_8799.n208 gnd 0.052275f
C5693 a_n7636_8799.t104 gnd 0.601377f
C5694 a_n7636_8799.n209 gnd 0.268587f
C5695 a_n7636_8799.n210 gnd 0.052275f
C5696 a_n7636_8799.t39 gnd 0.601377f
C5697 a_n7636_8799.t110 gnd 0.601377f
C5698 a_n7636_8799.n211 gnd 0.052275f
C5699 a_n7636_8799.t109 gnd 0.601377f
C5700 a_n7636_8799.n212 gnd 0.268587f
C5701 a_n7636_8799.n213 gnd 0.052275f
C5702 a_n7636_8799.t41 gnd 0.601377f
C5703 a_n7636_8799.t40 gnd 0.601377f
C5704 a_n7636_8799.n214 gnd 0.052275f
C5705 a_n7636_8799.t126 gnd 0.601377f
C5706 a_n7636_8799.n215 gnd 0.268587f
C5707 a_n7636_8799.n216 gnd 0.052275f
C5708 a_n7636_8799.t60 gnd 0.601377f
C5709 a_n7636_8799.t44 gnd 0.601377f
C5710 a_n7636_8799.n217 gnd 0.052275f
C5711 a_n7636_8799.t130 gnd 0.601377f
C5712 a_n7636_8799.n218 gnd 0.268587f
C5713 a_n7636_8799.t64 gnd 0.612759f
C5714 a_n7636_8799.n219 gnd 0.252102f
C5715 a_n7636_8799.t88 gnd 0.601377f
C5716 a_n7636_8799.n220 gnd 0.26488f
C5717 a_n7636_8799.n221 gnd 0.011862f
C5718 a_n7636_8799.n222 gnd 0.165151f
C5719 a_n7636_8799.n223 gnd 0.052275f
C5720 a_n7636_8799.n224 gnd 0.052275f
C5721 a_n7636_8799.n225 gnd 0.011862f
C5722 a_n7636_8799.n226 gnd 0.266492f
C5723 a_n7636_8799.n227 gnd 0.265202f
C5724 a_n7636_8799.n228 gnd 0.011862f
C5725 a_n7636_8799.n229 gnd 0.052275f
C5726 a_n7636_8799.n230 gnd 0.052275f
C5727 a_n7636_8799.n231 gnd 0.052275f
C5728 a_n7636_8799.n232 gnd 0.011862f
C5729 a_n7636_8799.n233 gnd 0.266169f
C5730 a_n7636_8799.n234 gnd 0.265525f
C5731 a_n7636_8799.n235 gnd 0.011862f
C5732 a_n7636_8799.n236 gnd 0.052275f
C5733 a_n7636_8799.n237 gnd 0.052275f
C5734 a_n7636_8799.n238 gnd 0.052275f
C5735 a_n7636_8799.n239 gnd 0.011862f
C5736 a_n7636_8799.n240 gnd 0.265847f
C5737 a_n7636_8799.n241 gnd 0.265847f
C5738 a_n7636_8799.n242 gnd 0.011862f
C5739 a_n7636_8799.n243 gnd 0.052275f
C5740 a_n7636_8799.n244 gnd 0.052275f
C5741 a_n7636_8799.n245 gnd 0.052275f
C5742 a_n7636_8799.n246 gnd 0.011862f
C5743 a_n7636_8799.n247 gnd 0.265525f
C5744 a_n7636_8799.n248 gnd 0.266169f
C5745 a_n7636_8799.n249 gnd 0.011862f
C5746 a_n7636_8799.n250 gnd 0.052275f
C5747 a_n7636_8799.n251 gnd 0.052275f
C5748 a_n7636_8799.n252 gnd 0.052275f
C5749 a_n7636_8799.n253 gnd 0.011862f
C5750 a_n7636_8799.n254 gnd 0.265202f
C5751 a_n7636_8799.n255 gnd 0.266492f
C5752 a_n7636_8799.n256 gnd 0.011862f
C5753 a_n7636_8799.n257 gnd 0.052275f
C5754 a_n7636_8799.n258 gnd 0.052275f
C5755 a_n7636_8799.n259 gnd 0.052275f
C5756 a_n7636_8799.n260 gnd 0.011862f
C5757 a_n7636_8799.n261 gnd 0.26488f
C5758 a_n7636_8799.n262 gnd 0.263108f
C5759 a_n7636_8799.n263 gnd 0.296385f
C5760 a_n7636_8799.n264 gnd 0.052275f
C5761 a_n7636_8799.t96 gnd 0.601377f
C5762 a_n7636_8799.t95 gnd 0.601377f
C5763 a_n7636_8799.t73 gnd 0.601377f
C5764 a_n7636_8799.n265 gnd 0.268587f
C5765 a_n7636_8799.n266 gnd 0.052275f
C5766 a_n7636_8799.t149 gnd 0.601377f
C5767 a_n7636_8799.t102 gnd 0.601377f
C5768 a_n7636_8799.n267 gnd 0.052275f
C5769 a_n7636_8799.t75 gnd 0.601377f
C5770 a_n7636_8799.n268 gnd 0.268587f
C5771 a_n7636_8799.n269 gnd 0.052275f
C5772 a_n7636_8799.t155 gnd 0.601377f
C5773 a_n7636_8799.t119 gnd 0.601377f
C5774 a_n7636_8799.n270 gnd 0.052275f
C5775 a_n7636_8799.t118 gnd 0.601377f
C5776 a_n7636_8799.n271 gnd 0.268587f
C5777 a_n7636_8799.n272 gnd 0.052275f
C5778 a_n7636_8799.t49 gnd 0.601377f
C5779 a_n7636_8799.t122 gnd 0.601377f
C5780 a_n7636_8799.n273 gnd 0.052275f
C5781 a_n7636_8799.t121 gnd 0.601377f
C5782 a_n7636_8799.n274 gnd 0.268587f
C5783 a_n7636_8799.n275 gnd 0.052275f
C5784 a_n7636_8799.t53 gnd 0.601377f
C5785 a_n7636_8799.t52 gnd 0.601377f
C5786 a_n7636_8799.n276 gnd 0.052275f
C5787 a_n7636_8799.t143 gnd 0.601377f
C5788 a_n7636_8799.n277 gnd 0.268587f
C5789 a_n7636_8799.n278 gnd 0.052275f
C5790 a_n7636_8799.t74 gnd 0.601377f
C5791 a_n7636_8799.t56 gnd 0.601377f
C5792 a_n7636_8799.n279 gnd 0.052275f
C5793 a_n7636_8799.t144 gnd 0.601377f
C5794 a_n7636_8799.n280 gnd 0.268587f
C5795 a_n7636_8799.t76 gnd 0.612759f
C5796 a_n7636_8799.n281 gnd 0.252102f
C5797 a_n7636_8799.t103 gnd 0.601377f
C5798 a_n7636_8799.n282 gnd 0.26488f
C5799 a_n7636_8799.n283 gnd 0.011862f
C5800 a_n7636_8799.n284 gnd 0.165151f
C5801 a_n7636_8799.n285 gnd 0.052275f
C5802 a_n7636_8799.n286 gnd 0.052275f
C5803 a_n7636_8799.n287 gnd 0.011862f
C5804 a_n7636_8799.n288 gnd 0.266492f
C5805 a_n7636_8799.n289 gnd 0.265202f
C5806 a_n7636_8799.n290 gnd 0.011862f
C5807 a_n7636_8799.n291 gnd 0.052275f
C5808 a_n7636_8799.n292 gnd 0.052275f
C5809 a_n7636_8799.n293 gnd 0.052275f
C5810 a_n7636_8799.n294 gnd 0.011862f
C5811 a_n7636_8799.n295 gnd 0.266169f
C5812 a_n7636_8799.n296 gnd 0.265525f
C5813 a_n7636_8799.n297 gnd 0.011862f
C5814 a_n7636_8799.n298 gnd 0.052275f
C5815 a_n7636_8799.n299 gnd 0.052275f
C5816 a_n7636_8799.n300 gnd 0.052275f
C5817 a_n7636_8799.n301 gnd 0.011862f
C5818 a_n7636_8799.n302 gnd 0.265847f
C5819 a_n7636_8799.n303 gnd 0.265847f
C5820 a_n7636_8799.n304 gnd 0.011862f
C5821 a_n7636_8799.n305 gnd 0.052275f
C5822 a_n7636_8799.n306 gnd 0.052275f
C5823 a_n7636_8799.n307 gnd 0.052275f
C5824 a_n7636_8799.n308 gnd 0.011862f
C5825 a_n7636_8799.n309 gnd 0.265525f
C5826 a_n7636_8799.n310 gnd 0.266169f
C5827 a_n7636_8799.n311 gnd 0.011862f
C5828 a_n7636_8799.n312 gnd 0.052275f
C5829 a_n7636_8799.n313 gnd 0.052275f
C5830 a_n7636_8799.n314 gnd 0.052275f
C5831 a_n7636_8799.n315 gnd 0.011862f
C5832 a_n7636_8799.n316 gnd 0.265202f
C5833 a_n7636_8799.n317 gnd 0.266492f
C5834 a_n7636_8799.n318 gnd 0.011862f
C5835 a_n7636_8799.n319 gnd 0.052275f
C5836 a_n7636_8799.n320 gnd 0.052275f
C5837 a_n7636_8799.n321 gnd 0.052275f
C5838 a_n7636_8799.n322 gnd 0.011862f
C5839 a_n7636_8799.n323 gnd 0.26488f
C5840 a_n7636_8799.n324 gnd 0.263108f
C5841 a_n7636_8799.n325 gnd 0.130296f
C5842 a_n7636_8799.n326 gnd 0.904087f
C5843 a_n7636_8799.n327 gnd 0.052275f
C5844 a_n7636_8799.t154 gnd 0.601377f
C5845 a_n7636_8799.t51 gnd 0.601377f
C5846 a_n7636_8799.t101 gnd 0.601377f
C5847 a_n7636_8799.n328 gnd 0.268587f
C5848 a_n7636_8799.n329 gnd 0.052275f
C5849 a_n7636_8799.t38 gnd 0.601377f
C5850 a_n7636_8799.t125 gnd 0.601377f
C5851 a_n7636_8799.n330 gnd 0.052275f
C5852 a_n7636_8799.t62 gnd 0.601377f
C5853 a_n7636_8799.n331 gnd 0.268587f
C5854 a_n7636_8799.n332 gnd 0.052275f
C5855 a_n7636_8799.t108 gnd 0.601377f
C5856 a_n7636_8799.t43 gnd 0.601377f
C5857 a_n7636_8799.n333 gnd 0.052275f
C5858 a_n7636_8799.t68 gnd 0.601377f
C5859 a_n7636_8799.n334 gnd 0.268587f
C5860 a_n7636_8799.n335 gnd 0.052275f
C5861 a_n7636_8799.t148 gnd 0.601377f
C5862 a_n7636_8799.t117 gnd 0.601377f
C5863 a_n7636_8799.n336 gnd 0.052275f
C5864 a_n7636_8799.t142 gnd 0.601377f
C5865 a_n7636_8799.n337 gnd 0.268587f
C5866 a_n7636_8799.n338 gnd 0.052275f
C5867 a_n7636_8799.t99 gnd 0.601377f
C5868 a_n7636_8799.t120 gnd 0.601377f
C5869 a_n7636_8799.n339 gnd 0.052275f
C5870 a_n7636_8799.t55 gnd 0.601377f
C5871 a_n7636_8799.n340 gnd 0.268587f
C5872 a_n7636_8799.n341 gnd 0.052275f
C5873 a_n7636_8799.t139 gnd 0.601377f
C5874 a_n7636_8799.t80 gnd 0.601377f
C5875 a_n7636_8799.n342 gnd 0.052275f
C5876 a_n7636_8799.t131 gnd 0.601377f
C5877 a_n7636_8799.n343 gnd 0.268587f
C5878 a_n7636_8799.t113 gnd 0.612759f
C5879 a_n7636_8799.n344 gnd 0.252102f
C5880 a_n7636_8799.t67 gnd 0.601377f
C5881 a_n7636_8799.n345 gnd 0.26488f
C5882 a_n7636_8799.n346 gnd 0.011862f
C5883 a_n7636_8799.n347 gnd 0.165151f
C5884 a_n7636_8799.n348 gnd 0.052275f
C5885 a_n7636_8799.n349 gnd 0.052275f
C5886 a_n7636_8799.n350 gnd 0.011862f
C5887 a_n7636_8799.n351 gnd 0.266492f
C5888 a_n7636_8799.n352 gnd 0.265202f
C5889 a_n7636_8799.n353 gnd 0.011862f
C5890 a_n7636_8799.n354 gnd 0.052275f
C5891 a_n7636_8799.n355 gnd 0.052275f
C5892 a_n7636_8799.n356 gnd 0.052275f
C5893 a_n7636_8799.n357 gnd 0.011862f
C5894 a_n7636_8799.n358 gnd 0.266169f
C5895 a_n7636_8799.n359 gnd 0.265525f
C5896 a_n7636_8799.n360 gnd 0.011862f
C5897 a_n7636_8799.n361 gnd 0.052275f
C5898 a_n7636_8799.n362 gnd 0.052275f
C5899 a_n7636_8799.n363 gnd 0.052275f
C5900 a_n7636_8799.n364 gnd 0.011862f
C5901 a_n7636_8799.n365 gnd 0.265847f
C5902 a_n7636_8799.n366 gnd 0.265847f
C5903 a_n7636_8799.n367 gnd 0.011862f
C5904 a_n7636_8799.n368 gnd 0.052275f
C5905 a_n7636_8799.n369 gnd 0.052275f
C5906 a_n7636_8799.n370 gnd 0.052275f
C5907 a_n7636_8799.n371 gnd 0.011862f
C5908 a_n7636_8799.n372 gnd 0.265525f
C5909 a_n7636_8799.n373 gnd 0.266169f
C5910 a_n7636_8799.n374 gnd 0.011862f
C5911 a_n7636_8799.n375 gnd 0.052275f
C5912 a_n7636_8799.n376 gnd 0.052275f
C5913 a_n7636_8799.n377 gnd 0.052275f
C5914 a_n7636_8799.n378 gnd 0.011862f
C5915 a_n7636_8799.n379 gnd 0.265202f
C5916 a_n7636_8799.n380 gnd 0.266492f
C5917 a_n7636_8799.n381 gnd 0.011862f
C5918 a_n7636_8799.n382 gnd 0.052275f
C5919 a_n7636_8799.n383 gnd 0.052275f
C5920 a_n7636_8799.n384 gnd 0.052275f
C5921 a_n7636_8799.n385 gnd 0.011862f
C5922 a_n7636_8799.n386 gnd 0.26488f
C5923 a_n7636_8799.n387 gnd 0.263108f
C5924 a_n7636_8799.n388 gnd 0.130296f
C5925 a_n7636_8799.n389 gnd 1.11709f
C5926 a_n7636_8799.n390 gnd 12.302299f
C5927 a_n7636_8799.n391 gnd 4.40121f
C5928 a_n7636_8799.t13 gnd 0.112804f
C5929 a_n7636_8799.t14 gnd 0.112804f
C5930 a_n7636_8799.n392 gnd 0.998992f
C5931 a_n7636_8799.t7 gnd 0.112804f
C5932 a_n7636_8799.t8 gnd 0.112804f
C5933 a_n7636_8799.n393 gnd 0.996776f
C5934 a_n7636_8799.n394 gnd 0.793977f
C5935 a_n7636_8799.t6 gnd 0.112804f
C5936 a_n7636_8799.t24 gnd 0.112804f
C5937 a_n7636_8799.n395 gnd 0.996776f
C5938 a_n7636_8799.n396 gnd 0.331538f
C5939 a_n7636_8799.n397 gnd 0.47333f
C5940 a_n7636_8799.t26 gnd 0.112804f
C5941 a_n7636_8799.t19 gnd 0.112804f
C5942 a_n7636_8799.n398 gnd 0.996776f
C5943 a_n7636_8799.n399 gnd 0.331538f
C5944 a_n7636_8799.t21 gnd 0.112804f
C5945 a_n7636_8799.t5 gnd 0.112804f
C5946 a_n7636_8799.n400 gnd 0.996776f
C5947 a_n7636_8799.n401 gnd 0.389883f
C5948 a_n7636_8799.t23 gnd 0.112804f
C5949 a_n7636_8799.t25 gnd 0.112804f
C5950 a_n7636_8799.n402 gnd 0.996776f
C5951 a_n7636_8799.n403 gnd 2.87037f
C5952 a_n7636_8799.t20 gnd 0.112804f
C5953 a_n7636_8799.t18 gnd 0.112804f
C5954 a_n7636_8799.n404 gnd 0.998992f
C5955 a_n7636_8799.t9 gnd 0.112804f
C5956 a_n7636_8799.t15 gnd 0.112804f
C5957 a_n7636_8799.n405 gnd 0.996775f
C5958 a_n7636_8799.n406 gnd 0.793979f
C5959 a_n7636_8799.t27 gnd 0.112804f
C5960 a_n7636_8799.t10 gnd 0.112804f
C5961 a_n7636_8799.n407 gnd 0.996775f
C5962 a_n7636_8799.n408 gnd 0.331539f
C5963 a_n7636_8799.n409 gnd 2.41583f
C5964 a_n7636_8799.n410 gnd 0.331541f
C5965 a_n7636_8799.n411 gnd 0.996772f
C5966 a_n7636_8799.t28 gnd 0.112804f
C5967 a_n2903_n3924.n0 gnd 2.10908f
C5968 a_n2903_n3924.n1 gnd 2.29654f
C5969 a_n2903_n3924.n2 gnd 1.52909f
C5970 a_n2903_n3924.n3 gnd 1.39023f
C5971 a_n2903_n3924.n4 gnd 1.91428f
C5972 a_n2903_n3924.n5 gnd 1.87222f
C5973 a_n2903_n3924.n6 gnd 1.87222f
C5974 a_n2903_n3924.n7 gnd 2.19334f
C5975 a_n2903_n3924.n8 gnd 1.00796f
C5976 a_n2903_n3924.n9 gnd 0.764541f
C5977 a_n2903_n3924.n10 gnd 1.34454f
C5978 a_n2903_n3924.n11 gnd 1.6947f
C5979 a_n2903_n3924.t54 gnd 0.102925f
C5980 a_n2903_n3924.t13 gnd 0.102925f
C5981 a_n2903_n3924.t51 gnd 0.102925f
C5982 a_n2903_n3924.n12 gnd 0.840609f
C5983 a_n2903_n3924.t11 gnd 1.3291f
C5984 a_n2903_n3924.t50 gnd 0.102925f
C5985 a_n2903_n3924.t22 gnd 0.102925f
C5986 a_n2903_n3924.n13 gnd 0.840609f
C5987 a_n2903_n3924.t49 gnd 0.102925f
C5988 a_n2903_n3924.t17 gnd 0.102925f
C5989 a_n2903_n3924.n14 gnd 0.840609f
C5990 a_n2903_n3924.t3 gnd 0.102925f
C5991 a_n2903_n3924.t14 gnd 0.102925f
C5992 a_n2903_n3924.n15 gnd 0.840609f
C5993 a_n2903_n3924.t52 gnd 1.06972f
C5994 a_n2903_n3924.t21 gnd 1.32974f
C5995 a_n2903_n3924.t55 gnd 1.3291f
C5996 a_n2903_n3924.t9 gnd 1.3291f
C5997 a_n2903_n3924.t18 gnd 1.3291f
C5998 a_n2903_n3924.t10 gnd 1.3291f
C5999 a_n2903_n3924.t12 gnd 1.3291f
C6000 a_n2903_n3924.t48 gnd 1.3291f
C6001 a_n2903_n3924.n16 gnd 0.965474f
C6002 a_n2903_n3924.t46 gnd 1.06972f
C6003 a_n2903_n3924.t32 gnd 0.102925f
C6004 a_n2903_n3924.t35 gnd 0.102925f
C6005 a_n2903_n3924.n17 gnd 0.840607f
C6006 a_n2903_n3924.t41 gnd 0.102925f
C6007 a_n2903_n3924.t24 gnd 0.102925f
C6008 a_n2903_n3924.n18 gnd 0.840607f
C6009 a_n2903_n3924.t40 gnd 0.102925f
C6010 a_n2903_n3924.t33 gnd 0.102925f
C6011 a_n2903_n3924.n19 gnd 0.840607f
C6012 a_n2903_n3924.t31 gnd 0.102925f
C6013 a_n2903_n3924.t23 gnd 0.102925f
C6014 a_n2903_n3924.n20 gnd 0.840607f
C6015 a_n2903_n3924.t30 gnd 0.102925f
C6016 a_n2903_n3924.t27 gnd 0.102925f
C6017 a_n2903_n3924.n21 gnd 0.840607f
C6018 a_n2903_n3924.t38 gnd 1.06972f
C6019 a_n2903_n3924.t20 gnd 1.06972f
C6020 a_n2903_n3924.t15 gnd 0.102925f
C6021 a_n2903_n3924.t47 gnd 0.102925f
C6022 a_n2903_n3924.n22 gnd 0.840607f
C6023 a_n2903_n3924.t8 gnd 0.102925f
C6024 a_n2903_n3924.t2 gnd 0.102925f
C6025 a_n2903_n3924.n23 gnd 0.840607f
C6026 a_n2903_n3924.t1 gnd 0.102925f
C6027 a_n2903_n3924.t5 gnd 0.102925f
C6028 a_n2903_n3924.n24 gnd 0.840607f
C6029 a_n2903_n3924.t4 gnd 0.102925f
C6030 a_n2903_n3924.t6 gnd 0.102925f
C6031 a_n2903_n3924.n25 gnd 0.840607f
C6032 a_n2903_n3924.t19 gnd 0.102925f
C6033 a_n2903_n3924.t53 gnd 0.102925f
C6034 a_n2903_n3924.n26 gnd 0.840607f
C6035 a_n2903_n3924.t7 gnd 1.06972f
C6036 a_n2903_n3924.n27 gnd 1.02539f
C6037 a_n2903_n3924.t37 gnd 1.06972f
C6038 a_n2903_n3924.t43 gnd 0.102925f
C6039 a_n2903_n3924.t26 gnd 0.102925f
C6040 a_n2903_n3924.n28 gnd 0.840609f
C6041 a_n2903_n3924.t29 gnd 0.102925f
C6042 a_n2903_n3924.t34 gnd 0.102925f
C6043 a_n2903_n3924.n29 gnd 0.840609f
C6044 a_n2903_n3924.t39 gnd 0.102925f
C6045 a_n2903_n3924.t28 gnd 0.102925f
C6046 a_n2903_n3924.n30 gnd 0.840609f
C6047 a_n2903_n3924.t42 gnd 0.102925f
C6048 a_n2903_n3924.t45 gnd 0.102925f
C6049 a_n2903_n3924.n31 gnd 0.840609f
C6050 a_n2903_n3924.t25 gnd 0.102925f
C6051 a_n2903_n3924.t44 gnd 0.102925f
C6052 a_n2903_n3924.n32 gnd 0.840609f
C6053 a_n2903_n3924.t36 gnd 1.06972f
C6054 a_n2903_n3924.t16 gnd 1.06972f
C6055 a_n2903_n3924.n33 gnd 0.84061f
C6056 a_n2903_n3924.t0 gnd 0.102925f
C6057 plus.n0 gnd 0.02427f
C6058 plus.t21 gnd 0.343283f
C6059 plus.n1 gnd 0.02427f
C6060 plus.t22 gnd 0.343283f
C6061 plus.t16 gnd 0.343283f
C6062 plus.n2 gnd 0.152497f
C6063 plus.n3 gnd 0.02427f
C6064 plus.t17 gnd 0.343283f
C6065 plus.t11 gnd 0.343283f
C6066 plus.n4 gnd 0.152497f
C6067 plus.n5 gnd 0.02427f
C6068 plus.t5 gnd 0.343283f
C6069 plus.t6 gnd 0.343283f
C6070 plus.n6 gnd 0.152497f
C6071 plus.n7 gnd 0.02427f
C6072 plus.t23 gnd 0.343283f
C6073 plus.t24 gnd 0.343283f
C6074 plus.n8 gnd 0.152497f
C6075 plus.n9 gnd 0.02427f
C6076 plus.t18 gnd 0.343283f
C6077 plus.t13 gnd 0.343283f
C6078 plus.n10 gnd 0.157464f
C6079 plus.t15 gnd 0.355744f
C6080 plus.n11 gnd 0.141329f
C6081 plus.n12 gnd 0.104486f
C6082 plus.n13 gnd 0.005507f
C6083 plus.n14 gnd 0.152497f
C6084 plus.n15 gnd 0.005507f
C6085 plus.n16 gnd 0.02427f
C6086 plus.n17 gnd 0.02427f
C6087 plus.n18 gnd 0.02427f
C6088 plus.n19 gnd 0.005507f
C6089 plus.n20 gnd 0.152497f
C6090 plus.n21 gnd 0.005507f
C6091 plus.n22 gnd 0.02427f
C6092 plus.n23 gnd 0.02427f
C6093 plus.n24 gnd 0.02427f
C6094 plus.n25 gnd 0.005507f
C6095 plus.n26 gnd 0.152497f
C6096 plus.n27 gnd 0.005507f
C6097 plus.n28 gnd 0.02427f
C6098 plus.n29 gnd 0.02427f
C6099 plus.n30 gnd 0.02427f
C6100 plus.n31 gnd 0.005507f
C6101 plus.n32 gnd 0.152497f
C6102 plus.n33 gnd 0.005507f
C6103 plus.n34 gnd 0.02427f
C6104 plus.n35 gnd 0.02427f
C6105 plus.n36 gnd 0.02427f
C6106 plus.n37 gnd 0.005507f
C6107 plus.n38 gnd 0.152497f
C6108 plus.n39 gnd 0.005507f
C6109 plus.n40 gnd 0.152722f
C6110 plus.n41 gnd 0.274825f
C6111 plus.n42 gnd 0.02427f
C6112 plus.n43 gnd 0.005507f
C6113 plus.t10 gnd 0.343283f
C6114 plus.n44 gnd 0.02427f
C6115 plus.n45 gnd 0.005507f
C6116 plus.t12 gnd 0.343283f
C6117 plus.n46 gnd 0.02427f
C6118 plus.n47 gnd 0.005507f
C6119 plus.t7 gnd 0.343283f
C6120 plus.n48 gnd 0.02427f
C6121 plus.n49 gnd 0.005507f
C6122 plus.t27 gnd 0.343283f
C6123 plus.n50 gnd 0.02427f
C6124 plus.n51 gnd 0.005507f
C6125 plus.t26 gnd 0.343283f
C6126 plus.t20 gnd 0.355744f
C6127 plus.t19 gnd 0.343283f
C6128 plus.n52 gnd 0.157464f
C6129 plus.n53 gnd 0.141329f
C6130 plus.n54 gnd 0.104486f
C6131 plus.n55 gnd 0.02427f
C6132 plus.n56 gnd 0.152497f
C6133 plus.n57 gnd 0.005507f
C6134 plus.t25 gnd 0.343283f
C6135 plus.n58 gnd 0.152497f
C6136 plus.n59 gnd 0.02427f
C6137 plus.n60 gnd 0.02427f
C6138 plus.n61 gnd 0.02427f
C6139 plus.n62 gnd 0.152497f
C6140 plus.n63 gnd 0.005507f
C6141 plus.t9 gnd 0.343283f
C6142 plus.n64 gnd 0.152497f
C6143 plus.n65 gnd 0.02427f
C6144 plus.n66 gnd 0.02427f
C6145 plus.n67 gnd 0.02427f
C6146 plus.n68 gnd 0.152497f
C6147 plus.n69 gnd 0.005507f
C6148 plus.t14 gnd 0.343283f
C6149 plus.n70 gnd 0.152497f
C6150 plus.n71 gnd 0.02427f
C6151 plus.n72 gnd 0.02427f
C6152 plus.n73 gnd 0.02427f
C6153 plus.n74 gnd 0.152497f
C6154 plus.n75 gnd 0.005507f
C6155 plus.t28 gnd 0.343283f
C6156 plus.n76 gnd 0.152497f
C6157 plus.n77 gnd 0.02427f
C6158 plus.n78 gnd 0.02427f
C6159 plus.n79 gnd 0.02427f
C6160 plus.n80 gnd 0.152497f
C6161 plus.n81 gnd 0.005507f
C6162 plus.t8 gnd 0.343283f
C6163 plus.n82 gnd 0.152722f
C6164 plus.n83 gnd 0.803355f
C6165 plus.n84 gnd 1.20187f
C6166 plus.t2 gnd 0.041898f
C6167 plus.t0 gnd 0.007482f
C6168 plus.t3 gnd 0.007482f
C6169 plus.n85 gnd 0.024265f
C6170 plus.n86 gnd 0.188372f
C6171 plus.t1 gnd 0.007482f
C6172 plus.t4 gnd 0.007482f
C6173 plus.n87 gnd 0.024265f
C6174 plus.n88 gnd 0.141396f
C6175 plus.n89 gnd 2.59439f
.ends

