* NGSPICE file created from opamp633.ext - technology: sky130A

.subckt opamp633 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n1808_13878.t19 a_n1986_13878.t34 a_n1986_13878.t35 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X1 a_n1808_13878.t5 a_n1986_13878.t40 vdd.t188 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 CSoutput.t79 a_n5644_8799.t28 vdd.t118 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X3 CSoutput.t98 commonsourceibias.t64 gnd.t172 gnd.t103 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X4 CSoutput.t144 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X5 CSoutput.t99 commonsourceibias.t65 gnd.t171 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X6 a_n5644_8799.t3 plus.t5 a_n2903_n3924.t37 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X7 CSoutput.t117 commonsourceibias.t66 gnd.t170 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 gnd.t169 commonsourceibias.t67 CSoutput.t118 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 vdd.t91 vdd.t89 vdd.t90 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X10 minus.t4 gnd.t316 gnd.t318 gnd.t317 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X11 a_n1986_8322.t21 a_n1986_13878.t41 a_n5644_8799.t24 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X12 vdd.t125 CSoutput.t145 output.t18 gnd.t345 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X13 gnd.t168 commonsourceibias.t68 CSoutput.t132 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X14 CSoutput.t133 commonsourceibias.t69 gnd.t167 gnd.t92 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X15 CSoutput.t25 commonsourceibias.t70 gnd.t166 gnd.t92 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 CSoutput.t26 commonsourceibias.t71 gnd.t165 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 gnd.t164 commonsourceibias.t72 CSoutput.t100 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 gnd.t163 commonsourceibias.t73 CSoutput.t101 gnd.t73 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X19 commonsourceibias.t1 commonsourceibias.t0 gnd.t161 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 CSoutput.t80 commonsourceibias.t74 gnd.t162 gnd.t108 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X21 CSoutput.t81 commonsourceibias.t75 gnd.t160 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 a_n1986_13878.t1 minus.t5 a_n2903_n3924.t7 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X23 a_n5644_8799.t2 plus.t6 a_n2903_n3924.t36 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X24 CSoutput.t78 a_n5644_8799.t29 vdd.t111 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X25 vdd.t193 a_n5644_8799.t30 CSoutput.t77 vdd.t101 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X26 a_n1986_13878.t0 minus.t6 a_n2903_n3924.t6 gnd.t319 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X27 a_n5644_8799.t21 a_n1986_13878.t42 a_n1986_8322.t20 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X28 vdd.t119 a_n5644_8799.t31 CSoutput.t76 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X29 CSoutput.t146 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X30 CSoutput.t75 a_n5644_8799.t32 vdd.t121 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X31 CSoutput.t122 commonsourceibias.t76 gnd.t159 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 gnd.t158 commonsourceibias.t77 CSoutput.t123 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X33 CSoutput.t27 commonsourceibias.t78 gnd.t157 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X34 CSoutput.t28 commonsourceibias.t79 gnd.t156 gnd.t103 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 gnd.t315 gnd.t313 gnd.t314 gnd.t240 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X36 gnd.t312 gnd.t310 gnd.t311 gnd.t226 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X37 vdd.t88 vdd.t86 vdd.t87 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X38 a_n2903_n3924.t35 plus.t7 a_n5644_8799.t12 gnd.t329 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X39 CSoutput.t124 commonsourceibias.t80 gnd.t155 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 CSoutput.t74 a_n5644_8799.t33 vdd.t13 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X41 a_n2903_n3924.t10 minus.t7 a_n1986_13878.t4 gnd.t327 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X42 gnd.t154 commonsourceibias.t81 CSoutput.t125 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 a_n2903_n3924.t2 diffpairibias.t16 gnd.t178 gnd.t177 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X44 CSoutput.t91 commonsourceibias.t82 gnd.t153 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X45 gnd.t106 commonsourceibias.t44 commonsourceibias.t45 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X46 output.t2 outputibias.t8 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X47 CSoutput.t92 commonsourceibias.t83 gnd.t152 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X48 gnd.t151 commonsourceibias.t84 CSoutput.t0 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 a_n1808_13878.t18 a_n1986_13878.t32 a_n1986_13878.t33 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X50 a_n1986_13878.t21 a_n1986_13878.t20 a_n1808_13878.t17 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X51 CSoutput.t73 a_n5644_8799.t34 vdd.t190 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X52 vdd.t189 a_n5644_8799.t35 CSoutput.t72 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 CSoutput.t1 commonsourceibias.t85 gnd.t150 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X54 CSoutput.t5 commonsourceibias.t86 gnd.t149 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 vdd.t94 CSoutput.t147 output.t17 gnd.t344 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X56 gnd.t148 commonsourceibias.t87 CSoutput.t6 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X57 gnd.t306 gnd.t304 plus.t4 gnd.t305 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X58 gnd.t147 commonsourceibias.t88 CSoutput.t134 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X59 vdd.t85 vdd.t83 vdd.t84 vdd.t53 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X60 CSoutput.t135 commonsourceibias.t89 gnd.t146 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X61 a_n2903_n3924.t34 plus.t8 a_n5644_8799.t9 gnd.t321 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X62 gnd.t309 gnd.t307 gnd.t308 gnd.t240 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X63 gnd.t303 gnd.t300 gnd.t302 gnd.t301 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X64 CSoutput.t137 commonsourceibias.t90 gnd.t145 gnd.t92 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X65 gnd.t144 commonsourceibias.t28 commonsourceibias.t29 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X66 diffpairibias.t15 diffpairibias.t14 gnd.t12 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X67 gnd.t143 commonsourceibias.t91 CSoutput.t138 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 CSoutput.t104 commonsourceibias.t92 gnd.t142 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X69 CSoutput.t105 commonsourceibias.t93 gnd.t141 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X70 vdd.t82 vdd.t80 vdd.t81 vdd.t32 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X71 gnd.t140 commonsourceibias.t94 CSoutput.t106 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X72 gnd.t139 commonsourceibias.t95 CSoutput.t107 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X73 vdd.t110 a_n5644_8799.t36 CSoutput.t71 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 CSoutput.t70 a_n5644_8799.t37 vdd.t138 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X75 vdd.t9 a_n5644_8799.t38 CSoutput.t69 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X76 CSoutput.t22 commonsourceibias.t96 gnd.t138 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X77 diffpairibias.t13 diffpairibias.t12 gnd.t324 gnd.t323 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X78 gnd.t137 commonsourceibias.t60 commonsourceibias.t61 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 CSoutput.t82 commonsourceibias.t97 gnd.t136 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 CSoutput.t136 commonsourceibias.t98 gnd.t135 gnd.t108 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X81 gnd.t299 gnd.t297 gnd.t298 gnd.t222 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X82 gnd.t134 commonsourceibias.t99 CSoutput.t85 gnd.t73 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X83 CSoutput.t139 commonsourceibias.t100 gnd.t133 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 gnd.t132 commonsourceibias.t101 CSoutput.t86 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 CSoutput.t68 a_n5644_8799.t39 vdd.t139 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 vdd.t194 a_n5644_8799.t40 CSoutput.t67 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X87 gnd.t131 commonsourceibias.t102 CSoutput.t140 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 CSoutput.t66 a_n5644_8799.t41 vdd.t123 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X89 CSoutput.t65 a_n5644_8799.t42 vdd.t124 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X90 a_n2903_n3924.t17 minus.t8 a_n1986_13878.t11 gnd.t325 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X91 CSoutput.t148 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X92 vdd.t115 a_n5644_8799.t43 CSoutput.t64 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X93 a_n2903_n3924.t33 plus.t9 a_n5644_8799.t27 gnd.t328 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X94 gnd.t130 commonsourceibias.t8 commonsourceibias.t9 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X95 gnd.t129 commonsourceibias.t103 CSoutput.t93 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X96 output.t16 CSoutput.t149 vdd.t95 gnd.t343 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X97 a_n2903_n3924.t4 diffpairibias.t17 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X98 vdd.t102 a_n5644_8799.t44 CSoutput.t63 vdd.t101 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X99 a_n5644_8799.t23 a_n1986_13878.t43 a_n1986_8322.t19 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X100 a_n1986_13878.t39 a_n1986_13878.t38 a_n1808_13878.t16 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X101 a_n2903_n3924.t32 plus.t10 a_n5644_8799.t6 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X102 gnd.t128 commonsourceibias.t104 CSoutput.t7 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X103 gnd.t296 gnd.t294 gnd.t295 gnd.t218 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X104 a_n1986_13878.t17 a_n1986_13878.t16 a_n1808_13878.t15 vdd.t149 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X105 vdd.t198 a_n5644_8799.t45 CSoutput.t62 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X106 gnd.t293 gnd.t291 gnd.t292 gnd.t218 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X107 CSoutput.t126 commonsourceibias.t105 gnd.t127 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 vdd.t79 vdd.t77 vdd.t78 vdd.t32 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X109 gnd.t126 commonsourceibias.t106 CSoutput.t96 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X110 vdd.t116 a_n5644_8799.t46 CSoutput.t61 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X111 vdd.t76 vdd.t74 vdd.t75 vdd.t61 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X112 gnd.t125 commonsourceibias.t107 CSoutput.t127 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X113 output.t15 CSoutput.t150 vdd.t92 gnd.t342 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X114 gnd.t124 commonsourceibias.t62 commonsourceibias.t63 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X115 vdd.t73 vdd.t70 vdd.t72 vdd.t71 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X116 output.t19 outputibias.t9 gnd.t347 gnd.t346 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X117 vdd.t69 vdd.t67 vdd.t68 vdd.t57 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X118 vdd.t66 vdd.t64 vdd.t65 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X119 CSoutput.t151 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X120 a_n1986_8322.t9 a_n1986_13878.t44 vdd.t185 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X121 vdd.t183 a_n1986_13878.t45 a_n1986_8322.t8 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X122 gnd.t290 gnd.t288 minus.t3 gnd.t289 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X123 CSoutput.t60 a_n5644_8799.t47 vdd.t191 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X124 CSoutput.t108 commonsourceibias.t108 gnd.t123 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X125 gnd.t122 commonsourceibias.t109 CSoutput.t143 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X126 CSoutput.t114 commonsourceibias.t110 gnd.t121 gnd.t108 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X127 gnd.t120 commonsourceibias.t111 CSoutput.t109 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X128 vdd.t93 CSoutput.t152 output.t14 gnd.t341 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X129 output.t13 CSoutput.t153 vdd.t4 gnd.t340 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X130 a_n2903_n3924.t3 diffpairibias.t18 gnd.t183 gnd.t182 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X131 gnd.t119 commonsourceibias.t112 CSoutput.t87 gnd.t73 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X132 gnd.t118 commonsourceibias.t50 commonsourceibias.t51 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 vdd.t11 a_n5644_8799.t48 CSoutput.t59 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X134 CSoutput.t8 commonsourceibias.t113 gnd.t117 gnd.t103 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X135 gnd.t274 gnd.t272 gnd.t273 gnd.t236 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X136 CSoutput.t154 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X137 vdd.t181 a_n1986_13878.t46 a_n1808_13878.t2 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X138 vdd.t63 vdd.t60 vdd.t62 vdd.t61 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X139 vdd.t59 vdd.t56 vdd.t58 vdd.t57 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X140 vdd.t112 a_n5644_8799.t49 CSoutput.t58 vdd.t101 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X141 gnd.t287 gnd.t285 gnd.t286 gnd.t218 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X142 a_n5644_8799.t15 a_n1986_13878.t47 a_n1986_8322.t18 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X143 a_n1986_8322.t7 a_n1986_13878.t48 vdd.t179 vdd.t178 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X144 vdd.t55 vdd.t52 vdd.t54 vdd.t53 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X145 a_n5644_8799.t8 plus.t11 a_n2903_n3924.t31 gnd.t320 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X146 a_n1986_13878.t27 a_n1986_13878.t26 a_n1808_13878.t14 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X147 a_n5644_8799.t4 plus.t12 a_n2903_n3924.t30 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X148 diffpairibias.t11 diffpairibias.t10 gnd.t198 gnd.t197 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X149 a_n5644_8799.t25 a_n1986_13878.t49 a_n1986_8322.t17 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X150 CSoutput.t115 commonsourceibias.t114 gnd.t116 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X151 a_n1808_13878.t13 a_n1986_13878.t24 a_n1986_13878.t25 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X152 gnd.t284 gnd.t282 gnd.t283 gnd.t200 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X153 gnd.t115 commonsourceibias.t115 CSoutput.t31 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X154 output.t12 CSoutput.t155 vdd.t5 gnd.t339 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X155 commonsourceibias.t49 commonsourceibias.t48 gnd.t114 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X156 CSoutput.t128 commonsourceibias.t116 gnd.t113 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X157 gnd.t281 gnd.t278 gnd.t280 gnd.t279 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X158 vdd.t175 a_n1986_13878.t50 a_n1986_8322.t6 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X159 gnd.t271 gnd.t269 gnd.t270 gnd.t226 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X160 CSoutput.t141 commonsourceibias.t117 gnd.t112 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 output.t11 CSoutput.t156 vdd.t126 gnd.t338 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X162 vdd.t51 vdd.t49 vdd.t50 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X163 gnd.t111 commonsourceibias.t118 CSoutput.t129 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X164 gnd.t110 commonsourceibias.t119 CSoutput.t97 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 a_n2903_n3924.t29 plus.t13 a_n5644_8799.t1 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X166 a_n1986_13878.t3 minus.t9 a_n2903_n3924.t9 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X167 outputibias.t7 outputibias.t6 gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X168 commonsourceibias.t47 commonsourceibias.t46 gnd.t109 gnd.t108 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 CSoutput.t57 a_n5644_8799.t50 vdd.t114 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X170 vdd.t104 a_n5644_8799.t51 CSoutput.t56 vdd.t103 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X171 plus.t3 gnd.t275 gnd.t277 gnd.t276 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X172 gnd.t107 commonsourceibias.t120 CSoutput.t142 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X173 outputibias.t5 outputibias.t4 gnd.t357 gnd.t356 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X174 CSoutput.t130 commonsourceibias.t121 gnd.t105 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X175 gnd.t268 gnd.t266 minus.t2 gnd.t267 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X176 gnd.t265 gnd.t262 gnd.t264 gnd.t263 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X177 a_n2903_n3924.t1 diffpairibias.t19 gnd.t176 gnd.t175 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X178 a_n5644_8799.t0 plus.t14 a_n2903_n3924.t28 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X179 a_n2903_n3924.t0 diffpairibias.t20 gnd.t10 gnd.t9 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X180 commonsourceibias.t43 commonsourceibias.t42 gnd.t104 gnd.t103 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X181 vdd.t197 a_n5644_8799.t52 CSoutput.t55 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X182 gnd.t261 gnd.t259 gnd.t260 gnd.t240 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X183 gnd.t258 gnd.t256 gnd.t257 gnd.t226 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X184 a_n5644_8799.t7 plus.t15 a_n2903_n3924.t27 gnd.t319 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X185 CSoutput.t9 commonsourceibias.t122 gnd.t102 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X186 vdd.t127 CSoutput.t157 output.t10 gnd.t337 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X187 CSoutput.t29 commonsourceibias.t123 gnd.t101 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 CSoutput.t54 a_n5644_8799.t53 vdd.t144 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X189 commonsourceibias.t41 commonsourceibias.t40 gnd.t100 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X190 a_n1808_13878.t4 a_n1986_13878.t51 vdd.t173 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X191 vdd.t128 CSoutput.t158 output.t9 gnd.t336 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X192 gnd.t99 commonsourceibias.t38 commonsourceibias.t39 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 diffpairibias.t9 diffpairibias.t8 gnd.t355 gnd.t354 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X194 vdd.t48 vdd.t46 vdd.t47 vdd.t28 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X195 vdd.t171 a_n1986_13878.t52 a_n1808_13878.t3 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X196 CSoutput.t102 commonsourceibias.t124 gnd.t97 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X197 CSoutput.t88 commonsourceibias.t125 gnd.t96 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X198 a_n1986_13878.t2 minus.t10 a_n2903_n3924.t8 gnd.t326 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X199 a_n2903_n3924.t26 plus.t16 a_n5644_8799.t26 gnd.t327 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X200 gnd.t95 commonsourceibias.t36 commonsourceibias.t37 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 vdd.t45 vdd.t42 vdd.t44 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X202 commonsourceibias.t35 commonsourceibias.t34 gnd.t93 gnd.t92 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 outputibias.t3 outputibias.t2 gnd.t187 gnd.t186 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X204 CSoutput.t53 a_n5644_8799.t54 vdd.t143 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X205 vdd.t142 a_n5644_8799.t55 CSoutput.t52 vdd.t103 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X206 gnd.t91 commonsourceibias.t126 CSoutput.t30 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 commonsourceibias.t59 commonsourceibias.t58 gnd.t90 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X208 a_n1986_8322.t16 a_n1986_13878.t53 a_n5644_8799.t19 vdd.t145 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X209 a_n2903_n3924.t16 minus.t11 a_n1986_13878.t10 gnd.t322 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X210 gnd.t87 commonsourceibias.t54 commonsourceibias.t55 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X211 CSoutput.t51 a_n5644_8799.t56 vdd.t192 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X212 diffpairibias.t7 diffpairibias.t6 gnd.t180 gnd.t179 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X213 CSoutput.t131 commonsourceibias.t127 gnd.t89 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X214 commonsourceibias.t57 commonsourceibias.t56 gnd.t88 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 vdd.t136 a_n5644_8799.t57 CSoutput.t50 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X216 vdd.t166 a_n1986_13878.t54 a_n1986_8322.t5 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X217 vdd.t135 a_n5644_8799.t58 CSoutput.t49 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X218 gnd.t255 gnd.t253 minus.t1 gnd.t254 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X219 plus.t2 gnd.t250 gnd.t252 gnd.t251 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X220 gnd.t86 commonsourceibias.t128 CSoutput.t89 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X221 a_n1808_13878.t6 a_n1986_13878.t55 vdd.t169 vdd.t168 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X222 CSoutput.t90 commonsourceibias.t129 gnd.t85 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X223 gnd.t84 commonsourceibias.t52 commonsourceibias.t53 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X224 output.t8 CSoutput.t159 vdd.t129 gnd.t335 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X225 CSoutput.t48 a_n5644_8799.t59 vdd.t15 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X226 CSoutput.t47 a_n5644_8799.t60 vdd.t106 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X227 gnd.t82 commonsourceibias.t130 CSoutput.t103 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X228 vdd.t41 vdd.t39 vdd.t40 vdd.t28 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X229 gnd.t249 gnd.t246 gnd.t248 gnd.t247 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X230 a_n1986_8322.t15 a_n1986_13878.t56 a_n5644_8799.t20 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X231 vdd.t164 a_n1986_13878.t57 a_n1986_8322.t4 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X232 CSoutput.t46 a_n5644_8799.t61 vdd.t196 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X233 a_n2903_n3924.t39 diffpairibias.t21 gnd.t353 gnd.t352 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X234 vdd.t195 a_n5644_8799.t62 CSoutput.t45 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X235 a_n5644_8799.t5 plus.t17 a_n2903_n3924.t25 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X236 a_n1986_13878.t5 minus.t12 a_n2903_n3924.t11 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X237 gnd.t81 commonsourceibias.t4 commonsourceibias.t5 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X238 a_n2903_n3924.t15 minus.t13 a_n1986_13878.t9 gnd.t328 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X239 gnd.t245 gnd.t243 gnd.t244 gnd.t222 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X240 output.t0 outputibias.t10 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X241 vdd.t38 vdd.t35 vdd.t37 vdd.t36 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X242 vdd.t34 vdd.t31 vdd.t33 vdd.t32 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X243 a_n2903_n3924.t14 minus.t14 a_n1986_13878.t8 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X244 CSoutput.t10 commonsourceibias.t131 gnd.t80 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X245 gnd.t79 commonsourceibias.t2 commonsourceibias.t3 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 gnd.t234 gnd.t232 gnd.t233 gnd.t222 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X247 a_n1808_13878.t12 a_n1986_13878.t18 a_n1986_13878.t19 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X248 a_n2903_n3924.t18 minus.t15 a_n1986_13878.t12 gnd.t329 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X249 CSoutput.t23 commonsourceibias.t132 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X250 vdd.t130 CSoutput.t160 output.t7 gnd.t334 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X251 output.t1 outputibias.t11 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X252 a_n1986_8322.t14 a_n1986_13878.t58 a_n5644_8799.t18 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X253 diffpairibias.t5 diffpairibias.t4 gnd.t185 gnd.t184 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X254 gnd.t242 gnd.t239 gnd.t241 gnd.t240 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X255 CSoutput.t16 commonsourceibias.t133 gnd.t76 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X256 output.t6 CSoutput.t161 vdd.t131 gnd.t333 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X257 gnd.t74 commonsourceibias.t14 commonsourceibias.t15 gnd.t73 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X258 CSoutput.t44 a_n5644_8799.t63 vdd.t133 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X259 a_n1986_8322.t3 a_n1986_13878.t59 vdd.t161 vdd.t160 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X260 a_n2903_n3924.t21 minus.t16 a_n1986_13878.t15 gnd.t321 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X261 gnd.t72 commonsourceibias.t134 CSoutput.t121 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X262 vdd.t159 a_n1986_13878.t60 a_n1808_13878.t0 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X263 vdd.t30 vdd.t27 vdd.t29 vdd.t28 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X264 gnd.t238 gnd.t235 gnd.t237 gnd.t236 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X265 gnd.t231 gnd.t229 plus.t1 gnd.t230 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X266 gnd.t71 commonsourceibias.t135 CSoutput.t119 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X267 gnd.t70 commonsourceibias.t136 CSoutput.t111 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X268 vdd.t26 vdd.t24 vdd.t25 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X269 a_n5644_8799.t22 a_n1986_13878.t61 a_n1986_8322.t13 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X270 a_n1986_8322.t12 a_n1986_13878.t62 a_n5644_8799.t14 vdd.t152 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X271 CSoutput.t43 a_n5644_8799.t64 vdd.t141 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X272 vdd.t98 CSoutput.t162 output.t5 gnd.t332 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X273 output.t4 CSoutput.t163 vdd.t99 gnd.t331 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X274 commonsourceibias.t13 commonsourceibias.t12 gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 a_n1808_13878.t7 a_n1986_13878.t63 vdd.t156 vdd.t155 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X276 vdd.t7 a_n5644_8799.t65 CSoutput.t42 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X277 gnd.t67 commonsourceibias.t137 CSoutput.t2 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 commonsourceibias.t11 commonsourceibias.t10 gnd.t66 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X279 gnd.t228 gnd.t225 gnd.t227 gnd.t226 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X280 a_n2903_n3924.t24 plus.t18 a_n5644_8799.t11 gnd.t325 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X281 gnd.t64 commonsourceibias.t138 CSoutput.t12 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X282 a_n1986_13878.t7 minus.t17 a_n2903_n3924.t13 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X283 commonsourceibias.t25 commonsourceibias.t24 gnd.t62 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X284 CSoutput.t20 commonsourceibias.t139 gnd.t63 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X285 gnd.t60 commonsourceibias.t140 CSoutput.t110 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 gnd.t58 commonsourceibias.t22 commonsourceibias.t23 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 CSoutput.t41 a_n5644_8799.t66 vdd.t137 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 a_n1808_13878.t11 a_n1986_13878.t30 a_n1986_13878.t31 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X289 gnd.t224 gnd.t221 gnd.t223 gnd.t222 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X290 gnd.t56 commonsourceibias.t20 commonsourceibias.t21 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X291 commonsourceibias.t7 commonsourceibias.t6 gnd.t55 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 CSoutput.t40 a_n5644_8799.t67 vdd.t140 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 gnd.t53 commonsourceibias.t141 CSoutput.t94 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X294 vdd.t120 a_n5644_8799.t68 CSoutput.t39 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X295 a_n2903_n3924.t12 minus.t18 a_n1986_13878.t6 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X296 gnd.t52 commonsourceibias.t142 CSoutput.t95 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X297 CSoutput.t21 commonsourceibias.t143 gnd.t50 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X298 gnd.t49 commonsourceibias.t144 CSoutput.t112 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X299 a_n2903_n3924.t5 diffpairibias.t22 gnd.t196 gnd.t195 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X300 a_n5644_8799.t17 a_n1986_13878.t64 a_n1986_8322.t11 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X301 a_n1986_13878.t29 a_n1986_13878.t28 a_n1808_13878.t10 vdd.t152 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X302 gnd.t220 gnd.t217 gnd.t219 gnd.t218 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X303 CSoutput.t113 commonsourceibias.t145 gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X304 vdd.t100 CSoutput.t164 output.t3 gnd.t330 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X305 vdd.t1 a_n5644_8799.t69 CSoutput.t38 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X306 CSoutput.t120 commonsourceibias.t146 gnd.t45 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 gnd.t44 commonsourceibias.t147 CSoutput.t116 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X308 commonsourceibias.t27 commonsourceibias.t26 gnd.t42 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X309 vdd.t23 vdd.t20 vdd.t22 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X310 minus.t0 gnd.t214 gnd.t216 gnd.t215 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X311 gnd.t213 gnd.t211 plus.t0 gnd.t212 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X312 CSoutput.t165 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X313 diffpairibias.t3 diffpairibias.t2 gnd.t351 gnd.t350 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X314 gnd.t40 commonsourceibias.t148 CSoutput.t13 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 a_n1986_13878.t14 minus.t19 a_n2903_n3924.t20 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X316 gnd.t210 gnd.t207 gnd.t209 gnd.t208 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X317 gnd.t39 commonsourceibias.t149 CSoutput.t4 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X318 diffpairibias.t1 diffpairibias.t0 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X319 CSoutput.t83 commonsourceibias.t150 gnd.t37 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X320 gnd.t35 commonsourceibias.t151 CSoutput.t84 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X321 commonsourceibias.t33 commonsourceibias.t32 gnd.t34 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X322 vdd.t151 a_n1986_13878.t65 a_n1808_13878.t1 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X323 CSoutput.t37 a_n5644_8799.t70 vdd.t97 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X324 gnd.t33 commonsourceibias.t30 commonsourceibias.t31 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X325 gnd.t31 commonsourceibias.t152 CSoutput.t18 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 a_n5644_8799.t13 plus.t19 a_n2903_n3924.t23 gnd.t326 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X327 CSoutput.t36 a_n5644_8799.t71 vdd.t134 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X328 a_n1986_8322.t10 a_n1986_13878.t66 a_n5644_8799.t16 vdd.t149 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X329 a_n1986_13878.t13 minus.t20 a_n2903_n3924.t19 gnd.t320 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X330 gnd.t29 commonsourceibias.t153 CSoutput.t19 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X331 gnd.t27 commonsourceibias.t154 CSoutput.t3 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X332 commonsourceibias.t19 commonsourceibias.t18 gnd.t25 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X333 gnd.t206 gnd.t203 gnd.t205 gnd.t204 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X334 vdd.t108 a_n5644_8799.t72 CSoutput.t35 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X335 CSoutput.t34 a_n5644_8799.t73 vdd.t3 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X336 vdd.t132 a_n5644_8799.t74 CSoutput.t33 vdd.t103 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X337 gnd.t23 commonsourceibias.t155 CSoutput.t14 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X338 a_n1986_8322.t2 a_n1986_13878.t67 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X339 a_n1808_13878.t9 a_n1986_13878.t36 a_n1986_13878.t37 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X340 gnd.t22 commonsourceibias.t156 CSoutput.t17 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X341 gnd.t202 gnd.t199 gnd.t201 gnd.t200 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X342 vdd.t199 a_n5644_8799.t75 CSoutput.t32 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X343 CSoutput.t11 commonsourceibias.t157 gnd.t20 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X344 gnd.t18 commonsourceibias.t158 CSoutput.t24 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X345 CSoutput.t15 commonsourceibias.t159 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X346 a_n2903_n3924.t22 plus.t20 a_n5644_8799.t10 gnd.t322 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X347 outputibias.t1 outputibias.t0 gnd.t359 gnd.t358 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X348 commonsourceibias.t17 commonsourceibias.t16 gnd.t14 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X349 a_n1986_13878.t23 a_n1986_13878.t22 a_n1808_13878.t8 vdd.t145 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X350 vdd.t19 vdd.t16 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X351 a_n2903_n3924.t38 diffpairibias.t23 gnd.t349 gnd.t348 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
R0 a_n1986_13878.n6 a_n1986_13878.t66 539.01
R1 a_n1986_13878.n64 a_n1986_13878.t49 512.366
R2 a_n1986_13878.n63 a_n1986_13878.t53 512.366
R3 a_n1986_13878.n61 a_n1986_13878.t43 512.366
R4 a_n1986_13878.n62 a_n1986_13878.t58 512.366
R5 a_n1986_13878.n49 a_n1986_13878.t36 533.058
R6 a_n1986_13878.n8 a_n1986_13878.t28 539.01
R7 a_n1986_13878.n67 a_n1986_13878.t18 512.366
R8 a_n1986_13878.n66 a_n1986_13878.t38 512.366
R9 a_n1986_13878.n52 a_n1986_13878.t30 512.366
R10 a_n1986_13878.n65 a_n1986_13878.t26 512.366
R11 a_n1986_13878.n20 a_n1986_13878.t16 539.01
R12 a_n1986_13878.n88 a_n1986_13878.t34 512.366
R13 a_n1986_13878.n89 a_n1986_13878.t22 512.366
R14 a_n1986_13878.n50 a_n1986_13878.t24 512.366
R15 a_n1986_13878.n90 a_n1986_13878.t20 512.366
R16 a_n1986_13878.n24 a_n1986_13878.t62 539.01
R17 a_n1986_13878.n85 a_n1986_13878.t61 512.366
R18 a_n1986_13878.n86 a_n1986_13878.t41 512.366
R19 a_n1986_13878.n51 a_n1986_13878.t47 512.366
R20 a_n1986_13878.n87 a_n1986_13878.t56 512.366
R21 a_n1986_13878.n77 a_n1986_13878.t55 512.366
R22 a_n1986_13878.n76 a_n1986_13878.t46 512.366
R23 a_n1986_13878.n75 a_n1986_13878.t40 512.366
R24 a_n1986_13878.n79 a_n1986_13878.t63 512.366
R25 a_n1986_13878.n78 a_n1986_13878.t52 512.366
R26 a_n1986_13878.n74 a_n1986_13878.t51 512.366
R27 a_n1986_13878.n81 a_n1986_13878.t59 512.366
R28 a_n1986_13878.n80 a_n1986_13878.t45 512.366
R29 a_n1986_13878.n73 a_n1986_13878.t44 512.366
R30 a_n1986_13878.n83 a_n1986_13878.t48 512.366
R31 a_n1986_13878.n82 a_n1986_13878.t57 512.366
R32 a_n1986_13878.n72 a_n1986_13878.t67 512.366
R33 a_n1986_13878.n48 a_n1986_13878.n4 70.3058
R34 a_n1986_13878.n17 a_n1986_13878.n33 70.3058
R35 a_n1986_13878.n21 a_n1986_13878.n30 70.3058
R36 a_n1986_13878.n29 a_n1986_13878.n22 70.1674
R37 a_n1986_13878.n29 a_n1986_13878.n51 20.9683
R38 a_n1986_13878.n22 a_n1986_13878.n28 75.0448
R39 a_n1986_13878.n86 a_n1986_13878.n28 11.2134
R40 a_n1986_13878.n23 a_n1986_13878.n24 44.8194
R41 a_n1986_13878.n32 a_n1986_13878.n18 70.1674
R42 a_n1986_13878.n32 a_n1986_13878.n50 20.9683
R43 a_n1986_13878.n18 a_n1986_13878.n31 75.0448
R44 a_n1986_13878.n89 a_n1986_13878.n31 11.2134
R45 a_n1986_13878.n19 a_n1986_13878.n20 44.8194
R46 a_n1986_13878.n9 a_n1986_13878.n42 70.1674
R47 a_n1986_13878.n11 a_n1986_13878.n39 70.1674
R48 a_n1986_13878.n13 a_n1986_13878.n37 70.1674
R49 a_n1986_13878.n15 a_n1986_13878.n35 70.1674
R50 a_n1986_13878.n35 a_n1986_13878.n72 20.9683
R51 a_n1986_13878.n34 a_n1986_13878.n16 75.0448
R52 a_n1986_13878.n82 a_n1986_13878.n34 11.2134
R53 a_n1986_13878.n16 a_n1986_13878.n83 161.3
R54 a_n1986_13878.n37 a_n1986_13878.n73 20.9683
R55 a_n1986_13878.n36 a_n1986_13878.n14 75.0448
R56 a_n1986_13878.n80 a_n1986_13878.n36 11.2134
R57 a_n1986_13878.n14 a_n1986_13878.n81 161.3
R58 a_n1986_13878.n39 a_n1986_13878.n74 20.9683
R59 a_n1986_13878.n38 a_n1986_13878.n12 75.0448
R60 a_n1986_13878.n78 a_n1986_13878.n38 11.2134
R61 a_n1986_13878.n12 a_n1986_13878.n79 161.3
R62 a_n1986_13878.n42 a_n1986_13878.n75 20.9683
R63 a_n1986_13878.n40 a_n1986_13878.n10 75.0448
R64 a_n1986_13878.n76 a_n1986_13878.n40 11.2134
R65 a_n1986_13878.n10 a_n1986_13878.n77 161.3
R66 a_n1986_13878.n27 a_n1986_13878.n45 70.1674
R67 a_n1986_13878.n45 a_n1986_13878.n52 20.9683
R68 a_n1986_13878.n44 a_n1986_13878.n43 75.0448
R69 a_n1986_13878.n66 a_n1986_13878.n44 11.2134
R70 a_n1986_13878.n7 a_n1986_13878.n8 44.8194
R71 a_n1986_13878.n49 a_n1986_13878.n27 70.3058
R72 a_n1986_13878.n5 a_n1986_13878.n47 70.1674
R73 a_n1986_13878.n47 a_n1986_13878.n61 20.9683
R74 a_n1986_13878.n46 a_n1986_13878.n5 75.0448
R75 a_n1986_13878.n63 a_n1986_13878.n46 11.2134
R76 a_n1986_13878.n3 a_n1986_13878.n6 44.8194
R77 a_n1986_13878.n1 a_n1986_13878.n59 81.4626
R78 a_n1986_13878.n2 a_n1986_13878.n55 81.4626
R79 a_n1986_13878.n2 a_n1986_13878.n53 81.4626
R80 a_n1986_13878.n1 a_n1986_13878.n60 80.9324
R81 a_n1986_13878.n1 a_n1986_13878.n58 80.9324
R82 a_n1986_13878.n0 a_n1986_13878.n57 80.9324
R83 a_n1986_13878.n2 a_n1986_13878.n56 80.9324
R84 a_n1986_13878.n2 a_n1986_13878.n54 80.9324
R85 a_n1986_13878.n25 a_n1986_13878.t37 74.6477
R86 a_n1986_13878.t17 a_n1986_13878.n94 74.6477
R87 a_n1986_13878.n70 a_n1986_13878.t29 74.2899
R88 a_n1986_13878.n26 a_n1986_13878.t33 74.2897
R89 a_n1986_13878.n26 a_n1986_13878.n92 70.6783
R90 a_n1986_13878.n94 a_n1986_13878.n93 70.6783
R91 a_n1986_13878.n25 a_n1986_13878.n68 70.6783
R92 a_n1986_13878.n25 a_n1986_13878.n69 70.6783
R93 a_n1986_13878.n64 a_n1986_13878.n63 48.2005
R94 a_n1986_13878.n62 a_n1986_13878.n47 20.9683
R95 a_n1986_13878.n67 a_n1986_13878.n66 48.2005
R96 a_n1986_13878.n65 a_n1986_13878.n45 20.9683
R97 a_n1986_13878.n89 a_n1986_13878.n88 48.2005
R98 a_n1986_13878.n90 a_n1986_13878.n32 20.9683
R99 a_n1986_13878.n86 a_n1986_13878.n85 48.2005
R100 a_n1986_13878.n87 a_n1986_13878.n29 20.9683
R101 a_n1986_13878.n77 a_n1986_13878.n76 48.2005
R102 a_n1986_13878.t60 a_n1986_13878.n42 533.335
R103 a_n1986_13878.n79 a_n1986_13878.n78 48.2005
R104 a_n1986_13878.t65 a_n1986_13878.n39 533.335
R105 a_n1986_13878.n81 a_n1986_13878.n80 48.2005
R106 a_n1986_13878.t54 a_n1986_13878.n37 533.335
R107 a_n1986_13878.n83 a_n1986_13878.n82 48.2005
R108 a_n1986_13878.t50 a_n1986_13878.n35 533.335
R109 a_n1986_13878.n48 a_n1986_13878.t64 533.058
R110 a_n1986_13878.t32 a_n1986_13878.n33 533.058
R111 a_n1986_13878.t42 a_n1986_13878.n30 533.058
R112 a_n1986_13878.n46 a_n1986_13878.n61 35.3134
R113 a_n1986_13878.n44 a_n1986_13878.n52 35.3134
R114 a_n1986_13878.n50 a_n1986_13878.n31 35.3134
R115 a_n1986_13878.n51 a_n1986_13878.n28 35.3134
R116 a_n1986_13878.n40 a_n1986_13878.n75 35.3134
R117 a_n1986_13878.n38 a_n1986_13878.n74 35.3134
R118 a_n1986_13878.n36 a_n1986_13878.n73 35.3134
R119 a_n1986_13878.n34 a_n1986_13878.n72 35.3134
R120 a_n1986_13878.n0 a_n1986_13878.n2 32.5247
R121 a_n1986_13878.n27 a_n1986_13878.n1 23.891
R122 a_n1986_13878.n23 a_n1986_13878.n84 12.046
R123 a_n1986_13878.n4 a_n1986_13878.n41 11.8414
R124 a_n1986_13878.n71 a_n1986_13878.n7 10.5365
R125 a_n1986_13878.n26 a_n1986_13878.n91 9.50122
R126 a_n1986_13878.n9 a_n1986_13878.n41 7.47588
R127 a_n1986_13878.n84 a_n1986_13878.n16 7.47588
R128 a_n1986_13878.n91 a_n1986_13878.n17 6.70126
R129 a_n1986_13878.n71 a_n1986_13878.n70 5.65783
R130 a_n1986_13878.n91 a_n1986_13878.n41 5.3452
R131 a_n1986_13878.n19 a_n1986_13878.n21 3.95126
R132 a_n1986_13878.n27 a_n1986_13878.n3 3.95126
R133 a_n1986_13878.n92 a_n1986_13878.t25 3.61217
R134 a_n1986_13878.n92 a_n1986_13878.t21 3.61217
R135 a_n1986_13878.n93 a_n1986_13878.t35 3.61217
R136 a_n1986_13878.n93 a_n1986_13878.t23 3.61217
R137 a_n1986_13878.n68 a_n1986_13878.t31 3.61217
R138 a_n1986_13878.n68 a_n1986_13878.t27 3.61217
R139 a_n1986_13878.n69 a_n1986_13878.t19 3.61217
R140 a_n1986_13878.n69 a_n1986_13878.t39 3.61217
R141 a_n1986_13878.n59 a_n1986_13878.t15 2.82907
R142 a_n1986_13878.n59 a_n1986_13878.t13 2.82907
R143 a_n1986_13878.n60 a_n1986_13878.t10 2.82907
R144 a_n1986_13878.n60 a_n1986_13878.t2 2.82907
R145 a_n1986_13878.n58 a_n1986_13878.t4 2.82907
R146 a_n1986_13878.n58 a_n1986_13878.t0 2.82907
R147 a_n1986_13878.n57 a_n1986_13878.t12 2.82907
R148 a_n1986_13878.n57 a_n1986_13878.t5 2.82907
R149 a_n1986_13878.n55 a_n1986_13878.t8 2.82907
R150 a_n1986_13878.n55 a_n1986_13878.t7 2.82907
R151 a_n1986_13878.n56 a_n1986_13878.t6 2.82907
R152 a_n1986_13878.n56 a_n1986_13878.t14 2.82907
R153 a_n1986_13878.n54 a_n1986_13878.t11 2.82907
R154 a_n1986_13878.n54 a_n1986_13878.t1 2.82907
R155 a_n1986_13878.n53 a_n1986_13878.t9 2.82907
R156 a_n1986_13878.n53 a_n1986_13878.t3 2.82907
R157 a_n1986_13878.n84 a_n1986_13878.n71 1.30542
R158 a_n1986_13878.n13 a_n1986_13878.n12 1.04595
R159 a_n1986_13878.n6 a_n1986_13878.n64 13.657
R160 a_n1986_13878.n62 a_n1986_13878.n48 21.4216
R161 a_n1986_13878.n8 a_n1986_13878.n67 13.657
R162 a_n1986_13878.n65 a_n1986_13878.n49 21.4216
R163 a_n1986_13878.n88 a_n1986_13878.n20 13.657
R164 a_n1986_13878.n33 a_n1986_13878.n90 21.4216
R165 a_n1986_13878.n85 a_n1986_13878.n24 13.657
R166 a_n1986_13878.n30 a_n1986_13878.n87 21.4216
R167 a_n1986_13878.n1 a_n1986_13878.n0 1.06084
R168 a_n1986_13878.n23 a_n1986_13878.n22 0.758076
R169 a_n1986_13878.n22 a_n1986_13878.n21 0.758076
R170 a_n1986_13878.n19 a_n1986_13878.n18 0.758076
R171 a_n1986_13878.n18 a_n1986_13878.n17 0.758076
R172 a_n1986_13878.n16 a_n1986_13878.n15 0.758076
R173 a_n1986_13878.n14 a_n1986_13878.n13 0.758076
R174 a_n1986_13878.n12 a_n1986_13878.n11 0.758076
R175 a_n1986_13878.n10 a_n1986_13878.n9 0.758076
R176 a_n1986_13878.n43 a_n1986_13878.n7 0.758076
R177 a_n1986_13878.n5 a_n1986_13878.n3 0.758076
R178 a_n1986_13878.n5 a_n1986_13878.n4 0.758076
R179 a_n1986_13878.n43 a_n1986_13878.n27 0.720197
R180 a_n1986_13878.n94 a_n1986_13878.n26 0.716017
R181 a_n1986_13878.n70 a_n1986_13878.n25 0.716017
R182 a_n1986_13878.n15 a_n1986_13878.n14 0.67853
R183 a_n1986_13878.n11 a_n1986_13878.n10 0.67853
R184 a_n1808_13878.n2 a_n1808_13878.n0 98.9633
R185 a_n1808_13878.n5 a_n1808_13878.n3 98.7517
R186 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R187 a_n1808_13878.n7 a_n1808_13878.n6 98.6055
R188 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R189 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R190 a_n1808_13878.n9 a_n1808_13878.t7 74.6477
R191 a_n1808_13878.n14 a_n1808_13878.t0 74.2899
R192 a_n1808_13878.n11 a_n1808_13878.t6 74.2899
R193 a_n1808_13878.n10 a_n1808_13878.t1 74.2899
R194 a_n1808_13878.n13 a_n1808_13878.n12 70.6783
R195 a_n1808_13878.n9 a_n1808_13878.n8 70.6783
R196 a_n1808_13878.n15 a_n1808_13878.n7 13.5694
R197 a_n1808_13878.n16 a_n1808_13878.n15 11.5762
R198 a_n1808_13878.n15 a_n1808_13878.n14 6.2408
R199 a_n1808_13878.n1 a_n1808_13878.t8 3.61217
R200 a_n1808_13878.n1 a_n1808_13878.t13 3.61217
R201 a_n1808_13878.n0 a_n1808_13878.t15 3.61217
R202 a_n1808_13878.n0 a_n1808_13878.t19 3.61217
R203 a_n1808_13878.n12 a_n1808_13878.t2 3.61217
R204 a_n1808_13878.n12 a_n1808_13878.t5 3.61217
R205 a_n1808_13878.n8 a_n1808_13878.t3 3.61217
R206 a_n1808_13878.n8 a_n1808_13878.t4 3.61217
R207 a_n1808_13878.n6 a_n1808_13878.t14 3.61217
R208 a_n1808_13878.n6 a_n1808_13878.t9 3.61217
R209 a_n1808_13878.n4 a_n1808_13878.t16 3.61217
R210 a_n1808_13878.n4 a_n1808_13878.t11 3.61217
R211 a_n1808_13878.n3 a_n1808_13878.t10 3.61217
R212 a_n1808_13878.n3 a_n1808_13878.t12 3.61217
R213 a_n1808_13878.n17 a_n1808_13878.t17 3.61217
R214 a_n1808_13878.t18 a_n1808_13878.n17 3.61217
R215 a_n1808_13878.n10 a_n1808_13878.n9 0.358259
R216 a_n1808_13878.n13 a_n1808_13878.n11 0.358259
R217 a_n1808_13878.n14 a_n1808_13878.n13 0.358259
R218 a_n1808_13878.n16 a_n1808_13878.n2 0.358259
R219 a_n1808_13878.n7 a_n1808_13878.n5 0.146627
R220 a_n1808_13878.n11 a_n1808_13878.n10 0.101793
R221 vdd.n291 vdd.n255 756.745
R222 vdd.n244 vdd.n208 756.745
R223 vdd.n201 vdd.n165 756.745
R224 vdd.n154 vdd.n118 756.745
R225 vdd.n112 vdd.n76 756.745
R226 vdd.n65 vdd.n29 756.745
R227 vdd.n1106 vdd.n1070 756.745
R228 vdd.n1153 vdd.n1117 756.745
R229 vdd.n1016 vdd.n980 756.745
R230 vdd.n1063 vdd.n1027 756.745
R231 vdd.n927 vdd.n891 756.745
R232 vdd.n974 vdd.n938 756.745
R233 vdd.n1791 vdd.t64 640.208
R234 vdd.n755 vdd.t52 640.208
R235 vdd.n1765 vdd.t16 640.208
R236 vdd.n747 vdd.t83 640.208
R237 vdd.n2536 vdd.t35 640.208
R238 vdd.n2256 vdd.t74 640.208
R239 vdd.n622 vdd.t56 640.208
R240 vdd.n2253 vdd.t60 640.208
R241 vdd.n589 vdd.t67 640.208
R242 vdd.n817 vdd.t70 640.208
R243 vdd.n1320 vdd.t31 592.009
R244 vdd.n1358 vdd.t77 592.009
R245 vdd.n1254 vdd.t80 592.009
R246 vdd.n1947 vdd.t27 592.009
R247 vdd.n1584 vdd.t39 592.009
R248 vdd.n1544 vdd.t46 592.009
R249 vdd.n2908 vdd.t89 592.009
R250 vdd.n405 vdd.t42 592.009
R251 vdd.n365 vdd.t49 592.009
R252 vdd.n557 vdd.t20 592.009
R253 vdd.n2804 vdd.t24 592.009
R254 vdd.n2711 vdd.t86 592.009
R255 vdd.n292 vdd.n291 585
R256 vdd.n290 vdd.n257 585
R257 vdd.n289 vdd.n288 585
R258 vdd.n260 vdd.n258 585
R259 vdd.n283 vdd.n282 585
R260 vdd.n281 vdd.n280 585
R261 vdd.n264 vdd.n263 585
R262 vdd.n275 vdd.n274 585
R263 vdd.n273 vdd.n272 585
R264 vdd.n268 vdd.n267 585
R265 vdd.n245 vdd.n244 585
R266 vdd.n243 vdd.n210 585
R267 vdd.n242 vdd.n241 585
R268 vdd.n213 vdd.n211 585
R269 vdd.n236 vdd.n235 585
R270 vdd.n234 vdd.n233 585
R271 vdd.n217 vdd.n216 585
R272 vdd.n228 vdd.n227 585
R273 vdd.n226 vdd.n225 585
R274 vdd.n221 vdd.n220 585
R275 vdd.n202 vdd.n201 585
R276 vdd.n200 vdd.n167 585
R277 vdd.n199 vdd.n198 585
R278 vdd.n170 vdd.n168 585
R279 vdd.n193 vdd.n192 585
R280 vdd.n191 vdd.n190 585
R281 vdd.n174 vdd.n173 585
R282 vdd.n185 vdd.n184 585
R283 vdd.n183 vdd.n182 585
R284 vdd.n178 vdd.n177 585
R285 vdd.n155 vdd.n154 585
R286 vdd.n153 vdd.n120 585
R287 vdd.n152 vdd.n151 585
R288 vdd.n123 vdd.n121 585
R289 vdd.n146 vdd.n145 585
R290 vdd.n144 vdd.n143 585
R291 vdd.n127 vdd.n126 585
R292 vdd.n138 vdd.n137 585
R293 vdd.n136 vdd.n135 585
R294 vdd.n131 vdd.n130 585
R295 vdd.n113 vdd.n112 585
R296 vdd.n111 vdd.n78 585
R297 vdd.n110 vdd.n109 585
R298 vdd.n81 vdd.n79 585
R299 vdd.n104 vdd.n103 585
R300 vdd.n102 vdd.n101 585
R301 vdd.n85 vdd.n84 585
R302 vdd.n96 vdd.n95 585
R303 vdd.n94 vdd.n93 585
R304 vdd.n89 vdd.n88 585
R305 vdd.n66 vdd.n65 585
R306 vdd.n64 vdd.n31 585
R307 vdd.n63 vdd.n62 585
R308 vdd.n34 vdd.n32 585
R309 vdd.n57 vdd.n56 585
R310 vdd.n55 vdd.n54 585
R311 vdd.n38 vdd.n37 585
R312 vdd.n49 vdd.n48 585
R313 vdd.n47 vdd.n46 585
R314 vdd.n42 vdd.n41 585
R315 vdd.n1107 vdd.n1106 585
R316 vdd.n1105 vdd.n1072 585
R317 vdd.n1104 vdd.n1103 585
R318 vdd.n1075 vdd.n1073 585
R319 vdd.n1098 vdd.n1097 585
R320 vdd.n1096 vdd.n1095 585
R321 vdd.n1079 vdd.n1078 585
R322 vdd.n1090 vdd.n1089 585
R323 vdd.n1088 vdd.n1087 585
R324 vdd.n1083 vdd.n1082 585
R325 vdd.n1154 vdd.n1153 585
R326 vdd.n1152 vdd.n1119 585
R327 vdd.n1151 vdd.n1150 585
R328 vdd.n1122 vdd.n1120 585
R329 vdd.n1145 vdd.n1144 585
R330 vdd.n1143 vdd.n1142 585
R331 vdd.n1126 vdd.n1125 585
R332 vdd.n1137 vdd.n1136 585
R333 vdd.n1135 vdd.n1134 585
R334 vdd.n1130 vdd.n1129 585
R335 vdd.n1017 vdd.n1016 585
R336 vdd.n1015 vdd.n982 585
R337 vdd.n1014 vdd.n1013 585
R338 vdd.n985 vdd.n983 585
R339 vdd.n1008 vdd.n1007 585
R340 vdd.n1006 vdd.n1005 585
R341 vdd.n989 vdd.n988 585
R342 vdd.n1000 vdd.n999 585
R343 vdd.n998 vdd.n997 585
R344 vdd.n993 vdd.n992 585
R345 vdd.n1064 vdd.n1063 585
R346 vdd.n1062 vdd.n1029 585
R347 vdd.n1061 vdd.n1060 585
R348 vdd.n1032 vdd.n1030 585
R349 vdd.n1055 vdd.n1054 585
R350 vdd.n1053 vdd.n1052 585
R351 vdd.n1036 vdd.n1035 585
R352 vdd.n1047 vdd.n1046 585
R353 vdd.n1045 vdd.n1044 585
R354 vdd.n1040 vdd.n1039 585
R355 vdd.n928 vdd.n927 585
R356 vdd.n926 vdd.n893 585
R357 vdd.n925 vdd.n924 585
R358 vdd.n896 vdd.n894 585
R359 vdd.n919 vdd.n918 585
R360 vdd.n917 vdd.n916 585
R361 vdd.n900 vdd.n899 585
R362 vdd.n911 vdd.n910 585
R363 vdd.n909 vdd.n908 585
R364 vdd.n904 vdd.n903 585
R365 vdd.n975 vdd.n974 585
R366 vdd.n973 vdd.n940 585
R367 vdd.n972 vdd.n971 585
R368 vdd.n943 vdd.n941 585
R369 vdd.n966 vdd.n965 585
R370 vdd.n964 vdd.n963 585
R371 vdd.n947 vdd.n946 585
R372 vdd.n958 vdd.n957 585
R373 vdd.n956 vdd.n955 585
R374 vdd.n951 vdd.n950 585
R375 vdd.n3024 vdd.n330 515.122
R376 vdd.n2906 vdd.n328 515.122
R377 vdd.n515 vdd.n478 515.122
R378 vdd.n2842 vdd.n479 515.122
R379 vdd.n1942 vdd.n865 515.122
R380 vdd.n1945 vdd.n1944 515.122
R381 vdd.n1227 vdd.n1191 515.122
R382 vdd.n1423 vdd.n1192 515.122
R383 vdd.n269 vdd.t15 329.043
R384 vdd.n222 vdd.t104 329.043
R385 vdd.n179 vdd.t133 329.043
R386 vdd.n132 vdd.t142 329.043
R387 vdd.n90 vdd.t111 329.043
R388 vdd.n43 vdd.t132 329.043
R389 vdd.n1084 vdd.t121 329.043
R390 vdd.n1131 vdd.t102 329.043
R391 vdd.n994 vdd.t138 329.043
R392 vdd.n1041 vdd.t112 329.043
R393 vdd.n905 vdd.t3 329.043
R394 vdd.n952 vdd.t193 329.043
R395 vdd.n1320 vdd.t34 319.788
R396 vdd.n1358 vdd.t79 319.788
R397 vdd.n1254 vdd.t82 319.788
R398 vdd.n1947 vdd.t29 319.788
R399 vdd.n1584 vdd.t40 319.788
R400 vdd.n1544 vdd.t47 319.788
R401 vdd.n2908 vdd.t90 319.788
R402 vdd.n405 vdd.t44 319.788
R403 vdd.n365 vdd.t50 319.788
R404 vdd.n557 vdd.t23 319.788
R405 vdd.n2804 vdd.t26 319.788
R406 vdd.n2711 vdd.t88 319.788
R407 vdd.n1321 vdd.t33 303.69
R408 vdd.n1359 vdd.t78 303.69
R409 vdd.n1255 vdd.t81 303.69
R410 vdd.n1948 vdd.t30 303.69
R411 vdd.n1585 vdd.t41 303.69
R412 vdd.n1545 vdd.t48 303.69
R413 vdd.n2909 vdd.t91 303.69
R414 vdd.n406 vdd.t45 303.69
R415 vdd.n366 vdd.t51 303.69
R416 vdd.n558 vdd.t22 303.69
R417 vdd.n2805 vdd.t25 303.69
R418 vdd.n2712 vdd.t87 303.69
R419 vdd.n2479 vdd.n703 297.074
R420 vdd.n2672 vdd.n599 297.074
R421 vdd.n2609 vdd.n596 297.074
R422 vdd.n2402 vdd.n704 297.074
R423 vdd.n2217 vdd.n744 297.074
R424 vdd.n2148 vdd.n2147 297.074
R425 vdd.n1894 vdd.n840 297.074
R426 vdd.n1990 vdd.n838 297.074
R427 vdd.n2588 vdd.n597 297.074
R428 vdd.n2675 vdd.n2674 297.074
R429 vdd.n2251 vdd.n705 297.074
R430 vdd.n2477 vdd.n706 297.074
R431 vdd.n2145 vdd.n753 297.074
R432 vdd.n751 vdd.n726 297.074
R433 vdd.n1831 vdd.n841 297.074
R434 vdd.n1988 vdd.n842 297.074
R435 vdd.n2590 vdd.n597 185
R436 vdd.n2673 vdd.n597 185
R437 vdd.n2592 vdd.n2591 185
R438 vdd.n2591 vdd.n595 185
R439 vdd.n2593 vdd.n629 185
R440 vdd.n2603 vdd.n629 185
R441 vdd.n2594 vdd.n638 185
R442 vdd.n638 vdd.n636 185
R443 vdd.n2596 vdd.n2595 185
R444 vdd.n2597 vdd.n2596 185
R445 vdd.n2549 vdd.n637 185
R446 vdd.n637 vdd.n633 185
R447 vdd.n2548 vdd.n2547 185
R448 vdd.n2547 vdd.n2546 185
R449 vdd.n640 vdd.n639 185
R450 vdd.n641 vdd.n640 185
R451 vdd.n2539 vdd.n2538 185
R452 vdd.n2540 vdd.n2539 185
R453 vdd.n2535 vdd.n650 185
R454 vdd.n650 vdd.n647 185
R455 vdd.n2534 vdd.n2533 185
R456 vdd.n2533 vdd.n2532 185
R457 vdd.n652 vdd.n651 185
R458 vdd.n660 vdd.n652 185
R459 vdd.n2525 vdd.n2524 185
R460 vdd.n2526 vdd.n2525 185
R461 vdd.n2523 vdd.n661 185
R462 vdd.n2374 vdd.n661 185
R463 vdd.n2522 vdd.n2521 185
R464 vdd.n2521 vdd.n2520 185
R465 vdd.n663 vdd.n662 185
R466 vdd.n664 vdd.n663 185
R467 vdd.n2513 vdd.n2512 185
R468 vdd.n2514 vdd.n2513 185
R469 vdd.n2511 vdd.n673 185
R470 vdd.n673 vdd.n670 185
R471 vdd.n2510 vdd.n2509 185
R472 vdd.n2509 vdd.n2508 185
R473 vdd.n675 vdd.n674 185
R474 vdd.n683 vdd.n675 185
R475 vdd.n2501 vdd.n2500 185
R476 vdd.n2502 vdd.n2501 185
R477 vdd.n2499 vdd.n684 185
R478 vdd.n690 vdd.n684 185
R479 vdd.n2498 vdd.n2497 185
R480 vdd.n2497 vdd.n2496 185
R481 vdd.n686 vdd.n685 185
R482 vdd.n687 vdd.n686 185
R483 vdd.n2489 vdd.n2488 185
R484 vdd.n2490 vdd.n2489 185
R485 vdd.n2487 vdd.n696 185
R486 vdd.n2395 vdd.n696 185
R487 vdd.n2486 vdd.n2485 185
R488 vdd.n2485 vdd.n2484 185
R489 vdd.n698 vdd.n697 185
R490 vdd.t172 vdd.n698 185
R491 vdd.n2477 vdd.n2476 185
R492 vdd.n2478 vdd.n2477 185
R493 vdd.n2475 vdd.n706 185
R494 vdd.n2474 vdd.n2473 185
R495 vdd.n708 vdd.n707 185
R496 vdd.n2260 vdd.n2259 185
R497 vdd.n2262 vdd.n2261 185
R498 vdd.n2264 vdd.n2263 185
R499 vdd.n2266 vdd.n2265 185
R500 vdd.n2268 vdd.n2267 185
R501 vdd.n2270 vdd.n2269 185
R502 vdd.n2272 vdd.n2271 185
R503 vdd.n2274 vdd.n2273 185
R504 vdd.n2276 vdd.n2275 185
R505 vdd.n2278 vdd.n2277 185
R506 vdd.n2280 vdd.n2279 185
R507 vdd.n2282 vdd.n2281 185
R508 vdd.n2284 vdd.n2283 185
R509 vdd.n2286 vdd.n2285 185
R510 vdd.n2288 vdd.n2287 185
R511 vdd.n2290 vdd.n2289 185
R512 vdd.n2292 vdd.n2291 185
R513 vdd.n2294 vdd.n2293 185
R514 vdd.n2296 vdd.n2295 185
R515 vdd.n2298 vdd.n2297 185
R516 vdd.n2300 vdd.n2299 185
R517 vdd.n2302 vdd.n2301 185
R518 vdd.n2304 vdd.n2303 185
R519 vdd.n2306 vdd.n2305 185
R520 vdd.n2308 vdd.n2307 185
R521 vdd.n2310 vdd.n2309 185
R522 vdd.n2312 vdd.n2311 185
R523 vdd.n2314 vdd.n2313 185
R524 vdd.n2316 vdd.n2315 185
R525 vdd.n2318 vdd.n2317 185
R526 vdd.n2320 vdd.n2319 185
R527 vdd.n2321 vdd.n2251 185
R528 vdd.n2471 vdd.n2251 185
R529 vdd.n2676 vdd.n2675 185
R530 vdd.n2677 vdd.n588 185
R531 vdd.n2679 vdd.n2678 185
R532 vdd.n2681 vdd.n586 185
R533 vdd.n2683 vdd.n2682 185
R534 vdd.n2684 vdd.n585 185
R535 vdd.n2686 vdd.n2685 185
R536 vdd.n2688 vdd.n583 185
R537 vdd.n2690 vdd.n2689 185
R538 vdd.n2691 vdd.n582 185
R539 vdd.n2693 vdd.n2692 185
R540 vdd.n2695 vdd.n580 185
R541 vdd.n2697 vdd.n2696 185
R542 vdd.n2698 vdd.n579 185
R543 vdd.n2700 vdd.n2699 185
R544 vdd.n2702 vdd.n578 185
R545 vdd.n2703 vdd.n576 185
R546 vdd.n2706 vdd.n2705 185
R547 vdd.n577 vdd.n575 185
R548 vdd.n2562 vdd.n2561 185
R549 vdd.n2564 vdd.n2563 185
R550 vdd.n2566 vdd.n2558 185
R551 vdd.n2568 vdd.n2567 185
R552 vdd.n2569 vdd.n2557 185
R553 vdd.n2571 vdd.n2570 185
R554 vdd.n2573 vdd.n2555 185
R555 vdd.n2575 vdd.n2574 185
R556 vdd.n2576 vdd.n2554 185
R557 vdd.n2578 vdd.n2577 185
R558 vdd.n2580 vdd.n2552 185
R559 vdd.n2582 vdd.n2581 185
R560 vdd.n2583 vdd.n2551 185
R561 vdd.n2585 vdd.n2584 185
R562 vdd.n2587 vdd.n2550 185
R563 vdd.n2589 vdd.n2588 185
R564 vdd.n2588 vdd.n484 185
R565 vdd.n2674 vdd.n592 185
R566 vdd.n2674 vdd.n2673 185
R567 vdd.n2326 vdd.n594 185
R568 vdd.n595 vdd.n594 185
R569 vdd.n2327 vdd.n628 185
R570 vdd.n2603 vdd.n628 185
R571 vdd.n2329 vdd.n2328 185
R572 vdd.n2328 vdd.n636 185
R573 vdd.n2330 vdd.n635 185
R574 vdd.n2597 vdd.n635 185
R575 vdd.n2332 vdd.n2331 185
R576 vdd.n2331 vdd.n633 185
R577 vdd.n2333 vdd.n643 185
R578 vdd.n2546 vdd.n643 185
R579 vdd.n2335 vdd.n2334 185
R580 vdd.n2334 vdd.n641 185
R581 vdd.n2336 vdd.n649 185
R582 vdd.n2540 vdd.n649 185
R583 vdd.n2338 vdd.n2337 185
R584 vdd.n2337 vdd.n647 185
R585 vdd.n2339 vdd.n654 185
R586 vdd.n2532 vdd.n654 185
R587 vdd.n2341 vdd.n2340 185
R588 vdd.n2340 vdd.n660 185
R589 vdd.n2342 vdd.n659 185
R590 vdd.n2526 vdd.n659 185
R591 vdd.n2376 vdd.n2375 185
R592 vdd.n2375 vdd.n2374 185
R593 vdd.n2377 vdd.n666 185
R594 vdd.n2520 vdd.n666 185
R595 vdd.n2379 vdd.n2378 185
R596 vdd.n2378 vdd.n664 185
R597 vdd.n2380 vdd.n672 185
R598 vdd.n2514 vdd.n672 185
R599 vdd.n2382 vdd.n2381 185
R600 vdd.n2381 vdd.n670 185
R601 vdd.n2383 vdd.n677 185
R602 vdd.n2508 vdd.n677 185
R603 vdd.n2385 vdd.n2384 185
R604 vdd.n2384 vdd.n683 185
R605 vdd.n2386 vdd.n682 185
R606 vdd.n2502 vdd.n682 185
R607 vdd.n2388 vdd.n2387 185
R608 vdd.n2387 vdd.n690 185
R609 vdd.n2389 vdd.n689 185
R610 vdd.n2496 vdd.n689 185
R611 vdd.n2391 vdd.n2390 185
R612 vdd.n2390 vdd.n687 185
R613 vdd.n2392 vdd.n695 185
R614 vdd.n2490 vdd.n695 185
R615 vdd.n2394 vdd.n2393 185
R616 vdd.n2395 vdd.n2394 185
R617 vdd.n2325 vdd.n700 185
R618 vdd.n2484 vdd.n700 185
R619 vdd.n2324 vdd.n2323 185
R620 vdd.n2323 vdd.t172 185
R621 vdd.n2322 vdd.n705 185
R622 vdd.n2478 vdd.n705 185
R623 vdd.n1942 vdd.n1941 185
R624 vdd.n1943 vdd.n1942 185
R625 vdd.n866 vdd.n864 185
R626 vdd.n1508 vdd.n864 185
R627 vdd.n1511 vdd.n1510 185
R628 vdd.n1510 vdd.n1509 185
R629 vdd.n869 vdd.n868 185
R630 vdd.n870 vdd.n869 185
R631 vdd.n1497 vdd.n1496 185
R632 vdd.n1498 vdd.n1497 185
R633 vdd.n878 vdd.n877 185
R634 vdd.n1489 vdd.n877 185
R635 vdd.n1492 vdd.n1491 185
R636 vdd.n1491 vdd.n1490 185
R637 vdd.n881 vdd.n880 185
R638 vdd.n888 vdd.n881 185
R639 vdd.n1480 vdd.n1479 185
R640 vdd.n1481 vdd.n1480 185
R641 vdd.n890 vdd.n889 185
R642 vdd.n889 vdd.n887 185
R643 vdd.n1475 vdd.n1474 185
R644 vdd.n1474 vdd.n1473 185
R645 vdd.n1163 vdd.n1162 185
R646 vdd.n1164 vdd.n1163 185
R647 vdd.n1464 vdd.n1463 185
R648 vdd.n1465 vdd.n1464 185
R649 vdd.n1171 vdd.n1170 185
R650 vdd.n1455 vdd.n1170 185
R651 vdd.n1458 vdd.n1457 185
R652 vdd.n1457 vdd.n1456 185
R653 vdd.n1174 vdd.n1173 185
R654 vdd.n1180 vdd.n1174 185
R655 vdd.n1446 vdd.n1445 185
R656 vdd.n1447 vdd.n1446 185
R657 vdd.n1182 vdd.n1181 185
R658 vdd.n1438 vdd.n1181 185
R659 vdd.n1441 vdd.n1440 185
R660 vdd.n1440 vdd.n1439 185
R661 vdd.n1185 vdd.n1184 185
R662 vdd.n1186 vdd.n1185 185
R663 vdd.n1429 vdd.n1428 185
R664 vdd.n1430 vdd.n1429 185
R665 vdd.n1193 vdd.n1192 185
R666 vdd.n1228 vdd.n1192 185
R667 vdd.n1424 vdd.n1423 185
R668 vdd.n1196 vdd.n1195 185
R669 vdd.n1420 vdd.n1419 185
R670 vdd.n1421 vdd.n1420 185
R671 vdd.n1230 vdd.n1229 185
R672 vdd.n1415 vdd.n1232 185
R673 vdd.n1414 vdd.n1233 185
R674 vdd.n1413 vdd.n1234 185
R675 vdd.n1236 vdd.n1235 185
R676 vdd.n1409 vdd.n1238 185
R677 vdd.n1408 vdd.n1239 185
R678 vdd.n1407 vdd.n1240 185
R679 vdd.n1242 vdd.n1241 185
R680 vdd.n1403 vdd.n1244 185
R681 vdd.n1402 vdd.n1245 185
R682 vdd.n1401 vdd.n1246 185
R683 vdd.n1248 vdd.n1247 185
R684 vdd.n1397 vdd.n1250 185
R685 vdd.n1396 vdd.n1251 185
R686 vdd.n1395 vdd.n1252 185
R687 vdd.n1256 vdd.n1253 185
R688 vdd.n1391 vdd.n1258 185
R689 vdd.n1390 vdd.n1259 185
R690 vdd.n1389 vdd.n1260 185
R691 vdd.n1262 vdd.n1261 185
R692 vdd.n1385 vdd.n1264 185
R693 vdd.n1384 vdd.n1265 185
R694 vdd.n1383 vdd.n1266 185
R695 vdd.n1268 vdd.n1267 185
R696 vdd.n1379 vdd.n1270 185
R697 vdd.n1378 vdd.n1271 185
R698 vdd.n1377 vdd.n1272 185
R699 vdd.n1274 vdd.n1273 185
R700 vdd.n1373 vdd.n1276 185
R701 vdd.n1372 vdd.n1277 185
R702 vdd.n1371 vdd.n1278 185
R703 vdd.n1280 vdd.n1279 185
R704 vdd.n1367 vdd.n1282 185
R705 vdd.n1366 vdd.n1283 185
R706 vdd.n1365 vdd.n1284 185
R707 vdd.n1286 vdd.n1285 185
R708 vdd.n1361 vdd.n1288 185
R709 vdd.n1360 vdd.n1357 185
R710 vdd.n1356 vdd.n1289 185
R711 vdd.n1291 vdd.n1290 185
R712 vdd.n1352 vdd.n1293 185
R713 vdd.n1351 vdd.n1294 185
R714 vdd.n1350 vdd.n1295 185
R715 vdd.n1297 vdd.n1296 185
R716 vdd.n1346 vdd.n1299 185
R717 vdd.n1345 vdd.n1300 185
R718 vdd.n1344 vdd.n1301 185
R719 vdd.n1303 vdd.n1302 185
R720 vdd.n1340 vdd.n1305 185
R721 vdd.n1339 vdd.n1306 185
R722 vdd.n1338 vdd.n1307 185
R723 vdd.n1309 vdd.n1308 185
R724 vdd.n1334 vdd.n1311 185
R725 vdd.n1333 vdd.n1312 185
R726 vdd.n1332 vdd.n1313 185
R727 vdd.n1315 vdd.n1314 185
R728 vdd.n1328 vdd.n1317 185
R729 vdd.n1327 vdd.n1318 185
R730 vdd.n1326 vdd.n1319 185
R731 vdd.n1323 vdd.n1227 185
R732 vdd.n1421 vdd.n1227 185
R733 vdd.n1946 vdd.n1945 185
R734 vdd.n1950 vdd.n859 185
R735 vdd.n1613 vdd.n858 185
R736 vdd.n1616 vdd.n1615 185
R737 vdd.n1618 vdd.n1617 185
R738 vdd.n1621 vdd.n1620 185
R739 vdd.n1623 vdd.n1622 185
R740 vdd.n1625 vdd.n1611 185
R741 vdd.n1627 vdd.n1626 185
R742 vdd.n1628 vdd.n1605 185
R743 vdd.n1630 vdd.n1629 185
R744 vdd.n1632 vdd.n1603 185
R745 vdd.n1634 vdd.n1633 185
R746 vdd.n1635 vdd.n1598 185
R747 vdd.n1637 vdd.n1636 185
R748 vdd.n1639 vdd.n1596 185
R749 vdd.n1641 vdd.n1640 185
R750 vdd.n1642 vdd.n1592 185
R751 vdd.n1644 vdd.n1643 185
R752 vdd.n1646 vdd.n1589 185
R753 vdd.n1648 vdd.n1647 185
R754 vdd.n1590 vdd.n1583 185
R755 vdd.n1652 vdd.n1587 185
R756 vdd.n1653 vdd.n1579 185
R757 vdd.n1655 vdd.n1654 185
R758 vdd.n1657 vdd.n1577 185
R759 vdd.n1659 vdd.n1658 185
R760 vdd.n1660 vdd.n1572 185
R761 vdd.n1662 vdd.n1661 185
R762 vdd.n1664 vdd.n1570 185
R763 vdd.n1666 vdd.n1665 185
R764 vdd.n1667 vdd.n1565 185
R765 vdd.n1669 vdd.n1668 185
R766 vdd.n1671 vdd.n1563 185
R767 vdd.n1673 vdd.n1672 185
R768 vdd.n1674 vdd.n1558 185
R769 vdd.n1676 vdd.n1675 185
R770 vdd.n1678 vdd.n1556 185
R771 vdd.n1680 vdd.n1679 185
R772 vdd.n1681 vdd.n1552 185
R773 vdd.n1683 vdd.n1682 185
R774 vdd.n1685 vdd.n1549 185
R775 vdd.n1687 vdd.n1686 185
R776 vdd.n1550 vdd.n1543 185
R777 vdd.n1691 vdd.n1547 185
R778 vdd.n1692 vdd.n1539 185
R779 vdd.n1694 vdd.n1693 185
R780 vdd.n1696 vdd.n1537 185
R781 vdd.n1698 vdd.n1697 185
R782 vdd.n1699 vdd.n1532 185
R783 vdd.n1701 vdd.n1700 185
R784 vdd.n1703 vdd.n1530 185
R785 vdd.n1705 vdd.n1704 185
R786 vdd.n1706 vdd.n1525 185
R787 vdd.n1708 vdd.n1707 185
R788 vdd.n1710 vdd.n1524 185
R789 vdd.n1711 vdd.n1521 185
R790 vdd.n1714 vdd.n1713 185
R791 vdd.n1523 vdd.n1519 185
R792 vdd.n1931 vdd.n1517 185
R793 vdd.n1933 vdd.n1932 185
R794 vdd.n1935 vdd.n1515 185
R795 vdd.n1937 vdd.n1936 185
R796 vdd.n1938 vdd.n865 185
R797 vdd.n1944 vdd.n862 185
R798 vdd.n1944 vdd.n1943 185
R799 vdd.n873 vdd.n861 185
R800 vdd.n1508 vdd.n861 185
R801 vdd.n1507 vdd.n1506 185
R802 vdd.n1509 vdd.n1507 185
R803 vdd.n872 vdd.n871 185
R804 vdd.n871 vdd.n870 185
R805 vdd.n1500 vdd.n1499 185
R806 vdd.n1499 vdd.n1498 185
R807 vdd.n876 vdd.n875 185
R808 vdd.n1489 vdd.n876 185
R809 vdd.n1488 vdd.n1487 185
R810 vdd.n1490 vdd.n1488 185
R811 vdd.n883 vdd.n882 185
R812 vdd.n888 vdd.n882 185
R813 vdd.n1483 vdd.n1482 185
R814 vdd.n1482 vdd.n1481 185
R815 vdd.n886 vdd.n885 185
R816 vdd.n887 vdd.n886 185
R817 vdd.n1472 vdd.n1471 185
R818 vdd.n1473 vdd.n1472 185
R819 vdd.n1166 vdd.n1165 185
R820 vdd.n1165 vdd.n1164 185
R821 vdd.n1467 vdd.n1466 185
R822 vdd.n1466 vdd.n1465 185
R823 vdd.n1169 vdd.n1168 185
R824 vdd.n1455 vdd.n1169 185
R825 vdd.n1454 vdd.n1453 185
R826 vdd.n1456 vdd.n1454 185
R827 vdd.n1176 vdd.n1175 185
R828 vdd.n1180 vdd.n1175 185
R829 vdd.n1449 vdd.n1448 185
R830 vdd.n1448 vdd.n1447 185
R831 vdd.n1179 vdd.n1178 185
R832 vdd.n1438 vdd.n1179 185
R833 vdd.n1437 vdd.n1436 185
R834 vdd.n1439 vdd.n1437 185
R835 vdd.n1188 vdd.n1187 185
R836 vdd.n1187 vdd.n1186 185
R837 vdd.n1432 vdd.n1431 185
R838 vdd.n1431 vdd.n1430 185
R839 vdd.n1191 vdd.n1190 185
R840 vdd.n1228 vdd.n1191 185
R841 vdd.n746 vdd.n744 185
R842 vdd.n2146 vdd.n744 185
R843 vdd.n2068 vdd.n763 185
R844 vdd.n763 vdd.t182 185
R845 vdd.n2070 vdd.n2069 185
R846 vdd.n2071 vdd.n2070 185
R847 vdd.n2067 vdd.n762 185
R848 vdd.n1770 vdd.n762 185
R849 vdd.n2066 vdd.n2065 185
R850 vdd.n2065 vdd.n2064 185
R851 vdd.n765 vdd.n764 185
R852 vdd.n766 vdd.n765 185
R853 vdd.n2055 vdd.n2054 185
R854 vdd.n2056 vdd.n2055 185
R855 vdd.n2053 vdd.n776 185
R856 vdd.n776 vdd.n773 185
R857 vdd.n2052 vdd.n2051 185
R858 vdd.n2051 vdd.n2050 185
R859 vdd.n778 vdd.n777 185
R860 vdd.n779 vdd.n778 185
R861 vdd.n2043 vdd.n2042 185
R862 vdd.n2044 vdd.n2043 185
R863 vdd.n2041 vdd.n787 185
R864 vdd.n792 vdd.n787 185
R865 vdd.n2040 vdd.n2039 185
R866 vdd.n2039 vdd.n2038 185
R867 vdd.n789 vdd.n788 185
R868 vdd.n798 vdd.n789 185
R869 vdd.n2031 vdd.n2030 185
R870 vdd.n2032 vdd.n2031 185
R871 vdd.n2029 vdd.n799 185
R872 vdd.n1871 vdd.n799 185
R873 vdd.n2028 vdd.n2027 185
R874 vdd.n2027 vdd.n2026 185
R875 vdd.n801 vdd.n800 185
R876 vdd.n802 vdd.n801 185
R877 vdd.n2019 vdd.n2018 185
R878 vdd.n2020 vdd.n2019 185
R879 vdd.n2017 vdd.n811 185
R880 vdd.n811 vdd.n808 185
R881 vdd.n2016 vdd.n2015 185
R882 vdd.n2015 vdd.n2014 185
R883 vdd.n813 vdd.n812 185
R884 vdd.n823 vdd.n813 185
R885 vdd.n2006 vdd.n2005 185
R886 vdd.n2007 vdd.n2006 185
R887 vdd.n2004 vdd.n824 185
R888 vdd.n824 vdd.n820 185
R889 vdd.n2003 vdd.n2002 185
R890 vdd.n2002 vdd.n2001 185
R891 vdd.n826 vdd.n825 185
R892 vdd.n827 vdd.n826 185
R893 vdd.n1994 vdd.n1993 185
R894 vdd.n1995 vdd.n1994 185
R895 vdd.n1992 vdd.n836 185
R896 vdd.n836 vdd.n833 185
R897 vdd.n1991 vdd.n1990 185
R898 vdd.n1990 vdd.n1989 185
R899 vdd.n838 vdd.n837 185
R900 vdd.n1726 vdd.n1725 185
R901 vdd.n1727 vdd.n1723 185
R902 vdd.n1723 vdd.n839 185
R903 vdd.n1729 vdd.n1728 185
R904 vdd.n1731 vdd.n1722 185
R905 vdd.n1734 vdd.n1733 185
R906 vdd.n1735 vdd.n1721 185
R907 vdd.n1737 vdd.n1736 185
R908 vdd.n1739 vdd.n1720 185
R909 vdd.n1742 vdd.n1741 185
R910 vdd.n1743 vdd.n1719 185
R911 vdd.n1745 vdd.n1744 185
R912 vdd.n1747 vdd.n1718 185
R913 vdd.n1750 vdd.n1749 185
R914 vdd.n1751 vdd.n1717 185
R915 vdd.n1753 vdd.n1752 185
R916 vdd.n1755 vdd.n1716 185
R917 vdd.n1928 vdd.n1756 185
R918 vdd.n1927 vdd.n1926 185
R919 vdd.n1924 vdd.n1757 185
R920 vdd.n1922 vdd.n1921 185
R921 vdd.n1920 vdd.n1758 185
R922 vdd.n1919 vdd.n1918 185
R923 vdd.n1916 vdd.n1759 185
R924 vdd.n1914 vdd.n1913 185
R925 vdd.n1912 vdd.n1760 185
R926 vdd.n1911 vdd.n1910 185
R927 vdd.n1908 vdd.n1761 185
R928 vdd.n1906 vdd.n1905 185
R929 vdd.n1904 vdd.n1762 185
R930 vdd.n1903 vdd.n1902 185
R931 vdd.n1900 vdd.n1763 185
R932 vdd.n1898 vdd.n1897 185
R933 vdd.n1896 vdd.n1764 185
R934 vdd.n1895 vdd.n1894 185
R935 vdd.n2149 vdd.n2148 185
R936 vdd.n2151 vdd.n2150 185
R937 vdd.n2153 vdd.n2152 185
R938 vdd.n2156 vdd.n2155 185
R939 vdd.n2158 vdd.n2157 185
R940 vdd.n2160 vdd.n2159 185
R941 vdd.n2162 vdd.n2161 185
R942 vdd.n2164 vdd.n2163 185
R943 vdd.n2166 vdd.n2165 185
R944 vdd.n2168 vdd.n2167 185
R945 vdd.n2170 vdd.n2169 185
R946 vdd.n2172 vdd.n2171 185
R947 vdd.n2174 vdd.n2173 185
R948 vdd.n2176 vdd.n2175 185
R949 vdd.n2178 vdd.n2177 185
R950 vdd.n2180 vdd.n2179 185
R951 vdd.n2182 vdd.n2181 185
R952 vdd.n2184 vdd.n2183 185
R953 vdd.n2186 vdd.n2185 185
R954 vdd.n2188 vdd.n2187 185
R955 vdd.n2190 vdd.n2189 185
R956 vdd.n2192 vdd.n2191 185
R957 vdd.n2194 vdd.n2193 185
R958 vdd.n2196 vdd.n2195 185
R959 vdd.n2198 vdd.n2197 185
R960 vdd.n2200 vdd.n2199 185
R961 vdd.n2202 vdd.n2201 185
R962 vdd.n2204 vdd.n2203 185
R963 vdd.n2206 vdd.n2205 185
R964 vdd.n2208 vdd.n2207 185
R965 vdd.n2210 vdd.n2209 185
R966 vdd.n2212 vdd.n2211 185
R967 vdd.n2214 vdd.n2213 185
R968 vdd.n2215 vdd.n745 185
R969 vdd.n2217 vdd.n2216 185
R970 vdd.n2218 vdd.n2217 185
R971 vdd.n2147 vdd.n749 185
R972 vdd.n2147 vdd.n2146 185
R973 vdd.n1768 vdd.n750 185
R974 vdd.t182 vdd.n750 185
R975 vdd.n1769 vdd.n760 185
R976 vdd.n2071 vdd.n760 185
R977 vdd.n1772 vdd.n1771 185
R978 vdd.n1771 vdd.n1770 185
R979 vdd.n1773 vdd.n767 185
R980 vdd.n2064 vdd.n767 185
R981 vdd.n1775 vdd.n1774 185
R982 vdd.n1774 vdd.n766 185
R983 vdd.n1776 vdd.n774 185
R984 vdd.n2056 vdd.n774 185
R985 vdd.n1778 vdd.n1777 185
R986 vdd.n1777 vdd.n773 185
R987 vdd.n1779 vdd.n780 185
R988 vdd.n2050 vdd.n780 185
R989 vdd.n1781 vdd.n1780 185
R990 vdd.n1780 vdd.n779 185
R991 vdd.n1782 vdd.n785 185
R992 vdd.n2044 vdd.n785 185
R993 vdd.n1784 vdd.n1783 185
R994 vdd.n1783 vdd.n792 185
R995 vdd.n1785 vdd.n790 185
R996 vdd.n2038 vdd.n790 185
R997 vdd.n1787 vdd.n1786 185
R998 vdd.n1786 vdd.n798 185
R999 vdd.n1788 vdd.n796 185
R1000 vdd.n2032 vdd.n796 185
R1001 vdd.n1873 vdd.n1872 185
R1002 vdd.n1872 vdd.n1871 185
R1003 vdd.n1874 vdd.n803 185
R1004 vdd.n2026 vdd.n803 185
R1005 vdd.n1876 vdd.n1875 185
R1006 vdd.n1875 vdd.n802 185
R1007 vdd.n1877 vdd.n809 185
R1008 vdd.n2020 vdd.n809 185
R1009 vdd.n1879 vdd.n1878 185
R1010 vdd.n1878 vdd.n808 185
R1011 vdd.n1880 vdd.n814 185
R1012 vdd.n2014 vdd.n814 185
R1013 vdd.n1882 vdd.n1881 185
R1014 vdd.n1881 vdd.n823 185
R1015 vdd.n1883 vdd.n821 185
R1016 vdd.n2007 vdd.n821 185
R1017 vdd.n1885 vdd.n1884 185
R1018 vdd.n1884 vdd.n820 185
R1019 vdd.n1886 vdd.n828 185
R1020 vdd.n2001 vdd.n828 185
R1021 vdd.n1888 vdd.n1887 185
R1022 vdd.n1887 vdd.n827 185
R1023 vdd.n1889 vdd.n834 185
R1024 vdd.n1995 vdd.n834 185
R1025 vdd.n1891 vdd.n1890 185
R1026 vdd.n1890 vdd.n833 185
R1027 vdd.n1892 vdd.n840 185
R1028 vdd.n1989 vdd.n840 185
R1029 vdd.n3024 vdd.n3023 185
R1030 vdd.n3025 vdd.n3024 185
R1031 vdd.n325 vdd.n324 185
R1032 vdd.n3026 vdd.n325 185
R1033 vdd.n3029 vdd.n3028 185
R1034 vdd.n3028 vdd.n3027 185
R1035 vdd.n3030 vdd.n319 185
R1036 vdd.n319 vdd.n318 185
R1037 vdd.n3032 vdd.n3031 185
R1038 vdd.n3033 vdd.n3032 185
R1039 vdd.n314 vdd.n313 185
R1040 vdd.n3034 vdd.n314 185
R1041 vdd.n3037 vdd.n3036 185
R1042 vdd.n3036 vdd.n3035 185
R1043 vdd.n3038 vdd.n309 185
R1044 vdd.n309 vdd.n308 185
R1045 vdd.n3040 vdd.n3039 185
R1046 vdd.n3041 vdd.n3040 185
R1047 vdd.n303 vdd.n301 185
R1048 vdd.n3042 vdd.n303 185
R1049 vdd.n3045 vdd.n3044 185
R1050 vdd.n3044 vdd.n3043 185
R1051 vdd.n302 vdd.n300 185
R1052 vdd.n304 vdd.n302 185
R1053 vdd.n2881 vdd.n2880 185
R1054 vdd.n2882 vdd.n2881 185
R1055 vdd.n458 vdd.n457 185
R1056 vdd.n457 vdd.n456 185
R1057 vdd.n2876 vdd.n2875 185
R1058 vdd.n2875 vdd.n2874 185
R1059 vdd.n461 vdd.n460 185
R1060 vdd.n467 vdd.n461 185
R1061 vdd.n2865 vdd.n2864 185
R1062 vdd.n2866 vdd.n2865 185
R1063 vdd.n469 vdd.n468 185
R1064 vdd.n2857 vdd.n468 185
R1065 vdd.n2860 vdd.n2859 185
R1066 vdd.n2859 vdd.n2858 185
R1067 vdd.n472 vdd.n471 185
R1068 vdd.n473 vdd.n472 185
R1069 vdd.n2848 vdd.n2847 185
R1070 vdd.n2849 vdd.n2848 185
R1071 vdd.n480 vdd.n479 185
R1072 vdd.n516 vdd.n479 185
R1073 vdd.n2843 vdd.n2842 185
R1074 vdd.n483 vdd.n482 185
R1075 vdd.n2839 vdd.n2838 185
R1076 vdd.n2840 vdd.n2839 185
R1077 vdd.n518 vdd.n517 185
R1078 vdd.n522 vdd.n521 185
R1079 vdd.n2834 vdd.n523 185
R1080 vdd.n2833 vdd.n2832 185
R1081 vdd.n2831 vdd.n2830 185
R1082 vdd.n2829 vdd.n2828 185
R1083 vdd.n2827 vdd.n2826 185
R1084 vdd.n2825 vdd.n2824 185
R1085 vdd.n2823 vdd.n2822 185
R1086 vdd.n2821 vdd.n2820 185
R1087 vdd.n2819 vdd.n2818 185
R1088 vdd.n2817 vdd.n2816 185
R1089 vdd.n2815 vdd.n2814 185
R1090 vdd.n2813 vdd.n2812 185
R1091 vdd.n2811 vdd.n2810 185
R1092 vdd.n2809 vdd.n2808 185
R1093 vdd.n2807 vdd.n2806 185
R1094 vdd.n2798 vdd.n536 185
R1095 vdd.n2800 vdd.n2799 185
R1096 vdd.n2797 vdd.n2796 185
R1097 vdd.n2795 vdd.n2794 185
R1098 vdd.n2793 vdd.n2792 185
R1099 vdd.n2791 vdd.n2790 185
R1100 vdd.n2789 vdd.n2788 185
R1101 vdd.n2787 vdd.n2786 185
R1102 vdd.n2785 vdd.n2784 185
R1103 vdd.n2783 vdd.n2782 185
R1104 vdd.n2781 vdd.n2780 185
R1105 vdd.n2779 vdd.n2778 185
R1106 vdd.n2777 vdd.n2776 185
R1107 vdd.n2775 vdd.n2774 185
R1108 vdd.n2773 vdd.n2772 185
R1109 vdd.n2771 vdd.n2770 185
R1110 vdd.n2769 vdd.n2768 185
R1111 vdd.n2767 vdd.n2766 185
R1112 vdd.n2765 vdd.n2764 185
R1113 vdd.n2763 vdd.n2762 185
R1114 vdd.n2761 vdd.n2760 185
R1115 vdd.n2759 vdd.n2758 185
R1116 vdd.n2752 vdd.n556 185
R1117 vdd.n2754 vdd.n2753 185
R1118 vdd.n2751 vdd.n2750 185
R1119 vdd.n2749 vdd.n2748 185
R1120 vdd.n2747 vdd.n2746 185
R1121 vdd.n2745 vdd.n2744 185
R1122 vdd.n2743 vdd.n2742 185
R1123 vdd.n2741 vdd.n2740 185
R1124 vdd.n2739 vdd.n2738 185
R1125 vdd.n2737 vdd.n2736 185
R1126 vdd.n2735 vdd.n2734 185
R1127 vdd.n2733 vdd.n2732 185
R1128 vdd.n2731 vdd.n2730 185
R1129 vdd.n2729 vdd.n2728 185
R1130 vdd.n2727 vdd.n2726 185
R1131 vdd.n2725 vdd.n2724 185
R1132 vdd.n2723 vdd.n2722 185
R1133 vdd.n2721 vdd.n2720 185
R1134 vdd.n2719 vdd.n2718 185
R1135 vdd.n2717 vdd.n2716 185
R1136 vdd.n2715 vdd.n2714 185
R1137 vdd.n2710 vdd.n515 185
R1138 vdd.n2840 vdd.n515 185
R1139 vdd.n2907 vdd.n2906 185
R1140 vdd.n2911 vdd.n440 185
R1141 vdd.n2913 vdd.n2912 185
R1142 vdd.n2915 vdd.n438 185
R1143 vdd.n2917 vdd.n2916 185
R1144 vdd.n2918 vdd.n433 185
R1145 vdd.n2920 vdd.n2919 185
R1146 vdd.n2922 vdd.n431 185
R1147 vdd.n2924 vdd.n2923 185
R1148 vdd.n2925 vdd.n426 185
R1149 vdd.n2927 vdd.n2926 185
R1150 vdd.n2929 vdd.n424 185
R1151 vdd.n2931 vdd.n2930 185
R1152 vdd.n2932 vdd.n419 185
R1153 vdd.n2934 vdd.n2933 185
R1154 vdd.n2936 vdd.n417 185
R1155 vdd.n2938 vdd.n2937 185
R1156 vdd.n2939 vdd.n413 185
R1157 vdd.n2941 vdd.n2940 185
R1158 vdd.n2943 vdd.n410 185
R1159 vdd.n2945 vdd.n2944 185
R1160 vdd.n411 vdd.n404 185
R1161 vdd.n2949 vdd.n408 185
R1162 vdd.n2950 vdd.n400 185
R1163 vdd.n2952 vdd.n2951 185
R1164 vdd.n2954 vdd.n398 185
R1165 vdd.n2956 vdd.n2955 185
R1166 vdd.n2957 vdd.n393 185
R1167 vdd.n2959 vdd.n2958 185
R1168 vdd.n2961 vdd.n391 185
R1169 vdd.n2963 vdd.n2962 185
R1170 vdd.n2964 vdd.n386 185
R1171 vdd.n2966 vdd.n2965 185
R1172 vdd.n2968 vdd.n384 185
R1173 vdd.n2970 vdd.n2969 185
R1174 vdd.n2971 vdd.n379 185
R1175 vdd.n2973 vdd.n2972 185
R1176 vdd.n2975 vdd.n377 185
R1177 vdd.n2977 vdd.n2976 185
R1178 vdd.n2978 vdd.n373 185
R1179 vdd.n2980 vdd.n2979 185
R1180 vdd.n2982 vdd.n370 185
R1181 vdd.n2984 vdd.n2983 185
R1182 vdd.n371 vdd.n364 185
R1183 vdd.n2988 vdd.n368 185
R1184 vdd.n2989 vdd.n360 185
R1185 vdd.n2991 vdd.n2990 185
R1186 vdd.n2993 vdd.n358 185
R1187 vdd.n2995 vdd.n2994 185
R1188 vdd.n2996 vdd.n353 185
R1189 vdd.n2998 vdd.n2997 185
R1190 vdd.n3000 vdd.n351 185
R1191 vdd.n3002 vdd.n3001 185
R1192 vdd.n3003 vdd.n346 185
R1193 vdd.n3005 vdd.n3004 185
R1194 vdd.n3007 vdd.n344 185
R1195 vdd.n3009 vdd.n3008 185
R1196 vdd.n3010 vdd.n338 185
R1197 vdd.n3012 vdd.n3011 185
R1198 vdd.n3014 vdd.n337 185
R1199 vdd.n3015 vdd.n336 185
R1200 vdd.n3018 vdd.n3017 185
R1201 vdd.n3019 vdd.n334 185
R1202 vdd.n3020 vdd.n330 185
R1203 vdd.n2902 vdd.n328 185
R1204 vdd.n3025 vdd.n328 185
R1205 vdd.n2901 vdd.n327 185
R1206 vdd.n3026 vdd.n327 185
R1207 vdd.n2900 vdd.n326 185
R1208 vdd.n3027 vdd.n326 185
R1209 vdd.n446 vdd.n445 185
R1210 vdd.n445 vdd.n318 185
R1211 vdd.n2896 vdd.n317 185
R1212 vdd.n3033 vdd.n317 185
R1213 vdd.n2895 vdd.n316 185
R1214 vdd.n3034 vdd.n316 185
R1215 vdd.n2894 vdd.n315 185
R1216 vdd.n3035 vdd.n315 185
R1217 vdd.n449 vdd.n448 185
R1218 vdd.n448 vdd.n308 185
R1219 vdd.n2890 vdd.n307 185
R1220 vdd.n3041 vdd.n307 185
R1221 vdd.n2889 vdd.n306 185
R1222 vdd.n3042 vdd.n306 185
R1223 vdd.n2888 vdd.n305 185
R1224 vdd.n3043 vdd.n305 185
R1225 vdd.n455 vdd.n451 185
R1226 vdd.n455 vdd.n304 185
R1227 vdd.n2884 vdd.n2883 185
R1228 vdd.n2883 vdd.n2882 185
R1229 vdd.n454 vdd.n453 185
R1230 vdd.n456 vdd.n454 185
R1231 vdd.n2873 vdd.n2872 185
R1232 vdd.n2874 vdd.n2873 185
R1233 vdd.n463 vdd.n462 185
R1234 vdd.n467 vdd.n462 185
R1235 vdd.n2868 vdd.n2867 185
R1236 vdd.n2867 vdd.n2866 185
R1237 vdd.n466 vdd.n465 185
R1238 vdd.n2857 vdd.n466 185
R1239 vdd.n2856 vdd.n2855 185
R1240 vdd.n2858 vdd.n2856 185
R1241 vdd.n475 vdd.n474 185
R1242 vdd.n474 vdd.n473 185
R1243 vdd.n2851 vdd.n2850 185
R1244 vdd.n2850 vdd.n2849 185
R1245 vdd.n478 vdd.n477 185
R1246 vdd.n516 vdd.n478 185
R1247 vdd.n703 vdd.n702 185
R1248 vdd.n2469 vdd.n2468 185
R1249 vdd.n2467 vdd.n2252 185
R1250 vdd.n2471 vdd.n2252 185
R1251 vdd.n2466 vdd.n2465 185
R1252 vdd.n2464 vdd.n2463 185
R1253 vdd.n2462 vdd.n2461 185
R1254 vdd.n2460 vdd.n2459 185
R1255 vdd.n2458 vdd.n2457 185
R1256 vdd.n2456 vdd.n2455 185
R1257 vdd.n2454 vdd.n2453 185
R1258 vdd.n2452 vdd.n2451 185
R1259 vdd.n2450 vdd.n2449 185
R1260 vdd.n2448 vdd.n2447 185
R1261 vdd.n2446 vdd.n2445 185
R1262 vdd.n2444 vdd.n2443 185
R1263 vdd.n2442 vdd.n2441 185
R1264 vdd.n2440 vdd.n2439 185
R1265 vdd.n2438 vdd.n2437 185
R1266 vdd.n2436 vdd.n2435 185
R1267 vdd.n2434 vdd.n2433 185
R1268 vdd.n2432 vdd.n2431 185
R1269 vdd.n2430 vdd.n2429 185
R1270 vdd.n2428 vdd.n2427 185
R1271 vdd.n2426 vdd.n2425 185
R1272 vdd.n2424 vdd.n2423 185
R1273 vdd.n2422 vdd.n2421 185
R1274 vdd.n2420 vdd.n2419 185
R1275 vdd.n2418 vdd.n2417 185
R1276 vdd.n2416 vdd.n2415 185
R1277 vdd.n2414 vdd.n2413 185
R1278 vdd.n2412 vdd.n2411 185
R1279 vdd.n2410 vdd.n2409 185
R1280 vdd.n2407 vdd.n2406 185
R1281 vdd.n2405 vdd.n2404 185
R1282 vdd.n2403 vdd.n2402 185
R1283 vdd.n2609 vdd.n2608 185
R1284 vdd.n2611 vdd.n624 185
R1285 vdd.n2613 vdd.n2612 185
R1286 vdd.n2615 vdd.n621 185
R1287 vdd.n2617 vdd.n2616 185
R1288 vdd.n2619 vdd.n619 185
R1289 vdd.n2621 vdd.n2620 185
R1290 vdd.n2622 vdd.n618 185
R1291 vdd.n2624 vdd.n2623 185
R1292 vdd.n2626 vdd.n616 185
R1293 vdd.n2628 vdd.n2627 185
R1294 vdd.n2629 vdd.n615 185
R1295 vdd.n2631 vdd.n2630 185
R1296 vdd.n2633 vdd.n613 185
R1297 vdd.n2635 vdd.n2634 185
R1298 vdd.n2636 vdd.n612 185
R1299 vdd.n2638 vdd.n2637 185
R1300 vdd.n2640 vdd.n520 185
R1301 vdd.n2642 vdd.n2641 185
R1302 vdd.n2644 vdd.n610 185
R1303 vdd.n2646 vdd.n2645 185
R1304 vdd.n2647 vdd.n609 185
R1305 vdd.n2649 vdd.n2648 185
R1306 vdd.n2651 vdd.n607 185
R1307 vdd.n2653 vdd.n2652 185
R1308 vdd.n2654 vdd.n606 185
R1309 vdd.n2656 vdd.n2655 185
R1310 vdd.n2658 vdd.n604 185
R1311 vdd.n2660 vdd.n2659 185
R1312 vdd.n2661 vdd.n603 185
R1313 vdd.n2663 vdd.n2662 185
R1314 vdd.n2665 vdd.n602 185
R1315 vdd.n2666 vdd.n601 185
R1316 vdd.n2669 vdd.n2668 185
R1317 vdd.n2670 vdd.n599 185
R1318 vdd.n599 vdd.n484 185
R1319 vdd.n2607 vdd.n596 185
R1320 vdd.n2673 vdd.n596 185
R1321 vdd.n2606 vdd.n2605 185
R1322 vdd.n2605 vdd.n595 185
R1323 vdd.n2604 vdd.n626 185
R1324 vdd.n2604 vdd.n2603 185
R1325 vdd.n2358 vdd.n627 185
R1326 vdd.n636 vdd.n627 185
R1327 vdd.n2359 vdd.n634 185
R1328 vdd.n2597 vdd.n634 185
R1329 vdd.n2361 vdd.n2360 185
R1330 vdd.n2360 vdd.n633 185
R1331 vdd.n2362 vdd.n642 185
R1332 vdd.n2546 vdd.n642 185
R1333 vdd.n2364 vdd.n2363 185
R1334 vdd.n2363 vdd.n641 185
R1335 vdd.n2365 vdd.n648 185
R1336 vdd.n2540 vdd.n648 185
R1337 vdd.n2367 vdd.n2366 185
R1338 vdd.n2366 vdd.n647 185
R1339 vdd.n2368 vdd.n653 185
R1340 vdd.n2532 vdd.n653 185
R1341 vdd.n2370 vdd.n2369 185
R1342 vdd.n2369 vdd.n660 185
R1343 vdd.n2371 vdd.n658 185
R1344 vdd.n2526 vdd.n658 185
R1345 vdd.n2373 vdd.n2372 185
R1346 vdd.n2374 vdd.n2373 185
R1347 vdd.n2357 vdd.n665 185
R1348 vdd.n2520 vdd.n665 185
R1349 vdd.n2356 vdd.n2355 185
R1350 vdd.n2355 vdd.n664 185
R1351 vdd.n2354 vdd.n671 185
R1352 vdd.n2514 vdd.n671 185
R1353 vdd.n2353 vdd.n2352 185
R1354 vdd.n2352 vdd.n670 185
R1355 vdd.n2351 vdd.n676 185
R1356 vdd.n2508 vdd.n676 185
R1357 vdd.n2350 vdd.n2349 185
R1358 vdd.n2349 vdd.n683 185
R1359 vdd.n2348 vdd.n681 185
R1360 vdd.n2502 vdd.n681 185
R1361 vdd.n2347 vdd.n2346 185
R1362 vdd.n2346 vdd.n690 185
R1363 vdd.n2345 vdd.n688 185
R1364 vdd.n2496 vdd.n688 185
R1365 vdd.n2344 vdd.n2343 185
R1366 vdd.n2343 vdd.n687 185
R1367 vdd.n2255 vdd.n694 185
R1368 vdd.n2490 vdd.n694 185
R1369 vdd.n2397 vdd.n2396 185
R1370 vdd.n2396 vdd.n2395 185
R1371 vdd.n2398 vdd.n699 185
R1372 vdd.n2484 vdd.n699 185
R1373 vdd.n2400 vdd.n2399 185
R1374 vdd.n2399 vdd.t172 185
R1375 vdd.n2401 vdd.n704 185
R1376 vdd.n2478 vdd.n704 185
R1377 vdd.n2480 vdd.n2479 185
R1378 vdd.n2479 vdd.n2478 185
R1379 vdd.n2481 vdd.n701 185
R1380 vdd.n701 vdd.t172 185
R1381 vdd.n2483 vdd.n2482 185
R1382 vdd.n2484 vdd.n2483 185
R1383 vdd.n693 vdd.n692 185
R1384 vdd.n2395 vdd.n693 185
R1385 vdd.n2492 vdd.n2491 185
R1386 vdd.n2491 vdd.n2490 185
R1387 vdd.n2493 vdd.n691 185
R1388 vdd.n691 vdd.n687 185
R1389 vdd.n2495 vdd.n2494 185
R1390 vdd.n2496 vdd.n2495 185
R1391 vdd.n680 vdd.n679 185
R1392 vdd.n690 vdd.n680 185
R1393 vdd.n2504 vdd.n2503 185
R1394 vdd.n2503 vdd.n2502 185
R1395 vdd.n2505 vdd.n678 185
R1396 vdd.n683 vdd.n678 185
R1397 vdd.n2507 vdd.n2506 185
R1398 vdd.n2508 vdd.n2507 185
R1399 vdd.n669 vdd.n668 185
R1400 vdd.n670 vdd.n669 185
R1401 vdd.n2516 vdd.n2515 185
R1402 vdd.n2515 vdd.n2514 185
R1403 vdd.n2517 vdd.n667 185
R1404 vdd.n667 vdd.n664 185
R1405 vdd.n2519 vdd.n2518 185
R1406 vdd.n2520 vdd.n2519 185
R1407 vdd.n657 vdd.n656 185
R1408 vdd.n2374 vdd.n657 185
R1409 vdd.n2528 vdd.n2527 185
R1410 vdd.n2527 vdd.n2526 185
R1411 vdd.n2529 vdd.n655 185
R1412 vdd.n660 vdd.n655 185
R1413 vdd.n2531 vdd.n2530 185
R1414 vdd.n2532 vdd.n2531 185
R1415 vdd.n646 vdd.n645 185
R1416 vdd.n647 vdd.n646 185
R1417 vdd.n2542 vdd.n2541 185
R1418 vdd.n2541 vdd.n2540 185
R1419 vdd.n2543 vdd.n644 185
R1420 vdd.n644 vdd.n641 185
R1421 vdd.n2545 vdd.n2544 185
R1422 vdd.n2546 vdd.n2545 185
R1423 vdd.n632 vdd.n631 185
R1424 vdd.n633 vdd.n632 185
R1425 vdd.n2599 vdd.n2598 185
R1426 vdd.n2598 vdd.n2597 185
R1427 vdd.n2600 vdd.n630 185
R1428 vdd.n636 vdd.n630 185
R1429 vdd.n2602 vdd.n2601 185
R1430 vdd.n2603 vdd.n2602 185
R1431 vdd.n600 vdd.n598 185
R1432 vdd.n598 vdd.n595 185
R1433 vdd.n2672 vdd.n2671 185
R1434 vdd.n2673 vdd.n2672 185
R1435 vdd.n2145 vdd.n2144 185
R1436 vdd.n2146 vdd.n2145 185
R1437 vdd.n754 vdd.n752 185
R1438 vdd.n752 vdd.t182 185
R1439 vdd.n2060 vdd.n761 185
R1440 vdd.n2071 vdd.n761 185
R1441 vdd.n2061 vdd.n770 185
R1442 vdd.n1770 vdd.n770 185
R1443 vdd.n2063 vdd.n2062 185
R1444 vdd.n2064 vdd.n2063 185
R1445 vdd.n2059 vdd.n769 185
R1446 vdd.n769 vdd.n766 185
R1447 vdd.n2058 vdd.n2057 185
R1448 vdd.n2057 vdd.n2056 185
R1449 vdd.n772 vdd.n771 185
R1450 vdd.n773 vdd.n772 185
R1451 vdd.n2049 vdd.n2048 185
R1452 vdd.n2050 vdd.n2049 185
R1453 vdd.n2047 vdd.n782 185
R1454 vdd.n782 vdd.n779 185
R1455 vdd.n2046 vdd.n2045 185
R1456 vdd.n2045 vdd.n2044 185
R1457 vdd.n784 vdd.n783 185
R1458 vdd.n792 vdd.n784 185
R1459 vdd.n2037 vdd.n2036 185
R1460 vdd.n2038 vdd.n2037 185
R1461 vdd.n2035 vdd.n793 185
R1462 vdd.n798 vdd.n793 185
R1463 vdd.n2034 vdd.n2033 185
R1464 vdd.n2033 vdd.n2032 185
R1465 vdd.n795 vdd.n794 185
R1466 vdd.n1871 vdd.n795 185
R1467 vdd.n2025 vdd.n2024 185
R1468 vdd.n2026 vdd.n2025 185
R1469 vdd.n2023 vdd.n805 185
R1470 vdd.n805 vdd.n802 185
R1471 vdd.n2022 vdd.n2021 185
R1472 vdd.n2021 vdd.n2020 185
R1473 vdd.n807 vdd.n806 185
R1474 vdd.n808 vdd.n807 185
R1475 vdd.n2013 vdd.n2012 185
R1476 vdd.n2014 vdd.n2013 185
R1477 vdd.n2010 vdd.n816 185
R1478 vdd.n823 vdd.n816 185
R1479 vdd.n2009 vdd.n2008 185
R1480 vdd.n2008 vdd.n2007 185
R1481 vdd.n819 vdd.n818 185
R1482 vdd.n820 vdd.n819 185
R1483 vdd.n2000 vdd.n1999 185
R1484 vdd.n2001 vdd.n2000 185
R1485 vdd.n1998 vdd.n830 185
R1486 vdd.n830 vdd.n827 185
R1487 vdd.n1997 vdd.n1996 185
R1488 vdd.n1996 vdd.n1995 185
R1489 vdd.n832 vdd.n831 185
R1490 vdd.n833 vdd.n832 185
R1491 vdd.n1988 vdd.n1987 185
R1492 vdd.n1989 vdd.n1988 185
R1493 vdd.n2076 vdd.n726 185
R1494 vdd.n2218 vdd.n726 185
R1495 vdd.n2078 vdd.n2077 185
R1496 vdd.n2080 vdd.n2079 185
R1497 vdd.n2082 vdd.n2081 185
R1498 vdd.n2084 vdd.n2083 185
R1499 vdd.n2086 vdd.n2085 185
R1500 vdd.n2088 vdd.n2087 185
R1501 vdd.n2090 vdd.n2089 185
R1502 vdd.n2092 vdd.n2091 185
R1503 vdd.n2094 vdd.n2093 185
R1504 vdd.n2096 vdd.n2095 185
R1505 vdd.n2098 vdd.n2097 185
R1506 vdd.n2100 vdd.n2099 185
R1507 vdd.n2102 vdd.n2101 185
R1508 vdd.n2104 vdd.n2103 185
R1509 vdd.n2106 vdd.n2105 185
R1510 vdd.n2108 vdd.n2107 185
R1511 vdd.n2110 vdd.n2109 185
R1512 vdd.n2112 vdd.n2111 185
R1513 vdd.n2114 vdd.n2113 185
R1514 vdd.n2116 vdd.n2115 185
R1515 vdd.n2118 vdd.n2117 185
R1516 vdd.n2120 vdd.n2119 185
R1517 vdd.n2122 vdd.n2121 185
R1518 vdd.n2124 vdd.n2123 185
R1519 vdd.n2126 vdd.n2125 185
R1520 vdd.n2128 vdd.n2127 185
R1521 vdd.n2130 vdd.n2129 185
R1522 vdd.n2132 vdd.n2131 185
R1523 vdd.n2134 vdd.n2133 185
R1524 vdd.n2136 vdd.n2135 185
R1525 vdd.n2138 vdd.n2137 185
R1526 vdd.n2140 vdd.n2139 185
R1527 vdd.n2142 vdd.n2141 185
R1528 vdd.n2143 vdd.n753 185
R1529 vdd.n2075 vdd.n751 185
R1530 vdd.n2146 vdd.n751 185
R1531 vdd.n2074 vdd.n2073 185
R1532 vdd.n2073 vdd.t182 185
R1533 vdd.n2072 vdd.n758 185
R1534 vdd.n2072 vdd.n2071 185
R1535 vdd.n1852 vdd.n759 185
R1536 vdd.n1770 vdd.n759 185
R1537 vdd.n1853 vdd.n768 185
R1538 vdd.n2064 vdd.n768 185
R1539 vdd.n1855 vdd.n1854 185
R1540 vdd.n1854 vdd.n766 185
R1541 vdd.n1856 vdd.n775 185
R1542 vdd.n2056 vdd.n775 185
R1543 vdd.n1858 vdd.n1857 185
R1544 vdd.n1857 vdd.n773 185
R1545 vdd.n1859 vdd.n781 185
R1546 vdd.n2050 vdd.n781 185
R1547 vdd.n1861 vdd.n1860 185
R1548 vdd.n1860 vdd.n779 185
R1549 vdd.n1862 vdd.n786 185
R1550 vdd.n2044 vdd.n786 185
R1551 vdd.n1864 vdd.n1863 185
R1552 vdd.n1863 vdd.n792 185
R1553 vdd.n1865 vdd.n791 185
R1554 vdd.n2038 vdd.n791 185
R1555 vdd.n1867 vdd.n1866 185
R1556 vdd.n1866 vdd.n798 185
R1557 vdd.n1868 vdd.n797 185
R1558 vdd.n2032 vdd.n797 185
R1559 vdd.n1870 vdd.n1869 185
R1560 vdd.n1871 vdd.n1870 185
R1561 vdd.n1851 vdd.n804 185
R1562 vdd.n2026 vdd.n804 185
R1563 vdd.n1850 vdd.n1849 185
R1564 vdd.n1849 vdd.n802 185
R1565 vdd.n1848 vdd.n810 185
R1566 vdd.n2020 vdd.n810 185
R1567 vdd.n1847 vdd.n1846 185
R1568 vdd.n1846 vdd.n808 185
R1569 vdd.n1845 vdd.n815 185
R1570 vdd.n2014 vdd.n815 185
R1571 vdd.n1844 vdd.n1843 185
R1572 vdd.n1843 vdd.n823 185
R1573 vdd.n1842 vdd.n822 185
R1574 vdd.n2007 vdd.n822 185
R1575 vdd.n1841 vdd.n1840 185
R1576 vdd.n1840 vdd.n820 185
R1577 vdd.n1839 vdd.n829 185
R1578 vdd.n2001 vdd.n829 185
R1579 vdd.n1838 vdd.n1837 185
R1580 vdd.n1837 vdd.n827 185
R1581 vdd.n1836 vdd.n835 185
R1582 vdd.n1995 vdd.n835 185
R1583 vdd.n1835 vdd.n1834 185
R1584 vdd.n1834 vdd.n833 185
R1585 vdd.n1833 vdd.n841 185
R1586 vdd.n1989 vdd.n841 185
R1587 vdd.n1986 vdd.n842 185
R1588 vdd.n1985 vdd.n1984 185
R1589 vdd.n1982 vdd.n843 185
R1590 vdd.n1980 vdd.n1979 185
R1591 vdd.n1978 vdd.n844 185
R1592 vdd.n1977 vdd.n1976 185
R1593 vdd.n1974 vdd.n845 185
R1594 vdd.n1972 vdd.n1971 185
R1595 vdd.n1970 vdd.n846 185
R1596 vdd.n1969 vdd.n1968 185
R1597 vdd.n1966 vdd.n847 185
R1598 vdd.n1964 vdd.n1963 185
R1599 vdd.n1962 vdd.n848 185
R1600 vdd.n1961 vdd.n1960 185
R1601 vdd.n1958 vdd.n849 185
R1602 vdd.n1956 vdd.n1955 185
R1603 vdd.n1954 vdd.n850 185
R1604 vdd.n1953 vdd.n852 185
R1605 vdd.n1798 vdd.n853 185
R1606 vdd.n1801 vdd.n1800 185
R1607 vdd.n1803 vdd.n1802 185
R1608 vdd.n1805 vdd.n1797 185
R1609 vdd.n1808 vdd.n1807 185
R1610 vdd.n1809 vdd.n1796 185
R1611 vdd.n1811 vdd.n1810 185
R1612 vdd.n1813 vdd.n1795 185
R1613 vdd.n1816 vdd.n1815 185
R1614 vdd.n1817 vdd.n1794 185
R1615 vdd.n1819 vdd.n1818 185
R1616 vdd.n1821 vdd.n1793 185
R1617 vdd.n1824 vdd.n1823 185
R1618 vdd.n1825 vdd.n1790 185
R1619 vdd.n1828 vdd.n1827 185
R1620 vdd.n1830 vdd.n1789 185
R1621 vdd.n1832 vdd.n1831 185
R1622 vdd.n1831 vdd.n839 185
R1623 vdd.n291 vdd.n290 171.744
R1624 vdd.n290 vdd.n289 171.744
R1625 vdd.n289 vdd.n258 171.744
R1626 vdd.n282 vdd.n258 171.744
R1627 vdd.n282 vdd.n281 171.744
R1628 vdd.n281 vdd.n263 171.744
R1629 vdd.n274 vdd.n263 171.744
R1630 vdd.n274 vdd.n273 171.744
R1631 vdd.n273 vdd.n267 171.744
R1632 vdd.n244 vdd.n243 171.744
R1633 vdd.n243 vdd.n242 171.744
R1634 vdd.n242 vdd.n211 171.744
R1635 vdd.n235 vdd.n211 171.744
R1636 vdd.n235 vdd.n234 171.744
R1637 vdd.n234 vdd.n216 171.744
R1638 vdd.n227 vdd.n216 171.744
R1639 vdd.n227 vdd.n226 171.744
R1640 vdd.n226 vdd.n220 171.744
R1641 vdd.n201 vdd.n200 171.744
R1642 vdd.n200 vdd.n199 171.744
R1643 vdd.n199 vdd.n168 171.744
R1644 vdd.n192 vdd.n168 171.744
R1645 vdd.n192 vdd.n191 171.744
R1646 vdd.n191 vdd.n173 171.744
R1647 vdd.n184 vdd.n173 171.744
R1648 vdd.n184 vdd.n183 171.744
R1649 vdd.n183 vdd.n177 171.744
R1650 vdd.n154 vdd.n153 171.744
R1651 vdd.n153 vdd.n152 171.744
R1652 vdd.n152 vdd.n121 171.744
R1653 vdd.n145 vdd.n121 171.744
R1654 vdd.n145 vdd.n144 171.744
R1655 vdd.n144 vdd.n126 171.744
R1656 vdd.n137 vdd.n126 171.744
R1657 vdd.n137 vdd.n136 171.744
R1658 vdd.n136 vdd.n130 171.744
R1659 vdd.n112 vdd.n111 171.744
R1660 vdd.n111 vdd.n110 171.744
R1661 vdd.n110 vdd.n79 171.744
R1662 vdd.n103 vdd.n79 171.744
R1663 vdd.n103 vdd.n102 171.744
R1664 vdd.n102 vdd.n84 171.744
R1665 vdd.n95 vdd.n84 171.744
R1666 vdd.n95 vdd.n94 171.744
R1667 vdd.n94 vdd.n88 171.744
R1668 vdd.n65 vdd.n64 171.744
R1669 vdd.n64 vdd.n63 171.744
R1670 vdd.n63 vdd.n32 171.744
R1671 vdd.n56 vdd.n32 171.744
R1672 vdd.n56 vdd.n55 171.744
R1673 vdd.n55 vdd.n37 171.744
R1674 vdd.n48 vdd.n37 171.744
R1675 vdd.n48 vdd.n47 171.744
R1676 vdd.n47 vdd.n41 171.744
R1677 vdd.n1106 vdd.n1105 171.744
R1678 vdd.n1105 vdd.n1104 171.744
R1679 vdd.n1104 vdd.n1073 171.744
R1680 vdd.n1097 vdd.n1073 171.744
R1681 vdd.n1097 vdd.n1096 171.744
R1682 vdd.n1096 vdd.n1078 171.744
R1683 vdd.n1089 vdd.n1078 171.744
R1684 vdd.n1089 vdd.n1088 171.744
R1685 vdd.n1088 vdd.n1082 171.744
R1686 vdd.n1153 vdd.n1152 171.744
R1687 vdd.n1152 vdd.n1151 171.744
R1688 vdd.n1151 vdd.n1120 171.744
R1689 vdd.n1144 vdd.n1120 171.744
R1690 vdd.n1144 vdd.n1143 171.744
R1691 vdd.n1143 vdd.n1125 171.744
R1692 vdd.n1136 vdd.n1125 171.744
R1693 vdd.n1136 vdd.n1135 171.744
R1694 vdd.n1135 vdd.n1129 171.744
R1695 vdd.n1016 vdd.n1015 171.744
R1696 vdd.n1015 vdd.n1014 171.744
R1697 vdd.n1014 vdd.n983 171.744
R1698 vdd.n1007 vdd.n983 171.744
R1699 vdd.n1007 vdd.n1006 171.744
R1700 vdd.n1006 vdd.n988 171.744
R1701 vdd.n999 vdd.n988 171.744
R1702 vdd.n999 vdd.n998 171.744
R1703 vdd.n998 vdd.n992 171.744
R1704 vdd.n1063 vdd.n1062 171.744
R1705 vdd.n1062 vdd.n1061 171.744
R1706 vdd.n1061 vdd.n1030 171.744
R1707 vdd.n1054 vdd.n1030 171.744
R1708 vdd.n1054 vdd.n1053 171.744
R1709 vdd.n1053 vdd.n1035 171.744
R1710 vdd.n1046 vdd.n1035 171.744
R1711 vdd.n1046 vdd.n1045 171.744
R1712 vdd.n1045 vdd.n1039 171.744
R1713 vdd.n927 vdd.n926 171.744
R1714 vdd.n926 vdd.n925 171.744
R1715 vdd.n925 vdd.n894 171.744
R1716 vdd.n918 vdd.n894 171.744
R1717 vdd.n918 vdd.n917 171.744
R1718 vdd.n917 vdd.n899 171.744
R1719 vdd.n910 vdd.n899 171.744
R1720 vdd.n910 vdd.n909 171.744
R1721 vdd.n909 vdd.n903 171.744
R1722 vdd.n974 vdd.n973 171.744
R1723 vdd.n973 vdd.n972 171.744
R1724 vdd.n972 vdd.n941 171.744
R1725 vdd.n965 vdd.n941 171.744
R1726 vdd.n965 vdd.n964 171.744
R1727 vdd.n964 vdd.n946 171.744
R1728 vdd.n957 vdd.n946 171.744
R1729 vdd.n957 vdd.n956 171.744
R1730 vdd.n956 vdd.n950 171.744
R1731 vdd.n3017 vdd.n334 146.341
R1732 vdd.n3015 vdd.n3014 146.341
R1733 vdd.n3012 vdd.n338 146.341
R1734 vdd.n3008 vdd.n3007 146.341
R1735 vdd.n3005 vdd.n346 146.341
R1736 vdd.n3001 vdd.n3000 146.341
R1737 vdd.n2998 vdd.n353 146.341
R1738 vdd.n2994 vdd.n2993 146.341
R1739 vdd.n2991 vdd.n360 146.341
R1740 vdd.n371 vdd.n368 146.341
R1741 vdd.n2983 vdd.n2982 146.341
R1742 vdd.n2980 vdd.n373 146.341
R1743 vdd.n2976 vdd.n2975 146.341
R1744 vdd.n2973 vdd.n379 146.341
R1745 vdd.n2969 vdd.n2968 146.341
R1746 vdd.n2966 vdd.n386 146.341
R1747 vdd.n2962 vdd.n2961 146.341
R1748 vdd.n2959 vdd.n393 146.341
R1749 vdd.n2955 vdd.n2954 146.341
R1750 vdd.n2952 vdd.n400 146.341
R1751 vdd.n411 vdd.n408 146.341
R1752 vdd.n2944 vdd.n2943 146.341
R1753 vdd.n2941 vdd.n413 146.341
R1754 vdd.n2937 vdd.n2936 146.341
R1755 vdd.n2934 vdd.n419 146.341
R1756 vdd.n2930 vdd.n2929 146.341
R1757 vdd.n2927 vdd.n426 146.341
R1758 vdd.n2923 vdd.n2922 146.341
R1759 vdd.n2920 vdd.n433 146.341
R1760 vdd.n2916 vdd.n2915 146.341
R1761 vdd.n2913 vdd.n440 146.341
R1762 vdd.n2850 vdd.n478 146.341
R1763 vdd.n2850 vdd.n474 146.341
R1764 vdd.n2856 vdd.n474 146.341
R1765 vdd.n2856 vdd.n466 146.341
R1766 vdd.n2867 vdd.n466 146.341
R1767 vdd.n2867 vdd.n462 146.341
R1768 vdd.n2873 vdd.n462 146.341
R1769 vdd.n2873 vdd.n454 146.341
R1770 vdd.n2883 vdd.n454 146.341
R1771 vdd.n2883 vdd.n455 146.341
R1772 vdd.n455 vdd.n305 146.341
R1773 vdd.n306 vdd.n305 146.341
R1774 vdd.n307 vdd.n306 146.341
R1775 vdd.n448 vdd.n307 146.341
R1776 vdd.n448 vdd.n315 146.341
R1777 vdd.n316 vdd.n315 146.341
R1778 vdd.n317 vdd.n316 146.341
R1779 vdd.n445 vdd.n317 146.341
R1780 vdd.n445 vdd.n326 146.341
R1781 vdd.n327 vdd.n326 146.341
R1782 vdd.n328 vdd.n327 146.341
R1783 vdd.n2839 vdd.n483 146.341
R1784 vdd.n2839 vdd.n517 146.341
R1785 vdd.n523 vdd.n522 146.341
R1786 vdd.n2832 vdd.n2831 146.341
R1787 vdd.n2828 vdd.n2827 146.341
R1788 vdd.n2824 vdd.n2823 146.341
R1789 vdd.n2820 vdd.n2819 146.341
R1790 vdd.n2816 vdd.n2815 146.341
R1791 vdd.n2812 vdd.n2811 146.341
R1792 vdd.n2808 vdd.n2807 146.341
R1793 vdd.n2799 vdd.n2798 146.341
R1794 vdd.n2796 vdd.n2795 146.341
R1795 vdd.n2792 vdd.n2791 146.341
R1796 vdd.n2788 vdd.n2787 146.341
R1797 vdd.n2784 vdd.n2783 146.341
R1798 vdd.n2780 vdd.n2779 146.341
R1799 vdd.n2776 vdd.n2775 146.341
R1800 vdd.n2772 vdd.n2771 146.341
R1801 vdd.n2768 vdd.n2767 146.341
R1802 vdd.n2764 vdd.n2763 146.341
R1803 vdd.n2760 vdd.n2759 146.341
R1804 vdd.n2753 vdd.n2752 146.341
R1805 vdd.n2750 vdd.n2749 146.341
R1806 vdd.n2746 vdd.n2745 146.341
R1807 vdd.n2742 vdd.n2741 146.341
R1808 vdd.n2738 vdd.n2737 146.341
R1809 vdd.n2734 vdd.n2733 146.341
R1810 vdd.n2730 vdd.n2729 146.341
R1811 vdd.n2726 vdd.n2725 146.341
R1812 vdd.n2722 vdd.n2721 146.341
R1813 vdd.n2718 vdd.n2717 146.341
R1814 vdd.n2714 vdd.n515 146.341
R1815 vdd.n2848 vdd.n479 146.341
R1816 vdd.n2848 vdd.n472 146.341
R1817 vdd.n2859 vdd.n472 146.341
R1818 vdd.n2859 vdd.n468 146.341
R1819 vdd.n2865 vdd.n468 146.341
R1820 vdd.n2865 vdd.n461 146.341
R1821 vdd.n2875 vdd.n461 146.341
R1822 vdd.n2875 vdd.n457 146.341
R1823 vdd.n2881 vdd.n457 146.341
R1824 vdd.n2881 vdd.n302 146.341
R1825 vdd.n3044 vdd.n302 146.341
R1826 vdd.n3044 vdd.n303 146.341
R1827 vdd.n3040 vdd.n303 146.341
R1828 vdd.n3040 vdd.n309 146.341
R1829 vdd.n3036 vdd.n309 146.341
R1830 vdd.n3036 vdd.n314 146.341
R1831 vdd.n3032 vdd.n314 146.341
R1832 vdd.n3032 vdd.n319 146.341
R1833 vdd.n3028 vdd.n319 146.341
R1834 vdd.n3028 vdd.n325 146.341
R1835 vdd.n3024 vdd.n325 146.341
R1836 vdd.n1936 vdd.n1935 146.341
R1837 vdd.n1933 vdd.n1517 146.341
R1838 vdd.n1713 vdd.n1523 146.341
R1839 vdd.n1711 vdd.n1710 146.341
R1840 vdd.n1708 vdd.n1525 146.341
R1841 vdd.n1704 vdd.n1703 146.341
R1842 vdd.n1701 vdd.n1532 146.341
R1843 vdd.n1697 vdd.n1696 146.341
R1844 vdd.n1694 vdd.n1539 146.341
R1845 vdd.n1550 vdd.n1547 146.341
R1846 vdd.n1686 vdd.n1685 146.341
R1847 vdd.n1683 vdd.n1552 146.341
R1848 vdd.n1679 vdd.n1678 146.341
R1849 vdd.n1676 vdd.n1558 146.341
R1850 vdd.n1672 vdd.n1671 146.341
R1851 vdd.n1669 vdd.n1565 146.341
R1852 vdd.n1665 vdd.n1664 146.341
R1853 vdd.n1662 vdd.n1572 146.341
R1854 vdd.n1658 vdd.n1657 146.341
R1855 vdd.n1655 vdd.n1579 146.341
R1856 vdd.n1590 vdd.n1587 146.341
R1857 vdd.n1647 vdd.n1646 146.341
R1858 vdd.n1644 vdd.n1592 146.341
R1859 vdd.n1640 vdd.n1639 146.341
R1860 vdd.n1637 vdd.n1598 146.341
R1861 vdd.n1633 vdd.n1632 146.341
R1862 vdd.n1630 vdd.n1605 146.341
R1863 vdd.n1626 vdd.n1625 146.341
R1864 vdd.n1623 vdd.n1620 146.341
R1865 vdd.n1618 vdd.n1615 146.341
R1866 vdd.n1613 vdd.n859 146.341
R1867 vdd.n1431 vdd.n1191 146.341
R1868 vdd.n1431 vdd.n1187 146.341
R1869 vdd.n1437 vdd.n1187 146.341
R1870 vdd.n1437 vdd.n1179 146.341
R1871 vdd.n1448 vdd.n1179 146.341
R1872 vdd.n1448 vdd.n1175 146.341
R1873 vdd.n1454 vdd.n1175 146.341
R1874 vdd.n1454 vdd.n1169 146.341
R1875 vdd.n1466 vdd.n1169 146.341
R1876 vdd.n1466 vdd.n1165 146.341
R1877 vdd.n1472 vdd.n1165 146.341
R1878 vdd.n1472 vdd.n886 146.341
R1879 vdd.n1482 vdd.n886 146.341
R1880 vdd.n1482 vdd.n882 146.341
R1881 vdd.n1488 vdd.n882 146.341
R1882 vdd.n1488 vdd.n876 146.341
R1883 vdd.n1499 vdd.n876 146.341
R1884 vdd.n1499 vdd.n871 146.341
R1885 vdd.n1507 vdd.n871 146.341
R1886 vdd.n1507 vdd.n861 146.341
R1887 vdd.n1944 vdd.n861 146.341
R1888 vdd.n1420 vdd.n1196 146.341
R1889 vdd.n1420 vdd.n1229 146.341
R1890 vdd.n1233 vdd.n1232 146.341
R1891 vdd.n1235 vdd.n1234 146.341
R1892 vdd.n1239 vdd.n1238 146.341
R1893 vdd.n1241 vdd.n1240 146.341
R1894 vdd.n1245 vdd.n1244 146.341
R1895 vdd.n1247 vdd.n1246 146.341
R1896 vdd.n1251 vdd.n1250 146.341
R1897 vdd.n1253 vdd.n1252 146.341
R1898 vdd.n1259 vdd.n1258 146.341
R1899 vdd.n1261 vdd.n1260 146.341
R1900 vdd.n1265 vdd.n1264 146.341
R1901 vdd.n1267 vdd.n1266 146.341
R1902 vdd.n1271 vdd.n1270 146.341
R1903 vdd.n1273 vdd.n1272 146.341
R1904 vdd.n1277 vdd.n1276 146.341
R1905 vdd.n1279 vdd.n1278 146.341
R1906 vdd.n1283 vdd.n1282 146.341
R1907 vdd.n1285 vdd.n1284 146.341
R1908 vdd.n1357 vdd.n1288 146.341
R1909 vdd.n1290 vdd.n1289 146.341
R1910 vdd.n1294 vdd.n1293 146.341
R1911 vdd.n1296 vdd.n1295 146.341
R1912 vdd.n1300 vdd.n1299 146.341
R1913 vdd.n1302 vdd.n1301 146.341
R1914 vdd.n1306 vdd.n1305 146.341
R1915 vdd.n1308 vdd.n1307 146.341
R1916 vdd.n1312 vdd.n1311 146.341
R1917 vdd.n1314 vdd.n1313 146.341
R1918 vdd.n1318 vdd.n1317 146.341
R1919 vdd.n1319 vdd.n1227 146.341
R1920 vdd.n1429 vdd.n1192 146.341
R1921 vdd.n1429 vdd.n1185 146.341
R1922 vdd.n1440 vdd.n1185 146.341
R1923 vdd.n1440 vdd.n1181 146.341
R1924 vdd.n1446 vdd.n1181 146.341
R1925 vdd.n1446 vdd.n1174 146.341
R1926 vdd.n1457 vdd.n1174 146.341
R1927 vdd.n1457 vdd.n1170 146.341
R1928 vdd.n1464 vdd.n1170 146.341
R1929 vdd.n1464 vdd.n1163 146.341
R1930 vdd.n1474 vdd.n1163 146.341
R1931 vdd.n1474 vdd.n889 146.341
R1932 vdd.n1480 vdd.n889 146.341
R1933 vdd.n1480 vdd.n881 146.341
R1934 vdd.n1491 vdd.n881 146.341
R1935 vdd.n1491 vdd.n877 146.341
R1936 vdd.n1497 vdd.n877 146.341
R1937 vdd.n1497 vdd.n869 146.341
R1938 vdd.n1510 vdd.n869 146.341
R1939 vdd.n1510 vdd.n864 146.341
R1940 vdd.n1942 vdd.n864 146.341
R1941 vdd.n863 vdd.n839 141.707
R1942 vdd.n2840 vdd.n484 141.707
R1943 vdd.n1791 vdd.t66 127.284
R1944 vdd.n755 vdd.t54 127.284
R1945 vdd.n1765 vdd.t19 127.284
R1946 vdd.n747 vdd.t84 127.284
R1947 vdd.n2536 vdd.t37 127.284
R1948 vdd.n2536 vdd.t38 127.284
R1949 vdd.n2256 vdd.t76 127.284
R1950 vdd.n622 vdd.t58 127.284
R1951 vdd.n2253 vdd.t63 127.284
R1952 vdd.n589 vdd.t68 127.284
R1953 vdd.n817 vdd.t72 127.284
R1954 vdd.n817 vdd.t73 127.284
R1955 vdd.n22 vdd.n20 117.314
R1956 vdd.n17 vdd.n15 117.314
R1957 vdd.n27 vdd.n26 116.927
R1958 vdd.n24 vdd.n23 116.927
R1959 vdd.n22 vdd.n21 116.927
R1960 vdd.n17 vdd.n16 116.927
R1961 vdd.n19 vdd.n18 116.927
R1962 vdd.n27 vdd.n25 116.927
R1963 vdd.n1792 vdd.t65 111.188
R1964 vdd.n756 vdd.t55 111.188
R1965 vdd.n1766 vdd.t18 111.188
R1966 vdd.n748 vdd.t85 111.188
R1967 vdd.n2257 vdd.t75 111.188
R1968 vdd.n623 vdd.t59 111.188
R1969 vdd.n2254 vdd.t62 111.188
R1970 vdd.n590 vdd.t69 111.188
R1971 vdd.n2479 vdd.n701 99.5127
R1972 vdd.n2483 vdd.n701 99.5127
R1973 vdd.n2483 vdd.n693 99.5127
R1974 vdd.n2491 vdd.n693 99.5127
R1975 vdd.n2491 vdd.n691 99.5127
R1976 vdd.n2495 vdd.n691 99.5127
R1977 vdd.n2495 vdd.n680 99.5127
R1978 vdd.n2503 vdd.n680 99.5127
R1979 vdd.n2503 vdd.n678 99.5127
R1980 vdd.n2507 vdd.n678 99.5127
R1981 vdd.n2507 vdd.n669 99.5127
R1982 vdd.n2515 vdd.n669 99.5127
R1983 vdd.n2515 vdd.n667 99.5127
R1984 vdd.n2519 vdd.n667 99.5127
R1985 vdd.n2519 vdd.n657 99.5127
R1986 vdd.n2527 vdd.n657 99.5127
R1987 vdd.n2527 vdd.n655 99.5127
R1988 vdd.n2531 vdd.n655 99.5127
R1989 vdd.n2531 vdd.n646 99.5127
R1990 vdd.n2541 vdd.n646 99.5127
R1991 vdd.n2541 vdd.n644 99.5127
R1992 vdd.n2545 vdd.n644 99.5127
R1993 vdd.n2545 vdd.n632 99.5127
R1994 vdd.n2598 vdd.n632 99.5127
R1995 vdd.n2598 vdd.n630 99.5127
R1996 vdd.n2602 vdd.n630 99.5127
R1997 vdd.n2602 vdd.n598 99.5127
R1998 vdd.n2672 vdd.n598 99.5127
R1999 vdd.n2668 vdd.n599 99.5127
R2000 vdd.n2666 vdd.n2665 99.5127
R2001 vdd.n2663 vdd.n603 99.5127
R2002 vdd.n2659 vdd.n2658 99.5127
R2003 vdd.n2656 vdd.n606 99.5127
R2004 vdd.n2652 vdd.n2651 99.5127
R2005 vdd.n2649 vdd.n609 99.5127
R2006 vdd.n2645 vdd.n2644 99.5127
R2007 vdd.n2642 vdd.n2640 99.5127
R2008 vdd.n2638 vdd.n612 99.5127
R2009 vdd.n2634 vdd.n2633 99.5127
R2010 vdd.n2631 vdd.n615 99.5127
R2011 vdd.n2627 vdd.n2626 99.5127
R2012 vdd.n2624 vdd.n618 99.5127
R2013 vdd.n2620 vdd.n2619 99.5127
R2014 vdd.n2617 vdd.n621 99.5127
R2015 vdd.n2612 vdd.n2611 99.5127
R2016 vdd.n2399 vdd.n704 99.5127
R2017 vdd.n2399 vdd.n699 99.5127
R2018 vdd.n2396 vdd.n699 99.5127
R2019 vdd.n2396 vdd.n694 99.5127
R2020 vdd.n2343 vdd.n694 99.5127
R2021 vdd.n2343 vdd.n688 99.5127
R2022 vdd.n2346 vdd.n688 99.5127
R2023 vdd.n2346 vdd.n681 99.5127
R2024 vdd.n2349 vdd.n681 99.5127
R2025 vdd.n2349 vdd.n676 99.5127
R2026 vdd.n2352 vdd.n676 99.5127
R2027 vdd.n2352 vdd.n671 99.5127
R2028 vdd.n2355 vdd.n671 99.5127
R2029 vdd.n2355 vdd.n665 99.5127
R2030 vdd.n2373 vdd.n665 99.5127
R2031 vdd.n2373 vdd.n658 99.5127
R2032 vdd.n2369 vdd.n658 99.5127
R2033 vdd.n2369 vdd.n653 99.5127
R2034 vdd.n2366 vdd.n653 99.5127
R2035 vdd.n2366 vdd.n648 99.5127
R2036 vdd.n2363 vdd.n648 99.5127
R2037 vdd.n2363 vdd.n642 99.5127
R2038 vdd.n2360 vdd.n642 99.5127
R2039 vdd.n2360 vdd.n634 99.5127
R2040 vdd.n634 vdd.n627 99.5127
R2041 vdd.n2604 vdd.n627 99.5127
R2042 vdd.n2605 vdd.n2604 99.5127
R2043 vdd.n2605 vdd.n596 99.5127
R2044 vdd.n2469 vdd.n2252 99.5127
R2045 vdd.n2465 vdd.n2252 99.5127
R2046 vdd.n2463 vdd.n2462 99.5127
R2047 vdd.n2459 vdd.n2458 99.5127
R2048 vdd.n2455 vdd.n2454 99.5127
R2049 vdd.n2451 vdd.n2450 99.5127
R2050 vdd.n2447 vdd.n2446 99.5127
R2051 vdd.n2443 vdd.n2442 99.5127
R2052 vdd.n2439 vdd.n2438 99.5127
R2053 vdd.n2435 vdd.n2434 99.5127
R2054 vdd.n2431 vdd.n2430 99.5127
R2055 vdd.n2427 vdd.n2426 99.5127
R2056 vdd.n2423 vdd.n2422 99.5127
R2057 vdd.n2419 vdd.n2418 99.5127
R2058 vdd.n2415 vdd.n2414 99.5127
R2059 vdd.n2411 vdd.n2410 99.5127
R2060 vdd.n2406 vdd.n2405 99.5127
R2061 vdd.n2217 vdd.n745 99.5127
R2062 vdd.n2213 vdd.n2212 99.5127
R2063 vdd.n2209 vdd.n2208 99.5127
R2064 vdd.n2205 vdd.n2204 99.5127
R2065 vdd.n2201 vdd.n2200 99.5127
R2066 vdd.n2197 vdd.n2196 99.5127
R2067 vdd.n2193 vdd.n2192 99.5127
R2068 vdd.n2189 vdd.n2188 99.5127
R2069 vdd.n2185 vdd.n2184 99.5127
R2070 vdd.n2181 vdd.n2180 99.5127
R2071 vdd.n2177 vdd.n2176 99.5127
R2072 vdd.n2173 vdd.n2172 99.5127
R2073 vdd.n2169 vdd.n2168 99.5127
R2074 vdd.n2165 vdd.n2164 99.5127
R2075 vdd.n2161 vdd.n2160 99.5127
R2076 vdd.n2157 vdd.n2156 99.5127
R2077 vdd.n2152 vdd.n2151 99.5127
R2078 vdd.n1890 vdd.n840 99.5127
R2079 vdd.n1890 vdd.n834 99.5127
R2080 vdd.n1887 vdd.n834 99.5127
R2081 vdd.n1887 vdd.n828 99.5127
R2082 vdd.n1884 vdd.n828 99.5127
R2083 vdd.n1884 vdd.n821 99.5127
R2084 vdd.n1881 vdd.n821 99.5127
R2085 vdd.n1881 vdd.n814 99.5127
R2086 vdd.n1878 vdd.n814 99.5127
R2087 vdd.n1878 vdd.n809 99.5127
R2088 vdd.n1875 vdd.n809 99.5127
R2089 vdd.n1875 vdd.n803 99.5127
R2090 vdd.n1872 vdd.n803 99.5127
R2091 vdd.n1872 vdd.n796 99.5127
R2092 vdd.n1786 vdd.n796 99.5127
R2093 vdd.n1786 vdd.n790 99.5127
R2094 vdd.n1783 vdd.n790 99.5127
R2095 vdd.n1783 vdd.n785 99.5127
R2096 vdd.n1780 vdd.n785 99.5127
R2097 vdd.n1780 vdd.n780 99.5127
R2098 vdd.n1777 vdd.n780 99.5127
R2099 vdd.n1777 vdd.n774 99.5127
R2100 vdd.n1774 vdd.n774 99.5127
R2101 vdd.n1774 vdd.n767 99.5127
R2102 vdd.n1771 vdd.n767 99.5127
R2103 vdd.n1771 vdd.n760 99.5127
R2104 vdd.n760 vdd.n750 99.5127
R2105 vdd.n2147 vdd.n750 99.5127
R2106 vdd.n1725 vdd.n1723 99.5127
R2107 vdd.n1729 vdd.n1723 99.5127
R2108 vdd.n1733 vdd.n1731 99.5127
R2109 vdd.n1737 vdd.n1721 99.5127
R2110 vdd.n1741 vdd.n1739 99.5127
R2111 vdd.n1745 vdd.n1719 99.5127
R2112 vdd.n1749 vdd.n1747 99.5127
R2113 vdd.n1753 vdd.n1717 99.5127
R2114 vdd.n1756 vdd.n1755 99.5127
R2115 vdd.n1926 vdd.n1924 99.5127
R2116 vdd.n1922 vdd.n1758 99.5127
R2117 vdd.n1918 vdd.n1916 99.5127
R2118 vdd.n1914 vdd.n1760 99.5127
R2119 vdd.n1910 vdd.n1908 99.5127
R2120 vdd.n1906 vdd.n1762 99.5127
R2121 vdd.n1902 vdd.n1900 99.5127
R2122 vdd.n1898 vdd.n1764 99.5127
R2123 vdd.n1990 vdd.n836 99.5127
R2124 vdd.n1994 vdd.n836 99.5127
R2125 vdd.n1994 vdd.n826 99.5127
R2126 vdd.n2002 vdd.n826 99.5127
R2127 vdd.n2002 vdd.n824 99.5127
R2128 vdd.n2006 vdd.n824 99.5127
R2129 vdd.n2006 vdd.n813 99.5127
R2130 vdd.n2015 vdd.n813 99.5127
R2131 vdd.n2015 vdd.n811 99.5127
R2132 vdd.n2019 vdd.n811 99.5127
R2133 vdd.n2019 vdd.n801 99.5127
R2134 vdd.n2027 vdd.n801 99.5127
R2135 vdd.n2027 vdd.n799 99.5127
R2136 vdd.n2031 vdd.n799 99.5127
R2137 vdd.n2031 vdd.n789 99.5127
R2138 vdd.n2039 vdd.n789 99.5127
R2139 vdd.n2039 vdd.n787 99.5127
R2140 vdd.n2043 vdd.n787 99.5127
R2141 vdd.n2043 vdd.n778 99.5127
R2142 vdd.n2051 vdd.n778 99.5127
R2143 vdd.n2051 vdd.n776 99.5127
R2144 vdd.n2055 vdd.n776 99.5127
R2145 vdd.n2055 vdd.n765 99.5127
R2146 vdd.n2065 vdd.n765 99.5127
R2147 vdd.n2065 vdd.n762 99.5127
R2148 vdd.n2070 vdd.n762 99.5127
R2149 vdd.n2070 vdd.n763 99.5127
R2150 vdd.n763 vdd.n744 99.5127
R2151 vdd.n2588 vdd.n2587 99.5127
R2152 vdd.n2585 vdd.n2551 99.5127
R2153 vdd.n2581 vdd.n2580 99.5127
R2154 vdd.n2578 vdd.n2554 99.5127
R2155 vdd.n2574 vdd.n2573 99.5127
R2156 vdd.n2571 vdd.n2557 99.5127
R2157 vdd.n2567 vdd.n2566 99.5127
R2158 vdd.n2564 vdd.n2561 99.5127
R2159 vdd.n2705 vdd.n577 99.5127
R2160 vdd.n2703 vdd.n2702 99.5127
R2161 vdd.n2700 vdd.n579 99.5127
R2162 vdd.n2696 vdd.n2695 99.5127
R2163 vdd.n2693 vdd.n582 99.5127
R2164 vdd.n2689 vdd.n2688 99.5127
R2165 vdd.n2686 vdd.n585 99.5127
R2166 vdd.n2682 vdd.n2681 99.5127
R2167 vdd.n2679 vdd.n588 99.5127
R2168 vdd.n2323 vdd.n705 99.5127
R2169 vdd.n2323 vdd.n700 99.5127
R2170 vdd.n2394 vdd.n700 99.5127
R2171 vdd.n2394 vdd.n695 99.5127
R2172 vdd.n2390 vdd.n695 99.5127
R2173 vdd.n2390 vdd.n689 99.5127
R2174 vdd.n2387 vdd.n689 99.5127
R2175 vdd.n2387 vdd.n682 99.5127
R2176 vdd.n2384 vdd.n682 99.5127
R2177 vdd.n2384 vdd.n677 99.5127
R2178 vdd.n2381 vdd.n677 99.5127
R2179 vdd.n2381 vdd.n672 99.5127
R2180 vdd.n2378 vdd.n672 99.5127
R2181 vdd.n2378 vdd.n666 99.5127
R2182 vdd.n2375 vdd.n666 99.5127
R2183 vdd.n2375 vdd.n659 99.5127
R2184 vdd.n2340 vdd.n659 99.5127
R2185 vdd.n2340 vdd.n654 99.5127
R2186 vdd.n2337 vdd.n654 99.5127
R2187 vdd.n2337 vdd.n649 99.5127
R2188 vdd.n2334 vdd.n649 99.5127
R2189 vdd.n2334 vdd.n643 99.5127
R2190 vdd.n2331 vdd.n643 99.5127
R2191 vdd.n2331 vdd.n635 99.5127
R2192 vdd.n2328 vdd.n635 99.5127
R2193 vdd.n2328 vdd.n628 99.5127
R2194 vdd.n628 vdd.n594 99.5127
R2195 vdd.n2674 vdd.n594 99.5127
R2196 vdd.n2473 vdd.n708 99.5127
R2197 vdd.n2261 vdd.n2260 99.5127
R2198 vdd.n2265 vdd.n2264 99.5127
R2199 vdd.n2269 vdd.n2268 99.5127
R2200 vdd.n2273 vdd.n2272 99.5127
R2201 vdd.n2277 vdd.n2276 99.5127
R2202 vdd.n2281 vdd.n2280 99.5127
R2203 vdd.n2285 vdd.n2284 99.5127
R2204 vdd.n2289 vdd.n2288 99.5127
R2205 vdd.n2293 vdd.n2292 99.5127
R2206 vdd.n2297 vdd.n2296 99.5127
R2207 vdd.n2301 vdd.n2300 99.5127
R2208 vdd.n2305 vdd.n2304 99.5127
R2209 vdd.n2309 vdd.n2308 99.5127
R2210 vdd.n2313 vdd.n2312 99.5127
R2211 vdd.n2317 vdd.n2316 99.5127
R2212 vdd.n2319 vdd.n2251 99.5127
R2213 vdd.n2477 vdd.n698 99.5127
R2214 vdd.n2485 vdd.n698 99.5127
R2215 vdd.n2485 vdd.n696 99.5127
R2216 vdd.n2489 vdd.n696 99.5127
R2217 vdd.n2489 vdd.n686 99.5127
R2218 vdd.n2497 vdd.n686 99.5127
R2219 vdd.n2497 vdd.n684 99.5127
R2220 vdd.n2501 vdd.n684 99.5127
R2221 vdd.n2501 vdd.n675 99.5127
R2222 vdd.n2509 vdd.n675 99.5127
R2223 vdd.n2509 vdd.n673 99.5127
R2224 vdd.n2513 vdd.n673 99.5127
R2225 vdd.n2513 vdd.n663 99.5127
R2226 vdd.n2521 vdd.n663 99.5127
R2227 vdd.n2521 vdd.n661 99.5127
R2228 vdd.n2525 vdd.n661 99.5127
R2229 vdd.n2525 vdd.n652 99.5127
R2230 vdd.n2533 vdd.n652 99.5127
R2231 vdd.n2533 vdd.n650 99.5127
R2232 vdd.n2539 vdd.n650 99.5127
R2233 vdd.n2539 vdd.n640 99.5127
R2234 vdd.n2547 vdd.n640 99.5127
R2235 vdd.n2547 vdd.n637 99.5127
R2236 vdd.n2596 vdd.n637 99.5127
R2237 vdd.n2596 vdd.n638 99.5127
R2238 vdd.n638 vdd.n629 99.5127
R2239 vdd.n2591 vdd.n629 99.5127
R2240 vdd.n2591 vdd.n597 99.5127
R2241 vdd.n2141 vdd.n2140 99.5127
R2242 vdd.n2137 vdd.n2136 99.5127
R2243 vdd.n2133 vdd.n2132 99.5127
R2244 vdd.n2129 vdd.n2128 99.5127
R2245 vdd.n2125 vdd.n2124 99.5127
R2246 vdd.n2121 vdd.n2120 99.5127
R2247 vdd.n2117 vdd.n2116 99.5127
R2248 vdd.n2113 vdd.n2112 99.5127
R2249 vdd.n2109 vdd.n2108 99.5127
R2250 vdd.n2105 vdd.n2104 99.5127
R2251 vdd.n2101 vdd.n2100 99.5127
R2252 vdd.n2097 vdd.n2096 99.5127
R2253 vdd.n2093 vdd.n2092 99.5127
R2254 vdd.n2089 vdd.n2088 99.5127
R2255 vdd.n2085 vdd.n2084 99.5127
R2256 vdd.n2081 vdd.n2080 99.5127
R2257 vdd.n2077 vdd.n726 99.5127
R2258 vdd.n1834 vdd.n841 99.5127
R2259 vdd.n1834 vdd.n835 99.5127
R2260 vdd.n1837 vdd.n835 99.5127
R2261 vdd.n1837 vdd.n829 99.5127
R2262 vdd.n1840 vdd.n829 99.5127
R2263 vdd.n1840 vdd.n822 99.5127
R2264 vdd.n1843 vdd.n822 99.5127
R2265 vdd.n1843 vdd.n815 99.5127
R2266 vdd.n1846 vdd.n815 99.5127
R2267 vdd.n1846 vdd.n810 99.5127
R2268 vdd.n1849 vdd.n810 99.5127
R2269 vdd.n1849 vdd.n804 99.5127
R2270 vdd.n1870 vdd.n804 99.5127
R2271 vdd.n1870 vdd.n797 99.5127
R2272 vdd.n1866 vdd.n797 99.5127
R2273 vdd.n1866 vdd.n791 99.5127
R2274 vdd.n1863 vdd.n791 99.5127
R2275 vdd.n1863 vdd.n786 99.5127
R2276 vdd.n1860 vdd.n786 99.5127
R2277 vdd.n1860 vdd.n781 99.5127
R2278 vdd.n1857 vdd.n781 99.5127
R2279 vdd.n1857 vdd.n775 99.5127
R2280 vdd.n1854 vdd.n775 99.5127
R2281 vdd.n1854 vdd.n768 99.5127
R2282 vdd.n768 vdd.n759 99.5127
R2283 vdd.n2072 vdd.n759 99.5127
R2284 vdd.n2073 vdd.n2072 99.5127
R2285 vdd.n2073 vdd.n751 99.5127
R2286 vdd.n1984 vdd.n1982 99.5127
R2287 vdd.n1980 vdd.n844 99.5127
R2288 vdd.n1976 vdd.n1974 99.5127
R2289 vdd.n1972 vdd.n846 99.5127
R2290 vdd.n1968 vdd.n1966 99.5127
R2291 vdd.n1964 vdd.n848 99.5127
R2292 vdd.n1960 vdd.n1958 99.5127
R2293 vdd.n1956 vdd.n850 99.5127
R2294 vdd.n1798 vdd.n852 99.5127
R2295 vdd.n1803 vdd.n1800 99.5127
R2296 vdd.n1807 vdd.n1805 99.5127
R2297 vdd.n1811 vdd.n1796 99.5127
R2298 vdd.n1815 vdd.n1813 99.5127
R2299 vdd.n1819 vdd.n1794 99.5127
R2300 vdd.n1823 vdd.n1821 99.5127
R2301 vdd.n1828 vdd.n1790 99.5127
R2302 vdd.n1831 vdd.n1830 99.5127
R2303 vdd.n1988 vdd.n832 99.5127
R2304 vdd.n1996 vdd.n832 99.5127
R2305 vdd.n1996 vdd.n830 99.5127
R2306 vdd.n2000 vdd.n830 99.5127
R2307 vdd.n2000 vdd.n819 99.5127
R2308 vdd.n2008 vdd.n819 99.5127
R2309 vdd.n2008 vdd.n816 99.5127
R2310 vdd.n2013 vdd.n816 99.5127
R2311 vdd.n2013 vdd.n807 99.5127
R2312 vdd.n2021 vdd.n807 99.5127
R2313 vdd.n2021 vdd.n805 99.5127
R2314 vdd.n2025 vdd.n805 99.5127
R2315 vdd.n2025 vdd.n795 99.5127
R2316 vdd.n2033 vdd.n795 99.5127
R2317 vdd.n2033 vdd.n793 99.5127
R2318 vdd.n2037 vdd.n793 99.5127
R2319 vdd.n2037 vdd.n784 99.5127
R2320 vdd.n2045 vdd.n784 99.5127
R2321 vdd.n2045 vdd.n782 99.5127
R2322 vdd.n2049 vdd.n782 99.5127
R2323 vdd.n2049 vdd.n772 99.5127
R2324 vdd.n2057 vdd.n772 99.5127
R2325 vdd.n2057 vdd.n769 99.5127
R2326 vdd.n2063 vdd.n769 99.5127
R2327 vdd.n2063 vdd.n770 99.5127
R2328 vdd.n770 vdd.n761 99.5127
R2329 vdd.n761 vdd.n752 99.5127
R2330 vdd.n2145 vdd.n752 99.5127
R2331 vdd.n9 vdd.n7 98.9633
R2332 vdd.n2 vdd.n0 98.9633
R2333 vdd.n9 vdd.n8 98.6055
R2334 vdd.n11 vdd.n10 98.6055
R2335 vdd.n13 vdd.n12 98.6055
R2336 vdd.n6 vdd.n5 98.6055
R2337 vdd.n4 vdd.n3 98.6055
R2338 vdd.n2 vdd.n1 98.6055
R2339 vdd.t15 vdd.n267 85.8723
R2340 vdd.t104 vdd.n220 85.8723
R2341 vdd.t133 vdd.n177 85.8723
R2342 vdd.t142 vdd.n130 85.8723
R2343 vdd.t111 vdd.n88 85.8723
R2344 vdd.t132 vdd.n41 85.8723
R2345 vdd.t121 vdd.n1082 85.8723
R2346 vdd.t102 vdd.n1129 85.8723
R2347 vdd.t138 vdd.n992 85.8723
R2348 vdd.t112 vdd.n1039 85.8723
R2349 vdd.t3 vdd.n903 85.8723
R2350 vdd.t193 vdd.n950 85.8723
R2351 vdd.n2537 vdd.n2536 78.546
R2352 vdd.n2011 vdd.n817 78.546
R2353 vdd.n254 vdd.n253 75.1835
R2354 vdd.n252 vdd.n251 75.1835
R2355 vdd.n250 vdd.n249 75.1835
R2356 vdd.n164 vdd.n163 75.1835
R2357 vdd.n162 vdd.n161 75.1835
R2358 vdd.n160 vdd.n159 75.1835
R2359 vdd.n75 vdd.n74 75.1835
R2360 vdd.n73 vdd.n72 75.1835
R2361 vdd.n71 vdd.n70 75.1835
R2362 vdd.n1112 vdd.n1111 75.1835
R2363 vdd.n1114 vdd.n1113 75.1835
R2364 vdd.n1116 vdd.n1115 75.1835
R2365 vdd.n1022 vdd.n1021 75.1835
R2366 vdd.n1024 vdd.n1023 75.1835
R2367 vdd.n1026 vdd.n1025 75.1835
R2368 vdd.n933 vdd.n932 75.1835
R2369 vdd.n935 vdd.n934 75.1835
R2370 vdd.n937 vdd.n936 75.1835
R2371 vdd.n2472 vdd.n2471 72.8958
R2372 vdd.n2471 vdd.n2235 72.8958
R2373 vdd.n2471 vdd.n2236 72.8958
R2374 vdd.n2471 vdd.n2237 72.8958
R2375 vdd.n2471 vdd.n2238 72.8958
R2376 vdd.n2471 vdd.n2239 72.8958
R2377 vdd.n2471 vdd.n2240 72.8958
R2378 vdd.n2471 vdd.n2241 72.8958
R2379 vdd.n2471 vdd.n2242 72.8958
R2380 vdd.n2471 vdd.n2243 72.8958
R2381 vdd.n2471 vdd.n2244 72.8958
R2382 vdd.n2471 vdd.n2245 72.8958
R2383 vdd.n2471 vdd.n2246 72.8958
R2384 vdd.n2471 vdd.n2247 72.8958
R2385 vdd.n2471 vdd.n2248 72.8958
R2386 vdd.n2471 vdd.n2249 72.8958
R2387 vdd.n2471 vdd.n2250 72.8958
R2388 vdd.n593 vdd.n484 72.8958
R2389 vdd.n2680 vdd.n484 72.8958
R2390 vdd.n587 vdd.n484 72.8958
R2391 vdd.n2687 vdd.n484 72.8958
R2392 vdd.n584 vdd.n484 72.8958
R2393 vdd.n2694 vdd.n484 72.8958
R2394 vdd.n581 vdd.n484 72.8958
R2395 vdd.n2701 vdd.n484 72.8958
R2396 vdd.n2704 vdd.n484 72.8958
R2397 vdd.n2560 vdd.n484 72.8958
R2398 vdd.n2565 vdd.n484 72.8958
R2399 vdd.n2559 vdd.n484 72.8958
R2400 vdd.n2572 vdd.n484 72.8958
R2401 vdd.n2556 vdd.n484 72.8958
R2402 vdd.n2579 vdd.n484 72.8958
R2403 vdd.n2553 vdd.n484 72.8958
R2404 vdd.n2586 vdd.n484 72.8958
R2405 vdd.n1724 vdd.n839 72.8958
R2406 vdd.n1730 vdd.n839 72.8958
R2407 vdd.n1732 vdd.n839 72.8958
R2408 vdd.n1738 vdd.n839 72.8958
R2409 vdd.n1740 vdd.n839 72.8958
R2410 vdd.n1746 vdd.n839 72.8958
R2411 vdd.n1748 vdd.n839 72.8958
R2412 vdd.n1754 vdd.n839 72.8958
R2413 vdd.n1925 vdd.n839 72.8958
R2414 vdd.n1923 vdd.n839 72.8958
R2415 vdd.n1917 vdd.n839 72.8958
R2416 vdd.n1915 vdd.n839 72.8958
R2417 vdd.n1909 vdd.n839 72.8958
R2418 vdd.n1907 vdd.n839 72.8958
R2419 vdd.n1901 vdd.n839 72.8958
R2420 vdd.n1899 vdd.n839 72.8958
R2421 vdd.n1893 vdd.n839 72.8958
R2422 vdd.n2218 vdd.n727 72.8958
R2423 vdd.n2218 vdd.n728 72.8958
R2424 vdd.n2218 vdd.n729 72.8958
R2425 vdd.n2218 vdd.n730 72.8958
R2426 vdd.n2218 vdd.n731 72.8958
R2427 vdd.n2218 vdd.n732 72.8958
R2428 vdd.n2218 vdd.n733 72.8958
R2429 vdd.n2218 vdd.n734 72.8958
R2430 vdd.n2218 vdd.n735 72.8958
R2431 vdd.n2218 vdd.n736 72.8958
R2432 vdd.n2218 vdd.n737 72.8958
R2433 vdd.n2218 vdd.n738 72.8958
R2434 vdd.n2218 vdd.n739 72.8958
R2435 vdd.n2218 vdd.n740 72.8958
R2436 vdd.n2218 vdd.n741 72.8958
R2437 vdd.n2218 vdd.n742 72.8958
R2438 vdd.n2218 vdd.n743 72.8958
R2439 vdd.n2471 vdd.n2470 72.8958
R2440 vdd.n2471 vdd.n2219 72.8958
R2441 vdd.n2471 vdd.n2220 72.8958
R2442 vdd.n2471 vdd.n2221 72.8958
R2443 vdd.n2471 vdd.n2222 72.8958
R2444 vdd.n2471 vdd.n2223 72.8958
R2445 vdd.n2471 vdd.n2224 72.8958
R2446 vdd.n2471 vdd.n2225 72.8958
R2447 vdd.n2471 vdd.n2226 72.8958
R2448 vdd.n2471 vdd.n2227 72.8958
R2449 vdd.n2471 vdd.n2228 72.8958
R2450 vdd.n2471 vdd.n2229 72.8958
R2451 vdd.n2471 vdd.n2230 72.8958
R2452 vdd.n2471 vdd.n2231 72.8958
R2453 vdd.n2471 vdd.n2232 72.8958
R2454 vdd.n2471 vdd.n2233 72.8958
R2455 vdd.n2471 vdd.n2234 72.8958
R2456 vdd.n2610 vdd.n484 72.8958
R2457 vdd.n625 vdd.n484 72.8958
R2458 vdd.n2618 vdd.n484 72.8958
R2459 vdd.n620 vdd.n484 72.8958
R2460 vdd.n2625 vdd.n484 72.8958
R2461 vdd.n617 vdd.n484 72.8958
R2462 vdd.n2632 vdd.n484 72.8958
R2463 vdd.n614 vdd.n484 72.8958
R2464 vdd.n2639 vdd.n484 72.8958
R2465 vdd.n2643 vdd.n484 72.8958
R2466 vdd.n611 vdd.n484 72.8958
R2467 vdd.n2650 vdd.n484 72.8958
R2468 vdd.n608 vdd.n484 72.8958
R2469 vdd.n2657 vdd.n484 72.8958
R2470 vdd.n605 vdd.n484 72.8958
R2471 vdd.n2664 vdd.n484 72.8958
R2472 vdd.n2667 vdd.n484 72.8958
R2473 vdd.n2218 vdd.n725 72.8958
R2474 vdd.n2218 vdd.n724 72.8958
R2475 vdd.n2218 vdd.n723 72.8958
R2476 vdd.n2218 vdd.n722 72.8958
R2477 vdd.n2218 vdd.n721 72.8958
R2478 vdd.n2218 vdd.n720 72.8958
R2479 vdd.n2218 vdd.n719 72.8958
R2480 vdd.n2218 vdd.n718 72.8958
R2481 vdd.n2218 vdd.n717 72.8958
R2482 vdd.n2218 vdd.n716 72.8958
R2483 vdd.n2218 vdd.n715 72.8958
R2484 vdd.n2218 vdd.n714 72.8958
R2485 vdd.n2218 vdd.n713 72.8958
R2486 vdd.n2218 vdd.n712 72.8958
R2487 vdd.n2218 vdd.n711 72.8958
R2488 vdd.n2218 vdd.n710 72.8958
R2489 vdd.n2218 vdd.n709 72.8958
R2490 vdd.n1983 vdd.n839 72.8958
R2491 vdd.n1981 vdd.n839 72.8958
R2492 vdd.n1975 vdd.n839 72.8958
R2493 vdd.n1973 vdd.n839 72.8958
R2494 vdd.n1967 vdd.n839 72.8958
R2495 vdd.n1965 vdd.n839 72.8958
R2496 vdd.n1959 vdd.n839 72.8958
R2497 vdd.n1957 vdd.n839 72.8958
R2498 vdd.n851 vdd.n839 72.8958
R2499 vdd.n1799 vdd.n839 72.8958
R2500 vdd.n1804 vdd.n839 72.8958
R2501 vdd.n1806 vdd.n839 72.8958
R2502 vdd.n1812 vdd.n839 72.8958
R2503 vdd.n1814 vdd.n839 72.8958
R2504 vdd.n1820 vdd.n839 72.8958
R2505 vdd.n1822 vdd.n839 72.8958
R2506 vdd.n1829 vdd.n839 72.8958
R2507 vdd.n1422 vdd.n1421 66.2847
R2508 vdd.n1421 vdd.n1197 66.2847
R2509 vdd.n1421 vdd.n1198 66.2847
R2510 vdd.n1421 vdd.n1199 66.2847
R2511 vdd.n1421 vdd.n1200 66.2847
R2512 vdd.n1421 vdd.n1201 66.2847
R2513 vdd.n1421 vdd.n1202 66.2847
R2514 vdd.n1421 vdd.n1203 66.2847
R2515 vdd.n1421 vdd.n1204 66.2847
R2516 vdd.n1421 vdd.n1205 66.2847
R2517 vdd.n1421 vdd.n1206 66.2847
R2518 vdd.n1421 vdd.n1207 66.2847
R2519 vdd.n1421 vdd.n1208 66.2847
R2520 vdd.n1421 vdd.n1209 66.2847
R2521 vdd.n1421 vdd.n1210 66.2847
R2522 vdd.n1421 vdd.n1211 66.2847
R2523 vdd.n1421 vdd.n1212 66.2847
R2524 vdd.n1421 vdd.n1213 66.2847
R2525 vdd.n1421 vdd.n1214 66.2847
R2526 vdd.n1421 vdd.n1215 66.2847
R2527 vdd.n1421 vdd.n1216 66.2847
R2528 vdd.n1421 vdd.n1217 66.2847
R2529 vdd.n1421 vdd.n1218 66.2847
R2530 vdd.n1421 vdd.n1219 66.2847
R2531 vdd.n1421 vdd.n1220 66.2847
R2532 vdd.n1421 vdd.n1221 66.2847
R2533 vdd.n1421 vdd.n1222 66.2847
R2534 vdd.n1421 vdd.n1223 66.2847
R2535 vdd.n1421 vdd.n1224 66.2847
R2536 vdd.n1421 vdd.n1225 66.2847
R2537 vdd.n1421 vdd.n1226 66.2847
R2538 vdd.n863 vdd.n860 66.2847
R2539 vdd.n1614 vdd.n863 66.2847
R2540 vdd.n1619 vdd.n863 66.2847
R2541 vdd.n1624 vdd.n863 66.2847
R2542 vdd.n1612 vdd.n863 66.2847
R2543 vdd.n1631 vdd.n863 66.2847
R2544 vdd.n1604 vdd.n863 66.2847
R2545 vdd.n1638 vdd.n863 66.2847
R2546 vdd.n1597 vdd.n863 66.2847
R2547 vdd.n1645 vdd.n863 66.2847
R2548 vdd.n1591 vdd.n863 66.2847
R2549 vdd.n1586 vdd.n863 66.2847
R2550 vdd.n1656 vdd.n863 66.2847
R2551 vdd.n1578 vdd.n863 66.2847
R2552 vdd.n1663 vdd.n863 66.2847
R2553 vdd.n1571 vdd.n863 66.2847
R2554 vdd.n1670 vdd.n863 66.2847
R2555 vdd.n1564 vdd.n863 66.2847
R2556 vdd.n1677 vdd.n863 66.2847
R2557 vdd.n1557 vdd.n863 66.2847
R2558 vdd.n1684 vdd.n863 66.2847
R2559 vdd.n1551 vdd.n863 66.2847
R2560 vdd.n1546 vdd.n863 66.2847
R2561 vdd.n1695 vdd.n863 66.2847
R2562 vdd.n1538 vdd.n863 66.2847
R2563 vdd.n1702 vdd.n863 66.2847
R2564 vdd.n1531 vdd.n863 66.2847
R2565 vdd.n1709 vdd.n863 66.2847
R2566 vdd.n1712 vdd.n863 66.2847
R2567 vdd.n1522 vdd.n863 66.2847
R2568 vdd.n1934 vdd.n863 66.2847
R2569 vdd.n1516 vdd.n863 66.2847
R2570 vdd.n2841 vdd.n2840 66.2847
R2571 vdd.n2840 vdd.n485 66.2847
R2572 vdd.n2840 vdd.n486 66.2847
R2573 vdd.n2840 vdd.n487 66.2847
R2574 vdd.n2840 vdd.n488 66.2847
R2575 vdd.n2840 vdd.n489 66.2847
R2576 vdd.n2840 vdd.n490 66.2847
R2577 vdd.n2840 vdd.n491 66.2847
R2578 vdd.n2840 vdd.n492 66.2847
R2579 vdd.n2840 vdd.n493 66.2847
R2580 vdd.n2840 vdd.n494 66.2847
R2581 vdd.n2840 vdd.n495 66.2847
R2582 vdd.n2840 vdd.n496 66.2847
R2583 vdd.n2840 vdd.n497 66.2847
R2584 vdd.n2840 vdd.n498 66.2847
R2585 vdd.n2840 vdd.n499 66.2847
R2586 vdd.n2840 vdd.n500 66.2847
R2587 vdd.n2840 vdd.n501 66.2847
R2588 vdd.n2840 vdd.n502 66.2847
R2589 vdd.n2840 vdd.n503 66.2847
R2590 vdd.n2840 vdd.n504 66.2847
R2591 vdd.n2840 vdd.n505 66.2847
R2592 vdd.n2840 vdd.n506 66.2847
R2593 vdd.n2840 vdd.n507 66.2847
R2594 vdd.n2840 vdd.n508 66.2847
R2595 vdd.n2840 vdd.n509 66.2847
R2596 vdd.n2840 vdd.n510 66.2847
R2597 vdd.n2840 vdd.n511 66.2847
R2598 vdd.n2840 vdd.n512 66.2847
R2599 vdd.n2840 vdd.n513 66.2847
R2600 vdd.n2840 vdd.n514 66.2847
R2601 vdd.n2905 vdd.n329 66.2847
R2602 vdd.n2914 vdd.n329 66.2847
R2603 vdd.n439 vdd.n329 66.2847
R2604 vdd.n2921 vdd.n329 66.2847
R2605 vdd.n432 vdd.n329 66.2847
R2606 vdd.n2928 vdd.n329 66.2847
R2607 vdd.n425 vdd.n329 66.2847
R2608 vdd.n2935 vdd.n329 66.2847
R2609 vdd.n418 vdd.n329 66.2847
R2610 vdd.n2942 vdd.n329 66.2847
R2611 vdd.n412 vdd.n329 66.2847
R2612 vdd.n407 vdd.n329 66.2847
R2613 vdd.n2953 vdd.n329 66.2847
R2614 vdd.n399 vdd.n329 66.2847
R2615 vdd.n2960 vdd.n329 66.2847
R2616 vdd.n392 vdd.n329 66.2847
R2617 vdd.n2967 vdd.n329 66.2847
R2618 vdd.n385 vdd.n329 66.2847
R2619 vdd.n2974 vdd.n329 66.2847
R2620 vdd.n378 vdd.n329 66.2847
R2621 vdd.n2981 vdd.n329 66.2847
R2622 vdd.n372 vdd.n329 66.2847
R2623 vdd.n367 vdd.n329 66.2847
R2624 vdd.n2992 vdd.n329 66.2847
R2625 vdd.n359 vdd.n329 66.2847
R2626 vdd.n2999 vdd.n329 66.2847
R2627 vdd.n352 vdd.n329 66.2847
R2628 vdd.n3006 vdd.n329 66.2847
R2629 vdd.n345 vdd.n329 66.2847
R2630 vdd.n3013 vdd.n329 66.2847
R2631 vdd.n3016 vdd.n329 66.2847
R2632 vdd.n333 vdd.n329 66.2847
R2633 vdd.n334 vdd.n333 52.4337
R2634 vdd.n3016 vdd.n3015 52.4337
R2635 vdd.n3013 vdd.n3012 52.4337
R2636 vdd.n3008 vdd.n345 52.4337
R2637 vdd.n3006 vdd.n3005 52.4337
R2638 vdd.n3001 vdd.n352 52.4337
R2639 vdd.n2999 vdd.n2998 52.4337
R2640 vdd.n2994 vdd.n359 52.4337
R2641 vdd.n2992 vdd.n2991 52.4337
R2642 vdd.n368 vdd.n367 52.4337
R2643 vdd.n2983 vdd.n372 52.4337
R2644 vdd.n2981 vdd.n2980 52.4337
R2645 vdd.n2976 vdd.n378 52.4337
R2646 vdd.n2974 vdd.n2973 52.4337
R2647 vdd.n2969 vdd.n385 52.4337
R2648 vdd.n2967 vdd.n2966 52.4337
R2649 vdd.n2962 vdd.n392 52.4337
R2650 vdd.n2960 vdd.n2959 52.4337
R2651 vdd.n2955 vdd.n399 52.4337
R2652 vdd.n2953 vdd.n2952 52.4337
R2653 vdd.n408 vdd.n407 52.4337
R2654 vdd.n2944 vdd.n412 52.4337
R2655 vdd.n2942 vdd.n2941 52.4337
R2656 vdd.n2937 vdd.n418 52.4337
R2657 vdd.n2935 vdd.n2934 52.4337
R2658 vdd.n2930 vdd.n425 52.4337
R2659 vdd.n2928 vdd.n2927 52.4337
R2660 vdd.n2923 vdd.n432 52.4337
R2661 vdd.n2921 vdd.n2920 52.4337
R2662 vdd.n2916 vdd.n439 52.4337
R2663 vdd.n2914 vdd.n2913 52.4337
R2664 vdd.n2906 vdd.n2905 52.4337
R2665 vdd.n2842 vdd.n2841 52.4337
R2666 vdd.n517 vdd.n485 52.4337
R2667 vdd.n523 vdd.n486 52.4337
R2668 vdd.n2831 vdd.n487 52.4337
R2669 vdd.n2827 vdd.n488 52.4337
R2670 vdd.n2823 vdd.n489 52.4337
R2671 vdd.n2819 vdd.n490 52.4337
R2672 vdd.n2815 vdd.n491 52.4337
R2673 vdd.n2811 vdd.n492 52.4337
R2674 vdd.n2807 vdd.n493 52.4337
R2675 vdd.n2799 vdd.n494 52.4337
R2676 vdd.n2795 vdd.n495 52.4337
R2677 vdd.n2791 vdd.n496 52.4337
R2678 vdd.n2787 vdd.n497 52.4337
R2679 vdd.n2783 vdd.n498 52.4337
R2680 vdd.n2779 vdd.n499 52.4337
R2681 vdd.n2775 vdd.n500 52.4337
R2682 vdd.n2771 vdd.n501 52.4337
R2683 vdd.n2767 vdd.n502 52.4337
R2684 vdd.n2763 vdd.n503 52.4337
R2685 vdd.n2759 vdd.n504 52.4337
R2686 vdd.n2753 vdd.n505 52.4337
R2687 vdd.n2749 vdd.n506 52.4337
R2688 vdd.n2745 vdd.n507 52.4337
R2689 vdd.n2741 vdd.n508 52.4337
R2690 vdd.n2737 vdd.n509 52.4337
R2691 vdd.n2733 vdd.n510 52.4337
R2692 vdd.n2729 vdd.n511 52.4337
R2693 vdd.n2725 vdd.n512 52.4337
R2694 vdd.n2721 vdd.n513 52.4337
R2695 vdd.n2717 vdd.n514 52.4337
R2696 vdd.n1936 vdd.n1516 52.4337
R2697 vdd.n1934 vdd.n1933 52.4337
R2698 vdd.n1523 vdd.n1522 52.4337
R2699 vdd.n1712 vdd.n1711 52.4337
R2700 vdd.n1709 vdd.n1708 52.4337
R2701 vdd.n1704 vdd.n1531 52.4337
R2702 vdd.n1702 vdd.n1701 52.4337
R2703 vdd.n1697 vdd.n1538 52.4337
R2704 vdd.n1695 vdd.n1694 52.4337
R2705 vdd.n1547 vdd.n1546 52.4337
R2706 vdd.n1686 vdd.n1551 52.4337
R2707 vdd.n1684 vdd.n1683 52.4337
R2708 vdd.n1679 vdd.n1557 52.4337
R2709 vdd.n1677 vdd.n1676 52.4337
R2710 vdd.n1672 vdd.n1564 52.4337
R2711 vdd.n1670 vdd.n1669 52.4337
R2712 vdd.n1665 vdd.n1571 52.4337
R2713 vdd.n1663 vdd.n1662 52.4337
R2714 vdd.n1658 vdd.n1578 52.4337
R2715 vdd.n1656 vdd.n1655 52.4337
R2716 vdd.n1587 vdd.n1586 52.4337
R2717 vdd.n1647 vdd.n1591 52.4337
R2718 vdd.n1645 vdd.n1644 52.4337
R2719 vdd.n1640 vdd.n1597 52.4337
R2720 vdd.n1638 vdd.n1637 52.4337
R2721 vdd.n1633 vdd.n1604 52.4337
R2722 vdd.n1631 vdd.n1630 52.4337
R2723 vdd.n1626 vdd.n1612 52.4337
R2724 vdd.n1624 vdd.n1623 52.4337
R2725 vdd.n1619 vdd.n1618 52.4337
R2726 vdd.n1614 vdd.n1613 52.4337
R2727 vdd.n1945 vdd.n860 52.4337
R2728 vdd.n1423 vdd.n1422 52.4337
R2729 vdd.n1229 vdd.n1197 52.4337
R2730 vdd.n1233 vdd.n1198 52.4337
R2731 vdd.n1235 vdd.n1199 52.4337
R2732 vdd.n1239 vdd.n1200 52.4337
R2733 vdd.n1241 vdd.n1201 52.4337
R2734 vdd.n1245 vdd.n1202 52.4337
R2735 vdd.n1247 vdd.n1203 52.4337
R2736 vdd.n1251 vdd.n1204 52.4337
R2737 vdd.n1253 vdd.n1205 52.4337
R2738 vdd.n1259 vdd.n1206 52.4337
R2739 vdd.n1261 vdd.n1207 52.4337
R2740 vdd.n1265 vdd.n1208 52.4337
R2741 vdd.n1267 vdd.n1209 52.4337
R2742 vdd.n1271 vdd.n1210 52.4337
R2743 vdd.n1273 vdd.n1211 52.4337
R2744 vdd.n1277 vdd.n1212 52.4337
R2745 vdd.n1279 vdd.n1213 52.4337
R2746 vdd.n1283 vdd.n1214 52.4337
R2747 vdd.n1285 vdd.n1215 52.4337
R2748 vdd.n1357 vdd.n1216 52.4337
R2749 vdd.n1290 vdd.n1217 52.4337
R2750 vdd.n1294 vdd.n1218 52.4337
R2751 vdd.n1296 vdd.n1219 52.4337
R2752 vdd.n1300 vdd.n1220 52.4337
R2753 vdd.n1302 vdd.n1221 52.4337
R2754 vdd.n1306 vdd.n1222 52.4337
R2755 vdd.n1308 vdd.n1223 52.4337
R2756 vdd.n1312 vdd.n1224 52.4337
R2757 vdd.n1314 vdd.n1225 52.4337
R2758 vdd.n1318 vdd.n1226 52.4337
R2759 vdd.n1422 vdd.n1196 52.4337
R2760 vdd.n1232 vdd.n1197 52.4337
R2761 vdd.n1234 vdd.n1198 52.4337
R2762 vdd.n1238 vdd.n1199 52.4337
R2763 vdd.n1240 vdd.n1200 52.4337
R2764 vdd.n1244 vdd.n1201 52.4337
R2765 vdd.n1246 vdd.n1202 52.4337
R2766 vdd.n1250 vdd.n1203 52.4337
R2767 vdd.n1252 vdd.n1204 52.4337
R2768 vdd.n1258 vdd.n1205 52.4337
R2769 vdd.n1260 vdd.n1206 52.4337
R2770 vdd.n1264 vdd.n1207 52.4337
R2771 vdd.n1266 vdd.n1208 52.4337
R2772 vdd.n1270 vdd.n1209 52.4337
R2773 vdd.n1272 vdd.n1210 52.4337
R2774 vdd.n1276 vdd.n1211 52.4337
R2775 vdd.n1278 vdd.n1212 52.4337
R2776 vdd.n1282 vdd.n1213 52.4337
R2777 vdd.n1284 vdd.n1214 52.4337
R2778 vdd.n1288 vdd.n1215 52.4337
R2779 vdd.n1289 vdd.n1216 52.4337
R2780 vdd.n1293 vdd.n1217 52.4337
R2781 vdd.n1295 vdd.n1218 52.4337
R2782 vdd.n1299 vdd.n1219 52.4337
R2783 vdd.n1301 vdd.n1220 52.4337
R2784 vdd.n1305 vdd.n1221 52.4337
R2785 vdd.n1307 vdd.n1222 52.4337
R2786 vdd.n1311 vdd.n1223 52.4337
R2787 vdd.n1313 vdd.n1224 52.4337
R2788 vdd.n1317 vdd.n1225 52.4337
R2789 vdd.n1319 vdd.n1226 52.4337
R2790 vdd.n860 vdd.n859 52.4337
R2791 vdd.n1615 vdd.n1614 52.4337
R2792 vdd.n1620 vdd.n1619 52.4337
R2793 vdd.n1625 vdd.n1624 52.4337
R2794 vdd.n1612 vdd.n1605 52.4337
R2795 vdd.n1632 vdd.n1631 52.4337
R2796 vdd.n1604 vdd.n1598 52.4337
R2797 vdd.n1639 vdd.n1638 52.4337
R2798 vdd.n1597 vdd.n1592 52.4337
R2799 vdd.n1646 vdd.n1645 52.4337
R2800 vdd.n1591 vdd.n1590 52.4337
R2801 vdd.n1586 vdd.n1579 52.4337
R2802 vdd.n1657 vdd.n1656 52.4337
R2803 vdd.n1578 vdd.n1572 52.4337
R2804 vdd.n1664 vdd.n1663 52.4337
R2805 vdd.n1571 vdd.n1565 52.4337
R2806 vdd.n1671 vdd.n1670 52.4337
R2807 vdd.n1564 vdd.n1558 52.4337
R2808 vdd.n1678 vdd.n1677 52.4337
R2809 vdd.n1557 vdd.n1552 52.4337
R2810 vdd.n1685 vdd.n1684 52.4337
R2811 vdd.n1551 vdd.n1550 52.4337
R2812 vdd.n1546 vdd.n1539 52.4337
R2813 vdd.n1696 vdd.n1695 52.4337
R2814 vdd.n1538 vdd.n1532 52.4337
R2815 vdd.n1703 vdd.n1702 52.4337
R2816 vdd.n1531 vdd.n1525 52.4337
R2817 vdd.n1710 vdd.n1709 52.4337
R2818 vdd.n1713 vdd.n1712 52.4337
R2819 vdd.n1522 vdd.n1517 52.4337
R2820 vdd.n1935 vdd.n1934 52.4337
R2821 vdd.n1516 vdd.n865 52.4337
R2822 vdd.n2841 vdd.n483 52.4337
R2823 vdd.n522 vdd.n485 52.4337
R2824 vdd.n2832 vdd.n486 52.4337
R2825 vdd.n2828 vdd.n487 52.4337
R2826 vdd.n2824 vdd.n488 52.4337
R2827 vdd.n2820 vdd.n489 52.4337
R2828 vdd.n2816 vdd.n490 52.4337
R2829 vdd.n2812 vdd.n491 52.4337
R2830 vdd.n2808 vdd.n492 52.4337
R2831 vdd.n2798 vdd.n493 52.4337
R2832 vdd.n2796 vdd.n494 52.4337
R2833 vdd.n2792 vdd.n495 52.4337
R2834 vdd.n2788 vdd.n496 52.4337
R2835 vdd.n2784 vdd.n497 52.4337
R2836 vdd.n2780 vdd.n498 52.4337
R2837 vdd.n2776 vdd.n499 52.4337
R2838 vdd.n2772 vdd.n500 52.4337
R2839 vdd.n2768 vdd.n501 52.4337
R2840 vdd.n2764 vdd.n502 52.4337
R2841 vdd.n2760 vdd.n503 52.4337
R2842 vdd.n2752 vdd.n504 52.4337
R2843 vdd.n2750 vdd.n505 52.4337
R2844 vdd.n2746 vdd.n506 52.4337
R2845 vdd.n2742 vdd.n507 52.4337
R2846 vdd.n2738 vdd.n508 52.4337
R2847 vdd.n2734 vdd.n509 52.4337
R2848 vdd.n2730 vdd.n510 52.4337
R2849 vdd.n2726 vdd.n511 52.4337
R2850 vdd.n2722 vdd.n512 52.4337
R2851 vdd.n2718 vdd.n513 52.4337
R2852 vdd.n2714 vdd.n514 52.4337
R2853 vdd.n2905 vdd.n440 52.4337
R2854 vdd.n2915 vdd.n2914 52.4337
R2855 vdd.n439 vdd.n433 52.4337
R2856 vdd.n2922 vdd.n2921 52.4337
R2857 vdd.n432 vdd.n426 52.4337
R2858 vdd.n2929 vdd.n2928 52.4337
R2859 vdd.n425 vdd.n419 52.4337
R2860 vdd.n2936 vdd.n2935 52.4337
R2861 vdd.n418 vdd.n413 52.4337
R2862 vdd.n2943 vdd.n2942 52.4337
R2863 vdd.n412 vdd.n411 52.4337
R2864 vdd.n407 vdd.n400 52.4337
R2865 vdd.n2954 vdd.n2953 52.4337
R2866 vdd.n399 vdd.n393 52.4337
R2867 vdd.n2961 vdd.n2960 52.4337
R2868 vdd.n392 vdd.n386 52.4337
R2869 vdd.n2968 vdd.n2967 52.4337
R2870 vdd.n385 vdd.n379 52.4337
R2871 vdd.n2975 vdd.n2974 52.4337
R2872 vdd.n378 vdd.n373 52.4337
R2873 vdd.n2982 vdd.n2981 52.4337
R2874 vdd.n372 vdd.n371 52.4337
R2875 vdd.n367 vdd.n360 52.4337
R2876 vdd.n2993 vdd.n2992 52.4337
R2877 vdd.n359 vdd.n353 52.4337
R2878 vdd.n3000 vdd.n2999 52.4337
R2879 vdd.n352 vdd.n346 52.4337
R2880 vdd.n3007 vdd.n3006 52.4337
R2881 vdd.n345 vdd.n338 52.4337
R2882 vdd.n3014 vdd.n3013 52.4337
R2883 vdd.n3017 vdd.n3016 52.4337
R2884 vdd.n333 vdd.n330 52.4337
R2885 vdd.t155 vdd.t165 51.4683
R2886 vdd.n250 vdd.n248 42.0461
R2887 vdd.n160 vdd.n158 42.0461
R2888 vdd.n71 vdd.n69 42.0461
R2889 vdd.n1112 vdd.n1110 42.0461
R2890 vdd.n1022 vdd.n1020 42.0461
R2891 vdd.n933 vdd.n931 42.0461
R2892 vdd.n296 vdd.n295 41.6884
R2893 vdd.n206 vdd.n205 41.6884
R2894 vdd.n117 vdd.n116 41.6884
R2895 vdd.n1158 vdd.n1157 41.6884
R2896 vdd.n1068 vdd.n1067 41.6884
R2897 vdd.n979 vdd.n978 41.6884
R2898 vdd.n1322 vdd.n1321 41.1157
R2899 vdd.n1360 vdd.n1359 41.1157
R2900 vdd.n1256 vdd.n1255 41.1157
R2901 vdd.n2910 vdd.n2909 41.1157
R2902 vdd.n2949 vdd.n406 41.1157
R2903 vdd.n2988 vdd.n366 41.1157
R2904 vdd.n2667 vdd.n2666 39.2114
R2905 vdd.n2664 vdd.n2663 39.2114
R2906 vdd.n2659 vdd.n605 39.2114
R2907 vdd.n2657 vdd.n2656 39.2114
R2908 vdd.n2652 vdd.n608 39.2114
R2909 vdd.n2650 vdd.n2649 39.2114
R2910 vdd.n2645 vdd.n611 39.2114
R2911 vdd.n2643 vdd.n2642 39.2114
R2912 vdd.n2639 vdd.n2638 39.2114
R2913 vdd.n2634 vdd.n614 39.2114
R2914 vdd.n2632 vdd.n2631 39.2114
R2915 vdd.n2627 vdd.n617 39.2114
R2916 vdd.n2625 vdd.n2624 39.2114
R2917 vdd.n2620 vdd.n620 39.2114
R2918 vdd.n2618 vdd.n2617 39.2114
R2919 vdd.n2612 vdd.n625 39.2114
R2920 vdd.n2610 vdd.n2609 39.2114
R2921 vdd.n2470 vdd.n703 39.2114
R2922 vdd.n2465 vdd.n2219 39.2114
R2923 vdd.n2462 vdd.n2220 39.2114
R2924 vdd.n2458 vdd.n2221 39.2114
R2925 vdd.n2454 vdd.n2222 39.2114
R2926 vdd.n2450 vdd.n2223 39.2114
R2927 vdd.n2446 vdd.n2224 39.2114
R2928 vdd.n2442 vdd.n2225 39.2114
R2929 vdd.n2438 vdd.n2226 39.2114
R2930 vdd.n2434 vdd.n2227 39.2114
R2931 vdd.n2430 vdd.n2228 39.2114
R2932 vdd.n2426 vdd.n2229 39.2114
R2933 vdd.n2422 vdd.n2230 39.2114
R2934 vdd.n2418 vdd.n2231 39.2114
R2935 vdd.n2414 vdd.n2232 39.2114
R2936 vdd.n2410 vdd.n2233 39.2114
R2937 vdd.n2405 vdd.n2234 39.2114
R2938 vdd.n2213 vdd.n743 39.2114
R2939 vdd.n2209 vdd.n742 39.2114
R2940 vdd.n2205 vdd.n741 39.2114
R2941 vdd.n2201 vdd.n740 39.2114
R2942 vdd.n2197 vdd.n739 39.2114
R2943 vdd.n2193 vdd.n738 39.2114
R2944 vdd.n2189 vdd.n737 39.2114
R2945 vdd.n2185 vdd.n736 39.2114
R2946 vdd.n2181 vdd.n735 39.2114
R2947 vdd.n2177 vdd.n734 39.2114
R2948 vdd.n2173 vdd.n733 39.2114
R2949 vdd.n2169 vdd.n732 39.2114
R2950 vdd.n2165 vdd.n731 39.2114
R2951 vdd.n2161 vdd.n730 39.2114
R2952 vdd.n2157 vdd.n729 39.2114
R2953 vdd.n2152 vdd.n728 39.2114
R2954 vdd.n2148 vdd.n727 39.2114
R2955 vdd.n1724 vdd.n838 39.2114
R2956 vdd.n1730 vdd.n1729 39.2114
R2957 vdd.n1733 vdd.n1732 39.2114
R2958 vdd.n1738 vdd.n1737 39.2114
R2959 vdd.n1741 vdd.n1740 39.2114
R2960 vdd.n1746 vdd.n1745 39.2114
R2961 vdd.n1749 vdd.n1748 39.2114
R2962 vdd.n1754 vdd.n1753 39.2114
R2963 vdd.n1925 vdd.n1756 39.2114
R2964 vdd.n1924 vdd.n1923 39.2114
R2965 vdd.n1917 vdd.n1758 39.2114
R2966 vdd.n1916 vdd.n1915 39.2114
R2967 vdd.n1909 vdd.n1760 39.2114
R2968 vdd.n1908 vdd.n1907 39.2114
R2969 vdd.n1901 vdd.n1762 39.2114
R2970 vdd.n1900 vdd.n1899 39.2114
R2971 vdd.n1893 vdd.n1764 39.2114
R2972 vdd.n2586 vdd.n2585 39.2114
R2973 vdd.n2581 vdd.n2553 39.2114
R2974 vdd.n2579 vdd.n2578 39.2114
R2975 vdd.n2574 vdd.n2556 39.2114
R2976 vdd.n2572 vdd.n2571 39.2114
R2977 vdd.n2567 vdd.n2559 39.2114
R2978 vdd.n2565 vdd.n2564 39.2114
R2979 vdd.n2560 vdd.n577 39.2114
R2980 vdd.n2704 vdd.n2703 39.2114
R2981 vdd.n2701 vdd.n2700 39.2114
R2982 vdd.n2696 vdd.n581 39.2114
R2983 vdd.n2694 vdd.n2693 39.2114
R2984 vdd.n2689 vdd.n584 39.2114
R2985 vdd.n2687 vdd.n2686 39.2114
R2986 vdd.n2682 vdd.n587 39.2114
R2987 vdd.n2680 vdd.n2679 39.2114
R2988 vdd.n2675 vdd.n593 39.2114
R2989 vdd.n2472 vdd.n706 39.2114
R2990 vdd.n2235 vdd.n708 39.2114
R2991 vdd.n2261 vdd.n2236 39.2114
R2992 vdd.n2265 vdd.n2237 39.2114
R2993 vdd.n2269 vdd.n2238 39.2114
R2994 vdd.n2273 vdd.n2239 39.2114
R2995 vdd.n2277 vdd.n2240 39.2114
R2996 vdd.n2281 vdd.n2241 39.2114
R2997 vdd.n2285 vdd.n2242 39.2114
R2998 vdd.n2289 vdd.n2243 39.2114
R2999 vdd.n2293 vdd.n2244 39.2114
R3000 vdd.n2297 vdd.n2245 39.2114
R3001 vdd.n2301 vdd.n2246 39.2114
R3002 vdd.n2305 vdd.n2247 39.2114
R3003 vdd.n2309 vdd.n2248 39.2114
R3004 vdd.n2313 vdd.n2249 39.2114
R3005 vdd.n2317 vdd.n2250 39.2114
R3006 vdd.n2473 vdd.n2472 39.2114
R3007 vdd.n2260 vdd.n2235 39.2114
R3008 vdd.n2264 vdd.n2236 39.2114
R3009 vdd.n2268 vdd.n2237 39.2114
R3010 vdd.n2272 vdd.n2238 39.2114
R3011 vdd.n2276 vdd.n2239 39.2114
R3012 vdd.n2280 vdd.n2240 39.2114
R3013 vdd.n2284 vdd.n2241 39.2114
R3014 vdd.n2288 vdd.n2242 39.2114
R3015 vdd.n2292 vdd.n2243 39.2114
R3016 vdd.n2296 vdd.n2244 39.2114
R3017 vdd.n2300 vdd.n2245 39.2114
R3018 vdd.n2304 vdd.n2246 39.2114
R3019 vdd.n2308 vdd.n2247 39.2114
R3020 vdd.n2312 vdd.n2248 39.2114
R3021 vdd.n2316 vdd.n2249 39.2114
R3022 vdd.n2319 vdd.n2250 39.2114
R3023 vdd.n593 vdd.n588 39.2114
R3024 vdd.n2681 vdd.n2680 39.2114
R3025 vdd.n587 vdd.n585 39.2114
R3026 vdd.n2688 vdd.n2687 39.2114
R3027 vdd.n584 vdd.n582 39.2114
R3028 vdd.n2695 vdd.n2694 39.2114
R3029 vdd.n581 vdd.n579 39.2114
R3030 vdd.n2702 vdd.n2701 39.2114
R3031 vdd.n2705 vdd.n2704 39.2114
R3032 vdd.n2561 vdd.n2560 39.2114
R3033 vdd.n2566 vdd.n2565 39.2114
R3034 vdd.n2559 vdd.n2557 39.2114
R3035 vdd.n2573 vdd.n2572 39.2114
R3036 vdd.n2556 vdd.n2554 39.2114
R3037 vdd.n2580 vdd.n2579 39.2114
R3038 vdd.n2553 vdd.n2551 39.2114
R3039 vdd.n2587 vdd.n2586 39.2114
R3040 vdd.n1725 vdd.n1724 39.2114
R3041 vdd.n1731 vdd.n1730 39.2114
R3042 vdd.n1732 vdd.n1721 39.2114
R3043 vdd.n1739 vdd.n1738 39.2114
R3044 vdd.n1740 vdd.n1719 39.2114
R3045 vdd.n1747 vdd.n1746 39.2114
R3046 vdd.n1748 vdd.n1717 39.2114
R3047 vdd.n1755 vdd.n1754 39.2114
R3048 vdd.n1926 vdd.n1925 39.2114
R3049 vdd.n1923 vdd.n1922 39.2114
R3050 vdd.n1918 vdd.n1917 39.2114
R3051 vdd.n1915 vdd.n1914 39.2114
R3052 vdd.n1910 vdd.n1909 39.2114
R3053 vdd.n1907 vdd.n1906 39.2114
R3054 vdd.n1902 vdd.n1901 39.2114
R3055 vdd.n1899 vdd.n1898 39.2114
R3056 vdd.n1894 vdd.n1893 39.2114
R3057 vdd.n2151 vdd.n727 39.2114
R3058 vdd.n2156 vdd.n728 39.2114
R3059 vdd.n2160 vdd.n729 39.2114
R3060 vdd.n2164 vdd.n730 39.2114
R3061 vdd.n2168 vdd.n731 39.2114
R3062 vdd.n2172 vdd.n732 39.2114
R3063 vdd.n2176 vdd.n733 39.2114
R3064 vdd.n2180 vdd.n734 39.2114
R3065 vdd.n2184 vdd.n735 39.2114
R3066 vdd.n2188 vdd.n736 39.2114
R3067 vdd.n2192 vdd.n737 39.2114
R3068 vdd.n2196 vdd.n738 39.2114
R3069 vdd.n2200 vdd.n739 39.2114
R3070 vdd.n2204 vdd.n740 39.2114
R3071 vdd.n2208 vdd.n741 39.2114
R3072 vdd.n2212 vdd.n742 39.2114
R3073 vdd.n745 vdd.n743 39.2114
R3074 vdd.n2470 vdd.n2469 39.2114
R3075 vdd.n2463 vdd.n2219 39.2114
R3076 vdd.n2459 vdd.n2220 39.2114
R3077 vdd.n2455 vdd.n2221 39.2114
R3078 vdd.n2451 vdd.n2222 39.2114
R3079 vdd.n2447 vdd.n2223 39.2114
R3080 vdd.n2443 vdd.n2224 39.2114
R3081 vdd.n2439 vdd.n2225 39.2114
R3082 vdd.n2435 vdd.n2226 39.2114
R3083 vdd.n2431 vdd.n2227 39.2114
R3084 vdd.n2427 vdd.n2228 39.2114
R3085 vdd.n2423 vdd.n2229 39.2114
R3086 vdd.n2419 vdd.n2230 39.2114
R3087 vdd.n2415 vdd.n2231 39.2114
R3088 vdd.n2411 vdd.n2232 39.2114
R3089 vdd.n2406 vdd.n2233 39.2114
R3090 vdd.n2402 vdd.n2234 39.2114
R3091 vdd.n2611 vdd.n2610 39.2114
R3092 vdd.n625 vdd.n621 39.2114
R3093 vdd.n2619 vdd.n2618 39.2114
R3094 vdd.n620 vdd.n618 39.2114
R3095 vdd.n2626 vdd.n2625 39.2114
R3096 vdd.n617 vdd.n615 39.2114
R3097 vdd.n2633 vdd.n2632 39.2114
R3098 vdd.n614 vdd.n612 39.2114
R3099 vdd.n2640 vdd.n2639 39.2114
R3100 vdd.n2644 vdd.n2643 39.2114
R3101 vdd.n611 vdd.n609 39.2114
R3102 vdd.n2651 vdd.n2650 39.2114
R3103 vdd.n608 vdd.n606 39.2114
R3104 vdd.n2658 vdd.n2657 39.2114
R3105 vdd.n605 vdd.n603 39.2114
R3106 vdd.n2665 vdd.n2664 39.2114
R3107 vdd.n2668 vdd.n2667 39.2114
R3108 vdd.n753 vdd.n709 39.2114
R3109 vdd.n2140 vdd.n710 39.2114
R3110 vdd.n2136 vdd.n711 39.2114
R3111 vdd.n2132 vdd.n712 39.2114
R3112 vdd.n2128 vdd.n713 39.2114
R3113 vdd.n2124 vdd.n714 39.2114
R3114 vdd.n2120 vdd.n715 39.2114
R3115 vdd.n2116 vdd.n716 39.2114
R3116 vdd.n2112 vdd.n717 39.2114
R3117 vdd.n2108 vdd.n718 39.2114
R3118 vdd.n2104 vdd.n719 39.2114
R3119 vdd.n2100 vdd.n720 39.2114
R3120 vdd.n2096 vdd.n721 39.2114
R3121 vdd.n2092 vdd.n722 39.2114
R3122 vdd.n2088 vdd.n723 39.2114
R3123 vdd.n2084 vdd.n724 39.2114
R3124 vdd.n2080 vdd.n725 39.2114
R3125 vdd.n1983 vdd.n842 39.2114
R3126 vdd.n1982 vdd.n1981 39.2114
R3127 vdd.n1975 vdd.n844 39.2114
R3128 vdd.n1974 vdd.n1973 39.2114
R3129 vdd.n1967 vdd.n846 39.2114
R3130 vdd.n1966 vdd.n1965 39.2114
R3131 vdd.n1959 vdd.n848 39.2114
R3132 vdd.n1958 vdd.n1957 39.2114
R3133 vdd.n851 vdd.n850 39.2114
R3134 vdd.n1799 vdd.n1798 39.2114
R3135 vdd.n1804 vdd.n1803 39.2114
R3136 vdd.n1807 vdd.n1806 39.2114
R3137 vdd.n1812 vdd.n1811 39.2114
R3138 vdd.n1815 vdd.n1814 39.2114
R3139 vdd.n1820 vdd.n1819 39.2114
R3140 vdd.n1823 vdd.n1822 39.2114
R3141 vdd.n1829 vdd.n1828 39.2114
R3142 vdd.n2077 vdd.n725 39.2114
R3143 vdd.n2081 vdd.n724 39.2114
R3144 vdd.n2085 vdd.n723 39.2114
R3145 vdd.n2089 vdd.n722 39.2114
R3146 vdd.n2093 vdd.n721 39.2114
R3147 vdd.n2097 vdd.n720 39.2114
R3148 vdd.n2101 vdd.n719 39.2114
R3149 vdd.n2105 vdd.n718 39.2114
R3150 vdd.n2109 vdd.n717 39.2114
R3151 vdd.n2113 vdd.n716 39.2114
R3152 vdd.n2117 vdd.n715 39.2114
R3153 vdd.n2121 vdd.n714 39.2114
R3154 vdd.n2125 vdd.n713 39.2114
R3155 vdd.n2129 vdd.n712 39.2114
R3156 vdd.n2133 vdd.n711 39.2114
R3157 vdd.n2137 vdd.n710 39.2114
R3158 vdd.n2141 vdd.n709 39.2114
R3159 vdd.n1984 vdd.n1983 39.2114
R3160 vdd.n1981 vdd.n1980 39.2114
R3161 vdd.n1976 vdd.n1975 39.2114
R3162 vdd.n1973 vdd.n1972 39.2114
R3163 vdd.n1968 vdd.n1967 39.2114
R3164 vdd.n1965 vdd.n1964 39.2114
R3165 vdd.n1960 vdd.n1959 39.2114
R3166 vdd.n1957 vdd.n1956 39.2114
R3167 vdd.n852 vdd.n851 39.2114
R3168 vdd.n1800 vdd.n1799 39.2114
R3169 vdd.n1805 vdd.n1804 39.2114
R3170 vdd.n1806 vdd.n1796 39.2114
R3171 vdd.n1813 vdd.n1812 39.2114
R3172 vdd.n1814 vdd.n1794 39.2114
R3173 vdd.n1821 vdd.n1820 39.2114
R3174 vdd.n1822 vdd.n1790 39.2114
R3175 vdd.n1830 vdd.n1829 39.2114
R3176 vdd.n1949 vdd.n1948 37.2369
R3177 vdd.n1652 vdd.n1585 37.2369
R3178 vdd.n1691 vdd.n1545 37.2369
R3179 vdd.n2758 vdd.n558 37.2369
R3180 vdd.n2806 vdd.n2805 37.2369
R3181 vdd.n2713 vdd.n2712 37.2369
R3182 vdd.n1991 vdd.n837 31.6883
R3183 vdd.n2216 vdd.n746 31.6883
R3184 vdd.n2149 vdd.n749 31.6883
R3185 vdd.n1895 vdd.n1892 31.6883
R3186 vdd.n2403 vdd.n2401 31.6883
R3187 vdd.n2608 vdd.n2607 31.6883
R3188 vdd.n2480 vdd.n702 31.6883
R3189 vdd.n2671 vdd.n2670 31.6883
R3190 vdd.n2590 vdd.n2589 31.6883
R3191 vdd.n2676 vdd.n592 31.6883
R3192 vdd.n2322 vdd.n2321 31.6883
R3193 vdd.n2476 vdd.n2475 31.6883
R3194 vdd.n1987 vdd.n1986 31.6883
R3195 vdd.n2144 vdd.n2143 31.6883
R3196 vdd.n2076 vdd.n2075 31.6883
R3197 vdd.n1833 vdd.n1832 31.6883
R3198 vdd.n1826 vdd.n1792 30.449
R3199 vdd.n757 vdd.n756 30.449
R3200 vdd.n1767 vdd.n1766 30.449
R3201 vdd.n2154 vdd.n748 30.449
R3202 vdd.n2258 vdd.n2257 30.449
R3203 vdd.n2614 vdd.n623 30.449
R3204 vdd.n2408 vdd.n2254 30.449
R3205 vdd.n591 vdd.n590 30.449
R3206 vdd.n1421 vdd.n1228 22.6735
R3207 vdd.n1943 vdd.n863 22.6735
R3208 vdd.n2840 vdd.n516 22.6735
R3209 vdd.n3025 vdd.n329 22.6735
R3210 vdd.n1432 vdd.n1190 19.3944
R3211 vdd.n1432 vdd.n1188 19.3944
R3212 vdd.n1436 vdd.n1188 19.3944
R3213 vdd.n1436 vdd.n1178 19.3944
R3214 vdd.n1449 vdd.n1178 19.3944
R3215 vdd.n1449 vdd.n1176 19.3944
R3216 vdd.n1453 vdd.n1176 19.3944
R3217 vdd.n1453 vdd.n1168 19.3944
R3218 vdd.n1467 vdd.n1168 19.3944
R3219 vdd.n1467 vdd.n1166 19.3944
R3220 vdd.n1471 vdd.n1166 19.3944
R3221 vdd.n1471 vdd.n885 19.3944
R3222 vdd.n1483 vdd.n885 19.3944
R3223 vdd.n1483 vdd.n883 19.3944
R3224 vdd.n1487 vdd.n883 19.3944
R3225 vdd.n1487 vdd.n875 19.3944
R3226 vdd.n1500 vdd.n875 19.3944
R3227 vdd.n1500 vdd.n872 19.3944
R3228 vdd.n1506 vdd.n872 19.3944
R3229 vdd.n1506 vdd.n873 19.3944
R3230 vdd.n873 vdd.n862 19.3944
R3231 vdd.n1356 vdd.n1291 19.3944
R3232 vdd.n1352 vdd.n1291 19.3944
R3233 vdd.n1352 vdd.n1351 19.3944
R3234 vdd.n1351 vdd.n1350 19.3944
R3235 vdd.n1350 vdd.n1297 19.3944
R3236 vdd.n1346 vdd.n1297 19.3944
R3237 vdd.n1346 vdd.n1345 19.3944
R3238 vdd.n1345 vdd.n1344 19.3944
R3239 vdd.n1344 vdd.n1303 19.3944
R3240 vdd.n1340 vdd.n1303 19.3944
R3241 vdd.n1340 vdd.n1339 19.3944
R3242 vdd.n1339 vdd.n1338 19.3944
R3243 vdd.n1338 vdd.n1309 19.3944
R3244 vdd.n1334 vdd.n1309 19.3944
R3245 vdd.n1334 vdd.n1333 19.3944
R3246 vdd.n1333 vdd.n1332 19.3944
R3247 vdd.n1332 vdd.n1315 19.3944
R3248 vdd.n1328 vdd.n1315 19.3944
R3249 vdd.n1328 vdd.n1327 19.3944
R3250 vdd.n1327 vdd.n1326 19.3944
R3251 vdd.n1391 vdd.n1390 19.3944
R3252 vdd.n1390 vdd.n1389 19.3944
R3253 vdd.n1389 vdd.n1262 19.3944
R3254 vdd.n1385 vdd.n1262 19.3944
R3255 vdd.n1385 vdd.n1384 19.3944
R3256 vdd.n1384 vdd.n1383 19.3944
R3257 vdd.n1383 vdd.n1268 19.3944
R3258 vdd.n1379 vdd.n1268 19.3944
R3259 vdd.n1379 vdd.n1378 19.3944
R3260 vdd.n1378 vdd.n1377 19.3944
R3261 vdd.n1377 vdd.n1274 19.3944
R3262 vdd.n1373 vdd.n1274 19.3944
R3263 vdd.n1373 vdd.n1372 19.3944
R3264 vdd.n1372 vdd.n1371 19.3944
R3265 vdd.n1371 vdd.n1280 19.3944
R3266 vdd.n1367 vdd.n1280 19.3944
R3267 vdd.n1367 vdd.n1366 19.3944
R3268 vdd.n1366 vdd.n1365 19.3944
R3269 vdd.n1365 vdd.n1286 19.3944
R3270 vdd.n1361 vdd.n1286 19.3944
R3271 vdd.n1424 vdd.n1195 19.3944
R3272 vdd.n1419 vdd.n1195 19.3944
R3273 vdd.n1419 vdd.n1230 19.3944
R3274 vdd.n1415 vdd.n1230 19.3944
R3275 vdd.n1415 vdd.n1414 19.3944
R3276 vdd.n1414 vdd.n1413 19.3944
R3277 vdd.n1413 vdd.n1236 19.3944
R3278 vdd.n1409 vdd.n1236 19.3944
R3279 vdd.n1409 vdd.n1408 19.3944
R3280 vdd.n1408 vdd.n1407 19.3944
R3281 vdd.n1407 vdd.n1242 19.3944
R3282 vdd.n1403 vdd.n1242 19.3944
R3283 vdd.n1403 vdd.n1402 19.3944
R3284 vdd.n1402 vdd.n1401 19.3944
R3285 vdd.n1401 vdd.n1248 19.3944
R3286 vdd.n1397 vdd.n1248 19.3944
R3287 vdd.n1397 vdd.n1396 19.3944
R3288 vdd.n1396 vdd.n1395 19.3944
R3289 vdd.n1648 vdd.n1583 19.3944
R3290 vdd.n1648 vdd.n1589 19.3944
R3291 vdd.n1643 vdd.n1589 19.3944
R3292 vdd.n1643 vdd.n1642 19.3944
R3293 vdd.n1642 vdd.n1641 19.3944
R3294 vdd.n1641 vdd.n1596 19.3944
R3295 vdd.n1636 vdd.n1596 19.3944
R3296 vdd.n1636 vdd.n1635 19.3944
R3297 vdd.n1635 vdd.n1634 19.3944
R3298 vdd.n1634 vdd.n1603 19.3944
R3299 vdd.n1629 vdd.n1603 19.3944
R3300 vdd.n1629 vdd.n1628 19.3944
R3301 vdd.n1628 vdd.n1627 19.3944
R3302 vdd.n1627 vdd.n1611 19.3944
R3303 vdd.n1622 vdd.n1611 19.3944
R3304 vdd.n1622 vdd.n1621 19.3944
R3305 vdd.n1617 vdd.n1616 19.3944
R3306 vdd.n1950 vdd.n858 19.3944
R3307 vdd.n1687 vdd.n1543 19.3944
R3308 vdd.n1687 vdd.n1549 19.3944
R3309 vdd.n1682 vdd.n1549 19.3944
R3310 vdd.n1682 vdd.n1681 19.3944
R3311 vdd.n1681 vdd.n1680 19.3944
R3312 vdd.n1680 vdd.n1556 19.3944
R3313 vdd.n1675 vdd.n1556 19.3944
R3314 vdd.n1675 vdd.n1674 19.3944
R3315 vdd.n1674 vdd.n1673 19.3944
R3316 vdd.n1673 vdd.n1563 19.3944
R3317 vdd.n1668 vdd.n1563 19.3944
R3318 vdd.n1668 vdd.n1667 19.3944
R3319 vdd.n1667 vdd.n1666 19.3944
R3320 vdd.n1666 vdd.n1570 19.3944
R3321 vdd.n1661 vdd.n1570 19.3944
R3322 vdd.n1661 vdd.n1660 19.3944
R3323 vdd.n1660 vdd.n1659 19.3944
R3324 vdd.n1659 vdd.n1577 19.3944
R3325 vdd.n1654 vdd.n1577 19.3944
R3326 vdd.n1654 vdd.n1653 19.3944
R3327 vdd.n1938 vdd.n1937 19.3944
R3328 vdd.n1937 vdd.n1515 19.3944
R3329 vdd.n1932 vdd.n1931 19.3944
R3330 vdd.n1714 vdd.n1519 19.3944
R3331 vdd.n1714 vdd.n1521 19.3944
R3332 vdd.n1524 vdd.n1521 19.3944
R3333 vdd.n1707 vdd.n1524 19.3944
R3334 vdd.n1707 vdd.n1706 19.3944
R3335 vdd.n1706 vdd.n1705 19.3944
R3336 vdd.n1705 vdd.n1530 19.3944
R3337 vdd.n1700 vdd.n1530 19.3944
R3338 vdd.n1700 vdd.n1699 19.3944
R3339 vdd.n1699 vdd.n1698 19.3944
R3340 vdd.n1698 vdd.n1537 19.3944
R3341 vdd.n1693 vdd.n1537 19.3944
R3342 vdd.n1693 vdd.n1692 19.3944
R3343 vdd.n1428 vdd.n1193 19.3944
R3344 vdd.n1428 vdd.n1184 19.3944
R3345 vdd.n1441 vdd.n1184 19.3944
R3346 vdd.n1441 vdd.n1182 19.3944
R3347 vdd.n1445 vdd.n1182 19.3944
R3348 vdd.n1445 vdd.n1173 19.3944
R3349 vdd.n1458 vdd.n1173 19.3944
R3350 vdd.n1458 vdd.n1171 19.3944
R3351 vdd.n1463 vdd.n1171 19.3944
R3352 vdd.n1463 vdd.n1162 19.3944
R3353 vdd.n1475 vdd.n1162 19.3944
R3354 vdd.n1475 vdd.n890 19.3944
R3355 vdd.n1479 vdd.n890 19.3944
R3356 vdd.n1479 vdd.n880 19.3944
R3357 vdd.n1492 vdd.n880 19.3944
R3358 vdd.n1492 vdd.n878 19.3944
R3359 vdd.n1496 vdd.n878 19.3944
R3360 vdd.n1496 vdd.n868 19.3944
R3361 vdd.n1511 vdd.n868 19.3944
R3362 vdd.n1511 vdd.n866 19.3944
R3363 vdd.n1941 vdd.n866 19.3944
R3364 vdd.n2851 vdd.n477 19.3944
R3365 vdd.n2851 vdd.n475 19.3944
R3366 vdd.n2855 vdd.n475 19.3944
R3367 vdd.n2855 vdd.n465 19.3944
R3368 vdd.n2868 vdd.n465 19.3944
R3369 vdd.n2868 vdd.n463 19.3944
R3370 vdd.n2872 vdd.n463 19.3944
R3371 vdd.n2872 vdd.n453 19.3944
R3372 vdd.n2884 vdd.n453 19.3944
R3373 vdd.n2884 vdd.n451 19.3944
R3374 vdd.n2888 vdd.n451 19.3944
R3375 vdd.n2889 vdd.n2888 19.3944
R3376 vdd.n2890 vdd.n2889 19.3944
R3377 vdd.n2890 vdd.n449 19.3944
R3378 vdd.n2894 vdd.n449 19.3944
R3379 vdd.n2895 vdd.n2894 19.3944
R3380 vdd.n2896 vdd.n2895 19.3944
R3381 vdd.n2896 vdd.n446 19.3944
R3382 vdd.n2900 vdd.n446 19.3944
R3383 vdd.n2901 vdd.n2900 19.3944
R3384 vdd.n2902 vdd.n2901 19.3944
R3385 vdd.n2945 vdd.n404 19.3944
R3386 vdd.n2945 vdd.n410 19.3944
R3387 vdd.n2940 vdd.n410 19.3944
R3388 vdd.n2940 vdd.n2939 19.3944
R3389 vdd.n2939 vdd.n2938 19.3944
R3390 vdd.n2938 vdd.n417 19.3944
R3391 vdd.n2933 vdd.n417 19.3944
R3392 vdd.n2933 vdd.n2932 19.3944
R3393 vdd.n2932 vdd.n2931 19.3944
R3394 vdd.n2931 vdd.n424 19.3944
R3395 vdd.n2926 vdd.n424 19.3944
R3396 vdd.n2926 vdd.n2925 19.3944
R3397 vdd.n2925 vdd.n2924 19.3944
R3398 vdd.n2924 vdd.n431 19.3944
R3399 vdd.n2919 vdd.n431 19.3944
R3400 vdd.n2919 vdd.n2918 19.3944
R3401 vdd.n2918 vdd.n2917 19.3944
R3402 vdd.n2917 vdd.n438 19.3944
R3403 vdd.n2912 vdd.n438 19.3944
R3404 vdd.n2912 vdd.n2911 19.3944
R3405 vdd.n2984 vdd.n364 19.3944
R3406 vdd.n2984 vdd.n370 19.3944
R3407 vdd.n2979 vdd.n370 19.3944
R3408 vdd.n2979 vdd.n2978 19.3944
R3409 vdd.n2978 vdd.n2977 19.3944
R3410 vdd.n2977 vdd.n377 19.3944
R3411 vdd.n2972 vdd.n377 19.3944
R3412 vdd.n2972 vdd.n2971 19.3944
R3413 vdd.n2971 vdd.n2970 19.3944
R3414 vdd.n2970 vdd.n384 19.3944
R3415 vdd.n2965 vdd.n384 19.3944
R3416 vdd.n2965 vdd.n2964 19.3944
R3417 vdd.n2964 vdd.n2963 19.3944
R3418 vdd.n2963 vdd.n391 19.3944
R3419 vdd.n2958 vdd.n391 19.3944
R3420 vdd.n2958 vdd.n2957 19.3944
R3421 vdd.n2957 vdd.n2956 19.3944
R3422 vdd.n2956 vdd.n398 19.3944
R3423 vdd.n2951 vdd.n398 19.3944
R3424 vdd.n2951 vdd.n2950 19.3944
R3425 vdd.n3020 vdd.n3019 19.3944
R3426 vdd.n3019 vdd.n3018 19.3944
R3427 vdd.n3018 vdd.n336 19.3944
R3428 vdd.n337 vdd.n336 19.3944
R3429 vdd.n3011 vdd.n337 19.3944
R3430 vdd.n3011 vdd.n3010 19.3944
R3431 vdd.n3010 vdd.n3009 19.3944
R3432 vdd.n3009 vdd.n344 19.3944
R3433 vdd.n3004 vdd.n344 19.3944
R3434 vdd.n3004 vdd.n3003 19.3944
R3435 vdd.n3003 vdd.n3002 19.3944
R3436 vdd.n3002 vdd.n351 19.3944
R3437 vdd.n2997 vdd.n351 19.3944
R3438 vdd.n2997 vdd.n2996 19.3944
R3439 vdd.n2996 vdd.n2995 19.3944
R3440 vdd.n2995 vdd.n358 19.3944
R3441 vdd.n2990 vdd.n358 19.3944
R3442 vdd.n2990 vdd.n2989 19.3944
R3443 vdd.n2847 vdd.n480 19.3944
R3444 vdd.n2847 vdd.n471 19.3944
R3445 vdd.n2860 vdd.n471 19.3944
R3446 vdd.n2860 vdd.n469 19.3944
R3447 vdd.n2864 vdd.n469 19.3944
R3448 vdd.n2864 vdd.n460 19.3944
R3449 vdd.n2876 vdd.n460 19.3944
R3450 vdd.n2876 vdd.n458 19.3944
R3451 vdd.n2880 vdd.n458 19.3944
R3452 vdd.n2880 vdd.n300 19.3944
R3453 vdd.n3045 vdd.n300 19.3944
R3454 vdd.n3045 vdd.n301 19.3944
R3455 vdd.n3039 vdd.n301 19.3944
R3456 vdd.n3039 vdd.n3038 19.3944
R3457 vdd.n3038 vdd.n3037 19.3944
R3458 vdd.n3037 vdd.n313 19.3944
R3459 vdd.n3031 vdd.n313 19.3944
R3460 vdd.n3031 vdd.n3030 19.3944
R3461 vdd.n3030 vdd.n3029 19.3944
R3462 vdd.n3029 vdd.n324 19.3944
R3463 vdd.n3023 vdd.n324 19.3944
R3464 vdd.n2800 vdd.n536 19.3944
R3465 vdd.n2800 vdd.n2797 19.3944
R3466 vdd.n2797 vdd.n2794 19.3944
R3467 vdd.n2794 vdd.n2793 19.3944
R3468 vdd.n2793 vdd.n2790 19.3944
R3469 vdd.n2790 vdd.n2789 19.3944
R3470 vdd.n2789 vdd.n2786 19.3944
R3471 vdd.n2786 vdd.n2785 19.3944
R3472 vdd.n2785 vdd.n2782 19.3944
R3473 vdd.n2782 vdd.n2781 19.3944
R3474 vdd.n2781 vdd.n2778 19.3944
R3475 vdd.n2778 vdd.n2777 19.3944
R3476 vdd.n2777 vdd.n2774 19.3944
R3477 vdd.n2774 vdd.n2773 19.3944
R3478 vdd.n2773 vdd.n2770 19.3944
R3479 vdd.n2770 vdd.n2769 19.3944
R3480 vdd.n2769 vdd.n2766 19.3944
R3481 vdd.n2766 vdd.n2765 19.3944
R3482 vdd.n2765 vdd.n2762 19.3944
R3483 vdd.n2762 vdd.n2761 19.3944
R3484 vdd.n2843 vdd.n482 19.3944
R3485 vdd.n2838 vdd.n482 19.3944
R3486 vdd.n521 vdd.n518 19.3944
R3487 vdd.n2834 vdd.n2833 19.3944
R3488 vdd.n2833 vdd.n2830 19.3944
R3489 vdd.n2830 vdd.n2829 19.3944
R3490 vdd.n2829 vdd.n2826 19.3944
R3491 vdd.n2826 vdd.n2825 19.3944
R3492 vdd.n2825 vdd.n2822 19.3944
R3493 vdd.n2822 vdd.n2821 19.3944
R3494 vdd.n2821 vdd.n2818 19.3944
R3495 vdd.n2818 vdd.n2817 19.3944
R3496 vdd.n2817 vdd.n2814 19.3944
R3497 vdd.n2814 vdd.n2813 19.3944
R3498 vdd.n2813 vdd.n2810 19.3944
R3499 vdd.n2810 vdd.n2809 19.3944
R3500 vdd.n2754 vdd.n556 19.3944
R3501 vdd.n2754 vdd.n2751 19.3944
R3502 vdd.n2751 vdd.n2748 19.3944
R3503 vdd.n2748 vdd.n2747 19.3944
R3504 vdd.n2747 vdd.n2744 19.3944
R3505 vdd.n2744 vdd.n2743 19.3944
R3506 vdd.n2743 vdd.n2740 19.3944
R3507 vdd.n2740 vdd.n2739 19.3944
R3508 vdd.n2739 vdd.n2736 19.3944
R3509 vdd.n2736 vdd.n2735 19.3944
R3510 vdd.n2735 vdd.n2732 19.3944
R3511 vdd.n2732 vdd.n2731 19.3944
R3512 vdd.n2731 vdd.n2728 19.3944
R3513 vdd.n2728 vdd.n2727 19.3944
R3514 vdd.n2727 vdd.n2724 19.3944
R3515 vdd.n2724 vdd.n2723 19.3944
R3516 vdd.n2720 vdd.n2719 19.3944
R3517 vdd.n2716 vdd.n2715 19.3944
R3518 vdd.n1360 vdd.n1356 19.0066
R3519 vdd.n1652 vdd.n1583 19.0066
R3520 vdd.n2949 vdd.n404 19.0066
R3521 vdd.n2758 vdd.n556 19.0066
R3522 vdd.n1792 vdd.n1791 16.0975
R3523 vdd.n756 vdd.n755 16.0975
R3524 vdd.n1321 vdd.n1320 16.0975
R3525 vdd.n1359 vdd.n1358 16.0975
R3526 vdd.n1255 vdd.n1254 16.0975
R3527 vdd.n1948 vdd.n1947 16.0975
R3528 vdd.n1585 vdd.n1584 16.0975
R3529 vdd.n1545 vdd.n1544 16.0975
R3530 vdd.n1766 vdd.n1765 16.0975
R3531 vdd.n748 vdd.n747 16.0975
R3532 vdd.n2257 vdd.n2256 16.0975
R3533 vdd.n2909 vdd.n2908 16.0975
R3534 vdd.n406 vdd.n405 16.0975
R3535 vdd.n366 vdd.n365 16.0975
R3536 vdd.n558 vdd.n557 16.0975
R3537 vdd.n2805 vdd.n2804 16.0975
R3538 vdd.n623 vdd.n622 16.0975
R3539 vdd.n2254 vdd.n2253 16.0975
R3540 vdd.n2712 vdd.n2711 16.0975
R3541 vdd.n590 vdd.n589 16.0975
R3542 vdd.t165 vdd.n2218 15.4182
R3543 vdd.n2471 vdd.t155 15.4182
R3544 vdd.n28 vdd.n27 14.5674
R3545 vdd.n1989 vdd.n839 14.5112
R3546 vdd.n2673 vdd.n484 14.5112
R3547 vdd.n292 vdd.n257 13.1884
R3548 vdd.n245 vdd.n210 13.1884
R3549 vdd.n202 vdd.n167 13.1884
R3550 vdd.n155 vdd.n120 13.1884
R3551 vdd.n113 vdd.n78 13.1884
R3552 vdd.n66 vdd.n31 13.1884
R3553 vdd.n1107 vdd.n1072 13.1884
R3554 vdd.n1154 vdd.n1119 13.1884
R3555 vdd.n1017 vdd.n982 13.1884
R3556 vdd.n1064 vdd.n1029 13.1884
R3557 vdd.n928 vdd.n893 13.1884
R3558 vdd.n975 vdd.n940 13.1884
R3559 vdd.n1391 vdd.n1256 12.9944
R3560 vdd.n1395 vdd.n1256 12.9944
R3561 vdd.n1691 vdd.n1543 12.9944
R3562 vdd.n1692 vdd.n1691 12.9944
R3563 vdd.n2988 vdd.n364 12.9944
R3564 vdd.n2989 vdd.n2988 12.9944
R3565 vdd.n2806 vdd.n536 12.9944
R3566 vdd.n2809 vdd.n2806 12.9944
R3567 vdd.n293 vdd.n255 12.8005
R3568 vdd.n288 vdd.n259 12.8005
R3569 vdd.n246 vdd.n208 12.8005
R3570 vdd.n241 vdd.n212 12.8005
R3571 vdd.n203 vdd.n165 12.8005
R3572 vdd.n198 vdd.n169 12.8005
R3573 vdd.n156 vdd.n118 12.8005
R3574 vdd.n151 vdd.n122 12.8005
R3575 vdd.n114 vdd.n76 12.8005
R3576 vdd.n109 vdd.n80 12.8005
R3577 vdd.n67 vdd.n29 12.8005
R3578 vdd.n62 vdd.n33 12.8005
R3579 vdd.n1108 vdd.n1070 12.8005
R3580 vdd.n1103 vdd.n1074 12.8005
R3581 vdd.n1155 vdd.n1117 12.8005
R3582 vdd.n1150 vdd.n1121 12.8005
R3583 vdd.n1018 vdd.n980 12.8005
R3584 vdd.n1013 vdd.n984 12.8005
R3585 vdd.n1065 vdd.n1027 12.8005
R3586 vdd.n1060 vdd.n1031 12.8005
R3587 vdd.n929 vdd.n891 12.8005
R3588 vdd.n924 vdd.n895 12.8005
R3589 vdd.n976 vdd.n938 12.8005
R3590 vdd.n971 vdd.n942 12.8005
R3591 vdd.n287 vdd.n260 12.0247
R3592 vdd.n240 vdd.n213 12.0247
R3593 vdd.n197 vdd.n170 12.0247
R3594 vdd.n150 vdd.n123 12.0247
R3595 vdd.n108 vdd.n81 12.0247
R3596 vdd.n61 vdd.n34 12.0247
R3597 vdd.n1102 vdd.n1075 12.0247
R3598 vdd.n1149 vdd.n1122 12.0247
R3599 vdd.n1012 vdd.n985 12.0247
R3600 vdd.n1059 vdd.n1032 12.0247
R3601 vdd.n923 vdd.n896 12.0247
R3602 vdd.n970 vdd.n943 12.0247
R3603 vdd.n1430 vdd.n1186 11.337
R3604 vdd.n1439 vdd.n1186 11.337
R3605 vdd.n1439 vdd.n1438 11.337
R3606 vdd.n1447 vdd.n1180 11.337
R3607 vdd.n1456 vdd.n1455 11.337
R3608 vdd.n1473 vdd.n1164 11.337
R3609 vdd.n1481 vdd.n887 11.337
R3610 vdd.n1490 vdd.n1489 11.337
R3611 vdd.n1498 vdd.n870 11.337
R3612 vdd.n1509 vdd.n870 11.337
R3613 vdd.n1509 vdd.n1508 11.337
R3614 vdd.n2849 vdd.n473 11.337
R3615 vdd.n2858 vdd.n473 11.337
R3616 vdd.n2858 vdd.n2857 11.337
R3617 vdd.n2866 vdd.n467 11.337
R3618 vdd.n2882 vdd.n456 11.337
R3619 vdd.n3043 vdd.n304 11.337
R3620 vdd.n3041 vdd.n308 11.337
R3621 vdd.n3035 vdd.n3034 11.337
R3622 vdd.n3033 vdd.n318 11.337
R3623 vdd.n3027 vdd.n318 11.337
R3624 vdd.n3027 vdd.n3026 11.337
R3625 vdd.n284 vdd.n283 11.249
R3626 vdd.n237 vdd.n236 11.249
R3627 vdd.n194 vdd.n193 11.249
R3628 vdd.n147 vdd.n146 11.249
R3629 vdd.n105 vdd.n104 11.249
R3630 vdd.n58 vdd.n57 11.249
R3631 vdd.n1099 vdd.n1098 11.249
R3632 vdd.n1146 vdd.n1145 11.249
R3633 vdd.n1009 vdd.n1008 11.249
R3634 vdd.n1056 vdd.n1055 11.249
R3635 vdd.n920 vdd.n919 11.249
R3636 vdd.n967 vdd.n966 11.249
R3637 vdd.n2146 vdd.t184 11.1103
R3638 vdd.n2478 vdd.t170 11.1103
R3639 vdd.n1228 vdd.t32 10.7702
R3640 vdd.t43 vdd.n3025 10.7702
R3641 vdd.n269 vdd.n268 10.7238
R3642 vdd.n222 vdd.n221 10.7238
R3643 vdd.n179 vdd.n178 10.7238
R3644 vdd.n132 vdd.n131 10.7238
R3645 vdd.n90 vdd.n89 10.7238
R3646 vdd.n43 vdd.n42 10.7238
R3647 vdd.n1084 vdd.n1083 10.7238
R3648 vdd.n1131 vdd.n1130 10.7238
R3649 vdd.n994 vdd.n993 10.7238
R3650 vdd.n1041 vdd.n1040 10.7238
R3651 vdd.n905 vdd.n904 10.7238
R3652 vdd.n952 vdd.n951 10.7238
R3653 vdd.n1992 vdd.n1991 10.6151
R3654 vdd.n1993 vdd.n1992 10.6151
R3655 vdd.n1993 vdd.n825 10.6151
R3656 vdd.n2003 vdd.n825 10.6151
R3657 vdd.n2004 vdd.n2003 10.6151
R3658 vdd.n2005 vdd.n2004 10.6151
R3659 vdd.n2005 vdd.n812 10.6151
R3660 vdd.n2016 vdd.n812 10.6151
R3661 vdd.n2017 vdd.n2016 10.6151
R3662 vdd.n2018 vdd.n2017 10.6151
R3663 vdd.n2018 vdd.n800 10.6151
R3664 vdd.n2028 vdd.n800 10.6151
R3665 vdd.n2029 vdd.n2028 10.6151
R3666 vdd.n2030 vdd.n2029 10.6151
R3667 vdd.n2030 vdd.n788 10.6151
R3668 vdd.n2040 vdd.n788 10.6151
R3669 vdd.n2041 vdd.n2040 10.6151
R3670 vdd.n2042 vdd.n2041 10.6151
R3671 vdd.n2042 vdd.n777 10.6151
R3672 vdd.n2052 vdd.n777 10.6151
R3673 vdd.n2053 vdd.n2052 10.6151
R3674 vdd.n2054 vdd.n2053 10.6151
R3675 vdd.n2054 vdd.n764 10.6151
R3676 vdd.n2066 vdd.n764 10.6151
R3677 vdd.n2067 vdd.n2066 10.6151
R3678 vdd.n2069 vdd.n2067 10.6151
R3679 vdd.n2069 vdd.n2068 10.6151
R3680 vdd.n2068 vdd.n746 10.6151
R3681 vdd.n2216 vdd.n2215 10.6151
R3682 vdd.n2215 vdd.n2214 10.6151
R3683 vdd.n2214 vdd.n2211 10.6151
R3684 vdd.n2211 vdd.n2210 10.6151
R3685 vdd.n2210 vdd.n2207 10.6151
R3686 vdd.n2207 vdd.n2206 10.6151
R3687 vdd.n2206 vdd.n2203 10.6151
R3688 vdd.n2203 vdd.n2202 10.6151
R3689 vdd.n2202 vdd.n2199 10.6151
R3690 vdd.n2199 vdd.n2198 10.6151
R3691 vdd.n2198 vdd.n2195 10.6151
R3692 vdd.n2195 vdd.n2194 10.6151
R3693 vdd.n2194 vdd.n2191 10.6151
R3694 vdd.n2191 vdd.n2190 10.6151
R3695 vdd.n2190 vdd.n2187 10.6151
R3696 vdd.n2187 vdd.n2186 10.6151
R3697 vdd.n2186 vdd.n2183 10.6151
R3698 vdd.n2183 vdd.n2182 10.6151
R3699 vdd.n2182 vdd.n2179 10.6151
R3700 vdd.n2179 vdd.n2178 10.6151
R3701 vdd.n2178 vdd.n2175 10.6151
R3702 vdd.n2175 vdd.n2174 10.6151
R3703 vdd.n2174 vdd.n2171 10.6151
R3704 vdd.n2171 vdd.n2170 10.6151
R3705 vdd.n2170 vdd.n2167 10.6151
R3706 vdd.n2167 vdd.n2166 10.6151
R3707 vdd.n2166 vdd.n2163 10.6151
R3708 vdd.n2163 vdd.n2162 10.6151
R3709 vdd.n2162 vdd.n2159 10.6151
R3710 vdd.n2159 vdd.n2158 10.6151
R3711 vdd.n2158 vdd.n2155 10.6151
R3712 vdd.n2153 vdd.n2150 10.6151
R3713 vdd.n2150 vdd.n2149 10.6151
R3714 vdd.n1892 vdd.n1891 10.6151
R3715 vdd.n1891 vdd.n1889 10.6151
R3716 vdd.n1889 vdd.n1888 10.6151
R3717 vdd.n1888 vdd.n1886 10.6151
R3718 vdd.n1886 vdd.n1885 10.6151
R3719 vdd.n1885 vdd.n1883 10.6151
R3720 vdd.n1883 vdd.n1882 10.6151
R3721 vdd.n1882 vdd.n1880 10.6151
R3722 vdd.n1880 vdd.n1879 10.6151
R3723 vdd.n1879 vdd.n1877 10.6151
R3724 vdd.n1877 vdd.n1876 10.6151
R3725 vdd.n1876 vdd.n1874 10.6151
R3726 vdd.n1874 vdd.n1873 10.6151
R3727 vdd.n1873 vdd.n1788 10.6151
R3728 vdd.n1788 vdd.n1787 10.6151
R3729 vdd.n1787 vdd.n1785 10.6151
R3730 vdd.n1785 vdd.n1784 10.6151
R3731 vdd.n1784 vdd.n1782 10.6151
R3732 vdd.n1782 vdd.n1781 10.6151
R3733 vdd.n1781 vdd.n1779 10.6151
R3734 vdd.n1779 vdd.n1778 10.6151
R3735 vdd.n1778 vdd.n1776 10.6151
R3736 vdd.n1776 vdd.n1775 10.6151
R3737 vdd.n1775 vdd.n1773 10.6151
R3738 vdd.n1773 vdd.n1772 10.6151
R3739 vdd.n1772 vdd.n1769 10.6151
R3740 vdd.n1769 vdd.n1768 10.6151
R3741 vdd.n1768 vdd.n749 10.6151
R3742 vdd.n1726 vdd.n837 10.6151
R3743 vdd.n1727 vdd.n1726 10.6151
R3744 vdd.n1728 vdd.n1727 10.6151
R3745 vdd.n1728 vdd.n1722 10.6151
R3746 vdd.n1734 vdd.n1722 10.6151
R3747 vdd.n1735 vdd.n1734 10.6151
R3748 vdd.n1736 vdd.n1735 10.6151
R3749 vdd.n1736 vdd.n1720 10.6151
R3750 vdd.n1742 vdd.n1720 10.6151
R3751 vdd.n1743 vdd.n1742 10.6151
R3752 vdd.n1744 vdd.n1743 10.6151
R3753 vdd.n1744 vdd.n1718 10.6151
R3754 vdd.n1750 vdd.n1718 10.6151
R3755 vdd.n1751 vdd.n1750 10.6151
R3756 vdd.n1752 vdd.n1751 10.6151
R3757 vdd.n1752 vdd.n1716 10.6151
R3758 vdd.n1928 vdd.n1716 10.6151
R3759 vdd.n1928 vdd.n1927 10.6151
R3760 vdd.n1927 vdd.n1757 10.6151
R3761 vdd.n1921 vdd.n1757 10.6151
R3762 vdd.n1921 vdd.n1920 10.6151
R3763 vdd.n1920 vdd.n1919 10.6151
R3764 vdd.n1919 vdd.n1759 10.6151
R3765 vdd.n1913 vdd.n1759 10.6151
R3766 vdd.n1913 vdd.n1912 10.6151
R3767 vdd.n1912 vdd.n1911 10.6151
R3768 vdd.n1911 vdd.n1761 10.6151
R3769 vdd.n1905 vdd.n1761 10.6151
R3770 vdd.n1905 vdd.n1904 10.6151
R3771 vdd.n1904 vdd.n1903 10.6151
R3772 vdd.n1903 vdd.n1763 10.6151
R3773 vdd.n1897 vdd.n1896 10.6151
R3774 vdd.n1896 vdd.n1895 10.6151
R3775 vdd.n2401 vdd.n2400 10.6151
R3776 vdd.n2400 vdd.n2398 10.6151
R3777 vdd.n2398 vdd.n2397 10.6151
R3778 vdd.n2397 vdd.n2255 10.6151
R3779 vdd.n2344 vdd.n2255 10.6151
R3780 vdd.n2345 vdd.n2344 10.6151
R3781 vdd.n2347 vdd.n2345 10.6151
R3782 vdd.n2348 vdd.n2347 10.6151
R3783 vdd.n2350 vdd.n2348 10.6151
R3784 vdd.n2351 vdd.n2350 10.6151
R3785 vdd.n2353 vdd.n2351 10.6151
R3786 vdd.n2354 vdd.n2353 10.6151
R3787 vdd.n2356 vdd.n2354 10.6151
R3788 vdd.n2357 vdd.n2356 10.6151
R3789 vdd.n2372 vdd.n2357 10.6151
R3790 vdd.n2372 vdd.n2371 10.6151
R3791 vdd.n2371 vdd.n2370 10.6151
R3792 vdd.n2370 vdd.n2368 10.6151
R3793 vdd.n2368 vdd.n2367 10.6151
R3794 vdd.n2367 vdd.n2365 10.6151
R3795 vdd.n2365 vdd.n2364 10.6151
R3796 vdd.n2364 vdd.n2362 10.6151
R3797 vdd.n2362 vdd.n2361 10.6151
R3798 vdd.n2361 vdd.n2359 10.6151
R3799 vdd.n2359 vdd.n2358 10.6151
R3800 vdd.n2358 vdd.n626 10.6151
R3801 vdd.n2606 vdd.n626 10.6151
R3802 vdd.n2607 vdd.n2606 10.6151
R3803 vdd.n2468 vdd.n702 10.6151
R3804 vdd.n2468 vdd.n2467 10.6151
R3805 vdd.n2467 vdd.n2466 10.6151
R3806 vdd.n2466 vdd.n2464 10.6151
R3807 vdd.n2464 vdd.n2461 10.6151
R3808 vdd.n2461 vdd.n2460 10.6151
R3809 vdd.n2460 vdd.n2457 10.6151
R3810 vdd.n2457 vdd.n2456 10.6151
R3811 vdd.n2456 vdd.n2453 10.6151
R3812 vdd.n2453 vdd.n2452 10.6151
R3813 vdd.n2452 vdd.n2449 10.6151
R3814 vdd.n2449 vdd.n2448 10.6151
R3815 vdd.n2448 vdd.n2445 10.6151
R3816 vdd.n2445 vdd.n2444 10.6151
R3817 vdd.n2444 vdd.n2441 10.6151
R3818 vdd.n2441 vdd.n2440 10.6151
R3819 vdd.n2440 vdd.n2437 10.6151
R3820 vdd.n2437 vdd.n2436 10.6151
R3821 vdd.n2436 vdd.n2433 10.6151
R3822 vdd.n2433 vdd.n2432 10.6151
R3823 vdd.n2432 vdd.n2429 10.6151
R3824 vdd.n2429 vdd.n2428 10.6151
R3825 vdd.n2428 vdd.n2425 10.6151
R3826 vdd.n2425 vdd.n2424 10.6151
R3827 vdd.n2424 vdd.n2421 10.6151
R3828 vdd.n2421 vdd.n2420 10.6151
R3829 vdd.n2420 vdd.n2417 10.6151
R3830 vdd.n2417 vdd.n2416 10.6151
R3831 vdd.n2416 vdd.n2413 10.6151
R3832 vdd.n2413 vdd.n2412 10.6151
R3833 vdd.n2412 vdd.n2409 10.6151
R3834 vdd.n2407 vdd.n2404 10.6151
R3835 vdd.n2404 vdd.n2403 10.6151
R3836 vdd.n2481 vdd.n2480 10.6151
R3837 vdd.n2482 vdd.n2481 10.6151
R3838 vdd.n2482 vdd.n692 10.6151
R3839 vdd.n2492 vdd.n692 10.6151
R3840 vdd.n2493 vdd.n2492 10.6151
R3841 vdd.n2494 vdd.n2493 10.6151
R3842 vdd.n2494 vdd.n679 10.6151
R3843 vdd.n2504 vdd.n679 10.6151
R3844 vdd.n2505 vdd.n2504 10.6151
R3845 vdd.n2506 vdd.n2505 10.6151
R3846 vdd.n2506 vdd.n668 10.6151
R3847 vdd.n2516 vdd.n668 10.6151
R3848 vdd.n2517 vdd.n2516 10.6151
R3849 vdd.n2518 vdd.n2517 10.6151
R3850 vdd.n2518 vdd.n656 10.6151
R3851 vdd.n2528 vdd.n656 10.6151
R3852 vdd.n2529 vdd.n2528 10.6151
R3853 vdd.n2530 vdd.n2529 10.6151
R3854 vdd.n2530 vdd.n645 10.6151
R3855 vdd.n2542 vdd.n645 10.6151
R3856 vdd.n2543 vdd.n2542 10.6151
R3857 vdd.n2544 vdd.n2543 10.6151
R3858 vdd.n2544 vdd.n631 10.6151
R3859 vdd.n2599 vdd.n631 10.6151
R3860 vdd.n2600 vdd.n2599 10.6151
R3861 vdd.n2601 vdd.n2600 10.6151
R3862 vdd.n2601 vdd.n600 10.6151
R3863 vdd.n2671 vdd.n600 10.6151
R3864 vdd.n2670 vdd.n2669 10.6151
R3865 vdd.n2669 vdd.n601 10.6151
R3866 vdd.n602 vdd.n601 10.6151
R3867 vdd.n2662 vdd.n602 10.6151
R3868 vdd.n2662 vdd.n2661 10.6151
R3869 vdd.n2661 vdd.n2660 10.6151
R3870 vdd.n2660 vdd.n604 10.6151
R3871 vdd.n2655 vdd.n604 10.6151
R3872 vdd.n2655 vdd.n2654 10.6151
R3873 vdd.n2654 vdd.n2653 10.6151
R3874 vdd.n2653 vdd.n607 10.6151
R3875 vdd.n2648 vdd.n607 10.6151
R3876 vdd.n2648 vdd.n2647 10.6151
R3877 vdd.n2647 vdd.n2646 10.6151
R3878 vdd.n2646 vdd.n610 10.6151
R3879 vdd.n2641 vdd.n610 10.6151
R3880 vdd.n2641 vdd.n520 10.6151
R3881 vdd.n2637 vdd.n520 10.6151
R3882 vdd.n2637 vdd.n2636 10.6151
R3883 vdd.n2636 vdd.n2635 10.6151
R3884 vdd.n2635 vdd.n613 10.6151
R3885 vdd.n2630 vdd.n613 10.6151
R3886 vdd.n2630 vdd.n2629 10.6151
R3887 vdd.n2629 vdd.n2628 10.6151
R3888 vdd.n2628 vdd.n616 10.6151
R3889 vdd.n2623 vdd.n616 10.6151
R3890 vdd.n2623 vdd.n2622 10.6151
R3891 vdd.n2622 vdd.n2621 10.6151
R3892 vdd.n2621 vdd.n619 10.6151
R3893 vdd.n2616 vdd.n619 10.6151
R3894 vdd.n2616 vdd.n2615 10.6151
R3895 vdd.n2613 vdd.n624 10.6151
R3896 vdd.n2608 vdd.n624 10.6151
R3897 vdd.n2589 vdd.n2550 10.6151
R3898 vdd.n2584 vdd.n2550 10.6151
R3899 vdd.n2584 vdd.n2583 10.6151
R3900 vdd.n2583 vdd.n2582 10.6151
R3901 vdd.n2582 vdd.n2552 10.6151
R3902 vdd.n2577 vdd.n2552 10.6151
R3903 vdd.n2577 vdd.n2576 10.6151
R3904 vdd.n2576 vdd.n2575 10.6151
R3905 vdd.n2575 vdd.n2555 10.6151
R3906 vdd.n2570 vdd.n2555 10.6151
R3907 vdd.n2570 vdd.n2569 10.6151
R3908 vdd.n2569 vdd.n2568 10.6151
R3909 vdd.n2568 vdd.n2558 10.6151
R3910 vdd.n2563 vdd.n2558 10.6151
R3911 vdd.n2563 vdd.n2562 10.6151
R3912 vdd.n2562 vdd.n575 10.6151
R3913 vdd.n2706 vdd.n575 10.6151
R3914 vdd.n2706 vdd.n576 10.6151
R3915 vdd.n578 vdd.n576 10.6151
R3916 vdd.n2699 vdd.n578 10.6151
R3917 vdd.n2699 vdd.n2698 10.6151
R3918 vdd.n2698 vdd.n2697 10.6151
R3919 vdd.n2697 vdd.n580 10.6151
R3920 vdd.n2692 vdd.n580 10.6151
R3921 vdd.n2692 vdd.n2691 10.6151
R3922 vdd.n2691 vdd.n2690 10.6151
R3923 vdd.n2690 vdd.n583 10.6151
R3924 vdd.n2685 vdd.n583 10.6151
R3925 vdd.n2685 vdd.n2684 10.6151
R3926 vdd.n2684 vdd.n2683 10.6151
R3927 vdd.n2683 vdd.n586 10.6151
R3928 vdd.n2678 vdd.n2677 10.6151
R3929 vdd.n2677 vdd.n2676 10.6151
R3930 vdd.n2324 vdd.n2322 10.6151
R3931 vdd.n2325 vdd.n2324 10.6151
R3932 vdd.n2393 vdd.n2325 10.6151
R3933 vdd.n2393 vdd.n2392 10.6151
R3934 vdd.n2392 vdd.n2391 10.6151
R3935 vdd.n2391 vdd.n2389 10.6151
R3936 vdd.n2389 vdd.n2388 10.6151
R3937 vdd.n2388 vdd.n2386 10.6151
R3938 vdd.n2386 vdd.n2385 10.6151
R3939 vdd.n2385 vdd.n2383 10.6151
R3940 vdd.n2383 vdd.n2382 10.6151
R3941 vdd.n2382 vdd.n2380 10.6151
R3942 vdd.n2380 vdd.n2379 10.6151
R3943 vdd.n2379 vdd.n2377 10.6151
R3944 vdd.n2377 vdd.n2376 10.6151
R3945 vdd.n2376 vdd.n2342 10.6151
R3946 vdd.n2342 vdd.n2341 10.6151
R3947 vdd.n2341 vdd.n2339 10.6151
R3948 vdd.n2339 vdd.n2338 10.6151
R3949 vdd.n2338 vdd.n2336 10.6151
R3950 vdd.n2336 vdd.n2335 10.6151
R3951 vdd.n2335 vdd.n2333 10.6151
R3952 vdd.n2333 vdd.n2332 10.6151
R3953 vdd.n2332 vdd.n2330 10.6151
R3954 vdd.n2330 vdd.n2329 10.6151
R3955 vdd.n2329 vdd.n2327 10.6151
R3956 vdd.n2327 vdd.n2326 10.6151
R3957 vdd.n2326 vdd.n592 10.6151
R3958 vdd.n2475 vdd.n2474 10.6151
R3959 vdd.n2474 vdd.n707 10.6151
R3960 vdd.n2259 vdd.n707 10.6151
R3961 vdd.n2262 vdd.n2259 10.6151
R3962 vdd.n2263 vdd.n2262 10.6151
R3963 vdd.n2266 vdd.n2263 10.6151
R3964 vdd.n2267 vdd.n2266 10.6151
R3965 vdd.n2270 vdd.n2267 10.6151
R3966 vdd.n2271 vdd.n2270 10.6151
R3967 vdd.n2274 vdd.n2271 10.6151
R3968 vdd.n2275 vdd.n2274 10.6151
R3969 vdd.n2278 vdd.n2275 10.6151
R3970 vdd.n2279 vdd.n2278 10.6151
R3971 vdd.n2282 vdd.n2279 10.6151
R3972 vdd.n2283 vdd.n2282 10.6151
R3973 vdd.n2286 vdd.n2283 10.6151
R3974 vdd.n2287 vdd.n2286 10.6151
R3975 vdd.n2290 vdd.n2287 10.6151
R3976 vdd.n2291 vdd.n2290 10.6151
R3977 vdd.n2294 vdd.n2291 10.6151
R3978 vdd.n2295 vdd.n2294 10.6151
R3979 vdd.n2298 vdd.n2295 10.6151
R3980 vdd.n2299 vdd.n2298 10.6151
R3981 vdd.n2302 vdd.n2299 10.6151
R3982 vdd.n2303 vdd.n2302 10.6151
R3983 vdd.n2306 vdd.n2303 10.6151
R3984 vdd.n2307 vdd.n2306 10.6151
R3985 vdd.n2310 vdd.n2307 10.6151
R3986 vdd.n2311 vdd.n2310 10.6151
R3987 vdd.n2314 vdd.n2311 10.6151
R3988 vdd.n2315 vdd.n2314 10.6151
R3989 vdd.n2320 vdd.n2318 10.6151
R3990 vdd.n2321 vdd.n2320 10.6151
R3991 vdd.n2476 vdd.n697 10.6151
R3992 vdd.n2486 vdd.n697 10.6151
R3993 vdd.n2487 vdd.n2486 10.6151
R3994 vdd.n2488 vdd.n2487 10.6151
R3995 vdd.n2488 vdd.n685 10.6151
R3996 vdd.n2498 vdd.n685 10.6151
R3997 vdd.n2499 vdd.n2498 10.6151
R3998 vdd.n2500 vdd.n2499 10.6151
R3999 vdd.n2500 vdd.n674 10.6151
R4000 vdd.n2510 vdd.n674 10.6151
R4001 vdd.n2511 vdd.n2510 10.6151
R4002 vdd.n2512 vdd.n2511 10.6151
R4003 vdd.n2512 vdd.n662 10.6151
R4004 vdd.n2522 vdd.n662 10.6151
R4005 vdd.n2523 vdd.n2522 10.6151
R4006 vdd.n2524 vdd.n2523 10.6151
R4007 vdd.n2524 vdd.n651 10.6151
R4008 vdd.n2534 vdd.n651 10.6151
R4009 vdd.n2535 vdd.n2534 10.6151
R4010 vdd.n2538 vdd.n2535 10.6151
R4011 vdd.n2548 vdd.n639 10.6151
R4012 vdd.n2549 vdd.n2548 10.6151
R4013 vdd.n2595 vdd.n2549 10.6151
R4014 vdd.n2595 vdd.n2594 10.6151
R4015 vdd.n2594 vdd.n2593 10.6151
R4016 vdd.n2593 vdd.n2592 10.6151
R4017 vdd.n2592 vdd.n2590 10.6151
R4018 vdd.n1987 vdd.n831 10.6151
R4019 vdd.n1997 vdd.n831 10.6151
R4020 vdd.n1998 vdd.n1997 10.6151
R4021 vdd.n1999 vdd.n1998 10.6151
R4022 vdd.n1999 vdd.n818 10.6151
R4023 vdd.n2009 vdd.n818 10.6151
R4024 vdd.n2010 vdd.n2009 10.6151
R4025 vdd.n2012 vdd.n806 10.6151
R4026 vdd.n2022 vdd.n806 10.6151
R4027 vdd.n2023 vdd.n2022 10.6151
R4028 vdd.n2024 vdd.n2023 10.6151
R4029 vdd.n2024 vdd.n794 10.6151
R4030 vdd.n2034 vdd.n794 10.6151
R4031 vdd.n2035 vdd.n2034 10.6151
R4032 vdd.n2036 vdd.n2035 10.6151
R4033 vdd.n2036 vdd.n783 10.6151
R4034 vdd.n2046 vdd.n783 10.6151
R4035 vdd.n2047 vdd.n2046 10.6151
R4036 vdd.n2048 vdd.n2047 10.6151
R4037 vdd.n2048 vdd.n771 10.6151
R4038 vdd.n2058 vdd.n771 10.6151
R4039 vdd.n2059 vdd.n2058 10.6151
R4040 vdd.n2062 vdd.n2059 10.6151
R4041 vdd.n2062 vdd.n2061 10.6151
R4042 vdd.n2061 vdd.n2060 10.6151
R4043 vdd.n2060 vdd.n754 10.6151
R4044 vdd.n2144 vdd.n754 10.6151
R4045 vdd.n2143 vdd.n2142 10.6151
R4046 vdd.n2142 vdd.n2139 10.6151
R4047 vdd.n2139 vdd.n2138 10.6151
R4048 vdd.n2138 vdd.n2135 10.6151
R4049 vdd.n2135 vdd.n2134 10.6151
R4050 vdd.n2134 vdd.n2131 10.6151
R4051 vdd.n2131 vdd.n2130 10.6151
R4052 vdd.n2130 vdd.n2127 10.6151
R4053 vdd.n2127 vdd.n2126 10.6151
R4054 vdd.n2126 vdd.n2123 10.6151
R4055 vdd.n2123 vdd.n2122 10.6151
R4056 vdd.n2122 vdd.n2119 10.6151
R4057 vdd.n2119 vdd.n2118 10.6151
R4058 vdd.n2118 vdd.n2115 10.6151
R4059 vdd.n2115 vdd.n2114 10.6151
R4060 vdd.n2114 vdd.n2111 10.6151
R4061 vdd.n2111 vdd.n2110 10.6151
R4062 vdd.n2110 vdd.n2107 10.6151
R4063 vdd.n2107 vdd.n2106 10.6151
R4064 vdd.n2106 vdd.n2103 10.6151
R4065 vdd.n2103 vdd.n2102 10.6151
R4066 vdd.n2102 vdd.n2099 10.6151
R4067 vdd.n2099 vdd.n2098 10.6151
R4068 vdd.n2098 vdd.n2095 10.6151
R4069 vdd.n2095 vdd.n2094 10.6151
R4070 vdd.n2094 vdd.n2091 10.6151
R4071 vdd.n2091 vdd.n2090 10.6151
R4072 vdd.n2090 vdd.n2087 10.6151
R4073 vdd.n2087 vdd.n2086 10.6151
R4074 vdd.n2086 vdd.n2083 10.6151
R4075 vdd.n2083 vdd.n2082 10.6151
R4076 vdd.n2079 vdd.n2078 10.6151
R4077 vdd.n2078 vdd.n2076 10.6151
R4078 vdd.n1835 vdd.n1833 10.6151
R4079 vdd.n1836 vdd.n1835 10.6151
R4080 vdd.n1838 vdd.n1836 10.6151
R4081 vdd.n1839 vdd.n1838 10.6151
R4082 vdd.n1841 vdd.n1839 10.6151
R4083 vdd.n1842 vdd.n1841 10.6151
R4084 vdd.n1844 vdd.n1842 10.6151
R4085 vdd.n1845 vdd.n1844 10.6151
R4086 vdd.n1847 vdd.n1845 10.6151
R4087 vdd.n1848 vdd.n1847 10.6151
R4088 vdd.n1850 vdd.n1848 10.6151
R4089 vdd.n1851 vdd.n1850 10.6151
R4090 vdd.n1869 vdd.n1851 10.6151
R4091 vdd.n1869 vdd.n1868 10.6151
R4092 vdd.n1868 vdd.n1867 10.6151
R4093 vdd.n1867 vdd.n1865 10.6151
R4094 vdd.n1865 vdd.n1864 10.6151
R4095 vdd.n1864 vdd.n1862 10.6151
R4096 vdd.n1862 vdd.n1861 10.6151
R4097 vdd.n1861 vdd.n1859 10.6151
R4098 vdd.n1859 vdd.n1858 10.6151
R4099 vdd.n1858 vdd.n1856 10.6151
R4100 vdd.n1856 vdd.n1855 10.6151
R4101 vdd.n1855 vdd.n1853 10.6151
R4102 vdd.n1853 vdd.n1852 10.6151
R4103 vdd.n1852 vdd.n758 10.6151
R4104 vdd.n2074 vdd.n758 10.6151
R4105 vdd.n2075 vdd.n2074 10.6151
R4106 vdd.n1986 vdd.n1985 10.6151
R4107 vdd.n1985 vdd.n843 10.6151
R4108 vdd.n1979 vdd.n843 10.6151
R4109 vdd.n1979 vdd.n1978 10.6151
R4110 vdd.n1978 vdd.n1977 10.6151
R4111 vdd.n1977 vdd.n845 10.6151
R4112 vdd.n1971 vdd.n845 10.6151
R4113 vdd.n1971 vdd.n1970 10.6151
R4114 vdd.n1970 vdd.n1969 10.6151
R4115 vdd.n1969 vdd.n847 10.6151
R4116 vdd.n1963 vdd.n847 10.6151
R4117 vdd.n1963 vdd.n1962 10.6151
R4118 vdd.n1962 vdd.n1961 10.6151
R4119 vdd.n1961 vdd.n849 10.6151
R4120 vdd.n1955 vdd.n849 10.6151
R4121 vdd.n1955 vdd.n1954 10.6151
R4122 vdd.n1954 vdd.n1953 10.6151
R4123 vdd.n1953 vdd.n853 10.6151
R4124 vdd.n1801 vdd.n853 10.6151
R4125 vdd.n1802 vdd.n1801 10.6151
R4126 vdd.n1802 vdd.n1797 10.6151
R4127 vdd.n1808 vdd.n1797 10.6151
R4128 vdd.n1809 vdd.n1808 10.6151
R4129 vdd.n1810 vdd.n1809 10.6151
R4130 vdd.n1810 vdd.n1795 10.6151
R4131 vdd.n1816 vdd.n1795 10.6151
R4132 vdd.n1817 vdd.n1816 10.6151
R4133 vdd.n1818 vdd.n1817 10.6151
R4134 vdd.n1818 vdd.n1793 10.6151
R4135 vdd.n1824 vdd.n1793 10.6151
R4136 vdd.n1825 vdd.n1824 10.6151
R4137 vdd.n1827 vdd.n1789 10.6151
R4138 vdd.n1832 vdd.n1789 10.6151
R4139 vdd.n280 vdd.n262 10.4732
R4140 vdd.n233 vdd.n215 10.4732
R4141 vdd.n190 vdd.n172 10.4732
R4142 vdd.n143 vdd.n125 10.4732
R4143 vdd.n101 vdd.n83 10.4732
R4144 vdd.n54 vdd.n36 10.4732
R4145 vdd.n1095 vdd.n1077 10.4732
R4146 vdd.n1142 vdd.n1124 10.4732
R4147 vdd.n1005 vdd.n987 10.4732
R4148 vdd.n1052 vdd.n1034 10.4732
R4149 vdd.n916 vdd.n898 10.4732
R4150 vdd.n963 vdd.n945 10.4732
R4151 vdd.t96 vdd.n888 10.3167
R4152 vdd.n2874 vdd.t109 10.3167
R4153 vdd.n1465 vdd.t107 10.09
R4154 vdd.n3042 vdd.t122 10.09
R4155 vdd.n279 vdd.n264 9.69747
R4156 vdd.n232 vdd.n217 9.69747
R4157 vdd.n189 vdd.n174 9.69747
R4158 vdd.n142 vdd.n127 9.69747
R4159 vdd.n100 vdd.n85 9.69747
R4160 vdd.n53 vdd.n38 9.69747
R4161 vdd.n1094 vdd.n1079 9.69747
R4162 vdd.n1141 vdd.n1126 9.69747
R4163 vdd.n1004 vdd.n989 9.69747
R4164 vdd.n1051 vdd.n1036 9.69747
R4165 vdd.n915 vdd.n900 9.69747
R4166 vdd.n962 vdd.n947 9.69747
R4167 vdd.n1929 vdd.n1928 9.67831
R4168 vdd.n2836 vdd.n520 9.67831
R4169 vdd.n2707 vdd.n2706 9.67831
R4170 vdd.n1953 vdd.n1952 9.67831
R4171 vdd.n295 vdd.n294 9.45567
R4172 vdd.n248 vdd.n247 9.45567
R4173 vdd.n205 vdd.n204 9.45567
R4174 vdd.n158 vdd.n157 9.45567
R4175 vdd.n116 vdd.n115 9.45567
R4176 vdd.n69 vdd.n68 9.45567
R4177 vdd.n1110 vdd.n1109 9.45567
R4178 vdd.n1157 vdd.n1156 9.45567
R4179 vdd.n1020 vdd.n1019 9.45567
R4180 vdd.n1067 vdd.n1066 9.45567
R4181 vdd.n931 vdd.n930 9.45567
R4182 vdd.n978 vdd.n977 9.45567
R4183 vdd.n1689 vdd.n1543 9.3005
R4184 vdd.n1688 vdd.n1687 9.3005
R4185 vdd.n1549 vdd.n1548 9.3005
R4186 vdd.n1682 vdd.n1553 9.3005
R4187 vdd.n1681 vdd.n1554 9.3005
R4188 vdd.n1680 vdd.n1555 9.3005
R4189 vdd.n1559 vdd.n1556 9.3005
R4190 vdd.n1675 vdd.n1560 9.3005
R4191 vdd.n1674 vdd.n1561 9.3005
R4192 vdd.n1673 vdd.n1562 9.3005
R4193 vdd.n1566 vdd.n1563 9.3005
R4194 vdd.n1668 vdd.n1567 9.3005
R4195 vdd.n1667 vdd.n1568 9.3005
R4196 vdd.n1666 vdd.n1569 9.3005
R4197 vdd.n1573 vdd.n1570 9.3005
R4198 vdd.n1661 vdd.n1574 9.3005
R4199 vdd.n1660 vdd.n1575 9.3005
R4200 vdd.n1659 vdd.n1576 9.3005
R4201 vdd.n1580 vdd.n1577 9.3005
R4202 vdd.n1654 vdd.n1581 9.3005
R4203 vdd.n1653 vdd.n1582 9.3005
R4204 vdd.n1652 vdd.n1651 9.3005
R4205 vdd.n1650 vdd.n1583 9.3005
R4206 vdd.n1649 vdd.n1648 9.3005
R4207 vdd.n1589 vdd.n1588 9.3005
R4208 vdd.n1643 vdd.n1593 9.3005
R4209 vdd.n1642 vdd.n1594 9.3005
R4210 vdd.n1641 vdd.n1595 9.3005
R4211 vdd.n1599 vdd.n1596 9.3005
R4212 vdd.n1636 vdd.n1600 9.3005
R4213 vdd.n1635 vdd.n1601 9.3005
R4214 vdd.n1634 vdd.n1602 9.3005
R4215 vdd.n1606 vdd.n1603 9.3005
R4216 vdd.n1629 vdd.n1607 9.3005
R4217 vdd.n1628 vdd.n1608 9.3005
R4218 vdd.n1627 vdd.n1609 9.3005
R4219 vdd.n1611 vdd.n1610 9.3005
R4220 vdd.n1622 vdd.n854 9.3005
R4221 vdd.n1691 vdd.n1690 9.3005
R4222 vdd.n1715 vdd.n1714 9.3005
R4223 vdd.n1521 vdd.n1520 9.3005
R4224 vdd.n1526 vdd.n1524 9.3005
R4225 vdd.n1707 vdd.n1527 9.3005
R4226 vdd.n1706 vdd.n1528 9.3005
R4227 vdd.n1705 vdd.n1529 9.3005
R4228 vdd.n1533 vdd.n1530 9.3005
R4229 vdd.n1700 vdd.n1534 9.3005
R4230 vdd.n1699 vdd.n1535 9.3005
R4231 vdd.n1698 vdd.n1536 9.3005
R4232 vdd.n1540 vdd.n1537 9.3005
R4233 vdd.n1693 vdd.n1541 9.3005
R4234 vdd.n1692 vdd.n1542 9.3005
R4235 vdd.n1937 vdd.n1514 9.3005
R4236 vdd.n1939 vdd.n1938 9.3005
R4237 vdd.n1476 vdd.n1475 9.3005
R4238 vdd.n1477 vdd.n890 9.3005
R4239 vdd.n1479 vdd.n1478 9.3005
R4240 vdd.n880 vdd.n879 9.3005
R4241 vdd.n1493 vdd.n1492 9.3005
R4242 vdd.n1494 vdd.n878 9.3005
R4243 vdd.n1496 vdd.n1495 9.3005
R4244 vdd.n868 vdd.n867 9.3005
R4245 vdd.n1512 vdd.n1511 9.3005
R4246 vdd.n1513 vdd.n866 9.3005
R4247 vdd.n1941 vdd.n1940 9.3005
R4248 vdd.n271 vdd.n270 9.3005
R4249 vdd.n266 vdd.n265 9.3005
R4250 vdd.n277 vdd.n276 9.3005
R4251 vdd.n279 vdd.n278 9.3005
R4252 vdd.n262 vdd.n261 9.3005
R4253 vdd.n285 vdd.n284 9.3005
R4254 vdd.n287 vdd.n286 9.3005
R4255 vdd.n259 vdd.n256 9.3005
R4256 vdd.n294 vdd.n293 9.3005
R4257 vdd.n224 vdd.n223 9.3005
R4258 vdd.n219 vdd.n218 9.3005
R4259 vdd.n230 vdd.n229 9.3005
R4260 vdd.n232 vdd.n231 9.3005
R4261 vdd.n215 vdd.n214 9.3005
R4262 vdd.n238 vdd.n237 9.3005
R4263 vdd.n240 vdd.n239 9.3005
R4264 vdd.n212 vdd.n209 9.3005
R4265 vdd.n247 vdd.n246 9.3005
R4266 vdd.n181 vdd.n180 9.3005
R4267 vdd.n176 vdd.n175 9.3005
R4268 vdd.n187 vdd.n186 9.3005
R4269 vdd.n189 vdd.n188 9.3005
R4270 vdd.n172 vdd.n171 9.3005
R4271 vdd.n195 vdd.n194 9.3005
R4272 vdd.n197 vdd.n196 9.3005
R4273 vdd.n169 vdd.n166 9.3005
R4274 vdd.n204 vdd.n203 9.3005
R4275 vdd.n134 vdd.n133 9.3005
R4276 vdd.n129 vdd.n128 9.3005
R4277 vdd.n140 vdd.n139 9.3005
R4278 vdd.n142 vdd.n141 9.3005
R4279 vdd.n125 vdd.n124 9.3005
R4280 vdd.n148 vdd.n147 9.3005
R4281 vdd.n150 vdd.n149 9.3005
R4282 vdd.n122 vdd.n119 9.3005
R4283 vdd.n157 vdd.n156 9.3005
R4284 vdd.n92 vdd.n91 9.3005
R4285 vdd.n87 vdd.n86 9.3005
R4286 vdd.n98 vdd.n97 9.3005
R4287 vdd.n100 vdd.n99 9.3005
R4288 vdd.n83 vdd.n82 9.3005
R4289 vdd.n106 vdd.n105 9.3005
R4290 vdd.n108 vdd.n107 9.3005
R4291 vdd.n80 vdd.n77 9.3005
R4292 vdd.n115 vdd.n114 9.3005
R4293 vdd.n45 vdd.n44 9.3005
R4294 vdd.n40 vdd.n39 9.3005
R4295 vdd.n51 vdd.n50 9.3005
R4296 vdd.n53 vdd.n52 9.3005
R4297 vdd.n36 vdd.n35 9.3005
R4298 vdd.n59 vdd.n58 9.3005
R4299 vdd.n61 vdd.n60 9.3005
R4300 vdd.n33 vdd.n30 9.3005
R4301 vdd.n68 vdd.n67 9.3005
R4302 vdd.n2758 vdd.n2757 9.3005
R4303 vdd.n2761 vdd.n555 9.3005
R4304 vdd.n2762 vdd.n554 9.3005
R4305 vdd.n2765 vdd.n553 9.3005
R4306 vdd.n2766 vdd.n552 9.3005
R4307 vdd.n2769 vdd.n551 9.3005
R4308 vdd.n2770 vdd.n550 9.3005
R4309 vdd.n2773 vdd.n549 9.3005
R4310 vdd.n2774 vdd.n548 9.3005
R4311 vdd.n2777 vdd.n547 9.3005
R4312 vdd.n2778 vdd.n546 9.3005
R4313 vdd.n2781 vdd.n545 9.3005
R4314 vdd.n2782 vdd.n544 9.3005
R4315 vdd.n2785 vdd.n543 9.3005
R4316 vdd.n2786 vdd.n542 9.3005
R4317 vdd.n2789 vdd.n541 9.3005
R4318 vdd.n2790 vdd.n540 9.3005
R4319 vdd.n2793 vdd.n539 9.3005
R4320 vdd.n2794 vdd.n538 9.3005
R4321 vdd.n2797 vdd.n537 9.3005
R4322 vdd.n2801 vdd.n2800 9.3005
R4323 vdd.n2802 vdd.n536 9.3005
R4324 vdd.n2806 vdd.n2803 9.3005
R4325 vdd.n2809 vdd.n535 9.3005
R4326 vdd.n2810 vdd.n534 9.3005
R4327 vdd.n2813 vdd.n533 9.3005
R4328 vdd.n2814 vdd.n532 9.3005
R4329 vdd.n2817 vdd.n531 9.3005
R4330 vdd.n2818 vdd.n530 9.3005
R4331 vdd.n2821 vdd.n529 9.3005
R4332 vdd.n2822 vdd.n528 9.3005
R4333 vdd.n2825 vdd.n527 9.3005
R4334 vdd.n2826 vdd.n526 9.3005
R4335 vdd.n2829 vdd.n525 9.3005
R4336 vdd.n2830 vdd.n524 9.3005
R4337 vdd.n2833 vdd.n519 9.3005
R4338 vdd.n482 vdd.n481 9.3005
R4339 vdd.n2844 vdd.n2843 9.3005
R4340 vdd.n2847 vdd.n2846 9.3005
R4341 vdd.n471 vdd.n470 9.3005
R4342 vdd.n2861 vdd.n2860 9.3005
R4343 vdd.n2862 vdd.n469 9.3005
R4344 vdd.n2864 vdd.n2863 9.3005
R4345 vdd.n460 vdd.n459 9.3005
R4346 vdd.n2877 vdd.n2876 9.3005
R4347 vdd.n2878 vdd.n458 9.3005
R4348 vdd.n2880 vdd.n2879 9.3005
R4349 vdd.n300 vdd.n298 9.3005
R4350 vdd.n2845 vdd.n480 9.3005
R4351 vdd.n3046 vdd.n3045 9.3005
R4352 vdd.n301 vdd.n299 9.3005
R4353 vdd.n3039 vdd.n310 9.3005
R4354 vdd.n3038 vdd.n311 9.3005
R4355 vdd.n3037 vdd.n312 9.3005
R4356 vdd.n320 vdd.n313 9.3005
R4357 vdd.n3031 vdd.n321 9.3005
R4358 vdd.n3030 vdd.n322 9.3005
R4359 vdd.n3029 vdd.n323 9.3005
R4360 vdd.n331 vdd.n324 9.3005
R4361 vdd.n3023 vdd.n3022 9.3005
R4362 vdd.n3019 vdd.n332 9.3005
R4363 vdd.n3018 vdd.n335 9.3005
R4364 vdd.n339 vdd.n336 9.3005
R4365 vdd.n340 vdd.n337 9.3005
R4366 vdd.n3011 vdd.n341 9.3005
R4367 vdd.n3010 vdd.n342 9.3005
R4368 vdd.n3009 vdd.n343 9.3005
R4369 vdd.n347 vdd.n344 9.3005
R4370 vdd.n3004 vdd.n348 9.3005
R4371 vdd.n3003 vdd.n349 9.3005
R4372 vdd.n3002 vdd.n350 9.3005
R4373 vdd.n354 vdd.n351 9.3005
R4374 vdd.n2997 vdd.n355 9.3005
R4375 vdd.n2996 vdd.n356 9.3005
R4376 vdd.n2995 vdd.n357 9.3005
R4377 vdd.n361 vdd.n358 9.3005
R4378 vdd.n2990 vdd.n362 9.3005
R4379 vdd.n2989 vdd.n363 9.3005
R4380 vdd.n2988 vdd.n2987 9.3005
R4381 vdd.n2986 vdd.n364 9.3005
R4382 vdd.n2985 vdd.n2984 9.3005
R4383 vdd.n370 vdd.n369 9.3005
R4384 vdd.n2979 vdd.n374 9.3005
R4385 vdd.n2978 vdd.n375 9.3005
R4386 vdd.n2977 vdd.n376 9.3005
R4387 vdd.n380 vdd.n377 9.3005
R4388 vdd.n2972 vdd.n381 9.3005
R4389 vdd.n2971 vdd.n382 9.3005
R4390 vdd.n2970 vdd.n383 9.3005
R4391 vdd.n387 vdd.n384 9.3005
R4392 vdd.n2965 vdd.n388 9.3005
R4393 vdd.n2964 vdd.n389 9.3005
R4394 vdd.n2963 vdd.n390 9.3005
R4395 vdd.n394 vdd.n391 9.3005
R4396 vdd.n2958 vdd.n395 9.3005
R4397 vdd.n2957 vdd.n396 9.3005
R4398 vdd.n2956 vdd.n397 9.3005
R4399 vdd.n401 vdd.n398 9.3005
R4400 vdd.n2951 vdd.n402 9.3005
R4401 vdd.n2950 vdd.n403 9.3005
R4402 vdd.n2949 vdd.n2948 9.3005
R4403 vdd.n2947 vdd.n404 9.3005
R4404 vdd.n2946 vdd.n2945 9.3005
R4405 vdd.n410 vdd.n409 9.3005
R4406 vdd.n2940 vdd.n414 9.3005
R4407 vdd.n2939 vdd.n415 9.3005
R4408 vdd.n2938 vdd.n416 9.3005
R4409 vdd.n420 vdd.n417 9.3005
R4410 vdd.n2933 vdd.n421 9.3005
R4411 vdd.n2932 vdd.n422 9.3005
R4412 vdd.n2931 vdd.n423 9.3005
R4413 vdd.n427 vdd.n424 9.3005
R4414 vdd.n2926 vdd.n428 9.3005
R4415 vdd.n2925 vdd.n429 9.3005
R4416 vdd.n2924 vdd.n430 9.3005
R4417 vdd.n434 vdd.n431 9.3005
R4418 vdd.n2919 vdd.n435 9.3005
R4419 vdd.n2918 vdd.n436 9.3005
R4420 vdd.n2917 vdd.n437 9.3005
R4421 vdd.n441 vdd.n438 9.3005
R4422 vdd.n2912 vdd.n442 9.3005
R4423 vdd.n2911 vdd.n443 9.3005
R4424 vdd.n2907 vdd.n2904 9.3005
R4425 vdd.n3021 vdd.n3020 9.3005
R4426 vdd.n2852 vdd.n2851 9.3005
R4427 vdd.n2853 vdd.n475 9.3005
R4428 vdd.n2855 vdd.n2854 9.3005
R4429 vdd.n465 vdd.n464 9.3005
R4430 vdd.n2869 vdd.n2868 9.3005
R4431 vdd.n2870 vdd.n463 9.3005
R4432 vdd.n2872 vdd.n2871 9.3005
R4433 vdd.n453 vdd.n452 9.3005
R4434 vdd.n2885 vdd.n2884 9.3005
R4435 vdd.n2886 vdd.n451 9.3005
R4436 vdd.n2888 vdd.n2887 9.3005
R4437 vdd.n2889 vdd.n450 9.3005
R4438 vdd.n2891 vdd.n2890 9.3005
R4439 vdd.n2892 vdd.n449 9.3005
R4440 vdd.n2894 vdd.n2893 9.3005
R4441 vdd.n2895 vdd.n447 9.3005
R4442 vdd.n2897 vdd.n2896 9.3005
R4443 vdd.n2898 vdd.n446 9.3005
R4444 vdd.n2900 vdd.n2899 9.3005
R4445 vdd.n2901 vdd.n444 9.3005
R4446 vdd.n2903 vdd.n2902 9.3005
R4447 vdd.n477 vdd.n476 9.3005
R4448 vdd.n2710 vdd.n2709 9.3005
R4449 vdd.n2715 vdd.n2708 9.3005
R4450 vdd.n2724 vdd.n572 9.3005
R4451 vdd.n2727 vdd.n571 9.3005
R4452 vdd.n2728 vdd.n570 9.3005
R4453 vdd.n2731 vdd.n569 9.3005
R4454 vdd.n2732 vdd.n568 9.3005
R4455 vdd.n2735 vdd.n567 9.3005
R4456 vdd.n2736 vdd.n566 9.3005
R4457 vdd.n2739 vdd.n565 9.3005
R4458 vdd.n2740 vdd.n564 9.3005
R4459 vdd.n2743 vdd.n563 9.3005
R4460 vdd.n2744 vdd.n562 9.3005
R4461 vdd.n2747 vdd.n561 9.3005
R4462 vdd.n2748 vdd.n560 9.3005
R4463 vdd.n2751 vdd.n559 9.3005
R4464 vdd.n2755 vdd.n2754 9.3005
R4465 vdd.n2756 vdd.n556 9.3005
R4466 vdd.n1951 vdd.n1950 9.3005
R4467 vdd.n1946 vdd.n857 9.3005
R4468 vdd.n1433 vdd.n1432 9.3005
R4469 vdd.n1434 vdd.n1188 9.3005
R4470 vdd.n1436 vdd.n1435 9.3005
R4471 vdd.n1178 vdd.n1177 9.3005
R4472 vdd.n1450 vdd.n1449 9.3005
R4473 vdd.n1451 vdd.n1176 9.3005
R4474 vdd.n1453 vdd.n1452 9.3005
R4475 vdd.n1168 vdd.n1167 9.3005
R4476 vdd.n1468 vdd.n1467 9.3005
R4477 vdd.n1469 vdd.n1166 9.3005
R4478 vdd.n1471 vdd.n1470 9.3005
R4479 vdd.n885 vdd.n884 9.3005
R4480 vdd.n1484 vdd.n1483 9.3005
R4481 vdd.n1485 vdd.n883 9.3005
R4482 vdd.n1487 vdd.n1486 9.3005
R4483 vdd.n875 vdd.n874 9.3005
R4484 vdd.n1501 vdd.n1500 9.3005
R4485 vdd.n1502 vdd.n872 9.3005
R4486 vdd.n1506 vdd.n1505 9.3005
R4487 vdd.n1504 vdd.n873 9.3005
R4488 vdd.n1503 vdd.n862 9.3005
R4489 vdd.n1190 vdd.n1189 9.3005
R4490 vdd.n1326 vdd.n1325 9.3005
R4491 vdd.n1327 vdd.n1316 9.3005
R4492 vdd.n1329 vdd.n1328 9.3005
R4493 vdd.n1330 vdd.n1315 9.3005
R4494 vdd.n1332 vdd.n1331 9.3005
R4495 vdd.n1333 vdd.n1310 9.3005
R4496 vdd.n1335 vdd.n1334 9.3005
R4497 vdd.n1336 vdd.n1309 9.3005
R4498 vdd.n1338 vdd.n1337 9.3005
R4499 vdd.n1339 vdd.n1304 9.3005
R4500 vdd.n1341 vdd.n1340 9.3005
R4501 vdd.n1342 vdd.n1303 9.3005
R4502 vdd.n1344 vdd.n1343 9.3005
R4503 vdd.n1345 vdd.n1298 9.3005
R4504 vdd.n1347 vdd.n1346 9.3005
R4505 vdd.n1348 vdd.n1297 9.3005
R4506 vdd.n1350 vdd.n1349 9.3005
R4507 vdd.n1351 vdd.n1292 9.3005
R4508 vdd.n1353 vdd.n1352 9.3005
R4509 vdd.n1354 vdd.n1291 9.3005
R4510 vdd.n1356 vdd.n1355 9.3005
R4511 vdd.n1360 vdd.n1287 9.3005
R4512 vdd.n1362 vdd.n1361 9.3005
R4513 vdd.n1363 vdd.n1286 9.3005
R4514 vdd.n1365 vdd.n1364 9.3005
R4515 vdd.n1366 vdd.n1281 9.3005
R4516 vdd.n1368 vdd.n1367 9.3005
R4517 vdd.n1369 vdd.n1280 9.3005
R4518 vdd.n1371 vdd.n1370 9.3005
R4519 vdd.n1372 vdd.n1275 9.3005
R4520 vdd.n1374 vdd.n1373 9.3005
R4521 vdd.n1375 vdd.n1274 9.3005
R4522 vdd.n1377 vdd.n1376 9.3005
R4523 vdd.n1378 vdd.n1269 9.3005
R4524 vdd.n1380 vdd.n1379 9.3005
R4525 vdd.n1381 vdd.n1268 9.3005
R4526 vdd.n1383 vdd.n1382 9.3005
R4527 vdd.n1384 vdd.n1263 9.3005
R4528 vdd.n1386 vdd.n1385 9.3005
R4529 vdd.n1387 vdd.n1262 9.3005
R4530 vdd.n1389 vdd.n1388 9.3005
R4531 vdd.n1390 vdd.n1257 9.3005
R4532 vdd.n1392 vdd.n1391 9.3005
R4533 vdd.n1393 vdd.n1256 9.3005
R4534 vdd.n1395 vdd.n1394 9.3005
R4535 vdd.n1396 vdd.n1249 9.3005
R4536 vdd.n1398 vdd.n1397 9.3005
R4537 vdd.n1399 vdd.n1248 9.3005
R4538 vdd.n1401 vdd.n1400 9.3005
R4539 vdd.n1402 vdd.n1243 9.3005
R4540 vdd.n1404 vdd.n1403 9.3005
R4541 vdd.n1405 vdd.n1242 9.3005
R4542 vdd.n1407 vdd.n1406 9.3005
R4543 vdd.n1408 vdd.n1237 9.3005
R4544 vdd.n1410 vdd.n1409 9.3005
R4545 vdd.n1411 vdd.n1236 9.3005
R4546 vdd.n1413 vdd.n1412 9.3005
R4547 vdd.n1414 vdd.n1231 9.3005
R4548 vdd.n1416 vdd.n1415 9.3005
R4549 vdd.n1417 vdd.n1230 9.3005
R4550 vdd.n1419 vdd.n1418 9.3005
R4551 vdd.n1195 vdd.n1194 9.3005
R4552 vdd.n1425 vdd.n1424 9.3005
R4553 vdd.n1324 vdd.n1323 9.3005
R4554 vdd.n1428 vdd.n1427 9.3005
R4555 vdd.n1184 vdd.n1183 9.3005
R4556 vdd.n1442 vdd.n1441 9.3005
R4557 vdd.n1443 vdd.n1182 9.3005
R4558 vdd.n1445 vdd.n1444 9.3005
R4559 vdd.n1173 vdd.n1172 9.3005
R4560 vdd.n1459 vdd.n1458 9.3005
R4561 vdd.n1460 vdd.n1171 9.3005
R4562 vdd.n1463 vdd.n1462 9.3005
R4563 vdd.n1461 vdd.n1162 9.3005
R4564 vdd.n1426 vdd.n1193 9.3005
R4565 vdd.n1086 vdd.n1085 9.3005
R4566 vdd.n1081 vdd.n1080 9.3005
R4567 vdd.n1092 vdd.n1091 9.3005
R4568 vdd.n1094 vdd.n1093 9.3005
R4569 vdd.n1077 vdd.n1076 9.3005
R4570 vdd.n1100 vdd.n1099 9.3005
R4571 vdd.n1102 vdd.n1101 9.3005
R4572 vdd.n1074 vdd.n1071 9.3005
R4573 vdd.n1109 vdd.n1108 9.3005
R4574 vdd.n1133 vdd.n1132 9.3005
R4575 vdd.n1128 vdd.n1127 9.3005
R4576 vdd.n1139 vdd.n1138 9.3005
R4577 vdd.n1141 vdd.n1140 9.3005
R4578 vdd.n1124 vdd.n1123 9.3005
R4579 vdd.n1147 vdd.n1146 9.3005
R4580 vdd.n1149 vdd.n1148 9.3005
R4581 vdd.n1121 vdd.n1118 9.3005
R4582 vdd.n1156 vdd.n1155 9.3005
R4583 vdd.n996 vdd.n995 9.3005
R4584 vdd.n991 vdd.n990 9.3005
R4585 vdd.n1002 vdd.n1001 9.3005
R4586 vdd.n1004 vdd.n1003 9.3005
R4587 vdd.n987 vdd.n986 9.3005
R4588 vdd.n1010 vdd.n1009 9.3005
R4589 vdd.n1012 vdd.n1011 9.3005
R4590 vdd.n984 vdd.n981 9.3005
R4591 vdd.n1019 vdd.n1018 9.3005
R4592 vdd.n1043 vdd.n1042 9.3005
R4593 vdd.n1038 vdd.n1037 9.3005
R4594 vdd.n1049 vdd.n1048 9.3005
R4595 vdd.n1051 vdd.n1050 9.3005
R4596 vdd.n1034 vdd.n1033 9.3005
R4597 vdd.n1057 vdd.n1056 9.3005
R4598 vdd.n1059 vdd.n1058 9.3005
R4599 vdd.n1031 vdd.n1028 9.3005
R4600 vdd.n1066 vdd.n1065 9.3005
R4601 vdd.n907 vdd.n906 9.3005
R4602 vdd.n902 vdd.n901 9.3005
R4603 vdd.n913 vdd.n912 9.3005
R4604 vdd.n915 vdd.n914 9.3005
R4605 vdd.n898 vdd.n897 9.3005
R4606 vdd.n921 vdd.n920 9.3005
R4607 vdd.n923 vdd.n922 9.3005
R4608 vdd.n895 vdd.n892 9.3005
R4609 vdd.n930 vdd.n929 9.3005
R4610 vdd.n954 vdd.n953 9.3005
R4611 vdd.n949 vdd.n948 9.3005
R4612 vdd.n960 vdd.n959 9.3005
R4613 vdd.n962 vdd.n961 9.3005
R4614 vdd.n945 vdd.n944 9.3005
R4615 vdd.n968 vdd.n967 9.3005
R4616 vdd.n970 vdd.n969 9.3005
R4617 vdd.n942 vdd.n939 9.3005
R4618 vdd.n977 vdd.n976 9.3005
R4619 vdd.n1438 vdd.t101 8.95635
R4620 vdd.t14 vdd.n3033 8.95635
R4621 vdd.n276 vdd.n275 8.92171
R4622 vdd.n229 vdd.n228 8.92171
R4623 vdd.n186 vdd.n185 8.92171
R4624 vdd.n139 vdd.n138 8.92171
R4625 vdd.n97 vdd.n96 8.92171
R4626 vdd.n50 vdd.n49 8.92171
R4627 vdd.n1091 vdd.n1090 8.92171
R4628 vdd.n1138 vdd.n1137 8.92171
R4629 vdd.n1001 vdd.n1000 8.92171
R4630 vdd.n1048 vdd.n1047 8.92171
R4631 vdd.n912 vdd.n911 8.92171
R4632 vdd.n959 vdd.n958 8.92171
R4633 vdd.n207 vdd.n117 8.81535
R4634 vdd.n1069 vdd.n979 8.81535
R4635 vdd.n1465 vdd.t12 8.72962
R4636 vdd.t6 vdd.n3042 8.72962
R4637 vdd.n888 vdd.t8 8.50289
R4638 vdd.n1943 vdd.t28 8.50289
R4639 vdd.n516 vdd.t21 8.50289
R4640 vdd.n2874 vdd.t113 8.50289
R4641 vdd.n28 vdd.n14 8.42249
R4642 vdd.n3048 vdd.n3047 8.16225
R4643 vdd.n1161 vdd.n1160 8.16225
R4644 vdd.n272 vdd.n266 8.14595
R4645 vdd.n225 vdd.n219 8.14595
R4646 vdd.n182 vdd.n176 8.14595
R4647 vdd.n135 vdd.n129 8.14595
R4648 vdd.n93 vdd.n87 8.14595
R4649 vdd.n46 vdd.n40 8.14595
R4650 vdd.n1087 vdd.n1081 8.14595
R4651 vdd.n1134 vdd.n1128 8.14595
R4652 vdd.n997 vdd.n991 8.14595
R4653 vdd.n1044 vdd.n1038 8.14595
R4654 vdd.n908 vdd.n902 8.14595
R4655 vdd.n955 vdd.n949 8.14595
R4656 vdd.n2537 vdd.n639 8.11757
R4657 vdd.n2011 vdd.n2010 8.11757
R4658 vdd.n1989 vdd.n833 7.70933
R4659 vdd.n1995 vdd.n833 7.70933
R4660 vdd.n2001 vdd.n827 7.70933
R4661 vdd.n2001 vdd.n820 7.70933
R4662 vdd.n2007 vdd.n820 7.70933
R4663 vdd.n2007 vdd.n823 7.70933
R4664 vdd.n2014 vdd.n808 7.70933
R4665 vdd.n2020 vdd.n808 7.70933
R4666 vdd.n2026 vdd.n802 7.70933
R4667 vdd.n2032 vdd.n798 7.70933
R4668 vdd.n2038 vdd.n792 7.70933
R4669 vdd.n2050 vdd.n779 7.70933
R4670 vdd.n2056 vdd.n773 7.70933
R4671 vdd.n2056 vdd.n766 7.70933
R4672 vdd.n2064 vdd.n766 7.70933
R4673 vdd.n2071 vdd.t182 7.70933
R4674 vdd.n2146 vdd.t182 7.70933
R4675 vdd.n2478 vdd.t172 7.70933
R4676 vdd.n2484 vdd.t172 7.70933
R4677 vdd.n2490 vdd.n687 7.70933
R4678 vdd.n2496 vdd.n687 7.70933
R4679 vdd.n2496 vdd.n690 7.70933
R4680 vdd.n2502 vdd.n683 7.70933
R4681 vdd.n2514 vdd.n670 7.70933
R4682 vdd.n2520 vdd.n664 7.70933
R4683 vdd.n2526 vdd.n660 7.70933
R4684 vdd.n2532 vdd.n647 7.70933
R4685 vdd.n2540 vdd.n647 7.70933
R4686 vdd.n2546 vdd.n641 7.70933
R4687 vdd.n2546 vdd.n633 7.70933
R4688 vdd.n2597 vdd.n633 7.70933
R4689 vdd.n2597 vdd.n636 7.70933
R4690 vdd.n2603 vdd.n595 7.70933
R4691 vdd.n2673 vdd.n595 7.70933
R4692 vdd.n271 vdd.n268 7.3702
R4693 vdd.n224 vdd.n221 7.3702
R4694 vdd.n181 vdd.n178 7.3702
R4695 vdd.n134 vdd.n131 7.3702
R4696 vdd.n92 vdd.n89 7.3702
R4697 vdd.n45 vdd.n42 7.3702
R4698 vdd.n1086 vdd.n1083 7.3702
R4699 vdd.n1133 vdd.n1130 7.3702
R4700 vdd.n996 vdd.n993 7.3702
R4701 vdd.n1043 vdd.n1040 7.3702
R4702 vdd.n907 vdd.n904 7.3702
R4703 vdd.n954 vdd.n951 7.3702
R4704 vdd.n1361 vdd.n1360 6.98232
R4705 vdd.n1653 vdd.n1652 6.98232
R4706 vdd.n2950 vdd.n2949 6.98232
R4707 vdd.n2761 vdd.n2758 6.98232
R4708 vdd.n1498 vdd.t2 6.68904
R4709 vdd.n2857 vdd.t103 6.68904
R4710 vdd.t10 vdd.n887 6.46231
R4711 vdd.n2882 vdd.t117 6.46231
R4712 vdd.n1456 vdd.t105 6.23558
R4713 vdd.t0 vdd.n308 6.23558
R4714 vdd.n3048 vdd.n297 6.22547
R4715 vdd.n1160 vdd.n1159 6.22547
R4716 vdd.n2026 vdd.t186 6.00885
R4717 vdd.n2526 vdd.t176 6.00885
R4718 vdd.n823 vdd.t71 5.89549
R4719 vdd.t36 vdd.n641 5.89549
R4720 vdd.n272 vdd.n271 5.81868
R4721 vdd.n225 vdd.n224 5.81868
R4722 vdd.n182 vdd.n181 5.81868
R4723 vdd.n135 vdd.n134 5.81868
R4724 vdd.n93 vdd.n92 5.81868
R4725 vdd.n46 vdd.n45 5.81868
R4726 vdd.n1087 vdd.n1086 5.81868
R4727 vdd.n1134 vdd.n1133 5.81868
R4728 vdd.n997 vdd.n996 5.81868
R4729 vdd.n1044 vdd.n1043 5.81868
R4730 vdd.n908 vdd.n907 5.81868
R4731 vdd.n955 vdd.n954 5.81868
R4732 vdd.t17 vdd.n827 5.78212
R4733 vdd.n1770 vdd.t53 5.78212
R4734 vdd.n2395 vdd.t61 5.78212
R4735 vdd.n636 vdd.t57 5.78212
R4736 vdd.n2154 vdd.n2153 5.77611
R4737 vdd.n1897 vdd.n1767 5.77611
R4738 vdd.n2408 vdd.n2407 5.77611
R4739 vdd.n2614 vdd.n2613 5.77611
R4740 vdd.n2678 vdd.n591 5.77611
R4741 vdd.n2318 vdd.n2258 5.77611
R4742 vdd.n2079 vdd.n757 5.77611
R4743 vdd.n1827 vdd.n1826 5.77611
R4744 vdd.n1323 vdd.n1322 5.62474
R4745 vdd.n1949 vdd.n1946 5.62474
R4746 vdd.n2910 vdd.n2907 5.62474
R4747 vdd.n2713 vdd.n2710 5.62474
R4748 vdd.t147 vdd.n779 5.44203
R4749 vdd.n683 vdd.t180 5.44203
R4750 vdd.n1180 vdd.t105 5.10193
R4751 vdd.t157 vdd.n802 5.10193
R4752 vdd.n792 vdd.t167 5.10193
R4753 vdd.t177 vdd.n670 5.10193
R4754 vdd.n660 vdd.t162 5.10193
R4755 vdd.n3035 vdd.t0 5.10193
R4756 vdd.n275 vdd.n266 5.04292
R4757 vdd.n228 vdd.n219 5.04292
R4758 vdd.n185 vdd.n176 5.04292
R4759 vdd.n138 vdd.n129 5.04292
R4760 vdd.n96 vdd.n87 5.04292
R4761 vdd.n49 vdd.n40 5.04292
R4762 vdd.n1090 vdd.n1081 5.04292
R4763 vdd.n1137 vdd.n1128 5.04292
R4764 vdd.n1000 vdd.n991 5.04292
R4765 vdd.n1047 vdd.n1038 5.04292
R4766 vdd.n911 vdd.n902 5.04292
R4767 vdd.n958 vdd.n949 5.04292
R4768 vdd.n1473 vdd.t10 4.8752
R4769 vdd.t154 vdd.t163 4.8752
R4770 vdd.t146 vdd.t174 4.8752
R4771 vdd.t168 vdd.t149 4.8752
R4772 vdd.t187 vdd.t145 4.8752
R4773 vdd.t117 vdd.n304 4.8752
R4774 vdd.n2155 vdd.n2154 4.83952
R4775 vdd.n1767 vdd.n1763 4.83952
R4776 vdd.n2409 vdd.n2408 4.83952
R4777 vdd.n2615 vdd.n2614 4.83952
R4778 vdd.n591 vdd.n586 4.83952
R4779 vdd.n2315 vdd.n2258 4.83952
R4780 vdd.n2082 vdd.n757 4.83952
R4781 vdd.n1826 vdd.n1825 4.83952
R4782 vdd.n1621 vdd.n855 4.74817
R4783 vdd.n1616 vdd.n856 4.74817
R4784 vdd.n1518 vdd.n1515 4.74817
R4785 vdd.n1930 vdd.n1519 4.74817
R4786 vdd.n1932 vdd.n1518 4.74817
R4787 vdd.n1931 vdd.n1930 4.74817
R4788 vdd.n2838 vdd.n2837 4.74817
R4789 vdd.n2835 vdd.n2834 4.74817
R4790 vdd.n2835 vdd.n521 4.74817
R4791 vdd.n2837 vdd.n518 4.74817
R4792 vdd.n2720 vdd.n573 4.74817
R4793 vdd.n2716 vdd.n574 4.74817
R4794 vdd.n2719 vdd.n574 4.74817
R4795 vdd.n2723 vdd.n573 4.74817
R4796 vdd.n1617 vdd.n855 4.74817
R4797 vdd.n858 vdd.n856 4.74817
R4798 vdd.n297 vdd.n296 4.7074
R4799 vdd.n207 vdd.n206 4.7074
R4800 vdd.n1159 vdd.n1158 4.7074
R4801 vdd.n1069 vdd.n1068 4.7074
R4802 vdd.n1489 vdd.t2 4.64847
R4803 vdd.n2866 vdd.t103 4.64847
R4804 vdd.n2032 vdd.t178 4.53511
R4805 vdd.n2520 vdd.t158 4.53511
R4806 vdd.n2064 vdd.t160 4.30838
R4807 vdd.n2490 vdd.t150 4.30838
R4808 vdd.n276 vdd.n264 4.26717
R4809 vdd.n229 vdd.n217 4.26717
R4810 vdd.n186 vdd.n174 4.26717
R4811 vdd.n139 vdd.n127 4.26717
R4812 vdd.n97 vdd.n85 4.26717
R4813 vdd.n50 vdd.n38 4.26717
R4814 vdd.n1091 vdd.n1079 4.26717
R4815 vdd.n1138 vdd.n1126 4.26717
R4816 vdd.n1001 vdd.n989 4.26717
R4817 vdd.n1048 vdd.n1036 4.26717
R4818 vdd.n912 vdd.n900 4.26717
R4819 vdd.n959 vdd.n947 4.26717
R4820 vdd.n297 vdd.n207 4.10845
R4821 vdd.n1159 vdd.n1069 4.10845
R4822 vdd.n253 vdd.t123 4.06363
R4823 vdd.n253 vdd.t1 4.06363
R4824 vdd.n251 vdd.t140 4.06363
R4825 vdd.n251 vdd.t197 4.06363
R4826 vdd.n249 vdd.t114 4.06363
R4827 vdd.n249 vdd.t110 4.06363
R4828 vdd.n163 vdd.t191 4.06363
R4829 vdd.n163 vdd.t199 4.06363
R4830 vdd.n161 vdd.t134 4.06363
R4831 vdd.n161 vdd.t136 4.06363
R4832 vdd.n159 vdd.t143 4.06363
R4833 vdd.n159 vdd.t116 4.06363
R4834 vdd.n74 vdd.t139 4.06363
R4835 vdd.n74 vdd.t195 4.06363
R4836 vdd.n72 vdd.t118 4.06363
R4837 vdd.n72 vdd.t7 4.06363
R4838 vdd.n70 vdd.t190 4.06363
R4839 vdd.n70 vdd.t135 4.06363
R4840 vdd.n1111 vdd.t137 4.06363
R4841 vdd.n1111 vdd.t119 4.06363
R4842 vdd.n1113 vdd.t13 4.06363
R4843 vdd.n1113 vdd.t115 4.06363
R4844 vdd.n1115 vdd.t144 4.06363
R4845 vdd.n1115 vdd.t120 4.06363
R4846 vdd.n1021 vdd.t97 4.06363
R4847 vdd.n1021 vdd.t9 4.06363
R4848 vdd.n1023 vdd.t124 4.06363
R4849 vdd.n1023 vdd.t11 4.06363
R4850 vdd.n1025 vdd.t106 4.06363
R4851 vdd.n1025 vdd.t108 4.06363
R4852 vdd.n932 vdd.t192 4.06363
R4853 vdd.n932 vdd.t189 4.06363
R4854 vdd.n934 vdd.t141 4.06363
R4855 vdd.n934 vdd.t198 4.06363
R4856 vdd.n936 vdd.t196 4.06363
R4857 vdd.n936 vdd.t194 4.06363
R4858 vdd.n26 vdd.t99 3.9605
R4859 vdd.n26 vdd.t93 3.9605
R4860 vdd.n23 vdd.t129 3.9605
R4861 vdd.n23 vdd.t130 3.9605
R4862 vdd.n21 vdd.t4 3.9605
R4863 vdd.n21 vdd.t94 3.9605
R4864 vdd.n20 vdd.t131 3.9605
R4865 vdd.n20 vdd.t128 3.9605
R4866 vdd.n15 vdd.t92 3.9605
R4867 vdd.n15 vdd.t98 3.9605
R4868 vdd.n16 vdd.t126 3.9605
R4869 vdd.n16 vdd.t127 3.9605
R4870 vdd.n18 vdd.t5 3.9605
R4871 vdd.n18 vdd.t100 3.9605
R4872 vdd.n25 vdd.t95 3.9605
R4873 vdd.n25 vdd.t125 3.9605
R4874 vdd.n7 vdd.t188 3.61217
R4875 vdd.n7 vdd.t159 3.61217
R4876 vdd.n8 vdd.t169 3.61217
R4877 vdd.n8 vdd.t181 3.61217
R4878 vdd.n10 vdd.t173 3.61217
R4879 vdd.n10 vdd.t151 3.61217
R4880 vdd.n12 vdd.t156 3.61217
R4881 vdd.n12 vdd.t171 3.61217
R4882 vdd.n5 vdd.t185 3.61217
R4883 vdd.n5 vdd.t166 3.61217
R4884 vdd.n3 vdd.t161 3.61217
R4885 vdd.n3 vdd.t183 3.61217
R4886 vdd.n1 vdd.t148 3.61217
R4887 vdd.n1 vdd.t175 3.61217
R4888 vdd.n0 vdd.t179 3.61217
R4889 vdd.n0 vdd.t164 3.61217
R4890 vdd.n280 vdd.n279 3.49141
R4891 vdd.n233 vdd.n232 3.49141
R4892 vdd.n190 vdd.n189 3.49141
R4893 vdd.n143 vdd.n142 3.49141
R4894 vdd.n101 vdd.n100 3.49141
R4895 vdd.n54 vdd.n53 3.49141
R4896 vdd.n1095 vdd.n1094 3.49141
R4897 vdd.n1142 vdd.n1141 3.49141
R4898 vdd.n1005 vdd.n1004 3.49141
R4899 vdd.n1052 vdd.n1051 3.49141
R4900 vdd.n916 vdd.n915 3.49141
R4901 vdd.n963 vdd.n962 3.49141
R4902 vdd.n1770 vdd.t160 3.40145
R4903 vdd.n2218 vdd.t184 3.40145
R4904 vdd.n2471 vdd.t170 3.40145
R4905 vdd.n2395 vdd.t150 3.40145
R4906 vdd.n1871 vdd.t178 3.17472
R4907 vdd.n2374 vdd.t158 3.17472
R4908 vdd.n1490 vdd.t8 2.83463
R4909 vdd.n1508 vdd.t28 2.83463
R4910 vdd.n2849 vdd.t21 2.83463
R4911 vdd.n467 vdd.t113 2.83463
R4912 vdd.n283 vdd.n262 2.71565
R4913 vdd.n236 vdd.n215 2.71565
R4914 vdd.n193 vdd.n172 2.71565
R4915 vdd.n146 vdd.n125 2.71565
R4916 vdd.n104 vdd.n83 2.71565
R4917 vdd.n57 vdd.n36 2.71565
R4918 vdd.n1098 vdd.n1077 2.71565
R4919 vdd.n1145 vdd.n1124 2.71565
R4920 vdd.n1008 vdd.n987 2.71565
R4921 vdd.n1055 vdd.n1034 2.71565
R4922 vdd.n919 vdd.n898 2.71565
R4923 vdd.n966 vdd.n945 2.71565
R4924 vdd.t12 vdd.n1164 2.6079
R4925 vdd.n2020 vdd.t157 2.6079
R4926 vdd.n2044 vdd.t167 2.6079
R4927 vdd.n2508 vdd.t177 2.6079
R4928 vdd.n2532 vdd.t162 2.6079
R4929 vdd.n3043 vdd.t6 2.6079
R4930 vdd.n2538 vdd.n2537 2.49806
R4931 vdd.n2012 vdd.n2011 2.49806
R4932 vdd.n270 vdd.n269 2.4129
R4933 vdd.n223 vdd.n222 2.4129
R4934 vdd.n180 vdd.n179 2.4129
R4935 vdd.n133 vdd.n132 2.4129
R4936 vdd.n91 vdd.n90 2.4129
R4937 vdd.n44 vdd.n43 2.4129
R4938 vdd.n1085 vdd.n1084 2.4129
R4939 vdd.n1132 vdd.n1131 2.4129
R4940 vdd.n995 vdd.n994 2.4129
R4941 vdd.n1042 vdd.n1041 2.4129
R4942 vdd.n906 vdd.n905 2.4129
R4943 vdd.n953 vdd.n952 2.4129
R4944 vdd.n1447 vdd.t101 2.38117
R4945 vdd.n3034 vdd.t14 2.38117
R4946 vdd.n1929 vdd.n1518 2.27742
R4947 vdd.n1930 vdd.n1929 2.27742
R4948 vdd.n2836 vdd.n2835 2.27742
R4949 vdd.n2837 vdd.n2836 2.27742
R4950 vdd.n2707 vdd.n574 2.27742
R4951 vdd.n2707 vdd.n573 2.27742
R4952 vdd.n1952 vdd.n855 2.27742
R4953 vdd.n1952 vdd.n856 2.27742
R4954 vdd.n2044 vdd.t147 2.2678
R4955 vdd.n2508 vdd.t180 2.2678
R4956 vdd.t174 vdd.n773 2.04107
R4957 vdd.n690 vdd.t168 2.04107
R4958 vdd.n284 vdd.n260 1.93989
R4959 vdd.n237 vdd.n213 1.93989
R4960 vdd.n194 vdd.n170 1.93989
R4961 vdd.n147 vdd.n123 1.93989
R4962 vdd.n105 vdd.n81 1.93989
R4963 vdd.n58 vdd.n34 1.93989
R4964 vdd.n1099 vdd.n1075 1.93989
R4965 vdd.n1146 vdd.n1122 1.93989
R4966 vdd.n1009 vdd.n985 1.93989
R4967 vdd.n1056 vdd.n1032 1.93989
R4968 vdd.n920 vdd.n896 1.93989
R4969 vdd.n967 vdd.n943 1.93989
R4970 vdd.n1995 vdd.t17 1.92771
R4971 vdd.n2071 vdd.t53 1.92771
R4972 vdd.n2484 vdd.t61 1.92771
R4973 vdd.n2603 vdd.t57 1.92771
R4974 vdd.n1871 vdd.t186 1.70098
R4975 vdd.n798 vdd.t154 1.70098
R4976 vdd.t145 vdd.n664 1.70098
R4977 vdd.n2374 vdd.t176 1.70098
R4978 vdd.n1455 vdd.t107 1.24752
R4979 vdd.t122 vdd.n3041 1.24752
R4980 vdd.n295 vdd.n255 1.16414
R4981 vdd.n288 vdd.n287 1.16414
R4982 vdd.n248 vdd.n208 1.16414
R4983 vdd.n241 vdd.n240 1.16414
R4984 vdd.n205 vdd.n165 1.16414
R4985 vdd.n198 vdd.n197 1.16414
R4986 vdd.n158 vdd.n118 1.16414
R4987 vdd.n151 vdd.n150 1.16414
R4988 vdd.n116 vdd.n76 1.16414
R4989 vdd.n109 vdd.n108 1.16414
R4990 vdd.n69 vdd.n29 1.16414
R4991 vdd.n62 vdd.n61 1.16414
R4992 vdd.n1110 vdd.n1070 1.16414
R4993 vdd.n1103 vdd.n1102 1.16414
R4994 vdd.n1157 vdd.n1117 1.16414
R4995 vdd.n1150 vdd.n1149 1.16414
R4996 vdd.n1020 vdd.n980 1.16414
R4997 vdd.n1013 vdd.n1012 1.16414
R4998 vdd.n1067 vdd.n1027 1.16414
R4999 vdd.n1060 vdd.n1059 1.16414
R5000 vdd.n931 vdd.n891 1.16414
R5001 vdd.n924 vdd.n923 1.16414
R5002 vdd.n978 vdd.n938 1.16414
R5003 vdd.n971 vdd.n970 1.16414
R5004 vdd.n2038 vdd.t163 1.13415
R5005 vdd.n2514 vdd.t187 1.13415
R5006 vdd.n1481 vdd.t96 1.02079
R5007 vdd.t71 vdd.t152 1.02079
R5008 vdd.t153 vdd.t36 1.02079
R5009 vdd.t109 vdd.n456 1.02079
R5010 vdd.n1326 vdd.n1322 0.970197
R5011 vdd.n1950 vdd.n1949 0.970197
R5012 vdd.n2911 vdd.n2910 0.970197
R5013 vdd.n2715 vdd.n2713 0.970197
R5014 vdd.n2014 vdd.t152 0.794056
R5015 vdd.n2050 vdd.t146 0.794056
R5016 vdd.n2502 vdd.t149 0.794056
R5017 vdd.n2540 vdd.t153 0.794056
R5018 vdd.n1160 vdd.n28 0.74827
R5019 vdd vdd.n3048 0.740437
R5020 vdd.n1430 vdd.t32 0.567326
R5021 vdd.n3026 vdd.t43 0.567326
R5022 vdd.n1940 vdd.n1939 0.537085
R5023 vdd.n2845 vdd.n2844 0.537085
R5024 vdd.n3022 vdd.n3021 0.537085
R5025 vdd.n2904 vdd.n2903 0.537085
R5026 vdd.n2709 vdd.n476 0.537085
R5027 vdd.n1503 vdd.n857 0.537085
R5028 vdd.n1324 vdd.n1189 0.537085
R5029 vdd.n1426 vdd.n1425 0.537085
R5030 vdd.n4 vdd.n2 0.459552
R5031 vdd.n11 vdd.n9 0.459552
R5032 vdd.n293 vdd.n292 0.388379
R5033 vdd.n259 vdd.n257 0.388379
R5034 vdd.n246 vdd.n245 0.388379
R5035 vdd.n212 vdd.n210 0.388379
R5036 vdd.n203 vdd.n202 0.388379
R5037 vdd.n169 vdd.n167 0.388379
R5038 vdd.n156 vdd.n155 0.388379
R5039 vdd.n122 vdd.n120 0.388379
R5040 vdd.n114 vdd.n113 0.388379
R5041 vdd.n80 vdd.n78 0.388379
R5042 vdd.n67 vdd.n66 0.388379
R5043 vdd.n33 vdd.n31 0.388379
R5044 vdd.n1108 vdd.n1107 0.388379
R5045 vdd.n1074 vdd.n1072 0.388379
R5046 vdd.n1155 vdd.n1154 0.388379
R5047 vdd.n1121 vdd.n1119 0.388379
R5048 vdd.n1018 vdd.n1017 0.388379
R5049 vdd.n984 vdd.n982 0.388379
R5050 vdd.n1065 vdd.n1064 0.388379
R5051 vdd.n1031 vdd.n1029 0.388379
R5052 vdd.n929 vdd.n928 0.388379
R5053 vdd.n895 vdd.n893 0.388379
R5054 vdd.n976 vdd.n975 0.388379
R5055 vdd.n942 vdd.n940 0.388379
R5056 vdd.n19 vdd.n17 0.387128
R5057 vdd.n24 vdd.n22 0.387128
R5058 vdd.n6 vdd.n4 0.358259
R5059 vdd.n13 vdd.n11 0.358259
R5060 vdd.n252 vdd.n250 0.358259
R5061 vdd.n254 vdd.n252 0.358259
R5062 vdd.n296 vdd.n254 0.358259
R5063 vdd.n162 vdd.n160 0.358259
R5064 vdd.n164 vdd.n162 0.358259
R5065 vdd.n206 vdd.n164 0.358259
R5066 vdd.n73 vdd.n71 0.358259
R5067 vdd.n75 vdd.n73 0.358259
R5068 vdd.n117 vdd.n75 0.358259
R5069 vdd.n1158 vdd.n1116 0.358259
R5070 vdd.n1116 vdd.n1114 0.358259
R5071 vdd.n1114 vdd.n1112 0.358259
R5072 vdd.n1068 vdd.n1026 0.358259
R5073 vdd.n1026 vdd.n1024 0.358259
R5074 vdd.n1024 vdd.n1022 0.358259
R5075 vdd.n979 vdd.n937 0.358259
R5076 vdd.n937 vdd.n935 0.358259
R5077 vdd.n935 vdd.n933 0.358259
R5078 vdd.n14 vdd.n6 0.334552
R5079 vdd.n14 vdd.n13 0.334552
R5080 vdd.n27 vdd.n19 0.21707
R5081 vdd.n27 vdd.n24 0.21707
R5082 vdd.n294 vdd.n256 0.155672
R5083 vdd.n286 vdd.n256 0.155672
R5084 vdd.n286 vdd.n285 0.155672
R5085 vdd.n285 vdd.n261 0.155672
R5086 vdd.n278 vdd.n261 0.155672
R5087 vdd.n278 vdd.n277 0.155672
R5088 vdd.n277 vdd.n265 0.155672
R5089 vdd.n270 vdd.n265 0.155672
R5090 vdd.n247 vdd.n209 0.155672
R5091 vdd.n239 vdd.n209 0.155672
R5092 vdd.n239 vdd.n238 0.155672
R5093 vdd.n238 vdd.n214 0.155672
R5094 vdd.n231 vdd.n214 0.155672
R5095 vdd.n231 vdd.n230 0.155672
R5096 vdd.n230 vdd.n218 0.155672
R5097 vdd.n223 vdd.n218 0.155672
R5098 vdd.n204 vdd.n166 0.155672
R5099 vdd.n196 vdd.n166 0.155672
R5100 vdd.n196 vdd.n195 0.155672
R5101 vdd.n195 vdd.n171 0.155672
R5102 vdd.n188 vdd.n171 0.155672
R5103 vdd.n188 vdd.n187 0.155672
R5104 vdd.n187 vdd.n175 0.155672
R5105 vdd.n180 vdd.n175 0.155672
R5106 vdd.n157 vdd.n119 0.155672
R5107 vdd.n149 vdd.n119 0.155672
R5108 vdd.n149 vdd.n148 0.155672
R5109 vdd.n148 vdd.n124 0.155672
R5110 vdd.n141 vdd.n124 0.155672
R5111 vdd.n141 vdd.n140 0.155672
R5112 vdd.n140 vdd.n128 0.155672
R5113 vdd.n133 vdd.n128 0.155672
R5114 vdd.n115 vdd.n77 0.155672
R5115 vdd.n107 vdd.n77 0.155672
R5116 vdd.n107 vdd.n106 0.155672
R5117 vdd.n106 vdd.n82 0.155672
R5118 vdd.n99 vdd.n82 0.155672
R5119 vdd.n99 vdd.n98 0.155672
R5120 vdd.n98 vdd.n86 0.155672
R5121 vdd.n91 vdd.n86 0.155672
R5122 vdd.n68 vdd.n30 0.155672
R5123 vdd.n60 vdd.n30 0.155672
R5124 vdd.n60 vdd.n59 0.155672
R5125 vdd.n59 vdd.n35 0.155672
R5126 vdd.n52 vdd.n35 0.155672
R5127 vdd.n52 vdd.n51 0.155672
R5128 vdd.n51 vdd.n39 0.155672
R5129 vdd.n44 vdd.n39 0.155672
R5130 vdd.n1109 vdd.n1071 0.155672
R5131 vdd.n1101 vdd.n1071 0.155672
R5132 vdd.n1101 vdd.n1100 0.155672
R5133 vdd.n1100 vdd.n1076 0.155672
R5134 vdd.n1093 vdd.n1076 0.155672
R5135 vdd.n1093 vdd.n1092 0.155672
R5136 vdd.n1092 vdd.n1080 0.155672
R5137 vdd.n1085 vdd.n1080 0.155672
R5138 vdd.n1156 vdd.n1118 0.155672
R5139 vdd.n1148 vdd.n1118 0.155672
R5140 vdd.n1148 vdd.n1147 0.155672
R5141 vdd.n1147 vdd.n1123 0.155672
R5142 vdd.n1140 vdd.n1123 0.155672
R5143 vdd.n1140 vdd.n1139 0.155672
R5144 vdd.n1139 vdd.n1127 0.155672
R5145 vdd.n1132 vdd.n1127 0.155672
R5146 vdd.n1019 vdd.n981 0.155672
R5147 vdd.n1011 vdd.n981 0.155672
R5148 vdd.n1011 vdd.n1010 0.155672
R5149 vdd.n1010 vdd.n986 0.155672
R5150 vdd.n1003 vdd.n986 0.155672
R5151 vdd.n1003 vdd.n1002 0.155672
R5152 vdd.n1002 vdd.n990 0.155672
R5153 vdd.n995 vdd.n990 0.155672
R5154 vdd.n1066 vdd.n1028 0.155672
R5155 vdd.n1058 vdd.n1028 0.155672
R5156 vdd.n1058 vdd.n1057 0.155672
R5157 vdd.n1057 vdd.n1033 0.155672
R5158 vdd.n1050 vdd.n1033 0.155672
R5159 vdd.n1050 vdd.n1049 0.155672
R5160 vdd.n1049 vdd.n1037 0.155672
R5161 vdd.n1042 vdd.n1037 0.155672
R5162 vdd.n930 vdd.n892 0.155672
R5163 vdd.n922 vdd.n892 0.155672
R5164 vdd.n922 vdd.n921 0.155672
R5165 vdd.n921 vdd.n897 0.155672
R5166 vdd.n914 vdd.n897 0.155672
R5167 vdd.n914 vdd.n913 0.155672
R5168 vdd.n913 vdd.n901 0.155672
R5169 vdd.n906 vdd.n901 0.155672
R5170 vdd.n977 vdd.n939 0.155672
R5171 vdd.n969 vdd.n939 0.155672
R5172 vdd.n969 vdd.n968 0.155672
R5173 vdd.n968 vdd.n944 0.155672
R5174 vdd.n961 vdd.n944 0.155672
R5175 vdd.n961 vdd.n960 0.155672
R5176 vdd.n960 vdd.n948 0.155672
R5177 vdd.n953 vdd.n948 0.155672
R5178 vdd.n1715 vdd.n1520 0.152939
R5179 vdd.n1526 vdd.n1520 0.152939
R5180 vdd.n1527 vdd.n1526 0.152939
R5181 vdd.n1528 vdd.n1527 0.152939
R5182 vdd.n1529 vdd.n1528 0.152939
R5183 vdd.n1533 vdd.n1529 0.152939
R5184 vdd.n1534 vdd.n1533 0.152939
R5185 vdd.n1535 vdd.n1534 0.152939
R5186 vdd.n1536 vdd.n1535 0.152939
R5187 vdd.n1540 vdd.n1536 0.152939
R5188 vdd.n1541 vdd.n1540 0.152939
R5189 vdd.n1542 vdd.n1541 0.152939
R5190 vdd.n1690 vdd.n1542 0.152939
R5191 vdd.n1690 vdd.n1689 0.152939
R5192 vdd.n1689 vdd.n1688 0.152939
R5193 vdd.n1688 vdd.n1548 0.152939
R5194 vdd.n1553 vdd.n1548 0.152939
R5195 vdd.n1554 vdd.n1553 0.152939
R5196 vdd.n1555 vdd.n1554 0.152939
R5197 vdd.n1559 vdd.n1555 0.152939
R5198 vdd.n1560 vdd.n1559 0.152939
R5199 vdd.n1561 vdd.n1560 0.152939
R5200 vdd.n1562 vdd.n1561 0.152939
R5201 vdd.n1566 vdd.n1562 0.152939
R5202 vdd.n1567 vdd.n1566 0.152939
R5203 vdd.n1568 vdd.n1567 0.152939
R5204 vdd.n1569 vdd.n1568 0.152939
R5205 vdd.n1573 vdd.n1569 0.152939
R5206 vdd.n1574 vdd.n1573 0.152939
R5207 vdd.n1575 vdd.n1574 0.152939
R5208 vdd.n1576 vdd.n1575 0.152939
R5209 vdd.n1580 vdd.n1576 0.152939
R5210 vdd.n1581 vdd.n1580 0.152939
R5211 vdd.n1582 vdd.n1581 0.152939
R5212 vdd.n1651 vdd.n1582 0.152939
R5213 vdd.n1651 vdd.n1650 0.152939
R5214 vdd.n1650 vdd.n1649 0.152939
R5215 vdd.n1649 vdd.n1588 0.152939
R5216 vdd.n1593 vdd.n1588 0.152939
R5217 vdd.n1594 vdd.n1593 0.152939
R5218 vdd.n1595 vdd.n1594 0.152939
R5219 vdd.n1599 vdd.n1595 0.152939
R5220 vdd.n1600 vdd.n1599 0.152939
R5221 vdd.n1601 vdd.n1600 0.152939
R5222 vdd.n1602 vdd.n1601 0.152939
R5223 vdd.n1606 vdd.n1602 0.152939
R5224 vdd.n1607 vdd.n1606 0.152939
R5225 vdd.n1608 vdd.n1607 0.152939
R5226 vdd.n1609 vdd.n1608 0.152939
R5227 vdd.n1610 vdd.n1609 0.152939
R5228 vdd.n1610 vdd.n854 0.152939
R5229 vdd.n1939 vdd.n1514 0.152939
R5230 vdd.n1477 vdd.n1476 0.152939
R5231 vdd.n1478 vdd.n1477 0.152939
R5232 vdd.n1478 vdd.n879 0.152939
R5233 vdd.n1493 vdd.n879 0.152939
R5234 vdd.n1494 vdd.n1493 0.152939
R5235 vdd.n1495 vdd.n1494 0.152939
R5236 vdd.n1495 vdd.n867 0.152939
R5237 vdd.n1512 vdd.n867 0.152939
R5238 vdd.n1513 vdd.n1512 0.152939
R5239 vdd.n1940 vdd.n1513 0.152939
R5240 vdd.n524 vdd.n519 0.152939
R5241 vdd.n525 vdd.n524 0.152939
R5242 vdd.n526 vdd.n525 0.152939
R5243 vdd.n527 vdd.n526 0.152939
R5244 vdd.n528 vdd.n527 0.152939
R5245 vdd.n529 vdd.n528 0.152939
R5246 vdd.n530 vdd.n529 0.152939
R5247 vdd.n531 vdd.n530 0.152939
R5248 vdd.n532 vdd.n531 0.152939
R5249 vdd.n533 vdd.n532 0.152939
R5250 vdd.n534 vdd.n533 0.152939
R5251 vdd.n535 vdd.n534 0.152939
R5252 vdd.n2803 vdd.n535 0.152939
R5253 vdd.n2803 vdd.n2802 0.152939
R5254 vdd.n2802 vdd.n2801 0.152939
R5255 vdd.n2801 vdd.n537 0.152939
R5256 vdd.n538 vdd.n537 0.152939
R5257 vdd.n539 vdd.n538 0.152939
R5258 vdd.n540 vdd.n539 0.152939
R5259 vdd.n541 vdd.n540 0.152939
R5260 vdd.n542 vdd.n541 0.152939
R5261 vdd.n543 vdd.n542 0.152939
R5262 vdd.n544 vdd.n543 0.152939
R5263 vdd.n545 vdd.n544 0.152939
R5264 vdd.n546 vdd.n545 0.152939
R5265 vdd.n547 vdd.n546 0.152939
R5266 vdd.n548 vdd.n547 0.152939
R5267 vdd.n549 vdd.n548 0.152939
R5268 vdd.n550 vdd.n549 0.152939
R5269 vdd.n551 vdd.n550 0.152939
R5270 vdd.n552 vdd.n551 0.152939
R5271 vdd.n553 vdd.n552 0.152939
R5272 vdd.n554 vdd.n553 0.152939
R5273 vdd.n555 vdd.n554 0.152939
R5274 vdd.n2757 vdd.n555 0.152939
R5275 vdd.n2757 vdd.n2756 0.152939
R5276 vdd.n2756 vdd.n2755 0.152939
R5277 vdd.n2755 vdd.n559 0.152939
R5278 vdd.n560 vdd.n559 0.152939
R5279 vdd.n561 vdd.n560 0.152939
R5280 vdd.n562 vdd.n561 0.152939
R5281 vdd.n563 vdd.n562 0.152939
R5282 vdd.n564 vdd.n563 0.152939
R5283 vdd.n565 vdd.n564 0.152939
R5284 vdd.n566 vdd.n565 0.152939
R5285 vdd.n567 vdd.n566 0.152939
R5286 vdd.n568 vdd.n567 0.152939
R5287 vdd.n569 vdd.n568 0.152939
R5288 vdd.n570 vdd.n569 0.152939
R5289 vdd.n571 vdd.n570 0.152939
R5290 vdd.n572 vdd.n571 0.152939
R5291 vdd.n2844 vdd.n481 0.152939
R5292 vdd.n2846 vdd.n2845 0.152939
R5293 vdd.n2846 vdd.n470 0.152939
R5294 vdd.n2861 vdd.n470 0.152939
R5295 vdd.n2862 vdd.n2861 0.152939
R5296 vdd.n2863 vdd.n2862 0.152939
R5297 vdd.n2863 vdd.n459 0.152939
R5298 vdd.n2877 vdd.n459 0.152939
R5299 vdd.n2878 vdd.n2877 0.152939
R5300 vdd.n2879 vdd.n2878 0.152939
R5301 vdd.n2879 vdd.n298 0.152939
R5302 vdd.n3046 vdd.n299 0.152939
R5303 vdd.n310 vdd.n299 0.152939
R5304 vdd.n311 vdd.n310 0.152939
R5305 vdd.n312 vdd.n311 0.152939
R5306 vdd.n320 vdd.n312 0.152939
R5307 vdd.n321 vdd.n320 0.152939
R5308 vdd.n322 vdd.n321 0.152939
R5309 vdd.n323 vdd.n322 0.152939
R5310 vdd.n331 vdd.n323 0.152939
R5311 vdd.n3022 vdd.n331 0.152939
R5312 vdd.n3021 vdd.n332 0.152939
R5313 vdd.n335 vdd.n332 0.152939
R5314 vdd.n339 vdd.n335 0.152939
R5315 vdd.n340 vdd.n339 0.152939
R5316 vdd.n341 vdd.n340 0.152939
R5317 vdd.n342 vdd.n341 0.152939
R5318 vdd.n343 vdd.n342 0.152939
R5319 vdd.n347 vdd.n343 0.152939
R5320 vdd.n348 vdd.n347 0.152939
R5321 vdd.n349 vdd.n348 0.152939
R5322 vdd.n350 vdd.n349 0.152939
R5323 vdd.n354 vdd.n350 0.152939
R5324 vdd.n355 vdd.n354 0.152939
R5325 vdd.n356 vdd.n355 0.152939
R5326 vdd.n357 vdd.n356 0.152939
R5327 vdd.n361 vdd.n357 0.152939
R5328 vdd.n362 vdd.n361 0.152939
R5329 vdd.n363 vdd.n362 0.152939
R5330 vdd.n2987 vdd.n363 0.152939
R5331 vdd.n2987 vdd.n2986 0.152939
R5332 vdd.n2986 vdd.n2985 0.152939
R5333 vdd.n2985 vdd.n369 0.152939
R5334 vdd.n374 vdd.n369 0.152939
R5335 vdd.n375 vdd.n374 0.152939
R5336 vdd.n376 vdd.n375 0.152939
R5337 vdd.n380 vdd.n376 0.152939
R5338 vdd.n381 vdd.n380 0.152939
R5339 vdd.n382 vdd.n381 0.152939
R5340 vdd.n383 vdd.n382 0.152939
R5341 vdd.n387 vdd.n383 0.152939
R5342 vdd.n388 vdd.n387 0.152939
R5343 vdd.n389 vdd.n388 0.152939
R5344 vdd.n390 vdd.n389 0.152939
R5345 vdd.n394 vdd.n390 0.152939
R5346 vdd.n395 vdd.n394 0.152939
R5347 vdd.n396 vdd.n395 0.152939
R5348 vdd.n397 vdd.n396 0.152939
R5349 vdd.n401 vdd.n397 0.152939
R5350 vdd.n402 vdd.n401 0.152939
R5351 vdd.n403 vdd.n402 0.152939
R5352 vdd.n2948 vdd.n403 0.152939
R5353 vdd.n2948 vdd.n2947 0.152939
R5354 vdd.n2947 vdd.n2946 0.152939
R5355 vdd.n2946 vdd.n409 0.152939
R5356 vdd.n414 vdd.n409 0.152939
R5357 vdd.n415 vdd.n414 0.152939
R5358 vdd.n416 vdd.n415 0.152939
R5359 vdd.n420 vdd.n416 0.152939
R5360 vdd.n421 vdd.n420 0.152939
R5361 vdd.n422 vdd.n421 0.152939
R5362 vdd.n423 vdd.n422 0.152939
R5363 vdd.n427 vdd.n423 0.152939
R5364 vdd.n428 vdd.n427 0.152939
R5365 vdd.n429 vdd.n428 0.152939
R5366 vdd.n430 vdd.n429 0.152939
R5367 vdd.n434 vdd.n430 0.152939
R5368 vdd.n435 vdd.n434 0.152939
R5369 vdd.n436 vdd.n435 0.152939
R5370 vdd.n437 vdd.n436 0.152939
R5371 vdd.n441 vdd.n437 0.152939
R5372 vdd.n442 vdd.n441 0.152939
R5373 vdd.n443 vdd.n442 0.152939
R5374 vdd.n2904 vdd.n443 0.152939
R5375 vdd.n2852 vdd.n476 0.152939
R5376 vdd.n2853 vdd.n2852 0.152939
R5377 vdd.n2854 vdd.n2853 0.152939
R5378 vdd.n2854 vdd.n464 0.152939
R5379 vdd.n2869 vdd.n464 0.152939
R5380 vdd.n2870 vdd.n2869 0.152939
R5381 vdd.n2871 vdd.n2870 0.152939
R5382 vdd.n2871 vdd.n452 0.152939
R5383 vdd.n2885 vdd.n452 0.152939
R5384 vdd.n2886 vdd.n2885 0.152939
R5385 vdd.n2887 vdd.n2886 0.152939
R5386 vdd.n2887 vdd.n450 0.152939
R5387 vdd.n2891 vdd.n450 0.152939
R5388 vdd.n2892 vdd.n2891 0.152939
R5389 vdd.n2893 vdd.n2892 0.152939
R5390 vdd.n2893 vdd.n447 0.152939
R5391 vdd.n2897 vdd.n447 0.152939
R5392 vdd.n2898 vdd.n2897 0.152939
R5393 vdd.n2899 vdd.n2898 0.152939
R5394 vdd.n2899 vdd.n444 0.152939
R5395 vdd.n2903 vdd.n444 0.152939
R5396 vdd.n2709 vdd.n2708 0.152939
R5397 vdd.n1951 vdd.n857 0.152939
R5398 vdd.n1433 vdd.n1189 0.152939
R5399 vdd.n1434 vdd.n1433 0.152939
R5400 vdd.n1435 vdd.n1434 0.152939
R5401 vdd.n1435 vdd.n1177 0.152939
R5402 vdd.n1450 vdd.n1177 0.152939
R5403 vdd.n1451 vdd.n1450 0.152939
R5404 vdd.n1452 vdd.n1451 0.152939
R5405 vdd.n1452 vdd.n1167 0.152939
R5406 vdd.n1468 vdd.n1167 0.152939
R5407 vdd.n1469 vdd.n1468 0.152939
R5408 vdd.n1470 vdd.n1469 0.152939
R5409 vdd.n1470 vdd.n884 0.152939
R5410 vdd.n1484 vdd.n884 0.152939
R5411 vdd.n1485 vdd.n1484 0.152939
R5412 vdd.n1486 vdd.n1485 0.152939
R5413 vdd.n1486 vdd.n874 0.152939
R5414 vdd.n1501 vdd.n874 0.152939
R5415 vdd.n1502 vdd.n1501 0.152939
R5416 vdd.n1505 vdd.n1502 0.152939
R5417 vdd.n1505 vdd.n1504 0.152939
R5418 vdd.n1504 vdd.n1503 0.152939
R5419 vdd.n1425 vdd.n1194 0.152939
R5420 vdd.n1418 vdd.n1194 0.152939
R5421 vdd.n1418 vdd.n1417 0.152939
R5422 vdd.n1417 vdd.n1416 0.152939
R5423 vdd.n1416 vdd.n1231 0.152939
R5424 vdd.n1412 vdd.n1231 0.152939
R5425 vdd.n1412 vdd.n1411 0.152939
R5426 vdd.n1411 vdd.n1410 0.152939
R5427 vdd.n1410 vdd.n1237 0.152939
R5428 vdd.n1406 vdd.n1237 0.152939
R5429 vdd.n1406 vdd.n1405 0.152939
R5430 vdd.n1405 vdd.n1404 0.152939
R5431 vdd.n1404 vdd.n1243 0.152939
R5432 vdd.n1400 vdd.n1243 0.152939
R5433 vdd.n1400 vdd.n1399 0.152939
R5434 vdd.n1399 vdd.n1398 0.152939
R5435 vdd.n1398 vdd.n1249 0.152939
R5436 vdd.n1394 vdd.n1249 0.152939
R5437 vdd.n1394 vdd.n1393 0.152939
R5438 vdd.n1393 vdd.n1392 0.152939
R5439 vdd.n1392 vdd.n1257 0.152939
R5440 vdd.n1388 vdd.n1257 0.152939
R5441 vdd.n1388 vdd.n1387 0.152939
R5442 vdd.n1387 vdd.n1386 0.152939
R5443 vdd.n1386 vdd.n1263 0.152939
R5444 vdd.n1382 vdd.n1263 0.152939
R5445 vdd.n1382 vdd.n1381 0.152939
R5446 vdd.n1381 vdd.n1380 0.152939
R5447 vdd.n1380 vdd.n1269 0.152939
R5448 vdd.n1376 vdd.n1269 0.152939
R5449 vdd.n1376 vdd.n1375 0.152939
R5450 vdd.n1375 vdd.n1374 0.152939
R5451 vdd.n1374 vdd.n1275 0.152939
R5452 vdd.n1370 vdd.n1275 0.152939
R5453 vdd.n1370 vdd.n1369 0.152939
R5454 vdd.n1369 vdd.n1368 0.152939
R5455 vdd.n1368 vdd.n1281 0.152939
R5456 vdd.n1364 vdd.n1281 0.152939
R5457 vdd.n1364 vdd.n1363 0.152939
R5458 vdd.n1363 vdd.n1362 0.152939
R5459 vdd.n1362 vdd.n1287 0.152939
R5460 vdd.n1355 vdd.n1287 0.152939
R5461 vdd.n1355 vdd.n1354 0.152939
R5462 vdd.n1354 vdd.n1353 0.152939
R5463 vdd.n1353 vdd.n1292 0.152939
R5464 vdd.n1349 vdd.n1292 0.152939
R5465 vdd.n1349 vdd.n1348 0.152939
R5466 vdd.n1348 vdd.n1347 0.152939
R5467 vdd.n1347 vdd.n1298 0.152939
R5468 vdd.n1343 vdd.n1298 0.152939
R5469 vdd.n1343 vdd.n1342 0.152939
R5470 vdd.n1342 vdd.n1341 0.152939
R5471 vdd.n1341 vdd.n1304 0.152939
R5472 vdd.n1337 vdd.n1304 0.152939
R5473 vdd.n1337 vdd.n1336 0.152939
R5474 vdd.n1336 vdd.n1335 0.152939
R5475 vdd.n1335 vdd.n1310 0.152939
R5476 vdd.n1331 vdd.n1310 0.152939
R5477 vdd.n1331 vdd.n1330 0.152939
R5478 vdd.n1330 vdd.n1329 0.152939
R5479 vdd.n1329 vdd.n1316 0.152939
R5480 vdd.n1325 vdd.n1316 0.152939
R5481 vdd.n1325 vdd.n1324 0.152939
R5482 vdd.n1427 vdd.n1426 0.152939
R5483 vdd.n1427 vdd.n1183 0.152939
R5484 vdd.n1442 vdd.n1183 0.152939
R5485 vdd.n1443 vdd.n1442 0.152939
R5486 vdd.n1444 vdd.n1443 0.152939
R5487 vdd.n1444 vdd.n1172 0.152939
R5488 vdd.n1459 vdd.n1172 0.152939
R5489 vdd.n1460 vdd.n1459 0.152939
R5490 vdd.n1462 vdd.n1460 0.152939
R5491 vdd.n1462 vdd.n1461 0.152939
R5492 vdd.n1929 vdd.n1514 0.110256
R5493 vdd.n2836 vdd.n481 0.110256
R5494 vdd.n2708 vdd.n2707 0.110256
R5495 vdd.n1952 vdd.n1951 0.110256
R5496 vdd.n1476 vdd.n1161 0.0695946
R5497 vdd.n3047 vdd.n298 0.0695946
R5498 vdd.n3047 vdd.n3046 0.0695946
R5499 vdd.n1461 vdd.n1161 0.0695946
R5500 vdd.n1929 vdd.n1715 0.0431829
R5501 vdd.n1952 vdd.n854 0.0431829
R5502 vdd.n2836 vdd.n519 0.0431829
R5503 vdd.n2707 vdd.n572 0.0431829
R5504 vdd vdd.n28 0.00833333
R5505 a_n5644_8799.n89 a_n5644_8799.t59 485.149
R5506 a_n5644_8799.n96 a_n5644_8799.t63 485.149
R5507 a_n5644_8799.n104 a_n5644_8799.t29 485.149
R5508 a_n5644_8799.n65 a_n5644_8799.t44 485.149
R5509 a_n5644_8799.n72 a_n5644_8799.t49 485.149
R5510 a_n5644_8799.n80 a_n5644_8799.t30 485.149
R5511 a_n5644_8799.n23 a_n5644_8799.t51 485.135
R5512 a_n5644_8799.n93 a_n5644_8799.t50 464.166
R5513 a_n5644_8799.n87 a_n5644_8799.t36 464.166
R5514 a_n5644_8799.n92 a_n5644_8799.t67 464.166
R5515 a_n5644_8799.n91 a_n5644_8799.t52 464.166
R5516 a_n5644_8799.n88 a_n5644_8799.t41 464.166
R5517 a_n5644_8799.n90 a_n5644_8799.t69 464.166
R5518 a_n5644_8799.n28 a_n5644_8799.t55 485.135
R5519 a_n5644_8799.n100 a_n5644_8799.t54 464.166
R5520 a_n5644_8799.n94 a_n5644_8799.t46 464.166
R5521 a_n5644_8799.n99 a_n5644_8799.t71 464.166
R5522 a_n5644_8799.n98 a_n5644_8799.t57 464.166
R5523 a_n5644_8799.n95 a_n5644_8799.t47 464.166
R5524 a_n5644_8799.n97 a_n5644_8799.t75 464.166
R5525 a_n5644_8799.n33 a_n5644_8799.t74 485.135
R5526 a_n5644_8799.n108 a_n5644_8799.t34 464.166
R5527 a_n5644_8799.n102 a_n5644_8799.t58 464.166
R5528 a_n5644_8799.n107 a_n5644_8799.t28 464.166
R5529 a_n5644_8799.n106 a_n5644_8799.t65 464.166
R5530 a_n5644_8799.n103 a_n5644_8799.t39 464.166
R5531 a_n5644_8799.n105 a_n5644_8799.t62 464.166
R5532 a_n5644_8799.n66 a_n5644_8799.t53 464.166
R5533 a_n5644_8799.n67 a_n5644_8799.t68 464.166
R5534 a_n5644_8799.n68 a_n5644_8799.t33 464.166
R5535 a_n5644_8799.n69 a_n5644_8799.t43 464.166
R5536 a_n5644_8799.n64 a_n5644_8799.t66 464.166
R5537 a_n5644_8799.n70 a_n5644_8799.t31 464.166
R5538 a_n5644_8799.n73 a_n5644_8799.t60 464.166
R5539 a_n5644_8799.n74 a_n5644_8799.t72 464.166
R5540 a_n5644_8799.n75 a_n5644_8799.t42 464.166
R5541 a_n5644_8799.n76 a_n5644_8799.t48 464.166
R5542 a_n5644_8799.n71 a_n5644_8799.t70 464.166
R5543 a_n5644_8799.n77 a_n5644_8799.t38 464.166
R5544 a_n5644_8799.n81 a_n5644_8799.t61 464.166
R5545 a_n5644_8799.n82 a_n5644_8799.t40 464.166
R5546 a_n5644_8799.n83 a_n5644_8799.t64 464.166
R5547 a_n5644_8799.n84 a_n5644_8799.t45 464.166
R5548 a_n5644_8799.n79 a_n5644_8799.t56 464.166
R5549 a_n5644_8799.n85 a_n5644_8799.t35 464.166
R5550 a_n5644_8799.n19 a_n5644_8799.n27 72.3034
R5551 a_n5644_8799.n27 a_n5644_8799.n88 16.6962
R5552 a_n5644_8799.n26 a_n5644_8799.n19 77.6622
R5553 a_n5644_8799.n91 a_n5644_8799.n26 5.97853
R5554 a_n5644_8799.n25 a_n5644_8799.n18 77.6622
R5555 a_n5644_8799.n18 a_n5644_8799.n24 72.3034
R5556 a_n5644_8799.n93 a_n5644_8799.n23 20.9683
R5557 a_n5644_8799.n20 a_n5644_8799.n23 70.1674
R5558 a_n5644_8799.n16 a_n5644_8799.n32 72.3034
R5559 a_n5644_8799.n32 a_n5644_8799.n95 16.6962
R5560 a_n5644_8799.n31 a_n5644_8799.n16 77.6622
R5561 a_n5644_8799.n98 a_n5644_8799.n31 5.97853
R5562 a_n5644_8799.n30 a_n5644_8799.n15 77.6622
R5563 a_n5644_8799.n15 a_n5644_8799.n29 72.3034
R5564 a_n5644_8799.n100 a_n5644_8799.n28 20.9683
R5565 a_n5644_8799.n17 a_n5644_8799.n28 70.1674
R5566 a_n5644_8799.n13 a_n5644_8799.n37 72.3034
R5567 a_n5644_8799.n37 a_n5644_8799.n103 16.6962
R5568 a_n5644_8799.n36 a_n5644_8799.n13 77.6622
R5569 a_n5644_8799.n106 a_n5644_8799.n36 5.97853
R5570 a_n5644_8799.n35 a_n5644_8799.n12 77.6622
R5571 a_n5644_8799.n12 a_n5644_8799.n34 72.3034
R5572 a_n5644_8799.n108 a_n5644_8799.n33 20.9683
R5573 a_n5644_8799.n14 a_n5644_8799.n33 70.1674
R5574 a_n5644_8799.n10 a_n5644_8799.n42 70.1674
R5575 a_n5644_8799.n70 a_n5644_8799.n42 20.9683
R5576 a_n5644_8799.n41 a_n5644_8799.n10 72.3034
R5577 a_n5644_8799.n41 a_n5644_8799.n64 16.6962
R5578 a_n5644_8799.n9 a_n5644_8799.n40 77.6622
R5579 a_n5644_8799.n69 a_n5644_8799.n40 5.97853
R5580 a_n5644_8799.n39 a_n5644_8799.n9 77.6622
R5581 a_n5644_8799.n38 a_n5644_8799.n67 16.6962
R5582 a_n5644_8799.n38 a_n5644_8799.n11 72.3034
R5583 a_n5644_8799.n7 a_n5644_8799.n47 70.1674
R5584 a_n5644_8799.n77 a_n5644_8799.n47 20.9683
R5585 a_n5644_8799.n46 a_n5644_8799.n7 72.3034
R5586 a_n5644_8799.n46 a_n5644_8799.n71 16.6962
R5587 a_n5644_8799.n6 a_n5644_8799.n45 77.6622
R5588 a_n5644_8799.n76 a_n5644_8799.n45 5.97853
R5589 a_n5644_8799.n44 a_n5644_8799.n6 77.6622
R5590 a_n5644_8799.n43 a_n5644_8799.n74 16.6962
R5591 a_n5644_8799.n43 a_n5644_8799.n8 72.3034
R5592 a_n5644_8799.n4 a_n5644_8799.n52 70.1674
R5593 a_n5644_8799.n85 a_n5644_8799.n52 20.9683
R5594 a_n5644_8799.n51 a_n5644_8799.n4 72.3034
R5595 a_n5644_8799.n51 a_n5644_8799.n79 16.6962
R5596 a_n5644_8799.n3 a_n5644_8799.n50 77.6622
R5597 a_n5644_8799.n84 a_n5644_8799.n50 5.97853
R5598 a_n5644_8799.n49 a_n5644_8799.n3 77.6622
R5599 a_n5644_8799.n48 a_n5644_8799.n82 16.6962
R5600 a_n5644_8799.n48 a_n5644_8799.n5 72.3034
R5601 a_n5644_8799.n21 a_n5644_8799.n53 98.9633
R5602 a_n5644_8799.n22 a_n5644_8799.n113 98.9631
R5603 a_n5644_8799.n22 a_n5644_8799.n114 98.6055
R5604 a_n5644_8799.n21 a_n5644_8799.n55 98.6055
R5605 a_n5644_8799.n21 a_n5644_8799.n54 98.6055
R5606 a_n5644_8799.n115 a_n5644_8799.n22 98.6054
R5607 a_n5644_8799.n1 a_n5644_8799.n56 81.4626
R5608 a_n5644_8799.n2 a_n5644_8799.n60 81.4626
R5609 a_n5644_8799.n2 a_n5644_8799.n58 81.4626
R5610 a_n5644_8799.n0 a_n5644_8799.n62 80.9324
R5611 a_n5644_8799.n1 a_n5644_8799.n63 80.9324
R5612 a_n5644_8799.n1 a_n5644_8799.n57 80.9324
R5613 a_n5644_8799.n2 a_n5644_8799.n61 80.9324
R5614 a_n5644_8799.n2 a_n5644_8799.n59 80.9324
R5615 a_n5644_8799.n19 a_n5644_8799.n89 70.4033
R5616 a_n5644_8799.n16 a_n5644_8799.n96 70.4033
R5617 a_n5644_8799.n13 a_n5644_8799.n104 70.4033
R5618 a_n5644_8799.n65 a_n5644_8799.n11 70.4033
R5619 a_n5644_8799.n72 a_n5644_8799.n8 70.4033
R5620 a_n5644_8799.n80 a_n5644_8799.n5 70.4033
R5621 a_n5644_8799.n92 a_n5644_8799.n91 48.2005
R5622 a_n5644_8799.n99 a_n5644_8799.n98 48.2005
R5623 a_n5644_8799.n107 a_n5644_8799.n106 48.2005
R5624 a_n5644_8799.n69 a_n5644_8799.n68 48.2005
R5625 a_n5644_8799.t32 a_n5644_8799.n42 485.135
R5626 a_n5644_8799.n76 a_n5644_8799.n75 48.2005
R5627 a_n5644_8799.t37 a_n5644_8799.n47 485.135
R5628 a_n5644_8799.n84 a_n5644_8799.n83 48.2005
R5629 a_n5644_8799.t73 a_n5644_8799.n52 485.135
R5630 a_n5644_8799.n24 a_n5644_8799.n87 16.6962
R5631 a_n5644_8799.n90 a_n5644_8799.n27 27.6507
R5632 a_n5644_8799.n29 a_n5644_8799.n94 16.6962
R5633 a_n5644_8799.n97 a_n5644_8799.n32 27.6507
R5634 a_n5644_8799.n34 a_n5644_8799.n102 16.6962
R5635 a_n5644_8799.n105 a_n5644_8799.n37 27.6507
R5636 a_n5644_8799.n70 a_n5644_8799.n41 27.6507
R5637 a_n5644_8799.n77 a_n5644_8799.n46 27.6507
R5638 a_n5644_8799.n85 a_n5644_8799.n51 27.6507
R5639 a_n5644_8799.n25 a_n5644_8799.n87 41.7634
R5640 a_n5644_8799.n30 a_n5644_8799.n94 41.7634
R5641 a_n5644_8799.n35 a_n5644_8799.n102 41.7634
R5642 a_n5644_8799.n67 a_n5644_8799.n39 41.7634
R5643 a_n5644_8799.n74 a_n5644_8799.n44 41.7634
R5644 a_n5644_8799.n82 a_n5644_8799.n49 41.7634
R5645 a_n5644_8799.n90 a_n5644_8799.n89 20.9576
R5646 a_n5644_8799.n97 a_n5644_8799.n96 20.9576
R5647 a_n5644_8799.n105 a_n5644_8799.n104 20.9576
R5648 a_n5644_8799.n66 a_n5644_8799.n65 20.9576
R5649 a_n5644_8799.n73 a_n5644_8799.n72 20.9576
R5650 a_n5644_8799.n81 a_n5644_8799.n80 20.9576
R5651 a_n5644_8799.n25 a_n5644_8799.n92 5.97853
R5652 a_n5644_8799.n26 a_n5644_8799.n88 41.7634
R5653 a_n5644_8799.n30 a_n5644_8799.n99 5.97853
R5654 a_n5644_8799.n31 a_n5644_8799.n95 41.7634
R5655 a_n5644_8799.n35 a_n5644_8799.n107 5.97853
R5656 a_n5644_8799.n36 a_n5644_8799.n103 41.7634
R5657 a_n5644_8799.n68 a_n5644_8799.n39 5.97853
R5658 a_n5644_8799.n64 a_n5644_8799.n40 41.7634
R5659 a_n5644_8799.n75 a_n5644_8799.n44 5.97853
R5660 a_n5644_8799.n71 a_n5644_8799.n45 41.7634
R5661 a_n5644_8799.n83 a_n5644_8799.n49 5.97853
R5662 a_n5644_8799.n79 a_n5644_8799.n50 41.7634
R5663 a_n5644_8799.n0 a_n5644_8799.n2 33.2634
R5664 a_n5644_8799.n22 a_n5644_8799.n112 31.0217
R5665 a_n5644_8799.n111 a_n5644_8799.n1 12.3339
R5666 a_n5644_8799.n112 a_n5644_8799.n111 11.4887
R5667 a_n5644_8799.n93 a_n5644_8799.n24 27.6507
R5668 a_n5644_8799.n100 a_n5644_8799.n29 27.6507
R5669 a_n5644_8799.n108 a_n5644_8799.n34 27.6507
R5670 a_n5644_8799.n38 a_n5644_8799.n66 27.6507
R5671 a_n5644_8799.n43 a_n5644_8799.n73 27.6507
R5672 a_n5644_8799.n48 a_n5644_8799.n81 27.6507
R5673 a_n5644_8799.n112 a_n5644_8799.n21 18.1434
R5674 a_n5644_8799.n101 a_n5644_8799.n20 9.05164
R5675 a_n5644_8799.n78 a_n5644_8799.n10 9.05164
R5676 a_n5644_8799.n110 a_n5644_8799.n86 6.86264
R5677 a_n5644_8799.n110 a_n5644_8799.n109 6.52017
R5678 a_n5644_8799.n101 a_n5644_8799.n17 4.94368
R5679 a_n5644_8799.n109 a_n5644_8799.n14 4.94368
R5680 a_n5644_8799.n78 a_n5644_8799.n7 4.94368
R5681 a_n5644_8799.n86 a_n5644_8799.n4 4.94368
R5682 a_n5644_8799.n109 a_n5644_8799.n101 4.10845
R5683 a_n5644_8799.n86 a_n5644_8799.n78 4.10845
R5684 a_n5644_8799.n113 a_n5644_8799.t20 3.61217
R5685 a_n5644_8799.n113 a_n5644_8799.t21 3.61217
R5686 a_n5644_8799.n114 a_n5644_8799.t24 3.61217
R5687 a_n5644_8799.n114 a_n5644_8799.t15 3.61217
R5688 a_n5644_8799.n55 a_n5644_8799.t18 3.61217
R5689 a_n5644_8799.n55 a_n5644_8799.t17 3.61217
R5690 a_n5644_8799.n54 a_n5644_8799.t19 3.61217
R5691 a_n5644_8799.n54 a_n5644_8799.t23 3.61217
R5692 a_n5644_8799.n53 a_n5644_8799.t16 3.61217
R5693 a_n5644_8799.n53 a_n5644_8799.t25 3.61217
R5694 a_n5644_8799.t14 a_n5644_8799.n115 3.61217
R5695 a_n5644_8799.n115 a_n5644_8799.t22 3.61217
R5696 a_n5644_8799.n111 a_n5644_8799.n110 3.4105
R5697 a_n5644_8799.n62 a_n5644_8799.t6 2.82907
R5698 a_n5644_8799.n62 a_n5644_8799.t4 2.82907
R5699 a_n5644_8799.n63 a_n5644_8799.t1 2.82907
R5700 a_n5644_8799.n63 a_n5644_8799.t0 2.82907
R5701 a_n5644_8799.n57 a_n5644_8799.t11 2.82907
R5702 a_n5644_8799.n57 a_n5644_8799.t5 2.82907
R5703 a_n5644_8799.n56 a_n5644_8799.t27 2.82907
R5704 a_n5644_8799.n56 a_n5644_8799.t3 2.82907
R5705 a_n5644_8799.n60 a_n5644_8799.t9 2.82907
R5706 a_n5644_8799.n60 a_n5644_8799.t8 2.82907
R5707 a_n5644_8799.n61 a_n5644_8799.t10 2.82907
R5708 a_n5644_8799.n61 a_n5644_8799.t13 2.82907
R5709 a_n5644_8799.n59 a_n5644_8799.t26 2.82907
R5710 a_n5644_8799.n59 a_n5644_8799.t7 2.82907
R5711 a_n5644_8799.n58 a_n5644_8799.t12 2.82907
R5712 a_n5644_8799.n58 a_n5644_8799.t2 2.82907
R5713 a_n5644_8799.n19 a_n5644_8799.n18 1.13686
R5714 a_n5644_8799.n16 a_n5644_8799.n15 1.13686
R5715 a_n5644_8799.n13 a_n5644_8799.n12 1.13686
R5716 a_n5644_8799.n10 a_n5644_8799.n9 1.13686
R5717 a_n5644_8799.n7 a_n5644_8799.n6 1.13686
R5718 a_n5644_8799.n4 a_n5644_8799.n3 1.13686
R5719 a_n5644_8799.n1 a_n5644_8799.n0 1.06084
R5720 a_n5644_8799.n3 a_n5644_8799.n5 0.568682
R5721 a_n5644_8799.n6 a_n5644_8799.n8 0.568682
R5722 a_n5644_8799.n9 a_n5644_8799.n11 0.568682
R5723 a_n5644_8799.n12 a_n5644_8799.n14 0.568682
R5724 a_n5644_8799.n15 a_n5644_8799.n17 0.568682
R5725 a_n5644_8799.n18 a_n5644_8799.n20 0.568682
R5726 CSoutput.n19 CSoutput.t161 184.661
R5727 CSoutput.n78 CSoutput.n77 165.8
R5728 CSoutput.n76 CSoutput.n0 165.8
R5729 CSoutput.n75 CSoutput.n74 165.8
R5730 CSoutput.n73 CSoutput.n72 165.8
R5731 CSoutput.n71 CSoutput.n2 165.8
R5732 CSoutput.n69 CSoutput.n68 165.8
R5733 CSoutput.n67 CSoutput.n3 165.8
R5734 CSoutput.n66 CSoutput.n65 165.8
R5735 CSoutput.n63 CSoutput.n4 165.8
R5736 CSoutput.n61 CSoutput.n60 165.8
R5737 CSoutput.n59 CSoutput.n5 165.8
R5738 CSoutput.n58 CSoutput.n57 165.8
R5739 CSoutput.n55 CSoutput.n6 165.8
R5740 CSoutput.n54 CSoutput.n53 165.8
R5741 CSoutput.n52 CSoutput.n51 165.8
R5742 CSoutput.n50 CSoutput.n8 165.8
R5743 CSoutput.n48 CSoutput.n47 165.8
R5744 CSoutput.n46 CSoutput.n9 165.8
R5745 CSoutput.n45 CSoutput.n44 165.8
R5746 CSoutput.n42 CSoutput.n10 165.8
R5747 CSoutput.n41 CSoutput.n40 165.8
R5748 CSoutput.n39 CSoutput.n38 165.8
R5749 CSoutput.n37 CSoutput.n12 165.8
R5750 CSoutput.n35 CSoutput.n34 165.8
R5751 CSoutput.n33 CSoutput.n13 165.8
R5752 CSoutput.n32 CSoutput.n31 165.8
R5753 CSoutput.n29 CSoutput.n14 165.8
R5754 CSoutput.n28 CSoutput.n27 165.8
R5755 CSoutput.n26 CSoutput.n25 165.8
R5756 CSoutput.n24 CSoutput.n16 165.8
R5757 CSoutput.n22 CSoutput.n21 165.8
R5758 CSoutput.n20 CSoutput.n17 165.8
R5759 CSoutput.n77 CSoutput.t162 162.194
R5760 CSoutput.n18 CSoutput.t158 120.501
R5761 CSoutput.n23 CSoutput.t153 120.501
R5762 CSoutput.n15 CSoutput.t147 120.501
R5763 CSoutput.n30 CSoutput.t159 120.501
R5764 CSoutput.n36 CSoutput.t160 120.501
R5765 CSoutput.n11 CSoutput.t149 120.501
R5766 CSoutput.n43 CSoutput.t145 120.501
R5767 CSoutput.n49 CSoutput.t163 120.501
R5768 CSoutput.n7 CSoutput.t152 120.501
R5769 CSoutput.n56 CSoutput.t155 120.501
R5770 CSoutput.n62 CSoutput.t164 120.501
R5771 CSoutput.n64 CSoutput.t156 120.501
R5772 CSoutput.n70 CSoutput.t157 120.501
R5773 CSoutput.n1 CSoutput.t150 120.501
R5774 CSoutput.n270 CSoutput.n268 103.469
R5775 CSoutput.n262 CSoutput.n260 103.469
R5776 CSoutput.n255 CSoutput.n253 103.469
R5777 CSoutput.n96 CSoutput.n94 103.469
R5778 CSoutput.n88 CSoutput.n86 103.469
R5779 CSoutput.n81 CSoutput.n79 103.469
R5780 CSoutput.n272 CSoutput.n271 103.111
R5781 CSoutput.n270 CSoutput.n269 103.111
R5782 CSoutput.n266 CSoutput.n265 103.111
R5783 CSoutput.n264 CSoutput.n263 103.111
R5784 CSoutput.n262 CSoutput.n261 103.111
R5785 CSoutput.n259 CSoutput.n258 103.111
R5786 CSoutput.n257 CSoutput.n256 103.111
R5787 CSoutput.n255 CSoutput.n254 103.111
R5788 CSoutput.n96 CSoutput.n95 103.111
R5789 CSoutput.n98 CSoutput.n97 103.111
R5790 CSoutput.n100 CSoutput.n99 103.111
R5791 CSoutput.n88 CSoutput.n87 103.111
R5792 CSoutput.n90 CSoutput.n89 103.111
R5793 CSoutput.n92 CSoutput.n91 103.111
R5794 CSoutput.n81 CSoutput.n80 103.111
R5795 CSoutput.n83 CSoutput.n82 103.111
R5796 CSoutput.n85 CSoutput.n84 103.111
R5797 CSoutput.n274 CSoutput.n273 103.111
R5798 CSoutput.n310 CSoutput.n308 81.5057
R5799 CSoutput.n294 CSoutput.n292 81.5057
R5800 CSoutput.n279 CSoutput.n277 81.5057
R5801 CSoutput.n358 CSoutput.n356 81.5057
R5802 CSoutput.n342 CSoutput.n340 81.5057
R5803 CSoutput.n327 CSoutput.n325 81.5057
R5804 CSoutput.n322 CSoutput.n321 80.9324
R5805 CSoutput.n320 CSoutput.n319 80.9324
R5806 CSoutput.n318 CSoutput.n317 80.9324
R5807 CSoutput.n316 CSoutput.n315 80.9324
R5808 CSoutput.n314 CSoutput.n313 80.9324
R5809 CSoutput.n312 CSoutput.n311 80.9324
R5810 CSoutput.n310 CSoutput.n309 80.9324
R5811 CSoutput.n306 CSoutput.n305 80.9324
R5812 CSoutput.n304 CSoutput.n303 80.9324
R5813 CSoutput.n302 CSoutput.n301 80.9324
R5814 CSoutput.n300 CSoutput.n299 80.9324
R5815 CSoutput.n298 CSoutput.n297 80.9324
R5816 CSoutput.n296 CSoutput.n295 80.9324
R5817 CSoutput.n294 CSoutput.n293 80.9324
R5818 CSoutput.n291 CSoutput.n290 80.9324
R5819 CSoutput.n289 CSoutput.n288 80.9324
R5820 CSoutput.n287 CSoutput.n286 80.9324
R5821 CSoutput.n285 CSoutput.n284 80.9324
R5822 CSoutput.n283 CSoutput.n282 80.9324
R5823 CSoutput.n281 CSoutput.n280 80.9324
R5824 CSoutput.n279 CSoutput.n278 80.9324
R5825 CSoutput.n358 CSoutput.n357 80.9324
R5826 CSoutput.n360 CSoutput.n359 80.9324
R5827 CSoutput.n362 CSoutput.n361 80.9324
R5828 CSoutput.n364 CSoutput.n363 80.9324
R5829 CSoutput.n366 CSoutput.n365 80.9324
R5830 CSoutput.n368 CSoutput.n367 80.9324
R5831 CSoutput.n370 CSoutput.n369 80.9324
R5832 CSoutput.n342 CSoutput.n341 80.9324
R5833 CSoutput.n344 CSoutput.n343 80.9324
R5834 CSoutput.n346 CSoutput.n345 80.9324
R5835 CSoutput.n348 CSoutput.n347 80.9324
R5836 CSoutput.n350 CSoutput.n349 80.9324
R5837 CSoutput.n352 CSoutput.n351 80.9324
R5838 CSoutput.n354 CSoutput.n353 80.9324
R5839 CSoutput.n327 CSoutput.n326 80.9324
R5840 CSoutput.n329 CSoutput.n328 80.9324
R5841 CSoutput.n331 CSoutput.n330 80.9324
R5842 CSoutput.n333 CSoutput.n332 80.9324
R5843 CSoutput.n335 CSoutput.n334 80.9324
R5844 CSoutput.n337 CSoutput.n336 80.9324
R5845 CSoutput.n339 CSoutput.n338 80.9324
R5846 CSoutput.n25 CSoutput.n24 48.1486
R5847 CSoutput.n69 CSoutput.n3 48.1486
R5848 CSoutput.n38 CSoutput.n37 48.1486
R5849 CSoutput.n42 CSoutput.n41 48.1486
R5850 CSoutput.n51 CSoutput.n50 48.1486
R5851 CSoutput.n55 CSoutput.n54 48.1486
R5852 CSoutput.n22 CSoutput.n17 46.462
R5853 CSoutput.n72 CSoutput.n71 46.462
R5854 CSoutput.n20 CSoutput.n19 44.9055
R5855 CSoutput.n29 CSoutput.n28 43.7635
R5856 CSoutput.n65 CSoutput.n63 43.7635
R5857 CSoutput.n35 CSoutput.n13 41.7396
R5858 CSoutput.n57 CSoutput.n5 41.7396
R5859 CSoutput.n44 CSoutput.n9 37.0171
R5860 CSoutput.n48 CSoutput.n9 37.0171
R5861 CSoutput.n76 CSoutput.n75 34.9932
R5862 CSoutput.n31 CSoutput.n13 32.2947
R5863 CSoutput.n61 CSoutput.n5 32.2947
R5864 CSoutput.n30 CSoutput.n29 29.6014
R5865 CSoutput.n63 CSoutput.n62 29.6014
R5866 CSoutput.n19 CSoutput.n18 28.4085
R5867 CSoutput.n18 CSoutput.n17 25.1176
R5868 CSoutput.n72 CSoutput.n1 25.1176
R5869 CSoutput.n43 CSoutput.n42 22.0922
R5870 CSoutput.n50 CSoutput.n49 22.0922
R5871 CSoutput.n77 CSoutput.n76 21.8586
R5872 CSoutput.n37 CSoutput.n36 18.9681
R5873 CSoutput.n56 CSoutput.n55 18.9681
R5874 CSoutput.n25 CSoutput.n15 17.6292
R5875 CSoutput.n64 CSoutput.n3 17.6292
R5876 CSoutput.n24 CSoutput.n23 15.844
R5877 CSoutput.n70 CSoutput.n69 15.844
R5878 CSoutput.n38 CSoutput.n11 14.5051
R5879 CSoutput.n54 CSoutput.n7 14.5051
R5880 CSoutput.n373 CSoutput.n78 11.4982
R5881 CSoutput.n41 CSoutput.n11 11.3811
R5882 CSoutput.n51 CSoutput.n7 11.3811
R5883 CSoutput.n23 CSoutput.n22 10.0422
R5884 CSoutput.n71 CSoutput.n70 10.0422
R5885 CSoutput.n267 CSoutput.n259 9.25285
R5886 CSoutput.n93 CSoutput.n85 9.25285
R5887 CSoutput.n324 CSoutput.n276 9.09499
R5888 CSoutput.n307 CSoutput.n291 8.98182
R5889 CSoutput.n355 CSoutput.n339 8.98182
R5890 CSoutput.n28 CSoutput.n15 8.25698
R5891 CSoutput.n65 CSoutput.n64 8.25698
R5892 CSoutput.n276 CSoutput.n275 7.12641
R5893 CSoutput.n102 CSoutput.n101 7.12641
R5894 CSoutput.n36 CSoutput.n35 6.91809
R5895 CSoutput.n57 CSoutput.n56 6.91809
R5896 CSoutput.n324 CSoutput.n323 6.02792
R5897 CSoutput.n372 CSoutput.n371 6.02792
R5898 CSoutput.n373 CSoutput.n102 5.50255
R5899 CSoutput.n323 CSoutput.n322 5.25266
R5900 CSoutput.n307 CSoutput.n306 5.25266
R5901 CSoutput.n371 CSoutput.n370 5.25266
R5902 CSoutput.n355 CSoutput.n354 5.25266
R5903 CSoutput.n275 CSoutput.n274 5.1449
R5904 CSoutput.n267 CSoutput.n266 5.1449
R5905 CSoutput.n101 CSoutput.n100 5.1449
R5906 CSoutput.n93 CSoutput.n92 5.1449
R5907 CSoutput.n193 CSoutput.n146 4.5005
R5908 CSoutput.n162 CSoutput.n146 4.5005
R5909 CSoutput.n157 CSoutput.n141 4.5005
R5910 CSoutput.n157 CSoutput.n143 4.5005
R5911 CSoutput.n157 CSoutput.n140 4.5005
R5912 CSoutput.n157 CSoutput.n144 4.5005
R5913 CSoutput.n157 CSoutput.n139 4.5005
R5914 CSoutput.n157 CSoutput.t165 4.5005
R5915 CSoutput.n157 CSoutput.n138 4.5005
R5916 CSoutput.n157 CSoutput.n145 4.5005
R5917 CSoutput.n157 CSoutput.n146 4.5005
R5918 CSoutput.n155 CSoutput.n141 4.5005
R5919 CSoutput.n155 CSoutput.n143 4.5005
R5920 CSoutput.n155 CSoutput.n140 4.5005
R5921 CSoutput.n155 CSoutput.n144 4.5005
R5922 CSoutput.n155 CSoutput.n139 4.5005
R5923 CSoutput.n155 CSoutput.t165 4.5005
R5924 CSoutput.n155 CSoutput.n138 4.5005
R5925 CSoutput.n155 CSoutput.n145 4.5005
R5926 CSoutput.n155 CSoutput.n146 4.5005
R5927 CSoutput.n154 CSoutput.n141 4.5005
R5928 CSoutput.n154 CSoutput.n143 4.5005
R5929 CSoutput.n154 CSoutput.n140 4.5005
R5930 CSoutput.n154 CSoutput.n144 4.5005
R5931 CSoutput.n154 CSoutput.n139 4.5005
R5932 CSoutput.n154 CSoutput.t165 4.5005
R5933 CSoutput.n154 CSoutput.n138 4.5005
R5934 CSoutput.n154 CSoutput.n145 4.5005
R5935 CSoutput.n154 CSoutput.n146 4.5005
R5936 CSoutput.n239 CSoutput.n141 4.5005
R5937 CSoutput.n239 CSoutput.n143 4.5005
R5938 CSoutput.n239 CSoutput.n140 4.5005
R5939 CSoutput.n239 CSoutput.n144 4.5005
R5940 CSoutput.n239 CSoutput.n139 4.5005
R5941 CSoutput.n239 CSoutput.t165 4.5005
R5942 CSoutput.n239 CSoutput.n138 4.5005
R5943 CSoutput.n239 CSoutput.n145 4.5005
R5944 CSoutput.n239 CSoutput.n146 4.5005
R5945 CSoutput.n237 CSoutput.n141 4.5005
R5946 CSoutput.n237 CSoutput.n143 4.5005
R5947 CSoutput.n237 CSoutput.n140 4.5005
R5948 CSoutput.n237 CSoutput.n144 4.5005
R5949 CSoutput.n237 CSoutput.n139 4.5005
R5950 CSoutput.n237 CSoutput.t165 4.5005
R5951 CSoutput.n237 CSoutput.n138 4.5005
R5952 CSoutput.n237 CSoutput.n145 4.5005
R5953 CSoutput.n235 CSoutput.n141 4.5005
R5954 CSoutput.n235 CSoutput.n143 4.5005
R5955 CSoutput.n235 CSoutput.n140 4.5005
R5956 CSoutput.n235 CSoutput.n144 4.5005
R5957 CSoutput.n235 CSoutput.n139 4.5005
R5958 CSoutput.n235 CSoutput.t165 4.5005
R5959 CSoutput.n235 CSoutput.n138 4.5005
R5960 CSoutput.n235 CSoutput.n145 4.5005
R5961 CSoutput.n165 CSoutput.n141 4.5005
R5962 CSoutput.n165 CSoutput.n143 4.5005
R5963 CSoutput.n165 CSoutput.n140 4.5005
R5964 CSoutput.n165 CSoutput.n144 4.5005
R5965 CSoutput.n165 CSoutput.n139 4.5005
R5966 CSoutput.n165 CSoutput.t165 4.5005
R5967 CSoutput.n165 CSoutput.n138 4.5005
R5968 CSoutput.n165 CSoutput.n145 4.5005
R5969 CSoutput.n165 CSoutput.n146 4.5005
R5970 CSoutput.n164 CSoutput.n141 4.5005
R5971 CSoutput.n164 CSoutput.n143 4.5005
R5972 CSoutput.n164 CSoutput.n140 4.5005
R5973 CSoutput.n164 CSoutput.n144 4.5005
R5974 CSoutput.n164 CSoutput.n139 4.5005
R5975 CSoutput.n164 CSoutput.t165 4.5005
R5976 CSoutput.n164 CSoutput.n138 4.5005
R5977 CSoutput.n164 CSoutput.n145 4.5005
R5978 CSoutput.n164 CSoutput.n146 4.5005
R5979 CSoutput.n168 CSoutput.n141 4.5005
R5980 CSoutput.n168 CSoutput.n143 4.5005
R5981 CSoutput.n168 CSoutput.n140 4.5005
R5982 CSoutput.n168 CSoutput.n144 4.5005
R5983 CSoutput.n168 CSoutput.n139 4.5005
R5984 CSoutput.n168 CSoutput.t165 4.5005
R5985 CSoutput.n168 CSoutput.n138 4.5005
R5986 CSoutput.n168 CSoutput.n145 4.5005
R5987 CSoutput.n168 CSoutput.n146 4.5005
R5988 CSoutput.n167 CSoutput.n141 4.5005
R5989 CSoutput.n167 CSoutput.n143 4.5005
R5990 CSoutput.n167 CSoutput.n140 4.5005
R5991 CSoutput.n167 CSoutput.n144 4.5005
R5992 CSoutput.n167 CSoutput.n139 4.5005
R5993 CSoutput.n167 CSoutput.t165 4.5005
R5994 CSoutput.n167 CSoutput.n138 4.5005
R5995 CSoutput.n167 CSoutput.n145 4.5005
R5996 CSoutput.n167 CSoutput.n146 4.5005
R5997 CSoutput.n150 CSoutput.n141 4.5005
R5998 CSoutput.n150 CSoutput.n143 4.5005
R5999 CSoutput.n150 CSoutput.n140 4.5005
R6000 CSoutput.n150 CSoutput.n144 4.5005
R6001 CSoutput.n150 CSoutput.n139 4.5005
R6002 CSoutput.n150 CSoutput.t165 4.5005
R6003 CSoutput.n150 CSoutput.n138 4.5005
R6004 CSoutput.n150 CSoutput.n145 4.5005
R6005 CSoutput.n150 CSoutput.n146 4.5005
R6006 CSoutput.n242 CSoutput.n141 4.5005
R6007 CSoutput.n242 CSoutput.n143 4.5005
R6008 CSoutput.n242 CSoutput.n140 4.5005
R6009 CSoutput.n242 CSoutput.n144 4.5005
R6010 CSoutput.n242 CSoutput.n139 4.5005
R6011 CSoutput.n242 CSoutput.t165 4.5005
R6012 CSoutput.n242 CSoutput.n138 4.5005
R6013 CSoutput.n242 CSoutput.n145 4.5005
R6014 CSoutput.n242 CSoutput.n146 4.5005
R6015 CSoutput.n229 CSoutput.n200 4.5005
R6016 CSoutput.n229 CSoutput.n206 4.5005
R6017 CSoutput.n187 CSoutput.n176 4.5005
R6018 CSoutput.n187 CSoutput.n178 4.5005
R6019 CSoutput.n187 CSoutput.n175 4.5005
R6020 CSoutput.n187 CSoutput.n179 4.5005
R6021 CSoutput.n187 CSoutput.n174 4.5005
R6022 CSoutput.n187 CSoutput.t144 4.5005
R6023 CSoutput.n187 CSoutput.n173 4.5005
R6024 CSoutput.n187 CSoutput.n180 4.5005
R6025 CSoutput.n229 CSoutput.n187 4.5005
R6026 CSoutput.n208 CSoutput.n176 4.5005
R6027 CSoutput.n208 CSoutput.n178 4.5005
R6028 CSoutput.n208 CSoutput.n175 4.5005
R6029 CSoutput.n208 CSoutput.n179 4.5005
R6030 CSoutput.n208 CSoutput.n174 4.5005
R6031 CSoutput.n208 CSoutput.t144 4.5005
R6032 CSoutput.n208 CSoutput.n173 4.5005
R6033 CSoutput.n208 CSoutput.n180 4.5005
R6034 CSoutput.n229 CSoutput.n208 4.5005
R6035 CSoutput.n186 CSoutput.n176 4.5005
R6036 CSoutput.n186 CSoutput.n178 4.5005
R6037 CSoutput.n186 CSoutput.n175 4.5005
R6038 CSoutput.n186 CSoutput.n179 4.5005
R6039 CSoutput.n186 CSoutput.n174 4.5005
R6040 CSoutput.n186 CSoutput.t144 4.5005
R6041 CSoutput.n186 CSoutput.n173 4.5005
R6042 CSoutput.n186 CSoutput.n180 4.5005
R6043 CSoutput.n229 CSoutput.n186 4.5005
R6044 CSoutput.n210 CSoutput.n176 4.5005
R6045 CSoutput.n210 CSoutput.n178 4.5005
R6046 CSoutput.n210 CSoutput.n175 4.5005
R6047 CSoutput.n210 CSoutput.n179 4.5005
R6048 CSoutput.n210 CSoutput.n174 4.5005
R6049 CSoutput.n210 CSoutput.t144 4.5005
R6050 CSoutput.n210 CSoutput.n173 4.5005
R6051 CSoutput.n210 CSoutput.n180 4.5005
R6052 CSoutput.n229 CSoutput.n210 4.5005
R6053 CSoutput.n176 CSoutput.n171 4.5005
R6054 CSoutput.n178 CSoutput.n171 4.5005
R6055 CSoutput.n175 CSoutput.n171 4.5005
R6056 CSoutput.n179 CSoutput.n171 4.5005
R6057 CSoutput.n174 CSoutput.n171 4.5005
R6058 CSoutput.t144 CSoutput.n171 4.5005
R6059 CSoutput.n173 CSoutput.n171 4.5005
R6060 CSoutput.n180 CSoutput.n171 4.5005
R6061 CSoutput.n232 CSoutput.n176 4.5005
R6062 CSoutput.n232 CSoutput.n178 4.5005
R6063 CSoutput.n232 CSoutput.n175 4.5005
R6064 CSoutput.n232 CSoutput.n179 4.5005
R6065 CSoutput.n232 CSoutput.n174 4.5005
R6066 CSoutput.n232 CSoutput.t144 4.5005
R6067 CSoutput.n232 CSoutput.n173 4.5005
R6068 CSoutput.n232 CSoutput.n180 4.5005
R6069 CSoutput.n230 CSoutput.n176 4.5005
R6070 CSoutput.n230 CSoutput.n178 4.5005
R6071 CSoutput.n230 CSoutput.n175 4.5005
R6072 CSoutput.n230 CSoutput.n179 4.5005
R6073 CSoutput.n230 CSoutput.n174 4.5005
R6074 CSoutput.n230 CSoutput.t144 4.5005
R6075 CSoutput.n230 CSoutput.n173 4.5005
R6076 CSoutput.n230 CSoutput.n180 4.5005
R6077 CSoutput.n230 CSoutput.n229 4.5005
R6078 CSoutput.n212 CSoutput.n176 4.5005
R6079 CSoutput.n212 CSoutput.n178 4.5005
R6080 CSoutput.n212 CSoutput.n175 4.5005
R6081 CSoutput.n212 CSoutput.n179 4.5005
R6082 CSoutput.n212 CSoutput.n174 4.5005
R6083 CSoutput.n212 CSoutput.t144 4.5005
R6084 CSoutput.n212 CSoutput.n173 4.5005
R6085 CSoutput.n212 CSoutput.n180 4.5005
R6086 CSoutput.n229 CSoutput.n212 4.5005
R6087 CSoutput.n184 CSoutput.n176 4.5005
R6088 CSoutput.n184 CSoutput.n178 4.5005
R6089 CSoutput.n184 CSoutput.n175 4.5005
R6090 CSoutput.n184 CSoutput.n179 4.5005
R6091 CSoutput.n184 CSoutput.n174 4.5005
R6092 CSoutput.n184 CSoutput.t144 4.5005
R6093 CSoutput.n184 CSoutput.n173 4.5005
R6094 CSoutput.n184 CSoutput.n180 4.5005
R6095 CSoutput.n229 CSoutput.n184 4.5005
R6096 CSoutput.n214 CSoutput.n176 4.5005
R6097 CSoutput.n214 CSoutput.n178 4.5005
R6098 CSoutput.n214 CSoutput.n175 4.5005
R6099 CSoutput.n214 CSoutput.n179 4.5005
R6100 CSoutput.n214 CSoutput.n174 4.5005
R6101 CSoutput.n214 CSoutput.t144 4.5005
R6102 CSoutput.n214 CSoutput.n173 4.5005
R6103 CSoutput.n214 CSoutput.n180 4.5005
R6104 CSoutput.n229 CSoutput.n214 4.5005
R6105 CSoutput.n183 CSoutput.n176 4.5005
R6106 CSoutput.n183 CSoutput.n178 4.5005
R6107 CSoutput.n183 CSoutput.n175 4.5005
R6108 CSoutput.n183 CSoutput.n179 4.5005
R6109 CSoutput.n183 CSoutput.n174 4.5005
R6110 CSoutput.n183 CSoutput.t144 4.5005
R6111 CSoutput.n183 CSoutput.n173 4.5005
R6112 CSoutput.n183 CSoutput.n180 4.5005
R6113 CSoutput.n229 CSoutput.n183 4.5005
R6114 CSoutput.n228 CSoutput.n176 4.5005
R6115 CSoutput.n228 CSoutput.n178 4.5005
R6116 CSoutput.n228 CSoutput.n175 4.5005
R6117 CSoutput.n228 CSoutput.n179 4.5005
R6118 CSoutput.n228 CSoutput.n174 4.5005
R6119 CSoutput.n228 CSoutput.t144 4.5005
R6120 CSoutput.n228 CSoutput.n173 4.5005
R6121 CSoutput.n228 CSoutput.n180 4.5005
R6122 CSoutput.n229 CSoutput.n228 4.5005
R6123 CSoutput.n227 CSoutput.n112 4.5005
R6124 CSoutput.n128 CSoutput.n112 4.5005
R6125 CSoutput.n123 CSoutput.n107 4.5005
R6126 CSoutput.n123 CSoutput.n109 4.5005
R6127 CSoutput.n123 CSoutput.n106 4.5005
R6128 CSoutput.n123 CSoutput.n110 4.5005
R6129 CSoutput.n123 CSoutput.n105 4.5005
R6130 CSoutput.n123 CSoutput.t151 4.5005
R6131 CSoutput.n123 CSoutput.n104 4.5005
R6132 CSoutput.n123 CSoutput.n111 4.5005
R6133 CSoutput.n123 CSoutput.n112 4.5005
R6134 CSoutput.n121 CSoutput.n107 4.5005
R6135 CSoutput.n121 CSoutput.n109 4.5005
R6136 CSoutput.n121 CSoutput.n106 4.5005
R6137 CSoutput.n121 CSoutput.n110 4.5005
R6138 CSoutput.n121 CSoutput.n105 4.5005
R6139 CSoutput.n121 CSoutput.t151 4.5005
R6140 CSoutput.n121 CSoutput.n104 4.5005
R6141 CSoutput.n121 CSoutput.n111 4.5005
R6142 CSoutput.n121 CSoutput.n112 4.5005
R6143 CSoutput.n120 CSoutput.n107 4.5005
R6144 CSoutput.n120 CSoutput.n109 4.5005
R6145 CSoutput.n120 CSoutput.n106 4.5005
R6146 CSoutput.n120 CSoutput.n110 4.5005
R6147 CSoutput.n120 CSoutput.n105 4.5005
R6148 CSoutput.n120 CSoutput.t151 4.5005
R6149 CSoutput.n120 CSoutput.n104 4.5005
R6150 CSoutput.n120 CSoutput.n111 4.5005
R6151 CSoutput.n120 CSoutput.n112 4.5005
R6152 CSoutput.n249 CSoutput.n107 4.5005
R6153 CSoutput.n249 CSoutput.n109 4.5005
R6154 CSoutput.n249 CSoutput.n106 4.5005
R6155 CSoutput.n249 CSoutput.n110 4.5005
R6156 CSoutput.n249 CSoutput.n105 4.5005
R6157 CSoutput.n249 CSoutput.t151 4.5005
R6158 CSoutput.n249 CSoutput.n104 4.5005
R6159 CSoutput.n249 CSoutput.n111 4.5005
R6160 CSoutput.n249 CSoutput.n112 4.5005
R6161 CSoutput.n247 CSoutput.n107 4.5005
R6162 CSoutput.n247 CSoutput.n109 4.5005
R6163 CSoutput.n247 CSoutput.n106 4.5005
R6164 CSoutput.n247 CSoutput.n110 4.5005
R6165 CSoutput.n247 CSoutput.n105 4.5005
R6166 CSoutput.n247 CSoutput.t151 4.5005
R6167 CSoutput.n247 CSoutput.n104 4.5005
R6168 CSoutput.n247 CSoutput.n111 4.5005
R6169 CSoutput.n245 CSoutput.n107 4.5005
R6170 CSoutput.n245 CSoutput.n109 4.5005
R6171 CSoutput.n245 CSoutput.n106 4.5005
R6172 CSoutput.n245 CSoutput.n110 4.5005
R6173 CSoutput.n245 CSoutput.n105 4.5005
R6174 CSoutput.n245 CSoutput.t151 4.5005
R6175 CSoutput.n245 CSoutput.n104 4.5005
R6176 CSoutput.n245 CSoutput.n111 4.5005
R6177 CSoutput.n131 CSoutput.n107 4.5005
R6178 CSoutput.n131 CSoutput.n109 4.5005
R6179 CSoutput.n131 CSoutput.n106 4.5005
R6180 CSoutput.n131 CSoutput.n110 4.5005
R6181 CSoutput.n131 CSoutput.n105 4.5005
R6182 CSoutput.n131 CSoutput.t151 4.5005
R6183 CSoutput.n131 CSoutput.n104 4.5005
R6184 CSoutput.n131 CSoutput.n111 4.5005
R6185 CSoutput.n131 CSoutput.n112 4.5005
R6186 CSoutput.n130 CSoutput.n107 4.5005
R6187 CSoutput.n130 CSoutput.n109 4.5005
R6188 CSoutput.n130 CSoutput.n106 4.5005
R6189 CSoutput.n130 CSoutput.n110 4.5005
R6190 CSoutput.n130 CSoutput.n105 4.5005
R6191 CSoutput.n130 CSoutput.t151 4.5005
R6192 CSoutput.n130 CSoutput.n104 4.5005
R6193 CSoutput.n130 CSoutput.n111 4.5005
R6194 CSoutput.n130 CSoutput.n112 4.5005
R6195 CSoutput.n134 CSoutput.n107 4.5005
R6196 CSoutput.n134 CSoutput.n109 4.5005
R6197 CSoutput.n134 CSoutput.n106 4.5005
R6198 CSoutput.n134 CSoutput.n110 4.5005
R6199 CSoutput.n134 CSoutput.n105 4.5005
R6200 CSoutput.n134 CSoutput.t151 4.5005
R6201 CSoutput.n134 CSoutput.n104 4.5005
R6202 CSoutput.n134 CSoutput.n111 4.5005
R6203 CSoutput.n134 CSoutput.n112 4.5005
R6204 CSoutput.n133 CSoutput.n107 4.5005
R6205 CSoutput.n133 CSoutput.n109 4.5005
R6206 CSoutput.n133 CSoutput.n106 4.5005
R6207 CSoutput.n133 CSoutput.n110 4.5005
R6208 CSoutput.n133 CSoutput.n105 4.5005
R6209 CSoutput.n133 CSoutput.t151 4.5005
R6210 CSoutput.n133 CSoutput.n104 4.5005
R6211 CSoutput.n133 CSoutput.n111 4.5005
R6212 CSoutput.n133 CSoutput.n112 4.5005
R6213 CSoutput.n116 CSoutput.n107 4.5005
R6214 CSoutput.n116 CSoutput.n109 4.5005
R6215 CSoutput.n116 CSoutput.n106 4.5005
R6216 CSoutput.n116 CSoutput.n110 4.5005
R6217 CSoutput.n116 CSoutput.n105 4.5005
R6218 CSoutput.n116 CSoutput.t151 4.5005
R6219 CSoutput.n116 CSoutput.n104 4.5005
R6220 CSoutput.n116 CSoutput.n111 4.5005
R6221 CSoutput.n116 CSoutput.n112 4.5005
R6222 CSoutput.n252 CSoutput.n107 4.5005
R6223 CSoutput.n252 CSoutput.n109 4.5005
R6224 CSoutput.n252 CSoutput.n106 4.5005
R6225 CSoutput.n252 CSoutput.n110 4.5005
R6226 CSoutput.n252 CSoutput.n105 4.5005
R6227 CSoutput.n252 CSoutput.t151 4.5005
R6228 CSoutput.n252 CSoutput.n104 4.5005
R6229 CSoutput.n252 CSoutput.n111 4.5005
R6230 CSoutput.n252 CSoutput.n112 4.5005
R6231 CSoutput.n275 CSoutput.n267 4.10845
R6232 CSoutput.n101 CSoutput.n93 4.10845
R6233 CSoutput.n273 CSoutput.t38 4.06363
R6234 CSoutput.n273 CSoutput.t48 4.06363
R6235 CSoutput.n271 CSoutput.t55 4.06363
R6236 CSoutput.n271 CSoutput.t66 4.06363
R6237 CSoutput.n269 CSoutput.t71 4.06363
R6238 CSoutput.n269 CSoutput.t40 4.06363
R6239 CSoutput.n268 CSoutput.t56 4.06363
R6240 CSoutput.n268 CSoutput.t57 4.06363
R6241 CSoutput.n265 CSoutput.t32 4.06363
R6242 CSoutput.n265 CSoutput.t44 4.06363
R6243 CSoutput.n263 CSoutput.t50 4.06363
R6244 CSoutput.n263 CSoutput.t60 4.06363
R6245 CSoutput.n261 CSoutput.t61 4.06363
R6246 CSoutput.n261 CSoutput.t36 4.06363
R6247 CSoutput.n260 CSoutput.t52 4.06363
R6248 CSoutput.n260 CSoutput.t53 4.06363
R6249 CSoutput.n258 CSoutput.t45 4.06363
R6250 CSoutput.n258 CSoutput.t78 4.06363
R6251 CSoutput.n256 CSoutput.t42 4.06363
R6252 CSoutput.n256 CSoutput.t68 4.06363
R6253 CSoutput.n254 CSoutput.t49 4.06363
R6254 CSoutput.n254 CSoutput.t79 4.06363
R6255 CSoutput.n253 CSoutput.t33 4.06363
R6256 CSoutput.n253 CSoutput.t73 4.06363
R6257 CSoutput.n94 CSoutput.t76 4.06363
R6258 CSoutput.n94 CSoutput.t75 4.06363
R6259 CSoutput.n95 CSoutput.t64 4.06363
R6260 CSoutput.n95 CSoutput.t41 4.06363
R6261 CSoutput.n97 CSoutput.t39 4.06363
R6262 CSoutput.n97 CSoutput.t74 4.06363
R6263 CSoutput.n99 CSoutput.t63 4.06363
R6264 CSoutput.n99 CSoutput.t54 4.06363
R6265 CSoutput.n86 CSoutput.t69 4.06363
R6266 CSoutput.n86 CSoutput.t70 4.06363
R6267 CSoutput.n87 CSoutput.t59 4.06363
R6268 CSoutput.n87 CSoutput.t37 4.06363
R6269 CSoutput.n89 CSoutput.t35 4.06363
R6270 CSoutput.n89 CSoutput.t65 4.06363
R6271 CSoutput.n91 CSoutput.t58 4.06363
R6272 CSoutput.n91 CSoutput.t47 4.06363
R6273 CSoutput.n79 CSoutput.t72 4.06363
R6274 CSoutput.n79 CSoutput.t34 4.06363
R6275 CSoutput.n80 CSoutput.t62 4.06363
R6276 CSoutput.n80 CSoutput.t51 4.06363
R6277 CSoutput.n82 CSoutput.t67 4.06363
R6278 CSoutput.n82 CSoutput.t43 4.06363
R6279 CSoutput.n84 CSoutput.t77 4.06363
R6280 CSoutput.n84 CSoutput.t46 4.06363
R6281 CSoutput.n44 CSoutput.n43 3.79402
R6282 CSoutput.n49 CSoutput.n48 3.79402
R6283 CSoutput.n323 CSoutput.n307 3.72967
R6284 CSoutput.n371 CSoutput.n355 3.72967
R6285 CSoutput.n373 CSoutput.n372 3.57343
R6286 CSoutput.n372 CSoutput.n324 3.08965
R6287 CSoutput.n321 CSoutput.t103 2.82907
R6288 CSoutput.n321 CSoutput.t20 2.82907
R6289 CSoutput.n319 CSoutput.t4 2.82907
R6290 CSoutput.n319 CSoutput.t122 2.82907
R6291 CSoutput.n317 CSoutput.t2 2.82907
R6292 CSoutput.n317 CSoutput.t16 2.82907
R6293 CSoutput.n315 CSoutput.t12 2.82907
R6294 CSoutput.n315 CSoutput.t98 2.82907
R6295 CSoutput.n313 CSoutput.t129 2.82907
R6296 CSoutput.n313 CSoutput.t120 2.82907
R6297 CSoutput.n311 CSoutput.t14 2.82907
R6298 CSoutput.n311 CSoutput.t135 2.82907
R6299 CSoutput.n309 CSoutput.t89 2.82907
R6300 CSoutput.n309 CSoutput.t102 2.82907
R6301 CSoutput.n308 CSoutput.t116 2.82907
R6302 CSoutput.n308 CSoutput.t81 2.82907
R6303 CSoutput.n305 CSoutput.t138 2.82907
R6304 CSoutput.n305 CSoutput.t108 2.82907
R6305 CSoutput.n303 CSoutput.t143 2.82907
R6306 CSoutput.n303 CSoutput.t126 2.82907
R6307 CSoutput.n301 CSoutput.t17 2.82907
R6308 CSoutput.n301 CSoutput.t104 2.82907
R6309 CSoutput.n299 CSoutput.t106 2.82907
R6310 CSoutput.n299 CSoutput.t8 2.82907
R6311 CSoutput.n297 CSoutput.t123 2.82907
R6312 CSoutput.n297 CSoutput.t11 2.82907
R6313 CSoutput.n295 CSoutput.t24 2.82907
R6314 CSoutput.n295 CSoutput.t1 2.82907
R6315 CSoutput.n293 CSoutput.t13 2.82907
R6316 CSoutput.n293 CSoutput.t27 2.82907
R6317 CSoutput.n292 CSoutput.t132 2.82907
R6318 CSoutput.n292 CSoutput.t15 2.82907
R6319 CSoutput.n290 CSoutput.t18 2.82907
R6320 CSoutput.n290 CSoutput.t90 2.82907
R6321 CSoutput.n288 CSoutput.t94 2.82907
R6322 CSoutput.n288 CSoutput.t128 2.82907
R6323 CSoutput.n286 CSoutput.t96 2.82907
R6324 CSoutput.n286 CSoutput.t22 2.82907
R6325 CSoutput.n284 CSoutput.t97 2.82907
R6326 CSoutput.n284 CSoutput.t28 2.82907
R6327 CSoutput.n282 CSoutput.t140 2.82907
R6328 CSoutput.n282 CSoutput.t88 2.82907
R6329 CSoutput.n280 CSoutput.t119 2.82907
R6330 CSoutput.n280 CSoutput.t141 2.82907
R6331 CSoutput.n278 CSoutput.t30 2.82907
R6332 CSoutput.n278 CSoutput.t130 2.82907
R6333 CSoutput.n277 CSoutput.t142 2.82907
R6334 CSoutput.n277 CSoutput.t99 2.82907
R6335 CSoutput.n356 CSoutput.t127 2.82907
R6336 CSoutput.n356 CSoutput.t91 2.82907
R6337 CSoutput.n357 CSoutput.t111 2.82907
R6338 CSoutput.n357 CSoutput.t9 2.82907
R6339 CSoutput.n359 CSoutput.t31 2.82907
R6340 CSoutput.n359 CSoutput.t82 2.82907
R6341 CSoutput.n361 CSoutput.t125 2.82907
R6342 CSoutput.n361 CSoutput.t114 2.82907
R6343 CSoutput.n363 CSoutput.t93 2.82907
R6344 CSoutput.n363 CSoutput.t133 2.82907
R6345 CSoutput.n365 CSoutput.t19 2.82907
R6346 CSoutput.n365 CSoutput.t23 2.82907
R6347 CSoutput.n367 CSoutput.t109 2.82907
R6348 CSoutput.n367 CSoutput.t5 2.82907
R6349 CSoutput.n369 CSoutput.t101 2.82907
R6350 CSoutput.n369 CSoutput.t113 2.82907
R6351 CSoutput.n340 CSoutput.t95 2.82907
R6352 CSoutput.n340 CSoutput.t83 2.82907
R6353 CSoutput.n341 CSoutput.t3 2.82907
R6354 CSoutput.n341 CSoutput.t117 2.82907
R6355 CSoutput.n343 CSoutput.t118 2.82907
R6356 CSoutput.n343 CSoutput.t21 2.82907
R6357 CSoutput.n345 CSoutput.t112 2.82907
R6358 CSoutput.n345 CSoutput.t136 2.82907
R6359 CSoutput.n347 CSoutput.t86 2.82907
R6360 CSoutput.n347 CSoutput.t25 2.82907
R6361 CSoutput.n349 CSoutput.t100 2.82907
R6362 CSoutput.n349 CSoutput.t124 2.82907
R6363 CSoutput.n351 CSoutput.t6 2.82907
R6364 CSoutput.n351 CSoutput.t139 2.82907
R6365 CSoutput.n353 CSoutput.t85 2.82907
R6366 CSoutput.n353 CSoutput.t26 2.82907
R6367 CSoutput.n325 CSoutput.t121 2.82907
R6368 CSoutput.n325 CSoutput.t105 2.82907
R6369 CSoutput.n326 CSoutput.t107 2.82907
R6370 CSoutput.n326 CSoutput.t115 2.82907
R6371 CSoutput.n328 CSoutput.t134 2.82907
R6372 CSoutput.n328 CSoutput.t29 2.82907
R6373 CSoutput.n330 CSoutput.t7 2.82907
R6374 CSoutput.n330 CSoutput.t80 2.82907
R6375 CSoutput.n332 CSoutput.t110 2.82907
R6376 CSoutput.n332 CSoutput.t137 2.82907
R6377 CSoutput.n334 CSoutput.t84 2.82907
R6378 CSoutput.n334 CSoutput.t92 2.82907
R6379 CSoutput.n336 CSoutput.t0 2.82907
R6380 CSoutput.n336 CSoutput.t131 2.82907
R6381 CSoutput.n338 CSoutput.t87 2.82907
R6382 CSoutput.n338 CSoutput.t10 2.82907
R6383 CSoutput.n75 CSoutput.n1 2.45513
R6384 CSoutput.n193 CSoutput.n191 2.251
R6385 CSoutput.n193 CSoutput.n190 2.251
R6386 CSoutput.n193 CSoutput.n189 2.251
R6387 CSoutput.n193 CSoutput.n188 2.251
R6388 CSoutput.n162 CSoutput.n161 2.251
R6389 CSoutput.n162 CSoutput.n160 2.251
R6390 CSoutput.n162 CSoutput.n159 2.251
R6391 CSoutput.n162 CSoutput.n158 2.251
R6392 CSoutput.n235 CSoutput.n234 2.251
R6393 CSoutput.n200 CSoutput.n198 2.251
R6394 CSoutput.n200 CSoutput.n197 2.251
R6395 CSoutput.n200 CSoutput.n196 2.251
R6396 CSoutput.n218 CSoutput.n200 2.251
R6397 CSoutput.n206 CSoutput.n205 2.251
R6398 CSoutput.n206 CSoutput.n204 2.251
R6399 CSoutput.n206 CSoutput.n203 2.251
R6400 CSoutput.n206 CSoutput.n202 2.251
R6401 CSoutput.n232 CSoutput.n172 2.251
R6402 CSoutput.n227 CSoutput.n225 2.251
R6403 CSoutput.n227 CSoutput.n224 2.251
R6404 CSoutput.n227 CSoutput.n223 2.251
R6405 CSoutput.n227 CSoutput.n222 2.251
R6406 CSoutput.n128 CSoutput.n127 2.251
R6407 CSoutput.n128 CSoutput.n126 2.251
R6408 CSoutput.n128 CSoutput.n125 2.251
R6409 CSoutput.n128 CSoutput.n124 2.251
R6410 CSoutput.n245 CSoutput.n244 2.251
R6411 CSoutput.n162 CSoutput.n142 2.2505
R6412 CSoutput.n157 CSoutput.n142 2.2505
R6413 CSoutput.n155 CSoutput.n142 2.2505
R6414 CSoutput.n154 CSoutput.n142 2.2505
R6415 CSoutput.n239 CSoutput.n142 2.2505
R6416 CSoutput.n237 CSoutput.n142 2.2505
R6417 CSoutput.n235 CSoutput.n142 2.2505
R6418 CSoutput.n165 CSoutput.n142 2.2505
R6419 CSoutput.n164 CSoutput.n142 2.2505
R6420 CSoutput.n168 CSoutput.n142 2.2505
R6421 CSoutput.n167 CSoutput.n142 2.2505
R6422 CSoutput.n150 CSoutput.n142 2.2505
R6423 CSoutput.n242 CSoutput.n142 2.2505
R6424 CSoutput.n242 CSoutput.n241 2.2505
R6425 CSoutput.n206 CSoutput.n177 2.2505
R6426 CSoutput.n187 CSoutput.n177 2.2505
R6427 CSoutput.n208 CSoutput.n177 2.2505
R6428 CSoutput.n186 CSoutput.n177 2.2505
R6429 CSoutput.n210 CSoutput.n177 2.2505
R6430 CSoutput.n177 CSoutput.n171 2.2505
R6431 CSoutput.n232 CSoutput.n177 2.2505
R6432 CSoutput.n230 CSoutput.n177 2.2505
R6433 CSoutput.n212 CSoutput.n177 2.2505
R6434 CSoutput.n184 CSoutput.n177 2.2505
R6435 CSoutput.n214 CSoutput.n177 2.2505
R6436 CSoutput.n183 CSoutput.n177 2.2505
R6437 CSoutput.n228 CSoutput.n177 2.2505
R6438 CSoutput.n228 CSoutput.n181 2.2505
R6439 CSoutput.n128 CSoutput.n108 2.2505
R6440 CSoutput.n123 CSoutput.n108 2.2505
R6441 CSoutput.n121 CSoutput.n108 2.2505
R6442 CSoutput.n120 CSoutput.n108 2.2505
R6443 CSoutput.n249 CSoutput.n108 2.2505
R6444 CSoutput.n247 CSoutput.n108 2.2505
R6445 CSoutput.n245 CSoutput.n108 2.2505
R6446 CSoutput.n131 CSoutput.n108 2.2505
R6447 CSoutput.n130 CSoutput.n108 2.2505
R6448 CSoutput.n134 CSoutput.n108 2.2505
R6449 CSoutput.n133 CSoutput.n108 2.2505
R6450 CSoutput.n116 CSoutput.n108 2.2505
R6451 CSoutput.n252 CSoutput.n108 2.2505
R6452 CSoutput.n252 CSoutput.n251 2.2505
R6453 CSoutput.n170 CSoutput.n163 2.25024
R6454 CSoutput.n170 CSoutput.n156 2.25024
R6455 CSoutput.n238 CSoutput.n170 2.25024
R6456 CSoutput.n170 CSoutput.n166 2.25024
R6457 CSoutput.n170 CSoutput.n169 2.25024
R6458 CSoutput.n170 CSoutput.n137 2.25024
R6459 CSoutput.n220 CSoutput.n217 2.25024
R6460 CSoutput.n220 CSoutput.n216 2.25024
R6461 CSoutput.n220 CSoutput.n215 2.25024
R6462 CSoutput.n220 CSoutput.n182 2.25024
R6463 CSoutput.n220 CSoutput.n219 2.25024
R6464 CSoutput.n221 CSoutput.n220 2.25024
R6465 CSoutput.n136 CSoutput.n129 2.25024
R6466 CSoutput.n136 CSoutput.n122 2.25024
R6467 CSoutput.n248 CSoutput.n136 2.25024
R6468 CSoutput.n136 CSoutput.n132 2.25024
R6469 CSoutput.n136 CSoutput.n135 2.25024
R6470 CSoutput.n136 CSoutput.n103 2.25024
R6471 CSoutput.n276 CSoutput.n102 1.95131
R6472 CSoutput.n237 CSoutput.n147 1.50111
R6473 CSoutput.n185 CSoutput.n171 1.50111
R6474 CSoutput.n247 CSoutput.n113 1.50111
R6475 CSoutput.n193 CSoutput.n192 1.501
R6476 CSoutput.n200 CSoutput.n199 1.501
R6477 CSoutput.n227 CSoutput.n226 1.501
R6478 CSoutput.n241 CSoutput.n152 1.12536
R6479 CSoutput.n241 CSoutput.n153 1.12536
R6480 CSoutput.n241 CSoutput.n240 1.12536
R6481 CSoutput.n201 CSoutput.n181 1.12536
R6482 CSoutput.n207 CSoutput.n181 1.12536
R6483 CSoutput.n209 CSoutput.n181 1.12536
R6484 CSoutput.n251 CSoutput.n118 1.12536
R6485 CSoutput.n251 CSoutput.n119 1.12536
R6486 CSoutput.n251 CSoutput.n250 1.12536
R6487 CSoutput.n241 CSoutput.n148 1.12536
R6488 CSoutput.n241 CSoutput.n149 1.12536
R6489 CSoutput.n241 CSoutput.n151 1.12536
R6490 CSoutput.n231 CSoutput.n181 1.12536
R6491 CSoutput.n211 CSoutput.n181 1.12536
R6492 CSoutput.n213 CSoutput.n181 1.12536
R6493 CSoutput.n251 CSoutput.n114 1.12536
R6494 CSoutput.n251 CSoutput.n115 1.12536
R6495 CSoutput.n251 CSoutput.n117 1.12536
R6496 CSoutput.n31 CSoutput.n30 0.669944
R6497 CSoutput.n62 CSoutput.n61 0.669944
R6498 CSoutput.n312 CSoutput.n310 0.573776
R6499 CSoutput.n314 CSoutput.n312 0.573776
R6500 CSoutput.n316 CSoutput.n314 0.573776
R6501 CSoutput.n318 CSoutput.n316 0.573776
R6502 CSoutput.n320 CSoutput.n318 0.573776
R6503 CSoutput.n322 CSoutput.n320 0.573776
R6504 CSoutput.n296 CSoutput.n294 0.573776
R6505 CSoutput.n298 CSoutput.n296 0.573776
R6506 CSoutput.n300 CSoutput.n298 0.573776
R6507 CSoutput.n302 CSoutput.n300 0.573776
R6508 CSoutput.n304 CSoutput.n302 0.573776
R6509 CSoutput.n306 CSoutput.n304 0.573776
R6510 CSoutput.n281 CSoutput.n279 0.573776
R6511 CSoutput.n283 CSoutput.n281 0.573776
R6512 CSoutput.n285 CSoutput.n283 0.573776
R6513 CSoutput.n287 CSoutput.n285 0.573776
R6514 CSoutput.n289 CSoutput.n287 0.573776
R6515 CSoutput.n291 CSoutput.n289 0.573776
R6516 CSoutput.n370 CSoutput.n368 0.573776
R6517 CSoutput.n368 CSoutput.n366 0.573776
R6518 CSoutput.n366 CSoutput.n364 0.573776
R6519 CSoutput.n364 CSoutput.n362 0.573776
R6520 CSoutput.n362 CSoutput.n360 0.573776
R6521 CSoutput.n360 CSoutput.n358 0.573776
R6522 CSoutput.n354 CSoutput.n352 0.573776
R6523 CSoutput.n352 CSoutput.n350 0.573776
R6524 CSoutput.n350 CSoutput.n348 0.573776
R6525 CSoutput.n348 CSoutput.n346 0.573776
R6526 CSoutput.n346 CSoutput.n344 0.573776
R6527 CSoutput.n344 CSoutput.n342 0.573776
R6528 CSoutput.n339 CSoutput.n337 0.573776
R6529 CSoutput.n337 CSoutput.n335 0.573776
R6530 CSoutput.n335 CSoutput.n333 0.573776
R6531 CSoutput.n333 CSoutput.n331 0.573776
R6532 CSoutput.n331 CSoutput.n329 0.573776
R6533 CSoutput.n329 CSoutput.n327 0.573776
R6534 CSoutput.n373 CSoutput.n252 0.53442
R6535 CSoutput.n272 CSoutput.n270 0.358259
R6536 CSoutput.n274 CSoutput.n272 0.358259
R6537 CSoutput.n264 CSoutput.n262 0.358259
R6538 CSoutput.n266 CSoutput.n264 0.358259
R6539 CSoutput.n257 CSoutput.n255 0.358259
R6540 CSoutput.n259 CSoutput.n257 0.358259
R6541 CSoutput.n100 CSoutput.n98 0.358259
R6542 CSoutput.n98 CSoutput.n96 0.358259
R6543 CSoutput.n92 CSoutput.n90 0.358259
R6544 CSoutput.n90 CSoutput.n88 0.358259
R6545 CSoutput.n85 CSoutput.n83 0.358259
R6546 CSoutput.n83 CSoutput.n81 0.358259
R6547 CSoutput.n21 CSoutput.n20 0.169105
R6548 CSoutput.n21 CSoutput.n16 0.169105
R6549 CSoutput.n26 CSoutput.n16 0.169105
R6550 CSoutput.n27 CSoutput.n26 0.169105
R6551 CSoutput.n27 CSoutput.n14 0.169105
R6552 CSoutput.n32 CSoutput.n14 0.169105
R6553 CSoutput.n33 CSoutput.n32 0.169105
R6554 CSoutput.n34 CSoutput.n33 0.169105
R6555 CSoutput.n34 CSoutput.n12 0.169105
R6556 CSoutput.n39 CSoutput.n12 0.169105
R6557 CSoutput.n40 CSoutput.n39 0.169105
R6558 CSoutput.n40 CSoutput.n10 0.169105
R6559 CSoutput.n45 CSoutput.n10 0.169105
R6560 CSoutput.n46 CSoutput.n45 0.169105
R6561 CSoutput.n47 CSoutput.n46 0.169105
R6562 CSoutput.n47 CSoutput.n8 0.169105
R6563 CSoutput.n52 CSoutput.n8 0.169105
R6564 CSoutput.n53 CSoutput.n52 0.169105
R6565 CSoutput.n53 CSoutput.n6 0.169105
R6566 CSoutput.n58 CSoutput.n6 0.169105
R6567 CSoutput.n59 CSoutput.n58 0.169105
R6568 CSoutput.n60 CSoutput.n59 0.169105
R6569 CSoutput.n60 CSoutput.n4 0.169105
R6570 CSoutput.n66 CSoutput.n4 0.169105
R6571 CSoutput.n67 CSoutput.n66 0.169105
R6572 CSoutput.n68 CSoutput.n67 0.169105
R6573 CSoutput.n68 CSoutput.n2 0.169105
R6574 CSoutput.n73 CSoutput.n2 0.169105
R6575 CSoutput.n74 CSoutput.n73 0.169105
R6576 CSoutput.n74 CSoutput.n0 0.169105
R6577 CSoutput.n78 CSoutput.n0 0.169105
R6578 CSoutput.n195 CSoutput.n194 0.0910737
R6579 CSoutput.n246 CSoutput.n243 0.0723685
R6580 CSoutput.n200 CSoutput.n195 0.0522944
R6581 CSoutput.n243 CSoutput.n242 0.0499135
R6582 CSoutput.n194 CSoutput.n193 0.0499135
R6583 CSoutput.n228 CSoutput.n227 0.0464294
R6584 CSoutput.n236 CSoutput.n233 0.0391444
R6585 CSoutput.n195 CSoutput.t154 0.023435
R6586 CSoutput.n243 CSoutput.t146 0.02262
R6587 CSoutput.n194 CSoutput.t148 0.02262
R6588 CSoutput CSoutput.n373 0.0052
R6589 CSoutput.n165 CSoutput.n148 0.00365111
R6590 CSoutput.n168 CSoutput.n149 0.00365111
R6591 CSoutput.n151 CSoutput.n150 0.00365111
R6592 CSoutput.n193 CSoutput.n152 0.00365111
R6593 CSoutput.n157 CSoutput.n153 0.00365111
R6594 CSoutput.n240 CSoutput.n154 0.00365111
R6595 CSoutput.n231 CSoutput.n230 0.00365111
R6596 CSoutput.n211 CSoutput.n184 0.00365111
R6597 CSoutput.n213 CSoutput.n183 0.00365111
R6598 CSoutput.n201 CSoutput.n200 0.00365111
R6599 CSoutput.n207 CSoutput.n187 0.00365111
R6600 CSoutput.n209 CSoutput.n186 0.00365111
R6601 CSoutput.n131 CSoutput.n114 0.00365111
R6602 CSoutput.n134 CSoutput.n115 0.00365111
R6603 CSoutput.n117 CSoutput.n116 0.00365111
R6604 CSoutput.n227 CSoutput.n118 0.00365111
R6605 CSoutput.n123 CSoutput.n119 0.00365111
R6606 CSoutput.n250 CSoutput.n120 0.00365111
R6607 CSoutput.n162 CSoutput.n152 0.00340054
R6608 CSoutput.n155 CSoutput.n153 0.00340054
R6609 CSoutput.n240 CSoutput.n239 0.00340054
R6610 CSoutput.n235 CSoutput.n148 0.00340054
R6611 CSoutput.n164 CSoutput.n149 0.00340054
R6612 CSoutput.n167 CSoutput.n151 0.00340054
R6613 CSoutput.n206 CSoutput.n201 0.00340054
R6614 CSoutput.n208 CSoutput.n207 0.00340054
R6615 CSoutput.n210 CSoutput.n209 0.00340054
R6616 CSoutput.n232 CSoutput.n231 0.00340054
R6617 CSoutput.n212 CSoutput.n211 0.00340054
R6618 CSoutput.n214 CSoutput.n213 0.00340054
R6619 CSoutput.n128 CSoutput.n118 0.00340054
R6620 CSoutput.n121 CSoutput.n119 0.00340054
R6621 CSoutput.n250 CSoutput.n249 0.00340054
R6622 CSoutput.n245 CSoutput.n114 0.00340054
R6623 CSoutput.n130 CSoutput.n115 0.00340054
R6624 CSoutput.n133 CSoutput.n117 0.00340054
R6625 CSoutput.n163 CSoutput.n157 0.00252698
R6626 CSoutput.n156 CSoutput.n154 0.00252698
R6627 CSoutput.n238 CSoutput.n237 0.00252698
R6628 CSoutput.n166 CSoutput.n164 0.00252698
R6629 CSoutput.n169 CSoutput.n167 0.00252698
R6630 CSoutput.n242 CSoutput.n137 0.00252698
R6631 CSoutput.n163 CSoutput.n162 0.00252698
R6632 CSoutput.n156 CSoutput.n155 0.00252698
R6633 CSoutput.n239 CSoutput.n238 0.00252698
R6634 CSoutput.n166 CSoutput.n165 0.00252698
R6635 CSoutput.n169 CSoutput.n168 0.00252698
R6636 CSoutput.n150 CSoutput.n137 0.00252698
R6637 CSoutput.n217 CSoutput.n187 0.00252698
R6638 CSoutput.n216 CSoutput.n186 0.00252698
R6639 CSoutput.n215 CSoutput.n171 0.00252698
R6640 CSoutput.n212 CSoutput.n182 0.00252698
R6641 CSoutput.n219 CSoutput.n214 0.00252698
R6642 CSoutput.n228 CSoutput.n221 0.00252698
R6643 CSoutput.n217 CSoutput.n206 0.00252698
R6644 CSoutput.n216 CSoutput.n208 0.00252698
R6645 CSoutput.n215 CSoutput.n210 0.00252698
R6646 CSoutput.n230 CSoutput.n182 0.00252698
R6647 CSoutput.n219 CSoutput.n184 0.00252698
R6648 CSoutput.n221 CSoutput.n183 0.00252698
R6649 CSoutput.n129 CSoutput.n123 0.00252698
R6650 CSoutput.n122 CSoutput.n120 0.00252698
R6651 CSoutput.n248 CSoutput.n247 0.00252698
R6652 CSoutput.n132 CSoutput.n130 0.00252698
R6653 CSoutput.n135 CSoutput.n133 0.00252698
R6654 CSoutput.n252 CSoutput.n103 0.00252698
R6655 CSoutput.n129 CSoutput.n128 0.00252698
R6656 CSoutput.n122 CSoutput.n121 0.00252698
R6657 CSoutput.n249 CSoutput.n248 0.00252698
R6658 CSoutput.n132 CSoutput.n131 0.00252698
R6659 CSoutput.n135 CSoutput.n134 0.00252698
R6660 CSoutput.n116 CSoutput.n103 0.00252698
R6661 CSoutput.n237 CSoutput.n236 0.0020275
R6662 CSoutput.n236 CSoutput.n235 0.0020275
R6663 CSoutput.n233 CSoutput.n171 0.0020275
R6664 CSoutput.n233 CSoutput.n232 0.0020275
R6665 CSoutput.n247 CSoutput.n246 0.0020275
R6666 CSoutput.n246 CSoutput.n245 0.0020275
R6667 CSoutput.n147 CSoutput.n146 0.00166668
R6668 CSoutput.n229 CSoutput.n185 0.00166668
R6669 CSoutput.n113 CSoutput.n112 0.00166668
R6670 CSoutput.n251 CSoutput.n113 0.00133328
R6671 CSoutput.n185 CSoutput.n181 0.00133328
R6672 CSoutput.n241 CSoutput.n147 0.00133328
R6673 CSoutput.n244 CSoutput.n136 0.001
R6674 CSoutput.n222 CSoutput.n136 0.001
R6675 CSoutput.n124 CSoutput.n104 0.001
R6676 CSoutput.n223 CSoutput.n104 0.001
R6677 CSoutput.n125 CSoutput.n105 0.001
R6678 CSoutput.n224 CSoutput.n105 0.001
R6679 CSoutput.n126 CSoutput.n106 0.001
R6680 CSoutput.n225 CSoutput.n106 0.001
R6681 CSoutput.n127 CSoutput.n107 0.001
R6682 CSoutput.n226 CSoutput.n107 0.001
R6683 CSoutput.n220 CSoutput.n172 0.001
R6684 CSoutput.n220 CSoutput.n218 0.001
R6685 CSoutput.n202 CSoutput.n173 0.001
R6686 CSoutput.n196 CSoutput.n173 0.001
R6687 CSoutput.n203 CSoutput.n174 0.001
R6688 CSoutput.n197 CSoutput.n174 0.001
R6689 CSoutput.n204 CSoutput.n175 0.001
R6690 CSoutput.n198 CSoutput.n175 0.001
R6691 CSoutput.n205 CSoutput.n176 0.001
R6692 CSoutput.n199 CSoutput.n176 0.001
R6693 CSoutput.n234 CSoutput.n170 0.001
R6694 CSoutput.n188 CSoutput.n170 0.001
R6695 CSoutput.n158 CSoutput.n138 0.001
R6696 CSoutput.n189 CSoutput.n138 0.001
R6697 CSoutput.n159 CSoutput.n139 0.001
R6698 CSoutput.n190 CSoutput.n139 0.001
R6699 CSoutput.n160 CSoutput.n140 0.001
R6700 CSoutput.n191 CSoutput.n140 0.001
R6701 CSoutput.n161 CSoutput.n141 0.001
R6702 CSoutput.n192 CSoutput.n141 0.001
R6703 CSoutput.n192 CSoutput.n142 0.001
R6704 CSoutput.n191 CSoutput.n143 0.001
R6705 CSoutput.n190 CSoutput.n144 0.001
R6706 CSoutput.n189 CSoutput.t165 0.001
R6707 CSoutput.n188 CSoutput.n145 0.001
R6708 CSoutput.n161 CSoutput.n143 0.001
R6709 CSoutput.n160 CSoutput.n144 0.001
R6710 CSoutput.n159 CSoutput.t165 0.001
R6711 CSoutput.n158 CSoutput.n145 0.001
R6712 CSoutput.n234 CSoutput.n146 0.001
R6713 CSoutput.n199 CSoutput.n177 0.001
R6714 CSoutput.n198 CSoutput.n178 0.001
R6715 CSoutput.n197 CSoutput.n179 0.001
R6716 CSoutput.n196 CSoutput.t144 0.001
R6717 CSoutput.n218 CSoutput.n180 0.001
R6718 CSoutput.n205 CSoutput.n178 0.001
R6719 CSoutput.n204 CSoutput.n179 0.001
R6720 CSoutput.n203 CSoutput.t144 0.001
R6721 CSoutput.n202 CSoutput.n180 0.001
R6722 CSoutput.n229 CSoutput.n172 0.001
R6723 CSoutput.n226 CSoutput.n108 0.001
R6724 CSoutput.n225 CSoutput.n109 0.001
R6725 CSoutput.n224 CSoutput.n110 0.001
R6726 CSoutput.n223 CSoutput.t151 0.001
R6727 CSoutput.n222 CSoutput.n111 0.001
R6728 CSoutput.n127 CSoutput.n109 0.001
R6729 CSoutput.n126 CSoutput.n110 0.001
R6730 CSoutput.n125 CSoutput.t151 0.001
R6731 CSoutput.n124 CSoutput.n111 0.001
R6732 CSoutput.n244 CSoutput.n112 0.001
R6733 commonsourceibias.n35 commonsourceibias.t16 223.028
R6734 commonsourceibias.n128 commonsourceibias.t129 223.028
R6735 commonsourceibias.n307 commonsourceibias.t139 223.028
R6736 commonsourceibias.n217 commonsourceibias.t108 223.028
R6737 commonsourceibias.n454 commonsourceibias.t14 223.028
R6738 commonsourceibias.n395 commonsourceibias.t112 223.028
R6739 commonsourceibias.n679 commonsourceibias.t73 223.028
R6740 commonsourceibias.n589 commonsourceibias.t99 223.028
R6741 commonsourceibias.n99 commonsourceibias.t20 207.983
R6742 commonsourceibias.n192 commonsourceibias.t120 207.983
R6743 commonsourceibias.n371 commonsourceibias.t147 207.983
R6744 commonsourceibias.n281 commonsourceibias.t68 207.983
R6745 commonsourceibias.n520 commonsourceibias.t58 207.983
R6746 commonsourceibias.n566 commonsourceibias.t93 207.983
R6747 commonsourceibias.n745 commonsourceibias.t82 207.983
R6748 commonsourceibias.n655 commonsourceibias.t150 207.983
R6749 commonsourceibias.n97 commonsourceibias.t48 168.701
R6750 commonsourceibias.n91 commonsourceibias.t30 168.701
R6751 commonsourceibias.n17 commonsourceibias.t6 168.701
R6752 commonsourceibias.n83 commonsourceibias.t28 168.701
R6753 commonsourceibias.n77 commonsourceibias.t24 168.701
R6754 commonsourceibias.n22 commonsourceibias.t52 168.701
R6755 commonsourceibias.n69 commonsourceibias.t32 168.701
R6756 commonsourceibias.n63 commonsourceibias.t22 168.701
R6757 commonsourceibias.n25 commonsourceibias.t42 168.701
R6758 commonsourceibias.n27 commonsourceibias.t2 168.701
R6759 commonsourceibias.n29 commonsourceibias.t56 168.701
R6760 commonsourceibias.n46 commonsourceibias.t8 168.701
R6761 commonsourceibias.n40 commonsourceibias.t10 168.701
R6762 commonsourceibias.n34 commonsourceibias.t50 168.701
R6763 commonsourceibias.n190 commonsourceibias.t65 168.701
R6764 commonsourceibias.n184 commonsourceibias.t126 168.701
R6765 commonsourceibias.n5 commonsourceibias.t121 168.701
R6766 commonsourceibias.n176 commonsourceibias.t135 168.701
R6767 commonsourceibias.n170 commonsourceibias.t117 168.701
R6768 commonsourceibias.n10 commonsourceibias.t102 168.701
R6769 commonsourceibias.n162 commonsourceibias.t125 168.701
R6770 commonsourceibias.n156 commonsourceibias.t119 168.701
R6771 commonsourceibias.n118 commonsourceibias.t79 168.701
R6772 commonsourceibias.n120 commonsourceibias.t106 168.701
R6773 commonsourceibias.n122 commonsourceibias.t96 168.701
R6774 commonsourceibias.n139 commonsourceibias.t141 168.701
R6775 commonsourceibias.n133 commonsourceibias.t116 168.701
R6776 commonsourceibias.n127 commonsourceibias.t152 168.701
R6777 commonsourceibias.n306 commonsourceibias.t130 168.701
R6778 commonsourceibias.n312 commonsourceibias.t76 168.701
R6779 commonsourceibias.n318 commonsourceibias.t149 168.701
R6780 commonsourceibias.n301 commonsourceibias.t133 168.701
R6781 commonsourceibias.n299 commonsourceibias.t137 168.701
R6782 commonsourceibias.n297 commonsourceibias.t64 168.701
R6783 commonsourceibias.n335 commonsourceibias.t138 168.701
R6784 commonsourceibias.n341 commonsourceibias.t146 168.701
R6785 commonsourceibias.n294 commonsourceibias.t118 168.701
R6786 commonsourceibias.n349 commonsourceibias.t89 168.701
R6787 commonsourceibias.n355 commonsourceibias.t155 168.701
R6788 commonsourceibias.n289 commonsourceibias.t124 168.701
R6789 commonsourceibias.n363 commonsourceibias.t128 168.701
R6790 commonsourceibias.n369 commonsourceibias.t75 168.701
R6791 commonsourceibias.n279 commonsourceibias.t159 168.701
R6792 commonsourceibias.n273 commonsourceibias.t148 168.701
R6793 commonsourceibias.n199 commonsourceibias.t78 168.701
R6794 commonsourceibias.n265 commonsourceibias.t158 168.701
R6795 commonsourceibias.n259 commonsourceibias.t85 168.701
R6796 commonsourceibias.n204 commonsourceibias.t77 168.701
R6797 commonsourceibias.n251 commonsourceibias.t157 168.701
R6798 commonsourceibias.n245 commonsourceibias.t94 168.701
R6799 commonsourceibias.n207 commonsourceibias.t113 168.701
R6800 commonsourceibias.n209 commonsourceibias.t156 168.701
R6801 commonsourceibias.n211 commonsourceibias.t92 168.701
R6802 commonsourceibias.n228 commonsourceibias.t109 168.701
R6803 commonsourceibias.n222 commonsourceibias.t105 168.701
R6804 commonsourceibias.n216 commonsourceibias.t91 168.701
R6805 commonsourceibias.n453 commonsourceibias.t0 168.701
R6806 commonsourceibias.n459 commonsourceibias.t38 168.701
R6807 commonsourceibias.n465 commonsourceibias.t18 168.701
R6808 commonsourceibias.n448 commonsourceibias.t62 168.701
R6809 commonsourceibias.n446 commonsourceibias.t40 168.701
R6810 commonsourceibias.n444 commonsourceibias.t60 168.701
R6811 commonsourceibias.n482 commonsourceibias.t34 168.701
R6812 commonsourceibias.n488 commonsourceibias.t4 168.701
R6813 commonsourceibias.n490 commonsourceibias.t46 168.701
R6814 commonsourceibias.n497 commonsourceibias.t36 168.701
R6815 commonsourceibias.n503 commonsourceibias.t26 168.701
R6816 commonsourceibias.n505 commonsourceibias.t54 168.701
R6817 commonsourceibias.n512 commonsourceibias.t12 168.701
R6818 commonsourceibias.n518 commonsourceibias.t44 168.701
R6819 commonsourceibias.n564 commonsourceibias.t134 168.701
R6820 commonsourceibias.n558 commonsourceibias.t114 168.701
R6821 commonsourceibias.n551 commonsourceibias.t95 168.701
R6822 commonsourceibias.n549 commonsourceibias.t123 168.701
R6823 commonsourceibias.n543 commonsourceibias.t88 168.701
R6824 commonsourceibias.n536 commonsourceibias.t74 168.701
R6825 commonsourceibias.n534 commonsourceibias.t104 168.701
R6826 commonsourceibias.n394 commonsourceibias.t131 168.701
R6827 commonsourceibias.n400 commonsourceibias.t84 168.701
R6828 commonsourceibias.n406 commonsourceibias.t127 168.701
R6829 commonsourceibias.n389 commonsourceibias.t151 168.701
R6830 commonsourceibias.n387 commonsourceibias.t83 168.701
R6831 commonsourceibias.n385 commonsourceibias.t140 168.701
R6832 commonsourceibias.n423 commonsourceibias.t90 168.701
R6833 commonsourceibias.n678 commonsourceibias.t145 168.701
R6834 commonsourceibias.n684 commonsourceibias.t111 168.701
R6835 commonsourceibias.n690 commonsourceibias.t86 168.701
R6836 commonsourceibias.n673 commonsourceibias.t153 168.701
R6837 commonsourceibias.n671 commonsourceibias.t132 168.701
R6838 commonsourceibias.n669 commonsourceibias.t103 168.701
R6839 commonsourceibias.n707 commonsourceibias.t69 168.701
R6840 commonsourceibias.n713 commonsourceibias.t81 168.701
R6841 commonsourceibias.n715 commonsourceibias.t110 168.701
R6842 commonsourceibias.n722 commonsourceibias.t115 168.701
R6843 commonsourceibias.n728 commonsourceibias.t97 168.701
R6844 commonsourceibias.n730 commonsourceibias.t136 168.701
R6845 commonsourceibias.n737 commonsourceibias.t122 168.701
R6846 commonsourceibias.n743 commonsourceibias.t107 168.701
R6847 commonsourceibias.n588 commonsourceibias.t71 168.701
R6848 commonsourceibias.n594 commonsourceibias.t87 168.701
R6849 commonsourceibias.n600 commonsourceibias.t100 168.701
R6850 commonsourceibias.n583 commonsourceibias.t72 168.701
R6851 commonsourceibias.n581 commonsourceibias.t80 168.701
R6852 commonsourceibias.n579 commonsourceibias.t101 168.701
R6853 commonsourceibias.n617 commonsourceibias.t70 168.701
R6854 commonsourceibias.n623 commonsourceibias.t144 168.701
R6855 commonsourceibias.n625 commonsourceibias.t98 168.701
R6856 commonsourceibias.n632 commonsourceibias.t67 168.701
R6857 commonsourceibias.n638 commonsourceibias.t143 168.701
R6858 commonsourceibias.n640 commonsourceibias.t154 168.701
R6859 commonsourceibias.n647 commonsourceibias.t66 168.701
R6860 commonsourceibias.n653 commonsourceibias.t142 168.701
R6861 commonsourceibias.n36 commonsourceibias.n33 161.3
R6862 commonsourceibias.n38 commonsourceibias.n37 161.3
R6863 commonsourceibias.n39 commonsourceibias.n32 161.3
R6864 commonsourceibias.n42 commonsourceibias.n41 161.3
R6865 commonsourceibias.n43 commonsourceibias.n31 161.3
R6866 commonsourceibias.n45 commonsourceibias.n44 161.3
R6867 commonsourceibias.n47 commonsourceibias.n30 161.3
R6868 commonsourceibias.n49 commonsourceibias.n48 161.3
R6869 commonsourceibias.n51 commonsourceibias.n50 161.3
R6870 commonsourceibias.n52 commonsourceibias.n28 161.3
R6871 commonsourceibias.n54 commonsourceibias.n53 161.3
R6872 commonsourceibias.n56 commonsourceibias.n55 161.3
R6873 commonsourceibias.n57 commonsourceibias.n26 161.3
R6874 commonsourceibias.n59 commonsourceibias.n58 161.3
R6875 commonsourceibias.n61 commonsourceibias.n60 161.3
R6876 commonsourceibias.n62 commonsourceibias.n24 161.3
R6877 commonsourceibias.n65 commonsourceibias.n64 161.3
R6878 commonsourceibias.n66 commonsourceibias.n23 161.3
R6879 commonsourceibias.n68 commonsourceibias.n67 161.3
R6880 commonsourceibias.n70 commonsourceibias.n21 161.3
R6881 commonsourceibias.n72 commonsourceibias.n71 161.3
R6882 commonsourceibias.n73 commonsourceibias.n20 161.3
R6883 commonsourceibias.n75 commonsourceibias.n74 161.3
R6884 commonsourceibias.n76 commonsourceibias.n19 161.3
R6885 commonsourceibias.n79 commonsourceibias.n78 161.3
R6886 commonsourceibias.n80 commonsourceibias.n18 161.3
R6887 commonsourceibias.n82 commonsourceibias.n81 161.3
R6888 commonsourceibias.n84 commonsourceibias.n16 161.3
R6889 commonsourceibias.n86 commonsourceibias.n85 161.3
R6890 commonsourceibias.n87 commonsourceibias.n15 161.3
R6891 commonsourceibias.n89 commonsourceibias.n88 161.3
R6892 commonsourceibias.n90 commonsourceibias.n14 161.3
R6893 commonsourceibias.n93 commonsourceibias.n92 161.3
R6894 commonsourceibias.n94 commonsourceibias.n13 161.3
R6895 commonsourceibias.n96 commonsourceibias.n95 161.3
R6896 commonsourceibias.n98 commonsourceibias.n12 161.3
R6897 commonsourceibias.n129 commonsourceibias.n126 161.3
R6898 commonsourceibias.n131 commonsourceibias.n130 161.3
R6899 commonsourceibias.n132 commonsourceibias.n125 161.3
R6900 commonsourceibias.n135 commonsourceibias.n134 161.3
R6901 commonsourceibias.n136 commonsourceibias.n124 161.3
R6902 commonsourceibias.n138 commonsourceibias.n137 161.3
R6903 commonsourceibias.n140 commonsourceibias.n123 161.3
R6904 commonsourceibias.n142 commonsourceibias.n141 161.3
R6905 commonsourceibias.n144 commonsourceibias.n143 161.3
R6906 commonsourceibias.n145 commonsourceibias.n121 161.3
R6907 commonsourceibias.n147 commonsourceibias.n146 161.3
R6908 commonsourceibias.n149 commonsourceibias.n148 161.3
R6909 commonsourceibias.n150 commonsourceibias.n119 161.3
R6910 commonsourceibias.n152 commonsourceibias.n151 161.3
R6911 commonsourceibias.n154 commonsourceibias.n153 161.3
R6912 commonsourceibias.n155 commonsourceibias.n117 161.3
R6913 commonsourceibias.n158 commonsourceibias.n157 161.3
R6914 commonsourceibias.n159 commonsourceibias.n11 161.3
R6915 commonsourceibias.n161 commonsourceibias.n160 161.3
R6916 commonsourceibias.n163 commonsourceibias.n9 161.3
R6917 commonsourceibias.n165 commonsourceibias.n164 161.3
R6918 commonsourceibias.n166 commonsourceibias.n8 161.3
R6919 commonsourceibias.n168 commonsourceibias.n167 161.3
R6920 commonsourceibias.n169 commonsourceibias.n7 161.3
R6921 commonsourceibias.n172 commonsourceibias.n171 161.3
R6922 commonsourceibias.n173 commonsourceibias.n6 161.3
R6923 commonsourceibias.n175 commonsourceibias.n174 161.3
R6924 commonsourceibias.n177 commonsourceibias.n4 161.3
R6925 commonsourceibias.n179 commonsourceibias.n178 161.3
R6926 commonsourceibias.n180 commonsourceibias.n3 161.3
R6927 commonsourceibias.n182 commonsourceibias.n181 161.3
R6928 commonsourceibias.n183 commonsourceibias.n2 161.3
R6929 commonsourceibias.n186 commonsourceibias.n185 161.3
R6930 commonsourceibias.n187 commonsourceibias.n1 161.3
R6931 commonsourceibias.n189 commonsourceibias.n188 161.3
R6932 commonsourceibias.n191 commonsourceibias.n0 161.3
R6933 commonsourceibias.n370 commonsourceibias.n284 161.3
R6934 commonsourceibias.n368 commonsourceibias.n367 161.3
R6935 commonsourceibias.n366 commonsourceibias.n285 161.3
R6936 commonsourceibias.n365 commonsourceibias.n364 161.3
R6937 commonsourceibias.n362 commonsourceibias.n286 161.3
R6938 commonsourceibias.n361 commonsourceibias.n360 161.3
R6939 commonsourceibias.n359 commonsourceibias.n287 161.3
R6940 commonsourceibias.n358 commonsourceibias.n357 161.3
R6941 commonsourceibias.n356 commonsourceibias.n288 161.3
R6942 commonsourceibias.n354 commonsourceibias.n353 161.3
R6943 commonsourceibias.n352 commonsourceibias.n290 161.3
R6944 commonsourceibias.n351 commonsourceibias.n350 161.3
R6945 commonsourceibias.n348 commonsourceibias.n291 161.3
R6946 commonsourceibias.n347 commonsourceibias.n346 161.3
R6947 commonsourceibias.n345 commonsourceibias.n292 161.3
R6948 commonsourceibias.n344 commonsourceibias.n343 161.3
R6949 commonsourceibias.n342 commonsourceibias.n293 161.3
R6950 commonsourceibias.n340 commonsourceibias.n339 161.3
R6951 commonsourceibias.n338 commonsourceibias.n295 161.3
R6952 commonsourceibias.n337 commonsourceibias.n336 161.3
R6953 commonsourceibias.n334 commonsourceibias.n296 161.3
R6954 commonsourceibias.n333 commonsourceibias.n332 161.3
R6955 commonsourceibias.n331 commonsourceibias.n330 161.3
R6956 commonsourceibias.n329 commonsourceibias.n298 161.3
R6957 commonsourceibias.n328 commonsourceibias.n327 161.3
R6958 commonsourceibias.n326 commonsourceibias.n325 161.3
R6959 commonsourceibias.n324 commonsourceibias.n300 161.3
R6960 commonsourceibias.n323 commonsourceibias.n322 161.3
R6961 commonsourceibias.n321 commonsourceibias.n320 161.3
R6962 commonsourceibias.n319 commonsourceibias.n302 161.3
R6963 commonsourceibias.n317 commonsourceibias.n316 161.3
R6964 commonsourceibias.n315 commonsourceibias.n303 161.3
R6965 commonsourceibias.n314 commonsourceibias.n313 161.3
R6966 commonsourceibias.n311 commonsourceibias.n304 161.3
R6967 commonsourceibias.n310 commonsourceibias.n309 161.3
R6968 commonsourceibias.n308 commonsourceibias.n305 161.3
R6969 commonsourceibias.n218 commonsourceibias.n215 161.3
R6970 commonsourceibias.n220 commonsourceibias.n219 161.3
R6971 commonsourceibias.n221 commonsourceibias.n214 161.3
R6972 commonsourceibias.n224 commonsourceibias.n223 161.3
R6973 commonsourceibias.n225 commonsourceibias.n213 161.3
R6974 commonsourceibias.n227 commonsourceibias.n226 161.3
R6975 commonsourceibias.n229 commonsourceibias.n212 161.3
R6976 commonsourceibias.n231 commonsourceibias.n230 161.3
R6977 commonsourceibias.n233 commonsourceibias.n232 161.3
R6978 commonsourceibias.n234 commonsourceibias.n210 161.3
R6979 commonsourceibias.n236 commonsourceibias.n235 161.3
R6980 commonsourceibias.n238 commonsourceibias.n237 161.3
R6981 commonsourceibias.n239 commonsourceibias.n208 161.3
R6982 commonsourceibias.n241 commonsourceibias.n240 161.3
R6983 commonsourceibias.n243 commonsourceibias.n242 161.3
R6984 commonsourceibias.n244 commonsourceibias.n206 161.3
R6985 commonsourceibias.n247 commonsourceibias.n246 161.3
R6986 commonsourceibias.n248 commonsourceibias.n205 161.3
R6987 commonsourceibias.n250 commonsourceibias.n249 161.3
R6988 commonsourceibias.n252 commonsourceibias.n203 161.3
R6989 commonsourceibias.n254 commonsourceibias.n253 161.3
R6990 commonsourceibias.n255 commonsourceibias.n202 161.3
R6991 commonsourceibias.n257 commonsourceibias.n256 161.3
R6992 commonsourceibias.n258 commonsourceibias.n201 161.3
R6993 commonsourceibias.n261 commonsourceibias.n260 161.3
R6994 commonsourceibias.n262 commonsourceibias.n200 161.3
R6995 commonsourceibias.n264 commonsourceibias.n263 161.3
R6996 commonsourceibias.n266 commonsourceibias.n198 161.3
R6997 commonsourceibias.n268 commonsourceibias.n267 161.3
R6998 commonsourceibias.n269 commonsourceibias.n197 161.3
R6999 commonsourceibias.n271 commonsourceibias.n270 161.3
R7000 commonsourceibias.n272 commonsourceibias.n196 161.3
R7001 commonsourceibias.n275 commonsourceibias.n274 161.3
R7002 commonsourceibias.n276 commonsourceibias.n195 161.3
R7003 commonsourceibias.n278 commonsourceibias.n277 161.3
R7004 commonsourceibias.n280 commonsourceibias.n194 161.3
R7005 commonsourceibias.n519 commonsourceibias.n433 161.3
R7006 commonsourceibias.n517 commonsourceibias.n516 161.3
R7007 commonsourceibias.n515 commonsourceibias.n434 161.3
R7008 commonsourceibias.n514 commonsourceibias.n513 161.3
R7009 commonsourceibias.n511 commonsourceibias.n435 161.3
R7010 commonsourceibias.n510 commonsourceibias.n509 161.3
R7011 commonsourceibias.n508 commonsourceibias.n436 161.3
R7012 commonsourceibias.n507 commonsourceibias.n506 161.3
R7013 commonsourceibias.n504 commonsourceibias.n437 161.3
R7014 commonsourceibias.n502 commonsourceibias.n501 161.3
R7015 commonsourceibias.n500 commonsourceibias.n438 161.3
R7016 commonsourceibias.n499 commonsourceibias.n498 161.3
R7017 commonsourceibias.n496 commonsourceibias.n439 161.3
R7018 commonsourceibias.n495 commonsourceibias.n494 161.3
R7019 commonsourceibias.n493 commonsourceibias.n440 161.3
R7020 commonsourceibias.n492 commonsourceibias.n491 161.3
R7021 commonsourceibias.n489 commonsourceibias.n441 161.3
R7022 commonsourceibias.n487 commonsourceibias.n486 161.3
R7023 commonsourceibias.n485 commonsourceibias.n442 161.3
R7024 commonsourceibias.n484 commonsourceibias.n483 161.3
R7025 commonsourceibias.n481 commonsourceibias.n443 161.3
R7026 commonsourceibias.n480 commonsourceibias.n479 161.3
R7027 commonsourceibias.n478 commonsourceibias.n477 161.3
R7028 commonsourceibias.n476 commonsourceibias.n445 161.3
R7029 commonsourceibias.n475 commonsourceibias.n474 161.3
R7030 commonsourceibias.n473 commonsourceibias.n472 161.3
R7031 commonsourceibias.n471 commonsourceibias.n447 161.3
R7032 commonsourceibias.n470 commonsourceibias.n469 161.3
R7033 commonsourceibias.n468 commonsourceibias.n467 161.3
R7034 commonsourceibias.n466 commonsourceibias.n449 161.3
R7035 commonsourceibias.n464 commonsourceibias.n463 161.3
R7036 commonsourceibias.n462 commonsourceibias.n450 161.3
R7037 commonsourceibias.n461 commonsourceibias.n460 161.3
R7038 commonsourceibias.n458 commonsourceibias.n451 161.3
R7039 commonsourceibias.n457 commonsourceibias.n456 161.3
R7040 commonsourceibias.n455 commonsourceibias.n452 161.3
R7041 commonsourceibias.n425 commonsourceibias.n424 161.3
R7042 commonsourceibias.n422 commonsourceibias.n384 161.3
R7043 commonsourceibias.n421 commonsourceibias.n420 161.3
R7044 commonsourceibias.n419 commonsourceibias.n418 161.3
R7045 commonsourceibias.n417 commonsourceibias.n386 161.3
R7046 commonsourceibias.n416 commonsourceibias.n415 161.3
R7047 commonsourceibias.n414 commonsourceibias.n413 161.3
R7048 commonsourceibias.n412 commonsourceibias.n388 161.3
R7049 commonsourceibias.n411 commonsourceibias.n410 161.3
R7050 commonsourceibias.n409 commonsourceibias.n408 161.3
R7051 commonsourceibias.n407 commonsourceibias.n390 161.3
R7052 commonsourceibias.n405 commonsourceibias.n404 161.3
R7053 commonsourceibias.n403 commonsourceibias.n391 161.3
R7054 commonsourceibias.n402 commonsourceibias.n401 161.3
R7055 commonsourceibias.n399 commonsourceibias.n392 161.3
R7056 commonsourceibias.n398 commonsourceibias.n397 161.3
R7057 commonsourceibias.n396 commonsourceibias.n393 161.3
R7058 commonsourceibias.n531 commonsourceibias.n383 161.3
R7059 commonsourceibias.n565 commonsourceibias.n374 161.3
R7060 commonsourceibias.n563 commonsourceibias.n562 161.3
R7061 commonsourceibias.n561 commonsourceibias.n375 161.3
R7062 commonsourceibias.n560 commonsourceibias.n559 161.3
R7063 commonsourceibias.n557 commonsourceibias.n376 161.3
R7064 commonsourceibias.n556 commonsourceibias.n555 161.3
R7065 commonsourceibias.n554 commonsourceibias.n377 161.3
R7066 commonsourceibias.n553 commonsourceibias.n552 161.3
R7067 commonsourceibias.n550 commonsourceibias.n378 161.3
R7068 commonsourceibias.n548 commonsourceibias.n547 161.3
R7069 commonsourceibias.n546 commonsourceibias.n379 161.3
R7070 commonsourceibias.n545 commonsourceibias.n544 161.3
R7071 commonsourceibias.n542 commonsourceibias.n380 161.3
R7072 commonsourceibias.n541 commonsourceibias.n540 161.3
R7073 commonsourceibias.n539 commonsourceibias.n381 161.3
R7074 commonsourceibias.n538 commonsourceibias.n537 161.3
R7075 commonsourceibias.n535 commonsourceibias.n382 161.3
R7076 commonsourceibias.n533 commonsourceibias.n532 161.3
R7077 commonsourceibias.n744 commonsourceibias.n658 161.3
R7078 commonsourceibias.n742 commonsourceibias.n741 161.3
R7079 commonsourceibias.n740 commonsourceibias.n659 161.3
R7080 commonsourceibias.n739 commonsourceibias.n738 161.3
R7081 commonsourceibias.n736 commonsourceibias.n660 161.3
R7082 commonsourceibias.n735 commonsourceibias.n734 161.3
R7083 commonsourceibias.n733 commonsourceibias.n661 161.3
R7084 commonsourceibias.n732 commonsourceibias.n731 161.3
R7085 commonsourceibias.n729 commonsourceibias.n662 161.3
R7086 commonsourceibias.n727 commonsourceibias.n726 161.3
R7087 commonsourceibias.n725 commonsourceibias.n663 161.3
R7088 commonsourceibias.n724 commonsourceibias.n723 161.3
R7089 commonsourceibias.n721 commonsourceibias.n664 161.3
R7090 commonsourceibias.n720 commonsourceibias.n719 161.3
R7091 commonsourceibias.n718 commonsourceibias.n665 161.3
R7092 commonsourceibias.n717 commonsourceibias.n716 161.3
R7093 commonsourceibias.n714 commonsourceibias.n666 161.3
R7094 commonsourceibias.n712 commonsourceibias.n711 161.3
R7095 commonsourceibias.n710 commonsourceibias.n667 161.3
R7096 commonsourceibias.n709 commonsourceibias.n708 161.3
R7097 commonsourceibias.n706 commonsourceibias.n668 161.3
R7098 commonsourceibias.n705 commonsourceibias.n704 161.3
R7099 commonsourceibias.n703 commonsourceibias.n702 161.3
R7100 commonsourceibias.n701 commonsourceibias.n670 161.3
R7101 commonsourceibias.n700 commonsourceibias.n699 161.3
R7102 commonsourceibias.n698 commonsourceibias.n697 161.3
R7103 commonsourceibias.n696 commonsourceibias.n672 161.3
R7104 commonsourceibias.n695 commonsourceibias.n694 161.3
R7105 commonsourceibias.n693 commonsourceibias.n692 161.3
R7106 commonsourceibias.n691 commonsourceibias.n674 161.3
R7107 commonsourceibias.n689 commonsourceibias.n688 161.3
R7108 commonsourceibias.n687 commonsourceibias.n675 161.3
R7109 commonsourceibias.n686 commonsourceibias.n685 161.3
R7110 commonsourceibias.n683 commonsourceibias.n676 161.3
R7111 commonsourceibias.n682 commonsourceibias.n681 161.3
R7112 commonsourceibias.n680 commonsourceibias.n677 161.3
R7113 commonsourceibias.n654 commonsourceibias.n568 161.3
R7114 commonsourceibias.n652 commonsourceibias.n651 161.3
R7115 commonsourceibias.n650 commonsourceibias.n569 161.3
R7116 commonsourceibias.n649 commonsourceibias.n648 161.3
R7117 commonsourceibias.n646 commonsourceibias.n570 161.3
R7118 commonsourceibias.n645 commonsourceibias.n644 161.3
R7119 commonsourceibias.n643 commonsourceibias.n571 161.3
R7120 commonsourceibias.n642 commonsourceibias.n641 161.3
R7121 commonsourceibias.n639 commonsourceibias.n572 161.3
R7122 commonsourceibias.n637 commonsourceibias.n636 161.3
R7123 commonsourceibias.n635 commonsourceibias.n573 161.3
R7124 commonsourceibias.n634 commonsourceibias.n633 161.3
R7125 commonsourceibias.n631 commonsourceibias.n574 161.3
R7126 commonsourceibias.n630 commonsourceibias.n629 161.3
R7127 commonsourceibias.n628 commonsourceibias.n575 161.3
R7128 commonsourceibias.n627 commonsourceibias.n626 161.3
R7129 commonsourceibias.n624 commonsourceibias.n576 161.3
R7130 commonsourceibias.n622 commonsourceibias.n621 161.3
R7131 commonsourceibias.n620 commonsourceibias.n577 161.3
R7132 commonsourceibias.n619 commonsourceibias.n618 161.3
R7133 commonsourceibias.n616 commonsourceibias.n578 161.3
R7134 commonsourceibias.n615 commonsourceibias.n614 161.3
R7135 commonsourceibias.n613 commonsourceibias.n612 161.3
R7136 commonsourceibias.n611 commonsourceibias.n580 161.3
R7137 commonsourceibias.n610 commonsourceibias.n609 161.3
R7138 commonsourceibias.n608 commonsourceibias.n607 161.3
R7139 commonsourceibias.n606 commonsourceibias.n582 161.3
R7140 commonsourceibias.n605 commonsourceibias.n604 161.3
R7141 commonsourceibias.n603 commonsourceibias.n602 161.3
R7142 commonsourceibias.n601 commonsourceibias.n584 161.3
R7143 commonsourceibias.n599 commonsourceibias.n598 161.3
R7144 commonsourceibias.n597 commonsourceibias.n585 161.3
R7145 commonsourceibias.n596 commonsourceibias.n595 161.3
R7146 commonsourceibias.n593 commonsourceibias.n586 161.3
R7147 commonsourceibias.n592 commonsourceibias.n591 161.3
R7148 commonsourceibias.n590 commonsourceibias.n587 161.3
R7149 commonsourceibias.n111 commonsourceibias.n109 81.5057
R7150 commonsourceibias.n428 commonsourceibias.n426 81.5057
R7151 commonsourceibias.n111 commonsourceibias.n110 80.9324
R7152 commonsourceibias.n113 commonsourceibias.n112 80.9324
R7153 commonsourceibias.n115 commonsourceibias.n114 80.9324
R7154 commonsourceibias.n108 commonsourceibias.n107 80.9324
R7155 commonsourceibias.n106 commonsourceibias.n105 80.9324
R7156 commonsourceibias.n104 commonsourceibias.n103 80.9324
R7157 commonsourceibias.n102 commonsourceibias.n101 80.9324
R7158 commonsourceibias.n523 commonsourceibias.n522 80.9324
R7159 commonsourceibias.n525 commonsourceibias.n524 80.9324
R7160 commonsourceibias.n527 commonsourceibias.n526 80.9324
R7161 commonsourceibias.n529 commonsourceibias.n528 80.9324
R7162 commonsourceibias.n432 commonsourceibias.n431 80.9324
R7163 commonsourceibias.n430 commonsourceibias.n429 80.9324
R7164 commonsourceibias.n428 commonsourceibias.n427 80.9324
R7165 commonsourceibias.n100 commonsourceibias.n99 80.6037
R7166 commonsourceibias.n193 commonsourceibias.n192 80.6037
R7167 commonsourceibias.n372 commonsourceibias.n371 80.6037
R7168 commonsourceibias.n282 commonsourceibias.n281 80.6037
R7169 commonsourceibias.n521 commonsourceibias.n520 80.6037
R7170 commonsourceibias.n567 commonsourceibias.n566 80.6037
R7171 commonsourceibias.n746 commonsourceibias.n745 80.6037
R7172 commonsourceibias.n656 commonsourceibias.n655 80.6037
R7173 commonsourceibias.n85 commonsourceibias.n84 56.5617
R7174 commonsourceibias.n71 commonsourceibias.n70 56.5617
R7175 commonsourceibias.n62 commonsourceibias.n61 56.5617
R7176 commonsourceibias.n48 commonsourceibias.n47 56.5617
R7177 commonsourceibias.n178 commonsourceibias.n177 56.5617
R7178 commonsourceibias.n164 commonsourceibias.n163 56.5617
R7179 commonsourceibias.n155 commonsourceibias.n154 56.5617
R7180 commonsourceibias.n141 commonsourceibias.n140 56.5617
R7181 commonsourceibias.n320 commonsourceibias.n319 56.5617
R7182 commonsourceibias.n334 commonsourceibias.n333 56.5617
R7183 commonsourceibias.n343 commonsourceibias.n342 56.5617
R7184 commonsourceibias.n357 commonsourceibias.n356 56.5617
R7185 commonsourceibias.n267 commonsourceibias.n266 56.5617
R7186 commonsourceibias.n253 commonsourceibias.n252 56.5617
R7187 commonsourceibias.n244 commonsourceibias.n243 56.5617
R7188 commonsourceibias.n230 commonsourceibias.n229 56.5617
R7189 commonsourceibias.n467 commonsourceibias.n466 56.5617
R7190 commonsourceibias.n481 commonsourceibias.n480 56.5617
R7191 commonsourceibias.n491 commonsourceibias.n489 56.5617
R7192 commonsourceibias.n506 commonsourceibias.n504 56.5617
R7193 commonsourceibias.n552 commonsourceibias.n550 56.5617
R7194 commonsourceibias.n537 commonsourceibias.n535 56.5617
R7195 commonsourceibias.n408 commonsourceibias.n407 56.5617
R7196 commonsourceibias.n422 commonsourceibias.n421 56.5617
R7197 commonsourceibias.n692 commonsourceibias.n691 56.5617
R7198 commonsourceibias.n706 commonsourceibias.n705 56.5617
R7199 commonsourceibias.n716 commonsourceibias.n714 56.5617
R7200 commonsourceibias.n731 commonsourceibias.n729 56.5617
R7201 commonsourceibias.n602 commonsourceibias.n601 56.5617
R7202 commonsourceibias.n616 commonsourceibias.n615 56.5617
R7203 commonsourceibias.n626 commonsourceibias.n624 56.5617
R7204 commonsourceibias.n641 commonsourceibias.n639 56.5617
R7205 commonsourceibias.n76 commonsourceibias.n75 56.0773
R7206 commonsourceibias.n57 commonsourceibias.n56 56.0773
R7207 commonsourceibias.n169 commonsourceibias.n168 56.0773
R7208 commonsourceibias.n150 commonsourceibias.n149 56.0773
R7209 commonsourceibias.n329 commonsourceibias.n328 56.0773
R7210 commonsourceibias.n348 commonsourceibias.n347 56.0773
R7211 commonsourceibias.n258 commonsourceibias.n257 56.0773
R7212 commonsourceibias.n239 commonsourceibias.n238 56.0773
R7213 commonsourceibias.n476 commonsourceibias.n475 56.0773
R7214 commonsourceibias.n496 commonsourceibias.n495 56.0773
R7215 commonsourceibias.n542 commonsourceibias.n541 56.0773
R7216 commonsourceibias.n417 commonsourceibias.n416 56.0773
R7217 commonsourceibias.n701 commonsourceibias.n700 56.0773
R7218 commonsourceibias.n721 commonsourceibias.n720 56.0773
R7219 commonsourceibias.n611 commonsourceibias.n610 56.0773
R7220 commonsourceibias.n631 commonsourceibias.n630 56.0773
R7221 commonsourceibias.n99 commonsourceibias.n98 55.3321
R7222 commonsourceibias.n192 commonsourceibias.n191 55.3321
R7223 commonsourceibias.n371 commonsourceibias.n370 55.3321
R7224 commonsourceibias.n281 commonsourceibias.n280 55.3321
R7225 commonsourceibias.n520 commonsourceibias.n519 55.3321
R7226 commonsourceibias.n566 commonsourceibias.n565 55.3321
R7227 commonsourceibias.n745 commonsourceibias.n744 55.3321
R7228 commonsourceibias.n655 commonsourceibias.n654 55.3321
R7229 commonsourceibias.n90 commonsourceibias.n89 55.1086
R7230 commonsourceibias.n41 commonsourceibias.n31 55.1086
R7231 commonsourceibias.n183 commonsourceibias.n182 55.1086
R7232 commonsourceibias.n134 commonsourceibias.n124 55.1086
R7233 commonsourceibias.n313 commonsourceibias.n303 55.1086
R7234 commonsourceibias.n362 commonsourceibias.n361 55.1086
R7235 commonsourceibias.n272 commonsourceibias.n271 55.1086
R7236 commonsourceibias.n223 commonsourceibias.n213 55.1086
R7237 commonsourceibias.n460 commonsourceibias.n450 55.1086
R7238 commonsourceibias.n511 commonsourceibias.n510 55.1086
R7239 commonsourceibias.n557 commonsourceibias.n556 55.1086
R7240 commonsourceibias.n401 commonsourceibias.n391 55.1086
R7241 commonsourceibias.n685 commonsourceibias.n675 55.1086
R7242 commonsourceibias.n736 commonsourceibias.n735 55.1086
R7243 commonsourceibias.n595 commonsourceibias.n585 55.1086
R7244 commonsourceibias.n646 commonsourceibias.n645 55.1086
R7245 commonsourceibias.n35 commonsourceibias.n34 47.4592
R7246 commonsourceibias.n128 commonsourceibias.n127 47.4592
R7247 commonsourceibias.n307 commonsourceibias.n306 47.4592
R7248 commonsourceibias.n217 commonsourceibias.n216 47.4592
R7249 commonsourceibias.n454 commonsourceibias.n453 47.4592
R7250 commonsourceibias.n395 commonsourceibias.n394 47.4592
R7251 commonsourceibias.n679 commonsourceibias.n678 47.4592
R7252 commonsourceibias.n589 commonsourceibias.n588 47.4592
R7253 commonsourceibias.n308 commonsourceibias.n307 44.0436
R7254 commonsourceibias.n455 commonsourceibias.n454 44.0436
R7255 commonsourceibias.n396 commonsourceibias.n395 44.0436
R7256 commonsourceibias.n680 commonsourceibias.n679 44.0436
R7257 commonsourceibias.n590 commonsourceibias.n589 44.0436
R7258 commonsourceibias.n36 commonsourceibias.n35 44.0436
R7259 commonsourceibias.n129 commonsourceibias.n128 44.0436
R7260 commonsourceibias.n218 commonsourceibias.n217 44.0436
R7261 commonsourceibias.n92 commonsourceibias.n13 42.5146
R7262 commonsourceibias.n39 commonsourceibias.n38 42.5146
R7263 commonsourceibias.n185 commonsourceibias.n1 42.5146
R7264 commonsourceibias.n132 commonsourceibias.n131 42.5146
R7265 commonsourceibias.n311 commonsourceibias.n310 42.5146
R7266 commonsourceibias.n364 commonsourceibias.n285 42.5146
R7267 commonsourceibias.n274 commonsourceibias.n195 42.5146
R7268 commonsourceibias.n221 commonsourceibias.n220 42.5146
R7269 commonsourceibias.n458 commonsourceibias.n457 42.5146
R7270 commonsourceibias.n513 commonsourceibias.n434 42.5146
R7271 commonsourceibias.n559 commonsourceibias.n375 42.5146
R7272 commonsourceibias.n399 commonsourceibias.n398 42.5146
R7273 commonsourceibias.n683 commonsourceibias.n682 42.5146
R7274 commonsourceibias.n738 commonsourceibias.n659 42.5146
R7275 commonsourceibias.n593 commonsourceibias.n592 42.5146
R7276 commonsourceibias.n648 commonsourceibias.n569 42.5146
R7277 commonsourceibias.n78 commonsourceibias.n18 41.5458
R7278 commonsourceibias.n53 commonsourceibias.n52 41.5458
R7279 commonsourceibias.n171 commonsourceibias.n6 41.5458
R7280 commonsourceibias.n146 commonsourceibias.n145 41.5458
R7281 commonsourceibias.n325 commonsourceibias.n324 41.5458
R7282 commonsourceibias.n350 commonsourceibias.n290 41.5458
R7283 commonsourceibias.n260 commonsourceibias.n200 41.5458
R7284 commonsourceibias.n235 commonsourceibias.n234 41.5458
R7285 commonsourceibias.n472 commonsourceibias.n471 41.5458
R7286 commonsourceibias.n498 commonsourceibias.n438 41.5458
R7287 commonsourceibias.n544 commonsourceibias.n379 41.5458
R7288 commonsourceibias.n413 commonsourceibias.n412 41.5458
R7289 commonsourceibias.n697 commonsourceibias.n696 41.5458
R7290 commonsourceibias.n723 commonsourceibias.n663 41.5458
R7291 commonsourceibias.n607 commonsourceibias.n606 41.5458
R7292 commonsourceibias.n633 commonsourceibias.n573 41.5458
R7293 commonsourceibias.n68 commonsourceibias.n23 40.577
R7294 commonsourceibias.n64 commonsourceibias.n23 40.577
R7295 commonsourceibias.n161 commonsourceibias.n11 40.577
R7296 commonsourceibias.n157 commonsourceibias.n11 40.577
R7297 commonsourceibias.n336 commonsourceibias.n295 40.577
R7298 commonsourceibias.n340 commonsourceibias.n295 40.577
R7299 commonsourceibias.n250 commonsourceibias.n205 40.577
R7300 commonsourceibias.n246 commonsourceibias.n205 40.577
R7301 commonsourceibias.n483 commonsourceibias.n442 40.577
R7302 commonsourceibias.n487 commonsourceibias.n442 40.577
R7303 commonsourceibias.n533 commonsourceibias.n383 40.577
R7304 commonsourceibias.n424 commonsourceibias.n383 40.577
R7305 commonsourceibias.n708 commonsourceibias.n667 40.577
R7306 commonsourceibias.n712 commonsourceibias.n667 40.577
R7307 commonsourceibias.n618 commonsourceibias.n577 40.577
R7308 commonsourceibias.n622 commonsourceibias.n577 40.577
R7309 commonsourceibias.n82 commonsourceibias.n18 39.6083
R7310 commonsourceibias.n52 commonsourceibias.n51 39.6083
R7311 commonsourceibias.n175 commonsourceibias.n6 39.6083
R7312 commonsourceibias.n145 commonsourceibias.n144 39.6083
R7313 commonsourceibias.n324 commonsourceibias.n323 39.6083
R7314 commonsourceibias.n354 commonsourceibias.n290 39.6083
R7315 commonsourceibias.n264 commonsourceibias.n200 39.6083
R7316 commonsourceibias.n234 commonsourceibias.n233 39.6083
R7317 commonsourceibias.n471 commonsourceibias.n470 39.6083
R7318 commonsourceibias.n502 commonsourceibias.n438 39.6083
R7319 commonsourceibias.n548 commonsourceibias.n379 39.6083
R7320 commonsourceibias.n412 commonsourceibias.n411 39.6083
R7321 commonsourceibias.n696 commonsourceibias.n695 39.6083
R7322 commonsourceibias.n727 commonsourceibias.n663 39.6083
R7323 commonsourceibias.n606 commonsourceibias.n605 39.6083
R7324 commonsourceibias.n637 commonsourceibias.n573 39.6083
R7325 commonsourceibias.n96 commonsourceibias.n13 38.6395
R7326 commonsourceibias.n38 commonsourceibias.n33 38.6395
R7327 commonsourceibias.n189 commonsourceibias.n1 38.6395
R7328 commonsourceibias.n131 commonsourceibias.n126 38.6395
R7329 commonsourceibias.n310 commonsourceibias.n305 38.6395
R7330 commonsourceibias.n368 commonsourceibias.n285 38.6395
R7331 commonsourceibias.n278 commonsourceibias.n195 38.6395
R7332 commonsourceibias.n220 commonsourceibias.n215 38.6395
R7333 commonsourceibias.n457 commonsourceibias.n452 38.6395
R7334 commonsourceibias.n517 commonsourceibias.n434 38.6395
R7335 commonsourceibias.n563 commonsourceibias.n375 38.6395
R7336 commonsourceibias.n398 commonsourceibias.n393 38.6395
R7337 commonsourceibias.n682 commonsourceibias.n677 38.6395
R7338 commonsourceibias.n742 commonsourceibias.n659 38.6395
R7339 commonsourceibias.n592 commonsourceibias.n587 38.6395
R7340 commonsourceibias.n652 commonsourceibias.n569 38.6395
R7341 commonsourceibias.n89 commonsourceibias.n15 26.0455
R7342 commonsourceibias.n45 commonsourceibias.n31 26.0455
R7343 commonsourceibias.n182 commonsourceibias.n3 26.0455
R7344 commonsourceibias.n138 commonsourceibias.n124 26.0455
R7345 commonsourceibias.n317 commonsourceibias.n303 26.0455
R7346 commonsourceibias.n361 commonsourceibias.n287 26.0455
R7347 commonsourceibias.n271 commonsourceibias.n197 26.0455
R7348 commonsourceibias.n227 commonsourceibias.n213 26.0455
R7349 commonsourceibias.n464 commonsourceibias.n450 26.0455
R7350 commonsourceibias.n510 commonsourceibias.n436 26.0455
R7351 commonsourceibias.n556 commonsourceibias.n377 26.0455
R7352 commonsourceibias.n405 commonsourceibias.n391 26.0455
R7353 commonsourceibias.n689 commonsourceibias.n675 26.0455
R7354 commonsourceibias.n735 commonsourceibias.n661 26.0455
R7355 commonsourceibias.n599 commonsourceibias.n585 26.0455
R7356 commonsourceibias.n645 commonsourceibias.n571 26.0455
R7357 commonsourceibias.n75 commonsourceibias.n20 25.0767
R7358 commonsourceibias.n58 commonsourceibias.n57 25.0767
R7359 commonsourceibias.n168 commonsourceibias.n8 25.0767
R7360 commonsourceibias.n151 commonsourceibias.n150 25.0767
R7361 commonsourceibias.n330 commonsourceibias.n329 25.0767
R7362 commonsourceibias.n347 commonsourceibias.n292 25.0767
R7363 commonsourceibias.n257 commonsourceibias.n202 25.0767
R7364 commonsourceibias.n240 commonsourceibias.n239 25.0767
R7365 commonsourceibias.n477 commonsourceibias.n476 25.0767
R7366 commonsourceibias.n495 commonsourceibias.n440 25.0767
R7367 commonsourceibias.n541 commonsourceibias.n381 25.0767
R7368 commonsourceibias.n418 commonsourceibias.n417 25.0767
R7369 commonsourceibias.n702 commonsourceibias.n701 25.0767
R7370 commonsourceibias.n720 commonsourceibias.n665 25.0767
R7371 commonsourceibias.n612 commonsourceibias.n611 25.0767
R7372 commonsourceibias.n630 commonsourceibias.n575 25.0767
R7373 commonsourceibias.n71 commonsourceibias.n22 24.3464
R7374 commonsourceibias.n61 commonsourceibias.n25 24.3464
R7375 commonsourceibias.n164 commonsourceibias.n10 24.3464
R7376 commonsourceibias.n154 commonsourceibias.n118 24.3464
R7377 commonsourceibias.n333 commonsourceibias.n297 24.3464
R7378 commonsourceibias.n343 commonsourceibias.n294 24.3464
R7379 commonsourceibias.n253 commonsourceibias.n204 24.3464
R7380 commonsourceibias.n243 commonsourceibias.n207 24.3464
R7381 commonsourceibias.n480 commonsourceibias.n444 24.3464
R7382 commonsourceibias.n491 commonsourceibias.n490 24.3464
R7383 commonsourceibias.n537 commonsourceibias.n536 24.3464
R7384 commonsourceibias.n421 commonsourceibias.n385 24.3464
R7385 commonsourceibias.n705 commonsourceibias.n669 24.3464
R7386 commonsourceibias.n716 commonsourceibias.n715 24.3464
R7387 commonsourceibias.n615 commonsourceibias.n579 24.3464
R7388 commonsourceibias.n626 commonsourceibias.n625 24.3464
R7389 commonsourceibias.n85 commonsourceibias.n17 23.8546
R7390 commonsourceibias.n47 commonsourceibias.n46 23.8546
R7391 commonsourceibias.n178 commonsourceibias.n5 23.8546
R7392 commonsourceibias.n140 commonsourceibias.n139 23.8546
R7393 commonsourceibias.n319 commonsourceibias.n318 23.8546
R7394 commonsourceibias.n357 commonsourceibias.n289 23.8546
R7395 commonsourceibias.n267 commonsourceibias.n199 23.8546
R7396 commonsourceibias.n229 commonsourceibias.n228 23.8546
R7397 commonsourceibias.n466 commonsourceibias.n465 23.8546
R7398 commonsourceibias.n506 commonsourceibias.n505 23.8546
R7399 commonsourceibias.n552 commonsourceibias.n551 23.8546
R7400 commonsourceibias.n407 commonsourceibias.n406 23.8546
R7401 commonsourceibias.n691 commonsourceibias.n690 23.8546
R7402 commonsourceibias.n731 commonsourceibias.n730 23.8546
R7403 commonsourceibias.n601 commonsourceibias.n600 23.8546
R7404 commonsourceibias.n641 commonsourceibias.n640 23.8546
R7405 commonsourceibias.n98 commonsourceibias.n97 17.4607
R7406 commonsourceibias.n191 commonsourceibias.n190 17.4607
R7407 commonsourceibias.n370 commonsourceibias.n369 17.4607
R7408 commonsourceibias.n280 commonsourceibias.n279 17.4607
R7409 commonsourceibias.n519 commonsourceibias.n518 17.4607
R7410 commonsourceibias.n565 commonsourceibias.n564 17.4607
R7411 commonsourceibias.n744 commonsourceibias.n743 17.4607
R7412 commonsourceibias.n654 commonsourceibias.n653 17.4607
R7413 commonsourceibias.n84 commonsourceibias.n83 16.9689
R7414 commonsourceibias.n48 commonsourceibias.n29 16.9689
R7415 commonsourceibias.n177 commonsourceibias.n176 16.9689
R7416 commonsourceibias.n141 commonsourceibias.n122 16.9689
R7417 commonsourceibias.n320 commonsourceibias.n301 16.9689
R7418 commonsourceibias.n356 commonsourceibias.n355 16.9689
R7419 commonsourceibias.n266 commonsourceibias.n265 16.9689
R7420 commonsourceibias.n230 commonsourceibias.n211 16.9689
R7421 commonsourceibias.n467 commonsourceibias.n448 16.9689
R7422 commonsourceibias.n504 commonsourceibias.n503 16.9689
R7423 commonsourceibias.n550 commonsourceibias.n549 16.9689
R7424 commonsourceibias.n408 commonsourceibias.n389 16.9689
R7425 commonsourceibias.n692 commonsourceibias.n673 16.9689
R7426 commonsourceibias.n729 commonsourceibias.n728 16.9689
R7427 commonsourceibias.n602 commonsourceibias.n583 16.9689
R7428 commonsourceibias.n639 commonsourceibias.n638 16.9689
R7429 commonsourceibias.n70 commonsourceibias.n69 16.477
R7430 commonsourceibias.n63 commonsourceibias.n62 16.477
R7431 commonsourceibias.n163 commonsourceibias.n162 16.477
R7432 commonsourceibias.n156 commonsourceibias.n155 16.477
R7433 commonsourceibias.n335 commonsourceibias.n334 16.477
R7434 commonsourceibias.n342 commonsourceibias.n341 16.477
R7435 commonsourceibias.n252 commonsourceibias.n251 16.477
R7436 commonsourceibias.n245 commonsourceibias.n244 16.477
R7437 commonsourceibias.n482 commonsourceibias.n481 16.477
R7438 commonsourceibias.n489 commonsourceibias.n488 16.477
R7439 commonsourceibias.n535 commonsourceibias.n534 16.477
R7440 commonsourceibias.n423 commonsourceibias.n422 16.477
R7441 commonsourceibias.n707 commonsourceibias.n706 16.477
R7442 commonsourceibias.n714 commonsourceibias.n713 16.477
R7443 commonsourceibias.n617 commonsourceibias.n616 16.477
R7444 commonsourceibias.n624 commonsourceibias.n623 16.477
R7445 commonsourceibias.n77 commonsourceibias.n76 15.9852
R7446 commonsourceibias.n56 commonsourceibias.n27 15.9852
R7447 commonsourceibias.n170 commonsourceibias.n169 15.9852
R7448 commonsourceibias.n149 commonsourceibias.n120 15.9852
R7449 commonsourceibias.n328 commonsourceibias.n299 15.9852
R7450 commonsourceibias.n349 commonsourceibias.n348 15.9852
R7451 commonsourceibias.n259 commonsourceibias.n258 15.9852
R7452 commonsourceibias.n238 commonsourceibias.n209 15.9852
R7453 commonsourceibias.n475 commonsourceibias.n446 15.9852
R7454 commonsourceibias.n497 commonsourceibias.n496 15.9852
R7455 commonsourceibias.n543 commonsourceibias.n542 15.9852
R7456 commonsourceibias.n416 commonsourceibias.n387 15.9852
R7457 commonsourceibias.n700 commonsourceibias.n671 15.9852
R7458 commonsourceibias.n722 commonsourceibias.n721 15.9852
R7459 commonsourceibias.n610 commonsourceibias.n581 15.9852
R7460 commonsourceibias.n632 commonsourceibias.n631 15.9852
R7461 commonsourceibias.n91 commonsourceibias.n90 15.4934
R7462 commonsourceibias.n41 commonsourceibias.n40 15.4934
R7463 commonsourceibias.n184 commonsourceibias.n183 15.4934
R7464 commonsourceibias.n134 commonsourceibias.n133 15.4934
R7465 commonsourceibias.n313 commonsourceibias.n312 15.4934
R7466 commonsourceibias.n363 commonsourceibias.n362 15.4934
R7467 commonsourceibias.n273 commonsourceibias.n272 15.4934
R7468 commonsourceibias.n223 commonsourceibias.n222 15.4934
R7469 commonsourceibias.n460 commonsourceibias.n459 15.4934
R7470 commonsourceibias.n512 commonsourceibias.n511 15.4934
R7471 commonsourceibias.n558 commonsourceibias.n557 15.4934
R7472 commonsourceibias.n401 commonsourceibias.n400 15.4934
R7473 commonsourceibias.n685 commonsourceibias.n684 15.4934
R7474 commonsourceibias.n737 commonsourceibias.n736 15.4934
R7475 commonsourceibias.n595 commonsourceibias.n594 15.4934
R7476 commonsourceibias.n647 commonsourceibias.n646 15.4934
R7477 commonsourceibias.n102 commonsourceibias.n100 13.2663
R7478 commonsourceibias.n523 commonsourceibias.n521 13.2663
R7479 commonsourceibias.n748 commonsourceibias.n373 10.122
R7480 commonsourceibias.n159 commonsourceibias.n116 9.50363
R7481 commonsourceibias.n531 commonsourceibias.n530 9.50363
R7482 commonsourceibias.n92 commonsourceibias.n91 9.09948
R7483 commonsourceibias.n40 commonsourceibias.n39 9.09948
R7484 commonsourceibias.n185 commonsourceibias.n184 9.09948
R7485 commonsourceibias.n133 commonsourceibias.n132 9.09948
R7486 commonsourceibias.n312 commonsourceibias.n311 9.09948
R7487 commonsourceibias.n364 commonsourceibias.n363 9.09948
R7488 commonsourceibias.n274 commonsourceibias.n273 9.09948
R7489 commonsourceibias.n222 commonsourceibias.n221 9.09948
R7490 commonsourceibias.n459 commonsourceibias.n458 9.09948
R7491 commonsourceibias.n513 commonsourceibias.n512 9.09948
R7492 commonsourceibias.n559 commonsourceibias.n558 9.09948
R7493 commonsourceibias.n400 commonsourceibias.n399 9.09948
R7494 commonsourceibias.n684 commonsourceibias.n683 9.09948
R7495 commonsourceibias.n738 commonsourceibias.n737 9.09948
R7496 commonsourceibias.n594 commonsourceibias.n593 9.09948
R7497 commonsourceibias.n648 commonsourceibias.n647 9.09948
R7498 commonsourceibias.n283 commonsourceibias.n193 8.79451
R7499 commonsourceibias.n657 commonsourceibias.n567 8.79451
R7500 commonsourceibias.n78 commonsourceibias.n77 8.60764
R7501 commonsourceibias.n53 commonsourceibias.n27 8.60764
R7502 commonsourceibias.n171 commonsourceibias.n170 8.60764
R7503 commonsourceibias.n146 commonsourceibias.n120 8.60764
R7504 commonsourceibias.n325 commonsourceibias.n299 8.60764
R7505 commonsourceibias.n350 commonsourceibias.n349 8.60764
R7506 commonsourceibias.n260 commonsourceibias.n259 8.60764
R7507 commonsourceibias.n235 commonsourceibias.n209 8.60764
R7508 commonsourceibias.n472 commonsourceibias.n446 8.60764
R7509 commonsourceibias.n498 commonsourceibias.n497 8.60764
R7510 commonsourceibias.n544 commonsourceibias.n543 8.60764
R7511 commonsourceibias.n413 commonsourceibias.n387 8.60764
R7512 commonsourceibias.n697 commonsourceibias.n671 8.60764
R7513 commonsourceibias.n723 commonsourceibias.n722 8.60764
R7514 commonsourceibias.n607 commonsourceibias.n581 8.60764
R7515 commonsourceibias.n633 commonsourceibias.n632 8.60764
R7516 commonsourceibias.n748 commonsourceibias.n747 8.46921
R7517 commonsourceibias.n69 commonsourceibias.n68 8.11581
R7518 commonsourceibias.n64 commonsourceibias.n63 8.11581
R7519 commonsourceibias.n162 commonsourceibias.n161 8.11581
R7520 commonsourceibias.n157 commonsourceibias.n156 8.11581
R7521 commonsourceibias.n336 commonsourceibias.n335 8.11581
R7522 commonsourceibias.n341 commonsourceibias.n340 8.11581
R7523 commonsourceibias.n251 commonsourceibias.n250 8.11581
R7524 commonsourceibias.n246 commonsourceibias.n245 8.11581
R7525 commonsourceibias.n483 commonsourceibias.n482 8.11581
R7526 commonsourceibias.n488 commonsourceibias.n487 8.11581
R7527 commonsourceibias.n534 commonsourceibias.n533 8.11581
R7528 commonsourceibias.n424 commonsourceibias.n423 8.11581
R7529 commonsourceibias.n708 commonsourceibias.n707 8.11581
R7530 commonsourceibias.n713 commonsourceibias.n712 8.11581
R7531 commonsourceibias.n618 commonsourceibias.n617 8.11581
R7532 commonsourceibias.n623 commonsourceibias.n622 8.11581
R7533 commonsourceibias.n83 commonsourceibias.n82 7.62397
R7534 commonsourceibias.n51 commonsourceibias.n29 7.62397
R7535 commonsourceibias.n176 commonsourceibias.n175 7.62397
R7536 commonsourceibias.n144 commonsourceibias.n122 7.62397
R7537 commonsourceibias.n323 commonsourceibias.n301 7.62397
R7538 commonsourceibias.n355 commonsourceibias.n354 7.62397
R7539 commonsourceibias.n265 commonsourceibias.n264 7.62397
R7540 commonsourceibias.n233 commonsourceibias.n211 7.62397
R7541 commonsourceibias.n470 commonsourceibias.n448 7.62397
R7542 commonsourceibias.n503 commonsourceibias.n502 7.62397
R7543 commonsourceibias.n549 commonsourceibias.n548 7.62397
R7544 commonsourceibias.n411 commonsourceibias.n389 7.62397
R7545 commonsourceibias.n695 commonsourceibias.n673 7.62397
R7546 commonsourceibias.n728 commonsourceibias.n727 7.62397
R7547 commonsourceibias.n605 commonsourceibias.n583 7.62397
R7548 commonsourceibias.n638 commonsourceibias.n637 7.62397
R7549 commonsourceibias.n97 commonsourceibias.n96 7.13213
R7550 commonsourceibias.n34 commonsourceibias.n33 7.13213
R7551 commonsourceibias.n190 commonsourceibias.n189 7.13213
R7552 commonsourceibias.n127 commonsourceibias.n126 7.13213
R7553 commonsourceibias.n306 commonsourceibias.n305 7.13213
R7554 commonsourceibias.n369 commonsourceibias.n368 7.13213
R7555 commonsourceibias.n279 commonsourceibias.n278 7.13213
R7556 commonsourceibias.n216 commonsourceibias.n215 7.13213
R7557 commonsourceibias.n453 commonsourceibias.n452 7.13213
R7558 commonsourceibias.n518 commonsourceibias.n517 7.13213
R7559 commonsourceibias.n564 commonsourceibias.n563 7.13213
R7560 commonsourceibias.n394 commonsourceibias.n393 7.13213
R7561 commonsourceibias.n678 commonsourceibias.n677 7.13213
R7562 commonsourceibias.n743 commonsourceibias.n742 7.13213
R7563 commonsourceibias.n588 commonsourceibias.n587 7.13213
R7564 commonsourceibias.n653 commonsourceibias.n652 7.13213
R7565 commonsourceibias.n373 commonsourceibias.n372 5.06534
R7566 commonsourceibias.n283 commonsourceibias.n282 5.06534
R7567 commonsourceibias.n747 commonsourceibias.n746 5.06534
R7568 commonsourceibias.n657 commonsourceibias.n656 5.06534
R7569 commonsourceibias commonsourceibias.n748 4.04308
R7570 commonsourceibias.n373 commonsourceibias.n283 3.72967
R7571 commonsourceibias.n747 commonsourceibias.n657 3.72967
R7572 commonsourceibias.n109 commonsourceibias.t51 2.82907
R7573 commonsourceibias.n109 commonsourceibias.t17 2.82907
R7574 commonsourceibias.n110 commonsourceibias.t9 2.82907
R7575 commonsourceibias.n110 commonsourceibias.t11 2.82907
R7576 commonsourceibias.n112 commonsourceibias.t3 2.82907
R7577 commonsourceibias.n112 commonsourceibias.t57 2.82907
R7578 commonsourceibias.n114 commonsourceibias.t23 2.82907
R7579 commonsourceibias.n114 commonsourceibias.t43 2.82907
R7580 commonsourceibias.n107 commonsourceibias.t53 2.82907
R7581 commonsourceibias.n107 commonsourceibias.t33 2.82907
R7582 commonsourceibias.n105 commonsourceibias.t29 2.82907
R7583 commonsourceibias.n105 commonsourceibias.t25 2.82907
R7584 commonsourceibias.n103 commonsourceibias.t31 2.82907
R7585 commonsourceibias.n103 commonsourceibias.t7 2.82907
R7586 commonsourceibias.n101 commonsourceibias.t21 2.82907
R7587 commonsourceibias.n101 commonsourceibias.t49 2.82907
R7588 commonsourceibias.n522 commonsourceibias.t45 2.82907
R7589 commonsourceibias.n522 commonsourceibias.t59 2.82907
R7590 commonsourceibias.n524 commonsourceibias.t55 2.82907
R7591 commonsourceibias.n524 commonsourceibias.t13 2.82907
R7592 commonsourceibias.n526 commonsourceibias.t37 2.82907
R7593 commonsourceibias.n526 commonsourceibias.t27 2.82907
R7594 commonsourceibias.n528 commonsourceibias.t5 2.82907
R7595 commonsourceibias.n528 commonsourceibias.t47 2.82907
R7596 commonsourceibias.n431 commonsourceibias.t61 2.82907
R7597 commonsourceibias.n431 commonsourceibias.t35 2.82907
R7598 commonsourceibias.n429 commonsourceibias.t63 2.82907
R7599 commonsourceibias.n429 commonsourceibias.t41 2.82907
R7600 commonsourceibias.n427 commonsourceibias.t39 2.82907
R7601 commonsourceibias.n427 commonsourceibias.t19 2.82907
R7602 commonsourceibias.n426 commonsourceibias.t15 2.82907
R7603 commonsourceibias.n426 commonsourceibias.t1 2.82907
R7604 commonsourceibias.n17 commonsourceibias.n15 0.738255
R7605 commonsourceibias.n46 commonsourceibias.n45 0.738255
R7606 commonsourceibias.n5 commonsourceibias.n3 0.738255
R7607 commonsourceibias.n139 commonsourceibias.n138 0.738255
R7608 commonsourceibias.n318 commonsourceibias.n317 0.738255
R7609 commonsourceibias.n289 commonsourceibias.n287 0.738255
R7610 commonsourceibias.n199 commonsourceibias.n197 0.738255
R7611 commonsourceibias.n228 commonsourceibias.n227 0.738255
R7612 commonsourceibias.n465 commonsourceibias.n464 0.738255
R7613 commonsourceibias.n505 commonsourceibias.n436 0.738255
R7614 commonsourceibias.n551 commonsourceibias.n377 0.738255
R7615 commonsourceibias.n406 commonsourceibias.n405 0.738255
R7616 commonsourceibias.n690 commonsourceibias.n689 0.738255
R7617 commonsourceibias.n730 commonsourceibias.n661 0.738255
R7618 commonsourceibias.n600 commonsourceibias.n599 0.738255
R7619 commonsourceibias.n640 commonsourceibias.n571 0.738255
R7620 commonsourceibias.n104 commonsourceibias.n102 0.573776
R7621 commonsourceibias.n106 commonsourceibias.n104 0.573776
R7622 commonsourceibias.n108 commonsourceibias.n106 0.573776
R7623 commonsourceibias.n115 commonsourceibias.n113 0.573776
R7624 commonsourceibias.n113 commonsourceibias.n111 0.573776
R7625 commonsourceibias.n430 commonsourceibias.n428 0.573776
R7626 commonsourceibias.n432 commonsourceibias.n430 0.573776
R7627 commonsourceibias.n529 commonsourceibias.n527 0.573776
R7628 commonsourceibias.n527 commonsourceibias.n525 0.573776
R7629 commonsourceibias.n525 commonsourceibias.n523 0.573776
R7630 commonsourceibias.n116 commonsourceibias.n108 0.287138
R7631 commonsourceibias.n116 commonsourceibias.n115 0.287138
R7632 commonsourceibias.n530 commonsourceibias.n432 0.287138
R7633 commonsourceibias.n530 commonsourceibias.n529 0.287138
R7634 commonsourceibias.n100 commonsourceibias.n12 0.285035
R7635 commonsourceibias.n193 commonsourceibias.n0 0.285035
R7636 commonsourceibias.n372 commonsourceibias.n284 0.285035
R7637 commonsourceibias.n282 commonsourceibias.n194 0.285035
R7638 commonsourceibias.n521 commonsourceibias.n433 0.285035
R7639 commonsourceibias.n567 commonsourceibias.n374 0.285035
R7640 commonsourceibias.n746 commonsourceibias.n658 0.285035
R7641 commonsourceibias.n656 commonsourceibias.n568 0.285035
R7642 commonsourceibias.n22 commonsourceibias.n20 0.246418
R7643 commonsourceibias.n58 commonsourceibias.n25 0.246418
R7644 commonsourceibias.n10 commonsourceibias.n8 0.246418
R7645 commonsourceibias.n151 commonsourceibias.n118 0.246418
R7646 commonsourceibias.n330 commonsourceibias.n297 0.246418
R7647 commonsourceibias.n294 commonsourceibias.n292 0.246418
R7648 commonsourceibias.n204 commonsourceibias.n202 0.246418
R7649 commonsourceibias.n240 commonsourceibias.n207 0.246418
R7650 commonsourceibias.n477 commonsourceibias.n444 0.246418
R7651 commonsourceibias.n490 commonsourceibias.n440 0.246418
R7652 commonsourceibias.n536 commonsourceibias.n381 0.246418
R7653 commonsourceibias.n418 commonsourceibias.n385 0.246418
R7654 commonsourceibias.n702 commonsourceibias.n669 0.246418
R7655 commonsourceibias.n715 commonsourceibias.n665 0.246418
R7656 commonsourceibias.n612 commonsourceibias.n579 0.246418
R7657 commonsourceibias.n625 commonsourceibias.n575 0.246418
R7658 commonsourceibias.n95 commonsourceibias.n12 0.189894
R7659 commonsourceibias.n95 commonsourceibias.n94 0.189894
R7660 commonsourceibias.n94 commonsourceibias.n93 0.189894
R7661 commonsourceibias.n93 commonsourceibias.n14 0.189894
R7662 commonsourceibias.n88 commonsourceibias.n14 0.189894
R7663 commonsourceibias.n88 commonsourceibias.n87 0.189894
R7664 commonsourceibias.n87 commonsourceibias.n86 0.189894
R7665 commonsourceibias.n86 commonsourceibias.n16 0.189894
R7666 commonsourceibias.n81 commonsourceibias.n16 0.189894
R7667 commonsourceibias.n81 commonsourceibias.n80 0.189894
R7668 commonsourceibias.n80 commonsourceibias.n79 0.189894
R7669 commonsourceibias.n79 commonsourceibias.n19 0.189894
R7670 commonsourceibias.n74 commonsourceibias.n19 0.189894
R7671 commonsourceibias.n74 commonsourceibias.n73 0.189894
R7672 commonsourceibias.n73 commonsourceibias.n72 0.189894
R7673 commonsourceibias.n72 commonsourceibias.n21 0.189894
R7674 commonsourceibias.n67 commonsourceibias.n21 0.189894
R7675 commonsourceibias.n67 commonsourceibias.n66 0.189894
R7676 commonsourceibias.n66 commonsourceibias.n65 0.189894
R7677 commonsourceibias.n65 commonsourceibias.n24 0.189894
R7678 commonsourceibias.n60 commonsourceibias.n24 0.189894
R7679 commonsourceibias.n60 commonsourceibias.n59 0.189894
R7680 commonsourceibias.n59 commonsourceibias.n26 0.189894
R7681 commonsourceibias.n55 commonsourceibias.n26 0.189894
R7682 commonsourceibias.n55 commonsourceibias.n54 0.189894
R7683 commonsourceibias.n54 commonsourceibias.n28 0.189894
R7684 commonsourceibias.n50 commonsourceibias.n28 0.189894
R7685 commonsourceibias.n50 commonsourceibias.n49 0.189894
R7686 commonsourceibias.n49 commonsourceibias.n30 0.189894
R7687 commonsourceibias.n44 commonsourceibias.n30 0.189894
R7688 commonsourceibias.n44 commonsourceibias.n43 0.189894
R7689 commonsourceibias.n43 commonsourceibias.n42 0.189894
R7690 commonsourceibias.n42 commonsourceibias.n32 0.189894
R7691 commonsourceibias.n37 commonsourceibias.n32 0.189894
R7692 commonsourceibias.n37 commonsourceibias.n36 0.189894
R7693 commonsourceibias.n158 commonsourceibias.n117 0.189894
R7694 commonsourceibias.n153 commonsourceibias.n117 0.189894
R7695 commonsourceibias.n153 commonsourceibias.n152 0.189894
R7696 commonsourceibias.n152 commonsourceibias.n119 0.189894
R7697 commonsourceibias.n148 commonsourceibias.n119 0.189894
R7698 commonsourceibias.n148 commonsourceibias.n147 0.189894
R7699 commonsourceibias.n147 commonsourceibias.n121 0.189894
R7700 commonsourceibias.n143 commonsourceibias.n121 0.189894
R7701 commonsourceibias.n143 commonsourceibias.n142 0.189894
R7702 commonsourceibias.n142 commonsourceibias.n123 0.189894
R7703 commonsourceibias.n137 commonsourceibias.n123 0.189894
R7704 commonsourceibias.n137 commonsourceibias.n136 0.189894
R7705 commonsourceibias.n136 commonsourceibias.n135 0.189894
R7706 commonsourceibias.n135 commonsourceibias.n125 0.189894
R7707 commonsourceibias.n130 commonsourceibias.n125 0.189894
R7708 commonsourceibias.n130 commonsourceibias.n129 0.189894
R7709 commonsourceibias.n188 commonsourceibias.n0 0.189894
R7710 commonsourceibias.n188 commonsourceibias.n187 0.189894
R7711 commonsourceibias.n187 commonsourceibias.n186 0.189894
R7712 commonsourceibias.n186 commonsourceibias.n2 0.189894
R7713 commonsourceibias.n181 commonsourceibias.n2 0.189894
R7714 commonsourceibias.n181 commonsourceibias.n180 0.189894
R7715 commonsourceibias.n180 commonsourceibias.n179 0.189894
R7716 commonsourceibias.n179 commonsourceibias.n4 0.189894
R7717 commonsourceibias.n174 commonsourceibias.n4 0.189894
R7718 commonsourceibias.n174 commonsourceibias.n173 0.189894
R7719 commonsourceibias.n173 commonsourceibias.n172 0.189894
R7720 commonsourceibias.n172 commonsourceibias.n7 0.189894
R7721 commonsourceibias.n167 commonsourceibias.n7 0.189894
R7722 commonsourceibias.n167 commonsourceibias.n166 0.189894
R7723 commonsourceibias.n166 commonsourceibias.n165 0.189894
R7724 commonsourceibias.n165 commonsourceibias.n9 0.189894
R7725 commonsourceibias.n160 commonsourceibias.n9 0.189894
R7726 commonsourceibias.n367 commonsourceibias.n284 0.189894
R7727 commonsourceibias.n367 commonsourceibias.n366 0.189894
R7728 commonsourceibias.n366 commonsourceibias.n365 0.189894
R7729 commonsourceibias.n365 commonsourceibias.n286 0.189894
R7730 commonsourceibias.n360 commonsourceibias.n286 0.189894
R7731 commonsourceibias.n360 commonsourceibias.n359 0.189894
R7732 commonsourceibias.n359 commonsourceibias.n358 0.189894
R7733 commonsourceibias.n358 commonsourceibias.n288 0.189894
R7734 commonsourceibias.n353 commonsourceibias.n288 0.189894
R7735 commonsourceibias.n353 commonsourceibias.n352 0.189894
R7736 commonsourceibias.n352 commonsourceibias.n351 0.189894
R7737 commonsourceibias.n351 commonsourceibias.n291 0.189894
R7738 commonsourceibias.n346 commonsourceibias.n291 0.189894
R7739 commonsourceibias.n346 commonsourceibias.n345 0.189894
R7740 commonsourceibias.n345 commonsourceibias.n344 0.189894
R7741 commonsourceibias.n344 commonsourceibias.n293 0.189894
R7742 commonsourceibias.n339 commonsourceibias.n293 0.189894
R7743 commonsourceibias.n339 commonsourceibias.n338 0.189894
R7744 commonsourceibias.n338 commonsourceibias.n337 0.189894
R7745 commonsourceibias.n337 commonsourceibias.n296 0.189894
R7746 commonsourceibias.n332 commonsourceibias.n296 0.189894
R7747 commonsourceibias.n332 commonsourceibias.n331 0.189894
R7748 commonsourceibias.n331 commonsourceibias.n298 0.189894
R7749 commonsourceibias.n327 commonsourceibias.n298 0.189894
R7750 commonsourceibias.n327 commonsourceibias.n326 0.189894
R7751 commonsourceibias.n326 commonsourceibias.n300 0.189894
R7752 commonsourceibias.n322 commonsourceibias.n300 0.189894
R7753 commonsourceibias.n322 commonsourceibias.n321 0.189894
R7754 commonsourceibias.n321 commonsourceibias.n302 0.189894
R7755 commonsourceibias.n316 commonsourceibias.n302 0.189894
R7756 commonsourceibias.n316 commonsourceibias.n315 0.189894
R7757 commonsourceibias.n315 commonsourceibias.n314 0.189894
R7758 commonsourceibias.n314 commonsourceibias.n304 0.189894
R7759 commonsourceibias.n309 commonsourceibias.n304 0.189894
R7760 commonsourceibias.n309 commonsourceibias.n308 0.189894
R7761 commonsourceibias.n277 commonsourceibias.n194 0.189894
R7762 commonsourceibias.n277 commonsourceibias.n276 0.189894
R7763 commonsourceibias.n276 commonsourceibias.n275 0.189894
R7764 commonsourceibias.n275 commonsourceibias.n196 0.189894
R7765 commonsourceibias.n270 commonsourceibias.n196 0.189894
R7766 commonsourceibias.n270 commonsourceibias.n269 0.189894
R7767 commonsourceibias.n269 commonsourceibias.n268 0.189894
R7768 commonsourceibias.n268 commonsourceibias.n198 0.189894
R7769 commonsourceibias.n263 commonsourceibias.n198 0.189894
R7770 commonsourceibias.n263 commonsourceibias.n262 0.189894
R7771 commonsourceibias.n262 commonsourceibias.n261 0.189894
R7772 commonsourceibias.n261 commonsourceibias.n201 0.189894
R7773 commonsourceibias.n256 commonsourceibias.n201 0.189894
R7774 commonsourceibias.n256 commonsourceibias.n255 0.189894
R7775 commonsourceibias.n255 commonsourceibias.n254 0.189894
R7776 commonsourceibias.n254 commonsourceibias.n203 0.189894
R7777 commonsourceibias.n249 commonsourceibias.n203 0.189894
R7778 commonsourceibias.n249 commonsourceibias.n248 0.189894
R7779 commonsourceibias.n248 commonsourceibias.n247 0.189894
R7780 commonsourceibias.n247 commonsourceibias.n206 0.189894
R7781 commonsourceibias.n242 commonsourceibias.n206 0.189894
R7782 commonsourceibias.n242 commonsourceibias.n241 0.189894
R7783 commonsourceibias.n241 commonsourceibias.n208 0.189894
R7784 commonsourceibias.n237 commonsourceibias.n208 0.189894
R7785 commonsourceibias.n237 commonsourceibias.n236 0.189894
R7786 commonsourceibias.n236 commonsourceibias.n210 0.189894
R7787 commonsourceibias.n232 commonsourceibias.n210 0.189894
R7788 commonsourceibias.n232 commonsourceibias.n231 0.189894
R7789 commonsourceibias.n231 commonsourceibias.n212 0.189894
R7790 commonsourceibias.n226 commonsourceibias.n212 0.189894
R7791 commonsourceibias.n226 commonsourceibias.n225 0.189894
R7792 commonsourceibias.n225 commonsourceibias.n224 0.189894
R7793 commonsourceibias.n224 commonsourceibias.n214 0.189894
R7794 commonsourceibias.n219 commonsourceibias.n214 0.189894
R7795 commonsourceibias.n219 commonsourceibias.n218 0.189894
R7796 commonsourceibias.n456 commonsourceibias.n455 0.189894
R7797 commonsourceibias.n456 commonsourceibias.n451 0.189894
R7798 commonsourceibias.n461 commonsourceibias.n451 0.189894
R7799 commonsourceibias.n462 commonsourceibias.n461 0.189894
R7800 commonsourceibias.n463 commonsourceibias.n462 0.189894
R7801 commonsourceibias.n463 commonsourceibias.n449 0.189894
R7802 commonsourceibias.n468 commonsourceibias.n449 0.189894
R7803 commonsourceibias.n469 commonsourceibias.n468 0.189894
R7804 commonsourceibias.n469 commonsourceibias.n447 0.189894
R7805 commonsourceibias.n473 commonsourceibias.n447 0.189894
R7806 commonsourceibias.n474 commonsourceibias.n473 0.189894
R7807 commonsourceibias.n474 commonsourceibias.n445 0.189894
R7808 commonsourceibias.n478 commonsourceibias.n445 0.189894
R7809 commonsourceibias.n479 commonsourceibias.n478 0.189894
R7810 commonsourceibias.n479 commonsourceibias.n443 0.189894
R7811 commonsourceibias.n484 commonsourceibias.n443 0.189894
R7812 commonsourceibias.n485 commonsourceibias.n484 0.189894
R7813 commonsourceibias.n486 commonsourceibias.n485 0.189894
R7814 commonsourceibias.n486 commonsourceibias.n441 0.189894
R7815 commonsourceibias.n492 commonsourceibias.n441 0.189894
R7816 commonsourceibias.n493 commonsourceibias.n492 0.189894
R7817 commonsourceibias.n494 commonsourceibias.n493 0.189894
R7818 commonsourceibias.n494 commonsourceibias.n439 0.189894
R7819 commonsourceibias.n499 commonsourceibias.n439 0.189894
R7820 commonsourceibias.n500 commonsourceibias.n499 0.189894
R7821 commonsourceibias.n501 commonsourceibias.n500 0.189894
R7822 commonsourceibias.n501 commonsourceibias.n437 0.189894
R7823 commonsourceibias.n507 commonsourceibias.n437 0.189894
R7824 commonsourceibias.n508 commonsourceibias.n507 0.189894
R7825 commonsourceibias.n509 commonsourceibias.n508 0.189894
R7826 commonsourceibias.n509 commonsourceibias.n435 0.189894
R7827 commonsourceibias.n514 commonsourceibias.n435 0.189894
R7828 commonsourceibias.n515 commonsourceibias.n514 0.189894
R7829 commonsourceibias.n516 commonsourceibias.n515 0.189894
R7830 commonsourceibias.n516 commonsourceibias.n433 0.189894
R7831 commonsourceibias.n397 commonsourceibias.n396 0.189894
R7832 commonsourceibias.n397 commonsourceibias.n392 0.189894
R7833 commonsourceibias.n402 commonsourceibias.n392 0.189894
R7834 commonsourceibias.n403 commonsourceibias.n402 0.189894
R7835 commonsourceibias.n404 commonsourceibias.n403 0.189894
R7836 commonsourceibias.n404 commonsourceibias.n390 0.189894
R7837 commonsourceibias.n409 commonsourceibias.n390 0.189894
R7838 commonsourceibias.n410 commonsourceibias.n409 0.189894
R7839 commonsourceibias.n410 commonsourceibias.n388 0.189894
R7840 commonsourceibias.n414 commonsourceibias.n388 0.189894
R7841 commonsourceibias.n415 commonsourceibias.n414 0.189894
R7842 commonsourceibias.n415 commonsourceibias.n386 0.189894
R7843 commonsourceibias.n419 commonsourceibias.n386 0.189894
R7844 commonsourceibias.n420 commonsourceibias.n419 0.189894
R7845 commonsourceibias.n420 commonsourceibias.n384 0.189894
R7846 commonsourceibias.n425 commonsourceibias.n384 0.189894
R7847 commonsourceibias.n532 commonsourceibias.n382 0.189894
R7848 commonsourceibias.n538 commonsourceibias.n382 0.189894
R7849 commonsourceibias.n539 commonsourceibias.n538 0.189894
R7850 commonsourceibias.n540 commonsourceibias.n539 0.189894
R7851 commonsourceibias.n540 commonsourceibias.n380 0.189894
R7852 commonsourceibias.n545 commonsourceibias.n380 0.189894
R7853 commonsourceibias.n546 commonsourceibias.n545 0.189894
R7854 commonsourceibias.n547 commonsourceibias.n546 0.189894
R7855 commonsourceibias.n547 commonsourceibias.n378 0.189894
R7856 commonsourceibias.n553 commonsourceibias.n378 0.189894
R7857 commonsourceibias.n554 commonsourceibias.n553 0.189894
R7858 commonsourceibias.n555 commonsourceibias.n554 0.189894
R7859 commonsourceibias.n555 commonsourceibias.n376 0.189894
R7860 commonsourceibias.n560 commonsourceibias.n376 0.189894
R7861 commonsourceibias.n561 commonsourceibias.n560 0.189894
R7862 commonsourceibias.n562 commonsourceibias.n561 0.189894
R7863 commonsourceibias.n562 commonsourceibias.n374 0.189894
R7864 commonsourceibias.n681 commonsourceibias.n680 0.189894
R7865 commonsourceibias.n681 commonsourceibias.n676 0.189894
R7866 commonsourceibias.n686 commonsourceibias.n676 0.189894
R7867 commonsourceibias.n687 commonsourceibias.n686 0.189894
R7868 commonsourceibias.n688 commonsourceibias.n687 0.189894
R7869 commonsourceibias.n688 commonsourceibias.n674 0.189894
R7870 commonsourceibias.n693 commonsourceibias.n674 0.189894
R7871 commonsourceibias.n694 commonsourceibias.n693 0.189894
R7872 commonsourceibias.n694 commonsourceibias.n672 0.189894
R7873 commonsourceibias.n698 commonsourceibias.n672 0.189894
R7874 commonsourceibias.n699 commonsourceibias.n698 0.189894
R7875 commonsourceibias.n699 commonsourceibias.n670 0.189894
R7876 commonsourceibias.n703 commonsourceibias.n670 0.189894
R7877 commonsourceibias.n704 commonsourceibias.n703 0.189894
R7878 commonsourceibias.n704 commonsourceibias.n668 0.189894
R7879 commonsourceibias.n709 commonsourceibias.n668 0.189894
R7880 commonsourceibias.n710 commonsourceibias.n709 0.189894
R7881 commonsourceibias.n711 commonsourceibias.n710 0.189894
R7882 commonsourceibias.n711 commonsourceibias.n666 0.189894
R7883 commonsourceibias.n717 commonsourceibias.n666 0.189894
R7884 commonsourceibias.n718 commonsourceibias.n717 0.189894
R7885 commonsourceibias.n719 commonsourceibias.n718 0.189894
R7886 commonsourceibias.n719 commonsourceibias.n664 0.189894
R7887 commonsourceibias.n724 commonsourceibias.n664 0.189894
R7888 commonsourceibias.n725 commonsourceibias.n724 0.189894
R7889 commonsourceibias.n726 commonsourceibias.n725 0.189894
R7890 commonsourceibias.n726 commonsourceibias.n662 0.189894
R7891 commonsourceibias.n732 commonsourceibias.n662 0.189894
R7892 commonsourceibias.n733 commonsourceibias.n732 0.189894
R7893 commonsourceibias.n734 commonsourceibias.n733 0.189894
R7894 commonsourceibias.n734 commonsourceibias.n660 0.189894
R7895 commonsourceibias.n739 commonsourceibias.n660 0.189894
R7896 commonsourceibias.n740 commonsourceibias.n739 0.189894
R7897 commonsourceibias.n741 commonsourceibias.n740 0.189894
R7898 commonsourceibias.n741 commonsourceibias.n658 0.189894
R7899 commonsourceibias.n591 commonsourceibias.n590 0.189894
R7900 commonsourceibias.n591 commonsourceibias.n586 0.189894
R7901 commonsourceibias.n596 commonsourceibias.n586 0.189894
R7902 commonsourceibias.n597 commonsourceibias.n596 0.189894
R7903 commonsourceibias.n598 commonsourceibias.n597 0.189894
R7904 commonsourceibias.n598 commonsourceibias.n584 0.189894
R7905 commonsourceibias.n603 commonsourceibias.n584 0.189894
R7906 commonsourceibias.n604 commonsourceibias.n603 0.189894
R7907 commonsourceibias.n604 commonsourceibias.n582 0.189894
R7908 commonsourceibias.n608 commonsourceibias.n582 0.189894
R7909 commonsourceibias.n609 commonsourceibias.n608 0.189894
R7910 commonsourceibias.n609 commonsourceibias.n580 0.189894
R7911 commonsourceibias.n613 commonsourceibias.n580 0.189894
R7912 commonsourceibias.n614 commonsourceibias.n613 0.189894
R7913 commonsourceibias.n614 commonsourceibias.n578 0.189894
R7914 commonsourceibias.n619 commonsourceibias.n578 0.189894
R7915 commonsourceibias.n620 commonsourceibias.n619 0.189894
R7916 commonsourceibias.n621 commonsourceibias.n620 0.189894
R7917 commonsourceibias.n621 commonsourceibias.n576 0.189894
R7918 commonsourceibias.n627 commonsourceibias.n576 0.189894
R7919 commonsourceibias.n628 commonsourceibias.n627 0.189894
R7920 commonsourceibias.n629 commonsourceibias.n628 0.189894
R7921 commonsourceibias.n629 commonsourceibias.n574 0.189894
R7922 commonsourceibias.n634 commonsourceibias.n574 0.189894
R7923 commonsourceibias.n635 commonsourceibias.n634 0.189894
R7924 commonsourceibias.n636 commonsourceibias.n635 0.189894
R7925 commonsourceibias.n636 commonsourceibias.n572 0.189894
R7926 commonsourceibias.n642 commonsourceibias.n572 0.189894
R7927 commonsourceibias.n643 commonsourceibias.n642 0.189894
R7928 commonsourceibias.n644 commonsourceibias.n643 0.189894
R7929 commonsourceibias.n644 commonsourceibias.n570 0.189894
R7930 commonsourceibias.n649 commonsourceibias.n570 0.189894
R7931 commonsourceibias.n650 commonsourceibias.n649 0.189894
R7932 commonsourceibias.n651 commonsourceibias.n650 0.189894
R7933 commonsourceibias.n651 commonsourceibias.n568 0.189894
R7934 commonsourceibias.n159 commonsourceibias.n158 0.170955
R7935 commonsourceibias.n160 commonsourceibias.n159 0.170955
R7936 commonsourceibias.n531 commonsourceibias.n425 0.170955
R7937 commonsourceibias.n532 commonsourceibias.n531 0.170955
R7938 gnd.n4039 gnd.n3725 939.716
R7939 gnd.n6505 gnd.n520 870.29
R7940 gnd.n211 gnd.n201 795.207
R7941 gnd.n6952 gnd.n6951 795.207
R7942 gnd.n5273 gnd.n1277 795.207
R7943 gnd.n5477 gnd.n5476 795.207
R7944 gnd.n979 gnd.n967 795.207
R7945 gnd.n4470 gnd.n4469 795.207
R7946 gnd.n3879 gnd.n3762 795.207
R7947 gnd.n3918 gnd.n2240 795.207
R7948 gnd.n1943 gnd.n1841 771.183
R7949 gnd.n5242 gnd.n1356 771.183
R7950 gnd.n4479 gnd.n1843 771.183
R7951 gnd.n5716 gnd.n1215 771.183
R7952 gnd.n3633 gnd.n2248 766.379
R7953 gnd.n3636 gnd.n3635 766.379
R7954 gnd.n2875 gnd.n2778 766.379
R7955 gnd.n2871 gnd.n2776 766.379
R7956 gnd.n3724 gnd.n2270 756.769
R7957 gnd.n3627 gnd.n3626 756.769
R7958 gnd.n2968 gnd.n2685 756.769
R7959 gnd.n2966 gnd.n2688 756.769
R7960 gnd.n7112 gnd.n205 739.952
R7961 gnd.n6988 gnd.n6987 739.952
R7962 gnd.n5272 gnd.n5271 739.952
R7963 gnd.n5706 gnd.n1281 739.952
R7964 gnd.n5952 gnd.n972 739.952
R7965 gnd.n2048 gnd.n1852 739.952
R7966 gnd.n4042 gnd.n4041 739.952
R7967 gnd.n4037 gnd.n2236 739.952
R7968 gnd.n6177 gnd.n712 655.866
R7969 gnd.n6504 gnd.n521 655.866
R7970 gnd.n6716 gnd.n6715 655.866
R7971 gnd.n6009 gnd.n882 655.866
R7972 gnd.n6178 gnd.n6177 585
R7973 gnd.n6177 gnd.n6176 585
R7974 gnd.n716 gnd.n715 585
R7975 gnd.n6175 gnd.n716 585
R7976 gnd.n6173 gnd.n6172 585
R7977 gnd.n6174 gnd.n6173 585
R7978 gnd.n6171 gnd.n718 585
R7979 gnd.n718 gnd.n717 585
R7980 gnd.n6170 gnd.n6169 585
R7981 gnd.n6169 gnd.n6168 585
R7982 gnd.n723 gnd.n722 585
R7983 gnd.n6167 gnd.n723 585
R7984 gnd.n6165 gnd.n6164 585
R7985 gnd.n6166 gnd.n6165 585
R7986 gnd.n6163 gnd.n725 585
R7987 gnd.n725 gnd.n724 585
R7988 gnd.n6162 gnd.n6161 585
R7989 gnd.n6161 gnd.n6160 585
R7990 gnd.n731 gnd.n730 585
R7991 gnd.n6159 gnd.n731 585
R7992 gnd.n6157 gnd.n6156 585
R7993 gnd.n6158 gnd.n6157 585
R7994 gnd.n6155 gnd.n733 585
R7995 gnd.n733 gnd.n732 585
R7996 gnd.n6154 gnd.n6153 585
R7997 gnd.n6153 gnd.n6152 585
R7998 gnd.n739 gnd.n738 585
R7999 gnd.n6151 gnd.n739 585
R8000 gnd.n6149 gnd.n6148 585
R8001 gnd.n6150 gnd.n6149 585
R8002 gnd.n6147 gnd.n741 585
R8003 gnd.n741 gnd.n740 585
R8004 gnd.n6146 gnd.n6145 585
R8005 gnd.n6145 gnd.n6144 585
R8006 gnd.n747 gnd.n746 585
R8007 gnd.n6143 gnd.n747 585
R8008 gnd.n6141 gnd.n6140 585
R8009 gnd.n6142 gnd.n6141 585
R8010 gnd.n6139 gnd.n749 585
R8011 gnd.n749 gnd.n748 585
R8012 gnd.n6138 gnd.n6137 585
R8013 gnd.n6137 gnd.n6136 585
R8014 gnd.n755 gnd.n754 585
R8015 gnd.n6135 gnd.n755 585
R8016 gnd.n6133 gnd.n6132 585
R8017 gnd.n6134 gnd.n6133 585
R8018 gnd.n6131 gnd.n757 585
R8019 gnd.n757 gnd.n756 585
R8020 gnd.n6130 gnd.n6129 585
R8021 gnd.n6129 gnd.n6128 585
R8022 gnd.n763 gnd.n762 585
R8023 gnd.n6127 gnd.n763 585
R8024 gnd.n6125 gnd.n6124 585
R8025 gnd.n6126 gnd.n6125 585
R8026 gnd.n6123 gnd.n765 585
R8027 gnd.n765 gnd.n764 585
R8028 gnd.n6122 gnd.n6121 585
R8029 gnd.n6121 gnd.n6120 585
R8030 gnd.n771 gnd.n770 585
R8031 gnd.n6119 gnd.n771 585
R8032 gnd.n6117 gnd.n6116 585
R8033 gnd.n6118 gnd.n6117 585
R8034 gnd.n6115 gnd.n773 585
R8035 gnd.n773 gnd.n772 585
R8036 gnd.n6114 gnd.n6113 585
R8037 gnd.n6113 gnd.n6112 585
R8038 gnd.n779 gnd.n778 585
R8039 gnd.n6111 gnd.n779 585
R8040 gnd.n6109 gnd.n6108 585
R8041 gnd.n6110 gnd.n6109 585
R8042 gnd.n6107 gnd.n781 585
R8043 gnd.n781 gnd.n780 585
R8044 gnd.n6106 gnd.n6105 585
R8045 gnd.n6105 gnd.n6104 585
R8046 gnd.n787 gnd.n786 585
R8047 gnd.n6103 gnd.n787 585
R8048 gnd.n6101 gnd.n6100 585
R8049 gnd.n6102 gnd.n6101 585
R8050 gnd.n6099 gnd.n789 585
R8051 gnd.n789 gnd.n788 585
R8052 gnd.n6098 gnd.n6097 585
R8053 gnd.n6097 gnd.n6096 585
R8054 gnd.n795 gnd.n794 585
R8055 gnd.n6095 gnd.n795 585
R8056 gnd.n6093 gnd.n6092 585
R8057 gnd.n6094 gnd.n6093 585
R8058 gnd.n6091 gnd.n797 585
R8059 gnd.n797 gnd.n796 585
R8060 gnd.n6090 gnd.n6089 585
R8061 gnd.n6089 gnd.n6088 585
R8062 gnd.n803 gnd.n802 585
R8063 gnd.n6087 gnd.n803 585
R8064 gnd.n6085 gnd.n6084 585
R8065 gnd.n6086 gnd.n6085 585
R8066 gnd.n6083 gnd.n805 585
R8067 gnd.n805 gnd.n804 585
R8068 gnd.n6082 gnd.n6081 585
R8069 gnd.n6081 gnd.n6080 585
R8070 gnd.n811 gnd.n810 585
R8071 gnd.n6079 gnd.n811 585
R8072 gnd.n6077 gnd.n6076 585
R8073 gnd.n6078 gnd.n6077 585
R8074 gnd.n6075 gnd.n813 585
R8075 gnd.n813 gnd.n812 585
R8076 gnd.n6074 gnd.n6073 585
R8077 gnd.n6073 gnd.n6072 585
R8078 gnd.n819 gnd.n818 585
R8079 gnd.n6071 gnd.n819 585
R8080 gnd.n6069 gnd.n6068 585
R8081 gnd.n6070 gnd.n6069 585
R8082 gnd.n6067 gnd.n821 585
R8083 gnd.n821 gnd.n820 585
R8084 gnd.n6066 gnd.n6065 585
R8085 gnd.n6065 gnd.n6064 585
R8086 gnd.n827 gnd.n826 585
R8087 gnd.n6063 gnd.n827 585
R8088 gnd.n6061 gnd.n6060 585
R8089 gnd.n6062 gnd.n6061 585
R8090 gnd.n6059 gnd.n829 585
R8091 gnd.n829 gnd.n828 585
R8092 gnd.n6058 gnd.n6057 585
R8093 gnd.n6057 gnd.n6056 585
R8094 gnd.n835 gnd.n834 585
R8095 gnd.n6055 gnd.n835 585
R8096 gnd.n6053 gnd.n6052 585
R8097 gnd.n6054 gnd.n6053 585
R8098 gnd.n6051 gnd.n837 585
R8099 gnd.n837 gnd.n836 585
R8100 gnd.n6050 gnd.n6049 585
R8101 gnd.n6049 gnd.n6048 585
R8102 gnd.n843 gnd.n842 585
R8103 gnd.n6047 gnd.n843 585
R8104 gnd.n6045 gnd.n6044 585
R8105 gnd.n6046 gnd.n6045 585
R8106 gnd.n6043 gnd.n845 585
R8107 gnd.n845 gnd.n844 585
R8108 gnd.n6042 gnd.n6041 585
R8109 gnd.n6041 gnd.n6040 585
R8110 gnd.n851 gnd.n850 585
R8111 gnd.n6039 gnd.n851 585
R8112 gnd.n6037 gnd.n6036 585
R8113 gnd.n6038 gnd.n6037 585
R8114 gnd.n6035 gnd.n853 585
R8115 gnd.n853 gnd.n852 585
R8116 gnd.n6034 gnd.n6033 585
R8117 gnd.n6033 gnd.n6032 585
R8118 gnd.n859 gnd.n858 585
R8119 gnd.n6031 gnd.n859 585
R8120 gnd.n6029 gnd.n6028 585
R8121 gnd.n6030 gnd.n6029 585
R8122 gnd.n6027 gnd.n861 585
R8123 gnd.n861 gnd.n860 585
R8124 gnd.n6026 gnd.n6025 585
R8125 gnd.n6025 gnd.n6024 585
R8126 gnd.n867 gnd.n866 585
R8127 gnd.n6023 gnd.n867 585
R8128 gnd.n6021 gnd.n6020 585
R8129 gnd.n6022 gnd.n6021 585
R8130 gnd.n6019 gnd.n869 585
R8131 gnd.n869 gnd.n868 585
R8132 gnd.n6018 gnd.n6017 585
R8133 gnd.n6017 gnd.n6016 585
R8134 gnd.n875 gnd.n874 585
R8135 gnd.n6015 gnd.n875 585
R8136 gnd.n6013 gnd.n6012 585
R8137 gnd.n6014 gnd.n6013 585
R8138 gnd.n6011 gnd.n877 585
R8139 gnd.n877 gnd.n876 585
R8140 gnd.n713 gnd.n712 585
R8141 gnd.n712 gnd.n711 585
R8142 gnd.n6183 gnd.n6182 585
R8143 gnd.n6184 gnd.n6183 585
R8144 gnd.n710 gnd.n709 585
R8145 gnd.n6185 gnd.n710 585
R8146 gnd.n6188 gnd.n6187 585
R8147 gnd.n6187 gnd.n6186 585
R8148 gnd.n707 gnd.n706 585
R8149 gnd.n706 gnd.n705 585
R8150 gnd.n6193 gnd.n6192 585
R8151 gnd.n6194 gnd.n6193 585
R8152 gnd.n704 gnd.n703 585
R8153 gnd.n6195 gnd.n704 585
R8154 gnd.n6198 gnd.n6197 585
R8155 gnd.n6197 gnd.n6196 585
R8156 gnd.n701 gnd.n700 585
R8157 gnd.n700 gnd.n699 585
R8158 gnd.n6203 gnd.n6202 585
R8159 gnd.n6204 gnd.n6203 585
R8160 gnd.n698 gnd.n697 585
R8161 gnd.n6205 gnd.n698 585
R8162 gnd.n6208 gnd.n6207 585
R8163 gnd.n6207 gnd.n6206 585
R8164 gnd.n695 gnd.n694 585
R8165 gnd.n694 gnd.n693 585
R8166 gnd.n6213 gnd.n6212 585
R8167 gnd.n6214 gnd.n6213 585
R8168 gnd.n692 gnd.n691 585
R8169 gnd.n6215 gnd.n692 585
R8170 gnd.n6218 gnd.n6217 585
R8171 gnd.n6217 gnd.n6216 585
R8172 gnd.n689 gnd.n688 585
R8173 gnd.n688 gnd.n687 585
R8174 gnd.n6223 gnd.n6222 585
R8175 gnd.n6224 gnd.n6223 585
R8176 gnd.n686 gnd.n685 585
R8177 gnd.n6225 gnd.n686 585
R8178 gnd.n6228 gnd.n6227 585
R8179 gnd.n6227 gnd.n6226 585
R8180 gnd.n683 gnd.n682 585
R8181 gnd.n682 gnd.n681 585
R8182 gnd.n6233 gnd.n6232 585
R8183 gnd.n6234 gnd.n6233 585
R8184 gnd.n680 gnd.n679 585
R8185 gnd.n6235 gnd.n680 585
R8186 gnd.n6238 gnd.n6237 585
R8187 gnd.n6237 gnd.n6236 585
R8188 gnd.n677 gnd.n676 585
R8189 gnd.n676 gnd.n675 585
R8190 gnd.n6243 gnd.n6242 585
R8191 gnd.n6244 gnd.n6243 585
R8192 gnd.n674 gnd.n673 585
R8193 gnd.n6245 gnd.n674 585
R8194 gnd.n6248 gnd.n6247 585
R8195 gnd.n6247 gnd.n6246 585
R8196 gnd.n671 gnd.n670 585
R8197 gnd.n670 gnd.n669 585
R8198 gnd.n6253 gnd.n6252 585
R8199 gnd.n6254 gnd.n6253 585
R8200 gnd.n668 gnd.n667 585
R8201 gnd.n6255 gnd.n668 585
R8202 gnd.n6258 gnd.n6257 585
R8203 gnd.n6257 gnd.n6256 585
R8204 gnd.n665 gnd.n664 585
R8205 gnd.n664 gnd.n663 585
R8206 gnd.n6263 gnd.n6262 585
R8207 gnd.n6264 gnd.n6263 585
R8208 gnd.n662 gnd.n661 585
R8209 gnd.n6265 gnd.n662 585
R8210 gnd.n6268 gnd.n6267 585
R8211 gnd.n6267 gnd.n6266 585
R8212 gnd.n659 gnd.n658 585
R8213 gnd.n658 gnd.n657 585
R8214 gnd.n6273 gnd.n6272 585
R8215 gnd.n6274 gnd.n6273 585
R8216 gnd.n656 gnd.n655 585
R8217 gnd.n6275 gnd.n656 585
R8218 gnd.n6278 gnd.n6277 585
R8219 gnd.n6277 gnd.n6276 585
R8220 gnd.n653 gnd.n652 585
R8221 gnd.n652 gnd.n651 585
R8222 gnd.n6283 gnd.n6282 585
R8223 gnd.n6284 gnd.n6283 585
R8224 gnd.n650 gnd.n649 585
R8225 gnd.n6285 gnd.n650 585
R8226 gnd.n6288 gnd.n6287 585
R8227 gnd.n6287 gnd.n6286 585
R8228 gnd.n647 gnd.n646 585
R8229 gnd.n646 gnd.n645 585
R8230 gnd.n6293 gnd.n6292 585
R8231 gnd.n6294 gnd.n6293 585
R8232 gnd.n644 gnd.n643 585
R8233 gnd.n6295 gnd.n644 585
R8234 gnd.n6298 gnd.n6297 585
R8235 gnd.n6297 gnd.n6296 585
R8236 gnd.n641 gnd.n640 585
R8237 gnd.n640 gnd.n639 585
R8238 gnd.n6303 gnd.n6302 585
R8239 gnd.n6304 gnd.n6303 585
R8240 gnd.n638 gnd.n637 585
R8241 gnd.n6305 gnd.n638 585
R8242 gnd.n6308 gnd.n6307 585
R8243 gnd.n6307 gnd.n6306 585
R8244 gnd.n635 gnd.n634 585
R8245 gnd.n634 gnd.n633 585
R8246 gnd.n6313 gnd.n6312 585
R8247 gnd.n6314 gnd.n6313 585
R8248 gnd.n632 gnd.n631 585
R8249 gnd.n6315 gnd.n632 585
R8250 gnd.n6318 gnd.n6317 585
R8251 gnd.n6317 gnd.n6316 585
R8252 gnd.n629 gnd.n628 585
R8253 gnd.n628 gnd.n627 585
R8254 gnd.n6323 gnd.n6322 585
R8255 gnd.n6324 gnd.n6323 585
R8256 gnd.n626 gnd.n625 585
R8257 gnd.n6325 gnd.n626 585
R8258 gnd.n6328 gnd.n6327 585
R8259 gnd.n6327 gnd.n6326 585
R8260 gnd.n623 gnd.n622 585
R8261 gnd.n622 gnd.n621 585
R8262 gnd.n6333 gnd.n6332 585
R8263 gnd.n6334 gnd.n6333 585
R8264 gnd.n620 gnd.n619 585
R8265 gnd.n6335 gnd.n620 585
R8266 gnd.n6338 gnd.n6337 585
R8267 gnd.n6337 gnd.n6336 585
R8268 gnd.n617 gnd.n616 585
R8269 gnd.n616 gnd.n615 585
R8270 gnd.n6343 gnd.n6342 585
R8271 gnd.n6344 gnd.n6343 585
R8272 gnd.n614 gnd.n613 585
R8273 gnd.n6345 gnd.n614 585
R8274 gnd.n6348 gnd.n6347 585
R8275 gnd.n6347 gnd.n6346 585
R8276 gnd.n611 gnd.n610 585
R8277 gnd.n610 gnd.n609 585
R8278 gnd.n6353 gnd.n6352 585
R8279 gnd.n6354 gnd.n6353 585
R8280 gnd.n608 gnd.n607 585
R8281 gnd.n6355 gnd.n608 585
R8282 gnd.n6358 gnd.n6357 585
R8283 gnd.n6357 gnd.n6356 585
R8284 gnd.n605 gnd.n604 585
R8285 gnd.n604 gnd.n603 585
R8286 gnd.n6363 gnd.n6362 585
R8287 gnd.n6364 gnd.n6363 585
R8288 gnd.n602 gnd.n601 585
R8289 gnd.n6365 gnd.n602 585
R8290 gnd.n6368 gnd.n6367 585
R8291 gnd.n6367 gnd.n6366 585
R8292 gnd.n599 gnd.n598 585
R8293 gnd.n598 gnd.n597 585
R8294 gnd.n6373 gnd.n6372 585
R8295 gnd.n6374 gnd.n6373 585
R8296 gnd.n596 gnd.n595 585
R8297 gnd.n6375 gnd.n596 585
R8298 gnd.n6378 gnd.n6377 585
R8299 gnd.n6377 gnd.n6376 585
R8300 gnd.n593 gnd.n592 585
R8301 gnd.n592 gnd.n591 585
R8302 gnd.n6383 gnd.n6382 585
R8303 gnd.n6384 gnd.n6383 585
R8304 gnd.n590 gnd.n589 585
R8305 gnd.n6385 gnd.n590 585
R8306 gnd.n6388 gnd.n6387 585
R8307 gnd.n6387 gnd.n6386 585
R8308 gnd.n587 gnd.n586 585
R8309 gnd.n586 gnd.n585 585
R8310 gnd.n6393 gnd.n6392 585
R8311 gnd.n6394 gnd.n6393 585
R8312 gnd.n584 gnd.n583 585
R8313 gnd.n6395 gnd.n584 585
R8314 gnd.n6398 gnd.n6397 585
R8315 gnd.n6397 gnd.n6396 585
R8316 gnd.n581 gnd.n580 585
R8317 gnd.n580 gnd.n579 585
R8318 gnd.n6403 gnd.n6402 585
R8319 gnd.n6404 gnd.n6403 585
R8320 gnd.n578 gnd.n577 585
R8321 gnd.n6405 gnd.n578 585
R8322 gnd.n6408 gnd.n6407 585
R8323 gnd.n6407 gnd.n6406 585
R8324 gnd.n575 gnd.n574 585
R8325 gnd.n574 gnd.n573 585
R8326 gnd.n6413 gnd.n6412 585
R8327 gnd.n6414 gnd.n6413 585
R8328 gnd.n572 gnd.n571 585
R8329 gnd.n6415 gnd.n572 585
R8330 gnd.n6418 gnd.n6417 585
R8331 gnd.n6417 gnd.n6416 585
R8332 gnd.n569 gnd.n568 585
R8333 gnd.n568 gnd.n567 585
R8334 gnd.n6423 gnd.n6422 585
R8335 gnd.n6424 gnd.n6423 585
R8336 gnd.n566 gnd.n565 585
R8337 gnd.n6425 gnd.n566 585
R8338 gnd.n6428 gnd.n6427 585
R8339 gnd.n6427 gnd.n6426 585
R8340 gnd.n563 gnd.n562 585
R8341 gnd.n562 gnd.n561 585
R8342 gnd.n6433 gnd.n6432 585
R8343 gnd.n6434 gnd.n6433 585
R8344 gnd.n560 gnd.n559 585
R8345 gnd.n6435 gnd.n560 585
R8346 gnd.n6438 gnd.n6437 585
R8347 gnd.n6437 gnd.n6436 585
R8348 gnd.n557 gnd.n556 585
R8349 gnd.n556 gnd.n555 585
R8350 gnd.n6443 gnd.n6442 585
R8351 gnd.n6444 gnd.n6443 585
R8352 gnd.n554 gnd.n553 585
R8353 gnd.n6445 gnd.n554 585
R8354 gnd.n6448 gnd.n6447 585
R8355 gnd.n6447 gnd.n6446 585
R8356 gnd.n551 gnd.n550 585
R8357 gnd.n550 gnd.n549 585
R8358 gnd.n6453 gnd.n6452 585
R8359 gnd.n6454 gnd.n6453 585
R8360 gnd.n548 gnd.n547 585
R8361 gnd.n6455 gnd.n548 585
R8362 gnd.n6458 gnd.n6457 585
R8363 gnd.n6457 gnd.n6456 585
R8364 gnd.n545 gnd.n544 585
R8365 gnd.n544 gnd.n543 585
R8366 gnd.n6463 gnd.n6462 585
R8367 gnd.n6464 gnd.n6463 585
R8368 gnd.n542 gnd.n541 585
R8369 gnd.n6465 gnd.n542 585
R8370 gnd.n6468 gnd.n6467 585
R8371 gnd.n6467 gnd.n6466 585
R8372 gnd.n539 gnd.n538 585
R8373 gnd.n538 gnd.n537 585
R8374 gnd.n6473 gnd.n6472 585
R8375 gnd.n6474 gnd.n6473 585
R8376 gnd.n536 gnd.n535 585
R8377 gnd.n6475 gnd.n536 585
R8378 gnd.n6478 gnd.n6477 585
R8379 gnd.n6477 gnd.n6476 585
R8380 gnd.n533 gnd.n532 585
R8381 gnd.n532 gnd.n531 585
R8382 gnd.n6483 gnd.n6482 585
R8383 gnd.n6484 gnd.n6483 585
R8384 gnd.n530 gnd.n529 585
R8385 gnd.n6485 gnd.n530 585
R8386 gnd.n6488 gnd.n6487 585
R8387 gnd.n6487 gnd.n6486 585
R8388 gnd.n527 gnd.n526 585
R8389 gnd.n526 gnd.n525 585
R8390 gnd.n6494 gnd.n6493 585
R8391 gnd.n6495 gnd.n6494 585
R8392 gnd.n524 gnd.n523 585
R8393 gnd.n6496 gnd.n524 585
R8394 gnd.n6499 gnd.n6498 585
R8395 gnd.n6498 gnd.n6497 585
R8396 gnd.n6500 gnd.n521 585
R8397 gnd.n521 gnd.n520 585
R8398 gnd.n396 gnd.n395 585
R8399 gnd.n6707 gnd.n395 585
R8400 gnd.n6710 gnd.n6709 585
R8401 gnd.n6709 gnd.n6708 585
R8402 gnd.n399 gnd.n398 585
R8403 gnd.n6706 gnd.n399 585
R8404 gnd.n6704 gnd.n6703 585
R8405 gnd.n6705 gnd.n6704 585
R8406 gnd.n402 gnd.n401 585
R8407 gnd.n401 gnd.n400 585
R8408 gnd.n6699 gnd.n6698 585
R8409 gnd.n6698 gnd.n6697 585
R8410 gnd.n405 gnd.n404 585
R8411 gnd.n6696 gnd.n405 585
R8412 gnd.n6694 gnd.n6693 585
R8413 gnd.n6695 gnd.n6694 585
R8414 gnd.n408 gnd.n407 585
R8415 gnd.n407 gnd.n406 585
R8416 gnd.n6689 gnd.n6688 585
R8417 gnd.n6688 gnd.n6687 585
R8418 gnd.n411 gnd.n410 585
R8419 gnd.n6686 gnd.n411 585
R8420 gnd.n6684 gnd.n6683 585
R8421 gnd.n6685 gnd.n6684 585
R8422 gnd.n414 gnd.n413 585
R8423 gnd.n413 gnd.n412 585
R8424 gnd.n6679 gnd.n6678 585
R8425 gnd.n6678 gnd.n6677 585
R8426 gnd.n417 gnd.n416 585
R8427 gnd.n6676 gnd.n417 585
R8428 gnd.n6674 gnd.n6673 585
R8429 gnd.n6675 gnd.n6674 585
R8430 gnd.n420 gnd.n419 585
R8431 gnd.n419 gnd.n418 585
R8432 gnd.n6669 gnd.n6668 585
R8433 gnd.n6668 gnd.n6667 585
R8434 gnd.n423 gnd.n422 585
R8435 gnd.n6666 gnd.n423 585
R8436 gnd.n6664 gnd.n6663 585
R8437 gnd.n6665 gnd.n6664 585
R8438 gnd.n426 gnd.n425 585
R8439 gnd.n425 gnd.n424 585
R8440 gnd.n6659 gnd.n6658 585
R8441 gnd.n6658 gnd.n6657 585
R8442 gnd.n429 gnd.n428 585
R8443 gnd.n6656 gnd.n429 585
R8444 gnd.n6654 gnd.n6653 585
R8445 gnd.n6655 gnd.n6654 585
R8446 gnd.n432 gnd.n431 585
R8447 gnd.n431 gnd.n430 585
R8448 gnd.n6649 gnd.n6648 585
R8449 gnd.n6648 gnd.n6647 585
R8450 gnd.n435 gnd.n434 585
R8451 gnd.n6646 gnd.n435 585
R8452 gnd.n6644 gnd.n6643 585
R8453 gnd.n6645 gnd.n6644 585
R8454 gnd.n438 gnd.n437 585
R8455 gnd.n437 gnd.n436 585
R8456 gnd.n6639 gnd.n6638 585
R8457 gnd.n6638 gnd.n6637 585
R8458 gnd.n441 gnd.n440 585
R8459 gnd.n6636 gnd.n441 585
R8460 gnd.n6634 gnd.n6633 585
R8461 gnd.n6635 gnd.n6634 585
R8462 gnd.n444 gnd.n443 585
R8463 gnd.n443 gnd.n442 585
R8464 gnd.n6629 gnd.n6628 585
R8465 gnd.n6628 gnd.n6627 585
R8466 gnd.n447 gnd.n446 585
R8467 gnd.n6626 gnd.n447 585
R8468 gnd.n6624 gnd.n6623 585
R8469 gnd.n6625 gnd.n6624 585
R8470 gnd.n450 gnd.n449 585
R8471 gnd.n449 gnd.n448 585
R8472 gnd.n6619 gnd.n6618 585
R8473 gnd.n6618 gnd.n6617 585
R8474 gnd.n453 gnd.n452 585
R8475 gnd.n6616 gnd.n453 585
R8476 gnd.n6614 gnd.n6613 585
R8477 gnd.n6615 gnd.n6614 585
R8478 gnd.n456 gnd.n455 585
R8479 gnd.n455 gnd.n454 585
R8480 gnd.n6609 gnd.n6608 585
R8481 gnd.n6608 gnd.n6607 585
R8482 gnd.n459 gnd.n458 585
R8483 gnd.n6606 gnd.n459 585
R8484 gnd.n6604 gnd.n6603 585
R8485 gnd.n6605 gnd.n6604 585
R8486 gnd.n462 gnd.n461 585
R8487 gnd.n461 gnd.n460 585
R8488 gnd.n6599 gnd.n6598 585
R8489 gnd.n6598 gnd.n6597 585
R8490 gnd.n465 gnd.n464 585
R8491 gnd.n6596 gnd.n465 585
R8492 gnd.n6594 gnd.n6593 585
R8493 gnd.n6595 gnd.n6594 585
R8494 gnd.n468 gnd.n467 585
R8495 gnd.n467 gnd.n466 585
R8496 gnd.n6589 gnd.n6588 585
R8497 gnd.n6588 gnd.n6587 585
R8498 gnd.n471 gnd.n470 585
R8499 gnd.n6586 gnd.n471 585
R8500 gnd.n6584 gnd.n6583 585
R8501 gnd.n6585 gnd.n6584 585
R8502 gnd.n474 gnd.n473 585
R8503 gnd.n473 gnd.n472 585
R8504 gnd.n6579 gnd.n6578 585
R8505 gnd.n6578 gnd.n6577 585
R8506 gnd.n477 gnd.n476 585
R8507 gnd.n6576 gnd.n477 585
R8508 gnd.n6574 gnd.n6573 585
R8509 gnd.n6575 gnd.n6574 585
R8510 gnd.n480 gnd.n479 585
R8511 gnd.n479 gnd.n478 585
R8512 gnd.n6569 gnd.n6568 585
R8513 gnd.n6568 gnd.n6567 585
R8514 gnd.n483 gnd.n482 585
R8515 gnd.n6566 gnd.n483 585
R8516 gnd.n6564 gnd.n6563 585
R8517 gnd.n6565 gnd.n6564 585
R8518 gnd.n486 gnd.n485 585
R8519 gnd.n485 gnd.n484 585
R8520 gnd.n6559 gnd.n6558 585
R8521 gnd.n6558 gnd.n6557 585
R8522 gnd.n489 gnd.n488 585
R8523 gnd.n6556 gnd.n489 585
R8524 gnd.n6554 gnd.n6553 585
R8525 gnd.n6555 gnd.n6554 585
R8526 gnd.n492 gnd.n491 585
R8527 gnd.n491 gnd.n490 585
R8528 gnd.n6549 gnd.n6548 585
R8529 gnd.n6548 gnd.n6547 585
R8530 gnd.n495 gnd.n494 585
R8531 gnd.n6546 gnd.n495 585
R8532 gnd.n6544 gnd.n6543 585
R8533 gnd.n6545 gnd.n6544 585
R8534 gnd.n498 gnd.n497 585
R8535 gnd.n497 gnd.n496 585
R8536 gnd.n6539 gnd.n6538 585
R8537 gnd.n6538 gnd.n6537 585
R8538 gnd.n501 gnd.n500 585
R8539 gnd.n6536 gnd.n501 585
R8540 gnd.n6534 gnd.n6533 585
R8541 gnd.n6535 gnd.n6534 585
R8542 gnd.n504 gnd.n503 585
R8543 gnd.n503 gnd.n502 585
R8544 gnd.n6529 gnd.n6528 585
R8545 gnd.n6528 gnd.n6527 585
R8546 gnd.n507 gnd.n506 585
R8547 gnd.n6526 gnd.n507 585
R8548 gnd.n6524 gnd.n6523 585
R8549 gnd.n6525 gnd.n6524 585
R8550 gnd.n510 gnd.n509 585
R8551 gnd.n509 gnd.n508 585
R8552 gnd.n6519 gnd.n6518 585
R8553 gnd.n6518 gnd.n6517 585
R8554 gnd.n513 gnd.n512 585
R8555 gnd.n6516 gnd.n513 585
R8556 gnd.n6514 gnd.n6513 585
R8557 gnd.n6515 gnd.n6514 585
R8558 gnd.n516 gnd.n515 585
R8559 gnd.n515 gnd.n514 585
R8560 gnd.n6509 gnd.n6508 585
R8561 gnd.n6508 gnd.n6507 585
R8562 gnd.n519 gnd.n518 585
R8563 gnd.n6506 gnd.n519 585
R8564 gnd.n6504 gnd.n6503 585
R8565 gnd.n6505 gnd.n6504 585
R8566 gnd.n967 gnd.n966 585
R8567 gnd.n4468 gnd.n967 585
R8568 gnd.n5961 gnd.n5960 585
R8569 gnd.n5960 gnd.n5959 585
R8570 gnd.n5962 gnd.n962 585
R8571 gnd.n4372 gnd.n962 585
R8572 gnd.n5964 gnd.n5963 585
R8573 gnd.n5965 gnd.n5964 585
R8574 gnd.n946 gnd.n945 585
R8575 gnd.n4362 gnd.n946 585
R8576 gnd.n5973 gnd.n5972 585
R8577 gnd.n5972 gnd.n5971 585
R8578 gnd.n5974 gnd.n941 585
R8579 gnd.n4355 gnd.n941 585
R8580 gnd.n5976 gnd.n5975 585
R8581 gnd.n5977 gnd.n5976 585
R8582 gnd.n927 gnd.n926 585
R8583 gnd.n4347 gnd.n927 585
R8584 gnd.n5985 gnd.n5984 585
R8585 gnd.n5984 gnd.n5983 585
R8586 gnd.n5986 gnd.n922 585
R8587 gnd.n4340 gnd.n922 585
R8588 gnd.n5988 gnd.n5987 585
R8589 gnd.n5989 gnd.n5988 585
R8590 gnd.n906 gnd.n905 585
R8591 gnd.n4283 gnd.n906 585
R8592 gnd.n5997 gnd.n5996 585
R8593 gnd.n5996 gnd.n5995 585
R8594 gnd.n5998 gnd.n900 585
R8595 gnd.n4294 gnd.n900 585
R8596 gnd.n6000 gnd.n5999 585
R8597 gnd.n6001 gnd.n6000 585
R8598 gnd.n901 gnd.n899 585
R8599 gnd.n4274 gnd.n899 585
R8600 gnd.n4249 gnd.n887 585
R8601 gnd.n6007 gnd.n887 585
R8602 gnd.n4251 gnd.n4250 585
R8603 gnd.n4250 gnd.n883 585
R8604 gnd.n4252 gnd.n2080 585
R8605 gnd.n4265 gnd.n2080 585
R8606 gnd.n4253 gnd.n2091 585
R8607 gnd.n2091 gnd.n2089 585
R8608 gnd.n4255 gnd.n4254 585
R8609 gnd.n4256 gnd.n4255 585
R8610 gnd.n2092 gnd.n2090 585
R8611 gnd.n2090 gnd.n2086 585
R8612 gnd.n4225 gnd.n2101 585
R8613 gnd.n4237 gnd.n2101 585
R8614 gnd.n4226 gnd.n2110 585
R8615 gnd.n2110 gnd.n2099 585
R8616 gnd.n4228 gnd.n4227 585
R8617 gnd.n4229 gnd.n4228 585
R8618 gnd.n2111 gnd.n2109 585
R8619 gnd.n4218 gnd.n2109 585
R8620 gnd.n4181 gnd.n4180 585
R8621 gnd.n4180 gnd.n2116 585
R8622 gnd.n4182 gnd.n2125 585
R8623 gnd.n4196 gnd.n2125 585
R8624 gnd.n4183 gnd.n2135 585
R8625 gnd.n2135 gnd.n2123 585
R8626 gnd.n4185 gnd.n4184 585
R8627 gnd.n4186 gnd.n4185 585
R8628 gnd.n2136 gnd.n2134 585
R8629 gnd.n4171 gnd.n2134 585
R8630 gnd.n4146 gnd.n4145 585
R8631 gnd.n4145 gnd.n2142 585
R8632 gnd.n4147 gnd.n2149 585
R8633 gnd.n4161 gnd.n2149 585
R8634 gnd.n4148 gnd.n2160 585
R8635 gnd.n2160 gnd.n2158 585
R8636 gnd.n4150 gnd.n4149 585
R8637 gnd.n4151 gnd.n4150 585
R8638 gnd.n2161 gnd.n2159 585
R8639 gnd.n4136 gnd.n2159 585
R8640 gnd.n4111 gnd.n4110 585
R8641 gnd.n4110 gnd.n2167 585
R8642 gnd.n4112 gnd.n2174 585
R8643 gnd.n4126 gnd.n2174 585
R8644 gnd.n4113 gnd.n2186 585
R8645 gnd.n2186 gnd.n2184 585
R8646 gnd.n4115 gnd.n4114 585
R8647 gnd.n4116 gnd.n4115 585
R8648 gnd.n2187 gnd.n2185 585
R8649 gnd.n2185 gnd.n2181 585
R8650 gnd.n4088 gnd.n2195 585
R8651 gnd.n4100 gnd.n2195 585
R8652 gnd.n4089 gnd.n2205 585
R8653 gnd.n2205 gnd.n2193 585
R8654 gnd.n4091 gnd.n4090 585
R8655 gnd.n4092 gnd.n4091 585
R8656 gnd.n2206 gnd.n2204 585
R8657 gnd.n2204 gnd.n2201 585
R8658 gnd.n4068 gnd.n2212 585
R8659 gnd.n4080 gnd.n2212 585
R8660 gnd.n4069 gnd.n2223 585
R8661 gnd.n2223 gnd.n2221 585
R8662 gnd.n4071 gnd.n4070 585
R8663 gnd.n4072 gnd.n4071 585
R8664 gnd.n2224 gnd.n2222 585
R8665 gnd.n2222 gnd.n2218 585
R8666 gnd.n4048 gnd.n2231 585
R8667 gnd.n4060 gnd.n2231 585
R8668 gnd.n4049 gnd.n2241 585
R8669 gnd.n2241 gnd.n2229 585
R8670 gnd.n4051 gnd.n4050 585
R8671 gnd.n4052 gnd.n4051 585
R8672 gnd.n2242 gnd.n2240 585
R8673 gnd.n2240 gnd.n2237 585
R8674 gnd.n3919 gnd.n3918 585
R8675 gnd.n3917 gnd.n3916 585
R8676 gnd.n3915 gnd.n3914 585
R8677 gnd.n3913 gnd.n3912 585
R8678 gnd.n3911 gnd.n3910 585
R8679 gnd.n3909 gnd.n3908 585
R8680 gnd.n3907 gnd.n3906 585
R8681 gnd.n3905 gnd.n3904 585
R8682 gnd.n3903 gnd.n3902 585
R8683 gnd.n3901 gnd.n3900 585
R8684 gnd.n3899 gnd.n3898 585
R8685 gnd.n3897 gnd.n3896 585
R8686 gnd.n3895 gnd.n3894 585
R8687 gnd.n3893 gnd.n3892 585
R8688 gnd.n3891 gnd.n3890 585
R8689 gnd.n3889 gnd.n3888 585
R8690 gnd.n3887 gnd.n3886 585
R8691 gnd.n3846 gnd.n3843 585
R8692 gnd.n3882 gnd.n3762 585
R8693 gnd.n4039 gnd.n3762 585
R8694 gnd.n4471 gnd.n4470 585
R8695 gnd.n4449 gnd.n1850 585
R8696 gnd.n4451 gnd.n4450 585
R8697 gnd.n4448 gnd.n1883 585
R8698 gnd.n1882 gnd.n1881 585
R8699 gnd.n4438 gnd.n4437 585
R8700 gnd.n4436 gnd.n4435 585
R8701 gnd.n4424 gnd.n1889 585
R8702 gnd.n4426 gnd.n4425 585
R8703 gnd.n4423 gnd.n1895 585
R8704 gnd.n1894 gnd.n1893 585
R8705 gnd.n4414 gnd.n4413 585
R8706 gnd.n4412 gnd.n4411 585
R8707 gnd.n4400 gnd.n1901 585
R8708 gnd.n4402 gnd.n4401 585
R8709 gnd.n4399 gnd.n1907 585
R8710 gnd.n1906 gnd.n1905 585
R8711 gnd.n4390 gnd.n4389 585
R8712 gnd.n4388 gnd.n979 585
R8713 gnd.n5951 gnd.n979 585
R8714 gnd.n4469 gnd.n1851 585
R8715 gnd.n4469 gnd.n4468 585
R8716 gnd.n2053 gnd.n970 585
R8717 gnd.n5959 gnd.n970 585
R8718 gnd.n4371 gnd.n4370 585
R8719 gnd.n4372 gnd.n4371 585
R8720 gnd.n2052 gnd.n960 585
R8721 gnd.n5965 gnd.n960 585
R8722 gnd.n4364 gnd.n4363 585
R8723 gnd.n4363 gnd.n4362 585
R8724 gnd.n2055 gnd.n949 585
R8725 gnd.n5971 gnd.n949 585
R8726 gnd.n4354 gnd.n4353 585
R8727 gnd.n4355 gnd.n4354 585
R8728 gnd.n2058 gnd.n940 585
R8729 gnd.n5977 gnd.n940 585
R8730 gnd.n4349 gnd.n4348 585
R8731 gnd.n4348 gnd.n4347 585
R8732 gnd.n2060 gnd.n929 585
R8733 gnd.n5983 gnd.n929 585
R8734 gnd.n4286 gnd.n2062 585
R8735 gnd.n4340 gnd.n2062 585
R8736 gnd.n4287 gnd.n920 585
R8737 gnd.n5989 gnd.n920 585
R8738 gnd.n4288 gnd.n4284 585
R8739 gnd.n4284 gnd.n4283 585
R8740 gnd.n2070 gnd.n909 585
R8741 gnd.n5995 gnd.n909 585
R8742 gnd.n4293 gnd.n4292 585
R8743 gnd.n4294 gnd.n4293 585
R8744 gnd.n2069 gnd.n898 585
R8745 gnd.n6001 gnd.n898 585
R8746 gnd.n4273 gnd.n4272 585
R8747 gnd.n4274 gnd.n4273 585
R8748 gnd.n2075 gnd.n885 585
R8749 gnd.n6007 gnd.n885 585
R8750 gnd.n4268 gnd.n4267 585
R8751 gnd.n4267 gnd.n883 585
R8752 gnd.n4266 gnd.n2077 585
R8753 gnd.n4266 gnd.n4265 585
R8754 gnd.n4206 gnd.n2078 585
R8755 gnd.n2089 gnd.n2078 585
R8756 gnd.n4205 gnd.n2088 585
R8757 gnd.n4256 gnd.n2088 585
R8758 gnd.n4210 gnd.n4204 585
R8759 gnd.n4204 gnd.n2086 585
R8760 gnd.n4211 gnd.n2100 585
R8761 gnd.n4237 gnd.n2100 585
R8762 gnd.n4212 gnd.n4203 585
R8763 gnd.n4203 gnd.n2099 585
R8764 gnd.n2119 gnd.n2108 585
R8765 gnd.n4229 gnd.n2108 585
R8766 gnd.n4217 gnd.n4216 585
R8767 gnd.n4218 gnd.n4217 585
R8768 gnd.n2118 gnd.n2117 585
R8769 gnd.n2117 gnd.n2116 585
R8770 gnd.n4198 gnd.n4197 585
R8771 gnd.n4197 gnd.n4196 585
R8772 gnd.n2122 gnd.n2121 585
R8773 gnd.n2123 gnd.n2122 585
R8774 gnd.n4168 gnd.n2133 585
R8775 gnd.n4186 gnd.n2133 585
R8776 gnd.n4170 gnd.n4169 585
R8777 gnd.n4171 gnd.n4170 585
R8778 gnd.n2144 gnd.n2143 585
R8779 gnd.n2143 gnd.n2142 585
R8780 gnd.n4163 gnd.n4162 585
R8781 gnd.n4162 gnd.n4161 585
R8782 gnd.n2147 gnd.n2146 585
R8783 gnd.n2158 gnd.n2147 585
R8784 gnd.n4133 gnd.n2157 585
R8785 gnd.n4151 gnd.n2157 585
R8786 gnd.n4135 gnd.n4134 585
R8787 gnd.n4136 gnd.n4135 585
R8788 gnd.n2169 gnd.n2168 585
R8789 gnd.n2168 gnd.n2167 585
R8790 gnd.n4128 gnd.n4127 585
R8791 gnd.n4127 gnd.n4126 585
R8792 gnd.n2172 gnd.n2171 585
R8793 gnd.n2184 gnd.n2172 585
R8794 gnd.n3860 gnd.n2183 585
R8795 gnd.n4116 gnd.n2183 585
R8796 gnd.n3862 gnd.n3861 585
R8797 gnd.n3861 gnd.n2181 585
R8798 gnd.n3863 gnd.n2194 585
R8799 gnd.n4100 gnd.n2194 585
R8800 gnd.n3865 gnd.n3864 585
R8801 gnd.n3864 gnd.n2193 585
R8802 gnd.n3866 gnd.n2203 585
R8803 gnd.n4092 gnd.n2203 585
R8804 gnd.n3868 gnd.n3867 585
R8805 gnd.n3867 gnd.n2201 585
R8806 gnd.n3869 gnd.n2211 585
R8807 gnd.n4080 gnd.n2211 585
R8808 gnd.n3871 gnd.n3870 585
R8809 gnd.n3870 gnd.n2221 585
R8810 gnd.n3872 gnd.n2220 585
R8811 gnd.n4072 gnd.n2220 585
R8812 gnd.n3874 gnd.n3873 585
R8813 gnd.n3873 gnd.n2218 585
R8814 gnd.n3875 gnd.n2230 585
R8815 gnd.n4060 gnd.n2230 585
R8816 gnd.n3877 gnd.n3876 585
R8817 gnd.n3876 gnd.n2229 585
R8818 gnd.n3878 gnd.n2239 585
R8819 gnd.n4052 gnd.n2239 585
R8820 gnd.n3880 gnd.n3879 585
R8821 gnd.n3879 gnd.n2237 585
R8822 gnd.n3633 gnd.n3632 585
R8823 gnd.n3634 gnd.n3633 585
R8824 gnd.n2324 gnd.n2323 585
R8825 gnd.n2330 gnd.n2323 585
R8826 gnd.n3608 gnd.n2342 585
R8827 gnd.n2342 gnd.n2329 585
R8828 gnd.n3610 gnd.n3609 585
R8829 gnd.n3611 gnd.n3610 585
R8830 gnd.n2343 gnd.n2341 585
R8831 gnd.n2341 gnd.n2337 585
R8832 gnd.n3342 gnd.n3341 585
R8833 gnd.n3341 gnd.n3340 585
R8834 gnd.n2348 gnd.n2347 585
R8835 gnd.n3311 gnd.n2348 585
R8836 gnd.n3331 gnd.n3330 585
R8837 gnd.n3330 gnd.n3329 585
R8838 gnd.n2355 gnd.n2354 585
R8839 gnd.n3317 gnd.n2355 585
R8840 gnd.n3287 gnd.n2375 585
R8841 gnd.n2375 gnd.n2374 585
R8842 gnd.n3289 gnd.n3288 585
R8843 gnd.n3290 gnd.n3289 585
R8844 gnd.n2376 gnd.n2373 585
R8845 gnd.n2384 gnd.n2373 585
R8846 gnd.n3265 gnd.n2396 585
R8847 gnd.n2396 gnd.n2383 585
R8848 gnd.n3267 gnd.n3266 585
R8849 gnd.n3268 gnd.n3267 585
R8850 gnd.n2397 gnd.n2395 585
R8851 gnd.n2395 gnd.n2391 585
R8852 gnd.n3253 gnd.n3252 585
R8853 gnd.n3252 gnd.n3251 585
R8854 gnd.n2402 gnd.n2401 585
R8855 gnd.n2412 gnd.n2402 585
R8856 gnd.n3242 gnd.n3241 585
R8857 gnd.n3241 gnd.n3240 585
R8858 gnd.n2409 gnd.n2408 585
R8859 gnd.n3228 gnd.n2409 585
R8860 gnd.n3202 gnd.n2430 585
R8861 gnd.n2430 gnd.n2419 585
R8862 gnd.n3204 gnd.n3203 585
R8863 gnd.n3205 gnd.n3204 585
R8864 gnd.n2431 gnd.n2429 585
R8865 gnd.n2439 gnd.n2429 585
R8866 gnd.n3180 gnd.n2451 585
R8867 gnd.n2451 gnd.n2438 585
R8868 gnd.n3182 gnd.n3181 585
R8869 gnd.n3183 gnd.n3182 585
R8870 gnd.n2452 gnd.n2450 585
R8871 gnd.n2450 gnd.n2446 585
R8872 gnd.n3168 gnd.n3167 585
R8873 gnd.n3167 gnd.n3166 585
R8874 gnd.n2457 gnd.n2456 585
R8875 gnd.n2466 gnd.n2457 585
R8876 gnd.n3157 gnd.n3156 585
R8877 gnd.n3156 gnd.n3155 585
R8878 gnd.n2464 gnd.n2463 585
R8879 gnd.n3143 gnd.n2464 585
R8880 gnd.n2581 gnd.n2580 585
R8881 gnd.n2581 gnd.n2473 585
R8882 gnd.n3100 gnd.n3099 585
R8883 gnd.n3099 gnd.n3098 585
R8884 gnd.n3101 gnd.n2575 585
R8885 gnd.n2586 gnd.n2575 585
R8886 gnd.n3103 gnd.n3102 585
R8887 gnd.n3104 gnd.n3103 585
R8888 gnd.n2576 gnd.n2574 585
R8889 gnd.n2599 gnd.n2574 585
R8890 gnd.n2559 gnd.n2558 585
R8891 gnd.n2562 gnd.n2559 585
R8892 gnd.n3114 gnd.n3113 585
R8893 gnd.n3113 gnd.n3112 585
R8894 gnd.n3115 gnd.n2553 585
R8895 gnd.n3074 gnd.n2553 585
R8896 gnd.n3117 gnd.n3116 585
R8897 gnd.n3118 gnd.n3117 585
R8898 gnd.n2554 gnd.n2552 585
R8899 gnd.n2613 gnd.n2552 585
R8900 gnd.n3066 gnd.n3065 585
R8901 gnd.n3065 gnd.n3064 585
R8902 gnd.n2610 gnd.n2609 585
R8903 gnd.n3048 gnd.n2610 585
R8904 gnd.n3035 gnd.n2629 585
R8905 gnd.n2629 gnd.n2628 585
R8906 gnd.n3037 gnd.n3036 585
R8907 gnd.n3038 gnd.n3037 585
R8908 gnd.n2630 gnd.n2627 585
R8909 gnd.n2636 gnd.n2627 585
R8910 gnd.n3016 gnd.n3015 585
R8911 gnd.n3017 gnd.n3016 585
R8912 gnd.n2647 gnd.n2646 585
R8913 gnd.n2646 gnd.n2642 585
R8914 gnd.n3006 gnd.n3005 585
R8915 gnd.n3007 gnd.n3006 585
R8916 gnd.n2657 gnd.n2656 585
R8917 gnd.n2662 gnd.n2656 585
R8918 gnd.n2984 gnd.n2675 585
R8919 gnd.n2675 gnd.n2661 585
R8920 gnd.n2986 gnd.n2985 585
R8921 gnd.n2987 gnd.n2986 585
R8922 gnd.n2676 gnd.n2674 585
R8923 gnd.n2674 gnd.n2670 585
R8924 gnd.n2975 gnd.n2974 585
R8925 gnd.n2976 gnd.n2975 585
R8926 gnd.n2683 gnd.n2682 585
R8927 gnd.n2687 gnd.n2682 585
R8928 gnd.n2952 gnd.n2704 585
R8929 gnd.n2704 gnd.n2686 585
R8930 gnd.n2954 gnd.n2953 585
R8931 gnd.n2955 gnd.n2954 585
R8932 gnd.n2705 gnd.n2703 585
R8933 gnd.n2703 gnd.n2694 585
R8934 gnd.n2947 gnd.n2946 585
R8935 gnd.n2946 gnd.n2945 585
R8936 gnd.n2752 gnd.n2751 585
R8937 gnd.n2753 gnd.n2752 585
R8938 gnd.n2906 gnd.n2905 585
R8939 gnd.n2907 gnd.n2906 585
R8940 gnd.n2762 gnd.n2761 585
R8941 gnd.n2761 gnd.n2760 585
R8942 gnd.n2901 gnd.n2900 585
R8943 gnd.n2900 gnd.n2899 585
R8944 gnd.n2765 gnd.n2764 585
R8945 gnd.n2766 gnd.n2765 585
R8946 gnd.n2890 gnd.n2889 585
R8947 gnd.n2891 gnd.n2890 585
R8948 gnd.n2773 gnd.n2772 585
R8949 gnd.n2882 gnd.n2772 585
R8950 gnd.n2885 gnd.n2884 585
R8951 gnd.n2884 gnd.n2883 585
R8952 gnd.n2776 gnd.n2775 585
R8953 gnd.n2777 gnd.n2776 585
R8954 gnd.n2871 gnd.n2870 585
R8955 gnd.n2869 gnd.n2795 585
R8956 gnd.n2868 gnd.n2794 585
R8957 gnd.n2873 gnd.n2794 585
R8958 gnd.n2867 gnd.n2866 585
R8959 gnd.n2865 gnd.n2864 585
R8960 gnd.n2863 gnd.n2862 585
R8961 gnd.n2861 gnd.n2860 585
R8962 gnd.n2859 gnd.n2858 585
R8963 gnd.n2857 gnd.n2856 585
R8964 gnd.n2855 gnd.n2854 585
R8965 gnd.n2853 gnd.n2852 585
R8966 gnd.n2851 gnd.n2850 585
R8967 gnd.n2849 gnd.n2848 585
R8968 gnd.n2847 gnd.n2846 585
R8969 gnd.n2845 gnd.n2844 585
R8970 gnd.n2843 gnd.n2842 585
R8971 gnd.n2841 gnd.n2840 585
R8972 gnd.n2839 gnd.n2838 585
R8973 gnd.n2837 gnd.n2836 585
R8974 gnd.n2835 gnd.n2834 585
R8975 gnd.n2833 gnd.n2832 585
R8976 gnd.n2831 gnd.n2830 585
R8977 gnd.n2829 gnd.n2828 585
R8978 gnd.n2827 gnd.n2826 585
R8979 gnd.n2825 gnd.n2824 585
R8980 gnd.n2782 gnd.n2781 585
R8981 gnd.n2876 gnd.n2875 585
R8982 gnd.n3637 gnd.n3636 585
R8983 gnd.n3639 gnd.n3638 585
R8984 gnd.n3641 gnd.n3640 585
R8985 gnd.n3643 gnd.n3642 585
R8986 gnd.n3645 gnd.n3644 585
R8987 gnd.n3647 gnd.n3646 585
R8988 gnd.n3649 gnd.n3648 585
R8989 gnd.n3651 gnd.n3650 585
R8990 gnd.n3653 gnd.n3652 585
R8991 gnd.n3655 gnd.n3654 585
R8992 gnd.n3657 gnd.n3656 585
R8993 gnd.n3659 gnd.n3658 585
R8994 gnd.n3661 gnd.n3660 585
R8995 gnd.n3663 gnd.n3662 585
R8996 gnd.n3665 gnd.n3664 585
R8997 gnd.n3667 gnd.n3666 585
R8998 gnd.n3669 gnd.n3668 585
R8999 gnd.n3671 gnd.n3670 585
R9000 gnd.n3673 gnd.n3672 585
R9001 gnd.n3675 gnd.n3674 585
R9002 gnd.n3677 gnd.n3676 585
R9003 gnd.n3679 gnd.n3678 585
R9004 gnd.n3681 gnd.n3680 585
R9005 gnd.n3683 gnd.n3682 585
R9006 gnd.n3685 gnd.n3684 585
R9007 gnd.n3686 gnd.n2290 585
R9008 gnd.n3687 gnd.n2248 585
R9009 gnd.n3725 gnd.n2248 585
R9010 gnd.n3635 gnd.n2320 585
R9011 gnd.n3635 gnd.n3634 585
R9012 gnd.n3304 gnd.n2319 585
R9013 gnd.n2330 gnd.n2319 585
R9014 gnd.n3306 gnd.n3305 585
R9015 gnd.n3305 gnd.n2329 585
R9016 gnd.n3307 gnd.n2339 585
R9017 gnd.n3611 gnd.n2339 585
R9018 gnd.n3309 gnd.n3308 585
R9019 gnd.n3308 gnd.n2337 585
R9020 gnd.n3310 gnd.n2350 585
R9021 gnd.n3340 gnd.n2350 585
R9022 gnd.n3313 gnd.n3312 585
R9023 gnd.n3312 gnd.n3311 585
R9024 gnd.n3314 gnd.n2357 585
R9025 gnd.n3329 gnd.n2357 585
R9026 gnd.n3316 gnd.n3315 585
R9027 gnd.n3317 gnd.n3316 585
R9028 gnd.n2367 gnd.n2366 585
R9029 gnd.n2374 gnd.n2366 585
R9030 gnd.n3292 gnd.n3291 585
R9031 gnd.n3291 gnd.n3290 585
R9032 gnd.n2370 gnd.n2369 585
R9033 gnd.n2384 gnd.n2370 585
R9034 gnd.n3218 gnd.n3217 585
R9035 gnd.n3217 gnd.n2383 585
R9036 gnd.n3219 gnd.n2393 585
R9037 gnd.n3268 gnd.n2393 585
R9038 gnd.n3221 gnd.n3220 585
R9039 gnd.n3220 gnd.n2391 585
R9040 gnd.n3222 gnd.n2404 585
R9041 gnd.n3251 gnd.n2404 585
R9042 gnd.n3224 gnd.n3223 585
R9043 gnd.n3223 gnd.n2412 585
R9044 gnd.n3225 gnd.n2411 585
R9045 gnd.n3240 gnd.n2411 585
R9046 gnd.n3227 gnd.n3226 585
R9047 gnd.n3228 gnd.n3227 585
R9048 gnd.n2423 gnd.n2422 585
R9049 gnd.n2422 gnd.n2419 585
R9050 gnd.n3207 gnd.n3206 585
R9051 gnd.n3206 gnd.n3205 585
R9052 gnd.n2426 gnd.n2425 585
R9053 gnd.n2439 gnd.n2426 585
R9054 gnd.n3131 gnd.n3130 585
R9055 gnd.n3130 gnd.n2438 585
R9056 gnd.n3132 gnd.n2448 585
R9057 gnd.n3183 gnd.n2448 585
R9058 gnd.n3134 gnd.n3133 585
R9059 gnd.n3133 gnd.n2446 585
R9060 gnd.n3135 gnd.n2459 585
R9061 gnd.n3166 gnd.n2459 585
R9062 gnd.n3137 gnd.n3136 585
R9063 gnd.n3136 gnd.n2466 585
R9064 gnd.n3138 gnd.n2465 585
R9065 gnd.n3155 gnd.n2465 585
R9066 gnd.n3140 gnd.n3139 585
R9067 gnd.n3143 gnd.n3140 585
R9068 gnd.n2476 gnd.n2475 585
R9069 gnd.n2475 gnd.n2473 585
R9070 gnd.n2583 gnd.n2582 585
R9071 gnd.n3098 gnd.n2582 585
R9072 gnd.n2585 gnd.n2584 585
R9073 gnd.n2586 gnd.n2585 585
R9074 gnd.n2596 gnd.n2572 585
R9075 gnd.n3104 gnd.n2572 585
R9076 gnd.n2598 gnd.n2597 585
R9077 gnd.n2599 gnd.n2598 585
R9078 gnd.n2595 gnd.n2594 585
R9079 gnd.n2595 gnd.n2562 585
R9080 gnd.n2593 gnd.n2560 585
R9081 gnd.n3112 gnd.n2560 585
R9082 gnd.n2549 gnd.n2547 585
R9083 gnd.n3074 gnd.n2549 585
R9084 gnd.n3120 gnd.n3119 585
R9085 gnd.n3119 gnd.n3118 585
R9086 gnd.n2548 gnd.n2546 585
R9087 gnd.n2613 gnd.n2548 585
R9088 gnd.n3045 gnd.n2612 585
R9089 gnd.n3064 gnd.n2612 585
R9090 gnd.n3047 gnd.n3046 585
R9091 gnd.n3048 gnd.n3047 585
R9092 gnd.n2622 gnd.n2621 585
R9093 gnd.n2628 gnd.n2621 585
R9094 gnd.n3040 gnd.n3039 585
R9095 gnd.n3039 gnd.n3038 585
R9096 gnd.n2625 gnd.n2624 585
R9097 gnd.n2636 gnd.n2625 585
R9098 gnd.n2925 gnd.n2644 585
R9099 gnd.n3017 gnd.n2644 585
R9100 gnd.n2927 gnd.n2926 585
R9101 gnd.n2926 gnd.n2642 585
R9102 gnd.n2928 gnd.n2655 585
R9103 gnd.n3007 gnd.n2655 585
R9104 gnd.n2930 gnd.n2929 585
R9105 gnd.n2930 gnd.n2662 585
R9106 gnd.n2932 gnd.n2931 585
R9107 gnd.n2931 gnd.n2661 585
R9108 gnd.n2933 gnd.n2672 585
R9109 gnd.n2987 gnd.n2672 585
R9110 gnd.n2935 gnd.n2934 585
R9111 gnd.n2934 gnd.n2670 585
R9112 gnd.n2936 gnd.n2681 585
R9113 gnd.n2976 gnd.n2681 585
R9114 gnd.n2938 gnd.n2937 585
R9115 gnd.n2938 gnd.n2687 585
R9116 gnd.n2940 gnd.n2939 585
R9117 gnd.n2939 gnd.n2686 585
R9118 gnd.n2941 gnd.n2702 585
R9119 gnd.n2955 gnd.n2702 585
R9120 gnd.n2942 gnd.n2755 585
R9121 gnd.n2755 gnd.n2694 585
R9122 gnd.n2944 gnd.n2943 585
R9123 gnd.n2945 gnd.n2944 585
R9124 gnd.n2756 gnd.n2754 585
R9125 gnd.n2754 gnd.n2753 585
R9126 gnd.n2909 gnd.n2908 585
R9127 gnd.n2908 gnd.n2907 585
R9128 gnd.n2759 gnd.n2758 585
R9129 gnd.n2760 gnd.n2759 585
R9130 gnd.n2898 gnd.n2897 585
R9131 gnd.n2899 gnd.n2898 585
R9132 gnd.n2768 gnd.n2767 585
R9133 gnd.n2767 gnd.n2766 585
R9134 gnd.n2893 gnd.n2892 585
R9135 gnd.n2892 gnd.n2891 585
R9136 gnd.n2771 gnd.n2770 585
R9137 gnd.n2882 gnd.n2771 585
R9138 gnd.n2881 gnd.n2880 585
R9139 gnd.n2883 gnd.n2881 585
R9140 gnd.n2779 gnd.n2778 585
R9141 gnd.n2778 gnd.n2777 585
R9142 gnd.n201 gnd.n200 585
R9143 gnd.n204 gnd.n201 585
R9144 gnd.n7121 gnd.n7120 585
R9145 gnd.n7120 gnd.n7119 585
R9146 gnd.n7122 gnd.n196 585
R9147 gnd.n196 gnd.n195 585
R9148 gnd.n7124 gnd.n7123 585
R9149 gnd.n7125 gnd.n7124 585
R9150 gnd.n181 gnd.n180 585
R9151 gnd.n185 gnd.n181 585
R9152 gnd.n7133 gnd.n7132 585
R9153 gnd.n7132 gnd.n7131 585
R9154 gnd.n7134 gnd.n176 585
R9155 gnd.n182 gnd.n176 585
R9156 gnd.n7136 gnd.n7135 585
R9157 gnd.n7137 gnd.n7136 585
R9158 gnd.n163 gnd.n162 585
R9159 gnd.n166 gnd.n163 585
R9160 gnd.n7145 gnd.n7144 585
R9161 gnd.n7144 gnd.n7143 585
R9162 gnd.n7146 gnd.n158 585
R9163 gnd.n6969 gnd.n158 585
R9164 gnd.n7148 gnd.n7147 585
R9165 gnd.n7149 gnd.n7148 585
R9166 gnd.n143 gnd.n142 585
R9167 gnd.n147 gnd.n143 585
R9168 gnd.n7157 gnd.n7156 585
R9169 gnd.n7156 gnd.n7155 585
R9170 gnd.n7158 gnd.n138 585
R9171 gnd.n144 gnd.n138 585
R9172 gnd.n7160 gnd.n7159 585
R9173 gnd.n7161 gnd.n7160 585
R9174 gnd.n125 gnd.n124 585
R9175 gnd.n128 gnd.n125 585
R9176 gnd.n7169 gnd.n7168 585
R9177 gnd.n7168 gnd.n7167 585
R9178 gnd.n7170 gnd.n120 585
R9179 gnd.n120 gnd.n119 585
R9180 gnd.n7172 gnd.n7171 585
R9181 gnd.n7173 gnd.n7172 585
R9182 gnd.n105 gnd.n104 585
R9183 gnd.n109 gnd.n105 585
R9184 gnd.n7181 gnd.n7180 585
R9185 gnd.n7180 gnd.n7179 585
R9186 gnd.n7182 gnd.n99 585
R9187 gnd.n106 gnd.n99 585
R9188 gnd.n7184 gnd.n7183 585
R9189 gnd.n7185 gnd.n7184 585
R9190 gnd.n100 gnd.n98 585
R9191 gnd.n98 gnd.n86 585
R9192 gnd.n6824 gnd.n87 585
R9193 gnd.n7191 gnd.n87 585
R9194 gnd.n6823 gnd.n6822 585
R9195 gnd.n6822 gnd.n6821 585
R9196 gnd.n312 gnd.n311 585
R9197 gnd.n313 gnd.n312 585
R9198 gnd.n6815 gnd.n6814 585
R9199 gnd.n6814 gnd.n6813 585
R9200 gnd.n318 gnd.n317 585
R9201 gnd.n319 gnd.n318 585
R9202 gnd.n6801 gnd.n6800 585
R9203 gnd.n6802 gnd.n6801 585
R9204 gnd.n332 gnd.n331 585
R9205 gnd.n6793 gnd.n331 585
R9206 gnd.n6764 gnd.n6763 585
R9207 gnd.n6763 gnd.n336 585
R9208 gnd.n6765 gnd.n344 585
R9209 gnd.n6779 gnd.n344 585
R9210 gnd.n6766 gnd.n356 585
R9211 gnd.n356 gnd.n354 585
R9212 gnd.n6768 gnd.n6767 585
R9213 gnd.n6769 gnd.n6768 585
R9214 gnd.n357 gnd.n355 585
R9215 gnd.n6754 gnd.n355 585
R9216 gnd.n6730 gnd.n6729 585
R9217 gnd.n6729 gnd.n6728 585
R9218 gnd.n6731 gnd.n372 585
R9219 gnd.n6745 gnd.n372 585
R9220 gnd.n6732 gnd.n384 585
R9221 gnd.n6722 gnd.n384 585
R9222 gnd.n6734 gnd.n6733 585
R9223 gnd.n6735 gnd.n6734 585
R9224 gnd.n385 gnd.n383 585
R9225 gnd.n5417 gnd.n383 585
R9226 gnd.n5445 gnd.n5444 585
R9227 gnd.n5444 gnd.n5443 585
R9228 gnd.n5446 gnd.n5330 585
R9229 gnd.n5426 gnd.n5330 585
R9230 gnd.n5448 gnd.n5447 585
R9231 gnd.n5449 gnd.n5448 585
R9232 gnd.n5316 gnd.n5315 585
R9233 gnd.n5408 gnd.n5316 585
R9234 gnd.n5457 gnd.n5456 585
R9235 gnd.n5456 gnd.n5455 585
R9236 gnd.n5458 gnd.n5310 585
R9237 gnd.n5400 gnd.n5310 585
R9238 gnd.n5460 gnd.n5459 585
R9239 gnd.n5461 gnd.n5460 585
R9240 gnd.n5311 gnd.n5309 585
R9241 gnd.n5380 gnd.n5309 585
R9242 gnd.n5364 gnd.n5290 585
R9243 gnd.n5467 gnd.n5290 585
R9244 gnd.n5363 gnd.n5362 585
R9245 gnd.n5362 gnd.n5286 585
R9246 gnd.n5361 gnd.n5268 585
R9247 gnd.n5274 gnd.n5268 585
R9248 gnd.n5476 gnd.n5269 585
R9249 gnd.n5476 gnd.n5475 585
R9250 gnd.n5478 gnd.n5477 585
R9251 gnd.n5584 gnd.n5479 585
R9252 gnd.n5583 gnd.n5480 585
R9253 gnd.n5487 gnd.n5481 585
R9254 gnd.n5576 gnd.n5488 585
R9255 gnd.n5575 gnd.n5489 585
R9256 gnd.n5491 gnd.n5490 585
R9257 gnd.n5568 gnd.n5499 585
R9258 gnd.n5567 gnd.n5500 585
R9259 gnd.n5507 gnd.n5501 585
R9260 gnd.n5560 gnd.n5508 585
R9261 gnd.n5559 gnd.n5509 585
R9262 gnd.n5511 gnd.n5510 585
R9263 gnd.n5552 gnd.n5519 585
R9264 gnd.n5551 gnd.n5520 585
R9265 gnd.n5529 gnd.n5521 585
R9266 gnd.n5544 gnd.n5530 585
R9267 gnd.n5543 gnd.n5540 585
R9268 gnd.n5531 gnd.n1277 585
R9269 gnd.n5708 gnd.n1277 585
R9270 gnd.n6951 gnd.n6950 585
R9271 gnd.n6944 gnd.n6897 585
R9272 gnd.n6946 gnd.n6945 585
R9273 gnd.n6943 gnd.n6942 585
R9274 gnd.n6941 gnd.n6940 585
R9275 gnd.n6934 gnd.n6899 585
R9276 gnd.n6936 gnd.n6935 585
R9277 gnd.n6933 gnd.n6932 585
R9278 gnd.n6931 gnd.n6930 585
R9279 gnd.n6924 gnd.n6901 585
R9280 gnd.n6926 gnd.n6925 585
R9281 gnd.n6923 gnd.n6922 585
R9282 gnd.n6921 gnd.n6920 585
R9283 gnd.n6914 gnd.n6903 585
R9284 gnd.n6916 gnd.n6915 585
R9285 gnd.n6913 gnd.n6912 585
R9286 gnd.n6911 gnd.n6910 585
R9287 gnd.n6907 gnd.n6906 585
R9288 gnd.n6905 gnd.n211 585
R9289 gnd.n7111 gnd.n211 585
R9290 gnd.n6953 gnd.n6952 585
R9291 gnd.n6952 gnd.n204 585
R9292 gnd.n6954 gnd.n203 585
R9293 gnd.n7119 gnd.n203 585
R9294 gnd.n6956 gnd.n6955 585
R9295 gnd.n6955 gnd.n195 585
R9296 gnd.n6957 gnd.n194 585
R9297 gnd.n7125 gnd.n194 585
R9298 gnd.n6959 gnd.n6958 585
R9299 gnd.n6958 gnd.n185 585
R9300 gnd.n6960 gnd.n184 585
R9301 gnd.n7131 gnd.n184 585
R9302 gnd.n6962 gnd.n6961 585
R9303 gnd.n6961 gnd.n182 585
R9304 gnd.n6963 gnd.n175 585
R9305 gnd.n7137 gnd.n175 585
R9306 gnd.n6965 gnd.n6964 585
R9307 gnd.n6964 gnd.n166 585
R9308 gnd.n6966 gnd.n165 585
R9309 gnd.n7143 gnd.n165 585
R9310 gnd.n6968 gnd.n6967 585
R9311 gnd.n6969 gnd.n6968 585
R9312 gnd.n6851 gnd.n156 585
R9313 gnd.n7149 gnd.n156 585
R9314 gnd.n6881 gnd.n6880 585
R9315 gnd.n6880 gnd.n147 585
R9316 gnd.n6879 gnd.n146 585
R9317 gnd.n7155 gnd.n146 585
R9318 gnd.n6878 gnd.n6877 585
R9319 gnd.n6877 gnd.n144 585
R9320 gnd.n6853 gnd.n137 585
R9321 gnd.n7161 gnd.n137 585
R9322 gnd.n6873 gnd.n6872 585
R9323 gnd.n6872 gnd.n128 585
R9324 gnd.n6871 gnd.n127 585
R9325 gnd.n7167 gnd.n127 585
R9326 gnd.n6870 gnd.n6869 585
R9327 gnd.n6869 gnd.n119 585
R9328 gnd.n6855 gnd.n118 585
R9329 gnd.n7173 gnd.n118 585
R9330 gnd.n6865 gnd.n6864 585
R9331 gnd.n6864 gnd.n109 585
R9332 gnd.n6863 gnd.n108 585
R9333 gnd.n7179 gnd.n108 585
R9334 gnd.n6862 gnd.n6861 585
R9335 gnd.n6861 gnd.n106 585
R9336 gnd.n6857 gnd.n97 585
R9337 gnd.n7185 gnd.n97 585
R9338 gnd.n84 gnd.n83 585
R9339 gnd.n86 gnd.n84 585
R9340 gnd.n7193 gnd.n7192 585
R9341 gnd.n7192 gnd.n7191 585
R9342 gnd.n7194 gnd.n82 585
R9343 gnd.n6821 gnd.n82 585
R9344 gnd.n321 gnd.n81 585
R9345 gnd.n321 gnd.n313 585
R9346 gnd.n6786 gnd.n322 585
R9347 gnd.n6813 gnd.n322 585
R9348 gnd.n6787 gnd.n6785 585
R9349 gnd.n6785 gnd.n319 585
R9350 gnd.n339 gnd.n330 585
R9351 gnd.n6802 gnd.n330 585
R9352 gnd.n6792 gnd.n6791 585
R9353 gnd.n6793 gnd.n6792 585
R9354 gnd.n338 gnd.n337 585
R9355 gnd.n337 gnd.n336 585
R9356 gnd.n6781 gnd.n6780 585
R9357 gnd.n6780 gnd.n6779 585
R9358 gnd.n342 gnd.n341 585
R9359 gnd.n354 gnd.n342 585
R9360 gnd.n366 gnd.n353 585
R9361 gnd.n6769 gnd.n353 585
R9362 gnd.n6753 gnd.n6752 585
R9363 gnd.n6754 gnd.n6753 585
R9364 gnd.n365 gnd.n364 585
R9365 gnd.n6728 gnd.n364 585
R9366 gnd.n6747 gnd.n6746 585
R9367 gnd.n6746 gnd.n6745 585
R9368 gnd.n369 gnd.n368 585
R9369 gnd.n6722 gnd.n369 585
R9370 gnd.n5419 gnd.n381 585
R9371 gnd.n6735 gnd.n381 585
R9372 gnd.n5420 gnd.n5418 585
R9373 gnd.n5418 gnd.n5417 585
R9374 gnd.n5345 gnd.n5336 585
R9375 gnd.n5443 gnd.n5336 585
R9376 gnd.n5425 gnd.n5424 585
R9377 gnd.n5426 gnd.n5425 585
R9378 gnd.n5344 gnd.n5329 585
R9379 gnd.n5449 gnd.n5329 585
R9380 gnd.n5407 gnd.n5406 585
R9381 gnd.n5408 gnd.n5407 585
R9382 gnd.n5350 gnd.n5318 585
R9383 gnd.n5455 gnd.n5318 585
R9384 gnd.n5402 gnd.n5401 585
R9385 gnd.n5401 gnd.n5400 585
R9386 gnd.n5352 gnd.n5307 585
R9387 gnd.n5461 gnd.n5307 585
R9388 gnd.n5379 gnd.n5378 585
R9389 gnd.n5380 gnd.n5379 585
R9390 gnd.n5367 gnd.n5288 585
R9391 gnd.n5467 gnd.n5288 585
R9392 gnd.n5374 gnd.n5373 585
R9393 gnd.n5373 gnd.n5286 585
R9394 gnd.n5372 gnd.n5371 585
R9395 gnd.n5372 gnd.n5274 585
R9396 gnd.n5370 gnd.n5273 585
R9397 gnd.n5475 gnd.n5273 585
R9398 gnd.n3620 gnd.n2270 585
R9399 gnd.n2322 gnd.n2270 585
R9400 gnd.n3621 gnd.n2332 585
R9401 gnd.n2332 gnd.n2321 585
R9402 gnd.n3623 gnd.n3622 585
R9403 gnd.n3624 gnd.n3623 585
R9404 gnd.n2333 gnd.n2331 585
R9405 gnd.n2340 gnd.n2331 585
R9406 gnd.n3614 gnd.n3613 585
R9407 gnd.n3613 gnd.n3612 585
R9408 gnd.n2336 gnd.n2335 585
R9409 gnd.n3339 gnd.n2336 585
R9410 gnd.n3325 gnd.n2359 585
R9411 gnd.n2359 gnd.n2349 585
R9412 gnd.n3327 gnd.n3326 585
R9413 gnd.n3328 gnd.n3327 585
R9414 gnd.n2360 gnd.n2358 585
R9415 gnd.n2358 gnd.n2356 585
R9416 gnd.n3320 gnd.n3319 585
R9417 gnd.n3319 gnd.n3318 585
R9418 gnd.n2363 gnd.n2362 585
R9419 gnd.n2372 gnd.n2363 585
R9420 gnd.n3276 gnd.n2386 585
R9421 gnd.n2386 gnd.n2371 585
R9422 gnd.n3278 gnd.n3277 585
R9423 gnd.n3279 gnd.n3278 585
R9424 gnd.n2387 gnd.n2385 585
R9425 gnd.n2394 gnd.n2385 585
R9426 gnd.n3271 gnd.n3270 585
R9427 gnd.n3270 gnd.n3269 585
R9428 gnd.n2390 gnd.n2389 585
R9429 gnd.n3250 gnd.n2390 585
R9430 gnd.n3236 gnd.n2414 585
R9431 gnd.n2414 gnd.n2403 585
R9432 gnd.n3238 gnd.n3237 585
R9433 gnd.n3239 gnd.n3238 585
R9434 gnd.n2415 gnd.n2413 585
R9435 gnd.n2413 gnd.n2410 585
R9436 gnd.n3231 gnd.n3230 585
R9437 gnd.n3230 gnd.n3229 585
R9438 gnd.n2418 gnd.n2417 585
R9439 gnd.n2428 gnd.n2418 585
R9440 gnd.n3191 gnd.n2441 585
R9441 gnd.n2441 gnd.n2427 585
R9442 gnd.n3193 gnd.n3192 585
R9443 gnd.n3194 gnd.n3193 585
R9444 gnd.n2442 gnd.n2440 585
R9445 gnd.n2449 gnd.n2440 585
R9446 gnd.n3186 gnd.n3185 585
R9447 gnd.n3185 gnd.n3184 585
R9448 gnd.n2445 gnd.n2444 585
R9449 gnd.n3165 gnd.n2445 585
R9450 gnd.n3151 gnd.n2468 585
R9451 gnd.n2468 gnd.n2458 585
R9452 gnd.n3153 gnd.n3152 585
R9453 gnd.n3154 gnd.n3153 585
R9454 gnd.n2469 gnd.n2467 585
R9455 gnd.n3142 gnd.n2467 585
R9456 gnd.n3146 gnd.n3145 585
R9457 gnd.n3145 gnd.n3144 585
R9458 gnd.n2472 gnd.n2471 585
R9459 gnd.n3097 gnd.n2472 585
R9460 gnd.n2590 gnd.n2589 585
R9461 gnd.n2591 gnd.n2590 585
R9462 gnd.n2570 gnd.n2569 585
R9463 gnd.n2573 gnd.n2570 585
R9464 gnd.n3107 gnd.n3106 585
R9465 gnd.n3106 gnd.n3105 585
R9466 gnd.n3108 gnd.n2564 585
R9467 gnd.n2600 gnd.n2564 585
R9468 gnd.n3110 gnd.n3109 585
R9469 gnd.n3111 gnd.n3110 585
R9470 gnd.n2565 gnd.n2563 585
R9471 gnd.n3075 gnd.n2563 585
R9472 gnd.n3059 gnd.n3058 585
R9473 gnd.n3058 gnd.n2551 585
R9474 gnd.n3060 gnd.n2615 585
R9475 gnd.n2615 gnd.n2550 585
R9476 gnd.n3062 gnd.n3061 585
R9477 gnd.n3063 gnd.n3062 585
R9478 gnd.n2616 gnd.n2614 585
R9479 gnd.n2614 gnd.n2611 585
R9480 gnd.n3051 gnd.n3050 585
R9481 gnd.n3050 gnd.n3049 585
R9482 gnd.n2619 gnd.n2618 585
R9483 gnd.n2626 gnd.n2619 585
R9484 gnd.n3025 gnd.n3024 585
R9485 gnd.n3026 gnd.n3025 585
R9486 gnd.n2638 gnd.n2637 585
R9487 gnd.n2645 gnd.n2637 585
R9488 gnd.n3020 gnd.n3019 585
R9489 gnd.n3019 gnd.n3018 585
R9490 gnd.n2641 gnd.n2640 585
R9491 gnd.n3008 gnd.n2641 585
R9492 gnd.n2995 gnd.n2665 585
R9493 gnd.n2665 gnd.n2664 585
R9494 gnd.n2997 gnd.n2996 585
R9495 gnd.n2998 gnd.n2997 585
R9496 gnd.n2666 gnd.n2663 585
R9497 gnd.n2673 gnd.n2663 585
R9498 gnd.n2990 gnd.n2989 585
R9499 gnd.n2989 gnd.n2988 585
R9500 gnd.n2669 gnd.n2668 585
R9501 gnd.n2977 gnd.n2669 585
R9502 gnd.n2964 gnd.n2690 585
R9503 gnd.n2690 gnd.n2689 585
R9504 gnd.n2966 gnd.n2965 585
R9505 gnd.n2967 gnd.n2966 585
R9506 gnd.n2960 gnd.n2688 585
R9507 gnd.n2959 gnd.n2958 585
R9508 gnd.n2693 gnd.n2692 585
R9509 gnd.n2956 gnd.n2693 585
R9510 gnd.n2715 gnd.n2714 585
R9511 gnd.n2718 gnd.n2717 585
R9512 gnd.n2716 gnd.n2711 585
R9513 gnd.n2723 gnd.n2722 585
R9514 gnd.n2725 gnd.n2724 585
R9515 gnd.n2728 gnd.n2727 585
R9516 gnd.n2726 gnd.n2709 585
R9517 gnd.n2733 gnd.n2732 585
R9518 gnd.n2735 gnd.n2734 585
R9519 gnd.n2738 gnd.n2737 585
R9520 gnd.n2736 gnd.n2707 585
R9521 gnd.n2743 gnd.n2742 585
R9522 gnd.n2747 gnd.n2744 585
R9523 gnd.n2748 gnd.n2685 585
R9524 gnd.n3626 gnd.n2285 585
R9525 gnd.n3693 gnd.n3692 585
R9526 gnd.n3695 gnd.n3694 585
R9527 gnd.n3697 gnd.n3696 585
R9528 gnd.n3699 gnd.n3698 585
R9529 gnd.n3701 gnd.n3700 585
R9530 gnd.n3703 gnd.n3702 585
R9531 gnd.n3705 gnd.n3704 585
R9532 gnd.n3707 gnd.n3706 585
R9533 gnd.n3709 gnd.n3708 585
R9534 gnd.n3711 gnd.n3710 585
R9535 gnd.n3713 gnd.n3712 585
R9536 gnd.n3715 gnd.n3714 585
R9537 gnd.n3718 gnd.n3717 585
R9538 gnd.n3716 gnd.n2273 585
R9539 gnd.n3722 gnd.n2271 585
R9540 gnd.n3724 gnd.n3723 585
R9541 gnd.n3725 gnd.n3724 585
R9542 gnd.n3627 gnd.n2327 585
R9543 gnd.n3627 gnd.n2322 585
R9544 gnd.n3629 gnd.n3628 585
R9545 gnd.n3628 gnd.n2321 585
R9546 gnd.n3625 gnd.n2326 585
R9547 gnd.n3625 gnd.n3624 585
R9548 gnd.n3604 gnd.n2328 585
R9549 gnd.n2340 gnd.n2328 585
R9550 gnd.n3603 gnd.n2338 585
R9551 gnd.n3612 gnd.n2338 585
R9552 gnd.n3338 gnd.n2345 585
R9553 gnd.n3339 gnd.n3338 585
R9554 gnd.n3337 gnd.n3336 585
R9555 gnd.n3337 gnd.n2349 585
R9556 gnd.n3335 gnd.n2351 585
R9557 gnd.n3328 gnd.n2351 585
R9558 gnd.n2364 gnd.n2352 585
R9559 gnd.n2364 gnd.n2356 585
R9560 gnd.n3284 gnd.n2365 585
R9561 gnd.n3318 gnd.n2365 585
R9562 gnd.n3283 gnd.n3282 585
R9563 gnd.n3282 gnd.n2372 585
R9564 gnd.n3281 gnd.n2380 585
R9565 gnd.n3281 gnd.n2371 585
R9566 gnd.n3280 gnd.n2382 585
R9567 gnd.n3280 gnd.n3279 585
R9568 gnd.n3259 gnd.n2381 585
R9569 gnd.n2394 gnd.n2381 585
R9570 gnd.n3258 gnd.n2392 585
R9571 gnd.n3269 gnd.n2392 585
R9572 gnd.n3249 gnd.n2399 585
R9573 gnd.n3250 gnd.n3249 585
R9574 gnd.n3248 gnd.n3247 585
R9575 gnd.n3248 gnd.n2403 585
R9576 gnd.n3246 gnd.n2405 585
R9577 gnd.n3239 gnd.n2405 585
R9578 gnd.n2420 gnd.n2406 585
R9579 gnd.n2420 gnd.n2410 585
R9580 gnd.n3199 gnd.n2421 585
R9581 gnd.n3229 gnd.n2421 585
R9582 gnd.n3198 gnd.n3197 585
R9583 gnd.n3197 gnd.n2428 585
R9584 gnd.n3196 gnd.n2435 585
R9585 gnd.n3196 gnd.n2427 585
R9586 gnd.n3195 gnd.n2437 585
R9587 gnd.n3195 gnd.n3194 585
R9588 gnd.n3174 gnd.n2436 585
R9589 gnd.n2449 gnd.n2436 585
R9590 gnd.n3173 gnd.n2447 585
R9591 gnd.n3184 gnd.n2447 585
R9592 gnd.n3164 gnd.n2454 585
R9593 gnd.n3165 gnd.n3164 585
R9594 gnd.n3163 gnd.n3162 585
R9595 gnd.n3163 gnd.n2458 585
R9596 gnd.n3161 gnd.n2460 585
R9597 gnd.n3154 gnd.n2460 585
R9598 gnd.n3141 gnd.n2461 585
R9599 gnd.n3142 gnd.n3141 585
R9600 gnd.n3094 gnd.n2474 585
R9601 gnd.n3144 gnd.n2474 585
R9602 gnd.n3096 gnd.n3095 585
R9603 gnd.n3097 gnd.n3096 585
R9604 gnd.n3089 gnd.n2592 585
R9605 gnd.n2592 gnd.n2591 585
R9606 gnd.n3087 gnd.n3086 585
R9607 gnd.n3086 gnd.n2573 585
R9608 gnd.n3084 gnd.n2571 585
R9609 gnd.n3105 gnd.n2571 585
R9610 gnd.n2602 gnd.n2601 585
R9611 gnd.n2601 gnd.n2600 585
R9612 gnd.n3078 gnd.n2561 585
R9613 gnd.n3111 gnd.n2561 585
R9614 gnd.n3077 gnd.n3076 585
R9615 gnd.n3076 gnd.n3075 585
R9616 gnd.n3073 gnd.n2604 585
R9617 gnd.n3073 gnd.n2551 585
R9618 gnd.n3072 gnd.n3071 585
R9619 gnd.n3072 gnd.n2550 585
R9620 gnd.n2607 gnd.n2606 585
R9621 gnd.n3063 gnd.n2606 585
R9622 gnd.n3031 gnd.n3030 585
R9623 gnd.n3030 gnd.n2611 585
R9624 gnd.n3032 gnd.n2620 585
R9625 gnd.n3049 gnd.n2620 585
R9626 gnd.n3029 gnd.n3028 585
R9627 gnd.n3028 gnd.n2626 585
R9628 gnd.n3027 gnd.n2634 585
R9629 gnd.n3027 gnd.n3026 585
R9630 gnd.n3012 gnd.n2635 585
R9631 gnd.n2645 gnd.n2635 585
R9632 gnd.n3011 gnd.n2643 585
R9633 gnd.n3018 gnd.n2643 585
R9634 gnd.n3010 gnd.n3009 585
R9635 gnd.n3009 gnd.n3008 585
R9636 gnd.n2654 gnd.n2651 585
R9637 gnd.n2664 gnd.n2654 585
R9638 gnd.n3000 gnd.n2999 585
R9639 gnd.n2999 gnd.n2998 585
R9640 gnd.n2660 gnd.n2659 585
R9641 gnd.n2673 gnd.n2660 585
R9642 gnd.n2980 gnd.n2671 585
R9643 gnd.n2988 gnd.n2671 585
R9644 gnd.n2979 gnd.n2978 585
R9645 gnd.n2978 gnd.n2977 585
R9646 gnd.n2680 gnd.n2678 585
R9647 gnd.n2689 gnd.n2680 585
R9648 gnd.n2969 gnd.n2968 585
R9649 gnd.n2968 gnd.n2967 585
R9650 gnd.n5182 gnd.n5181 585
R9651 gnd.n5183 gnd.n5182 585
R9652 gnd.n1408 gnd.n1406 585
R9653 gnd.n1406 gnd.n1402 585
R9654 gnd.n5055 gnd.n5054 585
R9655 gnd.n5056 gnd.n5055 585
R9656 gnd.n5053 gnd.n1481 585
R9657 gnd.n1486 gnd.n1481 585
R9658 gnd.n5052 gnd.n5051 585
R9659 gnd.n5051 gnd.n5050 585
R9660 gnd.n1483 gnd.n1482 585
R9661 gnd.n5027 gnd.n1483 585
R9662 gnd.n5039 gnd.n5038 585
R9663 gnd.n5040 gnd.n5039 585
R9664 gnd.n5037 gnd.n1497 585
R9665 gnd.n1497 gnd.n1493 585
R9666 gnd.n5036 gnd.n5035 585
R9667 gnd.n5035 gnd.n5034 585
R9668 gnd.n1499 gnd.n1498 585
R9669 gnd.n4967 gnd.n1499 585
R9670 gnd.n5020 gnd.n5019 585
R9671 gnd.n5021 gnd.n5020 585
R9672 gnd.n5018 gnd.n1506 585
R9673 gnd.n1506 gnd.n1505 585
R9674 gnd.n5017 gnd.n5016 585
R9675 gnd.n5016 gnd.n5015 585
R9676 gnd.n1508 gnd.n1507 585
R9677 gnd.n1521 gnd.n1508 585
R9678 gnd.n5002 gnd.n5001 585
R9679 gnd.n5003 gnd.n5002 585
R9680 gnd.n5000 gnd.n1522 585
R9681 gnd.n1522 gnd.n1518 585
R9682 gnd.n4999 gnd.n4998 585
R9683 gnd.n4998 gnd.n4997 585
R9684 gnd.n1524 gnd.n1523 585
R9685 gnd.n4875 gnd.n1524 585
R9686 gnd.n4942 gnd.n4941 585
R9687 gnd.n4942 gnd.n1532 585
R9688 gnd.n4944 gnd.n4943 585
R9689 gnd.n4943 gnd.t8 585
R9690 gnd.n4945 gnd.n1545 585
R9691 gnd.n1545 gnd.n1543 585
R9692 gnd.n4947 gnd.n4946 585
R9693 gnd.n4948 gnd.n4947 585
R9694 gnd.n4940 gnd.n1544 585
R9695 gnd.n1544 gnd.n1539 585
R9696 gnd.n4939 gnd.n4938 585
R9697 gnd.n4938 gnd.n4937 585
R9698 gnd.n1547 gnd.n1546 585
R9699 gnd.n4871 gnd.n1547 585
R9700 gnd.n4910 gnd.n4909 585
R9701 gnd.n4910 gnd.n1556 585
R9702 gnd.n4912 gnd.n4911 585
R9703 gnd.n4911 gnd.n1555 585
R9704 gnd.n4913 gnd.n1569 585
R9705 gnd.n4898 gnd.n1569 585
R9706 gnd.n4915 gnd.n4914 585
R9707 gnd.n4916 gnd.n4915 585
R9708 gnd.n4908 gnd.n1568 585
R9709 gnd.n1568 gnd.n1563 585
R9710 gnd.n4907 gnd.n4906 585
R9711 gnd.n4906 gnd.n4905 585
R9712 gnd.n1571 gnd.n1570 585
R9713 gnd.n1578 gnd.n1571 585
R9714 gnd.n4864 gnd.n4863 585
R9715 gnd.n4865 gnd.n4864 585
R9716 gnd.n4862 gnd.n1580 585
R9717 gnd.n1580 gnd.n1577 585
R9718 gnd.n4861 gnd.n4860 585
R9719 gnd.n4860 gnd.n4859 585
R9720 gnd.n1582 gnd.n1581 585
R9721 gnd.n1596 gnd.n1582 585
R9722 gnd.n4846 gnd.n4845 585
R9723 gnd.n4847 gnd.n4846 585
R9724 gnd.n4844 gnd.n1597 585
R9725 gnd.n1597 gnd.n1593 585
R9726 gnd.n4843 gnd.n4842 585
R9727 gnd.n4842 gnd.n4841 585
R9728 gnd.n1599 gnd.n1598 585
R9729 gnd.n1600 gnd.n1599 585
R9730 gnd.n4801 gnd.n4800 585
R9731 gnd.n4801 gnd.n1609 585
R9732 gnd.n4803 gnd.n4802 585
R9733 gnd.n4802 gnd.n1608 585
R9734 gnd.n4804 gnd.n1623 585
R9735 gnd.n1623 gnd.n1621 585
R9736 gnd.n4806 gnd.n4805 585
R9737 gnd.n4807 gnd.n4806 585
R9738 gnd.n4799 gnd.n1622 585
R9739 gnd.n4793 gnd.n1622 585
R9740 gnd.n4798 gnd.n4797 585
R9741 gnd.n4797 gnd.n4796 585
R9742 gnd.n1625 gnd.n1624 585
R9743 gnd.n1626 gnd.n1625 585
R9744 gnd.n4769 gnd.n4768 585
R9745 gnd.n4770 gnd.n4769 585
R9746 gnd.n4767 gnd.n1632 585
R9747 gnd.n4763 gnd.n1632 585
R9748 gnd.n4766 gnd.n4765 585
R9749 gnd.n4765 gnd.n4764 585
R9750 gnd.n1634 gnd.n1633 585
R9751 gnd.n4750 gnd.n1634 585
R9752 gnd.n4739 gnd.n1651 585
R9753 gnd.n1651 gnd.n1644 585
R9754 gnd.n4741 gnd.n4740 585
R9755 gnd.n4742 gnd.n4741 585
R9756 gnd.n4738 gnd.n1650 585
R9757 gnd.n1656 gnd.n1650 585
R9758 gnd.n4737 gnd.n4736 585
R9759 gnd.n4736 gnd.n4735 585
R9760 gnd.n1653 gnd.n1652 585
R9761 gnd.n4711 gnd.n1653 585
R9762 gnd.n4723 gnd.n4722 585
R9763 gnd.n4724 gnd.n4723 585
R9764 gnd.n4721 gnd.n1666 585
R9765 gnd.n1666 gnd.n1662 585
R9766 gnd.n4720 gnd.n4719 585
R9767 gnd.n4719 gnd.n4718 585
R9768 gnd.n1668 gnd.n1667 585
R9769 gnd.n1675 gnd.n1668 585
R9770 gnd.n4705 gnd.n4704 585
R9771 gnd.n4706 gnd.n4705 585
R9772 gnd.n4703 gnd.n1677 585
R9773 gnd.n1677 gnd.n1674 585
R9774 gnd.n4702 gnd.n4701 585
R9775 gnd.n4701 gnd.t327 585
R9776 gnd.n1679 gnd.n1678 585
R9777 gnd.n1692 gnd.n1679 585
R9778 gnd.n4688 gnd.n4687 585
R9779 gnd.n4689 gnd.n4688 585
R9780 gnd.n4686 gnd.n1693 585
R9781 gnd.n4681 gnd.n1693 585
R9782 gnd.n4685 gnd.n4684 585
R9783 gnd.n4684 gnd.n4683 585
R9784 gnd.n1695 gnd.n1694 585
R9785 gnd.n4671 gnd.n1695 585
R9786 gnd.n4669 gnd.n4668 585
R9787 gnd.n4670 gnd.n4669 585
R9788 gnd.n4667 gnd.n1703 585
R9789 gnd.n4633 gnd.n1703 585
R9790 gnd.n4666 gnd.n4665 585
R9791 gnd.n4665 gnd.n4664 585
R9792 gnd.n1705 gnd.n1704 585
R9793 gnd.n1706 gnd.n1705 585
R9794 gnd.n4648 gnd.n4647 585
R9795 gnd.n4649 gnd.n4648 585
R9796 gnd.n4646 gnd.n1716 585
R9797 gnd.n1716 gnd.n1713 585
R9798 gnd.n4645 gnd.n4644 585
R9799 gnd.n4644 gnd.n4643 585
R9800 gnd.n1718 gnd.n1717 585
R9801 gnd.n1718 gnd.n1126 585
R9802 gnd.n4625 gnd.n4623 585
R9803 gnd.n4623 gnd.n1124 585
R9804 gnd.n4627 gnd.n4626 585
R9805 gnd.n4628 gnd.n4627 585
R9806 gnd.n4624 gnd.n4622 585
R9807 gnd.n4622 gnd.n1114 585
R9808 gnd.n1109 gnd.n1108 585
R9809 gnd.n5826 gnd.n1109 585
R9810 gnd.n5829 gnd.n5828 585
R9811 gnd.n5828 gnd.n5827 585
R9812 gnd.n5830 gnd.n1087 585
R9813 gnd.n1787 gnd.n1087 585
R9814 gnd.n5895 gnd.n5894 585
R9815 gnd.n5893 gnd.n1086 585
R9816 gnd.n5892 gnd.n1085 585
R9817 gnd.n5897 gnd.n1085 585
R9818 gnd.n5891 gnd.n5890 585
R9819 gnd.n5889 gnd.n5888 585
R9820 gnd.n5887 gnd.n5886 585
R9821 gnd.n5885 gnd.n5884 585
R9822 gnd.n5883 gnd.n5882 585
R9823 gnd.n5881 gnd.n5880 585
R9824 gnd.n5879 gnd.n5878 585
R9825 gnd.n5877 gnd.n5876 585
R9826 gnd.n5875 gnd.n5874 585
R9827 gnd.n5873 gnd.n5872 585
R9828 gnd.n5871 gnd.n5870 585
R9829 gnd.n5869 gnd.n5868 585
R9830 gnd.n5867 gnd.n5866 585
R9831 gnd.n5865 gnd.n5864 585
R9832 gnd.n5863 gnd.n5862 585
R9833 gnd.n5861 gnd.n5860 585
R9834 gnd.n5859 gnd.n5858 585
R9835 gnd.n5857 gnd.n5856 585
R9836 gnd.n5855 gnd.n5854 585
R9837 gnd.n5853 gnd.n5852 585
R9838 gnd.n5851 gnd.n5850 585
R9839 gnd.n5849 gnd.n5848 585
R9840 gnd.n5847 gnd.n5846 585
R9841 gnd.n5845 gnd.n5844 585
R9842 gnd.n5843 gnd.n5842 585
R9843 gnd.n5841 gnd.n5840 585
R9844 gnd.n5839 gnd.n5838 585
R9845 gnd.n5837 gnd.n5836 585
R9846 gnd.n5835 gnd.n1049 585
R9847 gnd.n5900 gnd.n5899 585
R9848 gnd.n1051 gnd.n1048 585
R9849 gnd.n1725 gnd.n1724 585
R9850 gnd.n1727 gnd.n1726 585
R9851 gnd.n1730 gnd.n1729 585
R9852 gnd.n1732 gnd.n1731 585
R9853 gnd.n1734 gnd.n1733 585
R9854 gnd.n1736 gnd.n1735 585
R9855 gnd.n1738 gnd.n1737 585
R9856 gnd.n1740 gnd.n1739 585
R9857 gnd.n1742 gnd.n1741 585
R9858 gnd.n1744 gnd.n1743 585
R9859 gnd.n1746 gnd.n1745 585
R9860 gnd.n1748 gnd.n1747 585
R9861 gnd.n1750 gnd.n1749 585
R9862 gnd.n1752 gnd.n1751 585
R9863 gnd.n1754 gnd.n1753 585
R9864 gnd.n1756 gnd.n1755 585
R9865 gnd.n1758 gnd.n1757 585
R9866 gnd.n1760 gnd.n1759 585
R9867 gnd.n1762 gnd.n1761 585
R9868 gnd.n1764 gnd.n1763 585
R9869 gnd.n1766 gnd.n1765 585
R9870 gnd.n1768 gnd.n1767 585
R9871 gnd.n1770 gnd.n1769 585
R9872 gnd.n1772 gnd.n1771 585
R9873 gnd.n1774 gnd.n1773 585
R9874 gnd.n1776 gnd.n1775 585
R9875 gnd.n1778 gnd.n1777 585
R9876 gnd.n1780 gnd.n1779 585
R9877 gnd.n1782 gnd.n1781 585
R9878 gnd.n1784 gnd.n1783 585
R9879 gnd.n1786 gnd.n1785 585
R9880 gnd.n5063 gnd.n5062 585
R9881 gnd.n5064 gnd.n1477 585
R9882 gnd.n5066 gnd.n5065 585
R9883 gnd.n5068 gnd.n1475 585
R9884 gnd.n5070 gnd.n5069 585
R9885 gnd.n5071 gnd.n1474 585
R9886 gnd.n5073 gnd.n5072 585
R9887 gnd.n5075 gnd.n1472 585
R9888 gnd.n5077 gnd.n5076 585
R9889 gnd.n5078 gnd.n1471 585
R9890 gnd.n5080 gnd.n5079 585
R9891 gnd.n5082 gnd.n1469 585
R9892 gnd.n5084 gnd.n5083 585
R9893 gnd.n5085 gnd.n1468 585
R9894 gnd.n5087 gnd.n5086 585
R9895 gnd.n5089 gnd.n1466 585
R9896 gnd.n5091 gnd.n5090 585
R9897 gnd.n5092 gnd.n1465 585
R9898 gnd.n5094 gnd.n5093 585
R9899 gnd.n5096 gnd.n1463 585
R9900 gnd.n5098 gnd.n5097 585
R9901 gnd.n5099 gnd.n1462 585
R9902 gnd.n5101 gnd.n5100 585
R9903 gnd.n5103 gnd.n1460 585
R9904 gnd.n5105 gnd.n5104 585
R9905 gnd.n5106 gnd.n1459 585
R9906 gnd.n5108 gnd.n5107 585
R9907 gnd.n5110 gnd.n1457 585
R9908 gnd.n5112 gnd.n5111 585
R9909 gnd.n5114 gnd.n1454 585
R9910 gnd.n5116 gnd.n5115 585
R9911 gnd.n5118 gnd.n1453 585
R9912 gnd.n5119 gnd.n1394 585
R9913 gnd.n5122 gnd.n1310 585
R9914 gnd.n5124 gnd.n5123 585
R9915 gnd.n5126 gnd.n1451 585
R9916 gnd.n5128 gnd.n5127 585
R9917 gnd.n5130 gnd.n1448 585
R9918 gnd.n5132 gnd.n5131 585
R9919 gnd.n5134 gnd.n1446 585
R9920 gnd.n5136 gnd.n5135 585
R9921 gnd.n5137 gnd.n1445 585
R9922 gnd.n5139 gnd.n5138 585
R9923 gnd.n5141 gnd.n1443 585
R9924 gnd.n5143 gnd.n5142 585
R9925 gnd.n5144 gnd.n1442 585
R9926 gnd.n5146 gnd.n5145 585
R9927 gnd.n5148 gnd.n1440 585
R9928 gnd.n5150 gnd.n5149 585
R9929 gnd.n5151 gnd.n1439 585
R9930 gnd.n5153 gnd.n5152 585
R9931 gnd.n5155 gnd.n1437 585
R9932 gnd.n5157 gnd.n5156 585
R9933 gnd.n5158 gnd.n1436 585
R9934 gnd.n5160 gnd.n5159 585
R9935 gnd.n5162 gnd.n1434 585
R9936 gnd.n5164 gnd.n5163 585
R9937 gnd.n5165 gnd.n1433 585
R9938 gnd.n5167 gnd.n5166 585
R9939 gnd.n5169 gnd.n1431 585
R9940 gnd.n5171 gnd.n5170 585
R9941 gnd.n5172 gnd.n1430 585
R9942 gnd.n5174 gnd.n5173 585
R9943 gnd.n5176 gnd.n1428 585
R9944 gnd.n5178 gnd.n5177 585
R9945 gnd.n5179 gnd.n1407 585
R9946 gnd.n5060 gnd.n1404 585
R9947 gnd.n5183 gnd.n1404 585
R9948 gnd.n5059 gnd.n5058 585
R9949 gnd.n5058 gnd.n1402 585
R9950 gnd.n5057 gnd.n1478 585
R9951 gnd.n5057 gnd.n5056 585
R9952 gnd.n5025 gnd.n1479 585
R9953 gnd.n1486 gnd.n1479 585
R9954 gnd.n5026 gnd.n1484 585
R9955 gnd.n5050 gnd.n1484 585
R9956 gnd.n5029 gnd.n5028 585
R9957 gnd.n5028 gnd.n5027 585
R9958 gnd.n5030 gnd.n1495 585
R9959 gnd.n5040 gnd.n1495 585
R9960 gnd.n5031 gnd.n1502 585
R9961 gnd.n1502 gnd.n1493 585
R9962 gnd.n5033 gnd.n5032 585
R9963 gnd.n5034 gnd.n5033 585
R9964 gnd.n5024 gnd.n1501 585
R9965 gnd.n4967 gnd.n1501 585
R9966 gnd.n5023 gnd.n5022 585
R9967 gnd.n5022 gnd.n5021 585
R9968 gnd.n1504 gnd.n1503 585
R9969 gnd.n1505 gnd.n1504 585
R9970 gnd.n4877 gnd.n1510 585
R9971 gnd.n5015 gnd.n1510 585
R9972 gnd.n4879 gnd.n4878 585
R9973 gnd.n4878 gnd.n1521 585
R9974 gnd.n4880 gnd.n1520 585
R9975 gnd.n5003 gnd.n1520 585
R9976 gnd.n4882 gnd.n4881 585
R9977 gnd.n4881 gnd.n1518 585
R9978 gnd.n4883 gnd.n1525 585
R9979 gnd.n4997 gnd.n1525 585
R9980 gnd.n4884 gnd.n4876 585
R9981 gnd.n4876 gnd.n4875 585
R9982 gnd.n4886 gnd.n4885 585
R9983 gnd.n4886 gnd.n1532 585
R9984 gnd.n4887 gnd.n4873 585
R9985 gnd.n4887 gnd.t8 585
R9986 gnd.n4889 gnd.n4888 585
R9987 gnd.n4888 gnd.n1543 585
R9988 gnd.n4890 gnd.n1541 585
R9989 gnd.n4948 gnd.n1541 585
R9990 gnd.n4892 gnd.n4891 585
R9991 gnd.n4891 gnd.n1539 585
R9992 gnd.n4893 gnd.n1548 585
R9993 gnd.n4937 gnd.n1548 585
R9994 gnd.n4894 gnd.n4872 585
R9995 gnd.n4872 gnd.n4871 585
R9996 gnd.n4896 gnd.n4895 585
R9997 gnd.n4896 gnd.n1556 585
R9998 gnd.n4897 gnd.n4869 585
R9999 gnd.n4897 gnd.n1555 585
R10000 gnd.n4900 gnd.n4899 585
R10001 gnd.n4899 gnd.n4898 585
R10002 gnd.n4901 gnd.n1565 585
R10003 gnd.n4916 gnd.n1565 585
R10004 gnd.n4902 gnd.n1574 585
R10005 gnd.n1574 gnd.n1563 585
R10006 gnd.n4904 gnd.n4903 585
R10007 gnd.n4905 gnd.n4904 585
R10008 gnd.n4868 gnd.n1573 585
R10009 gnd.n1578 gnd.n1573 585
R10010 gnd.n4867 gnd.n4866 585
R10011 gnd.n4866 gnd.n4865 585
R10012 gnd.n1576 gnd.n1575 585
R10013 gnd.n1577 gnd.n1576 585
R10014 gnd.n4777 gnd.n1584 585
R10015 gnd.n4859 gnd.n1584 585
R10016 gnd.n4779 gnd.n4778 585
R10017 gnd.n4778 gnd.n1596 585
R10018 gnd.n4780 gnd.n1595 585
R10019 gnd.n4847 gnd.n1595 585
R10020 gnd.n4782 gnd.n4781 585
R10021 gnd.n4781 gnd.n1593 585
R10022 gnd.n4783 gnd.n1601 585
R10023 gnd.n4841 gnd.n1601 585
R10024 gnd.n4784 gnd.n4776 585
R10025 gnd.n4776 gnd.n1600 585
R10026 gnd.n4786 gnd.n4785 585
R10027 gnd.n4786 gnd.n1609 585
R10028 gnd.n4787 gnd.n4775 585
R10029 gnd.n4787 gnd.n1608 585
R10030 gnd.n4789 gnd.n4788 585
R10031 gnd.n4788 gnd.n1621 585
R10032 gnd.n4790 gnd.n1619 585
R10033 gnd.n4807 gnd.n1619 585
R10034 gnd.n4792 gnd.n4791 585
R10035 gnd.n4793 gnd.n4792 585
R10036 gnd.n4774 gnd.n1627 585
R10037 gnd.n4796 gnd.n1627 585
R10038 gnd.n4773 gnd.n4772 585
R10039 gnd.n4772 gnd.n1626 585
R10040 gnd.n4771 gnd.n1629 585
R10041 gnd.n4771 gnd.n4770 585
R10042 gnd.n4746 gnd.n1630 585
R10043 gnd.n4763 gnd.n1630 585
R10044 gnd.n4747 gnd.n1636 585
R10045 gnd.n4764 gnd.n1636 585
R10046 gnd.n4749 gnd.n4748 585
R10047 gnd.n4750 gnd.n4749 585
R10048 gnd.n4745 gnd.n1646 585
R10049 gnd.n1646 gnd.n1644 585
R10050 gnd.n4744 gnd.n4743 585
R10051 gnd.n4743 gnd.n4742 585
R10052 gnd.n1648 gnd.n1647 585
R10053 gnd.n1656 gnd.n1648 585
R10054 gnd.n4710 gnd.n1654 585
R10055 gnd.n4735 gnd.n1654 585
R10056 gnd.n4713 gnd.n4712 585
R10057 gnd.n4712 gnd.n4711 585
R10058 gnd.n4714 gnd.n1664 585
R10059 gnd.n4724 gnd.n1664 585
R10060 gnd.n4715 gnd.n1671 585
R10061 gnd.n1671 gnd.n1662 585
R10062 gnd.n4717 gnd.n4716 585
R10063 gnd.n4718 gnd.n4717 585
R10064 gnd.n4709 gnd.n1670 585
R10065 gnd.n1675 gnd.n1670 585
R10066 gnd.n4708 gnd.n4707 585
R10067 gnd.n4707 gnd.n4706 585
R10068 gnd.n1673 gnd.n1672 585
R10069 gnd.n1674 gnd.n1673 585
R10070 gnd.n4675 gnd.n1682 585
R10071 gnd.t327 gnd.n1682 585
R10072 gnd.n4677 gnd.n4676 585
R10073 gnd.n4676 gnd.n1692 585
R10074 gnd.n4678 gnd.n1691 585
R10075 gnd.n4689 gnd.n1691 585
R10076 gnd.n4680 gnd.n4679 585
R10077 gnd.n4681 gnd.n4680 585
R10078 gnd.n4674 gnd.n1697 585
R10079 gnd.n4683 gnd.n1697 585
R10080 gnd.n4673 gnd.n4672 585
R10081 gnd.n4672 gnd.n4671 585
R10082 gnd.n1700 gnd.n1699 585
R10083 gnd.n4670 gnd.n1700 585
R10084 gnd.n4635 gnd.n4634 585
R10085 gnd.n4634 gnd.n4633 585
R10086 gnd.n4636 gnd.n1707 585
R10087 gnd.n4664 gnd.n1707 585
R10088 gnd.n4638 gnd.n4637 585
R10089 gnd.n4637 gnd.n1706 585
R10090 gnd.n4639 gnd.n1715 585
R10091 gnd.n4649 gnd.n1715 585
R10092 gnd.n4640 gnd.n1720 585
R10093 gnd.n1720 gnd.n1713 585
R10094 gnd.n4642 gnd.n4641 585
R10095 gnd.n4643 gnd.n4642 585
R10096 gnd.n4632 gnd.n1719 585
R10097 gnd.n1719 gnd.n1126 585
R10098 gnd.n4631 gnd.n4630 585
R10099 gnd.n4630 gnd.n1124 585
R10100 gnd.n4629 gnd.n1721 585
R10101 gnd.n4629 gnd.n4628 585
R10102 gnd.n1793 gnd.n1792 585
R10103 gnd.n1793 gnd.n1114 585
R10104 gnd.n1791 gnd.n1112 585
R10105 gnd.n5826 gnd.n1112 585
R10106 gnd.n1790 gnd.n1111 585
R10107 gnd.n5827 gnd.n1111 585
R10108 gnd.n1789 gnd.n1788 585
R10109 gnd.n1788 gnd.n1787 585
R10110 gnd.n5956 gnd.n972 585
R10111 gnd.n4468 gnd.n972 585
R10112 gnd.n5958 gnd.n5957 585
R10113 gnd.n5959 gnd.n5958 585
R10114 gnd.n957 gnd.n956 585
R10115 gnd.n4372 gnd.n957 585
R10116 gnd.n5967 gnd.n5966 585
R10117 gnd.n5966 gnd.n5965 585
R10118 gnd.n5968 gnd.n951 585
R10119 gnd.n4362 gnd.n951 585
R10120 gnd.n5970 gnd.n5969 585
R10121 gnd.n5971 gnd.n5970 585
R10122 gnd.n937 gnd.n936 585
R10123 gnd.n4355 gnd.n937 585
R10124 gnd.n5979 gnd.n5978 585
R10125 gnd.n5978 gnd.n5977 585
R10126 gnd.n5980 gnd.n931 585
R10127 gnd.n4347 gnd.n931 585
R10128 gnd.n5982 gnd.n5981 585
R10129 gnd.n5983 gnd.n5982 585
R10130 gnd.n917 gnd.n916 585
R10131 gnd.n4340 gnd.n917 585
R10132 gnd.n5991 gnd.n5990 585
R10133 gnd.n5990 gnd.n5989 585
R10134 gnd.n5992 gnd.n911 585
R10135 gnd.n4283 gnd.n911 585
R10136 gnd.n5994 gnd.n5993 585
R10137 gnd.n5995 gnd.n5994 585
R10138 gnd.n895 gnd.n894 585
R10139 gnd.n4294 gnd.n895 585
R10140 gnd.n6003 gnd.n6002 585
R10141 gnd.n6002 gnd.n6001 585
R10142 gnd.n6004 gnd.n889 585
R10143 gnd.n4274 gnd.n889 585
R10144 gnd.n6006 gnd.n6005 585
R10145 gnd.n6007 gnd.n6006 585
R10146 gnd.n890 gnd.n888 585
R10147 gnd.n888 gnd.n883 585
R10148 gnd.n4264 gnd.n4263 585
R10149 gnd.n4265 gnd.n4264 585
R10150 gnd.n2082 gnd.n2081 585
R10151 gnd.n2089 gnd.n2081 585
R10152 gnd.n4258 gnd.n4257 585
R10153 gnd.n4257 gnd.n4256 585
R10154 gnd.n2085 gnd.n2084 585
R10155 gnd.n2086 gnd.n2085 585
R10156 gnd.n4236 gnd.n4235 585
R10157 gnd.n4237 gnd.n4236 585
R10158 gnd.n2103 gnd.n2102 585
R10159 gnd.n2102 gnd.n2099 585
R10160 gnd.n4231 gnd.n4230 585
R10161 gnd.n4230 gnd.n4229 585
R10162 gnd.n2106 gnd.n2105 585
R10163 gnd.n4218 gnd.n2106 585
R10164 gnd.n4193 gnd.n2127 585
R10165 gnd.n2127 gnd.n2116 585
R10166 gnd.n4195 gnd.n4194 585
R10167 gnd.n4196 gnd.n4195 585
R10168 gnd.n2128 gnd.n2126 585
R10169 gnd.n2126 gnd.n2123 585
R10170 gnd.n4188 gnd.n4187 585
R10171 gnd.n4187 gnd.n4186 585
R10172 gnd.n2131 gnd.n2130 585
R10173 gnd.n4171 gnd.n2131 585
R10174 gnd.n4158 gnd.n2151 585
R10175 gnd.n2151 gnd.n2142 585
R10176 gnd.n4160 gnd.n4159 585
R10177 gnd.n4161 gnd.n4160 585
R10178 gnd.n2152 gnd.n2150 585
R10179 gnd.n2158 gnd.n2150 585
R10180 gnd.n4153 gnd.n4152 585
R10181 gnd.n4152 gnd.n4151 585
R10182 gnd.n2155 gnd.n2154 585
R10183 gnd.n4136 gnd.n2155 585
R10184 gnd.n4123 gnd.n2176 585
R10185 gnd.n2176 gnd.n2167 585
R10186 gnd.n4125 gnd.n4124 585
R10187 gnd.n4126 gnd.n4125 585
R10188 gnd.n2177 gnd.n2175 585
R10189 gnd.n2184 gnd.n2175 585
R10190 gnd.n4118 gnd.n4117 585
R10191 gnd.n4117 gnd.n4116 585
R10192 gnd.n2180 gnd.n2179 585
R10193 gnd.n2181 gnd.n2180 585
R10194 gnd.n4099 gnd.n4098 585
R10195 gnd.n4100 gnd.n4099 585
R10196 gnd.n2197 gnd.n2196 585
R10197 gnd.n2196 gnd.n2193 585
R10198 gnd.n4094 gnd.n4093 585
R10199 gnd.n4093 gnd.n4092 585
R10200 gnd.n2200 gnd.n2199 585
R10201 gnd.n2201 gnd.n2200 585
R10202 gnd.n4079 gnd.n4078 585
R10203 gnd.n4080 gnd.n4079 585
R10204 gnd.n2214 gnd.n2213 585
R10205 gnd.n2221 gnd.n2213 585
R10206 gnd.n4074 gnd.n4073 585
R10207 gnd.n4073 gnd.n4072 585
R10208 gnd.n2217 gnd.n2216 585
R10209 gnd.n2218 gnd.n2217 585
R10210 gnd.n4059 gnd.n4058 585
R10211 gnd.n4060 gnd.n4059 585
R10212 gnd.n2233 gnd.n2232 585
R10213 gnd.n2232 gnd.n2229 585
R10214 gnd.n4054 gnd.n4053 585
R10215 gnd.n4053 gnd.n4052 585
R10216 gnd.n2236 gnd.n2235 585
R10217 gnd.n2237 gnd.n2236 585
R10218 gnd.n4037 gnd.n4036 585
R10219 gnd.n4035 gnd.n3764 585
R10220 gnd.n4034 gnd.n3763 585
R10221 gnd.n4039 gnd.n3763 585
R10222 gnd.n4033 gnd.n4032 585
R10223 gnd.n4031 gnd.n4030 585
R10224 gnd.n4029 gnd.n4028 585
R10225 gnd.n4027 gnd.n4026 585
R10226 gnd.n4025 gnd.n4024 585
R10227 gnd.n4023 gnd.n4022 585
R10228 gnd.n4021 gnd.n4020 585
R10229 gnd.n4019 gnd.n4018 585
R10230 gnd.n4017 gnd.n4016 585
R10231 gnd.n4015 gnd.n4014 585
R10232 gnd.n4013 gnd.n4012 585
R10233 gnd.n4011 gnd.n4010 585
R10234 gnd.n4009 gnd.n4008 585
R10235 gnd.n4007 gnd.n4006 585
R10236 gnd.n4005 gnd.n4004 585
R10237 gnd.n4002 gnd.n4001 585
R10238 gnd.n4000 gnd.n3999 585
R10239 gnd.n3998 gnd.n3997 585
R10240 gnd.n3996 gnd.n3995 585
R10241 gnd.n3994 gnd.n3993 585
R10242 gnd.n3992 gnd.n3991 585
R10243 gnd.n3990 gnd.n3989 585
R10244 gnd.n3988 gnd.n3987 585
R10245 gnd.n3986 gnd.n3985 585
R10246 gnd.n3984 gnd.n3983 585
R10247 gnd.n3982 gnd.n3981 585
R10248 gnd.n3980 gnd.n3979 585
R10249 gnd.n3978 gnd.n3977 585
R10250 gnd.n3976 gnd.n3975 585
R10251 gnd.n3974 gnd.n3973 585
R10252 gnd.n3972 gnd.n3971 585
R10253 gnd.n3970 gnd.n3969 585
R10254 gnd.n3968 gnd.n3967 585
R10255 gnd.n3966 gnd.n3965 585
R10256 gnd.n3964 gnd.n3963 585
R10257 gnd.n3962 gnd.n3961 585
R10258 gnd.n3960 gnd.n3959 585
R10259 gnd.n3958 gnd.n3957 585
R10260 gnd.n3956 gnd.n3955 585
R10261 gnd.n3954 gnd.n3953 585
R10262 gnd.n3952 gnd.n3951 585
R10263 gnd.n3950 gnd.n3949 585
R10264 gnd.n3948 gnd.n3947 585
R10265 gnd.n3946 gnd.n3945 585
R10266 gnd.n3944 gnd.n3943 585
R10267 gnd.n3942 gnd.n3941 585
R10268 gnd.n3940 gnd.n3939 585
R10269 gnd.n3938 gnd.n3937 585
R10270 gnd.n3936 gnd.n3935 585
R10271 gnd.n3934 gnd.n3933 585
R10272 gnd.n3932 gnd.n3931 585
R10273 gnd.n3930 gnd.n3929 585
R10274 gnd.n3928 gnd.n3927 585
R10275 gnd.n3926 gnd.n3925 585
R10276 gnd.n3924 gnd.n2246 585
R10277 gnd.n4041 gnd.n2245 585
R10278 gnd.n2049 gnd.n2048 585
R10279 gnd.n2047 gnd.n1958 585
R10280 gnd.n2046 gnd.n2045 585
R10281 gnd.n2039 gnd.n1959 585
R10282 gnd.n2041 gnd.n2040 585
R10283 gnd.n2038 gnd.n2037 585
R10284 gnd.n2036 gnd.n2035 585
R10285 gnd.n2029 gnd.n1961 585
R10286 gnd.n2031 gnd.n2030 585
R10287 gnd.n2028 gnd.n2027 585
R10288 gnd.n2026 gnd.n2025 585
R10289 gnd.n2019 gnd.n1963 585
R10290 gnd.n2021 gnd.n2020 585
R10291 gnd.n2018 gnd.n2017 585
R10292 gnd.n2016 gnd.n2015 585
R10293 gnd.n2009 gnd.n1965 585
R10294 gnd.n2011 gnd.n2010 585
R10295 gnd.n2008 gnd.n2007 585
R10296 gnd.n2006 gnd.n2005 585
R10297 gnd.n1999 gnd.n1967 585
R10298 gnd.n2001 gnd.n2000 585
R10299 gnd.n1998 gnd.n1971 585
R10300 gnd.n1997 gnd.n1996 585
R10301 gnd.n1990 gnd.n1972 585
R10302 gnd.n1992 gnd.n1991 585
R10303 gnd.n1989 gnd.n1988 585
R10304 gnd.n1987 gnd.n1986 585
R10305 gnd.n1980 gnd.n1974 585
R10306 gnd.n1982 gnd.n1981 585
R10307 gnd.n1979 gnd.n1978 585
R10308 gnd.n1977 gnd.n1045 585
R10309 gnd.n5903 gnd.n5902 585
R10310 gnd.n5905 gnd.n5904 585
R10311 gnd.n5907 gnd.n5906 585
R10312 gnd.n5909 gnd.n5908 585
R10313 gnd.n5911 gnd.n5910 585
R10314 gnd.n5913 gnd.n5912 585
R10315 gnd.n5915 gnd.n5914 585
R10316 gnd.n5917 gnd.n5916 585
R10317 gnd.n5920 gnd.n5919 585
R10318 gnd.n5922 gnd.n5921 585
R10319 gnd.n5924 gnd.n5923 585
R10320 gnd.n5926 gnd.n5925 585
R10321 gnd.n5928 gnd.n5927 585
R10322 gnd.n5930 gnd.n5929 585
R10323 gnd.n5932 gnd.n5931 585
R10324 gnd.n5934 gnd.n5933 585
R10325 gnd.n5936 gnd.n5935 585
R10326 gnd.n5938 gnd.n5937 585
R10327 gnd.n5940 gnd.n5939 585
R10328 gnd.n5942 gnd.n5941 585
R10329 gnd.n5944 gnd.n5943 585
R10330 gnd.n5946 gnd.n5945 585
R10331 gnd.n5947 gnd.n1018 585
R10332 gnd.n5949 gnd.n5948 585
R10333 gnd.n977 gnd.n976 585
R10334 gnd.n5953 gnd.n5952 585
R10335 gnd.n5952 gnd.n5951 585
R10336 gnd.n4376 gnd.n1852 585
R10337 gnd.n4468 gnd.n1852 585
R10338 gnd.n4375 gnd.n969 585
R10339 gnd.n5959 gnd.n969 585
R10340 gnd.n4374 gnd.n4373 585
R10341 gnd.n4373 gnd.n4372 585
R10342 gnd.n2051 gnd.n959 585
R10343 gnd.n5965 gnd.n959 585
R10344 gnd.n4361 gnd.n4360 585
R10345 gnd.n4362 gnd.n4361 585
R10346 gnd.n4358 gnd.n948 585
R10347 gnd.n5971 gnd.n948 585
R10348 gnd.n4357 gnd.n4356 585
R10349 gnd.n4356 gnd.n4355 585
R10350 gnd.n2056 gnd.n939 585
R10351 gnd.n5977 gnd.n939 585
R10352 gnd.n4346 gnd.n4345 585
R10353 gnd.n4347 gnd.n4346 585
R10354 gnd.n4343 gnd.n928 585
R10355 gnd.n5983 gnd.n928 585
R10356 gnd.n4342 gnd.n4341 585
R10357 gnd.n4341 gnd.n4340 585
R10358 gnd.n2061 gnd.n919 585
R10359 gnd.n5989 gnd.n919 585
R10360 gnd.n4282 gnd.n4281 585
R10361 gnd.n4283 gnd.n4282 585
R10362 gnd.n4279 gnd.n908 585
R10363 gnd.n5995 gnd.n908 585
R10364 gnd.n4278 gnd.n2068 585
R10365 gnd.n4294 gnd.n2068 585
R10366 gnd.n4277 gnd.n897 585
R10367 gnd.n6001 gnd.n897 585
R10368 gnd.n4276 gnd.n4275 585
R10369 gnd.n4275 gnd.n4274 585
R10370 gnd.n2073 gnd.n884 585
R10371 gnd.n6007 gnd.n884 585
R10372 gnd.n4246 gnd.n4245 585
R10373 gnd.n4245 gnd.n883 585
R10374 gnd.n4244 gnd.n2079 585
R10375 gnd.n4265 gnd.n2079 585
R10376 gnd.n4243 gnd.n4242 585
R10377 gnd.n4242 gnd.n2089 585
R10378 gnd.n4241 gnd.n2087 585
R10379 gnd.n4256 gnd.n2087 585
R10380 gnd.n4240 gnd.n4239 585
R10381 gnd.n4239 gnd.n2086 585
R10382 gnd.n4238 gnd.n2096 585
R10383 gnd.n4238 gnd.n4237 585
R10384 gnd.n4222 gnd.n2098 585
R10385 gnd.n2099 gnd.n2098 585
R10386 gnd.n4221 gnd.n2107 585
R10387 gnd.n4229 gnd.n2107 585
R10388 gnd.n4220 gnd.n4219 585
R10389 gnd.n4219 gnd.n4218 585
R10390 gnd.n2115 gnd.n2113 585
R10391 gnd.n2116 gnd.n2115 585
R10392 gnd.n4177 gnd.n2124 585
R10393 gnd.n4196 gnd.n2124 585
R10394 gnd.n4176 gnd.n4175 585
R10395 gnd.n4175 gnd.n2123 585
R10396 gnd.n4174 gnd.n2132 585
R10397 gnd.n4186 gnd.n2132 585
R10398 gnd.n4173 gnd.n4172 585
R10399 gnd.n4172 gnd.n4171 585
R10400 gnd.n2141 gnd.n2139 585
R10401 gnd.n2142 gnd.n2141 585
R10402 gnd.n4142 gnd.n2148 585
R10403 gnd.n4161 gnd.n2148 585
R10404 gnd.n4141 gnd.n4140 585
R10405 gnd.n4140 gnd.n2158 585
R10406 gnd.n4139 gnd.n2156 585
R10407 gnd.n4151 gnd.n2156 585
R10408 gnd.n4138 gnd.n4137 585
R10409 gnd.n4137 gnd.n4136 585
R10410 gnd.n2166 gnd.n2164 585
R10411 gnd.n2167 gnd.n2166 585
R10412 gnd.n4107 gnd.n2173 585
R10413 gnd.n4126 gnd.n2173 585
R10414 gnd.n4106 gnd.n4105 585
R10415 gnd.n4105 gnd.n2184 585
R10416 gnd.n4104 gnd.n2182 585
R10417 gnd.n4116 gnd.n2182 585
R10418 gnd.n4103 gnd.n4102 585
R10419 gnd.n4102 gnd.n2181 585
R10420 gnd.n4101 gnd.n2190 585
R10421 gnd.n4101 gnd.n4100 585
R10422 gnd.n4085 gnd.n2192 585
R10423 gnd.n2193 gnd.n2192 585
R10424 gnd.n4084 gnd.n2202 585
R10425 gnd.n4092 gnd.n2202 585
R10426 gnd.n4083 gnd.n4082 585
R10427 gnd.n4082 gnd.n2201 585
R10428 gnd.n4081 gnd.n2208 585
R10429 gnd.n4081 gnd.n4080 585
R10430 gnd.n4065 gnd.n2210 585
R10431 gnd.n2221 gnd.n2210 585
R10432 gnd.n4064 gnd.n2219 585
R10433 gnd.n4072 gnd.n2219 585
R10434 gnd.n4063 gnd.n4062 585
R10435 gnd.n4062 gnd.n2218 585
R10436 gnd.n4061 gnd.n2226 585
R10437 gnd.n4061 gnd.n4060 585
R10438 gnd.n4045 gnd.n2228 585
R10439 gnd.n2229 gnd.n2228 585
R10440 gnd.n4044 gnd.n2238 585
R10441 gnd.n4052 gnd.n2238 585
R10442 gnd.n4043 gnd.n4042 585
R10443 gnd.n4042 gnd.n2237 585
R10444 gnd.n7116 gnd.n205 585
R10445 gnd.n205 gnd.n204 585
R10446 gnd.n7118 gnd.n7117 585
R10447 gnd.n7119 gnd.n7118 585
R10448 gnd.n192 gnd.n191 585
R10449 gnd.n195 gnd.n192 585
R10450 gnd.n7127 gnd.n7126 585
R10451 gnd.n7126 gnd.n7125 585
R10452 gnd.n7128 gnd.n186 585
R10453 gnd.n186 gnd.n185 585
R10454 gnd.n7130 gnd.n7129 585
R10455 gnd.n7131 gnd.n7130 585
R10456 gnd.n173 gnd.n172 585
R10457 gnd.n182 gnd.n173 585
R10458 gnd.n7139 gnd.n7138 585
R10459 gnd.n7138 gnd.n7137 585
R10460 gnd.n7140 gnd.n167 585
R10461 gnd.n167 gnd.n166 585
R10462 gnd.n7142 gnd.n7141 585
R10463 gnd.n7143 gnd.n7142 585
R10464 gnd.n154 gnd.n153 585
R10465 gnd.n6969 gnd.n154 585
R10466 gnd.n7151 gnd.n7150 585
R10467 gnd.n7150 gnd.n7149 585
R10468 gnd.n7152 gnd.n148 585
R10469 gnd.n148 gnd.n147 585
R10470 gnd.n7154 gnd.n7153 585
R10471 gnd.n7155 gnd.n7154 585
R10472 gnd.n135 gnd.n134 585
R10473 gnd.n144 gnd.n135 585
R10474 gnd.n7163 gnd.n7162 585
R10475 gnd.n7162 gnd.n7161 585
R10476 gnd.n7164 gnd.n129 585
R10477 gnd.n129 gnd.n128 585
R10478 gnd.n7166 gnd.n7165 585
R10479 gnd.n7167 gnd.n7166 585
R10480 gnd.n116 gnd.n115 585
R10481 gnd.n119 gnd.n116 585
R10482 gnd.n7175 gnd.n7174 585
R10483 gnd.n7174 gnd.n7173 585
R10484 gnd.n7176 gnd.n110 585
R10485 gnd.n110 gnd.n109 585
R10486 gnd.n7178 gnd.n7177 585
R10487 gnd.n7179 gnd.n7178 585
R10488 gnd.n95 gnd.n94 585
R10489 gnd.n106 gnd.n95 585
R10490 gnd.n7187 gnd.n7186 585
R10491 gnd.n7186 gnd.n7185 585
R10492 gnd.n7188 gnd.n89 585
R10493 gnd.n89 gnd.n86 585
R10494 gnd.n7190 gnd.n7189 585
R10495 gnd.n7191 gnd.n7190 585
R10496 gnd.n90 gnd.n88 585
R10497 gnd.n6821 gnd.n88 585
R10498 gnd.n6810 gnd.n324 585
R10499 gnd.n324 gnd.n313 585
R10500 gnd.n6812 gnd.n6811 585
R10501 gnd.n6813 gnd.n6812 585
R10502 gnd.n325 gnd.n323 585
R10503 gnd.n323 gnd.n319 585
R10504 gnd.n6804 gnd.n6803 585
R10505 gnd.n6803 gnd.n6802 585
R10506 gnd.n328 gnd.n327 585
R10507 gnd.n6793 gnd.n328 585
R10508 gnd.n6776 gnd.n346 585
R10509 gnd.n346 gnd.n336 585
R10510 gnd.n6778 gnd.n6777 585
R10511 gnd.n6779 gnd.n6778 585
R10512 gnd.n347 gnd.n345 585
R10513 gnd.n354 gnd.n345 585
R10514 gnd.n6771 gnd.n6770 585
R10515 gnd.n6770 gnd.n6769 585
R10516 gnd.n350 gnd.n349 585
R10517 gnd.n6754 gnd.n350 585
R10518 gnd.n6742 gnd.n374 585
R10519 gnd.n6728 gnd.n374 585
R10520 gnd.n6744 gnd.n6743 585
R10521 gnd.n6745 gnd.n6744 585
R10522 gnd.n375 gnd.n373 585
R10523 gnd.n6722 gnd.n373 585
R10524 gnd.n6737 gnd.n6736 585
R10525 gnd.n6736 gnd.n6735 585
R10526 gnd.n378 gnd.n377 585
R10527 gnd.n5417 gnd.n378 585
R10528 gnd.n5442 gnd.n5441 585
R10529 gnd.n5443 gnd.n5442 585
R10530 gnd.n5326 gnd.n5325 585
R10531 gnd.n5426 gnd.n5326 585
R10532 gnd.n5451 gnd.n5450 585
R10533 gnd.n5450 gnd.n5449 585
R10534 gnd.n5452 gnd.n5320 585
R10535 gnd.n5408 gnd.n5320 585
R10536 gnd.n5454 gnd.n5453 585
R10537 gnd.n5455 gnd.n5454 585
R10538 gnd.n5304 gnd.n5303 585
R10539 gnd.n5400 gnd.n5304 585
R10540 gnd.n5463 gnd.n5462 585
R10541 gnd.n5462 gnd.n5461 585
R10542 gnd.n5464 gnd.n5292 585
R10543 gnd.n5380 gnd.n5292 585
R10544 gnd.n5466 gnd.n5465 585
R10545 gnd.n5467 gnd.n5466 585
R10546 gnd.n5293 gnd.n5291 585
R10547 gnd.n5291 gnd.n5286 585
R10548 gnd.n5297 gnd.n5296 585
R10549 gnd.n5296 gnd.n5274 585
R10550 gnd.n5295 gnd.n1281 585
R10551 gnd.n5475 gnd.n1281 585
R10552 gnd.n5706 gnd.n5705 585
R10553 gnd.n5704 gnd.n1280 585
R10554 gnd.n5703 gnd.n1279 585
R10555 gnd.n5708 gnd.n1279 585
R10556 gnd.n5702 gnd.n5701 585
R10557 gnd.n5700 gnd.n5699 585
R10558 gnd.n5698 gnd.n5697 585
R10559 gnd.n5696 gnd.n5695 585
R10560 gnd.n5694 gnd.n5693 585
R10561 gnd.n5692 gnd.n5691 585
R10562 gnd.n5690 gnd.n5689 585
R10563 gnd.n5688 gnd.n5687 585
R10564 gnd.n5686 gnd.n5685 585
R10565 gnd.n5684 gnd.n5683 585
R10566 gnd.n5682 gnd.n5681 585
R10567 gnd.n5680 gnd.n5679 585
R10568 gnd.n5678 gnd.n5677 585
R10569 gnd.n5676 gnd.n5675 585
R10570 gnd.n5674 gnd.n5673 585
R10571 gnd.n5671 gnd.n5670 585
R10572 gnd.n5669 gnd.n5668 585
R10573 gnd.n5667 gnd.n5666 585
R10574 gnd.n5665 gnd.n5664 585
R10575 gnd.n5663 gnd.n5662 585
R10576 gnd.n5661 gnd.n5660 585
R10577 gnd.n5659 gnd.n5658 585
R10578 gnd.n5657 gnd.n5656 585
R10579 gnd.n5654 gnd.n5653 585
R10580 gnd.n5652 gnd.n5651 585
R10581 gnd.n5650 gnd.n5649 585
R10582 gnd.n5648 gnd.n5647 585
R10583 gnd.n5646 gnd.n5645 585
R10584 gnd.n5644 gnd.n5643 585
R10585 gnd.n5642 gnd.n5641 585
R10586 gnd.n5640 gnd.n5639 585
R10587 gnd.n5638 gnd.n5637 585
R10588 gnd.n5636 gnd.n5635 585
R10589 gnd.n5634 gnd.n5633 585
R10590 gnd.n5632 gnd.n5631 585
R10591 gnd.n5630 gnd.n5629 585
R10592 gnd.n5628 gnd.n5627 585
R10593 gnd.n5626 gnd.n5625 585
R10594 gnd.n5624 gnd.n5623 585
R10595 gnd.n5622 gnd.n5621 585
R10596 gnd.n5620 gnd.n5619 585
R10597 gnd.n5618 gnd.n5617 585
R10598 gnd.n5616 gnd.n5615 585
R10599 gnd.n5614 gnd.n5613 585
R10600 gnd.n5612 gnd.n5611 585
R10601 gnd.n5610 gnd.n5609 585
R10602 gnd.n5608 gnd.n5607 585
R10603 gnd.n5606 gnd.n5605 585
R10604 gnd.n5604 gnd.n5603 585
R10605 gnd.n5602 gnd.n5601 585
R10606 gnd.n5600 gnd.n5599 585
R10607 gnd.n5598 gnd.n5597 585
R10608 gnd.n5596 gnd.n5595 585
R10609 gnd.n5271 gnd.n1344 585
R10610 gnd.n6987 gnd.n305 585
R10611 gnd.n6995 gnd.n6994 585
R10612 gnd.n6997 gnd.n6996 585
R10613 gnd.n6999 gnd.n6998 585
R10614 gnd.n7001 gnd.n7000 585
R10615 gnd.n7003 gnd.n7002 585
R10616 gnd.n7005 gnd.n7004 585
R10617 gnd.n7007 gnd.n7006 585
R10618 gnd.n7009 gnd.n7008 585
R10619 gnd.n7011 gnd.n7010 585
R10620 gnd.n7013 gnd.n7012 585
R10621 gnd.n7015 gnd.n7014 585
R10622 gnd.n7017 gnd.n7016 585
R10623 gnd.n7019 gnd.n7018 585
R10624 gnd.n7021 gnd.n7020 585
R10625 gnd.n7023 gnd.n7022 585
R10626 gnd.n7025 gnd.n7024 585
R10627 gnd.n7027 gnd.n7026 585
R10628 gnd.n7029 gnd.n7028 585
R10629 gnd.n7032 gnd.n7031 585
R10630 gnd.n7030 gnd.n285 585
R10631 gnd.n7037 gnd.n7036 585
R10632 gnd.n7039 gnd.n7038 585
R10633 gnd.n7041 gnd.n7040 585
R10634 gnd.n7043 gnd.n7042 585
R10635 gnd.n7045 gnd.n7044 585
R10636 gnd.n7047 gnd.n7046 585
R10637 gnd.n7049 gnd.n7048 585
R10638 gnd.n7051 gnd.n7050 585
R10639 gnd.n7053 gnd.n7052 585
R10640 gnd.n7055 gnd.n7054 585
R10641 gnd.n7057 gnd.n7056 585
R10642 gnd.n7059 gnd.n7058 585
R10643 gnd.n7061 gnd.n7060 585
R10644 gnd.n7063 gnd.n7062 585
R10645 gnd.n7065 gnd.n7064 585
R10646 gnd.n7067 gnd.n7066 585
R10647 gnd.n7069 gnd.n7068 585
R10648 gnd.n7071 gnd.n7070 585
R10649 gnd.n7073 gnd.n7072 585
R10650 gnd.n7075 gnd.n7074 585
R10651 gnd.n7080 gnd.n7079 585
R10652 gnd.n7082 gnd.n7081 585
R10653 gnd.n7084 gnd.n7083 585
R10654 gnd.n7086 gnd.n7085 585
R10655 gnd.n7088 gnd.n7087 585
R10656 gnd.n7090 gnd.n7089 585
R10657 gnd.n7092 gnd.n7091 585
R10658 gnd.n7094 gnd.n7093 585
R10659 gnd.n7096 gnd.n7095 585
R10660 gnd.n7098 gnd.n7097 585
R10661 gnd.n7100 gnd.n7099 585
R10662 gnd.n7102 gnd.n7101 585
R10663 gnd.n7104 gnd.n7103 585
R10664 gnd.n7106 gnd.n7105 585
R10665 gnd.n7107 gnd.n249 585
R10666 gnd.n7109 gnd.n7108 585
R10667 gnd.n210 gnd.n209 585
R10668 gnd.n7113 gnd.n7112 585
R10669 gnd.n7112 gnd.n7111 585
R10670 gnd.n6989 gnd.n6988 585
R10671 gnd.n6988 gnd.n204 585
R10672 gnd.n6986 gnd.n202 585
R10673 gnd.n7119 gnd.n202 585
R10674 gnd.n6985 gnd.n6984 585
R10675 gnd.n6984 gnd.n195 585
R10676 gnd.n6983 gnd.n193 585
R10677 gnd.n7125 gnd.n193 585
R10678 gnd.n6982 gnd.n6981 585
R10679 gnd.n6981 gnd.n185 585
R10680 gnd.n6979 gnd.n183 585
R10681 gnd.n7131 gnd.n183 585
R10682 gnd.n6978 gnd.n6977 585
R10683 gnd.n6977 gnd.n182 585
R10684 gnd.n6976 gnd.n174 585
R10685 gnd.n7137 gnd.n174 585
R10686 gnd.n6975 gnd.n6974 585
R10687 gnd.n6974 gnd.n166 585
R10688 gnd.n6972 gnd.n164 585
R10689 gnd.n7143 gnd.n164 585
R10690 gnd.n6971 gnd.n6970 585
R10691 gnd.n6970 gnd.n6969 585
R10692 gnd.n6850 gnd.n155 585
R10693 gnd.n7149 gnd.n155 585
R10694 gnd.n6849 gnd.n6848 585
R10695 gnd.n6848 gnd.n147 585
R10696 gnd.n6846 gnd.n145 585
R10697 gnd.n7155 gnd.n145 585
R10698 gnd.n6845 gnd.n6844 585
R10699 gnd.n6844 gnd.n144 585
R10700 gnd.n6843 gnd.n136 585
R10701 gnd.n7161 gnd.n136 585
R10702 gnd.n6842 gnd.n6841 585
R10703 gnd.n6841 gnd.n128 585
R10704 gnd.n6839 gnd.n126 585
R10705 gnd.n7167 gnd.n126 585
R10706 gnd.n6838 gnd.n6837 585
R10707 gnd.n6837 gnd.n119 585
R10708 gnd.n6836 gnd.n117 585
R10709 gnd.n7173 gnd.n117 585
R10710 gnd.n6835 gnd.n6834 585
R10711 gnd.n6834 gnd.n109 585
R10712 gnd.n6832 gnd.n107 585
R10713 gnd.n7179 gnd.n107 585
R10714 gnd.n6831 gnd.n6830 585
R10715 gnd.n6830 gnd.n106 585
R10716 gnd.n6829 gnd.n96 585
R10717 gnd.n7185 gnd.n96 585
R10718 gnd.n6828 gnd.n6827 585
R10719 gnd.n6827 gnd.n86 585
R10720 gnd.n309 gnd.n85 585
R10721 gnd.n7191 gnd.n85 585
R10722 gnd.n6820 gnd.n6819 585
R10723 gnd.n6821 gnd.n6820 585
R10724 gnd.n6818 gnd.n314 585
R10725 gnd.n314 gnd.n313 585
R10726 gnd.n320 gnd.n315 585
R10727 gnd.n6813 gnd.n320 585
R10728 gnd.n6797 gnd.n6796 585
R10729 gnd.n6796 gnd.n319 585
R10730 gnd.n6798 gnd.n329 585
R10731 gnd.n6802 gnd.n329 585
R10732 gnd.n6795 gnd.n6794 585
R10733 gnd.n6794 gnd.n6793 585
R10734 gnd.n335 gnd.n334 585
R10735 gnd.n336 gnd.n335 585
R10736 gnd.n6760 gnd.n343 585
R10737 gnd.n6779 gnd.n343 585
R10738 gnd.n6759 gnd.n6758 585
R10739 gnd.n6758 gnd.n354 585
R10740 gnd.n6757 gnd.n352 585
R10741 gnd.n6769 gnd.n352 585
R10742 gnd.n6756 gnd.n6755 585
R10743 gnd.n6755 gnd.n6754 585
R10744 gnd.n362 gnd.n360 585
R10745 gnd.n6728 gnd.n362 585
R10746 gnd.n6725 gnd.n370 585
R10747 gnd.n6745 gnd.n370 585
R10748 gnd.n6724 gnd.n6723 585
R10749 gnd.n6723 gnd.n6722 585
R10750 gnd.n388 gnd.n380 585
R10751 gnd.n6735 gnd.n380 585
R10752 gnd.n5416 gnd.n5415 585
R10753 gnd.n5417 gnd.n5416 585
R10754 gnd.n5413 gnd.n5335 585
R10755 gnd.n5443 gnd.n5335 585
R10756 gnd.n5412 gnd.n5343 585
R10757 gnd.n5426 gnd.n5343 585
R10758 gnd.n5411 gnd.n5328 585
R10759 gnd.n5449 gnd.n5328 585
R10760 gnd.n5410 gnd.n5409 585
R10761 gnd.n5409 gnd.n5408 585
R10762 gnd.n5348 gnd.n5317 585
R10763 gnd.n5455 gnd.n5317 585
R10764 gnd.n5385 gnd.n5384 585
R10765 gnd.n5400 gnd.n5385 585
R10766 gnd.n5383 gnd.n5306 585
R10767 gnd.n5461 gnd.n5306 585
R10768 gnd.n5382 gnd.n5381 585
R10769 gnd.n5381 gnd.n5380 585
R10770 gnd.n5353 gnd.n5287 585
R10771 gnd.n5467 gnd.n5287 585
R10772 gnd.n5358 gnd.n5357 585
R10773 gnd.n5357 gnd.n5286 585
R10774 gnd.n5359 gnd.n5356 585
R10775 gnd.n5356 gnd.n5274 585
R10776 gnd.n5355 gnd.n5272 585
R10777 gnd.n5475 gnd.n5272 585
R10778 gnd.n6010 gnd.n6009 585
R10779 gnd.n6009 gnd.n6008 585
R10780 gnd.n6715 gnd.n6714 585
R10781 gnd.n6715 gnd.n351 585
R10782 gnd.n6717 gnd.n6716 585
R10783 gnd.n6716 gnd.n363 585
R10784 gnd.n6718 gnd.n390 585
R10785 gnd.n390 gnd.n371 585
R10786 gnd.n6720 gnd.n6719 585
R10787 gnd.n6721 gnd.n6720 585
R10788 gnd.n391 gnd.n389 585
R10789 gnd.n389 gnd.n382 585
R10790 gnd.n5435 gnd.n5338 585
R10791 gnd.n5338 gnd.n379 585
R10792 gnd.n5437 gnd.n5436 585
R10793 gnd.n5438 gnd.n5437 585
R10794 gnd.n5339 gnd.n5337 585
R10795 gnd.n5337 gnd.n5334 585
R10796 gnd.n5429 gnd.n5428 585
R10797 gnd.n5428 gnd.n5427 585
R10798 gnd.n5342 gnd.n5341 585
R10799 gnd.n5342 gnd.n5327 585
R10800 gnd.n5396 gnd.n5387 585
R10801 gnd.n5387 gnd.n5319 585
R10802 gnd.n5398 gnd.n5397 585
R10803 gnd.n5399 gnd.n5398 585
R10804 gnd.n5388 gnd.n5386 585
R10805 gnd.n5386 gnd.n5308 585
R10806 gnd.n5391 gnd.n5390 585
R10807 gnd.n5390 gnd.n5305 585
R10808 gnd.n5284 gnd.n5283 585
R10809 gnd.n5289 gnd.n5284 585
R10810 gnd.n5470 gnd.n5469 585
R10811 gnd.n5469 gnd.n5468 585
R10812 gnd.n5471 gnd.n5276 585
R10813 gnd.n5285 gnd.n5276 585
R10814 gnd.n5473 gnd.n5472 585
R10815 gnd.n5474 gnd.n5473 585
R10816 gnd.n5277 gnd.n5275 585
R10817 gnd.n5275 gnd.n5270 585
R10818 gnd.n1239 gnd.n1238 585
R10819 gnd.n1278 gnd.n1239 585
R10820 gnd.n5711 gnd.n5710 585
R10821 gnd.n5710 gnd.n5709 585
R10822 gnd.n5712 gnd.n1233 585
R10823 gnd.n1233 gnd.n1231 585
R10824 gnd.n5714 gnd.n5713 585
R10825 gnd.n5715 gnd.n5714 585
R10826 gnd.n1234 gnd.n1232 585
R10827 gnd.n1232 gnd.n1216 585
R10828 gnd.n5240 gnd.n5239 585
R10829 gnd.n5241 gnd.n5240 585
R10830 gnd.n1359 gnd.n1358 585
R10831 gnd.n1358 gnd.n1357 585
R10832 gnd.n5234 gnd.n5233 585
R10833 gnd.n5233 gnd.n5232 585
R10834 gnd.n1362 gnd.n1361 585
R10835 gnd.n1363 gnd.n1362 585
R10836 gnd.n5223 gnd.n5222 585
R10837 gnd.n5224 gnd.n5223 585
R10838 gnd.n1372 gnd.n1371 585
R10839 gnd.n1371 gnd.n1369 585
R10840 gnd.n5218 gnd.n5217 585
R10841 gnd.n5217 gnd.n5216 585
R10842 gnd.n1375 gnd.n1374 585
R10843 gnd.n1382 gnd.n1375 585
R10844 gnd.n5207 gnd.n5206 585
R10845 gnd.n5208 gnd.n5207 585
R10846 gnd.n1385 gnd.n1384 585
R10847 gnd.n1384 gnd.n1381 585
R10848 gnd.n5202 gnd.n5201 585
R10849 gnd.n5201 gnd.n5200 585
R10850 gnd.n1388 gnd.n1387 585
R10851 gnd.n1395 gnd.n1388 585
R10852 gnd.n5191 gnd.n5190 585
R10853 gnd.n5192 gnd.n5191 585
R10854 gnd.n1398 gnd.n1397 585
R10855 gnd.n1405 gnd.n1397 585
R10856 gnd.n5186 gnd.n5185 585
R10857 gnd.n5185 gnd.n5184 585
R10858 gnd.n1401 gnd.n1400 585
R10859 gnd.n1480 gnd.n1401 585
R10860 gnd.n5048 gnd.n5047 585
R10861 gnd.n5049 gnd.n5048 585
R10862 gnd.n1489 gnd.n1488 585
R10863 gnd.n1496 gnd.n1488 585
R10864 gnd.n5043 gnd.n5042 585
R10865 gnd.n5042 gnd.n5041 585
R10866 gnd.n1492 gnd.n1491 585
R10867 gnd.n1500 gnd.n1492 585
R10868 gnd.n5011 gnd.n1513 585
R10869 gnd.n4969 gnd.n1513 585
R10870 gnd.n5013 gnd.n5012 585
R10871 gnd.n5014 gnd.n5013 585
R10872 gnd.n1514 gnd.n1512 585
R10873 gnd.n1512 gnd.n1509 585
R10874 gnd.n5006 gnd.n5005 585
R10875 gnd.n5005 gnd.n5004 585
R10876 gnd.n1517 gnd.n1516 585
R10877 gnd.n4996 gnd.n1517 585
R10878 gnd.n4957 gnd.n1534 585
R10879 gnd.n4874 gnd.n1534 585
R10880 gnd.n4959 gnd.n4958 585
R10881 gnd.n4960 gnd.n4959 585
R10882 gnd.n1535 gnd.n1533 585
R10883 gnd.n1542 gnd.n1533 585
R10884 gnd.n4952 gnd.n4951 585
R10885 gnd.n4951 gnd.n4950 585
R10886 gnd.n1538 gnd.n1537 585
R10887 gnd.n4936 gnd.n1538 585
R10888 gnd.n4924 gnd.n1558 585
R10889 gnd.n4870 gnd.n1558 585
R10890 gnd.n4926 gnd.n4925 585
R10891 gnd.n4927 gnd.n4926 585
R10892 gnd.n1559 gnd.n1557 585
R10893 gnd.n1567 gnd.n1557 585
R10894 gnd.n4919 gnd.n4918 585
R10895 gnd.n4918 gnd.n4917 585
R10896 gnd.n1562 gnd.n1561 585
R10897 gnd.n1572 gnd.n1562 585
R10898 gnd.n4855 gnd.n1588 585
R10899 gnd.n1588 gnd.n1579 585
R10900 gnd.n4857 gnd.n4856 585
R10901 gnd.n4858 gnd.n4857 585
R10902 gnd.n1589 gnd.n1587 585
R10903 gnd.n1587 gnd.n1583 585
R10904 gnd.n4850 gnd.n4849 585
R10905 gnd.n4849 gnd.n4848 585
R10906 gnd.n1592 gnd.n1591 585
R10907 gnd.n4840 gnd.n1592 585
R10908 gnd.n4815 gnd.n1613 585
R10909 gnd.n1613 gnd.n1612 585
R10910 gnd.n4817 gnd.n4816 585
R10911 gnd.n4818 gnd.n4817 585
R10912 gnd.n1614 gnd.n1610 585
R10913 gnd.n1620 gnd.n1610 585
R10914 gnd.n4810 gnd.n4809 585
R10915 gnd.n4809 gnd.n4808 585
R10916 gnd.n1617 gnd.n1616 585
R10917 gnd.n4795 gnd.n1617 585
R10918 gnd.n4759 gnd.n1639 585
R10919 gnd.n1639 gnd.n1631 585
R10920 gnd.n4761 gnd.n4760 585
R10921 gnd.n4762 gnd.n4761 585
R10922 gnd.n1640 gnd.n1638 585
R10923 gnd.n1638 gnd.n1635 585
R10924 gnd.n4754 gnd.n4753 585
R10925 gnd.n4753 gnd.n4752 585
R10926 gnd.n1643 gnd.n1642 585
R10927 gnd.n1649 gnd.n1643 585
R10928 gnd.n4733 gnd.n4732 585
R10929 gnd.n4734 gnd.n4733 585
R10930 gnd.n1658 gnd.n1657 585
R10931 gnd.n1665 gnd.n1657 585
R10932 gnd.n4728 gnd.n4727 585
R10933 gnd.n4727 gnd.n4726 585
R10934 gnd.n1661 gnd.n1660 585
R10935 gnd.n1669 gnd.n1661 585
R10936 gnd.n4697 gnd.n1685 585
R10937 gnd.n1685 gnd.n1676 585
R10938 gnd.n4699 gnd.n4698 585
R10939 gnd.n4700 gnd.n4699 585
R10940 gnd.n1686 gnd.n1684 585
R10941 gnd.n1684 gnd.n1681 585
R10942 gnd.n4692 gnd.n4691 585
R10943 gnd.n4691 gnd.n4690 585
R10944 gnd.n1689 gnd.n1688 585
R10945 gnd.n4682 gnd.n1689 585
R10946 gnd.n4659 gnd.n4658 585
R10947 gnd.n4658 gnd.n1696 585
R10948 gnd.n4660 gnd.n1710 585
R10949 gnd.n1710 gnd.n1702 585
R10950 gnd.n4662 gnd.n4661 585
R10951 gnd.n4663 gnd.n4662 585
R10952 gnd.n1711 gnd.n1709 585
R10953 gnd.n4563 gnd.n1709 585
R10954 gnd.n4652 gnd.n4651 585
R10955 gnd.n4651 gnd.n4650 585
R10956 gnd.n1123 gnd.n1122 585
R10957 gnd.n4561 gnd.n1123 585
R10958 gnd.n5821 gnd.n5820 585
R10959 gnd.n5820 gnd.n5819 585
R10960 gnd.n5822 gnd.n1117 585
R10961 gnd.n4621 gnd.n1117 585
R10962 gnd.n5824 gnd.n5823 585
R10963 gnd.n5825 gnd.n5824 585
R10964 gnd.n1118 gnd.n1116 585
R10965 gnd.n1116 gnd.n1110 585
R10966 gnd.n4541 gnd.n4540 585
R10967 gnd.n4541 gnd.n1084 585
R10968 gnd.n4543 gnd.n4542 585
R10969 gnd.n4542 gnd.n1052 585
R10970 gnd.n4544 gnd.n1806 585
R10971 gnd.n4510 gnd.n1806 585
R10972 gnd.n4546 gnd.n4545 585
R10973 gnd.n4547 gnd.n4546 585
R10974 gnd.n1807 gnd.n1805 585
R10975 gnd.n1805 gnd.n1803 585
R10976 gnd.n4532 gnd.n4531 585
R10977 gnd.n4531 gnd.n4530 585
R10978 gnd.n1810 gnd.n1809 585
R10979 gnd.n1811 gnd.n1810 585
R10980 gnd.n4503 gnd.n4502 585
R10981 gnd.n4504 gnd.n4503 585
R10982 gnd.n1823 gnd.n1822 585
R10983 gnd.n1822 gnd.n1820 585
R10984 gnd.n4498 gnd.n4497 585
R10985 gnd.n4497 gnd.n4496 585
R10986 gnd.n1826 gnd.n1825 585
R10987 gnd.n1827 gnd.n1826 585
R10988 gnd.n4487 gnd.n4486 585
R10989 gnd.n4488 gnd.n4487 585
R10990 gnd.n1836 gnd.n1835 585
R10991 gnd.n1842 gnd.n1835 585
R10992 gnd.n4482 gnd.n4481 585
R10993 gnd.n4481 gnd.n4480 585
R10994 gnd.n1839 gnd.n1838 585
R10995 gnd.n1840 gnd.n1839 585
R10996 gnd.n1863 gnd.n1862 585
R10997 gnd.n4459 gnd.n1863 585
R10998 gnd.n4461 gnd.n1859 585
R10999 gnd.n4461 gnd.n4460 585
R11000 gnd.n4463 gnd.n4462 585
R11001 gnd.n4462 gnd.n989 585
R11002 gnd.n4464 gnd.n1854 585
R11003 gnd.n1854 gnd.n978 585
R11004 gnd.n4466 gnd.n4465 585
R11005 gnd.n4467 gnd.n4466 585
R11006 gnd.n1855 gnd.n1853 585
R11007 gnd.n1853 gnd.n971 585
R11008 gnd.n4326 gnd.n4325 585
R11009 gnd.n4326 gnd.n968 585
R11010 gnd.n4327 gnd.n4321 585
R11011 gnd.n4327 gnd.n961 585
R11012 gnd.n4329 gnd.n4328 585
R11013 gnd.n4328 gnd.n958 585
R11014 gnd.n4330 gnd.n4316 585
R11015 gnd.n4316 gnd.n950 585
R11016 gnd.n4332 gnd.n4331 585
R11017 gnd.n4332 gnd.n947 585
R11018 gnd.n4333 gnd.n4315 585
R11019 gnd.n4333 gnd.n2057 585
R11020 gnd.n4335 gnd.n4334 585
R11021 gnd.n4334 gnd.n938 585
R11022 gnd.n4336 gnd.n2064 585
R11023 gnd.n2064 gnd.n930 585
R11024 gnd.n4338 gnd.n4337 585
R11025 gnd.n4339 gnd.n4338 585
R11026 gnd.n2065 gnd.n2063 585
R11027 gnd.n2063 gnd.n921 585
R11028 gnd.n4309 gnd.n4308 585
R11029 gnd.n4308 gnd.n918 585
R11030 gnd.n4307 gnd.n2067 585
R11031 gnd.n4307 gnd.n910 585
R11032 gnd.n4306 gnd.n4305 585
R11033 gnd.n4306 gnd.n907 585
R11034 gnd.n4297 gnd.n4296 585
R11035 gnd.n4296 gnd.n4295 585
R11036 gnd.n4301 gnd.n4300 585
R11037 gnd.n4300 gnd.n896 585
R11038 gnd.n4299 gnd.n882 585
R11039 gnd.n886 gnd.n882 585
R11040 gnd.n5243 gnd.n5242 585
R11041 gnd.n5242 gnd.n5241 585
R11042 gnd.n1355 gnd.n1354 585
R11043 gnd.n1357 gnd.n1355 585
R11044 gnd.n5231 gnd.n5230 585
R11045 gnd.n5232 gnd.n5231 585
R11046 gnd.n1365 gnd.n1364 585
R11047 gnd.n1364 gnd.n1363 585
R11048 gnd.n5226 gnd.n5225 585
R11049 gnd.n5225 gnd.n5224 585
R11050 gnd.n1368 gnd.n1367 585
R11051 gnd.n1369 gnd.n1368 585
R11052 gnd.n5215 gnd.n5214 585
R11053 gnd.n5216 gnd.n5215 585
R11054 gnd.n1377 gnd.n1376 585
R11055 gnd.n1382 gnd.n1376 585
R11056 gnd.n5210 gnd.n5209 585
R11057 gnd.n5209 gnd.n5208 585
R11058 gnd.n1380 gnd.n1379 585
R11059 gnd.n1381 gnd.n1380 585
R11060 gnd.n5199 gnd.n5198 585
R11061 gnd.n5200 gnd.n5199 585
R11062 gnd.n1390 gnd.n1389 585
R11063 gnd.n1395 gnd.n1389 585
R11064 gnd.n5194 gnd.n5193 585
R11065 gnd.n5193 gnd.n5192 585
R11066 gnd.n1393 gnd.n1392 585
R11067 gnd.n1405 gnd.n1393 585
R11068 gnd.n4977 gnd.n1403 585
R11069 gnd.n5184 gnd.n1403 585
R11070 gnd.n4976 gnd.n4975 585
R11071 gnd.n4975 gnd.n1480 585
R11072 gnd.n4981 gnd.n1485 585
R11073 gnd.n5049 gnd.n1485 585
R11074 gnd.n4982 gnd.n4974 585
R11075 gnd.n4974 gnd.n1496 585
R11076 gnd.n4983 gnd.n1494 585
R11077 gnd.n5041 gnd.n1494 585
R11078 gnd.n4972 gnd.n4971 585
R11079 gnd.n4971 gnd.n1500 585
R11080 gnd.n4987 gnd.n4970 585
R11081 gnd.n4970 gnd.n4969 585
R11082 gnd.n4988 gnd.n1511 585
R11083 gnd.n5014 gnd.n1511 585
R11084 gnd.n4989 gnd.n4966 585
R11085 gnd.n4966 gnd.n1509 585
R11086 gnd.n1528 gnd.n1519 585
R11087 gnd.n5004 gnd.n1519 585
R11088 gnd.n4994 gnd.n4993 585
R11089 gnd.n4996 gnd.n4994 585
R11090 gnd.n1527 gnd.n1526 585
R11091 gnd.n4874 gnd.n1526 585
R11092 gnd.n4962 gnd.n4961 585
R11093 gnd.n4961 gnd.n4960 585
R11094 gnd.n1531 gnd.n1530 585
R11095 gnd.n1542 gnd.n1531 585
R11096 gnd.n1551 gnd.n1540 585
R11097 gnd.n4950 gnd.n1540 585
R11098 gnd.n4935 gnd.n4934 585
R11099 gnd.n4936 gnd.n4935 585
R11100 gnd.n1550 gnd.n1549 585
R11101 gnd.n4870 gnd.n1549 585
R11102 gnd.n4929 gnd.n4928 585
R11103 gnd.n4928 gnd.n4927 585
R11104 gnd.n1554 gnd.n1553 585
R11105 gnd.n1567 gnd.n1554 585
R11106 gnd.n4828 gnd.n1564 585
R11107 gnd.n4917 gnd.n1564 585
R11108 gnd.n4827 gnd.n4826 585
R11109 gnd.n4826 gnd.n1572 585
R11110 gnd.n4832 gnd.n4825 585
R11111 gnd.n4825 gnd.n1579 585
R11112 gnd.n4833 gnd.n1585 585
R11113 gnd.n4858 gnd.n1585 585
R11114 gnd.n4834 gnd.n4824 585
R11115 gnd.n4824 gnd.n1583 585
R11116 gnd.n1604 gnd.n1594 585
R11117 gnd.n4848 gnd.n1594 585
R11118 gnd.n4839 gnd.n4838 585
R11119 gnd.n4840 gnd.n4839 585
R11120 gnd.n1603 gnd.n1602 585
R11121 gnd.n1612 gnd.n1602 585
R11122 gnd.n4820 gnd.n4819 585
R11123 gnd.n4819 gnd.n4818 585
R11124 gnd.n1607 gnd.n1606 585
R11125 gnd.n1620 gnd.n1607 585
R11126 gnd.n4584 gnd.n1618 585
R11127 gnd.n4808 gnd.n1618 585
R11128 gnd.n4585 gnd.n1628 585
R11129 gnd.n4795 gnd.n1628 585
R11130 gnd.n4582 gnd.n4581 585
R11131 gnd.n4581 gnd.n1631 585
R11132 gnd.n4589 gnd.n1637 585
R11133 gnd.n4762 gnd.n1637 585
R11134 gnd.n4590 gnd.n4580 585
R11135 gnd.n4580 gnd.n1635 585
R11136 gnd.n4591 gnd.n1645 585
R11137 gnd.n4752 gnd.n1645 585
R11138 gnd.n4578 gnd.n4577 585
R11139 gnd.n4577 gnd.n1649 585
R11140 gnd.n4595 gnd.n1655 585
R11141 gnd.n4734 gnd.n1655 585
R11142 gnd.n4596 gnd.n4576 585
R11143 gnd.n4576 gnd.n1665 585
R11144 gnd.n4597 gnd.n1663 585
R11145 gnd.n4726 gnd.n1663 585
R11146 gnd.n4574 gnd.n4573 585
R11147 gnd.n4573 gnd.n1669 585
R11148 gnd.n4601 gnd.n4572 585
R11149 gnd.n4572 gnd.n1676 585
R11150 gnd.n4602 gnd.n1683 585
R11151 gnd.n4700 gnd.n1683 585
R11152 gnd.n4603 gnd.n4571 585
R11153 gnd.n4571 gnd.n1681 585
R11154 gnd.n4569 gnd.n1690 585
R11155 gnd.n4690 gnd.n1690 585
R11156 gnd.n4607 gnd.n1698 585
R11157 gnd.n4682 gnd.n1698 585
R11158 gnd.n4608 gnd.n4568 585
R11159 gnd.n4568 gnd.n1696 585
R11160 gnd.n4609 gnd.n4567 585
R11161 gnd.n4567 gnd.n1702 585
R11162 gnd.n4565 gnd.n1708 585
R11163 gnd.n4663 gnd.n1708 585
R11164 gnd.n4613 gnd.n4564 585
R11165 gnd.n4564 gnd.n4563 585
R11166 gnd.n4614 gnd.n1714 585
R11167 gnd.n4650 gnd.n1714 585
R11168 gnd.n4615 gnd.n4562 585
R11169 gnd.n4562 gnd.n4561 585
R11170 gnd.n1795 gnd.n1125 585
R11171 gnd.n5819 gnd.n1125 585
R11172 gnd.n4620 gnd.n4619 585
R11173 gnd.n4621 gnd.n4620 585
R11174 gnd.n1794 gnd.n1113 585
R11175 gnd.n5825 gnd.n1113 585
R11176 gnd.n4557 gnd.n4556 585
R11177 gnd.n4556 gnd.n1110 585
R11178 gnd.n4555 gnd.n1797 585
R11179 gnd.n4555 gnd.n1084 585
R11180 gnd.n4554 gnd.n4553 585
R11181 gnd.n4554 gnd.n1052 585
R11182 gnd.n1799 gnd.n1798 585
R11183 gnd.n4510 gnd.n1798 585
R11184 gnd.n4549 gnd.n4548 585
R11185 gnd.n4548 gnd.n4547 585
R11186 gnd.n1802 gnd.n1801 585
R11187 gnd.n1803 gnd.n1802 585
R11188 gnd.n1929 gnd.n1812 585
R11189 gnd.n4530 gnd.n1812 585
R11190 gnd.n1928 gnd.n1927 585
R11191 gnd.n1927 gnd.n1811 585
R11192 gnd.n1933 gnd.n1821 585
R11193 gnd.n4504 gnd.n1821 585
R11194 gnd.n1934 gnd.n1926 585
R11195 gnd.n1926 gnd.n1820 585
R11196 gnd.n1935 gnd.n1828 585
R11197 gnd.n4496 gnd.n1828 585
R11198 gnd.n1924 gnd.n1923 585
R11199 gnd.n1923 gnd.n1827 585
R11200 gnd.n1939 gnd.n1834 585
R11201 gnd.n4488 gnd.n1834 585
R11202 gnd.n1940 gnd.n1922 585
R11203 gnd.n1922 gnd.n1842 585
R11204 gnd.n1941 gnd.n1841 585
R11205 gnd.n4480 gnd.n1841 585
R11206 gnd.n1944 gnd.n1943 585
R11207 gnd.n1919 gnd.n1918 585
R11208 gnd.n1948 gnd.n1920 585
R11209 gnd.n1950 gnd.n1949 585
R11210 gnd.n1952 gnd.n1951 585
R11211 gnd.n1915 gnd.n1914 585
R11212 gnd.n4381 gnd.n1916 585
R11213 gnd.n4383 gnd.n4382 585
R11214 gnd.n4385 gnd.n4384 585
R11215 gnd.n1910 gnd.n1909 585
R11216 gnd.n4393 gnd.n1911 585
R11217 gnd.n4396 gnd.n4395 585
R11218 gnd.n4394 gnd.n1903 585
R11219 gnd.n4406 gnd.n4405 585
R11220 gnd.n4408 gnd.n4407 585
R11221 gnd.n1898 gnd.n1897 585
R11222 gnd.n4417 gnd.n1899 585
R11223 gnd.n4420 gnd.n4419 585
R11224 gnd.n4418 gnd.n1891 585
R11225 gnd.n4430 gnd.n4429 585
R11226 gnd.n4432 gnd.n4431 585
R11227 gnd.n1886 gnd.n1885 585
R11228 gnd.n4441 gnd.n1887 585
R11229 gnd.n4445 gnd.n4442 585
R11230 gnd.n4444 gnd.n4443 585
R11231 gnd.n4456 gnd.n4455 585
R11232 gnd.n4457 gnd.n1845 585
R11233 gnd.n4474 gnd.n1846 585
R11234 gnd.n4475 gnd.n1843 585
R11235 gnd.n4459 gnd.n1843 585
R11236 gnd.n1215 gnd.n1211 585
R11237 gnd.n5241 gnd.n1215 585
R11238 gnd.n5721 gnd.n1210 585
R11239 gnd.n1357 gnd.n1210 585
R11240 gnd.n5722 gnd.n1209 585
R11241 gnd.n5232 gnd.n1209 585
R11242 gnd.n5723 gnd.n1208 585
R11243 gnd.n1363 gnd.n1208 585
R11244 gnd.n1370 gnd.n1206 585
R11245 gnd.n5224 gnd.n1370 585
R11246 gnd.n5727 gnd.n1205 585
R11247 gnd.n1369 gnd.n1205 585
R11248 gnd.n5728 gnd.n1204 585
R11249 gnd.n5216 gnd.n1204 585
R11250 gnd.n5729 gnd.n1203 585
R11251 gnd.n1382 gnd.n1203 585
R11252 gnd.n1383 gnd.n1201 585
R11253 gnd.n5208 gnd.n1383 585
R11254 gnd.n5733 gnd.n1200 585
R11255 gnd.n1381 gnd.n1200 585
R11256 gnd.n5734 gnd.n1199 585
R11257 gnd.n5200 gnd.n1199 585
R11258 gnd.n5735 gnd.n1198 585
R11259 gnd.n1395 gnd.n1198 585
R11260 gnd.n1396 gnd.n1196 585
R11261 gnd.n5192 gnd.n1396 585
R11262 gnd.n5739 gnd.n1195 585
R11263 gnd.n1405 gnd.n1195 585
R11264 gnd.n5740 gnd.n1194 585
R11265 gnd.n5184 gnd.n1194 585
R11266 gnd.n5741 gnd.n1193 585
R11267 gnd.n1480 gnd.n1193 585
R11268 gnd.n1487 gnd.n1191 585
R11269 gnd.n5049 gnd.n1487 585
R11270 gnd.n5745 gnd.n1190 585
R11271 gnd.n1496 gnd.n1190 585
R11272 gnd.n5746 gnd.n1189 585
R11273 gnd.n5041 gnd.n1189 585
R11274 gnd.n5747 gnd.n1188 585
R11275 gnd.n1500 gnd.n1188 585
R11276 gnd.n4968 gnd.n1186 585
R11277 gnd.n4969 gnd.n4968 585
R11278 gnd.n5751 gnd.n1185 585
R11279 gnd.n5014 gnd.n1185 585
R11280 gnd.n5752 gnd.n1184 585
R11281 gnd.n1509 gnd.n1184 585
R11282 gnd.n5753 gnd.n1183 585
R11283 gnd.n5004 gnd.n1183 585
R11284 gnd.n4995 gnd.n1181 585
R11285 gnd.n4996 gnd.n4995 585
R11286 gnd.n5757 gnd.n1180 585
R11287 gnd.n4874 gnd.n1180 585
R11288 gnd.n5758 gnd.n1179 585
R11289 gnd.n4960 gnd.n1179 585
R11290 gnd.n5759 gnd.n1178 585
R11291 gnd.n1542 gnd.n1178 585
R11292 gnd.n4949 gnd.n1176 585
R11293 gnd.n4950 gnd.n4949 585
R11294 gnd.n5763 gnd.n1175 585
R11295 gnd.n4936 gnd.n1175 585
R11296 gnd.n5764 gnd.n1174 585
R11297 gnd.n4870 gnd.n1174 585
R11298 gnd.n5765 gnd.n1173 585
R11299 gnd.n4927 gnd.n1173 585
R11300 gnd.n1566 gnd.n1171 585
R11301 gnd.n1567 gnd.n1566 585
R11302 gnd.n5769 gnd.n1170 585
R11303 gnd.n4917 gnd.n1170 585
R11304 gnd.n5770 gnd.n1169 585
R11305 gnd.n1572 gnd.n1169 585
R11306 gnd.n5771 gnd.n1168 585
R11307 gnd.n1579 gnd.n1168 585
R11308 gnd.n1586 gnd.n1166 585
R11309 gnd.n4858 gnd.n1586 585
R11310 gnd.n5775 gnd.n1165 585
R11311 gnd.n1583 gnd.n1165 585
R11312 gnd.n5776 gnd.n1164 585
R11313 gnd.n4848 gnd.n1164 585
R11314 gnd.n5777 gnd.n1163 585
R11315 gnd.n4840 gnd.n1163 585
R11316 gnd.n1611 gnd.n1161 585
R11317 gnd.n1612 gnd.n1611 585
R11318 gnd.n5781 gnd.n1160 585
R11319 gnd.n4818 gnd.n1160 585
R11320 gnd.n5782 gnd.n1159 585
R11321 gnd.n1620 gnd.n1159 585
R11322 gnd.n5783 gnd.n1158 585
R11323 gnd.n4808 gnd.n1158 585
R11324 gnd.n4794 gnd.n1156 585
R11325 gnd.n4795 gnd.n4794 585
R11326 gnd.n5787 gnd.n1155 585
R11327 gnd.n1631 gnd.n1155 585
R11328 gnd.n5788 gnd.n1154 585
R11329 gnd.n4762 gnd.n1154 585
R11330 gnd.n5789 gnd.n1153 585
R11331 gnd.n1635 gnd.n1153 585
R11332 gnd.n4751 gnd.n1151 585
R11333 gnd.n4752 gnd.n4751 585
R11334 gnd.n5793 gnd.n1150 585
R11335 gnd.n1649 gnd.n1150 585
R11336 gnd.n5794 gnd.n1149 585
R11337 gnd.n4734 gnd.n1149 585
R11338 gnd.n5795 gnd.n1148 585
R11339 gnd.n1665 gnd.n1148 585
R11340 gnd.n4725 gnd.n1146 585
R11341 gnd.n4726 gnd.n4725 585
R11342 gnd.n5799 gnd.n1145 585
R11343 gnd.n1669 gnd.n1145 585
R11344 gnd.n5800 gnd.n1144 585
R11345 gnd.n1676 gnd.n1144 585
R11346 gnd.n5801 gnd.n1143 585
R11347 gnd.n4700 gnd.n1143 585
R11348 gnd.n1680 gnd.n1141 585
R11349 gnd.n1681 gnd.n1680 585
R11350 gnd.n5805 gnd.n1140 585
R11351 gnd.n4690 gnd.n1140 585
R11352 gnd.n5806 gnd.n1139 585
R11353 gnd.n4682 gnd.n1139 585
R11354 gnd.n5807 gnd.n1138 585
R11355 gnd.n1696 gnd.n1138 585
R11356 gnd.n1701 gnd.n1136 585
R11357 gnd.n1702 gnd.n1701 585
R11358 gnd.n5811 gnd.n1135 585
R11359 gnd.n4663 gnd.n1135 585
R11360 gnd.n5812 gnd.n1134 585
R11361 gnd.n4563 gnd.n1134 585
R11362 gnd.n5813 gnd.n1133 585
R11363 gnd.n4650 gnd.n1133 585
R11364 gnd.n1130 gnd.n1128 585
R11365 gnd.n4561 gnd.n1128 585
R11366 gnd.n5818 gnd.n5817 585
R11367 gnd.n5819 gnd.n5818 585
R11368 gnd.n1129 gnd.n1127 585
R11369 gnd.n4621 gnd.n1127 585
R11370 gnd.n4517 gnd.n1115 585
R11371 gnd.n5825 gnd.n1115 585
R11372 gnd.n4518 gnd.n4516 585
R11373 gnd.n4516 gnd.n1110 585
R11374 gnd.n4515 gnd.n4513 585
R11375 gnd.n4515 gnd.n1084 585
R11376 gnd.n4522 gnd.n4512 585
R11377 gnd.n4512 gnd.n1052 585
R11378 gnd.n4523 gnd.n4511 585
R11379 gnd.n4511 gnd.n4510 585
R11380 gnd.n4524 gnd.n1804 585
R11381 gnd.n4547 gnd.n1804 585
R11382 gnd.n1816 gnd.n1814 585
R11383 gnd.n1814 gnd.n1803 585
R11384 gnd.n4529 gnd.n4528 585
R11385 gnd.n4530 gnd.n4529 585
R11386 gnd.n1815 gnd.n1813 585
R11387 gnd.n1813 gnd.n1811 585
R11388 gnd.n4506 gnd.n4505 585
R11389 gnd.n4505 gnd.n4504 585
R11390 gnd.n1819 gnd.n1818 585
R11391 gnd.n1820 gnd.n1819 585
R11392 gnd.n4495 gnd.n4494 585
R11393 gnd.n4496 gnd.n4495 585
R11394 gnd.n1830 gnd.n1829 585
R11395 gnd.n1829 gnd.n1827 585
R11396 gnd.n4490 gnd.n4489 585
R11397 gnd.n4489 gnd.n4488 585
R11398 gnd.n1833 gnd.n1832 585
R11399 gnd.n1842 gnd.n1833 585
R11400 gnd.n4479 gnd.n4478 585
R11401 gnd.n4480 gnd.n4479 585
R11402 gnd.n5547 gnd.n5524 585
R11403 gnd.n5548 gnd.n5523 585
R11404 gnd.n5517 gnd.n5516 585
R11405 gnd.n5555 gnd.n5515 585
R11406 gnd.n5556 gnd.n5514 585
R11407 gnd.n5513 gnd.n5505 585
R11408 gnd.n5563 gnd.n5504 585
R11409 gnd.n5564 gnd.n5503 585
R11410 gnd.n5497 gnd.n5496 585
R11411 gnd.n5571 gnd.n5495 585
R11412 gnd.n5572 gnd.n5494 585
R11413 gnd.n5493 gnd.n5485 585
R11414 gnd.n5579 gnd.n5484 585
R11415 gnd.n5580 gnd.n5483 585
R11416 gnd.n5265 gnd.n5264 585
R11417 gnd.n5587 gnd.n5263 585
R11418 gnd.n5588 gnd.n5262 585
R11419 gnd.n5589 gnd.n5261 585
R11420 gnd.n5260 gnd.n5259 585
R11421 gnd.n5258 gnd.n5257 585
R11422 gnd.n5251 gnd.n1350 585
R11423 gnd.n5253 gnd.n5252 585
R11424 gnd.n5250 gnd.n5249 585
R11425 gnd.n5248 gnd.n5247 585
R11426 gnd.n1356 gnd.n1352 585
R11427 gnd.n5717 gnd.n5716 585
R11428 gnd.n5716 gnd.n5715 585
R11429 gnd.n1214 gnd.n1213 585
R11430 gnd.n5537 gnd.n5536 585
R11431 gnd.n5535 gnd.n5534 585
R11432 gnd.n5182 gnd.n1407 511.721
R11433 gnd.n5062 gnd.n1404 511.721
R11434 gnd.n1788 gnd.n1786 511.721
R11435 gnd.n5895 gnd.n1087 511.721
R11436 gnd.n1722 gnd.t282 389.64
R11437 gnd.n1455 gnd.t235 389.64
R11438 gnd.n5832 gnd.t199 389.64
R11439 gnd.n1449 gnd.t272 389.64
R11440 gnd.n1877 gnd.t262 371.625
R11441 gnd.n5541 gnd.t294 371.625
R11442 gnd.n306 gnd.t310 371.625
R11443 gnd.n286 gnd.t225 371.625
R11444 gnd.n7076 gnd.t269 371.625
R11445 gnd.n1300 gnd.t291 371.625
R11446 gnd.n1323 gnd.t285 371.625
R11447 gnd.n1345 gnd.t217 371.625
R11448 gnd.n6895 gnd.t256 371.625
R11449 gnd.n1848 gnd.t313 371.625
R11450 gnd.n3844 gnd.t297 371.625
R11451 gnd.n3783 gnd.t243 371.625
R11452 gnd.n3805 gnd.t232 371.625
R11453 gnd.n3826 gnd.t221 371.625
R11454 gnd.n1035 gnd.t307 371.625
R11455 gnd.n1956 gnd.t239 371.625
R11456 gnd.n1969 gnd.t259 371.625
R11457 gnd.n5525 gnd.t246 371.625
R11458 gnd.n6176 gnd.n711 345.092
R11459 gnd.n2745 gnd.t278 323.425
R11460 gnd.n2286 gnd.t300 323.425
R11461 gnd.n3593 gnd.n3567 289.615
R11462 gnd.n3561 gnd.n3535 289.615
R11463 gnd.n3529 gnd.n3503 289.615
R11464 gnd.n3498 gnd.n3472 289.615
R11465 gnd.n3466 gnd.n3440 289.615
R11466 gnd.n3434 gnd.n3408 289.615
R11467 gnd.n3402 gnd.n3376 289.615
R11468 gnd.n3371 gnd.n3345 289.615
R11469 gnd.n2819 gnd.t207 279.217
R11470 gnd.n2312 gnd.t203 279.217
R11471 gnd.n1094 gnd.t213 260.649
R11472 gnd.n1420 gnd.t255 260.649
R11473 gnd.n5897 gnd.n5896 256.663
R11474 gnd.n5897 gnd.n1053 256.663
R11475 gnd.n5897 gnd.n1054 256.663
R11476 gnd.n5897 gnd.n1055 256.663
R11477 gnd.n5897 gnd.n1056 256.663
R11478 gnd.n5897 gnd.n1057 256.663
R11479 gnd.n5897 gnd.n1058 256.663
R11480 gnd.n5897 gnd.n1059 256.663
R11481 gnd.n5897 gnd.n1060 256.663
R11482 gnd.n5897 gnd.n1061 256.663
R11483 gnd.n5897 gnd.n1062 256.663
R11484 gnd.n5897 gnd.n1063 256.663
R11485 gnd.n5897 gnd.n1064 256.663
R11486 gnd.n5897 gnd.n1065 256.663
R11487 gnd.n5897 gnd.n1066 256.663
R11488 gnd.n5897 gnd.n1067 256.663
R11489 gnd.n5900 gnd.n1050 256.663
R11490 gnd.n5898 gnd.n5897 256.663
R11491 gnd.n5897 gnd.n1068 256.663
R11492 gnd.n5897 gnd.n1069 256.663
R11493 gnd.n5897 gnd.n1070 256.663
R11494 gnd.n5897 gnd.n1071 256.663
R11495 gnd.n5897 gnd.n1072 256.663
R11496 gnd.n5897 gnd.n1073 256.663
R11497 gnd.n5897 gnd.n1074 256.663
R11498 gnd.n5897 gnd.n1075 256.663
R11499 gnd.n5897 gnd.n1076 256.663
R11500 gnd.n5897 gnd.n1077 256.663
R11501 gnd.n5897 gnd.n1078 256.663
R11502 gnd.n5897 gnd.n1079 256.663
R11503 gnd.n5897 gnd.n1080 256.663
R11504 gnd.n5897 gnd.n1081 256.663
R11505 gnd.n5897 gnd.n1082 256.663
R11506 gnd.n5897 gnd.n1083 256.663
R11507 gnd.n5061 gnd.n1394 256.663
R11508 gnd.n5067 gnd.n1394 256.663
R11509 gnd.n1476 gnd.n1394 256.663
R11510 gnd.n5074 gnd.n1394 256.663
R11511 gnd.n1473 gnd.n1394 256.663
R11512 gnd.n5081 gnd.n1394 256.663
R11513 gnd.n1470 gnd.n1394 256.663
R11514 gnd.n5088 gnd.n1394 256.663
R11515 gnd.n1467 gnd.n1394 256.663
R11516 gnd.n5095 gnd.n1394 256.663
R11517 gnd.n1464 gnd.n1394 256.663
R11518 gnd.n5102 gnd.n1394 256.663
R11519 gnd.n1461 gnd.n1394 256.663
R11520 gnd.n5109 gnd.n1394 256.663
R11521 gnd.n1458 gnd.n1394 256.663
R11522 gnd.n5117 gnd.n1394 256.663
R11523 gnd.n5120 gnd.n1310 256.663
R11524 gnd.n5121 gnd.n1394 256.663
R11525 gnd.n5125 gnd.n1394 256.663
R11526 gnd.n1452 gnd.n1394 256.663
R11527 gnd.n5133 gnd.n1394 256.663
R11528 gnd.n1447 gnd.n1394 256.663
R11529 gnd.n5140 gnd.n1394 256.663
R11530 gnd.n1444 gnd.n1394 256.663
R11531 gnd.n5147 gnd.n1394 256.663
R11532 gnd.n1441 gnd.n1394 256.663
R11533 gnd.n5154 gnd.n1394 256.663
R11534 gnd.n1438 gnd.n1394 256.663
R11535 gnd.n5161 gnd.n1394 256.663
R11536 gnd.n1435 gnd.n1394 256.663
R11537 gnd.n5168 gnd.n1394 256.663
R11538 gnd.n1432 gnd.n1394 256.663
R11539 gnd.n5175 gnd.n1394 256.663
R11540 gnd.n1429 gnd.n1394 256.663
R11541 gnd.n4039 gnd.n3753 242.672
R11542 gnd.n4039 gnd.n3754 242.672
R11543 gnd.n4039 gnd.n3755 242.672
R11544 gnd.n4039 gnd.n3756 242.672
R11545 gnd.n4039 gnd.n3757 242.672
R11546 gnd.n4039 gnd.n3758 242.672
R11547 gnd.n4039 gnd.n3759 242.672
R11548 gnd.n4039 gnd.n3760 242.672
R11549 gnd.n4039 gnd.n3761 242.672
R11550 gnd.n5951 gnd.n988 242.672
R11551 gnd.n5951 gnd.n987 242.672
R11552 gnd.n5951 gnd.n986 242.672
R11553 gnd.n5951 gnd.n985 242.672
R11554 gnd.n5951 gnd.n984 242.672
R11555 gnd.n5951 gnd.n983 242.672
R11556 gnd.n5951 gnd.n982 242.672
R11557 gnd.n5951 gnd.n981 242.672
R11558 gnd.n5951 gnd.n980 242.672
R11559 gnd.n2873 gnd.n2872 242.672
R11560 gnd.n2873 gnd.n2783 242.672
R11561 gnd.n2873 gnd.n2784 242.672
R11562 gnd.n2873 gnd.n2785 242.672
R11563 gnd.n2873 gnd.n2786 242.672
R11564 gnd.n2873 gnd.n2787 242.672
R11565 gnd.n2873 gnd.n2788 242.672
R11566 gnd.n2873 gnd.n2789 242.672
R11567 gnd.n2873 gnd.n2790 242.672
R11568 gnd.n2873 gnd.n2791 242.672
R11569 gnd.n2873 gnd.n2792 242.672
R11570 gnd.n2873 gnd.n2793 242.672
R11571 gnd.n2874 gnd.n2873 242.672
R11572 gnd.n3725 gnd.n2261 242.672
R11573 gnd.n3725 gnd.n2260 242.672
R11574 gnd.n3725 gnd.n2259 242.672
R11575 gnd.n3725 gnd.n2258 242.672
R11576 gnd.n3725 gnd.n2257 242.672
R11577 gnd.n3725 gnd.n2256 242.672
R11578 gnd.n3725 gnd.n2255 242.672
R11579 gnd.n3725 gnd.n2254 242.672
R11580 gnd.n3725 gnd.n2253 242.672
R11581 gnd.n3725 gnd.n2252 242.672
R11582 gnd.n3725 gnd.n2251 242.672
R11583 gnd.n3725 gnd.n2250 242.672
R11584 gnd.n3725 gnd.n2249 242.672
R11585 gnd.n5708 gnd.n1268 242.672
R11586 gnd.n5708 gnd.n1269 242.672
R11587 gnd.n5708 gnd.n1270 242.672
R11588 gnd.n5708 gnd.n1271 242.672
R11589 gnd.n5708 gnd.n1272 242.672
R11590 gnd.n5708 gnd.n1273 242.672
R11591 gnd.n5708 gnd.n1274 242.672
R11592 gnd.n5708 gnd.n1275 242.672
R11593 gnd.n5708 gnd.n1276 242.672
R11594 gnd.n7111 gnd.n220 242.672
R11595 gnd.n7111 gnd.n219 242.672
R11596 gnd.n7111 gnd.n218 242.672
R11597 gnd.n7111 gnd.n217 242.672
R11598 gnd.n7111 gnd.n216 242.672
R11599 gnd.n7111 gnd.n215 242.672
R11600 gnd.n7111 gnd.n214 242.672
R11601 gnd.n7111 gnd.n213 242.672
R11602 gnd.n7111 gnd.n212 242.672
R11603 gnd.n2957 gnd.n2956 242.672
R11604 gnd.n2956 gnd.n2695 242.672
R11605 gnd.n2956 gnd.n2696 242.672
R11606 gnd.n2956 gnd.n2697 242.672
R11607 gnd.n2956 gnd.n2698 242.672
R11608 gnd.n2956 gnd.n2699 242.672
R11609 gnd.n2956 gnd.n2700 242.672
R11610 gnd.n2956 gnd.n2701 242.672
R11611 gnd.n3725 gnd.n2262 242.672
R11612 gnd.n3725 gnd.n2263 242.672
R11613 gnd.n3725 gnd.n2264 242.672
R11614 gnd.n3725 gnd.n2265 242.672
R11615 gnd.n3725 gnd.n2266 242.672
R11616 gnd.n3725 gnd.n2267 242.672
R11617 gnd.n3725 gnd.n2268 242.672
R11618 gnd.n3725 gnd.n2269 242.672
R11619 gnd.n4039 gnd.n4038 242.672
R11620 gnd.n4039 gnd.n3726 242.672
R11621 gnd.n4039 gnd.n3727 242.672
R11622 gnd.n4039 gnd.n3728 242.672
R11623 gnd.n4039 gnd.n3729 242.672
R11624 gnd.n4039 gnd.n3730 242.672
R11625 gnd.n4039 gnd.n3731 242.672
R11626 gnd.n4039 gnd.n3732 242.672
R11627 gnd.n4039 gnd.n3733 242.672
R11628 gnd.n4039 gnd.n3734 242.672
R11629 gnd.n4039 gnd.n3735 242.672
R11630 gnd.n4039 gnd.n3736 242.672
R11631 gnd.n4039 gnd.n3737 242.672
R11632 gnd.n4039 gnd.n3738 242.672
R11633 gnd.n4039 gnd.n3739 242.672
R11634 gnd.n4039 gnd.n3740 242.672
R11635 gnd.n4039 gnd.n3741 242.672
R11636 gnd.n4039 gnd.n3742 242.672
R11637 gnd.n4039 gnd.n3743 242.672
R11638 gnd.n4039 gnd.n3744 242.672
R11639 gnd.n4039 gnd.n3745 242.672
R11640 gnd.n4039 gnd.n3746 242.672
R11641 gnd.n4039 gnd.n3747 242.672
R11642 gnd.n4039 gnd.n3748 242.672
R11643 gnd.n4039 gnd.n3749 242.672
R11644 gnd.n4039 gnd.n3750 242.672
R11645 gnd.n4039 gnd.n3751 242.672
R11646 gnd.n4039 gnd.n3752 242.672
R11647 gnd.n4040 gnd.n4039 242.672
R11648 gnd.n5951 gnd.n990 242.672
R11649 gnd.n5951 gnd.n991 242.672
R11650 gnd.n5951 gnd.n992 242.672
R11651 gnd.n5951 gnd.n993 242.672
R11652 gnd.n5951 gnd.n994 242.672
R11653 gnd.n5951 gnd.n995 242.672
R11654 gnd.n5951 gnd.n996 242.672
R11655 gnd.n5951 gnd.n997 242.672
R11656 gnd.n5951 gnd.n998 242.672
R11657 gnd.n5951 gnd.n999 242.672
R11658 gnd.n5951 gnd.n1000 242.672
R11659 gnd.n5951 gnd.n1001 242.672
R11660 gnd.n5951 gnd.n1002 242.672
R11661 gnd.n5951 gnd.n1003 242.672
R11662 gnd.n5951 gnd.n1004 242.672
R11663 gnd.n5951 gnd.n1005 242.672
R11664 gnd.n5901 gnd.n1046 242.672
R11665 gnd.n5951 gnd.n1006 242.672
R11666 gnd.n5951 gnd.n1007 242.672
R11667 gnd.n5951 gnd.n1008 242.672
R11668 gnd.n5951 gnd.n1009 242.672
R11669 gnd.n5951 gnd.n1010 242.672
R11670 gnd.n5951 gnd.n1011 242.672
R11671 gnd.n5951 gnd.n1012 242.672
R11672 gnd.n5951 gnd.n1013 242.672
R11673 gnd.n5951 gnd.n1014 242.672
R11674 gnd.n5951 gnd.n1015 242.672
R11675 gnd.n5951 gnd.n1016 242.672
R11676 gnd.n5951 gnd.n1017 242.672
R11677 gnd.n5951 gnd.n5950 242.672
R11678 gnd.n5708 gnd.n5707 242.672
R11679 gnd.n5708 gnd.n1240 242.672
R11680 gnd.n5708 gnd.n1241 242.672
R11681 gnd.n5708 gnd.n1242 242.672
R11682 gnd.n5708 gnd.n1243 242.672
R11683 gnd.n5708 gnd.n1244 242.672
R11684 gnd.n5708 gnd.n1245 242.672
R11685 gnd.n5708 gnd.n1246 242.672
R11686 gnd.n5708 gnd.n1247 242.672
R11687 gnd.n5708 gnd.n1248 242.672
R11688 gnd.n5708 gnd.n1249 242.672
R11689 gnd.n5708 gnd.n1250 242.672
R11690 gnd.n5708 gnd.n1251 242.672
R11691 gnd.n5655 gnd.n1311 242.672
R11692 gnd.n5708 gnd.n1252 242.672
R11693 gnd.n5708 gnd.n1253 242.672
R11694 gnd.n5708 gnd.n1254 242.672
R11695 gnd.n5708 gnd.n1255 242.672
R11696 gnd.n5708 gnd.n1256 242.672
R11697 gnd.n5708 gnd.n1257 242.672
R11698 gnd.n5708 gnd.n1258 242.672
R11699 gnd.n5708 gnd.n1259 242.672
R11700 gnd.n5708 gnd.n1260 242.672
R11701 gnd.n5708 gnd.n1261 242.672
R11702 gnd.n5708 gnd.n1262 242.672
R11703 gnd.n5708 gnd.n1263 242.672
R11704 gnd.n5708 gnd.n1264 242.672
R11705 gnd.n5708 gnd.n1265 242.672
R11706 gnd.n5708 gnd.n1266 242.672
R11707 gnd.n5708 gnd.n1267 242.672
R11708 gnd.n7111 gnd.n221 242.672
R11709 gnd.n7111 gnd.n222 242.672
R11710 gnd.n7111 gnd.n223 242.672
R11711 gnd.n7111 gnd.n224 242.672
R11712 gnd.n7111 gnd.n225 242.672
R11713 gnd.n7111 gnd.n226 242.672
R11714 gnd.n7111 gnd.n227 242.672
R11715 gnd.n7111 gnd.n228 242.672
R11716 gnd.n7111 gnd.n229 242.672
R11717 gnd.n7111 gnd.n230 242.672
R11718 gnd.n7111 gnd.n231 242.672
R11719 gnd.n7111 gnd.n232 242.672
R11720 gnd.n7111 gnd.n233 242.672
R11721 gnd.n7111 gnd.n234 242.672
R11722 gnd.n7111 gnd.n235 242.672
R11723 gnd.n7111 gnd.n236 242.672
R11724 gnd.n7111 gnd.n237 242.672
R11725 gnd.n7111 gnd.n238 242.672
R11726 gnd.n7111 gnd.n239 242.672
R11727 gnd.n7111 gnd.n240 242.672
R11728 gnd.n7111 gnd.n241 242.672
R11729 gnd.n7111 gnd.n242 242.672
R11730 gnd.n7111 gnd.n243 242.672
R11731 gnd.n7111 gnd.n244 242.672
R11732 gnd.n7111 gnd.n245 242.672
R11733 gnd.n7111 gnd.n246 242.672
R11734 gnd.n7111 gnd.n247 242.672
R11735 gnd.n7111 gnd.n248 242.672
R11736 gnd.n7111 gnd.n7110 242.672
R11737 gnd.n4459 gnd.n1864 242.672
R11738 gnd.n4459 gnd.n1865 242.672
R11739 gnd.n4459 gnd.n1866 242.672
R11740 gnd.n4459 gnd.n1867 242.672
R11741 gnd.n4459 gnd.n1868 242.672
R11742 gnd.n4459 gnd.n1869 242.672
R11743 gnd.n4459 gnd.n1870 242.672
R11744 gnd.n4459 gnd.n1871 242.672
R11745 gnd.n4459 gnd.n1872 242.672
R11746 gnd.n4459 gnd.n1873 242.672
R11747 gnd.n4459 gnd.n1874 242.672
R11748 gnd.n4459 gnd.n1875 242.672
R11749 gnd.n4459 gnd.n1876 242.672
R11750 gnd.n4459 gnd.n4458 242.672
R11751 gnd.n5715 gnd.n1229 242.672
R11752 gnd.n5715 gnd.n1228 242.672
R11753 gnd.n5715 gnd.n1227 242.672
R11754 gnd.n5715 gnd.n1226 242.672
R11755 gnd.n5715 gnd.n1225 242.672
R11756 gnd.n5715 gnd.n1224 242.672
R11757 gnd.n5715 gnd.n1223 242.672
R11758 gnd.n5715 gnd.n1222 242.672
R11759 gnd.n5715 gnd.n1221 242.672
R11760 gnd.n5715 gnd.n1220 242.672
R11761 gnd.n5715 gnd.n1219 242.672
R11762 gnd.n5715 gnd.n1218 242.672
R11763 gnd.n5715 gnd.n1217 242.672
R11764 gnd.n5715 gnd.n1230 242.672
R11765 gnd.n7112 gnd.n210 240.244
R11766 gnd.n7109 gnd.n249 240.244
R11767 gnd.n7105 gnd.n7104 240.244
R11768 gnd.n7101 gnd.n7100 240.244
R11769 gnd.n7097 gnd.n7096 240.244
R11770 gnd.n7093 gnd.n7092 240.244
R11771 gnd.n7089 gnd.n7088 240.244
R11772 gnd.n7085 gnd.n7084 240.244
R11773 gnd.n7081 gnd.n7080 240.244
R11774 gnd.n7074 gnd.n7073 240.244
R11775 gnd.n7070 gnd.n7069 240.244
R11776 gnd.n7066 gnd.n7065 240.244
R11777 gnd.n7062 gnd.n7061 240.244
R11778 gnd.n7058 gnd.n7057 240.244
R11779 gnd.n7054 gnd.n7053 240.244
R11780 gnd.n7050 gnd.n7049 240.244
R11781 gnd.n7046 gnd.n7045 240.244
R11782 gnd.n7042 gnd.n7041 240.244
R11783 gnd.n7038 gnd.n7037 240.244
R11784 gnd.n7031 gnd.n7030 240.244
R11785 gnd.n7028 gnd.n7027 240.244
R11786 gnd.n7024 gnd.n7023 240.244
R11787 gnd.n7020 gnd.n7019 240.244
R11788 gnd.n7016 gnd.n7015 240.244
R11789 gnd.n7012 gnd.n7011 240.244
R11790 gnd.n7008 gnd.n7007 240.244
R11791 gnd.n7004 gnd.n7003 240.244
R11792 gnd.n7000 gnd.n6999 240.244
R11793 gnd.n6996 gnd.n6995 240.244
R11794 gnd.n5356 gnd.n5272 240.244
R11795 gnd.n5357 gnd.n5356 240.244
R11796 gnd.n5357 gnd.n5287 240.244
R11797 gnd.n5381 gnd.n5287 240.244
R11798 gnd.n5381 gnd.n5306 240.244
R11799 gnd.n5385 gnd.n5306 240.244
R11800 gnd.n5385 gnd.n5317 240.244
R11801 gnd.n5409 gnd.n5317 240.244
R11802 gnd.n5409 gnd.n5328 240.244
R11803 gnd.n5343 gnd.n5328 240.244
R11804 gnd.n5343 gnd.n5335 240.244
R11805 gnd.n5416 gnd.n5335 240.244
R11806 gnd.n5416 gnd.n380 240.244
R11807 gnd.n6723 gnd.n380 240.244
R11808 gnd.n6723 gnd.n370 240.244
R11809 gnd.n370 gnd.n362 240.244
R11810 gnd.n6755 gnd.n362 240.244
R11811 gnd.n6755 gnd.n352 240.244
R11812 gnd.n6758 gnd.n352 240.244
R11813 gnd.n6758 gnd.n343 240.244
R11814 gnd.n343 gnd.n335 240.244
R11815 gnd.n6794 gnd.n335 240.244
R11816 gnd.n6794 gnd.n329 240.244
R11817 gnd.n6796 gnd.n329 240.244
R11818 gnd.n6796 gnd.n320 240.244
R11819 gnd.n320 gnd.n314 240.244
R11820 gnd.n6820 gnd.n314 240.244
R11821 gnd.n6820 gnd.n85 240.244
R11822 gnd.n6827 gnd.n85 240.244
R11823 gnd.n6827 gnd.n96 240.244
R11824 gnd.n6830 gnd.n96 240.244
R11825 gnd.n6830 gnd.n107 240.244
R11826 gnd.n6834 gnd.n107 240.244
R11827 gnd.n6834 gnd.n117 240.244
R11828 gnd.n6837 gnd.n117 240.244
R11829 gnd.n6837 gnd.n126 240.244
R11830 gnd.n6841 gnd.n126 240.244
R11831 gnd.n6841 gnd.n136 240.244
R11832 gnd.n6844 gnd.n136 240.244
R11833 gnd.n6844 gnd.n145 240.244
R11834 gnd.n6848 gnd.n145 240.244
R11835 gnd.n6848 gnd.n155 240.244
R11836 gnd.n6970 gnd.n155 240.244
R11837 gnd.n6970 gnd.n164 240.244
R11838 gnd.n6974 gnd.n164 240.244
R11839 gnd.n6974 gnd.n174 240.244
R11840 gnd.n6977 gnd.n174 240.244
R11841 gnd.n6977 gnd.n183 240.244
R11842 gnd.n6981 gnd.n183 240.244
R11843 gnd.n6981 gnd.n193 240.244
R11844 gnd.n6984 gnd.n193 240.244
R11845 gnd.n6984 gnd.n202 240.244
R11846 gnd.n6988 gnd.n202 240.244
R11847 gnd.n1280 gnd.n1279 240.244
R11848 gnd.n5701 gnd.n1279 240.244
R11849 gnd.n5699 gnd.n5698 240.244
R11850 gnd.n5695 gnd.n5694 240.244
R11851 gnd.n5691 gnd.n5690 240.244
R11852 gnd.n5687 gnd.n5686 240.244
R11853 gnd.n5683 gnd.n5682 240.244
R11854 gnd.n5679 gnd.n5678 240.244
R11855 gnd.n5675 gnd.n5674 240.244
R11856 gnd.n5670 gnd.n5669 240.244
R11857 gnd.n5666 gnd.n5665 240.244
R11858 gnd.n5662 gnd.n5661 240.244
R11859 gnd.n5658 gnd.n5657 240.244
R11860 gnd.n5653 gnd.n5652 240.244
R11861 gnd.n5649 gnd.n5648 240.244
R11862 gnd.n5645 gnd.n5644 240.244
R11863 gnd.n5641 gnd.n5640 240.244
R11864 gnd.n5637 gnd.n5636 240.244
R11865 gnd.n5633 gnd.n5632 240.244
R11866 gnd.n5629 gnd.n5628 240.244
R11867 gnd.n5625 gnd.n5624 240.244
R11868 gnd.n5621 gnd.n5620 240.244
R11869 gnd.n5617 gnd.n5616 240.244
R11870 gnd.n5613 gnd.n5612 240.244
R11871 gnd.n5609 gnd.n5608 240.244
R11872 gnd.n5605 gnd.n5604 240.244
R11873 gnd.n5601 gnd.n5600 240.244
R11874 gnd.n5597 gnd.n5596 240.244
R11875 gnd.n5296 gnd.n1281 240.244
R11876 gnd.n5296 gnd.n5291 240.244
R11877 gnd.n5466 gnd.n5291 240.244
R11878 gnd.n5466 gnd.n5292 240.244
R11879 gnd.n5462 gnd.n5292 240.244
R11880 gnd.n5462 gnd.n5304 240.244
R11881 gnd.n5454 gnd.n5304 240.244
R11882 gnd.n5454 gnd.n5320 240.244
R11883 gnd.n5450 gnd.n5320 240.244
R11884 gnd.n5450 gnd.n5326 240.244
R11885 gnd.n5442 gnd.n5326 240.244
R11886 gnd.n5442 gnd.n378 240.244
R11887 gnd.n6736 gnd.n378 240.244
R11888 gnd.n6736 gnd.n373 240.244
R11889 gnd.n6744 gnd.n373 240.244
R11890 gnd.n6744 gnd.n374 240.244
R11891 gnd.n374 gnd.n350 240.244
R11892 gnd.n6770 gnd.n350 240.244
R11893 gnd.n6770 gnd.n345 240.244
R11894 gnd.n6778 gnd.n345 240.244
R11895 gnd.n6778 gnd.n346 240.244
R11896 gnd.n346 gnd.n328 240.244
R11897 gnd.n6803 gnd.n328 240.244
R11898 gnd.n6803 gnd.n323 240.244
R11899 gnd.n6812 gnd.n323 240.244
R11900 gnd.n6812 gnd.n324 240.244
R11901 gnd.n324 gnd.n88 240.244
R11902 gnd.n7190 gnd.n88 240.244
R11903 gnd.n7190 gnd.n89 240.244
R11904 gnd.n7186 gnd.n89 240.244
R11905 gnd.n7186 gnd.n95 240.244
R11906 gnd.n7178 gnd.n95 240.244
R11907 gnd.n7178 gnd.n110 240.244
R11908 gnd.n7174 gnd.n110 240.244
R11909 gnd.n7174 gnd.n116 240.244
R11910 gnd.n7166 gnd.n116 240.244
R11911 gnd.n7166 gnd.n129 240.244
R11912 gnd.n7162 gnd.n129 240.244
R11913 gnd.n7162 gnd.n135 240.244
R11914 gnd.n7154 gnd.n135 240.244
R11915 gnd.n7154 gnd.n148 240.244
R11916 gnd.n7150 gnd.n148 240.244
R11917 gnd.n7150 gnd.n154 240.244
R11918 gnd.n7142 gnd.n154 240.244
R11919 gnd.n7142 gnd.n167 240.244
R11920 gnd.n7138 gnd.n167 240.244
R11921 gnd.n7138 gnd.n173 240.244
R11922 gnd.n7130 gnd.n173 240.244
R11923 gnd.n7130 gnd.n186 240.244
R11924 gnd.n7126 gnd.n186 240.244
R11925 gnd.n7126 gnd.n192 240.244
R11926 gnd.n7118 gnd.n192 240.244
R11927 gnd.n7118 gnd.n205 240.244
R11928 gnd.n5952 gnd.n977 240.244
R11929 gnd.n5949 gnd.n1018 240.244
R11930 gnd.n5945 gnd.n5944 240.244
R11931 gnd.n5941 gnd.n5940 240.244
R11932 gnd.n5937 gnd.n5936 240.244
R11933 gnd.n5933 gnd.n5932 240.244
R11934 gnd.n5929 gnd.n5928 240.244
R11935 gnd.n5925 gnd.n5924 240.244
R11936 gnd.n5921 gnd.n5920 240.244
R11937 gnd.n5916 gnd.n5915 240.244
R11938 gnd.n5912 gnd.n5911 240.244
R11939 gnd.n5908 gnd.n5907 240.244
R11940 gnd.n5904 gnd.n5903 240.244
R11941 gnd.n1978 gnd.n1977 240.244
R11942 gnd.n1981 gnd.n1980 240.244
R11943 gnd.n1988 gnd.n1987 240.244
R11944 gnd.n1991 gnd.n1990 240.244
R11945 gnd.n1996 gnd.n1971 240.244
R11946 gnd.n2000 gnd.n1999 240.244
R11947 gnd.n2007 gnd.n2006 240.244
R11948 gnd.n2010 gnd.n2009 240.244
R11949 gnd.n2017 gnd.n2016 240.244
R11950 gnd.n2020 gnd.n2019 240.244
R11951 gnd.n2027 gnd.n2026 240.244
R11952 gnd.n2030 gnd.n2029 240.244
R11953 gnd.n2037 gnd.n2036 240.244
R11954 gnd.n2040 gnd.n2039 240.244
R11955 gnd.n2045 gnd.n1958 240.244
R11956 gnd.n4042 gnd.n2238 240.244
R11957 gnd.n2238 gnd.n2228 240.244
R11958 gnd.n4061 gnd.n2228 240.244
R11959 gnd.n4062 gnd.n4061 240.244
R11960 gnd.n4062 gnd.n2219 240.244
R11961 gnd.n2219 gnd.n2210 240.244
R11962 gnd.n4081 gnd.n2210 240.244
R11963 gnd.n4082 gnd.n4081 240.244
R11964 gnd.n4082 gnd.n2202 240.244
R11965 gnd.n2202 gnd.n2192 240.244
R11966 gnd.n4101 gnd.n2192 240.244
R11967 gnd.n4102 gnd.n4101 240.244
R11968 gnd.n4102 gnd.n2182 240.244
R11969 gnd.n4105 gnd.n2182 240.244
R11970 gnd.n4105 gnd.n2173 240.244
R11971 gnd.n2173 gnd.n2166 240.244
R11972 gnd.n4137 gnd.n2166 240.244
R11973 gnd.n4137 gnd.n2156 240.244
R11974 gnd.n4140 gnd.n2156 240.244
R11975 gnd.n4140 gnd.n2148 240.244
R11976 gnd.n2148 gnd.n2141 240.244
R11977 gnd.n4172 gnd.n2141 240.244
R11978 gnd.n4172 gnd.n2132 240.244
R11979 gnd.n4175 gnd.n2132 240.244
R11980 gnd.n4175 gnd.n2124 240.244
R11981 gnd.n2124 gnd.n2115 240.244
R11982 gnd.n4219 gnd.n2115 240.244
R11983 gnd.n4219 gnd.n2107 240.244
R11984 gnd.n2107 gnd.n2098 240.244
R11985 gnd.n4238 gnd.n2098 240.244
R11986 gnd.n4239 gnd.n4238 240.244
R11987 gnd.n4239 gnd.n2087 240.244
R11988 gnd.n4242 gnd.n2087 240.244
R11989 gnd.n4242 gnd.n2079 240.244
R11990 gnd.n4245 gnd.n2079 240.244
R11991 gnd.n4245 gnd.n884 240.244
R11992 gnd.n4275 gnd.n884 240.244
R11993 gnd.n4275 gnd.n897 240.244
R11994 gnd.n2068 gnd.n897 240.244
R11995 gnd.n2068 gnd.n908 240.244
R11996 gnd.n4282 gnd.n908 240.244
R11997 gnd.n4282 gnd.n919 240.244
R11998 gnd.n4341 gnd.n919 240.244
R11999 gnd.n4341 gnd.n928 240.244
R12000 gnd.n4346 gnd.n928 240.244
R12001 gnd.n4346 gnd.n939 240.244
R12002 gnd.n4356 gnd.n939 240.244
R12003 gnd.n4356 gnd.n948 240.244
R12004 gnd.n4361 gnd.n948 240.244
R12005 gnd.n4361 gnd.n959 240.244
R12006 gnd.n4373 gnd.n959 240.244
R12007 gnd.n4373 gnd.n969 240.244
R12008 gnd.n1852 gnd.n969 240.244
R12009 gnd.n3764 gnd.n3763 240.244
R12010 gnd.n4032 gnd.n3763 240.244
R12011 gnd.n4030 gnd.n4029 240.244
R12012 gnd.n4026 gnd.n4025 240.244
R12013 gnd.n4022 gnd.n4021 240.244
R12014 gnd.n4018 gnd.n4017 240.244
R12015 gnd.n4014 gnd.n4013 240.244
R12016 gnd.n4010 gnd.n4009 240.244
R12017 gnd.n4006 gnd.n4005 240.244
R12018 gnd.n4001 gnd.n4000 240.244
R12019 gnd.n3997 gnd.n3996 240.244
R12020 gnd.n3993 gnd.n3992 240.244
R12021 gnd.n3989 gnd.n3988 240.244
R12022 gnd.n3985 gnd.n3984 240.244
R12023 gnd.n3981 gnd.n3980 240.244
R12024 gnd.n3977 gnd.n3976 240.244
R12025 gnd.n3973 gnd.n3972 240.244
R12026 gnd.n3969 gnd.n3968 240.244
R12027 gnd.n3965 gnd.n3964 240.244
R12028 gnd.n3961 gnd.n3960 240.244
R12029 gnd.n3957 gnd.n3956 240.244
R12030 gnd.n3953 gnd.n3952 240.244
R12031 gnd.n3949 gnd.n3948 240.244
R12032 gnd.n3945 gnd.n3944 240.244
R12033 gnd.n3941 gnd.n3940 240.244
R12034 gnd.n3937 gnd.n3936 240.244
R12035 gnd.n3933 gnd.n3932 240.244
R12036 gnd.n3929 gnd.n3928 240.244
R12037 gnd.n3925 gnd.n2246 240.244
R12038 gnd.n4053 gnd.n2236 240.244
R12039 gnd.n4053 gnd.n2232 240.244
R12040 gnd.n4059 gnd.n2232 240.244
R12041 gnd.n4059 gnd.n2217 240.244
R12042 gnd.n4073 gnd.n2217 240.244
R12043 gnd.n4073 gnd.n2213 240.244
R12044 gnd.n4079 gnd.n2213 240.244
R12045 gnd.n4079 gnd.n2200 240.244
R12046 gnd.n4093 gnd.n2200 240.244
R12047 gnd.n4093 gnd.n2196 240.244
R12048 gnd.n4099 gnd.n2196 240.244
R12049 gnd.n4099 gnd.n2180 240.244
R12050 gnd.n4117 gnd.n2180 240.244
R12051 gnd.n4117 gnd.n2175 240.244
R12052 gnd.n4125 gnd.n2175 240.244
R12053 gnd.n4125 gnd.n2176 240.244
R12054 gnd.n2176 gnd.n2155 240.244
R12055 gnd.n4152 gnd.n2155 240.244
R12056 gnd.n4152 gnd.n2150 240.244
R12057 gnd.n4160 gnd.n2150 240.244
R12058 gnd.n4160 gnd.n2151 240.244
R12059 gnd.n2151 gnd.n2131 240.244
R12060 gnd.n4187 gnd.n2131 240.244
R12061 gnd.n4187 gnd.n2126 240.244
R12062 gnd.n4195 gnd.n2126 240.244
R12063 gnd.n4195 gnd.n2127 240.244
R12064 gnd.n2127 gnd.n2106 240.244
R12065 gnd.n4230 gnd.n2106 240.244
R12066 gnd.n4230 gnd.n2102 240.244
R12067 gnd.n4236 gnd.n2102 240.244
R12068 gnd.n4236 gnd.n2085 240.244
R12069 gnd.n4257 gnd.n2085 240.244
R12070 gnd.n4257 gnd.n2081 240.244
R12071 gnd.n4264 gnd.n2081 240.244
R12072 gnd.n4264 gnd.n888 240.244
R12073 gnd.n6006 gnd.n888 240.244
R12074 gnd.n6006 gnd.n889 240.244
R12075 gnd.n6002 gnd.n889 240.244
R12076 gnd.n6002 gnd.n895 240.244
R12077 gnd.n5994 gnd.n895 240.244
R12078 gnd.n5994 gnd.n911 240.244
R12079 gnd.n5990 gnd.n911 240.244
R12080 gnd.n5990 gnd.n917 240.244
R12081 gnd.n5982 gnd.n917 240.244
R12082 gnd.n5982 gnd.n931 240.244
R12083 gnd.n5978 gnd.n931 240.244
R12084 gnd.n5978 gnd.n937 240.244
R12085 gnd.n5970 gnd.n937 240.244
R12086 gnd.n5970 gnd.n951 240.244
R12087 gnd.n5966 gnd.n951 240.244
R12088 gnd.n5966 gnd.n957 240.244
R12089 gnd.n5958 gnd.n957 240.244
R12090 gnd.n5958 gnd.n972 240.244
R12091 gnd.n3724 gnd.n2271 240.244
R12092 gnd.n3717 gnd.n3716 240.244
R12093 gnd.n3714 gnd.n3713 240.244
R12094 gnd.n3710 gnd.n3709 240.244
R12095 gnd.n3706 gnd.n3705 240.244
R12096 gnd.n3702 gnd.n3701 240.244
R12097 gnd.n3698 gnd.n3697 240.244
R12098 gnd.n3694 gnd.n3693 240.244
R12099 gnd.n2968 gnd.n2680 240.244
R12100 gnd.n2978 gnd.n2680 240.244
R12101 gnd.n2978 gnd.n2671 240.244
R12102 gnd.n2671 gnd.n2660 240.244
R12103 gnd.n2999 gnd.n2660 240.244
R12104 gnd.n2999 gnd.n2654 240.244
R12105 gnd.n3009 gnd.n2654 240.244
R12106 gnd.n3009 gnd.n2643 240.244
R12107 gnd.n2643 gnd.n2635 240.244
R12108 gnd.n3027 gnd.n2635 240.244
R12109 gnd.n3028 gnd.n3027 240.244
R12110 gnd.n3028 gnd.n2620 240.244
R12111 gnd.n3030 gnd.n2620 240.244
R12112 gnd.n3030 gnd.n2606 240.244
R12113 gnd.n3072 gnd.n2606 240.244
R12114 gnd.n3073 gnd.n3072 240.244
R12115 gnd.n3076 gnd.n3073 240.244
R12116 gnd.n3076 gnd.n2561 240.244
R12117 gnd.n2601 gnd.n2561 240.244
R12118 gnd.n2601 gnd.n2571 240.244
R12119 gnd.n3086 gnd.n2571 240.244
R12120 gnd.n3086 gnd.n2592 240.244
R12121 gnd.n3096 gnd.n2592 240.244
R12122 gnd.n3096 gnd.n2474 240.244
R12123 gnd.n3141 gnd.n2474 240.244
R12124 gnd.n3141 gnd.n2460 240.244
R12125 gnd.n3163 gnd.n2460 240.244
R12126 gnd.n3164 gnd.n3163 240.244
R12127 gnd.n3164 gnd.n2447 240.244
R12128 gnd.n2447 gnd.n2436 240.244
R12129 gnd.n3195 gnd.n2436 240.244
R12130 gnd.n3196 gnd.n3195 240.244
R12131 gnd.n3197 gnd.n3196 240.244
R12132 gnd.n3197 gnd.n2421 240.244
R12133 gnd.n2421 gnd.n2420 240.244
R12134 gnd.n2420 gnd.n2405 240.244
R12135 gnd.n3248 gnd.n2405 240.244
R12136 gnd.n3249 gnd.n3248 240.244
R12137 gnd.n3249 gnd.n2392 240.244
R12138 gnd.n2392 gnd.n2381 240.244
R12139 gnd.n3280 gnd.n2381 240.244
R12140 gnd.n3281 gnd.n3280 240.244
R12141 gnd.n3282 gnd.n3281 240.244
R12142 gnd.n3282 gnd.n2365 240.244
R12143 gnd.n2365 gnd.n2364 240.244
R12144 gnd.n2364 gnd.n2351 240.244
R12145 gnd.n3337 gnd.n2351 240.244
R12146 gnd.n3338 gnd.n3337 240.244
R12147 gnd.n3338 gnd.n2338 240.244
R12148 gnd.n2338 gnd.n2328 240.244
R12149 gnd.n3625 gnd.n2328 240.244
R12150 gnd.n3628 gnd.n3625 240.244
R12151 gnd.n3628 gnd.n3627 240.244
R12152 gnd.n2958 gnd.n2693 240.244
R12153 gnd.n2714 gnd.n2693 240.244
R12154 gnd.n2717 gnd.n2716 240.244
R12155 gnd.n2724 gnd.n2723 240.244
R12156 gnd.n2727 gnd.n2726 240.244
R12157 gnd.n2734 gnd.n2733 240.244
R12158 gnd.n2737 gnd.n2736 240.244
R12159 gnd.n2744 gnd.n2743 240.244
R12160 gnd.n2966 gnd.n2690 240.244
R12161 gnd.n2690 gnd.n2669 240.244
R12162 gnd.n2989 gnd.n2669 240.244
R12163 gnd.n2989 gnd.n2663 240.244
R12164 gnd.n2997 gnd.n2663 240.244
R12165 gnd.n2997 gnd.n2665 240.244
R12166 gnd.n2665 gnd.n2641 240.244
R12167 gnd.n3019 gnd.n2641 240.244
R12168 gnd.n3019 gnd.n2637 240.244
R12169 gnd.n3025 gnd.n2637 240.244
R12170 gnd.n3025 gnd.n2619 240.244
R12171 gnd.n3050 gnd.n2619 240.244
R12172 gnd.n3050 gnd.n2614 240.244
R12173 gnd.n3062 gnd.n2614 240.244
R12174 gnd.n3062 gnd.n2615 240.244
R12175 gnd.n3058 gnd.n2615 240.244
R12176 gnd.n3058 gnd.n2563 240.244
R12177 gnd.n3110 gnd.n2563 240.244
R12178 gnd.n3110 gnd.n2564 240.244
R12179 gnd.n3106 gnd.n2564 240.244
R12180 gnd.n3106 gnd.n2570 240.244
R12181 gnd.n2590 gnd.n2570 240.244
R12182 gnd.n2590 gnd.n2472 240.244
R12183 gnd.n3145 gnd.n2472 240.244
R12184 gnd.n3145 gnd.n2467 240.244
R12185 gnd.n3153 gnd.n2467 240.244
R12186 gnd.n3153 gnd.n2468 240.244
R12187 gnd.n2468 gnd.n2445 240.244
R12188 gnd.n3185 gnd.n2445 240.244
R12189 gnd.n3185 gnd.n2440 240.244
R12190 gnd.n3193 gnd.n2440 240.244
R12191 gnd.n3193 gnd.n2441 240.244
R12192 gnd.n2441 gnd.n2418 240.244
R12193 gnd.n3230 gnd.n2418 240.244
R12194 gnd.n3230 gnd.n2413 240.244
R12195 gnd.n3238 gnd.n2413 240.244
R12196 gnd.n3238 gnd.n2414 240.244
R12197 gnd.n2414 gnd.n2390 240.244
R12198 gnd.n3270 gnd.n2390 240.244
R12199 gnd.n3270 gnd.n2385 240.244
R12200 gnd.n3278 gnd.n2385 240.244
R12201 gnd.n3278 gnd.n2386 240.244
R12202 gnd.n2386 gnd.n2363 240.244
R12203 gnd.n3319 gnd.n2363 240.244
R12204 gnd.n3319 gnd.n2358 240.244
R12205 gnd.n3327 gnd.n2358 240.244
R12206 gnd.n3327 gnd.n2359 240.244
R12207 gnd.n2359 gnd.n2336 240.244
R12208 gnd.n3613 gnd.n2336 240.244
R12209 gnd.n3613 gnd.n2331 240.244
R12210 gnd.n3623 gnd.n2331 240.244
R12211 gnd.n3623 gnd.n2332 240.244
R12212 gnd.n2332 gnd.n2270 240.244
R12213 gnd.n6906 gnd.n211 240.244
R12214 gnd.n6912 gnd.n6911 240.244
R12215 gnd.n6915 gnd.n6914 240.244
R12216 gnd.n6922 gnd.n6921 240.244
R12217 gnd.n6925 gnd.n6924 240.244
R12218 gnd.n6932 gnd.n6931 240.244
R12219 gnd.n6935 gnd.n6934 240.244
R12220 gnd.n6942 gnd.n6941 240.244
R12221 gnd.n6945 gnd.n6944 240.244
R12222 gnd.n5372 gnd.n5273 240.244
R12223 gnd.n5373 gnd.n5372 240.244
R12224 gnd.n5373 gnd.n5288 240.244
R12225 gnd.n5379 gnd.n5288 240.244
R12226 gnd.n5379 gnd.n5307 240.244
R12227 gnd.n5401 gnd.n5307 240.244
R12228 gnd.n5401 gnd.n5318 240.244
R12229 gnd.n5407 gnd.n5318 240.244
R12230 gnd.n5407 gnd.n5329 240.244
R12231 gnd.n5425 gnd.n5329 240.244
R12232 gnd.n5425 gnd.n5336 240.244
R12233 gnd.n5418 gnd.n5336 240.244
R12234 gnd.n5418 gnd.n381 240.244
R12235 gnd.n381 gnd.n369 240.244
R12236 gnd.n6746 gnd.n369 240.244
R12237 gnd.n6746 gnd.n364 240.244
R12238 gnd.n6753 gnd.n364 240.244
R12239 gnd.n6753 gnd.n353 240.244
R12240 gnd.n353 gnd.n342 240.244
R12241 gnd.n6780 gnd.n342 240.244
R12242 gnd.n6780 gnd.n337 240.244
R12243 gnd.n6792 gnd.n337 240.244
R12244 gnd.n6792 gnd.n330 240.244
R12245 gnd.n6785 gnd.n330 240.244
R12246 gnd.n6785 gnd.n322 240.244
R12247 gnd.n322 gnd.n321 240.244
R12248 gnd.n321 gnd.n82 240.244
R12249 gnd.n7192 gnd.n82 240.244
R12250 gnd.n7192 gnd.n84 240.244
R12251 gnd.n97 gnd.n84 240.244
R12252 gnd.n6861 gnd.n97 240.244
R12253 gnd.n6861 gnd.n108 240.244
R12254 gnd.n6864 gnd.n108 240.244
R12255 gnd.n6864 gnd.n118 240.244
R12256 gnd.n6869 gnd.n118 240.244
R12257 gnd.n6869 gnd.n127 240.244
R12258 gnd.n6872 gnd.n127 240.244
R12259 gnd.n6872 gnd.n137 240.244
R12260 gnd.n6877 gnd.n137 240.244
R12261 gnd.n6877 gnd.n146 240.244
R12262 gnd.n6880 gnd.n146 240.244
R12263 gnd.n6880 gnd.n156 240.244
R12264 gnd.n6968 gnd.n156 240.244
R12265 gnd.n6968 gnd.n165 240.244
R12266 gnd.n6964 gnd.n165 240.244
R12267 gnd.n6964 gnd.n175 240.244
R12268 gnd.n6961 gnd.n175 240.244
R12269 gnd.n6961 gnd.n184 240.244
R12270 gnd.n6958 gnd.n184 240.244
R12271 gnd.n6958 gnd.n194 240.244
R12272 gnd.n6955 gnd.n194 240.244
R12273 gnd.n6955 gnd.n203 240.244
R12274 gnd.n6952 gnd.n203 240.244
R12275 gnd.n5480 gnd.n5479 240.244
R12276 gnd.n5488 gnd.n5487 240.244
R12277 gnd.n5490 gnd.n5489 240.244
R12278 gnd.n5500 gnd.n5499 240.244
R12279 gnd.n5508 gnd.n5507 240.244
R12280 gnd.n5510 gnd.n5509 240.244
R12281 gnd.n5520 gnd.n5519 240.244
R12282 gnd.n5530 gnd.n5529 240.244
R12283 gnd.n5540 gnd.n1277 240.244
R12284 gnd.n5476 gnd.n5268 240.244
R12285 gnd.n5362 gnd.n5268 240.244
R12286 gnd.n5362 gnd.n5290 240.244
R12287 gnd.n5309 gnd.n5290 240.244
R12288 gnd.n5460 gnd.n5309 240.244
R12289 gnd.n5460 gnd.n5310 240.244
R12290 gnd.n5456 gnd.n5310 240.244
R12291 gnd.n5456 gnd.n5316 240.244
R12292 gnd.n5448 gnd.n5316 240.244
R12293 gnd.n5448 gnd.n5330 240.244
R12294 gnd.n5444 gnd.n5330 240.244
R12295 gnd.n5444 gnd.n383 240.244
R12296 gnd.n6734 gnd.n383 240.244
R12297 gnd.n6734 gnd.n384 240.244
R12298 gnd.n384 gnd.n372 240.244
R12299 gnd.n6729 gnd.n372 240.244
R12300 gnd.n6729 gnd.n355 240.244
R12301 gnd.n6768 gnd.n355 240.244
R12302 gnd.n6768 gnd.n356 240.244
R12303 gnd.n356 gnd.n344 240.244
R12304 gnd.n6763 gnd.n344 240.244
R12305 gnd.n6763 gnd.n331 240.244
R12306 gnd.n6801 gnd.n331 240.244
R12307 gnd.n6801 gnd.n318 240.244
R12308 gnd.n6814 gnd.n318 240.244
R12309 gnd.n6814 gnd.n312 240.244
R12310 gnd.n6822 gnd.n312 240.244
R12311 gnd.n6822 gnd.n87 240.244
R12312 gnd.n98 gnd.n87 240.244
R12313 gnd.n7184 gnd.n98 240.244
R12314 gnd.n7184 gnd.n99 240.244
R12315 gnd.n7180 gnd.n99 240.244
R12316 gnd.n7180 gnd.n105 240.244
R12317 gnd.n7172 gnd.n105 240.244
R12318 gnd.n7172 gnd.n120 240.244
R12319 gnd.n7168 gnd.n120 240.244
R12320 gnd.n7168 gnd.n125 240.244
R12321 gnd.n7160 gnd.n125 240.244
R12322 gnd.n7160 gnd.n138 240.244
R12323 gnd.n7156 gnd.n138 240.244
R12324 gnd.n7156 gnd.n143 240.244
R12325 gnd.n7148 gnd.n143 240.244
R12326 gnd.n7148 gnd.n158 240.244
R12327 gnd.n7144 gnd.n158 240.244
R12328 gnd.n7144 gnd.n163 240.244
R12329 gnd.n7136 gnd.n163 240.244
R12330 gnd.n7136 gnd.n176 240.244
R12331 gnd.n7132 gnd.n176 240.244
R12332 gnd.n7132 gnd.n181 240.244
R12333 gnd.n7124 gnd.n181 240.244
R12334 gnd.n7124 gnd.n196 240.244
R12335 gnd.n7120 gnd.n196 240.244
R12336 gnd.n7120 gnd.n201 240.244
R12337 gnd.n2290 gnd.n2248 240.244
R12338 gnd.n3684 gnd.n3683 240.244
R12339 gnd.n3680 gnd.n3679 240.244
R12340 gnd.n3676 gnd.n3675 240.244
R12341 gnd.n3672 gnd.n3671 240.244
R12342 gnd.n3668 gnd.n3667 240.244
R12343 gnd.n3664 gnd.n3663 240.244
R12344 gnd.n3660 gnd.n3659 240.244
R12345 gnd.n3656 gnd.n3655 240.244
R12346 gnd.n3652 gnd.n3651 240.244
R12347 gnd.n3648 gnd.n3647 240.244
R12348 gnd.n3644 gnd.n3643 240.244
R12349 gnd.n3640 gnd.n3639 240.244
R12350 gnd.n2881 gnd.n2778 240.244
R12351 gnd.n2881 gnd.n2771 240.244
R12352 gnd.n2892 gnd.n2771 240.244
R12353 gnd.n2892 gnd.n2767 240.244
R12354 gnd.n2898 gnd.n2767 240.244
R12355 gnd.n2898 gnd.n2759 240.244
R12356 gnd.n2908 gnd.n2759 240.244
R12357 gnd.n2908 gnd.n2754 240.244
R12358 gnd.n2944 gnd.n2754 240.244
R12359 gnd.n2944 gnd.n2755 240.244
R12360 gnd.n2755 gnd.n2702 240.244
R12361 gnd.n2939 gnd.n2702 240.244
R12362 gnd.n2939 gnd.n2938 240.244
R12363 gnd.n2938 gnd.n2681 240.244
R12364 gnd.n2934 gnd.n2681 240.244
R12365 gnd.n2934 gnd.n2672 240.244
R12366 gnd.n2931 gnd.n2672 240.244
R12367 gnd.n2931 gnd.n2930 240.244
R12368 gnd.n2930 gnd.n2655 240.244
R12369 gnd.n2926 gnd.n2655 240.244
R12370 gnd.n2926 gnd.n2644 240.244
R12371 gnd.n2644 gnd.n2625 240.244
R12372 gnd.n3039 gnd.n2625 240.244
R12373 gnd.n3039 gnd.n2621 240.244
R12374 gnd.n3047 gnd.n2621 240.244
R12375 gnd.n3047 gnd.n2612 240.244
R12376 gnd.n2612 gnd.n2548 240.244
R12377 gnd.n3119 gnd.n2548 240.244
R12378 gnd.n3119 gnd.n2549 240.244
R12379 gnd.n2560 gnd.n2549 240.244
R12380 gnd.n2595 gnd.n2560 240.244
R12381 gnd.n2598 gnd.n2595 240.244
R12382 gnd.n2598 gnd.n2572 240.244
R12383 gnd.n2585 gnd.n2572 240.244
R12384 gnd.n2585 gnd.n2582 240.244
R12385 gnd.n2582 gnd.n2475 240.244
R12386 gnd.n3140 gnd.n2475 240.244
R12387 gnd.n3140 gnd.n2465 240.244
R12388 gnd.n3136 gnd.n2465 240.244
R12389 gnd.n3136 gnd.n2459 240.244
R12390 gnd.n3133 gnd.n2459 240.244
R12391 gnd.n3133 gnd.n2448 240.244
R12392 gnd.n3130 gnd.n2448 240.244
R12393 gnd.n3130 gnd.n2426 240.244
R12394 gnd.n3206 gnd.n2426 240.244
R12395 gnd.n3206 gnd.n2422 240.244
R12396 gnd.n3227 gnd.n2422 240.244
R12397 gnd.n3227 gnd.n2411 240.244
R12398 gnd.n3223 gnd.n2411 240.244
R12399 gnd.n3223 gnd.n2404 240.244
R12400 gnd.n3220 gnd.n2404 240.244
R12401 gnd.n3220 gnd.n2393 240.244
R12402 gnd.n3217 gnd.n2393 240.244
R12403 gnd.n3217 gnd.n2370 240.244
R12404 gnd.n3291 gnd.n2370 240.244
R12405 gnd.n3291 gnd.n2366 240.244
R12406 gnd.n3316 gnd.n2366 240.244
R12407 gnd.n3316 gnd.n2357 240.244
R12408 gnd.n3312 gnd.n2357 240.244
R12409 gnd.n3312 gnd.n2350 240.244
R12410 gnd.n3308 gnd.n2350 240.244
R12411 gnd.n3308 gnd.n2339 240.244
R12412 gnd.n3305 gnd.n2339 240.244
R12413 gnd.n3305 gnd.n2319 240.244
R12414 gnd.n3635 gnd.n2319 240.244
R12415 gnd.n2795 gnd.n2794 240.244
R12416 gnd.n2866 gnd.n2794 240.244
R12417 gnd.n2864 gnd.n2863 240.244
R12418 gnd.n2860 gnd.n2859 240.244
R12419 gnd.n2856 gnd.n2855 240.244
R12420 gnd.n2852 gnd.n2851 240.244
R12421 gnd.n2848 gnd.n2847 240.244
R12422 gnd.n2844 gnd.n2843 240.244
R12423 gnd.n2840 gnd.n2839 240.244
R12424 gnd.n2836 gnd.n2835 240.244
R12425 gnd.n2832 gnd.n2831 240.244
R12426 gnd.n2828 gnd.n2827 240.244
R12427 gnd.n2824 gnd.n2782 240.244
R12428 gnd.n2884 gnd.n2776 240.244
R12429 gnd.n2884 gnd.n2772 240.244
R12430 gnd.n2890 gnd.n2772 240.244
R12431 gnd.n2890 gnd.n2765 240.244
R12432 gnd.n2900 gnd.n2765 240.244
R12433 gnd.n2900 gnd.n2761 240.244
R12434 gnd.n2906 gnd.n2761 240.244
R12435 gnd.n2906 gnd.n2752 240.244
R12436 gnd.n2946 gnd.n2752 240.244
R12437 gnd.n2946 gnd.n2703 240.244
R12438 gnd.n2954 gnd.n2703 240.244
R12439 gnd.n2954 gnd.n2704 240.244
R12440 gnd.n2704 gnd.n2682 240.244
R12441 gnd.n2975 gnd.n2682 240.244
R12442 gnd.n2975 gnd.n2674 240.244
R12443 gnd.n2986 gnd.n2674 240.244
R12444 gnd.n2986 gnd.n2675 240.244
R12445 gnd.n2675 gnd.n2656 240.244
R12446 gnd.n3006 gnd.n2656 240.244
R12447 gnd.n3006 gnd.n2646 240.244
R12448 gnd.n3016 gnd.n2646 240.244
R12449 gnd.n3016 gnd.n2627 240.244
R12450 gnd.n3037 gnd.n2627 240.244
R12451 gnd.n3037 gnd.n2629 240.244
R12452 gnd.n2629 gnd.n2610 240.244
R12453 gnd.n3065 gnd.n2610 240.244
R12454 gnd.n3065 gnd.n2552 240.244
R12455 gnd.n3117 gnd.n2552 240.244
R12456 gnd.n3117 gnd.n2553 240.244
R12457 gnd.n3113 gnd.n2553 240.244
R12458 gnd.n3113 gnd.n2559 240.244
R12459 gnd.n2574 gnd.n2559 240.244
R12460 gnd.n3103 gnd.n2574 240.244
R12461 gnd.n3103 gnd.n2575 240.244
R12462 gnd.n3099 gnd.n2575 240.244
R12463 gnd.n3099 gnd.n2581 240.244
R12464 gnd.n2581 gnd.n2464 240.244
R12465 gnd.n3156 gnd.n2464 240.244
R12466 gnd.n3156 gnd.n2457 240.244
R12467 gnd.n3167 gnd.n2457 240.244
R12468 gnd.n3167 gnd.n2450 240.244
R12469 gnd.n3182 gnd.n2450 240.244
R12470 gnd.n3182 gnd.n2451 240.244
R12471 gnd.n2451 gnd.n2429 240.244
R12472 gnd.n3204 gnd.n2429 240.244
R12473 gnd.n3204 gnd.n2430 240.244
R12474 gnd.n2430 gnd.n2409 240.244
R12475 gnd.n3241 gnd.n2409 240.244
R12476 gnd.n3241 gnd.n2402 240.244
R12477 gnd.n3252 gnd.n2402 240.244
R12478 gnd.n3252 gnd.n2395 240.244
R12479 gnd.n3267 gnd.n2395 240.244
R12480 gnd.n3267 gnd.n2396 240.244
R12481 gnd.n2396 gnd.n2373 240.244
R12482 gnd.n3289 gnd.n2373 240.244
R12483 gnd.n3289 gnd.n2375 240.244
R12484 gnd.n2375 gnd.n2355 240.244
R12485 gnd.n3330 gnd.n2355 240.244
R12486 gnd.n3330 gnd.n2348 240.244
R12487 gnd.n3341 gnd.n2348 240.244
R12488 gnd.n3341 gnd.n2341 240.244
R12489 gnd.n3610 gnd.n2341 240.244
R12490 gnd.n3610 gnd.n2342 240.244
R12491 gnd.n2342 gnd.n2323 240.244
R12492 gnd.n3633 gnd.n2323 240.244
R12493 gnd.n4389 gnd.n979 240.244
R12494 gnd.n1907 gnd.n1906 240.244
R12495 gnd.n4401 gnd.n4400 240.244
R12496 gnd.n4413 gnd.n4412 240.244
R12497 gnd.n1895 gnd.n1894 240.244
R12498 gnd.n4425 gnd.n4424 240.244
R12499 gnd.n4437 gnd.n4436 240.244
R12500 gnd.n1883 gnd.n1882 240.244
R12501 gnd.n4450 gnd.n4449 240.244
R12502 gnd.n3879 gnd.n2239 240.244
R12503 gnd.n3876 gnd.n2239 240.244
R12504 gnd.n3876 gnd.n2230 240.244
R12505 gnd.n3873 gnd.n2230 240.244
R12506 gnd.n3873 gnd.n2220 240.244
R12507 gnd.n3870 gnd.n2220 240.244
R12508 gnd.n3870 gnd.n2211 240.244
R12509 gnd.n3867 gnd.n2211 240.244
R12510 gnd.n3867 gnd.n2203 240.244
R12511 gnd.n3864 gnd.n2203 240.244
R12512 gnd.n3864 gnd.n2194 240.244
R12513 gnd.n3861 gnd.n2194 240.244
R12514 gnd.n3861 gnd.n2183 240.244
R12515 gnd.n2183 gnd.n2172 240.244
R12516 gnd.n4127 gnd.n2172 240.244
R12517 gnd.n4127 gnd.n2168 240.244
R12518 gnd.n4135 gnd.n2168 240.244
R12519 gnd.n4135 gnd.n2157 240.244
R12520 gnd.n2157 gnd.n2147 240.244
R12521 gnd.n4162 gnd.n2147 240.244
R12522 gnd.n4162 gnd.n2143 240.244
R12523 gnd.n4170 gnd.n2143 240.244
R12524 gnd.n4170 gnd.n2133 240.244
R12525 gnd.n2133 gnd.n2122 240.244
R12526 gnd.n4197 gnd.n2122 240.244
R12527 gnd.n4197 gnd.n2117 240.244
R12528 gnd.n4217 gnd.n2117 240.244
R12529 gnd.n4217 gnd.n2108 240.244
R12530 gnd.n4203 gnd.n2108 240.244
R12531 gnd.n4203 gnd.n2100 240.244
R12532 gnd.n4204 gnd.n2100 240.244
R12533 gnd.n4204 gnd.n2088 240.244
R12534 gnd.n2088 gnd.n2078 240.244
R12535 gnd.n4266 gnd.n2078 240.244
R12536 gnd.n4267 gnd.n4266 240.244
R12537 gnd.n4267 gnd.n885 240.244
R12538 gnd.n4273 gnd.n885 240.244
R12539 gnd.n4273 gnd.n898 240.244
R12540 gnd.n4293 gnd.n898 240.244
R12541 gnd.n4293 gnd.n909 240.244
R12542 gnd.n4284 gnd.n909 240.244
R12543 gnd.n4284 gnd.n920 240.244
R12544 gnd.n2062 gnd.n920 240.244
R12545 gnd.n2062 gnd.n929 240.244
R12546 gnd.n4348 gnd.n929 240.244
R12547 gnd.n4348 gnd.n940 240.244
R12548 gnd.n4354 gnd.n940 240.244
R12549 gnd.n4354 gnd.n949 240.244
R12550 gnd.n4363 gnd.n949 240.244
R12551 gnd.n4363 gnd.n960 240.244
R12552 gnd.n4371 gnd.n960 240.244
R12553 gnd.n4371 gnd.n970 240.244
R12554 gnd.n4469 gnd.n970 240.244
R12555 gnd.n3916 gnd.n3915 240.244
R12556 gnd.n3912 gnd.n3911 240.244
R12557 gnd.n3908 gnd.n3907 240.244
R12558 gnd.n3904 gnd.n3903 240.244
R12559 gnd.n3900 gnd.n3899 240.244
R12560 gnd.n3896 gnd.n3895 240.244
R12561 gnd.n3892 gnd.n3891 240.244
R12562 gnd.n3888 gnd.n3887 240.244
R12563 gnd.n3843 gnd.n3762 240.244
R12564 gnd.n4051 gnd.n2240 240.244
R12565 gnd.n4051 gnd.n2241 240.244
R12566 gnd.n2241 gnd.n2231 240.244
R12567 gnd.n2231 gnd.n2222 240.244
R12568 gnd.n4071 gnd.n2222 240.244
R12569 gnd.n4071 gnd.n2223 240.244
R12570 gnd.n2223 gnd.n2212 240.244
R12571 gnd.n2212 gnd.n2204 240.244
R12572 gnd.n4091 gnd.n2204 240.244
R12573 gnd.n4091 gnd.n2205 240.244
R12574 gnd.n2205 gnd.n2195 240.244
R12575 gnd.n2195 gnd.n2185 240.244
R12576 gnd.n4115 gnd.n2185 240.244
R12577 gnd.n4115 gnd.n2186 240.244
R12578 gnd.n2186 gnd.n2174 240.244
R12579 gnd.n4110 gnd.n2174 240.244
R12580 gnd.n4110 gnd.n2159 240.244
R12581 gnd.n4150 gnd.n2159 240.244
R12582 gnd.n4150 gnd.n2160 240.244
R12583 gnd.n2160 gnd.n2149 240.244
R12584 gnd.n4145 gnd.n2149 240.244
R12585 gnd.n4145 gnd.n2134 240.244
R12586 gnd.n4185 gnd.n2134 240.244
R12587 gnd.n4185 gnd.n2135 240.244
R12588 gnd.n2135 gnd.n2125 240.244
R12589 gnd.n4180 gnd.n2125 240.244
R12590 gnd.n4180 gnd.n2109 240.244
R12591 gnd.n4228 gnd.n2109 240.244
R12592 gnd.n4228 gnd.n2110 240.244
R12593 gnd.n2110 gnd.n2101 240.244
R12594 gnd.n2101 gnd.n2090 240.244
R12595 gnd.n4255 gnd.n2090 240.244
R12596 gnd.n4255 gnd.n2091 240.244
R12597 gnd.n2091 gnd.n2080 240.244
R12598 gnd.n4250 gnd.n2080 240.244
R12599 gnd.n4250 gnd.n887 240.244
R12600 gnd.n899 gnd.n887 240.244
R12601 gnd.n6000 gnd.n899 240.244
R12602 gnd.n6000 gnd.n900 240.244
R12603 gnd.n5996 gnd.n900 240.244
R12604 gnd.n5996 gnd.n906 240.244
R12605 gnd.n5988 gnd.n906 240.244
R12606 gnd.n5988 gnd.n922 240.244
R12607 gnd.n5984 gnd.n922 240.244
R12608 gnd.n5984 gnd.n927 240.244
R12609 gnd.n5976 gnd.n927 240.244
R12610 gnd.n5976 gnd.n941 240.244
R12611 gnd.n5972 gnd.n941 240.244
R12612 gnd.n5972 gnd.n946 240.244
R12613 gnd.n5964 gnd.n946 240.244
R12614 gnd.n5964 gnd.n962 240.244
R12615 gnd.n5960 gnd.n962 240.244
R12616 gnd.n5960 gnd.n967 240.244
R12617 gnd.n6183 gnd.n712 240.244
R12618 gnd.n6183 gnd.n710 240.244
R12619 gnd.n6187 gnd.n710 240.244
R12620 gnd.n6187 gnd.n706 240.244
R12621 gnd.n6193 gnd.n706 240.244
R12622 gnd.n6193 gnd.n704 240.244
R12623 gnd.n6197 gnd.n704 240.244
R12624 gnd.n6197 gnd.n700 240.244
R12625 gnd.n6203 gnd.n700 240.244
R12626 gnd.n6203 gnd.n698 240.244
R12627 gnd.n6207 gnd.n698 240.244
R12628 gnd.n6207 gnd.n694 240.244
R12629 gnd.n6213 gnd.n694 240.244
R12630 gnd.n6213 gnd.n692 240.244
R12631 gnd.n6217 gnd.n692 240.244
R12632 gnd.n6217 gnd.n688 240.244
R12633 gnd.n6223 gnd.n688 240.244
R12634 gnd.n6223 gnd.n686 240.244
R12635 gnd.n6227 gnd.n686 240.244
R12636 gnd.n6227 gnd.n682 240.244
R12637 gnd.n6233 gnd.n682 240.244
R12638 gnd.n6233 gnd.n680 240.244
R12639 gnd.n6237 gnd.n680 240.244
R12640 gnd.n6237 gnd.n676 240.244
R12641 gnd.n6243 gnd.n676 240.244
R12642 gnd.n6243 gnd.n674 240.244
R12643 gnd.n6247 gnd.n674 240.244
R12644 gnd.n6247 gnd.n670 240.244
R12645 gnd.n6253 gnd.n670 240.244
R12646 gnd.n6253 gnd.n668 240.244
R12647 gnd.n6257 gnd.n668 240.244
R12648 gnd.n6257 gnd.n664 240.244
R12649 gnd.n6263 gnd.n664 240.244
R12650 gnd.n6263 gnd.n662 240.244
R12651 gnd.n6267 gnd.n662 240.244
R12652 gnd.n6267 gnd.n658 240.244
R12653 gnd.n6273 gnd.n658 240.244
R12654 gnd.n6273 gnd.n656 240.244
R12655 gnd.n6277 gnd.n656 240.244
R12656 gnd.n6277 gnd.n652 240.244
R12657 gnd.n6283 gnd.n652 240.244
R12658 gnd.n6283 gnd.n650 240.244
R12659 gnd.n6287 gnd.n650 240.244
R12660 gnd.n6287 gnd.n646 240.244
R12661 gnd.n6293 gnd.n646 240.244
R12662 gnd.n6293 gnd.n644 240.244
R12663 gnd.n6297 gnd.n644 240.244
R12664 gnd.n6297 gnd.n640 240.244
R12665 gnd.n6303 gnd.n640 240.244
R12666 gnd.n6303 gnd.n638 240.244
R12667 gnd.n6307 gnd.n638 240.244
R12668 gnd.n6307 gnd.n634 240.244
R12669 gnd.n6313 gnd.n634 240.244
R12670 gnd.n6313 gnd.n632 240.244
R12671 gnd.n6317 gnd.n632 240.244
R12672 gnd.n6317 gnd.n628 240.244
R12673 gnd.n6323 gnd.n628 240.244
R12674 gnd.n6323 gnd.n626 240.244
R12675 gnd.n6327 gnd.n626 240.244
R12676 gnd.n6327 gnd.n622 240.244
R12677 gnd.n6333 gnd.n622 240.244
R12678 gnd.n6333 gnd.n620 240.244
R12679 gnd.n6337 gnd.n620 240.244
R12680 gnd.n6337 gnd.n616 240.244
R12681 gnd.n6343 gnd.n616 240.244
R12682 gnd.n6343 gnd.n614 240.244
R12683 gnd.n6347 gnd.n614 240.244
R12684 gnd.n6347 gnd.n610 240.244
R12685 gnd.n6353 gnd.n610 240.244
R12686 gnd.n6353 gnd.n608 240.244
R12687 gnd.n6357 gnd.n608 240.244
R12688 gnd.n6357 gnd.n604 240.244
R12689 gnd.n6363 gnd.n604 240.244
R12690 gnd.n6363 gnd.n602 240.244
R12691 gnd.n6367 gnd.n602 240.244
R12692 gnd.n6367 gnd.n598 240.244
R12693 gnd.n6373 gnd.n598 240.244
R12694 gnd.n6373 gnd.n596 240.244
R12695 gnd.n6377 gnd.n596 240.244
R12696 gnd.n6377 gnd.n592 240.244
R12697 gnd.n6383 gnd.n592 240.244
R12698 gnd.n6383 gnd.n590 240.244
R12699 gnd.n6387 gnd.n590 240.244
R12700 gnd.n6387 gnd.n586 240.244
R12701 gnd.n6393 gnd.n586 240.244
R12702 gnd.n6393 gnd.n584 240.244
R12703 gnd.n6397 gnd.n584 240.244
R12704 gnd.n6397 gnd.n580 240.244
R12705 gnd.n6403 gnd.n580 240.244
R12706 gnd.n6403 gnd.n578 240.244
R12707 gnd.n6407 gnd.n578 240.244
R12708 gnd.n6407 gnd.n574 240.244
R12709 gnd.n6413 gnd.n574 240.244
R12710 gnd.n6413 gnd.n572 240.244
R12711 gnd.n6417 gnd.n572 240.244
R12712 gnd.n6417 gnd.n568 240.244
R12713 gnd.n6423 gnd.n568 240.244
R12714 gnd.n6423 gnd.n566 240.244
R12715 gnd.n6427 gnd.n566 240.244
R12716 gnd.n6427 gnd.n562 240.244
R12717 gnd.n6433 gnd.n562 240.244
R12718 gnd.n6433 gnd.n560 240.244
R12719 gnd.n6437 gnd.n560 240.244
R12720 gnd.n6437 gnd.n556 240.244
R12721 gnd.n6443 gnd.n556 240.244
R12722 gnd.n6443 gnd.n554 240.244
R12723 gnd.n6447 gnd.n554 240.244
R12724 gnd.n6447 gnd.n550 240.244
R12725 gnd.n6453 gnd.n550 240.244
R12726 gnd.n6453 gnd.n548 240.244
R12727 gnd.n6457 gnd.n548 240.244
R12728 gnd.n6457 gnd.n544 240.244
R12729 gnd.n6463 gnd.n544 240.244
R12730 gnd.n6463 gnd.n542 240.244
R12731 gnd.n6467 gnd.n542 240.244
R12732 gnd.n6467 gnd.n538 240.244
R12733 gnd.n6473 gnd.n538 240.244
R12734 gnd.n6473 gnd.n536 240.244
R12735 gnd.n6477 gnd.n536 240.244
R12736 gnd.n6477 gnd.n532 240.244
R12737 gnd.n6483 gnd.n532 240.244
R12738 gnd.n6483 gnd.n530 240.244
R12739 gnd.n6487 gnd.n530 240.244
R12740 gnd.n6487 gnd.n526 240.244
R12741 gnd.n6494 gnd.n526 240.244
R12742 gnd.n6494 gnd.n524 240.244
R12743 gnd.n6498 gnd.n524 240.244
R12744 gnd.n6498 gnd.n521 240.244
R12745 gnd.n6504 gnd.n519 240.244
R12746 gnd.n6508 gnd.n519 240.244
R12747 gnd.n6508 gnd.n515 240.244
R12748 gnd.n6514 gnd.n515 240.244
R12749 gnd.n6514 gnd.n513 240.244
R12750 gnd.n6518 gnd.n513 240.244
R12751 gnd.n6518 gnd.n509 240.244
R12752 gnd.n6524 gnd.n509 240.244
R12753 gnd.n6524 gnd.n507 240.244
R12754 gnd.n6528 gnd.n507 240.244
R12755 gnd.n6528 gnd.n503 240.244
R12756 gnd.n6534 gnd.n503 240.244
R12757 gnd.n6534 gnd.n501 240.244
R12758 gnd.n6538 gnd.n501 240.244
R12759 gnd.n6538 gnd.n497 240.244
R12760 gnd.n6544 gnd.n497 240.244
R12761 gnd.n6544 gnd.n495 240.244
R12762 gnd.n6548 gnd.n495 240.244
R12763 gnd.n6548 gnd.n491 240.244
R12764 gnd.n6554 gnd.n491 240.244
R12765 gnd.n6554 gnd.n489 240.244
R12766 gnd.n6558 gnd.n489 240.244
R12767 gnd.n6558 gnd.n485 240.244
R12768 gnd.n6564 gnd.n485 240.244
R12769 gnd.n6564 gnd.n483 240.244
R12770 gnd.n6568 gnd.n483 240.244
R12771 gnd.n6568 gnd.n479 240.244
R12772 gnd.n6574 gnd.n479 240.244
R12773 gnd.n6574 gnd.n477 240.244
R12774 gnd.n6578 gnd.n477 240.244
R12775 gnd.n6578 gnd.n473 240.244
R12776 gnd.n6584 gnd.n473 240.244
R12777 gnd.n6584 gnd.n471 240.244
R12778 gnd.n6588 gnd.n471 240.244
R12779 gnd.n6588 gnd.n467 240.244
R12780 gnd.n6594 gnd.n467 240.244
R12781 gnd.n6594 gnd.n465 240.244
R12782 gnd.n6598 gnd.n465 240.244
R12783 gnd.n6598 gnd.n461 240.244
R12784 gnd.n6604 gnd.n461 240.244
R12785 gnd.n6604 gnd.n459 240.244
R12786 gnd.n6608 gnd.n459 240.244
R12787 gnd.n6608 gnd.n455 240.244
R12788 gnd.n6614 gnd.n455 240.244
R12789 gnd.n6614 gnd.n453 240.244
R12790 gnd.n6618 gnd.n453 240.244
R12791 gnd.n6618 gnd.n449 240.244
R12792 gnd.n6624 gnd.n449 240.244
R12793 gnd.n6624 gnd.n447 240.244
R12794 gnd.n6628 gnd.n447 240.244
R12795 gnd.n6628 gnd.n443 240.244
R12796 gnd.n6634 gnd.n443 240.244
R12797 gnd.n6634 gnd.n441 240.244
R12798 gnd.n6638 gnd.n441 240.244
R12799 gnd.n6638 gnd.n437 240.244
R12800 gnd.n6644 gnd.n437 240.244
R12801 gnd.n6644 gnd.n435 240.244
R12802 gnd.n6648 gnd.n435 240.244
R12803 gnd.n6648 gnd.n431 240.244
R12804 gnd.n6654 gnd.n431 240.244
R12805 gnd.n6654 gnd.n429 240.244
R12806 gnd.n6658 gnd.n429 240.244
R12807 gnd.n6658 gnd.n425 240.244
R12808 gnd.n6664 gnd.n425 240.244
R12809 gnd.n6664 gnd.n423 240.244
R12810 gnd.n6668 gnd.n423 240.244
R12811 gnd.n6668 gnd.n419 240.244
R12812 gnd.n6674 gnd.n419 240.244
R12813 gnd.n6674 gnd.n417 240.244
R12814 gnd.n6678 gnd.n417 240.244
R12815 gnd.n6678 gnd.n413 240.244
R12816 gnd.n6684 gnd.n413 240.244
R12817 gnd.n6684 gnd.n411 240.244
R12818 gnd.n6688 gnd.n411 240.244
R12819 gnd.n6688 gnd.n407 240.244
R12820 gnd.n6694 gnd.n407 240.244
R12821 gnd.n6694 gnd.n405 240.244
R12822 gnd.n6698 gnd.n405 240.244
R12823 gnd.n6698 gnd.n401 240.244
R12824 gnd.n6704 gnd.n401 240.244
R12825 gnd.n6704 gnd.n399 240.244
R12826 gnd.n6709 gnd.n399 240.244
R12827 gnd.n6709 gnd.n395 240.244
R12828 gnd.n6715 gnd.n395 240.244
R12829 gnd.n4300 gnd.n882 240.244
R12830 gnd.n4300 gnd.n4296 240.244
R12831 gnd.n4306 gnd.n4296 240.244
R12832 gnd.n4307 gnd.n4306 240.244
R12833 gnd.n4308 gnd.n4307 240.244
R12834 gnd.n4308 gnd.n2063 240.244
R12835 gnd.n4338 gnd.n2063 240.244
R12836 gnd.n4338 gnd.n2064 240.244
R12837 gnd.n4334 gnd.n2064 240.244
R12838 gnd.n4334 gnd.n4333 240.244
R12839 gnd.n4333 gnd.n4332 240.244
R12840 gnd.n4332 gnd.n4316 240.244
R12841 gnd.n4328 gnd.n4316 240.244
R12842 gnd.n4328 gnd.n4327 240.244
R12843 gnd.n4327 gnd.n4326 240.244
R12844 gnd.n4326 gnd.n1853 240.244
R12845 gnd.n4466 gnd.n1853 240.244
R12846 gnd.n4466 gnd.n1854 240.244
R12847 gnd.n4462 gnd.n1854 240.244
R12848 gnd.n4462 gnd.n4461 240.244
R12849 gnd.n4461 gnd.n1863 240.244
R12850 gnd.n1863 gnd.n1839 240.244
R12851 gnd.n4481 gnd.n1839 240.244
R12852 gnd.n4481 gnd.n1835 240.244
R12853 gnd.n4487 gnd.n1835 240.244
R12854 gnd.n4487 gnd.n1826 240.244
R12855 gnd.n4497 gnd.n1826 240.244
R12856 gnd.n4497 gnd.n1822 240.244
R12857 gnd.n4503 gnd.n1822 240.244
R12858 gnd.n4503 gnd.n1810 240.244
R12859 gnd.n4531 gnd.n1810 240.244
R12860 gnd.n4531 gnd.n1805 240.244
R12861 gnd.n4546 gnd.n1805 240.244
R12862 gnd.n4546 gnd.n1806 240.244
R12863 gnd.n4542 gnd.n1806 240.244
R12864 gnd.n4542 gnd.n4541 240.244
R12865 gnd.n4541 gnd.n1116 240.244
R12866 gnd.n5824 gnd.n1116 240.244
R12867 gnd.n5824 gnd.n1117 240.244
R12868 gnd.n5820 gnd.n1117 240.244
R12869 gnd.n5820 gnd.n1123 240.244
R12870 gnd.n4651 gnd.n1123 240.244
R12871 gnd.n4651 gnd.n1709 240.244
R12872 gnd.n4662 gnd.n1709 240.244
R12873 gnd.n4662 gnd.n1710 240.244
R12874 gnd.n4658 gnd.n1710 240.244
R12875 gnd.n4658 gnd.n1689 240.244
R12876 gnd.n4691 gnd.n1689 240.244
R12877 gnd.n4691 gnd.n1684 240.244
R12878 gnd.n4699 gnd.n1684 240.244
R12879 gnd.n4699 gnd.n1685 240.244
R12880 gnd.n1685 gnd.n1661 240.244
R12881 gnd.n4727 gnd.n1661 240.244
R12882 gnd.n4727 gnd.n1657 240.244
R12883 gnd.n4733 gnd.n1657 240.244
R12884 gnd.n4733 gnd.n1643 240.244
R12885 gnd.n4753 gnd.n1643 240.244
R12886 gnd.n4753 gnd.n1638 240.244
R12887 gnd.n4761 gnd.n1638 240.244
R12888 gnd.n4761 gnd.n1639 240.244
R12889 gnd.n1639 gnd.n1617 240.244
R12890 gnd.n4809 gnd.n1617 240.244
R12891 gnd.n4809 gnd.n1610 240.244
R12892 gnd.n4817 gnd.n1610 240.244
R12893 gnd.n4817 gnd.n1613 240.244
R12894 gnd.n1613 gnd.n1592 240.244
R12895 gnd.n4849 gnd.n1592 240.244
R12896 gnd.n4849 gnd.n1587 240.244
R12897 gnd.n4857 gnd.n1587 240.244
R12898 gnd.n4857 gnd.n1588 240.244
R12899 gnd.n1588 gnd.n1562 240.244
R12900 gnd.n4918 gnd.n1562 240.244
R12901 gnd.n4918 gnd.n1557 240.244
R12902 gnd.n4926 gnd.n1557 240.244
R12903 gnd.n4926 gnd.n1558 240.244
R12904 gnd.n1558 gnd.n1538 240.244
R12905 gnd.n4951 gnd.n1538 240.244
R12906 gnd.n4951 gnd.n1533 240.244
R12907 gnd.n4959 gnd.n1533 240.244
R12908 gnd.n4959 gnd.n1534 240.244
R12909 gnd.n1534 gnd.n1517 240.244
R12910 gnd.n5005 gnd.n1517 240.244
R12911 gnd.n5005 gnd.n1512 240.244
R12912 gnd.n5013 gnd.n1512 240.244
R12913 gnd.n5013 gnd.n1513 240.244
R12914 gnd.n1513 gnd.n1492 240.244
R12915 gnd.n5042 gnd.n1492 240.244
R12916 gnd.n5042 gnd.n1488 240.244
R12917 gnd.n5048 gnd.n1488 240.244
R12918 gnd.n5048 gnd.n1401 240.244
R12919 gnd.n5185 gnd.n1401 240.244
R12920 gnd.n5185 gnd.n1397 240.244
R12921 gnd.n5191 gnd.n1397 240.244
R12922 gnd.n5191 gnd.n1388 240.244
R12923 gnd.n5201 gnd.n1388 240.244
R12924 gnd.n5201 gnd.n1384 240.244
R12925 gnd.n5207 gnd.n1384 240.244
R12926 gnd.n5207 gnd.n1375 240.244
R12927 gnd.n5217 gnd.n1375 240.244
R12928 gnd.n5217 gnd.n1371 240.244
R12929 gnd.n5223 gnd.n1371 240.244
R12930 gnd.n5223 gnd.n1362 240.244
R12931 gnd.n5233 gnd.n1362 240.244
R12932 gnd.n5233 gnd.n1358 240.244
R12933 gnd.n5240 gnd.n1358 240.244
R12934 gnd.n5240 gnd.n1232 240.244
R12935 gnd.n5714 gnd.n1232 240.244
R12936 gnd.n5714 gnd.n1233 240.244
R12937 gnd.n5710 gnd.n1233 240.244
R12938 gnd.n5710 gnd.n1239 240.244
R12939 gnd.n5275 gnd.n1239 240.244
R12940 gnd.n5473 gnd.n5275 240.244
R12941 gnd.n5473 gnd.n5276 240.244
R12942 gnd.n5469 gnd.n5276 240.244
R12943 gnd.n5469 gnd.n5284 240.244
R12944 gnd.n5390 gnd.n5284 240.244
R12945 gnd.n5390 gnd.n5386 240.244
R12946 gnd.n5398 gnd.n5386 240.244
R12947 gnd.n5398 gnd.n5387 240.244
R12948 gnd.n5387 gnd.n5342 240.244
R12949 gnd.n5428 gnd.n5342 240.244
R12950 gnd.n5428 gnd.n5337 240.244
R12951 gnd.n5437 gnd.n5337 240.244
R12952 gnd.n5437 gnd.n5338 240.244
R12953 gnd.n5338 gnd.n389 240.244
R12954 gnd.n6720 gnd.n389 240.244
R12955 gnd.n6720 gnd.n390 240.244
R12956 gnd.n6716 gnd.n390 240.244
R12957 gnd.n6177 gnd.n716 240.244
R12958 gnd.n6173 gnd.n716 240.244
R12959 gnd.n6173 gnd.n718 240.244
R12960 gnd.n6169 gnd.n718 240.244
R12961 gnd.n6169 gnd.n723 240.244
R12962 gnd.n6165 gnd.n723 240.244
R12963 gnd.n6165 gnd.n725 240.244
R12964 gnd.n6161 gnd.n725 240.244
R12965 gnd.n6161 gnd.n731 240.244
R12966 gnd.n6157 gnd.n731 240.244
R12967 gnd.n6157 gnd.n733 240.244
R12968 gnd.n6153 gnd.n733 240.244
R12969 gnd.n6153 gnd.n739 240.244
R12970 gnd.n6149 gnd.n739 240.244
R12971 gnd.n6149 gnd.n741 240.244
R12972 gnd.n6145 gnd.n741 240.244
R12973 gnd.n6145 gnd.n747 240.244
R12974 gnd.n6141 gnd.n747 240.244
R12975 gnd.n6141 gnd.n749 240.244
R12976 gnd.n6137 gnd.n749 240.244
R12977 gnd.n6137 gnd.n755 240.244
R12978 gnd.n6133 gnd.n755 240.244
R12979 gnd.n6133 gnd.n757 240.244
R12980 gnd.n6129 gnd.n757 240.244
R12981 gnd.n6129 gnd.n763 240.244
R12982 gnd.n6125 gnd.n763 240.244
R12983 gnd.n6125 gnd.n765 240.244
R12984 gnd.n6121 gnd.n765 240.244
R12985 gnd.n6121 gnd.n771 240.244
R12986 gnd.n6117 gnd.n771 240.244
R12987 gnd.n6117 gnd.n773 240.244
R12988 gnd.n6113 gnd.n773 240.244
R12989 gnd.n6113 gnd.n779 240.244
R12990 gnd.n6109 gnd.n779 240.244
R12991 gnd.n6109 gnd.n781 240.244
R12992 gnd.n6105 gnd.n781 240.244
R12993 gnd.n6105 gnd.n787 240.244
R12994 gnd.n6101 gnd.n787 240.244
R12995 gnd.n6101 gnd.n789 240.244
R12996 gnd.n6097 gnd.n789 240.244
R12997 gnd.n6097 gnd.n795 240.244
R12998 gnd.n6093 gnd.n795 240.244
R12999 gnd.n6093 gnd.n797 240.244
R13000 gnd.n6089 gnd.n797 240.244
R13001 gnd.n6089 gnd.n803 240.244
R13002 gnd.n6085 gnd.n803 240.244
R13003 gnd.n6085 gnd.n805 240.244
R13004 gnd.n6081 gnd.n805 240.244
R13005 gnd.n6081 gnd.n811 240.244
R13006 gnd.n6077 gnd.n811 240.244
R13007 gnd.n6077 gnd.n813 240.244
R13008 gnd.n6073 gnd.n813 240.244
R13009 gnd.n6073 gnd.n819 240.244
R13010 gnd.n6069 gnd.n819 240.244
R13011 gnd.n6069 gnd.n821 240.244
R13012 gnd.n6065 gnd.n821 240.244
R13013 gnd.n6065 gnd.n827 240.244
R13014 gnd.n6061 gnd.n827 240.244
R13015 gnd.n6061 gnd.n829 240.244
R13016 gnd.n6057 gnd.n829 240.244
R13017 gnd.n6057 gnd.n835 240.244
R13018 gnd.n6053 gnd.n835 240.244
R13019 gnd.n6053 gnd.n837 240.244
R13020 gnd.n6049 gnd.n837 240.244
R13021 gnd.n6049 gnd.n843 240.244
R13022 gnd.n6045 gnd.n843 240.244
R13023 gnd.n6045 gnd.n845 240.244
R13024 gnd.n6041 gnd.n845 240.244
R13025 gnd.n6041 gnd.n851 240.244
R13026 gnd.n6037 gnd.n851 240.244
R13027 gnd.n6037 gnd.n853 240.244
R13028 gnd.n6033 gnd.n853 240.244
R13029 gnd.n6033 gnd.n859 240.244
R13030 gnd.n6029 gnd.n859 240.244
R13031 gnd.n6029 gnd.n861 240.244
R13032 gnd.n6025 gnd.n861 240.244
R13033 gnd.n6025 gnd.n867 240.244
R13034 gnd.n6021 gnd.n867 240.244
R13035 gnd.n6021 gnd.n869 240.244
R13036 gnd.n6017 gnd.n869 240.244
R13037 gnd.n6017 gnd.n875 240.244
R13038 gnd.n6013 gnd.n875 240.244
R13039 gnd.n6013 gnd.n877 240.244
R13040 gnd.n6009 gnd.n877 240.244
R13041 gnd.n1922 gnd.n1841 240.244
R13042 gnd.n1922 gnd.n1834 240.244
R13043 gnd.n1923 gnd.n1834 240.244
R13044 gnd.n1923 gnd.n1828 240.244
R13045 gnd.n1926 gnd.n1828 240.244
R13046 gnd.n1926 gnd.n1821 240.244
R13047 gnd.n1927 gnd.n1821 240.244
R13048 gnd.n1927 gnd.n1812 240.244
R13049 gnd.n1812 gnd.n1802 240.244
R13050 gnd.n4548 gnd.n1802 240.244
R13051 gnd.n4548 gnd.n1798 240.244
R13052 gnd.n4554 gnd.n1798 240.244
R13053 gnd.n4555 gnd.n4554 240.244
R13054 gnd.n4556 gnd.n4555 240.244
R13055 gnd.n4556 gnd.n1113 240.244
R13056 gnd.n4620 gnd.n1113 240.244
R13057 gnd.n4620 gnd.n1125 240.244
R13058 gnd.n4562 gnd.n1125 240.244
R13059 gnd.n4562 gnd.n1714 240.244
R13060 gnd.n4564 gnd.n1714 240.244
R13061 gnd.n4564 gnd.n1708 240.244
R13062 gnd.n4567 gnd.n1708 240.244
R13063 gnd.n4568 gnd.n4567 240.244
R13064 gnd.n4568 gnd.n1698 240.244
R13065 gnd.n1698 gnd.n1690 240.244
R13066 gnd.n4571 gnd.n1690 240.244
R13067 gnd.n4571 gnd.n1683 240.244
R13068 gnd.n4572 gnd.n1683 240.244
R13069 gnd.n4573 gnd.n4572 240.244
R13070 gnd.n4573 gnd.n1663 240.244
R13071 gnd.n4576 gnd.n1663 240.244
R13072 gnd.n4576 gnd.n1655 240.244
R13073 gnd.n4577 gnd.n1655 240.244
R13074 gnd.n4577 gnd.n1645 240.244
R13075 gnd.n4580 gnd.n1645 240.244
R13076 gnd.n4580 gnd.n1637 240.244
R13077 gnd.n4581 gnd.n1637 240.244
R13078 gnd.n4581 gnd.n1628 240.244
R13079 gnd.n1628 gnd.n1618 240.244
R13080 gnd.n1618 gnd.n1607 240.244
R13081 gnd.n4819 gnd.n1607 240.244
R13082 gnd.n4819 gnd.n1602 240.244
R13083 gnd.n4839 gnd.n1602 240.244
R13084 gnd.n4839 gnd.n1594 240.244
R13085 gnd.n4824 gnd.n1594 240.244
R13086 gnd.n4824 gnd.n1585 240.244
R13087 gnd.n4825 gnd.n1585 240.244
R13088 gnd.n4826 gnd.n4825 240.244
R13089 gnd.n4826 gnd.n1564 240.244
R13090 gnd.n1564 gnd.n1554 240.244
R13091 gnd.n4928 gnd.n1554 240.244
R13092 gnd.n4928 gnd.n1549 240.244
R13093 gnd.n4935 gnd.n1549 240.244
R13094 gnd.n4935 gnd.n1540 240.244
R13095 gnd.n1540 gnd.n1531 240.244
R13096 gnd.n4961 gnd.n1531 240.244
R13097 gnd.n4961 gnd.n1526 240.244
R13098 gnd.n4994 gnd.n1526 240.244
R13099 gnd.n4994 gnd.n1519 240.244
R13100 gnd.n4966 gnd.n1519 240.244
R13101 gnd.n4966 gnd.n1511 240.244
R13102 gnd.n4970 gnd.n1511 240.244
R13103 gnd.n4971 gnd.n4970 240.244
R13104 gnd.n4971 gnd.n1494 240.244
R13105 gnd.n4974 gnd.n1494 240.244
R13106 gnd.n4974 gnd.n1485 240.244
R13107 gnd.n4975 gnd.n1485 240.244
R13108 gnd.n4975 gnd.n1403 240.244
R13109 gnd.n1403 gnd.n1393 240.244
R13110 gnd.n5193 gnd.n1393 240.244
R13111 gnd.n5193 gnd.n1389 240.244
R13112 gnd.n5199 gnd.n1389 240.244
R13113 gnd.n5199 gnd.n1380 240.244
R13114 gnd.n5209 gnd.n1380 240.244
R13115 gnd.n5209 gnd.n1376 240.244
R13116 gnd.n5215 gnd.n1376 240.244
R13117 gnd.n5215 gnd.n1368 240.244
R13118 gnd.n5225 gnd.n1368 240.244
R13119 gnd.n5225 gnd.n1364 240.244
R13120 gnd.n5231 gnd.n1364 240.244
R13121 gnd.n5231 gnd.n1355 240.244
R13122 gnd.n5242 gnd.n1355 240.244
R13123 gnd.n1920 gnd.n1919 240.244
R13124 gnd.n1951 gnd.n1950 240.244
R13125 gnd.n1916 gnd.n1915 240.244
R13126 gnd.n4384 gnd.n4383 240.244
R13127 gnd.n1911 gnd.n1910 240.244
R13128 gnd.n4395 gnd.n4394 240.244
R13129 gnd.n4407 gnd.n4406 240.244
R13130 gnd.n1899 gnd.n1898 240.244
R13131 gnd.n4419 gnd.n4418 240.244
R13132 gnd.n4431 gnd.n4430 240.244
R13133 gnd.n1887 gnd.n1886 240.244
R13134 gnd.n4443 gnd.n4442 240.244
R13135 gnd.n4457 gnd.n4456 240.244
R13136 gnd.n1846 gnd.n1843 240.244
R13137 gnd.n4479 gnd.n1833 240.244
R13138 gnd.n4489 gnd.n1833 240.244
R13139 gnd.n4489 gnd.n1829 240.244
R13140 gnd.n4495 gnd.n1829 240.244
R13141 gnd.n4495 gnd.n1819 240.244
R13142 gnd.n4505 gnd.n1819 240.244
R13143 gnd.n4505 gnd.n1813 240.244
R13144 gnd.n4529 gnd.n1813 240.244
R13145 gnd.n4529 gnd.n1814 240.244
R13146 gnd.n1814 gnd.n1804 240.244
R13147 gnd.n4511 gnd.n1804 240.244
R13148 gnd.n4512 gnd.n4511 240.244
R13149 gnd.n4515 gnd.n4512 240.244
R13150 gnd.n4516 gnd.n4515 240.244
R13151 gnd.n4516 gnd.n1115 240.244
R13152 gnd.n1127 gnd.n1115 240.244
R13153 gnd.n5818 gnd.n1127 240.244
R13154 gnd.n5818 gnd.n1128 240.244
R13155 gnd.n1133 gnd.n1128 240.244
R13156 gnd.n1134 gnd.n1133 240.244
R13157 gnd.n1135 gnd.n1134 240.244
R13158 gnd.n1701 gnd.n1135 240.244
R13159 gnd.n1701 gnd.n1138 240.244
R13160 gnd.n1139 gnd.n1138 240.244
R13161 gnd.n1140 gnd.n1139 240.244
R13162 gnd.n1680 gnd.n1140 240.244
R13163 gnd.n1680 gnd.n1143 240.244
R13164 gnd.n1144 gnd.n1143 240.244
R13165 gnd.n1145 gnd.n1144 240.244
R13166 gnd.n4725 gnd.n1145 240.244
R13167 gnd.n4725 gnd.n1148 240.244
R13168 gnd.n1149 gnd.n1148 240.244
R13169 gnd.n1150 gnd.n1149 240.244
R13170 gnd.n4751 gnd.n1150 240.244
R13171 gnd.n4751 gnd.n1153 240.244
R13172 gnd.n1154 gnd.n1153 240.244
R13173 gnd.n1155 gnd.n1154 240.244
R13174 gnd.n4794 gnd.n1155 240.244
R13175 gnd.n4794 gnd.n1158 240.244
R13176 gnd.n1159 gnd.n1158 240.244
R13177 gnd.n1160 gnd.n1159 240.244
R13178 gnd.n1611 gnd.n1160 240.244
R13179 gnd.n1611 gnd.n1163 240.244
R13180 gnd.n1164 gnd.n1163 240.244
R13181 gnd.n1165 gnd.n1164 240.244
R13182 gnd.n1586 gnd.n1165 240.244
R13183 gnd.n1586 gnd.n1168 240.244
R13184 gnd.n1169 gnd.n1168 240.244
R13185 gnd.n1170 gnd.n1169 240.244
R13186 gnd.n1566 gnd.n1170 240.244
R13187 gnd.n1566 gnd.n1173 240.244
R13188 gnd.n1174 gnd.n1173 240.244
R13189 gnd.n1175 gnd.n1174 240.244
R13190 gnd.n4949 gnd.n1175 240.244
R13191 gnd.n4949 gnd.n1178 240.244
R13192 gnd.n1179 gnd.n1178 240.244
R13193 gnd.n1180 gnd.n1179 240.244
R13194 gnd.n4995 gnd.n1180 240.244
R13195 gnd.n4995 gnd.n1183 240.244
R13196 gnd.n1184 gnd.n1183 240.244
R13197 gnd.n1185 gnd.n1184 240.244
R13198 gnd.n4968 gnd.n1185 240.244
R13199 gnd.n4968 gnd.n1188 240.244
R13200 gnd.n1189 gnd.n1188 240.244
R13201 gnd.n1190 gnd.n1189 240.244
R13202 gnd.n1487 gnd.n1190 240.244
R13203 gnd.n1487 gnd.n1193 240.244
R13204 gnd.n1194 gnd.n1193 240.244
R13205 gnd.n1195 gnd.n1194 240.244
R13206 gnd.n1396 gnd.n1195 240.244
R13207 gnd.n1396 gnd.n1198 240.244
R13208 gnd.n1199 gnd.n1198 240.244
R13209 gnd.n1200 gnd.n1199 240.244
R13210 gnd.n1383 gnd.n1200 240.244
R13211 gnd.n1383 gnd.n1203 240.244
R13212 gnd.n1204 gnd.n1203 240.244
R13213 gnd.n1205 gnd.n1204 240.244
R13214 gnd.n1370 gnd.n1205 240.244
R13215 gnd.n1370 gnd.n1208 240.244
R13216 gnd.n1209 gnd.n1208 240.244
R13217 gnd.n1210 gnd.n1209 240.244
R13218 gnd.n1215 gnd.n1210 240.244
R13219 gnd.n5249 gnd.n5248 240.244
R13220 gnd.n5252 gnd.n5251 240.244
R13221 gnd.n5259 gnd.n5258 240.244
R13222 gnd.n5262 gnd.n5261 240.244
R13223 gnd.n5264 gnd.n5263 240.244
R13224 gnd.n5484 gnd.n5483 240.244
R13225 gnd.n5494 gnd.n5493 240.244
R13226 gnd.n5496 gnd.n5495 240.244
R13227 gnd.n5504 gnd.n5503 240.244
R13228 gnd.n5514 gnd.n5513 240.244
R13229 gnd.n5516 gnd.n5515 240.244
R13230 gnd.n5524 gnd.n5523 240.244
R13231 gnd.n5536 gnd.n5535 240.244
R13232 gnd.n5716 gnd.n1214 240.244
R13233 gnd.n1094 gnd.n1093 240.132
R13234 gnd.n1420 gnd.n1419 240.132
R13235 gnd.n6184 gnd.n711 225.874
R13236 gnd.n6185 gnd.n6184 225.874
R13237 gnd.n6186 gnd.n6185 225.874
R13238 gnd.n6186 gnd.n705 225.874
R13239 gnd.n6194 gnd.n705 225.874
R13240 gnd.n6195 gnd.n6194 225.874
R13241 gnd.n6196 gnd.n6195 225.874
R13242 gnd.n6196 gnd.n699 225.874
R13243 gnd.n6204 gnd.n699 225.874
R13244 gnd.n6205 gnd.n6204 225.874
R13245 gnd.n6206 gnd.n6205 225.874
R13246 gnd.n6206 gnd.n693 225.874
R13247 gnd.n6214 gnd.n693 225.874
R13248 gnd.n6215 gnd.n6214 225.874
R13249 gnd.n6216 gnd.n6215 225.874
R13250 gnd.n6216 gnd.n687 225.874
R13251 gnd.n6224 gnd.n687 225.874
R13252 gnd.n6225 gnd.n6224 225.874
R13253 gnd.n6226 gnd.n6225 225.874
R13254 gnd.n6226 gnd.n681 225.874
R13255 gnd.n6234 gnd.n681 225.874
R13256 gnd.n6235 gnd.n6234 225.874
R13257 gnd.n6236 gnd.n6235 225.874
R13258 gnd.n6236 gnd.n675 225.874
R13259 gnd.n6244 gnd.n675 225.874
R13260 gnd.n6245 gnd.n6244 225.874
R13261 gnd.n6246 gnd.n6245 225.874
R13262 gnd.n6246 gnd.n669 225.874
R13263 gnd.n6254 gnd.n669 225.874
R13264 gnd.n6255 gnd.n6254 225.874
R13265 gnd.n6256 gnd.n6255 225.874
R13266 gnd.n6256 gnd.n663 225.874
R13267 gnd.n6264 gnd.n663 225.874
R13268 gnd.n6265 gnd.n6264 225.874
R13269 gnd.n6266 gnd.n6265 225.874
R13270 gnd.n6266 gnd.n657 225.874
R13271 gnd.n6274 gnd.n657 225.874
R13272 gnd.n6275 gnd.n6274 225.874
R13273 gnd.n6276 gnd.n6275 225.874
R13274 gnd.n6276 gnd.n651 225.874
R13275 gnd.n6284 gnd.n651 225.874
R13276 gnd.n6285 gnd.n6284 225.874
R13277 gnd.n6286 gnd.n6285 225.874
R13278 gnd.n6286 gnd.n645 225.874
R13279 gnd.n6294 gnd.n645 225.874
R13280 gnd.n6295 gnd.n6294 225.874
R13281 gnd.n6296 gnd.n6295 225.874
R13282 gnd.n6296 gnd.n639 225.874
R13283 gnd.n6304 gnd.n639 225.874
R13284 gnd.n6305 gnd.n6304 225.874
R13285 gnd.n6306 gnd.n6305 225.874
R13286 gnd.n6306 gnd.n633 225.874
R13287 gnd.n6314 gnd.n633 225.874
R13288 gnd.n6315 gnd.n6314 225.874
R13289 gnd.n6316 gnd.n6315 225.874
R13290 gnd.n6316 gnd.n627 225.874
R13291 gnd.n6324 gnd.n627 225.874
R13292 gnd.n6325 gnd.n6324 225.874
R13293 gnd.n6326 gnd.n6325 225.874
R13294 gnd.n6326 gnd.n621 225.874
R13295 gnd.n6334 gnd.n621 225.874
R13296 gnd.n6335 gnd.n6334 225.874
R13297 gnd.n6336 gnd.n6335 225.874
R13298 gnd.n6336 gnd.n615 225.874
R13299 gnd.n6344 gnd.n615 225.874
R13300 gnd.n6345 gnd.n6344 225.874
R13301 gnd.n6346 gnd.n6345 225.874
R13302 gnd.n6346 gnd.n609 225.874
R13303 gnd.n6354 gnd.n609 225.874
R13304 gnd.n6355 gnd.n6354 225.874
R13305 gnd.n6356 gnd.n6355 225.874
R13306 gnd.n6356 gnd.n603 225.874
R13307 gnd.n6364 gnd.n603 225.874
R13308 gnd.n6365 gnd.n6364 225.874
R13309 gnd.n6366 gnd.n6365 225.874
R13310 gnd.n6366 gnd.n597 225.874
R13311 gnd.n6374 gnd.n597 225.874
R13312 gnd.n6375 gnd.n6374 225.874
R13313 gnd.n6376 gnd.n6375 225.874
R13314 gnd.n6376 gnd.n591 225.874
R13315 gnd.n6384 gnd.n591 225.874
R13316 gnd.n6385 gnd.n6384 225.874
R13317 gnd.n6386 gnd.n6385 225.874
R13318 gnd.n6386 gnd.n585 225.874
R13319 gnd.n6394 gnd.n585 225.874
R13320 gnd.n6395 gnd.n6394 225.874
R13321 gnd.n6396 gnd.n6395 225.874
R13322 gnd.n6396 gnd.n579 225.874
R13323 gnd.n6404 gnd.n579 225.874
R13324 gnd.n6405 gnd.n6404 225.874
R13325 gnd.n6406 gnd.n6405 225.874
R13326 gnd.n6406 gnd.n573 225.874
R13327 gnd.n6414 gnd.n573 225.874
R13328 gnd.n6415 gnd.n6414 225.874
R13329 gnd.n6416 gnd.n6415 225.874
R13330 gnd.n6416 gnd.n567 225.874
R13331 gnd.n6424 gnd.n567 225.874
R13332 gnd.n6425 gnd.n6424 225.874
R13333 gnd.n6426 gnd.n6425 225.874
R13334 gnd.n6426 gnd.n561 225.874
R13335 gnd.n6434 gnd.n561 225.874
R13336 gnd.n6435 gnd.n6434 225.874
R13337 gnd.n6436 gnd.n6435 225.874
R13338 gnd.n6436 gnd.n555 225.874
R13339 gnd.n6444 gnd.n555 225.874
R13340 gnd.n6445 gnd.n6444 225.874
R13341 gnd.n6446 gnd.n6445 225.874
R13342 gnd.n6446 gnd.n549 225.874
R13343 gnd.n6454 gnd.n549 225.874
R13344 gnd.n6455 gnd.n6454 225.874
R13345 gnd.n6456 gnd.n6455 225.874
R13346 gnd.n6456 gnd.n543 225.874
R13347 gnd.n6464 gnd.n543 225.874
R13348 gnd.n6465 gnd.n6464 225.874
R13349 gnd.n6466 gnd.n6465 225.874
R13350 gnd.n6466 gnd.n537 225.874
R13351 gnd.n6474 gnd.n537 225.874
R13352 gnd.n6475 gnd.n6474 225.874
R13353 gnd.n6476 gnd.n6475 225.874
R13354 gnd.n6476 gnd.n531 225.874
R13355 gnd.n6484 gnd.n531 225.874
R13356 gnd.n6485 gnd.n6484 225.874
R13357 gnd.n6486 gnd.n6485 225.874
R13358 gnd.n6486 gnd.n525 225.874
R13359 gnd.n6495 gnd.n525 225.874
R13360 gnd.n6496 gnd.n6495 225.874
R13361 gnd.n6497 gnd.n6496 225.874
R13362 gnd.n6497 gnd.n520 225.874
R13363 gnd.n2819 gnd.t210 224.174
R13364 gnd.n2312 gnd.t205 224.174
R13365 gnd.n1311 gnd.n1251 199.319
R13366 gnd.n1311 gnd.n1252 199.319
R13367 gnd.n1046 gnd.n1006 199.319
R13368 gnd.n1046 gnd.n1005 199.319
R13369 gnd.n1095 gnd.n1092 186.49
R13370 gnd.n1421 gnd.n1418 186.49
R13371 gnd.n3594 gnd.n3593 185
R13372 gnd.n3592 gnd.n3591 185
R13373 gnd.n3571 gnd.n3570 185
R13374 gnd.n3586 gnd.n3585 185
R13375 gnd.n3584 gnd.n3583 185
R13376 gnd.n3575 gnd.n3574 185
R13377 gnd.n3578 gnd.n3577 185
R13378 gnd.n3562 gnd.n3561 185
R13379 gnd.n3560 gnd.n3559 185
R13380 gnd.n3539 gnd.n3538 185
R13381 gnd.n3554 gnd.n3553 185
R13382 gnd.n3552 gnd.n3551 185
R13383 gnd.n3543 gnd.n3542 185
R13384 gnd.n3546 gnd.n3545 185
R13385 gnd.n3530 gnd.n3529 185
R13386 gnd.n3528 gnd.n3527 185
R13387 gnd.n3507 gnd.n3506 185
R13388 gnd.n3522 gnd.n3521 185
R13389 gnd.n3520 gnd.n3519 185
R13390 gnd.n3511 gnd.n3510 185
R13391 gnd.n3514 gnd.n3513 185
R13392 gnd.n3499 gnd.n3498 185
R13393 gnd.n3497 gnd.n3496 185
R13394 gnd.n3476 gnd.n3475 185
R13395 gnd.n3491 gnd.n3490 185
R13396 gnd.n3489 gnd.n3488 185
R13397 gnd.n3480 gnd.n3479 185
R13398 gnd.n3483 gnd.n3482 185
R13399 gnd.n3467 gnd.n3466 185
R13400 gnd.n3465 gnd.n3464 185
R13401 gnd.n3444 gnd.n3443 185
R13402 gnd.n3459 gnd.n3458 185
R13403 gnd.n3457 gnd.n3456 185
R13404 gnd.n3448 gnd.n3447 185
R13405 gnd.n3451 gnd.n3450 185
R13406 gnd.n3435 gnd.n3434 185
R13407 gnd.n3433 gnd.n3432 185
R13408 gnd.n3412 gnd.n3411 185
R13409 gnd.n3427 gnd.n3426 185
R13410 gnd.n3425 gnd.n3424 185
R13411 gnd.n3416 gnd.n3415 185
R13412 gnd.n3419 gnd.n3418 185
R13413 gnd.n3403 gnd.n3402 185
R13414 gnd.n3401 gnd.n3400 185
R13415 gnd.n3380 gnd.n3379 185
R13416 gnd.n3395 gnd.n3394 185
R13417 gnd.n3393 gnd.n3392 185
R13418 gnd.n3384 gnd.n3383 185
R13419 gnd.n3387 gnd.n3386 185
R13420 gnd.n3372 gnd.n3371 185
R13421 gnd.n3370 gnd.n3369 185
R13422 gnd.n3349 gnd.n3348 185
R13423 gnd.n3364 gnd.n3363 185
R13424 gnd.n3362 gnd.n3361 185
R13425 gnd.n3353 gnd.n3352 185
R13426 gnd.n3356 gnd.n3355 185
R13427 gnd.n2820 gnd.t209 178.987
R13428 gnd.n2313 gnd.t206 178.987
R13429 gnd.n1 gnd.t353 170.774
R13430 gnd.n7 gnd.t183 170.103
R13431 gnd.n6 gnd.t196 170.103
R13432 gnd.n5 gnd.t10 170.103
R13433 gnd.n4 gnd.t349 170.103
R13434 gnd.n3 gnd.t176 170.103
R13435 gnd.n2 gnd.t178 170.103
R13436 gnd.n1 gnd.t191 170.103
R13437 gnd.n5177 gnd.n5176 163.367
R13438 gnd.n5174 gnd.n1430 163.367
R13439 gnd.n5170 gnd.n5169 163.367
R13440 gnd.n5167 gnd.n1433 163.367
R13441 gnd.n5163 gnd.n5162 163.367
R13442 gnd.n5160 gnd.n1436 163.367
R13443 gnd.n5156 gnd.n5155 163.367
R13444 gnd.n5153 gnd.n1439 163.367
R13445 gnd.n5149 gnd.n5148 163.367
R13446 gnd.n5146 gnd.n1442 163.367
R13447 gnd.n5142 gnd.n5141 163.367
R13448 gnd.n5139 gnd.n1445 163.367
R13449 gnd.n5135 gnd.n5134 163.367
R13450 gnd.n5132 gnd.n1448 163.367
R13451 gnd.n5127 gnd.n5126 163.367
R13452 gnd.n5124 gnd.n5122 163.367
R13453 gnd.n5119 gnd.n5118 163.367
R13454 gnd.n5116 gnd.n1454 163.367
R13455 gnd.n5111 gnd.n5110 163.367
R13456 gnd.n5108 gnd.n1459 163.367
R13457 gnd.n5104 gnd.n5103 163.367
R13458 gnd.n5101 gnd.n1462 163.367
R13459 gnd.n5097 gnd.n5096 163.367
R13460 gnd.n5094 gnd.n1465 163.367
R13461 gnd.n5090 gnd.n5089 163.367
R13462 gnd.n5087 gnd.n1468 163.367
R13463 gnd.n5083 gnd.n5082 163.367
R13464 gnd.n5080 gnd.n1471 163.367
R13465 gnd.n5076 gnd.n5075 163.367
R13466 gnd.n5073 gnd.n1474 163.367
R13467 gnd.n5069 gnd.n5068 163.367
R13468 gnd.n5066 gnd.n1477 163.367
R13469 gnd.n1788 gnd.n1111 163.367
R13470 gnd.n1112 gnd.n1111 163.367
R13471 gnd.n1793 gnd.n1112 163.367
R13472 gnd.n4629 gnd.n1793 163.367
R13473 gnd.n4630 gnd.n4629 163.367
R13474 gnd.n4630 gnd.n1719 163.367
R13475 gnd.n4642 gnd.n1719 163.367
R13476 gnd.n4642 gnd.n1720 163.367
R13477 gnd.n1720 gnd.n1715 163.367
R13478 gnd.n4637 gnd.n1715 163.367
R13479 gnd.n4637 gnd.n1707 163.367
R13480 gnd.n4634 gnd.n1707 163.367
R13481 gnd.n4634 gnd.n1700 163.367
R13482 gnd.n4672 gnd.n1700 163.367
R13483 gnd.n4672 gnd.n1697 163.367
R13484 gnd.n4680 gnd.n1697 163.367
R13485 gnd.n4680 gnd.n1691 163.367
R13486 gnd.n4676 gnd.n1691 163.367
R13487 gnd.n4676 gnd.n1682 163.367
R13488 gnd.n1682 gnd.n1673 163.367
R13489 gnd.n4707 gnd.n1673 163.367
R13490 gnd.n4707 gnd.n1670 163.367
R13491 gnd.n4717 gnd.n1670 163.367
R13492 gnd.n4717 gnd.n1671 163.367
R13493 gnd.n1671 gnd.n1664 163.367
R13494 gnd.n4712 gnd.n1664 163.367
R13495 gnd.n4712 gnd.n1654 163.367
R13496 gnd.n1654 gnd.n1648 163.367
R13497 gnd.n4743 gnd.n1648 163.367
R13498 gnd.n4743 gnd.n1646 163.367
R13499 gnd.n4749 gnd.n1646 163.367
R13500 gnd.n4749 gnd.n1636 163.367
R13501 gnd.n1636 gnd.n1630 163.367
R13502 gnd.n4771 gnd.n1630 163.367
R13503 gnd.n4772 gnd.n4771 163.367
R13504 gnd.n4772 gnd.n1627 163.367
R13505 gnd.n4792 gnd.n1627 163.367
R13506 gnd.n4792 gnd.n1619 163.367
R13507 gnd.n4788 gnd.n1619 163.367
R13508 gnd.n4788 gnd.n4787 163.367
R13509 gnd.n4787 gnd.n4786 163.367
R13510 gnd.n4786 gnd.n4776 163.367
R13511 gnd.n4776 gnd.n1601 163.367
R13512 gnd.n4781 gnd.n1601 163.367
R13513 gnd.n4781 gnd.n1595 163.367
R13514 gnd.n4778 gnd.n1595 163.367
R13515 gnd.n4778 gnd.n1584 163.367
R13516 gnd.n1584 gnd.n1576 163.367
R13517 gnd.n4866 gnd.n1576 163.367
R13518 gnd.n4866 gnd.n1573 163.367
R13519 gnd.n4904 gnd.n1573 163.367
R13520 gnd.n4904 gnd.n1574 163.367
R13521 gnd.n1574 gnd.n1565 163.367
R13522 gnd.n4899 gnd.n1565 163.367
R13523 gnd.n4899 gnd.n4897 163.367
R13524 gnd.n4897 gnd.n4896 163.367
R13525 gnd.n4896 gnd.n4872 163.367
R13526 gnd.n4872 gnd.n1548 163.367
R13527 gnd.n4891 gnd.n1548 163.367
R13528 gnd.n4891 gnd.n1541 163.367
R13529 gnd.n4888 gnd.n1541 163.367
R13530 gnd.n4888 gnd.n4887 163.367
R13531 gnd.n4887 gnd.n4886 163.367
R13532 gnd.n4886 gnd.n4876 163.367
R13533 gnd.n4876 gnd.n1525 163.367
R13534 gnd.n4881 gnd.n1525 163.367
R13535 gnd.n4881 gnd.n1520 163.367
R13536 gnd.n4878 gnd.n1520 163.367
R13537 gnd.n4878 gnd.n1510 163.367
R13538 gnd.n1510 gnd.n1504 163.367
R13539 gnd.n5022 gnd.n1504 163.367
R13540 gnd.n5022 gnd.n1501 163.367
R13541 gnd.n5033 gnd.n1501 163.367
R13542 gnd.n5033 gnd.n1502 163.367
R13543 gnd.n1502 gnd.n1495 163.367
R13544 gnd.n5028 gnd.n1495 163.367
R13545 gnd.n5028 gnd.n1484 163.367
R13546 gnd.n1484 gnd.n1479 163.367
R13547 gnd.n5057 gnd.n1479 163.367
R13548 gnd.n5058 gnd.n5057 163.367
R13549 gnd.n5058 gnd.n1404 163.367
R13550 gnd.n1086 gnd.n1085 163.367
R13551 gnd.n5890 gnd.n1085 163.367
R13552 gnd.n5888 gnd.n5887 163.367
R13553 gnd.n5884 gnd.n5883 163.367
R13554 gnd.n5880 gnd.n5879 163.367
R13555 gnd.n5876 gnd.n5875 163.367
R13556 gnd.n5872 gnd.n5871 163.367
R13557 gnd.n5868 gnd.n5867 163.367
R13558 gnd.n5864 gnd.n5863 163.367
R13559 gnd.n5860 gnd.n5859 163.367
R13560 gnd.n5856 gnd.n5855 163.367
R13561 gnd.n5852 gnd.n5851 163.367
R13562 gnd.n5848 gnd.n5847 163.367
R13563 gnd.n5844 gnd.n5843 163.367
R13564 gnd.n5840 gnd.n5839 163.367
R13565 gnd.n5836 gnd.n5835 163.367
R13566 gnd.n5899 gnd.n1051 163.367
R13567 gnd.n1726 gnd.n1725 163.367
R13568 gnd.n1731 gnd.n1730 163.367
R13569 gnd.n1735 gnd.n1734 163.367
R13570 gnd.n1739 gnd.n1738 163.367
R13571 gnd.n1743 gnd.n1742 163.367
R13572 gnd.n1747 gnd.n1746 163.367
R13573 gnd.n1751 gnd.n1750 163.367
R13574 gnd.n1755 gnd.n1754 163.367
R13575 gnd.n1759 gnd.n1758 163.367
R13576 gnd.n1763 gnd.n1762 163.367
R13577 gnd.n1767 gnd.n1766 163.367
R13578 gnd.n1771 gnd.n1770 163.367
R13579 gnd.n1775 gnd.n1774 163.367
R13580 gnd.n1779 gnd.n1778 163.367
R13581 gnd.n1783 gnd.n1782 163.367
R13582 gnd.n5828 gnd.n1087 163.367
R13583 gnd.n5828 gnd.n1109 163.367
R13584 gnd.n4622 gnd.n1109 163.367
R13585 gnd.n4627 gnd.n4622 163.367
R13586 gnd.n4627 gnd.n4623 163.367
R13587 gnd.n4623 gnd.n1718 163.367
R13588 gnd.n4644 gnd.n1718 163.367
R13589 gnd.n4644 gnd.n1716 163.367
R13590 gnd.n4648 gnd.n1716 163.367
R13591 gnd.n4648 gnd.n1705 163.367
R13592 gnd.n4665 gnd.n1705 163.367
R13593 gnd.n4665 gnd.n1703 163.367
R13594 gnd.n4669 gnd.n1703 163.367
R13595 gnd.n4669 gnd.n1695 163.367
R13596 gnd.n4684 gnd.n1695 163.367
R13597 gnd.n4684 gnd.n1693 163.367
R13598 gnd.n4688 gnd.n1693 163.367
R13599 gnd.n4688 gnd.n1679 163.367
R13600 gnd.n4701 gnd.n1679 163.367
R13601 gnd.n4701 gnd.n1677 163.367
R13602 gnd.n4705 gnd.n1677 163.367
R13603 gnd.n4705 gnd.n1668 163.367
R13604 gnd.n4719 gnd.n1668 163.367
R13605 gnd.n4719 gnd.n1666 163.367
R13606 gnd.n4723 gnd.n1666 163.367
R13607 gnd.n4723 gnd.n1653 163.367
R13608 gnd.n4736 gnd.n1653 163.367
R13609 gnd.n4736 gnd.n1650 163.367
R13610 gnd.n4741 gnd.n1650 163.367
R13611 gnd.n4741 gnd.n1651 163.367
R13612 gnd.n1651 gnd.n1634 163.367
R13613 gnd.n4765 gnd.n1634 163.367
R13614 gnd.n4765 gnd.n1632 163.367
R13615 gnd.n4769 gnd.n1632 163.367
R13616 gnd.n4769 gnd.n1625 163.367
R13617 gnd.n4797 gnd.n1625 163.367
R13618 gnd.n4797 gnd.n1622 163.367
R13619 gnd.n4806 gnd.n1622 163.367
R13620 gnd.n4806 gnd.n1623 163.367
R13621 gnd.n4802 gnd.n1623 163.367
R13622 gnd.n4802 gnd.n4801 163.367
R13623 gnd.n4801 gnd.n1599 163.367
R13624 gnd.n4842 gnd.n1599 163.367
R13625 gnd.n4842 gnd.n1597 163.367
R13626 gnd.n4846 gnd.n1597 163.367
R13627 gnd.n4846 gnd.n1582 163.367
R13628 gnd.n4860 gnd.n1582 163.367
R13629 gnd.n4860 gnd.n1580 163.367
R13630 gnd.n4864 gnd.n1580 163.367
R13631 gnd.n4864 gnd.n1571 163.367
R13632 gnd.n4906 gnd.n1571 163.367
R13633 gnd.n4906 gnd.n1568 163.367
R13634 gnd.n4915 gnd.n1568 163.367
R13635 gnd.n4915 gnd.n1569 163.367
R13636 gnd.n4911 gnd.n1569 163.367
R13637 gnd.n4911 gnd.n4910 163.367
R13638 gnd.n4910 gnd.n1547 163.367
R13639 gnd.n4938 gnd.n1547 163.367
R13640 gnd.n4938 gnd.n1544 163.367
R13641 gnd.n4947 gnd.n1544 163.367
R13642 gnd.n4947 gnd.n1545 163.367
R13643 gnd.n4943 gnd.n1545 163.367
R13644 gnd.n4943 gnd.n4942 163.367
R13645 gnd.n4942 gnd.n1524 163.367
R13646 gnd.n4998 gnd.n1524 163.367
R13647 gnd.n4998 gnd.n1522 163.367
R13648 gnd.n5002 gnd.n1522 163.367
R13649 gnd.n5002 gnd.n1508 163.367
R13650 gnd.n5016 gnd.n1508 163.367
R13651 gnd.n5016 gnd.n1506 163.367
R13652 gnd.n5020 gnd.n1506 163.367
R13653 gnd.n5020 gnd.n1499 163.367
R13654 gnd.n5035 gnd.n1499 163.367
R13655 gnd.n5035 gnd.n1497 163.367
R13656 gnd.n5039 gnd.n1497 163.367
R13657 gnd.n5039 gnd.n1483 163.367
R13658 gnd.n5051 gnd.n1483 163.367
R13659 gnd.n5051 gnd.n1481 163.367
R13660 gnd.n5055 gnd.n1481 163.367
R13661 gnd.n5055 gnd.n1406 163.367
R13662 gnd.n5182 gnd.n1406 163.367
R13663 gnd.n1427 gnd.n1426 156.462
R13664 gnd.n3534 gnd.n3502 153.042
R13665 gnd.n3598 gnd.n3597 152.079
R13666 gnd.n3566 gnd.n3565 152.079
R13667 gnd.n3534 gnd.n3533 152.079
R13668 gnd.n1100 gnd.n1099 152
R13669 gnd.n1101 gnd.n1090 152
R13670 gnd.n1103 gnd.n1102 152
R13671 gnd.n1105 gnd.n1088 152
R13672 gnd.n1107 gnd.n1106 152
R13673 gnd.n1425 gnd.n1409 152
R13674 gnd.n1417 gnd.n1410 152
R13675 gnd.n1416 gnd.n1415 152
R13676 gnd.n1414 gnd.n1411 152
R13677 gnd.n1412 gnd.t253 150.546
R13678 gnd.t1 gnd.n3576 147.661
R13679 gnd.t347 gnd.n3544 147.661
R13680 gnd.t5 gnd.n3512 147.661
R13681 gnd.t3 gnd.n3481 147.661
R13682 gnd.t7 gnd.n3449 147.661
R13683 gnd.t359 gnd.n3417 147.661
R13684 gnd.t187 gnd.n3385 147.661
R13685 gnd.t357 gnd.n3354 147.661
R13686 gnd.n5121 gnd.n5120 143.351
R13687 gnd.n1067 gnd.n1050 143.351
R13688 gnd.n5898 gnd.n1050 143.351
R13689 gnd.n1097 gnd.t304 130.484
R13690 gnd.n1106 gnd.t211 126.766
R13691 gnd.n1104 gnd.t275 126.766
R13692 gnd.n1090 gnd.t229 126.766
R13693 gnd.n1098 gnd.t250 126.766
R13694 gnd.n1413 gnd.t316 126.766
R13695 gnd.n1415 gnd.t266 126.766
R13696 gnd.n1424 gnd.t214 126.766
R13697 gnd.n1426 gnd.t288 126.766
R13698 gnd.n5655 gnd.n1310 108.609
R13699 gnd.n5901 gnd.n5900 108.609
R13700 gnd.n3593 gnd.n3592 104.615
R13701 gnd.n3592 gnd.n3570 104.615
R13702 gnd.n3585 gnd.n3570 104.615
R13703 gnd.n3585 gnd.n3584 104.615
R13704 gnd.n3584 gnd.n3574 104.615
R13705 gnd.n3577 gnd.n3574 104.615
R13706 gnd.n3561 gnd.n3560 104.615
R13707 gnd.n3560 gnd.n3538 104.615
R13708 gnd.n3553 gnd.n3538 104.615
R13709 gnd.n3553 gnd.n3552 104.615
R13710 gnd.n3552 gnd.n3542 104.615
R13711 gnd.n3545 gnd.n3542 104.615
R13712 gnd.n3529 gnd.n3528 104.615
R13713 gnd.n3528 gnd.n3506 104.615
R13714 gnd.n3521 gnd.n3506 104.615
R13715 gnd.n3521 gnd.n3520 104.615
R13716 gnd.n3520 gnd.n3510 104.615
R13717 gnd.n3513 gnd.n3510 104.615
R13718 gnd.n3498 gnd.n3497 104.615
R13719 gnd.n3497 gnd.n3475 104.615
R13720 gnd.n3490 gnd.n3475 104.615
R13721 gnd.n3490 gnd.n3489 104.615
R13722 gnd.n3489 gnd.n3479 104.615
R13723 gnd.n3482 gnd.n3479 104.615
R13724 gnd.n3466 gnd.n3465 104.615
R13725 gnd.n3465 gnd.n3443 104.615
R13726 gnd.n3458 gnd.n3443 104.615
R13727 gnd.n3458 gnd.n3457 104.615
R13728 gnd.n3457 gnd.n3447 104.615
R13729 gnd.n3450 gnd.n3447 104.615
R13730 gnd.n3434 gnd.n3433 104.615
R13731 gnd.n3433 gnd.n3411 104.615
R13732 gnd.n3426 gnd.n3411 104.615
R13733 gnd.n3426 gnd.n3425 104.615
R13734 gnd.n3425 gnd.n3415 104.615
R13735 gnd.n3418 gnd.n3415 104.615
R13736 gnd.n3402 gnd.n3401 104.615
R13737 gnd.n3401 gnd.n3379 104.615
R13738 gnd.n3394 gnd.n3379 104.615
R13739 gnd.n3394 gnd.n3393 104.615
R13740 gnd.n3393 gnd.n3383 104.615
R13741 gnd.n3386 gnd.n3383 104.615
R13742 gnd.n3371 gnd.n3370 104.615
R13743 gnd.n3370 gnd.n3348 104.615
R13744 gnd.n3363 gnd.n3348 104.615
R13745 gnd.n3363 gnd.n3362 104.615
R13746 gnd.n3362 gnd.n3352 104.615
R13747 gnd.n3355 gnd.n3352 104.615
R13748 gnd.n2745 gnd.t281 100.632
R13749 gnd.n2286 gnd.t302 100.632
R13750 gnd.n7110 gnd.n7109 99.6594
R13751 gnd.n7105 gnd.n248 99.6594
R13752 gnd.n7101 gnd.n247 99.6594
R13753 gnd.n7097 gnd.n246 99.6594
R13754 gnd.n7093 gnd.n245 99.6594
R13755 gnd.n7089 gnd.n244 99.6594
R13756 gnd.n7085 gnd.n243 99.6594
R13757 gnd.n7081 gnd.n242 99.6594
R13758 gnd.n7074 gnd.n241 99.6594
R13759 gnd.n7070 gnd.n240 99.6594
R13760 gnd.n7066 gnd.n239 99.6594
R13761 gnd.n7062 gnd.n238 99.6594
R13762 gnd.n7058 gnd.n237 99.6594
R13763 gnd.n7054 gnd.n236 99.6594
R13764 gnd.n7050 gnd.n235 99.6594
R13765 gnd.n7046 gnd.n234 99.6594
R13766 gnd.n7042 gnd.n233 99.6594
R13767 gnd.n7038 gnd.n232 99.6594
R13768 gnd.n7030 gnd.n231 99.6594
R13769 gnd.n7028 gnd.n230 99.6594
R13770 gnd.n7024 gnd.n229 99.6594
R13771 gnd.n7020 gnd.n228 99.6594
R13772 gnd.n7016 gnd.n227 99.6594
R13773 gnd.n7012 gnd.n226 99.6594
R13774 gnd.n7008 gnd.n225 99.6594
R13775 gnd.n7004 gnd.n224 99.6594
R13776 gnd.n7000 gnd.n223 99.6594
R13777 gnd.n6996 gnd.n222 99.6594
R13778 gnd.n6987 gnd.n221 99.6594
R13779 gnd.n5707 gnd.n5706 99.6594
R13780 gnd.n5701 gnd.n1240 99.6594
R13781 gnd.n5698 gnd.n1241 99.6594
R13782 gnd.n5694 gnd.n1242 99.6594
R13783 gnd.n5690 gnd.n1243 99.6594
R13784 gnd.n5686 gnd.n1244 99.6594
R13785 gnd.n5682 gnd.n1245 99.6594
R13786 gnd.n5678 gnd.n1246 99.6594
R13787 gnd.n5674 gnd.n1247 99.6594
R13788 gnd.n5669 gnd.n1248 99.6594
R13789 gnd.n5665 gnd.n1249 99.6594
R13790 gnd.n5661 gnd.n1250 99.6594
R13791 gnd.n5657 gnd.n1251 99.6594
R13792 gnd.n5652 gnd.n1253 99.6594
R13793 gnd.n5648 gnd.n1254 99.6594
R13794 gnd.n5644 gnd.n1255 99.6594
R13795 gnd.n5640 gnd.n1256 99.6594
R13796 gnd.n5636 gnd.n1257 99.6594
R13797 gnd.n5632 gnd.n1258 99.6594
R13798 gnd.n5628 gnd.n1259 99.6594
R13799 gnd.n5624 gnd.n1260 99.6594
R13800 gnd.n5620 gnd.n1261 99.6594
R13801 gnd.n5616 gnd.n1262 99.6594
R13802 gnd.n5612 gnd.n1263 99.6594
R13803 gnd.n5608 gnd.n1264 99.6594
R13804 gnd.n5604 gnd.n1265 99.6594
R13805 gnd.n5600 gnd.n1266 99.6594
R13806 gnd.n5596 gnd.n1267 99.6594
R13807 gnd.n5950 gnd.n5949 99.6594
R13808 gnd.n5945 gnd.n1017 99.6594
R13809 gnd.n5941 gnd.n1016 99.6594
R13810 gnd.n5937 gnd.n1015 99.6594
R13811 gnd.n5933 gnd.n1014 99.6594
R13812 gnd.n5929 gnd.n1013 99.6594
R13813 gnd.n5925 gnd.n1012 99.6594
R13814 gnd.n5921 gnd.n1011 99.6594
R13815 gnd.n5916 gnd.n1010 99.6594
R13816 gnd.n5912 gnd.n1009 99.6594
R13817 gnd.n5908 gnd.n1008 99.6594
R13818 gnd.n5904 gnd.n1007 99.6594
R13819 gnd.n1977 gnd.n1005 99.6594
R13820 gnd.n1981 gnd.n1004 99.6594
R13821 gnd.n1987 gnd.n1003 99.6594
R13822 gnd.n1991 gnd.n1002 99.6594
R13823 gnd.n1996 gnd.n1001 99.6594
R13824 gnd.n2000 gnd.n1000 99.6594
R13825 gnd.n2006 gnd.n999 99.6594
R13826 gnd.n2010 gnd.n998 99.6594
R13827 gnd.n2016 gnd.n997 99.6594
R13828 gnd.n2020 gnd.n996 99.6594
R13829 gnd.n2026 gnd.n995 99.6594
R13830 gnd.n2030 gnd.n994 99.6594
R13831 gnd.n2036 gnd.n993 99.6594
R13832 gnd.n2040 gnd.n992 99.6594
R13833 gnd.n2045 gnd.n991 99.6594
R13834 gnd.n2048 gnd.n990 99.6594
R13835 gnd.n4038 gnd.n4037 99.6594
R13836 gnd.n4032 gnd.n3726 99.6594
R13837 gnd.n4029 gnd.n3727 99.6594
R13838 gnd.n4025 gnd.n3728 99.6594
R13839 gnd.n4021 gnd.n3729 99.6594
R13840 gnd.n4017 gnd.n3730 99.6594
R13841 gnd.n4013 gnd.n3731 99.6594
R13842 gnd.n4009 gnd.n3732 99.6594
R13843 gnd.n4005 gnd.n3733 99.6594
R13844 gnd.n4000 gnd.n3734 99.6594
R13845 gnd.n3996 gnd.n3735 99.6594
R13846 gnd.n3992 gnd.n3736 99.6594
R13847 gnd.n3988 gnd.n3737 99.6594
R13848 gnd.n3984 gnd.n3738 99.6594
R13849 gnd.n3980 gnd.n3739 99.6594
R13850 gnd.n3976 gnd.n3740 99.6594
R13851 gnd.n3972 gnd.n3741 99.6594
R13852 gnd.n3968 gnd.n3742 99.6594
R13853 gnd.n3964 gnd.n3743 99.6594
R13854 gnd.n3960 gnd.n3744 99.6594
R13855 gnd.n3956 gnd.n3745 99.6594
R13856 gnd.n3952 gnd.n3746 99.6594
R13857 gnd.n3948 gnd.n3747 99.6594
R13858 gnd.n3944 gnd.n3748 99.6594
R13859 gnd.n3940 gnd.n3749 99.6594
R13860 gnd.n3936 gnd.n3750 99.6594
R13861 gnd.n3932 gnd.n3751 99.6594
R13862 gnd.n3928 gnd.n3752 99.6594
R13863 gnd.n4040 gnd.n2246 99.6594
R13864 gnd.n3716 gnd.n2269 99.6594
R13865 gnd.n3714 gnd.n2268 99.6594
R13866 gnd.n3710 gnd.n2267 99.6594
R13867 gnd.n3706 gnd.n2266 99.6594
R13868 gnd.n3702 gnd.n2265 99.6594
R13869 gnd.n3698 gnd.n2264 99.6594
R13870 gnd.n3694 gnd.n2263 99.6594
R13871 gnd.n3626 gnd.n2262 99.6594
R13872 gnd.n2957 gnd.n2688 99.6594
R13873 gnd.n2714 gnd.n2695 99.6594
R13874 gnd.n2716 gnd.n2696 99.6594
R13875 gnd.n2724 gnd.n2697 99.6594
R13876 gnd.n2726 gnd.n2698 99.6594
R13877 gnd.n2734 gnd.n2699 99.6594
R13878 gnd.n2736 gnd.n2700 99.6594
R13879 gnd.n2744 gnd.n2701 99.6594
R13880 gnd.n6911 gnd.n212 99.6594
R13881 gnd.n6915 gnd.n213 99.6594
R13882 gnd.n6921 gnd.n214 99.6594
R13883 gnd.n6925 gnd.n215 99.6594
R13884 gnd.n6931 gnd.n216 99.6594
R13885 gnd.n6935 gnd.n217 99.6594
R13886 gnd.n6941 gnd.n218 99.6594
R13887 gnd.n6945 gnd.n219 99.6594
R13888 gnd.n6951 gnd.n220 99.6594
R13889 gnd.n5477 gnd.n1268 99.6594
R13890 gnd.n5480 gnd.n1269 99.6594
R13891 gnd.n5488 gnd.n1270 99.6594
R13892 gnd.n5490 gnd.n1271 99.6594
R13893 gnd.n5500 gnd.n1272 99.6594
R13894 gnd.n5508 gnd.n1273 99.6594
R13895 gnd.n5510 gnd.n1274 99.6594
R13896 gnd.n5520 gnd.n1275 99.6594
R13897 gnd.n5530 gnd.n1276 99.6594
R13898 gnd.n3684 gnd.n2249 99.6594
R13899 gnd.n3680 gnd.n2250 99.6594
R13900 gnd.n3676 gnd.n2251 99.6594
R13901 gnd.n3672 gnd.n2252 99.6594
R13902 gnd.n3668 gnd.n2253 99.6594
R13903 gnd.n3664 gnd.n2254 99.6594
R13904 gnd.n3660 gnd.n2255 99.6594
R13905 gnd.n3656 gnd.n2256 99.6594
R13906 gnd.n3652 gnd.n2257 99.6594
R13907 gnd.n3648 gnd.n2258 99.6594
R13908 gnd.n3644 gnd.n2259 99.6594
R13909 gnd.n3640 gnd.n2260 99.6594
R13910 gnd.n3636 gnd.n2261 99.6594
R13911 gnd.n2872 gnd.n2871 99.6594
R13912 gnd.n2866 gnd.n2783 99.6594
R13913 gnd.n2863 gnd.n2784 99.6594
R13914 gnd.n2859 gnd.n2785 99.6594
R13915 gnd.n2855 gnd.n2786 99.6594
R13916 gnd.n2851 gnd.n2787 99.6594
R13917 gnd.n2847 gnd.n2788 99.6594
R13918 gnd.n2843 gnd.n2789 99.6594
R13919 gnd.n2839 gnd.n2790 99.6594
R13920 gnd.n2835 gnd.n2791 99.6594
R13921 gnd.n2831 gnd.n2792 99.6594
R13922 gnd.n2827 gnd.n2793 99.6594
R13923 gnd.n2874 gnd.n2782 99.6594
R13924 gnd.n1906 gnd.n980 99.6594
R13925 gnd.n4401 gnd.n981 99.6594
R13926 gnd.n4412 gnd.n982 99.6594
R13927 gnd.n1894 gnd.n983 99.6594
R13928 gnd.n4425 gnd.n984 99.6594
R13929 gnd.n4436 gnd.n985 99.6594
R13930 gnd.n1882 gnd.n986 99.6594
R13931 gnd.n4450 gnd.n987 99.6594
R13932 gnd.n4470 gnd.n988 99.6594
R13933 gnd.n3918 gnd.n3753 99.6594
R13934 gnd.n3915 gnd.n3754 99.6594
R13935 gnd.n3911 gnd.n3755 99.6594
R13936 gnd.n3907 gnd.n3756 99.6594
R13937 gnd.n3903 gnd.n3757 99.6594
R13938 gnd.n3899 gnd.n3758 99.6594
R13939 gnd.n3895 gnd.n3759 99.6594
R13940 gnd.n3891 gnd.n3760 99.6594
R13941 gnd.n3887 gnd.n3761 99.6594
R13942 gnd.n3916 gnd.n3753 99.6594
R13943 gnd.n3912 gnd.n3754 99.6594
R13944 gnd.n3908 gnd.n3755 99.6594
R13945 gnd.n3904 gnd.n3756 99.6594
R13946 gnd.n3900 gnd.n3757 99.6594
R13947 gnd.n3896 gnd.n3758 99.6594
R13948 gnd.n3892 gnd.n3759 99.6594
R13949 gnd.n3888 gnd.n3760 99.6594
R13950 gnd.n3843 gnd.n3761 99.6594
R13951 gnd.n4449 gnd.n988 99.6594
R13952 gnd.n1883 gnd.n987 99.6594
R13953 gnd.n4437 gnd.n986 99.6594
R13954 gnd.n4424 gnd.n985 99.6594
R13955 gnd.n1895 gnd.n984 99.6594
R13956 gnd.n4413 gnd.n983 99.6594
R13957 gnd.n4400 gnd.n982 99.6594
R13958 gnd.n1907 gnd.n981 99.6594
R13959 gnd.n4389 gnd.n980 99.6594
R13960 gnd.n2872 gnd.n2795 99.6594
R13961 gnd.n2864 gnd.n2783 99.6594
R13962 gnd.n2860 gnd.n2784 99.6594
R13963 gnd.n2856 gnd.n2785 99.6594
R13964 gnd.n2852 gnd.n2786 99.6594
R13965 gnd.n2848 gnd.n2787 99.6594
R13966 gnd.n2844 gnd.n2788 99.6594
R13967 gnd.n2840 gnd.n2789 99.6594
R13968 gnd.n2836 gnd.n2790 99.6594
R13969 gnd.n2832 gnd.n2791 99.6594
R13970 gnd.n2828 gnd.n2792 99.6594
R13971 gnd.n2824 gnd.n2793 99.6594
R13972 gnd.n2875 gnd.n2874 99.6594
R13973 gnd.n3639 gnd.n2261 99.6594
R13974 gnd.n3643 gnd.n2260 99.6594
R13975 gnd.n3647 gnd.n2259 99.6594
R13976 gnd.n3651 gnd.n2258 99.6594
R13977 gnd.n3655 gnd.n2257 99.6594
R13978 gnd.n3659 gnd.n2256 99.6594
R13979 gnd.n3663 gnd.n2255 99.6594
R13980 gnd.n3667 gnd.n2254 99.6594
R13981 gnd.n3671 gnd.n2253 99.6594
R13982 gnd.n3675 gnd.n2252 99.6594
R13983 gnd.n3679 gnd.n2251 99.6594
R13984 gnd.n3683 gnd.n2250 99.6594
R13985 gnd.n2290 gnd.n2249 99.6594
R13986 gnd.n5479 gnd.n1268 99.6594
R13987 gnd.n5487 gnd.n1269 99.6594
R13988 gnd.n5489 gnd.n1270 99.6594
R13989 gnd.n5499 gnd.n1271 99.6594
R13990 gnd.n5507 gnd.n1272 99.6594
R13991 gnd.n5509 gnd.n1273 99.6594
R13992 gnd.n5519 gnd.n1274 99.6594
R13993 gnd.n5529 gnd.n1275 99.6594
R13994 gnd.n5540 gnd.n1276 99.6594
R13995 gnd.n6944 gnd.n220 99.6594
R13996 gnd.n6942 gnd.n219 99.6594
R13997 gnd.n6934 gnd.n218 99.6594
R13998 gnd.n6932 gnd.n217 99.6594
R13999 gnd.n6924 gnd.n216 99.6594
R14000 gnd.n6922 gnd.n215 99.6594
R14001 gnd.n6914 gnd.n214 99.6594
R14002 gnd.n6912 gnd.n213 99.6594
R14003 gnd.n6906 gnd.n212 99.6594
R14004 gnd.n2958 gnd.n2957 99.6594
R14005 gnd.n2717 gnd.n2695 99.6594
R14006 gnd.n2723 gnd.n2696 99.6594
R14007 gnd.n2727 gnd.n2697 99.6594
R14008 gnd.n2733 gnd.n2698 99.6594
R14009 gnd.n2737 gnd.n2699 99.6594
R14010 gnd.n2743 gnd.n2700 99.6594
R14011 gnd.n2701 gnd.n2685 99.6594
R14012 gnd.n3693 gnd.n2262 99.6594
R14013 gnd.n3697 gnd.n2263 99.6594
R14014 gnd.n3701 gnd.n2264 99.6594
R14015 gnd.n3705 gnd.n2265 99.6594
R14016 gnd.n3709 gnd.n2266 99.6594
R14017 gnd.n3713 gnd.n2267 99.6594
R14018 gnd.n3717 gnd.n2268 99.6594
R14019 gnd.n2271 gnd.n2269 99.6594
R14020 gnd.n4038 gnd.n3764 99.6594
R14021 gnd.n4030 gnd.n3726 99.6594
R14022 gnd.n4026 gnd.n3727 99.6594
R14023 gnd.n4022 gnd.n3728 99.6594
R14024 gnd.n4018 gnd.n3729 99.6594
R14025 gnd.n4014 gnd.n3730 99.6594
R14026 gnd.n4010 gnd.n3731 99.6594
R14027 gnd.n4006 gnd.n3732 99.6594
R14028 gnd.n4001 gnd.n3733 99.6594
R14029 gnd.n3997 gnd.n3734 99.6594
R14030 gnd.n3993 gnd.n3735 99.6594
R14031 gnd.n3989 gnd.n3736 99.6594
R14032 gnd.n3985 gnd.n3737 99.6594
R14033 gnd.n3981 gnd.n3738 99.6594
R14034 gnd.n3977 gnd.n3739 99.6594
R14035 gnd.n3973 gnd.n3740 99.6594
R14036 gnd.n3969 gnd.n3741 99.6594
R14037 gnd.n3965 gnd.n3742 99.6594
R14038 gnd.n3961 gnd.n3743 99.6594
R14039 gnd.n3957 gnd.n3744 99.6594
R14040 gnd.n3953 gnd.n3745 99.6594
R14041 gnd.n3949 gnd.n3746 99.6594
R14042 gnd.n3945 gnd.n3747 99.6594
R14043 gnd.n3941 gnd.n3748 99.6594
R14044 gnd.n3937 gnd.n3749 99.6594
R14045 gnd.n3933 gnd.n3750 99.6594
R14046 gnd.n3929 gnd.n3751 99.6594
R14047 gnd.n3925 gnd.n3752 99.6594
R14048 gnd.n4041 gnd.n4040 99.6594
R14049 gnd.n1958 gnd.n990 99.6594
R14050 gnd.n2039 gnd.n991 99.6594
R14051 gnd.n2037 gnd.n992 99.6594
R14052 gnd.n2029 gnd.n993 99.6594
R14053 gnd.n2027 gnd.n994 99.6594
R14054 gnd.n2019 gnd.n995 99.6594
R14055 gnd.n2017 gnd.n996 99.6594
R14056 gnd.n2009 gnd.n997 99.6594
R14057 gnd.n2007 gnd.n998 99.6594
R14058 gnd.n1999 gnd.n999 99.6594
R14059 gnd.n1971 gnd.n1000 99.6594
R14060 gnd.n1990 gnd.n1001 99.6594
R14061 gnd.n1988 gnd.n1002 99.6594
R14062 gnd.n1980 gnd.n1003 99.6594
R14063 gnd.n1978 gnd.n1004 99.6594
R14064 gnd.n5903 gnd.n1006 99.6594
R14065 gnd.n5907 gnd.n1007 99.6594
R14066 gnd.n5911 gnd.n1008 99.6594
R14067 gnd.n5915 gnd.n1009 99.6594
R14068 gnd.n5920 gnd.n1010 99.6594
R14069 gnd.n5924 gnd.n1011 99.6594
R14070 gnd.n5928 gnd.n1012 99.6594
R14071 gnd.n5932 gnd.n1013 99.6594
R14072 gnd.n5936 gnd.n1014 99.6594
R14073 gnd.n5940 gnd.n1015 99.6594
R14074 gnd.n5944 gnd.n1016 99.6594
R14075 gnd.n1018 gnd.n1017 99.6594
R14076 gnd.n5950 gnd.n977 99.6594
R14077 gnd.n5707 gnd.n1280 99.6594
R14078 gnd.n5699 gnd.n1240 99.6594
R14079 gnd.n5695 gnd.n1241 99.6594
R14080 gnd.n5691 gnd.n1242 99.6594
R14081 gnd.n5687 gnd.n1243 99.6594
R14082 gnd.n5683 gnd.n1244 99.6594
R14083 gnd.n5679 gnd.n1245 99.6594
R14084 gnd.n5675 gnd.n1246 99.6594
R14085 gnd.n5670 gnd.n1247 99.6594
R14086 gnd.n5666 gnd.n1248 99.6594
R14087 gnd.n5662 gnd.n1249 99.6594
R14088 gnd.n5658 gnd.n1250 99.6594
R14089 gnd.n5653 gnd.n1252 99.6594
R14090 gnd.n5649 gnd.n1253 99.6594
R14091 gnd.n5645 gnd.n1254 99.6594
R14092 gnd.n5641 gnd.n1255 99.6594
R14093 gnd.n5637 gnd.n1256 99.6594
R14094 gnd.n5633 gnd.n1257 99.6594
R14095 gnd.n5629 gnd.n1258 99.6594
R14096 gnd.n5625 gnd.n1259 99.6594
R14097 gnd.n5621 gnd.n1260 99.6594
R14098 gnd.n5617 gnd.n1261 99.6594
R14099 gnd.n5613 gnd.n1262 99.6594
R14100 gnd.n5609 gnd.n1263 99.6594
R14101 gnd.n5605 gnd.n1264 99.6594
R14102 gnd.n5601 gnd.n1265 99.6594
R14103 gnd.n5597 gnd.n1266 99.6594
R14104 gnd.n5271 gnd.n1267 99.6594
R14105 gnd.n6995 gnd.n221 99.6594
R14106 gnd.n6999 gnd.n222 99.6594
R14107 gnd.n7003 gnd.n223 99.6594
R14108 gnd.n7007 gnd.n224 99.6594
R14109 gnd.n7011 gnd.n225 99.6594
R14110 gnd.n7015 gnd.n226 99.6594
R14111 gnd.n7019 gnd.n227 99.6594
R14112 gnd.n7023 gnd.n228 99.6594
R14113 gnd.n7027 gnd.n229 99.6594
R14114 gnd.n7031 gnd.n230 99.6594
R14115 gnd.n7037 gnd.n231 99.6594
R14116 gnd.n7041 gnd.n232 99.6594
R14117 gnd.n7045 gnd.n233 99.6594
R14118 gnd.n7049 gnd.n234 99.6594
R14119 gnd.n7053 gnd.n235 99.6594
R14120 gnd.n7057 gnd.n236 99.6594
R14121 gnd.n7061 gnd.n237 99.6594
R14122 gnd.n7065 gnd.n238 99.6594
R14123 gnd.n7069 gnd.n239 99.6594
R14124 gnd.n7073 gnd.n240 99.6594
R14125 gnd.n7080 gnd.n241 99.6594
R14126 gnd.n7084 gnd.n242 99.6594
R14127 gnd.n7088 gnd.n243 99.6594
R14128 gnd.n7092 gnd.n244 99.6594
R14129 gnd.n7096 gnd.n245 99.6594
R14130 gnd.n7100 gnd.n246 99.6594
R14131 gnd.n7104 gnd.n247 99.6594
R14132 gnd.n249 gnd.n248 99.6594
R14133 gnd.n7110 gnd.n210 99.6594
R14134 gnd.n1943 gnd.n1864 99.6594
R14135 gnd.n1920 gnd.n1865 99.6594
R14136 gnd.n1951 gnd.n1866 99.6594
R14137 gnd.n1916 gnd.n1867 99.6594
R14138 gnd.n4384 gnd.n1868 99.6594
R14139 gnd.n1911 gnd.n1869 99.6594
R14140 gnd.n4394 gnd.n1870 99.6594
R14141 gnd.n4407 gnd.n1871 99.6594
R14142 gnd.n1899 gnd.n1872 99.6594
R14143 gnd.n4418 gnd.n1873 99.6594
R14144 gnd.n4431 gnd.n1874 99.6594
R14145 gnd.n1887 gnd.n1875 99.6594
R14146 gnd.n4443 gnd.n1876 99.6594
R14147 gnd.n4458 gnd.n4457 99.6594
R14148 gnd.n1919 gnd.n1864 99.6594
R14149 gnd.n1950 gnd.n1865 99.6594
R14150 gnd.n1915 gnd.n1866 99.6594
R14151 gnd.n4383 gnd.n1867 99.6594
R14152 gnd.n1910 gnd.n1868 99.6594
R14153 gnd.n4395 gnd.n1869 99.6594
R14154 gnd.n4406 gnd.n1870 99.6594
R14155 gnd.n1898 gnd.n1871 99.6594
R14156 gnd.n4419 gnd.n1872 99.6594
R14157 gnd.n4430 gnd.n1873 99.6594
R14158 gnd.n1886 gnd.n1874 99.6594
R14159 gnd.n4442 gnd.n1875 99.6594
R14160 gnd.n4456 gnd.n1876 99.6594
R14161 gnd.n4458 gnd.n1846 99.6594
R14162 gnd.n1356 gnd.n1217 99.6594
R14163 gnd.n5249 gnd.n1218 99.6594
R14164 gnd.n5251 gnd.n1219 99.6594
R14165 gnd.n5259 gnd.n1220 99.6594
R14166 gnd.n5262 gnd.n1221 99.6594
R14167 gnd.n5264 gnd.n1222 99.6594
R14168 gnd.n5484 gnd.n1223 99.6594
R14169 gnd.n5494 gnd.n1224 99.6594
R14170 gnd.n5496 gnd.n1225 99.6594
R14171 gnd.n5504 gnd.n1226 99.6594
R14172 gnd.n5514 gnd.n1227 99.6594
R14173 gnd.n5516 gnd.n1228 99.6594
R14174 gnd.n5524 gnd.n1229 99.6594
R14175 gnd.n5536 gnd.n1230 99.6594
R14176 gnd.n5523 gnd.n1228 99.6594
R14177 gnd.n5515 gnd.n1227 99.6594
R14178 gnd.n5513 gnd.n1226 99.6594
R14179 gnd.n5503 gnd.n1225 99.6594
R14180 gnd.n5495 gnd.n1224 99.6594
R14181 gnd.n5493 gnd.n1223 99.6594
R14182 gnd.n5483 gnd.n1222 99.6594
R14183 gnd.n5263 gnd.n1221 99.6594
R14184 gnd.n5261 gnd.n1220 99.6594
R14185 gnd.n5258 gnd.n1219 99.6594
R14186 gnd.n5252 gnd.n1218 99.6594
R14187 gnd.n5248 gnd.n1217 99.6594
R14188 gnd.n1230 gnd.n1214 99.6594
R14189 gnd.n5535 gnd.n1229 99.6594
R14190 gnd.n1877 gnd.t265 98.63
R14191 gnd.n5541 gnd.t296 98.63
R14192 gnd.n306 gnd.t311 98.63
R14193 gnd.n286 gnd.t227 98.63
R14194 gnd.n7076 gnd.t270 98.63
R14195 gnd.n1300 gnd.t293 98.63
R14196 gnd.n1323 gnd.t287 98.63
R14197 gnd.n1345 gnd.t220 98.63
R14198 gnd.n6895 gnd.t257 98.63
R14199 gnd.n1848 gnd.t314 98.63
R14200 gnd.n3844 gnd.t299 98.63
R14201 gnd.n3783 gnd.t245 98.63
R14202 gnd.n3805 gnd.t234 98.63
R14203 gnd.n3826 gnd.t224 98.63
R14204 gnd.n1035 gnd.t308 98.63
R14205 gnd.n1956 gnd.t241 98.63
R14206 gnd.n1969 gnd.t260 98.63
R14207 gnd.n5525 gnd.t248 98.63
R14208 gnd.n1722 gnd.t284 96.6984
R14209 gnd.n1455 gnd.t237 96.6984
R14210 gnd.n5832 gnd.t202 96.6906
R14211 gnd.n1449 gnd.t273 96.6906
R14212 gnd.n6506 gnd.n6505 84.828
R14213 gnd.n6507 gnd.n6506 84.828
R14214 gnd.n6507 gnd.n514 84.828
R14215 gnd.n6515 gnd.n514 84.828
R14216 gnd.n6516 gnd.n6515 84.828
R14217 gnd.n6517 gnd.n6516 84.828
R14218 gnd.n6517 gnd.n508 84.828
R14219 gnd.n6525 gnd.n508 84.828
R14220 gnd.n6526 gnd.n6525 84.828
R14221 gnd.n6527 gnd.n6526 84.828
R14222 gnd.n6527 gnd.n502 84.828
R14223 gnd.n6535 gnd.n502 84.828
R14224 gnd.n6536 gnd.n6535 84.828
R14225 gnd.n6537 gnd.n6536 84.828
R14226 gnd.n6537 gnd.n496 84.828
R14227 gnd.n6545 gnd.n496 84.828
R14228 gnd.n6546 gnd.n6545 84.828
R14229 gnd.n6547 gnd.n6546 84.828
R14230 gnd.n6547 gnd.n490 84.828
R14231 gnd.n6555 gnd.n490 84.828
R14232 gnd.n6556 gnd.n6555 84.828
R14233 gnd.n6557 gnd.n6556 84.828
R14234 gnd.n6557 gnd.n484 84.828
R14235 gnd.n6565 gnd.n484 84.828
R14236 gnd.n6566 gnd.n6565 84.828
R14237 gnd.n6567 gnd.n6566 84.828
R14238 gnd.n6567 gnd.n478 84.828
R14239 gnd.n6575 gnd.n478 84.828
R14240 gnd.n6576 gnd.n6575 84.828
R14241 gnd.n6577 gnd.n6576 84.828
R14242 gnd.n6577 gnd.n472 84.828
R14243 gnd.n6585 gnd.n472 84.828
R14244 gnd.n6586 gnd.n6585 84.828
R14245 gnd.n6587 gnd.n6586 84.828
R14246 gnd.n6587 gnd.n466 84.828
R14247 gnd.n6595 gnd.n466 84.828
R14248 gnd.n6596 gnd.n6595 84.828
R14249 gnd.n6597 gnd.n6596 84.828
R14250 gnd.n6597 gnd.n460 84.828
R14251 gnd.n6605 gnd.n460 84.828
R14252 gnd.n6606 gnd.n6605 84.828
R14253 gnd.n6607 gnd.n6606 84.828
R14254 gnd.n6607 gnd.n454 84.828
R14255 gnd.n6615 gnd.n454 84.828
R14256 gnd.n6616 gnd.n6615 84.828
R14257 gnd.n6617 gnd.n6616 84.828
R14258 gnd.n6617 gnd.n448 84.828
R14259 gnd.n6625 gnd.n448 84.828
R14260 gnd.n6626 gnd.n6625 84.828
R14261 gnd.n6627 gnd.n6626 84.828
R14262 gnd.n6627 gnd.n442 84.828
R14263 gnd.n6635 gnd.n442 84.828
R14264 gnd.n6636 gnd.n6635 84.828
R14265 gnd.n6637 gnd.n6636 84.828
R14266 gnd.n6637 gnd.n436 84.828
R14267 gnd.n6645 gnd.n436 84.828
R14268 gnd.n6646 gnd.n6645 84.828
R14269 gnd.n6647 gnd.n6646 84.828
R14270 gnd.n6647 gnd.n430 84.828
R14271 gnd.n6655 gnd.n430 84.828
R14272 gnd.n6656 gnd.n6655 84.828
R14273 gnd.n6657 gnd.n6656 84.828
R14274 gnd.n6657 gnd.n424 84.828
R14275 gnd.n6665 gnd.n424 84.828
R14276 gnd.n6666 gnd.n6665 84.828
R14277 gnd.n6667 gnd.n6666 84.828
R14278 gnd.n6667 gnd.n418 84.828
R14279 gnd.n6675 gnd.n418 84.828
R14280 gnd.n6676 gnd.n6675 84.828
R14281 gnd.n6677 gnd.n6676 84.828
R14282 gnd.n6677 gnd.n412 84.828
R14283 gnd.n6685 gnd.n412 84.828
R14284 gnd.n6686 gnd.n6685 84.828
R14285 gnd.n6687 gnd.n6686 84.828
R14286 gnd.n6687 gnd.n406 84.828
R14287 gnd.n6695 gnd.n406 84.828
R14288 gnd.n6696 gnd.n6695 84.828
R14289 gnd.n6697 gnd.n6696 84.828
R14290 gnd.n6697 gnd.n400 84.828
R14291 gnd.n6705 gnd.n400 84.828
R14292 gnd.n6706 gnd.n6705 84.828
R14293 gnd.n6708 gnd.n6706 84.828
R14294 gnd.n6708 gnd.n6707 84.828
R14295 gnd.n1097 gnd.n1096 81.8399
R14296 gnd.n2746 gnd.t280 74.8376
R14297 gnd.n2287 gnd.t303 74.8376
R14298 gnd.n1723 gnd.t283 72.8438
R14299 gnd.n1456 gnd.t238 72.8438
R14300 gnd.n1098 gnd.n1091 72.8411
R14301 gnd.n1104 gnd.n1089 72.8411
R14302 gnd.n1424 gnd.n1423 72.8411
R14303 gnd.n1878 gnd.t264 72.836
R14304 gnd.n5833 gnd.t201 72.836
R14305 gnd.n1450 gnd.t274 72.836
R14306 gnd.n5542 gnd.t295 72.836
R14307 gnd.n307 gnd.t312 72.836
R14308 gnd.n287 gnd.t228 72.836
R14309 gnd.n7077 gnd.t271 72.836
R14310 gnd.n1301 gnd.t292 72.836
R14311 gnd.n1324 gnd.t286 72.836
R14312 gnd.n1346 gnd.t219 72.836
R14313 gnd.n6896 gnd.t258 72.836
R14314 gnd.n1849 gnd.t315 72.836
R14315 gnd.n3845 gnd.t298 72.836
R14316 gnd.n3784 gnd.t244 72.836
R14317 gnd.n3806 gnd.t233 72.836
R14318 gnd.n3827 gnd.t223 72.836
R14319 gnd.n1036 gnd.t309 72.836
R14320 gnd.n1957 gnd.t242 72.836
R14321 gnd.n1970 gnd.t261 72.836
R14322 gnd.n5526 gnd.t249 72.836
R14323 gnd.n5177 gnd.n1429 71.676
R14324 gnd.n5175 gnd.n5174 71.676
R14325 gnd.n5170 gnd.n1432 71.676
R14326 gnd.n5168 gnd.n5167 71.676
R14327 gnd.n5163 gnd.n1435 71.676
R14328 gnd.n5161 gnd.n5160 71.676
R14329 gnd.n5156 gnd.n1438 71.676
R14330 gnd.n5154 gnd.n5153 71.676
R14331 gnd.n5149 gnd.n1441 71.676
R14332 gnd.n5147 gnd.n5146 71.676
R14333 gnd.n5142 gnd.n1444 71.676
R14334 gnd.n5140 gnd.n5139 71.676
R14335 gnd.n5135 gnd.n1447 71.676
R14336 gnd.n5133 gnd.n5132 71.676
R14337 gnd.n5127 gnd.n1452 71.676
R14338 gnd.n5125 gnd.n5124 71.676
R14339 gnd.n5120 gnd.n5119 71.676
R14340 gnd.n5117 gnd.n5116 71.676
R14341 gnd.n5111 gnd.n1458 71.676
R14342 gnd.n5109 gnd.n5108 71.676
R14343 gnd.n5104 gnd.n1461 71.676
R14344 gnd.n5102 gnd.n5101 71.676
R14345 gnd.n5097 gnd.n1464 71.676
R14346 gnd.n5095 gnd.n5094 71.676
R14347 gnd.n5090 gnd.n1467 71.676
R14348 gnd.n5088 gnd.n5087 71.676
R14349 gnd.n5083 gnd.n1470 71.676
R14350 gnd.n5081 gnd.n5080 71.676
R14351 gnd.n5076 gnd.n1473 71.676
R14352 gnd.n5074 gnd.n5073 71.676
R14353 gnd.n5069 gnd.n1476 71.676
R14354 gnd.n5067 gnd.n5066 71.676
R14355 gnd.n5062 gnd.n5061 71.676
R14356 gnd.n5896 gnd.n5895 71.676
R14357 gnd.n5890 gnd.n1053 71.676
R14358 gnd.n5887 gnd.n1054 71.676
R14359 gnd.n5883 gnd.n1055 71.676
R14360 gnd.n5879 gnd.n1056 71.676
R14361 gnd.n5875 gnd.n1057 71.676
R14362 gnd.n5871 gnd.n1058 71.676
R14363 gnd.n5867 gnd.n1059 71.676
R14364 gnd.n5863 gnd.n1060 71.676
R14365 gnd.n5859 gnd.n1061 71.676
R14366 gnd.n5855 gnd.n1062 71.676
R14367 gnd.n5851 gnd.n1063 71.676
R14368 gnd.n5847 gnd.n1064 71.676
R14369 gnd.n5843 gnd.n1065 71.676
R14370 gnd.n5839 gnd.n1066 71.676
R14371 gnd.n5835 gnd.n1067 71.676
R14372 gnd.n1068 gnd.n1051 71.676
R14373 gnd.n1726 gnd.n1069 71.676
R14374 gnd.n1731 gnd.n1070 71.676
R14375 gnd.n1735 gnd.n1071 71.676
R14376 gnd.n1739 gnd.n1072 71.676
R14377 gnd.n1743 gnd.n1073 71.676
R14378 gnd.n1747 gnd.n1074 71.676
R14379 gnd.n1751 gnd.n1075 71.676
R14380 gnd.n1755 gnd.n1076 71.676
R14381 gnd.n1759 gnd.n1077 71.676
R14382 gnd.n1763 gnd.n1078 71.676
R14383 gnd.n1767 gnd.n1079 71.676
R14384 gnd.n1771 gnd.n1080 71.676
R14385 gnd.n1775 gnd.n1081 71.676
R14386 gnd.n1779 gnd.n1082 71.676
R14387 gnd.n1783 gnd.n1083 71.676
R14388 gnd.n5896 gnd.n1086 71.676
R14389 gnd.n5888 gnd.n1053 71.676
R14390 gnd.n5884 gnd.n1054 71.676
R14391 gnd.n5880 gnd.n1055 71.676
R14392 gnd.n5876 gnd.n1056 71.676
R14393 gnd.n5872 gnd.n1057 71.676
R14394 gnd.n5868 gnd.n1058 71.676
R14395 gnd.n5864 gnd.n1059 71.676
R14396 gnd.n5860 gnd.n1060 71.676
R14397 gnd.n5856 gnd.n1061 71.676
R14398 gnd.n5852 gnd.n1062 71.676
R14399 gnd.n5848 gnd.n1063 71.676
R14400 gnd.n5844 gnd.n1064 71.676
R14401 gnd.n5840 gnd.n1065 71.676
R14402 gnd.n5836 gnd.n1066 71.676
R14403 gnd.n5899 gnd.n5898 71.676
R14404 gnd.n1725 gnd.n1068 71.676
R14405 gnd.n1730 gnd.n1069 71.676
R14406 gnd.n1734 gnd.n1070 71.676
R14407 gnd.n1738 gnd.n1071 71.676
R14408 gnd.n1742 gnd.n1072 71.676
R14409 gnd.n1746 gnd.n1073 71.676
R14410 gnd.n1750 gnd.n1074 71.676
R14411 gnd.n1754 gnd.n1075 71.676
R14412 gnd.n1758 gnd.n1076 71.676
R14413 gnd.n1762 gnd.n1077 71.676
R14414 gnd.n1766 gnd.n1078 71.676
R14415 gnd.n1770 gnd.n1079 71.676
R14416 gnd.n1774 gnd.n1080 71.676
R14417 gnd.n1778 gnd.n1081 71.676
R14418 gnd.n1782 gnd.n1082 71.676
R14419 gnd.n1786 gnd.n1083 71.676
R14420 gnd.n5061 gnd.n1477 71.676
R14421 gnd.n5068 gnd.n5067 71.676
R14422 gnd.n1476 gnd.n1474 71.676
R14423 gnd.n5075 gnd.n5074 71.676
R14424 gnd.n1473 gnd.n1471 71.676
R14425 gnd.n5082 gnd.n5081 71.676
R14426 gnd.n1470 gnd.n1468 71.676
R14427 gnd.n5089 gnd.n5088 71.676
R14428 gnd.n1467 gnd.n1465 71.676
R14429 gnd.n5096 gnd.n5095 71.676
R14430 gnd.n1464 gnd.n1462 71.676
R14431 gnd.n5103 gnd.n5102 71.676
R14432 gnd.n1461 gnd.n1459 71.676
R14433 gnd.n5110 gnd.n5109 71.676
R14434 gnd.n1458 gnd.n1454 71.676
R14435 gnd.n5118 gnd.n5117 71.676
R14436 gnd.n5122 gnd.n5121 71.676
R14437 gnd.n5126 gnd.n5125 71.676
R14438 gnd.n1452 gnd.n1448 71.676
R14439 gnd.n5134 gnd.n5133 71.676
R14440 gnd.n1447 gnd.n1445 71.676
R14441 gnd.n5141 gnd.n5140 71.676
R14442 gnd.n1444 gnd.n1442 71.676
R14443 gnd.n5148 gnd.n5147 71.676
R14444 gnd.n1441 gnd.n1439 71.676
R14445 gnd.n5155 gnd.n5154 71.676
R14446 gnd.n1438 gnd.n1436 71.676
R14447 gnd.n5162 gnd.n5161 71.676
R14448 gnd.n1435 gnd.n1433 71.676
R14449 gnd.n5169 gnd.n5168 71.676
R14450 gnd.n1432 gnd.n1430 71.676
R14451 gnd.n5176 gnd.n5175 71.676
R14452 gnd.n1429 gnd.n1407 71.676
R14453 gnd.n8 gnd.t12 69.1507
R14454 gnd.n14 gnd.t193 68.4792
R14455 gnd.n13 gnd.t355 68.4792
R14456 gnd.n12 gnd.t198 68.4792
R14457 gnd.n11 gnd.t180 68.4792
R14458 gnd.n10 gnd.t351 68.4792
R14459 gnd.n9 gnd.t324 68.4792
R14460 gnd.n8 gnd.t185 68.4792
R14461 gnd.n2873 gnd.n2777 64.369
R14462 gnd.n1728 gnd.n1723 59.5399
R14463 gnd.n5113 gnd.n1456 59.5399
R14464 gnd.n5834 gnd.n5833 59.5399
R14465 gnd.n5129 gnd.n1450 59.5399
R14466 gnd.n5831 gnd.n1107 59.1804
R14467 gnd.n4039 gnd.n2237 57.3586
R14468 gnd.n7111 gnd.n204 57.3586
R14469 gnd.n2528 gnd.t90 56.407
R14470 gnd.n2481 gnd.t153 56.407
R14471 gnd.n2496 gnd.t37 56.407
R14472 gnd.n2512 gnd.t141 56.407
R14473 gnd.n64 gnd.t56 56.407
R14474 gnd.n17 gnd.t44 56.407
R14475 gnd.n32 gnd.t168 56.407
R14476 gnd.n48 gnd.t107 56.407
R14477 gnd.n2541 gnd.t74 55.8337
R14478 gnd.n2494 gnd.t163 55.8337
R14479 gnd.n2509 gnd.t134 55.8337
R14480 gnd.n2525 gnd.t119 55.8337
R14481 gnd.n77 gnd.t14 55.8337
R14482 gnd.n30 gnd.t63 55.8337
R14483 gnd.n45 gnd.t123 55.8337
R14484 gnd.n61 gnd.t85 55.8337
R14485 gnd.n1095 gnd.n1094 54.358
R14486 gnd.n1421 gnd.n1420 54.358
R14487 gnd.n2528 gnd.n2527 53.0052
R14488 gnd.n2530 gnd.n2529 53.0052
R14489 gnd.n2532 gnd.n2531 53.0052
R14490 gnd.n2534 gnd.n2533 53.0052
R14491 gnd.n2536 gnd.n2535 53.0052
R14492 gnd.n2538 gnd.n2537 53.0052
R14493 gnd.n2540 gnd.n2539 53.0052
R14494 gnd.n2481 gnd.n2480 53.0052
R14495 gnd.n2483 gnd.n2482 53.0052
R14496 gnd.n2485 gnd.n2484 53.0052
R14497 gnd.n2487 gnd.n2486 53.0052
R14498 gnd.n2489 gnd.n2488 53.0052
R14499 gnd.n2491 gnd.n2490 53.0052
R14500 gnd.n2493 gnd.n2492 53.0052
R14501 gnd.n2496 gnd.n2495 53.0052
R14502 gnd.n2498 gnd.n2497 53.0052
R14503 gnd.n2500 gnd.n2499 53.0052
R14504 gnd.n2502 gnd.n2501 53.0052
R14505 gnd.n2504 gnd.n2503 53.0052
R14506 gnd.n2506 gnd.n2505 53.0052
R14507 gnd.n2508 gnd.n2507 53.0052
R14508 gnd.n2512 gnd.n2511 53.0052
R14509 gnd.n2514 gnd.n2513 53.0052
R14510 gnd.n2516 gnd.n2515 53.0052
R14511 gnd.n2518 gnd.n2517 53.0052
R14512 gnd.n2520 gnd.n2519 53.0052
R14513 gnd.n2522 gnd.n2521 53.0052
R14514 gnd.n2524 gnd.n2523 53.0052
R14515 gnd.n76 gnd.n75 53.0052
R14516 gnd.n74 gnd.n73 53.0052
R14517 gnd.n72 gnd.n71 53.0052
R14518 gnd.n70 gnd.n69 53.0052
R14519 gnd.n68 gnd.n67 53.0052
R14520 gnd.n66 gnd.n65 53.0052
R14521 gnd.n64 gnd.n63 53.0052
R14522 gnd.n29 gnd.n28 53.0052
R14523 gnd.n27 gnd.n26 53.0052
R14524 gnd.n25 gnd.n24 53.0052
R14525 gnd.n23 gnd.n22 53.0052
R14526 gnd.n21 gnd.n20 53.0052
R14527 gnd.n19 gnd.n18 53.0052
R14528 gnd.n17 gnd.n16 53.0052
R14529 gnd.n44 gnd.n43 53.0052
R14530 gnd.n42 gnd.n41 53.0052
R14531 gnd.n40 gnd.n39 53.0052
R14532 gnd.n38 gnd.n37 53.0052
R14533 gnd.n36 gnd.n35 53.0052
R14534 gnd.n34 gnd.n33 53.0052
R14535 gnd.n32 gnd.n31 53.0052
R14536 gnd.n60 gnd.n59 53.0052
R14537 gnd.n58 gnd.n57 53.0052
R14538 gnd.n56 gnd.n55 53.0052
R14539 gnd.n54 gnd.n53 53.0052
R14540 gnd.n52 gnd.n51 53.0052
R14541 gnd.n50 gnd.n49 53.0052
R14542 gnd.n48 gnd.n47 53.0052
R14543 gnd.n1412 gnd.n1411 52.4801
R14544 gnd.n3577 gnd.t1 52.3082
R14545 gnd.n3545 gnd.t347 52.3082
R14546 gnd.n3513 gnd.t5 52.3082
R14547 gnd.n3482 gnd.t3 52.3082
R14548 gnd.n3450 gnd.t7 52.3082
R14549 gnd.n3418 gnd.t359 52.3082
R14550 gnd.n3386 gnd.t187 52.3082
R14551 gnd.n3355 gnd.t357 52.3082
R14552 gnd.n3407 gnd.n3375 51.4173
R14553 gnd.n6707 gnd.n157 50.897
R14554 gnd.n3471 gnd.n3470 50.455
R14555 gnd.n3439 gnd.n3438 50.455
R14556 gnd.n3407 gnd.n3406 50.455
R14557 gnd.n2820 gnd.n2819 45.1884
R14558 gnd.n2313 gnd.n2312 45.1884
R14559 gnd.n5180 gnd.n1427 44.3322
R14560 gnd.n1098 gnd.n1097 44.3189
R14561 gnd.n1879 gnd.n1878 42.2793
R14562 gnd.n5543 gnd.n5542 42.2793
R14563 gnd.n6994 gnd.n307 42.2793
R14564 gnd.n7036 gnd.n287 42.2793
R14565 gnd.n7078 gnd.n7077 42.2793
R14566 gnd.n5672 gnd.n1301 42.2793
R14567 gnd.n5635 gnd.n1324 42.2793
R14568 gnd.n5595 gnd.n1346 42.2793
R14569 gnd.n6897 gnd.n6896 42.2793
R14570 gnd.n2821 gnd.n2820 42.2793
R14571 gnd.n2314 gnd.n2313 42.2793
R14572 gnd.n2747 gnd.n2746 42.2793
R14573 gnd.n3692 gnd.n2287 42.2793
R14574 gnd.n1850 gnd.n1849 42.2793
R14575 gnd.n3846 gnd.n3845 42.2793
R14576 gnd.n4003 gnd.n3784 42.2793
R14577 gnd.n3963 gnd.n3806 42.2793
R14578 gnd.n3924 gnd.n3827 42.2793
R14579 gnd.n5918 gnd.n1036 42.2793
R14580 gnd.n2047 gnd.n1957 42.2793
R14581 gnd.n1998 gnd.n1970 42.2793
R14582 gnd.n5527 gnd.n5526 42.2793
R14583 gnd.n1096 gnd.n1095 41.6274
R14584 gnd.n1422 gnd.n1421 41.6274
R14585 gnd.n1105 gnd.n1104 40.8975
R14586 gnd.n1425 gnd.n1424 40.8975
R14587 gnd.n1104 gnd.n1103 35.055
R14588 gnd.n1099 gnd.n1098 35.055
R14589 gnd.n1414 gnd.n1413 35.055
R14590 gnd.n1424 gnd.n1410 35.055
R14591 gnd.n5063 gnd.n5060 33.2493
R14592 gnd.n1789 gnd.n1785 33.2493
R14593 gnd.n6176 gnd.n6175 31.9912
R14594 gnd.n6175 gnd.n6174 31.9912
R14595 gnd.n6174 gnd.n717 31.9912
R14596 gnd.n6168 gnd.n717 31.9912
R14597 gnd.n6168 gnd.n6167 31.9912
R14598 gnd.n6167 gnd.n6166 31.9912
R14599 gnd.n6166 gnd.n724 31.9912
R14600 gnd.n6160 gnd.n724 31.9912
R14601 gnd.n6160 gnd.n6159 31.9912
R14602 gnd.n6159 gnd.n6158 31.9912
R14603 gnd.n6158 gnd.n732 31.9912
R14604 gnd.n6152 gnd.n732 31.9912
R14605 gnd.n6152 gnd.n6151 31.9912
R14606 gnd.n6151 gnd.n6150 31.9912
R14607 gnd.n6150 gnd.n740 31.9912
R14608 gnd.n6144 gnd.n740 31.9912
R14609 gnd.n6144 gnd.n6143 31.9912
R14610 gnd.n6143 gnd.n6142 31.9912
R14611 gnd.n6142 gnd.n748 31.9912
R14612 gnd.n6136 gnd.n748 31.9912
R14613 gnd.n6136 gnd.n6135 31.9912
R14614 gnd.n6135 gnd.n6134 31.9912
R14615 gnd.n6134 gnd.n756 31.9912
R14616 gnd.n6128 gnd.n756 31.9912
R14617 gnd.n6128 gnd.n6127 31.9912
R14618 gnd.n6127 gnd.n6126 31.9912
R14619 gnd.n6126 gnd.n764 31.9912
R14620 gnd.n6120 gnd.n764 31.9912
R14621 gnd.n6120 gnd.n6119 31.9912
R14622 gnd.n6119 gnd.n6118 31.9912
R14623 gnd.n6118 gnd.n772 31.9912
R14624 gnd.n6112 gnd.n772 31.9912
R14625 gnd.n6112 gnd.n6111 31.9912
R14626 gnd.n6111 gnd.n6110 31.9912
R14627 gnd.n6110 gnd.n780 31.9912
R14628 gnd.n6104 gnd.n780 31.9912
R14629 gnd.n6104 gnd.n6103 31.9912
R14630 gnd.n6103 gnd.n6102 31.9912
R14631 gnd.n6102 gnd.n788 31.9912
R14632 gnd.n6096 gnd.n788 31.9912
R14633 gnd.n6096 gnd.n6095 31.9912
R14634 gnd.n6095 gnd.n6094 31.9912
R14635 gnd.n6094 gnd.n796 31.9912
R14636 gnd.n6088 gnd.n796 31.9912
R14637 gnd.n6088 gnd.n6087 31.9912
R14638 gnd.n6087 gnd.n6086 31.9912
R14639 gnd.n6086 gnd.n804 31.9912
R14640 gnd.n6080 gnd.n804 31.9912
R14641 gnd.n6080 gnd.n6079 31.9912
R14642 gnd.n6079 gnd.n6078 31.9912
R14643 gnd.n6078 gnd.n812 31.9912
R14644 gnd.n6072 gnd.n812 31.9912
R14645 gnd.n6072 gnd.n6071 31.9912
R14646 gnd.n6071 gnd.n6070 31.9912
R14647 gnd.n6070 gnd.n820 31.9912
R14648 gnd.n6064 gnd.n820 31.9912
R14649 gnd.n6064 gnd.n6063 31.9912
R14650 gnd.n6063 gnd.n6062 31.9912
R14651 gnd.n6062 gnd.n828 31.9912
R14652 gnd.n6056 gnd.n828 31.9912
R14653 gnd.n6056 gnd.n6055 31.9912
R14654 gnd.n6055 gnd.n6054 31.9912
R14655 gnd.n6054 gnd.n836 31.9912
R14656 gnd.n6048 gnd.n836 31.9912
R14657 gnd.n6048 gnd.n6047 31.9912
R14658 gnd.n6047 gnd.n6046 31.9912
R14659 gnd.n6046 gnd.n844 31.9912
R14660 gnd.n6040 gnd.n844 31.9912
R14661 gnd.n6040 gnd.n6039 31.9912
R14662 gnd.n6039 gnd.n6038 31.9912
R14663 gnd.n6038 gnd.n852 31.9912
R14664 gnd.n6032 gnd.n852 31.9912
R14665 gnd.n6032 gnd.n6031 31.9912
R14666 gnd.n6031 gnd.n6030 31.9912
R14667 gnd.n6030 gnd.n860 31.9912
R14668 gnd.n6024 gnd.n860 31.9912
R14669 gnd.n6024 gnd.n6023 31.9912
R14670 gnd.n6023 gnd.n6022 31.9912
R14671 gnd.n6022 gnd.n868 31.9912
R14672 gnd.n6016 gnd.n868 31.9912
R14673 gnd.n6016 gnd.n6015 31.9912
R14674 gnd.n6015 gnd.n6014 31.9912
R14675 gnd.n6014 gnd.n876 31.9912
R14676 gnd.n2883 gnd.n2777 31.8661
R14677 gnd.n2883 gnd.n2882 31.8661
R14678 gnd.n2891 gnd.n2766 31.8661
R14679 gnd.n2899 gnd.n2766 31.8661
R14680 gnd.n2899 gnd.n2760 31.8661
R14681 gnd.n2907 gnd.n2760 31.8661
R14682 gnd.n2907 gnd.n2753 31.8661
R14683 gnd.n2945 gnd.n2753 31.8661
R14684 gnd.n2955 gnd.n2686 31.8661
R14685 gnd.n4052 gnd.n2237 31.8661
R14686 gnd.n4060 gnd.n2229 31.8661
R14687 gnd.n4060 gnd.n2218 31.8661
R14688 gnd.n4072 gnd.n2218 31.8661
R14689 gnd.n4072 gnd.n2221 31.8661
R14690 gnd.n4080 gnd.n2201 31.8661
R14691 gnd.n4092 gnd.n2201 31.8661
R14692 gnd.n4100 gnd.n2193 31.8661
R14693 gnd.n4116 gnd.n2181 31.8661
R14694 gnd.n4116 gnd.n2184 31.8661
R14695 gnd.n4126 gnd.n2167 31.8661
R14696 gnd.n4136 gnd.n2167 31.8661
R14697 gnd.n4151 gnd.n2158 31.8661
R14698 gnd.n4161 gnd.n2142 31.8661
R14699 gnd.n4171 gnd.n2142 31.8661
R14700 gnd.n4186 gnd.n2123 31.8661
R14701 gnd.n4196 gnd.n2123 31.8661
R14702 gnd.n4218 gnd.n2116 31.8661
R14703 gnd.n4229 gnd.n2099 31.8661
R14704 gnd.n4237 gnd.n2099 31.8661
R14705 gnd.n4256 gnd.n2086 31.8661
R14706 gnd.n4256 gnd.n2089 31.8661
R14707 gnd.n4265 gnd.n883 31.8661
R14708 gnd.n4467 gnd.n978 31.8661
R14709 gnd.n4460 gnd.n989 31.8661
R14710 gnd.n4460 gnd.n4459 31.8661
R14711 gnd.n4459 gnd.n1840 31.8661
R14712 gnd.n4480 gnd.n1840 31.8661
R14713 gnd.n4480 gnd.n1842 31.8661
R14714 gnd.n4488 gnd.n1827 31.8661
R14715 gnd.n4496 gnd.n1827 31.8661
R14716 gnd.n4496 gnd.n1820 31.8661
R14717 gnd.n4504 gnd.n1820 31.8661
R14718 gnd.n4530 gnd.n1811 31.8661
R14719 gnd.n4530 gnd.n1803 31.8661
R14720 gnd.n4547 gnd.n1803 31.8661
R14721 gnd.n4510 gnd.n1052 31.8661
R14722 gnd.n5200 gnd.n1381 31.8661
R14723 gnd.n5208 gnd.n1381 31.8661
R14724 gnd.n5208 gnd.n1382 31.8661
R14725 gnd.n5216 gnd.n1369 31.8661
R14726 gnd.n5224 gnd.n1369 31.8661
R14727 gnd.n5224 gnd.n1363 31.8661
R14728 gnd.n5232 gnd.n1363 31.8661
R14729 gnd.n5241 gnd.n1357 31.8661
R14730 gnd.n5241 gnd.n1216 31.8661
R14731 gnd.n5715 gnd.n1216 31.8661
R14732 gnd.n5715 gnd.n1231 31.8661
R14733 gnd.n5709 gnd.n1231 31.8661
R14734 gnd.n5270 gnd.n1278 31.8661
R14735 gnd.n6769 gnd.n354 31.8661
R14736 gnd.n6779 gnd.n336 31.8661
R14737 gnd.n6793 gnd.n336 31.8661
R14738 gnd.n6802 gnd.n319 31.8661
R14739 gnd.n6813 gnd.n319 31.8661
R14740 gnd.n6821 gnd.n313 31.8661
R14741 gnd.n7191 gnd.n86 31.8661
R14742 gnd.n7185 gnd.n86 31.8661
R14743 gnd.n7179 gnd.n106 31.8661
R14744 gnd.n7179 gnd.n109 31.8661
R14745 gnd.n7173 gnd.n119 31.8661
R14746 gnd.n7167 gnd.n128 31.8661
R14747 gnd.n7161 gnd.n128 31.8661
R14748 gnd.n7155 gnd.n144 31.8661
R14749 gnd.n7155 gnd.n147 31.8661
R14750 gnd.n7143 gnd.n166 31.8661
R14751 gnd.n7137 gnd.n166 31.8661
R14752 gnd.n7131 gnd.n182 31.8661
R14753 gnd.n7131 gnd.n185 31.8661
R14754 gnd.n7125 gnd.n185 31.8661
R14755 gnd.n7125 gnd.n195 31.8661
R14756 gnd.n7119 gnd.n204 31.8661
R14757 gnd.n4547 gnd.t11 30.9101
R14758 gnd.n5200 gnd.t182 30.9101
R14759 gnd.t289 gnd.n1395 30.5915
R14760 gnd.n3725 gnd.n2247 29.9541
R14761 gnd.n5897 gnd.n1084 28.3609
R14762 gnd.n1405 gnd.n1394 28.3609
R14763 gnd.n4100 gnd.t98 27.7236
R14764 gnd.n7149 gnd.t65 27.7236
R14765 gnd.n2322 gnd.n2247 27.4049
R14766 gnd.n5951 gnd.n989 27.4049
R14767 gnd.n5709 gnd.n5708 27.4049
R14768 gnd.n2158 gnd.t77 27.0862
R14769 gnd.n4265 gnd.t94 27.0862
R14770 gnd.n354 gnd.t61 27.0862
R14771 gnd.n7173 gnd.t21 27.0862
R14772 gnd.t92 gnd.n2116 26.4489
R14773 gnd.n4218 gnd.t48 26.4489
R14774 gnd.t19 gnd.n313 26.4489
R14775 gnd.n6821 gnd.t57 26.4489
R14776 gnd.n4151 gnd.t28 25.8116
R14777 gnd.t75 gnd.n119 25.8116
R14778 gnd.n1878 gnd.n1877 25.7944
R14779 gnd.n5542 gnd.n5541 25.7944
R14780 gnd.n307 gnd.n306 25.7944
R14781 gnd.n287 gnd.n286 25.7944
R14782 gnd.n7077 gnd.n7076 25.7944
R14783 gnd.n1301 gnd.n1300 25.7944
R14784 gnd.n1324 gnd.n1323 25.7944
R14785 gnd.n1346 gnd.n1345 25.7944
R14786 gnd.n6896 gnd.n6895 25.7944
R14787 gnd.n2746 gnd.n2745 25.7944
R14788 gnd.n2287 gnd.n2286 25.7944
R14789 gnd.n1849 gnd.n1848 25.7944
R14790 gnd.n3845 gnd.n3844 25.7944
R14791 gnd.n3784 gnd.n3783 25.7944
R14792 gnd.n3806 gnd.n3805 25.7944
R14793 gnd.n3827 gnd.n3826 25.7944
R14794 gnd.n1036 gnd.n1035 25.7944
R14795 gnd.n1957 gnd.n1956 25.7944
R14796 gnd.n1970 gnd.n1969 25.7944
R14797 gnd.n5526 gnd.n5525 25.7944
R14798 gnd.t46 gnd.n2193 25.1743
R14799 gnd.n6969 gnd.t30 25.1743
R14800 gnd.n2967 gnd.n2687 24.8557
R14801 gnd.n2977 gnd.n2670 24.8557
R14802 gnd.n2673 gnd.n2661 24.8557
R14803 gnd.n2998 gnd.n2662 24.8557
R14804 gnd.n3008 gnd.n2642 24.8557
R14805 gnd.n3018 gnd.n3017 24.8557
R14806 gnd.n2628 gnd.n2626 24.8557
R14807 gnd.n3049 gnd.n3048 24.8557
R14808 gnd.n3064 gnd.n2611 24.8557
R14809 gnd.n3118 gnd.n2550 24.8557
R14810 gnd.n3074 gnd.n2551 24.8557
R14811 gnd.n3111 gnd.n2562 24.8557
R14812 gnd.n2600 gnd.n2599 24.8557
R14813 gnd.n3105 gnd.n3104 24.8557
R14814 gnd.n2586 gnd.n2573 24.8557
R14815 gnd.n3144 gnd.n3143 24.8557
R14816 gnd.n3154 gnd.n2466 24.8557
R14817 gnd.n3166 gnd.n2458 24.8557
R14818 gnd.n3165 gnd.n2446 24.8557
R14819 gnd.n3184 gnd.n3183 24.8557
R14820 gnd.n3194 gnd.n2439 24.8557
R14821 gnd.n3205 gnd.n2427 24.8557
R14822 gnd.n3229 gnd.n3228 24.8557
R14823 gnd.n3240 gnd.n2410 24.8557
R14824 gnd.n3239 gnd.n2412 24.8557
R14825 gnd.n3251 gnd.n2403 24.8557
R14826 gnd.n3269 gnd.n3268 24.8557
R14827 gnd.n2394 gnd.n2383 24.8557
R14828 gnd.n3290 gnd.n2371 24.8557
R14829 gnd.n3318 gnd.n3317 24.8557
R14830 gnd.n3329 gnd.n2356 24.8557
R14831 gnd.n3340 gnd.n2349 24.8557
R14832 gnd.n3339 gnd.n2337 24.8557
R14833 gnd.n3612 gnd.n3611 24.8557
R14834 gnd.n3634 gnd.n2321 24.8557
R14835 gnd.n1723 gnd.n1722 23.855
R14836 gnd.n1456 gnd.n1455 23.855
R14837 gnd.n5833 gnd.n5832 23.855
R14838 gnd.n1450 gnd.n1449 23.855
R14839 gnd.n2988 gnd.t356 23.2624
R14840 gnd.n2689 gnd.t279 22.6251
R14841 gnd.n4052 gnd.t222 22.6251
R14842 gnd.n7119 gnd.t226 22.6251
R14843 gnd.n6008 gnd.t41 21.6691
R14844 gnd.n4643 gnd.n1713 21.6691
R14845 gnd.n4664 gnd.n1706 21.6691
R14846 gnd.n4671 gnd.n4670 21.6691
R14847 gnd.n4689 gnd.n1692 21.6691
R14848 gnd.n4706 gnd.n1674 21.6691
R14849 gnd.n4764 gnd.n4763 21.6691
R14850 gnd.n4796 gnd.n1626 21.6691
R14851 gnd.n4807 gnd.n1621 21.6691
R14852 gnd.n4841 gnd.n1600 21.6691
R14853 gnd.n4847 gnd.n1596 21.6691
R14854 gnd.n4865 gnd.n1577 21.6691
R14855 gnd.n4948 gnd.n1543 21.6691
R14856 gnd.n4875 gnd.n1532 21.6691
R14857 gnd.n5003 gnd.n1521 21.6691
R14858 gnd.n5021 gnd.n1505 21.6691
R14859 gnd.n5056 gnd.n1402 21.6691
R14860 gnd.t17 gnd.n351 21.6691
R14861 gnd.t2 gnd.n2694 21.3504
R14862 gnd.n5831 gnd.n5830 21.0737
R14863 gnd.n5181 gnd.n5180 21.0737
R14864 gnd.n6007 gnd.n886 21.0318
R14865 gnd.n4274 gnd.n896 21.0318
R14866 gnd.n4294 gnd.n907 21.0318
R14867 gnd.n5995 gnd.n910 21.0318
R14868 gnd.n5989 gnd.n921 21.0318
R14869 gnd.n4340 gnd.n4339 21.0318
R14870 gnd.n5983 gnd.n930 21.0318
R14871 gnd.n4347 gnd.n938 21.0318
R14872 gnd.n4355 gnd.n947 21.0318
R14873 gnd.n5971 gnd.n950 21.0318
R14874 gnd.n4362 gnd.n958 21.0318
R14875 gnd.n5965 gnd.n961 21.0318
R14876 gnd.n5959 gnd.n971 21.0318
R14877 gnd.n4468 gnd.n4467 21.0318
R14878 gnd.n4683 gnd.n1696 21.0318
R14879 gnd.n1620 gnd.n1608 21.0318
R14880 gnd.n1612 gnd.n1609 21.0318
R14881 gnd.n5004 gnd.n1518 21.0318
R14882 gnd.n5475 gnd.n5270 21.0318
R14883 gnd.n5474 gnd.n5274 21.0318
R14884 gnd.n5468 gnd.n5467 21.0318
R14885 gnd.n5380 gnd.n5289 21.0318
R14886 gnd.n5461 gnd.n5305 21.0318
R14887 gnd.n5400 gnd.n5308 21.0318
R14888 gnd.n5408 gnd.n5319 21.0318
R14889 gnd.n5449 gnd.n5327 21.0318
R14890 gnd.n5427 gnd.n5426 21.0318
R14891 gnd.n5443 gnd.n5334 21.0318
R14892 gnd.n6735 gnd.n379 21.0318
R14893 gnd.n6722 gnd.n382 21.0318
R14894 gnd.n6728 gnd.n371 21.0318
R14895 gnd.n6754 gnd.n363 21.0318
R14896 gnd.t337 gnd.n2384 20.7131
R14897 gnd.t352 gnd.n1811 20.7131
R14898 gnd.n1382 gnd.t192 20.7131
R14899 gnd.n5050 gnd.t236 20.3945
R14900 gnd.t339 gnd.n2419 20.0758
R14901 gnd.n1093 gnd.t277 19.8005
R14902 gnd.n1093 gnd.t231 19.8005
R14903 gnd.n1092 gnd.t252 19.8005
R14904 gnd.n1092 gnd.t306 19.8005
R14905 gnd.n1419 gnd.t318 19.8005
R14906 gnd.n1419 gnd.t268 19.8005
R14907 gnd.n1418 gnd.t216 19.8005
R14908 gnd.n1418 gnd.t290 19.8005
R14909 gnd.n5827 gnd.t276 19.7572
R14910 gnd.t327 gnd.n4700 19.7572
R14911 gnd.n4795 gnd.n4793 19.7572
R14912 gnd.n4848 gnd.n1593 19.7572
R14913 gnd.n1542 gnd.t8 19.7572
R14914 gnd.n1089 gnd.n1088 19.5087
R14915 gnd.n1102 gnd.n1089 19.5087
R14916 gnd.n1100 gnd.n1091 19.5087
R14917 gnd.n1423 gnd.n1417 19.5087
R14918 gnd.n3155 gnd.t345 19.4385
R14919 gnd.n4478 gnd.n1832 19.3944
R14920 gnd.n4490 gnd.n1832 19.3944
R14921 gnd.n4490 gnd.n1830 19.3944
R14922 gnd.n4494 gnd.n1830 19.3944
R14923 gnd.n4494 gnd.n1818 19.3944
R14924 gnd.n4506 gnd.n1818 19.3944
R14925 gnd.n4506 gnd.n1815 19.3944
R14926 gnd.n4528 gnd.n1815 19.3944
R14927 gnd.n4528 gnd.n1816 19.3944
R14928 gnd.n4524 gnd.n1816 19.3944
R14929 gnd.n4524 gnd.n4523 19.3944
R14930 gnd.n4523 gnd.n4522 19.3944
R14931 gnd.n4522 gnd.n4513 19.3944
R14932 gnd.n4518 gnd.n4513 19.3944
R14933 gnd.n4518 gnd.n4517 19.3944
R14934 gnd.n4517 gnd.n1129 19.3944
R14935 gnd.n5817 gnd.n1129 19.3944
R14936 gnd.n5817 gnd.n1130 19.3944
R14937 gnd.n5813 gnd.n1130 19.3944
R14938 gnd.n5813 gnd.n5812 19.3944
R14939 gnd.n5812 gnd.n5811 19.3944
R14940 gnd.n5811 gnd.n1136 19.3944
R14941 gnd.n5807 gnd.n1136 19.3944
R14942 gnd.n5807 gnd.n5806 19.3944
R14943 gnd.n5806 gnd.n5805 19.3944
R14944 gnd.n5805 gnd.n1141 19.3944
R14945 gnd.n5801 gnd.n1141 19.3944
R14946 gnd.n5801 gnd.n5800 19.3944
R14947 gnd.n5800 gnd.n5799 19.3944
R14948 gnd.n5799 gnd.n1146 19.3944
R14949 gnd.n5795 gnd.n1146 19.3944
R14950 gnd.n5795 gnd.n5794 19.3944
R14951 gnd.n5794 gnd.n5793 19.3944
R14952 gnd.n5793 gnd.n1151 19.3944
R14953 gnd.n5789 gnd.n1151 19.3944
R14954 gnd.n5789 gnd.n5788 19.3944
R14955 gnd.n5788 gnd.n5787 19.3944
R14956 gnd.n5787 gnd.n1156 19.3944
R14957 gnd.n5783 gnd.n1156 19.3944
R14958 gnd.n5783 gnd.n5782 19.3944
R14959 gnd.n5782 gnd.n5781 19.3944
R14960 gnd.n5781 gnd.n1161 19.3944
R14961 gnd.n5777 gnd.n1161 19.3944
R14962 gnd.n5777 gnd.n5776 19.3944
R14963 gnd.n5776 gnd.n5775 19.3944
R14964 gnd.n5775 gnd.n1166 19.3944
R14965 gnd.n5771 gnd.n1166 19.3944
R14966 gnd.n5771 gnd.n5770 19.3944
R14967 gnd.n5770 gnd.n5769 19.3944
R14968 gnd.n5769 gnd.n1171 19.3944
R14969 gnd.n5765 gnd.n1171 19.3944
R14970 gnd.n5765 gnd.n5764 19.3944
R14971 gnd.n5764 gnd.n5763 19.3944
R14972 gnd.n5763 gnd.n1176 19.3944
R14973 gnd.n5759 gnd.n1176 19.3944
R14974 gnd.n5759 gnd.n5758 19.3944
R14975 gnd.n5758 gnd.n5757 19.3944
R14976 gnd.n5757 gnd.n1181 19.3944
R14977 gnd.n5753 gnd.n1181 19.3944
R14978 gnd.n5753 gnd.n5752 19.3944
R14979 gnd.n5752 gnd.n5751 19.3944
R14980 gnd.n5751 gnd.n1186 19.3944
R14981 gnd.n5747 gnd.n1186 19.3944
R14982 gnd.n5747 gnd.n5746 19.3944
R14983 gnd.n5746 gnd.n5745 19.3944
R14984 gnd.n5745 gnd.n1191 19.3944
R14985 gnd.n5741 gnd.n1191 19.3944
R14986 gnd.n5741 gnd.n5740 19.3944
R14987 gnd.n5740 gnd.n5739 19.3944
R14988 gnd.n5739 gnd.n1196 19.3944
R14989 gnd.n5735 gnd.n1196 19.3944
R14990 gnd.n5735 gnd.n5734 19.3944
R14991 gnd.n5734 gnd.n5733 19.3944
R14992 gnd.n5733 gnd.n1201 19.3944
R14993 gnd.n5729 gnd.n1201 19.3944
R14994 gnd.n5729 gnd.n5728 19.3944
R14995 gnd.n5728 gnd.n5727 19.3944
R14996 gnd.n5727 gnd.n1206 19.3944
R14997 gnd.n5723 gnd.n1206 19.3944
R14998 gnd.n5723 gnd.n5722 19.3944
R14999 gnd.n5722 gnd.n5721 19.3944
R15000 gnd.n5721 gnd.n1211 19.3944
R15001 gnd.n4455 gnd.n1845 19.3944
R15002 gnd.n4474 gnd.n1845 19.3944
R15003 gnd.n4475 gnd.n4474 19.3944
R15004 gnd.n1944 gnd.n1918 19.3944
R15005 gnd.n1948 gnd.n1918 19.3944
R15006 gnd.n1949 gnd.n1948 19.3944
R15007 gnd.n1952 gnd.n1949 19.3944
R15008 gnd.n1952 gnd.n1914 19.3944
R15009 gnd.n4381 gnd.n1914 19.3944
R15010 gnd.n4382 gnd.n4381 19.3944
R15011 gnd.n4385 gnd.n4382 19.3944
R15012 gnd.n4385 gnd.n1909 19.3944
R15013 gnd.n4393 gnd.n1909 19.3944
R15014 gnd.n4396 gnd.n4393 19.3944
R15015 gnd.n4396 gnd.n1903 19.3944
R15016 gnd.n4405 gnd.n1903 19.3944
R15017 gnd.n4408 gnd.n4405 19.3944
R15018 gnd.n4408 gnd.n1897 19.3944
R15019 gnd.n4417 gnd.n1897 19.3944
R15020 gnd.n4420 gnd.n4417 19.3944
R15021 gnd.n4420 gnd.n1891 19.3944
R15022 gnd.n4429 gnd.n1891 19.3944
R15023 gnd.n4432 gnd.n4429 19.3944
R15024 gnd.n4432 gnd.n1885 19.3944
R15025 gnd.n4441 gnd.n1885 19.3944
R15026 gnd.n4445 gnd.n4441 19.3944
R15027 gnd.n4445 gnd.n4444 19.3944
R15028 gnd.n5584 gnd.n5478 19.3944
R15029 gnd.n5584 gnd.n5583 19.3944
R15030 gnd.n5583 gnd.n5481 19.3944
R15031 gnd.n5576 gnd.n5481 19.3944
R15032 gnd.n5576 gnd.n5575 19.3944
R15033 gnd.n5575 gnd.n5491 19.3944
R15034 gnd.n5568 gnd.n5491 19.3944
R15035 gnd.n5568 gnd.n5567 19.3944
R15036 gnd.n5567 gnd.n5501 19.3944
R15037 gnd.n5560 gnd.n5501 19.3944
R15038 gnd.n5560 gnd.n5559 19.3944
R15039 gnd.n5559 gnd.n5511 19.3944
R15040 gnd.n5552 gnd.n5511 19.3944
R15041 gnd.n5552 gnd.n5551 19.3944
R15042 gnd.n5551 gnd.n5521 19.3944
R15043 gnd.n5544 gnd.n5521 19.3944
R15044 gnd.n5359 gnd.n5355 19.3944
R15045 gnd.n5359 gnd.n5358 19.3944
R15046 gnd.n5358 gnd.n5353 19.3944
R15047 gnd.n5382 gnd.n5353 19.3944
R15048 gnd.n5383 gnd.n5382 19.3944
R15049 gnd.n5384 gnd.n5383 19.3944
R15050 gnd.n5384 gnd.n5348 19.3944
R15051 gnd.n5410 gnd.n5348 19.3944
R15052 gnd.n5411 gnd.n5410 19.3944
R15053 gnd.n5412 gnd.n5411 19.3944
R15054 gnd.n5413 gnd.n5412 19.3944
R15055 gnd.n5415 gnd.n5413 19.3944
R15056 gnd.n5415 gnd.n388 19.3944
R15057 gnd.n6724 gnd.n388 19.3944
R15058 gnd.n6725 gnd.n6724 19.3944
R15059 gnd.n6725 gnd.n360 19.3944
R15060 gnd.n6756 gnd.n360 19.3944
R15061 gnd.n6757 gnd.n6756 19.3944
R15062 gnd.n6759 gnd.n6757 19.3944
R15063 gnd.n6760 gnd.n6759 19.3944
R15064 gnd.n6760 gnd.n334 19.3944
R15065 gnd.n6795 gnd.n334 19.3944
R15066 gnd.n6798 gnd.n6795 19.3944
R15067 gnd.n6798 gnd.n6797 19.3944
R15068 gnd.n6797 gnd.n315 19.3944
R15069 gnd.n6818 gnd.n315 19.3944
R15070 gnd.n6819 gnd.n6818 19.3944
R15071 gnd.n6819 gnd.n309 19.3944
R15072 gnd.n6828 gnd.n309 19.3944
R15073 gnd.n6829 gnd.n6828 19.3944
R15074 gnd.n6831 gnd.n6829 19.3944
R15075 gnd.n6832 gnd.n6831 19.3944
R15076 gnd.n6835 gnd.n6832 19.3944
R15077 gnd.n6836 gnd.n6835 19.3944
R15078 gnd.n6838 gnd.n6836 19.3944
R15079 gnd.n6839 gnd.n6838 19.3944
R15080 gnd.n6842 gnd.n6839 19.3944
R15081 gnd.n6843 gnd.n6842 19.3944
R15082 gnd.n6845 gnd.n6843 19.3944
R15083 gnd.n6846 gnd.n6845 19.3944
R15084 gnd.n6849 gnd.n6846 19.3944
R15085 gnd.n6850 gnd.n6849 19.3944
R15086 gnd.n6971 gnd.n6850 19.3944
R15087 gnd.n6972 gnd.n6971 19.3944
R15088 gnd.n6975 gnd.n6972 19.3944
R15089 gnd.n6976 gnd.n6975 19.3944
R15090 gnd.n6978 gnd.n6976 19.3944
R15091 gnd.n6979 gnd.n6978 19.3944
R15092 gnd.n6982 gnd.n6979 19.3944
R15093 gnd.n6983 gnd.n6982 19.3944
R15094 gnd.n6985 gnd.n6983 19.3944
R15095 gnd.n6986 gnd.n6985 19.3944
R15096 gnd.n6989 gnd.n6986 19.3944
R15097 gnd.n7032 gnd.n285 19.3944
R15098 gnd.n7032 gnd.n7029 19.3944
R15099 gnd.n7029 gnd.n7026 19.3944
R15100 gnd.n7026 gnd.n7025 19.3944
R15101 gnd.n7025 gnd.n7022 19.3944
R15102 gnd.n7022 gnd.n7021 19.3944
R15103 gnd.n7021 gnd.n7018 19.3944
R15104 gnd.n7018 gnd.n7017 19.3944
R15105 gnd.n7017 gnd.n7014 19.3944
R15106 gnd.n7014 gnd.n7013 19.3944
R15107 gnd.n7013 gnd.n7010 19.3944
R15108 gnd.n7010 gnd.n7009 19.3944
R15109 gnd.n7009 gnd.n7006 19.3944
R15110 gnd.n7006 gnd.n7005 19.3944
R15111 gnd.n7005 gnd.n7002 19.3944
R15112 gnd.n7002 gnd.n7001 19.3944
R15113 gnd.n7001 gnd.n6998 19.3944
R15114 gnd.n6998 gnd.n6997 19.3944
R15115 gnd.n7075 gnd.n7072 19.3944
R15116 gnd.n7072 gnd.n7071 19.3944
R15117 gnd.n7071 gnd.n7068 19.3944
R15118 gnd.n7068 gnd.n7067 19.3944
R15119 gnd.n7067 gnd.n7064 19.3944
R15120 gnd.n7064 gnd.n7063 19.3944
R15121 gnd.n7063 gnd.n7060 19.3944
R15122 gnd.n7060 gnd.n7059 19.3944
R15123 gnd.n7059 gnd.n7056 19.3944
R15124 gnd.n7056 gnd.n7055 19.3944
R15125 gnd.n7055 gnd.n7052 19.3944
R15126 gnd.n7052 gnd.n7051 19.3944
R15127 gnd.n7051 gnd.n7048 19.3944
R15128 gnd.n7048 gnd.n7047 19.3944
R15129 gnd.n7047 gnd.n7044 19.3944
R15130 gnd.n7044 gnd.n7043 19.3944
R15131 gnd.n7043 gnd.n7040 19.3944
R15132 gnd.n7040 gnd.n7039 19.3944
R15133 gnd.n7113 gnd.n209 19.3944
R15134 gnd.n7108 gnd.n209 19.3944
R15135 gnd.n7108 gnd.n7107 19.3944
R15136 gnd.n7107 gnd.n7106 19.3944
R15137 gnd.n7106 gnd.n7103 19.3944
R15138 gnd.n7103 gnd.n7102 19.3944
R15139 gnd.n7102 gnd.n7099 19.3944
R15140 gnd.n7099 gnd.n7098 19.3944
R15141 gnd.n7098 gnd.n7095 19.3944
R15142 gnd.n7095 gnd.n7094 19.3944
R15143 gnd.n7094 gnd.n7091 19.3944
R15144 gnd.n7091 gnd.n7090 19.3944
R15145 gnd.n7090 gnd.n7087 19.3944
R15146 gnd.n7087 gnd.n7086 19.3944
R15147 gnd.n7086 gnd.n7083 19.3944
R15148 gnd.n7083 gnd.n7082 19.3944
R15149 gnd.n7082 gnd.n7079 19.3944
R15150 gnd.n5297 gnd.n5295 19.3944
R15151 gnd.n5297 gnd.n5293 19.3944
R15152 gnd.n5465 gnd.n5293 19.3944
R15153 gnd.n5465 gnd.n5464 19.3944
R15154 gnd.n5464 gnd.n5463 19.3944
R15155 gnd.n5463 gnd.n5303 19.3944
R15156 gnd.n5453 gnd.n5303 19.3944
R15157 gnd.n5453 gnd.n5452 19.3944
R15158 gnd.n5452 gnd.n5451 19.3944
R15159 gnd.n5451 gnd.n5325 19.3944
R15160 gnd.n5441 gnd.n5325 19.3944
R15161 gnd.n5441 gnd.n377 19.3944
R15162 gnd.n6737 gnd.n377 19.3944
R15163 gnd.n6737 gnd.n375 19.3944
R15164 gnd.n6743 gnd.n375 19.3944
R15165 gnd.n6743 gnd.n6742 19.3944
R15166 gnd.n6742 gnd.n349 19.3944
R15167 gnd.n6771 gnd.n349 19.3944
R15168 gnd.n6771 gnd.n347 19.3944
R15169 gnd.n6777 gnd.n347 19.3944
R15170 gnd.n6777 gnd.n6776 19.3944
R15171 gnd.n6776 gnd.n327 19.3944
R15172 gnd.n6804 gnd.n327 19.3944
R15173 gnd.n6804 gnd.n325 19.3944
R15174 gnd.n6811 gnd.n325 19.3944
R15175 gnd.n6811 gnd.n6810 19.3944
R15176 gnd.n6810 gnd.n90 19.3944
R15177 gnd.n7189 gnd.n90 19.3944
R15178 gnd.n7189 gnd.n7188 19.3944
R15179 gnd.n7188 gnd.n7187 19.3944
R15180 gnd.n7187 gnd.n94 19.3944
R15181 gnd.n7177 gnd.n94 19.3944
R15182 gnd.n7177 gnd.n7176 19.3944
R15183 gnd.n7176 gnd.n7175 19.3944
R15184 gnd.n7175 gnd.n115 19.3944
R15185 gnd.n7165 gnd.n115 19.3944
R15186 gnd.n7165 gnd.n7164 19.3944
R15187 gnd.n7164 gnd.n7163 19.3944
R15188 gnd.n7163 gnd.n134 19.3944
R15189 gnd.n7153 gnd.n134 19.3944
R15190 gnd.n7153 gnd.n7152 19.3944
R15191 gnd.n7152 gnd.n7151 19.3944
R15192 gnd.n7151 gnd.n153 19.3944
R15193 gnd.n7141 gnd.n153 19.3944
R15194 gnd.n7141 gnd.n7140 19.3944
R15195 gnd.n7140 gnd.n7139 19.3944
R15196 gnd.n7139 gnd.n172 19.3944
R15197 gnd.n7129 gnd.n172 19.3944
R15198 gnd.n7129 gnd.n7128 19.3944
R15199 gnd.n7128 gnd.n7127 19.3944
R15200 gnd.n7127 gnd.n191 19.3944
R15201 gnd.n7117 gnd.n191 19.3944
R15202 gnd.n7117 gnd.n7116 19.3944
R15203 gnd.n5705 gnd.n5704 19.3944
R15204 gnd.n5704 gnd.n5703 19.3944
R15205 gnd.n5703 gnd.n5702 19.3944
R15206 gnd.n5702 gnd.n5700 19.3944
R15207 gnd.n5700 gnd.n5697 19.3944
R15208 gnd.n5697 gnd.n5696 19.3944
R15209 gnd.n5696 gnd.n5693 19.3944
R15210 gnd.n5693 gnd.n5692 19.3944
R15211 gnd.n5692 gnd.n5689 19.3944
R15212 gnd.n5689 gnd.n5688 19.3944
R15213 gnd.n5688 gnd.n5685 19.3944
R15214 gnd.n5685 gnd.n5684 19.3944
R15215 gnd.n5684 gnd.n5681 19.3944
R15216 gnd.n5681 gnd.n5680 19.3944
R15217 gnd.n5680 gnd.n5677 19.3944
R15218 gnd.n5677 gnd.n5676 19.3944
R15219 gnd.n5676 gnd.n5673 19.3944
R15220 gnd.n5671 gnd.n5668 19.3944
R15221 gnd.n5668 gnd.n5667 19.3944
R15222 gnd.n5667 gnd.n5664 19.3944
R15223 gnd.n5664 gnd.n5663 19.3944
R15224 gnd.n5663 gnd.n5660 19.3944
R15225 gnd.n5660 gnd.n5659 19.3944
R15226 gnd.n5659 gnd.n5656 19.3944
R15227 gnd.n5654 gnd.n5651 19.3944
R15228 gnd.n5651 gnd.n5650 19.3944
R15229 gnd.n5650 gnd.n5647 19.3944
R15230 gnd.n5647 gnd.n5646 19.3944
R15231 gnd.n5646 gnd.n5643 19.3944
R15232 gnd.n5643 gnd.n5642 19.3944
R15233 gnd.n5642 gnd.n5639 19.3944
R15234 gnd.n5639 gnd.n5638 19.3944
R15235 gnd.n5634 gnd.n5631 19.3944
R15236 gnd.n5631 gnd.n5630 19.3944
R15237 gnd.n5630 gnd.n5627 19.3944
R15238 gnd.n5627 gnd.n5626 19.3944
R15239 gnd.n5626 gnd.n5623 19.3944
R15240 gnd.n5623 gnd.n5622 19.3944
R15241 gnd.n5622 gnd.n5619 19.3944
R15242 gnd.n5619 gnd.n5618 19.3944
R15243 gnd.n5618 gnd.n5615 19.3944
R15244 gnd.n5615 gnd.n5614 19.3944
R15245 gnd.n5614 gnd.n5611 19.3944
R15246 gnd.n5611 gnd.n5610 19.3944
R15247 gnd.n5610 gnd.n5607 19.3944
R15248 gnd.n5607 gnd.n5606 19.3944
R15249 gnd.n5606 gnd.n5603 19.3944
R15250 gnd.n5603 gnd.n5602 19.3944
R15251 gnd.n5602 gnd.n5599 19.3944
R15252 gnd.n5599 gnd.n5598 19.3944
R15253 gnd.n6907 gnd.n6905 19.3944
R15254 gnd.n6910 gnd.n6907 19.3944
R15255 gnd.n6913 gnd.n6910 19.3944
R15256 gnd.n6916 gnd.n6913 19.3944
R15257 gnd.n6916 gnd.n6903 19.3944
R15258 gnd.n6920 gnd.n6903 19.3944
R15259 gnd.n6923 gnd.n6920 19.3944
R15260 gnd.n6926 gnd.n6923 19.3944
R15261 gnd.n6926 gnd.n6901 19.3944
R15262 gnd.n6930 gnd.n6901 19.3944
R15263 gnd.n6933 gnd.n6930 19.3944
R15264 gnd.n6936 gnd.n6933 19.3944
R15265 gnd.n6936 gnd.n6899 19.3944
R15266 gnd.n6940 gnd.n6899 19.3944
R15267 gnd.n6943 gnd.n6940 19.3944
R15268 gnd.n6946 gnd.n6943 19.3944
R15269 gnd.n5371 gnd.n5370 19.3944
R15270 gnd.n5374 gnd.n5371 19.3944
R15271 gnd.n5374 gnd.n5367 19.3944
R15272 gnd.n5378 gnd.n5367 19.3944
R15273 gnd.n5378 gnd.n5352 19.3944
R15274 gnd.n5402 gnd.n5352 19.3944
R15275 gnd.n5402 gnd.n5350 19.3944
R15276 gnd.n5406 gnd.n5350 19.3944
R15277 gnd.n5406 gnd.n5344 19.3944
R15278 gnd.n5424 gnd.n5344 19.3944
R15279 gnd.n5424 gnd.n5345 19.3944
R15280 gnd.n5420 gnd.n5345 19.3944
R15281 gnd.n5420 gnd.n5419 19.3944
R15282 gnd.n5419 gnd.n368 19.3944
R15283 gnd.n6747 gnd.n368 19.3944
R15284 gnd.n6747 gnd.n365 19.3944
R15285 gnd.n6752 gnd.n365 19.3944
R15286 gnd.n6752 gnd.n366 19.3944
R15287 gnd.n366 gnd.n341 19.3944
R15288 gnd.n6781 gnd.n341 19.3944
R15289 gnd.n6781 gnd.n338 19.3944
R15290 gnd.n6791 gnd.n338 19.3944
R15291 gnd.n6791 gnd.n339 19.3944
R15292 gnd.n6787 gnd.n339 19.3944
R15293 gnd.n6787 gnd.n6786 19.3944
R15294 gnd.n6786 gnd.n81 19.3944
R15295 gnd.n7194 gnd.n81 19.3944
R15296 gnd.n7194 gnd.n7193 19.3944
R15297 gnd.n7193 gnd.n83 19.3944
R15298 gnd.n6857 gnd.n83 19.3944
R15299 gnd.n6862 gnd.n6857 19.3944
R15300 gnd.n6863 gnd.n6862 19.3944
R15301 gnd.n6865 gnd.n6863 19.3944
R15302 gnd.n6865 gnd.n6855 19.3944
R15303 gnd.n6870 gnd.n6855 19.3944
R15304 gnd.n6871 gnd.n6870 19.3944
R15305 gnd.n6873 gnd.n6871 19.3944
R15306 gnd.n6873 gnd.n6853 19.3944
R15307 gnd.n6878 gnd.n6853 19.3944
R15308 gnd.n6879 gnd.n6878 19.3944
R15309 gnd.n6881 gnd.n6879 19.3944
R15310 gnd.n6881 gnd.n6851 19.3944
R15311 gnd.n6967 gnd.n6851 19.3944
R15312 gnd.n6967 gnd.n6966 19.3944
R15313 gnd.n6966 gnd.n6965 19.3944
R15314 gnd.n6965 gnd.n6963 19.3944
R15315 gnd.n6963 gnd.n6962 19.3944
R15316 gnd.n6962 gnd.n6960 19.3944
R15317 gnd.n6960 gnd.n6959 19.3944
R15318 gnd.n6959 gnd.n6957 19.3944
R15319 gnd.n6957 gnd.n6956 19.3944
R15320 gnd.n6956 gnd.n6954 19.3944
R15321 gnd.n6954 gnd.n6953 19.3944
R15322 gnd.n5361 gnd.n5269 19.3944
R15323 gnd.n5363 gnd.n5361 19.3944
R15324 gnd.n5364 gnd.n5363 19.3944
R15325 gnd.n5364 gnd.n5311 19.3944
R15326 gnd.n5459 gnd.n5311 19.3944
R15327 gnd.n5459 gnd.n5458 19.3944
R15328 gnd.n5458 gnd.n5457 19.3944
R15329 gnd.n5457 gnd.n5315 19.3944
R15330 gnd.n5447 gnd.n5315 19.3944
R15331 gnd.n5447 gnd.n5446 19.3944
R15332 gnd.n5446 gnd.n5445 19.3944
R15333 gnd.n5445 gnd.n385 19.3944
R15334 gnd.n6733 gnd.n385 19.3944
R15335 gnd.n6733 gnd.n6732 19.3944
R15336 gnd.n6732 gnd.n6731 19.3944
R15337 gnd.n6731 gnd.n6730 19.3944
R15338 gnd.n6730 gnd.n357 19.3944
R15339 gnd.n6767 gnd.n357 19.3944
R15340 gnd.n6767 gnd.n6766 19.3944
R15341 gnd.n6766 gnd.n6765 19.3944
R15342 gnd.n6765 gnd.n6764 19.3944
R15343 gnd.n6764 gnd.n332 19.3944
R15344 gnd.n6800 gnd.n332 19.3944
R15345 gnd.n6800 gnd.n317 19.3944
R15346 gnd.n6815 gnd.n317 19.3944
R15347 gnd.n6815 gnd.n311 19.3944
R15348 gnd.n6823 gnd.n311 19.3944
R15349 gnd.n6824 gnd.n6823 19.3944
R15350 gnd.n6824 gnd.n100 19.3944
R15351 gnd.n7183 gnd.n100 19.3944
R15352 gnd.n7183 gnd.n7182 19.3944
R15353 gnd.n7182 gnd.n7181 19.3944
R15354 gnd.n7181 gnd.n104 19.3944
R15355 gnd.n7171 gnd.n104 19.3944
R15356 gnd.n7171 gnd.n7170 19.3944
R15357 gnd.n7170 gnd.n7169 19.3944
R15358 gnd.n7169 gnd.n124 19.3944
R15359 gnd.n7159 gnd.n124 19.3944
R15360 gnd.n7159 gnd.n7158 19.3944
R15361 gnd.n7158 gnd.n7157 19.3944
R15362 gnd.n7157 gnd.n142 19.3944
R15363 gnd.n7147 gnd.n142 19.3944
R15364 gnd.n7147 gnd.n7146 19.3944
R15365 gnd.n7146 gnd.n7145 19.3944
R15366 gnd.n7145 gnd.n162 19.3944
R15367 gnd.n7135 gnd.n162 19.3944
R15368 gnd.n7135 gnd.n7134 19.3944
R15369 gnd.n7134 gnd.n7133 19.3944
R15370 gnd.n7133 gnd.n180 19.3944
R15371 gnd.n7123 gnd.n180 19.3944
R15372 gnd.n7123 gnd.n7122 19.3944
R15373 gnd.n7122 gnd.n7121 19.3944
R15374 gnd.n7121 gnd.n200 19.3944
R15375 gnd.n2870 gnd.n2869 19.3944
R15376 gnd.n2869 gnd.n2868 19.3944
R15377 gnd.n2868 gnd.n2867 19.3944
R15378 gnd.n2867 gnd.n2865 19.3944
R15379 gnd.n2865 gnd.n2862 19.3944
R15380 gnd.n2862 gnd.n2861 19.3944
R15381 gnd.n2861 gnd.n2858 19.3944
R15382 gnd.n2858 gnd.n2857 19.3944
R15383 gnd.n2857 gnd.n2854 19.3944
R15384 gnd.n2854 gnd.n2853 19.3944
R15385 gnd.n2853 gnd.n2850 19.3944
R15386 gnd.n2850 gnd.n2849 19.3944
R15387 gnd.n2849 gnd.n2846 19.3944
R15388 gnd.n2846 gnd.n2845 19.3944
R15389 gnd.n2845 gnd.n2842 19.3944
R15390 gnd.n2842 gnd.n2841 19.3944
R15391 gnd.n2841 gnd.n2838 19.3944
R15392 gnd.n2838 gnd.n2837 19.3944
R15393 gnd.n2837 gnd.n2834 19.3944
R15394 gnd.n2834 gnd.n2833 19.3944
R15395 gnd.n2833 gnd.n2830 19.3944
R15396 gnd.n2830 gnd.n2829 19.3944
R15397 gnd.n2826 gnd.n2825 19.3944
R15398 gnd.n2825 gnd.n2781 19.3944
R15399 gnd.n2876 gnd.n2781 19.3944
R15400 gnd.n3642 gnd.n3641 19.3944
R15401 gnd.n3641 gnd.n3638 19.3944
R15402 gnd.n3638 gnd.n3637 19.3944
R15403 gnd.n3687 gnd.n3686 19.3944
R15404 gnd.n3686 gnd.n3685 19.3944
R15405 gnd.n3685 gnd.n3682 19.3944
R15406 gnd.n3682 gnd.n3681 19.3944
R15407 gnd.n3681 gnd.n3678 19.3944
R15408 gnd.n3678 gnd.n3677 19.3944
R15409 gnd.n3677 gnd.n3674 19.3944
R15410 gnd.n3674 gnd.n3673 19.3944
R15411 gnd.n3673 gnd.n3670 19.3944
R15412 gnd.n3670 gnd.n3669 19.3944
R15413 gnd.n3669 gnd.n3666 19.3944
R15414 gnd.n3666 gnd.n3665 19.3944
R15415 gnd.n3665 gnd.n3662 19.3944
R15416 gnd.n3662 gnd.n3661 19.3944
R15417 gnd.n3661 gnd.n3658 19.3944
R15418 gnd.n3658 gnd.n3657 19.3944
R15419 gnd.n3657 gnd.n3654 19.3944
R15420 gnd.n3654 gnd.n3653 19.3944
R15421 gnd.n3653 gnd.n3650 19.3944
R15422 gnd.n3650 gnd.n3649 19.3944
R15423 gnd.n3649 gnd.n3646 19.3944
R15424 gnd.n3646 gnd.n3645 19.3944
R15425 gnd.n2969 gnd.n2678 19.3944
R15426 gnd.n2979 gnd.n2678 19.3944
R15427 gnd.n2980 gnd.n2979 19.3944
R15428 gnd.n2980 gnd.n2659 19.3944
R15429 gnd.n3000 gnd.n2659 19.3944
R15430 gnd.n3000 gnd.n2651 19.3944
R15431 gnd.n3010 gnd.n2651 19.3944
R15432 gnd.n3011 gnd.n3010 19.3944
R15433 gnd.n3012 gnd.n3011 19.3944
R15434 gnd.n3012 gnd.n2634 19.3944
R15435 gnd.n3029 gnd.n2634 19.3944
R15436 gnd.n3032 gnd.n3029 19.3944
R15437 gnd.n3032 gnd.n3031 19.3944
R15438 gnd.n3031 gnd.n2607 19.3944
R15439 gnd.n3071 gnd.n2607 19.3944
R15440 gnd.n3071 gnd.n2604 19.3944
R15441 gnd.n3077 gnd.n2604 19.3944
R15442 gnd.n3078 gnd.n3077 19.3944
R15443 gnd.n3078 gnd.n2602 19.3944
R15444 gnd.n3084 gnd.n2602 19.3944
R15445 gnd.n3087 gnd.n3084 19.3944
R15446 gnd.n3089 gnd.n3087 19.3944
R15447 gnd.n3095 gnd.n3089 19.3944
R15448 gnd.n3095 gnd.n3094 19.3944
R15449 gnd.n3094 gnd.n2461 19.3944
R15450 gnd.n3161 gnd.n2461 19.3944
R15451 gnd.n3162 gnd.n3161 19.3944
R15452 gnd.n3162 gnd.n2454 19.3944
R15453 gnd.n3173 gnd.n2454 19.3944
R15454 gnd.n3174 gnd.n3173 19.3944
R15455 gnd.n3174 gnd.n2437 19.3944
R15456 gnd.n2437 gnd.n2435 19.3944
R15457 gnd.n3198 gnd.n2435 19.3944
R15458 gnd.n3199 gnd.n3198 19.3944
R15459 gnd.n3199 gnd.n2406 19.3944
R15460 gnd.n3246 gnd.n2406 19.3944
R15461 gnd.n3247 gnd.n3246 19.3944
R15462 gnd.n3247 gnd.n2399 19.3944
R15463 gnd.n3258 gnd.n2399 19.3944
R15464 gnd.n3259 gnd.n3258 19.3944
R15465 gnd.n3259 gnd.n2382 19.3944
R15466 gnd.n2382 gnd.n2380 19.3944
R15467 gnd.n3283 gnd.n2380 19.3944
R15468 gnd.n3284 gnd.n3283 19.3944
R15469 gnd.n3284 gnd.n2352 19.3944
R15470 gnd.n3335 gnd.n2352 19.3944
R15471 gnd.n3336 gnd.n3335 19.3944
R15472 gnd.n3336 gnd.n2345 19.3944
R15473 gnd.n3603 gnd.n2345 19.3944
R15474 gnd.n3604 gnd.n3603 19.3944
R15475 gnd.n3604 gnd.n2326 19.3944
R15476 gnd.n3629 gnd.n2326 19.3944
R15477 gnd.n3629 gnd.n2327 19.3944
R15478 gnd.n2960 gnd.n2959 19.3944
R15479 gnd.n2959 gnd.n2692 19.3944
R15480 gnd.n2715 gnd.n2692 19.3944
R15481 gnd.n2718 gnd.n2715 19.3944
R15482 gnd.n2718 gnd.n2711 19.3944
R15483 gnd.n2722 gnd.n2711 19.3944
R15484 gnd.n2725 gnd.n2722 19.3944
R15485 gnd.n2728 gnd.n2725 19.3944
R15486 gnd.n2728 gnd.n2709 19.3944
R15487 gnd.n2732 gnd.n2709 19.3944
R15488 gnd.n2735 gnd.n2732 19.3944
R15489 gnd.n2738 gnd.n2735 19.3944
R15490 gnd.n2738 gnd.n2707 19.3944
R15491 gnd.n2742 gnd.n2707 19.3944
R15492 gnd.n2965 gnd.n2964 19.3944
R15493 gnd.n2964 gnd.n2668 19.3944
R15494 gnd.n2990 gnd.n2668 19.3944
R15495 gnd.n2990 gnd.n2666 19.3944
R15496 gnd.n2996 gnd.n2666 19.3944
R15497 gnd.n2996 gnd.n2995 19.3944
R15498 gnd.n2995 gnd.n2640 19.3944
R15499 gnd.n3020 gnd.n2640 19.3944
R15500 gnd.n3020 gnd.n2638 19.3944
R15501 gnd.n3024 gnd.n2638 19.3944
R15502 gnd.n3024 gnd.n2618 19.3944
R15503 gnd.n3051 gnd.n2618 19.3944
R15504 gnd.n3051 gnd.n2616 19.3944
R15505 gnd.n3061 gnd.n2616 19.3944
R15506 gnd.n3061 gnd.n3060 19.3944
R15507 gnd.n3060 gnd.n3059 19.3944
R15508 gnd.n3059 gnd.n2565 19.3944
R15509 gnd.n3109 gnd.n2565 19.3944
R15510 gnd.n3109 gnd.n3108 19.3944
R15511 gnd.n3108 gnd.n3107 19.3944
R15512 gnd.n3107 gnd.n2569 19.3944
R15513 gnd.n2589 gnd.n2569 19.3944
R15514 gnd.n2589 gnd.n2471 19.3944
R15515 gnd.n3146 gnd.n2471 19.3944
R15516 gnd.n3146 gnd.n2469 19.3944
R15517 gnd.n3152 gnd.n2469 19.3944
R15518 gnd.n3152 gnd.n3151 19.3944
R15519 gnd.n3151 gnd.n2444 19.3944
R15520 gnd.n3186 gnd.n2444 19.3944
R15521 gnd.n3186 gnd.n2442 19.3944
R15522 gnd.n3192 gnd.n2442 19.3944
R15523 gnd.n3192 gnd.n3191 19.3944
R15524 gnd.n3191 gnd.n2417 19.3944
R15525 gnd.n3231 gnd.n2417 19.3944
R15526 gnd.n3231 gnd.n2415 19.3944
R15527 gnd.n3237 gnd.n2415 19.3944
R15528 gnd.n3237 gnd.n3236 19.3944
R15529 gnd.n3236 gnd.n2389 19.3944
R15530 gnd.n3271 gnd.n2389 19.3944
R15531 gnd.n3271 gnd.n2387 19.3944
R15532 gnd.n3277 gnd.n2387 19.3944
R15533 gnd.n3277 gnd.n3276 19.3944
R15534 gnd.n3276 gnd.n2362 19.3944
R15535 gnd.n3320 gnd.n2362 19.3944
R15536 gnd.n3320 gnd.n2360 19.3944
R15537 gnd.n3326 gnd.n2360 19.3944
R15538 gnd.n3326 gnd.n3325 19.3944
R15539 gnd.n3325 gnd.n2335 19.3944
R15540 gnd.n3614 gnd.n2335 19.3944
R15541 gnd.n3614 gnd.n2333 19.3944
R15542 gnd.n3622 gnd.n2333 19.3944
R15543 gnd.n3622 gnd.n3621 19.3944
R15544 gnd.n3621 gnd.n3620 19.3944
R15545 gnd.n3723 gnd.n3722 19.3944
R15546 gnd.n3722 gnd.n2273 19.3944
R15547 gnd.n3718 gnd.n2273 19.3944
R15548 gnd.n3718 gnd.n3715 19.3944
R15549 gnd.n3715 gnd.n3712 19.3944
R15550 gnd.n3712 gnd.n3711 19.3944
R15551 gnd.n3711 gnd.n3708 19.3944
R15552 gnd.n3708 gnd.n3707 19.3944
R15553 gnd.n3707 gnd.n3704 19.3944
R15554 gnd.n3704 gnd.n3703 19.3944
R15555 gnd.n3703 gnd.n3700 19.3944
R15556 gnd.n3700 gnd.n3699 19.3944
R15557 gnd.n3699 gnd.n3696 19.3944
R15558 gnd.n3696 gnd.n3695 19.3944
R15559 gnd.n2880 gnd.n2779 19.3944
R15560 gnd.n2880 gnd.n2770 19.3944
R15561 gnd.n2893 gnd.n2770 19.3944
R15562 gnd.n2893 gnd.n2768 19.3944
R15563 gnd.n2897 gnd.n2768 19.3944
R15564 gnd.n2897 gnd.n2758 19.3944
R15565 gnd.n2909 gnd.n2758 19.3944
R15566 gnd.n2909 gnd.n2756 19.3944
R15567 gnd.n2943 gnd.n2756 19.3944
R15568 gnd.n2943 gnd.n2942 19.3944
R15569 gnd.n2942 gnd.n2941 19.3944
R15570 gnd.n2941 gnd.n2940 19.3944
R15571 gnd.n2940 gnd.n2937 19.3944
R15572 gnd.n2937 gnd.n2936 19.3944
R15573 gnd.n2936 gnd.n2935 19.3944
R15574 gnd.n2935 gnd.n2933 19.3944
R15575 gnd.n2933 gnd.n2932 19.3944
R15576 gnd.n2932 gnd.n2929 19.3944
R15577 gnd.n2929 gnd.n2928 19.3944
R15578 gnd.n2928 gnd.n2927 19.3944
R15579 gnd.n2927 gnd.n2925 19.3944
R15580 gnd.n2925 gnd.n2624 19.3944
R15581 gnd.n3040 gnd.n2624 19.3944
R15582 gnd.n3040 gnd.n2622 19.3944
R15583 gnd.n3046 gnd.n2622 19.3944
R15584 gnd.n3046 gnd.n3045 19.3944
R15585 gnd.n3045 gnd.n2546 19.3944
R15586 gnd.n3120 gnd.n2546 19.3944
R15587 gnd.n3120 gnd.n2547 19.3944
R15588 gnd.n2594 gnd.n2593 19.3944
R15589 gnd.n2597 gnd.n2596 19.3944
R15590 gnd.n2584 gnd.n2583 19.3944
R15591 gnd.n3139 gnd.n2476 19.3944
R15592 gnd.n3139 gnd.n3138 19.3944
R15593 gnd.n3138 gnd.n3137 19.3944
R15594 gnd.n3137 gnd.n3135 19.3944
R15595 gnd.n3135 gnd.n3134 19.3944
R15596 gnd.n3134 gnd.n3132 19.3944
R15597 gnd.n3132 gnd.n3131 19.3944
R15598 gnd.n3131 gnd.n2425 19.3944
R15599 gnd.n3207 gnd.n2425 19.3944
R15600 gnd.n3207 gnd.n2423 19.3944
R15601 gnd.n3226 gnd.n2423 19.3944
R15602 gnd.n3226 gnd.n3225 19.3944
R15603 gnd.n3225 gnd.n3224 19.3944
R15604 gnd.n3224 gnd.n3222 19.3944
R15605 gnd.n3222 gnd.n3221 19.3944
R15606 gnd.n3221 gnd.n3219 19.3944
R15607 gnd.n3219 gnd.n3218 19.3944
R15608 gnd.n3218 gnd.n2369 19.3944
R15609 gnd.n3292 gnd.n2369 19.3944
R15610 gnd.n3292 gnd.n2367 19.3944
R15611 gnd.n3315 gnd.n2367 19.3944
R15612 gnd.n3315 gnd.n3314 19.3944
R15613 gnd.n3314 gnd.n3313 19.3944
R15614 gnd.n3313 gnd.n3310 19.3944
R15615 gnd.n3310 gnd.n3309 19.3944
R15616 gnd.n3309 gnd.n3307 19.3944
R15617 gnd.n3307 gnd.n3306 19.3944
R15618 gnd.n3306 gnd.n3304 19.3944
R15619 gnd.n3304 gnd.n2320 19.3944
R15620 gnd.n2885 gnd.n2775 19.3944
R15621 gnd.n2885 gnd.n2773 19.3944
R15622 gnd.n2889 gnd.n2773 19.3944
R15623 gnd.n2889 gnd.n2764 19.3944
R15624 gnd.n2901 gnd.n2764 19.3944
R15625 gnd.n2901 gnd.n2762 19.3944
R15626 gnd.n2905 gnd.n2762 19.3944
R15627 gnd.n2905 gnd.n2751 19.3944
R15628 gnd.n2947 gnd.n2751 19.3944
R15629 gnd.n2947 gnd.n2705 19.3944
R15630 gnd.n2953 gnd.n2705 19.3944
R15631 gnd.n2953 gnd.n2952 19.3944
R15632 gnd.n2952 gnd.n2683 19.3944
R15633 gnd.n2974 gnd.n2683 19.3944
R15634 gnd.n2974 gnd.n2676 19.3944
R15635 gnd.n2985 gnd.n2676 19.3944
R15636 gnd.n2985 gnd.n2984 19.3944
R15637 gnd.n2984 gnd.n2657 19.3944
R15638 gnd.n3005 gnd.n2657 19.3944
R15639 gnd.n3005 gnd.n2647 19.3944
R15640 gnd.n3015 gnd.n2647 19.3944
R15641 gnd.n3015 gnd.n2630 19.3944
R15642 gnd.n3036 gnd.n2630 19.3944
R15643 gnd.n3036 gnd.n3035 19.3944
R15644 gnd.n3035 gnd.n2609 19.3944
R15645 gnd.n3066 gnd.n2609 19.3944
R15646 gnd.n3066 gnd.n2554 19.3944
R15647 gnd.n3116 gnd.n2554 19.3944
R15648 gnd.n3116 gnd.n3115 19.3944
R15649 gnd.n3115 gnd.n3114 19.3944
R15650 gnd.n3114 gnd.n2558 19.3944
R15651 gnd.n2576 gnd.n2558 19.3944
R15652 gnd.n3102 gnd.n2576 19.3944
R15653 gnd.n3102 gnd.n3101 19.3944
R15654 gnd.n3101 gnd.n3100 19.3944
R15655 gnd.n3100 gnd.n2580 19.3944
R15656 gnd.n2580 gnd.n2463 19.3944
R15657 gnd.n3157 gnd.n2463 19.3944
R15658 gnd.n3157 gnd.n2456 19.3944
R15659 gnd.n3168 gnd.n2456 19.3944
R15660 gnd.n3168 gnd.n2452 19.3944
R15661 gnd.n3181 gnd.n2452 19.3944
R15662 gnd.n3181 gnd.n3180 19.3944
R15663 gnd.n3180 gnd.n2431 19.3944
R15664 gnd.n3203 gnd.n2431 19.3944
R15665 gnd.n3203 gnd.n3202 19.3944
R15666 gnd.n3202 gnd.n2408 19.3944
R15667 gnd.n3242 gnd.n2408 19.3944
R15668 gnd.n3242 gnd.n2401 19.3944
R15669 gnd.n3253 gnd.n2401 19.3944
R15670 gnd.n3253 gnd.n2397 19.3944
R15671 gnd.n3266 gnd.n2397 19.3944
R15672 gnd.n3266 gnd.n3265 19.3944
R15673 gnd.n3265 gnd.n2376 19.3944
R15674 gnd.n3288 gnd.n2376 19.3944
R15675 gnd.n3288 gnd.n3287 19.3944
R15676 gnd.n3287 gnd.n2354 19.3944
R15677 gnd.n3331 gnd.n2354 19.3944
R15678 gnd.n3331 gnd.n2347 19.3944
R15679 gnd.n3342 gnd.n2347 19.3944
R15680 gnd.n3342 gnd.n2343 19.3944
R15681 gnd.n3609 gnd.n2343 19.3944
R15682 gnd.n3609 gnd.n3608 19.3944
R15683 gnd.n3608 gnd.n2324 19.3944
R15684 gnd.n3632 gnd.n2324 19.3944
R15685 gnd.n4390 gnd.n4388 19.3944
R15686 gnd.n4390 gnd.n1905 19.3944
R15687 gnd.n4399 gnd.n1905 19.3944
R15688 gnd.n4402 gnd.n4399 19.3944
R15689 gnd.n4402 gnd.n1901 19.3944
R15690 gnd.n4411 gnd.n1901 19.3944
R15691 gnd.n4414 gnd.n4411 19.3944
R15692 gnd.n4414 gnd.n1893 19.3944
R15693 gnd.n4423 gnd.n1893 19.3944
R15694 gnd.n4426 gnd.n4423 19.3944
R15695 gnd.n4426 gnd.n1889 19.3944
R15696 gnd.n4435 gnd.n1889 19.3944
R15697 gnd.n4438 gnd.n4435 19.3944
R15698 gnd.n4438 gnd.n1881 19.3944
R15699 gnd.n4448 gnd.n1881 19.3944
R15700 gnd.n4451 gnd.n4448 19.3944
R15701 gnd.n4044 gnd.n4043 19.3944
R15702 gnd.n4045 gnd.n4044 19.3944
R15703 gnd.n4045 gnd.n2226 19.3944
R15704 gnd.n4063 gnd.n2226 19.3944
R15705 gnd.n4064 gnd.n4063 19.3944
R15706 gnd.n4065 gnd.n4064 19.3944
R15707 gnd.n4065 gnd.n2208 19.3944
R15708 gnd.n4083 gnd.n2208 19.3944
R15709 gnd.n4084 gnd.n4083 19.3944
R15710 gnd.n4085 gnd.n4084 19.3944
R15711 gnd.n4085 gnd.n2190 19.3944
R15712 gnd.n4103 gnd.n2190 19.3944
R15713 gnd.n4104 gnd.n4103 19.3944
R15714 gnd.n4106 gnd.n4104 19.3944
R15715 gnd.n4107 gnd.n4106 19.3944
R15716 gnd.n4107 gnd.n2164 19.3944
R15717 gnd.n4138 gnd.n2164 19.3944
R15718 gnd.n4139 gnd.n4138 19.3944
R15719 gnd.n4141 gnd.n4139 19.3944
R15720 gnd.n4142 gnd.n4141 19.3944
R15721 gnd.n4142 gnd.n2139 19.3944
R15722 gnd.n4173 gnd.n2139 19.3944
R15723 gnd.n4174 gnd.n4173 19.3944
R15724 gnd.n4176 gnd.n4174 19.3944
R15725 gnd.n4177 gnd.n4176 19.3944
R15726 gnd.n4177 gnd.n2113 19.3944
R15727 gnd.n4220 gnd.n2113 19.3944
R15728 gnd.n4221 gnd.n4220 19.3944
R15729 gnd.n4222 gnd.n4221 19.3944
R15730 gnd.n4222 gnd.n2096 19.3944
R15731 gnd.n4240 gnd.n2096 19.3944
R15732 gnd.n4241 gnd.n4240 19.3944
R15733 gnd.n4243 gnd.n4241 19.3944
R15734 gnd.n4244 gnd.n4243 19.3944
R15735 gnd.n4246 gnd.n4244 19.3944
R15736 gnd.n4246 gnd.n2073 19.3944
R15737 gnd.n4276 gnd.n2073 19.3944
R15738 gnd.n4277 gnd.n4276 19.3944
R15739 gnd.n4278 gnd.n4277 19.3944
R15740 gnd.n4279 gnd.n4278 19.3944
R15741 gnd.n4281 gnd.n4279 19.3944
R15742 gnd.n4281 gnd.n2061 19.3944
R15743 gnd.n4342 gnd.n2061 19.3944
R15744 gnd.n4343 gnd.n4342 19.3944
R15745 gnd.n4345 gnd.n4343 19.3944
R15746 gnd.n4345 gnd.n2056 19.3944
R15747 gnd.n4357 gnd.n2056 19.3944
R15748 gnd.n4358 gnd.n4357 19.3944
R15749 gnd.n4360 gnd.n4358 19.3944
R15750 gnd.n4360 gnd.n2051 19.3944
R15751 gnd.n4374 gnd.n2051 19.3944
R15752 gnd.n4375 gnd.n4374 19.3944
R15753 gnd.n4376 gnd.n4375 19.3944
R15754 gnd.n3919 gnd.n3917 19.3944
R15755 gnd.n3917 gnd.n3914 19.3944
R15756 gnd.n3914 gnd.n3913 19.3944
R15757 gnd.n3913 gnd.n3910 19.3944
R15758 gnd.n3910 gnd.n3909 19.3944
R15759 gnd.n3909 gnd.n3906 19.3944
R15760 gnd.n3906 gnd.n3905 19.3944
R15761 gnd.n3905 gnd.n3902 19.3944
R15762 gnd.n3902 gnd.n3901 19.3944
R15763 gnd.n3901 gnd.n3898 19.3944
R15764 gnd.n3898 gnd.n3897 19.3944
R15765 gnd.n3897 gnd.n3894 19.3944
R15766 gnd.n3894 gnd.n3893 19.3944
R15767 gnd.n3893 gnd.n3890 19.3944
R15768 gnd.n3890 gnd.n3889 19.3944
R15769 gnd.n3889 gnd.n3886 19.3944
R15770 gnd.n3880 gnd.n3878 19.3944
R15771 gnd.n3878 gnd.n3877 19.3944
R15772 gnd.n3877 gnd.n3875 19.3944
R15773 gnd.n3875 gnd.n3874 19.3944
R15774 gnd.n3874 gnd.n3872 19.3944
R15775 gnd.n3872 gnd.n3871 19.3944
R15776 gnd.n3871 gnd.n3869 19.3944
R15777 gnd.n3869 gnd.n3868 19.3944
R15778 gnd.n3868 gnd.n3866 19.3944
R15779 gnd.n3866 gnd.n3865 19.3944
R15780 gnd.n3865 gnd.n3863 19.3944
R15781 gnd.n3863 gnd.n3862 19.3944
R15782 gnd.n3862 gnd.n3860 19.3944
R15783 gnd.n3860 gnd.n2171 19.3944
R15784 gnd.n4128 gnd.n2171 19.3944
R15785 gnd.n4128 gnd.n2169 19.3944
R15786 gnd.n4134 gnd.n2169 19.3944
R15787 gnd.n4134 gnd.n4133 19.3944
R15788 gnd.n4133 gnd.n2146 19.3944
R15789 gnd.n4163 gnd.n2146 19.3944
R15790 gnd.n4163 gnd.n2144 19.3944
R15791 gnd.n4169 gnd.n2144 19.3944
R15792 gnd.n4169 gnd.n4168 19.3944
R15793 gnd.n4168 gnd.n2121 19.3944
R15794 gnd.n4198 gnd.n2121 19.3944
R15795 gnd.n4198 gnd.n2118 19.3944
R15796 gnd.n4216 gnd.n2118 19.3944
R15797 gnd.n4216 gnd.n2119 19.3944
R15798 gnd.n4212 gnd.n2119 19.3944
R15799 gnd.n4212 gnd.n4211 19.3944
R15800 gnd.n4211 gnd.n4210 19.3944
R15801 gnd.n4210 gnd.n4205 19.3944
R15802 gnd.n4206 gnd.n4205 19.3944
R15803 gnd.n4206 gnd.n2077 19.3944
R15804 gnd.n4268 gnd.n2077 19.3944
R15805 gnd.n4268 gnd.n2075 19.3944
R15806 gnd.n4272 gnd.n2075 19.3944
R15807 gnd.n4272 gnd.n2069 19.3944
R15808 gnd.n4292 gnd.n2069 19.3944
R15809 gnd.n4292 gnd.n2070 19.3944
R15810 gnd.n4288 gnd.n2070 19.3944
R15811 gnd.n4288 gnd.n4287 19.3944
R15812 gnd.n4287 gnd.n4286 19.3944
R15813 gnd.n4286 gnd.n2060 19.3944
R15814 gnd.n4349 gnd.n2060 19.3944
R15815 gnd.n4349 gnd.n2058 19.3944
R15816 gnd.n4353 gnd.n2058 19.3944
R15817 gnd.n4353 gnd.n2055 19.3944
R15818 gnd.n4364 gnd.n2055 19.3944
R15819 gnd.n4364 gnd.n2052 19.3944
R15820 gnd.n4370 gnd.n2052 19.3944
R15821 gnd.n4370 gnd.n2053 19.3944
R15822 gnd.n2053 gnd.n1851 19.3944
R15823 gnd.n4036 gnd.n4035 19.3944
R15824 gnd.n4035 gnd.n4034 19.3944
R15825 gnd.n4034 gnd.n4033 19.3944
R15826 gnd.n4033 gnd.n4031 19.3944
R15827 gnd.n4031 gnd.n4028 19.3944
R15828 gnd.n4028 gnd.n4027 19.3944
R15829 gnd.n4027 gnd.n4024 19.3944
R15830 gnd.n4024 gnd.n4023 19.3944
R15831 gnd.n4023 gnd.n4020 19.3944
R15832 gnd.n4020 gnd.n4019 19.3944
R15833 gnd.n4019 gnd.n4016 19.3944
R15834 gnd.n4016 gnd.n4015 19.3944
R15835 gnd.n4015 gnd.n4012 19.3944
R15836 gnd.n4012 gnd.n4011 19.3944
R15837 gnd.n4011 gnd.n4008 19.3944
R15838 gnd.n4008 gnd.n4007 19.3944
R15839 gnd.n4007 gnd.n4004 19.3944
R15840 gnd.n4002 gnd.n3999 19.3944
R15841 gnd.n3999 gnd.n3998 19.3944
R15842 gnd.n3998 gnd.n3995 19.3944
R15843 gnd.n3995 gnd.n3994 19.3944
R15844 gnd.n3994 gnd.n3991 19.3944
R15845 gnd.n3991 gnd.n3990 19.3944
R15846 gnd.n3990 gnd.n3987 19.3944
R15847 gnd.n3987 gnd.n3986 19.3944
R15848 gnd.n3986 gnd.n3983 19.3944
R15849 gnd.n3983 gnd.n3982 19.3944
R15850 gnd.n3982 gnd.n3979 19.3944
R15851 gnd.n3979 gnd.n3978 19.3944
R15852 gnd.n3978 gnd.n3975 19.3944
R15853 gnd.n3975 gnd.n3974 19.3944
R15854 gnd.n3974 gnd.n3971 19.3944
R15855 gnd.n3971 gnd.n3970 19.3944
R15856 gnd.n3970 gnd.n3967 19.3944
R15857 gnd.n3967 gnd.n3966 19.3944
R15858 gnd.n3962 gnd.n3959 19.3944
R15859 gnd.n3959 gnd.n3958 19.3944
R15860 gnd.n3958 gnd.n3955 19.3944
R15861 gnd.n3955 gnd.n3954 19.3944
R15862 gnd.n3954 gnd.n3951 19.3944
R15863 gnd.n3951 gnd.n3950 19.3944
R15864 gnd.n3950 gnd.n3947 19.3944
R15865 gnd.n3947 gnd.n3946 19.3944
R15866 gnd.n3946 gnd.n3943 19.3944
R15867 gnd.n3943 gnd.n3942 19.3944
R15868 gnd.n3942 gnd.n3939 19.3944
R15869 gnd.n3939 gnd.n3938 19.3944
R15870 gnd.n3938 gnd.n3935 19.3944
R15871 gnd.n3935 gnd.n3934 19.3944
R15872 gnd.n3934 gnd.n3931 19.3944
R15873 gnd.n3931 gnd.n3930 19.3944
R15874 gnd.n3930 gnd.n3927 19.3944
R15875 gnd.n3927 gnd.n3926 19.3944
R15876 gnd.n4054 gnd.n2235 19.3944
R15877 gnd.n4054 gnd.n2233 19.3944
R15878 gnd.n4058 gnd.n2233 19.3944
R15879 gnd.n4058 gnd.n2216 19.3944
R15880 gnd.n4074 gnd.n2216 19.3944
R15881 gnd.n4074 gnd.n2214 19.3944
R15882 gnd.n4078 gnd.n2214 19.3944
R15883 gnd.n4078 gnd.n2199 19.3944
R15884 gnd.n4094 gnd.n2199 19.3944
R15885 gnd.n4094 gnd.n2197 19.3944
R15886 gnd.n4098 gnd.n2197 19.3944
R15887 gnd.n4098 gnd.n2179 19.3944
R15888 gnd.n4118 gnd.n2179 19.3944
R15889 gnd.n4118 gnd.n2177 19.3944
R15890 gnd.n4124 gnd.n2177 19.3944
R15891 gnd.n4124 gnd.n4123 19.3944
R15892 gnd.n4123 gnd.n2154 19.3944
R15893 gnd.n4153 gnd.n2154 19.3944
R15894 gnd.n4153 gnd.n2152 19.3944
R15895 gnd.n4159 gnd.n2152 19.3944
R15896 gnd.n4159 gnd.n4158 19.3944
R15897 gnd.n4158 gnd.n2130 19.3944
R15898 gnd.n4188 gnd.n2130 19.3944
R15899 gnd.n4188 gnd.n2128 19.3944
R15900 gnd.n4194 gnd.n2128 19.3944
R15901 gnd.n4194 gnd.n4193 19.3944
R15902 gnd.n4193 gnd.n2105 19.3944
R15903 gnd.n4231 gnd.n2105 19.3944
R15904 gnd.n4231 gnd.n2103 19.3944
R15905 gnd.n4235 gnd.n2103 19.3944
R15906 gnd.n4235 gnd.n2084 19.3944
R15907 gnd.n4258 gnd.n2084 19.3944
R15908 gnd.n4258 gnd.n2082 19.3944
R15909 gnd.n4263 gnd.n2082 19.3944
R15910 gnd.n4263 gnd.n890 19.3944
R15911 gnd.n6005 gnd.n890 19.3944
R15912 gnd.n6005 gnd.n6004 19.3944
R15913 gnd.n6004 gnd.n6003 19.3944
R15914 gnd.n6003 gnd.n894 19.3944
R15915 gnd.n5993 gnd.n894 19.3944
R15916 gnd.n5993 gnd.n5992 19.3944
R15917 gnd.n5992 gnd.n5991 19.3944
R15918 gnd.n5991 gnd.n916 19.3944
R15919 gnd.n5981 gnd.n916 19.3944
R15920 gnd.n5981 gnd.n5980 19.3944
R15921 gnd.n5980 gnd.n5979 19.3944
R15922 gnd.n5979 gnd.n936 19.3944
R15923 gnd.n5969 gnd.n936 19.3944
R15924 gnd.n5969 gnd.n5968 19.3944
R15925 gnd.n5968 gnd.n5967 19.3944
R15926 gnd.n5967 gnd.n956 19.3944
R15927 gnd.n5957 gnd.n956 19.3944
R15928 gnd.n5957 gnd.n5956 19.3944
R15929 gnd.n5953 gnd.n976 19.3944
R15930 gnd.n5948 gnd.n976 19.3944
R15931 gnd.n5948 gnd.n5947 19.3944
R15932 gnd.n5947 gnd.n5946 19.3944
R15933 gnd.n5946 gnd.n5943 19.3944
R15934 gnd.n5943 gnd.n5942 19.3944
R15935 gnd.n5942 gnd.n5939 19.3944
R15936 gnd.n5939 gnd.n5938 19.3944
R15937 gnd.n5938 gnd.n5935 19.3944
R15938 gnd.n5935 gnd.n5934 19.3944
R15939 gnd.n5934 gnd.n5931 19.3944
R15940 gnd.n5931 gnd.n5930 19.3944
R15941 gnd.n5930 gnd.n5927 19.3944
R15942 gnd.n5927 gnd.n5926 19.3944
R15943 gnd.n5926 gnd.n5923 19.3944
R15944 gnd.n5923 gnd.n5922 19.3944
R15945 gnd.n5922 gnd.n5919 19.3944
R15946 gnd.n2001 gnd.n1967 19.3944
R15947 gnd.n2005 gnd.n1967 19.3944
R15948 gnd.n2008 gnd.n2005 19.3944
R15949 gnd.n2011 gnd.n2008 19.3944
R15950 gnd.n2011 gnd.n1965 19.3944
R15951 gnd.n2015 gnd.n1965 19.3944
R15952 gnd.n2018 gnd.n2015 19.3944
R15953 gnd.n2021 gnd.n2018 19.3944
R15954 gnd.n2021 gnd.n1963 19.3944
R15955 gnd.n2025 gnd.n1963 19.3944
R15956 gnd.n2028 gnd.n2025 19.3944
R15957 gnd.n2031 gnd.n2028 19.3944
R15958 gnd.n2031 gnd.n1961 19.3944
R15959 gnd.n2035 gnd.n1961 19.3944
R15960 gnd.n2038 gnd.n2035 19.3944
R15961 gnd.n2041 gnd.n2038 19.3944
R15962 gnd.n2041 gnd.n1959 19.3944
R15963 gnd.n2046 gnd.n1959 19.3944
R15964 gnd.n1979 gnd.n1045 19.3944
R15965 gnd.n1982 gnd.n1979 19.3944
R15966 gnd.n1982 gnd.n1974 19.3944
R15967 gnd.n1986 gnd.n1974 19.3944
R15968 gnd.n1989 gnd.n1986 19.3944
R15969 gnd.n1992 gnd.n1989 19.3944
R15970 gnd.n1992 gnd.n1972 19.3944
R15971 gnd.n1997 gnd.n1972 19.3944
R15972 gnd.n5917 gnd.n5914 19.3944
R15973 gnd.n5914 gnd.n5913 19.3944
R15974 gnd.n5913 gnd.n5910 19.3944
R15975 gnd.n5910 gnd.n5909 19.3944
R15976 gnd.n5909 gnd.n5906 19.3944
R15977 gnd.n5906 gnd.n5905 19.3944
R15978 gnd.n5905 gnd.n5902 19.3944
R15979 gnd.n4050 gnd.n2242 19.3944
R15980 gnd.n4050 gnd.n4049 19.3944
R15981 gnd.n4049 gnd.n4048 19.3944
R15982 gnd.n4048 gnd.n2224 19.3944
R15983 gnd.n4070 gnd.n2224 19.3944
R15984 gnd.n4070 gnd.n4069 19.3944
R15985 gnd.n4069 gnd.n4068 19.3944
R15986 gnd.n4068 gnd.n2206 19.3944
R15987 gnd.n4090 gnd.n2206 19.3944
R15988 gnd.n4090 gnd.n4089 19.3944
R15989 gnd.n4089 gnd.n4088 19.3944
R15990 gnd.n4088 gnd.n2187 19.3944
R15991 gnd.n4114 gnd.n2187 19.3944
R15992 gnd.n4114 gnd.n4113 19.3944
R15993 gnd.n4113 gnd.n4112 19.3944
R15994 gnd.n4112 gnd.n4111 19.3944
R15995 gnd.n4111 gnd.n2161 19.3944
R15996 gnd.n4149 gnd.n2161 19.3944
R15997 gnd.n4149 gnd.n4148 19.3944
R15998 gnd.n4148 gnd.n4147 19.3944
R15999 gnd.n4147 gnd.n4146 19.3944
R16000 gnd.n4146 gnd.n2136 19.3944
R16001 gnd.n4184 gnd.n2136 19.3944
R16002 gnd.n4184 gnd.n4183 19.3944
R16003 gnd.n4183 gnd.n4182 19.3944
R16004 gnd.n4182 gnd.n4181 19.3944
R16005 gnd.n4181 gnd.n2111 19.3944
R16006 gnd.n4227 gnd.n2111 19.3944
R16007 gnd.n4227 gnd.n4226 19.3944
R16008 gnd.n4226 gnd.n4225 19.3944
R16009 gnd.n4225 gnd.n2092 19.3944
R16010 gnd.n4254 gnd.n2092 19.3944
R16011 gnd.n4254 gnd.n4253 19.3944
R16012 gnd.n4253 gnd.n4252 19.3944
R16013 gnd.n4252 gnd.n4251 19.3944
R16014 gnd.n4251 gnd.n4249 19.3944
R16015 gnd.n4249 gnd.n901 19.3944
R16016 gnd.n5999 gnd.n901 19.3944
R16017 gnd.n5999 gnd.n5998 19.3944
R16018 gnd.n5998 gnd.n5997 19.3944
R16019 gnd.n5997 gnd.n905 19.3944
R16020 gnd.n5987 gnd.n905 19.3944
R16021 gnd.n5987 gnd.n5986 19.3944
R16022 gnd.n5986 gnd.n5985 19.3944
R16023 gnd.n5985 gnd.n926 19.3944
R16024 gnd.n5975 gnd.n926 19.3944
R16025 gnd.n5975 gnd.n5974 19.3944
R16026 gnd.n5974 gnd.n5973 19.3944
R16027 gnd.n5973 gnd.n945 19.3944
R16028 gnd.n5963 gnd.n945 19.3944
R16029 gnd.n5963 gnd.n5962 19.3944
R16030 gnd.n5962 gnd.n5961 19.3944
R16031 gnd.n5961 gnd.n966 19.3944
R16032 gnd.n4301 gnd.n4299 19.3944
R16033 gnd.n4301 gnd.n4297 19.3944
R16034 gnd.n4305 gnd.n4297 19.3944
R16035 gnd.n4305 gnd.n2067 19.3944
R16036 gnd.n4309 gnd.n2067 19.3944
R16037 gnd.n4309 gnd.n2065 19.3944
R16038 gnd.n4337 gnd.n2065 19.3944
R16039 gnd.n4337 gnd.n4336 19.3944
R16040 gnd.n4336 gnd.n4335 19.3944
R16041 gnd.n4335 gnd.n4315 19.3944
R16042 gnd.n4331 gnd.n4315 19.3944
R16043 gnd.n4331 gnd.n4330 19.3944
R16044 gnd.n4330 gnd.n4329 19.3944
R16045 gnd.n4329 gnd.n4321 19.3944
R16046 gnd.n4325 gnd.n4321 19.3944
R16047 gnd.n4325 gnd.n1855 19.3944
R16048 gnd.n4465 gnd.n1855 19.3944
R16049 gnd.n4465 gnd.n4464 19.3944
R16050 gnd.n4464 gnd.n4463 19.3944
R16051 gnd.n4463 gnd.n1859 19.3944
R16052 gnd.n1862 gnd.n1859 19.3944
R16053 gnd.n1862 gnd.n1838 19.3944
R16054 gnd.n4482 gnd.n1838 19.3944
R16055 gnd.n4482 gnd.n1836 19.3944
R16056 gnd.n4486 gnd.n1836 19.3944
R16057 gnd.n4486 gnd.n1825 19.3944
R16058 gnd.n4498 gnd.n1825 19.3944
R16059 gnd.n4498 gnd.n1823 19.3944
R16060 gnd.n4502 gnd.n1823 19.3944
R16061 gnd.n4502 gnd.n1809 19.3944
R16062 gnd.n4532 gnd.n1809 19.3944
R16063 gnd.n4532 gnd.n1807 19.3944
R16064 gnd.n4545 gnd.n1807 19.3944
R16065 gnd.n4545 gnd.n4544 19.3944
R16066 gnd.n4544 gnd.n4543 19.3944
R16067 gnd.n4543 gnd.n4540 19.3944
R16068 gnd.n4540 gnd.n1118 19.3944
R16069 gnd.n5823 gnd.n1118 19.3944
R16070 gnd.n5823 gnd.n5822 19.3944
R16071 gnd.n5822 gnd.n5821 19.3944
R16072 gnd.n5821 gnd.n1122 19.3944
R16073 gnd.n4652 gnd.n1122 19.3944
R16074 gnd.n4652 gnd.n1711 19.3944
R16075 gnd.n4661 gnd.n1711 19.3944
R16076 gnd.n4661 gnd.n4660 19.3944
R16077 gnd.n4660 gnd.n4659 19.3944
R16078 gnd.n4659 gnd.n1688 19.3944
R16079 gnd.n4692 gnd.n1688 19.3944
R16080 gnd.n4692 gnd.n1686 19.3944
R16081 gnd.n4698 gnd.n1686 19.3944
R16082 gnd.n4698 gnd.n4697 19.3944
R16083 gnd.n4697 gnd.n1660 19.3944
R16084 gnd.n4728 gnd.n1660 19.3944
R16085 gnd.n4728 gnd.n1658 19.3944
R16086 gnd.n4732 gnd.n1658 19.3944
R16087 gnd.n4732 gnd.n1642 19.3944
R16088 gnd.n4754 gnd.n1642 19.3944
R16089 gnd.n4754 gnd.n1640 19.3944
R16090 gnd.n4760 gnd.n1640 19.3944
R16091 gnd.n4760 gnd.n4759 19.3944
R16092 gnd.n4759 gnd.n1616 19.3944
R16093 gnd.n4810 gnd.n1616 19.3944
R16094 gnd.n4810 gnd.n1614 19.3944
R16095 gnd.n4816 gnd.n1614 19.3944
R16096 gnd.n4816 gnd.n4815 19.3944
R16097 gnd.n4815 gnd.n1591 19.3944
R16098 gnd.n4850 gnd.n1591 19.3944
R16099 gnd.n4850 gnd.n1589 19.3944
R16100 gnd.n4856 gnd.n1589 19.3944
R16101 gnd.n4856 gnd.n4855 19.3944
R16102 gnd.n4855 gnd.n1561 19.3944
R16103 gnd.n4919 gnd.n1561 19.3944
R16104 gnd.n4919 gnd.n1559 19.3944
R16105 gnd.n4925 gnd.n1559 19.3944
R16106 gnd.n4925 gnd.n4924 19.3944
R16107 gnd.n4924 gnd.n1537 19.3944
R16108 gnd.n4952 gnd.n1537 19.3944
R16109 gnd.n4952 gnd.n1535 19.3944
R16110 gnd.n4958 gnd.n1535 19.3944
R16111 gnd.n4958 gnd.n4957 19.3944
R16112 gnd.n4957 gnd.n1516 19.3944
R16113 gnd.n5006 gnd.n1516 19.3944
R16114 gnd.n5006 gnd.n1514 19.3944
R16115 gnd.n5012 gnd.n1514 19.3944
R16116 gnd.n5012 gnd.n5011 19.3944
R16117 gnd.n5011 gnd.n1491 19.3944
R16118 gnd.n5043 gnd.n1491 19.3944
R16119 gnd.n5043 gnd.n1489 19.3944
R16120 gnd.n5047 gnd.n1489 19.3944
R16121 gnd.n5047 gnd.n1400 19.3944
R16122 gnd.n5186 gnd.n1400 19.3944
R16123 gnd.n5186 gnd.n1398 19.3944
R16124 gnd.n5190 gnd.n1398 19.3944
R16125 gnd.n5190 gnd.n1387 19.3944
R16126 gnd.n5202 gnd.n1387 19.3944
R16127 gnd.n5202 gnd.n1385 19.3944
R16128 gnd.n5206 gnd.n1385 19.3944
R16129 gnd.n5206 gnd.n1374 19.3944
R16130 gnd.n5218 gnd.n1374 19.3944
R16131 gnd.n5218 gnd.n1372 19.3944
R16132 gnd.n5222 gnd.n1372 19.3944
R16133 gnd.n5222 gnd.n1361 19.3944
R16134 gnd.n5234 gnd.n1361 19.3944
R16135 gnd.n5234 gnd.n1359 19.3944
R16136 gnd.n5239 gnd.n1359 19.3944
R16137 gnd.n5239 gnd.n1234 19.3944
R16138 gnd.n5713 gnd.n1234 19.3944
R16139 gnd.n5713 gnd.n5712 19.3944
R16140 gnd.n5712 gnd.n5711 19.3944
R16141 gnd.n5711 gnd.n1238 19.3944
R16142 gnd.n5277 gnd.n1238 19.3944
R16143 gnd.n5472 gnd.n5277 19.3944
R16144 gnd.n5472 gnd.n5471 19.3944
R16145 gnd.n5471 gnd.n5470 19.3944
R16146 gnd.n5470 gnd.n5283 19.3944
R16147 gnd.n5391 gnd.n5283 19.3944
R16148 gnd.n5391 gnd.n5388 19.3944
R16149 gnd.n5397 gnd.n5388 19.3944
R16150 gnd.n5397 gnd.n5396 19.3944
R16151 gnd.n5396 gnd.n5341 19.3944
R16152 gnd.n5429 gnd.n5341 19.3944
R16153 gnd.n5429 gnd.n5339 19.3944
R16154 gnd.n5436 gnd.n5339 19.3944
R16155 gnd.n5436 gnd.n5435 19.3944
R16156 gnd.n5435 gnd.n391 19.3944
R16157 gnd.n6719 gnd.n391 19.3944
R16158 gnd.n6719 gnd.n6718 19.3944
R16159 gnd.n6718 gnd.n6717 19.3944
R16160 gnd.n6503 gnd.n518 19.3944
R16161 gnd.n6509 gnd.n518 19.3944
R16162 gnd.n6509 gnd.n516 19.3944
R16163 gnd.n6513 gnd.n516 19.3944
R16164 gnd.n6513 gnd.n512 19.3944
R16165 gnd.n6519 gnd.n512 19.3944
R16166 gnd.n6519 gnd.n510 19.3944
R16167 gnd.n6523 gnd.n510 19.3944
R16168 gnd.n6523 gnd.n506 19.3944
R16169 gnd.n6529 gnd.n506 19.3944
R16170 gnd.n6529 gnd.n504 19.3944
R16171 gnd.n6533 gnd.n504 19.3944
R16172 gnd.n6533 gnd.n500 19.3944
R16173 gnd.n6539 gnd.n500 19.3944
R16174 gnd.n6539 gnd.n498 19.3944
R16175 gnd.n6543 gnd.n498 19.3944
R16176 gnd.n6543 gnd.n494 19.3944
R16177 gnd.n6549 gnd.n494 19.3944
R16178 gnd.n6549 gnd.n492 19.3944
R16179 gnd.n6553 gnd.n492 19.3944
R16180 gnd.n6553 gnd.n488 19.3944
R16181 gnd.n6559 gnd.n488 19.3944
R16182 gnd.n6559 gnd.n486 19.3944
R16183 gnd.n6563 gnd.n486 19.3944
R16184 gnd.n6563 gnd.n482 19.3944
R16185 gnd.n6569 gnd.n482 19.3944
R16186 gnd.n6569 gnd.n480 19.3944
R16187 gnd.n6573 gnd.n480 19.3944
R16188 gnd.n6573 gnd.n476 19.3944
R16189 gnd.n6579 gnd.n476 19.3944
R16190 gnd.n6579 gnd.n474 19.3944
R16191 gnd.n6583 gnd.n474 19.3944
R16192 gnd.n6583 gnd.n470 19.3944
R16193 gnd.n6589 gnd.n470 19.3944
R16194 gnd.n6589 gnd.n468 19.3944
R16195 gnd.n6593 gnd.n468 19.3944
R16196 gnd.n6593 gnd.n464 19.3944
R16197 gnd.n6599 gnd.n464 19.3944
R16198 gnd.n6599 gnd.n462 19.3944
R16199 gnd.n6603 gnd.n462 19.3944
R16200 gnd.n6603 gnd.n458 19.3944
R16201 gnd.n6609 gnd.n458 19.3944
R16202 gnd.n6609 gnd.n456 19.3944
R16203 gnd.n6613 gnd.n456 19.3944
R16204 gnd.n6613 gnd.n452 19.3944
R16205 gnd.n6619 gnd.n452 19.3944
R16206 gnd.n6619 gnd.n450 19.3944
R16207 gnd.n6623 gnd.n450 19.3944
R16208 gnd.n6623 gnd.n446 19.3944
R16209 gnd.n6629 gnd.n446 19.3944
R16210 gnd.n6629 gnd.n444 19.3944
R16211 gnd.n6633 gnd.n444 19.3944
R16212 gnd.n6633 gnd.n440 19.3944
R16213 gnd.n6639 gnd.n440 19.3944
R16214 gnd.n6639 gnd.n438 19.3944
R16215 gnd.n6643 gnd.n438 19.3944
R16216 gnd.n6643 gnd.n434 19.3944
R16217 gnd.n6649 gnd.n434 19.3944
R16218 gnd.n6649 gnd.n432 19.3944
R16219 gnd.n6653 gnd.n432 19.3944
R16220 gnd.n6653 gnd.n428 19.3944
R16221 gnd.n6659 gnd.n428 19.3944
R16222 gnd.n6659 gnd.n426 19.3944
R16223 gnd.n6663 gnd.n426 19.3944
R16224 gnd.n6663 gnd.n422 19.3944
R16225 gnd.n6669 gnd.n422 19.3944
R16226 gnd.n6669 gnd.n420 19.3944
R16227 gnd.n6673 gnd.n420 19.3944
R16228 gnd.n6673 gnd.n416 19.3944
R16229 gnd.n6679 gnd.n416 19.3944
R16230 gnd.n6679 gnd.n414 19.3944
R16231 gnd.n6683 gnd.n414 19.3944
R16232 gnd.n6683 gnd.n410 19.3944
R16233 gnd.n6689 gnd.n410 19.3944
R16234 gnd.n6689 gnd.n408 19.3944
R16235 gnd.n6693 gnd.n408 19.3944
R16236 gnd.n6693 gnd.n404 19.3944
R16237 gnd.n6699 gnd.n404 19.3944
R16238 gnd.n6699 gnd.n402 19.3944
R16239 gnd.n6703 gnd.n402 19.3944
R16240 gnd.n6703 gnd.n398 19.3944
R16241 gnd.n6710 gnd.n398 19.3944
R16242 gnd.n6710 gnd.n396 19.3944
R16243 gnd.n6714 gnd.n396 19.3944
R16244 gnd.n6182 gnd.n713 19.3944
R16245 gnd.n6182 gnd.n709 19.3944
R16246 gnd.n6188 gnd.n709 19.3944
R16247 gnd.n6188 gnd.n707 19.3944
R16248 gnd.n6192 gnd.n707 19.3944
R16249 gnd.n6192 gnd.n703 19.3944
R16250 gnd.n6198 gnd.n703 19.3944
R16251 gnd.n6198 gnd.n701 19.3944
R16252 gnd.n6202 gnd.n701 19.3944
R16253 gnd.n6202 gnd.n697 19.3944
R16254 gnd.n6208 gnd.n697 19.3944
R16255 gnd.n6208 gnd.n695 19.3944
R16256 gnd.n6212 gnd.n695 19.3944
R16257 gnd.n6212 gnd.n691 19.3944
R16258 gnd.n6218 gnd.n691 19.3944
R16259 gnd.n6218 gnd.n689 19.3944
R16260 gnd.n6222 gnd.n689 19.3944
R16261 gnd.n6222 gnd.n685 19.3944
R16262 gnd.n6228 gnd.n685 19.3944
R16263 gnd.n6228 gnd.n683 19.3944
R16264 gnd.n6232 gnd.n683 19.3944
R16265 gnd.n6232 gnd.n679 19.3944
R16266 gnd.n6238 gnd.n679 19.3944
R16267 gnd.n6238 gnd.n677 19.3944
R16268 gnd.n6242 gnd.n677 19.3944
R16269 gnd.n6242 gnd.n673 19.3944
R16270 gnd.n6248 gnd.n673 19.3944
R16271 gnd.n6248 gnd.n671 19.3944
R16272 gnd.n6252 gnd.n671 19.3944
R16273 gnd.n6252 gnd.n667 19.3944
R16274 gnd.n6258 gnd.n667 19.3944
R16275 gnd.n6258 gnd.n665 19.3944
R16276 gnd.n6262 gnd.n665 19.3944
R16277 gnd.n6262 gnd.n661 19.3944
R16278 gnd.n6268 gnd.n661 19.3944
R16279 gnd.n6268 gnd.n659 19.3944
R16280 gnd.n6272 gnd.n659 19.3944
R16281 gnd.n6272 gnd.n655 19.3944
R16282 gnd.n6278 gnd.n655 19.3944
R16283 gnd.n6278 gnd.n653 19.3944
R16284 gnd.n6282 gnd.n653 19.3944
R16285 gnd.n6282 gnd.n649 19.3944
R16286 gnd.n6288 gnd.n649 19.3944
R16287 gnd.n6288 gnd.n647 19.3944
R16288 gnd.n6292 gnd.n647 19.3944
R16289 gnd.n6292 gnd.n643 19.3944
R16290 gnd.n6298 gnd.n643 19.3944
R16291 gnd.n6298 gnd.n641 19.3944
R16292 gnd.n6302 gnd.n641 19.3944
R16293 gnd.n6302 gnd.n637 19.3944
R16294 gnd.n6308 gnd.n637 19.3944
R16295 gnd.n6308 gnd.n635 19.3944
R16296 gnd.n6312 gnd.n635 19.3944
R16297 gnd.n6312 gnd.n631 19.3944
R16298 gnd.n6318 gnd.n631 19.3944
R16299 gnd.n6318 gnd.n629 19.3944
R16300 gnd.n6322 gnd.n629 19.3944
R16301 gnd.n6322 gnd.n625 19.3944
R16302 gnd.n6328 gnd.n625 19.3944
R16303 gnd.n6328 gnd.n623 19.3944
R16304 gnd.n6332 gnd.n623 19.3944
R16305 gnd.n6332 gnd.n619 19.3944
R16306 gnd.n6338 gnd.n619 19.3944
R16307 gnd.n6338 gnd.n617 19.3944
R16308 gnd.n6342 gnd.n617 19.3944
R16309 gnd.n6342 gnd.n613 19.3944
R16310 gnd.n6348 gnd.n613 19.3944
R16311 gnd.n6348 gnd.n611 19.3944
R16312 gnd.n6352 gnd.n611 19.3944
R16313 gnd.n6352 gnd.n607 19.3944
R16314 gnd.n6358 gnd.n607 19.3944
R16315 gnd.n6358 gnd.n605 19.3944
R16316 gnd.n6362 gnd.n605 19.3944
R16317 gnd.n6362 gnd.n601 19.3944
R16318 gnd.n6368 gnd.n601 19.3944
R16319 gnd.n6368 gnd.n599 19.3944
R16320 gnd.n6372 gnd.n599 19.3944
R16321 gnd.n6372 gnd.n595 19.3944
R16322 gnd.n6378 gnd.n595 19.3944
R16323 gnd.n6378 gnd.n593 19.3944
R16324 gnd.n6382 gnd.n593 19.3944
R16325 gnd.n6382 gnd.n589 19.3944
R16326 gnd.n6388 gnd.n589 19.3944
R16327 gnd.n6388 gnd.n587 19.3944
R16328 gnd.n6392 gnd.n587 19.3944
R16329 gnd.n6392 gnd.n583 19.3944
R16330 gnd.n6398 gnd.n583 19.3944
R16331 gnd.n6398 gnd.n581 19.3944
R16332 gnd.n6402 gnd.n581 19.3944
R16333 gnd.n6402 gnd.n577 19.3944
R16334 gnd.n6408 gnd.n577 19.3944
R16335 gnd.n6408 gnd.n575 19.3944
R16336 gnd.n6412 gnd.n575 19.3944
R16337 gnd.n6412 gnd.n571 19.3944
R16338 gnd.n6418 gnd.n571 19.3944
R16339 gnd.n6418 gnd.n569 19.3944
R16340 gnd.n6422 gnd.n569 19.3944
R16341 gnd.n6422 gnd.n565 19.3944
R16342 gnd.n6428 gnd.n565 19.3944
R16343 gnd.n6428 gnd.n563 19.3944
R16344 gnd.n6432 gnd.n563 19.3944
R16345 gnd.n6432 gnd.n559 19.3944
R16346 gnd.n6438 gnd.n559 19.3944
R16347 gnd.n6438 gnd.n557 19.3944
R16348 gnd.n6442 gnd.n557 19.3944
R16349 gnd.n6442 gnd.n553 19.3944
R16350 gnd.n6448 gnd.n553 19.3944
R16351 gnd.n6448 gnd.n551 19.3944
R16352 gnd.n6452 gnd.n551 19.3944
R16353 gnd.n6452 gnd.n547 19.3944
R16354 gnd.n6458 gnd.n547 19.3944
R16355 gnd.n6458 gnd.n545 19.3944
R16356 gnd.n6462 gnd.n545 19.3944
R16357 gnd.n6462 gnd.n541 19.3944
R16358 gnd.n6468 gnd.n541 19.3944
R16359 gnd.n6468 gnd.n539 19.3944
R16360 gnd.n6472 gnd.n539 19.3944
R16361 gnd.n6472 gnd.n535 19.3944
R16362 gnd.n6478 gnd.n535 19.3944
R16363 gnd.n6478 gnd.n533 19.3944
R16364 gnd.n6482 gnd.n533 19.3944
R16365 gnd.n6482 gnd.n529 19.3944
R16366 gnd.n6488 gnd.n529 19.3944
R16367 gnd.n6488 gnd.n527 19.3944
R16368 gnd.n6493 gnd.n527 19.3944
R16369 gnd.n6493 gnd.n523 19.3944
R16370 gnd.n6499 gnd.n523 19.3944
R16371 gnd.n6500 gnd.n6499 19.3944
R16372 gnd.n6178 gnd.n715 19.3944
R16373 gnd.n6172 gnd.n715 19.3944
R16374 gnd.n6172 gnd.n6171 19.3944
R16375 gnd.n6171 gnd.n6170 19.3944
R16376 gnd.n6170 gnd.n722 19.3944
R16377 gnd.n6164 gnd.n722 19.3944
R16378 gnd.n6164 gnd.n6163 19.3944
R16379 gnd.n6163 gnd.n6162 19.3944
R16380 gnd.n6162 gnd.n730 19.3944
R16381 gnd.n6156 gnd.n730 19.3944
R16382 gnd.n6156 gnd.n6155 19.3944
R16383 gnd.n6155 gnd.n6154 19.3944
R16384 gnd.n6154 gnd.n738 19.3944
R16385 gnd.n6148 gnd.n738 19.3944
R16386 gnd.n6148 gnd.n6147 19.3944
R16387 gnd.n6147 gnd.n6146 19.3944
R16388 gnd.n6146 gnd.n746 19.3944
R16389 gnd.n6140 gnd.n746 19.3944
R16390 gnd.n6140 gnd.n6139 19.3944
R16391 gnd.n6139 gnd.n6138 19.3944
R16392 gnd.n6138 gnd.n754 19.3944
R16393 gnd.n6132 gnd.n754 19.3944
R16394 gnd.n6132 gnd.n6131 19.3944
R16395 gnd.n6131 gnd.n6130 19.3944
R16396 gnd.n6130 gnd.n762 19.3944
R16397 gnd.n6124 gnd.n762 19.3944
R16398 gnd.n6124 gnd.n6123 19.3944
R16399 gnd.n6123 gnd.n6122 19.3944
R16400 gnd.n6122 gnd.n770 19.3944
R16401 gnd.n6116 gnd.n770 19.3944
R16402 gnd.n6116 gnd.n6115 19.3944
R16403 gnd.n6115 gnd.n6114 19.3944
R16404 gnd.n6114 gnd.n778 19.3944
R16405 gnd.n6108 gnd.n778 19.3944
R16406 gnd.n6108 gnd.n6107 19.3944
R16407 gnd.n6107 gnd.n6106 19.3944
R16408 gnd.n6106 gnd.n786 19.3944
R16409 gnd.n6100 gnd.n786 19.3944
R16410 gnd.n6100 gnd.n6099 19.3944
R16411 gnd.n6099 gnd.n6098 19.3944
R16412 gnd.n6098 gnd.n794 19.3944
R16413 gnd.n6092 gnd.n794 19.3944
R16414 gnd.n6092 gnd.n6091 19.3944
R16415 gnd.n6091 gnd.n6090 19.3944
R16416 gnd.n6090 gnd.n802 19.3944
R16417 gnd.n6084 gnd.n802 19.3944
R16418 gnd.n6084 gnd.n6083 19.3944
R16419 gnd.n6083 gnd.n6082 19.3944
R16420 gnd.n6082 gnd.n810 19.3944
R16421 gnd.n6076 gnd.n810 19.3944
R16422 gnd.n6076 gnd.n6075 19.3944
R16423 gnd.n6075 gnd.n6074 19.3944
R16424 gnd.n6074 gnd.n818 19.3944
R16425 gnd.n6068 gnd.n818 19.3944
R16426 gnd.n6068 gnd.n6067 19.3944
R16427 gnd.n6067 gnd.n6066 19.3944
R16428 gnd.n6066 gnd.n826 19.3944
R16429 gnd.n6060 gnd.n826 19.3944
R16430 gnd.n6060 gnd.n6059 19.3944
R16431 gnd.n6059 gnd.n6058 19.3944
R16432 gnd.n6058 gnd.n834 19.3944
R16433 gnd.n6052 gnd.n834 19.3944
R16434 gnd.n6052 gnd.n6051 19.3944
R16435 gnd.n6051 gnd.n6050 19.3944
R16436 gnd.n6050 gnd.n842 19.3944
R16437 gnd.n6044 gnd.n842 19.3944
R16438 gnd.n6044 gnd.n6043 19.3944
R16439 gnd.n6043 gnd.n6042 19.3944
R16440 gnd.n6042 gnd.n850 19.3944
R16441 gnd.n6036 gnd.n850 19.3944
R16442 gnd.n6036 gnd.n6035 19.3944
R16443 gnd.n6035 gnd.n6034 19.3944
R16444 gnd.n6034 gnd.n858 19.3944
R16445 gnd.n6028 gnd.n858 19.3944
R16446 gnd.n6028 gnd.n6027 19.3944
R16447 gnd.n6027 gnd.n6026 19.3944
R16448 gnd.n6026 gnd.n866 19.3944
R16449 gnd.n6020 gnd.n866 19.3944
R16450 gnd.n6020 gnd.n6019 19.3944
R16451 gnd.n6019 gnd.n6018 19.3944
R16452 gnd.n6018 gnd.n874 19.3944
R16453 gnd.n6012 gnd.n874 19.3944
R16454 gnd.n6012 gnd.n6011 19.3944
R16455 gnd.n6011 gnd.n6010 19.3944
R16456 gnd.n1941 gnd.n1940 19.3944
R16457 gnd.n1940 gnd.n1939 19.3944
R16458 gnd.n1939 gnd.n1924 19.3944
R16459 gnd.n1935 gnd.n1924 19.3944
R16460 gnd.n1935 gnd.n1934 19.3944
R16461 gnd.n1934 gnd.n1933 19.3944
R16462 gnd.n1933 gnd.n1928 19.3944
R16463 gnd.n1929 gnd.n1928 19.3944
R16464 gnd.n1929 gnd.n1801 19.3944
R16465 gnd.n4549 gnd.n1801 19.3944
R16466 gnd.n4549 gnd.n1799 19.3944
R16467 gnd.n4553 gnd.n1799 19.3944
R16468 gnd.n4553 gnd.n1797 19.3944
R16469 gnd.n4557 gnd.n1797 19.3944
R16470 gnd.n4557 gnd.n1794 19.3944
R16471 gnd.n4619 gnd.n1794 19.3944
R16472 gnd.n4619 gnd.n1795 19.3944
R16473 gnd.n4615 gnd.n1795 19.3944
R16474 gnd.n4615 gnd.n4614 19.3944
R16475 gnd.n4614 gnd.n4613 19.3944
R16476 gnd.n4613 gnd.n4565 19.3944
R16477 gnd.n4609 gnd.n4565 19.3944
R16478 gnd.n4609 gnd.n4608 19.3944
R16479 gnd.n4608 gnd.n4607 19.3944
R16480 gnd.n4607 gnd.n4569 19.3944
R16481 gnd.n4603 gnd.n4569 19.3944
R16482 gnd.n4603 gnd.n4602 19.3944
R16483 gnd.n4602 gnd.n4601 19.3944
R16484 gnd.n4601 gnd.n4574 19.3944
R16485 gnd.n4597 gnd.n4574 19.3944
R16486 gnd.n4597 gnd.n4596 19.3944
R16487 gnd.n4596 gnd.n4595 19.3944
R16488 gnd.n4595 gnd.n4578 19.3944
R16489 gnd.n4591 gnd.n4578 19.3944
R16490 gnd.n4591 gnd.n4590 19.3944
R16491 gnd.n4590 gnd.n4589 19.3944
R16492 gnd.n4589 gnd.n4582 19.3944
R16493 gnd.n4585 gnd.n4582 19.3944
R16494 gnd.n4585 gnd.n4584 19.3944
R16495 gnd.n4584 gnd.n1606 19.3944
R16496 gnd.n4820 gnd.n1606 19.3944
R16497 gnd.n4820 gnd.n1603 19.3944
R16498 gnd.n4838 gnd.n1603 19.3944
R16499 gnd.n4838 gnd.n1604 19.3944
R16500 gnd.n4834 gnd.n1604 19.3944
R16501 gnd.n4834 gnd.n4833 19.3944
R16502 gnd.n4833 gnd.n4832 19.3944
R16503 gnd.n4832 gnd.n4827 19.3944
R16504 gnd.n4828 gnd.n4827 19.3944
R16505 gnd.n4828 gnd.n1553 19.3944
R16506 gnd.n4929 gnd.n1553 19.3944
R16507 gnd.n4929 gnd.n1550 19.3944
R16508 gnd.n4934 gnd.n1550 19.3944
R16509 gnd.n4934 gnd.n1551 19.3944
R16510 gnd.n1551 gnd.n1530 19.3944
R16511 gnd.n4962 gnd.n1530 19.3944
R16512 gnd.n4962 gnd.n1527 19.3944
R16513 gnd.n4993 gnd.n1527 19.3944
R16514 gnd.n4993 gnd.n1528 19.3944
R16515 gnd.n4989 gnd.n1528 19.3944
R16516 gnd.n4989 gnd.n4988 19.3944
R16517 gnd.n4988 gnd.n4987 19.3944
R16518 gnd.n4987 gnd.n4972 19.3944
R16519 gnd.n4983 gnd.n4972 19.3944
R16520 gnd.n4983 gnd.n4982 19.3944
R16521 gnd.n4982 gnd.n4981 19.3944
R16522 gnd.n4981 gnd.n4976 19.3944
R16523 gnd.n4977 gnd.n4976 19.3944
R16524 gnd.n4977 gnd.n1392 19.3944
R16525 gnd.n5194 gnd.n1392 19.3944
R16526 gnd.n5194 gnd.n1390 19.3944
R16527 gnd.n5198 gnd.n1390 19.3944
R16528 gnd.n5198 gnd.n1379 19.3944
R16529 gnd.n5210 gnd.n1379 19.3944
R16530 gnd.n5210 gnd.n1377 19.3944
R16531 gnd.n5214 gnd.n1377 19.3944
R16532 gnd.n5214 gnd.n1367 19.3944
R16533 gnd.n5226 gnd.n1367 19.3944
R16534 gnd.n5226 gnd.n1365 19.3944
R16535 gnd.n5230 gnd.n1365 19.3944
R16536 gnd.n5230 gnd.n1354 19.3944
R16537 gnd.n5243 gnd.n1354 19.3944
R16538 gnd.n5247 gnd.n1352 19.3944
R16539 gnd.n5250 gnd.n5247 19.3944
R16540 gnd.n5253 gnd.n5250 19.3944
R16541 gnd.n5253 gnd.n1350 19.3944
R16542 gnd.n5257 gnd.n1350 19.3944
R16543 gnd.n5260 gnd.n5257 19.3944
R16544 gnd.n5589 gnd.n5260 19.3944
R16545 gnd.n5589 gnd.n5588 19.3944
R16546 gnd.n5588 gnd.n5587 19.3944
R16547 gnd.n5587 gnd.n5265 19.3944
R16548 gnd.n5580 gnd.n5265 19.3944
R16549 gnd.n5580 gnd.n5579 19.3944
R16550 gnd.n5579 gnd.n5485 19.3944
R16551 gnd.n5572 gnd.n5485 19.3944
R16552 gnd.n5572 gnd.n5571 19.3944
R16553 gnd.n5571 gnd.n5497 19.3944
R16554 gnd.n5564 gnd.n5497 19.3944
R16555 gnd.n5564 gnd.n5563 19.3944
R16556 gnd.n5563 gnd.n5505 19.3944
R16557 gnd.n5556 gnd.n5505 19.3944
R16558 gnd.n5556 gnd.n5555 19.3944
R16559 gnd.n5555 gnd.n5517 19.3944
R16560 gnd.n5548 gnd.n5517 19.3944
R16561 gnd.n5548 gnd.n5547 19.3944
R16562 gnd.n5537 gnd.n5534 19.3944
R16563 gnd.n5537 gnd.n1213 19.3944
R16564 gnd.n5717 gnd.n1213 19.3944
R16565 gnd.n2247 gnd.n876 19.1949
R16566 gnd.n6969 gnd.n157 19.1199
R16567 gnd.n3112 gnd.t335 18.8012
R16568 gnd.n3097 gnd.t346 18.8012
R16569 gnd.n2956 gnd.n2955 18.4825
R16570 gnd.n4650 gnd.n4649 18.4825
R16571 gnd.n4742 gnd.t326 18.4825
R16572 gnd.t325 gnd.n1563 18.4825
R16573 gnd.n4967 gnd.n1500 18.4825
R16574 gnd.n5656 gnd.n5655 18.4247
R16575 gnd.n5902 gnd.n5901 18.4247
R16576 gnd.n5544 gnd.n5543 18.2308
R16577 gnd.n6946 gnd.n6897 18.2308
R16578 gnd.n4451 gnd.n1850 18.2308
R16579 gnd.n3886 gnd.n3846 18.2308
R16580 gnd.t336 gnd.n2636 18.1639
R16581 gnd.n2664 gnd.t333 17.5266
R16582 gnd.n2221 gnd.t73 17.5266
R16583 gnd.n182 gnd.t13 17.5266
R16584 gnd.n1787 gnd.n1110 17.2079
R16585 gnd.n5819 gnd.n1126 17.2079
R16586 gnd.n4724 gnd.n1665 17.2079
R16587 gnd.n4927 gnd.n1556 17.2079
R16588 gnd.n5040 gnd.n1496 17.2079
R16589 gnd.n3063 gnd.t344 16.8893
R16590 gnd.n2184 gnd.t24 16.8893
R16591 gnd.t68 gnd.n918 16.8893
R16592 gnd.n5438 gnd.t32 16.8893
R16593 gnd.n144 gnd.t38 16.8893
R16594 gnd.n7039 gnd.n7036 16.6793
R16595 gnd.n5638 gnd.n5635 16.6793
R16596 gnd.n3966 gnd.n3963 16.6793
R16597 gnd.n1998 gnd.n1997 16.6793
R16598 gnd.n4735 gnd.t322 16.5706
R16599 gnd.n4898 gnd.t189 16.5706
R16600 gnd.n2891 gnd.t208 16.2519
R16601 gnd.n2591 gnd.t343 16.2519
R16602 gnd.n4171 gnd.t59 16.2519
R16603 gnd.t108 gnd.n2086 16.2519
R16604 gnd.n1842 gnd.t263 16.2519
R16605 gnd.t247 gnd.n1357 16.2519
R16606 gnd.n6793 gnd.t83 16.2519
R16607 gnd.n106 gnd.t103 16.2519
R16608 gnd.n5825 gnd.n1114 15.9333
R16609 gnd.n4734 gnd.n1656 15.9333
R16610 gnd.n1656 gnd.n1649 15.9333
R16611 gnd.n4917 gnd.n4916 15.9333
R16612 gnd.n4916 gnd.n1567 15.9333
R16613 gnd.n3578 gnd.n3576 15.6674
R16614 gnd.n3546 gnd.n3544 15.6674
R16615 gnd.n3514 gnd.n3512 15.6674
R16616 gnd.n3483 gnd.n3481 15.6674
R16617 gnd.n3451 gnd.n3449 15.6674
R16618 gnd.n3419 gnd.n3417 15.6674
R16619 gnd.n3387 gnd.n3385 15.6674
R16620 gnd.n3356 gnd.n3354 15.6674
R16621 gnd.n2882 gnd.t208 15.6146
R16622 gnd.t204 gnd.n2329 15.6146
R16623 gnd.t301 gnd.n2330 15.6146
R16624 gnd.n4186 gnd.t59 15.6146
R16625 gnd.n4237 gnd.t108 15.6146
R16626 gnd.n4488 gnd.t263 15.6146
R16627 gnd.n4681 gnd.t177 15.6146
R16628 gnd.n4997 gnd.t197 15.6146
R16629 gnd.n5232 gnd.t247 15.6146
R16630 gnd.n6802 gnd.t83 15.6146
R16631 gnd.n7185 gnd.t103 15.6146
R16632 gnd.n6994 gnd.n305 15.3217
R16633 gnd.n5595 gnd.n1344 15.3217
R16634 gnd.n3924 gnd.n2245 15.3217
R16635 gnd.n2049 gnd.n2047 15.3217
R16636 gnd.n1413 gnd.n1412 15.0827
R16637 gnd.n1096 gnd.n1091 15.0481
R16638 gnd.n1423 gnd.n1422 15.0481
R16639 gnd.n3250 gnd.t338 14.9773
R16640 gnd.n4126 gnd.t24 14.9773
R16641 gnd.n6001 gnd.t26 14.9773
R16642 gnd.t175 gnd.n4750 14.9773
R16643 gnd.n1578 gnd.t179 14.9773
R16644 gnd.n6745 gnd.t54 14.9773
R16645 gnd.n7161 gnd.t38 14.9773
R16646 gnd.n4561 gnd.n1126 14.6587
R16647 gnd.n4663 gnd.t329 14.6587
R16648 gnd.n4726 gnd.n4724 14.6587
R16649 gnd.n4750 gnd.n1635 14.6587
R16650 gnd.n1579 gnd.n1578 14.6587
R16651 gnd.n4870 gnd.n1556 14.6587
R16652 gnd.t188 gnd.n5014 14.6587
R16653 gnd.n5041 gnd.n5040 14.6587
R16654 gnd.n5183 gnd.n1405 14.6587
R16655 gnd.t6 gnd.n2372 14.34
R16656 gnd.n3328 gnd.t332 14.34
R16657 gnd.n4080 gnd.t73 14.34
R16658 gnd.n5977 gnd.t36 14.34
R16659 gnd.n5455 gnd.t43 14.34
R16660 gnd.n7137 gnd.t13 14.34
R16661 gnd.n3038 gnd.t4 13.7027
R16662 gnd.n2748 gnd.n2747 13.5763
R16663 gnd.n3692 gnd.n2285 13.5763
R16664 gnd.n2956 gnd.n2694 13.384
R16665 gnd.n1676 gnd.n1675 13.384
R16666 gnd.n1675 gnd.t319 13.384
R16667 gnd.n4770 gnd.n1631 13.384
R16668 gnd.n4859 gnd.n1583 13.384
R16669 gnd.t173 gnd.n1539 13.384
R16670 gnd.n4950 gnd.n1539 13.384
R16671 gnd.n4969 gnd.n4967 13.384
R16672 gnd.n1107 gnd.n1088 13.1884
R16673 gnd.n1102 gnd.n1101 13.1884
R16674 gnd.n1101 gnd.n1100 13.1884
R16675 gnd.n1416 gnd.n1411 13.1884
R16676 gnd.n1417 gnd.n1416 13.1884
R16677 gnd.n1103 gnd.n1090 13.146
R16678 gnd.n1099 gnd.n1090 13.146
R16679 gnd.n1415 gnd.n1414 13.146
R16680 gnd.n1415 gnd.n1410 13.146
R16681 gnd.n4621 gnd.t190 13.0654
R16682 gnd.n5049 gnd.t354 13.0654
R16683 gnd.n3579 gnd.n3575 12.8005
R16684 gnd.n3547 gnd.n3543 12.8005
R16685 gnd.n3515 gnd.n3511 12.8005
R16686 gnd.n3484 gnd.n3480 12.8005
R16687 gnd.n3452 gnd.n3448 12.8005
R16688 gnd.n3420 gnd.n3416 12.8005
R16689 gnd.n3388 gnd.n3384 12.8005
R16690 gnd.n3357 gnd.n3353 12.8005
R16691 gnd.t230 gnd.t200 12.7467
R16692 gnd.n7149 gnd.n157 12.7467
R16693 gnd.n2747 gnd.n2742 12.4126
R16694 gnd.n3695 gnd.n3692 12.4126
R16695 gnd.n5894 gnd.n5831 12.1761
R16696 gnd.n5180 gnd.n5179 12.1761
R16697 gnd.n4633 gnd.n1702 12.1094
R16698 gnd.t327 gnd.n1681 12.1094
R16699 gnd.n4960 gnd.t8 12.1094
R16700 gnd.n5015 gnd.n1509 12.1094
R16701 gnd.t254 gnd.n1493 12.1094
R16702 gnd.n5184 gnd.t215 12.1094
R16703 gnd.n3583 gnd.n3582 12.0247
R16704 gnd.n3551 gnd.n3550 12.0247
R16705 gnd.n3519 gnd.n3518 12.0247
R16706 gnd.n3488 gnd.n3487 12.0247
R16707 gnd.n3456 gnd.n3455 12.0247
R16708 gnd.n3424 gnd.n3423 12.0247
R16709 gnd.n3392 gnd.n3391 12.0247
R16710 gnd.n3361 gnd.n3360 12.0247
R16711 gnd.t240 gnd.n968 11.7908
R16712 gnd.t218 gnd.n5285 11.7908
R16713 gnd.n1787 gnd.t212 11.4721
R16714 gnd.n4770 gnd.t321 11.4721
R16715 gnd.n4859 gnd.t181 11.4721
R16716 gnd.n3586 gnd.n3573 11.249
R16717 gnd.n3554 gnd.n3541 11.249
R16718 gnd.n3522 gnd.n3509 11.249
R16719 gnd.n3491 gnd.n3478 11.249
R16720 gnd.n3459 gnd.n3446 11.249
R16721 gnd.n3427 gnd.n3414 11.249
R16722 gnd.n3395 gnd.n3382 11.249
R16723 gnd.n3364 gnd.n3351 11.249
R16724 gnd.n3026 gnd.t4 11.1535
R16725 gnd.n4504 gnd.t352 11.1535
R16726 gnd.n4718 gnd.t323 11.1535
R16727 gnd.n4937 gnd.t9 11.1535
R16728 gnd.n5216 gnd.t192 11.1535
R16729 gnd.n4274 gnd.n886 10.8348
R16730 gnd.n6001 gnd.n896 10.8348
R16731 gnd.n4295 gnd.n4294 10.8348
R16732 gnd.n5995 gnd.n907 10.8348
R16733 gnd.n4283 gnd.n910 10.8348
R16734 gnd.n5989 gnd.n918 10.8348
R16735 gnd.n4340 gnd.n921 10.8348
R16736 gnd.n4347 gnd.n930 10.8348
R16737 gnd.n5977 gnd.n938 10.8348
R16738 gnd.n4355 gnd.n2057 10.8348
R16739 gnd.n5971 gnd.n947 10.8348
R16740 gnd.n4362 gnd.n950 10.8348
R16741 gnd.n5965 gnd.n958 10.8348
R16742 gnd.n4372 gnd.n961 10.8348
R16743 gnd.n5959 gnd.n968 10.8348
R16744 gnd.n4468 gnd.n971 10.8348
R16745 gnd.n4682 gnd.n4681 10.8348
R16746 gnd.n4818 gnd.n1608 10.8348
R16747 gnd.n4818 gnd.n1609 10.8348
R16748 gnd.n4997 gnd.n4996 10.8348
R16749 gnd.n5475 gnd.n5474 10.8348
R16750 gnd.n5285 gnd.n5274 10.8348
R16751 gnd.n5468 gnd.n5286 10.8348
R16752 gnd.n5467 gnd.n5289 10.8348
R16753 gnd.n5380 gnd.n5305 10.8348
R16754 gnd.n5461 gnd.n5308 10.8348
R16755 gnd.n5400 gnd.n5399 10.8348
R16756 gnd.n5455 gnd.n5319 10.8348
R16757 gnd.n5408 gnd.n5327 10.8348
R16758 gnd.n5426 gnd.n5334 10.8348
R16759 gnd.n5443 gnd.n5438 10.8348
R16760 gnd.n5417 gnd.n379 10.8348
R16761 gnd.n6735 gnd.n382 10.8348
R16762 gnd.n6722 gnd.n6721 10.8348
R16763 gnd.n6745 gnd.n371 10.8348
R16764 gnd.n6728 gnd.n363 10.8348
R16765 gnd.n6997 gnd.n6994 10.6672
R16766 gnd.n5598 gnd.n5595 10.6672
R16767 gnd.n3926 gnd.n3924 10.6672
R16768 gnd.n2047 gnd.n2046 10.6672
R16769 gnd.n5115 gnd.n1453 10.6151
R16770 gnd.n5115 gnd.n5114 10.6151
R16771 gnd.n5112 gnd.n1457 10.6151
R16772 gnd.n5107 gnd.n1457 10.6151
R16773 gnd.n5107 gnd.n5106 10.6151
R16774 gnd.n5106 gnd.n5105 10.6151
R16775 gnd.n5105 gnd.n1460 10.6151
R16776 gnd.n5100 gnd.n1460 10.6151
R16777 gnd.n5100 gnd.n5099 10.6151
R16778 gnd.n5099 gnd.n5098 10.6151
R16779 gnd.n5098 gnd.n1463 10.6151
R16780 gnd.n5093 gnd.n1463 10.6151
R16781 gnd.n5093 gnd.n5092 10.6151
R16782 gnd.n5092 gnd.n5091 10.6151
R16783 gnd.n5091 gnd.n1466 10.6151
R16784 gnd.n5086 gnd.n1466 10.6151
R16785 gnd.n5086 gnd.n5085 10.6151
R16786 gnd.n5085 gnd.n5084 10.6151
R16787 gnd.n5084 gnd.n1469 10.6151
R16788 gnd.n5079 gnd.n1469 10.6151
R16789 gnd.n5079 gnd.n5078 10.6151
R16790 gnd.n5078 gnd.n5077 10.6151
R16791 gnd.n5077 gnd.n1472 10.6151
R16792 gnd.n5072 gnd.n1472 10.6151
R16793 gnd.n5072 gnd.n5071 10.6151
R16794 gnd.n5071 gnd.n5070 10.6151
R16795 gnd.n5070 gnd.n1475 10.6151
R16796 gnd.n5065 gnd.n1475 10.6151
R16797 gnd.n5065 gnd.n5064 10.6151
R16798 gnd.n5064 gnd.n5063 10.6151
R16799 gnd.n1790 gnd.n1789 10.6151
R16800 gnd.n1791 gnd.n1790 10.6151
R16801 gnd.n1792 gnd.n1791 10.6151
R16802 gnd.n1792 gnd.n1721 10.6151
R16803 gnd.n4631 gnd.n1721 10.6151
R16804 gnd.n4632 gnd.n4631 10.6151
R16805 gnd.n4641 gnd.n4632 10.6151
R16806 gnd.n4641 gnd.n4640 10.6151
R16807 gnd.n4640 gnd.n4639 10.6151
R16808 gnd.n4639 gnd.n4638 10.6151
R16809 gnd.n4638 gnd.n4636 10.6151
R16810 gnd.n4636 gnd.n4635 10.6151
R16811 gnd.n4635 gnd.n1699 10.6151
R16812 gnd.n4673 gnd.n1699 10.6151
R16813 gnd.n4674 gnd.n4673 10.6151
R16814 gnd.n4679 gnd.n4674 10.6151
R16815 gnd.n4679 gnd.n4678 10.6151
R16816 gnd.n4678 gnd.n4677 10.6151
R16817 gnd.n4677 gnd.n4675 10.6151
R16818 gnd.n4675 gnd.n1672 10.6151
R16819 gnd.n4708 gnd.n1672 10.6151
R16820 gnd.n4709 gnd.n4708 10.6151
R16821 gnd.n4716 gnd.n4709 10.6151
R16822 gnd.n4716 gnd.n4715 10.6151
R16823 gnd.n4715 gnd.n4714 10.6151
R16824 gnd.n4714 gnd.n4713 10.6151
R16825 gnd.n4713 gnd.n4710 10.6151
R16826 gnd.n4710 gnd.n1647 10.6151
R16827 gnd.n4744 gnd.n1647 10.6151
R16828 gnd.n4745 gnd.n4744 10.6151
R16829 gnd.n4748 gnd.n4745 10.6151
R16830 gnd.n4748 gnd.n4747 10.6151
R16831 gnd.n4747 gnd.n4746 10.6151
R16832 gnd.n4746 gnd.n1629 10.6151
R16833 gnd.n4773 gnd.n1629 10.6151
R16834 gnd.n4774 gnd.n4773 10.6151
R16835 gnd.n4791 gnd.n4774 10.6151
R16836 gnd.n4791 gnd.n4790 10.6151
R16837 gnd.n4790 gnd.n4789 10.6151
R16838 gnd.n4789 gnd.n4775 10.6151
R16839 gnd.n4785 gnd.n4775 10.6151
R16840 gnd.n4785 gnd.n4784 10.6151
R16841 gnd.n4784 gnd.n4783 10.6151
R16842 gnd.n4783 gnd.n4782 10.6151
R16843 gnd.n4782 gnd.n4780 10.6151
R16844 gnd.n4780 gnd.n4779 10.6151
R16845 gnd.n4779 gnd.n4777 10.6151
R16846 gnd.n4777 gnd.n1575 10.6151
R16847 gnd.n4867 gnd.n1575 10.6151
R16848 gnd.n4868 gnd.n4867 10.6151
R16849 gnd.n4903 gnd.n4868 10.6151
R16850 gnd.n4903 gnd.n4902 10.6151
R16851 gnd.n4902 gnd.n4901 10.6151
R16852 gnd.n4901 gnd.n4900 10.6151
R16853 gnd.n4900 gnd.n4869 10.6151
R16854 gnd.n4895 gnd.n4869 10.6151
R16855 gnd.n4895 gnd.n4894 10.6151
R16856 gnd.n4894 gnd.n4893 10.6151
R16857 gnd.n4893 gnd.n4892 10.6151
R16858 gnd.n4892 gnd.n4890 10.6151
R16859 gnd.n4890 gnd.n4889 10.6151
R16860 gnd.n4889 gnd.n4873 10.6151
R16861 gnd.n4885 gnd.n4873 10.6151
R16862 gnd.n4885 gnd.n4884 10.6151
R16863 gnd.n4884 gnd.n4883 10.6151
R16864 gnd.n4883 gnd.n4882 10.6151
R16865 gnd.n4882 gnd.n4880 10.6151
R16866 gnd.n4880 gnd.n4879 10.6151
R16867 gnd.n4879 gnd.n4877 10.6151
R16868 gnd.n4877 gnd.n1503 10.6151
R16869 gnd.n5023 gnd.n1503 10.6151
R16870 gnd.n5024 gnd.n5023 10.6151
R16871 gnd.n5032 gnd.n5024 10.6151
R16872 gnd.n5032 gnd.n5031 10.6151
R16873 gnd.n5031 gnd.n5030 10.6151
R16874 gnd.n5030 gnd.n5029 10.6151
R16875 gnd.n5029 gnd.n5026 10.6151
R16876 gnd.n5026 gnd.n5025 10.6151
R16877 gnd.n5025 gnd.n1478 10.6151
R16878 gnd.n5059 gnd.n1478 10.6151
R16879 gnd.n5060 gnd.n5059 10.6151
R16880 gnd.n1724 gnd.n1048 10.6151
R16881 gnd.n1727 gnd.n1724 10.6151
R16882 gnd.n1732 gnd.n1729 10.6151
R16883 gnd.n1733 gnd.n1732 10.6151
R16884 gnd.n1736 gnd.n1733 10.6151
R16885 gnd.n1737 gnd.n1736 10.6151
R16886 gnd.n1740 gnd.n1737 10.6151
R16887 gnd.n1741 gnd.n1740 10.6151
R16888 gnd.n1744 gnd.n1741 10.6151
R16889 gnd.n1745 gnd.n1744 10.6151
R16890 gnd.n1748 gnd.n1745 10.6151
R16891 gnd.n1749 gnd.n1748 10.6151
R16892 gnd.n1752 gnd.n1749 10.6151
R16893 gnd.n1753 gnd.n1752 10.6151
R16894 gnd.n1756 gnd.n1753 10.6151
R16895 gnd.n1757 gnd.n1756 10.6151
R16896 gnd.n1760 gnd.n1757 10.6151
R16897 gnd.n1761 gnd.n1760 10.6151
R16898 gnd.n1764 gnd.n1761 10.6151
R16899 gnd.n1765 gnd.n1764 10.6151
R16900 gnd.n1768 gnd.n1765 10.6151
R16901 gnd.n1769 gnd.n1768 10.6151
R16902 gnd.n1772 gnd.n1769 10.6151
R16903 gnd.n1773 gnd.n1772 10.6151
R16904 gnd.n1776 gnd.n1773 10.6151
R16905 gnd.n1777 gnd.n1776 10.6151
R16906 gnd.n1780 gnd.n1777 10.6151
R16907 gnd.n1781 gnd.n1780 10.6151
R16908 gnd.n1784 gnd.n1781 10.6151
R16909 gnd.n1785 gnd.n1784 10.6151
R16910 gnd.n5894 gnd.n5893 10.6151
R16911 gnd.n5893 gnd.n5892 10.6151
R16912 gnd.n5892 gnd.n5891 10.6151
R16913 gnd.n5891 gnd.n5889 10.6151
R16914 gnd.n5889 gnd.n5886 10.6151
R16915 gnd.n5886 gnd.n5885 10.6151
R16916 gnd.n5885 gnd.n5882 10.6151
R16917 gnd.n5882 gnd.n5881 10.6151
R16918 gnd.n5881 gnd.n5878 10.6151
R16919 gnd.n5878 gnd.n5877 10.6151
R16920 gnd.n5877 gnd.n5874 10.6151
R16921 gnd.n5874 gnd.n5873 10.6151
R16922 gnd.n5873 gnd.n5870 10.6151
R16923 gnd.n5870 gnd.n5869 10.6151
R16924 gnd.n5869 gnd.n5866 10.6151
R16925 gnd.n5866 gnd.n5865 10.6151
R16926 gnd.n5865 gnd.n5862 10.6151
R16927 gnd.n5862 gnd.n5861 10.6151
R16928 gnd.n5861 gnd.n5858 10.6151
R16929 gnd.n5858 gnd.n5857 10.6151
R16930 gnd.n5857 gnd.n5854 10.6151
R16931 gnd.n5854 gnd.n5853 10.6151
R16932 gnd.n5853 gnd.n5850 10.6151
R16933 gnd.n5850 gnd.n5849 10.6151
R16934 gnd.n5849 gnd.n5846 10.6151
R16935 gnd.n5846 gnd.n5845 10.6151
R16936 gnd.n5845 gnd.n5842 10.6151
R16937 gnd.n5842 gnd.n5841 10.6151
R16938 gnd.n5838 gnd.n5837 10.6151
R16939 gnd.n5837 gnd.n1049 10.6151
R16940 gnd.n5179 gnd.n5178 10.6151
R16941 gnd.n5178 gnd.n1428 10.6151
R16942 gnd.n5173 gnd.n1428 10.6151
R16943 gnd.n5173 gnd.n5172 10.6151
R16944 gnd.n5172 gnd.n5171 10.6151
R16945 gnd.n5171 gnd.n1431 10.6151
R16946 gnd.n5166 gnd.n1431 10.6151
R16947 gnd.n5166 gnd.n5165 10.6151
R16948 gnd.n5165 gnd.n5164 10.6151
R16949 gnd.n5164 gnd.n1434 10.6151
R16950 gnd.n5159 gnd.n1434 10.6151
R16951 gnd.n5159 gnd.n5158 10.6151
R16952 gnd.n5158 gnd.n5157 10.6151
R16953 gnd.n5157 gnd.n1437 10.6151
R16954 gnd.n5152 gnd.n1437 10.6151
R16955 gnd.n5152 gnd.n5151 10.6151
R16956 gnd.n5151 gnd.n5150 10.6151
R16957 gnd.n5150 gnd.n1440 10.6151
R16958 gnd.n5145 gnd.n1440 10.6151
R16959 gnd.n5145 gnd.n5144 10.6151
R16960 gnd.n5144 gnd.n5143 10.6151
R16961 gnd.n5143 gnd.n1443 10.6151
R16962 gnd.n5138 gnd.n1443 10.6151
R16963 gnd.n5138 gnd.n5137 10.6151
R16964 gnd.n5137 gnd.n5136 10.6151
R16965 gnd.n5136 gnd.n1446 10.6151
R16966 gnd.n5131 gnd.n1446 10.6151
R16967 gnd.n5131 gnd.n5130 10.6151
R16968 gnd.n5128 gnd.n1451 10.6151
R16969 gnd.n5123 gnd.n1451 10.6151
R16970 gnd.n5830 gnd.n5829 10.6151
R16971 gnd.n5829 gnd.n1108 10.6151
R16972 gnd.n4624 gnd.n1108 10.6151
R16973 gnd.n4626 gnd.n4624 10.6151
R16974 gnd.n4626 gnd.n4625 10.6151
R16975 gnd.n4625 gnd.n1717 10.6151
R16976 gnd.n4645 gnd.n1717 10.6151
R16977 gnd.n4646 gnd.n4645 10.6151
R16978 gnd.n4647 gnd.n4646 10.6151
R16979 gnd.n4647 gnd.n1704 10.6151
R16980 gnd.n4666 gnd.n1704 10.6151
R16981 gnd.n4667 gnd.n4666 10.6151
R16982 gnd.n4668 gnd.n4667 10.6151
R16983 gnd.n4668 gnd.n1694 10.6151
R16984 gnd.n4685 gnd.n1694 10.6151
R16985 gnd.n4686 gnd.n4685 10.6151
R16986 gnd.n4687 gnd.n4686 10.6151
R16987 gnd.n4687 gnd.n1678 10.6151
R16988 gnd.n4702 gnd.n1678 10.6151
R16989 gnd.n4703 gnd.n4702 10.6151
R16990 gnd.n4704 gnd.n4703 10.6151
R16991 gnd.n4704 gnd.n1667 10.6151
R16992 gnd.n4720 gnd.n1667 10.6151
R16993 gnd.n4721 gnd.n4720 10.6151
R16994 gnd.n4722 gnd.n4721 10.6151
R16995 gnd.n4722 gnd.n1652 10.6151
R16996 gnd.n4737 gnd.n1652 10.6151
R16997 gnd.n4738 gnd.n4737 10.6151
R16998 gnd.n4740 gnd.n4738 10.6151
R16999 gnd.n4740 gnd.n4739 10.6151
R17000 gnd.n4739 gnd.n1633 10.6151
R17001 gnd.n4766 gnd.n1633 10.6151
R17002 gnd.n4767 gnd.n4766 10.6151
R17003 gnd.n4768 gnd.n4767 10.6151
R17004 gnd.n4768 gnd.n1624 10.6151
R17005 gnd.n4798 gnd.n1624 10.6151
R17006 gnd.n4799 gnd.n4798 10.6151
R17007 gnd.n4805 gnd.n4799 10.6151
R17008 gnd.n4805 gnd.n4804 10.6151
R17009 gnd.n4804 gnd.n4803 10.6151
R17010 gnd.n4803 gnd.n4800 10.6151
R17011 gnd.n4800 gnd.n1598 10.6151
R17012 gnd.n4843 gnd.n1598 10.6151
R17013 gnd.n4844 gnd.n4843 10.6151
R17014 gnd.n4845 gnd.n4844 10.6151
R17015 gnd.n4845 gnd.n1581 10.6151
R17016 gnd.n4861 gnd.n1581 10.6151
R17017 gnd.n4862 gnd.n4861 10.6151
R17018 gnd.n4863 gnd.n4862 10.6151
R17019 gnd.n4863 gnd.n1570 10.6151
R17020 gnd.n4907 gnd.n1570 10.6151
R17021 gnd.n4908 gnd.n4907 10.6151
R17022 gnd.n4914 gnd.n4908 10.6151
R17023 gnd.n4914 gnd.n4913 10.6151
R17024 gnd.n4913 gnd.n4912 10.6151
R17025 gnd.n4912 gnd.n4909 10.6151
R17026 gnd.n4909 gnd.n1546 10.6151
R17027 gnd.n4939 gnd.n1546 10.6151
R17028 gnd.n4940 gnd.n4939 10.6151
R17029 gnd.n4946 gnd.n4940 10.6151
R17030 gnd.n4946 gnd.n4945 10.6151
R17031 gnd.n4945 gnd.n4944 10.6151
R17032 gnd.n4944 gnd.n4941 10.6151
R17033 gnd.n4941 gnd.n1523 10.6151
R17034 gnd.n4999 gnd.n1523 10.6151
R17035 gnd.n5000 gnd.n4999 10.6151
R17036 gnd.n5001 gnd.n5000 10.6151
R17037 gnd.n5001 gnd.n1507 10.6151
R17038 gnd.n5017 gnd.n1507 10.6151
R17039 gnd.n5018 gnd.n5017 10.6151
R17040 gnd.n5019 gnd.n5018 10.6151
R17041 gnd.n5019 gnd.n1498 10.6151
R17042 gnd.n5036 gnd.n1498 10.6151
R17043 gnd.n5037 gnd.n5036 10.6151
R17044 gnd.n5038 gnd.n5037 10.6151
R17045 gnd.n5038 gnd.n1482 10.6151
R17046 gnd.n5052 gnd.n1482 10.6151
R17047 gnd.n5053 gnd.n5052 10.6151
R17048 gnd.n5054 gnd.n5053 10.6151
R17049 gnd.n5054 gnd.n1408 10.6151
R17050 gnd.n5181 gnd.n1408 10.6151
R17051 gnd.n2945 gnd.t2 10.5161
R17052 gnd.n2374 gnd.t6 10.5161
R17053 gnd.n3311 gnd.t332 10.5161
R17054 gnd.t323 gnd.n1662 10.5161
R17055 gnd.n4871 gnd.t9 10.5161
R17056 gnd.n3587 gnd.n3571 10.4732
R17057 gnd.n3555 gnd.n3539 10.4732
R17058 gnd.n3523 gnd.n3507 10.4732
R17059 gnd.n3492 gnd.n3476 10.4732
R17060 gnd.n3460 gnd.n3444 10.4732
R17061 gnd.n3428 gnd.n3412 10.4732
R17062 gnd.n3396 gnd.n3380 10.4732
R17063 gnd.n3365 gnd.n3349 10.4732
R17064 gnd.t338 gnd.n2391 9.87883
R17065 gnd.n4808 gnd.t350 9.87883
R17066 gnd.n4840 gnd.t348 9.87883
R17067 gnd.n3591 gnd.n3590 9.69747
R17068 gnd.n3559 gnd.n3558 9.69747
R17069 gnd.n3527 gnd.n3526 9.69747
R17070 gnd.n3496 gnd.n3495 9.69747
R17071 gnd.n3464 gnd.n3463 9.69747
R17072 gnd.n3432 gnd.n3431 9.69747
R17073 gnd.n3400 gnd.n3399 9.69747
R17074 gnd.n3369 gnd.n3368 9.69747
R17075 gnd.n4670 gnd.n1702 9.56018
R17076 gnd.n1692 gnd.n1681 9.56018
R17077 gnd.n4808 gnd.n4807 9.56018
R17078 gnd.n4841 gnd.n4840 9.56018
R17079 gnd.n4960 gnd.n1532 9.56018
R17080 gnd.n1521 gnd.n1509 9.56018
R17081 gnd.n5034 gnd.t254 9.56018
R17082 gnd.n3597 gnd.n3596 9.45567
R17083 gnd.n3565 gnd.n3564 9.45567
R17084 gnd.n3533 gnd.n3532 9.45567
R17085 gnd.n3502 gnd.n3501 9.45567
R17086 gnd.n3470 gnd.n3469 9.45567
R17087 gnd.n3438 gnd.n3437 9.45567
R17088 gnd.n3406 gnd.n3405 9.45567
R17089 gnd.n3375 gnd.n3374 9.45567
R17090 gnd.n7036 gnd.n285 9.30959
R17091 gnd.n5635 gnd.n5634 9.30959
R17092 gnd.n3963 gnd.n3962 9.30959
R17093 gnd.n2001 gnd.n1998 9.30959
R17094 gnd.n5595 gnd.n5594 9.3005
R17095 gnd.n5598 gnd.n1343 9.3005
R17096 gnd.n5599 gnd.n1342 9.3005
R17097 gnd.n5602 gnd.n1341 9.3005
R17098 gnd.n5603 gnd.n1340 9.3005
R17099 gnd.n5606 gnd.n1339 9.3005
R17100 gnd.n5607 gnd.n1338 9.3005
R17101 gnd.n5610 gnd.n1337 9.3005
R17102 gnd.n5611 gnd.n1336 9.3005
R17103 gnd.n5614 gnd.n1335 9.3005
R17104 gnd.n5615 gnd.n1334 9.3005
R17105 gnd.n5618 gnd.n1333 9.3005
R17106 gnd.n5619 gnd.n1332 9.3005
R17107 gnd.n5622 gnd.n1331 9.3005
R17108 gnd.n5623 gnd.n1330 9.3005
R17109 gnd.n5626 gnd.n1329 9.3005
R17110 gnd.n5627 gnd.n1328 9.3005
R17111 gnd.n5630 gnd.n1327 9.3005
R17112 gnd.n5631 gnd.n1326 9.3005
R17113 gnd.n5634 gnd.n1325 9.3005
R17114 gnd.n5638 gnd.n1321 9.3005
R17115 gnd.n5639 gnd.n1320 9.3005
R17116 gnd.n5642 gnd.n1319 9.3005
R17117 gnd.n5643 gnd.n1318 9.3005
R17118 gnd.n5646 gnd.n1317 9.3005
R17119 gnd.n5647 gnd.n1316 9.3005
R17120 gnd.n5650 gnd.n1315 9.3005
R17121 gnd.n5651 gnd.n1314 9.3005
R17122 gnd.n5654 gnd.n1313 9.3005
R17123 gnd.n5656 gnd.n1309 9.3005
R17124 gnd.n5659 gnd.n1308 9.3005
R17125 gnd.n5660 gnd.n1307 9.3005
R17126 gnd.n5663 gnd.n1306 9.3005
R17127 gnd.n5664 gnd.n1305 9.3005
R17128 gnd.n5667 gnd.n1304 9.3005
R17129 gnd.n5668 gnd.n1303 9.3005
R17130 gnd.n5671 gnd.n1302 9.3005
R17131 gnd.n5673 gnd.n1299 9.3005
R17132 gnd.n5676 gnd.n1298 9.3005
R17133 gnd.n5677 gnd.n1297 9.3005
R17134 gnd.n5680 gnd.n1296 9.3005
R17135 gnd.n5681 gnd.n1295 9.3005
R17136 gnd.n5684 gnd.n1294 9.3005
R17137 gnd.n5685 gnd.n1293 9.3005
R17138 gnd.n5688 gnd.n1292 9.3005
R17139 gnd.n5689 gnd.n1291 9.3005
R17140 gnd.n5692 gnd.n1290 9.3005
R17141 gnd.n5693 gnd.n1289 9.3005
R17142 gnd.n5696 gnd.n1288 9.3005
R17143 gnd.n5697 gnd.n1287 9.3005
R17144 gnd.n5700 gnd.n1286 9.3005
R17145 gnd.n5702 gnd.n1285 9.3005
R17146 gnd.n5703 gnd.n1284 9.3005
R17147 gnd.n5704 gnd.n1283 9.3005
R17148 gnd.n5705 gnd.n1282 9.3005
R17149 gnd.n5635 gnd.n1322 9.3005
R17150 gnd.n5593 gnd.n1344 9.3005
R17151 gnd.n5298 gnd.n5297 9.3005
R17152 gnd.n5299 gnd.n5293 9.3005
R17153 gnd.n5465 gnd.n5300 9.3005
R17154 gnd.n5464 gnd.n5301 9.3005
R17155 gnd.n5463 gnd.n5302 9.3005
R17156 gnd.n5321 gnd.n5303 9.3005
R17157 gnd.n5453 gnd.n5322 9.3005
R17158 gnd.n5452 gnd.n5323 9.3005
R17159 gnd.n5451 gnd.n5324 9.3005
R17160 gnd.n5439 gnd.n5325 9.3005
R17161 gnd.n5441 gnd.n5440 9.3005
R17162 gnd.n377 gnd.n376 9.3005
R17163 gnd.n6738 gnd.n6737 9.3005
R17164 gnd.n6739 gnd.n375 9.3005
R17165 gnd.n6743 gnd.n6740 9.3005
R17166 gnd.n6742 gnd.n6741 9.3005
R17167 gnd.n349 gnd.n348 9.3005
R17168 gnd.n6772 gnd.n6771 9.3005
R17169 gnd.n6773 gnd.n347 9.3005
R17170 gnd.n6777 gnd.n6774 9.3005
R17171 gnd.n6776 gnd.n6775 9.3005
R17172 gnd.n5295 gnd.n5294 9.3005
R17173 gnd.n327 gnd.n326 9.3005
R17174 gnd.n6805 gnd.n6804 9.3005
R17175 gnd.n6806 gnd.n325 9.3005
R17176 gnd.n6811 gnd.n6807 9.3005
R17177 gnd.n6810 gnd.n6809 9.3005
R17178 gnd.n6808 gnd.n90 9.3005
R17179 gnd.n7189 gnd.n91 9.3005
R17180 gnd.n7188 gnd.n92 9.3005
R17181 gnd.n7187 gnd.n93 9.3005
R17182 gnd.n111 gnd.n94 9.3005
R17183 gnd.n7177 gnd.n112 9.3005
R17184 gnd.n7176 gnd.n113 9.3005
R17185 gnd.n7175 gnd.n114 9.3005
R17186 gnd.n130 gnd.n115 9.3005
R17187 gnd.n7165 gnd.n131 9.3005
R17188 gnd.n7164 gnd.n132 9.3005
R17189 gnd.n7163 gnd.n133 9.3005
R17190 gnd.n149 gnd.n134 9.3005
R17191 gnd.n7153 gnd.n150 9.3005
R17192 gnd.n7152 gnd.n151 9.3005
R17193 gnd.n7151 gnd.n152 9.3005
R17194 gnd.n168 gnd.n153 9.3005
R17195 gnd.n7141 gnd.n169 9.3005
R17196 gnd.n7140 gnd.n170 9.3005
R17197 gnd.n7139 gnd.n171 9.3005
R17198 gnd.n187 gnd.n172 9.3005
R17199 gnd.n7129 gnd.n188 9.3005
R17200 gnd.n7128 gnd.n189 9.3005
R17201 gnd.n7127 gnd.n190 9.3005
R17202 gnd.n206 gnd.n191 9.3005
R17203 gnd.n7117 gnd.n207 9.3005
R17204 gnd.n7116 gnd.n7115 9.3005
R17205 gnd.n7195 gnd.n7194 9.3005
R17206 gnd.n7193 gnd.n80 9.3005
R17207 gnd.n6858 gnd.n83 9.3005
R17208 gnd.n6859 gnd.n6857 9.3005
R17209 gnd.n6862 gnd.n6860 9.3005
R17210 gnd.n6863 gnd.n6856 9.3005
R17211 gnd.n6866 gnd.n6865 9.3005
R17212 gnd.n6867 gnd.n6855 9.3005
R17213 gnd.n6870 gnd.n6868 9.3005
R17214 gnd.n6871 gnd.n6854 9.3005
R17215 gnd.n6874 gnd.n6873 9.3005
R17216 gnd.n6875 gnd.n6853 9.3005
R17217 gnd.n6878 gnd.n6876 9.3005
R17218 gnd.n6879 gnd.n6852 9.3005
R17219 gnd.n6882 gnd.n6881 9.3005
R17220 gnd.n6883 gnd.n6851 9.3005
R17221 gnd.n6967 gnd.n6884 9.3005
R17222 gnd.n6966 gnd.n6885 9.3005
R17223 gnd.n6965 gnd.n6886 9.3005
R17224 gnd.n6963 gnd.n6887 9.3005
R17225 gnd.n6962 gnd.n6888 9.3005
R17226 gnd.n6960 gnd.n6889 9.3005
R17227 gnd.n6959 gnd.n6890 9.3005
R17228 gnd.n6957 gnd.n6891 9.3005
R17229 gnd.n6956 gnd.n6892 9.3005
R17230 gnd.n6954 gnd.n6893 9.3005
R17231 gnd.n6953 gnd.n6894 9.3005
R17232 gnd.n6908 gnd.n6907 9.3005
R17233 gnd.n6910 gnd.n6909 9.3005
R17234 gnd.n6913 gnd.n6904 9.3005
R17235 gnd.n6917 gnd.n6916 9.3005
R17236 gnd.n6918 gnd.n6903 9.3005
R17237 gnd.n6920 gnd.n6919 9.3005
R17238 gnd.n6923 gnd.n6902 9.3005
R17239 gnd.n6927 gnd.n6926 9.3005
R17240 gnd.n6928 gnd.n6901 9.3005
R17241 gnd.n6930 gnd.n6929 9.3005
R17242 gnd.n6933 gnd.n6900 9.3005
R17243 gnd.n6937 gnd.n6936 9.3005
R17244 gnd.n6938 gnd.n6899 9.3005
R17245 gnd.n6940 gnd.n6939 9.3005
R17246 gnd.n6943 gnd.n6898 9.3005
R17247 gnd.n6947 gnd.n6946 9.3005
R17248 gnd.n6948 gnd.n6897 9.3005
R17249 gnd.n6950 gnd.n6949 9.3005
R17250 gnd.n6905 gnd.n308 9.3005
R17251 gnd.n209 gnd.n208 9.3005
R17252 gnd.n7108 gnd.n250 9.3005
R17253 gnd.n7107 gnd.n251 9.3005
R17254 gnd.n7106 gnd.n252 9.3005
R17255 gnd.n7103 gnd.n253 9.3005
R17256 gnd.n7102 gnd.n254 9.3005
R17257 gnd.n7099 gnd.n255 9.3005
R17258 gnd.n7098 gnd.n256 9.3005
R17259 gnd.n7095 gnd.n257 9.3005
R17260 gnd.n7094 gnd.n258 9.3005
R17261 gnd.n7091 gnd.n259 9.3005
R17262 gnd.n7090 gnd.n260 9.3005
R17263 gnd.n7087 gnd.n261 9.3005
R17264 gnd.n7086 gnd.n262 9.3005
R17265 gnd.n7083 gnd.n263 9.3005
R17266 gnd.n7082 gnd.n264 9.3005
R17267 gnd.n7079 gnd.n265 9.3005
R17268 gnd.n7075 gnd.n266 9.3005
R17269 gnd.n7072 gnd.n267 9.3005
R17270 gnd.n7071 gnd.n268 9.3005
R17271 gnd.n7068 gnd.n269 9.3005
R17272 gnd.n7067 gnd.n270 9.3005
R17273 gnd.n7064 gnd.n271 9.3005
R17274 gnd.n7063 gnd.n272 9.3005
R17275 gnd.n7060 gnd.n273 9.3005
R17276 gnd.n7059 gnd.n274 9.3005
R17277 gnd.n7056 gnd.n275 9.3005
R17278 gnd.n7055 gnd.n276 9.3005
R17279 gnd.n7052 gnd.n277 9.3005
R17280 gnd.n7051 gnd.n278 9.3005
R17281 gnd.n7048 gnd.n279 9.3005
R17282 gnd.n7047 gnd.n280 9.3005
R17283 gnd.n7044 gnd.n281 9.3005
R17284 gnd.n7043 gnd.n282 9.3005
R17285 gnd.n7040 gnd.n283 9.3005
R17286 gnd.n7039 gnd.n284 9.3005
R17287 gnd.n7036 gnd.n7035 9.3005
R17288 gnd.n7034 gnd.n285 9.3005
R17289 gnd.n7033 gnd.n7032 9.3005
R17290 gnd.n7029 gnd.n288 9.3005
R17291 gnd.n7026 gnd.n289 9.3005
R17292 gnd.n7025 gnd.n290 9.3005
R17293 gnd.n7022 gnd.n291 9.3005
R17294 gnd.n7021 gnd.n292 9.3005
R17295 gnd.n7018 gnd.n293 9.3005
R17296 gnd.n7017 gnd.n294 9.3005
R17297 gnd.n7014 gnd.n295 9.3005
R17298 gnd.n7013 gnd.n296 9.3005
R17299 gnd.n7010 gnd.n297 9.3005
R17300 gnd.n7009 gnd.n298 9.3005
R17301 gnd.n7006 gnd.n299 9.3005
R17302 gnd.n7005 gnd.n300 9.3005
R17303 gnd.n7002 gnd.n301 9.3005
R17304 gnd.n7001 gnd.n302 9.3005
R17305 gnd.n6998 gnd.n303 9.3005
R17306 gnd.n6997 gnd.n304 9.3005
R17307 gnd.n6994 gnd.n6993 9.3005
R17308 gnd.n6992 gnd.n305 9.3005
R17309 gnd.n7114 gnd.n7113 9.3005
R17310 gnd.n5360 gnd.n5359 9.3005
R17311 gnd.n5358 gnd.n5354 9.3005
R17312 gnd.n5365 gnd.n5353 9.3005
R17313 gnd.n5382 gnd.n5366 9.3005
R17314 gnd.n5383 gnd.n5312 9.3005
R17315 gnd.n5384 gnd.n5313 9.3005
R17316 gnd.n5348 gnd.n5314 9.3005
R17317 gnd.n5410 gnd.n5349 9.3005
R17318 gnd.n5411 gnd.n5331 9.3005
R17319 gnd.n5412 gnd.n5332 9.3005
R17320 gnd.n5413 gnd.n5333 9.3005
R17321 gnd.n5415 gnd.n5414 9.3005
R17322 gnd.n388 gnd.n386 9.3005
R17323 gnd.n6724 gnd.n387 9.3005
R17324 gnd.n6726 gnd.n6725 9.3005
R17325 gnd.n6727 gnd.n360 9.3005
R17326 gnd.n6756 gnd.n361 9.3005
R17327 gnd.n6757 gnd.n358 9.3005
R17328 gnd.n6759 gnd.n359 9.3005
R17329 gnd.n6761 gnd.n6760 9.3005
R17330 gnd.n6762 gnd.n334 9.3005
R17331 gnd.n6795 gnd.n333 9.3005
R17332 gnd.n6799 gnd.n6798 9.3005
R17333 gnd.n6797 gnd.n316 9.3005
R17334 gnd.n6816 gnd.n315 9.3005
R17335 gnd.n6818 gnd.n6817 9.3005
R17336 gnd.n6819 gnd.n310 9.3005
R17337 gnd.n6825 gnd.n309 9.3005
R17338 gnd.n6828 gnd.n6826 9.3005
R17339 gnd.n6829 gnd.n101 9.3005
R17340 gnd.n6831 gnd.n102 9.3005
R17341 gnd.n6832 gnd.n103 9.3005
R17342 gnd.n6835 gnd.n6833 9.3005
R17343 gnd.n6836 gnd.n121 9.3005
R17344 gnd.n6838 gnd.n122 9.3005
R17345 gnd.n6839 gnd.n123 9.3005
R17346 gnd.n6842 gnd.n6840 9.3005
R17347 gnd.n6843 gnd.n139 9.3005
R17348 gnd.n6845 gnd.n140 9.3005
R17349 gnd.n6846 gnd.n141 9.3005
R17350 gnd.n6849 gnd.n6847 9.3005
R17351 gnd.n6850 gnd.n159 9.3005
R17352 gnd.n6971 gnd.n160 9.3005
R17353 gnd.n6972 gnd.n161 9.3005
R17354 gnd.n6975 gnd.n6973 9.3005
R17355 gnd.n6976 gnd.n177 9.3005
R17356 gnd.n6978 gnd.n178 9.3005
R17357 gnd.n6979 gnd.n179 9.3005
R17358 gnd.n6982 gnd.n6980 9.3005
R17359 gnd.n6983 gnd.n197 9.3005
R17360 gnd.n6985 gnd.n198 9.3005
R17361 gnd.n6986 gnd.n199 9.3005
R17362 gnd.n6990 gnd.n6989 9.3005
R17363 gnd.n5355 gnd.n1347 9.3005
R17364 gnd.n5361 gnd.n5360 9.3005
R17365 gnd.n5363 gnd.n5354 9.3005
R17366 gnd.n5365 gnd.n5364 9.3005
R17367 gnd.n5366 gnd.n5311 9.3005
R17368 gnd.n5459 gnd.n5312 9.3005
R17369 gnd.n5458 gnd.n5313 9.3005
R17370 gnd.n5457 gnd.n5314 9.3005
R17371 gnd.n5349 gnd.n5315 9.3005
R17372 gnd.n5447 gnd.n5331 9.3005
R17373 gnd.n5446 gnd.n5332 9.3005
R17374 gnd.n5445 gnd.n5333 9.3005
R17375 gnd.n5414 gnd.n385 9.3005
R17376 gnd.n6733 gnd.n386 9.3005
R17377 gnd.n6732 gnd.n387 9.3005
R17378 gnd.n6731 gnd.n6726 9.3005
R17379 gnd.n6730 gnd.n6727 9.3005
R17380 gnd.n361 gnd.n357 9.3005
R17381 gnd.n6767 gnd.n358 9.3005
R17382 gnd.n6766 gnd.n359 9.3005
R17383 gnd.n6765 gnd.n6761 9.3005
R17384 gnd.n6764 gnd.n6762 9.3005
R17385 gnd.n333 gnd.n332 9.3005
R17386 gnd.n6800 gnd.n6799 9.3005
R17387 gnd.n317 gnd.n316 9.3005
R17388 gnd.n6816 gnd.n6815 9.3005
R17389 gnd.n6817 gnd.n311 9.3005
R17390 gnd.n6823 gnd.n310 9.3005
R17391 gnd.n6825 gnd.n6824 9.3005
R17392 gnd.n6826 gnd.n100 9.3005
R17393 gnd.n7183 gnd.n101 9.3005
R17394 gnd.n7182 gnd.n102 9.3005
R17395 gnd.n7181 gnd.n103 9.3005
R17396 gnd.n6833 gnd.n104 9.3005
R17397 gnd.n7171 gnd.n121 9.3005
R17398 gnd.n7170 gnd.n122 9.3005
R17399 gnd.n7169 gnd.n123 9.3005
R17400 gnd.n6840 gnd.n124 9.3005
R17401 gnd.n7159 gnd.n139 9.3005
R17402 gnd.n7158 gnd.n140 9.3005
R17403 gnd.n7157 gnd.n141 9.3005
R17404 gnd.n6847 gnd.n142 9.3005
R17405 gnd.n7147 gnd.n159 9.3005
R17406 gnd.n7146 gnd.n160 9.3005
R17407 gnd.n7145 gnd.n161 9.3005
R17408 gnd.n6973 gnd.n162 9.3005
R17409 gnd.n7135 gnd.n177 9.3005
R17410 gnd.n7134 gnd.n178 9.3005
R17411 gnd.n7133 gnd.n179 9.3005
R17412 gnd.n6980 gnd.n180 9.3005
R17413 gnd.n7123 gnd.n197 9.3005
R17414 gnd.n7122 gnd.n198 9.3005
R17415 gnd.n7121 gnd.n199 9.3005
R17416 gnd.n6990 gnd.n200 9.3005
R17417 gnd.n5269 gnd.n1347 9.3005
R17418 gnd.n3596 gnd.n3595 9.3005
R17419 gnd.n3569 gnd.n3568 9.3005
R17420 gnd.n3590 gnd.n3589 9.3005
R17421 gnd.n3588 gnd.n3587 9.3005
R17422 gnd.n3573 gnd.n3572 9.3005
R17423 gnd.n3582 gnd.n3581 9.3005
R17424 gnd.n3580 gnd.n3579 9.3005
R17425 gnd.n3564 gnd.n3563 9.3005
R17426 gnd.n3537 gnd.n3536 9.3005
R17427 gnd.n3558 gnd.n3557 9.3005
R17428 gnd.n3556 gnd.n3555 9.3005
R17429 gnd.n3541 gnd.n3540 9.3005
R17430 gnd.n3550 gnd.n3549 9.3005
R17431 gnd.n3548 gnd.n3547 9.3005
R17432 gnd.n3532 gnd.n3531 9.3005
R17433 gnd.n3505 gnd.n3504 9.3005
R17434 gnd.n3526 gnd.n3525 9.3005
R17435 gnd.n3524 gnd.n3523 9.3005
R17436 gnd.n3509 gnd.n3508 9.3005
R17437 gnd.n3518 gnd.n3517 9.3005
R17438 gnd.n3516 gnd.n3515 9.3005
R17439 gnd.n3501 gnd.n3500 9.3005
R17440 gnd.n3474 gnd.n3473 9.3005
R17441 gnd.n3495 gnd.n3494 9.3005
R17442 gnd.n3493 gnd.n3492 9.3005
R17443 gnd.n3478 gnd.n3477 9.3005
R17444 gnd.n3487 gnd.n3486 9.3005
R17445 gnd.n3485 gnd.n3484 9.3005
R17446 gnd.n3469 gnd.n3468 9.3005
R17447 gnd.n3442 gnd.n3441 9.3005
R17448 gnd.n3463 gnd.n3462 9.3005
R17449 gnd.n3461 gnd.n3460 9.3005
R17450 gnd.n3446 gnd.n3445 9.3005
R17451 gnd.n3455 gnd.n3454 9.3005
R17452 gnd.n3453 gnd.n3452 9.3005
R17453 gnd.n3437 gnd.n3436 9.3005
R17454 gnd.n3410 gnd.n3409 9.3005
R17455 gnd.n3431 gnd.n3430 9.3005
R17456 gnd.n3429 gnd.n3428 9.3005
R17457 gnd.n3414 gnd.n3413 9.3005
R17458 gnd.n3423 gnd.n3422 9.3005
R17459 gnd.n3421 gnd.n3420 9.3005
R17460 gnd.n3405 gnd.n3404 9.3005
R17461 gnd.n3378 gnd.n3377 9.3005
R17462 gnd.n3399 gnd.n3398 9.3005
R17463 gnd.n3397 gnd.n3396 9.3005
R17464 gnd.n3382 gnd.n3381 9.3005
R17465 gnd.n3391 gnd.n3390 9.3005
R17466 gnd.n3389 gnd.n3388 9.3005
R17467 gnd.n3374 gnd.n3373 9.3005
R17468 gnd.n3347 gnd.n3346 9.3005
R17469 gnd.n3368 gnd.n3367 9.3005
R17470 gnd.n3366 gnd.n3365 9.3005
R17471 gnd.n3351 gnd.n3350 9.3005
R17472 gnd.n3360 gnd.n3359 9.3005
R17473 gnd.n3358 gnd.n3357 9.3005
R17474 gnd.n3722 gnd.n3721 9.3005
R17475 gnd.n3720 gnd.n2273 9.3005
R17476 gnd.n3719 gnd.n3718 9.3005
R17477 gnd.n3715 gnd.n2274 9.3005
R17478 gnd.n3712 gnd.n2275 9.3005
R17479 gnd.n3711 gnd.n2276 9.3005
R17480 gnd.n3708 gnd.n2277 9.3005
R17481 gnd.n3707 gnd.n2278 9.3005
R17482 gnd.n3704 gnd.n2279 9.3005
R17483 gnd.n3703 gnd.n2280 9.3005
R17484 gnd.n3700 gnd.n2281 9.3005
R17485 gnd.n3699 gnd.n2282 9.3005
R17486 gnd.n3696 gnd.n2283 9.3005
R17487 gnd.n3695 gnd.n2284 9.3005
R17488 gnd.n3692 gnd.n3691 9.3005
R17489 gnd.n3690 gnd.n2285 9.3005
R17490 gnd.n3723 gnd.n2272 9.3005
R17491 gnd.n2964 gnd.n2963 9.3005
R17492 gnd.n2668 gnd.n2667 9.3005
R17493 gnd.n2991 gnd.n2990 9.3005
R17494 gnd.n2992 gnd.n2666 9.3005
R17495 gnd.n2996 gnd.n2993 9.3005
R17496 gnd.n2995 gnd.n2994 9.3005
R17497 gnd.n2640 gnd.n2639 9.3005
R17498 gnd.n3021 gnd.n3020 9.3005
R17499 gnd.n3022 gnd.n2638 9.3005
R17500 gnd.n3024 gnd.n3023 9.3005
R17501 gnd.n2618 gnd.n2617 9.3005
R17502 gnd.n3052 gnd.n3051 9.3005
R17503 gnd.n3053 gnd.n2616 9.3005
R17504 gnd.n3061 gnd.n3054 9.3005
R17505 gnd.n3060 gnd.n3055 9.3005
R17506 gnd.n3059 gnd.n3057 9.3005
R17507 gnd.n3056 gnd.n2565 9.3005
R17508 gnd.n3109 gnd.n2566 9.3005
R17509 gnd.n3108 gnd.n2567 9.3005
R17510 gnd.n3107 gnd.n2568 9.3005
R17511 gnd.n2587 gnd.n2569 9.3005
R17512 gnd.n2589 gnd.n2588 9.3005
R17513 gnd.n2471 gnd.n2470 9.3005
R17514 gnd.n3147 gnd.n3146 9.3005
R17515 gnd.n3148 gnd.n2469 9.3005
R17516 gnd.n3152 gnd.n3149 9.3005
R17517 gnd.n3151 gnd.n3150 9.3005
R17518 gnd.n2444 gnd.n2443 9.3005
R17519 gnd.n3187 gnd.n3186 9.3005
R17520 gnd.n3188 gnd.n2442 9.3005
R17521 gnd.n3192 gnd.n3189 9.3005
R17522 gnd.n3191 gnd.n3190 9.3005
R17523 gnd.n2417 gnd.n2416 9.3005
R17524 gnd.n3232 gnd.n3231 9.3005
R17525 gnd.n3233 gnd.n2415 9.3005
R17526 gnd.n3237 gnd.n3234 9.3005
R17527 gnd.n3236 gnd.n3235 9.3005
R17528 gnd.n2389 gnd.n2388 9.3005
R17529 gnd.n3272 gnd.n3271 9.3005
R17530 gnd.n3273 gnd.n2387 9.3005
R17531 gnd.n3277 gnd.n3274 9.3005
R17532 gnd.n3276 gnd.n3275 9.3005
R17533 gnd.n2362 gnd.n2361 9.3005
R17534 gnd.n3321 gnd.n3320 9.3005
R17535 gnd.n3322 gnd.n2360 9.3005
R17536 gnd.n3326 gnd.n3323 9.3005
R17537 gnd.n3325 gnd.n3324 9.3005
R17538 gnd.n2335 gnd.n2334 9.3005
R17539 gnd.n3615 gnd.n3614 9.3005
R17540 gnd.n3616 gnd.n2333 9.3005
R17541 gnd.n3622 gnd.n3617 9.3005
R17542 gnd.n3621 gnd.n3618 9.3005
R17543 gnd.n3620 gnd.n3619 9.3005
R17544 gnd.n2965 gnd.n2962 9.3005
R17545 gnd.n2747 gnd.n2706 9.3005
R17546 gnd.n2742 gnd.n2741 9.3005
R17547 gnd.n2740 gnd.n2707 9.3005
R17548 gnd.n2739 gnd.n2738 9.3005
R17549 gnd.n2735 gnd.n2708 9.3005
R17550 gnd.n2732 gnd.n2731 9.3005
R17551 gnd.n2730 gnd.n2709 9.3005
R17552 gnd.n2729 gnd.n2728 9.3005
R17553 gnd.n2725 gnd.n2710 9.3005
R17554 gnd.n2722 gnd.n2721 9.3005
R17555 gnd.n2720 gnd.n2711 9.3005
R17556 gnd.n2719 gnd.n2718 9.3005
R17557 gnd.n2715 gnd.n2713 9.3005
R17558 gnd.n2712 gnd.n2692 9.3005
R17559 gnd.n2959 gnd.n2691 9.3005
R17560 gnd.n2961 gnd.n2960 9.3005
R17561 gnd.n2749 gnd.n2748 9.3005
R17562 gnd.n2972 gnd.n2678 9.3005
R17563 gnd.n2979 gnd.n2679 9.3005
R17564 gnd.n2981 gnd.n2980 9.3005
R17565 gnd.n2982 gnd.n2659 9.3005
R17566 gnd.n3001 gnd.n3000 9.3005
R17567 gnd.n3003 gnd.n2651 9.3005
R17568 gnd.n3010 gnd.n2653 9.3005
R17569 gnd.n3011 gnd.n2648 9.3005
R17570 gnd.n3013 gnd.n3012 9.3005
R17571 gnd.n2649 gnd.n2634 9.3005
R17572 gnd.n3029 gnd.n2632 9.3005
R17573 gnd.n3033 gnd.n3032 9.3005
R17574 gnd.n3031 gnd.n2608 9.3005
R17575 gnd.n3068 gnd.n2607 9.3005
R17576 gnd.n3071 gnd.n3070 9.3005
R17577 gnd.n2604 gnd.n2603 9.3005
R17578 gnd.n3077 gnd.n2605 9.3005
R17579 gnd.n3079 gnd.n3078 9.3005
R17580 gnd.n3081 gnd.n2602 9.3005
R17581 gnd.n3084 gnd.n3083 9.3005
R17582 gnd.n3087 gnd.n3085 9.3005
R17583 gnd.n3089 gnd.n3088 9.3005
R17584 gnd.n3095 gnd.n3090 9.3005
R17585 gnd.n3094 gnd.n3093 9.3005
R17586 gnd.n2462 gnd.n2461 9.3005
R17587 gnd.n3161 gnd.n3160 9.3005
R17588 gnd.n3162 gnd.n2455 9.3005
R17589 gnd.n3170 gnd.n2454 9.3005
R17590 gnd.n3173 gnd.n3172 9.3005
R17591 gnd.n3175 gnd.n3174 9.3005
R17592 gnd.n3178 gnd.n2437 9.3005
R17593 gnd.n3176 gnd.n2435 9.3005
R17594 gnd.n3198 gnd.n2433 9.3005
R17595 gnd.n3200 gnd.n3199 9.3005
R17596 gnd.n2407 gnd.n2406 9.3005
R17597 gnd.n3246 gnd.n3245 9.3005
R17598 gnd.n3247 gnd.n2400 9.3005
R17599 gnd.n3255 gnd.n2399 9.3005
R17600 gnd.n3258 gnd.n3257 9.3005
R17601 gnd.n3260 gnd.n3259 9.3005
R17602 gnd.n3263 gnd.n2382 9.3005
R17603 gnd.n3261 gnd.n2380 9.3005
R17604 gnd.n3283 gnd.n2378 9.3005
R17605 gnd.n3285 gnd.n3284 9.3005
R17606 gnd.n2353 gnd.n2352 9.3005
R17607 gnd.n3335 gnd.n3334 9.3005
R17608 gnd.n3336 gnd.n2346 9.3005
R17609 gnd.n3344 gnd.n2345 9.3005
R17610 gnd.n3603 gnd.n3602 9.3005
R17611 gnd.n3605 gnd.n3604 9.3005
R17612 gnd.n3606 gnd.n2326 9.3005
R17613 gnd.n3630 gnd.n3629 9.3005
R17614 gnd.n2327 gnd.n2288 9.3005
R17615 gnd.n2970 gnd.n2969 9.3005
R17616 gnd.n3686 gnd.n2289 9.3005
R17617 gnd.n3685 gnd.n2291 9.3005
R17618 gnd.n3682 gnd.n2292 9.3005
R17619 gnd.n3681 gnd.n2293 9.3005
R17620 gnd.n3678 gnd.n2294 9.3005
R17621 gnd.n3677 gnd.n2295 9.3005
R17622 gnd.n3674 gnd.n2296 9.3005
R17623 gnd.n3673 gnd.n2297 9.3005
R17624 gnd.n3670 gnd.n2298 9.3005
R17625 gnd.n3669 gnd.n2299 9.3005
R17626 gnd.n3666 gnd.n2300 9.3005
R17627 gnd.n3665 gnd.n2301 9.3005
R17628 gnd.n3662 gnd.n2302 9.3005
R17629 gnd.n3661 gnd.n2303 9.3005
R17630 gnd.n3658 gnd.n2304 9.3005
R17631 gnd.n3657 gnd.n2305 9.3005
R17632 gnd.n3654 gnd.n2306 9.3005
R17633 gnd.n3653 gnd.n2307 9.3005
R17634 gnd.n3650 gnd.n2308 9.3005
R17635 gnd.n3649 gnd.n2309 9.3005
R17636 gnd.n3646 gnd.n2310 9.3005
R17637 gnd.n3645 gnd.n2311 9.3005
R17638 gnd.n3642 gnd.n2315 9.3005
R17639 gnd.n3641 gnd.n2316 9.3005
R17640 gnd.n3638 gnd.n2317 9.3005
R17641 gnd.n3637 gnd.n2318 9.3005
R17642 gnd.n3688 gnd.n3687 9.3005
R17643 gnd.n3139 gnd.n3123 9.3005
R17644 gnd.n3138 gnd.n3124 9.3005
R17645 gnd.n3137 gnd.n3125 9.3005
R17646 gnd.n3135 gnd.n3126 9.3005
R17647 gnd.n3134 gnd.n3127 9.3005
R17648 gnd.n3132 gnd.n3128 9.3005
R17649 gnd.n3131 gnd.n3129 9.3005
R17650 gnd.n2425 gnd.n2424 9.3005
R17651 gnd.n3208 gnd.n3207 9.3005
R17652 gnd.n3209 gnd.n2423 9.3005
R17653 gnd.n3226 gnd.n3210 9.3005
R17654 gnd.n3225 gnd.n3211 9.3005
R17655 gnd.n3224 gnd.n3212 9.3005
R17656 gnd.n3222 gnd.n3213 9.3005
R17657 gnd.n3221 gnd.n3214 9.3005
R17658 gnd.n3219 gnd.n3215 9.3005
R17659 gnd.n3218 gnd.n3216 9.3005
R17660 gnd.n2369 gnd.n2368 9.3005
R17661 gnd.n3293 gnd.n3292 9.3005
R17662 gnd.n3294 gnd.n2367 9.3005
R17663 gnd.n3315 gnd.n3295 9.3005
R17664 gnd.n3314 gnd.n3296 9.3005
R17665 gnd.n3313 gnd.n3297 9.3005
R17666 gnd.n3310 gnd.n3298 9.3005
R17667 gnd.n3309 gnd.n3299 9.3005
R17668 gnd.n3307 gnd.n3300 9.3005
R17669 gnd.n3306 gnd.n3301 9.3005
R17670 gnd.n3304 gnd.n3303 9.3005
R17671 gnd.n3302 gnd.n2320 9.3005
R17672 gnd.n2880 gnd.n2879 9.3005
R17673 gnd.n2770 gnd.n2769 9.3005
R17674 gnd.n2894 gnd.n2893 9.3005
R17675 gnd.n2895 gnd.n2768 9.3005
R17676 gnd.n2897 gnd.n2896 9.3005
R17677 gnd.n2758 gnd.n2757 9.3005
R17678 gnd.n2910 gnd.n2909 9.3005
R17679 gnd.n2911 gnd.n2756 9.3005
R17680 gnd.n2943 gnd.n2912 9.3005
R17681 gnd.n2942 gnd.n2913 9.3005
R17682 gnd.n2941 gnd.n2914 9.3005
R17683 gnd.n2940 gnd.n2915 9.3005
R17684 gnd.n2937 gnd.n2916 9.3005
R17685 gnd.n2936 gnd.n2917 9.3005
R17686 gnd.n2935 gnd.n2918 9.3005
R17687 gnd.n2933 gnd.n2919 9.3005
R17688 gnd.n2932 gnd.n2920 9.3005
R17689 gnd.n2929 gnd.n2921 9.3005
R17690 gnd.n2928 gnd.n2922 9.3005
R17691 gnd.n2927 gnd.n2923 9.3005
R17692 gnd.n2925 gnd.n2924 9.3005
R17693 gnd.n2624 gnd.n2623 9.3005
R17694 gnd.n3041 gnd.n3040 9.3005
R17695 gnd.n3042 gnd.n2622 9.3005
R17696 gnd.n3046 gnd.n3043 9.3005
R17697 gnd.n3045 gnd.n3044 9.3005
R17698 gnd.n2546 gnd.n2545 9.3005
R17699 gnd.n3121 gnd.n3120 9.3005
R17700 gnd.n2878 gnd.n2779 9.3005
R17701 gnd.n2781 gnd.n2780 9.3005
R17702 gnd.n2825 gnd.n2823 9.3005
R17703 gnd.n2826 gnd.n2822 9.3005
R17704 gnd.n2829 gnd.n2818 9.3005
R17705 gnd.n2830 gnd.n2817 9.3005
R17706 gnd.n2833 gnd.n2816 9.3005
R17707 gnd.n2834 gnd.n2815 9.3005
R17708 gnd.n2837 gnd.n2814 9.3005
R17709 gnd.n2838 gnd.n2813 9.3005
R17710 gnd.n2841 gnd.n2812 9.3005
R17711 gnd.n2842 gnd.n2811 9.3005
R17712 gnd.n2845 gnd.n2810 9.3005
R17713 gnd.n2846 gnd.n2809 9.3005
R17714 gnd.n2849 gnd.n2808 9.3005
R17715 gnd.n2850 gnd.n2807 9.3005
R17716 gnd.n2853 gnd.n2806 9.3005
R17717 gnd.n2854 gnd.n2805 9.3005
R17718 gnd.n2857 gnd.n2804 9.3005
R17719 gnd.n2858 gnd.n2803 9.3005
R17720 gnd.n2861 gnd.n2802 9.3005
R17721 gnd.n2862 gnd.n2801 9.3005
R17722 gnd.n2865 gnd.n2800 9.3005
R17723 gnd.n2867 gnd.n2799 9.3005
R17724 gnd.n2868 gnd.n2798 9.3005
R17725 gnd.n2869 gnd.n2797 9.3005
R17726 gnd.n2870 gnd.n2796 9.3005
R17727 gnd.n2877 gnd.n2876 9.3005
R17728 gnd.n2886 gnd.n2885 9.3005
R17729 gnd.n2887 gnd.n2773 9.3005
R17730 gnd.n2889 gnd.n2888 9.3005
R17731 gnd.n2764 gnd.n2763 9.3005
R17732 gnd.n2902 gnd.n2901 9.3005
R17733 gnd.n2903 gnd.n2762 9.3005
R17734 gnd.n2905 gnd.n2904 9.3005
R17735 gnd.n2751 gnd.n2750 9.3005
R17736 gnd.n2948 gnd.n2947 9.3005
R17737 gnd.n2949 gnd.n2705 9.3005
R17738 gnd.n2953 gnd.n2951 9.3005
R17739 gnd.n2952 gnd.n2684 9.3005
R17740 gnd.n2971 gnd.n2683 9.3005
R17741 gnd.n2974 gnd.n2973 9.3005
R17742 gnd.n2677 gnd.n2676 9.3005
R17743 gnd.n2985 gnd.n2983 9.3005
R17744 gnd.n2984 gnd.n2658 9.3005
R17745 gnd.n3002 gnd.n2657 9.3005
R17746 gnd.n3005 gnd.n3004 9.3005
R17747 gnd.n2652 gnd.n2647 9.3005
R17748 gnd.n3015 gnd.n3014 9.3005
R17749 gnd.n2650 gnd.n2630 9.3005
R17750 gnd.n3036 gnd.n2631 9.3005
R17751 gnd.n3035 gnd.n3034 9.3005
R17752 gnd.n2633 gnd.n2609 9.3005
R17753 gnd.n3067 gnd.n3066 9.3005
R17754 gnd.n3069 gnd.n2554 9.3005
R17755 gnd.n3116 gnd.n2555 9.3005
R17756 gnd.n3115 gnd.n2556 9.3005
R17757 gnd.n3114 gnd.n2557 9.3005
R17758 gnd.n3080 gnd.n2558 9.3005
R17759 gnd.n3082 gnd.n2576 9.3005
R17760 gnd.n3102 gnd.n2577 9.3005
R17761 gnd.n3101 gnd.n2578 9.3005
R17762 gnd.n3100 gnd.n2579 9.3005
R17763 gnd.n3091 gnd.n2580 9.3005
R17764 gnd.n3092 gnd.n2463 9.3005
R17765 gnd.n3158 gnd.n3157 9.3005
R17766 gnd.n3159 gnd.n2456 9.3005
R17767 gnd.n3169 gnd.n3168 9.3005
R17768 gnd.n3171 gnd.n2452 9.3005
R17769 gnd.n3181 gnd.n2453 9.3005
R17770 gnd.n3180 gnd.n3179 9.3005
R17771 gnd.n3177 gnd.n2431 9.3005
R17772 gnd.n3203 gnd.n2432 9.3005
R17773 gnd.n3202 gnd.n3201 9.3005
R17774 gnd.n2434 gnd.n2408 9.3005
R17775 gnd.n3243 gnd.n3242 9.3005
R17776 gnd.n3244 gnd.n2401 9.3005
R17777 gnd.n3254 gnd.n3253 9.3005
R17778 gnd.n3256 gnd.n2397 9.3005
R17779 gnd.n3266 gnd.n2398 9.3005
R17780 gnd.n3265 gnd.n3264 9.3005
R17781 gnd.n3262 gnd.n2376 9.3005
R17782 gnd.n3288 gnd.n2377 9.3005
R17783 gnd.n3287 gnd.n3286 9.3005
R17784 gnd.n2379 gnd.n2354 9.3005
R17785 gnd.n3332 gnd.n3331 9.3005
R17786 gnd.n3333 gnd.n2347 9.3005
R17787 gnd.n3343 gnd.n3342 9.3005
R17788 gnd.n3601 gnd.n2343 9.3005
R17789 gnd.n3609 gnd.n2344 9.3005
R17790 gnd.n3608 gnd.n3607 9.3005
R17791 gnd.n2325 gnd.n2324 9.3005
R17792 gnd.n3632 gnd.n3631 9.3005
R17793 gnd.n2775 gnd.n2774 9.3005
R17794 gnd.n3878 gnd.n3847 9.3005
R17795 gnd.n3877 gnd.n3848 9.3005
R17796 gnd.n3875 gnd.n3849 9.3005
R17797 gnd.n3874 gnd.n3850 9.3005
R17798 gnd.n3872 gnd.n3851 9.3005
R17799 gnd.n3871 gnd.n3852 9.3005
R17800 gnd.n3869 gnd.n3853 9.3005
R17801 gnd.n3868 gnd.n3854 9.3005
R17802 gnd.n3866 gnd.n3855 9.3005
R17803 gnd.n3865 gnd.n3856 9.3005
R17804 gnd.n3863 gnd.n3857 9.3005
R17805 gnd.n3862 gnd.n3858 9.3005
R17806 gnd.n3860 gnd.n3859 9.3005
R17807 gnd.n2171 gnd.n2170 9.3005
R17808 gnd.n4129 gnd.n4128 9.3005
R17809 gnd.n4130 gnd.n2169 9.3005
R17810 gnd.n4134 gnd.n4131 9.3005
R17811 gnd.n4133 gnd.n4132 9.3005
R17812 gnd.n2146 gnd.n2145 9.3005
R17813 gnd.n4164 gnd.n4163 9.3005
R17814 gnd.n4165 gnd.n2144 9.3005
R17815 gnd.n4169 gnd.n4166 9.3005
R17816 gnd.n4168 gnd.n4167 9.3005
R17817 gnd.n2121 gnd.n2120 9.3005
R17818 gnd.n4199 gnd.n4198 9.3005
R17819 gnd.n4200 gnd.n2118 9.3005
R17820 gnd.n3881 gnd.n3880 9.3005
R17821 gnd.n5902 gnd.n1044 9.3005
R17822 gnd.n5905 gnd.n1043 9.3005
R17823 gnd.n5906 gnd.n1042 9.3005
R17824 gnd.n5909 gnd.n1041 9.3005
R17825 gnd.n5910 gnd.n1040 9.3005
R17826 gnd.n5913 gnd.n1039 9.3005
R17827 gnd.n5914 gnd.n1038 9.3005
R17828 gnd.n5917 gnd.n1037 9.3005
R17829 gnd.n5919 gnd.n1034 9.3005
R17830 gnd.n5922 gnd.n1033 9.3005
R17831 gnd.n5923 gnd.n1032 9.3005
R17832 gnd.n5926 gnd.n1031 9.3005
R17833 gnd.n5927 gnd.n1030 9.3005
R17834 gnd.n5930 gnd.n1029 9.3005
R17835 gnd.n5931 gnd.n1028 9.3005
R17836 gnd.n5934 gnd.n1027 9.3005
R17837 gnd.n5935 gnd.n1026 9.3005
R17838 gnd.n5938 gnd.n1025 9.3005
R17839 gnd.n5939 gnd.n1024 9.3005
R17840 gnd.n5942 gnd.n1023 9.3005
R17841 gnd.n5943 gnd.n1022 9.3005
R17842 gnd.n5946 gnd.n1021 9.3005
R17843 gnd.n5947 gnd.n1020 9.3005
R17844 gnd.n5948 gnd.n1019 9.3005
R17845 gnd.n976 gnd.n975 9.3005
R17846 gnd.n5954 gnd.n5953 9.3005
R17847 gnd.n1979 gnd.n1976 9.3005
R17848 gnd.n1983 gnd.n1982 9.3005
R17849 gnd.n1984 gnd.n1974 9.3005
R17850 gnd.n1986 gnd.n1985 9.3005
R17851 gnd.n1989 gnd.n1973 9.3005
R17852 gnd.n1993 gnd.n1992 9.3005
R17853 gnd.n1994 gnd.n1972 9.3005
R17854 gnd.n1997 gnd.n1995 9.3005
R17855 gnd.n1998 gnd.n1968 9.3005
R17856 gnd.n2002 gnd.n2001 9.3005
R17857 gnd.n2003 gnd.n1967 9.3005
R17858 gnd.n2005 gnd.n2004 9.3005
R17859 gnd.n2008 gnd.n1966 9.3005
R17860 gnd.n2012 gnd.n2011 9.3005
R17861 gnd.n2013 gnd.n1965 9.3005
R17862 gnd.n2015 gnd.n2014 9.3005
R17863 gnd.n2018 gnd.n1964 9.3005
R17864 gnd.n2022 gnd.n2021 9.3005
R17865 gnd.n2023 gnd.n1963 9.3005
R17866 gnd.n2025 gnd.n2024 9.3005
R17867 gnd.n2028 gnd.n1962 9.3005
R17868 gnd.n2032 gnd.n2031 9.3005
R17869 gnd.n2033 gnd.n1961 9.3005
R17870 gnd.n2035 gnd.n2034 9.3005
R17871 gnd.n2038 gnd.n1960 9.3005
R17872 gnd.n2042 gnd.n2041 9.3005
R17873 gnd.n2043 gnd.n1959 9.3005
R17874 gnd.n2046 gnd.n2044 9.3005
R17875 gnd.n2047 gnd.n1955 9.3005
R17876 gnd.n2050 gnd.n2049 9.3005
R17877 gnd.n1975 gnd.n1045 9.3005
R17878 gnd.n4259 gnd.n4258 9.3005
R17879 gnd.n4260 gnd.n2082 9.3005
R17880 gnd.n4263 gnd.n4262 9.3005
R17881 gnd.n4261 gnd.n890 9.3005
R17882 gnd.n6005 gnd.n891 9.3005
R17883 gnd.n6004 gnd.n892 9.3005
R17884 gnd.n6003 gnd.n893 9.3005
R17885 gnd.n912 gnd.n894 9.3005
R17886 gnd.n5993 gnd.n913 9.3005
R17887 gnd.n5992 gnd.n914 9.3005
R17888 gnd.n5991 gnd.n915 9.3005
R17889 gnd.n932 gnd.n916 9.3005
R17890 gnd.n5981 gnd.n933 9.3005
R17891 gnd.n5980 gnd.n934 9.3005
R17892 gnd.n5979 gnd.n935 9.3005
R17893 gnd.n952 gnd.n936 9.3005
R17894 gnd.n5969 gnd.n953 9.3005
R17895 gnd.n5968 gnd.n954 9.3005
R17896 gnd.n5967 gnd.n955 9.3005
R17897 gnd.n973 gnd.n956 9.3005
R17898 gnd.n5957 gnd.n974 9.3005
R17899 gnd.n5956 gnd.n5955 9.3005
R17900 gnd.n2130 gnd.n2129 9.3005
R17901 gnd.n4189 gnd.n4188 9.3005
R17902 gnd.n4190 gnd.n2128 9.3005
R17903 gnd.n4194 gnd.n4191 9.3005
R17904 gnd.n4193 gnd.n4192 9.3005
R17905 gnd.n2105 gnd.n2104 9.3005
R17906 gnd.n4232 gnd.n4231 9.3005
R17907 gnd.n4233 gnd.n2103 9.3005
R17908 gnd.n4235 gnd.n4234 9.3005
R17909 gnd.n2084 gnd.n2083 9.3005
R17910 gnd.n4055 gnd.n4054 9.3005
R17911 gnd.n4056 gnd.n2233 9.3005
R17912 gnd.n4058 gnd.n4057 9.3005
R17913 gnd.n2216 gnd.n2215 9.3005
R17914 gnd.n4075 gnd.n4074 9.3005
R17915 gnd.n4076 gnd.n2214 9.3005
R17916 gnd.n4078 gnd.n4077 9.3005
R17917 gnd.n2199 gnd.n2198 9.3005
R17918 gnd.n4095 gnd.n4094 9.3005
R17919 gnd.n4096 gnd.n2197 9.3005
R17920 gnd.n4098 gnd.n4097 9.3005
R17921 gnd.n2179 gnd.n2178 9.3005
R17922 gnd.n4119 gnd.n4118 9.3005
R17923 gnd.n4120 gnd.n2177 9.3005
R17924 gnd.n4124 gnd.n4121 9.3005
R17925 gnd.n4123 gnd.n4122 9.3005
R17926 gnd.n2154 gnd.n2153 9.3005
R17927 gnd.n4154 gnd.n4153 9.3005
R17928 gnd.n4155 gnd.n2152 9.3005
R17929 gnd.n4159 gnd.n4156 9.3005
R17930 gnd.n4158 gnd.n4157 9.3005
R17931 gnd.n2235 gnd.n2234 9.3005
R17932 gnd.n3924 gnd.n3923 9.3005
R17933 gnd.n3926 gnd.n3825 9.3005
R17934 gnd.n3927 gnd.n3824 9.3005
R17935 gnd.n3930 gnd.n3823 9.3005
R17936 gnd.n3931 gnd.n3822 9.3005
R17937 gnd.n3934 gnd.n3821 9.3005
R17938 gnd.n3935 gnd.n3820 9.3005
R17939 gnd.n3938 gnd.n3819 9.3005
R17940 gnd.n3939 gnd.n3818 9.3005
R17941 gnd.n3942 gnd.n3817 9.3005
R17942 gnd.n3943 gnd.n3816 9.3005
R17943 gnd.n3946 gnd.n3815 9.3005
R17944 gnd.n3947 gnd.n3814 9.3005
R17945 gnd.n3950 gnd.n3813 9.3005
R17946 gnd.n3951 gnd.n3812 9.3005
R17947 gnd.n3954 gnd.n3811 9.3005
R17948 gnd.n3955 gnd.n3810 9.3005
R17949 gnd.n3958 gnd.n3809 9.3005
R17950 gnd.n3959 gnd.n3808 9.3005
R17951 gnd.n3962 gnd.n3807 9.3005
R17952 gnd.n3966 gnd.n3803 9.3005
R17953 gnd.n3967 gnd.n3802 9.3005
R17954 gnd.n3970 gnd.n3801 9.3005
R17955 gnd.n3971 gnd.n3800 9.3005
R17956 gnd.n3974 gnd.n3799 9.3005
R17957 gnd.n3975 gnd.n3798 9.3005
R17958 gnd.n3978 gnd.n3797 9.3005
R17959 gnd.n3979 gnd.n3796 9.3005
R17960 gnd.n3982 gnd.n3795 9.3005
R17961 gnd.n3983 gnd.n3794 9.3005
R17962 gnd.n3986 gnd.n3793 9.3005
R17963 gnd.n3987 gnd.n3792 9.3005
R17964 gnd.n3990 gnd.n3791 9.3005
R17965 gnd.n3991 gnd.n3790 9.3005
R17966 gnd.n3994 gnd.n3789 9.3005
R17967 gnd.n3995 gnd.n3788 9.3005
R17968 gnd.n3998 gnd.n3787 9.3005
R17969 gnd.n3999 gnd.n3786 9.3005
R17970 gnd.n4002 gnd.n3785 9.3005
R17971 gnd.n4004 gnd.n3782 9.3005
R17972 gnd.n4007 gnd.n3781 9.3005
R17973 gnd.n4008 gnd.n3780 9.3005
R17974 gnd.n4011 gnd.n3779 9.3005
R17975 gnd.n4012 gnd.n3778 9.3005
R17976 gnd.n4015 gnd.n3777 9.3005
R17977 gnd.n4016 gnd.n3776 9.3005
R17978 gnd.n4019 gnd.n3775 9.3005
R17979 gnd.n4020 gnd.n3774 9.3005
R17980 gnd.n4023 gnd.n3773 9.3005
R17981 gnd.n4024 gnd.n3772 9.3005
R17982 gnd.n4027 gnd.n3771 9.3005
R17983 gnd.n4028 gnd.n3770 9.3005
R17984 gnd.n4031 gnd.n3769 9.3005
R17985 gnd.n4033 gnd.n3768 9.3005
R17986 gnd.n4034 gnd.n3767 9.3005
R17987 gnd.n4035 gnd.n3766 9.3005
R17988 gnd.n4036 gnd.n3765 9.3005
R17989 gnd.n3963 gnd.n3804 9.3005
R17990 gnd.n3922 gnd.n2245 9.3005
R17991 gnd.n3886 gnd.n3885 9.3005
R17992 gnd.n3889 gnd.n3842 9.3005
R17993 gnd.n3890 gnd.n3841 9.3005
R17994 gnd.n3893 gnd.n3840 9.3005
R17995 gnd.n3894 gnd.n3839 9.3005
R17996 gnd.n3897 gnd.n3838 9.3005
R17997 gnd.n3898 gnd.n3837 9.3005
R17998 gnd.n3901 gnd.n3836 9.3005
R17999 gnd.n3902 gnd.n3835 9.3005
R18000 gnd.n3905 gnd.n3834 9.3005
R18001 gnd.n3906 gnd.n3833 9.3005
R18002 gnd.n3909 gnd.n3832 9.3005
R18003 gnd.n3910 gnd.n3831 9.3005
R18004 gnd.n3913 gnd.n3830 9.3005
R18005 gnd.n3914 gnd.n3829 9.3005
R18006 gnd.n3917 gnd.n3828 9.3005
R18007 gnd.n3920 gnd.n3919 9.3005
R18008 gnd.n3884 gnd.n3846 9.3005
R18009 gnd.n3883 gnd.n3882 9.3005
R18010 gnd.n4044 gnd.n2243 9.3005
R18011 gnd.n4046 gnd.n4045 9.3005
R18012 gnd.n4047 gnd.n2226 9.3005
R18013 gnd.n4063 gnd.n2227 9.3005
R18014 gnd.n4064 gnd.n2225 9.3005
R18015 gnd.n4066 gnd.n4065 9.3005
R18016 gnd.n4067 gnd.n2208 9.3005
R18017 gnd.n4083 gnd.n2209 9.3005
R18018 gnd.n4084 gnd.n2207 9.3005
R18019 gnd.n4086 gnd.n4085 9.3005
R18020 gnd.n4087 gnd.n2190 9.3005
R18021 gnd.n4103 gnd.n2191 9.3005
R18022 gnd.n4104 gnd.n2188 9.3005
R18023 gnd.n4106 gnd.n2189 9.3005
R18024 gnd.n4108 gnd.n4107 9.3005
R18025 gnd.n4109 gnd.n2164 9.3005
R18026 gnd.n4138 gnd.n2165 9.3005
R18027 gnd.n4139 gnd.n2162 9.3005
R18028 gnd.n4141 gnd.n2163 9.3005
R18029 gnd.n4143 gnd.n4142 9.3005
R18030 gnd.n4144 gnd.n2139 9.3005
R18031 gnd.n4173 gnd.n2140 9.3005
R18032 gnd.n4174 gnd.n2137 9.3005
R18033 gnd.n4176 gnd.n2138 9.3005
R18034 gnd.n4178 gnd.n4177 9.3005
R18035 gnd.n4179 gnd.n2113 9.3005
R18036 gnd.n4220 gnd.n2114 9.3005
R18037 gnd.n4221 gnd.n2112 9.3005
R18038 gnd.n4223 gnd.n4222 9.3005
R18039 gnd.n4224 gnd.n2096 9.3005
R18040 gnd.n4240 gnd.n2097 9.3005
R18041 gnd.n4241 gnd.n2093 9.3005
R18042 gnd.n4243 gnd.n2094 9.3005
R18043 gnd.n4244 gnd.n2095 9.3005
R18044 gnd.n4247 gnd.n4246 9.3005
R18045 gnd.n4248 gnd.n2073 9.3005
R18046 gnd.n4276 gnd.n2074 9.3005
R18047 gnd.n4277 gnd.n902 9.3005
R18048 gnd.n4278 gnd.n903 9.3005
R18049 gnd.n4279 gnd.n904 9.3005
R18050 gnd.n4281 gnd.n4280 9.3005
R18051 gnd.n2061 gnd.n923 9.3005
R18052 gnd.n4342 gnd.n924 9.3005
R18053 gnd.n4343 gnd.n925 9.3005
R18054 gnd.n4345 gnd.n4344 9.3005
R18055 gnd.n2056 gnd.n942 9.3005
R18056 gnd.n4357 gnd.n943 9.3005
R18057 gnd.n4358 gnd.n944 9.3005
R18058 gnd.n4360 gnd.n4359 9.3005
R18059 gnd.n2051 gnd.n963 9.3005
R18060 gnd.n4374 gnd.n964 9.3005
R18061 gnd.n4375 gnd.n965 9.3005
R18062 gnd.n4377 gnd.n4376 9.3005
R18063 gnd.n4043 gnd.n2244 9.3005
R18064 gnd.n4050 gnd.n2243 9.3005
R18065 gnd.n4049 gnd.n4046 9.3005
R18066 gnd.n4048 gnd.n4047 9.3005
R18067 gnd.n2227 gnd.n2224 9.3005
R18068 gnd.n4070 gnd.n2225 9.3005
R18069 gnd.n4069 gnd.n4066 9.3005
R18070 gnd.n4068 gnd.n4067 9.3005
R18071 gnd.n2209 gnd.n2206 9.3005
R18072 gnd.n4090 gnd.n2207 9.3005
R18073 gnd.n4089 gnd.n4086 9.3005
R18074 gnd.n4088 gnd.n4087 9.3005
R18075 gnd.n2191 gnd.n2187 9.3005
R18076 gnd.n4114 gnd.n2188 9.3005
R18077 gnd.n4113 gnd.n2189 9.3005
R18078 gnd.n4112 gnd.n4108 9.3005
R18079 gnd.n4111 gnd.n4109 9.3005
R18080 gnd.n2165 gnd.n2161 9.3005
R18081 gnd.n4149 gnd.n2162 9.3005
R18082 gnd.n4148 gnd.n2163 9.3005
R18083 gnd.n4147 gnd.n4143 9.3005
R18084 gnd.n4146 gnd.n4144 9.3005
R18085 gnd.n2140 gnd.n2136 9.3005
R18086 gnd.n4184 gnd.n2137 9.3005
R18087 gnd.n4183 gnd.n2138 9.3005
R18088 gnd.n4182 gnd.n4178 9.3005
R18089 gnd.n4181 gnd.n4179 9.3005
R18090 gnd.n2114 gnd.n2111 9.3005
R18091 gnd.n4227 gnd.n2112 9.3005
R18092 gnd.n4226 gnd.n4223 9.3005
R18093 gnd.n4225 gnd.n4224 9.3005
R18094 gnd.n2097 gnd.n2092 9.3005
R18095 gnd.n4254 gnd.n2093 9.3005
R18096 gnd.n4253 gnd.n2094 9.3005
R18097 gnd.n4252 gnd.n2095 9.3005
R18098 gnd.n4251 gnd.n4247 9.3005
R18099 gnd.n4249 gnd.n4248 9.3005
R18100 gnd.n2074 gnd.n901 9.3005
R18101 gnd.n5999 gnd.n902 9.3005
R18102 gnd.n5998 gnd.n903 9.3005
R18103 gnd.n5997 gnd.n904 9.3005
R18104 gnd.n4280 gnd.n905 9.3005
R18105 gnd.n5987 gnd.n923 9.3005
R18106 gnd.n5986 gnd.n924 9.3005
R18107 gnd.n5985 gnd.n925 9.3005
R18108 gnd.n4344 gnd.n926 9.3005
R18109 gnd.n5975 gnd.n942 9.3005
R18110 gnd.n5974 gnd.n943 9.3005
R18111 gnd.n5973 gnd.n944 9.3005
R18112 gnd.n4359 gnd.n945 9.3005
R18113 gnd.n5963 gnd.n963 9.3005
R18114 gnd.n5962 gnd.n964 9.3005
R18115 gnd.n5961 gnd.n965 9.3005
R18116 gnd.n4377 gnd.n966 9.3005
R18117 gnd.n2244 gnd.n2242 9.3005
R18118 gnd.n6180 gnd.n713 9.3005
R18119 gnd.n6182 gnd.n6181 9.3005
R18120 gnd.n709 gnd.n708 9.3005
R18121 gnd.n6189 gnd.n6188 9.3005
R18122 gnd.n6190 gnd.n707 9.3005
R18123 gnd.n6192 gnd.n6191 9.3005
R18124 gnd.n703 gnd.n702 9.3005
R18125 gnd.n6199 gnd.n6198 9.3005
R18126 gnd.n6200 gnd.n701 9.3005
R18127 gnd.n6202 gnd.n6201 9.3005
R18128 gnd.n697 gnd.n696 9.3005
R18129 gnd.n6209 gnd.n6208 9.3005
R18130 gnd.n6210 gnd.n695 9.3005
R18131 gnd.n6212 gnd.n6211 9.3005
R18132 gnd.n691 gnd.n690 9.3005
R18133 gnd.n6219 gnd.n6218 9.3005
R18134 gnd.n6220 gnd.n689 9.3005
R18135 gnd.n6222 gnd.n6221 9.3005
R18136 gnd.n685 gnd.n684 9.3005
R18137 gnd.n6229 gnd.n6228 9.3005
R18138 gnd.n6230 gnd.n683 9.3005
R18139 gnd.n6232 gnd.n6231 9.3005
R18140 gnd.n679 gnd.n678 9.3005
R18141 gnd.n6239 gnd.n6238 9.3005
R18142 gnd.n6240 gnd.n677 9.3005
R18143 gnd.n6242 gnd.n6241 9.3005
R18144 gnd.n673 gnd.n672 9.3005
R18145 gnd.n6249 gnd.n6248 9.3005
R18146 gnd.n6250 gnd.n671 9.3005
R18147 gnd.n6252 gnd.n6251 9.3005
R18148 gnd.n667 gnd.n666 9.3005
R18149 gnd.n6259 gnd.n6258 9.3005
R18150 gnd.n6260 gnd.n665 9.3005
R18151 gnd.n6262 gnd.n6261 9.3005
R18152 gnd.n661 gnd.n660 9.3005
R18153 gnd.n6269 gnd.n6268 9.3005
R18154 gnd.n6270 gnd.n659 9.3005
R18155 gnd.n6272 gnd.n6271 9.3005
R18156 gnd.n655 gnd.n654 9.3005
R18157 gnd.n6279 gnd.n6278 9.3005
R18158 gnd.n6280 gnd.n653 9.3005
R18159 gnd.n6282 gnd.n6281 9.3005
R18160 gnd.n649 gnd.n648 9.3005
R18161 gnd.n6289 gnd.n6288 9.3005
R18162 gnd.n6290 gnd.n647 9.3005
R18163 gnd.n6292 gnd.n6291 9.3005
R18164 gnd.n643 gnd.n642 9.3005
R18165 gnd.n6299 gnd.n6298 9.3005
R18166 gnd.n6300 gnd.n641 9.3005
R18167 gnd.n6302 gnd.n6301 9.3005
R18168 gnd.n637 gnd.n636 9.3005
R18169 gnd.n6309 gnd.n6308 9.3005
R18170 gnd.n6310 gnd.n635 9.3005
R18171 gnd.n6312 gnd.n6311 9.3005
R18172 gnd.n631 gnd.n630 9.3005
R18173 gnd.n6319 gnd.n6318 9.3005
R18174 gnd.n6320 gnd.n629 9.3005
R18175 gnd.n6322 gnd.n6321 9.3005
R18176 gnd.n625 gnd.n624 9.3005
R18177 gnd.n6329 gnd.n6328 9.3005
R18178 gnd.n6330 gnd.n623 9.3005
R18179 gnd.n6332 gnd.n6331 9.3005
R18180 gnd.n619 gnd.n618 9.3005
R18181 gnd.n6339 gnd.n6338 9.3005
R18182 gnd.n6340 gnd.n617 9.3005
R18183 gnd.n6342 gnd.n6341 9.3005
R18184 gnd.n613 gnd.n612 9.3005
R18185 gnd.n6349 gnd.n6348 9.3005
R18186 gnd.n6350 gnd.n611 9.3005
R18187 gnd.n6352 gnd.n6351 9.3005
R18188 gnd.n607 gnd.n606 9.3005
R18189 gnd.n6359 gnd.n6358 9.3005
R18190 gnd.n6360 gnd.n605 9.3005
R18191 gnd.n6362 gnd.n6361 9.3005
R18192 gnd.n601 gnd.n600 9.3005
R18193 gnd.n6369 gnd.n6368 9.3005
R18194 gnd.n6370 gnd.n599 9.3005
R18195 gnd.n6372 gnd.n6371 9.3005
R18196 gnd.n595 gnd.n594 9.3005
R18197 gnd.n6379 gnd.n6378 9.3005
R18198 gnd.n6380 gnd.n593 9.3005
R18199 gnd.n6382 gnd.n6381 9.3005
R18200 gnd.n589 gnd.n588 9.3005
R18201 gnd.n6389 gnd.n6388 9.3005
R18202 gnd.n6390 gnd.n587 9.3005
R18203 gnd.n6392 gnd.n6391 9.3005
R18204 gnd.n583 gnd.n582 9.3005
R18205 gnd.n6399 gnd.n6398 9.3005
R18206 gnd.n6400 gnd.n581 9.3005
R18207 gnd.n6402 gnd.n6401 9.3005
R18208 gnd.n577 gnd.n576 9.3005
R18209 gnd.n6409 gnd.n6408 9.3005
R18210 gnd.n6410 gnd.n575 9.3005
R18211 gnd.n6412 gnd.n6411 9.3005
R18212 gnd.n571 gnd.n570 9.3005
R18213 gnd.n6419 gnd.n6418 9.3005
R18214 gnd.n6420 gnd.n569 9.3005
R18215 gnd.n6422 gnd.n6421 9.3005
R18216 gnd.n565 gnd.n564 9.3005
R18217 gnd.n6429 gnd.n6428 9.3005
R18218 gnd.n6430 gnd.n563 9.3005
R18219 gnd.n6432 gnd.n6431 9.3005
R18220 gnd.n559 gnd.n558 9.3005
R18221 gnd.n6439 gnd.n6438 9.3005
R18222 gnd.n6440 gnd.n557 9.3005
R18223 gnd.n6442 gnd.n6441 9.3005
R18224 gnd.n553 gnd.n552 9.3005
R18225 gnd.n6449 gnd.n6448 9.3005
R18226 gnd.n6450 gnd.n551 9.3005
R18227 gnd.n6452 gnd.n6451 9.3005
R18228 gnd.n547 gnd.n546 9.3005
R18229 gnd.n6459 gnd.n6458 9.3005
R18230 gnd.n6460 gnd.n545 9.3005
R18231 gnd.n6462 gnd.n6461 9.3005
R18232 gnd.n541 gnd.n540 9.3005
R18233 gnd.n6469 gnd.n6468 9.3005
R18234 gnd.n6470 gnd.n539 9.3005
R18235 gnd.n6472 gnd.n6471 9.3005
R18236 gnd.n535 gnd.n534 9.3005
R18237 gnd.n6479 gnd.n6478 9.3005
R18238 gnd.n6480 gnd.n533 9.3005
R18239 gnd.n6482 gnd.n6481 9.3005
R18240 gnd.n529 gnd.n528 9.3005
R18241 gnd.n6489 gnd.n6488 9.3005
R18242 gnd.n6490 gnd.n527 9.3005
R18243 gnd.n6493 gnd.n6492 9.3005
R18244 gnd.n6491 gnd.n523 9.3005
R18245 gnd.n6499 gnd.n522 9.3005
R18246 gnd.n6501 gnd.n6500 9.3005
R18247 gnd.n518 gnd.n517 9.3005
R18248 gnd.n6510 gnd.n6509 9.3005
R18249 gnd.n6511 gnd.n516 9.3005
R18250 gnd.n6513 gnd.n6512 9.3005
R18251 gnd.n512 gnd.n511 9.3005
R18252 gnd.n6520 gnd.n6519 9.3005
R18253 gnd.n6521 gnd.n510 9.3005
R18254 gnd.n6523 gnd.n6522 9.3005
R18255 gnd.n506 gnd.n505 9.3005
R18256 gnd.n6530 gnd.n6529 9.3005
R18257 gnd.n6531 gnd.n504 9.3005
R18258 gnd.n6533 gnd.n6532 9.3005
R18259 gnd.n500 gnd.n499 9.3005
R18260 gnd.n6540 gnd.n6539 9.3005
R18261 gnd.n6541 gnd.n498 9.3005
R18262 gnd.n6543 gnd.n6542 9.3005
R18263 gnd.n494 gnd.n493 9.3005
R18264 gnd.n6550 gnd.n6549 9.3005
R18265 gnd.n6551 gnd.n492 9.3005
R18266 gnd.n6553 gnd.n6552 9.3005
R18267 gnd.n488 gnd.n487 9.3005
R18268 gnd.n6560 gnd.n6559 9.3005
R18269 gnd.n6561 gnd.n486 9.3005
R18270 gnd.n6563 gnd.n6562 9.3005
R18271 gnd.n482 gnd.n481 9.3005
R18272 gnd.n6570 gnd.n6569 9.3005
R18273 gnd.n6571 gnd.n480 9.3005
R18274 gnd.n6573 gnd.n6572 9.3005
R18275 gnd.n476 gnd.n475 9.3005
R18276 gnd.n6580 gnd.n6579 9.3005
R18277 gnd.n6581 gnd.n474 9.3005
R18278 gnd.n6583 gnd.n6582 9.3005
R18279 gnd.n470 gnd.n469 9.3005
R18280 gnd.n6590 gnd.n6589 9.3005
R18281 gnd.n6591 gnd.n468 9.3005
R18282 gnd.n6593 gnd.n6592 9.3005
R18283 gnd.n464 gnd.n463 9.3005
R18284 gnd.n6600 gnd.n6599 9.3005
R18285 gnd.n6601 gnd.n462 9.3005
R18286 gnd.n6603 gnd.n6602 9.3005
R18287 gnd.n458 gnd.n457 9.3005
R18288 gnd.n6610 gnd.n6609 9.3005
R18289 gnd.n6611 gnd.n456 9.3005
R18290 gnd.n6613 gnd.n6612 9.3005
R18291 gnd.n452 gnd.n451 9.3005
R18292 gnd.n6620 gnd.n6619 9.3005
R18293 gnd.n6621 gnd.n450 9.3005
R18294 gnd.n6623 gnd.n6622 9.3005
R18295 gnd.n446 gnd.n445 9.3005
R18296 gnd.n6630 gnd.n6629 9.3005
R18297 gnd.n6631 gnd.n444 9.3005
R18298 gnd.n6633 gnd.n6632 9.3005
R18299 gnd.n440 gnd.n439 9.3005
R18300 gnd.n6640 gnd.n6639 9.3005
R18301 gnd.n6641 gnd.n438 9.3005
R18302 gnd.n6643 gnd.n6642 9.3005
R18303 gnd.n434 gnd.n433 9.3005
R18304 gnd.n6650 gnd.n6649 9.3005
R18305 gnd.n6651 gnd.n432 9.3005
R18306 gnd.n6653 gnd.n6652 9.3005
R18307 gnd.n428 gnd.n427 9.3005
R18308 gnd.n6660 gnd.n6659 9.3005
R18309 gnd.n6661 gnd.n426 9.3005
R18310 gnd.n6663 gnd.n6662 9.3005
R18311 gnd.n422 gnd.n421 9.3005
R18312 gnd.n6670 gnd.n6669 9.3005
R18313 gnd.n6671 gnd.n420 9.3005
R18314 gnd.n6673 gnd.n6672 9.3005
R18315 gnd.n416 gnd.n415 9.3005
R18316 gnd.n6680 gnd.n6679 9.3005
R18317 gnd.n6681 gnd.n414 9.3005
R18318 gnd.n6683 gnd.n6682 9.3005
R18319 gnd.n410 gnd.n409 9.3005
R18320 gnd.n6690 gnd.n6689 9.3005
R18321 gnd.n6691 gnd.n408 9.3005
R18322 gnd.n6693 gnd.n6692 9.3005
R18323 gnd.n404 gnd.n403 9.3005
R18324 gnd.n6700 gnd.n6699 9.3005
R18325 gnd.n6701 gnd.n402 9.3005
R18326 gnd.n6703 gnd.n6702 9.3005
R18327 gnd.n398 gnd.n397 9.3005
R18328 gnd.n6711 gnd.n6710 9.3005
R18329 gnd.n6712 gnd.n396 9.3005
R18330 gnd.n6714 gnd.n6713 9.3005
R18331 gnd.n6503 gnd.n6502 9.3005
R18332 gnd.n4302 gnd.n4301 9.3005
R18333 gnd.n4303 gnd.n4297 9.3005
R18334 gnd.n4305 gnd.n4304 9.3005
R18335 gnd.n2067 gnd.n2066 9.3005
R18336 gnd.n4310 gnd.n4309 9.3005
R18337 gnd.n4311 gnd.n2065 9.3005
R18338 gnd.n4337 gnd.n4312 9.3005
R18339 gnd.n4336 gnd.n4313 9.3005
R18340 gnd.n4335 gnd.n4314 9.3005
R18341 gnd.n4317 gnd.n4315 9.3005
R18342 gnd.n4331 gnd.n4318 9.3005
R18343 gnd.n4330 gnd.n4319 9.3005
R18344 gnd.n4329 gnd.n4320 9.3005
R18345 gnd.n4322 gnd.n4321 9.3005
R18346 gnd.n4325 gnd.n4324 9.3005
R18347 gnd.n4323 gnd.n1855 9.3005
R18348 gnd.n4465 gnd.n1856 9.3005
R18349 gnd.n4464 gnd.n1857 9.3005
R18350 gnd.n4463 gnd.n1858 9.3005
R18351 gnd.n1860 gnd.n1859 9.3005
R18352 gnd.n1862 gnd.n1861 9.3005
R18353 gnd.n1838 gnd.n1837 9.3005
R18354 gnd.n4483 gnd.n4482 9.3005
R18355 gnd.n4484 gnd.n1836 9.3005
R18356 gnd.n4486 gnd.n4485 9.3005
R18357 gnd.n1825 gnd.n1824 9.3005
R18358 gnd.n4499 gnd.n4498 9.3005
R18359 gnd.n4500 gnd.n1823 9.3005
R18360 gnd.n4502 gnd.n4501 9.3005
R18361 gnd.n1809 gnd.n1808 9.3005
R18362 gnd.n4533 gnd.n4532 9.3005
R18363 gnd.n4534 gnd.n1807 9.3005
R18364 gnd.n4545 gnd.n4535 9.3005
R18365 gnd.n4544 gnd.n4536 9.3005
R18366 gnd.n4543 gnd.n4537 9.3005
R18367 gnd.n4540 gnd.n4539 9.3005
R18368 gnd.n4538 gnd.n1118 9.3005
R18369 gnd.n5823 gnd.n1119 9.3005
R18370 gnd.n5822 gnd.n1120 9.3005
R18371 gnd.n5821 gnd.n1121 9.3005
R18372 gnd.n1712 gnd.n1122 9.3005
R18373 gnd.n4653 gnd.n4652 9.3005
R18374 gnd.n4654 gnd.n1711 9.3005
R18375 gnd.n4661 gnd.n4655 9.3005
R18376 gnd.n4660 gnd.n4656 9.3005
R18377 gnd.n4659 gnd.n4657 9.3005
R18378 gnd.n1688 gnd.n1687 9.3005
R18379 gnd.n4693 gnd.n4692 9.3005
R18380 gnd.n4694 gnd.n1686 9.3005
R18381 gnd.n4698 gnd.n4695 9.3005
R18382 gnd.n4697 gnd.n4696 9.3005
R18383 gnd.n1660 gnd.n1659 9.3005
R18384 gnd.n4729 gnd.n4728 9.3005
R18385 gnd.n4730 gnd.n1658 9.3005
R18386 gnd.n4732 gnd.n4731 9.3005
R18387 gnd.n1642 gnd.n1641 9.3005
R18388 gnd.n4755 gnd.n4754 9.3005
R18389 gnd.n4756 gnd.n1640 9.3005
R18390 gnd.n4760 gnd.n4757 9.3005
R18391 gnd.n4759 gnd.n4758 9.3005
R18392 gnd.n1616 gnd.n1615 9.3005
R18393 gnd.n4811 gnd.n4810 9.3005
R18394 gnd.n4812 gnd.n1614 9.3005
R18395 gnd.n4816 gnd.n4813 9.3005
R18396 gnd.n4815 gnd.n4814 9.3005
R18397 gnd.n1591 gnd.n1590 9.3005
R18398 gnd.n4851 gnd.n4850 9.3005
R18399 gnd.n4852 gnd.n1589 9.3005
R18400 gnd.n4856 gnd.n4853 9.3005
R18401 gnd.n4855 gnd.n4854 9.3005
R18402 gnd.n1561 gnd.n1560 9.3005
R18403 gnd.n4920 gnd.n4919 9.3005
R18404 gnd.n4921 gnd.n1559 9.3005
R18405 gnd.n4925 gnd.n4922 9.3005
R18406 gnd.n4924 gnd.n4923 9.3005
R18407 gnd.n1537 gnd.n1536 9.3005
R18408 gnd.n4953 gnd.n4952 9.3005
R18409 gnd.n4954 gnd.n1535 9.3005
R18410 gnd.n4958 gnd.n4955 9.3005
R18411 gnd.n4957 gnd.n4956 9.3005
R18412 gnd.n1516 gnd.n1515 9.3005
R18413 gnd.n5007 gnd.n5006 9.3005
R18414 gnd.n5008 gnd.n1514 9.3005
R18415 gnd.n5012 gnd.n5009 9.3005
R18416 gnd.n5011 gnd.n5010 9.3005
R18417 gnd.n1491 gnd.n1490 9.3005
R18418 gnd.n5044 gnd.n5043 9.3005
R18419 gnd.n5045 gnd.n1489 9.3005
R18420 gnd.n5047 gnd.n5046 9.3005
R18421 gnd.n1400 gnd.n1399 9.3005
R18422 gnd.n5187 gnd.n5186 9.3005
R18423 gnd.n5188 gnd.n1398 9.3005
R18424 gnd.n5190 gnd.n5189 9.3005
R18425 gnd.n1387 gnd.n1386 9.3005
R18426 gnd.n5203 gnd.n5202 9.3005
R18427 gnd.n5204 gnd.n1385 9.3005
R18428 gnd.n5206 gnd.n5205 9.3005
R18429 gnd.n1374 gnd.n1373 9.3005
R18430 gnd.n5219 gnd.n5218 9.3005
R18431 gnd.n5220 gnd.n1372 9.3005
R18432 gnd.n5222 gnd.n5221 9.3005
R18433 gnd.n1361 gnd.n1360 9.3005
R18434 gnd.n5235 gnd.n5234 9.3005
R18435 gnd.n5236 gnd.n1359 9.3005
R18436 gnd.n5239 gnd.n5238 9.3005
R18437 gnd.n5237 gnd.n1234 9.3005
R18438 gnd.n5713 gnd.n1235 9.3005
R18439 gnd.n5712 gnd.n1236 9.3005
R18440 gnd.n5711 gnd.n1237 9.3005
R18441 gnd.n5278 gnd.n1238 9.3005
R18442 gnd.n5279 gnd.n5277 9.3005
R18443 gnd.n5472 gnd.n5280 9.3005
R18444 gnd.n5471 gnd.n5281 9.3005
R18445 gnd.n5470 gnd.n5282 9.3005
R18446 gnd.n5389 gnd.n5283 9.3005
R18447 gnd.n5392 gnd.n5391 9.3005
R18448 gnd.n5393 gnd.n5388 9.3005
R18449 gnd.n5397 gnd.n5394 9.3005
R18450 gnd.n5396 gnd.n5395 9.3005
R18451 gnd.n5341 gnd.n5340 9.3005
R18452 gnd.n5430 gnd.n5429 9.3005
R18453 gnd.n5431 gnd.n5339 9.3005
R18454 gnd.n5436 gnd.n5432 9.3005
R18455 gnd.n5435 gnd.n5434 9.3005
R18456 gnd.n5433 gnd.n391 9.3005
R18457 gnd.n6719 gnd.n392 9.3005
R18458 gnd.n6718 gnd.n393 9.3005
R18459 gnd.n6717 gnd.n394 9.3005
R18460 gnd.n4299 gnd.n4298 9.3005
R18461 gnd.n6011 gnd.n880 9.3005
R18462 gnd.n6012 gnd.n879 9.3005
R18463 gnd.n878 gnd.n874 9.3005
R18464 gnd.n6018 gnd.n873 9.3005
R18465 gnd.n6019 gnd.n872 9.3005
R18466 gnd.n6020 gnd.n871 9.3005
R18467 gnd.n870 gnd.n866 9.3005
R18468 gnd.n6026 gnd.n865 9.3005
R18469 gnd.n6027 gnd.n864 9.3005
R18470 gnd.n6028 gnd.n863 9.3005
R18471 gnd.n862 gnd.n858 9.3005
R18472 gnd.n6034 gnd.n857 9.3005
R18473 gnd.n6035 gnd.n856 9.3005
R18474 gnd.n6036 gnd.n855 9.3005
R18475 gnd.n854 gnd.n850 9.3005
R18476 gnd.n6042 gnd.n849 9.3005
R18477 gnd.n6043 gnd.n848 9.3005
R18478 gnd.n6044 gnd.n847 9.3005
R18479 gnd.n846 gnd.n842 9.3005
R18480 gnd.n6050 gnd.n841 9.3005
R18481 gnd.n6051 gnd.n840 9.3005
R18482 gnd.n6052 gnd.n839 9.3005
R18483 gnd.n838 gnd.n834 9.3005
R18484 gnd.n6058 gnd.n833 9.3005
R18485 gnd.n6059 gnd.n832 9.3005
R18486 gnd.n6060 gnd.n831 9.3005
R18487 gnd.n830 gnd.n826 9.3005
R18488 gnd.n6066 gnd.n825 9.3005
R18489 gnd.n6067 gnd.n824 9.3005
R18490 gnd.n6068 gnd.n823 9.3005
R18491 gnd.n822 gnd.n818 9.3005
R18492 gnd.n6074 gnd.n817 9.3005
R18493 gnd.n6075 gnd.n816 9.3005
R18494 gnd.n6076 gnd.n815 9.3005
R18495 gnd.n814 gnd.n810 9.3005
R18496 gnd.n6082 gnd.n809 9.3005
R18497 gnd.n6083 gnd.n808 9.3005
R18498 gnd.n6084 gnd.n807 9.3005
R18499 gnd.n806 gnd.n802 9.3005
R18500 gnd.n6090 gnd.n801 9.3005
R18501 gnd.n6091 gnd.n800 9.3005
R18502 gnd.n6092 gnd.n799 9.3005
R18503 gnd.n798 gnd.n794 9.3005
R18504 gnd.n6098 gnd.n793 9.3005
R18505 gnd.n6099 gnd.n792 9.3005
R18506 gnd.n6100 gnd.n791 9.3005
R18507 gnd.n790 gnd.n786 9.3005
R18508 gnd.n6106 gnd.n785 9.3005
R18509 gnd.n6107 gnd.n784 9.3005
R18510 gnd.n6108 gnd.n783 9.3005
R18511 gnd.n782 gnd.n778 9.3005
R18512 gnd.n6114 gnd.n777 9.3005
R18513 gnd.n6115 gnd.n776 9.3005
R18514 gnd.n6116 gnd.n775 9.3005
R18515 gnd.n774 gnd.n770 9.3005
R18516 gnd.n6122 gnd.n769 9.3005
R18517 gnd.n6123 gnd.n768 9.3005
R18518 gnd.n6124 gnd.n767 9.3005
R18519 gnd.n766 gnd.n762 9.3005
R18520 gnd.n6130 gnd.n761 9.3005
R18521 gnd.n6131 gnd.n760 9.3005
R18522 gnd.n6132 gnd.n759 9.3005
R18523 gnd.n758 gnd.n754 9.3005
R18524 gnd.n6138 gnd.n753 9.3005
R18525 gnd.n6139 gnd.n752 9.3005
R18526 gnd.n6140 gnd.n751 9.3005
R18527 gnd.n750 gnd.n746 9.3005
R18528 gnd.n6146 gnd.n745 9.3005
R18529 gnd.n6147 gnd.n744 9.3005
R18530 gnd.n6148 gnd.n743 9.3005
R18531 gnd.n742 gnd.n738 9.3005
R18532 gnd.n6154 gnd.n737 9.3005
R18533 gnd.n6155 gnd.n736 9.3005
R18534 gnd.n6156 gnd.n735 9.3005
R18535 gnd.n734 gnd.n730 9.3005
R18536 gnd.n6162 gnd.n729 9.3005
R18537 gnd.n6163 gnd.n728 9.3005
R18538 gnd.n6164 gnd.n727 9.3005
R18539 gnd.n726 gnd.n722 9.3005
R18540 gnd.n6170 gnd.n721 9.3005
R18541 gnd.n6171 gnd.n720 9.3005
R18542 gnd.n6172 gnd.n719 9.3005
R18543 gnd.n715 gnd.n714 9.3005
R18544 gnd.n6179 gnd.n6178 9.3005
R18545 gnd.n6010 gnd.n881 9.3005
R18546 gnd.n5718 gnd.n5717 9.3005
R18547 gnd.n1832 gnd.n1831 9.3005
R18548 gnd.n4491 gnd.n4490 9.3005
R18549 gnd.n4492 gnd.n1830 9.3005
R18550 gnd.n4494 gnd.n4493 9.3005
R18551 gnd.n1818 gnd.n1817 9.3005
R18552 gnd.n4507 gnd.n4506 9.3005
R18553 gnd.n4508 gnd.n1815 9.3005
R18554 gnd.n4528 gnd.n4527 9.3005
R18555 gnd.n4526 gnd.n1816 9.3005
R18556 gnd.n4525 gnd.n4524 9.3005
R18557 gnd.n4523 gnd.n4509 9.3005
R18558 gnd.n4522 gnd.n4521 9.3005
R18559 gnd.n4520 gnd.n4513 9.3005
R18560 gnd.n4519 gnd.n4518 9.3005
R18561 gnd.n4517 gnd.n4514 9.3005
R18562 gnd.n1131 gnd.n1129 9.3005
R18563 gnd.n5817 gnd.n5816 9.3005
R18564 gnd.n5815 gnd.n1130 9.3005
R18565 gnd.n5814 gnd.n5813 9.3005
R18566 gnd.n5812 gnd.n1132 9.3005
R18567 gnd.n5811 gnd.n5810 9.3005
R18568 gnd.n5809 gnd.n1136 9.3005
R18569 gnd.n5808 gnd.n5807 9.3005
R18570 gnd.n5806 gnd.n1137 9.3005
R18571 gnd.n5805 gnd.n5804 9.3005
R18572 gnd.n5803 gnd.n1141 9.3005
R18573 gnd.n5802 gnd.n5801 9.3005
R18574 gnd.n5800 gnd.n1142 9.3005
R18575 gnd.n5799 gnd.n5798 9.3005
R18576 gnd.n5797 gnd.n1146 9.3005
R18577 gnd.n5796 gnd.n5795 9.3005
R18578 gnd.n5794 gnd.n1147 9.3005
R18579 gnd.n5793 gnd.n5792 9.3005
R18580 gnd.n5791 gnd.n1151 9.3005
R18581 gnd.n5790 gnd.n5789 9.3005
R18582 gnd.n5788 gnd.n1152 9.3005
R18583 gnd.n5787 gnd.n5786 9.3005
R18584 gnd.n5785 gnd.n1156 9.3005
R18585 gnd.n5784 gnd.n5783 9.3005
R18586 gnd.n5782 gnd.n1157 9.3005
R18587 gnd.n5781 gnd.n5780 9.3005
R18588 gnd.n5779 gnd.n1161 9.3005
R18589 gnd.n5778 gnd.n5777 9.3005
R18590 gnd.n5776 gnd.n1162 9.3005
R18591 gnd.n5775 gnd.n5774 9.3005
R18592 gnd.n5773 gnd.n1166 9.3005
R18593 gnd.n5772 gnd.n5771 9.3005
R18594 gnd.n5770 gnd.n1167 9.3005
R18595 gnd.n5769 gnd.n5768 9.3005
R18596 gnd.n5767 gnd.n1171 9.3005
R18597 gnd.n5766 gnd.n5765 9.3005
R18598 gnd.n5764 gnd.n1172 9.3005
R18599 gnd.n5763 gnd.n5762 9.3005
R18600 gnd.n5761 gnd.n1176 9.3005
R18601 gnd.n5760 gnd.n5759 9.3005
R18602 gnd.n5758 gnd.n1177 9.3005
R18603 gnd.n5757 gnd.n5756 9.3005
R18604 gnd.n5755 gnd.n1181 9.3005
R18605 gnd.n5754 gnd.n5753 9.3005
R18606 gnd.n5752 gnd.n1182 9.3005
R18607 gnd.n5751 gnd.n5750 9.3005
R18608 gnd.n5749 gnd.n1186 9.3005
R18609 gnd.n5748 gnd.n5747 9.3005
R18610 gnd.n5746 gnd.n1187 9.3005
R18611 gnd.n5745 gnd.n5744 9.3005
R18612 gnd.n5743 gnd.n1191 9.3005
R18613 gnd.n5742 gnd.n5741 9.3005
R18614 gnd.n5740 gnd.n1192 9.3005
R18615 gnd.n5739 gnd.n5738 9.3005
R18616 gnd.n5737 gnd.n1196 9.3005
R18617 gnd.n5736 gnd.n5735 9.3005
R18618 gnd.n5734 gnd.n1197 9.3005
R18619 gnd.n5733 gnd.n5732 9.3005
R18620 gnd.n5731 gnd.n1201 9.3005
R18621 gnd.n5730 gnd.n5729 9.3005
R18622 gnd.n5728 gnd.n1202 9.3005
R18623 gnd.n5727 gnd.n5726 9.3005
R18624 gnd.n5725 gnd.n1206 9.3005
R18625 gnd.n5724 gnd.n5723 9.3005
R18626 gnd.n5722 gnd.n1207 9.3005
R18627 gnd.n5721 gnd.n5720 9.3005
R18628 gnd.n5719 gnd.n1211 9.3005
R18629 gnd.n4478 gnd.n4477 9.3005
R18630 gnd.n4476 gnd.n4475 9.3005
R18631 gnd.n4216 gnd.n4215 9.3005
R18632 gnd.n4214 gnd.n2119 9.3005
R18633 gnd.n4213 gnd.n4212 9.3005
R18634 gnd.n4211 gnd.n4202 9.3005
R18635 gnd.n4210 gnd.n4209 9.3005
R18636 gnd.n4208 gnd.n4205 9.3005
R18637 gnd.n4207 gnd.n4206 9.3005
R18638 gnd.n2077 gnd.n2076 9.3005
R18639 gnd.n4269 gnd.n4268 9.3005
R18640 gnd.n4270 gnd.n2075 9.3005
R18641 gnd.n4272 gnd.n4271 9.3005
R18642 gnd.n2071 gnd.n2069 9.3005
R18643 gnd.n4292 gnd.n4291 9.3005
R18644 gnd.n4290 gnd.n2070 9.3005
R18645 gnd.n4289 gnd.n4288 9.3005
R18646 gnd.n4287 gnd.n2072 9.3005
R18647 gnd.n4286 gnd.n4285 9.3005
R18648 gnd.n2060 gnd.n2059 9.3005
R18649 gnd.n4350 gnd.n4349 9.3005
R18650 gnd.n4351 gnd.n2058 9.3005
R18651 gnd.n4353 gnd.n4352 9.3005
R18652 gnd.n2055 gnd.n2054 9.3005
R18653 gnd.n4365 gnd.n4364 9.3005
R18654 gnd.n4366 gnd.n2052 9.3005
R18655 gnd.n4370 gnd.n4369 9.3005
R18656 gnd.n4368 gnd.n2053 9.3005
R18657 gnd.n4367 gnd.n1851 9.3005
R18658 gnd.n4391 gnd.n4390 9.3005
R18659 gnd.n1908 gnd.n1905 9.3005
R18660 gnd.n4399 gnd.n4398 9.3005
R18661 gnd.n4403 gnd.n4402 9.3005
R18662 gnd.n1902 gnd.n1901 9.3005
R18663 gnd.n4411 gnd.n4410 9.3005
R18664 gnd.n4415 gnd.n4414 9.3005
R18665 gnd.n1896 gnd.n1893 9.3005
R18666 gnd.n4423 gnd.n4422 9.3005
R18667 gnd.n4427 gnd.n4426 9.3005
R18668 gnd.n1890 gnd.n1889 9.3005
R18669 gnd.n4435 gnd.n4434 9.3005
R18670 gnd.n4439 gnd.n4438 9.3005
R18671 gnd.n1884 gnd.n1881 9.3005
R18672 gnd.n4448 gnd.n4447 9.3005
R18673 gnd.n4452 gnd.n4451 9.3005
R18674 gnd.n4453 gnd.n1850 9.3005
R18675 gnd.n4472 gnd.n4471 9.3005
R18676 gnd.n4388 gnd.n4387 9.3005
R18677 gnd.n4474 gnd.n4473 9.3005
R18678 gnd.n1847 gnd.n1845 9.3005
R18679 gnd.n4455 gnd.n4454 9.3005
R18680 gnd.n4444 gnd.n1880 9.3005
R18681 gnd.n4446 gnd.n4445 9.3005
R18682 gnd.n4441 gnd.n4440 9.3005
R18683 gnd.n1888 gnd.n1885 9.3005
R18684 gnd.n4433 gnd.n4432 9.3005
R18685 gnd.n4429 gnd.n4428 9.3005
R18686 gnd.n1892 gnd.n1891 9.3005
R18687 gnd.n4421 gnd.n4420 9.3005
R18688 gnd.n4417 gnd.n4416 9.3005
R18689 gnd.n1900 gnd.n1897 9.3005
R18690 gnd.n4409 gnd.n4408 9.3005
R18691 gnd.n4405 gnd.n4404 9.3005
R18692 gnd.n1904 gnd.n1903 9.3005
R18693 gnd.n4397 gnd.n4396 9.3005
R18694 gnd.n4393 gnd.n4392 9.3005
R18695 gnd.n1912 gnd.n1909 9.3005
R18696 gnd.n4386 gnd.n4385 9.3005
R18697 gnd.n4382 gnd.n1913 9.3005
R18698 gnd.n4381 gnd.n4380 9.3005
R18699 gnd.n1954 gnd.n1914 9.3005
R18700 gnd.n1953 gnd.n1952 9.3005
R18701 gnd.n1949 gnd.n1917 9.3005
R18702 gnd.n1948 gnd.n1947 9.3005
R18703 gnd.n1946 gnd.n1918 9.3005
R18704 gnd.n1945 gnd.n1944 9.3005
R18705 gnd.n1940 gnd.n1921 9.3005
R18706 gnd.n1939 gnd.n1938 9.3005
R18707 gnd.n1937 gnd.n1924 9.3005
R18708 gnd.n1936 gnd.n1935 9.3005
R18709 gnd.n1934 gnd.n1925 9.3005
R18710 gnd.n1933 gnd.n1932 9.3005
R18711 gnd.n1931 gnd.n1928 9.3005
R18712 gnd.n1930 gnd.n1929 9.3005
R18713 gnd.n1801 gnd.n1800 9.3005
R18714 gnd.n4550 gnd.n4549 9.3005
R18715 gnd.n4551 gnd.n1799 9.3005
R18716 gnd.n4553 gnd.n4552 9.3005
R18717 gnd.n1797 gnd.n1796 9.3005
R18718 gnd.n4558 gnd.n4557 9.3005
R18719 gnd.n4559 gnd.n1794 9.3005
R18720 gnd.n4619 gnd.n4618 9.3005
R18721 gnd.n4617 gnd.n1795 9.3005
R18722 gnd.n4616 gnd.n4615 9.3005
R18723 gnd.n4614 gnd.n4560 9.3005
R18724 gnd.n4613 gnd.n4612 9.3005
R18725 gnd.n4611 gnd.n4565 9.3005
R18726 gnd.n4610 gnd.n4609 9.3005
R18727 gnd.n4608 gnd.n4566 9.3005
R18728 gnd.n4607 gnd.n4606 9.3005
R18729 gnd.n4605 gnd.n4569 9.3005
R18730 gnd.n4604 gnd.n4603 9.3005
R18731 gnd.n4602 gnd.n4570 9.3005
R18732 gnd.n4601 gnd.n4600 9.3005
R18733 gnd.n4599 gnd.n4574 9.3005
R18734 gnd.n4598 gnd.n4597 9.3005
R18735 gnd.n4596 gnd.n4575 9.3005
R18736 gnd.n4595 gnd.n4594 9.3005
R18737 gnd.n4593 gnd.n4578 9.3005
R18738 gnd.n4592 gnd.n4591 9.3005
R18739 gnd.n4590 gnd.n4579 9.3005
R18740 gnd.n4589 gnd.n4588 9.3005
R18741 gnd.n4587 gnd.n4582 9.3005
R18742 gnd.n4586 gnd.n4585 9.3005
R18743 gnd.n4584 gnd.n4583 9.3005
R18744 gnd.n1606 gnd.n1605 9.3005
R18745 gnd.n4821 gnd.n4820 9.3005
R18746 gnd.n4822 gnd.n1603 9.3005
R18747 gnd.n4838 gnd.n4837 9.3005
R18748 gnd.n4836 gnd.n1604 9.3005
R18749 gnd.n4835 gnd.n4834 9.3005
R18750 gnd.n4833 gnd.n4823 9.3005
R18751 gnd.n4832 gnd.n4831 9.3005
R18752 gnd.n4830 gnd.n4827 9.3005
R18753 gnd.n4829 gnd.n4828 9.3005
R18754 gnd.n1553 gnd.n1552 9.3005
R18755 gnd.n4930 gnd.n4929 9.3005
R18756 gnd.n4931 gnd.n1550 9.3005
R18757 gnd.n4934 gnd.n4933 9.3005
R18758 gnd.n4932 gnd.n1551 9.3005
R18759 gnd.n1530 gnd.n1529 9.3005
R18760 gnd.n4963 gnd.n4962 9.3005
R18761 gnd.n4964 gnd.n1527 9.3005
R18762 gnd.n4993 gnd.n4992 9.3005
R18763 gnd.n4991 gnd.n1528 9.3005
R18764 gnd.n4990 gnd.n4989 9.3005
R18765 gnd.n4988 gnd.n4965 9.3005
R18766 gnd.n4987 gnd.n4986 9.3005
R18767 gnd.n4985 gnd.n4972 9.3005
R18768 gnd.n4984 gnd.n4983 9.3005
R18769 gnd.n4982 gnd.n4973 9.3005
R18770 gnd.n4981 gnd.n4980 9.3005
R18771 gnd.n4979 gnd.n4976 9.3005
R18772 gnd.n4978 gnd.n4977 9.3005
R18773 gnd.n1392 gnd.n1391 9.3005
R18774 gnd.n5195 gnd.n5194 9.3005
R18775 gnd.n5196 gnd.n1390 9.3005
R18776 gnd.n5198 gnd.n5197 9.3005
R18777 gnd.n1379 gnd.n1378 9.3005
R18778 gnd.n5211 gnd.n5210 9.3005
R18779 gnd.n5212 gnd.n1377 9.3005
R18780 gnd.n5214 gnd.n5213 9.3005
R18781 gnd.n1367 gnd.n1366 9.3005
R18782 gnd.n5227 gnd.n5226 9.3005
R18783 gnd.n5228 gnd.n1365 9.3005
R18784 gnd.n5230 gnd.n5229 9.3005
R18785 gnd.n1354 gnd.n1353 9.3005
R18786 gnd.n5244 gnd.n5243 9.3005
R18787 gnd.n1942 gnd.n1941 9.3005
R18788 gnd.n5247 gnd.n5246 9.3005
R18789 gnd.n5250 gnd.n1351 9.3005
R18790 gnd.n5254 gnd.n5253 9.3005
R18791 gnd.n5255 gnd.n1350 9.3005
R18792 gnd.n5257 gnd.n5256 9.3005
R18793 gnd.n5260 gnd.n1348 9.3005
R18794 gnd.n5245 gnd.n1352 9.3005
R18795 gnd.n5545 gnd.n5544 9.3005
R18796 gnd.n5522 gnd.n5521 9.3005
R18797 gnd.n5551 gnd.n5550 9.3005
R18798 gnd.n5553 gnd.n5552 9.3005
R18799 gnd.n5512 gnd.n5511 9.3005
R18800 gnd.n5559 gnd.n5558 9.3005
R18801 gnd.n5561 gnd.n5560 9.3005
R18802 gnd.n5502 gnd.n5501 9.3005
R18803 gnd.n5567 gnd.n5566 9.3005
R18804 gnd.n5569 gnd.n5568 9.3005
R18805 gnd.n5492 gnd.n5491 9.3005
R18806 gnd.n5575 gnd.n5574 9.3005
R18807 gnd.n5577 gnd.n5576 9.3005
R18808 gnd.n5482 gnd.n5481 9.3005
R18809 gnd.n5583 gnd.n5582 9.3005
R18810 gnd.n5585 gnd.n5584 9.3005
R18811 gnd.n5478 gnd.n5266 9.3005
R18812 gnd.n5543 gnd.n5539 9.3005
R18813 gnd.n5533 gnd.n5531 9.3005
R18814 gnd.n5590 gnd.n5589 9.3005
R18815 gnd.n5588 gnd.n1349 9.3005
R18816 gnd.n5587 gnd.n5586 9.3005
R18817 gnd.n5267 gnd.n5265 9.3005
R18818 gnd.n5581 gnd.n5580 9.3005
R18819 gnd.n5579 gnd.n5578 9.3005
R18820 gnd.n5486 gnd.n5485 9.3005
R18821 gnd.n5573 gnd.n5572 9.3005
R18822 gnd.n5571 gnd.n5570 9.3005
R18823 gnd.n5498 gnd.n5497 9.3005
R18824 gnd.n5565 gnd.n5564 9.3005
R18825 gnd.n5563 gnd.n5562 9.3005
R18826 gnd.n5506 gnd.n5505 9.3005
R18827 gnd.n5557 gnd.n5556 9.3005
R18828 gnd.n5555 gnd.n5554 9.3005
R18829 gnd.n5518 gnd.n5517 9.3005
R18830 gnd.n5549 gnd.n5548 9.3005
R18831 gnd.n5547 gnd.n5546 9.3005
R18832 gnd.n5534 gnd.n5528 9.3005
R18833 gnd.n5538 gnd.n5537 9.3005
R18834 gnd.n5532 gnd.n1213 9.3005
R18835 gnd.n5371 gnd.n5368 9.3005
R18836 gnd.n5375 gnd.n5374 9.3005
R18837 gnd.n5376 gnd.n5367 9.3005
R18838 gnd.n5378 gnd.n5377 9.3005
R18839 gnd.n5352 gnd.n5351 9.3005
R18840 gnd.n5403 gnd.n5402 9.3005
R18841 gnd.n5404 gnd.n5350 9.3005
R18842 gnd.n5406 gnd.n5405 9.3005
R18843 gnd.n5346 gnd.n5344 9.3005
R18844 gnd.n5424 gnd.n5423 9.3005
R18845 gnd.n5422 gnd.n5345 9.3005
R18846 gnd.n5421 gnd.n5420 9.3005
R18847 gnd.n5419 gnd.n5347 9.3005
R18848 gnd.n368 gnd.n367 9.3005
R18849 gnd.n6748 gnd.n6747 9.3005
R18850 gnd.n6749 gnd.n365 9.3005
R18851 gnd.n6752 gnd.n6751 9.3005
R18852 gnd.n6750 gnd.n366 9.3005
R18853 gnd.n341 gnd.n340 9.3005
R18854 gnd.n6782 gnd.n6781 9.3005
R18855 gnd.n6783 gnd.n338 9.3005
R18856 gnd.n6791 gnd.n6790 9.3005
R18857 gnd.n6789 gnd.n339 9.3005
R18858 gnd.n6788 gnd.n6787 9.3005
R18859 gnd.n6786 gnd.n6784 9.3005
R18860 gnd.n81 gnd.n79 9.3005
R18861 gnd.n5370 gnd.n5369 9.3005
R18862 gnd.t341 gnd.n2438 9.24152
R18863 gnd.n2340 gnd.t204 9.24152
R18864 gnd.n3624 gnd.t301 9.24152
R18865 gnd.t222 gnd.n2229 9.24152
R18866 gnd.n4372 gnd.t240 9.24152
R18867 gnd.n5286 gnd.t218 9.24152
R18868 gnd.t226 gnd.n195 9.24152
R18869 gnd.t358 gnd.t341 8.92286
R18870 gnd.t267 gnd.n1480 8.92286
R18871 gnd.n3594 gnd.n3569 8.92171
R18872 gnd.n3562 gnd.n3537 8.92171
R18873 gnd.n3530 gnd.n3505 8.92171
R18874 gnd.n3499 gnd.n3474 8.92171
R18875 gnd.n3467 gnd.n3442 8.92171
R18876 gnd.n3435 gnd.n3410 8.92171
R18877 gnd.n3403 gnd.n3378 8.92171
R18878 gnd.n3372 gnd.n3347 8.92171
R18879 gnd.n1427 gnd.n1409 8.72777
R18880 gnd.n3098 gnd.t343 8.60421
R18881 gnd.n2510 gnd.n2494 8.43656
R18882 gnd.n46 gnd.n30 8.43656
R18883 gnd.n4563 gnd.t305 8.28555
R18884 gnd.n4683 gnd.t174 8.28555
R18885 gnd.n4706 gnd.n1676 8.28555
R18886 gnd.n1631 gnd.n1626 8.28555
R18887 gnd.n1596 gnd.n1583 8.28555
R18888 gnd.n4950 gnd.n4948 8.28555
R18889 gnd.t194 gnd.n1518 8.28555
R18890 gnd.n3595 gnd.n3567 8.14595
R18891 gnd.n3563 gnd.n3535 8.14595
R18892 gnd.n3531 gnd.n3503 8.14595
R18893 gnd.n3500 gnd.n3472 8.14595
R18894 gnd.n3468 gnd.n3440 8.14595
R18895 gnd.n3436 gnd.n3408 8.14595
R18896 gnd.n3404 gnd.n3376 8.14595
R18897 gnd.n3373 gnd.n3345 8.14595
R18898 gnd.n4201 gnd.n0 8.10675
R18899 gnd.n7197 gnd.n7196 8.10675
R18900 gnd.n3600 gnd.n3599 7.97301
R18901 gnd.t344 gnd.n2613 7.9669
R18902 gnd.n7197 gnd.n78 7.86902
R18903 gnd.n5543 gnd.n5531 7.75808
R18904 gnd.n6950 gnd.n6897 7.75808
R18905 gnd.n4471 gnd.n1850 7.75808
R18906 gnd.n3882 gnd.n3846 7.75808
R18907 gnd.n4628 gnd.t230 7.64824
R18908 gnd.n2543 gnd.n2542 7.53171
R18909 gnd.n3007 gnd.t333 7.32958
R18910 gnd.n1106 gnd.n1105 7.30353
R18911 gnd.n1426 gnd.n1425 7.30353
R18912 gnd.n2967 gnd.n2686 7.01093
R18913 gnd.n2689 gnd.n2687 7.01093
R18914 gnd.n2977 gnd.n2976 7.01093
R18915 gnd.n2988 gnd.n2670 7.01093
R18916 gnd.n2987 gnd.n2673 7.01093
R18917 gnd.n2998 gnd.n2661 7.01093
R18918 gnd.n2664 gnd.n2662 7.01093
R18919 gnd.n3008 gnd.n3007 7.01093
R18920 gnd.n3018 gnd.n2642 7.01093
R18921 gnd.n3017 gnd.n2645 7.01093
R18922 gnd.n3026 gnd.n2636 7.01093
R18923 gnd.n3038 gnd.n2626 7.01093
R18924 gnd.n3048 gnd.n2611 7.01093
R18925 gnd.n3064 gnd.n3063 7.01093
R18926 gnd.n2613 gnd.n2550 7.01093
R18927 gnd.n3118 gnd.n2551 7.01093
R18928 gnd.n3112 gnd.n3111 7.01093
R18929 gnd.n2600 gnd.n2562 7.01093
R18930 gnd.n3104 gnd.n2573 7.01093
R18931 gnd.n2591 gnd.n2586 7.01093
R18932 gnd.n3098 gnd.n3097 7.01093
R18933 gnd.n3144 gnd.n2473 7.01093
R18934 gnd.n3143 gnd.n3142 7.01093
R18935 gnd.n3155 gnd.n3154 7.01093
R18936 gnd.n2466 gnd.n2458 7.01093
R18937 gnd.n3184 gnd.n2446 7.01093
R18938 gnd.n3183 gnd.n2449 7.01093
R18939 gnd.n3194 gnd.n2438 7.01093
R18940 gnd.n2439 gnd.n2427 7.01093
R18941 gnd.n3205 gnd.n2428 7.01093
R18942 gnd.n3229 gnd.n2419 7.01093
R18943 gnd.n3228 gnd.n2410 7.01093
R18944 gnd.n3251 gnd.n3250 7.01093
R18945 gnd.n3269 gnd.n2391 7.01093
R18946 gnd.n3268 gnd.n2394 7.01093
R18947 gnd.n3279 gnd.n2383 7.01093
R18948 gnd.n2384 gnd.n2371 7.01093
R18949 gnd.n3290 gnd.n2372 7.01093
R18950 gnd.n3317 gnd.n2356 7.01093
R18951 gnd.n3329 gnd.n3328 7.01093
R18952 gnd.n3311 gnd.n2349 7.01093
R18953 gnd.n3340 gnd.n3339 7.01093
R18954 gnd.n3612 gnd.n2337 7.01093
R18955 gnd.n3611 gnd.n2340 7.01093
R18956 gnd.n3624 gnd.n2329 7.01093
R18957 gnd.n2330 gnd.n2321 7.01093
R18958 gnd.n3634 gnd.n2322 7.01093
R18959 gnd.n4726 gnd.n1662 7.01093
R18960 gnd.n4764 gnd.n1635 7.01093
R18961 gnd.n4762 gnd.t321 7.01093
R18962 gnd.t181 gnd.n4858 7.01093
R18963 gnd.n4865 gnd.n1579 7.01093
R18964 gnd.n4871 gnd.n4870 7.01093
R18965 gnd.n5041 gnd.n1493 7.01093
R18966 gnd.n1486 gnd.t267 7.01093
R18967 gnd.n2645 gnd.t336 6.69227
R18968 gnd.n2449 gnd.t358 6.69227
R18969 gnd.n3318 gnd.t342 6.69227
R18970 gnd.n4092 gnd.t46 6.69227
R18971 gnd.n5983 gnd.t51 6.69227
R18972 gnd.n2057 gnd.t36 6.69227
R18973 gnd.n4563 gnd.t184 6.69227
R18974 gnd.n4969 gnd.t195 6.69227
R18975 gnd.n5399 gnd.t43 6.69227
R18976 gnd.n5449 gnd.t15 6.69227
R18977 gnd.n7143 gnd.t30 6.69227
R18978 gnd.n5114 gnd.n5113 6.5566
R18979 gnd.n1728 gnd.n1727 6.5566
R18980 gnd.n5838 gnd.n5834 6.5566
R18981 gnd.n5129 gnd.n5128 6.5566
R18982 gnd.n4455 gnd.n1879 6.20656
R18983 gnd.n5534 gnd.n5527 6.20656
R18984 gnd.t186 gnd.n3074 6.05496
R18985 gnd.n3075 gnd.t335 6.05496
R18986 gnd.t346 gnd.n2473 6.05496
R18987 gnd.t330 gnd.n3239 6.05496
R18988 gnd.n4136 gnd.t28 6.05496
R18989 gnd.t41 gnd.n6007 6.05496
R18990 gnd.n4295 gnd.t26 6.05496
R18991 gnd.n6721 gnd.t54 6.05496
R18992 gnd.n6754 gnd.t17 6.05496
R18993 gnd.n7167 gnd.t75 6.05496
R18994 gnd.n3597 gnd.n3567 5.81868
R18995 gnd.n3565 gnd.n3535 5.81868
R18996 gnd.n3533 gnd.n3503 5.81868
R18997 gnd.n3502 gnd.n3472 5.81868
R18998 gnd.n3470 gnd.n3440 5.81868
R18999 gnd.n3438 gnd.n3408 5.81868
R19000 gnd.n3406 gnd.n3376 5.81868
R19001 gnd.n3375 gnd.n3345 5.81868
R19002 gnd.n5826 gnd.n5825 5.73631
R19003 gnd.n4628 gnd.n4621 5.73631
R19004 gnd.n4735 gnd.n4734 5.73631
R19005 gnd.n4742 gnd.n1649 5.73631
R19006 gnd.n4917 gnd.n1563 5.73631
R19007 gnd.n4898 gnd.n1567 5.73631
R19008 gnd.n5050 gnd.n5049 5.73631
R19009 gnd.n5056 gnd.n1480 5.73631
R19010 gnd.n1453 gnd.n1310 5.62001
R19011 gnd.n5900 gnd.n1048 5.62001
R19012 gnd.n5900 gnd.n1049 5.62001
R19013 gnd.n5123 gnd.n1310 5.62001
R19014 gnd.n2826 gnd.n2821 5.4308
R19015 gnd.n3642 gnd.n2314 5.4308
R19016 gnd.n3142 gnd.t345 5.41765
R19017 gnd.t331 gnd.n3165 5.41765
R19018 gnd.t0 gnd.n2403 5.41765
R19019 gnd.n4196 gnd.t92 5.41765
R19020 gnd.n4229 gnd.t48 5.41765
R19021 gnd.n4690 gnd.t177 5.41765
R19022 gnd.n4874 gnd.t197 5.41765
R19023 gnd.n6813 gnd.t19 5.41765
R19024 gnd.n7191 gnd.t57 5.41765
R19025 gnd.n4649 gnd.t305 5.09899
R19026 gnd.n4633 gnd.t329 5.09899
R19027 gnd.t319 gnd.n1669 5.09899
R19028 gnd.n4711 gnd.t322 5.09899
R19029 gnd.t189 gnd.n1555 5.09899
R19030 gnd.n4936 gnd.t173 5.09899
R19031 gnd.n5015 gnd.t188 5.09899
R19032 gnd.t215 gnd.n5183 5.09899
R19033 gnd.n3595 gnd.n3594 5.04292
R19034 gnd.n3563 gnd.n3562 5.04292
R19035 gnd.n3531 gnd.n3530 5.04292
R19036 gnd.n3500 gnd.n3499 5.04292
R19037 gnd.n3468 gnd.n3467 5.04292
R19038 gnd.n3436 gnd.n3435 5.04292
R19039 gnd.n3404 gnd.n3403 5.04292
R19040 gnd.n3373 gnd.n3372 5.04292
R19041 gnd.n3105 gnd.t334 4.78034
R19042 gnd.n2428 gnd.t339 4.78034
R19043 gnd.n4161 gnd.t77 4.78034
R19044 gnd.n2089 gnd.t94 4.78034
R19045 gnd.n6779 gnd.t61 4.78034
R19046 gnd.t21 gnd.n109 4.78034
R19047 gnd.n2547 gnd.n2544 4.74817
R19048 gnd.n2597 gnd.n2479 4.74817
R19049 gnd.n2584 gnd.n2478 4.74817
R19050 gnd.n2477 gnd.n2476 4.74817
R19051 gnd.n2593 gnd.n2544 4.74817
R19052 gnd.n2594 gnd.n2479 4.74817
R19053 gnd.n2596 gnd.n2478 4.74817
R19054 gnd.n2583 gnd.n2477 4.74817
R19055 gnd.n2542 gnd.n2541 4.74296
R19056 gnd.n78 gnd.n77 4.74296
R19057 gnd.n2510 gnd.n2509 4.7074
R19058 gnd.n2526 gnd.n2525 4.7074
R19059 gnd.n46 gnd.n45 4.7074
R19060 gnd.n62 gnd.n61 4.7074
R19061 gnd.n2542 gnd.n2526 4.65959
R19062 gnd.n78 gnd.n62 4.65959
R19063 gnd.n5655 gnd.n1312 4.6132
R19064 gnd.n5901 gnd.n1047 4.6132
R19065 gnd.n5951 gnd.n978 4.46168
R19066 gnd.n5827 gnd.n1110 4.46168
R19067 gnd.n5819 gnd.n1124 4.46168
R19068 gnd.n4643 gnd.t251 4.46168
R19069 gnd.n4711 gnd.n1665 4.46168
R19070 gnd.n4752 gnd.n1644 4.46168
R19071 gnd.n4905 gnd.n1572 4.46168
R19072 gnd.n4927 gnd.n1555 4.46168
R19073 gnd.n5184 gnd.n1402 4.46168
R19074 gnd.n5708 gnd.n1278 4.46168
R19075 gnd.n1422 gnd.n1409 4.46111
R19076 gnd.n3580 gnd.n3576 4.38594
R19077 gnd.n3548 gnd.n3544 4.38594
R19078 gnd.n3516 gnd.n3512 4.38594
R19079 gnd.n3485 gnd.n3481 4.38594
R19080 gnd.n3453 gnd.n3449 4.38594
R19081 gnd.n3421 gnd.n3417 4.38594
R19082 gnd.n3389 gnd.n3385 4.38594
R19083 gnd.n3358 gnd.n3354 4.38594
R19084 gnd.n3591 gnd.n3569 4.26717
R19085 gnd.n3559 gnd.n3537 4.26717
R19086 gnd.n3527 gnd.n3505 4.26717
R19087 gnd.n3496 gnd.n3474 4.26717
R19088 gnd.n3464 gnd.n3442 4.26717
R19089 gnd.n3432 gnd.n3410 4.26717
R19090 gnd.n3400 gnd.n3378 4.26717
R19091 gnd.n3369 gnd.n3347 4.26717
R19092 gnd.n3049 gnd.t340 4.14303
R19093 gnd.n3279 gnd.t337 4.14303
R19094 gnd.t98 gnd.n2181 4.14303
R19095 gnd.n6008 gnd.n883 4.14303
R19096 gnd.n4283 gnd.t68 4.14303
R19097 gnd.n4339 gnd.t51 4.14303
R19098 gnd.n5427 gnd.t15 4.14303
R19099 gnd.n5417 gnd.t32 4.14303
R19100 gnd.n6769 gnd.n351 4.14303
R19101 gnd.t65 gnd.n147 4.14303
R19102 gnd.n3599 gnd.n3598 4.08274
R19103 gnd.n5113 gnd.n5112 4.05904
R19104 gnd.n1729 gnd.n1728 4.05904
R19105 gnd.n5841 gnd.n5834 4.05904
R19106 gnd.n5130 gnd.n5129 4.05904
R19107 gnd.n15 gnd.n7 3.99943
R19108 gnd.n3122 gnd.n2543 3.81325
R19109 gnd.n2526 gnd.n2510 3.72967
R19110 gnd.n62 gnd.n46 3.72967
R19111 gnd.n3599 gnd.n3471 3.70378
R19112 gnd.n15 gnd.n14 3.60163
R19113 gnd.n5897 gnd.n1052 3.50571
R19114 gnd.n5192 gnd.n1394 3.50571
R19115 gnd.n3590 gnd.n3571 3.49141
R19116 gnd.n3558 gnd.n3539 3.49141
R19117 gnd.n3526 gnd.n3507 3.49141
R19118 gnd.n3495 gnd.n3476 3.49141
R19119 gnd.n3463 gnd.n3444 3.49141
R19120 gnd.n3431 gnd.n3412 3.49141
R19121 gnd.n3399 gnd.n3380 3.49141
R19122 gnd.n3368 gnd.n3349 3.49141
R19123 gnd.n7078 gnd.n7075 3.29747
R19124 gnd.n7079 gnd.n7078 3.29747
R19125 gnd.n5673 gnd.n5672 3.29747
R19126 gnd.n5672 gnd.n5671 3.29747
R19127 gnd.n4004 gnd.n4003 3.29747
R19128 gnd.n4003 gnd.n4002 3.29747
R19129 gnd.n5919 gnd.n5918 3.29747
R19130 gnd.n5918 gnd.n5917 3.29747
R19131 gnd.t212 gnd.n1084 3.18706
R19132 gnd.n4650 gnd.n1713 3.18706
R19133 gnd.n4718 gnd.n1669 3.18706
R19134 gnd.t326 gnd.n1644 3.18706
R19135 gnd.n4763 gnd.n4762 3.18706
R19136 gnd.n4858 gnd.n1577 3.18706
R19137 gnd.n4905 gnd.t325 3.18706
R19138 gnd.n4937 gnd.n4936 3.18706
R19139 gnd.n5034 gnd.n1500 3.18706
R19140 gnd.n2628 gnd.t340 2.8684
R19141 gnd.t190 gnd.n1114 2.8684
R19142 gnd.t354 gnd.n1486 2.8684
R19143 gnd.n2527 gnd.t69 2.82907
R19144 gnd.n2527 gnd.t106 2.82907
R19145 gnd.n2529 gnd.t42 2.82907
R19146 gnd.n2529 gnd.t87 2.82907
R19147 gnd.n2531 gnd.t109 2.82907
R19148 gnd.n2531 gnd.t95 2.82907
R19149 gnd.n2533 gnd.t93 2.82907
R19150 gnd.n2533 gnd.t81 2.82907
R19151 gnd.n2535 gnd.t100 2.82907
R19152 gnd.n2535 gnd.t137 2.82907
R19153 gnd.n2537 gnd.t25 2.82907
R19154 gnd.n2537 gnd.t124 2.82907
R19155 gnd.n2539 gnd.t161 2.82907
R19156 gnd.n2539 gnd.t99 2.82907
R19157 gnd.n2480 gnd.t102 2.82907
R19158 gnd.n2480 gnd.t125 2.82907
R19159 gnd.n2482 gnd.t136 2.82907
R19160 gnd.n2482 gnd.t70 2.82907
R19161 gnd.n2484 gnd.t121 2.82907
R19162 gnd.n2484 gnd.t115 2.82907
R19163 gnd.n2486 gnd.t167 2.82907
R19164 gnd.n2486 gnd.t154 2.82907
R19165 gnd.n2488 gnd.t78 2.82907
R19166 gnd.n2488 gnd.t129 2.82907
R19167 gnd.n2490 gnd.t149 2.82907
R19168 gnd.n2490 gnd.t29 2.82907
R19169 gnd.n2492 gnd.t47 2.82907
R19170 gnd.n2492 gnd.t120 2.82907
R19171 gnd.n2495 gnd.t170 2.82907
R19172 gnd.n2495 gnd.t52 2.82907
R19173 gnd.n2497 gnd.t50 2.82907
R19174 gnd.n2497 gnd.t27 2.82907
R19175 gnd.n2499 gnd.t135 2.82907
R19176 gnd.n2499 gnd.t169 2.82907
R19177 gnd.n2501 gnd.t166 2.82907
R19178 gnd.n2501 gnd.t49 2.82907
R19179 gnd.n2503 gnd.t155 2.82907
R19180 gnd.n2503 gnd.t132 2.82907
R19181 gnd.n2505 gnd.t133 2.82907
R19182 gnd.n2505 gnd.t164 2.82907
R19183 gnd.n2507 gnd.t165 2.82907
R19184 gnd.n2507 gnd.t148 2.82907
R19185 gnd.n2511 gnd.t116 2.82907
R19186 gnd.n2511 gnd.t72 2.82907
R19187 gnd.n2513 gnd.t101 2.82907
R19188 gnd.n2513 gnd.t139 2.82907
R19189 gnd.n2515 gnd.t162 2.82907
R19190 gnd.n2515 gnd.t147 2.82907
R19191 gnd.n2517 gnd.t145 2.82907
R19192 gnd.n2517 gnd.t128 2.82907
R19193 gnd.n2519 gnd.t152 2.82907
R19194 gnd.n2519 gnd.t60 2.82907
R19195 gnd.n2521 gnd.t89 2.82907
R19196 gnd.n2521 gnd.t35 2.82907
R19197 gnd.n2523 gnd.t80 2.82907
R19198 gnd.n2523 gnd.t151 2.82907
R19199 gnd.n75 gnd.t66 2.82907
R19200 gnd.n75 gnd.t118 2.82907
R19201 gnd.n73 gnd.t88 2.82907
R19202 gnd.n73 gnd.t130 2.82907
R19203 gnd.n71 gnd.t104 2.82907
R19204 gnd.n71 gnd.t79 2.82907
R19205 gnd.n69 gnd.t34 2.82907
R19206 gnd.n69 gnd.t58 2.82907
R19207 gnd.n67 gnd.t62 2.82907
R19208 gnd.n67 gnd.t84 2.82907
R19209 gnd.n65 gnd.t55 2.82907
R19210 gnd.n65 gnd.t144 2.82907
R19211 gnd.n63 gnd.t114 2.82907
R19212 gnd.n63 gnd.t33 2.82907
R19213 gnd.n28 gnd.t159 2.82907
R19214 gnd.n28 gnd.t82 2.82907
R19215 gnd.n26 gnd.t76 2.82907
R19216 gnd.n26 gnd.t39 2.82907
R19217 gnd.n24 gnd.t172 2.82907
R19218 gnd.n24 gnd.t67 2.82907
R19219 gnd.n22 gnd.t45 2.82907
R19220 gnd.n22 gnd.t64 2.82907
R19221 gnd.n20 gnd.t146 2.82907
R19222 gnd.n20 gnd.t111 2.82907
R19223 gnd.n18 gnd.t97 2.82907
R19224 gnd.n18 gnd.t23 2.82907
R19225 gnd.n16 gnd.t160 2.82907
R19226 gnd.n16 gnd.t86 2.82907
R19227 gnd.n43 gnd.t127 2.82907
R19228 gnd.n43 gnd.t143 2.82907
R19229 gnd.n41 gnd.t142 2.82907
R19230 gnd.n41 gnd.t122 2.82907
R19231 gnd.n39 gnd.t117 2.82907
R19232 gnd.n39 gnd.t22 2.82907
R19233 gnd.n37 gnd.t20 2.82907
R19234 gnd.n37 gnd.t140 2.82907
R19235 gnd.n35 gnd.t150 2.82907
R19236 gnd.n35 gnd.t158 2.82907
R19237 gnd.n33 gnd.t157 2.82907
R19238 gnd.n33 gnd.t18 2.82907
R19239 gnd.n31 gnd.t16 2.82907
R19240 gnd.n31 gnd.t40 2.82907
R19241 gnd.n59 gnd.t113 2.82907
R19242 gnd.n59 gnd.t31 2.82907
R19243 gnd.n57 gnd.t138 2.82907
R19244 gnd.n57 gnd.t53 2.82907
R19245 gnd.n55 gnd.t156 2.82907
R19246 gnd.n55 gnd.t126 2.82907
R19247 gnd.n53 gnd.t96 2.82907
R19248 gnd.n53 gnd.t110 2.82907
R19249 gnd.n51 gnd.t112 2.82907
R19250 gnd.n51 gnd.t131 2.82907
R19251 gnd.n49 gnd.t105 2.82907
R19252 gnd.n49 gnd.t71 2.82907
R19253 gnd.n47 gnd.t171 2.82907
R19254 gnd.n47 gnd.t91 2.82907
R19255 gnd.n3587 gnd.n3586 2.71565
R19256 gnd.n3555 gnd.n3554 2.71565
R19257 gnd.n3523 gnd.n3522 2.71565
R19258 gnd.n3492 gnd.n3491 2.71565
R19259 gnd.n3460 gnd.n3459 2.71565
R19260 gnd.n3428 gnd.n3427 2.71565
R19261 gnd.n3396 gnd.n3395 2.71565
R19262 gnd.n3365 gnd.n3364 2.71565
R19263 gnd.n4561 gnd.t251 2.54975
R19264 gnd.t174 gnd.n4682 2.54975
R19265 gnd.n4996 gnd.t194 2.54975
R19266 gnd.n5027 gnd.t317 2.54975
R19267 gnd.n3122 gnd.n2544 2.27742
R19268 gnd.n3122 gnd.n2479 2.27742
R19269 gnd.n3122 gnd.n2478 2.27742
R19270 gnd.n3122 gnd.n2477 2.27742
R19271 gnd.n2976 gnd.t279 2.23109
R19272 gnd.n2599 gnd.t334 2.23109
R19273 gnd.n4752 gnd.t175 2.23109
R19274 gnd.t179 gnd.n1572 2.23109
R19275 gnd.n3583 gnd.n3573 1.93989
R19276 gnd.n3551 gnd.n3541 1.93989
R19277 gnd.n3519 gnd.n3509 1.93989
R19278 gnd.n3488 gnd.n3478 1.93989
R19279 gnd.n3456 gnd.n3446 1.93989
R19280 gnd.n3424 gnd.n3414 1.93989
R19281 gnd.n3392 gnd.n3382 1.93989
R19282 gnd.n3361 gnd.n3351 1.93989
R19283 gnd.t276 gnd.n5826 1.91244
R19284 gnd.n4664 gnd.n4663 1.91244
R19285 gnd.n4700 gnd.n1674 1.91244
R19286 gnd.n4796 gnd.n4795 1.91244
R19287 gnd.n4793 gnd.t320 1.91244
R19288 gnd.t328 gnd.n1593 1.91244
R19289 gnd.n4848 gnd.n4847 1.91244
R19290 gnd.n1543 gnd.n1542 1.91244
R19291 gnd.n5014 gnd.n1505 1.91244
R19292 gnd.t317 gnd.n1496 1.91244
R19293 gnd.t356 gnd.n2987 1.59378
R19294 gnd.n3166 gnd.t331 1.59378
R19295 gnd.n2412 gnd.t0 1.59378
R19296 gnd.t184 gnd.n1706 1.59378
R19297 gnd.n5021 gnd.t195 1.59378
R19298 gnd.t200 gnd.n1124 1.27512
R19299 gnd.n5027 gnd.t236 1.27512
R19300 gnd.n5192 gnd.t289 1.27512
R19301 gnd.n2829 gnd.n2821 1.16414
R19302 gnd.n3645 gnd.n2314 1.16414
R19303 gnd.n3582 gnd.n3575 1.16414
R19304 gnd.n3550 gnd.n3543 1.16414
R19305 gnd.n3518 gnd.n3511 1.16414
R19306 gnd.n3487 gnd.n3480 1.16414
R19307 gnd.n3455 gnd.n3448 1.16414
R19308 gnd.n3423 gnd.n3416 1.16414
R19309 gnd.n3391 gnd.n3384 1.16414
R19310 gnd.n3360 gnd.n3353 1.16414
R19311 gnd.n5655 gnd.n5654 0.970197
R19312 gnd.n5901 gnd.n1045 0.970197
R19313 gnd.n3566 gnd.n3534 0.962709
R19314 gnd.n3598 gnd.n3566 0.962709
R19315 gnd.n3439 gnd.n3407 0.962709
R19316 gnd.n3471 gnd.n3439 0.962709
R19317 gnd.n3075 gnd.t186 0.956468
R19318 gnd.n3240 gnd.t330 0.956468
R19319 gnd.n4510 gnd.t11 0.956468
R19320 gnd.n1395 gnd.t182 0.956468
R19321 gnd.n2 gnd.n1 0.672012
R19322 gnd.n3 gnd.n2 0.672012
R19323 gnd.n4 gnd.n3 0.672012
R19324 gnd.n5 gnd.n4 0.672012
R19325 gnd.n6 gnd.n5 0.672012
R19326 gnd.n7 gnd.n6 0.672012
R19327 gnd.n9 gnd.n8 0.672012
R19328 gnd.n10 gnd.n9 0.672012
R19329 gnd.n11 gnd.n10 0.672012
R19330 gnd.n12 gnd.n11 0.672012
R19331 gnd.n13 gnd.n12 0.672012
R19332 gnd.n14 gnd.n13 0.672012
R19333 gnd.n4671 gnd.n1696 0.637812
R19334 gnd.n4690 gnd.n4689 0.637812
R19335 gnd.n1621 gnd.n1620 0.637812
R19336 gnd.n1612 gnd.n1600 0.637812
R19337 gnd.n4875 gnd.n4874 0.637812
R19338 gnd.n5004 gnd.n5003 0.637812
R19339 gnd gnd.n0 0.59317
R19340 gnd.n2541 gnd.n2540 0.573776
R19341 gnd.n2540 gnd.n2538 0.573776
R19342 gnd.n2538 gnd.n2536 0.573776
R19343 gnd.n2536 gnd.n2534 0.573776
R19344 gnd.n2534 gnd.n2532 0.573776
R19345 gnd.n2532 gnd.n2530 0.573776
R19346 gnd.n2530 gnd.n2528 0.573776
R19347 gnd.n2494 gnd.n2493 0.573776
R19348 gnd.n2493 gnd.n2491 0.573776
R19349 gnd.n2491 gnd.n2489 0.573776
R19350 gnd.n2489 gnd.n2487 0.573776
R19351 gnd.n2487 gnd.n2485 0.573776
R19352 gnd.n2485 gnd.n2483 0.573776
R19353 gnd.n2483 gnd.n2481 0.573776
R19354 gnd.n2509 gnd.n2508 0.573776
R19355 gnd.n2508 gnd.n2506 0.573776
R19356 gnd.n2506 gnd.n2504 0.573776
R19357 gnd.n2504 gnd.n2502 0.573776
R19358 gnd.n2502 gnd.n2500 0.573776
R19359 gnd.n2500 gnd.n2498 0.573776
R19360 gnd.n2498 gnd.n2496 0.573776
R19361 gnd.n2525 gnd.n2524 0.573776
R19362 gnd.n2524 gnd.n2522 0.573776
R19363 gnd.n2522 gnd.n2520 0.573776
R19364 gnd.n2520 gnd.n2518 0.573776
R19365 gnd.n2518 gnd.n2516 0.573776
R19366 gnd.n2516 gnd.n2514 0.573776
R19367 gnd.n2514 gnd.n2512 0.573776
R19368 gnd.n66 gnd.n64 0.573776
R19369 gnd.n68 gnd.n66 0.573776
R19370 gnd.n70 gnd.n68 0.573776
R19371 gnd.n72 gnd.n70 0.573776
R19372 gnd.n74 gnd.n72 0.573776
R19373 gnd.n76 gnd.n74 0.573776
R19374 gnd.n77 gnd.n76 0.573776
R19375 gnd.n19 gnd.n17 0.573776
R19376 gnd.n21 gnd.n19 0.573776
R19377 gnd.n23 gnd.n21 0.573776
R19378 gnd.n25 gnd.n23 0.573776
R19379 gnd.n27 gnd.n25 0.573776
R19380 gnd.n29 gnd.n27 0.573776
R19381 gnd.n30 gnd.n29 0.573776
R19382 gnd.n34 gnd.n32 0.573776
R19383 gnd.n36 gnd.n34 0.573776
R19384 gnd.n38 gnd.n36 0.573776
R19385 gnd.n40 gnd.n38 0.573776
R19386 gnd.n42 gnd.n40 0.573776
R19387 gnd.n44 gnd.n42 0.573776
R19388 gnd.n45 gnd.n44 0.573776
R19389 gnd.n50 gnd.n48 0.573776
R19390 gnd.n52 gnd.n50 0.573776
R19391 gnd.n54 gnd.n52 0.573776
R19392 gnd.n56 gnd.n54 0.573776
R19393 gnd.n58 gnd.n56 0.573776
R19394 gnd.n60 gnd.n58 0.573776
R19395 gnd.n61 gnd.n60 0.573776
R19396 gnd.n7198 gnd.n7197 0.553533
R19397 gnd.n6949 gnd.n6894 0.505073
R19398 gnd.n3883 gnd.n3881 0.505073
R19399 gnd.n5719 gnd.n5718 0.489829
R19400 gnd.n4477 gnd.n4476 0.489829
R19401 gnd.n1945 gnd.n1942 0.489829
R19402 gnd.n5245 gnd.n5244 0.489829
R19403 gnd.n3302 gnd.n2318 0.486781
R19404 gnd.n2878 gnd.n2877 0.48678
R19405 gnd.n3619 gnd.n2272 0.480683
R19406 gnd.n2962 gnd.n2961 0.480683
R19407 gnd.n5294 gnd.n1282 0.470012
R19408 gnd.n7115 gnd.n7114 0.470012
R19409 gnd.n5955 gnd.n5954 0.470012
R19410 gnd.n3765 gnd.n2234 0.470012
R19411 gnd.n6180 gnd.n6179 0.416659
R19412 gnd.n6502 gnd.n6501 0.416659
R19413 gnd.n6713 gnd.n394 0.416659
R19414 gnd.n4298 gnd.n881 0.416659
R19415 gnd.n4444 gnd.n1879 0.388379
R19416 gnd.n3579 gnd.n3578 0.388379
R19417 gnd.n3547 gnd.n3546 0.388379
R19418 gnd.n3515 gnd.n3514 0.388379
R19419 gnd.n3484 gnd.n3483 0.388379
R19420 gnd.n3452 gnd.n3451 0.388379
R19421 gnd.n3420 gnd.n3419 0.388379
R19422 gnd.n3388 gnd.n3387 0.388379
R19423 gnd.n3357 gnd.n3356 0.388379
R19424 gnd.n5547 gnd.n5527 0.388379
R19425 gnd.n7198 gnd.n15 0.374463
R19426 gnd.n2374 gnd.t342 0.319156
R19427 gnd.t320 gnd.t350 0.319156
R19428 gnd.t348 gnd.t328 0.319156
R19429 gnd.n2796 gnd.n2774 0.311721
R19430 gnd gnd.n7198 0.295112
R19431 gnd.n6991 gnd.n308 0.293183
R19432 gnd.n3921 gnd.n3920 0.293183
R19433 gnd.n4367 gnd.n1844 0.27489
R19434 gnd.n5369 gnd.n1212 0.27489
R19435 gnd.n3690 gnd.n3689 0.268793
R19436 gnd.n5593 gnd.n5592 0.258122
R19437 gnd.n6992 gnd.n6991 0.258122
R19438 gnd.n4378 gnd.n2050 0.258122
R19439 gnd.n3922 gnd.n3921 0.258122
R19440 gnd.n3689 gnd.n3688 0.241354
R19441 gnd.n1312 gnd.n1309 0.229039
R19442 gnd.n1313 gnd.n1312 0.229039
R19443 gnd.n1047 gnd.n1044 0.229039
R19444 gnd.n1975 gnd.n1047 0.229039
R19445 gnd.n2950 gnd.n2749 0.206293
R19446 gnd.n2543 gnd.n0 0.169152
R19447 gnd.n3596 gnd.n3568 0.155672
R19448 gnd.n3589 gnd.n3568 0.155672
R19449 gnd.n3589 gnd.n3588 0.155672
R19450 gnd.n3588 gnd.n3572 0.155672
R19451 gnd.n3581 gnd.n3572 0.155672
R19452 gnd.n3581 gnd.n3580 0.155672
R19453 gnd.n3564 gnd.n3536 0.155672
R19454 gnd.n3557 gnd.n3536 0.155672
R19455 gnd.n3557 gnd.n3556 0.155672
R19456 gnd.n3556 gnd.n3540 0.155672
R19457 gnd.n3549 gnd.n3540 0.155672
R19458 gnd.n3549 gnd.n3548 0.155672
R19459 gnd.n3532 gnd.n3504 0.155672
R19460 gnd.n3525 gnd.n3504 0.155672
R19461 gnd.n3525 gnd.n3524 0.155672
R19462 gnd.n3524 gnd.n3508 0.155672
R19463 gnd.n3517 gnd.n3508 0.155672
R19464 gnd.n3517 gnd.n3516 0.155672
R19465 gnd.n3501 gnd.n3473 0.155672
R19466 gnd.n3494 gnd.n3473 0.155672
R19467 gnd.n3494 gnd.n3493 0.155672
R19468 gnd.n3493 gnd.n3477 0.155672
R19469 gnd.n3486 gnd.n3477 0.155672
R19470 gnd.n3486 gnd.n3485 0.155672
R19471 gnd.n3469 gnd.n3441 0.155672
R19472 gnd.n3462 gnd.n3441 0.155672
R19473 gnd.n3462 gnd.n3461 0.155672
R19474 gnd.n3461 gnd.n3445 0.155672
R19475 gnd.n3454 gnd.n3445 0.155672
R19476 gnd.n3454 gnd.n3453 0.155672
R19477 gnd.n3437 gnd.n3409 0.155672
R19478 gnd.n3430 gnd.n3409 0.155672
R19479 gnd.n3430 gnd.n3429 0.155672
R19480 gnd.n3429 gnd.n3413 0.155672
R19481 gnd.n3422 gnd.n3413 0.155672
R19482 gnd.n3422 gnd.n3421 0.155672
R19483 gnd.n3405 gnd.n3377 0.155672
R19484 gnd.n3398 gnd.n3377 0.155672
R19485 gnd.n3398 gnd.n3397 0.155672
R19486 gnd.n3397 gnd.n3381 0.155672
R19487 gnd.n3390 gnd.n3381 0.155672
R19488 gnd.n3390 gnd.n3389 0.155672
R19489 gnd.n3374 gnd.n3346 0.155672
R19490 gnd.n3367 gnd.n3346 0.155672
R19491 gnd.n3367 gnd.n3366 0.155672
R19492 gnd.n3366 gnd.n3350 0.155672
R19493 gnd.n3359 gnd.n3350 0.155672
R19494 gnd.n3359 gnd.n3358 0.155672
R19495 gnd.n1283 gnd.n1282 0.152939
R19496 gnd.n1284 gnd.n1283 0.152939
R19497 gnd.n1285 gnd.n1284 0.152939
R19498 gnd.n1286 gnd.n1285 0.152939
R19499 gnd.n1287 gnd.n1286 0.152939
R19500 gnd.n1288 gnd.n1287 0.152939
R19501 gnd.n1289 gnd.n1288 0.152939
R19502 gnd.n1290 gnd.n1289 0.152939
R19503 gnd.n1291 gnd.n1290 0.152939
R19504 gnd.n1292 gnd.n1291 0.152939
R19505 gnd.n1293 gnd.n1292 0.152939
R19506 gnd.n1294 gnd.n1293 0.152939
R19507 gnd.n1295 gnd.n1294 0.152939
R19508 gnd.n1296 gnd.n1295 0.152939
R19509 gnd.n1297 gnd.n1296 0.152939
R19510 gnd.n1298 gnd.n1297 0.152939
R19511 gnd.n1299 gnd.n1298 0.152939
R19512 gnd.n1302 gnd.n1299 0.152939
R19513 gnd.n1303 gnd.n1302 0.152939
R19514 gnd.n1304 gnd.n1303 0.152939
R19515 gnd.n1305 gnd.n1304 0.152939
R19516 gnd.n1306 gnd.n1305 0.152939
R19517 gnd.n1307 gnd.n1306 0.152939
R19518 gnd.n1308 gnd.n1307 0.152939
R19519 gnd.n1309 gnd.n1308 0.152939
R19520 gnd.n1314 gnd.n1313 0.152939
R19521 gnd.n1315 gnd.n1314 0.152939
R19522 gnd.n1316 gnd.n1315 0.152939
R19523 gnd.n1317 gnd.n1316 0.152939
R19524 gnd.n1318 gnd.n1317 0.152939
R19525 gnd.n1319 gnd.n1318 0.152939
R19526 gnd.n1320 gnd.n1319 0.152939
R19527 gnd.n1321 gnd.n1320 0.152939
R19528 gnd.n1322 gnd.n1321 0.152939
R19529 gnd.n1325 gnd.n1322 0.152939
R19530 gnd.n1326 gnd.n1325 0.152939
R19531 gnd.n1327 gnd.n1326 0.152939
R19532 gnd.n1328 gnd.n1327 0.152939
R19533 gnd.n1329 gnd.n1328 0.152939
R19534 gnd.n1330 gnd.n1329 0.152939
R19535 gnd.n1331 gnd.n1330 0.152939
R19536 gnd.n1332 gnd.n1331 0.152939
R19537 gnd.n1333 gnd.n1332 0.152939
R19538 gnd.n1334 gnd.n1333 0.152939
R19539 gnd.n1335 gnd.n1334 0.152939
R19540 gnd.n1336 gnd.n1335 0.152939
R19541 gnd.n1337 gnd.n1336 0.152939
R19542 gnd.n1338 gnd.n1337 0.152939
R19543 gnd.n1339 gnd.n1338 0.152939
R19544 gnd.n1340 gnd.n1339 0.152939
R19545 gnd.n1341 gnd.n1340 0.152939
R19546 gnd.n1342 gnd.n1341 0.152939
R19547 gnd.n1343 gnd.n1342 0.152939
R19548 gnd.n5594 gnd.n1343 0.152939
R19549 gnd.n5594 gnd.n5593 0.152939
R19550 gnd.n5298 gnd.n5294 0.152939
R19551 gnd.n5299 gnd.n5298 0.152939
R19552 gnd.n5300 gnd.n5299 0.152939
R19553 gnd.n5301 gnd.n5300 0.152939
R19554 gnd.n5302 gnd.n5301 0.152939
R19555 gnd.n5321 gnd.n5302 0.152939
R19556 gnd.n5322 gnd.n5321 0.152939
R19557 gnd.n5323 gnd.n5322 0.152939
R19558 gnd.n5324 gnd.n5323 0.152939
R19559 gnd.n5439 gnd.n5324 0.152939
R19560 gnd.n5440 gnd.n5439 0.152939
R19561 gnd.n5440 gnd.n376 0.152939
R19562 gnd.n6738 gnd.n376 0.152939
R19563 gnd.n6739 gnd.n6738 0.152939
R19564 gnd.n6740 gnd.n6739 0.152939
R19565 gnd.n6741 gnd.n6740 0.152939
R19566 gnd.n6741 gnd.n348 0.152939
R19567 gnd.n6772 gnd.n348 0.152939
R19568 gnd.n6773 gnd.n6772 0.152939
R19569 gnd.n6774 gnd.n6773 0.152939
R19570 gnd.n6775 gnd.n6774 0.152939
R19571 gnd.n113 gnd.n112 0.152939
R19572 gnd.n114 gnd.n113 0.152939
R19573 gnd.n130 gnd.n114 0.152939
R19574 gnd.n131 gnd.n130 0.152939
R19575 gnd.n132 gnd.n131 0.152939
R19576 gnd.n133 gnd.n132 0.152939
R19577 gnd.n149 gnd.n133 0.152939
R19578 gnd.n150 gnd.n149 0.152939
R19579 gnd.n151 gnd.n150 0.152939
R19580 gnd.n152 gnd.n151 0.152939
R19581 gnd.n168 gnd.n152 0.152939
R19582 gnd.n169 gnd.n168 0.152939
R19583 gnd.n170 gnd.n169 0.152939
R19584 gnd.n171 gnd.n170 0.152939
R19585 gnd.n187 gnd.n171 0.152939
R19586 gnd.n188 gnd.n187 0.152939
R19587 gnd.n189 gnd.n188 0.152939
R19588 gnd.n190 gnd.n189 0.152939
R19589 gnd.n206 gnd.n190 0.152939
R19590 gnd.n207 gnd.n206 0.152939
R19591 gnd.n7115 gnd.n207 0.152939
R19592 gnd.n7195 gnd.n80 0.152939
R19593 gnd.n6858 gnd.n80 0.152939
R19594 gnd.n6859 gnd.n6858 0.152939
R19595 gnd.n6860 gnd.n6859 0.152939
R19596 gnd.n6860 gnd.n6856 0.152939
R19597 gnd.n6866 gnd.n6856 0.152939
R19598 gnd.n6867 gnd.n6866 0.152939
R19599 gnd.n6868 gnd.n6867 0.152939
R19600 gnd.n6868 gnd.n6854 0.152939
R19601 gnd.n6874 gnd.n6854 0.152939
R19602 gnd.n6875 gnd.n6874 0.152939
R19603 gnd.n6876 gnd.n6875 0.152939
R19604 gnd.n6876 gnd.n6852 0.152939
R19605 gnd.n6882 gnd.n6852 0.152939
R19606 gnd.n6883 gnd.n6882 0.152939
R19607 gnd.n6884 gnd.n6883 0.152939
R19608 gnd.n6885 gnd.n6884 0.152939
R19609 gnd.n6886 gnd.n6885 0.152939
R19610 gnd.n6887 gnd.n6886 0.152939
R19611 gnd.n6888 gnd.n6887 0.152939
R19612 gnd.n6889 gnd.n6888 0.152939
R19613 gnd.n6890 gnd.n6889 0.152939
R19614 gnd.n6891 gnd.n6890 0.152939
R19615 gnd.n6892 gnd.n6891 0.152939
R19616 gnd.n6893 gnd.n6892 0.152939
R19617 gnd.n6894 gnd.n6893 0.152939
R19618 gnd.n6908 gnd.n308 0.152939
R19619 gnd.n6909 gnd.n6908 0.152939
R19620 gnd.n6909 gnd.n6904 0.152939
R19621 gnd.n6917 gnd.n6904 0.152939
R19622 gnd.n6918 gnd.n6917 0.152939
R19623 gnd.n6919 gnd.n6918 0.152939
R19624 gnd.n6919 gnd.n6902 0.152939
R19625 gnd.n6927 gnd.n6902 0.152939
R19626 gnd.n6928 gnd.n6927 0.152939
R19627 gnd.n6929 gnd.n6928 0.152939
R19628 gnd.n6929 gnd.n6900 0.152939
R19629 gnd.n6937 gnd.n6900 0.152939
R19630 gnd.n6938 gnd.n6937 0.152939
R19631 gnd.n6939 gnd.n6938 0.152939
R19632 gnd.n6939 gnd.n6898 0.152939
R19633 gnd.n6947 gnd.n6898 0.152939
R19634 gnd.n6948 gnd.n6947 0.152939
R19635 gnd.n6949 gnd.n6948 0.152939
R19636 gnd.n7114 gnd.n208 0.152939
R19637 gnd.n250 gnd.n208 0.152939
R19638 gnd.n251 gnd.n250 0.152939
R19639 gnd.n252 gnd.n251 0.152939
R19640 gnd.n253 gnd.n252 0.152939
R19641 gnd.n254 gnd.n253 0.152939
R19642 gnd.n255 gnd.n254 0.152939
R19643 gnd.n256 gnd.n255 0.152939
R19644 gnd.n257 gnd.n256 0.152939
R19645 gnd.n258 gnd.n257 0.152939
R19646 gnd.n259 gnd.n258 0.152939
R19647 gnd.n260 gnd.n259 0.152939
R19648 gnd.n261 gnd.n260 0.152939
R19649 gnd.n262 gnd.n261 0.152939
R19650 gnd.n263 gnd.n262 0.152939
R19651 gnd.n264 gnd.n263 0.152939
R19652 gnd.n265 gnd.n264 0.152939
R19653 gnd.n266 gnd.n265 0.152939
R19654 gnd.n267 gnd.n266 0.152939
R19655 gnd.n268 gnd.n267 0.152939
R19656 gnd.n269 gnd.n268 0.152939
R19657 gnd.n270 gnd.n269 0.152939
R19658 gnd.n271 gnd.n270 0.152939
R19659 gnd.n272 gnd.n271 0.152939
R19660 gnd.n273 gnd.n272 0.152939
R19661 gnd.n274 gnd.n273 0.152939
R19662 gnd.n275 gnd.n274 0.152939
R19663 gnd.n276 gnd.n275 0.152939
R19664 gnd.n277 gnd.n276 0.152939
R19665 gnd.n278 gnd.n277 0.152939
R19666 gnd.n279 gnd.n278 0.152939
R19667 gnd.n280 gnd.n279 0.152939
R19668 gnd.n281 gnd.n280 0.152939
R19669 gnd.n282 gnd.n281 0.152939
R19670 gnd.n283 gnd.n282 0.152939
R19671 gnd.n284 gnd.n283 0.152939
R19672 gnd.n7035 gnd.n284 0.152939
R19673 gnd.n7035 gnd.n7034 0.152939
R19674 gnd.n7034 gnd.n7033 0.152939
R19675 gnd.n7033 gnd.n288 0.152939
R19676 gnd.n289 gnd.n288 0.152939
R19677 gnd.n290 gnd.n289 0.152939
R19678 gnd.n291 gnd.n290 0.152939
R19679 gnd.n292 gnd.n291 0.152939
R19680 gnd.n293 gnd.n292 0.152939
R19681 gnd.n294 gnd.n293 0.152939
R19682 gnd.n295 gnd.n294 0.152939
R19683 gnd.n296 gnd.n295 0.152939
R19684 gnd.n297 gnd.n296 0.152939
R19685 gnd.n298 gnd.n297 0.152939
R19686 gnd.n299 gnd.n298 0.152939
R19687 gnd.n300 gnd.n299 0.152939
R19688 gnd.n301 gnd.n300 0.152939
R19689 gnd.n302 gnd.n301 0.152939
R19690 gnd.n303 gnd.n302 0.152939
R19691 gnd.n304 gnd.n303 0.152939
R19692 gnd.n6993 gnd.n304 0.152939
R19693 gnd.n6993 gnd.n6992 0.152939
R19694 gnd.n3721 gnd.n2272 0.152939
R19695 gnd.n3721 gnd.n3720 0.152939
R19696 gnd.n3720 gnd.n3719 0.152939
R19697 gnd.n3719 gnd.n2274 0.152939
R19698 gnd.n2275 gnd.n2274 0.152939
R19699 gnd.n2276 gnd.n2275 0.152939
R19700 gnd.n2277 gnd.n2276 0.152939
R19701 gnd.n2278 gnd.n2277 0.152939
R19702 gnd.n2279 gnd.n2278 0.152939
R19703 gnd.n2280 gnd.n2279 0.152939
R19704 gnd.n2281 gnd.n2280 0.152939
R19705 gnd.n2282 gnd.n2281 0.152939
R19706 gnd.n2283 gnd.n2282 0.152939
R19707 gnd.n2284 gnd.n2283 0.152939
R19708 gnd.n3691 gnd.n2284 0.152939
R19709 gnd.n3691 gnd.n3690 0.152939
R19710 gnd.n2963 gnd.n2962 0.152939
R19711 gnd.n2963 gnd.n2667 0.152939
R19712 gnd.n2991 gnd.n2667 0.152939
R19713 gnd.n2992 gnd.n2991 0.152939
R19714 gnd.n2993 gnd.n2992 0.152939
R19715 gnd.n2994 gnd.n2993 0.152939
R19716 gnd.n2994 gnd.n2639 0.152939
R19717 gnd.n3021 gnd.n2639 0.152939
R19718 gnd.n3022 gnd.n3021 0.152939
R19719 gnd.n3023 gnd.n3022 0.152939
R19720 gnd.n3023 gnd.n2617 0.152939
R19721 gnd.n3052 gnd.n2617 0.152939
R19722 gnd.n3053 gnd.n3052 0.152939
R19723 gnd.n3054 gnd.n3053 0.152939
R19724 gnd.n3055 gnd.n3054 0.152939
R19725 gnd.n3057 gnd.n3055 0.152939
R19726 gnd.n3057 gnd.n3056 0.152939
R19727 gnd.n3056 gnd.n2566 0.152939
R19728 gnd.n2567 gnd.n2566 0.152939
R19729 gnd.n2568 gnd.n2567 0.152939
R19730 gnd.n2587 gnd.n2568 0.152939
R19731 gnd.n2588 gnd.n2587 0.152939
R19732 gnd.n2588 gnd.n2470 0.152939
R19733 gnd.n3147 gnd.n2470 0.152939
R19734 gnd.n3148 gnd.n3147 0.152939
R19735 gnd.n3149 gnd.n3148 0.152939
R19736 gnd.n3150 gnd.n3149 0.152939
R19737 gnd.n3150 gnd.n2443 0.152939
R19738 gnd.n3187 gnd.n2443 0.152939
R19739 gnd.n3188 gnd.n3187 0.152939
R19740 gnd.n3189 gnd.n3188 0.152939
R19741 gnd.n3190 gnd.n3189 0.152939
R19742 gnd.n3190 gnd.n2416 0.152939
R19743 gnd.n3232 gnd.n2416 0.152939
R19744 gnd.n3233 gnd.n3232 0.152939
R19745 gnd.n3234 gnd.n3233 0.152939
R19746 gnd.n3235 gnd.n3234 0.152939
R19747 gnd.n3235 gnd.n2388 0.152939
R19748 gnd.n3272 gnd.n2388 0.152939
R19749 gnd.n3273 gnd.n3272 0.152939
R19750 gnd.n3274 gnd.n3273 0.152939
R19751 gnd.n3275 gnd.n3274 0.152939
R19752 gnd.n3275 gnd.n2361 0.152939
R19753 gnd.n3321 gnd.n2361 0.152939
R19754 gnd.n3322 gnd.n3321 0.152939
R19755 gnd.n3323 gnd.n3322 0.152939
R19756 gnd.n3324 gnd.n3323 0.152939
R19757 gnd.n3324 gnd.n2334 0.152939
R19758 gnd.n3615 gnd.n2334 0.152939
R19759 gnd.n3616 gnd.n3615 0.152939
R19760 gnd.n3617 gnd.n3616 0.152939
R19761 gnd.n3618 gnd.n3617 0.152939
R19762 gnd.n3619 gnd.n3618 0.152939
R19763 gnd.n2961 gnd.n2691 0.152939
R19764 gnd.n2712 gnd.n2691 0.152939
R19765 gnd.n2713 gnd.n2712 0.152939
R19766 gnd.n2719 gnd.n2713 0.152939
R19767 gnd.n2720 gnd.n2719 0.152939
R19768 gnd.n2721 gnd.n2720 0.152939
R19769 gnd.n2721 gnd.n2710 0.152939
R19770 gnd.n2729 gnd.n2710 0.152939
R19771 gnd.n2730 gnd.n2729 0.152939
R19772 gnd.n2731 gnd.n2730 0.152939
R19773 gnd.n2731 gnd.n2708 0.152939
R19774 gnd.n2739 gnd.n2708 0.152939
R19775 gnd.n2740 gnd.n2739 0.152939
R19776 gnd.n2741 gnd.n2740 0.152939
R19777 gnd.n2741 gnd.n2706 0.152939
R19778 gnd.n2749 gnd.n2706 0.152939
R19779 gnd.n3688 gnd.n2289 0.152939
R19780 gnd.n2291 gnd.n2289 0.152939
R19781 gnd.n2292 gnd.n2291 0.152939
R19782 gnd.n2293 gnd.n2292 0.152939
R19783 gnd.n2294 gnd.n2293 0.152939
R19784 gnd.n2295 gnd.n2294 0.152939
R19785 gnd.n2296 gnd.n2295 0.152939
R19786 gnd.n2297 gnd.n2296 0.152939
R19787 gnd.n2298 gnd.n2297 0.152939
R19788 gnd.n2299 gnd.n2298 0.152939
R19789 gnd.n2300 gnd.n2299 0.152939
R19790 gnd.n2301 gnd.n2300 0.152939
R19791 gnd.n2302 gnd.n2301 0.152939
R19792 gnd.n2303 gnd.n2302 0.152939
R19793 gnd.n2304 gnd.n2303 0.152939
R19794 gnd.n2305 gnd.n2304 0.152939
R19795 gnd.n2306 gnd.n2305 0.152939
R19796 gnd.n2307 gnd.n2306 0.152939
R19797 gnd.n2308 gnd.n2307 0.152939
R19798 gnd.n2309 gnd.n2308 0.152939
R19799 gnd.n2310 gnd.n2309 0.152939
R19800 gnd.n2311 gnd.n2310 0.152939
R19801 gnd.n2315 gnd.n2311 0.152939
R19802 gnd.n2316 gnd.n2315 0.152939
R19803 gnd.n2317 gnd.n2316 0.152939
R19804 gnd.n2318 gnd.n2317 0.152939
R19805 gnd.n3124 gnd.n3123 0.152939
R19806 gnd.n3125 gnd.n3124 0.152939
R19807 gnd.n3126 gnd.n3125 0.152939
R19808 gnd.n3127 gnd.n3126 0.152939
R19809 gnd.n3128 gnd.n3127 0.152939
R19810 gnd.n3129 gnd.n3128 0.152939
R19811 gnd.n3129 gnd.n2424 0.152939
R19812 gnd.n3208 gnd.n2424 0.152939
R19813 gnd.n3209 gnd.n3208 0.152939
R19814 gnd.n3210 gnd.n3209 0.152939
R19815 gnd.n3211 gnd.n3210 0.152939
R19816 gnd.n3212 gnd.n3211 0.152939
R19817 gnd.n3213 gnd.n3212 0.152939
R19818 gnd.n3214 gnd.n3213 0.152939
R19819 gnd.n3215 gnd.n3214 0.152939
R19820 gnd.n3216 gnd.n3215 0.152939
R19821 gnd.n3216 gnd.n2368 0.152939
R19822 gnd.n3293 gnd.n2368 0.152939
R19823 gnd.n3294 gnd.n3293 0.152939
R19824 gnd.n3295 gnd.n3294 0.152939
R19825 gnd.n3296 gnd.n3295 0.152939
R19826 gnd.n3297 gnd.n3296 0.152939
R19827 gnd.n3298 gnd.n3297 0.152939
R19828 gnd.n3299 gnd.n3298 0.152939
R19829 gnd.n3300 gnd.n3299 0.152939
R19830 gnd.n3301 gnd.n3300 0.152939
R19831 gnd.n3303 gnd.n3301 0.152939
R19832 gnd.n3303 gnd.n3302 0.152939
R19833 gnd.n2879 gnd.n2878 0.152939
R19834 gnd.n2879 gnd.n2769 0.152939
R19835 gnd.n2894 gnd.n2769 0.152939
R19836 gnd.n2895 gnd.n2894 0.152939
R19837 gnd.n2896 gnd.n2895 0.152939
R19838 gnd.n2896 gnd.n2757 0.152939
R19839 gnd.n2910 gnd.n2757 0.152939
R19840 gnd.n2911 gnd.n2910 0.152939
R19841 gnd.n2912 gnd.n2911 0.152939
R19842 gnd.n2913 gnd.n2912 0.152939
R19843 gnd.n2914 gnd.n2913 0.152939
R19844 gnd.n2915 gnd.n2914 0.152939
R19845 gnd.n2916 gnd.n2915 0.152939
R19846 gnd.n2917 gnd.n2916 0.152939
R19847 gnd.n2918 gnd.n2917 0.152939
R19848 gnd.n2919 gnd.n2918 0.152939
R19849 gnd.n2920 gnd.n2919 0.152939
R19850 gnd.n2921 gnd.n2920 0.152939
R19851 gnd.n2922 gnd.n2921 0.152939
R19852 gnd.n2923 gnd.n2922 0.152939
R19853 gnd.n2924 gnd.n2923 0.152939
R19854 gnd.n2924 gnd.n2623 0.152939
R19855 gnd.n3041 gnd.n2623 0.152939
R19856 gnd.n3042 gnd.n3041 0.152939
R19857 gnd.n3043 gnd.n3042 0.152939
R19858 gnd.n3044 gnd.n3043 0.152939
R19859 gnd.n3044 gnd.n2545 0.152939
R19860 gnd.n3121 gnd.n2545 0.152939
R19861 gnd.n2797 gnd.n2796 0.152939
R19862 gnd.n2798 gnd.n2797 0.152939
R19863 gnd.n2799 gnd.n2798 0.152939
R19864 gnd.n2800 gnd.n2799 0.152939
R19865 gnd.n2801 gnd.n2800 0.152939
R19866 gnd.n2802 gnd.n2801 0.152939
R19867 gnd.n2803 gnd.n2802 0.152939
R19868 gnd.n2804 gnd.n2803 0.152939
R19869 gnd.n2805 gnd.n2804 0.152939
R19870 gnd.n2806 gnd.n2805 0.152939
R19871 gnd.n2807 gnd.n2806 0.152939
R19872 gnd.n2808 gnd.n2807 0.152939
R19873 gnd.n2809 gnd.n2808 0.152939
R19874 gnd.n2810 gnd.n2809 0.152939
R19875 gnd.n2811 gnd.n2810 0.152939
R19876 gnd.n2812 gnd.n2811 0.152939
R19877 gnd.n2813 gnd.n2812 0.152939
R19878 gnd.n2814 gnd.n2813 0.152939
R19879 gnd.n2815 gnd.n2814 0.152939
R19880 gnd.n2816 gnd.n2815 0.152939
R19881 gnd.n2817 gnd.n2816 0.152939
R19882 gnd.n2818 gnd.n2817 0.152939
R19883 gnd.n2822 gnd.n2818 0.152939
R19884 gnd.n2823 gnd.n2822 0.152939
R19885 gnd.n2823 gnd.n2780 0.152939
R19886 gnd.n2877 gnd.n2780 0.152939
R19887 gnd.n3881 gnd.n3847 0.152939
R19888 gnd.n3848 gnd.n3847 0.152939
R19889 gnd.n3849 gnd.n3848 0.152939
R19890 gnd.n3850 gnd.n3849 0.152939
R19891 gnd.n3851 gnd.n3850 0.152939
R19892 gnd.n3852 gnd.n3851 0.152939
R19893 gnd.n3853 gnd.n3852 0.152939
R19894 gnd.n3854 gnd.n3853 0.152939
R19895 gnd.n3855 gnd.n3854 0.152939
R19896 gnd.n3856 gnd.n3855 0.152939
R19897 gnd.n3857 gnd.n3856 0.152939
R19898 gnd.n3858 gnd.n3857 0.152939
R19899 gnd.n3859 gnd.n3858 0.152939
R19900 gnd.n3859 gnd.n2170 0.152939
R19901 gnd.n4129 gnd.n2170 0.152939
R19902 gnd.n4130 gnd.n4129 0.152939
R19903 gnd.n4131 gnd.n4130 0.152939
R19904 gnd.n4132 gnd.n4131 0.152939
R19905 gnd.n4132 gnd.n2145 0.152939
R19906 gnd.n4164 gnd.n2145 0.152939
R19907 gnd.n4165 gnd.n4164 0.152939
R19908 gnd.n4166 gnd.n4165 0.152939
R19909 gnd.n4167 gnd.n4166 0.152939
R19910 gnd.n4167 gnd.n2120 0.152939
R19911 gnd.n4199 gnd.n2120 0.152939
R19912 gnd.n4200 gnd.n4199 0.152939
R19913 gnd.n5954 gnd.n975 0.152939
R19914 gnd.n1019 gnd.n975 0.152939
R19915 gnd.n1020 gnd.n1019 0.152939
R19916 gnd.n1021 gnd.n1020 0.152939
R19917 gnd.n1022 gnd.n1021 0.152939
R19918 gnd.n1023 gnd.n1022 0.152939
R19919 gnd.n1024 gnd.n1023 0.152939
R19920 gnd.n1025 gnd.n1024 0.152939
R19921 gnd.n1026 gnd.n1025 0.152939
R19922 gnd.n1027 gnd.n1026 0.152939
R19923 gnd.n1028 gnd.n1027 0.152939
R19924 gnd.n1029 gnd.n1028 0.152939
R19925 gnd.n1030 gnd.n1029 0.152939
R19926 gnd.n1031 gnd.n1030 0.152939
R19927 gnd.n1032 gnd.n1031 0.152939
R19928 gnd.n1033 gnd.n1032 0.152939
R19929 gnd.n1034 gnd.n1033 0.152939
R19930 gnd.n1037 gnd.n1034 0.152939
R19931 gnd.n1038 gnd.n1037 0.152939
R19932 gnd.n1039 gnd.n1038 0.152939
R19933 gnd.n1040 gnd.n1039 0.152939
R19934 gnd.n1041 gnd.n1040 0.152939
R19935 gnd.n1042 gnd.n1041 0.152939
R19936 gnd.n1043 gnd.n1042 0.152939
R19937 gnd.n1044 gnd.n1043 0.152939
R19938 gnd.n1976 gnd.n1975 0.152939
R19939 gnd.n1983 gnd.n1976 0.152939
R19940 gnd.n1984 gnd.n1983 0.152939
R19941 gnd.n1985 gnd.n1984 0.152939
R19942 gnd.n1985 gnd.n1973 0.152939
R19943 gnd.n1993 gnd.n1973 0.152939
R19944 gnd.n1994 gnd.n1993 0.152939
R19945 gnd.n1995 gnd.n1994 0.152939
R19946 gnd.n1995 gnd.n1968 0.152939
R19947 gnd.n2002 gnd.n1968 0.152939
R19948 gnd.n2003 gnd.n2002 0.152939
R19949 gnd.n2004 gnd.n2003 0.152939
R19950 gnd.n2004 gnd.n1966 0.152939
R19951 gnd.n2012 gnd.n1966 0.152939
R19952 gnd.n2013 gnd.n2012 0.152939
R19953 gnd.n2014 gnd.n2013 0.152939
R19954 gnd.n2014 gnd.n1964 0.152939
R19955 gnd.n2022 gnd.n1964 0.152939
R19956 gnd.n2023 gnd.n2022 0.152939
R19957 gnd.n2024 gnd.n2023 0.152939
R19958 gnd.n2024 gnd.n1962 0.152939
R19959 gnd.n2032 gnd.n1962 0.152939
R19960 gnd.n2033 gnd.n2032 0.152939
R19961 gnd.n2034 gnd.n2033 0.152939
R19962 gnd.n2034 gnd.n1960 0.152939
R19963 gnd.n2042 gnd.n1960 0.152939
R19964 gnd.n2043 gnd.n2042 0.152939
R19965 gnd.n2044 gnd.n2043 0.152939
R19966 gnd.n2044 gnd.n1955 0.152939
R19967 gnd.n2050 gnd.n1955 0.152939
R19968 gnd.n4260 gnd.n4259 0.152939
R19969 gnd.n4262 gnd.n4260 0.152939
R19970 gnd.n4262 gnd.n4261 0.152939
R19971 gnd.n4261 gnd.n891 0.152939
R19972 gnd.n892 gnd.n891 0.152939
R19973 gnd.n893 gnd.n892 0.152939
R19974 gnd.n912 gnd.n893 0.152939
R19975 gnd.n913 gnd.n912 0.152939
R19976 gnd.n914 gnd.n913 0.152939
R19977 gnd.n915 gnd.n914 0.152939
R19978 gnd.n932 gnd.n915 0.152939
R19979 gnd.n933 gnd.n932 0.152939
R19980 gnd.n934 gnd.n933 0.152939
R19981 gnd.n935 gnd.n934 0.152939
R19982 gnd.n952 gnd.n935 0.152939
R19983 gnd.n953 gnd.n952 0.152939
R19984 gnd.n954 gnd.n953 0.152939
R19985 gnd.n955 gnd.n954 0.152939
R19986 gnd.n973 gnd.n955 0.152939
R19987 gnd.n974 gnd.n973 0.152939
R19988 gnd.n5955 gnd.n974 0.152939
R19989 gnd.n4055 gnd.n2234 0.152939
R19990 gnd.n4056 gnd.n4055 0.152939
R19991 gnd.n4057 gnd.n4056 0.152939
R19992 gnd.n4057 gnd.n2215 0.152939
R19993 gnd.n4075 gnd.n2215 0.152939
R19994 gnd.n4076 gnd.n4075 0.152939
R19995 gnd.n4077 gnd.n4076 0.152939
R19996 gnd.n4077 gnd.n2198 0.152939
R19997 gnd.n4095 gnd.n2198 0.152939
R19998 gnd.n4096 gnd.n4095 0.152939
R19999 gnd.n4097 gnd.n4096 0.152939
R20000 gnd.n4097 gnd.n2178 0.152939
R20001 gnd.n4119 gnd.n2178 0.152939
R20002 gnd.n4120 gnd.n4119 0.152939
R20003 gnd.n4121 gnd.n4120 0.152939
R20004 gnd.n4122 gnd.n4121 0.152939
R20005 gnd.n4122 gnd.n2153 0.152939
R20006 gnd.n4154 gnd.n2153 0.152939
R20007 gnd.n4155 gnd.n4154 0.152939
R20008 gnd.n4156 gnd.n4155 0.152939
R20009 gnd.n4157 gnd.n4156 0.152939
R20010 gnd.n3766 gnd.n3765 0.152939
R20011 gnd.n3767 gnd.n3766 0.152939
R20012 gnd.n3768 gnd.n3767 0.152939
R20013 gnd.n3769 gnd.n3768 0.152939
R20014 gnd.n3770 gnd.n3769 0.152939
R20015 gnd.n3771 gnd.n3770 0.152939
R20016 gnd.n3772 gnd.n3771 0.152939
R20017 gnd.n3773 gnd.n3772 0.152939
R20018 gnd.n3774 gnd.n3773 0.152939
R20019 gnd.n3775 gnd.n3774 0.152939
R20020 gnd.n3776 gnd.n3775 0.152939
R20021 gnd.n3777 gnd.n3776 0.152939
R20022 gnd.n3778 gnd.n3777 0.152939
R20023 gnd.n3779 gnd.n3778 0.152939
R20024 gnd.n3780 gnd.n3779 0.152939
R20025 gnd.n3781 gnd.n3780 0.152939
R20026 gnd.n3782 gnd.n3781 0.152939
R20027 gnd.n3785 gnd.n3782 0.152939
R20028 gnd.n3786 gnd.n3785 0.152939
R20029 gnd.n3787 gnd.n3786 0.152939
R20030 gnd.n3788 gnd.n3787 0.152939
R20031 gnd.n3789 gnd.n3788 0.152939
R20032 gnd.n3790 gnd.n3789 0.152939
R20033 gnd.n3791 gnd.n3790 0.152939
R20034 gnd.n3792 gnd.n3791 0.152939
R20035 gnd.n3793 gnd.n3792 0.152939
R20036 gnd.n3794 gnd.n3793 0.152939
R20037 gnd.n3795 gnd.n3794 0.152939
R20038 gnd.n3796 gnd.n3795 0.152939
R20039 gnd.n3797 gnd.n3796 0.152939
R20040 gnd.n3798 gnd.n3797 0.152939
R20041 gnd.n3799 gnd.n3798 0.152939
R20042 gnd.n3800 gnd.n3799 0.152939
R20043 gnd.n3801 gnd.n3800 0.152939
R20044 gnd.n3802 gnd.n3801 0.152939
R20045 gnd.n3803 gnd.n3802 0.152939
R20046 gnd.n3804 gnd.n3803 0.152939
R20047 gnd.n3807 gnd.n3804 0.152939
R20048 gnd.n3808 gnd.n3807 0.152939
R20049 gnd.n3809 gnd.n3808 0.152939
R20050 gnd.n3810 gnd.n3809 0.152939
R20051 gnd.n3811 gnd.n3810 0.152939
R20052 gnd.n3812 gnd.n3811 0.152939
R20053 gnd.n3813 gnd.n3812 0.152939
R20054 gnd.n3814 gnd.n3813 0.152939
R20055 gnd.n3815 gnd.n3814 0.152939
R20056 gnd.n3816 gnd.n3815 0.152939
R20057 gnd.n3817 gnd.n3816 0.152939
R20058 gnd.n3818 gnd.n3817 0.152939
R20059 gnd.n3819 gnd.n3818 0.152939
R20060 gnd.n3820 gnd.n3819 0.152939
R20061 gnd.n3821 gnd.n3820 0.152939
R20062 gnd.n3822 gnd.n3821 0.152939
R20063 gnd.n3823 gnd.n3822 0.152939
R20064 gnd.n3824 gnd.n3823 0.152939
R20065 gnd.n3825 gnd.n3824 0.152939
R20066 gnd.n3923 gnd.n3825 0.152939
R20067 gnd.n3923 gnd.n3922 0.152939
R20068 gnd.n3920 gnd.n3828 0.152939
R20069 gnd.n3829 gnd.n3828 0.152939
R20070 gnd.n3830 gnd.n3829 0.152939
R20071 gnd.n3831 gnd.n3830 0.152939
R20072 gnd.n3832 gnd.n3831 0.152939
R20073 gnd.n3833 gnd.n3832 0.152939
R20074 gnd.n3834 gnd.n3833 0.152939
R20075 gnd.n3835 gnd.n3834 0.152939
R20076 gnd.n3836 gnd.n3835 0.152939
R20077 gnd.n3837 gnd.n3836 0.152939
R20078 gnd.n3838 gnd.n3837 0.152939
R20079 gnd.n3839 gnd.n3838 0.152939
R20080 gnd.n3840 gnd.n3839 0.152939
R20081 gnd.n3841 gnd.n3840 0.152939
R20082 gnd.n3842 gnd.n3841 0.152939
R20083 gnd.n3885 gnd.n3842 0.152939
R20084 gnd.n3885 gnd.n3884 0.152939
R20085 gnd.n3884 gnd.n3883 0.152939
R20086 gnd.n6181 gnd.n6180 0.152939
R20087 gnd.n6181 gnd.n708 0.152939
R20088 gnd.n6189 gnd.n708 0.152939
R20089 gnd.n6190 gnd.n6189 0.152939
R20090 gnd.n6191 gnd.n6190 0.152939
R20091 gnd.n6191 gnd.n702 0.152939
R20092 gnd.n6199 gnd.n702 0.152939
R20093 gnd.n6200 gnd.n6199 0.152939
R20094 gnd.n6201 gnd.n6200 0.152939
R20095 gnd.n6201 gnd.n696 0.152939
R20096 gnd.n6209 gnd.n696 0.152939
R20097 gnd.n6210 gnd.n6209 0.152939
R20098 gnd.n6211 gnd.n6210 0.152939
R20099 gnd.n6211 gnd.n690 0.152939
R20100 gnd.n6219 gnd.n690 0.152939
R20101 gnd.n6220 gnd.n6219 0.152939
R20102 gnd.n6221 gnd.n6220 0.152939
R20103 gnd.n6221 gnd.n684 0.152939
R20104 gnd.n6229 gnd.n684 0.152939
R20105 gnd.n6230 gnd.n6229 0.152939
R20106 gnd.n6231 gnd.n6230 0.152939
R20107 gnd.n6231 gnd.n678 0.152939
R20108 gnd.n6239 gnd.n678 0.152939
R20109 gnd.n6240 gnd.n6239 0.152939
R20110 gnd.n6241 gnd.n6240 0.152939
R20111 gnd.n6241 gnd.n672 0.152939
R20112 gnd.n6249 gnd.n672 0.152939
R20113 gnd.n6250 gnd.n6249 0.152939
R20114 gnd.n6251 gnd.n6250 0.152939
R20115 gnd.n6251 gnd.n666 0.152939
R20116 gnd.n6259 gnd.n666 0.152939
R20117 gnd.n6260 gnd.n6259 0.152939
R20118 gnd.n6261 gnd.n6260 0.152939
R20119 gnd.n6261 gnd.n660 0.152939
R20120 gnd.n6269 gnd.n660 0.152939
R20121 gnd.n6270 gnd.n6269 0.152939
R20122 gnd.n6271 gnd.n6270 0.152939
R20123 gnd.n6271 gnd.n654 0.152939
R20124 gnd.n6279 gnd.n654 0.152939
R20125 gnd.n6280 gnd.n6279 0.152939
R20126 gnd.n6281 gnd.n6280 0.152939
R20127 gnd.n6281 gnd.n648 0.152939
R20128 gnd.n6289 gnd.n648 0.152939
R20129 gnd.n6290 gnd.n6289 0.152939
R20130 gnd.n6291 gnd.n6290 0.152939
R20131 gnd.n6291 gnd.n642 0.152939
R20132 gnd.n6299 gnd.n642 0.152939
R20133 gnd.n6300 gnd.n6299 0.152939
R20134 gnd.n6301 gnd.n6300 0.152939
R20135 gnd.n6301 gnd.n636 0.152939
R20136 gnd.n6309 gnd.n636 0.152939
R20137 gnd.n6310 gnd.n6309 0.152939
R20138 gnd.n6311 gnd.n6310 0.152939
R20139 gnd.n6311 gnd.n630 0.152939
R20140 gnd.n6319 gnd.n630 0.152939
R20141 gnd.n6320 gnd.n6319 0.152939
R20142 gnd.n6321 gnd.n6320 0.152939
R20143 gnd.n6321 gnd.n624 0.152939
R20144 gnd.n6329 gnd.n624 0.152939
R20145 gnd.n6330 gnd.n6329 0.152939
R20146 gnd.n6331 gnd.n6330 0.152939
R20147 gnd.n6331 gnd.n618 0.152939
R20148 gnd.n6339 gnd.n618 0.152939
R20149 gnd.n6340 gnd.n6339 0.152939
R20150 gnd.n6341 gnd.n6340 0.152939
R20151 gnd.n6341 gnd.n612 0.152939
R20152 gnd.n6349 gnd.n612 0.152939
R20153 gnd.n6350 gnd.n6349 0.152939
R20154 gnd.n6351 gnd.n6350 0.152939
R20155 gnd.n6351 gnd.n606 0.152939
R20156 gnd.n6359 gnd.n606 0.152939
R20157 gnd.n6360 gnd.n6359 0.152939
R20158 gnd.n6361 gnd.n6360 0.152939
R20159 gnd.n6361 gnd.n600 0.152939
R20160 gnd.n6369 gnd.n600 0.152939
R20161 gnd.n6370 gnd.n6369 0.152939
R20162 gnd.n6371 gnd.n6370 0.152939
R20163 gnd.n6371 gnd.n594 0.152939
R20164 gnd.n6379 gnd.n594 0.152939
R20165 gnd.n6380 gnd.n6379 0.152939
R20166 gnd.n6381 gnd.n6380 0.152939
R20167 gnd.n6381 gnd.n588 0.152939
R20168 gnd.n6389 gnd.n588 0.152939
R20169 gnd.n6390 gnd.n6389 0.152939
R20170 gnd.n6391 gnd.n6390 0.152939
R20171 gnd.n6391 gnd.n582 0.152939
R20172 gnd.n6399 gnd.n582 0.152939
R20173 gnd.n6400 gnd.n6399 0.152939
R20174 gnd.n6401 gnd.n6400 0.152939
R20175 gnd.n6401 gnd.n576 0.152939
R20176 gnd.n6409 gnd.n576 0.152939
R20177 gnd.n6410 gnd.n6409 0.152939
R20178 gnd.n6411 gnd.n6410 0.152939
R20179 gnd.n6411 gnd.n570 0.152939
R20180 gnd.n6419 gnd.n570 0.152939
R20181 gnd.n6420 gnd.n6419 0.152939
R20182 gnd.n6421 gnd.n6420 0.152939
R20183 gnd.n6421 gnd.n564 0.152939
R20184 gnd.n6429 gnd.n564 0.152939
R20185 gnd.n6430 gnd.n6429 0.152939
R20186 gnd.n6431 gnd.n6430 0.152939
R20187 gnd.n6431 gnd.n558 0.152939
R20188 gnd.n6439 gnd.n558 0.152939
R20189 gnd.n6440 gnd.n6439 0.152939
R20190 gnd.n6441 gnd.n6440 0.152939
R20191 gnd.n6441 gnd.n552 0.152939
R20192 gnd.n6449 gnd.n552 0.152939
R20193 gnd.n6450 gnd.n6449 0.152939
R20194 gnd.n6451 gnd.n6450 0.152939
R20195 gnd.n6451 gnd.n546 0.152939
R20196 gnd.n6459 gnd.n546 0.152939
R20197 gnd.n6460 gnd.n6459 0.152939
R20198 gnd.n6461 gnd.n6460 0.152939
R20199 gnd.n6461 gnd.n540 0.152939
R20200 gnd.n6469 gnd.n540 0.152939
R20201 gnd.n6470 gnd.n6469 0.152939
R20202 gnd.n6471 gnd.n6470 0.152939
R20203 gnd.n6471 gnd.n534 0.152939
R20204 gnd.n6479 gnd.n534 0.152939
R20205 gnd.n6480 gnd.n6479 0.152939
R20206 gnd.n6481 gnd.n6480 0.152939
R20207 gnd.n6481 gnd.n528 0.152939
R20208 gnd.n6489 gnd.n528 0.152939
R20209 gnd.n6490 gnd.n6489 0.152939
R20210 gnd.n6492 gnd.n6490 0.152939
R20211 gnd.n6492 gnd.n6491 0.152939
R20212 gnd.n6491 gnd.n522 0.152939
R20213 gnd.n6501 gnd.n522 0.152939
R20214 gnd.n6502 gnd.n517 0.152939
R20215 gnd.n6510 gnd.n517 0.152939
R20216 gnd.n6511 gnd.n6510 0.152939
R20217 gnd.n6512 gnd.n6511 0.152939
R20218 gnd.n6512 gnd.n511 0.152939
R20219 gnd.n6520 gnd.n511 0.152939
R20220 gnd.n6521 gnd.n6520 0.152939
R20221 gnd.n6522 gnd.n6521 0.152939
R20222 gnd.n6522 gnd.n505 0.152939
R20223 gnd.n6530 gnd.n505 0.152939
R20224 gnd.n6531 gnd.n6530 0.152939
R20225 gnd.n6532 gnd.n6531 0.152939
R20226 gnd.n6532 gnd.n499 0.152939
R20227 gnd.n6540 gnd.n499 0.152939
R20228 gnd.n6541 gnd.n6540 0.152939
R20229 gnd.n6542 gnd.n6541 0.152939
R20230 gnd.n6542 gnd.n493 0.152939
R20231 gnd.n6550 gnd.n493 0.152939
R20232 gnd.n6551 gnd.n6550 0.152939
R20233 gnd.n6552 gnd.n6551 0.152939
R20234 gnd.n6552 gnd.n487 0.152939
R20235 gnd.n6560 gnd.n487 0.152939
R20236 gnd.n6561 gnd.n6560 0.152939
R20237 gnd.n6562 gnd.n6561 0.152939
R20238 gnd.n6562 gnd.n481 0.152939
R20239 gnd.n6570 gnd.n481 0.152939
R20240 gnd.n6571 gnd.n6570 0.152939
R20241 gnd.n6572 gnd.n6571 0.152939
R20242 gnd.n6572 gnd.n475 0.152939
R20243 gnd.n6580 gnd.n475 0.152939
R20244 gnd.n6581 gnd.n6580 0.152939
R20245 gnd.n6582 gnd.n6581 0.152939
R20246 gnd.n6582 gnd.n469 0.152939
R20247 gnd.n6590 gnd.n469 0.152939
R20248 gnd.n6591 gnd.n6590 0.152939
R20249 gnd.n6592 gnd.n6591 0.152939
R20250 gnd.n6592 gnd.n463 0.152939
R20251 gnd.n6600 gnd.n463 0.152939
R20252 gnd.n6601 gnd.n6600 0.152939
R20253 gnd.n6602 gnd.n6601 0.152939
R20254 gnd.n6602 gnd.n457 0.152939
R20255 gnd.n6610 gnd.n457 0.152939
R20256 gnd.n6611 gnd.n6610 0.152939
R20257 gnd.n6612 gnd.n6611 0.152939
R20258 gnd.n6612 gnd.n451 0.152939
R20259 gnd.n6620 gnd.n451 0.152939
R20260 gnd.n6621 gnd.n6620 0.152939
R20261 gnd.n6622 gnd.n6621 0.152939
R20262 gnd.n6622 gnd.n445 0.152939
R20263 gnd.n6630 gnd.n445 0.152939
R20264 gnd.n6631 gnd.n6630 0.152939
R20265 gnd.n6632 gnd.n6631 0.152939
R20266 gnd.n6632 gnd.n439 0.152939
R20267 gnd.n6640 gnd.n439 0.152939
R20268 gnd.n6641 gnd.n6640 0.152939
R20269 gnd.n6642 gnd.n6641 0.152939
R20270 gnd.n6642 gnd.n433 0.152939
R20271 gnd.n6650 gnd.n433 0.152939
R20272 gnd.n6651 gnd.n6650 0.152939
R20273 gnd.n6652 gnd.n6651 0.152939
R20274 gnd.n6652 gnd.n427 0.152939
R20275 gnd.n6660 gnd.n427 0.152939
R20276 gnd.n6661 gnd.n6660 0.152939
R20277 gnd.n6662 gnd.n6661 0.152939
R20278 gnd.n6662 gnd.n421 0.152939
R20279 gnd.n6670 gnd.n421 0.152939
R20280 gnd.n6671 gnd.n6670 0.152939
R20281 gnd.n6672 gnd.n6671 0.152939
R20282 gnd.n6672 gnd.n415 0.152939
R20283 gnd.n6680 gnd.n415 0.152939
R20284 gnd.n6681 gnd.n6680 0.152939
R20285 gnd.n6682 gnd.n6681 0.152939
R20286 gnd.n6682 gnd.n409 0.152939
R20287 gnd.n6690 gnd.n409 0.152939
R20288 gnd.n6691 gnd.n6690 0.152939
R20289 gnd.n6692 gnd.n6691 0.152939
R20290 gnd.n6692 gnd.n403 0.152939
R20291 gnd.n6700 gnd.n403 0.152939
R20292 gnd.n6701 gnd.n6700 0.152939
R20293 gnd.n6702 gnd.n6701 0.152939
R20294 gnd.n6702 gnd.n397 0.152939
R20295 gnd.n6711 gnd.n397 0.152939
R20296 gnd.n6712 gnd.n6711 0.152939
R20297 gnd.n6713 gnd.n6712 0.152939
R20298 gnd.n4302 gnd.n4298 0.152939
R20299 gnd.n4303 gnd.n4302 0.152939
R20300 gnd.n4304 gnd.n4303 0.152939
R20301 gnd.n4304 gnd.n2066 0.152939
R20302 gnd.n4310 gnd.n2066 0.152939
R20303 gnd.n4311 gnd.n4310 0.152939
R20304 gnd.n4312 gnd.n4311 0.152939
R20305 gnd.n4313 gnd.n4312 0.152939
R20306 gnd.n4314 gnd.n4313 0.152939
R20307 gnd.n4317 gnd.n4314 0.152939
R20308 gnd.n4318 gnd.n4317 0.152939
R20309 gnd.n4319 gnd.n4318 0.152939
R20310 gnd.n4320 gnd.n4319 0.152939
R20311 gnd.n4322 gnd.n4320 0.152939
R20312 gnd.n4324 gnd.n4322 0.152939
R20313 gnd.n4324 gnd.n4323 0.152939
R20314 gnd.n4323 gnd.n1856 0.152939
R20315 gnd.n1857 gnd.n1856 0.152939
R20316 gnd.n1858 gnd.n1857 0.152939
R20317 gnd.n1860 gnd.n1858 0.152939
R20318 gnd.n1861 gnd.n1860 0.152939
R20319 gnd.n1861 gnd.n1837 0.152939
R20320 gnd.n4483 gnd.n1837 0.152939
R20321 gnd.n4484 gnd.n4483 0.152939
R20322 gnd.n4485 gnd.n4484 0.152939
R20323 gnd.n4485 gnd.n1824 0.152939
R20324 gnd.n4499 gnd.n1824 0.152939
R20325 gnd.n4500 gnd.n4499 0.152939
R20326 gnd.n4501 gnd.n4500 0.152939
R20327 gnd.n4501 gnd.n1808 0.152939
R20328 gnd.n4533 gnd.n1808 0.152939
R20329 gnd.n4534 gnd.n4533 0.152939
R20330 gnd.n4535 gnd.n4534 0.152939
R20331 gnd.n4536 gnd.n4535 0.152939
R20332 gnd.n4537 gnd.n4536 0.152939
R20333 gnd.n4539 gnd.n4537 0.152939
R20334 gnd.n4539 gnd.n4538 0.152939
R20335 gnd.n4538 gnd.n1119 0.152939
R20336 gnd.n1120 gnd.n1119 0.152939
R20337 gnd.n1121 gnd.n1120 0.152939
R20338 gnd.n1712 gnd.n1121 0.152939
R20339 gnd.n4653 gnd.n1712 0.152939
R20340 gnd.n4654 gnd.n4653 0.152939
R20341 gnd.n4655 gnd.n4654 0.152939
R20342 gnd.n4656 gnd.n4655 0.152939
R20343 gnd.n4657 gnd.n4656 0.152939
R20344 gnd.n4657 gnd.n1687 0.152939
R20345 gnd.n4693 gnd.n1687 0.152939
R20346 gnd.n4694 gnd.n4693 0.152939
R20347 gnd.n4695 gnd.n4694 0.152939
R20348 gnd.n4696 gnd.n4695 0.152939
R20349 gnd.n4696 gnd.n1659 0.152939
R20350 gnd.n4729 gnd.n1659 0.152939
R20351 gnd.n4730 gnd.n4729 0.152939
R20352 gnd.n4731 gnd.n4730 0.152939
R20353 gnd.n4731 gnd.n1641 0.152939
R20354 gnd.n4755 gnd.n1641 0.152939
R20355 gnd.n4756 gnd.n4755 0.152939
R20356 gnd.n4757 gnd.n4756 0.152939
R20357 gnd.n4758 gnd.n4757 0.152939
R20358 gnd.n4758 gnd.n1615 0.152939
R20359 gnd.n4811 gnd.n1615 0.152939
R20360 gnd.n4812 gnd.n4811 0.152939
R20361 gnd.n4813 gnd.n4812 0.152939
R20362 gnd.n4814 gnd.n4813 0.152939
R20363 gnd.n4814 gnd.n1590 0.152939
R20364 gnd.n4851 gnd.n1590 0.152939
R20365 gnd.n4852 gnd.n4851 0.152939
R20366 gnd.n4853 gnd.n4852 0.152939
R20367 gnd.n4854 gnd.n4853 0.152939
R20368 gnd.n4854 gnd.n1560 0.152939
R20369 gnd.n4920 gnd.n1560 0.152939
R20370 gnd.n4921 gnd.n4920 0.152939
R20371 gnd.n4922 gnd.n4921 0.152939
R20372 gnd.n4923 gnd.n4922 0.152939
R20373 gnd.n4923 gnd.n1536 0.152939
R20374 gnd.n4953 gnd.n1536 0.152939
R20375 gnd.n4954 gnd.n4953 0.152939
R20376 gnd.n4955 gnd.n4954 0.152939
R20377 gnd.n4956 gnd.n4955 0.152939
R20378 gnd.n4956 gnd.n1515 0.152939
R20379 gnd.n5007 gnd.n1515 0.152939
R20380 gnd.n5008 gnd.n5007 0.152939
R20381 gnd.n5009 gnd.n5008 0.152939
R20382 gnd.n5010 gnd.n5009 0.152939
R20383 gnd.n5010 gnd.n1490 0.152939
R20384 gnd.n5044 gnd.n1490 0.152939
R20385 gnd.n5045 gnd.n5044 0.152939
R20386 gnd.n5046 gnd.n5045 0.152939
R20387 gnd.n5046 gnd.n1399 0.152939
R20388 gnd.n5187 gnd.n1399 0.152939
R20389 gnd.n5188 gnd.n5187 0.152939
R20390 gnd.n5189 gnd.n5188 0.152939
R20391 gnd.n5189 gnd.n1386 0.152939
R20392 gnd.n5203 gnd.n1386 0.152939
R20393 gnd.n5204 gnd.n5203 0.152939
R20394 gnd.n5205 gnd.n5204 0.152939
R20395 gnd.n5205 gnd.n1373 0.152939
R20396 gnd.n5219 gnd.n1373 0.152939
R20397 gnd.n5220 gnd.n5219 0.152939
R20398 gnd.n5221 gnd.n5220 0.152939
R20399 gnd.n5221 gnd.n1360 0.152939
R20400 gnd.n5235 gnd.n1360 0.152939
R20401 gnd.n5236 gnd.n5235 0.152939
R20402 gnd.n5238 gnd.n5236 0.152939
R20403 gnd.n5238 gnd.n5237 0.152939
R20404 gnd.n5237 gnd.n1235 0.152939
R20405 gnd.n1236 gnd.n1235 0.152939
R20406 gnd.n1237 gnd.n1236 0.152939
R20407 gnd.n5278 gnd.n1237 0.152939
R20408 gnd.n5279 gnd.n5278 0.152939
R20409 gnd.n5280 gnd.n5279 0.152939
R20410 gnd.n5281 gnd.n5280 0.152939
R20411 gnd.n5282 gnd.n5281 0.152939
R20412 gnd.n5389 gnd.n5282 0.152939
R20413 gnd.n5392 gnd.n5389 0.152939
R20414 gnd.n5393 gnd.n5392 0.152939
R20415 gnd.n5394 gnd.n5393 0.152939
R20416 gnd.n5395 gnd.n5394 0.152939
R20417 gnd.n5395 gnd.n5340 0.152939
R20418 gnd.n5430 gnd.n5340 0.152939
R20419 gnd.n5431 gnd.n5430 0.152939
R20420 gnd.n5432 gnd.n5431 0.152939
R20421 gnd.n5434 gnd.n5432 0.152939
R20422 gnd.n5434 gnd.n5433 0.152939
R20423 gnd.n5433 gnd.n392 0.152939
R20424 gnd.n393 gnd.n392 0.152939
R20425 gnd.n394 gnd.n393 0.152939
R20426 gnd.n6179 gnd.n714 0.152939
R20427 gnd.n719 gnd.n714 0.152939
R20428 gnd.n720 gnd.n719 0.152939
R20429 gnd.n721 gnd.n720 0.152939
R20430 gnd.n726 gnd.n721 0.152939
R20431 gnd.n727 gnd.n726 0.152939
R20432 gnd.n728 gnd.n727 0.152939
R20433 gnd.n729 gnd.n728 0.152939
R20434 gnd.n734 gnd.n729 0.152939
R20435 gnd.n735 gnd.n734 0.152939
R20436 gnd.n736 gnd.n735 0.152939
R20437 gnd.n737 gnd.n736 0.152939
R20438 gnd.n742 gnd.n737 0.152939
R20439 gnd.n743 gnd.n742 0.152939
R20440 gnd.n744 gnd.n743 0.152939
R20441 gnd.n745 gnd.n744 0.152939
R20442 gnd.n750 gnd.n745 0.152939
R20443 gnd.n751 gnd.n750 0.152939
R20444 gnd.n752 gnd.n751 0.152939
R20445 gnd.n753 gnd.n752 0.152939
R20446 gnd.n758 gnd.n753 0.152939
R20447 gnd.n759 gnd.n758 0.152939
R20448 gnd.n760 gnd.n759 0.152939
R20449 gnd.n761 gnd.n760 0.152939
R20450 gnd.n766 gnd.n761 0.152939
R20451 gnd.n767 gnd.n766 0.152939
R20452 gnd.n768 gnd.n767 0.152939
R20453 gnd.n769 gnd.n768 0.152939
R20454 gnd.n774 gnd.n769 0.152939
R20455 gnd.n775 gnd.n774 0.152939
R20456 gnd.n776 gnd.n775 0.152939
R20457 gnd.n777 gnd.n776 0.152939
R20458 gnd.n782 gnd.n777 0.152939
R20459 gnd.n783 gnd.n782 0.152939
R20460 gnd.n784 gnd.n783 0.152939
R20461 gnd.n785 gnd.n784 0.152939
R20462 gnd.n790 gnd.n785 0.152939
R20463 gnd.n791 gnd.n790 0.152939
R20464 gnd.n792 gnd.n791 0.152939
R20465 gnd.n793 gnd.n792 0.152939
R20466 gnd.n798 gnd.n793 0.152939
R20467 gnd.n799 gnd.n798 0.152939
R20468 gnd.n800 gnd.n799 0.152939
R20469 gnd.n801 gnd.n800 0.152939
R20470 gnd.n806 gnd.n801 0.152939
R20471 gnd.n807 gnd.n806 0.152939
R20472 gnd.n808 gnd.n807 0.152939
R20473 gnd.n809 gnd.n808 0.152939
R20474 gnd.n814 gnd.n809 0.152939
R20475 gnd.n815 gnd.n814 0.152939
R20476 gnd.n816 gnd.n815 0.152939
R20477 gnd.n817 gnd.n816 0.152939
R20478 gnd.n822 gnd.n817 0.152939
R20479 gnd.n823 gnd.n822 0.152939
R20480 gnd.n824 gnd.n823 0.152939
R20481 gnd.n825 gnd.n824 0.152939
R20482 gnd.n830 gnd.n825 0.152939
R20483 gnd.n831 gnd.n830 0.152939
R20484 gnd.n832 gnd.n831 0.152939
R20485 gnd.n833 gnd.n832 0.152939
R20486 gnd.n838 gnd.n833 0.152939
R20487 gnd.n839 gnd.n838 0.152939
R20488 gnd.n840 gnd.n839 0.152939
R20489 gnd.n841 gnd.n840 0.152939
R20490 gnd.n846 gnd.n841 0.152939
R20491 gnd.n847 gnd.n846 0.152939
R20492 gnd.n848 gnd.n847 0.152939
R20493 gnd.n849 gnd.n848 0.152939
R20494 gnd.n854 gnd.n849 0.152939
R20495 gnd.n855 gnd.n854 0.152939
R20496 gnd.n856 gnd.n855 0.152939
R20497 gnd.n857 gnd.n856 0.152939
R20498 gnd.n862 gnd.n857 0.152939
R20499 gnd.n863 gnd.n862 0.152939
R20500 gnd.n864 gnd.n863 0.152939
R20501 gnd.n865 gnd.n864 0.152939
R20502 gnd.n870 gnd.n865 0.152939
R20503 gnd.n871 gnd.n870 0.152939
R20504 gnd.n872 gnd.n871 0.152939
R20505 gnd.n873 gnd.n872 0.152939
R20506 gnd.n878 gnd.n873 0.152939
R20507 gnd.n879 gnd.n878 0.152939
R20508 gnd.n880 gnd.n879 0.152939
R20509 gnd.n881 gnd.n880 0.152939
R20510 gnd.n4477 gnd.n1831 0.152939
R20511 gnd.n4491 gnd.n1831 0.152939
R20512 gnd.n4492 gnd.n4491 0.152939
R20513 gnd.n4493 gnd.n4492 0.152939
R20514 gnd.n4493 gnd.n1817 0.152939
R20515 gnd.n4507 gnd.n1817 0.152939
R20516 gnd.n4508 gnd.n4507 0.152939
R20517 gnd.n4527 gnd.n4508 0.152939
R20518 gnd.n4527 gnd.n4526 0.152939
R20519 gnd.n4526 gnd.n4525 0.152939
R20520 gnd.n4525 gnd.n4509 0.152939
R20521 gnd.n4521 gnd.n4509 0.152939
R20522 gnd.n4521 gnd.n4520 0.152939
R20523 gnd.n4520 gnd.n4519 0.152939
R20524 gnd.n4519 gnd.n4514 0.152939
R20525 gnd.n4514 gnd.n1131 0.152939
R20526 gnd.n5816 gnd.n1131 0.152939
R20527 gnd.n5816 gnd.n5815 0.152939
R20528 gnd.n5815 gnd.n5814 0.152939
R20529 gnd.n5814 gnd.n1132 0.152939
R20530 gnd.n5810 gnd.n1132 0.152939
R20531 gnd.n5810 gnd.n5809 0.152939
R20532 gnd.n5809 gnd.n5808 0.152939
R20533 gnd.n5808 gnd.n1137 0.152939
R20534 gnd.n5804 gnd.n1137 0.152939
R20535 gnd.n5804 gnd.n5803 0.152939
R20536 gnd.n5803 gnd.n5802 0.152939
R20537 gnd.n5802 gnd.n1142 0.152939
R20538 gnd.n5798 gnd.n1142 0.152939
R20539 gnd.n5798 gnd.n5797 0.152939
R20540 gnd.n5797 gnd.n5796 0.152939
R20541 gnd.n5796 gnd.n1147 0.152939
R20542 gnd.n5792 gnd.n1147 0.152939
R20543 gnd.n5792 gnd.n5791 0.152939
R20544 gnd.n5791 gnd.n5790 0.152939
R20545 gnd.n5790 gnd.n1152 0.152939
R20546 gnd.n5786 gnd.n1152 0.152939
R20547 gnd.n5786 gnd.n5785 0.152939
R20548 gnd.n5785 gnd.n5784 0.152939
R20549 gnd.n5784 gnd.n1157 0.152939
R20550 gnd.n5780 gnd.n1157 0.152939
R20551 gnd.n5780 gnd.n5779 0.152939
R20552 gnd.n5779 gnd.n5778 0.152939
R20553 gnd.n5778 gnd.n1162 0.152939
R20554 gnd.n5774 gnd.n1162 0.152939
R20555 gnd.n5774 gnd.n5773 0.152939
R20556 gnd.n5773 gnd.n5772 0.152939
R20557 gnd.n5772 gnd.n1167 0.152939
R20558 gnd.n5768 gnd.n1167 0.152939
R20559 gnd.n5768 gnd.n5767 0.152939
R20560 gnd.n5767 gnd.n5766 0.152939
R20561 gnd.n5766 gnd.n1172 0.152939
R20562 gnd.n5762 gnd.n1172 0.152939
R20563 gnd.n5762 gnd.n5761 0.152939
R20564 gnd.n5761 gnd.n5760 0.152939
R20565 gnd.n5760 gnd.n1177 0.152939
R20566 gnd.n5756 gnd.n1177 0.152939
R20567 gnd.n5756 gnd.n5755 0.152939
R20568 gnd.n5755 gnd.n5754 0.152939
R20569 gnd.n5754 gnd.n1182 0.152939
R20570 gnd.n5750 gnd.n1182 0.152939
R20571 gnd.n5750 gnd.n5749 0.152939
R20572 gnd.n5749 gnd.n5748 0.152939
R20573 gnd.n5748 gnd.n1187 0.152939
R20574 gnd.n5744 gnd.n1187 0.152939
R20575 gnd.n5744 gnd.n5743 0.152939
R20576 gnd.n5743 gnd.n5742 0.152939
R20577 gnd.n5742 gnd.n1192 0.152939
R20578 gnd.n5738 gnd.n1192 0.152939
R20579 gnd.n5738 gnd.n5737 0.152939
R20580 gnd.n5737 gnd.n5736 0.152939
R20581 gnd.n5736 gnd.n1197 0.152939
R20582 gnd.n5732 gnd.n1197 0.152939
R20583 gnd.n5732 gnd.n5731 0.152939
R20584 gnd.n5731 gnd.n5730 0.152939
R20585 gnd.n5730 gnd.n1202 0.152939
R20586 gnd.n5726 gnd.n1202 0.152939
R20587 gnd.n5726 gnd.n5725 0.152939
R20588 gnd.n5725 gnd.n5724 0.152939
R20589 gnd.n5724 gnd.n1207 0.152939
R20590 gnd.n5720 gnd.n1207 0.152939
R20591 gnd.n5720 gnd.n5719 0.152939
R20592 gnd.n4215 gnd.n4214 0.152939
R20593 gnd.n4214 gnd.n4213 0.152939
R20594 gnd.n4213 gnd.n4202 0.152939
R20595 gnd.n4209 gnd.n4202 0.152939
R20596 gnd.n4209 gnd.n4208 0.152939
R20597 gnd.n4208 gnd.n4207 0.152939
R20598 gnd.n4207 gnd.n2076 0.152939
R20599 gnd.n4269 gnd.n2076 0.152939
R20600 gnd.n4270 gnd.n4269 0.152939
R20601 gnd.n4271 gnd.n4270 0.152939
R20602 gnd.n4271 gnd.n2071 0.152939
R20603 gnd.n4291 gnd.n2071 0.152939
R20604 gnd.n4291 gnd.n4290 0.152939
R20605 gnd.n4290 gnd.n4289 0.152939
R20606 gnd.n4289 gnd.n2072 0.152939
R20607 gnd.n4285 gnd.n2072 0.152939
R20608 gnd.n4285 gnd.n2059 0.152939
R20609 gnd.n4350 gnd.n2059 0.152939
R20610 gnd.n4351 gnd.n4350 0.152939
R20611 gnd.n4352 gnd.n4351 0.152939
R20612 gnd.n4352 gnd.n2054 0.152939
R20613 gnd.n4365 gnd.n2054 0.152939
R20614 gnd.n4366 gnd.n4365 0.152939
R20615 gnd.n4369 gnd.n4366 0.152939
R20616 gnd.n4369 gnd.n4368 0.152939
R20617 gnd.n4368 gnd.n4367 0.152939
R20618 gnd.n1946 gnd.n1945 0.152939
R20619 gnd.n1947 gnd.n1946 0.152939
R20620 gnd.n1947 gnd.n1917 0.152939
R20621 gnd.n1953 gnd.n1917 0.152939
R20622 gnd.n1954 gnd.n1953 0.152939
R20623 gnd.n4380 gnd.n1954 0.152939
R20624 gnd.n1942 gnd.n1921 0.152939
R20625 gnd.n1938 gnd.n1921 0.152939
R20626 gnd.n1938 gnd.n1937 0.152939
R20627 gnd.n1937 gnd.n1936 0.152939
R20628 gnd.n1936 gnd.n1925 0.152939
R20629 gnd.n1932 gnd.n1925 0.152939
R20630 gnd.n1932 gnd.n1931 0.152939
R20631 gnd.n1931 gnd.n1930 0.152939
R20632 gnd.n1930 gnd.n1800 0.152939
R20633 gnd.n4550 gnd.n1800 0.152939
R20634 gnd.n4551 gnd.n4550 0.152939
R20635 gnd.n4552 gnd.n4551 0.152939
R20636 gnd.n4552 gnd.n1796 0.152939
R20637 gnd.n4558 gnd.n1796 0.152939
R20638 gnd.n4559 gnd.n4558 0.152939
R20639 gnd.n4618 gnd.n4559 0.152939
R20640 gnd.n4618 gnd.n4617 0.152939
R20641 gnd.n4617 gnd.n4616 0.152939
R20642 gnd.n4616 gnd.n4560 0.152939
R20643 gnd.n4612 gnd.n4560 0.152939
R20644 gnd.n4612 gnd.n4611 0.152939
R20645 gnd.n4611 gnd.n4610 0.152939
R20646 gnd.n4610 gnd.n4566 0.152939
R20647 gnd.n4606 gnd.n4566 0.152939
R20648 gnd.n4606 gnd.n4605 0.152939
R20649 gnd.n4605 gnd.n4604 0.152939
R20650 gnd.n4604 gnd.n4570 0.152939
R20651 gnd.n4600 gnd.n4570 0.152939
R20652 gnd.n4600 gnd.n4599 0.152939
R20653 gnd.n4599 gnd.n4598 0.152939
R20654 gnd.n4598 gnd.n4575 0.152939
R20655 gnd.n4594 gnd.n4575 0.152939
R20656 gnd.n4594 gnd.n4593 0.152939
R20657 gnd.n4593 gnd.n4592 0.152939
R20658 gnd.n4592 gnd.n4579 0.152939
R20659 gnd.n4588 gnd.n4579 0.152939
R20660 gnd.n4588 gnd.n4587 0.152939
R20661 gnd.n4587 gnd.n4586 0.152939
R20662 gnd.n4586 gnd.n4583 0.152939
R20663 gnd.n4583 gnd.n1605 0.152939
R20664 gnd.n4821 gnd.n1605 0.152939
R20665 gnd.n4822 gnd.n4821 0.152939
R20666 gnd.n4837 gnd.n4822 0.152939
R20667 gnd.n4837 gnd.n4836 0.152939
R20668 gnd.n4836 gnd.n4835 0.152939
R20669 gnd.n4835 gnd.n4823 0.152939
R20670 gnd.n4831 gnd.n4823 0.152939
R20671 gnd.n4831 gnd.n4830 0.152939
R20672 gnd.n4830 gnd.n4829 0.152939
R20673 gnd.n4829 gnd.n1552 0.152939
R20674 gnd.n4930 gnd.n1552 0.152939
R20675 gnd.n4931 gnd.n4930 0.152939
R20676 gnd.n4933 gnd.n4931 0.152939
R20677 gnd.n4933 gnd.n4932 0.152939
R20678 gnd.n4932 gnd.n1529 0.152939
R20679 gnd.n4963 gnd.n1529 0.152939
R20680 gnd.n4964 gnd.n4963 0.152939
R20681 gnd.n4992 gnd.n4964 0.152939
R20682 gnd.n4992 gnd.n4991 0.152939
R20683 gnd.n4991 gnd.n4990 0.152939
R20684 gnd.n4990 gnd.n4965 0.152939
R20685 gnd.n4986 gnd.n4965 0.152939
R20686 gnd.n4986 gnd.n4985 0.152939
R20687 gnd.n4985 gnd.n4984 0.152939
R20688 gnd.n4984 gnd.n4973 0.152939
R20689 gnd.n4980 gnd.n4973 0.152939
R20690 gnd.n4980 gnd.n4979 0.152939
R20691 gnd.n4979 gnd.n4978 0.152939
R20692 gnd.n4978 gnd.n1391 0.152939
R20693 gnd.n5195 gnd.n1391 0.152939
R20694 gnd.n5196 gnd.n5195 0.152939
R20695 gnd.n5197 gnd.n5196 0.152939
R20696 gnd.n5197 gnd.n1378 0.152939
R20697 gnd.n5211 gnd.n1378 0.152939
R20698 gnd.n5212 gnd.n5211 0.152939
R20699 gnd.n5213 gnd.n5212 0.152939
R20700 gnd.n5213 gnd.n1366 0.152939
R20701 gnd.n5227 gnd.n1366 0.152939
R20702 gnd.n5228 gnd.n5227 0.152939
R20703 gnd.n5229 gnd.n5228 0.152939
R20704 gnd.n5229 gnd.n1353 0.152939
R20705 gnd.n5244 gnd.n1353 0.152939
R20706 gnd.n5246 gnd.n5245 0.152939
R20707 gnd.n5246 gnd.n1351 0.152939
R20708 gnd.n5254 gnd.n1351 0.152939
R20709 gnd.n5255 gnd.n5254 0.152939
R20710 gnd.n5256 gnd.n5255 0.152939
R20711 gnd.n5256 gnd.n1348 0.152939
R20712 gnd.n5369 gnd.n5368 0.152939
R20713 gnd.n5375 gnd.n5368 0.152939
R20714 gnd.n5376 gnd.n5375 0.152939
R20715 gnd.n5377 gnd.n5376 0.152939
R20716 gnd.n5377 gnd.n5351 0.152939
R20717 gnd.n5403 gnd.n5351 0.152939
R20718 gnd.n5404 gnd.n5403 0.152939
R20719 gnd.n5405 gnd.n5404 0.152939
R20720 gnd.n5405 gnd.n5346 0.152939
R20721 gnd.n5423 gnd.n5346 0.152939
R20722 gnd.n5423 gnd.n5422 0.152939
R20723 gnd.n5422 gnd.n5421 0.152939
R20724 gnd.n5421 gnd.n5347 0.152939
R20725 gnd.n5347 gnd.n367 0.152939
R20726 gnd.n6748 gnd.n367 0.152939
R20727 gnd.n6749 gnd.n6748 0.152939
R20728 gnd.n6751 gnd.n6749 0.152939
R20729 gnd.n6751 gnd.n6750 0.152939
R20730 gnd.n6750 gnd.n340 0.152939
R20731 gnd.n6782 gnd.n340 0.152939
R20732 gnd.n6783 gnd.n6782 0.152939
R20733 gnd.n6790 gnd.n6783 0.152939
R20734 gnd.n6790 gnd.n6789 0.152939
R20735 gnd.n6789 gnd.n6788 0.152939
R20736 gnd.n6788 gnd.n6784 0.152939
R20737 gnd.n6784 gnd.n79 0.152939
R20738 gnd.n4380 gnd.n4379 0.128549
R20739 gnd.n5591 gnd.n1348 0.128549
R20740 gnd.n6775 gnd.n326 0.0785577
R20741 gnd.n112 gnd.n111 0.0785577
R20742 gnd.n4259 gnd.n2083 0.0785577
R20743 gnd.n4157 gnd.n2129 0.0785577
R20744 gnd.n3123 gnd.n3122 0.0767195
R20745 gnd.n3122 gnd.n3121 0.0767195
R20746 gnd.n7196 gnd.n7195 0.0695946
R20747 gnd.n4201 gnd.n4200 0.0695946
R20748 gnd.n4215 gnd.n4201 0.0695946
R20749 gnd.n7196 gnd.n79 0.0695946
R20750 gnd.n4379 gnd.n4378 0.063
R20751 gnd.n5592 gnd.n5591 0.063
R20752 gnd.n5592 gnd.n1347 0.0477147
R20753 gnd.n6991 gnd.n6990 0.0477147
R20754 gnd.n3689 gnd.n2288 0.0477147
R20755 gnd.n3921 gnd.n2244 0.0477147
R20756 gnd.n4378 gnd.n4377 0.0477147
R20757 gnd.n2886 gnd.n2774 0.0442063
R20758 gnd.n2887 gnd.n2886 0.0442063
R20759 gnd.n2888 gnd.n2887 0.0442063
R20760 gnd.n2888 gnd.n2763 0.0442063
R20761 gnd.n2902 gnd.n2763 0.0442063
R20762 gnd.n2903 gnd.n2902 0.0442063
R20763 gnd.n2904 gnd.n2903 0.0442063
R20764 gnd.n2904 gnd.n2750 0.0442063
R20765 gnd.n2948 gnd.n2750 0.0442063
R20766 gnd.n2949 gnd.n2948 0.0442063
R20767 gnd.n5360 gnd.n1347 0.0344674
R20768 gnd.n5360 gnd.n5354 0.0344674
R20769 gnd.n5365 gnd.n5354 0.0344674
R20770 gnd.n5366 gnd.n5365 0.0344674
R20771 gnd.n5366 gnd.n5312 0.0344674
R20772 gnd.n5313 gnd.n5312 0.0344674
R20773 gnd.n5314 gnd.n5313 0.0344674
R20774 gnd.n5349 gnd.n5314 0.0344674
R20775 gnd.n5349 gnd.n5331 0.0344674
R20776 gnd.n5332 gnd.n5331 0.0344674
R20777 gnd.n5333 gnd.n5332 0.0344674
R20778 gnd.n5414 gnd.n5333 0.0344674
R20779 gnd.n5414 gnd.n386 0.0344674
R20780 gnd.n387 gnd.n386 0.0344674
R20781 gnd.n6726 gnd.n387 0.0344674
R20782 gnd.n6727 gnd.n6726 0.0344674
R20783 gnd.n6727 gnd.n361 0.0344674
R20784 gnd.n361 gnd.n358 0.0344674
R20785 gnd.n359 gnd.n358 0.0344674
R20786 gnd.n6761 gnd.n359 0.0344674
R20787 gnd.n6762 gnd.n6761 0.0344674
R20788 gnd.n6762 gnd.n333 0.0344674
R20789 gnd.n6799 gnd.n333 0.0344674
R20790 gnd.n6799 gnd.n316 0.0344674
R20791 gnd.n6816 gnd.n316 0.0344674
R20792 gnd.n6817 gnd.n6816 0.0344674
R20793 gnd.n6817 gnd.n310 0.0344674
R20794 gnd.n6825 gnd.n310 0.0344674
R20795 gnd.n6826 gnd.n6825 0.0344674
R20796 gnd.n6826 gnd.n101 0.0344674
R20797 gnd.n102 gnd.n101 0.0344674
R20798 gnd.n103 gnd.n102 0.0344674
R20799 gnd.n6833 gnd.n103 0.0344674
R20800 gnd.n6833 gnd.n121 0.0344674
R20801 gnd.n122 gnd.n121 0.0344674
R20802 gnd.n123 gnd.n122 0.0344674
R20803 gnd.n6840 gnd.n123 0.0344674
R20804 gnd.n6840 gnd.n139 0.0344674
R20805 gnd.n140 gnd.n139 0.0344674
R20806 gnd.n141 gnd.n140 0.0344674
R20807 gnd.n6847 gnd.n141 0.0344674
R20808 gnd.n6847 gnd.n159 0.0344674
R20809 gnd.n160 gnd.n159 0.0344674
R20810 gnd.n161 gnd.n160 0.0344674
R20811 gnd.n6973 gnd.n161 0.0344674
R20812 gnd.n6973 gnd.n177 0.0344674
R20813 gnd.n178 gnd.n177 0.0344674
R20814 gnd.n179 gnd.n178 0.0344674
R20815 gnd.n6980 gnd.n179 0.0344674
R20816 gnd.n6980 gnd.n197 0.0344674
R20817 gnd.n198 gnd.n197 0.0344674
R20818 gnd.n199 gnd.n198 0.0344674
R20819 gnd.n6990 gnd.n199 0.0344674
R20820 gnd.n2951 gnd.n2684 0.0344674
R20821 gnd.n2244 gnd.n2243 0.0344674
R20822 gnd.n4046 gnd.n2243 0.0344674
R20823 gnd.n4047 gnd.n4046 0.0344674
R20824 gnd.n4047 gnd.n2227 0.0344674
R20825 gnd.n2227 gnd.n2225 0.0344674
R20826 gnd.n4066 gnd.n2225 0.0344674
R20827 gnd.n4067 gnd.n4066 0.0344674
R20828 gnd.n4067 gnd.n2209 0.0344674
R20829 gnd.n2209 gnd.n2207 0.0344674
R20830 gnd.n4086 gnd.n2207 0.0344674
R20831 gnd.n4087 gnd.n4086 0.0344674
R20832 gnd.n4087 gnd.n2191 0.0344674
R20833 gnd.n2191 gnd.n2188 0.0344674
R20834 gnd.n2189 gnd.n2188 0.0344674
R20835 gnd.n4108 gnd.n2189 0.0344674
R20836 gnd.n4109 gnd.n4108 0.0344674
R20837 gnd.n4109 gnd.n2165 0.0344674
R20838 gnd.n2165 gnd.n2162 0.0344674
R20839 gnd.n2163 gnd.n2162 0.0344674
R20840 gnd.n4143 gnd.n2163 0.0344674
R20841 gnd.n4144 gnd.n4143 0.0344674
R20842 gnd.n4144 gnd.n2140 0.0344674
R20843 gnd.n2140 gnd.n2137 0.0344674
R20844 gnd.n2138 gnd.n2137 0.0344674
R20845 gnd.n4178 gnd.n2138 0.0344674
R20846 gnd.n4179 gnd.n4178 0.0344674
R20847 gnd.n4179 gnd.n2114 0.0344674
R20848 gnd.n2114 gnd.n2112 0.0344674
R20849 gnd.n4223 gnd.n2112 0.0344674
R20850 gnd.n4224 gnd.n4223 0.0344674
R20851 gnd.n4224 gnd.n2097 0.0344674
R20852 gnd.n2097 gnd.n2093 0.0344674
R20853 gnd.n2094 gnd.n2093 0.0344674
R20854 gnd.n2095 gnd.n2094 0.0344674
R20855 gnd.n4247 gnd.n2095 0.0344674
R20856 gnd.n4248 gnd.n4247 0.0344674
R20857 gnd.n4248 gnd.n2074 0.0344674
R20858 gnd.n2074 gnd.n902 0.0344674
R20859 gnd.n903 gnd.n902 0.0344674
R20860 gnd.n904 gnd.n903 0.0344674
R20861 gnd.n4280 gnd.n904 0.0344674
R20862 gnd.n4280 gnd.n923 0.0344674
R20863 gnd.n924 gnd.n923 0.0344674
R20864 gnd.n925 gnd.n924 0.0344674
R20865 gnd.n4344 gnd.n925 0.0344674
R20866 gnd.n4344 gnd.n942 0.0344674
R20867 gnd.n943 gnd.n942 0.0344674
R20868 gnd.n944 gnd.n943 0.0344674
R20869 gnd.n4359 gnd.n944 0.0344674
R20870 gnd.n4359 gnd.n963 0.0344674
R20871 gnd.n964 gnd.n963 0.0344674
R20872 gnd.n965 gnd.n964 0.0344674
R20873 gnd.n4377 gnd.n965 0.0344674
R20874 gnd.n4386 gnd.n1913 0.0344674
R20875 gnd.n5590 gnd.n1349 0.0344674
R20876 gnd.n4473 gnd.n1844 0.029712
R20877 gnd.n5532 gnd.n1212 0.029712
R20878 gnd.n2971 gnd.n2970 0.0269946
R20879 gnd.n2973 gnd.n2972 0.0269946
R20880 gnd.n2679 gnd.n2677 0.0269946
R20881 gnd.n2983 gnd.n2981 0.0269946
R20882 gnd.n2982 gnd.n2658 0.0269946
R20883 gnd.n3002 gnd.n3001 0.0269946
R20884 gnd.n3004 gnd.n3003 0.0269946
R20885 gnd.n2653 gnd.n2652 0.0269946
R20886 gnd.n3014 gnd.n2648 0.0269946
R20887 gnd.n3013 gnd.n2650 0.0269946
R20888 gnd.n2649 gnd.n2631 0.0269946
R20889 gnd.n3034 gnd.n2632 0.0269946
R20890 gnd.n3033 gnd.n2633 0.0269946
R20891 gnd.n3067 gnd.n2608 0.0269946
R20892 gnd.n3069 gnd.n3068 0.0269946
R20893 gnd.n3070 gnd.n2555 0.0269946
R20894 gnd.n2603 gnd.n2556 0.0269946
R20895 gnd.n2605 gnd.n2557 0.0269946
R20896 gnd.n3080 gnd.n3079 0.0269946
R20897 gnd.n3082 gnd.n3081 0.0269946
R20898 gnd.n3083 gnd.n2577 0.0269946
R20899 gnd.n3085 gnd.n2578 0.0269946
R20900 gnd.n3088 gnd.n2579 0.0269946
R20901 gnd.n3091 gnd.n3090 0.0269946
R20902 gnd.n3093 gnd.n3092 0.0269946
R20903 gnd.n3158 gnd.n2462 0.0269946
R20904 gnd.n3160 gnd.n3159 0.0269946
R20905 gnd.n3169 gnd.n2455 0.0269946
R20906 gnd.n3171 gnd.n3170 0.0269946
R20907 gnd.n3172 gnd.n2453 0.0269946
R20908 gnd.n3179 gnd.n3175 0.0269946
R20909 gnd.n3178 gnd.n3177 0.0269946
R20910 gnd.n3176 gnd.n2432 0.0269946
R20911 gnd.n3201 gnd.n2433 0.0269946
R20912 gnd.n3200 gnd.n2434 0.0269946
R20913 gnd.n3243 gnd.n2407 0.0269946
R20914 gnd.n3245 gnd.n3244 0.0269946
R20915 gnd.n3254 gnd.n2400 0.0269946
R20916 gnd.n3256 gnd.n3255 0.0269946
R20917 gnd.n3257 gnd.n2398 0.0269946
R20918 gnd.n3264 gnd.n3260 0.0269946
R20919 gnd.n3263 gnd.n3262 0.0269946
R20920 gnd.n3261 gnd.n2377 0.0269946
R20921 gnd.n3286 gnd.n2378 0.0269946
R20922 gnd.n3285 gnd.n2379 0.0269946
R20923 gnd.n3332 gnd.n2353 0.0269946
R20924 gnd.n3334 gnd.n3333 0.0269946
R20925 gnd.n3343 gnd.n2346 0.0269946
R20926 gnd.n3602 gnd.n2344 0.0269946
R20927 gnd.n3607 gnd.n3605 0.0269946
R20928 gnd.n3606 gnd.n2325 0.0269946
R20929 gnd.n3631 gnd.n3630 0.0269946
R20930 gnd.n4387 gnd.n1912 0.0225788
R20931 gnd.n4392 gnd.n4391 0.0225788
R20932 gnd.n4397 gnd.n1908 0.0225788
R20933 gnd.n4398 gnd.n1904 0.0225788
R20934 gnd.n4404 gnd.n4403 0.0225788
R20935 gnd.n4409 gnd.n1902 0.0225788
R20936 gnd.n4410 gnd.n1900 0.0225788
R20937 gnd.n4416 gnd.n4415 0.0225788
R20938 gnd.n4421 gnd.n1896 0.0225788
R20939 gnd.n4422 gnd.n1892 0.0225788
R20940 gnd.n4428 gnd.n4427 0.0225788
R20941 gnd.n4433 gnd.n1890 0.0225788
R20942 gnd.n4434 gnd.n1888 0.0225788
R20943 gnd.n4440 gnd.n4439 0.0225788
R20944 gnd.n4446 gnd.n1884 0.0225788
R20945 gnd.n4447 gnd.n1880 0.0225788
R20946 gnd.n4454 gnd.n4452 0.0225788
R20947 gnd.n4453 gnd.n1847 0.0225788
R20948 gnd.n4473 gnd.n4472 0.0225788
R20949 gnd.n5586 gnd.n5266 0.0225788
R20950 gnd.n5585 gnd.n5267 0.0225788
R20951 gnd.n5582 gnd.n5581 0.0225788
R20952 gnd.n5578 gnd.n5482 0.0225788
R20953 gnd.n5577 gnd.n5486 0.0225788
R20954 gnd.n5574 gnd.n5573 0.0225788
R20955 gnd.n5570 gnd.n5492 0.0225788
R20956 gnd.n5569 gnd.n5498 0.0225788
R20957 gnd.n5566 gnd.n5565 0.0225788
R20958 gnd.n5562 gnd.n5502 0.0225788
R20959 gnd.n5561 gnd.n5506 0.0225788
R20960 gnd.n5558 gnd.n5557 0.0225788
R20961 gnd.n5554 gnd.n5512 0.0225788
R20962 gnd.n5553 gnd.n5518 0.0225788
R20963 gnd.n5550 gnd.n5549 0.0225788
R20964 gnd.n5546 gnd.n5522 0.0225788
R20965 gnd.n5545 gnd.n5528 0.0225788
R20966 gnd.n5539 gnd.n5538 0.0225788
R20967 gnd.n5533 gnd.n5532 0.0225788
R20968 gnd.n5718 gnd.n1212 0.0218415
R20969 gnd.n4476 gnd.n1844 0.0218415
R20970 gnd.n2951 gnd.n2950 0.0202011
R20971 gnd.n2950 gnd.n2949 0.0148637
R20972 gnd.n3600 gnd.n3344 0.0144266
R20973 gnd.n3601 gnd.n3600 0.0130679
R20974 gnd.n4387 gnd.n4386 0.0123886
R20975 gnd.n4391 gnd.n1912 0.0123886
R20976 gnd.n4392 gnd.n1908 0.0123886
R20977 gnd.n4398 gnd.n4397 0.0123886
R20978 gnd.n4403 gnd.n1904 0.0123886
R20979 gnd.n4404 gnd.n1902 0.0123886
R20980 gnd.n4410 gnd.n4409 0.0123886
R20981 gnd.n4415 gnd.n1900 0.0123886
R20982 gnd.n4416 gnd.n1896 0.0123886
R20983 gnd.n4422 gnd.n4421 0.0123886
R20984 gnd.n4427 gnd.n1892 0.0123886
R20985 gnd.n4428 gnd.n1890 0.0123886
R20986 gnd.n4434 gnd.n4433 0.0123886
R20987 gnd.n4439 gnd.n1888 0.0123886
R20988 gnd.n4440 gnd.n1884 0.0123886
R20989 gnd.n4447 gnd.n4446 0.0123886
R20990 gnd.n4452 gnd.n1880 0.0123886
R20991 gnd.n4454 gnd.n4453 0.0123886
R20992 gnd.n4472 gnd.n1847 0.0123886
R20993 gnd.n5266 gnd.n1349 0.0123886
R20994 gnd.n5586 gnd.n5585 0.0123886
R20995 gnd.n5582 gnd.n5267 0.0123886
R20996 gnd.n5581 gnd.n5482 0.0123886
R20997 gnd.n5578 gnd.n5577 0.0123886
R20998 gnd.n5574 gnd.n5486 0.0123886
R20999 gnd.n5573 gnd.n5492 0.0123886
R21000 gnd.n5570 gnd.n5569 0.0123886
R21001 gnd.n5566 gnd.n5498 0.0123886
R21002 gnd.n5565 gnd.n5502 0.0123886
R21003 gnd.n5562 gnd.n5561 0.0123886
R21004 gnd.n5558 gnd.n5506 0.0123886
R21005 gnd.n5557 gnd.n5512 0.0123886
R21006 gnd.n5554 gnd.n5553 0.0123886
R21007 gnd.n5550 gnd.n5518 0.0123886
R21008 gnd.n5549 gnd.n5522 0.0123886
R21009 gnd.n5546 gnd.n5545 0.0123886
R21010 gnd.n5539 gnd.n5528 0.0123886
R21011 gnd.n5538 gnd.n5533 0.0123886
R21012 gnd.n2970 gnd.n2684 0.00797283
R21013 gnd.n2972 gnd.n2971 0.00797283
R21014 gnd.n2973 gnd.n2679 0.00797283
R21015 gnd.n2981 gnd.n2677 0.00797283
R21016 gnd.n2983 gnd.n2982 0.00797283
R21017 gnd.n3001 gnd.n2658 0.00797283
R21018 gnd.n3003 gnd.n3002 0.00797283
R21019 gnd.n3004 gnd.n2653 0.00797283
R21020 gnd.n2652 gnd.n2648 0.00797283
R21021 gnd.n3014 gnd.n3013 0.00797283
R21022 gnd.n2650 gnd.n2649 0.00797283
R21023 gnd.n2632 gnd.n2631 0.00797283
R21024 gnd.n3034 gnd.n3033 0.00797283
R21025 gnd.n2633 gnd.n2608 0.00797283
R21026 gnd.n3068 gnd.n3067 0.00797283
R21027 gnd.n3070 gnd.n3069 0.00797283
R21028 gnd.n2603 gnd.n2555 0.00797283
R21029 gnd.n2605 gnd.n2556 0.00797283
R21030 gnd.n3079 gnd.n2557 0.00797283
R21031 gnd.n3081 gnd.n3080 0.00797283
R21032 gnd.n3083 gnd.n3082 0.00797283
R21033 gnd.n3085 gnd.n2577 0.00797283
R21034 gnd.n3088 gnd.n2578 0.00797283
R21035 gnd.n3090 gnd.n2579 0.00797283
R21036 gnd.n3093 gnd.n3091 0.00797283
R21037 gnd.n3092 gnd.n2462 0.00797283
R21038 gnd.n3160 gnd.n3158 0.00797283
R21039 gnd.n3159 gnd.n2455 0.00797283
R21040 gnd.n3170 gnd.n3169 0.00797283
R21041 gnd.n3172 gnd.n3171 0.00797283
R21042 gnd.n3175 gnd.n2453 0.00797283
R21043 gnd.n3179 gnd.n3178 0.00797283
R21044 gnd.n3177 gnd.n3176 0.00797283
R21045 gnd.n2433 gnd.n2432 0.00797283
R21046 gnd.n3201 gnd.n3200 0.00797283
R21047 gnd.n2434 gnd.n2407 0.00797283
R21048 gnd.n3245 gnd.n3243 0.00797283
R21049 gnd.n3244 gnd.n2400 0.00797283
R21050 gnd.n3255 gnd.n3254 0.00797283
R21051 gnd.n3257 gnd.n3256 0.00797283
R21052 gnd.n3260 gnd.n2398 0.00797283
R21053 gnd.n3264 gnd.n3263 0.00797283
R21054 gnd.n3262 gnd.n3261 0.00797283
R21055 gnd.n2378 gnd.n2377 0.00797283
R21056 gnd.n3286 gnd.n3285 0.00797283
R21057 gnd.n2379 gnd.n2353 0.00797283
R21058 gnd.n3334 gnd.n3332 0.00797283
R21059 gnd.n3333 gnd.n2346 0.00797283
R21060 gnd.n3344 gnd.n3343 0.00797283
R21061 gnd.n3602 gnd.n3601 0.00797283
R21062 gnd.n3605 gnd.n2344 0.00797283
R21063 gnd.n3607 gnd.n3606 0.00797283
R21064 gnd.n3630 gnd.n2325 0.00797283
R21065 gnd.n3631 gnd.n2288 0.00797283
R21066 gnd.n4379 gnd.n1913 0.00593478
R21067 gnd.n5591 gnd.n5590 0.00593478
R21068 gnd.n6805 gnd.n326 0.00417647
R21069 gnd.n6806 gnd.n6805 0.00417647
R21070 gnd.n6807 gnd.n6806 0.00417647
R21071 gnd.n6809 gnd.n6807 0.00417647
R21072 gnd.n6809 gnd.n6808 0.00417647
R21073 gnd.n6808 gnd.n91 0.00417647
R21074 gnd.n92 gnd.n91 0.00417647
R21075 gnd.n93 gnd.n92 0.00417647
R21076 gnd.n111 gnd.n93 0.00417647
R21077 gnd.n4189 gnd.n2129 0.00417647
R21078 gnd.n4190 gnd.n4189 0.00417647
R21079 gnd.n4191 gnd.n4190 0.00417647
R21080 gnd.n4192 gnd.n4191 0.00417647
R21081 gnd.n4192 gnd.n2104 0.00417647
R21082 gnd.n4232 gnd.n2104 0.00417647
R21083 gnd.n4233 gnd.n4232 0.00417647
R21084 gnd.n4234 gnd.n4233 0.00417647
R21085 gnd.n4234 gnd.n2083 0.00417647
R21086 a_n1986_8322.n6 a_n1986_8322.t5 74.6477
R21087 a_n1986_8322.n1 a_n1986_8322.t11 74.6477
R21088 a_n1986_8322.t20 a_n1986_8322.n18 74.6476
R21089 a_n1986_8322.n14 a_n1986_8322.t12 74.2899
R21090 a_n1986_8322.n7 a_n1986_8322.t3 74.2899
R21091 a_n1986_8322.n8 a_n1986_8322.t6 74.2899
R21092 a_n1986_8322.n11 a_n1986_8322.t7 74.2899
R21093 a_n1986_8322.n4 a_n1986_8322.t10 74.2899
R21094 a_n1986_8322.n18 a_n1986_8322.n17 70.6783
R21095 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R21096 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R21097 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R21098 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R21099 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R21100 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R21101 a_n1986_8322.n13 a_n1986_8322.t1 9.96389
R21102 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R21103 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R21104 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R21105 a_n1986_8322.n17 a_n1986_8322.t18 3.61217
R21106 a_n1986_8322.n17 a_n1986_8322.t15 3.61217
R21107 a_n1986_8322.n15 a_n1986_8322.t13 3.61217
R21108 a_n1986_8322.n15 a_n1986_8322.t21 3.61217
R21109 a_n1986_8322.n5 a_n1986_8322.t8 3.61217
R21110 a_n1986_8322.n5 a_n1986_8322.t9 3.61217
R21111 a_n1986_8322.n9 a_n1986_8322.t4 3.61217
R21112 a_n1986_8322.n9 a_n1986_8322.t2 3.61217
R21113 a_n1986_8322.n0 a_n1986_8322.t19 3.61217
R21114 a_n1986_8322.n0 a_n1986_8322.t14 3.61217
R21115 a_n1986_8322.n2 a_n1986_8322.t17 3.61217
R21116 a_n1986_8322.n2 a_n1986_8322.t16 3.61217
R21117 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R21118 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R21119 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R21120 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R21121 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R21122 a_n1986_8322.n16 a_n1986_8322.n14 0.358259
R21123 a_n1986_8322.n18 a_n1986_8322.n16 0.358259
R21124 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R21125 a_n1986_8322.t1 a_n1986_8322.t0 0.057021
R21126 plus.n46 plus.t9 252.611
R21127 plus.n9 plus.t11 252.611
R21128 plus.n76 plus.t4 243.97
R21129 plus.n72 plus.t12 231.093
R21130 plus.n35 plus.t7 231.093
R21131 plus.n76 plus.n75 223.454
R21132 plus.n78 plus.n77 223.454
R21133 plus.n47 plus.t5 187.445
R21134 plus.n44 plus.t18 187.445
R21135 plus.n42 plus.t17 187.445
R21136 plus.n59 plus.t13 187.445
R21137 plus.n65 plus.t14 187.445
R21138 plus.n38 plus.t10 187.445
R21139 plus.n1 plus.t6 187.445
R21140 plus.n28 plus.t16 187.445
R21141 plus.n22 plus.t15 187.445
R21142 plus.n5 plus.t20 187.445
R21143 plus.n7 plus.t19 187.445
R21144 plus.n10 plus.t8 187.445
R21145 plus.n73 plus.n72 161.3
R21146 plus.n71 plus.n37 161.3
R21147 plus.n70 plus.n69 161.3
R21148 plus.n68 plus.n67 161.3
R21149 plus.n66 plus.n39 161.3
R21150 plus.n64 plus.n63 161.3
R21151 plus.n62 plus.n40 161.3
R21152 plus.n61 plus.n60 161.3
R21153 plus.n58 plus.n41 161.3
R21154 plus.n57 plus.n56 161.3
R21155 plus.n55 plus.n54 161.3
R21156 plus.n53 plus.n43 161.3
R21157 plus.n52 plus.n51 161.3
R21158 plus.n50 plus.n49 161.3
R21159 plus.n48 plus.n45 161.3
R21160 plus.n11 plus.n8 161.3
R21161 plus.n13 plus.n12 161.3
R21162 plus.n15 plus.n14 161.3
R21163 plus.n16 plus.n6 161.3
R21164 plus.n18 plus.n17 161.3
R21165 plus.n20 plus.n19 161.3
R21166 plus.n21 plus.n4 161.3
R21167 plus.n24 plus.n23 161.3
R21168 plus.n25 plus.n3 161.3
R21169 plus.n27 plus.n26 161.3
R21170 plus.n29 plus.n2 161.3
R21171 plus.n31 plus.n30 161.3
R21172 plus.n33 plus.n32 161.3
R21173 plus.n34 plus.n0 161.3
R21174 plus.n36 plus.n35 161.3
R21175 plus.n49 plus.n48 56.5617
R21176 plus.n58 plus.n57 56.5617
R21177 plus.n67 plus.n66 56.5617
R21178 plus.n30 plus.n29 56.5617
R21179 plus.n21 plus.n20 56.5617
R21180 plus.n12 plus.n11 56.5617
R21181 plus.n71 plus.n70 46.3896
R21182 plus.n34 plus.n33 46.3896
R21183 plus.n46 plus.n45 42.8164
R21184 plus.n9 plus.n8 42.8164
R21185 plus.n54 plus.n53 42.5146
R21186 plus.n60 plus.n40 42.5146
R21187 plus.n23 plus.n3 42.5146
R21188 plus.n17 plus.n16 42.5146
R21189 plus.n53 plus.n52 38.6395
R21190 plus.n64 plus.n40 38.6395
R21191 plus.n27 plus.n3 38.6395
R21192 plus.n16 plus.n15 38.6395
R21193 plus.n47 plus.n46 38.2514
R21194 plus.n10 plus.n9 38.2514
R21195 plus.n74 plus.n73 31.491
R21196 plus.n49 plus.n44 19.9199
R21197 plus.n66 plus.n65 19.9199
R21198 plus.n29 plus.n28 19.9199
R21199 plus.n12 plus.n7 19.9199
R21200 plus.n75 plus.t1 19.8005
R21201 plus.n75 plus.t2 19.8005
R21202 plus.n77 plus.t0 19.8005
R21203 plus.n77 plus.t3 19.8005
R21204 plus.n57 plus.n42 17.9525
R21205 plus.n59 plus.n58 17.9525
R21206 plus.n22 plus.n21 17.9525
R21207 plus.n20 plus.n5 17.9525
R21208 plus.n48 plus.n47 15.9852
R21209 plus.n67 plus.n38 15.9852
R21210 plus.n30 plus.n1 15.9852
R21211 plus.n11 plus.n10 15.9852
R21212 plus.n72 plus.n71 15.3369
R21213 plus.n35 plus.n34 15.3369
R21214 plus plus.n79 14.4284
R21215 plus.n74 plus.n36 11.9494
R21216 plus.n70 plus.n38 8.60764
R21217 plus.n33 plus.n1 8.60764
R21218 plus.n54 plus.n42 6.6403
R21219 plus.n60 plus.n59 6.6403
R21220 plus.n23 plus.n22 6.6403
R21221 plus.n17 plus.n5 6.6403
R21222 plus.n79 plus.n78 5.40567
R21223 plus.n52 plus.n44 4.67295
R21224 plus.n65 plus.n64 4.67295
R21225 plus.n28 plus.n27 4.67295
R21226 plus.n15 plus.n7 4.67295
R21227 plus.n79 plus.n74 1.188
R21228 plus.n78 plus.n76 0.716017
R21229 plus.n50 plus.n45 0.189894
R21230 plus.n51 plus.n50 0.189894
R21231 plus.n51 plus.n43 0.189894
R21232 plus.n55 plus.n43 0.189894
R21233 plus.n56 plus.n55 0.189894
R21234 plus.n56 plus.n41 0.189894
R21235 plus.n61 plus.n41 0.189894
R21236 plus.n62 plus.n61 0.189894
R21237 plus.n63 plus.n62 0.189894
R21238 plus.n63 plus.n39 0.189894
R21239 plus.n68 plus.n39 0.189894
R21240 plus.n69 plus.n68 0.189894
R21241 plus.n69 plus.n37 0.189894
R21242 plus.n73 plus.n37 0.189894
R21243 plus.n36 plus.n0 0.189894
R21244 plus.n32 plus.n0 0.189894
R21245 plus.n32 plus.n31 0.189894
R21246 plus.n31 plus.n2 0.189894
R21247 plus.n26 plus.n2 0.189894
R21248 plus.n26 plus.n25 0.189894
R21249 plus.n25 plus.n24 0.189894
R21250 plus.n24 plus.n4 0.189894
R21251 plus.n19 plus.n4 0.189894
R21252 plus.n19 plus.n18 0.189894
R21253 plus.n18 plus.n6 0.189894
R21254 plus.n14 plus.n6 0.189894
R21255 plus.n14 plus.n13 0.189894
R21256 plus.n13 plus.n8 0.189894
R21257 a_n2903_n3924.n0 a_n2903_n3924.t39 214.981
R21258 a_n2903_n3924.n2 a_n2903_n3924.t3 214.452
R21259 a_n2903_n3924.n11 a_n2903_n3924.t5 214.321
R21260 a_n2903_n3924.n12 a_n2903_n3924.t0 214.321
R21261 a_n2903_n3924.n13 a_n2903_n3924.t38 214.321
R21262 a_n2903_n3924.n14 a_n2903_n3924.t1 214.321
R21263 a_n2903_n3924.n15 a_n2903_n3924.t2 214.321
R21264 a_n2903_n3924.n0 a_n2903_n3924.t4 214.321
R21265 a_n2903_n3924.n1 a_n2903_n3924.t33 55.8337
R21266 a_n2903_n3924.n3 a_n2903_n3924.t19 55.8337
R21267 a_n2903_n3924.n10 a_n2903_n3924.t18 55.8337
R21268 a_n2903_n3924.n34 a_n2903_n3924.t30 55.8335
R21269 a_n2903_n3924.n32 a_n2903_n3924.t13 55.8335
R21270 a_n2903_n3924.n25 a_n2903_n3924.t15 55.8335
R21271 a_n2903_n3924.n24 a_n2903_n3924.t31 55.8335
R21272 a_n2903_n3924.n17 a_n2903_n3924.t35 55.8335
R21273 a_n2903_n3924.n36 a_n2903_n3924.n35 53.0052
R21274 a_n2903_n3924.n38 a_n2903_n3924.n37 53.0052
R21275 a_n2903_n3924.n5 a_n2903_n3924.n4 53.0052
R21276 a_n2903_n3924.n7 a_n2903_n3924.n6 53.0052
R21277 a_n2903_n3924.n9 a_n2903_n3924.n8 53.0052
R21278 a_n2903_n3924.n31 a_n2903_n3924.n30 53.0051
R21279 a_n2903_n3924.n29 a_n2903_n3924.n28 53.0051
R21280 a_n2903_n3924.n27 a_n2903_n3924.n26 53.0051
R21281 a_n2903_n3924.n23 a_n2903_n3924.n22 53.0051
R21282 a_n2903_n3924.n21 a_n2903_n3924.n20 53.0051
R21283 a_n2903_n3924.n19 a_n2903_n3924.n18 53.0051
R21284 a_n2903_n3924.n40 a_n2903_n3924.n39 53.0051
R21285 a_n2903_n3924.n16 a_n2903_n3924.n10 12.2417
R21286 a_n2903_n3924.n34 a_n2903_n3924.n33 12.2417
R21287 a_n2903_n3924.n17 a_n2903_n3924.n16 5.16214
R21288 a_n2903_n3924.n33 a_n2903_n3924.n32 5.16214
R21289 a_n2903_n3924.n35 a_n2903_n3924.t28 2.82907
R21290 a_n2903_n3924.n35 a_n2903_n3924.t32 2.82907
R21291 a_n2903_n3924.n37 a_n2903_n3924.t25 2.82907
R21292 a_n2903_n3924.n37 a_n2903_n3924.t29 2.82907
R21293 a_n2903_n3924.n4 a_n2903_n3924.t8 2.82907
R21294 a_n2903_n3924.n4 a_n2903_n3924.t21 2.82907
R21295 a_n2903_n3924.n6 a_n2903_n3924.t6 2.82907
R21296 a_n2903_n3924.n6 a_n2903_n3924.t16 2.82907
R21297 a_n2903_n3924.n8 a_n2903_n3924.t11 2.82907
R21298 a_n2903_n3924.n8 a_n2903_n3924.t10 2.82907
R21299 a_n2903_n3924.n30 a_n2903_n3924.t20 2.82907
R21300 a_n2903_n3924.n30 a_n2903_n3924.t14 2.82907
R21301 a_n2903_n3924.n28 a_n2903_n3924.t7 2.82907
R21302 a_n2903_n3924.n28 a_n2903_n3924.t12 2.82907
R21303 a_n2903_n3924.n26 a_n2903_n3924.t9 2.82907
R21304 a_n2903_n3924.n26 a_n2903_n3924.t17 2.82907
R21305 a_n2903_n3924.n22 a_n2903_n3924.t23 2.82907
R21306 a_n2903_n3924.n22 a_n2903_n3924.t34 2.82907
R21307 a_n2903_n3924.n20 a_n2903_n3924.t27 2.82907
R21308 a_n2903_n3924.n20 a_n2903_n3924.t22 2.82907
R21309 a_n2903_n3924.n18 a_n2903_n3924.t36 2.82907
R21310 a_n2903_n3924.n18 a_n2903_n3924.t26 2.82907
R21311 a_n2903_n3924.t37 a_n2903_n3924.n40 2.82907
R21312 a_n2903_n3924.n40 a_n2903_n3924.t24 2.82907
R21313 a_n2903_n3924.n33 a_n2903_n3924.n2 1.95694
R21314 a_n2903_n3924.n16 a_n2903_n3924.n0 1.95694
R21315 a_n2903_n3924.n0 a_n2903_n3924.n15 0.684366
R21316 a_n2903_n3924.n15 a_n2903_n3924.n14 0.672012
R21317 a_n2903_n3924.n14 a_n2903_n3924.n13 0.672012
R21318 a_n2903_n3924.n13 a_n2903_n3924.n12 0.672012
R21319 a_n2903_n3924.n12 a_n2903_n3924.n11 0.672012
R21320 a_n2903_n3924.n11 a_n2903_n3924.n2 0.541924
R21321 a_n2903_n3924.n19 a_n2903_n3924.n17 0.530672
R21322 a_n2903_n3924.n21 a_n2903_n3924.n19 0.530672
R21323 a_n2903_n3924.n23 a_n2903_n3924.n21 0.530672
R21324 a_n2903_n3924.n24 a_n2903_n3924.n23 0.530672
R21325 a_n2903_n3924.n27 a_n2903_n3924.n25 0.530672
R21326 a_n2903_n3924.n29 a_n2903_n3924.n27 0.530672
R21327 a_n2903_n3924.n31 a_n2903_n3924.n29 0.530672
R21328 a_n2903_n3924.n32 a_n2903_n3924.n31 0.530672
R21329 a_n2903_n3924.n10 a_n2903_n3924.n9 0.530672
R21330 a_n2903_n3924.n9 a_n2903_n3924.n7 0.530672
R21331 a_n2903_n3924.n7 a_n2903_n3924.n5 0.530672
R21332 a_n2903_n3924.n5 a_n2903_n3924.n3 0.530672
R21333 a_n2903_n3924.n39 a_n2903_n3924.n1 0.530672
R21334 a_n2903_n3924.n39 a_n2903_n3924.n38 0.530672
R21335 a_n2903_n3924.n38 a_n2903_n3924.n36 0.530672
R21336 a_n2903_n3924.n36 a_n2903_n3924.n34 0.530672
R21337 a_n2903_n3924.n25 a_n2903_n3924.n24 0.235414
R21338 a_n2903_n3924.n3 a_n2903_n3924.n1 0.235414
R21339 minus.n46 minus.t20 252.611
R21340 minus.n9 minus.t13 252.611
R21341 minus.n78 minus.t3 243.255
R21342 minus.n72 minus.t15 231.093
R21343 minus.n35 minus.t17 231.093
R21344 minus.n77 minus.n75 224.169
R21345 minus.n77 minus.n76 223.454
R21346 minus.n38 minus.t12 187.445
R21347 minus.n65 minus.t7 187.445
R21348 minus.n59 minus.t6 187.445
R21349 minus.n42 minus.t11 187.445
R21350 minus.n44 minus.t10 187.445
R21351 minus.n47 minus.t16 187.445
R21352 minus.n10 minus.t9 187.445
R21353 minus.n7 minus.t8 187.445
R21354 minus.n5 minus.t5 187.445
R21355 minus.n22 minus.t18 187.445
R21356 minus.n28 minus.t19 187.445
R21357 minus.n1 minus.t14 187.445
R21358 minus.n48 minus.n45 161.3
R21359 minus.n50 minus.n49 161.3
R21360 minus.n52 minus.n51 161.3
R21361 minus.n53 minus.n43 161.3
R21362 minus.n55 minus.n54 161.3
R21363 minus.n57 minus.n56 161.3
R21364 minus.n58 minus.n41 161.3
R21365 minus.n61 minus.n60 161.3
R21366 minus.n62 minus.n40 161.3
R21367 minus.n64 minus.n63 161.3
R21368 minus.n66 minus.n39 161.3
R21369 minus.n68 minus.n67 161.3
R21370 minus.n70 minus.n69 161.3
R21371 minus.n71 minus.n37 161.3
R21372 minus.n73 minus.n72 161.3
R21373 minus.n36 minus.n35 161.3
R21374 minus.n34 minus.n0 161.3
R21375 minus.n33 minus.n32 161.3
R21376 minus.n31 minus.n30 161.3
R21377 minus.n29 minus.n2 161.3
R21378 minus.n27 minus.n26 161.3
R21379 minus.n25 minus.n3 161.3
R21380 minus.n24 minus.n23 161.3
R21381 minus.n21 minus.n4 161.3
R21382 minus.n20 minus.n19 161.3
R21383 minus.n18 minus.n17 161.3
R21384 minus.n16 minus.n6 161.3
R21385 minus.n15 minus.n14 161.3
R21386 minus.n13 minus.n12 161.3
R21387 minus.n11 minus.n8 161.3
R21388 minus.n67 minus.n66 56.5617
R21389 minus.n58 minus.n57 56.5617
R21390 minus.n49 minus.n48 56.5617
R21391 minus.n12 minus.n11 56.5617
R21392 minus.n21 minus.n20 56.5617
R21393 minus.n30 minus.n29 56.5617
R21394 minus.n71 minus.n70 46.3896
R21395 minus.n34 minus.n33 46.3896
R21396 minus.n46 minus.n45 42.8164
R21397 minus.n9 minus.n8 42.8164
R21398 minus.n60 minus.n40 42.5146
R21399 minus.n54 minus.n53 42.5146
R21400 minus.n17 minus.n16 42.5146
R21401 minus.n23 minus.n3 42.5146
R21402 minus.n64 minus.n40 38.6395
R21403 minus.n53 minus.n52 38.6395
R21404 minus.n16 minus.n15 38.6395
R21405 minus.n27 minus.n3 38.6395
R21406 minus.n47 minus.n46 38.2514
R21407 minus.n10 minus.n9 38.2514
R21408 minus.n74 minus.n73 31.7069
R21409 minus.n66 minus.n65 19.9199
R21410 minus.n49 minus.n44 19.9199
R21411 minus.n12 minus.n7 19.9199
R21412 minus.n29 minus.n28 19.9199
R21413 minus.n76 minus.t2 19.8005
R21414 minus.n76 minus.t0 19.8005
R21415 minus.n75 minus.t1 19.8005
R21416 minus.n75 minus.t4 19.8005
R21417 minus.n59 minus.n58 17.9525
R21418 minus.n57 minus.n42 17.9525
R21419 minus.n20 minus.n5 17.9525
R21420 minus.n22 minus.n21 17.9525
R21421 minus.n67 minus.n38 15.9852
R21422 minus.n48 minus.n47 15.9852
R21423 minus.n11 minus.n10 15.9852
R21424 minus.n30 minus.n1 15.9852
R21425 minus.n72 minus.n71 15.3369
R21426 minus.n35 minus.n34 15.3369
R21427 minus.n74 minus.n36 12.1653
R21428 minus minus.n79 11.5562
R21429 minus.n70 minus.n38 8.60764
R21430 minus.n33 minus.n1 8.60764
R21431 minus.n60 minus.n59 6.6403
R21432 minus.n54 minus.n42 6.6403
R21433 minus.n17 minus.n5 6.6403
R21434 minus.n23 minus.n22 6.6403
R21435 minus.n79 minus.n78 4.80222
R21436 minus.n65 minus.n64 4.67295
R21437 minus.n52 minus.n44 4.67295
R21438 minus.n15 minus.n7 4.67295
R21439 minus.n28 minus.n27 4.67295
R21440 minus.n79 minus.n74 0.972091
R21441 minus.n78 minus.n77 0.716017
R21442 minus.n73 minus.n37 0.189894
R21443 minus.n69 minus.n37 0.189894
R21444 minus.n69 minus.n68 0.189894
R21445 minus.n68 minus.n39 0.189894
R21446 minus.n63 minus.n39 0.189894
R21447 minus.n63 minus.n62 0.189894
R21448 minus.n62 minus.n61 0.189894
R21449 minus.n61 minus.n41 0.189894
R21450 minus.n56 minus.n41 0.189894
R21451 minus.n56 minus.n55 0.189894
R21452 minus.n55 minus.n43 0.189894
R21453 minus.n51 minus.n43 0.189894
R21454 minus.n51 minus.n50 0.189894
R21455 minus.n50 minus.n45 0.189894
R21456 minus.n13 minus.n8 0.189894
R21457 minus.n14 minus.n13 0.189894
R21458 minus.n14 minus.n6 0.189894
R21459 minus.n18 minus.n6 0.189894
R21460 minus.n19 minus.n18 0.189894
R21461 minus.n19 minus.n4 0.189894
R21462 minus.n24 minus.n4 0.189894
R21463 minus.n25 minus.n24 0.189894
R21464 minus.n26 minus.n25 0.189894
R21465 minus.n26 minus.n2 0.189894
R21466 minus.n31 minus.n2 0.189894
R21467 minus.n32 minus.n31 0.189894
R21468 minus.n32 minus.n0 0.189894
R21469 minus.n36 minus.n0 0.189894
R21470 output.n41 output.n15 289.615
R21471 output.n72 output.n46 289.615
R21472 output.n104 output.n78 289.615
R21473 output.n136 output.n110 289.615
R21474 output.n77 output.n45 197.26
R21475 output.n77 output.n76 196.298
R21476 output.n109 output.n108 196.298
R21477 output.n141 output.n140 196.298
R21478 output.n42 output.n41 185
R21479 output.n40 output.n39 185
R21480 output.n19 output.n18 185
R21481 output.n34 output.n33 185
R21482 output.n32 output.n31 185
R21483 output.n23 output.n22 185
R21484 output.n26 output.n25 185
R21485 output.n73 output.n72 185
R21486 output.n71 output.n70 185
R21487 output.n50 output.n49 185
R21488 output.n65 output.n64 185
R21489 output.n63 output.n62 185
R21490 output.n54 output.n53 185
R21491 output.n57 output.n56 185
R21492 output.n105 output.n104 185
R21493 output.n103 output.n102 185
R21494 output.n82 output.n81 185
R21495 output.n97 output.n96 185
R21496 output.n95 output.n94 185
R21497 output.n86 output.n85 185
R21498 output.n89 output.n88 185
R21499 output.n137 output.n136 185
R21500 output.n135 output.n134 185
R21501 output.n114 output.n113 185
R21502 output.n129 output.n128 185
R21503 output.n127 output.n126 185
R21504 output.n118 output.n117 185
R21505 output.n121 output.n120 185
R21506 output.t0 output.n24 147.661
R21507 output.t19 output.n55 147.661
R21508 output.t2 output.n87 147.661
R21509 output.t1 output.n119 147.661
R21510 output.n41 output.n40 104.615
R21511 output.n40 output.n18 104.615
R21512 output.n33 output.n18 104.615
R21513 output.n33 output.n32 104.615
R21514 output.n32 output.n22 104.615
R21515 output.n25 output.n22 104.615
R21516 output.n72 output.n71 104.615
R21517 output.n71 output.n49 104.615
R21518 output.n64 output.n49 104.615
R21519 output.n64 output.n63 104.615
R21520 output.n63 output.n53 104.615
R21521 output.n56 output.n53 104.615
R21522 output.n104 output.n103 104.615
R21523 output.n103 output.n81 104.615
R21524 output.n96 output.n81 104.615
R21525 output.n96 output.n95 104.615
R21526 output.n95 output.n85 104.615
R21527 output.n88 output.n85 104.615
R21528 output.n136 output.n135 104.615
R21529 output.n135 output.n113 104.615
R21530 output.n128 output.n113 104.615
R21531 output.n128 output.n127 104.615
R21532 output.n127 output.n117 104.615
R21533 output.n120 output.n117 104.615
R21534 output.n1 output.t5 77.056
R21535 output.n14 output.t6 76.6694
R21536 output.n1 output.n0 72.7095
R21537 output.n3 output.n2 72.7095
R21538 output.n5 output.n4 72.7095
R21539 output.n7 output.n6 72.7095
R21540 output.n9 output.n8 72.7095
R21541 output.n11 output.n10 72.7095
R21542 output.n13 output.n12 72.7095
R21543 output.n25 output.t0 52.3082
R21544 output.n56 output.t19 52.3082
R21545 output.n88 output.t2 52.3082
R21546 output.n120 output.t1 52.3082
R21547 output.n26 output.n24 15.6674
R21548 output.n57 output.n55 15.6674
R21549 output.n89 output.n87 15.6674
R21550 output.n121 output.n119 15.6674
R21551 output.n27 output.n23 12.8005
R21552 output.n58 output.n54 12.8005
R21553 output.n90 output.n86 12.8005
R21554 output.n122 output.n118 12.8005
R21555 output.n31 output.n30 12.0247
R21556 output.n62 output.n61 12.0247
R21557 output.n94 output.n93 12.0247
R21558 output.n126 output.n125 12.0247
R21559 output.n34 output.n21 11.249
R21560 output.n65 output.n52 11.249
R21561 output.n97 output.n84 11.249
R21562 output.n129 output.n116 11.249
R21563 output.n35 output.n19 10.4732
R21564 output.n66 output.n50 10.4732
R21565 output.n98 output.n82 10.4732
R21566 output.n130 output.n114 10.4732
R21567 output.n39 output.n38 9.69747
R21568 output.n70 output.n69 9.69747
R21569 output.n102 output.n101 9.69747
R21570 output.n134 output.n133 9.69747
R21571 output.n45 output.n44 9.45567
R21572 output.n76 output.n75 9.45567
R21573 output.n108 output.n107 9.45567
R21574 output.n140 output.n139 9.45567
R21575 output.n44 output.n43 9.3005
R21576 output.n17 output.n16 9.3005
R21577 output.n38 output.n37 9.3005
R21578 output.n36 output.n35 9.3005
R21579 output.n21 output.n20 9.3005
R21580 output.n30 output.n29 9.3005
R21581 output.n28 output.n27 9.3005
R21582 output.n75 output.n74 9.3005
R21583 output.n48 output.n47 9.3005
R21584 output.n69 output.n68 9.3005
R21585 output.n67 output.n66 9.3005
R21586 output.n52 output.n51 9.3005
R21587 output.n61 output.n60 9.3005
R21588 output.n59 output.n58 9.3005
R21589 output.n107 output.n106 9.3005
R21590 output.n80 output.n79 9.3005
R21591 output.n101 output.n100 9.3005
R21592 output.n99 output.n98 9.3005
R21593 output.n84 output.n83 9.3005
R21594 output.n93 output.n92 9.3005
R21595 output.n91 output.n90 9.3005
R21596 output.n139 output.n138 9.3005
R21597 output.n112 output.n111 9.3005
R21598 output.n133 output.n132 9.3005
R21599 output.n131 output.n130 9.3005
R21600 output.n116 output.n115 9.3005
R21601 output.n125 output.n124 9.3005
R21602 output.n123 output.n122 9.3005
R21603 output.n42 output.n17 8.92171
R21604 output.n73 output.n48 8.92171
R21605 output.n105 output.n80 8.92171
R21606 output.n137 output.n112 8.92171
R21607 output output.n141 8.15037
R21608 output.n43 output.n15 8.14595
R21609 output.n74 output.n46 8.14595
R21610 output.n106 output.n78 8.14595
R21611 output.n138 output.n110 8.14595
R21612 output.n45 output.n15 5.81868
R21613 output.n76 output.n46 5.81868
R21614 output.n108 output.n78 5.81868
R21615 output.n140 output.n110 5.81868
R21616 output.n43 output.n42 5.04292
R21617 output.n74 output.n73 5.04292
R21618 output.n106 output.n105 5.04292
R21619 output.n138 output.n137 5.04292
R21620 output.n28 output.n24 4.38594
R21621 output.n59 output.n55 4.38594
R21622 output.n91 output.n87 4.38594
R21623 output.n123 output.n119 4.38594
R21624 output.n39 output.n17 4.26717
R21625 output.n70 output.n48 4.26717
R21626 output.n102 output.n80 4.26717
R21627 output.n134 output.n112 4.26717
R21628 output.n0 output.t10 3.9605
R21629 output.n0 output.t15 3.9605
R21630 output.n2 output.t3 3.9605
R21631 output.n2 output.t11 3.9605
R21632 output.n4 output.t14 3.9605
R21633 output.n4 output.t12 3.9605
R21634 output.n6 output.t18 3.9605
R21635 output.n6 output.t4 3.9605
R21636 output.n8 output.t7 3.9605
R21637 output.n8 output.t16 3.9605
R21638 output.n10 output.t17 3.9605
R21639 output.n10 output.t8 3.9605
R21640 output.n12 output.t9 3.9605
R21641 output.n12 output.t13 3.9605
R21642 output.n38 output.n19 3.49141
R21643 output.n69 output.n50 3.49141
R21644 output.n101 output.n82 3.49141
R21645 output.n133 output.n114 3.49141
R21646 output.n35 output.n34 2.71565
R21647 output.n66 output.n65 2.71565
R21648 output.n98 output.n97 2.71565
R21649 output.n130 output.n129 2.71565
R21650 output.n31 output.n21 1.93989
R21651 output.n62 output.n52 1.93989
R21652 output.n94 output.n84 1.93989
R21653 output.n126 output.n116 1.93989
R21654 output.n30 output.n23 1.16414
R21655 output.n61 output.n54 1.16414
R21656 output.n93 output.n86 1.16414
R21657 output.n125 output.n118 1.16414
R21658 output.n141 output.n109 0.962709
R21659 output.n109 output.n77 0.962709
R21660 output.n27 output.n26 0.388379
R21661 output.n58 output.n57 0.388379
R21662 output.n90 output.n89 0.388379
R21663 output.n122 output.n121 0.388379
R21664 output.n14 output.n13 0.387128
R21665 output.n13 output.n11 0.387128
R21666 output.n11 output.n9 0.387128
R21667 output.n9 output.n7 0.387128
R21668 output.n7 output.n5 0.387128
R21669 output.n5 output.n3 0.387128
R21670 output.n3 output.n1 0.387128
R21671 output.n44 output.n16 0.155672
R21672 output.n37 output.n16 0.155672
R21673 output.n37 output.n36 0.155672
R21674 output.n36 output.n20 0.155672
R21675 output.n29 output.n20 0.155672
R21676 output.n29 output.n28 0.155672
R21677 output.n75 output.n47 0.155672
R21678 output.n68 output.n47 0.155672
R21679 output.n68 output.n67 0.155672
R21680 output.n67 output.n51 0.155672
R21681 output.n60 output.n51 0.155672
R21682 output.n60 output.n59 0.155672
R21683 output.n107 output.n79 0.155672
R21684 output.n100 output.n79 0.155672
R21685 output.n100 output.n99 0.155672
R21686 output.n99 output.n83 0.155672
R21687 output.n92 output.n83 0.155672
R21688 output.n92 output.n91 0.155672
R21689 output.n139 output.n111 0.155672
R21690 output.n132 output.n111 0.155672
R21691 output.n132 output.n131 0.155672
R21692 output.n131 output.n115 0.155672
R21693 output.n124 output.n115 0.155672
R21694 output.n124 output.n123 0.155672
R21695 output output.n14 0.126227
R21696 diffpairibias.n0 diffpairibias.t18 436.822
R21697 diffpairibias.n21 diffpairibias.t19 435.479
R21698 diffpairibias.n20 diffpairibias.t16 435.479
R21699 diffpairibias.n19 diffpairibias.t17 435.479
R21700 diffpairibias.n18 diffpairibias.t21 435.479
R21701 diffpairibias.n0 diffpairibias.t22 435.479
R21702 diffpairibias.n1 diffpairibias.t20 435.479
R21703 diffpairibias.n2 diffpairibias.t23 435.479
R21704 diffpairibias.n10 diffpairibias.t0 377.536
R21705 diffpairibias.n10 diffpairibias.t8 376.193
R21706 diffpairibias.n11 diffpairibias.t10 376.193
R21707 diffpairibias.n12 diffpairibias.t6 376.193
R21708 diffpairibias.n13 diffpairibias.t2 376.193
R21709 diffpairibias.n14 diffpairibias.t12 376.193
R21710 diffpairibias.n15 diffpairibias.t4 376.193
R21711 diffpairibias.n16 diffpairibias.t14 376.193
R21712 diffpairibias.n3 diffpairibias.t1 113.368
R21713 diffpairibias.n3 diffpairibias.t9 112.698
R21714 diffpairibias.n4 diffpairibias.t11 112.698
R21715 diffpairibias.n5 diffpairibias.t7 112.698
R21716 diffpairibias.n6 diffpairibias.t3 112.698
R21717 diffpairibias.n7 diffpairibias.t13 112.698
R21718 diffpairibias.n8 diffpairibias.t5 112.698
R21719 diffpairibias.n9 diffpairibias.t15 112.698
R21720 diffpairibias.n17 diffpairibias.n16 4.77242
R21721 diffpairibias.n17 diffpairibias.n9 4.30807
R21722 diffpairibias.n18 diffpairibias.n17 4.13945
R21723 diffpairibias.n16 diffpairibias.n15 1.34352
R21724 diffpairibias.n15 diffpairibias.n14 1.34352
R21725 diffpairibias.n14 diffpairibias.n13 1.34352
R21726 diffpairibias.n13 diffpairibias.n12 1.34352
R21727 diffpairibias.n12 diffpairibias.n11 1.34352
R21728 diffpairibias.n11 diffpairibias.n10 1.34352
R21729 diffpairibias.n2 diffpairibias.n1 1.34352
R21730 diffpairibias.n1 diffpairibias.n0 1.34352
R21731 diffpairibias.n19 diffpairibias.n18 1.34352
R21732 diffpairibias.n20 diffpairibias.n19 1.34352
R21733 diffpairibias.n21 diffpairibias.n20 1.34352
R21734 diffpairibias.n22 diffpairibias.n21 0.862419
R21735 diffpairibias diffpairibias.n22 0.684875
R21736 diffpairibias.n9 diffpairibias.n8 0.672012
R21737 diffpairibias.n8 diffpairibias.n7 0.672012
R21738 diffpairibias.n7 diffpairibias.n6 0.672012
R21739 diffpairibias.n6 diffpairibias.n5 0.672012
R21740 diffpairibias.n5 diffpairibias.n4 0.672012
R21741 diffpairibias.n4 diffpairibias.n3 0.672012
R21742 diffpairibias.n22 diffpairibias.n2 0.190907
R21743 outputibias.n27 outputibias.n1 289.615
R21744 outputibias.n58 outputibias.n32 289.615
R21745 outputibias.n90 outputibias.n64 289.615
R21746 outputibias.n122 outputibias.n96 289.615
R21747 outputibias.n28 outputibias.n27 185
R21748 outputibias.n26 outputibias.n25 185
R21749 outputibias.n5 outputibias.n4 185
R21750 outputibias.n20 outputibias.n19 185
R21751 outputibias.n18 outputibias.n17 185
R21752 outputibias.n9 outputibias.n8 185
R21753 outputibias.n12 outputibias.n11 185
R21754 outputibias.n59 outputibias.n58 185
R21755 outputibias.n57 outputibias.n56 185
R21756 outputibias.n36 outputibias.n35 185
R21757 outputibias.n51 outputibias.n50 185
R21758 outputibias.n49 outputibias.n48 185
R21759 outputibias.n40 outputibias.n39 185
R21760 outputibias.n43 outputibias.n42 185
R21761 outputibias.n91 outputibias.n90 185
R21762 outputibias.n89 outputibias.n88 185
R21763 outputibias.n68 outputibias.n67 185
R21764 outputibias.n83 outputibias.n82 185
R21765 outputibias.n81 outputibias.n80 185
R21766 outputibias.n72 outputibias.n71 185
R21767 outputibias.n75 outputibias.n74 185
R21768 outputibias.n123 outputibias.n122 185
R21769 outputibias.n121 outputibias.n120 185
R21770 outputibias.n100 outputibias.n99 185
R21771 outputibias.n115 outputibias.n114 185
R21772 outputibias.n113 outputibias.n112 185
R21773 outputibias.n104 outputibias.n103 185
R21774 outputibias.n107 outputibias.n106 185
R21775 outputibias.n0 outputibias.t10 178.945
R21776 outputibias.n133 outputibias.t8 177.018
R21777 outputibias.n132 outputibias.t11 177.018
R21778 outputibias.n0 outputibias.t9 177.018
R21779 outputibias.t7 outputibias.n10 147.661
R21780 outputibias.t1 outputibias.n41 147.661
R21781 outputibias.t3 outputibias.n73 147.661
R21782 outputibias.t5 outputibias.n105 147.661
R21783 outputibias.n128 outputibias.t6 132.363
R21784 outputibias.n128 outputibias.t0 130.436
R21785 outputibias.n129 outputibias.t2 130.436
R21786 outputibias.n130 outputibias.t4 130.436
R21787 outputibias.n27 outputibias.n26 104.615
R21788 outputibias.n26 outputibias.n4 104.615
R21789 outputibias.n19 outputibias.n4 104.615
R21790 outputibias.n19 outputibias.n18 104.615
R21791 outputibias.n18 outputibias.n8 104.615
R21792 outputibias.n11 outputibias.n8 104.615
R21793 outputibias.n58 outputibias.n57 104.615
R21794 outputibias.n57 outputibias.n35 104.615
R21795 outputibias.n50 outputibias.n35 104.615
R21796 outputibias.n50 outputibias.n49 104.615
R21797 outputibias.n49 outputibias.n39 104.615
R21798 outputibias.n42 outputibias.n39 104.615
R21799 outputibias.n90 outputibias.n89 104.615
R21800 outputibias.n89 outputibias.n67 104.615
R21801 outputibias.n82 outputibias.n67 104.615
R21802 outputibias.n82 outputibias.n81 104.615
R21803 outputibias.n81 outputibias.n71 104.615
R21804 outputibias.n74 outputibias.n71 104.615
R21805 outputibias.n122 outputibias.n121 104.615
R21806 outputibias.n121 outputibias.n99 104.615
R21807 outputibias.n114 outputibias.n99 104.615
R21808 outputibias.n114 outputibias.n113 104.615
R21809 outputibias.n113 outputibias.n103 104.615
R21810 outputibias.n106 outputibias.n103 104.615
R21811 outputibias.n63 outputibias.n31 95.6354
R21812 outputibias.n63 outputibias.n62 94.6732
R21813 outputibias.n95 outputibias.n94 94.6732
R21814 outputibias.n127 outputibias.n126 94.6732
R21815 outputibias.n11 outputibias.t7 52.3082
R21816 outputibias.n42 outputibias.t1 52.3082
R21817 outputibias.n74 outputibias.t3 52.3082
R21818 outputibias.n106 outputibias.t5 52.3082
R21819 outputibias.n12 outputibias.n10 15.6674
R21820 outputibias.n43 outputibias.n41 15.6674
R21821 outputibias.n75 outputibias.n73 15.6674
R21822 outputibias.n107 outputibias.n105 15.6674
R21823 outputibias.n13 outputibias.n9 12.8005
R21824 outputibias.n44 outputibias.n40 12.8005
R21825 outputibias.n76 outputibias.n72 12.8005
R21826 outputibias.n108 outputibias.n104 12.8005
R21827 outputibias.n17 outputibias.n16 12.0247
R21828 outputibias.n48 outputibias.n47 12.0247
R21829 outputibias.n80 outputibias.n79 12.0247
R21830 outputibias.n112 outputibias.n111 12.0247
R21831 outputibias.n20 outputibias.n7 11.249
R21832 outputibias.n51 outputibias.n38 11.249
R21833 outputibias.n83 outputibias.n70 11.249
R21834 outputibias.n115 outputibias.n102 11.249
R21835 outputibias.n21 outputibias.n5 10.4732
R21836 outputibias.n52 outputibias.n36 10.4732
R21837 outputibias.n84 outputibias.n68 10.4732
R21838 outputibias.n116 outputibias.n100 10.4732
R21839 outputibias.n25 outputibias.n24 9.69747
R21840 outputibias.n56 outputibias.n55 9.69747
R21841 outputibias.n88 outputibias.n87 9.69747
R21842 outputibias.n120 outputibias.n119 9.69747
R21843 outputibias.n31 outputibias.n30 9.45567
R21844 outputibias.n62 outputibias.n61 9.45567
R21845 outputibias.n94 outputibias.n93 9.45567
R21846 outputibias.n126 outputibias.n125 9.45567
R21847 outputibias.n30 outputibias.n29 9.3005
R21848 outputibias.n3 outputibias.n2 9.3005
R21849 outputibias.n24 outputibias.n23 9.3005
R21850 outputibias.n22 outputibias.n21 9.3005
R21851 outputibias.n7 outputibias.n6 9.3005
R21852 outputibias.n16 outputibias.n15 9.3005
R21853 outputibias.n14 outputibias.n13 9.3005
R21854 outputibias.n61 outputibias.n60 9.3005
R21855 outputibias.n34 outputibias.n33 9.3005
R21856 outputibias.n55 outputibias.n54 9.3005
R21857 outputibias.n53 outputibias.n52 9.3005
R21858 outputibias.n38 outputibias.n37 9.3005
R21859 outputibias.n47 outputibias.n46 9.3005
R21860 outputibias.n45 outputibias.n44 9.3005
R21861 outputibias.n93 outputibias.n92 9.3005
R21862 outputibias.n66 outputibias.n65 9.3005
R21863 outputibias.n87 outputibias.n86 9.3005
R21864 outputibias.n85 outputibias.n84 9.3005
R21865 outputibias.n70 outputibias.n69 9.3005
R21866 outputibias.n79 outputibias.n78 9.3005
R21867 outputibias.n77 outputibias.n76 9.3005
R21868 outputibias.n125 outputibias.n124 9.3005
R21869 outputibias.n98 outputibias.n97 9.3005
R21870 outputibias.n119 outputibias.n118 9.3005
R21871 outputibias.n117 outputibias.n116 9.3005
R21872 outputibias.n102 outputibias.n101 9.3005
R21873 outputibias.n111 outputibias.n110 9.3005
R21874 outputibias.n109 outputibias.n108 9.3005
R21875 outputibias.n28 outputibias.n3 8.92171
R21876 outputibias.n59 outputibias.n34 8.92171
R21877 outputibias.n91 outputibias.n66 8.92171
R21878 outputibias.n123 outputibias.n98 8.92171
R21879 outputibias.n29 outputibias.n1 8.14595
R21880 outputibias.n60 outputibias.n32 8.14595
R21881 outputibias.n92 outputibias.n64 8.14595
R21882 outputibias.n124 outputibias.n96 8.14595
R21883 outputibias.n31 outputibias.n1 5.81868
R21884 outputibias.n62 outputibias.n32 5.81868
R21885 outputibias.n94 outputibias.n64 5.81868
R21886 outputibias.n126 outputibias.n96 5.81868
R21887 outputibias.n131 outputibias.n130 5.20947
R21888 outputibias.n29 outputibias.n28 5.04292
R21889 outputibias.n60 outputibias.n59 5.04292
R21890 outputibias.n92 outputibias.n91 5.04292
R21891 outputibias.n124 outputibias.n123 5.04292
R21892 outputibias.n131 outputibias.n127 4.42209
R21893 outputibias.n14 outputibias.n10 4.38594
R21894 outputibias.n45 outputibias.n41 4.38594
R21895 outputibias.n77 outputibias.n73 4.38594
R21896 outputibias.n109 outputibias.n105 4.38594
R21897 outputibias.n132 outputibias.n131 4.28454
R21898 outputibias.n25 outputibias.n3 4.26717
R21899 outputibias.n56 outputibias.n34 4.26717
R21900 outputibias.n88 outputibias.n66 4.26717
R21901 outputibias.n120 outputibias.n98 4.26717
R21902 outputibias.n24 outputibias.n5 3.49141
R21903 outputibias.n55 outputibias.n36 3.49141
R21904 outputibias.n87 outputibias.n68 3.49141
R21905 outputibias.n119 outputibias.n100 3.49141
R21906 outputibias.n21 outputibias.n20 2.71565
R21907 outputibias.n52 outputibias.n51 2.71565
R21908 outputibias.n84 outputibias.n83 2.71565
R21909 outputibias.n116 outputibias.n115 2.71565
R21910 outputibias.n17 outputibias.n7 1.93989
R21911 outputibias.n48 outputibias.n38 1.93989
R21912 outputibias.n80 outputibias.n70 1.93989
R21913 outputibias.n112 outputibias.n102 1.93989
R21914 outputibias.n130 outputibias.n129 1.9266
R21915 outputibias.n129 outputibias.n128 1.9266
R21916 outputibias.n133 outputibias.n132 1.92658
R21917 outputibias.n134 outputibias.n133 1.29913
R21918 outputibias.n16 outputibias.n9 1.16414
R21919 outputibias.n47 outputibias.n40 1.16414
R21920 outputibias.n79 outputibias.n72 1.16414
R21921 outputibias.n111 outputibias.n104 1.16414
R21922 outputibias.n127 outputibias.n95 0.962709
R21923 outputibias.n95 outputibias.n63 0.962709
R21924 outputibias.n13 outputibias.n12 0.388379
R21925 outputibias.n44 outputibias.n43 0.388379
R21926 outputibias.n76 outputibias.n75 0.388379
R21927 outputibias.n108 outputibias.n107 0.388379
R21928 outputibias.n134 outputibias.n0 0.337251
R21929 outputibias outputibias.n134 0.302375
R21930 outputibias.n30 outputibias.n2 0.155672
R21931 outputibias.n23 outputibias.n2 0.155672
R21932 outputibias.n23 outputibias.n22 0.155672
R21933 outputibias.n22 outputibias.n6 0.155672
R21934 outputibias.n15 outputibias.n6 0.155672
R21935 outputibias.n15 outputibias.n14 0.155672
R21936 outputibias.n61 outputibias.n33 0.155672
R21937 outputibias.n54 outputibias.n33 0.155672
R21938 outputibias.n54 outputibias.n53 0.155672
R21939 outputibias.n53 outputibias.n37 0.155672
R21940 outputibias.n46 outputibias.n37 0.155672
R21941 outputibias.n46 outputibias.n45 0.155672
R21942 outputibias.n93 outputibias.n65 0.155672
R21943 outputibias.n86 outputibias.n65 0.155672
R21944 outputibias.n86 outputibias.n85 0.155672
R21945 outputibias.n85 outputibias.n69 0.155672
R21946 outputibias.n78 outputibias.n69 0.155672
R21947 outputibias.n78 outputibias.n77 0.155672
R21948 outputibias.n125 outputibias.n97 0.155672
R21949 outputibias.n118 outputibias.n97 0.155672
R21950 outputibias.n118 outputibias.n117 0.155672
R21951 outputibias.n117 outputibias.n101 0.155672
R21952 outputibias.n110 outputibias.n101 0.155672
R21953 outputibias.n110 outputibias.n109 0.155672
C0 commonsourceibias diffpairibias 0.06482f
C1 minus plus 9.171639f
C2 CSoutput commonsourceibias 54.0646f
C3 minus commonsourceibias 0.323289f
C4 plus commonsourceibias 0.277692f
C5 output outputibias 2.34152f
C6 vdd output 7.23429f
C7 CSoutput output 6.13881f
C8 CSoutput outputibias 0.032386f
C9 vdd CSoutput 67.6707f
C10 minus diffpairibias 3.46e-19
C11 commonsourceibias output 0.006808f
C12 vdd plus 0.065956f
C13 CSoutput minus 2.77524f
C14 plus diffpairibias 2.47e-19
C15 commonsourceibias outputibias 0.003832f
C16 vdd commonsourceibias 0.004218f
C17 CSoutput plus 0.856907f
C18 diffpairibias gnd 48.980137f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.183542p
C22 plus gnd 32.72864f
C23 minus gnd 27.03175f
C24 CSoutput gnd 0.12555p
C25 vdd gnd 0.345104p
C26 outputibias.t9 gnd 0.11477f
C27 outputibias.t10 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t7 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t1 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t3 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t5 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t4 gnd 0.108319f
C161 outputibias.t2 gnd 0.108319f
C162 outputibias.t0 gnd 0.108319f
C163 outputibias.t6 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t11 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t8 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 diffpairibias.t18 gnd 0.087401f
C174 diffpairibias.t22 gnd 0.087239f
C175 diffpairibias.n0 gnd 0.102784f
C176 diffpairibias.t20 gnd 0.087239f
C177 diffpairibias.n1 gnd 0.050171f
C178 diffpairibias.t23 gnd 0.087239f
C179 diffpairibias.n2 gnd 0.039841f
C180 diffpairibias.t1 gnd 0.083757f
C181 diffpairibias.t9 gnd 0.083392f
C182 diffpairibias.n3 gnd 0.131682f
C183 diffpairibias.t11 gnd 0.083392f
C184 diffpairibias.n4 gnd 0.07027f
C185 diffpairibias.t7 gnd 0.083392f
C186 diffpairibias.n5 gnd 0.07027f
C187 diffpairibias.t3 gnd 0.083392f
C188 diffpairibias.n6 gnd 0.07027f
C189 diffpairibias.t13 gnd 0.083392f
C190 diffpairibias.n7 gnd 0.07027f
C191 diffpairibias.t5 gnd 0.083392f
C192 diffpairibias.n8 gnd 0.07027f
C193 diffpairibias.t15 gnd 0.083392f
C194 diffpairibias.n9 gnd 0.099771f
C195 diffpairibias.t0 gnd 0.08427f
C196 diffpairibias.t8 gnd 0.084123f
C197 diffpairibias.n10 gnd 0.091784f
C198 diffpairibias.t10 gnd 0.084123f
C199 diffpairibias.n11 gnd 0.050681f
C200 diffpairibias.t6 gnd 0.084123f
C201 diffpairibias.n12 gnd 0.050681f
C202 diffpairibias.t2 gnd 0.084123f
C203 diffpairibias.n13 gnd 0.050681f
C204 diffpairibias.t12 gnd 0.084123f
C205 diffpairibias.n14 gnd 0.050681f
C206 diffpairibias.t4 gnd 0.084123f
C207 diffpairibias.n15 gnd 0.050681f
C208 diffpairibias.t14 gnd 0.084123f
C209 diffpairibias.n16 gnd 0.059977f
C210 diffpairibias.n17 gnd 0.226448f
C211 diffpairibias.t21 gnd 0.087239f
C212 diffpairibias.n18 gnd 0.050181f
C213 diffpairibias.t17 gnd 0.087239f
C214 diffpairibias.n19 gnd 0.050171f
C215 diffpairibias.t16 gnd 0.087239f
C216 diffpairibias.n20 gnd 0.050171f
C217 diffpairibias.t19 gnd 0.087239f
C218 diffpairibias.n21 gnd 0.045859f
C219 diffpairibias.n22 gnd 0.046268f
C220 output.t5 gnd 0.464308f
C221 output.t10 gnd 0.044422f
C222 output.t15 gnd 0.044422f
C223 output.n0 gnd 0.364624f
C224 output.n1 gnd 0.614102f
C225 output.t3 gnd 0.044422f
C226 output.t11 gnd 0.044422f
C227 output.n2 gnd 0.364624f
C228 output.n3 gnd 0.350265f
C229 output.t14 gnd 0.044422f
C230 output.t12 gnd 0.044422f
C231 output.n4 gnd 0.364624f
C232 output.n5 gnd 0.350265f
C233 output.t18 gnd 0.044422f
C234 output.t4 gnd 0.044422f
C235 output.n6 gnd 0.364624f
C236 output.n7 gnd 0.350265f
C237 output.t7 gnd 0.044422f
C238 output.t16 gnd 0.044422f
C239 output.n8 gnd 0.364624f
C240 output.n9 gnd 0.350265f
C241 output.t17 gnd 0.044422f
C242 output.t8 gnd 0.044422f
C243 output.n10 gnd 0.364624f
C244 output.n11 gnd 0.350265f
C245 output.t9 gnd 0.044422f
C246 output.t13 gnd 0.044422f
C247 output.n12 gnd 0.364624f
C248 output.n13 gnd 0.350265f
C249 output.t6 gnd 0.462979f
C250 output.n14 gnd 0.28994f
C251 output.n15 gnd 0.015803f
C252 output.n16 gnd 0.011243f
C253 output.n17 gnd 0.006041f
C254 output.n18 gnd 0.01428f
C255 output.n19 gnd 0.006397f
C256 output.n20 gnd 0.011243f
C257 output.n21 gnd 0.006041f
C258 output.n22 gnd 0.01428f
C259 output.n23 gnd 0.006397f
C260 output.n24 gnd 0.048111f
C261 output.t0 gnd 0.023274f
C262 output.n25 gnd 0.01071f
C263 output.n26 gnd 0.008435f
C264 output.n27 gnd 0.006041f
C265 output.n28 gnd 0.267512f
C266 output.n29 gnd 0.011243f
C267 output.n30 gnd 0.006041f
C268 output.n31 gnd 0.006397f
C269 output.n32 gnd 0.01428f
C270 output.n33 gnd 0.01428f
C271 output.n34 gnd 0.006397f
C272 output.n35 gnd 0.006041f
C273 output.n36 gnd 0.011243f
C274 output.n37 gnd 0.011243f
C275 output.n38 gnd 0.006041f
C276 output.n39 gnd 0.006397f
C277 output.n40 gnd 0.01428f
C278 output.n41 gnd 0.030913f
C279 output.n42 gnd 0.006397f
C280 output.n43 gnd 0.006041f
C281 output.n44 gnd 0.025987f
C282 output.n45 gnd 0.097665f
C283 output.n46 gnd 0.015803f
C284 output.n47 gnd 0.011243f
C285 output.n48 gnd 0.006041f
C286 output.n49 gnd 0.01428f
C287 output.n50 gnd 0.006397f
C288 output.n51 gnd 0.011243f
C289 output.n52 gnd 0.006041f
C290 output.n53 gnd 0.01428f
C291 output.n54 gnd 0.006397f
C292 output.n55 gnd 0.048111f
C293 output.t19 gnd 0.023274f
C294 output.n56 gnd 0.01071f
C295 output.n57 gnd 0.008435f
C296 output.n58 gnd 0.006041f
C297 output.n59 gnd 0.267512f
C298 output.n60 gnd 0.011243f
C299 output.n61 gnd 0.006041f
C300 output.n62 gnd 0.006397f
C301 output.n63 gnd 0.01428f
C302 output.n64 gnd 0.01428f
C303 output.n65 gnd 0.006397f
C304 output.n66 gnd 0.006041f
C305 output.n67 gnd 0.011243f
C306 output.n68 gnd 0.011243f
C307 output.n69 gnd 0.006041f
C308 output.n70 gnd 0.006397f
C309 output.n71 gnd 0.01428f
C310 output.n72 gnd 0.030913f
C311 output.n73 gnd 0.006397f
C312 output.n74 gnd 0.006041f
C313 output.n75 gnd 0.025987f
C314 output.n76 gnd 0.09306f
C315 output.n77 gnd 1.65264f
C316 output.n78 gnd 0.015803f
C317 output.n79 gnd 0.011243f
C318 output.n80 gnd 0.006041f
C319 output.n81 gnd 0.01428f
C320 output.n82 gnd 0.006397f
C321 output.n83 gnd 0.011243f
C322 output.n84 gnd 0.006041f
C323 output.n85 gnd 0.01428f
C324 output.n86 gnd 0.006397f
C325 output.n87 gnd 0.048111f
C326 output.t2 gnd 0.023274f
C327 output.n88 gnd 0.01071f
C328 output.n89 gnd 0.008435f
C329 output.n90 gnd 0.006041f
C330 output.n91 gnd 0.267512f
C331 output.n92 gnd 0.011243f
C332 output.n93 gnd 0.006041f
C333 output.n94 gnd 0.006397f
C334 output.n95 gnd 0.01428f
C335 output.n96 gnd 0.01428f
C336 output.n97 gnd 0.006397f
C337 output.n98 gnd 0.006041f
C338 output.n99 gnd 0.011243f
C339 output.n100 gnd 0.011243f
C340 output.n101 gnd 0.006041f
C341 output.n102 gnd 0.006397f
C342 output.n103 gnd 0.01428f
C343 output.n104 gnd 0.030913f
C344 output.n105 gnd 0.006397f
C345 output.n106 gnd 0.006041f
C346 output.n107 gnd 0.025987f
C347 output.n108 gnd 0.09306f
C348 output.n109 gnd 0.713089f
C349 output.n110 gnd 0.015803f
C350 output.n111 gnd 0.011243f
C351 output.n112 gnd 0.006041f
C352 output.n113 gnd 0.01428f
C353 output.n114 gnd 0.006397f
C354 output.n115 gnd 0.011243f
C355 output.n116 gnd 0.006041f
C356 output.n117 gnd 0.01428f
C357 output.n118 gnd 0.006397f
C358 output.n119 gnd 0.048111f
C359 output.t1 gnd 0.023274f
C360 output.n120 gnd 0.01071f
C361 output.n121 gnd 0.008435f
C362 output.n122 gnd 0.006041f
C363 output.n123 gnd 0.267512f
C364 output.n124 gnd 0.011243f
C365 output.n125 gnd 0.006041f
C366 output.n126 gnd 0.006397f
C367 output.n127 gnd 0.01428f
C368 output.n128 gnd 0.01428f
C369 output.n129 gnd 0.006397f
C370 output.n130 gnd 0.006041f
C371 output.n131 gnd 0.011243f
C372 output.n132 gnd 0.011243f
C373 output.n133 gnd 0.006041f
C374 output.n134 gnd 0.006397f
C375 output.n135 gnd 0.01428f
C376 output.n136 gnd 0.030913f
C377 output.n137 gnd 0.006397f
C378 output.n138 gnd 0.006041f
C379 output.n139 gnd 0.025987f
C380 output.n140 gnd 0.09306f
C381 output.n141 gnd 1.67353f
C382 minus.n0 gnd 0.030059f
C383 minus.t14 gnd 0.505432f
C384 minus.n1 gnd 0.204419f
C385 minus.n2 gnd 0.030059f
C386 minus.t19 gnd 0.505432f
C387 minus.n3 gnd 0.024431f
C388 minus.n4 gnd 0.030059f
C389 minus.t18 gnd 0.505432f
C390 minus.t5 gnd 0.505432f
C391 minus.n5 gnd 0.204419f
C392 minus.n6 gnd 0.030059f
C393 minus.t8 gnd 0.505432f
C394 minus.n7 gnd 0.204419f
C395 minus.n8 gnd 0.12903f
C396 minus.t9 gnd 0.505432f
C397 minus.t13 gnd 0.567467f
C398 minus.n9 gnd 0.237182f
C399 minus.n10 gnd 0.236072f
C400 minus.n11 gnd 0.03739f
C401 minus.n12 gnd 0.03514f
C402 minus.n13 gnd 0.030059f
C403 minus.n14 gnd 0.030059f
C404 minus.n15 gnd 0.037653f
C405 minus.n16 gnd 0.024431f
C406 minus.n17 gnd 0.038669f
C407 minus.n18 gnd 0.030059f
C408 minus.n19 gnd 0.030059f
C409 minus.n20 gnd 0.036265f
C410 minus.n21 gnd 0.036265f
C411 minus.n22 gnd 0.204419f
C412 minus.n23 gnd 0.038669f
C413 minus.n24 gnd 0.030059f
C414 minus.n25 gnd 0.030059f
C415 minus.n26 gnd 0.030059f
C416 minus.n27 gnd 0.037653f
C417 minus.n28 gnd 0.204419f
C418 minus.n29 gnd 0.03514f
C419 minus.n30 gnd 0.03739f
C420 minus.n31 gnd 0.030059f
C421 minus.n32 gnd 0.030059f
C422 minus.n33 gnd 0.039147f
C423 minus.n34 gnd 0.01245f
C424 minus.t17 gnd 0.546625f
C425 minus.n35 gnd 0.237424f
C426 minus.n36 gnd 0.353195f
C427 minus.n37 gnd 0.030059f
C428 minus.t15 gnd 0.546625f
C429 minus.t12 gnd 0.505432f
C430 minus.n38 gnd 0.204419f
C431 minus.n39 gnd 0.030059f
C432 minus.t7 gnd 0.505432f
C433 minus.n40 gnd 0.024431f
C434 minus.n41 gnd 0.030059f
C435 minus.t6 gnd 0.505432f
C436 minus.t11 gnd 0.505432f
C437 minus.n42 gnd 0.204419f
C438 minus.n43 gnd 0.030059f
C439 minus.t10 gnd 0.505432f
C440 minus.n44 gnd 0.204419f
C441 minus.n45 gnd 0.12903f
C442 minus.t16 gnd 0.505432f
C443 minus.t20 gnd 0.567467f
C444 minus.n46 gnd 0.237182f
C445 minus.n47 gnd 0.236072f
C446 minus.n48 gnd 0.03739f
C447 minus.n49 gnd 0.03514f
C448 minus.n50 gnd 0.030059f
C449 minus.n51 gnd 0.030059f
C450 minus.n52 gnd 0.037653f
C451 minus.n53 gnd 0.024431f
C452 minus.n54 gnd 0.038669f
C453 minus.n55 gnd 0.030059f
C454 minus.n56 gnd 0.030059f
C455 minus.n57 gnd 0.036265f
C456 minus.n58 gnd 0.036265f
C457 minus.n59 gnd 0.204419f
C458 minus.n60 gnd 0.038669f
C459 minus.n61 gnd 0.030059f
C460 minus.n62 gnd 0.030059f
C461 minus.n63 gnd 0.030059f
C462 minus.n64 gnd 0.037653f
C463 minus.n65 gnd 0.204419f
C464 minus.n66 gnd 0.03514f
C465 minus.n67 gnd 0.03739f
C466 minus.n68 gnd 0.030059f
C467 minus.n69 gnd 0.030059f
C468 minus.n70 gnd 0.039147f
C469 minus.n71 gnd 0.01245f
C470 minus.n72 gnd 0.237424f
C471 minus.n73 gnd 0.936615f
C472 minus.n74 gnd 1.40781f
C473 minus.t1 gnd 0.009266f
C474 minus.t4 gnd 0.009266f
C475 minus.n75 gnd 0.030469f
C476 minus.t2 gnd 0.009266f
C477 minus.t0 gnd 0.009266f
C478 minus.n76 gnd 0.030052f
C479 minus.n77 gnd 0.25648f
C480 minus.t3 gnd 0.051575f
C481 minus.n78 gnd 0.139959f
C482 minus.n79 gnd 1.89864f
C483 a_n2903_n3924.n0 gnd 1.45586f
C484 a_n2903_n3924.t24 gnd 0.088483f
C485 a_n2903_n3924.t33 gnd 0.919619f
C486 a_n2903_n3924.n1 gnd 0.347657f
C487 a_n2903_n3924.t3 gnd 1.14306f
C488 a_n2903_n3924.n2 gnd 1.19083f
C489 a_n2903_n3924.t19 gnd 0.919619f
C490 a_n2903_n3924.n3 gnd 0.347657f
C491 a_n2903_n3924.t8 gnd 0.088483f
C492 a_n2903_n3924.t21 gnd 0.088483f
C493 a_n2903_n3924.n4 gnd 0.722655f
C494 a_n2903_n3924.n5 gnd 0.364177f
C495 a_n2903_n3924.t6 gnd 0.088483f
C496 a_n2903_n3924.t16 gnd 0.088483f
C497 a_n2903_n3924.n6 gnd 0.722655f
C498 a_n2903_n3924.n7 gnd 0.364177f
C499 a_n2903_n3924.t11 gnd 0.088483f
C500 a_n2903_n3924.t10 gnd 0.088483f
C501 a_n2903_n3924.n8 gnd 0.722655f
C502 a_n2903_n3924.n9 gnd 0.364177f
C503 a_n2903_n3924.t18 gnd 0.919619f
C504 a_n2903_n3924.n10 gnd 0.860834f
C505 a_n2903_n3924.t39 gnd 1.14419f
C506 a_n2903_n3924.t5 gnd 1.14261f
C507 a_n2903_n3924.n11 gnd 0.745791f
C508 a_n2903_n3924.t0 gnd 1.14261f
C509 a_n2903_n3924.n12 gnd 0.804757f
C510 a_n2903_n3924.t38 gnd 1.14261f
C511 a_n2903_n3924.n13 gnd 0.804757f
C512 a_n2903_n3924.t1 gnd 1.14261f
C513 a_n2903_n3924.n14 gnd 0.804757f
C514 a_n2903_n3924.t2 gnd 1.14261f
C515 a_n2903_n3924.n15 gnd 0.804757f
C516 a_n2903_n3924.t4 gnd 1.14261f
C517 a_n2903_n3924.n16 gnd 0.834168f
C518 a_n2903_n3924.t35 gnd 0.919616f
C519 a_n2903_n3924.n17 gnd 0.571219f
C520 a_n2903_n3924.t36 gnd 0.088483f
C521 a_n2903_n3924.t26 gnd 0.088483f
C522 a_n2903_n3924.n18 gnd 0.722654f
C523 a_n2903_n3924.n19 gnd 0.364178f
C524 a_n2903_n3924.t27 gnd 0.088483f
C525 a_n2903_n3924.t22 gnd 0.088483f
C526 a_n2903_n3924.n20 gnd 0.722654f
C527 a_n2903_n3924.n21 gnd 0.364178f
C528 a_n2903_n3924.t23 gnd 0.088483f
C529 a_n2903_n3924.t34 gnd 0.088483f
C530 a_n2903_n3924.n22 gnd 0.722654f
C531 a_n2903_n3924.n23 gnd 0.364178f
C532 a_n2903_n3924.t31 gnd 0.919616f
C533 a_n2903_n3924.n24 gnd 0.347661f
C534 a_n2903_n3924.t15 gnd 0.919616f
C535 a_n2903_n3924.n25 gnd 0.347661f
C536 a_n2903_n3924.t9 gnd 0.088483f
C537 a_n2903_n3924.t17 gnd 0.088483f
C538 a_n2903_n3924.n26 gnd 0.722654f
C539 a_n2903_n3924.n27 gnd 0.364178f
C540 a_n2903_n3924.t7 gnd 0.088483f
C541 a_n2903_n3924.t12 gnd 0.088483f
C542 a_n2903_n3924.n28 gnd 0.722654f
C543 a_n2903_n3924.n29 gnd 0.364178f
C544 a_n2903_n3924.t20 gnd 0.088483f
C545 a_n2903_n3924.t14 gnd 0.088483f
C546 a_n2903_n3924.n30 gnd 0.722654f
C547 a_n2903_n3924.n31 gnd 0.364178f
C548 a_n2903_n3924.t13 gnd 0.919616f
C549 a_n2903_n3924.n32 gnd 0.571219f
C550 a_n2903_n3924.n33 gnd 0.834168f
C551 a_n2903_n3924.t30 gnd 0.919616f
C552 a_n2903_n3924.n34 gnd 0.860837f
C553 a_n2903_n3924.t28 gnd 0.088483f
C554 a_n2903_n3924.t32 gnd 0.088483f
C555 a_n2903_n3924.n35 gnd 0.722655f
C556 a_n2903_n3924.n36 gnd 0.364177f
C557 a_n2903_n3924.t25 gnd 0.088483f
C558 a_n2903_n3924.t29 gnd 0.088483f
C559 a_n2903_n3924.n37 gnd 0.722655f
C560 a_n2903_n3924.n38 gnd 0.364177f
C561 a_n2903_n3924.n39 gnd 0.364176f
C562 a_n2903_n3924.n40 gnd 0.722656f
C563 a_n2903_n3924.t37 gnd 0.088483f
C564 plus.n0 gnd 0.022051f
C565 plus.t7 gnd 0.401003f
C566 plus.t6 gnd 0.370784f
C567 plus.n1 gnd 0.149962f
C568 plus.n2 gnd 0.022051f
C569 plus.t16 gnd 0.370784f
C570 plus.n3 gnd 0.017923f
C571 plus.n4 gnd 0.022051f
C572 plus.t15 gnd 0.370784f
C573 plus.t20 gnd 0.370784f
C574 plus.n5 gnd 0.149962f
C575 plus.n6 gnd 0.022051f
C576 plus.t19 gnd 0.370784f
C577 plus.n7 gnd 0.149962f
C578 plus.n8 gnd 0.094656f
C579 plus.t8 gnd 0.370784f
C580 plus.t11 gnd 0.416293f
C581 plus.n9 gnd 0.173997f
C582 plus.n10 gnd 0.173182f
C583 plus.n11 gnd 0.02743f
C584 plus.n12 gnd 0.025779f
C585 plus.n13 gnd 0.022051f
C586 plus.n14 gnd 0.022051f
C587 plus.n15 gnd 0.027622f
C588 plus.n16 gnd 0.017923f
C589 plus.n17 gnd 0.028368f
C590 plus.n18 gnd 0.022051f
C591 plus.n19 gnd 0.022051f
C592 plus.n20 gnd 0.026604f
C593 plus.n21 gnd 0.026604f
C594 plus.n22 gnd 0.149962f
C595 plus.n23 gnd 0.028368f
C596 plus.n24 gnd 0.022051f
C597 plus.n25 gnd 0.022051f
C598 plus.n26 gnd 0.022051f
C599 plus.n27 gnd 0.027622f
C600 plus.n28 gnd 0.149962f
C601 plus.n29 gnd 0.025779f
C602 plus.n30 gnd 0.02743f
C603 plus.n31 gnd 0.022051f
C604 plus.n32 gnd 0.022051f
C605 plus.n33 gnd 0.028719f
C606 plus.n34 gnd 0.009133f
C607 plus.n35 gnd 0.174174f
C608 plus.n36 gnd 0.253432f
C609 plus.n37 gnd 0.022051f
C610 plus.t10 gnd 0.370784f
C611 plus.n38 gnd 0.149962f
C612 plus.n39 gnd 0.022051f
C613 plus.t14 gnd 0.370784f
C614 plus.n40 gnd 0.017923f
C615 plus.n41 gnd 0.022051f
C616 plus.t13 gnd 0.370784f
C617 plus.t17 gnd 0.370784f
C618 plus.n42 gnd 0.149962f
C619 plus.n43 gnd 0.022051f
C620 plus.t18 gnd 0.370784f
C621 plus.n44 gnd 0.149962f
C622 plus.n45 gnd 0.094656f
C623 plus.t5 gnd 0.370784f
C624 plus.t9 gnd 0.416293f
C625 plus.n46 gnd 0.173997f
C626 plus.n47 gnd 0.173182f
C627 plus.n48 gnd 0.02743f
C628 plus.n49 gnd 0.025779f
C629 plus.n50 gnd 0.022051f
C630 plus.n51 gnd 0.022051f
C631 plus.n52 gnd 0.027622f
C632 plus.n53 gnd 0.017923f
C633 plus.n54 gnd 0.028368f
C634 plus.n55 gnd 0.022051f
C635 plus.n56 gnd 0.022051f
C636 plus.n57 gnd 0.026604f
C637 plus.n58 gnd 0.026604f
C638 plus.n59 gnd 0.149962f
C639 plus.n60 gnd 0.028368f
C640 plus.n61 gnd 0.022051f
C641 plus.n62 gnd 0.022051f
C642 plus.n63 gnd 0.022051f
C643 plus.n64 gnd 0.027622f
C644 plus.n65 gnd 0.149962f
C645 plus.n66 gnd 0.025779f
C646 plus.n67 gnd 0.02743f
C647 plus.n68 gnd 0.022051f
C648 plus.n69 gnd 0.022051f
C649 plus.n70 gnd 0.028719f
C650 plus.n71 gnd 0.009133f
C651 plus.t12 gnd 0.401003f
C652 plus.n72 gnd 0.174174f
C653 plus.n73 gnd 0.678265f
C654 plus.n74 gnd 1.02402f
C655 plus.t4 gnd 0.038066f
C656 plus.t1 gnd 0.006798f
C657 plus.t2 gnd 0.006798f
C658 plus.n75 gnd 0.022046f
C659 plus.n76 gnd 0.171146f
C660 plus.t0 gnd 0.006798f
C661 plus.t3 gnd 0.006798f
C662 plus.n77 gnd 0.022046f
C663 plus.n78 gnd 0.128466f
C664 plus.n79 gnd 2.48089f
C665 a_n1986_8322.t0 gnd 49.3562f
C666 a_n1986_8322.t1 gnd 75.4844f
C667 a_n1986_8322.t11 gnd 0.875761f
C668 a_n1986_8322.t19 gnd 0.093529f
C669 a_n1986_8322.t14 gnd 0.093529f
C670 a_n1986_8322.n0 gnd 0.65882f
C671 a_n1986_8322.n1 gnd 0.736135f
C672 a_n1986_8322.t17 gnd 0.093529f
C673 a_n1986_8322.t16 gnd 0.093529f
C674 a_n1986_8322.n2 gnd 0.65882f
C675 a_n1986_8322.n3 gnd 0.374021f
C676 a_n1986_8322.t10 gnd 0.874017f
C677 a_n1986_8322.n4 gnd 1.39891f
C678 a_n1986_8322.t5 gnd 0.875761f
C679 a_n1986_8322.t8 gnd 0.093529f
C680 a_n1986_8322.t9 gnd 0.093529f
C681 a_n1986_8322.n5 gnd 0.65882f
C682 a_n1986_8322.n6 gnd 0.736135f
C683 a_n1986_8322.t3 gnd 0.874017f
C684 a_n1986_8322.n7 gnd 0.370433f
C685 a_n1986_8322.t6 gnd 0.874017f
C686 a_n1986_8322.n8 gnd 0.370433f
C687 a_n1986_8322.t4 gnd 0.093529f
C688 a_n1986_8322.t2 gnd 0.093529f
C689 a_n1986_8322.n9 gnd 0.65882f
C690 a_n1986_8322.n10 gnd 0.374021f
C691 a_n1986_8322.t7 gnd 0.874017f
C692 a_n1986_8322.n11 gnd 0.872286f
C693 a_n1986_8322.n12 gnd 1.59065f
C694 a_n1986_8322.n13 gnd 3.48702f
C695 a_n1986_8322.t12 gnd 0.874017f
C696 a_n1986_8322.n14 gnd 0.766493f
C697 a_n1986_8322.t13 gnd 0.093529f
C698 a_n1986_8322.t21 gnd 0.093529f
C699 a_n1986_8322.n15 gnd 0.65882f
C700 a_n1986_8322.n16 gnd 0.374021f
C701 a_n1986_8322.t18 gnd 0.093529f
C702 a_n1986_8322.t15 gnd 0.093529f
C703 a_n1986_8322.n17 gnd 0.65882f
C704 a_n1986_8322.n18 gnd 0.736133f
C705 a_n1986_8322.t20 gnd 0.875763f
C706 commonsourceibias.n0 gnd 0.012624f
C707 commonsourceibias.t120 gnd 0.191163f
C708 commonsourceibias.t65 gnd 0.176757f
C709 commonsourceibias.n1 gnd 0.00769f
C710 commonsourceibias.n2 gnd 0.009461f
C711 commonsourceibias.t126 gnd 0.176757f
C712 commonsourceibias.n3 gnd 0.009597f
C713 commonsourceibias.n4 gnd 0.009461f
C714 commonsourceibias.t121 gnd 0.176757f
C715 commonsourceibias.n5 gnd 0.070526f
C716 commonsourceibias.t135 gnd 0.176757f
C717 commonsourceibias.n6 gnd 0.007653f
C718 commonsourceibias.n7 gnd 0.009461f
C719 commonsourceibias.t117 gnd 0.176757f
C720 commonsourceibias.n8 gnd 0.009134f
C721 commonsourceibias.n9 gnd 0.009461f
C722 commonsourceibias.t102 gnd 0.176757f
C723 commonsourceibias.n10 gnd 0.070526f
C724 commonsourceibias.t125 gnd 0.176757f
C725 commonsourceibias.n11 gnd 0.007641f
C726 commonsourceibias.n12 gnd 0.012624f
C727 commonsourceibias.t20 gnd 0.191163f
C728 commonsourceibias.t48 gnd 0.176757f
C729 commonsourceibias.n13 gnd 0.00769f
C730 commonsourceibias.n14 gnd 0.009461f
C731 commonsourceibias.t30 gnd 0.176757f
C732 commonsourceibias.n15 gnd 0.009597f
C733 commonsourceibias.n16 gnd 0.009461f
C734 commonsourceibias.t6 gnd 0.176757f
C735 commonsourceibias.n17 gnd 0.070526f
C736 commonsourceibias.t28 gnd 0.176757f
C737 commonsourceibias.n18 gnd 0.007653f
C738 commonsourceibias.n19 gnd 0.009461f
C739 commonsourceibias.t24 gnd 0.176757f
C740 commonsourceibias.n20 gnd 0.009134f
C741 commonsourceibias.n21 gnd 0.009461f
C742 commonsourceibias.t52 gnd 0.176757f
C743 commonsourceibias.n22 gnd 0.070526f
C744 commonsourceibias.t32 gnd 0.176757f
C745 commonsourceibias.n23 gnd 0.007641f
C746 commonsourceibias.n24 gnd 0.009461f
C747 commonsourceibias.t22 gnd 0.176757f
C748 commonsourceibias.t42 gnd 0.176757f
C749 commonsourceibias.n25 gnd 0.070526f
C750 commonsourceibias.n26 gnd 0.009461f
C751 commonsourceibias.t2 gnd 0.176757f
C752 commonsourceibias.n27 gnd 0.070526f
C753 commonsourceibias.n28 gnd 0.009461f
C754 commonsourceibias.t56 gnd 0.176757f
C755 commonsourceibias.n29 gnd 0.070526f
C756 commonsourceibias.n30 gnd 0.009461f
C757 commonsourceibias.t8 gnd 0.176757f
C758 commonsourceibias.n31 gnd 0.010754f
C759 commonsourceibias.n32 gnd 0.009461f
C760 commonsourceibias.t10 gnd 0.176757f
C761 commonsourceibias.n33 gnd 0.012717f
C762 commonsourceibias.t16 gnd 0.196904f
C763 commonsourceibias.t50 gnd 0.176757f
C764 commonsourceibias.n34 gnd 0.078584f
C765 commonsourceibias.n35 gnd 0.084191f
C766 commonsourceibias.n36 gnd 0.04027f
C767 commonsourceibias.n37 gnd 0.009461f
C768 commonsourceibias.n38 gnd 0.00769f
C769 commonsourceibias.n39 gnd 0.013037f
C770 commonsourceibias.n40 gnd 0.070526f
C771 commonsourceibias.n41 gnd 0.013093f
C772 commonsourceibias.n42 gnd 0.009461f
C773 commonsourceibias.n43 gnd 0.009461f
C774 commonsourceibias.n44 gnd 0.009461f
C775 commonsourceibias.n45 gnd 0.009597f
C776 commonsourceibias.n46 gnd 0.070526f
C777 commonsourceibias.n47 gnd 0.011661f
C778 commonsourceibias.n48 gnd 0.0129f
C779 commonsourceibias.n49 gnd 0.009461f
C780 commonsourceibias.n50 gnd 0.009461f
C781 commonsourceibias.n51 gnd 0.012816f
C782 commonsourceibias.n52 gnd 0.007653f
C783 commonsourceibias.n53 gnd 0.012975f
C784 commonsourceibias.n54 gnd 0.009461f
C785 commonsourceibias.n55 gnd 0.009461f
C786 commonsourceibias.n56 gnd 0.013054f
C787 commonsourceibias.n57 gnd 0.011256f
C788 commonsourceibias.n58 gnd 0.009134f
C789 commonsourceibias.n59 gnd 0.009461f
C790 commonsourceibias.n60 gnd 0.009461f
C791 commonsourceibias.n61 gnd 0.011572f
C792 commonsourceibias.n62 gnd 0.012989f
C793 commonsourceibias.n63 gnd 0.070526f
C794 commonsourceibias.n64 gnd 0.012901f
C795 commonsourceibias.n65 gnd 0.009461f
C796 commonsourceibias.n66 gnd 0.009461f
C797 commonsourceibias.n67 gnd 0.009461f
C798 commonsourceibias.n68 gnd 0.012901f
C799 commonsourceibias.n69 gnd 0.070526f
C800 commonsourceibias.n70 gnd 0.012989f
C801 commonsourceibias.n71 gnd 0.011572f
C802 commonsourceibias.n72 gnd 0.009461f
C803 commonsourceibias.n73 gnd 0.009461f
C804 commonsourceibias.n74 gnd 0.009461f
C805 commonsourceibias.n75 gnd 0.011256f
C806 commonsourceibias.n76 gnd 0.013054f
C807 commonsourceibias.n77 gnd 0.070526f
C808 commonsourceibias.n78 gnd 0.012975f
C809 commonsourceibias.n79 gnd 0.009461f
C810 commonsourceibias.n80 gnd 0.009461f
C811 commonsourceibias.n81 gnd 0.009461f
C812 commonsourceibias.n82 gnd 0.012816f
C813 commonsourceibias.n83 gnd 0.070526f
C814 commonsourceibias.n84 gnd 0.0129f
C815 commonsourceibias.n85 gnd 0.011661f
C816 commonsourceibias.n86 gnd 0.009461f
C817 commonsourceibias.n87 gnd 0.009461f
C818 commonsourceibias.n88 gnd 0.009461f
C819 commonsourceibias.n89 gnd 0.010754f
C820 commonsourceibias.n90 gnd 0.013093f
C821 commonsourceibias.n91 gnd 0.070526f
C822 commonsourceibias.n92 gnd 0.013037f
C823 commonsourceibias.n93 gnd 0.009461f
C824 commonsourceibias.n94 gnd 0.009461f
C825 commonsourceibias.n95 gnd 0.009461f
C826 commonsourceibias.n96 gnd 0.012717f
C827 commonsourceibias.n97 gnd 0.070526f
C828 commonsourceibias.n98 gnd 0.012748f
C829 commonsourceibias.n99 gnd 0.085044f
C830 commonsourceibias.n100 gnd 0.095092f
C831 commonsourceibias.t21 gnd 0.020415f
C832 commonsourceibias.t49 gnd 0.020415f
C833 commonsourceibias.n101 gnd 0.180398f
C834 commonsourceibias.n102 gnd 0.156264f
C835 commonsourceibias.t31 gnd 0.020415f
C836 commonsourceibias.t7 gnd 0.020415f
C837 commonsourceibias.n103 gnd 0.180398f
C838 commonsourceibias.n104 gnd 0.082864f
C839 commonsourceibias.t29 gnd 0.020415f
C840 commonsourceibias.t25 gnd 0.020415f
C841 commonsourceibias.n105 gnd 0.180398f
C842 commonsourceibias.n106 gnd 0.082864f
C843 commonsourceibias.t53 gnd 0.020415f
C844 commonsourceibias.t33 gnd 0.020415f
C845 commonsourceibias.n107 gnd 0.180398f
C846 commonsourceibias.n108 gnd 0.069229f
C847 commonsourceibias.t51 gnd 0.020415f
C848 commonsourceibias.t17 gnd 0.020415f
C849 commonsourceibias.n109 gnd 0.181002f
C850 commonsourceibias.t9 gnd 0.020415f
C851 commonsourceibias.t11 gnd 0.020415f
C852 commonsourceibias.n110 gnd 0.180398f
C853 commonsourceibias.n111 gnd 0.168097f
C854 commonsourceibias.t3 gnd 0.020415f
C855 commonsourceibias.t57 gnd 0.020415f
C856 commonsourceibias.n112 gnd 0.180398f
C857 commonsourceibias.n113 gnd 0.082864f
C858 commonsourceibias.t23 gnd 0.020415f
C859 commonsourceibias.t43 gnd 0.020415f
C860 commonsourceibias.n114 gnd 0.180398f
C861 commonsourceibias.n115 gnd 0.069229f
C862 commonsourceibias.n116 gnd 0.083829f
C863 commonsourceibias.n117 gnd 0.009461f
C864 commonsourceibias.t119 gnd 0.176757f
C865 commonsourceibias.t79 gnd 0.176757f
C866 commonsourceibias.n118 gnd 0.070526f
C867 commonsourceibias.n119 gnd 0.009461f
C868 commonsourceibias.t106 gnd 0.176757f
C869 commonsourceibias.n120 gnd 0.070526f
C870 commonsourceibias.n121 gnd 0.009461f
C871 commonsourceibias.t96 gnd 0.176757f
C872 commonsourceibias.n122 gnd 0.070526f
C873 commonsourceibias.n123 gnd 0.009461f
C874 commonsourceibias.t141 gnd 0.176757f
C875 commonsourceibias.n124 gnd 0.010754f
C876 commonsourceibias.n125 gnd 0.009461f
C877 commonsourceibias.t116 gnd 0.176757f
C878 commonsourceibias.n126 gnd 0.012717f
C879 commonsourceibias.t129 gnd 0.196904f
C880 commonsourceibias.t152 gnd 0.176757f
C881 commonsourceibias.n127 gnd 0.078584f
C882 commonsourceibias.n128 gnd 0.084191f
C883 commonsourceibias.n129 gnd 0.04027f
C884 commonsourceibias.n130 gnd 0.009461f
C885 commonsourceibias.n131 gnd 0.00769f
C886 commonsourceibias.n132 gnd 0.013037f
C887 commonsourceibias.n133 gnd 0.070526f
C888 commonsourceibias.n134 gnd 0.013093f
C889 commonsourceibias.n135 gnd 0.009461f
C890 commonsourceibias.n136 gnd 0.009461f
C891 commonsourceibias.n137 gnd 0.009461f
C892 commonsourceibias.n138 gnd 0.009597f
C893 commonsourceibias.n139 gnd 0.070526f
C894 commonsourceibias.n140 gnd 0.011661f
C895 commonsourceibias.n141 gnd 0.0129f
C896 commonsourceibias.n142 gnd 0.009461f
C897 commonsourceibias.n143 gnd 0.009461f
C898 commonsourceibias.n144 gnd 0.012816f
C899 commonsourceibias.n145 gnd 0.007653f
C900 commonsourceibias.n146 gnd 0.012975f
C901 commonsourceibias.n147 gnd 0.009461f
C902 commonsourceibias.n148 gnd 0.009461f
C903 commonsourceibias.n149 gnd 0.013054f
C904 commonsourceibias.n150 gnd 0.011256f
C905 commonsourceibias.n151 gnd 0.009134f
C906 commonsourceibias.n152 gnd 0.009461f
C907 commonsourceibias.n153 gnd 0.009461f
C908 commonsourceibias.n154 gnd 0.011572f
C909 commonsourceibias.n155 gnd 0.012989f
C910 commonsourceibias.n156 gnd 0.070526f
C911 commonsourceibias.n157 gnd 0.012901f
C912 commonsourceibias.n158 gnd 0.009415f
C913 commonsourceibias.n159 gnd 0.06839f
C914 commonsourceibias.n160 gnd 0.009415f
C915 commonsourceibias.n161 gnd 0.012901f
C916 commonsourceibias.n162 gnd 0.070526f
C917 commonsourceibias.n163 gnd 0.012989f
C918 commonsourceibias.n164 gnd 0.011572f
C919 commonsourceibias.n165 gnd 0.009461f
C920 commonsourceibias.n166 gnd 0.009461f
C921 commonsourceibias.n167 gnd 0.009461f
C922 commonsourceibias.n168 gnd 0.011256f
C923 commonsourceibias.n169 gnd 0.013054f
C924 commonsourceibias.n170 gnd 0.070526f
C925 commonsourceibias.n171 gnd 0.012975f
C926 commonsourceibias.n172 gnd 0.009461f
C927 commonsourceibias.n173 gnd 0.009461f
C928 commonsourceibias.n174 gnd 0.009461f
C929 commonsourceibias.n175 gnd 0.012816f
C930 commonsourceibias.n176 gnd 0.070526f
C931 commonsourceibias.n177 gnd 0.0129f
C932 commonsourceibias.n178 gnd 0.011661f
C933 commonsourceibias.n179 gnd 0.009461f
C934 commonsourceibias.n180 gnd 0.009461f
C935 commonsourceibias.n181 gnd 0.009461f
C936 commonsourceibias.n182 gnd 0.010754f
C937 commonsourceibias.n183 gnd 0.013093f
C938 commonsourceibias.n184 gnd 0.070526f
C939 commonsourceibias.n185 gnd 0.013037f
C940 commonsourceibias.n186 gnd 0.009461f
C941 commonsourceibias.n187 gnd 0.009461f
C942 commonsourceibias.n188 gnd 0.009461f
C943 commonsourceibias.n189 gnd 0.012717f
C944 commonsourceibias.n190 gnd 0.070526f
C945 commonsourceibias.n191 gnd 0.012748f
C946 commonsourceibias.n192 gnd 0.085044f
C947 commonsourceibias.n193 gnd 0.056182f
C948 commonsourceibias.n194 gnd 0.012624f
C949 commonsourceibias.t68 gnd 0.191163f
C950 commonsourceibias.t159 gnd 0.176757f
C951 commonsourceibias.n195 gnd 0.00769f
C952 commonsourceibias.n196 gnd 0.009461f
C953 commonsourceibias.t148 gnd 0.176757f
C954 commonsourceibias.n197 gnd 0.009597f
C955 commonsourceibias.n198 gnd 0.009461f
C956 commonsourceibias.t78 gnd 0.176757f
C957 commonsourceibias.n199 gnd 0.070526f
C958 commonsourceibias.t158 gnd 0.176757f
C959 commonsourceibias.n200 gnd 0.007653f
C960 commonsourceibias.n201 gnd 0.009461f
C961 commonsourceibias.t85 gnd 0.176757f
C962 commonsourceibias.n202 gnd 0.009134f
C963 commonsourceibias.n203 gnd 0.009461f
C964 commonsourceibias.t77 gnd 0.176757f
C965 commonsourceibias.n204 gnd 0.070526f
C966 commonsourceibias.t157 gnd 0.176757f
C967 commonsourceibias.n205 gnd 0.007641f
C968 commonsourceibias.n206 gnd 0.009461f
C969 commonsourceibias.t94 gnd 0.176757f
C970 commonsourceibias.t113 gnd 0.176757f
C971 commonsourceibias.n207 gnd 0.070526f
C972 commonsourceibias.n208 gnd 0.009461f
C973 commonsourceibias.t156 gnd 0.176757f
C974 commonsourceibias.n209 gnd 0.070526f
C975 commonsourceibias.n210 gnd 0.009461f
C976 commonsourceibias.t92 gnd 0.176757f
C977 commonsourceibias.n211 gnd 0.070526f
C978 commonsourceibias.n212 gnd 0.009461f
C979 commonsourceibias.t109 gnd 0.176757f
C980 commonsourceibias.n213 gnd 0.010754f
C981 commonsourceibias.n214 gnd 0.009461f
C982 commonsourceibias.t105 gnd 0.176757f
C983 commonsourceibias.n215 gnd 0.012717f
C984 commonsourceibias.t108 gnd 0.196904f
C985 commonsourceibias.t91 gnd 0.176757f
C986 commonsourceibias.n216 gnd 0.078584f
C987 commonsourceibias.n217 gnd 0.084191f
C988 commonsourceibias.n218 gnd 0.04027f
C989 commonsourceibias.n219 gnd 0.009461f
C990 commonsourceibias.n220 gnd 0.00769f
C991 commonsourceibias.n221 gnd 0.013037f
C992 commonsourceibias.n222 gnd 0.070526f
C993 commonsourceibias.n223 gnd 0.013093f
C994 commonsourceibias.n224 gnd 0.009461f
C995 commonsourceibias.n225 gnd 0.009461f
C996 commonsourceibias.n226 gnd 0.009461f
C997 commonsourceibias.n227 gnd 0.009597f
C998 commonsourceibias.n228 gnd 0.070526f
C999 commonsourceibias.n229 gnd 0.011661f
C1000 commonsourceibias.n230 gnd 0.0129f
C1001 commonsourceibias.n231 gnd 0.009461f
C1002 commonsourceibias.n232 gnd 0.009461f
C1003 commonsourceibias.n233 gnd 0.012816f
C1004 commonsourceibias.n234 gnd 0.007653f
C1005 commonsourceibias.n235 gnd 0.012975f
C1006 commonsourceibias.n236 gnd 0.009461f
C1007 commonsourceibias.n237 gnd 0.009461f
C1008 commonsourceibias.n238 gnd 0.013054f
C1009 commonsourceibias.n239 gnd 0.011256f
C1010 commonsourceibias.n240 gnd 0.009134f
C1011 commonsourceibias.n241 gnd 0.009461f
C1012 commonsourceibias.n242 gnd 0.009461f
C1013 commonsourceibias.n243 gnd 0.011572f
C1014 commonsourceibias.n244 gnd 0.012989f
C1015 commonsourceibias.n245 gnd 0.070526f
C1016 commonsourceibias.n246 gnd 0.012901f
C1017 commonsourceibias.n247 gnd 0.009461f
C1018 commonsourceibias.n248 gnd 0.009461f
C1019 commonsourceibias.n249 gnd 0.009461f
C1020 commonsourceibias.n250 gnd 0.012901f
C1021 commonsourceibias.n251 gnd 0.070526f
C1022 commonsourceibias.n252 gnd 0.012989f
C1023 commonsourceibias.n253 gnd 0.011572f
C1024 commonsourceibias.n254 gnd 0.009461f
C1025 commonsourceibias.n255 gnd 0.009461f
C1026 commonsourceibias.n256 gnd 0.009461f
C1027 commonsourceibias.n257 gnd 0.011256f
C1028 commonsourceibias.n258 gnd 0.013054f
C1029 commonsourceibias.n259 gnd 0.070526f
C1030 commonsourceibias.n260 gnd 0.012975f
C1031 commonsourceibias.n261 gnd 0.009461f
C1032 commonsourceibias.n262 gnd 0.009461f
C1033 commonsourceibias.n263 gnd 0.009461f
C1034 commonsourceibias.n264 gnd 0.012816f
C1035 commonsourceibias.n265 gnd 0.070526f
C1036 commonsourceibias.n266 gnd 0.0129f
C1037 commonsourceibias.n267 gnd 0.011661f
C1038 commonsourceibias.n268 gnd 0.009461f
C1039 commonsourceibias.n269 gnd 0.009461f
C1040 commonsourceibias.n270 gnd 0.009461f
C1041 commonsourceibias.n271 gnd 0.010754f
C1042 commonsourceibias.n272 gnd 0.013093f
C1043 commonsourceibias.n273 gnd 0.070526f
C1044 commonsourceibias.n274 gnd 0.013037f
C1045 commonsourceibias.n275 gnd 0.009461f
C1046 commonsourceibias.n276 gnd 0.009461f
C1047 commonsourceibias.n277 gnd 0.009461f
C1048 commonsourceibias.n278 gnd 0.012717f
C1049 commonsourceibias.n279 gnd 0.070526f
C1050 commonsourceibias.n280 gnd 0.012748f
C1051 commonsourceibias.n281 gnd 0.085044f
C1052 commonsourceibias.n282 gnd 0.030348f
C1053 commonsourceibias.n283 gnd 0.15151f
C1054 commonsourceibias.n284 gnd 0.012624f
C1055 commonsourceibias.t75 gnd 0.176757f
C1056 commonsourceibias.n285 gnd 0.00769f
C1057 commonsourceibias.n286 gnd 0.009461f
C1058 commonsourceibias.t128 gnd 0.176757f
C1059 commonsourceibias.n287 gnd 0.009597f
C1060 commonsourceibias.n288 gnd 0.009461f
C1061 commonsourceibias.t124 gnd 0.176757f
C1062 commonsourceibias.n289 gnd 0.070526f
C1063 commonsourceibias.t155 gnd 0.176757f
C1064 commonsourceibias.n290 gnd 0.007653f
C1065 commonsourceibias.n291 gnd 0.009461f
C1066 commonsourceibias.t89 gnd 0.176757f
C1067 commonsourceibias.n292 gnd 0.009134f
C1068 commonsourceibias.n293 gnd 0.009461f
C1069 commonsourceibias.t118 gnd 0.176757f
C1070 commonsourceibias.n294 gnd 0.070526f
C1071 commonsourceibias.t146 gnd 0.176757f
C1072 commonsourceibias.n295 gnd 0.007641f
C1073 commonsourceibias.n296 gnd 0.009461f
C1074 commonsourceibias.t138 gnd 0.176757f
C1075 commonsourceibias.t64 gnd 0.176757f
C1076 commonsourceibias.n297 gnd 0.070526f
C1077 commonsourceibias.n298 gnd 0.009461f
C1078 commonsourceibias.t137 gnd 0.176757f
C1079 commonsourceibias.n299 gnd 0.070526f
C1080 commonsourceibias.n300 gnd 0.009461f
C1081 commonsourceibias.t133 gnd 0.176757f
C1082 commonsourceibias.n301 gnd 0.070526f
C1083 commonsourceibias.n302 gnd 0.009461f
C1084 commonsourceibias.t149 gnd 0.176757f
C1085 commonsourceibias.n303 gnd 0.010754f
C1086 commonsourceibias.n304 gnd 0.009461f
C1087 commonsourceibias.t76 gnd 0.176757f
C1088 commonsourceibias.n305 gnd 0.012717f
C1089 commonsourceibias.t139 gnd 0.196904f
C1090 commonsourceibias.t130 gnd 0.176757f
C1091 commonsourceibias.n306 gnd 0.078584f
C1092 commonsourceibias.n307 gnd 0.084191f
C1093 commonsourceibias.n308 gnd 0.04027f
C1094 commonsourceibias.n309 gnd 0.009461f
C1095 commonsourceibias.n310 gnd 0.00769f
C1096 commonsourceibias.n311 gnd 0.013037f
C1097 commonsourceibias.n312 gnd 0.070526f
C1098 commonsourceibias.n313 gnd 0.013093f
C1099 commonsourceibias.n314 gnd 0.009461f
C1100 commonsourceibias.n315 gnd 0.009461f
C1101 commonsourceibias.n316 gnd 0.009461f
C1102 commonsourceibias.n317 gnd 0.009597f
C1103 commonsourceibias.n318 gnd 0.070526f
C1104 commonsourceibias.n319 gnd 0.011661f
C1105 commonsourceibias.n320 gnd 0.0129f
C1106 commonsourceibias.n321 gnd 0.009461f
C1107 commonsourceibias.n322 gnd 0.009461f
C1108 commonsourceibias.n323 gnd 0.012816f
C1109 commonsourceibias.n324 gnd 0.007653f
C1110 commonsourceibias.n325 gnd 0.012975f
C1111 commonsourceibias.n326 gnd 0.009461f
C1112 commonsourceibias.n327 gnd 0.009461f
C1113 commonsourceibias.n328 gnd 0.013054f
C1114 commonsourceibias.n329 gnd 0.011256f
C1115 commonsourceibias.n330 gnd 0.009134f
C1116 commonsourceibias.n331 gnd 0.009461f
C1117 commonsourceibias.n332 gnd 0.009461f
C1118 commonsourceibias.n333 gnd 0.011572f
C1119 commonsourceibias.n334 gnd 0.012989f
C1120 commonsourceibias.n335 gnd 0.070526f
C1121 commonsourceibias.n336 gnd 0.012901f
C1122 commonsourceibias.n337 gnd 0.009461f
C1123 commonsourceibias.n338 gnd 0.009461f
C1124 commonsourceibias.n339 gnd 0.009461f
C1125 commonsourceibias.n340 gnd 0.012901f
C1126 commonsourceibias.n341 gnd 0.070526f
C1127 commonsourceibias.n342 gnd 0.012989f
C1128 commonsourceibias.n343 gnd 0.011572f
C1129 commonsourceibias.n344 gnd 0.009461f
C1130 commonsourceibias.n345 gnd 0.009461f
C1131 commonsourceibias.n346 gnd 0.009461f
C1132 commonsourceibias.n347 gnd 0.011256f
C1133 commonsourceibias.n348 gnd 0.013054f
C1134 commonsourceibias.n349 gnd 0.070526f
C1135 commonsourceibias.n350 gnd 0.012975f
C1136 commonsourceibias.n351 gnd 0.009461f
C1137 commonsourceibias.n352 gnd 0.009461f
C1138 commonsourceibias.n353 gnd 0.009461f
C1139 commonsourceibias.n354 gnd 0.012816f
C1140 commonsourceibias.n355 gnd 0.070526f
C1141 commonsourceibias.n356 gnd 0.0129f
C1142 commonsourceibias.n357 gnd 0.011661f
C1143 commonsourceibias.n358 gnd 0.009461f
C1144 commonsourceibias.n359 gnd 0.009461f
C1145 commonsourceibias.n360 gnd 0.009461f
C1146 commonsourceibias.n361 gnd 0.010754f
C1147 commonsourceibias.n362 gnd 0.013093f
C1148 commonsourceibias.n363 gnd 0.070526f
C1149 commonsourceibias.n364 gnd 0.013037f
C1150 commonsourceibias.n365 gnd 0.009461f
C1151 commonsourceibias.n366 gnd 0.009461f
C1152 commonsourceibias.n367 gnd 0.009461f
C1153 commonsourceibias.n368 gnd 0.012717f
C1154 commonsourceibias.n369 gnd 0.070526f
C1155 commonsourceibias.n370 gnd 0.012748f
C1156 commonsourceibias.t147 gnd 0.191163f
C1157 commonsourceibias.n371 gnd 0.085044f
C1158 commonsourceibias.n372 gnd 0.030348f
C1159 commonsourceibias.n373 gnd 0.449685f
C1160 commonsourceibias.n374 gnd 0.012624f
C1161 commonsourceibias.t93 gnd 0.191163f
C1162 commonsourceibias.t134 gnd 0.176757f
C1163 commonsourceibias.n375 gnd 0.00769f
C1164 commonsourceibias.n376 gnd 0.009461f
C1165 commonsourceibias.t114 gnd 0.176757f
C1166 commonsourceibias.n377 gnd 0.009597f
C1167 commonsourceibias.n378 gnd 0.009461f
C1168 commonsourceibias.t123 gnd 0.176757f
C1169 commonsourceibias.n379 gnd 0.007653f
C1170 commonsourceibias.n380 gnd 0.009461f
C1171 commonsourceibias.t88 gnd 0.176757f
C1172 commonsourceibias.n381 gnd 0.009134f
C1173 commonsourceibias.n382 gnd 0.009461f
C1174 commonsourceibias.t104 gnd 0.176757f
C1175 commonsourceibias.n383 gnd 0.007641f
C1176 commonsourceibias.n384 gnd 0.009461f
C1177 commonsourceibias.t90 gnd 0.176757f
C1178 commonsourceibias.t140 gnd 0.176757f
C1179 commonsourceibias.n385 gnd 0.070526f
C1180 commonsourceibias.n386 gnd 0.009461f
C1181 commonsourceibias.t83 gnd 0.176757f
C1182 commonsourceibias.n387 gnd 0.070526f
C1183 commonsourceibias.n388 gnd 0.009461f
C1184 commonsourceibias.t151 gnd 0.176757f
C1185 commonsourceibias.n389 gnd 0.070526f
C1186 commonsourceibias.n390 gnd 0.009461f
C1187 commonsourceibias.t127 gnd 0.176757f
C1188 commonsourceibias.n391 gnd 0.010754f
C1189 commonsourceibias.n392 gnd 0.009461f
C1190 commonsourceibias.t84 gnd 0.176757f
C1191 commonsourceibias.n393 gnd 0.012717f
C1192 commonsourceibias.t112 gnd 0.196904f
C1193 commonsourceibias.t131 gnd 0.176757f
C1194 commonsourceibias.n394 gnd 0.078584f
C1195 commonsourceibias.n395 gnd 0.084191f
C1196 commonsourceibias.n396 gnd 0.04027f
C1197 commonsourceibias.n397 gnd 0.009461f
C1198 commonsourceibias.n398 gnd 0.00769f
C1199 commonsourceibias.n399 gnd 0.013037f
C1200 commonsourceibias.n400 gnd 0.070526f
C1201 commonsourceibias.n401 gnd 0.013093f
C1202 commonsourceibias.n402 gnd 0.009461f
C1203 commonsourceibias.n403 gnd 0.009461f
C1204 commonsourceibias.n404 gnd 0.009461f
C1205 commonsourceibias.n405 gnd 0.009597f
C1206 commonsourceibias.n406 gnd 0.070526f
C1207 commonsourceibias.n407 gnd 0.011661f
C1208 commonsourceibias.n408 gnd 0.0129f
C1209 commonsourceibias.n409 gnd 0.009461f
C1210 commonsourceibias.n410 gnd 0.009461f
C1211 commonsourceibias.n411 gnd 0.012816f
C1212 commonsourceibias.n412 gnd 0.007653f
C1213 commonsourceibias.n413 gnd 0.012975f
C1214 commonsourceibias.n414 gnd 0.009461f
C1215 commonsourceibias.n415 gnd 0.009461f
C1216 commonsourceibias.n416 gnd 0.013054f
C1217 commonsourceibias.n417 gnd 0.011256f
C1218 commonsourceibias.n418 gnd 0.009134f
C1219 commonsourceibias.n419 gnd 0.009461f
C1220 commonsourceibias.n420 gnd 0.009461f
C1221 commonsourceibias.n421 gnd 0.011572f
C1222 commonsourceibias.n422 gnd 0.012989f
C1223 commonsourceibias.n423 gnd 0.070526f
C1224 commonsourceibias.n424 gnd 0.012901f
C1225 commonsourceibias.n425 gnd 0.009415f
C1226 commonsourceibias.t15 gnd 0.020415f
C1227 commonsourceibias.t1 gnd 0.020415f
C1228 commonsourceibias.n426 gnd 0.181002f
C1229 commonsourceibias.t39 gnd 0.020415f
C1230 commonsourceibias.t19 gnd 0.020415f
C1231 commonsourceibias.n427 gnd 0.180398f
C1232 commonsourceibias.n428 gnd 0.168097f
C1233 commonsourceibias.t63 gnd 0.020415f
C1234 commonsourceibias.t41 gnd 0.020415f
C1235 commonsourceibias.n429 gnd 0.180398f
C1236 commonsourceibias.n430 gnd 0.082864f
C1237 commonsourceibias.t61 gnd 0.020415f
C1238 commonsourceibias.t35 gnd 0.020415f
C1239 commonsourceibias.n431 gnd 0.180398f
C1240 commonsourceibias.n432 gnd 0.069229f
C1241 commonsourceibias.n433 gnd 0.012624f
C1242 commonsourceibias.t44 gnd 0.176757f
C1243 commonsourceibias.n434 gnd 0.00769f
C1244 commonsourceibias.n435 gnd 0.009461f
C1245 commonsourceibias.t12 gnd 0.176757f
C1246 commonsourceibias.n436 gnd 0.009597f
C1247 commonsourceibias.n437 gnd 0.009461f
C1248 commonsourceibias.t26 gnd 0.176757f
C1249 commonsourceibias.n438 gnd 0.007653f
C1250 commonsourceibias.n439 gnd 0.009461f
C1251 commonsourceibias.t36 gnd 0.176757f
C1252 commonsourceibias.n440 gnd 0.009134f
C1253 commonsourceibias.n441 gnd 0.009461f
C1254 commonsourceibias.t4 gnd 0.176757f
C1255 commonsourceibias.n442 gnd 0.007641f
C1256 commonsourceibias.n443 gnd 0.009461f
C1257 commonsourceibias.t34 gnd 0.176757f
C1258 commonsourceibias.t60 gnd 0.176757f
C1259 commonsourceibias.n444 gnd 0.070526f
C1260 commonsourceibias.n445 gnd 0.009461f
C1261 commonsourceibias.t40 gnd 0.176757f
C1262 commonsourceibias.n446 gnd 0.070526f
C1263 commonsourceibias.n447 gnd 0.009461f
C1264 commonsourceibias.t62 gnd 0.176757f
C1265 commonsourceibias.n448 gnd 0.070526f
C1266 commonsourceibias.n449 gnd 0.009461f
C1267 commonsourceibias.t18 gnd 0.176757f
C1268 commonsourceibias.n450 gnd 0.010754f
C1269 commonsourceibias.n451 gnd 0.009461f
C1270 commonsourceibias.t38 gnd 0.176757f
C1271 commonsourceibias.n452 gnd 0.012717f
C1272 commonsourceibias.t14 gnd 0.196904f
C1273 commonsourceibias.t0 gnd 0.176757f
C1274 commonsourceibias.n453 gnd 0.078584f
C1275 commonsourceibias.n454 gnd 0.084191f
C1276 commonsourceibias.n455 gnd 0.04027f
C1277 commonsourceibias.n456 gnd 0.009461f
C1278 commonsourceibias.n457 gnd 0.00769f
C1279 commonsourceibias.n458 gnd 0.013037f
C1280 commonsourceibias.n459 gnd 0.070526f
C1281 commonsourceibias.n460 gnd 0.013093f
C1282 commonsourceibias.n461 gnd 0.009461f
C1283 commonsourceibias.n462 gnd 0.009461f
C1284 commonsourceibias.n463 gnd 0.009461f
C1285 commonsourceibias.n464 gnd 0.009597f
C1286 commonsourceibias.n465 gnd 0.070526f
C1287 commonsourceibias.n466 gnd 0.011661f
C1288 commonsourceibias.n467 gnd 0.0129f
C1289 commonsourceibias.n468 gnd 0.009461f
C1290 commonsourceibias.n469 gnd 0.009461f
C1291 commonsourceibias.n470 gnd 0.012816f
C1292 commonsourceibias.n471 gnd 0.007653f
C1293 commonsourceibias.n472 gnd 0.012975f
C1294 commonsourceibias.n473 gnd 0.009461f
C1295 commonsourceibias.n474 gnd 0.009461f
C1296 commonsourceibias.n475 gnd 0.013054f
C1297 commonsourceibias.n476 gnd 0.011256f
C1298 commonsourceibias.n477 gnd 0.009134f
C1299 commonsourceibias.n478 gnd 0.009461f
C1300 commonsourceibias.n479 gnd 0.009461f
C1301 commonsourceibias.n480 gnd 0.011572f
C1302 commonsourceibias.n481 gnd 0.012989f
C1303 commonsourceibias.n482 gnd 0.070526f
C1304 commonsourceibias.n483 gnd 0.012901f
C1305 commonsourceibias.n484 gnd 0.009461f
C1306 commonsourceibias.n485 gnd 0.009461f
C1307 commonsourceibias.n486 gnd 0.009461f
C1308 commonsourceibias.n487 gnd 0.012901f
C1309 commonsourceibias.n488 gnd 0.070526f
C1310 commonsourceibias.n489 gnd 0.012989f
C1311 commonsourceibias.t46 gnd 0.176757f
C1312 commonsourceibias.n490 gnd 0.070526f
C1313 commonsourceibias.n491 gnd 0.011572f
C1314 commonsourceibias.n492 gnd 0.009461f
C1315 commonsourceibias.n493 gnd 0.009461f
C1316 commonsourceibias.n494 gnd 0.009461f
C1317 commonsourceibias.n495 gnd 0.011256f
C1318 commonsourceibias.n496 gnd 0.013054f
C1319 commonsourceibias.n497 gnd 0.070526f
C1320 commonsourceibias.n498 gnd 0.012975f
C1321 commonsourceibias.n499 gnd 0.009461f
C1322 commonsourceibias.n500 gnd 0.009461f
C1323 commonsourceibias.n501 gnd 0.009461f
C1324 commonsourceibias.n502 gnd 0.012816f
C1325 commonsourceibias.n503 gnd 0.070526f
C1326 commonsourceibias.n504 gnd 0.0129f
C1327 commonsourceibias.t54 gnd 0.176757f
C1328 commonsourceibias.n505 gnd 0.070526f
C1329 commonsourceibias.n506 gnd 0.011661f
C1330 commonsourceibias.n507 gnd 0.009461f
C1331 commonsourceibias.n508 gnd 0.009461f
C1332 commonsourceibias.n509 gnd 0.009461f
C1333 commonsourceibias.n510 gnd 0.010754f
C1334 commonsourceibias.n511 gnd 0.013093f
C1335 commonsourceibias.n512 gnd 0.070526f
C1336 commonsourceibias.n513 gnd 0.013037f
C1337 commonsourceibias.n514 gnd 0.009461f
C1338 commonsourceibias.n515 gnd 0.009461f
C1339 commonsourceibias.n516 gnd 0.009461f
C1340 commonsourceibias.n517 gnd 0.012717f
C1341 commonsourceibias.n518 gnd 0.070526f
C1342 commonsourceibias.n519 gnd 0.012748f
C1343 commonsourceibias.t58 gnd 0.191163f
C1344 commonsourceibias.n520 gnd 0.085044f
C1345 commonsourceibias.n521 gnd 0.095092f
C1346 commonsourceibias.t45 gnd 0.020415f
C1347 commonsourceibias.t59 gnd 0.020415f
C1348 commonsourceibias.n522 gnd 0.180398f
C1349 commonsourceibias.n523 gnd 0.156264f
C1350 commonsourceibias.t55 gnd 0.020415f
C1351 commonsourceibias.t13 gnd 0.020415f
C1352 commonsourceibias.n524 gnd 0.180398f
C1353 commonsourceibias.n525 gnd 0.082864f
C1354 commonsourceibias.t37 gnd 0.020415f
C1355 commonsourceibias.t27 gnd 0.020415f
C1356 commonsourceibias.n526 gnd 0.180398f
C1357 commonsourceibias.n527 gnd 0.082864f
C1358 commonsourceibias.t5 gnd 0.020415f
C1359 commonsourceibias.t47 gnd 0.020415f
C1360 commonsourceibias.n528 gnd 0.180398f
C1361 commonsourceibias.n529 gnd 0.069229f
C1362 commonsourceibias.n530 gnd 0.083829f
C1363 commonsourceibias.n531 gnd 0.06839f
C1364 commonsourceibias.n532 gnd 0.009415f
C1365 commonsourceibias.n533 gnd 0.012901f
C1366 commonsourceibias.n534 gnd 0.070526f
C1367 commonsourceibias.n535 gnd 0.012989f
C1368 commonsourceibias.t74 gnd 0.176757f
C1369 commonsourceibias.n536 gnd 0.070526f
C1370 commonsourceibias.n537 gnd 0.011572f
C1371 commonsourceibias.n538 gnd 0.009461f
C1372 commonsourceibias.n539 gnd 0.009461f
C1373 commonsourceibias.n540 gnd 0.009461f
C1374 commonsourceibias.n541 gnd 0.011256f
C1375 commonsourceibias.n542 gnd 0.013054f
C1376 commonsourceibias.n543 gnd 0.070526f
C1377 commonsourceibias.n544 gnd 0.012975f
C1378 commonsourceibias.n545 gnd 0.009461f
C1379 commonsourceibias.n546 gnd 0.009461f
C1380 commonsourceibias.n547 gnd 0.009461f
C1381 commonsourceibias.n548 gnd 0.012816f
C1382 commonsourceibias.n549 gnd 0.070526f
C1383 commonsourceibias.n550 gnd 0.0129f
C1384 commonsourceibias.t95 gnd 0.176757f
C1385 commonsourceibias.n551 gnd 0.070526f
C1386 commonsourceibias.n552 gnd 0.011661f
C1387 commonsourceibias.n553 gnd 0.009461f
C1388 commonsourceibias.n554 gnd 0.009461f
C1389 commonsourceibias.n555 gnd 0.009461f
C1390 commonsourceibias.n556 gnd 0.010754f
C1391 commonsourceibias.n557 gnd 0.013093f
C1392 commonsourceibias.n558 gnd 0.070526f
C1393 commonsourceibias.n559 gnd 0.013037f
C1394 commonsourceibias.n560 gnd 0.009461f
C1395 commonsourceibias.n561 gnd 0.009461f
C1396 commonsourceibias.n562 gnd 0.009461f
C1397 commonsourceibias.n563 gnd 0.012717f
C1398 commonsourceibias.n564 gnd 0.070526f
C1399 commonsourceibias.n565 gnd 0.012748f
C1400 commonsourceibias.n566 gnd 0.085044f
C1401 commonsourceibias.n567 gnd 0.056182f
C1402 commonsourceibias.n568 gnd 0.012624f
C1403 commonsourceibias.t142 gnd 0.176757f
C1404 commonsourceibias.n569 gnd 0.00769f
C1405 commonsourceibias.n570 gnd 0.009461f
C1406 commonsourceibias.t66 gnd 0.176757f
C1407 commonsourceibias.n571 gnd 0.009597f
C1408 commonsourceibias.n572 gnd 0.009461f
C1409 commonsourceibias.t143 gnd 0.176757f
C1410 commonsourceibias.n573 gnd 0.007653f
C1411 commonsourceibias.n574 gnd 0.009461f
C1412 commonsourceibias.t67 gnd 0.176757f
C1413 commonsourceibias.n575 gnd 0.009134f
C1414 commonsourceibias.n576 gnd 0.009461f
C1415 commonsourceibias.t144 gnd 0.176757f
C1416 commonsourceibias.n577 gnd 0.007641f
C1417 commonsourceibias.n578 gnd 0.009461f
C1418 commonsourceibias.t70 gnd 0.176757f
C1419 commonsourceibias.t101 gnd 0.176757f
C1420 commonsourceibias.n579 gnd 0.070526f
C1421 commonsourceibias.n580 gnd 0.009461f
C1422 commonsourceibias.t80 gnd 0.176757f
C1423 commonsourceibias.n581 gnd 0.070526f
C1424 commonsourceibias.n582 gnd 0.009461f
C1425 commonsourceibias.t72 gnd 0.176757f
C1426 commonsourceibias.n583 gnd 0.070526f
C1427 commonsourceibias.n584 gnd 0.009461f
C1428 commonsourceibias.t100 gnd 0.176757f
C1429 commonsourceibias.n585 gnd 0.010754f
C1430 commonsourceibias.n586 gnd 0.009461f
C1431 commonsourceibias.t87 gnd 0.176757f
C1432 commonsourceibias.n587 gnd 0.012717f
C1433 commonsourceibias.t99 gnd 0.196904f
C1434 commonsourceibias.t71 gnd 0.176757f
C1435 commonsourceibias.n588 gnd 0.078584f
C1436 commonsourceibias.n589 gnd 0.084191f
C1437 commonsourceibias.n590 gnd 0.04027f
C1438 commonsourceibias.n591 gnd 0.009461f
C1439 commonsourceibias.n592 gnd 0.00769f
C1440 commonsourceibias.n593 gnd 0.013037f
C1441 commonsourceibias.n594 gnd 0.070526f
C1442 commonsourceibias.n595 gnd 0.013093f
C1443 commonsourceibias.n596 gnd 0.009461f
C1444 commonsourceibias.n597 gnd 0.009461f
C1445 commonsourceibias.n598 gnd 0.009461f
C1446 commonsourceibias.n599 gnd 0.009597f
C1447 commonsourceibias.n600 gnd 0.070526f
C1448 commonsourceibias.n601 gnd 0.011661f
C1449 commonsourceibias.n602 gnd 0.0129f
C1450 commonsourceibias.n603 gnd 0.009461f
C1451 commonsourceibias.n604 gnd 0.009461f
C1452 commonsourceibias.n605 gnd 0.012816f
C1453 commonsourceibias.n606 gnd 0.007653f
C1454 commonsourceibias.n607 gnd 0.012975f
C1455 commonsourceibias.n608 gnd 0.009461f
C1456 commonsourceibias.n609 gnd 0.009461f
C1457 commonsourceibias.n610 gnd 0.013054f
C1458 commonsourceibias.n611 gnd 0.011256f
C1459 commonsourceibias.n612 gnd 0.009134f
C1460 commonsourceibias.n613 gnd 0.009461f
C1461 commonsourceibias.n614 gnd 0.009461f
C1462 commonsourceibias.n615 gnd 0.011572f
C1463 commonsourceibias.n616 gnd 0.012989f
C1464 commonsourceibias.n617 gnd 0.070526f
C1465 commonsourceibias.n618 gnd 0.012901f
C1466 commonsourceibias.n619 gnd 0.009461f
C1467 commonsourceibias.n620 gnd 0.009461f
C1468 commonsourceibias.n621 gnd 0.009461f
C1469 commonsourceibias.n622 gnd 0.012901f
C1470 commonsourceibias.n623 gnd 0.070526f
C1471 commonsourceibias.n624 gnd 0.012989f
C1472 commonsourceibias.t98 gnd 0.176757f
C1473 commonsourceibias.n625 gnd 0.070526f
C1474 commonsourceibias.n626 gnd 0.011572f
C1475 commonsourceibias.n627 gnd 0.009461f
C1476 commonsourceibias.n628 gnd 0.009461f
C1477 commonsourceibias.n629 gnd 0.009461f
C1478 commonsourceibias.n630 gnd 0.011256f
C1479 commonsourceibias.n631 gnd 0.013054f
C1480 commonsourceibias.n632 gnd 0.070526f
C1481 commonsourceibias.n633 gnd 0.012975f
C1482 commonsourceibias.n634 gnd 0.009461f
C1483 commonsourceibias.n635 gnd 0.009461f
C1484 commonsourceibias.n636 gnd 0.009461f
C1485 commonsourceibias.n637 gnd 0.012816f
C1486 commonsourceibias.n638 gnd 0.070526f
C1487 commonsourceibias.n639 gnd 0.0129f
C1488 commonsourceibias.t154 gnd 0.176757f
C1489 commonsourceibias.n640 gnd 0.070526f
C1490 commonsourceibias.n641 gnd 0.011661f
C1491 commonsourceibias.n642 gnd 0.009461f
C1492 commonsourceibias.n643 gnd 0.009461f
C1493 commonsourceibias.n644 gnd 0.009461f
C1494 commonsourceibias.n645 gnd 0.010754f
C1495 commonsourceibias.n646 gnd 0.013093f
C1496 commonsourceibias.n647 gnd 0.070526f
C1497 commonsourceibias.n648 gnd 0.013037f
C1498 commonsourceibias.n649 gnd 0.009461f
C1499 commonsourceibias.n650 gnd 0.009461f
C1500 commonsourceibias.n651 gnd 0.009461f
C1501 commonsourceibias.n652 gnd 0.012717f
C1502 commonsourceibias.n653 gnd 0.070526f
C1503 commonsourceibias.n654 gnd 0.012748f
C1504 commonsourceibias.t150 gnd 0.191163f
C1505 commonsourceibias.n655 gnd 0.085044f
C1506 commonsourceibias.n656 gnd 0.030348f
C1507 commonsourceibias.n657 gnd 0.15151f
C1508 commonsourceibias.n658 gnd 0.012624f
C1509 commonsourceibias.t107 gnd 0.176757f
C1510 commonsourceibias.n659 gnd 0.00769f
C1511 commonsourceibias.n660 gnd 0.009461f
C1512 commonsourceibias.t122 gnd 0.176757f
C1513 commonsourceibias.n661 gnd 0.009597f
C1514 commonsourceibias.n662 gnd 0.009461f
C1515 commonsourceibias.t97 gnd 0.176757f
C1516 commonsourceibias.n663 gnd 0.007653f
C1517 commonsourceibias.n664 gnd 0.009461f
C1518 commonsourceibias.t115 gnd 0.176757f
C1519 commonsourceibias.n665 gnd 0.009134f
C1520 commonsourceibias.n666 gnd 0.009461f
C1521 commonsourceibias.t81 gnd 0.176757f
C1522 commonsourceibias.n667 gnd 0.007641f
C1523 commonsourceibias.n668 gnd 0.009461f
C1524 commonsourceibias.t69 gnd 0.176757f
C1525 commonsourceibias.t103 gnd 0.176757f
C1526 commonsourceibias.n669 gnd 0.070526f
C1527 commonsourceibias.n670 gnd 0.009461f
C1528 commonsourceibias.t132 gnd 0.176757f
C1529 commonsourceibias.n671 gnd 0.070526f
C1530 commonsourceibias.n672 gnd 0.009461f
C1531 commonsourceibias.t153 gnd 0.176757f
C1532 commonsourceibias.n673 gnd 0.070526f
C1533 commonsourceibias.n674 gnd 0.009461f
C1534 commonsourceibias.t86 gnd 0.176757f
C1535 commonsourceibias.n675 gnd 0.010754f
C1536 commonsourceibias.n676 gnd 0.009461f
C1537 commonsourceibias.t111 gnd 0.176757f
C1538 commonsourceibias.n677 gnd 0.012717f
C1539 commonsourceibias.t73 gnd 0.196904f
C1540 commonsourceibias.t145 gnd 0.176757f
C1541 commonsourceibias.n678 gnd 0.078584f
C1542 commonsourceibias.n679 gnd 0.084191f
C1543 commonsourceibias.n680 gnd 0.04027f
C1544 commonsourceibias.n681 gnd 0.009461f
C1545 commonsourceibias.n682 gnd 0.00769f
C1546 commonsourceibias.n683 gnd 0.013037f
C1547 commonsourceibias.n684 gnd 0.070526f
C1548 commonsourceibias.n685 gnd 0.013093f
C1549 commonsourceibias.n686 gnd 0.009461f
C1550 commonsourceibias.n687 gnd 0.009461f
C1551 commonsourceibias.n688 gnd 0.009461f
C1552 commonsourceibias.n689 gnd 0.009597f
C1553 commonsourceibias.n690 gnd 0.070526f
C1554 commonsourceibias.n691 gnd 0.011661f
C1555 commonsourceibias.n692 gnd 0.0129f
C1556 commonsourceibias.n693 gnd 0.009461f
C1557 commonsourceibias.n694 gnd 0.009461f
C1558 commonsourceibias.n695 gnd 0.012816f
C1559 commonsourceibias.n696 gnd 0.007653f
C1560 commonsourceibias.n697 gnd 0.012975f
C1561 commonsourceibias.n698 gnd 0.009461f
C1562 commonsourceibias.n699 gnd 0.009461f
C1563 commonsourceibias.n700 gnd 0.013054f
C1564 commonsourceibias.n701 gnd 0.011256f
C1565 commonsourceibias.n702 gnd 0.009134f
C1566 commonsourceibias.n703 gnd 0.009461f
C1567 commonsourceibias.n704 gnd 0.009461f
C1568 commonsourceibias.n705 gnd 0.011572f
C1569 commonsourceibias.n706 gnd 0.012989f
C1570 commonsourceibias.n707 gnd 0.070526f
C1571 commonsourceibias.n708 gnd 0.012901f
C1572 commonsourceibias.n709 gnd 0.009461f
C1573 commonsourceibias.n710 gnd 0.009461f
C1574 commonsourceibias.n711 gnd 0.009461f
C1575 commonsourceibias.n712 gnd 0.012901f
C1576 commonsourceibias.n713 gnd 0.070526f
C1577 commonsourceibias.n714 gnd 0.012989f
C1578 commonsourceibias.t110 gnd 0.176757f
C1579 commonsourceibias.n715 gnd 0.070526f
C1580 commonsourceibias.n716 gnd 0.011572f
C1581 commonsourceibias.n717 gnd 0.009461f
C1582 commonsourceibias.n718 gnd 0.009461f
C1583 commonsourceibias.n719 gnd 0.009461f
C1584 commonsourceibias.n720 gnd 0.011256f
C1585 commonsourceibias.n721 gnd 0.013054f
C1586 commonsourceibias.n722 gnd 0.070526f
C1587 commonsourceibias.n723 gnd 0.012975f
C1588 commonsourceibias.n724 gnd 0.009461f
C1589 commonsourceibias.n725 gnd 0.009461f
C1590 commonsourceibias.n726 gnd 0.009461f
C1591 commonsourceibias.n727 gnd 0.012816f
C1592 commonsourceibias.n728 gnd 0.070526f
C1593 commonsourceibias.n729 gnd 0.0129f
C1594 commonsourceibias.t136 gnd 0.176757f
C1595 commonsourceibias.n730 gnd 0.070526f
C1596 commonsourceibias.n731 gnd 0.011661f
C1597 commonsourceibias.n732 gnd 0.009461f
C1598 commonsourceibias.n733 gnd 0.009461f
C1599 commonsourceibias.n734 gnd 0.009461f
C1600 commonsourceibias.n735 gnd 0.010754f
C1601 commonsourceibias.n736 gnd 0.013093f
C1602 commonsourceibias.n737 gnd 0.070526f
C1603 commonsourceibias.n738 gnd 0.013037f
C1604 commonsourceibias.n739 gnd 0.009461f
C1605 commonsourceibias.n740 gnd 0.009461f
C1606 commonsourceibias.n741 gnd 0.009461f
C1607 commonsourceibias.n742 gnd 0.012717f
C1608 commonsourceibias.n743 gnd 0.070526f
C1609 commonsourceibias.n744 gnd 0.012748f
C1610 commonsourceibias.t82 gnd 0.191163f
C1611 commonsourceibias.n745 gnd 0.085044f
C1612 commonsourceibias.n746 gnd 0.030348f
C1613 commonsourceibias.n747 gnd 0.199656f
C1614 commonsourceibias.n748 gnd 5.01419f
C1615 CSoutput.n0 gnd 0.037845f
C1616 CSoutput.t150 gnd 0.250336f
C1617 CSoutput.n1 gnd 0.113039f
C1618 CSoutput.n2 gnd 0.037845f
C1619 CSoutput.t157 gnd 0.250336f
C1620 CSoutput.n3 gnd 0.029995f
C1621 CSoutput.n4 gnd 0.037845f
C1622 CSoutput.t164 gnd 0.250336f
C1623 CSoutput.n5 gnd 0.025865f
C1624 CSoutput.n6 gnd 0.037845f
C1625 CSoutput.t155 gnd 0.250336f
C1626 CSoutput.t152 gnd 0.250336f
C1627 CSoutput.n7 gnd 0.111807f
C1628 CSoutput.n8 gnd 0.037845f
C1629 CSoutput.t163 gnd 0.250336f
C1630 CSoutput.n9 gnd 0.024661f
C1631 CSoutput.n10 gnd 0.037845f
C1632 CSoutput.t145 gnd 0.250336f
C1633 CSoutput.t149 gnd 0.250336f
C1634 CSoutput.n11 gnd 0.111807f
C1635 CSoutput.n12 gnd 0.037845f
C1636 CSoutput.t160 gnd 0.250336f
C1637 CSoutput.n13 gnd 0.025865f
C1638 CSoutput.n14 gnd 0.037845f
C1639 CSoutput.t159 gnd 0.250336f
C1640 CSoutput.t147 gnd 0.250336f
C1641 CSoutput.n15 gnd 0.111807f
C1642 CSoutput.n16 gnd 0.037845f
C1643 CSoutput.t153 gnd 0.250336f
C1644 CSoutput.n17 gnd 0.027625f
C1645 CSoutput.t161 gnd 0.299159f
C1646 CSoutput.t158 gnd 0.250336f
C1647 CSoutput.n18 gnd 0.142735f
C1648 CSoutput.n19 gnd 0.138502f
C1649 CSoutput.n20 gnd 0.160679f
C1650 CSoutput.n21 gnd 0.037845f
C1651 CSoutput.n22 gnd 0.031586f
C1652 CSoutput.n23 gnd 0.111807f
C1653 CSoutput.n24 gnd 0.030448f
C1654 CSoutput.n25 gnd 0.029995f
C1655 CSoutput.n26 gnd 0.037845f
C1656 CSoutput.n27 gnd 0.037845f
C1657 CSoutput.n28 gnd 0.031343f
C1658 CSoutput.n29 gnd 0.026611f
C1659 CSoutput.n30 gnd 0.114296f
C1660 CSoutput.n31 gnd 0.026978f
C1661 CSoutput.n32 gnd 0.037845f
C1662 CSoutput.n33 gnd 0.037845f
C1663 CSoutput.n34 gnd 0.037845f
C1664 CSoutput.n35 gnd 0.031009f
C1665 CSoutput.n36 gnd 0.111807f
C1666 CSoutput.n37 gnd 0.029656f
C1667 CSoutput.n38 gnd 0.030787f
C1668 CSoutput.n39 gnd 0.037845f
C1669 CSoutput.n40 gnd 0.037845f
C1670 CSoutput.n41 gnd 0.031579f
C1671 CSoutput.n42 gnd 0.028864f
C1672 CSoutput.n43 gnd 0.111807f
C1673 CSoutput.n44 gnd 0.029595f
C1674 CSoutput.n45 gnd 0.037845f
C1675 CSoutput.n46 gnd 0.037845f
C1676 CSoutput.n47 gnd 0.037845f
C1677 CSoutput.n48 gnd 0.029595f
C1678 CSoutput.n49 gnd 0.111807f
C1679 CSoutput.n50 gnd 0.028864f
C1680 CSoutput.n51 gnd 0.031579f
C1681 CSoutput.n52 gnd 0.037845f
C1682 CSoutput.n53 gnd 0.037845f
C1683 CSoutput.n54 gnd 0.030787f
C1684 CSoutput.n55 gnd 0.029656f
C1685 CSoutput.n56 gnd 0.111807f
C1686 CSoutput.n57 gnd 0.031009f
C1687 CSoutput.n58 gnd 0.037845f
C1688 CSoutput.n59 gnd 0.037845f
C1689 CSoutput.n60 gnd 0.037845f
C1690 CSoutput.n61 gnd 0.026978f
C1691 CSoutput.n62 gnd 0.114296f
C1692 CSoutput.n63 gnd 0.026611f
C1693 CSoutput.t156 gnd 0.250336f
C1694 CSoutput.n64 gnd 0.111807f
C1695 CSoutput.n65 gnd 0.031343f
C1696 CSoutput.n66 gnd 0.037845f
C1697 CSoutput.n67 gnd 0.037845f
C1698 CSoutput.n68 gnd 0.037845f
C1699 CSoutput.n69 gnd 0.030448f
C1700 CSoutput.n70 gnd 0.111807f
C1701 CSoutput.n71 gnd 0.031586f
C1702 CSoutput.n72 gnd 0.027625f
C1703 CSoutput.n73 gnd 0.037845f
C1704 CSoutput.n74 gnd 0.037845f
C1705 CSoutput.n75 gnd 0.028649f
C1706 CSoutput.n76 gnd 0.017015f
C1707 CSoutput.t162 gnd 0.281271f
C1708 CSoutput.n77 gnd 0.139724f
C1709 CSoutput.n78 gnd 0.571604f
C1710 CSoutput.t72 gnd 0.047206f
C1711 CSoutput.t34 gnd 0.047206f
C1712 CSoutput.n79 gnd 0.365487f
C1713 CSoutput.t62 gnd 0.047206f
C1714 CSoutput.t51 gnd 0.047206f
C1715 CSoutput.n80 gnd 0.364835f
C1716 CSoutput.n81 gnd 0.370307f
C1717 CSoutput.t67 gnd 0.047206f
C1718 CSoutput.t43 gnd 0.047206f
C1719 CSoutput.n82 gnd 0.364835f
C1720 CSoutput.n83 gnd 0.182472f
C1721 CSoutput.t77 gnd 0.047206f
C1722 CSoutput.t46 gnd 0.047206f
C1723 CSoutput.n84 gnd 0.364835f
C1724 CSoutput.n85 gnd 0.334611f
C1725 CSoutput.t69 gnd 0.047206f
C1726 CSoutput.t70 gnd 0.047206f
C1727 CSoutput.n86 gnd 0.365487f
C1728 CSoutput.t59 gnd 0.047206f
C1729 CSoutput.t37 gnd 0.047206f
C1730 CSoutput.n87 gnd 0.364835f
C1731 CSoutput.n88 gnd 0.370307f
C1732 CSoutput.t35 gnd 0.047206f
C1733 CSoutput.t65 gnd 0.047206f
C1734 CSoutput.n89 gnd 0.364835f
C1735 CSoutput.n90 gnd 0.182472f
C1736 CSoutput.t58 gnd 0.047206f
C1737 CSoutput.t47 gnd 0.047206f
C1738 CSoutput.n91 gnd 0.364835f
C1739 CSoutput.n92 gnd 0.272111f
C1740 CSoutput.n93 gnd 0.343131f
C1741 CSoutput.t76 gnd 0.047206f
C1742 CSoutput.t75 gnd 0.047206f
C1743 CSoutput.n94 gnd 0.365487f
C1744 CSoutput.t64 gnd 0.047206f
C1745 CSoutput.t41 gnd 0.047206f
C1746 CSoutput.n95 gnd 0.364835f
C1747 CSoutput.n96 gnd 0.370307f
C1748 CSoutput.t39 gnd 0.047206f
C1749 CSoutput.t74 gnd 0.047206f
C1750 CSoutput.n97 gnd 0.364835f
C1751 CSoutput.n98 gnd 0.182472f
C1752 CSoutput.t63 gnd 0.047206f
C1753 CSoutput.t54 gnd 0.047206f
C1754 CSoutput.n99 gnd 0.364835f
C1755 CSoutput.n100 gnd 0.272111f
C1756 CSoutput.n101 gnd 0.383532f
C1757 CSoutput.n102 gnd 6.9206f
C1758 CSoutput.n104 gnd 0.669471f
C1759 CSoutput.n105 gnd 0.502103f
C1760 CSoutput.n106 gnd 0.669471f
C1761 CSoutput.n107 gnd 0.669471f
C1762 CSoutput.n108 gnd 1.80242f
C1763 CSoutput.n109 gnd 0.669471f
C1764 CSoutput.n110 gnd 0.669471f
C1765 CSoutput.t151 gnd 0.836839f
C1766 CSoutput.n111 gnd 0.669471f
C1767 CSoutput.n112 gnd 0.669471f
C1768 CSoutput.n116 gnd 0.669471f
C1769 CSoutput.n120 gnd 0.669471f
C1770 CSoutput.n121 gnd 0.669471f
C1771 CSoutput.n123 gnd 0.669471f
C1772 CSoutput.n128 gnd 0.669471f
C1773 CSoutput.n130 gnd 0.669471f
C1774 CSoutput.n131 gnd 0.669471f
C1775 CSoutput.n133 gnd 0.669471f
C1776 CSoutput.n134 gnd 0.669471f
C1777 CSoutput.n136 gnd 0.669471f
C1778 CSoutput.t146 gnd 11.1868f
C1779 CSoutput.n138 gnd 0.669471f
C1780 CSoutput.n139 gnd 0.502103f
C1781 CSoutput.n140 gnd 0.669471f
C1782 CSoutput.n141 gnd 0.669471f
C1783 CSoutput.n142 gnd 1.80242f
C1784 CSoutput.n143 gnd 0.669471f
C1785 CSoutput.n144 gnd 0.669471f
C1786 CSoutput.t165 gnd 0.836839f
C1787 CSoutput.n145 gnd 0.669471f
C1788 CSoutput.n146 gnd 0.669471f
C1789 CSoutput.n150 gnd 0.669471f
C1790 CSoutput.n154 gnd 0.669471f
C1791 CSoutput.n155 gnd 0.669471f
C1792 CSoutput.n157 gnd 0.669471f
C1793 CSoutput.n162 gnd 0.669471f
C1794 CSoutput.n164 gnd 0.669471f
C1795 CSoutput.n165 gnd 0.669471f
C1796 CSoutput.n167 gnd 0.669471f
C1797 CSoutput.n168 gnd 0.669471f
C1798 CSoutput.n170 gnd 0.669471f
C1799 CSoutput.n171 gnd 0.502103f
C1800 CSoutput.n173 gnd 0.669471f
C1801 CSoutput.n174 gnd 0.502103f
C1802 CSoutput.n175 gnd 0.669471f
C1803 CSoutput.n176 gnd 0.669471f
C1804 CSoutput.n177 gnd 1.80242f
C1805 CSoutput.n178 gnd 0.669471f
C1806 CSoutput.n179 gnd 0.669471f
C1807 CSoutput.t144 gnd 0.836839f
C1808 CSoutput.n180 gnd 0.669471f
C1809 CSoutput.n181 gnd 1.80242f
C1810 CSoutput.n183 gnd 0.669471f
C1811 CSoutput.n184 gnd 0.669471f
C1812 CSoutput.n186 gnd 0.669471f
C1813 CSoutput.n187 gnd 0.669471f
C1814 CSoutput.t154 gnd 11.004499f
C1815 CSoutput.t148 gnd 11.1868f
C1816 CSoutput.n193 gnd 2.10023f
C1817 CSoutput.n194 gnd 8.555571f
C1818 CSoutput.n195 gnd 8.91357f
C1819 CSoutput.n200 gnd 2.27511f
C1820 CSoutput.n206 gnd 0.669471f
C1821 CSoutput.n208 gnd 0.669471f
C1822 CSoutput.n210 gnd 0.669471f
C1823 CSoutput.n212 gnd 0.669471f
C1824 CSoutput.n214 gnd 0.669471f
C1825 CSoutput.n220 gnd 0.669471f
C1826 CSoutput.n227 gnd 1.22822f
C1827 CSoutput.n228 gnd 1.22822f
C1828 CSoutput.n229 gnd 0.669471f
C1829 CSoutput.n230 gnd 0.669471f
C1830 CSoutput.n232 gnd 0.502103f
C1831 CSoutput.n233 gnd 0.430006f
C1832 CSoutput.n235 gnd 0.502103f
C1833 CSoutput.n236 gnd 0.430006f
C1834 CSoutput.n237 gnd 0.502103f
C1835 CSoutput.n239 gnd 0.669471f
C1836 CSoutput.n241 gnd 1.80242f
C1837 CSoutput.n242 gnd 2.10023f
C1838 CSoutput.n243 gnd 7.86892f
C1839 CSoutput.n245 gnd 0.502103f
C1840 CSoutput.n246 gnd 1.29194f
C1841 CSoutput.n247 gnd 0.502103f
C1842 CSoutput.n249 gnd 0.669471f
C1843 CSoutput.n251 gnd 1.80242f
C1844 CSoutput.n252 gnd 3.92597f
C1845 CSoutput.t33 gnd 0.047206f
C1846 CSoutput.t73 gnd 0.047206f
C1847 CSoutput.n253 gnd 0.365487f
C1848 CSoutput.t49 gnd 0.047206f
C1849 CSoutput.t79 gnd 0.047206f
C1850 CSoutput.n254 gnd 0.364835f
C1851 CSoutput.n255 gnd 0.370307f
C1852 CSoutput.t42 gnd 0.047206f
C1853 CSoutput.t68 gnd 0.047206f
C1854 CSoutput.n256 gnd 0.364835f
C1855 CSoutput.n257 gnd 0.182472f
C1856 CSoutput.t45 gnd 0.047206f
C1857 CSoutput.t78 gnd 0.047206f
C1858 CSoutput.n258 gnd 0.364835f
C1859 CSoutput.n259 gnd 0.334611f
C1860 CSoutput.t52 gnd 0.047206f
C1861 CSoutput.t53 gnd 0.047206f
C1862 CSoutput.n260 gnd 0.365487f
C1863 CSoutput.t61 gnd 0.047206f
C1864 CSoutput.t36 gnd 0.047206f
C1865 CSoutput.n261 gnd 0.364835f
C1866 CSoutput.n262 gnd 0.370307f
C1867 CSoutput.t50 gnd 0.047206f
C1868 CSoutput.t60 gnd 0.047206f
C1869 CSoutput.n263 gnd 0.364835f
C1870 CSoutput.n264 gnd 0.182472f
C1871 CSoutput.t32 gnd 0.047206f
C1872 CSoutput.t44 gnd 0.047206f
C1873 CSoutput.n265 gnd 0.364835f
C1874 CSoutput.n266 gnd 0.272111f
C1875 CSoutput.n267 gnd 0.343131f
C1876 CSoutput.t56 gnd 0.047206f
C1877 CSoutput.t57 gnd 0.047206f
C1878 CSoutput.n268 gnd 0.365487f
C1879 CSoutput.t71 gnd 0.047206f
C1880 CSoutput.t40 gnd 0.047206f
C1881 CSoutput.n269 gnd 0.364835f
C1882 CSoutput.n270 gnd 0.370307f
C1883 CSoutput.t55 gnd 0.047206f
C1884 CSoutput.t66 gnd 0.047206f
C1885 CSoutput.n271 gnd 0.364835f
C1886 CSoutput.n272 gnd 0.182472f
C1887 CSoutput.t38 gnd 0.047206f
C1888 CSoutput.t48 gnd 0.047206f
C1889 CSoutput.n273 gnd 0.364834f
C1890 CSoutput.n274 gnd 0.272113f
C1891 CSoutput.n275 gnd 0.383532f
C1892 CSoutput.n276 gnd 9.9266f
C1893 CSoutput.t142 gnd 0.041305f
C1894 CSoutput.t99 gnd 0.041305f
C1895 CSoutput.n277 gnd 0.366211f
C1896 CSoutput.t30 gnd 0.041305f
C1897 CSoutput.t130 gnd 0.041305f
C1898 CSoutput.n278 gnd 0.36499f
C1899 CSoutput.n279 gnd 0.340103f
C1900 CSoutput.t119 gnd 0.041305f
C1901 CSoutput.t141 gnd 0.041305f
C1902 CSoutput.n280 gnd 0.36499f
C1903 CSoutput.n281 gnd 0.167654f
C1904 CSoutput.t140 gnd 0.041305f
C1905 CSoutput.t88 gnd 0.041305f
C1906 CSoutput.n282 gnd 0.36499f
C1907 CSoutput.n283 gnd 0.167654f
C1908 CSoutput.t97 gnd 0.041305f
C1909 CSoutput.t28 gnd 0.041305f
C1910 CSoutput.n284 gnd 0.36499f
C1911 CSoutput.n285 gnd 0.167654f
C1912 CSoutput.t96 gnd 0.041305f
C1913 CSoutput.t22 gnd 0.041305f
C1914 CSoutput.n286 gnd 0.36499f
C1915 CSoutput.n287 gnd 0.167654f
C1916 CSoutput.t94 gnd 0.041305f
C1917 CSoutput.t128 gnd 0.041305f
C1918 CSoutput.n288 gnd 0.36499f
C1919 CSoutput.n289 gnd 0.167654f
C1920 CSoutput.t18 gnd 0.041305f
C1921 CSoutput.t90 gnd 0.041305f
C1922 CSoutput.n290 gnd 0.36499f
C1923 CSoutput.n291 gnd 0.30923f
C1924 CSoutput.t132 gnd 0.041305f
C1925 CSoutput.t15 gnd 0.041305f
C1926 CSoutput.n292 gnd 0.366211f
C1927 CSoutput.t13 gnd 0.041305f
C1928 CSoutput.t27 gnd 0.041305f
C1929 CSoutput.n293 gnd 0.36499f
C1930 CSoutput.n294 gnd 0.340103f
C1931 CSoutput.t24 gnd 0.041305f
C1932 CSoutput.t1 gnd 0.041305f
C1933 CSoutput.n295 gnd 0.36499f
C1934 CSoutput.n296 gnd 0.167654f
C1935 CSoutput.t123 gnd 0.041305f
C1936 CSoutput.t11 gnd 0.041305f
C1937 CSoutput.n297 gnd 0.36499f
C1938 CSoutput.n298 gnd 0.167654f
C1939 CSoutput.t106 gnd 0.041305f
C1940 CSoutput.t8 gnd 0.041305f
C1941 CSoutput.n299 gnd 0.36499f
C1942 CSoutput.n300 gnd 0.167654f
C1943 CSoutput.t17 gnd 0.041305f
C1944 CSoutput.t104 gnd 0.041305f
C1945 CSoutput.n301 gnd 0.36499f
C1946 CSoutput.n302 gnd 0.167654f
C1947 CSoutput.t143 gnd 0.041305f
C1948 CSoutput.t126 gnd 0.041305f
C1949 CSoutput.n303 gnd 0.36499f
C1950 CSoutput.n304 gnd 0.167654f
C1951 CSoutput.t138 gnd 0.041305f
C1952 CSoutput.t108 gnd 0.041305f
C1953 CSoutput.n305 gnd 0.36499f
C1954 CSoutput.n306 gnd 0.254535f
C1955 CSoutput.n307 gnd 0.321048f
C1956 CSoutput.t116 gnd 0.041305f
C1957 CSoutput.t81 gnd 0.041305f
C1958 CSoutput.n308 gnd 0.366211f
C1959 CSoutput.t89 gnd 0.041305f
C1960 CSoutput.t102 gnd 0.041305f
C1961 CSoutput.n309 gnd 0.36499f
C1962 CSoutput.n310 gnd 0.340103f
C1963 CSoutput.t14 gnd 0.041305f
C1964 CSoutput.t135 gnd 0.041305f
C1965 CSoutput.n311 gnd 0.36499f
C1966 CSoutput.n312 gnd 0.167654f
C1967 CSoutput.t129 gnd 0.041305f
C1968 CSoutput.t120 gnd 0.041305f
C1969 CSoutput.n313 gnd 0.36499f
C1970 CSoutput.n314 gnd 0.167654f
C1971 CSoutput.t12 gnd 0.041305f
C1972 CSoutput.t98 gnd 0.041305f
C1973 CSoutput.n315 gnd 0.36499f
C1974 CSoutput.n316 gnd 0.167654f
C1975 CSoutput.t2 gnd 0.041305f
C1976 CSoutput.t16 gnd 0.041305f
C1977 CSoutput.n317 gnd 0.36499f
C1978 CSoutput.n318 gnd 0.167654f
C1979 CSoutput.t4 gnd 0.041305f
C1980 CSoutput.t122 gnd 0.041305f
C1981 CSoutput.n319 gnd 0.36499f
C1982 CSoutput.n320 gnd 0.167654f
C1983 CSoutput.t103 gnd 0.041305f
C1984 CSoutput.t20 gnd 0.041305f
C1985 CSoutput.n321 gnd 0.36499f
C1986 CSoutput.n322 gnd 0.254535f
C1987 CSoutput.n323 gnd 0.344755f
C1988 CSoutput.n324 gnd 10.6183f
C1989 CSoutput.t121 gnd 0.041305f
C1990 CSoutput.t105 gnd 0.041305f
C1991 CSoutput.n325 gnd 0.366211f
C1992 CSoutput.t107 gnd 0.041305f
C1993 CSoutput.t115 gnd 0.041305f
C1994 CSoutput.n326 gnd 0.36499f
C1995 CSoutput.n327 gnd 0.340103f
C1996 CSoutput.t134 gnd 0.041305f
C1997 CSoutput.t29 gnd 0.041305f
C1998 CSoutput.n328 gnd 0.36499f
C1999 CSoutput.n329 gnd 0.167654f
C2000 CSoutput.t7 gnd 0.041305f
C2001 CSoutput.t80 gnd 0.041305f
C2002 CSoutput.n330 gnd 0.36499f
C2003 CSoutput.n331 gnd 0.167654f
C2004 CSoutput.t110 gnd 0.041305f
C2005 CSoutput.t137 gnd 0.041305f
C2006 CSoutput.n332 gnd 0.36499f
C2007 CSoutput.n333 gnd 0.167654f
C2008 CSoutput.t84 gnd 0.041305f
C2009 CSoutput.t92 gnd 0.041305f
C2010 CSoutput.n334 gnd 0.36499f
C2011 CSoutput.n335 gnd 0.167654f
C2012 CSoutput.t0 gnd 0.041305f
C2013 CSoutput.t131 gnd 0.041305f
C2014 CSoutput.n336 gnd 0.36499f
C2015 CSoutput.n337 gnd 0.167654f
C2016 CSoutput.t87 gnd 0.041305f
C2017 CSoutput.t10 gnd 0.041305f
C2018 CSoutput.n338 gnd 0.36499f
C2019 CSoutput.n339 gnd 0.30923f
C2020 CSoutput.t95 gnd 0.041305f
C2021 CSoutput.t83 gnd 0.041305f
C2022 CSoutput.n340 gnd 0.366211f
C2023 CSoutput.t3 gnd 0.041305f
C2024 CSoutput.t117 gnd 0.041305f
C2025 CSoutput.n341 gnd 0.36499f
C2026 CSoutput.n342 gnd 0.340103f
C2027 CSoutput.t118 gnd 0.041305f
C2028 CSoutput.t21 gnd 0.041305f
C2029 CSoutput.n343 gnd 0.36499f
C2030 CSoutput.n344 gnd 0.167654f
C2031 CSoutput.t112 gnd 0.041305f
C2032 CSoutput.t136 gnd 0.041305f
C2033 CSoutput.n345 gnd 0.36499f
C2034 CSoutput.n346 gnd 0.167654f
C2035 CSoutput.t86 gnd 0.041305f
C2036 CSoutput.t25 gnd 0.041305f
C2037 CSoutput.n347 gnd 0.36499f
C2038 CSoutput.n348 gnd 0.167654f
C2039 CSoutput.t100 gnd 0.041305f
C2040 CSoutput.t124 gnd 0.041305f
C2041 CSoutput.n349 gnd 0.36499f
C2042 CSoutput.n350 gnd 0.167654f
C2043 CSoutput.t6 gnd 0.041305f
C2044 CSoutput.t139 gnd 0.041305f
C2045 CSoutput.n351 gnd 0.36499f
C2046 CSoutput.n352 gnd 0.167654f
C2047 CSoutput.t85 gnd 0.041305f
C2048 CSoutput.t26 gnd 0.041305f
C2049 CSoutput.n353 gnd 0.36499f
C2050 CSoutput.n354 gnd 0.254535f
C2051 CSoutput.n355 gnd 0.321048f
C2052 CSoutput.t127 gnd 0.041305f
C2053 CSoutput.t91 gnd 0.041305f
C2054 CSoutput.n356 gnd 0.366211f
C2055 CSoutput.t111 gnd 0.041305f
C2056 CSoutput.t9 gnd 0.041305f
C2057 CSoutput.n357 gnd 0.36499f
C2058 CSoutput.n358 gnd 0.340103f
C2059 CSoutput.t31 gnd 0.041305f
C2060 CSoutput.t82 gnd 0.041305f
C2061 CSoutput.n359 gnd 0.36499f
C2062 CSoutput.n360 gnd 0.167654f
C2063 CSoutput.t125 gnd 0.041305f
C2064 CSoutput.t114 gnd 0.041305f
C2065 CSoutput.n361 gnd 0.36499f
C2066 CSoutput.n362 gnd 0.167654f
C2067 CSoutput.t93 gnd 0.041305f
C2068 CSoutput.t133 gnd 0.041305f
C2069 CSoutput.n363 gnd 0.36499f
C2070 CSoutput.n364 gnd 0.167654f
C2071 CSoutput.t19 gnd 0.041305f
C2072 CSoutput.t23 gnd 0.041305f
C2073 CSoutput.n365 gnd 0.36499f
C2074 CSoutput.n366 gnd 0.167654f
C2075 CSoutput.t109 gnd 0.041305f
C2076 CSoutput.t5 gnd 0.041305f
C2077 CSoutput.n367 gnd 0.36499f
C2078 CSoutput.n368 gnd 0.167654f
C2079 CSoutput.t101 gnd 0.041305f
C2080 CSoutput.t113 gnd 0.041305f
C2081 CSoutput.n369 gnd 0.36499f
C2082 CSoutput.n370 gnd 0.254535f
C2083 CSoutput.n371 gnd 0.344755f
C2084 CSoutput.n372 gnd 6.01389f
C2085 CSoutput.n373 gnd 11.6587f
C2086 a_n5644_8799.n0 gnd 2.69839f
C2087 a_n5644_8799.n1 gnd 1.63488f
C2088 a_n5644_8799.n2 gnd 3.74044f
C2089 a_n5644_8799.n3 gnd 0.204003f
C2090 a_n5644_8799.n4 gnd 0.281239f
C2091 a_n5644_8799.n5 gnd 0.213379f
C2092 a_n5644_8799.n6 gnd 0.204003f
C2093 a_n5644_8799.n7 gnd 0.281239f
C2094 a_n5644_8799.n8 gnd 0.213379f
C2095 a_n5644_8799.n9 gnd 0.204003f
C2096 a_n5644_8799.n10 gnd 0.443208f
C2097 a_n5644_8799.n11 gnd 0.213379f
C2098 a_n5644_8799.n12 gnd 0.204003f
C2099 a_n5644_8799.n13 gnd 0.315381f
C2100 a_n5644_8799.n14 gnd 0.179237f
C2101 a_n5644_8799.n15 gnd 0.204003f
C2102 a_n5644_8799.n16 gnd 0.315381f
C2103 a_n5644_8799.n17 gnd 0.179237f
C2104 a_n5644_8799.n18 gnd 0.204003f
C2105 a_n5644_8799.n19 gnd 0.315381f
C2106 a_n5644_8799.n20 gnd 0.341207f
C2107 a_n5644_8799.n21 gnd 2.78513f
C2108 a_n5644_8799.n22 gnd 3.89483f
C2109 a_n5644_8799.n23 gnd 0.2456f
C2110 a_n5644_8799.n24 gnd 0.004585f
C2111 a_n5644_8799.n25 gnd 0.009917f
C2112 a_n5644_8799.n26 gnd 0.009917f
C2113 a_n5644_8799.n27 gnd 0.004585f
C2114 a_n5644_8799.n28 gnd 0.2456f
C2115 a_n5644_8799.n29 gnd 0.004585f
C2116 a_n5644_8799.n30 gnd 0.009917f
C2117 a_n5644_8799.n31 gnd 0.009917f
C2118 a_n5644_8799.n32 gnd 0.004585f
C2119 a_n5644_8799.n33 gnd 0.2456f
C2120 a_n5644_8799.n34 gnd 0.004585f
C2121 a_n5644_8799.n35 gnd 0.009917f
C2122 a_n5644_8799.n36 gnd 0.009917f
C2123 a_n5644_8799.n37 gnd 0.004585f
C2124 a_n5644_8799.n38 gnd 0.004585f
C2125 a_n5644_8799.n39 gnd 0.009917f
C2126 a_n5644_8799.n40 gnd 0.009917f
C2127 a_n5644_8799.n41 gnd 0.004585f
C2128 a_n5644_8799.n42 gnd 0.2456f
C2129 a_n5644_8799.n43 gnd 0.004585f
C2130 a_n5644_8799.n44 gnd 0.009917f
C2131 a_n5644_8799.n45 gnd 0.009917f
C2132 a_n5644_8799.n46 gnd 0.004585f
C2133 a_n5644_8799.n47 gnd 0.2456f
C2134 a_n5644_8799.n48 gnd 0.004585f
C2135 a_n5644_8799.n49 gnd 0.009917f
C2136 a_n5644_8799.n50 gnd 0.009917f
C2137 a_n5644_8799.n51 gnd 0.004585f
C2138 a_n5644_8799.n52 gnd 0.2456f
C2139 a_n5644_8799.t22 gnd 0.141499f
C2140 a_n5644_8799.t16 gnd 0.141499f
C2141 a_n5644_8799.t25 gnd 0.141499f
C2142 a_n5644_8799.n53 gnd 1.11602f
C2143 a_n5644_8799.t19 gnd 0.141499f
C2144 a_n5644_8799.t23 gnd 0.141499f
C2145 a_n5644_8799.n54 gnd 1.11418f
C2146 a_n5644_8799.t18 gnd 0.141499f
C2147 a_n5644_8799.t17 gnd 0.141499f
C2148 a_n5644_8799.n55 gnd 1.11418f
C2149 a_n5644_8799.t27 gnd 0.110055f
C2150 a_n5644_8799.t3 gnd 0.110055f
C2151 a_n5644_8799.n56 gnd 0.975348f
C2152 a_n5644_8799.t11 gnd 0.110055f
C2153 a_n5644_8799.t5 gnd 0.110055f
C2154 a_n5644_8799.n57 gnd 0.972481f
C2155 a_n5644_8799.t12 gnd 0.110055f
C2156 a_n5644_8799.t2 gnd 0.110055f
C2157 a_n5644_8799.n58 gnd 0.975348f
C2158 a_n5644_8799.t26 gnd 0.110055f
C2159 a_n5644_8799.t7 gnd 0.110055f
C2160 a_n5644_8799.n59 gnd 0.97248f
C2161 a_n5644_8799.t9 gnd 0.110055f
C2162 a_n5644_8799.t8 gnd 0.110055f
C2163 a_n5644_8799.n60 gnd 0.975348f
C2164 a_n5644_8799.t10 gnd 0.110055f
C2165 a_n5644_8799.t13 gnd 0.110055f
C2166 a_n5644_8799.n61 gnd 0.97248f
C2167 a_n5644_8799.t6 gnd 0.110055f
C2168 a_n5644_8799.t4 gnd 0.110055f
C2169 a_n5644_8799.n62 gnd 0.972481f
C2170 a_n5644_8799.t1 gnd 0.110055f
C2171 a_n5644_8799.t0 gnd 0.110055f
C2172 a_n5644_8799.n63 gnd 0.972481f
C2173 a_n5644_8799.t66 gnd 0.58672f
C2174 a_n5644_8799.n64 gnd 0.263697f
C2175 a_n5644_8799.t33 gnd 0.58672f
C2176 a_n5644_8799.t53 gnd 0.58672f
C2177 a_n5644_8799.t44 gnd 0.597824f
C2178 a_n5644_8799.n65 gnd 0.245962f
C2179 a_n5644_8799.n66 gnd 0.266041f
C2180 a_n5644_8799.t68 gnd 0.58672f
C2181 a_n5644_8799.n67 gnd 0.263697f
C2182 a_n5644_8799.n68 gnd 0.259367f
C2183 a_n5644_8799.t43 gnd 0.58672f
C2184 a_n5644_8799.n69 gnd 0.259367f
C2185 a_n5644_8799.t31 gnd 0.58672f
C2186 a_n5644_8799.n70 gnd 0.266041f
C2187 a_n5644_8799.t32 gnd 0.597814f
C2188 a_n5644_8799.t70 gnd 0.58672f
C2189 a_n5644_8799.n71 gnd 0.263697f
C2190 a_n5644_8799.t42 gnd 0.58672f
C2191 a_n5644_8799.t60 gnd 0.58672f
C2192 a_n5644_8799.t49 gnd 0.597824f
C2193 a_n5644_8799.n72 gnd 0.245962f
C2194 a_n5644_8799.n73 gnd 0.266041f
C2195 a_n5644_8799.t72 gnd 0.58672f
C2196 a_n5644_8799.n74 gnd 0.263697f
C2197 a_n5644_8799.n75 gnd 0.259367f
C2198 a_n5644_8799.t48 gnd 0.58672f
C2199 a_n5644_8799.n76 gnd 0.259367f
C2200 a_n5644_8799.t38 gnd 0.58672f
C2201 a_n5644_8799.n77 gnd 0.266041f
C2202 a_n5644_8799.t37 gnd 0.597814f
C2203 a_n5644_8799.n78 gnd 0.882406f
C2204 a_n5644_8799.t56 gnd 0.58672f
C2205 a_n5644_8799.n79 gnd 0.263697f
C2206 a_n5644_8799.t64 gnd 0.58672f
C2207 a_n5644_8799.t61 gnd 0.58672f
C2208 a_n5644_8799.t30 gnd 0.597824f
C2209 a_n5644_8799.n80 gnd 0.245962f
C2210 a_n5644_8799.n81 gnd 0.266041f
C2211 a_n5644_8799.t40 gnd 0.58672f
C2212 a_n5644_8799.n82 gnd 0.263697f
C2213 a_n5644_8799.n83 gnd 0.259367f
C2214 a_n5644_8799.t45 gnd 0.58672f
C2215 a_n5644_8799.n84 gnd 0.259367f
C2216 a_n5644_8799.t35 gnd 0.58672f
C2217 a_n5644_8799.n85 gnd 0.266041f
C2218 a_n5644_8799.t73 gnd 0.597814f
C2219 a_n5644_8799.n86 gnd 1.42454f
C2220 a_n5644_8799.t51 gnd 0.597814f
C2221 a_n5644_8799.t50 gnd 0.58672f
C2222 a_n5644_8799.t36 gnd 0.58672f
C2223 a_n5644_8799.n87 gnd 0.263697f
C2224 a_n5644_8799.t67 gnd 0.58672f
C2225 a_n5644_8799.t52 gnd 0.58672f
C2226 a_n5644_8799.t41 gnd 0.58672f
C2227 a_n5644_8799.n88 gnd 0.263697f
C2228 a_n5644_8799.t59 gnd 0.597824f
C2229 a_n5644_8799.n89 gnd 0.245962f
C2230 a_n5644_8799.t69 gnd 0.58672f
C2231 a_n5644_8799.n90 gnd 0.266041f
C2232 a_n5644_8799.n91 gnd 0.259367f
C2233 a_n5644_8799.n92 gnd 0.259367f
C2234 a_n5644_8799.n93 gnd 0.266041f
C2235 a_n5644_8799.t55 gnd 0.597814f
C2236 a_n5644_8799.t54 gnd 0.58672f
C2237 a_n5644_8799.t46 gnd 0.58672f
C2238 a_n5644_8799.n94 gnd 0.263697f
C2239 a_n5644_8799.t71 gnd 0.58672f
C2240 a_n5644_8799.t57 gnd 0.58672f
C2241 a_n5644_8799.t47 gnd 0.58672f
C2242 a_n5644_8799.n95 gnd 0.263697f
C2243 a_n5644_8799.t63 gnd 0.597824f
C2244 a_n5644_8799.n96 gnd 0.245962f
C2245 a_n5644_8799.t75 gnd 0.58672f
C2246 a_n5644_8799.n97 gnd 0.266041f
C2247 a_n5644_8799.n98 gnd 0.259367f
C2248 a_n5644_8799.n99 gnd 0.259367f
C2249 a_n5644_8799.n100 gnd 0.266041f
C2250 a_n5644_8799.n101 gnd 0.882406f
C2251 a_n5644_8799.t74 gnd 0.597814f
C2252 a_n5644_8799.t34 gnd 0.58672f
C2253 a_n5644_8799.t58 gnd 0.58672f
C2254 a_n5644_8799.n102 gnd 0.263697f
C2255 a_n5644_8799.t28 gnd 0.58672f
C2256 a_n5644_8799.t65 gnd 0.58672f
C2257 a_n5644_8799.t39 gnd 0.58672f
C2258 a_n5644_8799.n103 gnd 0.263697f
C2259 a_n5644_8799.t29 gnd 0.597824f
C2260 a_n5644_8799.n104 gnd 0.245962f
C2261 a_n5644_8799.t62 gnd 0.58672f
C2262 a_n5644_8799.n105 gnd 0.266041f
C2263 a_n5644_8799.n106 gnd 0.259367f
C2264 a_n5644_8799.n107 gnd 0.259367f
C2265 a_n5644_8799.n108 gnd 0.266041f
C2266 a_n5644_8799.n109 gnd 1.11694f
C2267 a_n5644_8799.n110 gnd 12.019f
C2268 a_n5644_8799.n111 gnd 4.29394f
C2269 a_n5644_8799.n112 gnd 5.58701f
C2270 a_n5644_8799.t20 gnd 0.141499f
C2271 a_n5644_8799.t21 gnd 0.141499f
C2272 a_n5644_8799.n113 gnd 1.11602f
C2273 a_n5644_8799.t24 gnd 0.141499f
C2274 a_n5644_8799.t15 gnd 0.141499f
C2275 a_n5644_8799.n114 gnd 1.11418f
C2276 a_n5644_8799.n115 gnd 1.11418f
C2277 a_n5644_8799.t14 gnd 0.141499f
C2278 vdd.t179 gnd 0.032956f
C2279 vdd.t164 gnd 0.032956f
C2280 vdd.n0 gnd 0.259932f
C2281 vdd.t148 gnd 0.032956f
C2282 vdd.t175 gnd 0.032956f
C2283 vdd.n1 gnd 0.259503f
C2284 vdd.n2 gnd 0.239312f
C2285 vdd.t161 gnd 0.032956f
C2286 vdd.t183 gnd 0.032956f
C2287 vdd.n3 gnd 0.259503f
C2288 vdd.n4 gnd 0.121029f
C2289 vdd.t185 gnd 0.032956f
C2290 vdd.t166 gnd 0.032956f
C2291 vdd.n5 gnd 0.259503f
C2292 vdd.n6 gnd 0.113563f
C2293 vdd.t188 gnd 0.032956f
C2294 vdd.t159 gnd 0.032956f
C2295 vdd.n7 gnd 0.259932f
C2296 vdd.t169 gnd 0.032956f
C2297 vdd.t181 gnd 0.032956f
C2298 vdd.n8 gnd 0.259503f
C2299 vdd.n9 gnd 0.239312f
C2300 vdd.t173 gnd 0.032956f
C2301 vdd.t151 gnd 0.032956f
C2302 vdd.n10 gnd 0.259503f
C2303 vdd.n11 gnd 0.121029f
C2304 vdd.t156 gnd 0.032956f
C2305 vdd.t171 gnd 0.032956f
C2306 vdd.n12 gnd 0.259503f
C2307 vdd.n13 gnd 0.113563f
C2308 vdd.n14 gnd 0.080287f
C2309 vdd.t92 gnd 0.018309f
C2310 vdd.t98 gnd 0.018309f
C2311 vdd.n15 gnd 0.168528f
C2312 vdd.t126 gnd 0.018309f
C2313 vdd.t127 gnd 0.018309f
C2314 vdd.n16 gnd 0.168034f
C2315 vdd.n17 gnd 0.292432f
C2316 vdd.t5 gnd 0.018309f
C2317 vdd.t100 gnd 0.018309f
C2318 vdd.n18 gnd 0.168034f
C2319 vdd.n19 gnd 0.120983f
C2320 vdd.t131 gnd 0.018309f
C2321 vdd.t128 gnd 0.018309f
C2322 vdd.n20 gnd 0.168528f
C2323 vdd.t4 gnd 0.018309f
C2324 vdd.t94 gnd 0.018309f
C2325 vdd.n21 gnd 0.168034f
C2326 vdd.n22 gnd 0.292432f
C2327 vdd.t129 gnd 0.018309f
C2328 vdd.t130 gnd 0.018309f
C2329 vdd.n23 gnd 0.168034f
C2330 vdd.n24 gnd 0.120983f
C2331 vdd.t95 gnd 0.018309f
C2332 vdd.t125 gnd 0.018309f
C2333 vdd.n25 gnd 0.168034f
C2334 vdd.t99 gnd 0.018309f
C2335 vdd.t93 gnd 0.018309f
C2336 vdd.n26 gnd 0.168034f
C2337 vdd.n27 gnd 18.423f
C2338 vdd.n28 gnd 6.88036f
C2339 vdd.n29 gnd 0.004994f
C2340 vdd.n30 gnd 0.004634f
C2341 vdd.n31 gnd 0.002563f
C2342 vdd.n32 gnd 0.005886f
C2343 vdd.n33 gnd 0.00249f
C2344 vdd.n34 gnd 0.002637f
C2345 vdd.n35 gnd 0.004634f
C2346 vdd.n36 gnd 0.00249f
C2347 vdd.n37 gnd 0.005886f
C2348 vdd.n38 gnd 0.002637f
C2349 vdd.n39 gnd 0.004634f
C2350 vdd.n40 gnd 0.00249f
C2351 vdd.n41 gnd 0.004414f
C2352 vdd.n42 gnd 0.004427f
C2353 vdd.t132 gnd 0.012645f
C2354 vdd.n43 gnd 0.028134f
C2355 vdd.n44 gnd 0.146416f
C2356 vdd.n45 gnd 0.00249f
C2357 vdd.n46 gnd 0.002637f
C2358 vdd.n47 gnd 0.005886f
C2359 vdd.n48 gnd 0.005886f
C2360 vdd.n49 gnd 0.002637f
C2361 vdd.n50 gnd 0.00249f
C2362 vdd.n51 gnd 0.004634f
C2363 vdd.n52 gnd 0.004634f
C2364 vdd.n53 gnd 0.00249f
C2365 vdd.n54 gnd 0.002637f
C2366 vdd.n55 gnd 0.005886f
C2367 vdd.n56 gnd 0.005886f
C2368 vdd.n57 gnd 0.002637f
C2369 vdd.n58 gnd 0.00249f
C2370 vdd.n59 gnd 0.004634f
C2371 vdd.n60 gnd 0.004634f
C2372 vdd.n61 gnd 0.00249f
C2373 vdd.n62 gnd 0.002637f
C2374 vdd.n63 gnd 0.005886f
C2375 vdd.n64 gnd 0.005886f
C2376 vdd.n65 gnd 0.013915f
C2377 vdd.n66 gnd 0.002563f
C2378 vdd.n67 gnd 0.00249f
C2379 vdd.n68 gnd 0.011977f
C2380 vdd.n69 gnd 0.008362f
C2381 vdd.t190 gnd 0.029295f
C2382 vdd.t135 gnd 0.029295f
C2383 vdd.n70 gnd 0.201332f
C2384 vdd.n71 gnd 0.158317f
C2385 vdd.t118 gnd 0.029295f
C2386 vdd.t7 gnd 0.029295f
C2387 vdd.n72 gnd 0.201332f
C2388 vdd.n73 gnd 0.127761f
C2389 vdd.t139 gnd 0.029295f
C2390 vdd.t195 gnd 0.029295f
C2391 vdd.n74 gnd 0.201332f
C2392 vdd.n75 gnd 0.127761f
C2393 vdd.n76 gnd 0.004994f
C2394 vdd.n77 gnd 0.004634f
C2395 vdd.n78 gnd 0.002563f
C2396 vdd.n79 gnd 0.005886f
C2397 vdd.n80 gnd 0.00249f
C2398 vdd.n81 gnd 0.002637f
C2399 vdd.n82 gnd 0.004634f
C2400 vdd.n83 gnd 0.00249f
C2401 vdd.n84 gnd 0.005886f
C2402 vdd.n85 gnd 0.002637f
C2403 vdd.n86 gnd 0.004634f
C2404 vdd.n87 gnd 0.00249f
C2405 vdd.n88 gnd 0.004414f
C2406 vdd.n89 gnd 0.004427f
C2407 vdd.t111 gnd 0.012645f
C2408 vdd.n90 gnd 0.028134f
C2409 vdd.n91 gnd 0.146416f
C2410 vdd.n92 gnd 0.00249f
C2411 vdd.n93 gnd 0.002637f
C2412 vdd.n94 gnd 0.005886f
C2413 vdd.n95 gnd 0.005886f
C2414 vdd.n96 gnd 0.002637f
C2415 vdd.n97 gnd 0.00249f
C2416 vdd.n98 gnd 0.004634f
C2417 vdd.n99 gnd 0.004634f
C2418 vdd.n100 gnd 0.00249f
C2419 vdd.n101 gnd 0.002637f
C2420 vdd.n102 gnd 0.005886f
C2421 vdd.n103 gnd 0.005886f
C2422 vdd.n104 gnd 0.002637f
C2423 vdd.n105 gnd 0.00249f
C2424 vdd.n106 gnd 0.004634f
C2425 vdd.n107 gnd 0.004634f
C2426 vdd.n108 gnd 0.00249f
C2427 vdd.n109 gnd 0.002637f
C2428 vdd.n110 gnd 0.005886f
C2429 vdd.n111 gnd 0.005886f
C2430 vdd.n112 gnd 0.013915f
C2431 vdd.n113 gnd 0.002563f
C2432 vdd.n114 gnd 0.00249f
C2433 vdd.n115 gnd 0.011977f
C2434 vdd.n116 gnd 0.008099f
C2435 vdd.n117 gnd 0.095055f
C2436 vdd.n118 gnd 0.004994f
C2437 vdd.n119 gnd 0.004634f
C2438 vdd.n120 gnd 0.002563f
C2439 vdd.n121 gnd 0.005886f
C2440 vdd.n122 gnd 0.00249f
C2441 vdd.n123 gnd 0.002637f
C2442 vdd.n124 gnd 0.004634f
C2443 vdd.n125 gnd 0.00249f
C2444 vdd.n126 gnd 0.005886f
C2445 vdd.n127 gnd 0.002637f
C2446 vdd.n128 gnd 0.004634f
C2447 vdd.n129 gnd 0.00249f
C2448 vdd.n130 gnd 0.004414f
C2449 vdd.n131 gnd 0.004427f
C2450 vdd.t142 gnd 0.012645f
C2451 vdd.n132 gnd 0.028134f
C2452 vdd.n133 gnd 0.146416f
C2453 vdd.n134 gnd 0.00249f
C2454 vdd.n135 gnd 0.002637f
C2455 vdd.n136 gnd 0.005886f
C2456 vdd.n137 gnd 0.005886f
C2457 vdd.n138 gnd 0.002637f
C2458 vdd.n139 gnd 0.00249f
C2459 vdd.n140 gnd 0.004634f
C2460 vdd.n141 gnd 0.004634f
C2461 vdd.n142 gnd 0.00249f
C2462 vdd.n143 gnd 0.002637f
C2463 vdd.n144 gnd 0.005886f
C2464 vdd.n145 gnd 0.005886f
C2465 vdd.n146 gnd 0.002637f
C2466 vdd.n147 gnd 0.00249f
C2467 vdd.n148 gnd 0.004634f
C2468 vdd.n149 gnd 0.004634f
C2469 vdd.n150 gnd 0.00249f
C2470 vdd.n151 gnd 0.002637f
C2471 vdd.n152 gnd 0.005886f
C2472 vdd.n153 gnd 0.005886f
C2473 vdd.n154 gnd 0.013915f
C2474 vdd.n155 gnd 0.002563f
C2475 vdd.n156 gnd 0.00249f
C2476 vdd.n157 gnd 0.011977f
C2477 vdd.n158 gnd 0.008362f
C2478 vdd.t143 gnd 0.029295f
C2479 vdd.t116 gnd 0.029295f
C2480 vdd.n159 gnd 0.201332f
C2481 vdd.n160 gnd 0.158317f
C2482 vdd.t134 gnd 0.029295f
C2483 vdd.t136 gnd 0.029295f
C2484 vdd.n161 gnd 0.201332f
C2485 vdd.n162 gnd 0.127761f
C2486 vdd.t191 gnd 0.029295f
C2487 vdd.t199 gnd 0.029295f
C2488 vdd.n163 gnd 0.201332f
C2489 vdd.n164 gnd 0.127761f
C2490 vdd.n165 gnd 0.004994f
C2491 vdd.n166 gnd 0.004634f
C2492 vdd.n167 gnd 0.002563f
C2493 vdd.n168 gnd 0.005886f
C2494 vdd.n169 gnd 0.00249f
C2495 vdd.n170 gnd 0.002637f
C2496 vdd.n171 gnd 0.004634f
C2497 vdd.n172 gnd 0.00249f
C2498 vdd.n173 gnd 0.005886f
C2499 vdd.n174 gnd 0.002637f
C2500 vdd.n175 gnd 0.004634f
C2501 vdd.n176 gnd 0.00249f
C2502 vdd.n177 gnd 0.004414f
C2503 vdd.n178 gnd 0.004427f
C2504 vdd.t133 gnd 0.012645f
C2505 vdd.n179 gnd 0.028134f
C2506 vdd.n180 gnd 0.146416f
C2507 vdd.n181 gnd 0.00249f
C2508 vdd.n182 gnd 0.002637f
C2509 vdd.n183 gnd 0.005886f
C2510 vdd.n184 gnd 0.005886f
C2511 vdd.n185 gnd 0.002637f
C2512 vdd.n186 gnd 0.00249f
C2513 vdd.n187 gnd 0.004634f
C2514 vdd.n188 gnd 0.004634f
C2515 vdd.n189 gnd 0.00249f
C2516 vdd.n190 gnd 0.002637f
C2517 vdd.n191 gnd 0.005886f
C2518 vdd.n192 gnd 0.005886f
C2519 vdd.n193 gnd 0.002637f
C2520 vdd.n194 gnd 0.00249f
C2521 vdd.n195 gnd 0.004634f
C2522 vdd.n196 gnd 0.004634f
C2523 vdd.n197 gnd 0.00249f
C2524 vdd.n198 gnd 0.002637f
C2525 vdd.n199 gnd 0.005886f
C2526 vdd.n200 gnd 0.005886f
C2527 vdd.n201 gnd 0.013915f
C2528 vdd.n202 gnd 0.002563f
C2529 vdd.n203 gnd 0.00249f
C2530 vdd.n204 gnd 0.011977f
C2531 vdd.n205 gnd 0.008099f
C2532 vdd.n206 gnd 0.056548f
C2533 vdd.n207 gnd 0.203758f
C2534 vdd.n208 gnd 0.004994f
C2535 vdd.n209 gnd 0.004634f
C2536 vdd.n210 gnd 0.002563f
C2537 vdd.n211 gnd 0.005886f
C2538 vdd.n212 gnd 0.00249f
C2539 vdd.n213 gnd 0.002637f
C2540 vdd.n214 gnd 0.004634f
C2541 vdd.n215 gnd 0.00249f
C2542 vdd.n216 gnd 0.005886f
C2543 vdd.n217 gnd 0.002637f
C2544 vdd.n218 gnd 0.004634f
C2545 vdd.n219 gnd 0.00249f
C2546 vdd.n220 gnd 0.004414f
C2547 vdd.n221 gnd 0.004427f
C2548 vdd.t104 gnd 0.012645f
C2549 vdd.n222 gnd 0.028134f
C2550 vdd.n223 gnd 0.146416f
C2551 vdd.n224 gnd 0.00249f
C2552 vdd.n225 gnd 0.002637f
C2553 vdd.n226 gnd 0.005886f
C2554 vdd.n227 gnd 0.005886f
C2555 vdd.n228 gnd 0.002637f
C2556 vdd.n229 gnd 0.00249f
C2557 vdd.n230 gnd 0.004634f
C2558 vdd.n231 gnd 0.004634f
C2559 vdd.n232 gnd 0.00249f
C2560 vdd.n233 gnd 0.002637f
C2561 vdd.n234 gnd 0.005886f
C2562 vdd.n235 gnd 0.005886f
C2563 vdd.n236 gnd 0.002637f
C2564 vdd.n237 gnd 0.00249f
C2565 vdd.n238 gnd 0.004634f
C2566 vdd.n239 gnd 0.004634f
C2567 vdd.n240 gnd 0.00249f
C2568 vdd.n241 gnd 0.002637f
C2569 vdd.n242 gnd 0.005886f
C2570 vdd.n243 gnd 0.005886f
C2571 vdd.n244 gnd 0.013915f
C2572 vdd.n245 gnd 0.002563f
C2573 vdd.n246 gnd 0.00249f
C2574 vdd.n247 gnd 0.011977f
C2575 vdd.n248 gnd 0.008362f
C2576 vdd.t114 gnd 0.029295f
C2577 vdd.t110 gnd 0.029295f
C2578 vdd.n249 gnd 0.201332f
C2579 vdd.n250 gnd 0.158317f
C2580 vdd.t140 gnd 0.029295f
C2581 vdd.t197 gnd 0.029295f
C2582 vdd.n251 gnd 0.201332f
C2583 vdd.n252 gnd 0.127761f
C2584 vdd.t123 gnd 0.029295f
C2585 vdd.t1 gnd 0.029295f
C2586 vdd.n253 gnd 0.201332f
C2587 vdd.n254 gnd 0.127761f
C2588 vdd.n255 gnd 0.004994f
C2589 vdd.n256 gnd 0.004634f
C2590 vdd.n257 gnd 0.002563f
C2591 vdd.n258 gnd 0.005886f
C2592 vdd.n259 gnd 0.00249f
C2593 vdd.n260 gnd 0.002637f
C2594 vdd.n261 gnd 0.004634f
C2595 vdd.n262 gnd 0.00249f
C2596 vdd.n263 gnd 0.005886f
C2597 vdd.n264 gnd 0.002637f
C2598 vdd.n265 gnd 0.004634f
C2599 vdd.n266 gnd 0.00249f
C2600 vdd.n267 gnd 0.004414f
C2601 vdd.n268 gnd 0.004427f
C2602 vdd.t15 gnd 0.012645f
C2603 vdd.n269 gnd 0.028134f
C2604 vdd.n270 gnd 0.146416f
C2605 vdd.n271 gnd 0.00249f
C2606 vdd.n272 gnd 0.002637f
C2607 vdd.n273 gnd 0.005886f
C2608 vdd.n274 gnd 0.005886f
C2609 vdd.n275 gnd 0.002637f
C2610 vdd.n276 gnd 0.00249f
C2611 vdd.n277 gnd 0.004634f
C2612 vdd.n278 gnd 0.004634f
C2613 vdd.n279 gnd 0.00249f
C2614 vdd.n280 gnd 0.002637f
C2615 vdd.n281 gnd 0.005886f
C2616 vdd.n282 gnd 0.005886f
C2617 vdd.n283 gnd 0.002637f
C2618 vdd.n284 gnd 0.00249f
C2619 vdd.n285 gnd 0.004634f
C2620 vdd.n286 gnd 0.004634f
C2621 vdd.n287 gnd 0.00249f
C2622 vdd.n288 gnd 0.002637f
C2623 vdd.n289 gnd 0.005886f
C2624 vdd.n290 gnd 0.005886f
C2625 vdd.n291 gnd 0.013915f
C2626 vdd.n292 gnd 0.002563f
C2627 vdd.n293 gnd 0.00249f
C2628 vdd.n294 gnd 0.011977f
C2629 vdd.n295 gnd 0.008099f
C2630 vdd.n296 gnd 0.056548f
C2631 vdd.n297 gnd 0.220543f
C2632 vdd.n298 gnd 0.006993f
C2633 vdd.n299 gnd 0.009099f
C2634 vdd.n300 gnd 0.007324f
C2635 vdd.n301 gnd 0.007324f
C2636 vdd.n302 gnd 0.009099f
C2637 vdd.n303 gnd 0.009099f
C2638 vdd.n304 gnd 0.664865f
C2639 vdd.n305 gnd 0.009099f
C2640 vdd.n306 gnd 0.009099f
C2641 vdd.n307 gnd 0.009099f
C2642 vdd.n308 gnd 0.720658f
C2643 vdd.n309 gnd 0.009099f
C2644 vdd.n310 gnd 0.009099f
C2645 vdd.n311 gnd 0.009099f
C2646 vdd.n312 gnd 0.009099f
C2647 vdd.n313 gnd 0.007324f
C2648 vdd.n314 gnd 0.009099f
C2649 vdd.t0 gnd 0.46494f
C2650 vdd.n315 gnd 0.009099f
C2651 vdd.n316 gnd 0.009099f
C2652 vdd.n317 gnd 0.009099f
C2653 vdd.n318 gnd 0.929881f
C2654 vdd.n319 gnd 0.009099f
C2655 vdd.n320 gnd 0.009099f
C2656 vdd.n321 gnd 0.009099f
C2657 vdd.n322 gnd 0.009099f
C2658 vdd.n323 gnd 0.009099f
C2659 vdd.n324 gnd 0.007324f
C2660 vdd.n325 gnd 0.009099f
C2661 vdd.n326 gnd 0.009099f
C2662 vdd.n327 gnd 0.009099f
C2663 vdd.n328 gnd 0.022175f
C2664 vdd.n329 gnd 2.22242f
C2665 vdd.n330 gnd 0.022684f
C2666 vdd.n331 gnd 0.009099f
C2667 vdd.n332 gnd 0.009099f
C2668 vdd.n334 gnd 0.009099f
C2669 vdd.n335 gnd 0.009099f
C2670 vdd.n336 gnd 0.007324f
C2671 vdd.n337 gnd 0.007324f
C2672 vdd.n338 gnd 0.009099f
C2673 vdd.n339 gnd 0.009099f
C2674 vdd.n340 gnd 0.009099f
C2675 vdd.n341 gnd 0.009099f
C2676 vdd.n342 gnd 0.009099f
C2677 vdd.n343 gnd 0.009099f
C2678 vdd.n344 gnd 0.007324f
C2679 vdd.n346 gnd 0.009099f
C2680 vdd.n347 gnd 0.009099f
C2681 vdd.n348 gnd 0.009099f
C2682 vdd.n349 gnd 0.009099f
C2683 vdd.n350 gnd 0.009099f
C2684 vdd.n351 gnd 0.007324f
C2685 vdd.n353 gnd 0.009099f
C2686 vdd.n354 gnd 0.009099f
C2687 vdd.n355 gnd 0.009099f
C2688 vdd.n356 gnd 0.009099f
C2689 vdd.n357 gnd 0.009099f
C2690 vdd.n358 gnd 0.007324f
C2691 vdd.n360 gnd 0.009099f
C2692 vdd.n361 gnd 0.009099f
C2693 vdd.n362 gnd 0.009099f
C2694 vdd.n363 gnd 0.009099f
C2695 vdd.n364 gnd 0.006115f
C2696 vdd.t51 gnd 0.111942f
C2697 vdd.t50 gnd 0.119636f
C2698 vdd.t49 gnd 0.146195f
C2699 vdd.n365 gnd 0.187402f
C2700 vdd.n366 gnd 0.158184f
C2701 vdd.n368 gnd 0.009099f
C2702 vdd.n369 gnd 0.009099f
C2703 vdd.n370 gnd 0.007324f
C2704 vdd.n371 gnd 0.009099f
C2705 vdd.n373 gnd 0.009099f
C2706 vdd.n374 gnd 0.009099f
C2707 vdd.n375 gnd 0.009099f
C2708 vdd.n376 gnd 0.009099f
C2709 vdd.n377 gnd 0.007324f
C2710 vdd.n379 gnd 0.009099f
C2711 vdd.n380 gnd 0.009099f
C2712 vdd.n381 gnd 0.009099f
C2713 vdd.n382 gnd 0.009099f
C2714 vdd.n383 gnd 0.009099f
C2715 vdd.n384 gnd 0.007324f
C2716 vdd.n386 gnd 0.009099f
C2717 vdd.n387 gnd 0.009099f
C2718 vdd.n388 gnd 0.009099f
C2719 vdd.n389 gnd 0.009099f
C2720 vdd.n390 gnd 0.009099f
C2721 vdd.n391 gnd 0.007324f
C2722 vdd.n393 gnd 0.009099f
C2723 vdd.n394 gnd 0.009099f
C2724 vdd.n395 gnd 0.009099f
C2725 vdd.n396 gnd 0.009099f
C2726 vdd.n397 gnd 0.009099f
C2727 vdd.n398 gnd 0.007324f
C2728 vdd.n400 gnd 0.009099f
C2729 vdd.n401 gnd 0.009099f
C2730 vdd.n402 gnd 0.009099f
C2731 vdd.n403 gnd 0.009099f
C2732 vdd.n404 gnd 0.00725f
C2733 vdd.t45 gnd 0.111942f
C2734 vdd.t44 gnd 0.119636f
C2735 vdd.t42 gnd 0.146195f
C2736 vdd.n405 gnd 0.187402f
C2737 vdd.n406 gnd 0.158184f
C2738 vdd.n408 gnd 0.009099f
C2739 vdd.n409 gnd 0.009099f
C2740 vdd.n410 gnd 0.007324f
C2741 vdd.n411 gnd 0.009099f
C2742 vdd.n413 gnd 0.009099f
C2743 vdd.n414 gnd 0.009099f
C2744 vdd.n415 gnd 0.009099f
C2745 vdd.n416 gnd 0.009099f
C2746 vdd.n417 gnd 0.007324f
C2747 vdd.n419 gnd 0.009099f
C2748 vdd.n420 gnd 0.009099f
C2749 vdd.n421 gnd 0.009099f
C2750 vdd.n422 gnd 0.009099f
C2751 vdd.n423 gnd 0.009099f
C2752 vdd.n424 gnd 0.007324f
C2753 vdd.n426 gnd 0.009099f
C2754 vdd.n427 gnd 0.009099f
C2755 vdd.n428 gnd 0.009099f
C2756 vdd.n429 gnd 0.009099f
C2757 vdd.n430 gnd 0.009099f
C2758 vdd.n431 gnd 0.007324f
C2759 vdd.n433 gnd 0.009099f
C2760 vdd.n434 gnd 0.009099f
C2761 vdd.n435 gnd 0.009099f
C2762 vdd.n436 gnd 0.009099f
C2763 vdd.n437 gnd 0.009099f
C2764 vdd.n438 gnd 0.007324f
C2765 vdd.n440 gnd 0.009099f
C2766 vdd.n441 gnd 0.009099f
C2767 vdd.n442 gnd 0.009099f
C2768 vdd.n443 gnd 0.009099f
C2769 vdd.n444 gnd 0.009099f
C2770 vdd.n445 gnd 0.009099f
C2771 vdd.n446 gnd 0.007324f
C2772 vdd.n447 gnd 0.009099f
C2773 vdd.n448 gnd 0.009099f
C2774 vdd.n449 gnd 0.007324f
C2775 vdd.n450 gnd 0.009099f
C2776 vdd.n451 gnd 0.007324f
C2777 vdd.n452 gnd 0.009099f
C2778 vdd.n453 gnd 0.007324f
C2779 vdd.n454 gnd 0.009099f
C2780 vdd.n455 gnd 0.009099f
C2781 vdd.n456 gnd 0.506785f
C2782 vdd.t117 gnd 0.46494f
C2783 vdd.n457 gnd 0.009099f
C2784 vdd.n458 gnd 0.007324f
C2785 vdd.n459 gnd 0.009099f
C2786 vdd.n460 gnd 0.007324f
C2787 vdd.n461 gnd 0.009099f
C2788 vdd.t113 gnd 0.46494f
C2789 vdd.n462 gnd 0.009099f
C2790 vdd.n463 gnd 0.007324f
C2791 vdd.n464 gnd 0.009099f
C2792 vdd.n465 gnd 0.007324f
C2793 vdd.n466 gnd 0.009099f
C2794 vdd.t103 gnd 0.46494f
C2795 vdd.n467 gnd 0.581176f
C2796 vdd.n468 gnd 0.009099f
C2797 vdd.n469 gnd 0.007324f
C2798 vdd.n470 gnd 0.009099f
C2799 vdd.n471 gnd 0.007324f
C2800 vdd.n472 gnd 0.009099f
C2801 vdd.n473 gnd 0.929881f
C2802 vdd.n474 gnd 0.009099f
C2803 vdd.n475 gnd 0.007324f
C2804 vdd.n476 gnd 0.022175f
C2805 vdd.n477 gnd 0.006079f
C2806 vdd.n478 gnd 0.022175f
C2807 vdd.t21 gnd 0.46494f
C2808 vdd.n479 gnd 0.022175f
C2809 vdd.n480 gnd 0.006079f
C2810 vdd.n481 gnd 0.007825f
C2811 vdd.n482 gnd 0.007324f
C2812 vdd.n483 gnd 0.009099f
C2813 vdd.n484 gnd 6.40688f
C2814 vdd.n515 gnd 0.022684f
C2815 vdd.n516 gnd 1.27859f
C2816 vdd.n517 gnd 0.009099f
C2817 vdd.n518 gnd 0.007324f
C2818 vdd.n519 gnd 0.005823f
C2819 vdd.n520 gnd 0.014868f
C2820 vdd.n521 gnd 0.007324f
C2821 vdd.n522 gnd 0.009099f
C2822 vdd.n523 gnd 0.009099f
C2823 vdd.n524 gnd 0.009099f
C2824 vdd.n525 gnd 0.009099f
C2825 vdd.n526 gnd 0.009099f
C2826 vdd.n527 gnd 0.009099f
C2827 vdd.n528 gnd 0.009099f
C2828 vdd.n529 gnd 0.009099f
C2829 vdd.n530 gnd 0.009099f
C2830 vdd.n531 gnd 0.009099f
C2831 vdd.n532 gnd 0.009099f
C2832 vdd.n533 gnd 0.009099f
C2833 vdd.n534 gnd 0.009099f
C2834 vdd.n535 gnd 0.009099f
C2835 vdd.n536 gnd 0.006115f
C2836 vdd.n537 gnd 0.009099f
C2837 vdd.n538 gnd 0.009099f
C2838 vdd.n539 gnd 0.009099f
C2839 vdd.n540 gnd 0.009099f
C2840 vdd.n541 gnd 0.009099f
C2841 vdd.n542 gnd 0.009099f
C2842 vdd.n543 gnd 0.009099f
C2843 vdd.n544 gnd 0.009099f
C2844 vdd.n545 gnd 0.009099f
C2845 vdd.n546 gnd 0.009099f
C2846 vdd.n547 gnd 0.009099f
C2847 vdd.n548 gnd 0.009099f
C2848 vdd.n549 gnd 0.009099f
C2849 vdd.n550 gnd 0.009099f
C2850 vdd.n551 gnd 0.009099f
C2851 vdd.n552 gnd 0.009099f
C2852 vdd.n553 gnd 0.009099f
C2853 vdd.n554 gnd 0.009099f
C2854 vdd.n555 gnd 0.009099f
C2855 vdd.n556 gnd 0.00725f
C2856 vdd.t22 gnd 0.111942f
C2857 vdd.t23 gnd 0.119636f
C2858 vdd.t20 gnd 0.146195f
C2859 vdd.n557 gnd 0.187402f
C2860 vdd.n558 gnd 0.157451f
C2861 vdd.n559 gnd 0.009099f
C2862 vdd.n560 gnd 0.009099f
C2863 vdd.n561 gnd 0.009099f
C2864 vdd.n562 gnd 0.009099f
C2865 vdd.n563 gnd 0.009099f
C2866 vdd.n564 gnd 0.009099f
C2867 vdd.n565 gnd 0.009099f
C2868 vdd.n566 gnd 0.009099f
C2869 vdd.n567 gnd 0.009099f
C2870 vdd.n568 gnd 0.009099f
C2871 vdd.n569 gnd 0.009099f
C2872 vdd.n570 gnd 0.009099f
C2873 vdd.n571 gnd 0.009099f
C2874 vdd.n572 gnd 0.005823f
C2875 vdd.n575 gnd 0.006187f
C2876 vdd.n576 gnd 0.006187f
C2877 vdd.n577 gnd 0.006187f
C2878 vdd.n578 gnd 0.006187f
C2879 vdd.n579 gnd 0.006187f
C2880 vdd.n580 gnd 0.006187f
C2881 vdd.n582 gnd 0.006187f
C2882 vdd.n583 gnd 0.006187f
C2883 vdd.n585 gnd 0.006187f
C2884 vdd.n586 gnd 0.004504f
C2885 vdd.n588 gnd 0.006187f
C2886 vdd.t69 gnd 0.25003f
C2887 vdd.t68 gnd 0.255937f
C2888 vdd.t67 gnd 0.163229f
C2889 vdd.n589 gnd 0.088216f
C2890 vdd.n590 gnd 0.050039f
C2891 vdd.n591 gnd 0.008843f
C2892 vdd.n592 gnd 0.014461f
C2893 vdd.n594 gnd 0.006187f
C2894 vdd.n595 gnd 0.632319f
C2895 vdd.n596 gnd 0.013708f
C2896 vdd.n597 gnd 0.013708f
C2897 vdd.n598 gnd 0.006187f
C2898 vdd.n599 gnd 0.014682f
C2899 vdd.n600 gnd 0.006187f
C2900 vdd.n601 gnd 0.006187f
C2901 vdd.n602 gnd 0.006187f
C2902 vdd.n603 gnd 0.006187f
C2903 vdd.n604 gnd 0.006187f
C2904 vdd.n606 gnd 0.006187f
C2905 vdd.n607 gnd 0.006187f
C2906 vdd.n609 gnd 0.006187f
C2907 vdd.n610 gnd 0.006187f
C2908 vdd.n612 gnd 0.006187f
C2909 vdd.n613 gnd 0.006187f
C2910 vdd.n615 gnd 0.006187f
C2911 vdd.n616 gnd 0.006187f
C2912 vdd.n618 gnd 0.006187f
C2913 vdd.n619 gnd 0.006187f
C2914 vdd.n621 gnd 0.006187f
C2915 vdd.t59 gnd 0.25003f
C2916 vdd.t58 gnd 0.255937f
C2917 vdd.t56 gnd 0.163229f
C2918 vdd.n622 gnd 0.088216f
C2919 vdd.n623 gnd 0.050039f
C2920 vdd.n624 gnd 0.006187f
C2921 vdd.n626 gnd 0.006187f
C2922 vdd.n627 gnd 0.006187f
C2923 vdd.t57 gnd 0.316159f
C2924 vdd.n628 gnd 0.006187f
C2925 vdd.n629 gnd 0.006187f
C2926 vdd.n630 gnd 0.006187f
C2927 vdd.n631 gnd 0.006187f
C2928 vdd.n632 gnd 0.006187f
C2929 vdd.n633 gnd 0.632319f
C2930 vdd.n634 gnd 0.006187f
C2931 vdd.n635 gnd 0.006187f
C2932 vdd.n636 gnd 0.553279f
C2933 vdd.n637 gnd 0.006187f
C2934 vdd.n638 gnd 0.006187f
C2935 vdd.n639 gnd 0.005459f
C2936 vdd.n640 gnd 0.006187f
C2937 vdd.n641 gnd 0.557929f
C2938 vdd.n642 gnd 0.006187f
C2939 vdd.n643 gnd 0.006187f
C2940 vdd.n644 gnd 0.006187f
C2941 vdd.n645 gnd 0.006187f
C2942 vdd.n646 gnd 0.006187f
C2943 vdd.n647 gnd 0.632319f
C2944 vdd.n648 gnd 0.006187f
C2945 vdd.n649 gnd 0.006187f
C2946 vdd.t36 gnd 0.283614f
C2947 vdd.t153 gnd 0.074391f
C2948 vdd.n650 gnd 0.006187f
C2949 vdd.n651 gnd 0.006187f
C2950 vdd.n652 gnd 0.006187f
C2951 vdd.t162 gnd 0.316159f
C2952 vdd.n653 gnd 0.006187f
C2953 vdd.n654 gnd 0.006187f
C2954 vdd.n655 gnd 0.006187f
C2955 vdd.n656 gnd 0.006187f
C2956 vdd.n657 gnd 0.006187f
C2957 vdd.t176 gnd 0.316159f
C2958 vdd.n658 gnd 0.006187f
C2959 vdd.n659 gnd 0.006187f
C2960 vdd.n660 gnd 0.525383f
C2961 vdd.n661 gnd 0.006187f
C2962 vdd.n662 gnd 0.006187f
C2963 vdd.n663 gnd 0.006187f
C2964 vdd.n664 gnd 0.385901f
C2965 vdd.n665 gnd 0.006187f
C2966 vdd.n666 gnd 0.006187f
C2967 vdd.t158 gnd 0.316159f
C2968 vdd.n667 gnd 0.006187f
C2969 vdd.n668 gnd 0.006187f
C2970 vdd.n669 gnd 0.006187f
C2971 vdd.n670 gnd 0.525383f
C2972 vdd.n671 gnd 0.006187f
C2973 vdd.n672 gnd 0.006187f
C2974 vdd.t145 gnd 0.269665f
C2975 vdd.t187 gnd 0.246418f
C2976 vdd.n673 gnd 0.006187f
C2977 vdd.n674 gnd 0.006187f
C2978 vdd.n675 gnd 0.006187f
C2979 vdd.t180 gnd 0.316159f
C2980 vdd.n676 gnd 0.006187f
C2981 vdd.n677 gnd 0.006187f
C2982 vdd.t177 gnd 0.316159f
C2983 vdd.n678 gnd 0.006187f
C2984 vdd.n679 gnd 0.006187f
C2985 vdd.n680 gnd 0.006187f
C2986 vdd.t149 gnd 0.23247f
C2987 vdd.n681 gnd 0.006187f
C2988 vdd.n682 gnd 0.006187f
C2989 vdd.n683 gnd 0.539331f
C2990 vdd.n684 gnd 0.006187f
C2991 vdd.n685 gnd 0.006187f
C2992 vdd.n686 gnd 0.006187f
C2993 vdd.n687 gnd 0.632319f
C2994 vdd.n688 gnd 0.006187f
C2995 vdd.n689 gnd 0.006187f
C2996 vdd.t168 gnd 0.283614f
C2997 vdd.n690 gnd 0.399849f
C2998 vdd.n691 gnd 0.006187f
C2999 vdd.n692 gnd 0.006187f
C3000 vdd.n693 gnd 0.006187f
C3001 vdd.t150 gnd 0.316159f
C3002 vdd.n694 gnd 0.006187f
C3003 vdd.n695 gnd 0.006187f
C3004 vdd.n696 gnd 0.006187f
C3005 vdd.n697 gnd 0.006187f
C3006 vdd.n698 gnd 0.006187f
C3007 vdd.t172 gnd 0.632319f
C3008 vdd.n699 gnd 0.006187f
C3009 vdd.n700 gnd 0.006187f
C3010 vdd.t61 gnd 0.316159f
C3011 vdd.n701 gnd 0.006187f
C3012 vdd.n702 gnd 0.014682f
C3013 vdd.n703 gnd 0.014682f
C3014 vdd.t170 gnd 0.595124f
C3015 vdd.n704 gnd 0.013708f
C3016 vdd.n705 gnd 0.013708f
C3017 vdd.n706 gnd 0.014682f
C3018 vdd.n707 gnd 0.006187f
C3019 vdd.n708 gnd 0.006187f
C3020 vdd.t184 gnd 0.595124f
C3021 vdd.n726 gnd 0.014682f
C3022 vdd.n744 gnd 0.013708f
C3023 vdd.n745 gnd 0.006187f
C3024 vdd.n746 gnd 0.013708f
C3025 vdd.t85 gnd 0.25003f
C3026 vdd.t84 gnd 0.255937f
C3027 vdd.t83 gnd 0.163229f
C3028 vdd.n747 gnd 0.088216f
C3029 vdd.n748 gnd 0.050039f
C3030 vdd.n749 gnd 0.014461f
C3031 vdd.n750 gnd 0.006187f
C3032 vdd.t182 gnd 0.632319f
C3033 vdd.n751 gnd 0.013708f
C3034 vdd.n752 gnd 0.006187f
C3035 vdd.n753 gnd 0.014682f
C3036 vdd.n754 gnd 0.006187f
C3037 vdd.t55 gnd 0.25003f
C3038 vdd.t54 gnd 0.255937f
C3039 vdd.t52 gnd 0.163229f
C3040 vdd.n755 gnd 0.088216f
C3041 vdd.n756 gnd 0.050039f
C3042 vdd.n757 gnd 0.008843f
C3043 vdd.n758 gnd 0.006187f
C3044 vdd.n759 gnd 0.006187f
C3045 vdd.t53 gnd 0.316159f
C3046 vdd.n760 gnd 0.006187f
C3047 vdd.n761 gnd 0.006187f
C3048 vdd.n762 gnd 0.006187f
C3049 vdd.n763 gnd 0.006187f
C3050 vdd.n764 gnd 0.006187f
C3051 vdd.n765 gnd 0.006187f
C3052 vdd.n766 gnd 0.632319f
C3053 vdd.n767 gnd 0.006187f
C3054 vdd.n768 gnd 0.006187f
C3055 vdd.t160 gnd 0.316159f
C3056 vdd.n769 gnd 0.006187f
C3057 vdd.n770 gnd 0.006187f
C3058 vdd.n771 gnd 0.006187f
C3059 vdd.n772 gnd 0.006187f
C3060 vdd.n773 gnd 0.399849f
C3061 vdd.n774 gnd 0.006187f
C3062 vdd.n775 gnd 0.006187f
C3063 vdd.n776 gnd 0.006187f
C3064 vdd.n777 gnd 0.006187f
C3065 vdd.n778 gnd 0.006187f
C3066 vdd.n779 gnd 0.539331f
C3067 vdd.n780 gnd 0.006187f
C3068 vdd.n781 gnd 0.006187f
C3069 vdd.t174 gnd 0.283614f
C3070 vdd.t146 gnd 0.23247f
C3071 vdd.n782 gnd 0.006187f
C3072 vdd.n783 gnd 0.006187f
C3073 vdd.n784 gnd 0.006187f
C3074 vdd.t167 gnd 0.316159f
C3075 vdd.n785 gnd 0.006187f
C3076 vdd.n786 gnd 0.006187f
C3077 vdd.t147 gnd 0.316159f
C3078 vdd.n787 gnd 0.006187f
C3079 vdd.n788 gnd 0.006187f
C3080 vdd.n789 gnd 0.006187f
C3081 vdd.t163 gnd 0.246418f
C3082 vdd.n790 gnd 0.006187f
C3083 vdd.n791 gnd 0.006187f
C3084 vdd.n792 gnd 0.525383f
C3085 vdd.n793 gnd 0.006187f
C3086 vdd.n794 gnd 0.006187f
C3087 vdd.n795 gnd 0.006187f
C3088 vdd.t178 gnd 0.316159f
C3089 vdd.n796 gnd 0.006187f
C3090 vdd.n797 gnd 0.006187f
C3091 vdd.t154 gnd 0.269665f
C3092 vdd.n798 gnd 0.385901f
C3093 vdd.n799 gnd 0.006187f
C3094 vdd.n800 gnd 0.006187f
C3095 vdd.n801 gnd 0.006187f
C3096 vdd.n802 gnd 0.525383f
C3097 vdd.n803 gnd 0.006187f
C3098 vdd.n804 gnd 0.006187f
C3099 vdd.t186 gnd 0.316159f
C3100 vdd.n805 gnd 0.006187f
C3101 vdd.n806 gnd 0.006187f
C3102 vdd.n807 gnd 0.006187f
C3103 vdd.n808 gnd 0.632319f
C3104 vdd.n809 gnd 0.006187f
C3105 vdd.n810 gnd 0.006187f
C3106 vdd.t157 gnd 0.316159f
C3107 vdd.n811 gnd 0.006187f
C3108 vdd.n812 gnd 0.006187f
C3109 vdd.n813 gnd 0.006187f
C3110 vdd.t152 gnd 0.074391f
C3111 vdd.n814 gnd 0.006187f
C3112 vdd.n815 gnd 0.006187f
C3113 vdd.n816 gnd 0.006187f
C3114 vdd.t72 gnd 0.255937f
C3115 vdd.t70 gnd 0.163229f
C3116 vdd.t73 gnd 0.255937f
C3117 vdd.n817 gnd 0.143847f
C3118 vdd.n818 gnd 0.006187f
C3119 vdd.n819 gnd 0.006187f
C3120 vdd.n820 gnd 0.632319f
C3121 vdd.n821 gnd 0.006187f
C3122 vdd.n822 gnd 0.006187f
C3123 vdd.t71 gnd 0.283614f
C3124 vdd.n823 gnd 0.557929f
C3125 vdd.n824 gnd 0.006187f
C3126 vdd.n825 gnd 0.006187f
C3127 vdd.n826 gnd 0.006187f
C3128 vdd.n827 gnd 0.553279f
C3129 vdd.n828 gnd 0.006187f
C3130 vdd.n829 gnd 0.006187f
C3131 vdd.n830 gnd 0.006187f
C3132 vdd.n831 gnd 0.006187f
C3133 vdd.n832 gnd 0.006187f
C3134 vdd.n833 gnd 0.632319f
C3135 vdd.n834 gnd 0.006187f
C3136 vdd.n835 gnd 0.006187f
C3137 vdd.t17 gnd 0.316159f
C3138 vdd.n836 gnd 0.006187f
C3139 vdd.n837 gnd 0.014682f
C3140 vdd.n838 gnd 0.014682f
C3141 vdd.n839 gnd 6.40688f
C3142 vdd.n840 gnd 0.013708f
C3143 vdd.n841 gnd 0.013708f
C3144 vdd.n842 gnd 0.014682f
C3145 vdd.n843 gnd 0.006187f
C3146 vdd.n844 gnd 0.006187f
C3147 vdd.n845 gnd 0.006187f
C3148 vdd.n846 gnd 0.006187f
C3149 vdd.n847 gnd 0.006187f
C3150 vdd.n848 gnd 0.006187f
C3151 vdd.n849 gnd 0.006187f
C3152 vdd.n850 gnd 0.006187f
C3153 vdd.n852 gnd 0.006187f
C3154 vdd.n853 gnd 0.006187f
C3155 vdd.n854 gnd 0.005823f
C3156 vdd.n857 gnd 0.022684f
C3157 vdd.n858 gnd 0.007324f
C3158 vdd.n859 gnd 0.009099f
C3159 vdd.n861 gnd 0.009099f
C3160 vdd.n862 gnd 0.006079f
C3161 vdd.t28 gnd 0.46494f
C3162 vdd.n863 gnd 6.74164f
C3163 vdd.n864 gnd 0.009099f
C3164 vdd.n865 gnd 0.022684f
C3165 vdd.n866 gnd 0.007324f
C3166 vdd.n867 gnd 0.009099f
C3167 vdd.n868 gnd 0.007324f
C3168 vdd.n869 gnd 0.009099f
C3169 vdd.n870 gnd 0.929881f
C3170 vdd.n871 gnd 0.009099f
C3171 vdd.n872 gnd 0.007324f
C3172 vdd.n873 gnd 0.007324f
C3173 vdd.n874 gnd 0.009099f
C3174 vdd.n875 gnd 0.007324f
C3175 vdd.n876 gnd 0.009099f
C3176 vdd.t2 gnd 0.46494f
C3177 vdd.n877 gnd 0.009099f
C3178 vdd.n878 gnd 0.007324f
C3179 vdd.n879 gnd 0.009099f
C3180 vdd.n880 gnd 0.007324f
C3181 vdd.n881 gnd 0.009099f
C3182 vdd.t8 gnd 0.46494f
C3183 vdd.n882 gnd 0.009099f
C3184 vdd.n883 gnd 0.007324f
C3185 vdd.n884 gnd 0.009099f
C3186 vdd.n885 gnd 0.007324f
C3187 vdd.n886 gnd 0.009099f
C3188 vdd.n887 gnd 0.729956f
C3189 vdd.n888 gnd 0.771801f
C3190 vdd.t96 gnd 0.46494f
C3191 vdd.n889 gnd 0.009099f
C3192 vdd.n890 gnd 0.007324f
C3193 vdd.n891 gnd 0.004994f
C3194 vdd.n892 gnd 0.004634f
C3195 vdd.n893 gnd 0.002563f
C3196 vdd.n894 gnd 0.005886f
C3197 vdd.n895 gnd 0.00249f
C3198 vdd.n896 gnd 0.002637f
C3199 vdd.n897 gnd 0.004634f
C3200 vdd.n898 gnd 0.00249f
C3201 vdd.n899 gnd 0.005886f
C3202 vdd.n900 gnd 0.002637f
C3203 vdd.n901 gnd 0.004634f
C3204 vdd.n902 gnd 0.00249f
C3205 vdd.n903 gnd 0.004414f
C3206 vdd.n904 gnd 0.004427f
C3207 vdd.t3 gnd 0.012645f
C3208 vdd.n905 gnd 0.028134f
C3209 vdd.n906 gnd 0.146416f
C3210 vdd.n907 gnd 0.00249f
C3211 vdd.n908 gnd 0.002637f
C3212 vdd.n909 gnd 0.005886f
C3213 vdd.n910 gnd 0.005886f
C3214 vdd.n911 gnd 0.002637f
C3215 vdd.n912 gnd 0.00249f
C3216 vdd.n913 gnd 0.004634f
C3217 vdd.n914 gnd 0.004634f
C3218 vdd.n915 gnd 0.00249f
C3219 vdd.n916 gnd 0.002637f
C3220 vdd.n917 gnd 0.005886f
C3221 vdd.n918 gnd 0.005886f
C3222 vdd.n919 gnd 0.002637f
C3223 vdd.n920 gnd 0.00249f
C3224 vdd.n921 gnd 0.004634f
C3225 vdd.n922 gnd 0.004634f
C3226 vdd.n923 gnd 0.00249f
C3227 vdd.n924 gnd 0.002637f
C3228 vdd.n925 gnd 0.005886f
C3229 vdd.n926 gnd 0.005886f
C3230 vdd.n927 gnd 0.013915f
C3231 vdd.n928 gnd 0.002563f
C3232 vdd.n929 gnd 0.00249f
C3233 vdd.n930 gnd 0.011977f
C3234 vdd.n931 gnd 0.008362f
C3235 vdd.t192 gnd 0.029295f
C3236 vdd.t189 gnd 0.029295f
C3237 vdd.n932 gnd 0.201332f
C3238 vdd.n933 gnd 0.158317f
C3239 vdd.t141 gnd 0.029295f
C3240 vdd.t198 gnd 0.029295f
C3241 vdd.n934 gnd 0.201332f
C3242 vdd.n935 gnd 0.127761f
C3243 vdd.t196 gnd 0.029295f
C3244 vdd.t194 gnd 0.029295f
C3245 vdd.n936 gnd 0.201332f
C3246 vdd.n937 gnd 0.127761f
C3247 vdd.n938 gnd 0.004994f
C3248 vdd.n939 gnd 0.004634f
C3249 vdd.n940 gnd 0.002563f
C3250 vdd.n941 gnd 0.005886f
C3251 vdd.n942 gnd 0.00249f
C3252 vdd.n943 gnd 0.002637f
C3253 vdd.n944 gnd 0.004634f
C3254 vdd.n945 gnd 0.00249f
C3255 vdd.n946 gnd 0.005886f
C3256 vdd.n947 gnd 0.002637f
C3257 vdd.n948 gnd 0.004634f
C3258 vdd.n949 gnd 0.00249f
C3259 vdd.n950 gnd 0.004414f
C3260 vdd.n951 gnd 0.004427f
C3261 vdd.t193 gnd 0.012645f
C3262 vdd.n952 gnd 0.028134f
C3263 vdd.n953 gnd 0.146416f
C3264 vdd.n954 gnd 0.00249f
C3265 vdd.n955 gnd 0.002637f
C3266 vdd.n956 gnd 0.005886f
C3267 vdd.n957 gnd 0.005886f
C3268 vdd.n958 gnd 0.002637f
C3269 vdd.n959 gnd 0.00249f
C3270 vdd.n960 gnd 0.004634f
C3271 vdd.n961 gnd 0.004634f
C3272 vdd.n962 gnd 0.00249f
C3273 vdd.n963 gnd 0.002637f
C3274 vdd.n964 gnd 0.005886f
C3275 vdd.n965 gnd 0.005886f
C3276 vdd.n966 gnd 0.002637f
C3277 vdd.n967 gnd 0.00249f
C3278 vdd.n968 gnd 0.004634f
C3279 vdd.n969 gnd 0.004634f
C3280 vdd.n970 gnd 0.00249f
C3281 vdd.n971 gnd 0.002637f
C3282 vdd.n972 gnd 0.005886f
C3283 vdd.n973 gnd 0.005886f
C3284 vdd.n974 gnd 0.013915f
C3285 vdd.n975 gnd 0.002563f
C3286 vdd.n976 gnd 0.00249f
C3287 vdd.n977 gnd 0.011977f
C3288 vdd.n978 gnd 0.008099f
C3289 vdd.n979 gnd 0.095055f
C3290 vdd.n980 gnd 0.004994f
C3291 vdd.n981 gnd 0.004634f
C3292 vdd.n982 gnd 0.002563f
C3293 vdd.n983 gnd 0.005886f
C3294 vdd.n984 gnd 0.00249f
C3295 vdd.n985 gnd 0.002637f
C3296 vdd.n986 gnd 0.004634f
C3297 vdd.n987 gnd 0.00249f
C3298 vdd.n988 gnd 0.005886f
C3299 vdd.n989 gnd 0.002637f
C3300 vdd.n990 gnd 0.004634f
C3301 vdd.n991 gnd 0.00249f
C3302 vdd.n992 gnd 0.004414f
C3303 vdd.n993 gnd 0.004427f
C3304 vdd.t138 gnd 0.012645f
C3305 vdd.n994 gnd 0.028134f
C3306 vdd.n995 gnd 0.146416f
C3307 vdd.n996 gnd 0.00249f
C3308 vdd.n997 gnd 0.002637f
C3309 vdd.n998 gnd 0.005886f
C3310 vdd.n999 gnd 0.005886f
C3311 vdd.n1000 gnd 0.002637f
C3312 vdd.n1001 gnd 0.00249f
C3313 vdd.n1002 gnd 0.004634f
C3314 vdd.n1003 gnd 0.004634f
C3315 vdd.n1004 gnd 0.00249f
C3316 vdd.n1005 gnd 0.002637f
C3317 vdd.n1006 gnd 0.005886f
C3318 vdd.n1007 gnd 0.005886f
C3319 vdd.n1008 gnd 0.002637f
C3320 vdd.n1009 gnd 0.00249f
C3321 vdd.n1010 gnd 0.004634f
C3322 vdd.n1011 gnd 0.004634f
C3323 vdd.n1012 gnd 0.00249f
C3324 vdd.n1013 gnd 0.002637f
C3325 vdd.n1014 gnd 0.005886f
C3326 vdd.n1015 gnd 0.005886f
C3327 vdd.n1016 gnd 0.013915f
C3328 vdd.n1017 gnd 0.002563f
C3329 vdd.n1018 gnd 0.00249f
C3330 vdd.n1019 gnd 0.011977f
C3331 vdd.n1020 gnd 0.008362f
C3332 vdd.t97 gnd 0.029295f
C3333 vdd.t9 gnd 0.029295f
C3334 vdd.n1021 gnd 0.201332f
C3335 vdd.n1022 gnd 0.158317f
C3336 vdd.t124 gnd 0.029295f
C3337 vdd.t11 gnd 0.029295f
C3338 vdd.n1023 gnd 0.201332f
C3339 vdd.n1024 gnd 0.127761f
C3340 vdd.t106 gnd 0.029295f
C3341 vdd.t108 gnd 0.029295f
C3342 vdd.n1025 gnd 0.201332f
C3343 vdd.n1026 gnd 0.127761f
C3344 vdd.n1027 gnd 0.004994f
C3345 vdd.n1028 gnd 0.004634f
C3346 vdd.n1029 gnd 0.002563f
C3347 vdd.n1030 gnd 0.005886f
C3348 vdd.n1031 gnd 0.00249f
C3349 vdd.n1032 gnd 0.002637f
C3350 vdd.n1033 gnd 0.004634f
C3351 vdd.n1034 gnd 0.00249f
C3352 vdd.n1035 gnd 0.005886f
C3353 vdd.n1036 gnd 0.002637f
C3354 vdd.n1037 gnd 0.004634f
C3355 vdd.n1038 gnd 0.00249f
C3356 vdd.n1039 gnd 0.004414f
C3357 vdd.n1040 gnd 0.004427f
C3358 vdd.t112 gnd 0.012645f
C3359 vdd.n1041 gnd 0.028134f
C3360 vdd.n1042 gnd 0.146416f
C3361 vdd.n1043 gnd 0.00249f
C3362 vdd.n1044 gnd 0.002637f
C3363 vdd.n1045 gnd 0.005886f
C3364 vdd.n1046 gnd 0.005886f
C3365 vdd.n1047 gnd 0.002637f
C3366 vdd.n1048 gnd 0.00249f
C3367 vdd.n1049 gnd 0.004634f
C3368 vdd.n1050 gnd 0.004634f
C3369 vdd.n1051 gnd 0.00249f
C3370 vdd.n1052 gnd 0.002637f
C3371 vdd.n1053 gnd 0.005886f
C3372 vdd.n1054 gnd 0.005886f
C3373 vdd.n1055 gnd 0.002637f
C3374 vdd.n1056 gnd 0.00249f
C3375 vdd.n1057 gnd 0.004634f
C3376 vdd.n1058 gnd 0.004634f
C3377 vdd.n1059 gnd 0.00249f
C3378 vdd.n1060 gnd 0.002637f
C3379 vdd.n1061 gnd 0.005886f
C3380 vdd.n1062 gnd 0.005886f
C3381 vdd.n1063 gnd 0.013915f
C3382 vdd.n1064 gnd 0.002563f
C3383 vdd.n1065 gnd 0.00249f
C3384 vdd.n1066 gnd 0.011977f
C3385 vdd.n1067 gnd 0.008099f
C3386 vdd.n1068 gnd 0.056548f
C3387 vdd.n1069 gnd 0.203758f
C3388 vdd.n1070 gnd 0.004994f
C3389 vdd.n1071 gnd 0.004634f
C3390 vdd.n1072 gnd 0.002563f
C3391 vdd.n1073 gnd 0.005886f
C3392 vdd.n1074 gnd 0.00249f
C3393 vdd.n1075 gnd 0.002637f
C3394 vdd.n1076 gnd 0.004634f
C3395 vdd.n1077 gnd 0.00249f
C3396 vdd.n1078 gnd 0.005886f
C3397 vdd.n1079 gnd 0.002637f
C3398 vdd.n1080 gnd 0.004634f
C3399 vdd.n1081 gnd 0.00249f
C3400 vdd.n1082 gnd 0.004414f
C3401 vdd.n1083 gnd 0.004427f
C3402 vdd.t121 gnd 0.012645f
C3403 vdd.n1084 gnd 0.028134f
C3404 vdd.n1085 gnd 0.146416f
C3405 vdd.n1086 gnd 0.00249f
C3406 vdd.n1087 gnd 0.002637f
C3407 vdd.n1088 gnd 0.005886f
C3408 vdd.n1089 gnd 0.005886f
C3409 vdd.n1090 gnd 0.002637f
C3410 vdd.n1091 gnd 0.00249f
C3411 vdd.n1092 gnd 0.004634f
C3412 vdd.n1093 gnd 0.004634f
C3413 vdd.n1094 gnd 0.00249f
C3414 vdd.n1095 gnd 0.002637f
C3415 vdd.n1096 gnd 0.005886f
C3416 vdd.n1097 gnd 0.005886f
C3417 vdd.n1098 gnd 0.002637f
C3418 vdd.n1099 gnd 0.00249f
C3419 vdd.n1100 gnd 0.004634f
C3420 vdd.n1101 gnd 0.004634f
C3421 vdd.n1102 gnd 0.00249f
C3422 vdd.n1103 gnd 0.002637f
C3423 vdd.n1104 gnd 0.005886f
C3424 vdd.n1105 gnd 0.005886f
C3425 vdd.n1106 gnd 0.013915f
C3426 vdd.n1107 gnd 0.002563f
C3427 vdd.n1108 gnd 0.00249f
C3428 vdd.n1109 gnd 0.011977f
C3429 vdd.n1110 gnd 0.008362f
C3430 vdd.t137 gnd 0.029295f
C3431 vdd.t119 gnd 0.029295f
C3432 vdd.n1111 gnd 0.201332f
C3433 vdd.n1112 gnd 0.158317f
C3434 vdd.t13 gnd 0.029295f
C3435 vdd.t115 gnd 0.029295f
C3436 vdd.n1113 gnd 0.201332f
C3437 vdd.n1114 gnd 0.127761f
C3438 vdd.t144 gnd 0.029295f
C3439 vdd.t120 gnd 0.029295f
C3440 vdd.n1115 gnd 0.201332f
C3441 vdd.n1116 gnd 0.127761f
C3442 vdd.n1117 gnd 0.004994f
C3443 vdd.n1118 gnd 0.004634f
C3444 vdd.n1119 gnd 0.002563f
C3445 vdd.n1120 gnd 0.005886f
C3446 vdd.n1121 gnd 0.00249f
C3447 vdd.n1122 gnd 0.002637f
C3448 vdd.n1123 gnd 0.004634f
C3449 vdd.n1124 gnd 0.00249f
C3450 vdd.n1125 gnd 0.005886f
C3451 vdd.n1126 gnd 0.002637f
C3452 vdd.n1127 gnd 0.004634f
C3453 vdd.n1128 gnd 0.00249f
C3454 vdd.n1129 gnd 0.004414f
C3455 vdd.n1130 gnd 0.004427f
C3456 vdd.t102 gnd 0.012645f
C3457 vdd.n1131 gnd 0.028134f
C3458 vdd.n1132 gnd 0.146416f
C3459 vdd.n1133 gnd 0.00249f
C3460 vdd.n1134 gnd 0.002637f
C3461 vdd.n1135 gnd 0.005886f
C3462 vdd.n1136 gnd 0.005886f
C3463 vdd.n1137 gnd 0.002637f
C3464 vdd.n1138 gnd 0.00249f
C3465 vdd.n1139 gnd 0.004634f
C3466 vdd.n1140 gnd 0.004634f
C3467 vdd.n1141 gnd 0.00249f
C3468 vdd.n1142 gnd 0.002637f
C3469 vdd.n1143 gnd 0.005886f
C3470 vdd.n1144 gnd 0.005886f
C3471 vdd.n1145 gnd 0.002637f
C3472 vdd.n1146 gnd 0.00249f
C3473 vdd.n1147 gnd 0.004634f
C3474 vdd.n1148 gnd 0.004634f
C3475 vdd.n1149 gnd 0.00249f
C3476 vdd.n1150 gnd 0.002637f
C3477 vdd.n1151 gnd 0.005886f
C3478 vdd.n1152 gnd 0.005886f
C3479 vdd.n1153 gnd 0.013915f
C3480 vdd.n1154 gnd 0.002563f
C3481 vdd.n1155 gnd 0.00249f
C3482 vdd.n1156 gnd 0.011977f
C3483 vdd.n1157 gnd 0.008099f
C3484 vdd.n1158 gnd 0.056548f
C3485 vdd.n1159 gnd 0.220543f
C3486 vdd.n1160 gnd 1.8535f
C3487 vdd.n1161 gnd 0.536697f
C3488 vdd.n1162 gnd 0.007324f
C3489 vdd.n1163 gnd 0.009099f
C3490 vdd.n1164 gnd 0.571877f
C3491 vdd.n1165 gnd 0.009099f
C3492 vdd.n1166 gnd 0.007324f
C3493 vdd.n1167 gnd 0.009099f
C3494 vdd.n1168 gnd 0.007324f
C3495 vdd.n1169 gnd 0.009099f
C3496 vdd.t107 gnd 0.46494f
C3497 vdd.t12 gnd 0.46494f
C3498 vdd.n1170 gnd 0.009099f
C3499 vdd.n1171 gnd 0.007324f
C3500 vdd.n1172 gnd 0.009099f
C3501 vdd.n1173 gnd 0.007324f
C3502 vdd.n1174 gnd 0.009099f
C3503 vdd.t105 gnd 0.46494f
C3504 vdd.n1175 gnd 0.009099f
C3505 vdd.n1176 gnd 0.007324f
C3506 vdd.n1177 gnd 0.009099f
C3507 vdd.n1178 gnd 0.007324f
C3508 vdd.n1179 gnd 0.009099f
C3509 vdd.t101 gnd 0.46494f
C3510 vdd.n1180 gnd 0.674164f
C3511 vdd.n1181 gnd 0.009099f
C3512 vdd.n1182 gnd 0.007324f
C3513 vdd.n1183 gnd 0.009099f
C3514 vdd.n1184 gnd 0.007324f
C3515 vdd.n1185 gnd 0.009099f
C3516 vdd.n1186 gnd 0.929881f
C3517 vdd.n1187 gnd 0.009099f
C3518 vdd.n1188 gnd 0.007324f
C3519 vdd.n1189 gnd 0.022175f
C3520 vdd.n1190 gnd 0.006079f
C3521 vdd.n1191 gnd 0.022175f
C3522 vdd.t32 gnd 0.46494f
C3523 vdd.n1192 gnd 0.022175f
C3524 vdd.n1193 gnd 0.006079f
C3525 vdd.n1194 gnd 0.009099f
C3526 vdd.n1195 gnd 0.007324f
C3527 vdd.n1196 gnd 0.009099f
C3528 vdd.n1227 gnd 0.022684f
C3529 vdd.n1228 gnd 1.37157f
C3530 vdd.n1229 gnd 0.009099f
C3531 vdd.n1230 gnd 0.007324f
C3532 vdd.n1231 gnd 0.009099f
C3533 vdd.n1232 gnd 0.009099f
C3534 vdd.n1233 gnd 0.009099f
C3535 vdd.n1234 gnd 0.009099f
C3536 vdd.n1235 gnd 0.009099f
C3537 vdd.n1236 gnd 0.007324f
C3538 vdd.n1237 gnd 0.009099f
C3539 vdd.n1238 gnd 0.009099f
C3540 vdd.n1239 gnd 0.009099f
C3541 vdd.n1240 gnd 0.009099f
C3542 vdd.n1241 gnd 0.009099f
C3543 vdd.n1242 gnd 0.007324f
C3544 vdd.n1243 gnd 0.009099f
C3545 vdd.n1244 gnd 0.009099f
C3546 vdd.n1245 gnd 0.009099f
C3547 vdd.n1246 gnd 0.009099f
C3548 vdd.n1247 gnd 0.009099f
C3549 vdd.n1248 gnd 0.007324f
C3550 vdd.n1249 gnd 0.009099f
C3551 vdd.n1250 gnd 0.009099f
C3552 vdd.n1251 gnd 0.009099f
C3553 vdd.n1252 gnd 0.009099f
C3554 vdd.n1253 gnd 0.009099f
C3555 vdd.t81 gnd 0.111942f
C3556 vdd.t82 gnd 0.119636f
C3557 vdd.t80 gnd 0.146195f
C3558 vdd.n1254 gnd 0.187402f
C3559 vdd.n1255 gnd 0.158184f
C3560 vdd.n1256 gnd 0.015673f
C3561 vdd.n1257 gnd 0.009099f
C3562 vdd.n1258 gnd 0.009099f
C3563 vdd.n1259 gnd 0.009099f
C3564 vdd.n1260 gnd 0.009099f
C3565 vdd.n1261 gnd 0.009099f
C3566 vdd.n1262 gnd 0.007324f
C3567 vdd.n1263 gnd 0.009099f
C3568 vdd.n1264 gnd 0.009099f
C3569 vdd.n1265 gnd 0.009099f
C3570 vdd.n1266 gnd 0.009099f
C3571 vdd.n1267 gnd 0.009099f
C3572 vdd.n1268 gnd 0.007324f
C3573 vdd.n1269 gnd 0.009099f
C3574 vdd.n1270 gnd 0.009099f
C3575 vdd.n1271 gnd 0.009099f
C3576 vdd.n1272 gnd 0.009099f
C3577 vdd.n1273 gnd 0.009099f
C3578 vdd.n1274 gnd 0.007324f
C3579 vdd.n1275 gnd 0.009099f
C3580 vdd.n1276 gnd 0.009099f
C3581 vdd.n1277 gnd 0.009099f
C3582 vdd.n1278 gnd 0.009099f
C3583 vdd.n1279 gnd 0.009099f
C3584 vdd.n1280 gnd 0.007324f
C3585 vdd.n1281 gnd 0.009099f
C3586 vdd.n1282 gnd 0.009099f
C3587 vdd.n1283 gnd 0.009099f
C3588 vdd.n1284 gnd 0.009099f
C3589 vdd.n1285 gnd 0.009099f
C3590 vdd.n1286 gnd 0.007324f
C3591 vdd.n1287 gnd 0.009099f
C3592 vdd.n1288 gnd 0.009099f
C3593 vdd.n1289 gnd 0.009099f
C3594 vdd.n1290 gnd 0.009099f
C3595 vdd.n1291 gnd 0.007324f
C3596 vdd.n1292 gnd 0.009099f
C3597 vdd.n1293 gnd 0.009099f
C3598 vdd.n1294 gnd 0.009099f
C3599 vdd.n1295 gnd 0.009099f
C3600 vdd.n1296 gnd 0.009099f
C3601 vdd.n1297 gnd 0.007324f
C3602 vdd.n1298 gnd 0.009099f
C3603 vdd.n1299 gnd 0.009099f
C3604 vdd.n1300 gnd 0.009099f
C3605 vdd.n1301 gnd 0.009099f
C3606 vdd.n1302 gnd 0.009099f
C3607 vdd.n1303 gnd 0.007324f
C3608 vdd.n1304 gnd 0.009099f
C3609 vdd.n1305 gnd 0.009099f
C3610 vdd.n1306 gnd 0.009099f
C3611 vdd.n1307 gnd 0.009099f
C3612 vdd.n1308 gnd 0.009099f
C3613 vdd.n1309 gnd 0.007324f
C3614 vdd.n1310 gnd 0.009099f
C3615 vdd.n1311 gnd 0.009099f
C3616 vdd.n1312 gnd 0.009099f
C3617 vdd.n1313 gnd 0.009099f
C3618 vdd.n1314 gnd 0.009099f
C3619 vdd.n1315 gnd 0.007324f
C3620 vdd.n1316 gnd 0.009099f
C3621 vdd.n1317 gnd 0.009099f
C3622 vdd.n1318 gnd 0.009099f
C3623 vdd.n1319 gnd 0.009099f
C3624 vdd.t33 gnd 0.111942f
C3625 vdd.t34 gnd 0.119636f
C3626 vdd.t31 gnd 0.146195f
C3627 vdd.n1320 gnd 0.187402f
C3628 vdd.n1321 gnd 0.158184f
C3629 vdd.n1322 gnd 0.012011f
C3630 vdd.n1323 gnd 0.003479f
C3631 vdd.n1324 gnd 0.022684f
C3632 vdd.n1325 gnd 0.009099f
C3633 vdd.n1326 gnd 0.003845f
C3634 vdd.n1327 gnd 0.007324f
C3635 vdd.n1328 gnd 0.007324f
C3636 vdd.n1329 gnd 0.009099f
C3637 vdd.n1330 gnd 0.009099f
C3638 vdd.n1331 gnd 0.009099f
C3639 vdd.n1332 gnd 0.007324f
C3640 vdd.n1333 gnd 0.007324f
C3641 vdd.n1334 gnd 0.007324f
C3642 vdd.n1335 gnd 0.009099f
C3643 vdd.n1336 gnd 0.009099f
C3644 vdd.n1337 gnd 0.009099f
C3645 vdd.n1338 gnd 0.007324f
C3646 vdd.n1339 gnd 0.007324f
C3647 vdd.n1340 gnd 0.007324f
C3648 vdd.n1341 gnd 0.009099f
C3649 vdd.n1342 gnd 0.009099f
C3650 vdd.n1343 gnd 0.009099f
C3651 vdd.n1344 gnd 0.007324f
C3652 vdd.n1345 gnd 0.007324f
C3653 vdd.n1346 gnd 0.007324f
C3654 vdd.n1347 gnd 0.009099f
C3655 vdd.n1348 gnd 0.009099f
C3656 vdd.n1349 gnd 0.009099f
C3657 vdd.n1350 gnd 0.007324f
C3658 vdd.n1351 gnd 0.007324f
C3659 vdd.n1352 gnd 0.007324f
C3660 vdd.n1353 gnd 0.009099f
C3661 vdd.n1354 gnd 0.009099f
C3662 vdd.n1355 gnd 0.009099f
C3663 vdd.n1356 gnd 0.00725f
C3664 vdd.n1357 gnd 0.009099f
C3665 vdd.t78 gnd 0.111942f
C3666 vdd.t79 gnd 0.119636f
C3667 vdd.t77 gnd 0.146195f
C3668 vdd.n1358 gnd 0.187402f
C3669 vdd.n1359 gnd 0.158184f
C3670 vdd.n1360 gnd 0.015673f
C3671 vdd.n1361 gnd 0.00498f
C3672 vdd.n1362 gnd 0.009099f
C3673 vdd.n1363 gnd 0.009099f
C3674 vdd.n1364 gnd 0.009099f
C3675 vdd.n1365 gnd 0.007324f
C3676 vdd.n1366 gnd 0.007324f
C3677 vdd.n1367 gnd 0.007324f
C3678 vdd.n1368 gnd 0.009099f
C3679 vdd.n1369 gnd 0.009099f
C3680 vdd.n1370 gnd 0.009099f
C3681 vdd.n1371 gnd 0.007324f
C3682 vdd.n1372 gnd 0.007324f
C3683 vdd.n1373 gnd 0.007324f
C3684 vdd.n1374 gnd 0.009099f
C3685 vdd.n1375 gnd 0.009099f
C3686 vdd.n1376 gnd 0.009099f
C3687 vdd.n1377 gnd 0.007324f
C3688 vdd.n1378 gnd 0.007324f
C3689 vdd.n1379 gnd 0.007324f
C3690 vdd.n1380 gnd 0.009099f
C3691 vdd.n1381 gnd 0.009099f
C3692 vdd.n1382 gnd 0.009099f
C3693 vdd.n1383 gnd 0.007324f
C3694 vdd.n1384 gnd 0.007324f
C3695 vdd.n1385 gnd 0.007324f
C3696 vdd.n1386 gnd 0.009099f
C3697 vdd.n1387 gnd 0.009099f
C3698 vdd.n1388 gnd 0.009099f
C3699 vdd.n1389 gnd 0.007324f
C3700 vdd.n1390 gnd 0.007324f
C3701 vdd.n1391 gnd 0.006115f
C3702 vdd.n1392 gnd 0.009099f
C3703 vdd.n1393 gnd 0.009099f
C3704 vdd.n1394 gnd 0.009099f
C3705 vdd.n1395 gnd 0.006115f
C3706 vdd.n1396 gnd 0.007324f
C3707 vdd.n1397 gnd 0.007324f
C3708 vdd.n1398 gnd 0.009099f
C3709 vdd.n1399 gnd 0.009099f
C3710 vdd.n1400 gnd 0.009099f
C3711 vdd.n1401 gnd 0.007324f
C3712 vdd.n1402 gnd 0.007324f
C3713 vdd.n1403 gnd 0.007324f
C3714 vdd.n1404 gnd 0.009099f
C3715 vdd.n1405 gnd 0.009099f
C3716 vdd.n1406 gnd 0.009099f
C3717 vdd.n1407 gnd 0.007324f
C3718 vdd.n1408 gnd 0.007324f
C3719 vdd.n1409 gnd 0.007324f
C3720 vdd.n1410 gnd 0.009099f
C3721 vdd.n1411 gnd 0.009099f
C3722 vdd.n1412 gnd 0.009099f
C3723 vdd.n1413 gnd 0.007324f
C3724 vdd.n1414 gnd 0.007324f
C3725 vdd.n1415 gnd 0.007324f
C3726 vdd.n1416 gnd 0.009099f
C3727 vdd.n1417 gnd 0.009099f
C3728 vdd.n1418 gnd 0.009099f
C3729 vdd.n1419 gnd 0.007324f
C3730 vdd.n1420 gnd 0.009099f
C3731 vdd.n1421 gnd 2.22242f
C3732 vdd.n1423 gnd 0.022684f
C3733 vdd.n1424 gnd 0.006079f
C3734 vdd.n1425 gnd 0.022684f
C3735 vdd.n1426 gnd 0.022175f
C3736 vdd.n1427 gnd 0.009099f
C3737 vdd.n1428 gnd 0.007324f
C3738 vdd.n1429 gnd 0.009099f
C3739 vdd.n1430 gnd 0.488187f
C3740 vdd.n1431 gnd 0.009099f
C3741 vdd.n1432 gnd 0.007324f
C3742 vdd.n1433 gnd 0.009099f
C3743 vdd.n1434 gnd 0.009099f
C3744 vdd.n1435 gnd 0.009099f
C3745 vdd.n1436 gnd 0.007324f
C3746 vdd.n1437 gnd 0.009099f
C3747 vdd.n1438 gnd 0.832243f
C3748 vdd.n1439 gnd 0.929881f
C3749 vdd.n1440 gnd 0.009099f
C3750 vdd.n1441 gnd 0.007324f
C3751 vdd.n1442 gnd 0.009099f
C3752 vdd.n1443 gnd 0.009099f
C3753 vdd.n1444 gnd 0.009099f
C3754 vdd.n1445 gnd 0.007324f
C3755 vdd.n1446 gnd 0.009099f
C3756 vdd.n1447 gnd 0.562578f
C3757 vdd.n1448 gnd 0.009099f
C3758 vdd.n1449 gnd 0.007324f
C3759 vdd.n1450 gnd 0.009099f
C3760 vdd.n1451 gnd 0.009099f
C3761 vdd.n1452 gnd 0.009099f
C3762 vdd.n1453 gnd 0.007324f
C3763 vdd.n1454 gnd 0.009099f
C3764 vdd.n1455 gnd 0.516084f
C3765 vdd.n1456 gnd 0.720658f
C3766 vdd.n1457 gnd 0.009099f
C3767 vdd.n1458 gnd 0.007324f
C3768 vdd.n1459 gnd 0.009099f
C3769 vdd.n1460 gnd 0.009099f
C3770 vdd.n1461 gnd 0.006993f
C3771 vdd.n1462 gnd 0.009099f
C3772 vdd.n1463 gnd 0.007324f
C3773 vdd.n1464 gnd 0.009099f
C3774 vdd.n1465 gnd 0.771801f
C3775 vdd.n1466 gnd 0.009099f
C3776 vdd.n1467 gnd 0.007324f
C3777 vdd.n1468 gnd 0.009099f
C3778 vdd.n1469 gnd 0.009099f
C3779 vdd.n1470 gnd 0.009099f
C3780 vdd.n1471 gnd 0.007324f
C3781 vdd.n1472 gnd 0.009099f
C3782 vdd.t10 gnd 0.46494f
C3783 vdd.n1473 gnd 0.664865f
C3784 vdd.n1474 gnd 0.009099f
C3785 vdd.n1475 gnd 0.007324f
C3786 vdd.n1476 gnd 0.006993f
C3787 vdd.n1477 gnd 0.009099f
C3788 vdd.n1478 gnd 0.009099f
C3789 vdd.n1479 gnd 0.007324f
C3790 vdd.n1480 gnd 0.009099f
C3791 vdd.n1481 gnd 0.506785f
C3792 vdd.n1482 gnd 0.009099f
C3793 vdd.n1483 gnd 0.007324f
C3794 vdd.n1484 gnd 0.009099f
C3795 vdd.n1485 gnd 0.009099f
C3796 vdd.n1486 gnd 0.009099f
C3797 vdd.n1487 gnd 0.007324f
C3798 vdd.n1488 gnd 0.009099f
C3799 vdd.n1489 gnd 0.655566f
C3800 vdd.n1490 gnd 0.581176f
C3801 vdd.n1491 gnd 0.009099f
C3802 vdd.n1492 gnd 0.007324f
C3803 vdd.n1493 gnd 0.009099f
C3804 vdd.n1494 gnd 0.009099f
C3805 vdd.n1495 gnd 0.009099f
C3806 vdd.n1496 gnd 0.007324f
C3807 vdd.n1497 gnd 0.009099f
C3808 vdd.n1498 gnd 0.739255f
C3809 vdd.n1499 gnd 0.009099f
C3810 vdd.n1500 gnd 0.007324f
C3811 vdd.n1501 gnd 0.009099f
C3812 vdd.n1502 gnd 0.009099f
C3813 vdd.n1503 gnd 0.022175f
C3814 vdd.n1504 gnd 0.009099f
C3815 vdd.n1505 gnd 0.009099f
C3816 vdd.n1506 gnd 0.007324f
C3817 vdd.n1507 gnd 0.009099f
C3818 vdd.n1508 gnd 0.581176f
C3819 vdd.n1509 gnd 0.929881f
C3820 vdd.n1510 gnd 0.009099f
C3821 vdd.n1511 gnd 0.007324f
C3822 vdd.n1512 gnd 0.009099f
C3823 vdd.n1513 gnd 0.009099f
C3824 vdd.n1514 gnd 0.007825f
C3825 vdd.n1515 gnd 0.007324f
C3826 vdd.n1517 gnd 0.009099f
C3827 vdd.n1519 gnd 0.007324f
C3828 vdd.n1520 gnd 0.009099f
C3829 vdd.n1521 gnd 0.007324f
C3830 vdd.n1523 gnd 0.009099f
C3831 vdd.n1524 gnd 0.007324f
C3832 vdd.n1525 gnd 0.009099f
C3833 vdd.n1526 gnd 0.009099f
C3834 vdd.n1527 gnd 0.009099f
C3835 vdd.n1528 gnd 0.009099f
C3836 vdd.n1529 gnd 0.009099f
C3837 vdd.n1530 gnd 0.007324f
C3838 vdd.n1532 gnd 0.009099f
C3839 vdd.n1533 gnd 0.009099f
C3840 vdd.n1534 gnd 0.009099f
C3841 vdd.n1535 gnd 0.009099f
C3842 vdd.n1536 gnd 0.009099f
C3843 vdd.n1537 gnd 0.007324f
C3844 vdd.n1539 gnd 0.009099f
C3845 vdd.n1540 gnd 0.009099f
C3846 vdd.n1541 gnd 0.009099f
C3847 vdd.n1542 gnd 0.009099f
C3848 vdd.n1543 gnd 0.006115f
C3849 vdd.t48 gnd 0.111942f
C3850 vdd.t47 gnd 0.119636f
C3851 vdd.t46 gnd 0.146195f
C3852 vdd.n1544 gnd 0.187402f
C3853 vdd.n1545 gnd 0.157451f
C3854 vdd.n1547 gnd 0.009099f
C3855 vdd.n1548 gnd 0.009099f
C3856 vdd.n1549 gnd 0.007324f
C3857 vdd.n1550 gnd 0.009099f
C3858 vdd.n1552 gnd 0.009099f
C3859 vdd.n1553 gnd 0.009099f
C3860 vdd.n1554 gnd 0.009099f
C3861 vdd.n1555 gnd 0.009099f
C3862 vdd.n1556 gnd 0.007324f
C3863 vdd.n1558 gnd 0.009099f
C3864 vdd.n1559 gnd 0.009099f
C3865 vdd.n1560 gnd 0.009099f
C3866 vdd.n1561 gnd 0.009099f
C3867 vdd.n1562 gnd 0.009099f
C3868 vdd.n1563 gnd 0.007324f
C3869 vdd.n1565 gnd 0.009099f
C3870 vdd.n1566 gnd 0.009099f
C3871 vdd.n1567 gnd 0.009099f
C3872 vdd.n1568 gnd 0.009099f
C3873 vdd.n1569 gnd 0.009099f
C3874 vdd.n1570 gnd 0.007324f
C3875 vdd.n1572 gnd 0.009099f
C3876 vdd.n1573 gnd 0.009099f
C3877 vdd.n1574 gnd 0.009099f
C3878 vdd.n1575 gnd 0.009099f
C3879 vdd.n1576 gnd 0.009099f
C3880 vdd.n1577 gnd 0.007324f
C3881 vdd.n1579 gnd 0.009099f
C3882 vdd.n1580 gnd 0.009099f
C3883 vdd.n1581 gnd 0.009099f
C3884 vdd.n1582 gnd 0.009099f
C3885 vdd.n1583 gnd 0.00725f
C3886 vdd.t41 gnd 0.111942f
C3887 vdd.t40 gnd 0.119636f
C3888 vdd.t39 gnd 0.146195f
C3889 vdd.n1584 gnd 0.187402f
C3890 vdd.n1585 gnd 0.157451f
C3891 vdd.n1587 gnd 0.009099f
C3892 vdd.n1588 gnd 0.009099f
C3893 vdd.n1589 gnd 0.007324f
C3894 vdd.n1590 gnd 0.009099f
C3895 vdd.n1592 gnd 0.009099f
C3896 vdd.n1593 gnd 0.009099f
C3897 vdd.n1594 gnd 0.009099f
C3898 vdd.n1595 gnd 0.009099f
C3899 vdd.n1596 gnd 0.007324f
C3900 vdd.n1598 gnd 0.009099f
C3901 vdd.n1599 gnd 0.009099f
C3902 vdd.n1600 gnd 0.009099f
C3903 vdd.n1601 gnd 0.009099f
C3904 vdd.n1602 gnd 0.009099f
C3905 vdd.n1603 gnd 0.007324f
C3906 vdd.n1605 gnd 0.009099f
C3907 vdd.n1606 gnd 0.009099f
C3908 vdd.n1607 gnd 0.009099f
C3909 vdd.n1608 gnd 0.009099f
C3910 vdd.n1609 gnd 0.009099f
C3911 vdd.n1610 gnd 0.009099f
C3912 vdd.n1611 gnd 0.007324f
C3913 vdd.n1613 gnd 0.009099f
C3914 vdd.n1615 gnd 0.009099f
C3915 vdd.n1616 gnd 0.007324f
C3916 vdd.n1617 gnd 0.007324f
C3917 vdd.n1618 gnd 0.009099f
C3918 vdd.n1620 gnd 0.009099f
C3919 vdd.n1621 gnd 0.007324f
C3920 vdd.n1622 gnd 0.007324f
C3921 vdd.n1623 gnd 0.009099f
C3922 vdd.n1625 gnd 0.009099f
C3923 vdd.n1626 gnd 0.009099f
C3924 vdd.n1627 gnd 0.007324f
C3925 vdd.n1628 gnd 0.007324f
C3926 vdd.n1629 gnd 0.007324f
C3927 vdd.n1630 gnd 0.009099f
C3928 vdd.n1632 gnd 0.009099f
C3929 vdd.n1633 gnd 0.009099f
C3930 vdd.n1634 gnd 0.007324f
C3931 vdd.n1635 gnd 0.007324f
C3932 vdd.n1636 gnd 0.007324f
C3933 vdd.n1637 gnd 0.009099f
C3934 vdd.n1639 gnd 0.009099f
C3935 vdd.n1640 gnd 0.009099f
C3936 vdd.n1641 gnd 0.007324f
C3937 vdd.n1642 gnd 0.007324f
C3938 vdd.n1643 gnd 0.007324f
C3939 vdd.n1644 gnd 0.009099f
C3940 vdd.n1646 gnd 0.009099f
C3941 vdd.n1647 gnd 0.009099f
C3942 vdd.n1648 gnd 0.007324f
C3943 vdd.n1649 gnd 0.009099f
C3944 vdd.n1650 gnd 0.009099f
C3945 vdd.n1651 gnd 0.009099f
C3946 vdd.n1652 gnd 0.01494f
C3947 vdd.n1653 gnd 0.00498f
C3948 vdd.n1654 gnd 0.007324f
C3949 vdd.n1655 gnd 0.009099f
C3950 vdd.n1657 gnd 0.009099f
C3951 vdd.n1658 gnd 0.009099f
C3952 vdd.n1659 gnd 0.007324f
C3953 vdd.n1660 gnd 0.007324f
C3954 vdd.n1661 gnd 0.007324f
C3955 vdd.n1662 gnd 0.009099f
C3956 vdd.n1664 gnd 0.009099f
C3957 vdd.n1665 gnd 0.009099f
C3958 vdd.n1666 gnd 0.007324f
C3959 vdd.n1667 gnd 0.007324f
C3960 vdd.n1668 gnd 0.007324f
C3961 vdd.n1669 gnd 0.009099f
C3962 vdd.n1671 gnd 0.009099f
C3963 vdd.n1672 gnd 0.009099f
C3964 vdd.n1673 gnd 0.007324f
C3965 vdd.n1674 gnd 0.007324f
C3966 vdd.n1675 gnd 0.007324f
C3967 vdd.n1676 gnd 0.009099f
C3968 vdd.n1678 gnd 0.009099f
C3969 vdd.n1679 gnd 0.009099f
C3970 vdd.n1680 gnd 0.007324f
C3971 vdd.n1681 gnd 0.007324f
C3972 vdd.n1682 gnd 0.007324f
C3973 vdd.n1683 gnd 0.009099f
C3974 vdd.n1685 gnd 0.009099f
C3975 vdd.n1686 gnd 0.009099f
C3976 vdd.n1687 gnd 0.007324f
C3977 vdd.n1688 gnd 0.009099f
C3978 vdd.n1689 gnd 0.009099f
C3979 vdd.n1690 gnd 0.009099f
C3980 vdd.n1691 gnd 0.01494f
C3981 vdd.n1692 gnd 0.006115f
C3982 vdd.n1693 gnd 0.007324f
C3983 vdd.n1694 gnd 0.009099f
C3984 vdd.n1696 gnd 0.009099f
C3985 vdd.n1697 gnd 0.009099f
C3986 vdd.n1698 gnd 0.007324f
C3987 vdd.n1699 gnd 0.007324f
C3988 vdd.n1700 gnd 0.007324f
C3989 vdd.n1701 gnd 0.009099f
C3990 vdd.n1703 gnd 0.009099f
C3991 vdd.n1704 gnd 0.009099f
C3992 vdd.n1705 gnd 0.007324f
C3993 vdd.n1706 gnd 0.007324f
C3994 vdd.n1707 gnd 0.007324f
C3995 vdd.n1708 gnd 0.009099f
C3996 vdd.n1710 gnd 0.009099f
C3997 vdd.n1711 gnd 0.009099f
C3998 vdd.n1713 gnd 0.009099f
C3999 vdd.n1714 gnd 0.007324f
C4000 vdd.n1715 gnd 0.005823f
C4001 vdd.n1716 gnd 0.006187f
C4002 vdd.n1717 gnd 0.006187f
C4003 vdd.n1718 gnd 0.006187f
C4004 vdd.n1719 gnd 0.006187f
C4005 vdd.n1720 gnd 0.006187f
C4006 vdd.n1721 gnd 0.006187f
C4007 vdd.n1722 gnd 0.006187f
C4008 vdd.n1723 gnd 0.006187f
C4009 vdd.n1725 gnd 0.006187f
C4010 vdd.n1726 gnd 0.006187f
C4011 vdd.n1727 gnd 0.006187f
C4012 vdd.n1728 gnd 0.006187f
C4013 vdd.n1729 gnd 0.006187f
C4014 vdd.n1731 gnd 0.006187f
C4015 vdd.n1733 gnd 0.006187f
C4016 vdd.n1734 gnd 0.006187f
C4017 vdd.n1735 gnd 0.006187f
C4018 vdd.n1736 gnd 0.006187f
C4019 vdd.n1737 gnd 0.006187f
C4020 vdd.n1739 gnd 0.006187f
C4021 vdd.n1741 gnd 0.006187f
C4022 vdd.n1742 gnd 0.006187f
C4023 vdd.n1743 gnd 0.006187f
C4024 vdd.n1744 gnd 0.006187f
C4025 vdd.n1745 gnd 0.006187f
C4026 vdd.n1747 gnd 0.006187f
C4027 vdd.n1749 gnd 0.006187f
C4028 vdd.n1750 gnd 0.006187f
C4029 vdd.n1751 gnd 0.006187f
C4030 vdd.n1752 gnd 0.006187f
C4031 vdd.n1753 gnd 0.006187f
C4032 vdd.n1755 gnd 0.006187f
C4033 vdd.n1756 gnd 0.006187f
C4034 vdd.n1757 gnd 0.006187f
C4035 vdd.n1758 gnd 0.006187f
C4036 vdd.n1759 gnd 0.006187f
C4037 vdd.n1760 gnd 0.006187f
C4038 vdd.n1761 gnd 0.006187f
C4039 vdd.n1762 gnd 0.006187f
C4040 vdd.n1763 gnd 0.004504f
C4041 vdd.n1764 gnd 0.006187f
C4042 vdd.t18 gnd 0.25003f
C4043 vdd.t19 gnd 0.255937f
C4044 vdd.t16 gnd 0.163229f
C4045 vdd.n1765 gnd 0.088216f
C4046 vdd.n1766 gnd 0.050039f
C4047 vdd.n1767 gnd 0.008843f
C4048 vdd.n1768 gnd 0.006187f
C4049 vdd.n1769 gnd 0.006187f
C4050 vdd.n1770 gnd 0.376602f
C4051 vdd.n1771 gnd 0.006187f
C4052 vdd.n1772 gnd 0.006187f
C4053 vdd.n1773 gnd 0.006187f
C4054 vdd.n1774 gnd 0.006187f
C4055 vdd.n1775 gnd 0.006187f
C4056 vdd.n1776 gnd 0.006187f
C4057 vdd.n1777 gnd 0.006187f
C4058 vdd.n1778 gnd 0.006187f
C4059 vdd.n1779 gnd 0.006187f
C4060 vdd.n1780 gnd 0.006187f
C4061 vdd.n1781 gnd 0.006187f
C4062 vdd.n1782 gnd 0.006187f
C4063 vdd.n1783 gnd 0.006187f
C4064 vdd.n1784 gnd 0.006187f
C4065 vdd.n1785 gnd 0.006187f
C4066 vdd.n1786 gnd 0.006187f
C4067 vdd.n1787 gnd 0.006187f
C4068 vdd.n1788 gnd 0.006187f
C4069 vdd.n1789 gnd 0.006187f
C4070 vdd.n1790 gnd 0.006187f
C4071 vdd.t65 gnd 0.25003f
C4072 vdd.t66 gnd 0.255937f
C4073 vdd.t64 gnd 0.163229f
C4074 vdd.n1791 gnd 0.088216f
C4075 vdd.n1792 gnd 0.050039f
C4076 vdd.n1793 gnd 0.006187f
C4077 vdd.n1794 gnd 0.006187f
C4078 vdd.n1795 gnd 0.006187f
C4079 vdd.n1796 gnd 0.006187f
C4080 vdd.n1797 gnd 0.006187f
C4081 vdd.n1798 gnd 0.006187f
C4082 vdd.n1800 gnd 0.006187f
C4083 vdd.n1801 gnd 0.006187f
C4084 vdd.n1802 gnd 0.006187f
C4085 vdd.n1803 gnd 0.006187f
C4086 vdd.n1805 gnd 0.006187f
C4087 vdd.n1807 gnd 0.006187f
C4088 vdd.n1808 gnd 0.006187f
C4089 vdd.n1809 gnd 0.006187f
C4090 vdd.n1810 gnd 0.006187f
C4091 vdd.n1811 gnd 0.006187f
C4092 vdd.n1813 gnd 0.006187f
C4093 vdd.n1815 gnd 0.006187f
C4094 vdd.n1816 gnd 0.006187f
C4095 vdd.n1817 gnd 0.006187f
C4096 vdd.n1818 gnd 0.006187f
C4097 vdd.n1819 gnd 0.006187f
C4098 vdd.n1821 gnd 0.006187f
C4099 vdd.n1823 gnd 0.006187f
C4100 vdd.n1824 gnd 0.006187f
C4101 vdd.n1825 gnd 0.004504f
C4102 vdd.n1826 gnd 0.008843f
C4103 vdd.n1827 gnd 0.004777f
C4104 vdd.n1828 gnd 0.006187f
C4105 vdd.n1830 gnd 0.006187f
C4106 vdd.n1831 gnd 0.014682f
C4107 vdd.n1832 gnd 0.014682f
C4108 vdd.n1833 gnd 0.013708f
C4109 vdd.n1834 gnd 0.006187f
C4110 vdd.n1835 gnd 0.006187f
C4111 vdd.n1836 gnd 0.006187f
C4112 vdd.n1837 gnd 0.006187f
C4113 vdd.n1838 gnd 0.006187f
C4114 vdd.n1839 gnd 0.006187f
C4115 vdd.n1840 gnd 0.006187f
C4116 vdd.n1841 gnd 0.006187f
C4117 vdd.n1842 gnd 0.006187f
C4118 vdd.n1843 gnd 0.006187f
C4119 vdd.n1844 gnd 0.006187f
C4120 vdd.n1845 gnd 0.006187f
C4121 vdd.n1846 gnd 0.006187f
C4122 vdd.n1847 gnd 0.006187f
C4123 vdd.n1848 gnd 0.006187f
C4124 vdd.n1849 gnd 0.006187f
C4125 vdd.n1850 gnd 0.006187f
C4126 vdd.n1851 gnd 0.006187f
C4127 vdd.n1852 gnd 0.006187f
C4128 vdd.n1853 gnd 0.006187f
C4129 vdd.n1854 gnd 0.006187f
C4130 vdd.n1855 gnd 0.006187f
C4131 vdd.n1856 gnd 0.006187f
C4132 vdd.n1857 gnd 0.006187f
C4133 vdd.n1858 gnd 0.006187f
C4134 vdd.n1859 gnd 0.006187f
C4135 vdd.n1860 gnd 0.006187f
C4136 vdd.n1861 gnd 0.006187f
C4137 vdd.n1862 gnd 0.006187f
C4138 vdd.n1863 gnd 0.006187f
C4139 vdd.n1864 gnd 0.006187f
C4140 vdd.n1865 gnd 0.006187f
C4141 vdd.n1866 gnd 0.006187f
C4142 vdd.n1867 gnd 0.006187f
C4143 vdd.n1868 gnd 0.006187f
C4144 vdd.n1869 gnd 0.006187f
C4145 vdd.n1870 gnd 0.006187f
C4146 vdd.n1871 gnd 0.199924f
C4147 vdd.n1872 gnd 0.006187f
C4148 vdd.n1873 gnd 0.006187f
C4149 vdd.n1874 gnd 0.006187f
C4150 vdd.n1875 gnd 0.006187f
C4151 vdd.n1876 gnd 0.006187f
C4152 vdd.n1877 gnd 0.006187f
C4153 vdd.n1878 gnd 0.006187f
C4154 vdd.n1879 gnd 0.006187f
C4155 vdd.n1880 gnd 0.006187f
C4156 vdd.n1881 gnd 0.006187f
C4157 vdd.n1882 gnd 0.006187f
C4158 vdd.n1883 gnd 0.006187f
C4159 vdd.n1884 gnd 0.006187f
C4160 vdd.n1885 gnd 0.006187f
C4161 vdd.n1886 gnd 0.006187f
C4162 vdd.n1887 gnd 0.006187f
C4163 vdd.n1888 gnd 0.006187f
C4164 vdd.n1889 gnd 0.006187f
C4165 vdd.n1890 gnd 0.006187f
C4166 vdd.n1891 gnd 0.006187f
C4167 vdd.n1892 gnd 0.013708f
C4168 vdd.n1894 gnd 0.014682f
C4169 vdd.n1895 gnd 0.014682f
C4170 vdd.n1896 gnd 0.006187f
C4171 vdd.n1897 gnd 0.004777f
C4172 vdd.n1898 gnd 0.006187f
C4173 vdd.n1900 gnd 0.006187f
C4174 vdd.n1902 gnd 0.006187f
C4175 vdd.n1903 gnd 0.006187f
C4176 vdd.n1904 gnd 0.006187f
C4177 vdd.n1905 gnd 0.006187f
C4178 vdd.n1906 gnd 0.006187f
C4179 vdd.n1908 gnd 0.006187f
C4180 vdd.n1910 gnd 0.006187f
C4181 vdd.n1911 gnd 0.006187f
C4182 vdd.n1912 gnd 0.006187f
C4183 vdd.n1913 gnd 0.006187f
C4184 vdd.n1914 gnd 0.006187f
C4185 vdd.n1916 gnd 0.006187f
C4186 vdd.n1918 gnd 0.006187f
C4187 vdd.n1919 gnd 0.006187f
C4188 vdd.n1920 gnd 0.006187f
C4189 vdd.n1921 gnd 0.006187f
C4190 vdd.n1922 gnd 0.006187f
C4191 vdd.n1924 gnd 0.006187f
C4192 vdd.n1926 gnd 0.006187f
C4193 vdd.n1927 gnd 0.006187f
C4194 vdd.n1928 gnd 0.018456f
C4195 vdd.n1929 gnd 0.547103f
C4196 vdd.n1931 gnd 0.007324f
C4197 vdd.n1932 gnd 0.007324f
C4198 vdd.n1933 gnd 0.009099f
C4199 vdd.n1935 gnd 0.009099f
C4200 vdd.n1936 gnd 0.009099f
C4201 vdd.n1937 gnd 0.007324f
C4202 vdd.n1938 gnd 0.006079f
C4203 vdd.n1939 gnd 0.022684f
C4204 vdd.n1940 gnd 0.022175f
C4205 vdd.n1941 gnd 0.006079f
C4206 vdd.n1942 gnd 0.022175f
C4207 vdd.n1943 gnd 1.27859f
C4208 vdd.n1944 gnd 0.022175f
C4209 vdd.n1945 gnd 0.022684f
C4210 vdd.n1946 gnd 0.003479f
C4211 vdd.t30 gnd 0.111942f
C4212 vdd.t29 gnd 0.119636f
C4213 vdd.t27 gnd 0.146195f
C4214 vdd.n1947 gnd 0.187402f
C4215 vdd.n1948 gnd 0.157451f
C4216 vdd.n1949 gnd 0.011278f
C4217 vdd.n1950 gnd 0.003845f
C4218 vdd.n1951 gnd 0.007825f
C4219 vdd.n1952 gnd 0.547103f
C4220 vdd.n1953 gnd 0.018456f
C4221 vdd.n1954 gnd 0.006187f
C4222 vdd.n1955 gnd 0.006187f
C4223 vdd.n1956 gnd 0.006187f
C4224 vdd.n1958 gnd 0.006187f
C4225 vdd.n1960 gnd 0.006187f
C4226 vdd.n1961 gnd 0.006187f
C4227 vdd.n1962 gnd 0.006187f
C4228 vdd.n1963 gnd 0.006187f
C4229 vdd.n1964 gnd 0.006187f
C4230 vdd.n1966 gnd 0.006187f
C4231 vdd.n1968 gnd 0.006187f
C4232 vdd.n1969 gnd 0.006187f
C4233 vdd.n1970 gnd 0.006187f
C4234 vdd.n1971 gnd 0.006187f
C4235 vdd.n1972 gnd 0.006187f
C4236 vdd.n1974 gnd 0.006187f
C4237 vdd.n1976 gnd 0.006187f
C4238 vdd.n1977 gnd 0.006187f
C4239 vdd.n1978 gnd 0.006187f
C4240 vdd.n1979 gnd 0.006187f
C4241 vdd.n1980 gnd 0.006187f
C4242 vdd.n1982 gnd 0.006187f
C4243 vdd.n1984 gnd 0.006187f
C4244 vdd.n1985 gnd 0.006187f
C4245 vdd.n1986 gnd 0.014682f
C4246 vdd.n1987 gnd 0.013708f
C4247 vdd.n1988 gnd 0.013708f
C4248 vdd.n1989 gnd 0.911283f
C4249 vdd.n1990 gnd 0.013708f
C4250 vdd.n1991 gnd 0.013708f
C4251 vdd.n1992 gnd 0.006187f
C4252 vdd.n1993 gnd 0.006187f
C4253 vdd.n1994 gnd 0.006187f
C4254 vdd.n1995 gnd 0.395199f
C4255 vdd.n1996 gnd 0.006187f
C4256 vdd.n1997 gnd 0.006187f
C4257 vdd.n1998 gnd 0.006187f
C4258 vdd.n1999 gnd 0.006187f
C4259 vdd.n2000 gnd 0.006187f
C4260 vdd.n2001 gnd 0.632319f
C4261 vdd.n2002 gnd 0.006187f
C4262 vdd.n2003 gnd 0.006187f
C4263 vdd.n2004 gnd 0.006187f
C4264 vdd.n2005 gnd 0.006187f
C4265 vdd.n2006 gnd 0.006187f
C4266 vdd.n2007 gnd 0.632319f
C4267 vdd.n2008 gnd 0.006187f
C4268 vdd.n2009 gnd 0.006187f
C4269 vdd.n2010 gnd 0.005459f
C4270 vdd.n2011 gnd 0.017924f
C4271 vdd.n2012 gnd 0.003822f
C4272 vdd.n2013 gnd 0.006187f
C4273 vdd.n2014 gnd 0.348705f
C4274 vdd.n2015 gnd 0.006187f
C4275 vdd.n2016 gnd 0.006187f
C4276 vdd.n2017 gnd 0.006187f
C4277 vdd.n2018 gnd 0.006187f
C4278 vdd.n2019 gnd 0.006187f
C4279 vdd.n2020 gnd 0.423096f
C4280 vdd.n2021 gnd 0.006187f
C4281 vdd.n2022 gnd 0.006187f
C4282 vdd.n2023 gnd 0.006187f
C4283 vdd.n2024 gnd 0.006187f
C4284 vdd.n2025 gnd 0.006187f
C4285 vdd.n2026 gnd 0.562578f
C4286 vdd.n2027 gnd 0.006187f
C4287 vdd.n2028 gnd 0.006187f
C4288 vdd.n2029 gnd 0.006187f
C4289 vdd.n2030 gnd 0.006187f
C4290 vdd.n2031 gnd 0.006187f
C4291 vdd.n2032 gnd 0.502136f
C4292 vdd.n2033 gnd 0.006187f
C4293 vdd.n2034 gnd 0.006187f
C4294 vdd.n2035 gnd 0.006187f
C4295 vdd.n2036 gnd 0.006187f
C4296 vdd.n2037 gnd 0.006187f
C4297 vdd.n2038 gnd 0.362654f
C4298 vdd.n2039 gnd 0.006187f
C4299 vdd.n2040 gnd 0.006187f
C4300 vdd.n2041 gnd 0.006187f
C4301 vdd.n2042 gnd 0.006187f
C4302 vdd.n2043 gnd 0.006187f
C4303 vdd.n2044 gnd 0.199924f
C4304 vdd.n2045 gnd 0.006187f
C4305 vdd.n2046 gnd 0.006187f
C4306 vdd.n2047 gnd 0.006187f
C4307 vdd.n2048 gnd 0.006187f
C4308 vdd.n2049 gnd 0.006187f
C4309 vdd.n2050 gnd 0.348705f
C4310 vdd.n2051 gnd 0.006187f
C4311 vdd.n2052 gnd 0.006187f
C4312 vdd.n2053 gnd 0.006187f
C4313 vdd.n2054 gnd 0.006187f
C4314 vdd.n2055 gnd 0.006187f
C4315 vdd.n2056 gnd 0.632319f
C4316 vdd.n2057 gnd 0.006187f
C4317 vdd.n2058 gnd 0.006187f
C4318 vdd.n2059 gnd 0.006187f
C4319 vdd.n2060 gnd 0.006187f
C4320 vdd.n2061 gnd 0.006187f
C4321 vdd.n2062 gnd 0.006187f
C4322 vdd.n2063 gnd 0.006187f
C4323 vdd.n2064 gnd 0.492837f
C4324 vdd.n2065 gnd 0.006187f
C4325 vdd.n2066 gnd 0.006187f
C4326 vdd.n2067 gnd 0.006187f
C4327 vdd.n2068 gnd 0.006187f
C4328 vdd.n2069 gnd 0.006187f
C4329 vdd.n2070 gnd 0.006187f
C4330 vdd.n2071 gnd 0.395199f
C4331 vdd.n2072 gnd 0.006187f
C4332 vdd.n2073 gnd 0.006187f
C4333 vdd.n2074 gnd 0.006187f
C4334 vdd.n2075 gnd 0.014461f
C4335 vdd.n2076 gnd 0.013928f
C4336 vdd.n2077 gnd 0.006187f
C4337 vdd.n2078 gnd 0.006187f
C4338 vdd.n2079 gnd 0.004777f
C4339 vdd.n2080 gnd 0.006187f
C4340 vdd.n2081 gnd 0.006187f
C4341 vdd.n2082 gnd 0.004504f
C4342 vdd.n2083 gnd 0.006187f
C4343 vdd.n2084 gnd 0.006187f
C4344 vdd.n2085 gnd 0.006187f
C4345 vdd.n2086 gnd 0.006187f
C4346 vdd.n2087 gnd 0.006187f
C4347 vdd.n2088 gnd 0.006187f
C4348 vdd.n2089 gnd 0.006187f
C4349 vdd.n2090 gnd 0.006187f
C4350 vdd.n2091 gnd 0.006187f
C4351 vdd.n2092 gnd 0.006187f
C4352 vdd.n2093 gnd 0.006187f
C4353 vdd.n2094 gnd 0.006187f
C4354 vdd.n2095 gnd 0.006187f
C4355 vdd.n2096 gnd 0.006187f
C4356 vdd.n2097 gnd 0.006187f
C4357 vdd.n2098 gnd 0.006187f
C4358 vdd.n2099 gnd 0.006187f
C4359 vdd.n2100 gnd 0.006187f
C4360 vdd.n2101 gnd 0.006187f
C4361 vdd.n2102 gnd 0.006187f
C4362 vdd.n2103 gnd 0.006187f
C4363 vdd.n2104 gnd 0.006187f
C4364 vdd.n2105 gnd 0.006187f
C4365 vdd.n2106 gnd 0.006187f
C4366 vdd.n2107 gnd 0.006187f
C4367 vdd.n2108 gnd 0.006187f
C4368 vdd.n2109 gnd 0.006187f
C4369 vdd.n2110 gnd 0.006187f
C4370 vdd.n2111 gnd 0.006187f
C4371 vdd.n2112 gnd 0.006187f
C4372 vdd.n2113 gnd 0.006187f
C4373 vdd.n2114 gnd 0.006187f
C4374 vdd.n2115 gnd 0.006187f
C4375 vdd.n2116 gnd 0.006187f
C4376 vdd.n2117 gnd 0.006187f
C4377 vdd.n2118 gnd 0.006187f
C4378 vdd.n2119 gnd 0.006187f
C4379 vdd.n2120 gnd 0.006187f
C4380 vdd.n2121 gnd 0.006187f
C4381 vdd.n2122 gnd 0.006187f
C4382 vdd.n2123 gnd 0.006187f
C4383 vdd.n2124 gnd 0.006187f
C4384 vdd.n2125 gnd 0.006187f
C4385 vdd.n2126 gnd 0.006187f
C4386 vdd.n2127 gnd 0.006187f
C4387 vdd.n2128 gnd 0.006187f
C4388 vdd.n2129 gnd 0.006187f
C4389 vdd.n2130 gnd 0.006187f
C4390 vdd.n2131 gnd 0.006187f
C4391 vdd.n2132 gnd 0.006187f
C4392 vdd.n2133 gnd 0.006187f
C4393 vdd.n2134 gnd 0.006187f
C4394 vdd.n2135 gnd 0.006187f
C4395 vdd.n2136 gnd 0.006187f
C4396 vdd.n2137 gnd 0.006187f
C4397 vdd.n2138 gnd 0.006187f
C4398 vdd.n2139 gnd 0.006187f
C4399 vdd.n2140 gnd 0.006187f
C4400 vdd.n2141 gnd 0.006187f
C4401 vdd.n2142 gnd 0.006187f
C4402 vdd.n2143 gnd 0.014682f
C4403 vdd.n2144 gnd 0.013708f
C4404 vdd.n2145 gnd 0.013708f
C4405 vdd.n2146 gnd 0.771801f
C4406 vdd.n2147 gnd 0.013708f
C4407 vdd.n2148 gnd 0.014682f
C4408 vdd.n2149 gnd 0.013928f
C4409 vdd.n2150 gnd 0.006187f
C4410 vdd.n2151 gnd 0.006187f
C4411 vdd.n2152 gnd 0.006187f
C4412 vdd.n2153 gnd 0.004777f
C4413 vdd.n2154 gnd 0.008843f
C4414 vdd.n2155 gnd 0.004504f
C4415 vdd.n2156 gnd 0.006187f
C4416 vdd.n2157 gnd 0.006187f
C4417 vdd.n2158 gnd 0.006187f
C4418 vdd.n2159 gnd 0.006187f
C4419 vdd.n2160 gnd 0.006187f
C4420 vdd.n2161 gnd 0.006187f
C4421 vdd.n2162 gnd 0.006187f
C4422 vdd.n2163 gnd 0.006187f
C4423 vdd.n2164 gnd 0.006187f
C4424 vdd.n2165 gnd 0.006187f
C4425 vdd.n2166 gnd 0.006187f
C4426 vdd.n2167 gnd 0.006187f
C4427 vdd.n2168 gnd 0.006187f
C4428 vdd.n2169 gnd 0.006187f
C4429 vdd.n2170 gnd 0.006187f
C4430 vdd.n2171 gnd 0.006187f
C4431 vdd.n2172 gnd 0.006187f
C4432 vdd.n2173 gnd 0.006187f
C4433 vdd.n2174 gnd 0.006187f
C4434 vdd.n2175 gnd 0.006187f
C4435 vdd.n2176 gnd 0.006187f
C4436 vdd.n2177 gnd 0.006187f
C4437 vdd.n2178 gnd 0.006187f
C4438 vdd.n2179 gnd 0.006187f
C4439 vdd.n2180 gnd 0.006187f
C4440 vdd.n2181 gnd 0.006187f
C4441 vdd.n2182 gnd 0.006187f
C4442 vdd.n2183 gnd 0.006187f
C4443 vdd.n2184 gnd 0.006187f
C4444 vdd.n2185 gnd 0.006187f
C4445 vdd.n2186 gnd 0.006187f
C4446 vdd.n2187 gnd 0.006187f
C4447 vdd.n2188 gnd 0.006187f
C4448 vdd.n2189 gnd 0.006187f
C4449 vdd.n2190 gnd 0.006187f
C4450 vdd.n2191 gnd 0.006187f
C4451 vdd.n2192 gnd 0.006187f
C4452 vdd.n2193 gnd 0.006187f
C4453 vdd.n2194 gnd 0.006187f
C4454 vdd.n2195 gnd 0.006187f
C4455 vdd.n2196 gnd 0.006187f
C4456 vdd.n2197 gnd 0.006187f
C4457 vdd.n2198 gnd 0.006187f
C4458 vdd.n2199 gnd 0.006187f
C4459 vdd.n2200 gnd 0.006187f
C4460 vdd.n2201 gnd 0.006187f
C4461 vdd.n2202 gnd 0.006187f
C4462 vdd.n2203 gnd 0.006187f
C4463 vdd.n2204 gnd 0.006187f
C4464 vdd.n2205 gnd 0.006187f
C4465 vdd.n2206 gnd 0.006187f
C4466 vdd.n2207 gnd 0.006187f
C4467 vdd.n2208 gnd 0.006187f
C4468 vdd.n2209 gnd 0.006187f
C4469 vdd.n2210 gnd 0.006187f
C4470 vdd.n2211 gnd 0.006187f
C4471 vdd.n2212 gnd 0.006187f
C4472 vdd.n2213 gnd 0.006187f
C4473 vdd.n2214 gnd 0.006187f
C4474 vdd.n2215 gnd 0.006187f
C4475 vdd.n2216 gnd 0.014682f
C4476 vdd.n2217 gnd 0.014682f
C4477 vdd.n2218 gnd 0.771801f
C4478 vdd.t165 gnd 2.74315f
C4479 vdd.t155 gnd 2.74315f
C4480 vdd.n2251 gnd 0.014682f
C4481 vdd.n2252 gnd 0.006187f
C4482 vdd.t62 gnd 0.25003f
C4483 vdd.t63 gnd 0.255937f
C4484 vdd.t60 gnd 0.163229f
C4485 vdd.n2253 gnd 0.088216f
C4486 vdd.n2254 gnd 0.050039f
C4487 vdd.n2255 gnd 0.006187f
C4488 vdd.t75 gnd 0.25003f
C4489 vdd.t76 gnd 0.255937f
C4490 vdd.t74 gnd 0.163229f
C4491 vdd.n2256 gnd 0.088216f
C4492 vdd.n2257 gnd 0.050039f
C4493 vdd.n2258 gnd 0.008843f
C4494 vdd.n2259 gnd 0.006187f
C4495 vdd.n2260 gnd 0.006187f
C4496 vdd.n2261 gnd 0.006187f
C4497 vdd.n2262 gnd 0.006187f
C4498 vdd.n2263 gnd 0.006187f
C4499 vdd.n2264 gnd 0.006187f
C4500 vdd.n2265 gnd 0.006187f
C4501 vdd.n2266 gnd 0.006187f
C4502 vdd.n2267 gnd 0.006187f
C4503 vdd.n2268 gnd 0.006187f
C4504 vdd.n2269 gnd 0.006187f
C4505 vdd.n2270 gnd 0.006187f
C4506 vdd.n2271 gnd 0.006187f
C4507 vdd.n2272 gnd 0.006187f
C4508 vdd.n2273 gnd 0.006187f
C4509 vdd.n2274 gnd 0.006187f
C4510 vdd.n2275 gnd 0.006187f
C4511 vdd.n2276 gnd 0.006187f
C4512 vdd.n2277 gnd 0.006187f
C4513 vdd.n2278 gnd 0.006187f
C4514 vdd.n2279 gnd 0.006187f
C4515 vdd.n2280 gnd 0.006187f
C4516 vdd.n2281 gnd 0.006187f
C4517 vdd.n2282 gnd 0.006187f
C4518 vdd.n2283 gnd 0.006187f
C4519 vdd.n2284 gnd 0.006187f
C4520 vdd.n2285 gnd 0.006187f
C4521 vdd.n2286 gnd 0.006187f
C4522 vdd.n2287 gnd 0.006187f
C4523 vdd.n2288 gnd 0.006187f
C4524 vdd.n2289 gnd 0.006187f
C4525 vdd.n2290 gnd 0.006187f
C4526 vdd.n2291 gnd 0.006187f
C4527 vdd.n2292 gnd 0.006187f
C4528 vdd.n2293 gnd 0.006187f
C4529 vdd.n2294 gnd 0.006187f
C4530 vdd.n2295 gnd 0.006187f
C4531 vdd.n2296 gnd 0.006187f
C4532 vdd.n2297 gnd 0.006187f
C4533 vdd.n2298 gnd 0.006187f
C4534 vdd.n2299 gnd 0.006187f
C4535 vdd.n2300 gnd 0.006187f
C4536 vdd.n2301 gnd 0.006187f
C4537 vdd.n2302 gnd 0.006187f
C4538 vdd.n2303 gnd 0.006187f
C4539 vdd.n2304 gnd 0.006187f
C4540 vdd.n2305 gnd 0.006187f
C4541 vdd.n2306 gnd 0.006187f
C4542 vdd.n2307 gnd 0.006187f
C4543 vdd.n2308 gnd 0.006187f
C4544 vdd.n2309 gnd 0.006187f
C4545 vdd.n2310 gnd 0.006187f
C4546 vdd.n2311 gnd 0.006187f
C4547 vdd.n2312 gnd 0.006187f
C4548 vdd.n2313 gnd 0.006187f
C4549 vdd.n2314 gnd 0.006187f
C4550 vdd.n2315 gnd 0.004504f
C4551 vdd.n2316 gnd 0.006187f
C4552 vdd.n2317 gnd 0.006187f
C4553 vdd.n2318 gnd 0.004777f
C4554 vdd.n2319 gnd 0.006187f
C4555 vdd.n2320 gnd 0.006187f
C4556 vdd.n2321 gnd 0.014682f
C4557 vdd.n2322 gnd 0.013708f
C4558 vdd.n2323 gnd 0.006187f
C4559 vdd.n2324 gnd 0.006187f
C4560 vdd.n2325 gnd 0.006187f
C4561 vdd.n2326 gnd 0.006187f
C4562 vdd.n2327 gnd 0.006187f
C4563 vdd.n2328 gnd 0.006187f
C4564 vdd.n2329 gnd 0.006187f
C4565 vdd.n2330 gnd 0.006187f
C4566 vdd.n2331 gnd 0.006187f
C4567 vdd.n2332 gnd 0.006187f
C4568 vdd.n2333 gnd 0.006187f
C4569 vdd.n2334 gnd 0.006187f
C4570 vdd.n2335 gnd 0.006187f
C4571 vdd.n2336 gnd 0.006187f
C4572 vdd.n2337 gnd 0.006187f
C4573 vdd.n2338 gnd 0.006187f
C4574 vdd.n2339 gnd 0.006187f
C4575 vdd.n2340 gnd 0.006187f
C4576 vdd.n2341 gnd 0.006187f
C4577 vdd.n2342 gnd 0.006187f
C4578 vdd.n2343 gnd 0.006187f
C4579 vdd.n2344 gnd 0.006187f
C4580 vdd.n2345 gnd 0.006187f
C4581 vdd.n2346 gnd 0.006187f
C4582 vdd.n2347 gnd 0.006187f
C4583 vdd.n2348 gnd 0.006187f
C4584 vdd.n2349 gnd 0.006187f
C4585 vdd.n2350 gnd 0.006187f
C4586 vdd.n2351 gnd 0.006187f
C4587 vdd.n2352 gnd 0.006187f
C4588 vdd.n2353 gnd 0.006187f
C4589 vdd.n2354 gnd 0.006187f
C4590 vdd.n2355 gnd 0.006187f
C4591 vdd.n2356 gnd 0.006187f
C4592 vdd.n2357 gnd 0.006187f
C4593 vdd.n2358 gnd 0.006187f
C4594 vdd.n2359 gnd 0.006187f
C4595 vdd.n2360 gnd 0.006187f
C4596 vdd.n2361 gnd 0.006187f
C4597 vdd.n2362 gnd 0.006187f
C4598 vdd.n2363 gnd 0.006187f
C4599 vdd.n2364 gnd 0.006187f
C4600 vdd.n2365 gnd 0.006187f
C4601 vdd.n2366 gnd 0.006187f
C4602 vdd.n2367 gnd 0.006187f
C4603 vdd.n2368 gnd 0.006187f
C4604 vdd.n2369 gnd 0.006187f
C4605 vdd.n2370 gnd 0.006187f
C4606 vdd.n2371 gnd 0.006187f
C4607 vdd.n2372 gnd 0.006187f
C4608 vdd.n2373 gnd 0.006187f
C4609 vdd.n2374 gnd 0.199924f
C4610 vdd.n2375 gnd 0.006187f
C4611 vdd.n2376 gnd 0.006187f
C4612 vdd.n2377 gnd 0.006187f
C4613 vdd.n2378 gnd 0.006187f
C4614 vdd.n2379 gnd 0.006187f
C4615 vdd.n2380 gnd 0.006187f
C4616 vdd.n2381 gnd 0.006187f
C4617 vdd.n2382 gnd 0.006187f
C4618 vdd.n2383 gnd 0.006187f
C4619 vdd.n2384 gnd 0.006187f
C4620 vdd.n2385 gnd 0.006187f
C4621 vdd.n2386 gnd 0.006187f
C4622 vdd.n2387 gnd 0.006187f
C4623 vdd.n2388 gnd 0.006187f
C4624 vdd.n2389 gnd 0.006187f
C4625 vdd.n2390 gnd 0.006187f
C4626 vdd.n2391 gnd 0.006187f
C4627 vdd.n2392 gnd 0.006187f
C4628 vdd.n2393 gnd 0.006187f
C4629 vdd.n2394 gnd 0.006187f
C4630 vdd.n2395 gnd 0.376602f
C4631 vdd.n2396 gnd 0.006187f
C4632 vdd.n2397 gnd 0.006187f
C4633 vdd.n2398 gnd 0.006187f
C4634 vdd.n2399 gnd 0.006187f
C4635 vdd.n2400 gnd 0.006187f
C4636 vdd.n2401 gnd 0.013708f
C4637 vdd.n2402 gnd 0.014682f
C4638 vdd.n2403 gnd 0.014682f
C4639 vdd.n2404 gnd 0.006187f
C4640 vdd.n2405 gnd 0.006187f
C4641 vdd.n2406 gnd 0.006187f
C4642 vdd.n2407 gnd 0.004777f
C4643 vdd.n2408 gnd 0.008843f
C4644 vdd.n2409 gnd 0.004504f
C4645 vdd.n2410 gnd 0.006187f
C4646 vdd.n2411 gnd 0.006187f
C4647 vdd.n2412 gnd 0.006187f
C4648 vdd.n2413 gnd 0.006187f
C4649 vdd.n2414 gnd 0.006187f
C4650 vdd.n2415 gnd 0.006187f
C4651 vdd.n2416 gnd 0.006187f
C4652 vdd.n2417 gnd 0.006187f
C4653 vdd.n2418 gnd 0.006187f
C4654 vdd.n2419 gnd 0.006187f
C4655 vdd.n2420 gnd 0.006187f
C4656 vdd.n2421 gnd 0.006187f
C4657 vdd.n2422 gnd 0.006187f
C4658 vdd.n2423 gnd 0.006187f
C4659 vdd.n2424 gnd 0.006187f
C4660 vdd.n2425 gnd 0.006187f
C4661 vdd.n2426 gnd 0.006187f
C4662 vdd.n2427 gnd 0.006187f
C4663 vdd.n2428 gnd 0.006187f
C4664 vdd.n2429 gnd 0.006187f
C4665 vdd.n2430 gnd 0.006187f
C4666 vdd.n2431 gnd 0.006187f
C4667 vdd.n2432 gnd 0.006187f
C4668 vdd.n2433 gnd 0.006187f
C4669 vdd.n2434 gnd 0.006187f
C4670 vdd.n2435 gnd 0.006187f
C4671 vdd.n2436 gnd 0.006187f
C4672 vdd.n2437 gnd 0.006187f
C4673 vdd.n2438 gnd 0.006187f
C4674 vdd.n2439 gnd 0.006187f
C4675 vdd.n2440 gnd 0.006187f
C4676 vdd.n2441 gnd 0.006187f
C4677 vdd.n2442 gnd 0.006187f
C4678 vdd.n2443 gnd 0.006187f
C4679 vdd.n2444 gnd 0.006187f
C4680 vdd.n2445 gnd 0.006187f
C4681 vdd.n2446 gnd 0.006187f
C4682 vdd.n2447 gnd 0.006187f
C4683 vdd.n2448 gnd 0.006187f
C4684 vdd.n2449 gnd 0.006187f
C4685 vdd.n2450 gnd 0.006187f
C4686 vdd.n2451 gnd 0.006187f
C4687 vdd.n2452 gnd 0.006187f
C4688 vdd.n2453 gnd 0.006187f
C4689 vdd.n2454 gnd 0.006187f
C4690 vdd.n2455 gnd 0.006187f
C4691 vdd.n2456 gnd 0.006187f
C4692 vdd.n2457 gnd 0.006187f
C4693 vdd.n2458 gnd 0.006187f
C4694 vdd.n2459 gnd 0.006187f
C4695 vdd.n2460 gnd 0.006187f
C4696 vdd.n2461 gnd 0.006187f
C4697 vdd.n2462 gnd 0.006187f
C4698 vdd.n2463 gnd 0.006187f
C4699 vdd.n2464 gnd 0.006187f
C4700 vdd.n2465 gnd 0.006187f
C4701 vdd.n2466 gnd 0.006187f
C4702 vdd.n2467 gnd 0.006187f
C4703 vdd.n2468 gnd 0.006187f
C4704 vdd.n2469 gnd 0.006187f
C4705 vdd.n2471 gnd 0.771801f
C4706 vdd.n2473 gnd 0.006187f
C4707 vdd.n2474 gnd 0.006187f
C4708 vdd.n2475 gnd 0.014682f
C4709 vdd.n2476 gnd 0.013708f
C4710 vdd.n2477 gnd 0.013708f
C4711 vdd.n2478 gnd 0.771801f
C4712 vdd.n2479 gnd 0.013708f
C4713 vdd.n2480 gnd 0.013708f
C4714 vdd.n2481 gnd 0.006187f
C4715 vdd.n2482 gnd 0.006187f
C4716 vdd.n2483 gnd 0.006187f
C4717 vdd.n2484 gnd 0.395199f
C4718 vdd.n2485 gnd 0.006187f
C4719 vdd.n2486 gnd 0.006187f
C4720 vdd.n2487 gnd 0.006187f
C4721 vdd.n2488 gnd 0.006187f
C4722 vdd.n2489 gnd 0.006187f
C4723 vdd.n2490 gnd 0.492837f
C4724 vdd.n2491 gnd 0.006187f
C4725 vdd.n2492 gnd 0.006187f
C4726 vdd.n2493 gnd 0.006187f
C4727 vdd.n2494 gnd 0.006187f
C4728 vdd.n2495 gnd 0.006187f
C4729 vdd.n2496 gnd 0.632319f
C4730 vdd.n2497 gnd 0.006187f
C4731 vdd.n2498 gnd 0.006187f
C4732 vdd.n2499 gnd 0.006187f
C4733 vdd.n2500 gnd 0.006187f
C4734 vdd.n2501 gnd 0.006187f
C4735 vdd.n2502 gnd 0.348705f
C4736 vdd.n2503 gnd 0.006187f
C4737 vdd.n2504 gnd 0.006187f
C4738 vdd.n2505 gnd 0.006187f
C4739 vdd.n2506 gnd 0.006187f
C4740 vdd.n2507 gnd 0.006187f
C4741 vdd.n2508 gnd 0.199924f
C4742 vdd.n2509 gnd 0.006187f
C4743 vdd.n2510 gnd 0.006187f
C4744 vdd.n2511 gnd 0.006187f
C4745 vdd.n2512 gnd 0.006187f
C4746 vdd.n2513 gnd 0.006187f
C4747 vdd.n2514 gnd 0.362654f
C4748 vdd.n2515 gnd 0.006187f
C4749 vdd.n2516 gnd 0.006187f
C4750 vdd.n2517 gnd 0.006187f
C4751 vdd.n2518 gnd 0.006187f
C4752 vdd.n2519 gnd 0.006187f
C4753 vdd.n2520 gnd 0.502136f
C4754 vdd.n2521 gnd 0.006187f
C4755 vdd.n2522 gnd 0.006187f
C4756 vdd.n2523 gnd 0.006187f
C4757 vdd.n2524 gnd 0.006187f
C4758 vdd.n2525 gnd 0.006187f
C4759 vdd.n2526 gnd 0.562578f
C4760 vdd.n2527 gnd 0.006187f
C4761 vdd.n2528 gnd 0.006187f
C4762 vdd.n2529 gnd 0.006187f
C4763 vdd.n2530 gnd 0.006187f
C4764 vdd.n2531 gnd 0.006187f
C4765 vdd.n2532 gnd 0.423096f
C4766 vdd.n2533 gnd 0.006187f
C4767 vdd.n2534 gnd 0.006187f
C4768 vdd.n2535 gnd 0.006187f
C4769 vdd.t37 gnd 0.255937f
C4770 vdd.t35 gnd 0.163229f
C4771 vdd.t38 gnd 0.255937f
C4772 vdd.n2536 gnd 0.143847f
C4773 vdd.n2537 gnd 0.017924f
C4774 vdd.n2538 gnd 0.003822f
C4775 vdd.n2539 gnd 0.006187f
C4776 vdd.n2540 gnd 0.348705f
C4777 vdd.n2541 gnd 0.006187f
C4778 vdd.n2542 gnd 0.006187f
C4779 vdd.n2543 gnd 0.006187f
C4780 vdd.n2544 gnd 0.006187f
C4781 vdd.n2545 gnd 0.006187f
C4782 vdd.n2546 gnd 0.632319f
C4783 vdd.n2547 gnd 0.006187f
C4784 vdd.n2548 gnd 0.006187f
C4785 vdd.n2549 gnd 0.006187f
C4786 vdd.n2550 gnd 0.006187f
C4787 vdd.n2551 gnd 0.006187f
C4788 vdd.n2552 gnd 0.006187f
C4789 vdd.n2554 gnd 0.006187f
C4790 vdd.n2555 gnd 0.006187f
C4791 vdd.n2557 gnd 0.006187f
C4792 vdd.n2558 gnd 0.006187f
C4793 vdd.n2561 gnd 0.006187f
C4794 vdd.n2562 gnd 0.006187f
C4795 vdd.n2563 gnd 0.006187f
C4796 vdd.n2564 gnd 0.006187f
C4797 vdd.n2566 gnd 0.006187f
C4798 vdd.n2567 gnd 0.006187f
C4799 vdd.n2568 gnd 0.006187f
C4800 vdd.n2569 gnd 0.006187f
C4801 vdd.n2570 gnd 0.006187f
C4802 vdd.n2571 gnd 0.006187f
C4803 vdd.n2573 gnd 0.006187f
C4804 vdd.n2574 gnd 0.006187f
C4805 vdd.n2575 gnd 0.006187f
C4806 vdd.n2576 gnd 0.006187f
C4807 vdd.n2577 gnd 0.006187f
C4808 vdd.n2578 gnd 0.006187f
C4809 vdd.n2580 gnd 0.006187f
C4810 vdd.n2581 gnd 0.006187f
C4811 vdd.n2582 gnd 0.006187f
C4812 vdd.n2583 gnd 0.006187f
C4813 vdd.n2584 gnd 0.006187f
C4814 vdd.n2585 gnd 0.006187f
C4815 vdd.n2587 gnd 0.006187f
C4816 vdd.n2588 gnd 0.014682f
C4817 vdd.n2589 gnd 0.014682f
C4818 vdd.n2590 gnd 0.013708f
C4819 vdd.n2591 gnd 0.006187f
C4820 vdd.n2592 gnd 0.006187f
C4821 vdd.n2593 gnd 0.006187f
C4822 vdd.n2594 gnd 0.006187f
C4823 vdd.n2595 gnd 0.006187f
C4824 vdd.n2596 gnd 0.006187f
C4825 vdd.n2597 gnd 0.632319f
C4826 vdd.n2598 gnd 0.006187f
C4827 vdd.n2599 gnd 0.006187f
C4828 vdd.n2600 gnd 0.006187f
C4829 vdd.n2601 gnd 0.006187f
C4830 vdd.n2602 gnd 0.006187f
C4831 vdd.n2603 gnd 0.395199f
C4832 vdd.n2604 gnd 0.006187f
C4833 vdd.n2605 gnd 0.006187f
C4834 vdd.n2606 gnd 0.006187f
C4835 vdd.n2607 gnd 0.014461f
C4836 vdd.n2608 gnd 0.013928f
C4837 vdd.n2609 gnd 0.014682f
C4838 vdd.n2611 gnd 0.006187f
C4839 vdd.n2612 gnd 0.006187f
C4840 vdd.n2613 gnd 0.004777f
C4841 vdd.n2614 gnd 0.008843f
C4842 vdd.n2615 gnd 0.004504f
C4843 vdd.n2616 gnd 0.006187f
C4844 vdd.n2617 gnd 0.006187f
C4845 vdd.n2619 gnd 0.006187f
C4846 vdd.n2620 gnd 0.006187f
C4847 vdd.n2621 gnd 0.006187f
C4848 vdd.n2622 gnd 0.006187f
C4849 vdd.n2623 gnd 0.006187f
C4850 vdd.n2624 gnd 0.006187f
C4851 vdd.n2626 gnd 0.006187f
C4852 vdd.n2627 gnd 0.006187f
C4853 vdd.n2628 gnd 0.006187f
C4854 vdd.n2629 gnd 0.006187f
C4855 vdd.n2630 gnd 0.006187f
C4856 vdd.n2631 gnd 0.006187f
C4857 vdd.n2633 gnd 0.006187f
C4858 vdd.n2634 gnd 0.006187f
C4859 vdd.n2635 gnd 0.006187f
C4860 vdd.n2636 gnd 0.006187f
C4861 vdd.n2637 gnd 0.006187f
C4862 vdd.n2638 gnd 0.006187f
C4863 vdd.n2640 gnd 0.006187f
C4864 vdd.n2641 gnd 0.006187f
C4865 vdd.n2642 gnd 0.006187f
C4866 vdd.n2644 gnd 0.006187f
C4867 vdd.n2645 gnd 0.006187f
C4868 vdd.n2646 gnd 0.006187f
C4869 vdd.n2647 gnd 0.006187f
C4870 vdd.n2648 gnd 0.006187f
C4871 vdd.n2649 gnd 0.006187f
C4872 vdd.n2651 gnd 0.006187f
C4873 vdd.n2652 gnd 0.006187f
C4874 vdd.n2653 gnd 0.006187f
C4875 vdd.n2654 gnd 0.006187f
C4876 vdd.n2655 gnd 0.006187f
C4877 vdd.n2656 gnd 0.006187f
C4878 vdd.n2658 gnd 0.006187f
C4879 vdd.n2659 gnd 0.006187f
C4880 vdd.n2660 gnd 0.006187f
C4881 vdd.n2661 gnd 0.006187f
C4882 vdd.n2662 gnd 0.006187f
C4883 vdd.n2663 gnd 0.006187f
C4884 vdd.n2665 gnd 0.006187f
C4885 vdd.n2666 gnd 0.006187f
C4886 vdd.n2668 gnd 0.006187f
C4887 vdd.n2669 gnd 0.006187f
C4888 vdd.n2670 gnd 0.014682f
C4889 vdd.n2671 gnd 0.013708f
C4890 vdd.n2672 gnd 0.013708f
C4891 vdd.n2673 gnd 0.911283f
C4892 vdd.n2674 gnd 0.013708f
C4893 vdd.n2675 gnd 0.014682f
C4894 vdd.n2676 gnd 0.013928f
C4895 vdd.n2677 gnd 0.006187f
C4896 vdd.n2678 gnd 0.004777f
C4897 vdd.n2679 gnd 0.006187f
C4898 vdd.n2681 gnd 0.006187f
C4899 vdd.n2682 gnd 0.006187f
C4900 vdd.n2683 gnd 0.006187f
C4901 vdd.n2684 gnd 0.006187f
C4902 vdd.n2685 gnd 0.006187f
C4903 vdd.n2686 gnd 0.006187f
C4904 vdd.n2688 gnd 0.006187f
C4905 vdd.n2689 gnd 0.006187f
C4906 vdd.n2690 gnd 0.006187f
C4907 vdd.n2691 gnd 0.006187f
C4908 vdd.n2692 gnd 0.006187f
C4909 vdd.n2693 gnd 0.006187f
C4910 vdd.n2695 gnd 0.006187f
C4911 vdd.n2696 gnd 0.006187f
C4912 vdd.n2697 gnd 0.006187f
C4913 vdd.n2698 gnd 0.006187f
C4914 vdd.n2699 gnd 0.006187f
C4915 vdd.n2700 gnd 0.006187f
C4916 vdd.n2702 gnd 0.006187f
C4917 vdd.n2703 gnd 0.006187f
C4918 vdd.n2705 gnd 0.006187f
C4919 vdd.n2706 gnd 0.014868f
C4920 vdd.n2707 gnd 0.55069f
C4921 vdd.n2708 gnd 0.007825f
C4922 vdd.n2709 gnd 0.022684f
C4923 vdd.n2710 gnd 0.003479f
C4924 vdd.t87 gnd 0.111942f
C4925 vdd.t88 gnd 0.119636f
C4926 vdd.t86 gnd 0.146195f
C4927 vdd.n2711 gnd 0.187402f
C4928 vdd.n2712 gnd 0.157451f
C4929 vdd.n2713 gnd 0.011278f
C4930 vdd.n2714 gnd 0.009099f
C4931 vdd.n2715 gnd 0.003845f
C4932 vdd.n2716 gnd 0.007324f
C4933 vdd.n2717 gnd 0.009099f
C4934 vdd.n2718 gnd 0.009099f
C4935 vdd.n2719 gnd 0.007324f
C4936 vdd.n2720 gnd 0.007324f
C4937 vdd.n2721 gnd 0.009099f
C4938 vdd.n2722 gnd 0.009099f
C4939 vdd.n2723 gnd 0.007324f
C4940 vdd.n2724 gnd 0.007324f
C4941 vdd.n2725 gnd 0.009099f
C4942 vdd.n2726 gnd 0.009099f
C4943 vdd.n2727 gnd 0.007324f
C4944 vdd.n2728 gnd 0.007324f
C4945 vdd.n2729 gnd 0.009099f
C4946 vdd.n2730 gnd 0.009099f
C4947 vdd.n2731 gnd 0.007324f
C4948 vdd.n2732 gnd 0.007324f
C4949 vdd.n2733 gnd 0.009099f
C4950 vdd.n2734 gnd 0.009099f
C4951 vdd.n2735 gnd 0.007324f
C4952 vdd.n2736 gnd 0.007324f
C4953 vdd.n2737 gnd 0.009099f
C4954 vdd.n2738 gnd 0.009099f
C4955 vdd.n2739 gnd 0.007324f
C4956 vdd.n2740 gnd 0.007324f
C4957 vdd.n2741 gnd 0.009099f
C4958 vdd.n2742 gnd 0.009099f
C4959 vdd.n2743 gnd 0.007324f
C4960 vdd.n2744 gnd 0.007324f
C4961 vdd.n2745 gnd 0.009099f
C4962 vdd.n2746 gnd 0.009099f
C4963 vdd.n2747 gnd 0.007324f
C4964 vdd.n2748 gnd 0.007324f
C4965 vdd.n2749 gnd 0.009099f
C4966 vdd.n2750 gnd 0.009099f
C4967 vdd.n2751 gnd 0.007324f
C4968 vdd.n2752 gnd 0.009099f
C4969 vdd.n2753 gnd 0.009099f
C4970 vdd.n2754 gnd 0.007324f
C4971 vdd.n2755 gnd 0.009099f
C4972 vdd.n2756 gnd 0.009099f
C4973 vdd.n2757 gnd 0.009099f
C4974 vdd.n2758 gnd 0.01494f
C4975 vdd.n2759 gnd 0.009099f
C4976 vdd.n2760 gnd 0.009099f
C4977 vdd.n2761 gnd 0.00498f
C4978 vdd.n2762 gnd 0.007324f
C4979 vdd.n2763 gnd 0.009099f
C4980 vdd.n2764 gnd 0.009099f
C4981 vdd.n2765 gnd 0.007324f
C4982 vdd.n2766 gnd 0.007324f
C4983 vdd.n2767 gnd 0.009099f
C4984 vdd.n2768 gnd 0.009099f
C4985 vdd.n2769 gnd 0.007324f
C4986 vdd.n2770 gnd 0.007324f
C4987 vdd.n2771 gnd 0.009099f
C4988 vdd.n2772 gnd 0.009099f
C4989 vdd.n2773 gnd 0.007324f
C4990 vdd.n2774 gnd 0.007324f
C4991 vdd.n2775 gnd 0.009099f
C4992 vdd.n2776 gnd 0.009099f
C4993 vdd.n2777 gnd 0.007324f
C4994 vdd.n2778 gnd 0.007324f
C4995 vdd.n2779 gnd 0.009099f
C4996 vdd.n2780 gnd 0.009099f
C4997 vdd.n2781 gnd 0.007324f
C4998 vdd.n2782 gnd 0.007324f
C4999 vdd.n2783 gnd 0.009099f
C5000 vdd.n2784 gnd 0.009099f
C5001 vdd.n2785 gnd 0.007324f
C5002 vdd.n2786 gnd 0.007324f
C5003 vdd.n2787 gnd 0.009099f
C5004 vdd.n2788 gnd 0.009099f
C5005 vdd.n2789 gnd 0.007324f
C5006 vdd.n2790 gnd 0.007324f
C5007 vdd.n2791 gnd 0.009099f
C5008 vdd.n2792 gnd 0.009099f
C5009 vdd.n2793 gnd 0.007324f
C5010 vdd.n2794 gnd 0.007324f
C5011 vdd.n2795 gnd 0.009099f
C5012 vdd.n2796 gnd 0.009099f
C5013 vdd.n2797 gnd 0.007324f
C5014 vdd.n2798 gnd 0.009099f
C5015 vdd.n2799 gnd 0.009099f
C5016 vdd.n2800 gnd 0.007324f
C5017 vdd.n2801 gnd 0.009099f
C5018 vdd.n2802 gnd 0.009099f
C5019 vdd.n2803 gnd 0.009099f
C5020 vdd.t25 gnd 0.111942f
C5021 vdd.t26 gnd 0.119636f
C5022 vdd.t24 gnd 0.146195f
C5023 vdd.n2804 gnd 0.187402f
C5024 vdd.n2805 gnd 0.157451f
C5025 vdd.n2806 gnd 0.01494f
C5026 vdd.n2807 gnd 0.009099f
C5027 vdd.n2808 gnd 0.009099f
C5028 vdd.n2809 gnd 0.006115f
C5029 vdd.n2810 gnd 0.007324f
C5030 vdd.n2811 gnd 0.009099f
C5031 vdd.n2812 gnd 0.009099f
C5032 vdd.n2813 gnd 0.007324f
C5033 vdd.n2814 gnd 0.007324f
C5034 vdd.n2815 gnd 0.009099f
C5035 vdd.n2816 gnd 0.009099f
C5036 vdd.n2817 gnd 0.007324f
C5037 vdd.n2818 gnd 0.007324f
C5038 vdd.n2819 gnd 0.009099f
C5039 vdd.n2820 gnd 0.009099f
C5040 vdd.n2821 gnd 0.007324f
C5041 vdd.n2822 gnd 0.007324f
C5042 vdd.n2823 gnd 0.009099f
C5043 vdd.n2824 gnd 0.009099f
C5044 vdd.n2825 gnd 0.007324f
C5045 vdd.n2826 gnd 0.007324f
C5046 vdd.n2827 gnd 0.009099f
C5047 vdd.n2828 gnd 0.009099f
C5048 vdd.n2829 gnd 0.007324f
C5049 vdd.n2830 gnd 0.007324f
C5050 vdd.n2831 gnd 0.009099f
C5051 vdd.n2832 gnd 0.009099f
C5052 vdd.n2833 gnd 0.007324f
C5053 vdd.n2834 gnd 0.007324f
C5054 vdd.n2836 gnd 0.55069f
C5055 vdd.n2838 gnd 0.007324f
C5056 vdd.n2839 gnd 0.009099f
C5057 vdd.n2840 gnd 6.74164f
C5058 vdd.n2842 gnd 0.022684f
C5059 vdd.n2843 gnd 0.006079f
C5060 vdd.n2844 gnd 0.022684f
C5061 vdd.n2845 gnd 0.022175f
C5062 vdd.n2846 gnd 0.009099f
C5063 vdd.n2847 gnd 0.007324f
C5064 vdd.n2848 gnd 0.009099f
C5065 vdd.n2849 gnd 0.581176f
C5066 vdd.n2850 gnd 0.009099f
C5067 vdd.n2851 gnd 0.007324f
C5068 vdd.n2852 gnd 0.009099f
C5069 vdd.n2853 gnd 0.009099f
C5070 vdd.n2854 gnd 0.009099f
C5071 vdd.n2855 gnd 0.007324f
C5072 vdd.n2856 gnd 0.009099f
C5073 vdd.n2857 gnd 0.739255f
C5074 vdd.n2858 gnd 0.929881f
C5075 vdd.n2859 gnd 0.009099f
C5076 vdd.n2860 gnd 0.007324f
C5077 vdd.n2861 gnd 0.009099f
C5078 vdd.n2862 gnd 0.009099f
C5079 vdd.n2863 gnd 0.009099f
C5080 vdd.n2864 gnd 0.007324f
C5081 vdd.n2865 gnd 0.009099f
C5082 vdd.n2866 gnd 0.655566f
C5083 vdd.n2867 gnd 0.009099f
C5084 vdd.n2868 gnd 0.007324f
C5085 vdd.n2869 gnd 0.009099f
C5086 vdd.n2870 gnd 0.009099f
C5087 vdd.n2871 gnd 0.009099f
C5088 vdd.n2872 gnd 0.007324f
C5089 vdd.n2873 gnd 0.009099f
C5090 vdd.t109 gnd 0.46494f
C5091 vdd.n2874 gnd 0.771801f
C5092 vdd.n2875 gnd 0.009099f
C5093 vdd.n2876 gnd 0.007324f
C5094 vdd.n2877 gnd 0.009099f
C5095 vdd.n2878 gnd 0.009099f
C5096 vdd.n2879 gnd 0.009099f
C5097 vdd.n2880 gnd 0.007324f
C5098 vdd.n2881 gnd 0.009099f
C5099 vdd.n2882 gnd 0.729956f
C5100 vdd.n2883 gnd 0.009099f
C5101 vdd.n2884 gnd 0.007324f
C5102 vdd.n2885 gnd 0.009099f
C5103 vdd.n2886 gnd 0.009099f
C5104 vdd.n2887 gnd 0.009099f
C5105 vdd.n2888 gnd 0.007324f
C5106 vdd.n2889 gnd 0.007324f
C5107 vdd.n2890 gnd 0.007324f
C5108 vdd.n2891 gnd 0.009099f
C5109 vdd.n2892 gnd 0.009099f
C5110 vdd.n2893 gnd 0.009099f
C5111 vdd.n2894 gnd 0.007324f
C5112 vdd.n2895 gnd 0.007324f
C5113 vdd.n2896 gnd 0.007324f
C5114 vdd.n2897 gnd 0.009099f
C5115 vdd.n2898 gnd 0.009099f
C5116 vdd.n2899 gnd 0.009099f
C5117 vdd.n2900 gnd 0.007324f
C5118 vdd.n2901 gnd 0.007324f
C5119 vdd.n2902 gnd 0.006079f
C5120 vdd.n2903 gnd 0.022175f
C5121 vdd.n2904 gnd 0.022684f
C5122 vdd.n2906 gnd 0.022684f
C5123 vdd.n2907 gnd 0.003479f
C5124 vdd.t91 gnd 0.111942f
C5125 vdd.t90 gnd 0.119636f
C5126 vdd.t89 gnd 0.146195f
C5127 vdd.n2908 gnd 0.187402f
C5128 vdd.n2909 gnd 0.158184f
C5129 vdd.n2910 gnd 0.012011f
C5130 vdd.n2911 gnd 0.003845f
C5131 vdd.n2912 gnd 0.007324f
C5132 vdd.n2913 gnd 0.009099f
C5133 vdd.n2915 gnd 0.009099f
C5134 vdd.n2916 gnd 0.009099f
C5135 vdd.n2917 gnd 0.007324f
C5136 vdd.n2918 gnd 0.007324f
C5137 vdd.n2919 gnd 0.007324f
C5138 vdd.n2920 gnd 0.009099f
C5139 vdd.n2922 gnd 0.009099f
C5140 vdd.n2923 gnd 0.009099f
C5141 vdd.n2924 gnd 0.007324f
C5142 vdd.n2925 gnd 0.007324f
C5143 vdd.n2926 gnd 0.007324f
C5144 vdd.n2927 gnd 0.009099f
C5145 vdd.n2929 gnd 0.009099f
C5146 vdd.n2930 gnd 0.009099f
C5147 vdd.n2931 gnd 0.007324f
C5148 vdd.n2932 gnd 0.007324f
C5149 vdd.n2933 gnd 0.007324f
C5150 vdd.n2934 gnd 0.009099f
C5151 vdd.n2936 gnd 0.009099f
C5152 vdd.n2937 gnd 0.009099f
C5153 vdd.n2938 gnd 0.007324f
C5154 vdd.n2939 gnd 0.007324f
C5155 vdd.n2940 gnd 0.007324f
C5156 vdd.n2941 gnd 0.009099f
C5157 vdd.n2943 gnd 0.009099f
C5158 vdd.n2944 gnd 0.009099f
C5159 vdd.n2945 gnd 0.007324f
C5160 vdd.n2946 gnd 0.009099f
C5161 vdd.n2947 gnd 0.009099f
C5162 vdd.n2948 gnd 0.009099f
C5163 vdd.n2949 gnd 0.015673f
C5164 vdd.n2950 gnd 0.00498f
C5165 vdd.n2951 gnd 0.007324f
C5166 vdd.n2952 gnd 0.009099f
C5167 vdd.n2954 gnd 0.009099f
C5168 vdd.n2955 gnd 0.009099f
C5169 vdd.n2956 gnd 0.007324f
C5170 vdd.n2957 gnd 0.007324f
C5171 vdd.n2958 gnd 0.007324f
C5172 vdd.n2959 gnd 0.009099f
C5173 vdd.n2961 gnd 0.009099f
C5174 vdd.n2962 gnd 0.009099f
C5175 vdd.n2963 gnd 0.007324f
C5176 vdd.n2964 gnd 0.007324f
C5177 vdd.n2965 gnd 0.007324f
C5178 vdd.n2966 gnd 0.009099f
C5179 vdd.n2968 gnd 0.009099f
C5180 vdd.n2969 gnd 0.009099f
C5181 vdd.n2970 gnd 0.007324f
C5182 vdd.n2971 gnd 0.007324f
C5183 vdd.n2972 gnd 0.007324f
C5184 vdd.n2973 gnd 0.009099f
C5185 vdd.n2975 gnd 0.009099f
C5186 vdd.n2976 gnd 0.009099f
C5187 vdd.n2977 gnd 0.007324f
C5188 vdd.n2978 gnd 0.007324f
C5189 vdd.n2979 gnd 0.007324f
C5190 vdd.n2980 gnd 0.009099f
C5191 vdd.n2982 gnd 0.009099f
C5192 vdd.n2983 gnd 0.009099f
C5193 vdd.n2984 gnd 0.007324f
C5194 vdd.n2985 gnd 0.009099f
C5195 vdd.n2986 gnd 0.009099f
C5196 vdd.n2987 gnd 0.009099f
C5197 vdd.n2988 gnd 0.015673f
C5198 vdd.n2989 gnd 0.006115f
C5199 vdd.n2990 gnd 0.007324f
C5200 vdd.n2991 gnd 0.009099f
C5201 vdd.n2993 gnd 0.009099f
C5202 vdd.n2994 gnd 0.009099f
C5203 vdd.n2995 gnd 0.007324f
C5204 vdd.n2996 gnd 0.007324f
C5205 vdd.n2997 gnd 0.007324f
C5206 vdd.n2998 gnd 0.009099f
C5207 vdd.n3000 gnd 0.009099f
C5208 vdd.n3001 gnd 0.009099f
C5209 vdd.n3002 gnd 0.007324f
C5210 vdd.n3003 gnd 0.007324f
C5211 vdd.n3004 gnd 0.007324f
C5212 vdd.n3005 gnd 0.009099f
C5213 vdd.n3007 gnd 0.009099f
C5214 vdd.n3008 gnd 0.009099f
C5215 vdd.n3009 gnd 0.007324f
C5216 vdd.n3010 gnd 0.007324f
C5217 vdd.n3011 gnd 0.007324f
C5218 vdd.n3012 gnd 0.009099f
C5219 vdd.n3014 gnd 0.009099f
C5220 vdd.n3015 gnd 0.009099f
C5221 vdd.n3017 gnd 0.009099f
C5222 vdd.n3018 gnd 0.007324f
C5223 vdd.n3019 gnd 0.007324f
C5224 vdd.n3020 gnd 0.006079f
C5225 vdd.n3021 gnd 0.022684f
C5226 vdd.n3022 gnd 0.022175f
C5227 vdd.n3023 gnd 0.006079f
C5228 vdd.n3024 gnd 0.022175f
C5229 vdd.n3025 gnd 1.37157f
C5230 vdd.t43 gnd 0.46494f
C5231 vdd.n3026 gnd 0.488187f
C5232 vdd.n3027 gnd 0.929881f
C5233 vdd.n3028 gnd 0.009099f
C5234 vdd.n3029 gnd 0.007324f
C5235 vdd.n3030 gnd 0.007324f
C5236 vdd.n3031 gnd 0.007324f
C5237 vdd.n3032 gnd 0.009099f
C5238 vdd.n3033 gnd 0.832243f
C5239 vdd.t14 gnd 0.46494f
C5240 vdd.n3034 gnd 0.562578f
C5241 vdd.n3035 gnd 0.674164f
C5242 vdd.n3036 gnd 0.009099f
C5243 vdd.n3037 gnd 0.007324f
C5244 vdd.n3038 gnd 0.007324f
C5245 vdd.n3039 gnd 0.007324f
C5246 vdd.n3040 gnd 0.009099f
C5247 vdd.n3041 gnd 0.516084f
C5248 vdd.t122 gnd 0.46494f
C5249 vdd.n3042 gnd 0.771801f
C5250 vdd.t6 gnd 0.46494f
C5251 vdd.n3043 gnd 0.571877f
C5252 vdd.n3044 gnd 0.009099f
C5253 vdd.n3045 gnd 0.007324f
C5254 vdd.n3046 gnd 0.006993f
C5255 vdd.n3047 gnd 0.536697f
C5256 vdd.n3048 gnd 1.84287f
C5257 a_n1808_13878.t17 gnd 0.185683f
C5258 a_n1808_13878.t15 gnd 0.185683f
C5259 a_n1808_13878.t19 gnd 0.185683f
C5260 a_n1808_13878.n0 gnd 1.46451f
C5261 a_n1808_13878.t8 gnd 0.185683f
C5262 a_n1808_13878.t13 gnd 0.185683f
C5263 a_n1808_13878.n1 gnd 1.46209f
C5264 a_n1808_13878.n2 gnd 1.31424f
C5265 a_n1808_13878.t10 gnd 0.185683f
C5266 a_n1808_13878.t12 gnd 0.185683f
C5267 a_n1808_13878.n3 gnd 1.46364f
C5268 a_n1808_13878.t16 gnd 0.185683f
C5269 a_n1808_13878.t11 gnd 0.185683f
C5270 a_n1808_13878.n4 gnd 1.46209f
C5271 a_n1808_13878.n5 gnd 2.04299f
C5272 a_n1808_13878.t14 gnd 0.185683f
C5273 a_n1808_13878.t9 gnd 0.185683f
C5274 a_n1808_13878.n6 gnd 1.46209f
C5275 a_n1808_13878.n7 gnd 3.70273f
C5276 a_n1808_13878.t7 gnd 1.73864f
C5277 a_n1808_13878.t3 gnd 0.185683f
C5278 a_n1808_13878.t4 gnd 0.185683f
C5279 a_n1808_13878.n8 gnd 1.30795f
C5280 a_n1808_13878.n9 gnd 1.46144f
C5281 a_n1808_13878.t1 gnd 1.73518f
C5282 a_n1808_13878.n10 gnd 0.735417f
C5283 a_n1808_13878.t6 gnd 1.73518f
C5284 a_n1808_13878.n11 gnd 0.735417f
C5285 a_n1808_13878.t2 gnd 0.185683f
C5286 a_n1808_13878.t5 gnd 0.185683f
C5287 a_n1808_13878.n12 gnd 1.30795f
C5288 a_n1808_13878.n13 gnd 0.742539f
C5289 a_n1808_13878.t0 gnd 1.73518f
C5290 a_n1808_13878.n14 gnd 1.73174f
C5291 a_n1808_13878.n15 gnd 2.52099f
C5292 a_n1808_13878.n16 gnd 1.80498f
C5293 a_n1808_13878.n17 gnd 1.46209f
C5294 a_n1808_13878.t18 gnd 0.185683f
C5295 a_n1986_13878.n0 gnd 2.75605f
C5296 a_n1986_13878.n1 gnd 3.98159f
C5297 a_n1986_13878.n2 gnd 3.8498f
C5298 a_n1986_13878.n3 gnd 0.485058f
C5299 a_n1986_13878.n4 gnd 0.654433f
C5300 a_n1986_13878.n5 gnd 0.212692f
C5301 a_n1986_13878.n6 gnd 0.278259f
C5302 a_n1986_13878.n7 gnd 0.629578f
C5303 a_n1986_13878.n8 gnd 0.278259f
C5304 a_n1986_13878.n9 gnd 0.518119f
C5305 a_n1986_13878.n10 gnd 0.20181f
C5306 a_n1986_13878.n11 gnd 0.148637f
C5307 a_n1986_13878.n12 gnd 0.233609f
C5308 a_n1986_13878.n13 gnd 0.180436f
C5309 a_n1986_13878.n14 gnd 0.20181f
C5310 a_n1986_13878.n15 gnd 0.148637f
C5311 a_n1986_13878.n16 gnd 0.571292f
C5312 a_n1986_13878.n17 gnd 0.425782f
C5313 a_n1986_13878.n18 gnd 0.212692f
C5314 a_n1986_13878.n19 gnd 0.485058f
C5315 a_n1986_13878.n20 gnd 0.278259f
C5316 a_n1986_13878.n21 gnd 0.431885f
C5317 a_n1986_13878.n22 gnd 0.212692f
C5318 a_n1986_13878.n23 gnd 0.720523f
C5319 a_n1986_13878.n24 gnd 0.278259f
C5320 a_n1986_13878.n25 gnd 1.75107f
C5321 a_n1986_13878.n26 gnd 1.88685f
C5322 a_n1986_13878.n27 gnd 3.1659f
C5323 a_n1986_13878.n28 gnd 0.008235f
C5324 a_n1986_13878.n30 gnd 0.281365f
C5325 a_n1986_13878.n31 gnd 0.008235f
C5326 a_n1986_13878.n33 gnd 0.281365f
C5327 a_n1986_13878.n34 gnd 0.008235f
C5328 a_n1986_13878.n35 gnd 0.280966f
C5329 a_n1986_13878.n36 gnd 0.008235f
C5330 a_n1986_13878.n37 gnd 0.280966f
C5331 a_n1986_13878.n38 gnd 0.008235f
C5332 a_n1986_13878.n39 gnd 0.280966f
C5333 a_n1986_13878.n40 gnd 0.008235f
C5334 a_n1986_13878.n41 gnd 1.3183f
C5335 a_n1986_13878.n42 gnd 0.280966f
C5336 a_n1986_13878.n43 gnd 0.106346f
C5337 a_n1986_13878.n44 gnd 0.008235f
C5338 a_n1986_13878.n46 gnd 0.008235f
C5339 a_n1986_13878.n48 gnd 0.281365f
C5340 a_n1986_13878.n49 gnd 0.281365f
C5341 a_n1986_13878.t24 gnd 0.686217f
C5342 a_n1986_13878.n50 gnd 0.301704f
C5343 a_n1986_13878.t20 gnd 0.686217f
C5344 a_n1986_13878.t34 gnd 0.686217f
C5345 a_n1986_13878.t47 gnd 0.686217f
C5346 a_n1986_13878.n51 gnd 0.301704f
C5347 a_n1986_13878.t56 gnd 0.686217f
C5348 a_n1986_13878.t61 gnd 0.686217f
C5349 a_n1986_13878.t28 gnd 0.700669f
C5350 a_n1986_13878.t18 gnd 0.686217f
C5351 a_n1986_13878.t38 gnd 0.686217f
C5352 a_n1986_13878.t30 gnd 0.686217f
C5353 a_n1986_13878.n52 gnd 0.301704f
C5354 a_n1986_13878.t26 gnd 0.686217f
C5355 a_n1986_13878.t36 gnd 0.697562f
C5356 a_n1986_13878.t9 gnd 0.114742f
C5357 a_n1986_13878.t3 gnd 0.114742f
C5358 a_n1986_13878.n53 gnd 1.01689f
C5359 a_n1986_13878.t11 gnd 0.114742f
C5360 a_n1986_13878.t1 gnd 0.114742f
C5361 a_n1986_13878.n54 gnd 1.0139f
C5362 a_n1986_13878.t8 gnd 0.114742f
C5363 a_n1986_13878.t7 gnd 0.114742f
C5364 a_n1986_13878.n55 gnd 1.01689f
C5365 a_n1986_13878.t6 gnd 0.114742f
C5366 a_n1986_13878.t14 gnd 0.114742f
C5367 a_n1986_13878.n56 gnd 1.0139f
C5368 a_n1986_13878.t12 gnd 0.114742f
C5369 a_n1986_13878.t5 gnd 0.114742f
C5370 a_n1986_13878.n57 gnd 1.0139f
C5371 a_n1986_13878.t4 gnd 0.114742f
C5372 a_n1986_13878.t0 gnd 0.114742f
C5373 a_n1986_13878.n58 gnd 1.0139f
C5374 a_n1986_13878.t15 gnd 0.114742f
C5375 a_n1986_13878.t13 gnd 0.114742f
C5376 a_n1986_13878.n59 gnd 1.01689f
C5377 a_n1986_13878.t10 gnd 0.114742f
C5378 a_n1986_13878.t2 gnd 0.114742f
C5379 a_n1986_13878.n60 gnd 1.0139f
C5380 a_n1986_13878.t66 gnd 0.700669f
C5381 a_n1986_13878.t49 gnd 0.686217f
C5382 a_n1986_13878.t53 gnd 0.686217f
C5383 a_n1986_13878.t43 gnd 0.686217f
C5384 a_n1986_13878.n61 gnd 0.301704f
C5385 a_n1986_13878.t58 gnd 0.686217f
C5386 a_n1986_13878.t64 gnd 0.697562f
C5387 a_n1986_13878.n62 gnd 0.304282f
C5388 a_n1986_13878.n63 gnd 0.297873f
C5389 a_n1986_13878.n64 gnd 0.304282f
C5390 a_n1986_13878.n65 gnd 0.304282f
C5391 a_n1986_13878.n66 gnd 0.297873f
C5392 a_n1986_13878.n67 gnd 0.304282f
C5393 a_n1986_13878.t37 gnd 1.38135f
C5394 a_n1986_13878.t31 gnd 0.147525f
C5395 a_n1986_13878.t27 gnd 0.147525f
C5396 a_n1986_13878.n68 gnd 1.03917f
C5397 a_n1986_13878.t19 gnd 0.147525f
C5398 a_n1986_13878.t39 gnd 0.147525f
C5399 a_n1986_13878.n69 gnd 1.03917f
C5400 a_n1986_13878.t29 gnd 1.3786f
C5401 a_n1986_13878.n70 gnd 1.12735f
C5402 a_n1986_13878.n71 gnd 0.775089f
C5403 a_n1986_13878.t48 gnd 0.686217f
C5404 a_n1986_13878.t57 gnd 0.686217f
C5405 a_n1986_13878.t67 gnd 0.686217f
C5406 a_n1986_13878.n72 gnd 0.301704f
C5407 a_n1986_13878.t59 gnd 0.686217f
C5408 a_n1986_13878.t45 gnd 0.686217f
C5409 a_n1986_13878.t44 gnd 0.686217f
C5410 a_n1986_13878.n73 gnd 0.301704f
C5411 a_n1986_13878.t63 gnd 0.686217f
C5412 a_n1986_13878.t52 gnd 0.686217f
C5413 a_n1986_13878.t51 gnd 0.686217f
C5414 a_n1986_13878.n74 gnd 0.301704f
C5415 a_n1986_13878.t55 gnd 0.686217f
C5416 a_n1986_13878.t46 gnd 0.686217f
C5417 a_n1986_13878.t40 gnd 0.686217f
C5418 a_n1986_13878.n75 gnd 0.301704f
C5419 a_n1986_13878.t60 gnd 0.697715f
C5420 a_n1986_13878.n76 gnd 0.297873f
C5421 a_n1986_13878.n77 gnd 0.292464f
C5422 a_n1986_13878.t65 gnd 0.697715f
C5423 a_n1986_13878.n78 gnd 0.297873f
C5424 a_n1986_13878.n79 gnd 0.292464f
C5425 a_n1986_13878.t54 gnd 0.697715f
C5426 a_n1986_13878.n80 gnd 0.297873f
C5427 a_n1986_13878.n81 gnd 0.292464f
C5428 a_n1986_13878.t50 gnd 0.697715f
C5429 a_n1986_13878.n82 gnd 0.297873f
C5430 a_n1986_13878.n83 gnd 0.292464f
C5431 a_n1986_13878.n84 gnd 0.991153f
C5432 a_n1986_13878.t62 gnd 0.700669f
C5433 a_n1986_13878.n85 gnd 0.304282f
C5434 a_n1986_13878.t41 gnd 0.686217f
C5435 a_n1986_13878.n86 gnd 0.297873f
C5436 a_n1986_13878.n87 gnd 0.304282f
C5437 a_n1986_13878.t42 gnd 0.697562f
C5438 a_n1986_13878.t16 gnd 0.700669f
C5439 a_n1986_13878.n88 gnd 0.304282f
C5440 a_n1986_13878.t22 gnd 0.686217f
C5441 a_n1986_13878.n89 gnd 0.297873f
C5442 a_n1986_13878.n90 gnd 0.304282f
C5443 a_n1986_13878.t32 gnd 0.697562f
C5444 a_n1986_13878.n91 gnd 1.115f
C5445 a_n1986_13878.t33 gnd 1.3786f
C5446 a_n1986_13878.t25 gnd 0.147525f
C5447 a_n1986_13878.t21 gnd 0.147525f
C5448 a_n1986_13878.n92 gnd 1.03917f
C5449 a_n1986_13878.t35 gnd 0.147525f
C5450 a_n1986_13878.t23 gnd 0.147525f
C5451 a_n1986_13878.n93 gnd 1.03917f
C5452 a_n1986_13878.n94 gnd 1.16112f
C5453 a_n1986_13878.t17 gnd 1.38135f
.ends

