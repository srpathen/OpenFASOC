* NGSPICE file created from opamp112.ext - technology: sky130A

.subckt opamp112 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n8964_8799.t42 plus.t5 a_n3827_n3924.t31 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X1 a_n2804_13878.t31 a_n2982_13878.t72 vdd.t55 vdd.t54 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 a_n2804_13878.t23 a_n2982_13878.t29 a_n2982_13878.t30 vdd.t42 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 gnd.t286 gnd.t284 gnd.t285 gnd.t244 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X4 vdd.t183 a_n8964_8799.t48 CSoutput.t105 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X5 gnd.t283 gnd.t281 minus.t4 gnd.t282 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X6 CSoutput.t104 a_n8964_8799.t49 vdd.t182 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X7 gnd.t113 commonsourceibias.t64 CSoutput.t130 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 a_n3827_n3924.t6 diffpairibias.t20 gnd.t30 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X9 a_n3827_n3924.t43 plus.t6 a_n8964_8799.t41 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X10 commonsourceibias.t63 commonsourceibias.t62 gnd.t163 gnd.t118 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 gnd.t280 gnd.t278 gnd.t279 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X12 vdd.t181 a_n8964_8799.t50 CSoutput.t103 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X13 a_n3827_n3924.t9 minus.t5 a_n2982_13878.t53 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X14 vdd.t194 CSoutput.t160 output.t18 gnd.t147 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X15 a_n2982_8322.t23 a_n2982_13878.t73 a_n8964_8799.t4 vdd.t52 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X16 gnd.t277 gnd.t275 gnd.t276 gnd.t195 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X17 CSoutput.t131 commonsourceibias.t65 gnd.t115 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 CSoutput.t102 a_n8964_8799.t51 vdd.t176 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X19 vdd.t180 a_n8964_8799.t52 CSoutput.t101 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X20 CSoutput.t100 a_n8964_8799.t53 vdd.t179 vdd.t95 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 gnd.t168 commonsourceibias.t60 commonsourceibias.t61 gnd.t72 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X22 CSoutput.t150 commonsourceibias.t66 gnd.t162 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 vdd.t178 a_n8964_8799.t54 CSoutput.t99 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X24 vdd.t177 a_n8964_8799.t55 CSoutput.t98 vdd.t121 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X25 gnd.t274 gnd.t272 gnd.t273 gnd.t195 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X26 a_n2982_13878.t4 minus.t6 a_n3827_n3924.t5 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X27 commonsourceibias.t59 commonsourceibias.t58 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 a_n8964_8799.t18 a_n2982_13878.t74 a_n2982_8322.t22 vdd.t38 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X29 CSoutput.t117 commonsourceibias.t67 gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X30 vdd.t175 a_n8964_8799.t56 CSoutput.t97 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X31 a_n2982_13878.t68 minus.t7 a_n3827_n3924.t52 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X32 vdd.t174 a_n8964_8799.t57 CSoutput.t96 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X33 a_n8964_8799.t44 a_n2982_13878.t75 a_n2982_8322.t21 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X34 commonsourceibias.t57 commonsourceibias.t56 gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 a_n3827_n3924.t22 minus.t8 a_n2982_13878.t64 gnd.t151 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X36 gnd.t271 gnd.t269 gnd.t270 gnd.t187 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X37 CSoutput.t161 a_n2982_8322.t37 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X38 CSoutput.t120 commonsourceibias.t68 gnd.t77 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X39 a_n3827_n3924.t57 diffpairibias.t21 gnd.t331 gnd.t330 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X40 CSoutput.t95 a_n8964_8799.t58 vdd.t173 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X41 gnd.t268 gnd.t265 gnd.t267 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X42 gnd.t320 commonsourceibias.t69 CSoutput.t159 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 vdd.t172 a_n8964_8799.t59 CSoutput.t94 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X44 gnd.t169 commonsourceibias.t54 commonsourceibias.t55 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X45 output.t17 CSoutput.t162 vdd.t195 gnd.t148 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X46 commonsourceibias.t53 commonsourceibias.t52 gnd.t164 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X47 a_n3827_n3924.t42 plus.t7 a_n8964_8799.t40 gnd.t108 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X48 vdd.t171 a_n8964_8799.t60 CSoutput.t93 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X49 gnd.t112 commonsourceibias.t70 CSoutput.t129 gnd.t74 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X50 a_n2804_13878.t22 a_n2982_13878.t15 a_n2982_13878.t16 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X51 a_n8964_8799.t39 plus.t8 a_n3827_n3924.t45 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X52 a_n2982_13878.t8 a_n2982_13878.t7 a_n2804_13878.t21 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X53 CSoutput.t163 a_n2982_8322.t36 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X54 gnd.t44 commonsourceibias.t71 CSoutput.t108 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 a_n8964_8799.t38 plus.t9 a_n3827_n3924.t41 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X56 CSoutput.t92 a_n8964_8799.t61 vdd.t170 vdd.t95 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X57 output.t16 CSoutput.t164 vdd.t189 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X58 vdd.t271 vdd.t269 vdd.t270 vdd.t246 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X59 vdd.t169 a_n8964_8799.t62 CSoutput.t91 vdd.t121 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X60 vdd.t168 a_n8964_8799.t63 CSoutput.t90 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 gnd.t78 commonsourceibias.t50 commonsourceibias.t51 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X62 diffpairibias.t19 diffpairibias.t18 gnd.t154 gnd.t153 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X63 a_n3827_n3924.t33 plus.t10 a_n8964_8799.t37 gnd.t104 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X64 commonsourceibias.t49 commonsourceibias.t48 gnd.t135 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X65 a_n2982_13878.t60 minus.t9 a_n3827_n3924.t18 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X66 a_n2982_13878.t40 a_n2982_13878.t39 a_n2804_13878.t20 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X67 CSoutput.t89 a_n8964_8799.t64 vdd.t166 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X68 vdd.t165 a_n8964_8799.t65 CSoutput.t88 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X69 a_n8964_8799.t14 a_n2982_13878.t76 a_n2982_8322.t20 vdd.t34 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X70 CSoutput.t87 a_n8964_8799.t66 vdd.t164 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 commonsourceibias.t47 commonsourceibias.t46 gnd.t129 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X72 gnd.t264 gnd.t262 plus.t4 gnd.t263 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X73 a_n2982_13878.t12 a_n2982_13878.t11 a_n2804_13878.t19 vdd.t53 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X74 vdd.t163 a_n8964_8799.t67 CSoutput.t86 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X75 vdd.t162 a_n8964_8799.t68 CSoutput.t85 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X76 a_n8964_8799.t9 a_n2982_13878.t77 a_n2982_8322.t19 vdd.t32 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X77 gnd.t261 gnd.t259 gnd.t260 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X78 diffpairibias.t17 diffpairibias.t16 gnd.t309 gnd.t308 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X79 gnd.t165 commonsourceibias.t44 commonsourceibias.t45 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 CSoutput.t84 a_n8964_8799.t69 vdd.t161 vdd.t75 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 a_n8964_8799.t0 a_n2982_13878.t78 a_n2982_8322.t18 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X82 CSoutput.t134 commonsourceibias.t72 gnd.t123 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X83 output.t2 outputibias.t8 gnd.t150 gnd.t149 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X84 a_n2982_8322.t17 a_n2982_13878.t79 a_n8964_8799.t43 vdd.t53 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X85 CSoutput.t83 a_n8964_8799.t70 vdd.t160 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 vdd.t190 CSoutput.t165 output.t15 gnd.t89 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X87 vdd.t186 CSoutput.t166 output.t14 gnd.t79 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X88 gnd.t289 commonsourceibias.t42 commonsourceibias.t43 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 CSoutput.t135 commonsourceibias.t73 gnd.t124 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 CSoutput.t153 commonsourceibias.t74 gnd.t177 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 gnd.t258 gnd.t256 gnd.t257 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X92 gnd.t255 gnd.t253 plus.t3 gnd.t254 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X93 a_n3827_n3924.t35 plus.t11 a_n8964_8799.t36 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X94 CSoutput.t128 commonsourceibias.t75 gnd.t102 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X95 outputibias.t7 outputibias.t6 gnd.t111 gnd.t110 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X96 CSoutput.t149 commonsourceibias.t76 gnd.t161 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X97 vdd.t268 vdd.t266 vdd.t267 vdd.t242 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X98 a_n3827_n3924.t13 diffpairibias.t22 gnd.t85 gnd.t84 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X99 vdd.t159 a_n8964_8799.t71 CSoutput.t82 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X100 vdd.t158 a_n8964_8799.t72 CSoutput.t81 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X101 a_n2982_13878.t18 a_n2982_13878.t17 a_n2804_13878.t18 vdd.t52 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X102 vdd.t157 a_n8964_8799.t73 CSoutput.t80 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X103 a_n8964_8799.t47 a_n2982_13878.t80 a_n2982_8322.t16 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X104 a_n2982_13878.t28 a_n2982_13878.t27 a_n2804_13878.t17 vdd.t6 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X105 gnd.t130 commonsourceibias.t40 commonsourceibias.t41 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X106 gnd.t132 commonsourceibias.t38 commonsourceibias.t39 gnd.t131 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X107 CSoutput.t79 a_n8964_8799.t74 vdd.t156 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X108 diffpairibias.t15 diffpairibias.t14 gnd.t288 gnd.t287 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X109 a_n2982_13878.t71 minus.t10 a_n3827_n3924.t55 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X110 vdd.t265 vdd.t263 vdd.t264 vdd.t253 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X111 CSoutput.t78 a_n8964_8799.t75 vdd.t155 vdd.t75 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X112 gnd.t304 commonsourceibias.t77 CSoutput.t157 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X113 vdd.t262 vdd.t259 vdd.t261 vdd.t260 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X114 gnd.t20 commonsourceibias.t78 CSoutput.t5 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X115 gnd.t142 commonsourceibias.t79 CSoutput.t140 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X116 gnd.t75 commonsourceibias.t80 CSoutput.t119 gnd.t74 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 a_n2804_13878.t16 a_n2982_13878.t5 a_n2982_13878.t6 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X118 a_n3827_n3924.t53 minus.t11 a_n2982_13878.t69 gnd.t171 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X119 CSoutput.t77 a_n8964_8799.t76 vdd.t154 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X120 output.t13 CSoutput.t167 vdd.t187 gnd.t80 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X121 vdd.t153 a_n8964_8799.t77 CSoutput.t76 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X122 vdd.t188 CSoutput.t168 output.t12 gnd.t81 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X123 vdd.t51 a_n2982_13878.t81 a_n2982_8322.t31 vdd.t50 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X124 a_n2982_13878.t24 a_n2982_13878.t23 a_n2804_13878.t15 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X125 gnd.t160 commonsourceibias.t81 CSoutput.t148 gnd.t72 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X126 gnd.t252 gnd.t250 gnd.t251 gnd.t214 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X127 a_n2982_8322.t30 a_n2982_13878.t82 vdd.t49 vdd.t48 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X128 a_n3827_n3924.t8 diffpairibias.t23 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X129 CSoutput.t75 a_n8964_8799.t78 vdd.t152 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X130 a_n3827_n3924.t4 minus.t12 a_n2982_13878.t3 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X131 a_n3827_n3924.t1 minus.t13 a_n2982_13878.t0 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X132 vdd.t47 a_n2982_13878.t83 a_n2804_13878.t30 vdd.t46 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X133 a_n2982_13878.t1 minus.t14 a_n3827_n3924.t2 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X134 vdd.t258 vdd.t256 vdd.t257 vdd.t242 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X135 a_n3827_n3924.t37 plus.t12 a_n8964_8799.t35 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X136 a_n3827_n3924.t48 plus.t13 a_n8964_8799.t34 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X137 gnd.t101 commonsourceibias.t82 CSoutput.t127 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 vdd.t255 vdd.t252 vdd.t254 vdd.t253 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X139 a_n2982_13878.t63 minus.t15 a_n3827_n3924.t21 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X140 a_n2804_13878.t14 a_n2982_13878.t47 a_n2982_13878.t48 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X141 vdd.t151 a_n8964_8799.t79 CSoutput.t74 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X142 vdd.t149 a_n8964_8799.t80 CSoutput.t73 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X143 a_n2982_8322.t15 a_n2982_13878.t84 a_n8964_8799.t12 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X144 gnd.t249 gnd.t247 plus.t2 gnd.t248 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X145 a_n8964_8799.t33 plus.t14 a_n3827_n3924.t38 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X146 a_n8964_8799.t32 plus.t15 a_n3827_n3924.t29 gnd.t166 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X147 vdd.t251 vdd.t249 vdd.t250 vdd.t219 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X148 vdd.t248 vdd.t245 vdd.t247 vdd.t246 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X149 a_n2982_8322.t29 a_n2982_13878.t85 vdd.t44 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X150 a_n8964_8799.t46 a_n2982_13878.t86 a_n2982_8322.t14 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X151 CSoutput.t72 a_n8964_8799.t81 vdd.t148 vdd.t86 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X152 diffpairibias.t13 diffpairibias.t12 gnd.t126 gnd.t125 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X153 vdd.t147 a_n8964_8799.t82 CSoutput.t71 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X154 a_n2982_13878.t61 minus.t16 a_n3827_n3924.t19 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X155 a_n2982_13878.t34 a_n2982_13878.t33 a_n2804_13878.t13 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X156 a_n8964_8799.t8 a_n2982_13878.t87 a_n2982_8322.t13 vdd.t42 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X157 CSoutput.t70 a_n8964_8799.t83 vdd.t145 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X158 CSoutput.t69 a_n8964_8799.t84 vdd.t143 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 CSoutput.t116 commonsourceibias.t83 gnd.t59 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X160 commonsourceibias.t37 commonsourceibias.t36 gnd.t133 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 CSoutput.t115 commonsourceibias.t84 gnd.t57 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X162 a_n2804_13878.t12 a_n2982_13878.t37 a_n2982_13878.t38 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X163 a_n3827_n3924.t54 minus.t17 a_n2982_13878.t70 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X164 CSoutput.t4 commonsourceibias.t85 gnd.t18 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X165 vdd.t184 CSoutput.t169 output.t11 gnd.t65 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X166 vdd.t244 vdd.t241 vdd.t243 vdd.t242 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X167 vdd.t240 vdd.t238 vdd.t239 vdd.t215 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X168 CSoutput.t7 commonsourceibias.t86 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 vdd.t237 vdd.t235 vdd.t236 vdd.t201 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X170 gnd.t4 commonsourceibias.t87 CSoutput.t0 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X171 CSoutput.t68 a_n8964_8799.t85 vdd.t142 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X172 gnd.t290 commonsourceibias.t34 commonsourceibias.t35 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X173 gnd.t246 gnd.t243 gnd.t245 gnd.t244 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X174 vdd.t40 a_n2982_13878.t88 a_n2982_8322.t28 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X175 a_n2804_13878.t11 a_n2982_13878.t19 a_n2982_13878.t20 vdd.t38 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X176 vdd.t135 a_n8964_8799.t86 CSoutput.t67 vdd.t123 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X177 vdd.t141 a_n8964_8799.t87 CSoutput.t66 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X178 commonsourceibias.t33 commonsourceibias.t32 gnd.t321 gnd.t49 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X179 a_n2982_13878.t26 a_n2982_13878.t25 a_n2804_13878.t10 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X180 gnd.t296 commonsourceibias.t30 commonsourceibias.t31 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X181 minus.t3 gnd.t240 gnd.t242 gnd.t241 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X182 a_n3827_n3924.t47 plus.t16 a_n8964_8799.t31 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X183 vdd.t140 a_n8964_8799.t88 CSoutput.t65 vdd.t81 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X184 gnd.t325 commonsourceibias.t28 commonsourceibias.t29 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X185 a_n3827_n3924.t49 diffpairibias.t24 gnd.t294 gnd.t293 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X186 commonsourceibias.t27 commonsourceibias.t26 gnd.t295 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 a_n3827_n3924.t7 diffpairibias.t25 gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X188 outputibias.t5 outputibias.t4 gnd.t106 gnd.t105 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X189 gnd.t34 commonsourceibias.t88 CSoutput.t9 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X190 vdd.t139 a_n8964_8799.t89 CSoutput.t64 vdd.t123 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X191 vdd.t138 a_n8964_8799.t90 CSoutput.t63 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X192 a_n8964_8799.t30 plus.t17 a_n3827_n3924.t36 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X193 gnd.t303 commonsourceibias.t89 CSoutput.t156 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 CSoutput.t62 a_n8964_8799.t91 vdd.t137 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X195 gnd.t16 commonsourceibias.t90 CSoutput.t3 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 gnd.t141 commonsourceibias.t91 CSoutput.t139 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X197 vdd.t234 vdd.t232 vdd.t233 vdd.t219 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X198 gnd.t73 commonsourceibias.t92 CSoutput.t118 gnd.t72 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X199 a_n2804_13878.t9 a_n2982_13878.t9 a_n2982_13878.t10 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X200 a_n2982_8322.t12 a_n2982_13878.t89 a_n8964_8799.t16 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X201 CSoutput.t61 a_n8964_8799.t92 vdd.t136 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X202 CSoutput.t60 a_n8964_8799.t93 vdd.t134 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X203 commonsourceibias.t25 commonsourceibias.t24 gnd.t322 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X204 outputibias.t3 outputibias.t2 gnd.t307 gnd.t306 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X205 gnd.t28 commonsourceibias.t93 CSoutput.t8 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X206 CSoutput.t154 commonsourceibias.t94 gnd.t178 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 diffpairibias.t11 diffpairibias.t10 gnd.t8 gnd.t7 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X208 a_n2804_13878.t29 a_n2982_13878.t90 vdd.t5 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X209 gnd.t43 commonsourceibias.t95 CSoutput.t107 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 vdd.t36 a_n2982_13878.t91 a_n2804_13878.t28 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X211 gnd.t297 commonsourceibias.t22 commonsourceibias.t23 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 CSoutput.t59 a_n8964_8799.t94 vdd.t133 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X213 vdd.t124 a_n8964_8799.t95 CSoutput.t58 vdd.t123 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X214 vdd.t131 a_n8964_8799.t96 CSoutput.t57 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X215 commonsourceibias.t21 commonsourceibias.t20 gnd.t326 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X216 vdd.t129 a_n8964_8799.t97 CSoutput.t56 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 CSoutput.t142 commonsourceibias.t96 gnd.t146 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 CSoutput.t55 a_n8964_8799.t98 vdd.t125 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X219 plus.t1 gnd.t237 gnd.t239 gnd.t238 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X220 a_n2804_13878.t8 a_n2982_13878.t13 a_n2982_13878.t14 vdd.t34 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X221 diffpairibias.t9 diffpairibias.t8 gnd.t292 gnd.t291 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X222 a_n3827_n3924.t17 minus.t18 a_n2982_13878.t59 gnd.t108 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X223 vdd.t127 a_n8964_8799.t99 CSoutput.t54 vdd.t81 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X224 gnd.t327 commonsourceibias.t18 commonsourceibias.t19 gnd.t74 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X225 CSoutput.t141 commonsourceibias.t97 gnd.t145 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X226 a_n2982_13878.t67 minus.t19 a_n3827_n3924.t51 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X227 a_n2982_8322.t11 a_n2982_13878.t92 a_n8964_8799.t10 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X228 a_n2982_13878.t52 a_n2982_13878.t51 a_n2804_13878.t7 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X229 CSoutput.t53 a_n8964_8799.t100 vdd.t126 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X230 diffpairibias.t7 diffpairibias.t6 gnd.t324 gnd.t323 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X231 vdd.t122 a_n8964_8799.t101 CSoutput.t52 vdd.t121 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X232 a_n2804_13878.t6 a_n2982_13878.t31 a_n2982_13878.t32 vdd.t32 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X233 a_n2982_13878.t56 minus.t20 a_n3827_n3924.t12 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X234 a_n2982_13878.t58 minus.t21 a_n3827_n3924.t16 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X235 vdd.t31 a_n2982_13878.t93 a_n2982_8322.t27 vdd.t30 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X236 vdd.t120 a_n8964_8799.t102 CSoutput.t51 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X237 a_n3827_n3924.t15 minus.t22 a_n2982_13878.t57 gnd.t104 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X238 vdd.t185 CSoutput.t170 output.t10 gnd.t66 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X239 CSoutput.t171 a_n2982_8322.t35 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X240 CSoutput.t151 commonsourceibias.t98 gnd.t167 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X241 a_n8964_8799.t29 plus.t18 a_n3827_n3924.t27 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X242 CSoutput.t106 commonsourceibias.t99 gnd.t41 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 gnd.t302 commonsourceibias.t100 CSoutput.t155 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X244 a_n3827_n3924.t11 minus.t23 a_n2982_13878.t55 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X245 CSoutput.t50 a_n8964_8799.t103 vdd.t118 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X246 gnd.t236 gnd.t233 gnd.t235 gnd.t234 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X247 a_n2804_13878.t27 a_n2982_13878.t94 vdd.t29 vdd.t28 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X248 outputibias.t1 outputibias.t0 gnd.t87 gnd.t86 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X249 vdd.t231 vdd.t229 vdd.t230 vdd.t215 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X250 CSoutput.t158 commonsourceibias.t101 gnd.t314 gnd.t118 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X251 commonsourceibias.t17 commonsourceibias.t16 gnd.t328 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X252 vdd.t117 a_n8964_8799.t104 CSoutput.t49 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X253 CSoutput.t48 a_n8964_8799.t105 vdd.t115 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X254 CSoutput.t172 a_n2982_8322.t34 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X255 CSoutput.t47 a_n8964_8799.t106 vdd.t113 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X256 gnd.t232 gnd.t230 minus.t2 gnd.t231 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X257 gnd.t229 gnd.t227 gnd.t228 gnd.t214 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X258 gnd.t226 gnd.t223 gnd.t225 gnd.t224 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X259 vdd.t228 vdd.t226 vdd.t227 vdd.t205 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X260 vdd.t98 a_n8964_8799.t107 CSoutput.t46 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X261 a_n3827_n3924.t0 diffpairibias.t26 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X262 vdd.t27 a_n2982_13878.t95 a_n2982_8322.t26 vdd.t26 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X263 a_n2982_8322.t10 a_n2982_13878.t96 a_n8964_8799.t5 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X264 gnd.t140 commonsourceibias.t102 CSoutput.t138 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X265 vdd.t112 a_n8964_8799.t108 CSoutput.t45 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X266 a_n8964_8799.t28 plus.t19 a_n3827_n3924.t46 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X267 output.t1 outputibias.t9 gnd.t83 gnd.t82 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X268 gnd.t100 commonsourceibias.t103 CSoutput.t126 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 CSoutput.t125 commonsourceibias.t104 gnd.t99 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X270 vdd.t225 vdd.t222 vdd.t224 vdd.t223 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X271 a_n3827_n3924.t25 plus.t20 a_n8964_8799.t27 gnd.t151 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X272 vdd.t111 a_n8964_8799.t109 CSoutput.t44 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 CSoutput.t43 a_n8964_8799.t110 vdd.t110 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X274 gnd.t55 commonsourceibias.t105 CSoutput.t114 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 a_n2804_13878.t5 a_n2982_13878.t45 a_n2982_13878.t46 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X276 CSoutput.t42 a_n8964_8799.t111 vdd.t108 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X277 CSoutput.t41 a_n8964_8799.t112 vdd.t107 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X278 CSoutput.t136 commonsourceibias.t106 gnd.t128 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X279 a_n2982_8322.t9 a_n2982_13878.t97 a_n8964_8799.t17 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X280 diffpairibias.t5 diffpairibias.t4 gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X281 commonsourceibias.t15 commonsourceibias.t14 gnd.t329 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X282 gnd.t134 commonsourceibias.t107 CSoutput.t137 gnd.t131 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X283 gnd.t222 gnd.t220 gnd.t221 gnd.t187 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X284 CSoutput.t147 commonsourceibias.t108 gnd.t159 gnd.t49 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X285 gnd.t122 commonsourceibias.t12 commonsourceibias.t13 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 CSoutput.t40 a_n8964_8799.t113 vdd.t106 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X287 CSoutput.t39 a_n8964_8799.t114 vdd.t104 vdd.t86 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 a_n3827_n3924.t14 diffpairibias.t27 gnd.t91 gnd.t90 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X289 vdd.t221 vdd.t218 vdd.t220 vdd.t219 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X290 vdd.t217 vdd.t214 vdd.t216 vdd.t215 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X291 CSoutput.t146 commonsourceibias.t109 gnd.t158 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 a_n2982_8322.t25 a_n2982_13878.t98 vdd.t23 vdd.t22 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X293 CSoutput.t38 a_n8964_8799.t115 vdd.t103 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X294 CSoutput.t124 commonsourceibias.t110 gnd.t97 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X295 vdd.t101 a_n8964_8799.t116 CSoutput.t37 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X296 CSoutput.t36 a_n8964_8799.t117 vdd.t100 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X297 vdd.t21 a_n2982_13878.t99 a_n2804_13878.t26 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X298 gnd.t116 commonsourceibias.t10 commonsourceibias.t11 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X299 plus.t0 gnd.t217 gnd.t219 gnd.t218 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X300 vdd.t99 a_n8964_8799.t118 CSoutput.t35 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 CSoutput.t34 a_n8964_8799.t119 vdd.t96 vdd.t95 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X302 output.t9 CSoutput.t173 vdd.t272 gnd.t300 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X303 CSoutput.t113 commonsourceibias.t111 gnd.t54 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X304 gnd.t52 commonsourceibias.t112 CSoutput.t112 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X305 vdd.t94 a_n8964_8799.t120 CSoutput.t33 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X306 a_n3827_n3924.t26 plus.t21 a_n8964_8799.t26 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X307 CSoutput.t2 commonsourceibias.t113 gnd.t14 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X308 commonsourceibias.t9 commonsourceibias.t8 gnd.t117 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X309 a_n3827_n3924.t23 minus.t24 a_n2982_13878.t65 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X310 a_n2982_8322.t8 a_n2982_13878.t100 a_n8964_8799.t2 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X311 CSoutput.t132 commonsourceibias.t114 gnd.t119 gnd.t118 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X312 a_n8964_8799.t13 a_n2982_13878.t101 a_n2982_8322.t7 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X313 output.t8 CSoutput.t174 vdd.t273 gnd.t301 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X314 gnd.t143 commonsourceibias.t6 commonsourceibias.t7 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 a_n8964_8799.t25 plus.t22 a_n3827_n3924.t34 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X316 a_n2804_13878.t25 a_n2982_13878.t102 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X317 gnd.t120 commonsourceibias.t115 CSoutput.t133 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X318 vdd.t213 vdd.t211 vdd.t212 vdd.t197 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X319 vdd.t78 a_n8964_8799.t121 CSoutput.t32 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X320 a_n2982_13878.t54 minus.t25 a_n3827_n3924.t10 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X321 CSoutput.t31 a_n8964_8799.t122 vdd.t92 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 CSoutput.t30 a_n8964_8799.t123 vdd.t90 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X323 CSoutput.t29 a_n8964_8799.t124 vdd.t88 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X324 a_n2982_13878.t42 a_n2982_13878.t41 a_n2804_13878.t4 vdd.t7 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X325 gnd.t216 gnd.t213 gnd.t215 gnd.t214 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X326 a_n8964_8799.t11 a_n2982_13878.t103 a_n2982_8322.t6 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X327 commonsourceibias.t5 commonsourceibias.t4 gnd.t315 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X328 a_n8964_8799.t15 a_n2982_13878.t104 a_n2982_8322.t5 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X329 a_n8964_8799.t24 plus.t23 a_n3827_n3924.t28 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X330 gnd.t212 gnd.t209 gnd.t211 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X331 gnd.t208 gnd.t206 minus.t1 gnd.t207 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X332 a_n2982_8322.t4 a_n2982_13878.t105 a_n8964_8799.t1 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X333 CSoutput.t175 a_n2982_8322.t33 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X334 a_n3827_n3924.t20 minus.t26 a_n2982_13878.t62 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X335 vdd.t82 a_n8964_8799.t125 CSoutput.t28 vdd.t81 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X336 CSoutput.t27 a_n8964_8799.t126 vdd.t87 vdd.t86 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X337 CSoutput.t26 a_n8964_8799.t127 vdd.t85 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X338 gnd.t305 commonsourceibias.t2 commonsourceibias.t3 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X339 CSoutput.t25 a_n8964_8799.t128 vdd.t77 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 a_n2804_13878.t3 a_n2982_13878.t43 a_n2982_13878.t44 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X341 a_n3827_n3924.t30 plus.t24 a_n8964_8799.t23 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X342 vdd.t84 a_n8964_8799.t129 CSoutput.t24 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X343 gnd.t22 commonsourceibias.t116 CSoutput.t6 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X344 CSoutput.t152 commonsourceibias.t117 gnd.t176 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X345 output.t7 CSoutput.t176 vdd.t274 gnd.t312 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X346 gnd.t95 commonsourceibias.t118 CSoutput.t123 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X347 a_n3827_n3924.t56 diffpairibias.t28 gnd.t311 gnd.t310 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X348 vdd.t83 a_n8964_8799.t130 CSoutput.t23 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X349 gnd.t205 gnd.t202 gnd.t204 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X350 CSoutput.t22 a_n8964_8799.t131 vdd.t80 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X351 gnd.t201 gnd.t198 gnd.t200 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X352 a_n2982_13878.t36 a_n2982_13878.t35 a_n2804_13878.t2 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X353 gnd.t197 gnd.t194 gnd.t196 gnd.t195 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X354 a_n8964_8799.t3 a_n2982_13878.t106 a_n2982_8322.t3 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X355 output.t19 outputibias.t10 gnd.t319 gnd.t318 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X356 vdd.t79 a_n8964_8799.t132 CSoutput.t21 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X357 gnd.t157 commonsourceibias.t119 CSoutput.t145 gnd.t131 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X358 CSoutput.t20 a_n8964_8799.t133 vdd.t76 vdd.t75 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X359 a_n8964_8799.t22 plus.t25 a_n3827_n3924.t40 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X360 vdd.t210 vdd.t208 vdd.t209 vdd.t205 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X361 vdd.t275 CSoutput.t177 output.t6 gnd.t313 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X362 gnd.t193 gnd.t190 gnd.t192 gnd.t191 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X363 CSoutput.t122 commonsourceibias.t120 gnd.t93 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X364 CSoutput.t111 commonsourceibias.t121 gnd.t50 gnd.t49 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X365 diffpairibias.t3 diffpairibias.t2 gnd.t317 gnd.t316 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X366 CSoutput.t19 a_n8964_8799.t134 vdd.t74 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X367 output.t0 outputibias.t11 gnd.t71 gnd.t70 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X368 a_n2982_8322.t2 a_n2982_13878.t107 a_n8964_8799.t6 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X369 a_n3827_n3924.t39 plus.t26 a_n8964_8799.t21 gnd.t171 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X370 vdd.t73 a_n8964_8799.t135 CSoutput.t18 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X371 CSoutput.t17 a_n8964_8799.t136 vdd.t71 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X372 CSoutput.t16 a_n8964_8799.t137 vdd.t69 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X373 diffpairibias.t1 diffpairibias.t0 gnd.t6 gnd.t5 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X374 a_n3827_n3924.t44 plus.t27 a_n8964_8799.t20 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X375 CSoutput.t144 commonsourceibias.t122 gnd.t156 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X376 CSoutput.t178 a_n2982_8322.t32 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X377 vdd.t9 a_n2982_13878.t108 a_n2804_13878.t24 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X378 gnd.t155 commonsourceibias.t123 CSoutput.t143 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X379 a_n8964_8799.t19 plus.t28 a_n3827_n3924.t32 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X380 CSoutput.t15 a_n8964_8799.t138 vdd.t67 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X381 gnd.t189 gnd.t186 gnd.t188 gnd.t187 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X382 gnd.t185 gnd.t182 gnd.t184 gnd.t183 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X383 a_n3827_n3924.t3 minus.t27 a_n2982_13878.t2 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X384 vdd.t192 CSoutput.t179 output.t5 gnd.t136 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X385 vdd.t65 a_n8964_8799.t139 CSoutput.t14 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X386 CSoutput.t121 commonsourceibias.t124 gnd.t92 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X387 output.t4 CSoutput.t180 vdd.t193 gnd.t137 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X388 gnd.t48 commonsourceibias.t125 CSoutput.t110 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X389 a_n2982_8322.t1 a_n2982_13878.t109 a_n8964_8799.t45 vdd.t7 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X390 a_n2982_13878.t66 minus.t28 a_n3827_n3924.t24 gnd.t166 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X391 gnd.t46 commonsourceibias.t126 CSoutput.t109 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X392 a_n2982_8322.t0 a_n2982_13878.t110 a_n8964_8799.t7 vdd.t6 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X393 vdd.t63 a_n8964_8799.t140 CSoutput.t13 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X394 vdd.t61 a_n8964_8799.t141 CSoutput.t12 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X395 CSoutput.t11 a_n8964_8799.t142 vdd.t59 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X396 output.t3 CSoutput.t181 vdd.t191 gnd.t103 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X397 gnd.t12 commonsourceibias.t127 CSoutput.t1 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X398 vdd.t207 vdd.t204 vdd.t206 vdd.t205 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X399 a_n2982_8322.t24 a_n2982_13878.t111 vdd.t3 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X400 a_n2804_13878.t1 a_n2982_13878.t21 a_n2982_13878.t22 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X401 minus.t0 gnd.t179 gnd.t181 gnd.t180 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X402 vdd.t203 vdd.t200 vdd.t202 vdd.t201 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X403 commonsourceibias.t1 commonsourceibias.t0 gnd.t170 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X404 a_n3827_n3924.t50 diffpairibias.t29 gnd.t299 gnd.t298 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X405 vdd.t199 vdd.t196 vdd.t198 vdd.t197 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X406 CSoutput.t10 a_n8964_8799.t143 vdd.t57 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X407 a_n2982_13878.t50 a_n2982_13878.t49 a_n2804_13878.t0 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 plus.n53 plus.t20 323.478
R1 plus.n11 plus.t15 323.478
R2 plus.n52 plus.t19 297.12
R3 plus.n56 plus.t26 297.12
R4 plus.n58 plus.t25 297.12
R5 plus.n62 plus.t27 297.12
R6 plus.n64 plus.t9 297.12
R7 plus.n68 plus.t7 297.12
R8 plus.n70 plus.t14 297.12
R9 plus.n74 plus.t12 297.12
R10 plus.n76 plus.t28 297.12
R11 plus.n80 plus.t10 297.12
R12 plus.n82 plus.t8 297.12
R13 plus.n40 plus.t21 297.12
R14 plus.n38 plus.t22 297.12
R15 plus.n2 plus.t16 297.12
R16 plus.n32 plus.t17 297.12
R17 plus.n4 plus.t11 297.12
R18 plus.n26 plus.t5 297.12
R19 plus.n6 plus.t6 297.12
R20 plus.n20 plus.t23 297.12
R21 plus.n8 plus.t24 297.12
R22 plus.n14 plus.t18 297.12
R23 plus.n10 plus.t13 297.12
R24 plus.n86 plus.t2 243.97
R25 plus.n86 plus.n85 223.454
R26 plus.n88 plus.n87 223.454
R27 plus.n83 plus.n82 161.3
R28 plus.n81 plus.n42 161.3
R29 plus.n80 plus.n79 161.3
R30 plus.n78 plus.n43 161.3
R31 plus.n77 plus.n76 161.3
R32 plus.n75 plus.n44 161.3
R33 plus.n74 plus.n73 161.3
R34 plus.n72 plus.n45 161.3
R35 plus.n71 plus.n70 161.3
R36 plus.n69 plus.n46 161.3
R37 plus.n68 plus.n67 161.3
R38 plus.n66 plus.n47 161.3
R39 plus.n65 plus.n64 161.3
R40 plus.n63 plus.n48 161.3
R41 plus.n62 plus.n61 161.3
R42 plus.n60 plus.n49 161.3
R43 plus.n59 plus.n58 161.3
R44 plus.n57 plus.n50 161.3
R45 plus.n56 plus.n55 161.3
R46 plus.n54 plus.n51 161.3
R47 plus.n13 plus.n12 161.3
R48 plus.n14 plus.n9 161.3
R49 plus.n16 plus.n15 161.3
R50 plus.n17 plus.n8 161.3
R51 plus.n19 plus.n18 161.3
R52 plus.n20 plus.n7 161.3
R53 plus.n22 plus.n21 161.3
R54 plus.n23 plus.n6 161.3
R55 plus.n25 plus.n24 161.3
R56 plus.n26 plus.n5 161.3
R57 plus.n28 plus.n27 161.3
R58 plus.n29 plus.n4 161.3
R59 plus.n31 plus.n30 161.3
R60 plus.n32 plus.n3 161.3
R61 plus.n34 plus.n33 161.3
R62 plus.n35 plus.n2 161.3
R63 plus.n37 plus.n36 161.3
R64 plus.n38 plus.n1 161.3
R65 plus.n39 plus.n0 161.3
R66 plus.n41 plus.n40 161.3
R67 plus.n82 plus.n81 46.0096
R68 plus.n40 plus.n39 46.0096
R69 plus.n54 plus.n53 45.0871
R70 plus.n12 plus.n11 45.0871
R71 plus.n52 plus.n51 41.6278
R72 plus.n80 plus.n43 41.6278
R73 plus.n38 plus.n37 41.6278
R74 plus.n13 plus.n10 41.6278
R75 plus.n57 plus.n56 37.246
R76 plus.n76 plus.n75 37.246
R77 plus.n33 plus.n2 37.246
R78 plus.n15 plus.n14 37.246
R79 plus.n84 plus.n83 33.1766
R80 plus.n58 plus.n49 32.8641
R81 plus.n74 plus.n45 32.8641
R82 plus.n32 plus.n31 32.8641
R83 plus.n19 plus.n8 32.8641
R84 plus.n63 plus.n62 28.4823
R85 plus.n70 plus.n69 28.4823
R86 plus.n27 plus.n4 28.4823
R87 plus.n21 plus.n20 28.4823
R88 plus.n64 plus.n47 24.1005
R89 plus.n68 plus.n47 24.1005
R90 plus.n26 plus.n25 24.1005
R91 plus.n25 plus.n6 24.1005
R92 plus.n85 plus.t3 19.8005
R93 plus.n85 plus.t1 19.8005
R94 plus.n87 plus.t4 19.8005
R95 plus.n87 plus.t0 19.8005
R96 plus.n64 plus.n63 19.7187
R97 plus.n69 plus.n68 19.7187
R98 plus.n27 plus.n26 19.7187
R99 plus.n21 plus.n6 19.7187
R100 plus.n62 plus.n49 15.3369
R101 plus.n70 plus.n45 15.3369
R102 plus.n31 plus.n4 15.3369
R103 plus.n20 plus.n19 15.3369
R104 plus plus.n89 14.8628
R105 plus.n53 plus.n52 14.1472
R106 plus.n11 plus.n10 14.1472
R107 plus.n84 plus.n41 11.8774
R108 plus.n58 plus.n57 10.955
R109 plus.n75 plus.n74 10.955
R110 plus.n33 plus.n32 10.955
R111 plus.n15 plus.n8 10.955
R112 plus.n56 plus.n51 6.57323
R113 plus.n76 plus.n43 6.57323
R114 plus.n37 plus.n2 6.57323
R115 plus.n14 plus.n13 6.57323
R116 plus.n89 plus.n88 5.40567
R117 plus.n81 plus.n80 2.19141
R118 plus.n39 plus.n38 2.19141
R119 plus.n89 plus.n84 1.188
R120 plus.n88 plus.n86 0.716017
R121 plus.n55 plus.n54 0.189894
R122 plus.n55 plus.n50 0.189894
R123 plus.n59 plus.n50 0.189894
R124 plus.n60 plus.n59 0.189894
R125 plus.n61 plus.n60 0.189894
R126 plus.n61 plus.n48 0.189894
R127 plus.n65 plus.n48 0.189894
R128 plus.n66 plus.n65 0.189894
R129 plus.n67 plus.n66 0.189894
R130 plus.n67 plus.n46 0.189894
R131 plus.n71 plus.n46 0.189894
R132 plus.n72 plus.n71 0.189894
R133 plus.n73 plus.n72 0.189894
R134 plus.n73 plus.n44 0.189894
R135 plus.n77 plus.n44 0.189894
R136 plus.n78 plus.n77 0.189894
R137 plus.n79 plus.n78 0.189894
R138 plus.n79 plus.n42 0.189894
R139 plus.n83 plus.n42 0.189894
R140 plus.n41 plus.n0 0.189894
R141 plus.n1 plus.n0 0.189894
R142 plus.n36 plus.n1 0.189894
R143 plus.n36 plus.n35 0.189894
R144 plus.n35 plus.n34 0.189894
R145 plus.n34 plus.n3 0.189894
R146 plus.n30 plus.n3 0.189894
R147 plus.n30 plus.n29 0.189894
R148 plus.n29 plus.n28 0.189894
R149 plus.n28 plus.n5 0.189894
R150 plus.n24 plus.n5 0.189894
R151 plus.n24 plus.n23 0.189894
R152 plus.n23 plus.n22 0.189894
R153 plus.n22 plus.n7 0.189894
R154 plus.n18 plus.n7 0.189894
R155 plus.n18 plus.n17 0.189894
R156 plus.n17 plus.n16 0.189894
R157 plus.n16 plus.n9 0.189894
R158 plus.n12 plus.n9 0.189894
R159 a_n3827_n3924.n9 a_n3827_n3924.t6 214.994
R160 a_n3827_n3924.n6 a_n3827_n3924.t14 214.786
R161 a_n3827_n3924.n6 a_n3827_n3924.t8 214.321
R162 a_n3827_n3924.n6 a_n3827_n3924.t56 214.321
R163 a_n3827_n3924.n6 a_n3827_n3924.t7 214.321
R164 a_n3827_n3924.n8 a_n3827_n3924.t50 214.321
R165 a_n3827_n3924.n8 a_n3827_n3924.t49 214.321
R166 a_n3827_n3924.n7 a_n3827_n3924.t57 214.321
R167 a_n3827_n3924.n9 a_n3827_n3924.t13 214.321
R168 a_n3827_n3924.n9 a_n3827_n3924.t0 214.321
R169 a_n3827_n3924.n1 a_n3827_n3924.t25 55.8337
R170 a_n3827_n3924.n1 a_n3827_n3924.t24 55.8337
R171 a_n3827_n3924.t1 a_n3827_n3924.n12 55.8337
R172 a_n3827_n3924.n0 a_n3827_n3924.t45 55.8335
R173 a_n3827_n3924.n10 a_n3827_n3924.t51 55.8335
R174 a_n3827_n3924.n4 a_n3827_n3924.t22 55.8335
R175 a_n3827_n3924.n4 a_n3827_n3924.t29 55.8335
R176 a_n3827_n3924.n3 a_n3827_n3924.t26 55.8335
R177 a_n3827_n3924.n0 a_n3827_n3924.n24 53.0052
R178 a_n3827_n3924.n0 a_n3827_n3924.n25 53.0052
R179 a_n3827_n3924.n0 a_n3827_n3924.n26 53.0052
R180 a_n3827_n3924.n1 a_n3827_n3924.n27 53.0052
R181 a_n3827_n3924.n1 a_n3827_n3924.n28 53.0052
R182 a_n3827_n3924.n1 a_n3827_n3924.n29 53.0052
R183 a_n3827_n3924.n1 a_n3827_n3924.n30 53.0052
R184 a_n3827_n3924.n11 a_n3827_n3924.n31 53.0052
R185 a_n3827_n3924.n11 a_n3827_n3924.n32 53.0052
R186 a_n3827_n3924.n12 a_n3827_n3924.n33 53.0052
R187 a_n3827_n3924.n10 a_n3827_n3924.n22 53.0051
R188 a_n3827_n3924.n2 a_n3827_n3924.n21 53.0051
R189 a_n3827_n3924.n2 a_n3827_n3924.n20 53.0051
R190 a_n3827_n3924.n2 a_n3827_n3924.n19 53.0051
R191 a_n3827_n3924.n2 a_n3827_n3924.n18 53.0051
R192 a_n3827_n3924.n4 a_n3827_n3924.n17 53.0051
R193 a_n3827_n3924.n4 a_n3827_n3924.n16 53.0051
R194 a_n3827_n3924.n4 a_n3827_n3924.n15 53.0051
R195 a_n3827_n3924.n3 a_n3827_n3924.n14 53.0051
R196 a_n3827_n3924.n3 a_n3827_n3924.n13 53.0051
R197 a_n3827_n3924.n12 a_n3827_n3924.n5 12.1986
R198 a_n3827_n3924.n0 a_n3827_n3924.n23 12.1986
R199 a_n3827_n3924.n3 a_n3827_n3924.n5 5.11903
R200 a_n3827_n3924.n23 a_n3827_n3924.n10 5.11903
R201 a_n3827_n3924.n24 a_n3827_n3924.t32 2.82907
R202 a_n3827_n3924.n24 a_n3827_n3924.t33 2.82907
R203 a_n3827_n3924.n25 a_n3827_n3924.t38 2.82907
R204 a_n3827_n3924.n25 a_n3827_n3924.t37 2.82907
R205 a_n3827_n3924.n26 a_n3827_n3924.t41 2.82907
R206 a_n3827_n3924.n26 a_n3827_n3924.t42 2.82907
R207 a_n3827_n3924.n27 a_n3827_n3924.t40 2.82907
R208 a_n3827_n3924.n27 a_n3827_n3924.t44 2.82907
R209 a_n3827_n3924.n28 a_n3827_n3924.t46 2.82907
R210 a_n3827_n3924.n28 a_n3827_n3924.t39 2.82907
R211 a_n3827_n3924.n29 a_n3827_n3924.t18 2.82907
R212 a_n3827_n3924.n29 a_n3827_n3924.t3 2.82907
R213 a_n3827_n3924.n30 a_n3827_n3924.t19 2.82907
R214 a_n3827_n3924.n30 a_n3827_n3924.t54 2.82907
R215 a_n3827_n3924.n31 a_n3827_n3924.t16 2.82907
R216 a_n3827_n3924.n31 a_n3827_n3924.t11 2.82907
R217 a_n3827_n3924.n32 a_n3827_n3924.t5 2.82907
R218 a_n3827_n3924.n32 a_n3827_n3924.t20 2.82907
R219 a_n3827_n3924.n33 a_n3827_n3924.t21 2.82907
R220 a_n3827_n3924.n33 a_n3827_n3924.t9 2.82907
R221 a_n3827_n3924.n22 a_n3827_n3924.t2 2.82907
R222 a_n3827_n3924.n22 a_n3827_n3924.t15 2.82907
R223 a_n3827_n3924.n21 a_n3827_n3924.t10 2.82907
R224 a_n3827_n3924.n21 a_n3827_n3924.t23 2.82907
R225 a_n3827_n3924.n20 a_n3827_n3924.t12 2.82907
R226 a_n3827_n3924.n20 a_n3827_n3924.t17 2.82907
R227 a_n3827_n3924.n19 a_n3827_n3924.t55 2.82907
R228 a_n3827_n3924.n19 a_n3827_n3924.t4 2.82907
R229 a_n3827_n3924.n18 a_n3827_n3924.t52 2.82907
R230 a_n3827_n3924.n18 a_n3827_n3924.t53 2.82907
R231 a_n3827_n3924.n17 a_n3827_n3924.t27 2.82907
R232 a_n3827_n3924.n17 a_n3827_n3924.t48 2.82907
R233 a_n3827_n3924.n16 a_n3827_n3924.t28 2.82907
R234 a_n3827_n3924.n16 a_n3827_n3924.t30 2.82907
R235 a_n3827_n3924.n15 a_n3827_n3924.t31 2.82907
R236 a_n3827_n3924.n15 a_n3827_n3924.t43 2.82907
R237 a_n3827_n3924.n14 a_n3827_n3924.t36 2.82907
R238 a_n3827_n3924.n14 a_n3827_n3924.t35 2.82907
R239 a_n3827_n3924.n13 a_n3827_n3924.t34 2.82907
R240 a_n3827_n3924.n13 a_n3827_n3924.t47 2.82907
R241 a_n3827_n3924.n1 a_n3827_n3924.n0 2.66429
R242 a_n3827_n3924.n6 a_n3827_n3924.n8 2.22216
R243 a_n3827_n3924.n2 a_n3827_n3924.n4 2.01128
R244 a_n3827_n3924.n23 a_n3827_n3924.n6 1.95694
R245 a_n3827_n3924.n9 a_n3827_n3924.n5 1.95694
R246 a_n3827_n3924.n4 a_n3827_n3924.n3 1.77636
R247 a_n3827_n3924.n10 a_n3827_n3924.n2 1.77636
R248 a_n3827_n3924.n11 a_n3827_n3924.n1 1.56731
R249 a_n3827_n3924.n8 a_n3827_n3924.n7 1.34352
R250 a_n3827_n3924.n7 a_n3827_n3924.n9 1.34352
R251 a_n3827_n3924.n12 a_n3827_n3924.n11 1.3324
R252 a_n8964_8799.n186 a_n8964_8799.t124 485.149
R253 a_n8964_8799.n234 a_n8964_8799.t136 485.149
R254 a_n8964_8799.n283 a_n8964_8799.t91 485.149
R255 a_n8964_8799.n38 a_n8964_8799.t86 485.149
R256 a_n8964_8799.n86 a_n8964_8799.t95 485.149
R257 a_n8964_8799.n135 a_n8964_8799.t89 485.149
R258 a_n8964_8799.n218 a_n8964_8799.t55 464.166
R259 a_n8964_8799.n217 a_n8964_8799.t53 464.166
R260 a_n8964_8799.n173 a_n8964_8799.t121 464.166
R261 a_n8964_8799.n211 a_n8964_8799.t69 464.166
R262 a_n8964_8799.n210 a_n8964_8799.t57 464.166
R263 a_n8964_8799.n176 a_n8964_8799.t127 464.166
R264 a_n8964_8799.n204 a_n8964_8799.t90 464.166
R265 a_n8964_8799.n203 a_n8964_8799.t70 464.166
R266 a_n8964_8799.n179 a_n8964_8799.t141 464.166
R267 a_n8964_8799.n198 a_n8964_8799.t106 464.166
R268 a_n8964_8799.n196 a_n8964_8799.t72 464.166
R269 a_n8964_8799.n182 a_n8964_8799.t137 464.166
R270 a_n8964_8799.n191 a_n8964_8799.t108 464.166
R271 a_n8964_8799.n189 a_n8964_8799.t84 464.166
R272 a_n8964_8799.n185 a_n8964_8799.t54 464.166
R273 a_n8964_8799.n266 a_n8964_8799.t62 464.166
R274 a_n8964_8799.n265 a_n8964_8799.t61 464.166
R275 a_n8964_8799.n221 a_n8964_8799.t135 464.166
R276 a_n8964_8799.n259 a_n8964_8799.t75 464.166
R277 a_n8964_8799.n258 a_n8964_8799.t68 464.166
R278 a_n8964_8799.n224 a_n8964_8799.t138 464.166
R279 a_n8964_8799.n252 a_n8964_8799.t102 464.166
R280 a_n8964_8799.n251 a_n8964_8799.t78 464.166
R281 a_n8964_8799.n227 a_n8964_8799.t56 464.166
R282 a_n8964_8799.n246 a_n8964_8799.t115 464.166
R283 a_n8964_8799.n244 a_n8964_8799.t79 464.166
R284 a_n8964_8799.n230 a_n8964_8799.t49 464.166
R285 a_n8964_8799.n239 a_n8964_8799.t120 464.166
R286 a_n8964_8799.n237 a_n8964_8799.t92 464.166
R287 a_n8964_8799.n233 a_n8964_8799.t63 464.166
R288 a_n8964_8799.n315 a_n8964_8799.t101 464.166
R289 a_n8964_8799.n314 a_n8964_8799.t119 464.166
R290 a_n8964_8799.n270 a_n8964_8799.t67 464.166
R291 a_n8964_8799.n308 a_n8964_8799.t133 464.166
R292 a_n8964_8799.n307 a_n8964_8799.t82 464.166
R293 a_n8964_8799.n273 a_n8964_8799.t128 464.166
R294 a_n8964_8799.n301 a_n8964_8799.t71 464.166
R295 a_n8964_8799.n300 a_n8964_8799.t110 464.166
R296 a_n8964_8799.n276 a_n8964_8799.t59 464.166
R297 a_n8964_8799.n295 a_n8964_8799.t98 464.166
R298 a_n8964_8799.n293 a_n8964_8799.t77 464.166
R299 a_n8964_8799.n279 a_n8964_8799.t117 464.166
R300 a_n8964_8799.n288 a_n8964_8799.t65 464.166
R301 a_n8964_8799.n286 a_n8964_8799.t105 464.166
R302 a_n8964_8799.n282 a_n8964_8799.t52 464.166
R303 a_n8964_8799.n37 a_n8964_8799.t111 464.166
R304 a_n8964_8799.n41 a_n8964_8799.t50 464.166
R305 a_n8964_8799.n35 a_n8964_8799.t74 464.166
R306 a_n8964_8799.n46 a_n8964_8799.t107 464.166
R307 a_n8964_8799.n48 a_n8964_8799.t134 464.166
R308 a_n8964_8799.n52 a_n8964_8799.t73 464.166
R309 a_n8964_8799.n53 a_n8964_8799.t103 464.166
R310 a_n8964_8799.n31 a_n8964_8799.t130 464.166
R311 a_n8964_8799.n58 a_n8964_8799.t131 464.166
R312 a_n8964_8799.n60 a_n8964_8799.t88 464.166
R313 a_n8964_8799.n64 a_n8964_8799.t114 464.166
R314 a_n8964_8799.n65 a_n8964_8799.t129 464.166
R315 a_n8964_8799.n27 a_n8964_8799.t85 464.166
R316 a_n8964_8799.n71 a_n8964_8799.t87 464.166
R317 a_n8964_8799.n72 a_n8964_8799.t112 464.166
R318 a_n8964_8799.n85 a_n8964_8799.t122 464.166
R319 a_n8964_8799.n89 a_n8964_8799.t60 464.166
R320 a_n8964_8799.n83 a_n8964_8799.t83 464.166
R321 a_n8964_8799.n94 a_n8964_8799.t116 464.166
R322 a_n8964_8799.n96 a_n8964_8799.t143 464.166
R323 a_n8964_8799.n100 a_n8964_8799.t80 464.166
R324 a_n8964_8799.n101 a_n8964_8799.t113 464.166
R325 a_n8964_8799.n79 a_n8964_8799.t140 464.166
R326 a_n8964_8799.n106 a_n8964_8799.t142 464.166
R327 a_n8964_8799.n108 a_n8964_8799.t99 464.166
R328 a_n8964_8799.n112 a_n8964_8799.t126 464.166
R329 a_n8964_8799.n113 a_n8964_8799.t139 464.166
R330 a_n8964_8799.n75 a_n8964_8799.t94 464.166
R331 a_n8964_8799.n119 a_n8964_8799.t96 464.166
R332 a_n8964_8799.n120 a_n8964_8799.t123 464.166
R333 a_n8964_8799.n134 a_n8964_8799.t51 464.166
R334 a_n8964_8799.n138 a_n8964_8799.t104 464.166
R335 a_n8964_8799.n132 a_n8964_8799.t64 464.166
R336 a_n8964_8799.n143 a_n8964_8799.t118 464.166
R337 a_n8964_8799.n145 a_n8964_8799.t76 464.166
R338 a_n8964_8799.n149 a_n8964_8799.t97 464.166
R339 a_n8964_8799.n150 a_n8964_8799.t58 464.166
R340 a_n8964_8799.n128 a_n8964_8799.t109 464.166
R341 a_n8964_8799.n155 a_n8964_8799.t93 464.166
R342 a_n8964_8799.n157 a_n8964_8799.t125 464.166
R343 a_n8964_8799.n161 a_n8964_8799.t81 464.166
R344 a_n8964_8799.n162 a_n8964_8799.t132 464.166
R345 a_n8964_8799.n124 a_n8964_8799.t66 464.166
R346 a_n8964_8799.n168 a_n8964_8799.t48 464.166
R347 a_n8964_8799.n169 a_n8964_8799.t100 464.166
R348 a_n8964_8799.n188 a_n8964_8799.n187 161.3
R349 a_n8964_8799.n189 a_n8964_8799.n184 161.3
R350 a_n8964_8799.n190 a_n8964_8799.n183 161.3
R351 a_n8964_8799.n192 a_n8964_8799.n191 161.3
R352 a_n8964_8799.n193 a_n8964_8799.n182 161.3
R353 a_n8964_8799.n195 a_n8964_8799.n194 161.3
R354 a_n8964_8799.n196 a_n8964_8799.n181 161.3
R355 a_n8964_8799.n197 a_n8964_8799.n180 161.3
R356 a_n8964_8799.n199 a_n8964_8799.n198 161.3
R357 a_n8964_8799.n200 a_n8964_8799.n179 161.3
R358 a_n8964_8799.n202 a_n8964_8799.n201 161.3
R359 a_n8964_8799.n203 a_n8964_8799.n178 161.3
R360 a_n8964_8799.n204 a_n8964_8799.n177 161.3
R361 a_n8964_8799.n206 a_n8964_8799.n205 161.3
R362 a_n8964_8799.n207 a_n8964_8799.n176 161.3
R363 a_n8964_8799.n209 a_n8964_8799.n208 161.3
R364 a_n8964_8799.n210 a_n8964_8799.n175 161.3
R365 a_n8964_8799.n211 a_n8964_8799.n174 161.3
R366 a_n8964_8799.n213 a_n8964_8799.n212 161.3
R367 a_n8964_8799.n214 a_n8964_8799.n173 161.3
R368 a_n8964_8799.n216 a_n8964_8799.n215 161.3
R369 a_n8964_8799.n217 a_n8964_8799.n172 161.3
R370 a_n8964_8799.n219 a_n8964_8799.n218 161.3
R371 a_n8964_8799.n236 a_n8964_8799.n235 161.3
R372 a_n8964_8799.n237 a_n8964_8799.n232 161.3
R373 a_n8964_8799.n238 a_n8964_8799.n231 161.3
R374 a_n8964_8799.n240 a_n8964_8799.n239 161.3
R375 a_n8964_8799.n241 a_n8964_8799.n230 161.3
R376 a_n8964_8799.n243 a_n8964_8799.n242 161.3
R377 a_n8964_8799.n244 a_n8964_8799.n229 161.3
R378 a_n8964_8799.n245 a_n8964_8799.n228 161.3
R379 a_n8964_8799.n247 a_n8964_8799.n246 161.3
R380 a_n8964_8799.n248 a_n8964_8799.n227 161.3
R381 a_n8964_8799.n250 a_n8964_8799.n249 161.3
R382 a_n8964_8799.n251 a_n8964_8799.n226 161.3
R383 a_n8964_8799.n252 a_n8964_8799.n225 161.3
R384 a_n8964_8799.n254 a_n8964_8799.n253 161.3
R385 a_n8964_8799.n255 a_n8964_8799.n224 161.3
R386 a_n8964_8799.n257 a_n8964_8799.n256 161.3
R387 a_n8964_8799.n258 a_n8964_8799.n223 161.3
R388 a_n8964_8799.n259 a_n8964_8799.n222 161.3
R389 a_n8964_8799.n261 a_n8964_8799.n260 161.3
R390 a_n8964_8799.n262 a_n8964_8799.n221 161.3
R391 a_n8964_8799.n264 a_n8964_8799.n263 161.3
R392 a_n8964_8799.n265 a_n8964_8799.n220 161.3
R393 a_n8964_8799.n267 a_n8964_8799.n266 161.3
R394 a_n8964_8799.n285 a_n8964_8799.n284 161.3
R395 a_n8964_8799.n286 a_n8964_8799.n281 161.3
R396 a_n8964_8799.n287 a_n8964_8799.n280 161.3
R397 a_n8964_8799.n289 a_n8964_8799.n288 161.3
R398 a_n8964_8799.n290 a_n8964_8799.n279 161.3
R399 a_n8964_8799.n292 a_n8964_8799.n291 161.3
R400 a_n8964_8799.n293 a_n8964_8799.n278 161.3
R401 a_n8964_8799.n294 a_n8964_8799.n277 161.3
R402 a_n8964_8799.n296 a_n8964_8799.n295 161.3
R403 a_n8964_8799.n297 a_n8964_8799.n276 161.3
R404 a_n8964_8799.n299 a_n8964_8799.n298 161.3
R405 a_n8964_8799.n300 a_n8964_8799.n275 161.3
R406 a_n8964_8799.n301 a_n8964_8799.n274 161.3
R407 a_n8964_8799.n303 a_n8964_8799.n302 161.3
R408 a_n8964_8799.n304 a_n8964_8799.n273 161.3
R409 a_n8964_8799.n306 a_n8964_8799.n305 161.3
R410 a_n8964_8799.n307 a_n8964_8799.n272 161.3
R411 a_n8964_8799.n308 a_n8964_8799.n271 161.3
R412 a_n8964_8799.n310 a_n8964_8799.n309 161.3
R413 a_n8964_8799.n311 a_n8964_8799.n270 161.3
R414 a_n8964_8799.n313 a_n8964_8799.n312 161.3
R415 a_n8964_8799.n314 a_n8964_8799.n269 161.3
R416 a_n8964_8799.n316 a_n8964_8799.n315 161.3
R417 a_n8964_8799.n73 a_n8964_8799.n72 161.3
R418 a_n8964_8799.n71 a_n8964_8799.n26 161.3
R419 a_n8964_8799.n70 a_n8964_8799.n69 161.3
R420 a_n8964_8799.n68 a_n8964_8799.n27 161.3
R421 a_n8964_8799.n67 a_n8964_8799.n66 161.3
R422 a_n8964_8799.n65 a_n8964_8799.n28 161.3
R423 a_n8964_8799.n64 a_n8964_8799.n63 161.3
R424 a_n8964_8799.n62 a_n8964_8799.n29 161.3
R425 a_n8964_8799.n61 a_n8964_8799.n60 161.3
R426 a_n8964_8799.n59 a_n8964_8799.n30 161.3
R427 a_n8964_8799.n58 a_n8964_8799.n57 161.3
R428 a_n8964_8799.n56 a_n8964_8799.n31 161.3
R429 a_n8964_8799.n55 a_n8964_8799.n54 161.3
R430 a_n8964_8799.n53 a_n8964_8799.n32 161.3
R431 a_n8964_8799.n52 a_n8964_8799.n51 161.3
R432 a_n8964_8799.n50 a_n8964_8799.n33 161.3
R433 a_n8964_8799.n49 a_n8964_8799.n48 161.3
R434 a_n8964_8799.n47 a_n8964_8799.n34 161.3
R435 a_n8964_8799.n46 a_n8964_8799.n45 161.3
R436 a_n8964_8799.n44 a_n8964_8799.n35 161.3
R437 a_n8964_8799.n43 a_n8964_8799.n42 161.3
R438 a_n8964_8799.n41 a_n8964_8799.n36 161.3
R439 a_n8964_8799.n40 a_n8964_8799.n39 161.3
R440 a_n8964_8799.n121 a_n8964_8799.n120 161.3
R441 a_n8964_8799.n119 a_n8964_8799.n74 161.3
R442 a_n8964_8799.n118 a_n8964_8799.n117 161.3
R443 a_n8964_8799.n116 a_n8964_8799.n75 161.3
R444 a_n8964_8799.n115 a_n8964_8799.n114 161.3
R445 a_n8964_8799.n113 a_n8964_8799.n76 161.3
R446 a_n8964_8799.n112 a_n8964_8799.n111 161.3
R447 a_n8964_8799.n110 a_n8964_8799.n77 161.3
R448 a_n8964_8799.n109 a_n8964_8799.n108 161.3
R449 a_n8964_8799.n107 a_n8964_8799.n78 161.3
R450 a_n8964_8799.n106 a_n8964_8799.n105 161.3
R451 a_n8964_8799.n104 a_n8964_8799.n79 161.3
R452 a_n8964_8799.n103 a_n8964_8799.n102 161.3
R453 a_n8964_8799.n101 a_n8964_8799.n80 161.3
R454 a_n8964_8799.n100 a_n8964_8799.n99 161.3
R455 a_n8964_8799.n98 a_n8964_8799.n81 161.3
R456 a_n8964_8799.n97 a_n8964_8799.n96 161.3
R457 a_n8964_8799.n95 a_n8964_8799.n82 161.3
R458 a_n8964_8799.n94 a_n8964_8799.n93 161.3
R459 a_n8964_8799.n92 a_n8964_8799.n83 161.3
R460 a_n8964_8799.n91 a_n8964_8799.n90 161.3
R461 a_n8964_8799.n89 a_n8964_8799.n84 161.3
R462 a_n8964_8799.n88 a_n8964_8799.n87 161.3
R463 a_n8964_8799.n170 a_n8964_8799.n169 161.3
R464 a_n8964_8799.n168 a_n8964_8799.n123 161.3
R465 a_n8964_8799.n167 a_n8964_8799.n166 161.3
R466 a_n8964_8799.n165 a_n8964_8799.n124 161.3
R467 a_n8964_8799.n164 a_n8964_8799.n163 161.3
R468 a_n8964_8799.n162 a_n8964_8799.n125 161.3
R469 a_n8964_8799.n161 a_n8964_8799.n160 161.3
R470 a_n8964_8799.n159 a_n8964_8799.n126 161.3
R471 a_n8964_8799.n158 a_n8964_8799.n157 161.3
R472 a_n8964_8799.n156 a_n8964_8799.n127 161.3
R473 a_n8964_8799.n155 a_n8964_8799.n154 161.3
R474 a_n8964_8799.n153 a_n8964_8799.n128 161.3
R475 a_n8964_8799.n152 a_n8964_8799.n151 161.3
R476 a_n8964_8799.n150 a_n8964_8799.n129 161.3
R477 a_n8964_8799.n149 a_n8964_8799.n148 161.3
R478 a_n8964_8799.n147 a_n8964_8799.n130 161.3
R479 a_n8964_8799.n146 a_n8964_8799.n145 161.3
R480 a_n8964_8799.n144 a_n8964_8799.n131 161.3
R481 a_n8964_8799.n143 a_n8964_8799.n142 161.3
R482 a_n8964_8799.n141 a_n8964_8799.n132 161.3
R483 a_n8964_8799.n140 a_n8964_8799.n139 161.3
R484 a_n8964_8799.n138 a_n8964_8799.n133 161.3
R485 a_n8964_8799.n137 a_n8964_8799.n136 161.3
R486 a_n8964_8799.n16 a_n8964_8799.n14 98.9633
R487 a_n8964_8799.n5 a_n8964_8799.n3 98.9631
R488 a_n8964_8799.n24 a_n8964_8799.n23 98.6055
R489 a_n8964_8799.n22 a_n8964_8799.n21 98.6055
R490 a_n8964_8799.n20 a_n8964_8799.n19 98.6055
R491 a_n8964_8799.n18 a_n8964_8799.n17 98.6055
R492 a_n8964_8799.n16 a_n8964_8799.n15 98.6055
R493 a_n8964_8799.n5 a_n8964_8799.n4 98.6055
R494 a_n8964_8799.n7 a_n8964_8799.n6 98.6055
R495 a_n8964_8799.n9 a_n8964_8799.n8 98.6055
R496 a_n8964_8799.n11 a_n8964_8799.n10 98.6055
R497 a_n8964_8799.n13 a_n8964_8799.n12 98.6055
R498 a_n8964_8799.n322 a_n8964_8799.n320 81.3764
R499 a_n8964_8799.n334 a_n8964_8799.n332 81.3764
R500 a_n8964_8799.n2 a_n8964_8799.n0 81.3764
R501 a_n8964_8799.n339 a_n8964_8799.n338 80.9326
R502 a_n8964_8799.n331 a_n8964_8799.n330 80.9324
R503 a_n8964_8799.n329 a_n8964_8799.n328 80.9324
R504 a_n8964_8799.n327 a_n8964_8799.n326 80.9324
R505 a_n8964_8799.n324 a_n8964_8799.n323 80.9324
R506 a_n8964_8799.n322 a_n8964_8799.n321 80.9324
R507 a_n8964_8799.n334 a_n8964_8799.n333 80.9324
R508 a_n8964_8799.n336 a_n8964_8799.n335 80.9324
R509 a_n8964_8799.n2 a_n8964_8799.n1 80.9324
R510 a_n8964_8799.n187 a_n8964_8799.n186 70.4033
R511 a_n8964_8799.n235 a_n8964_8799.n234 70.4033
R512 a_n8964_8799.n284 a_n8964_8799.n283 70.4033
R513 a_n8964_8799.n39 a_n8964_8799.n38 70.4033
R514 a_n8964_8799.n87 a_n8964_8799.n86 70.4033
R515 a_n8964_8799.n136 a_n8964_8799.n135 70.4033
R516 a_n8964_8799.n218 a_n8964_8799.n217 48.2005
R517 a_n8964_8799.n211 a_n8964_8799.n210 48.2005
R518 a_n8964_8799.n204 a_n8964_8799.n203 48.2005
R519 a_n8964_8799.n198 a_n8964_8799.n179 48.2005
R520 a_n8964_8799.n191 a_n8964_8799.n182 48.2005
R521 a_n8964_8799.n266 a_n8964_8799.n265 48.2005
R522 a_n8964_8799.n259 a_n8964_8799.n258 48.2005
R523 a_n8964_8799.n252 a_n8964_8799.n251 48.2005
R524 a_n8964_8799.n246 a_n8964_8799.n227 48.2005
R525 a_n8964_8799.n239 a_n8964_8799.n230 48.2005
R526 a_n8964_8799.n315 a_n8964_8799.n314 48.2005
R527 a_n8964_8799.n308 a_n8964_8799.n307 48.2005
R528 a_n8964_8799.n301 a_n8964_8799.n300 48.2005
R529 a_n8964_8799.n295 a_n8964_8799.n276 48.2005
R530 a_n8964_8799.n288 a_n8964_8799.n279 48.2005
R531 a_n8964_8799.n46 a_n8964_8799.n35 48.2005
R532 a_n8964_8799.n53 a_n8964_8799.n52 48.2005
R533 a_n8964_8799.n58 a_n8964_8799.n31 48.2005
R534 a_n8964_8799.n65 a_n8964_8799.n64 48.2005
R535 a_n8964_8799.n72 a_n8964_8799.n71 48.2005
R536 a_n8964_8799.n94 a_n8964_8799.n83 48.2005
R537 a_n8964_8799.n101 a_n8964_8799.n100 48.2005
R538 a_n8964_8799.n106 a_n8964_8799.n79 48.2005
R539 a_n8964_8799.n113 a_n8964_8799.n112 48.2005
R540 a_n8964_8799.n120 a_n8964_8799.n119 48.2005
R541 a_n8964_8799.n143 a_n8964_8799.n132 48.2005
R542 a_n8964_8799.n150 a_n8964_8799.n149 48.2005
R543 a_n8964_8799.n155 a_n8964_8799.n128 48.2005
R544 a_n8964_8799.n162 a_n8964_8799.n161 48.2005
R545 a_n8964_8799.n169 a_n8964_8799.n168 48.2005
R546 a_n8964_8799.n205 a_n8964_8799.n176 47.4702
R547 a_n8964_8799.n197 a_n8964_8799.n196 47.4702
R548 a_n8964_8799.n253 a_n8964_8799.n224 47.4702
R549 a_n8964_8799.n245 a_n8964_8799.n244 47.4702
R550 a_n8964_8799.n302 a_n8964_8799.n273 47.4702
R551 a_n8964_8799.n294 a_n8964_8799.n293 47.4702
R552 a_n8964_8799.n48 a_n8964_8799.n33 47.4702
R553 a_n8964_8799.n60 a_n8964_8799.n59 47.4702
R554 a_n8964_8799.n96 a_n8964_8799.n81 47.4702
R555 a_n8964_8799.n108 a_n8964_8799.n107 47.4702
R556 a_n8964_8799.n145 a_n8964_8799.n130 47.4702
R557 a_n8964_8799.n157 a_n8964_8799.n156 47.4702
R558 a_n8964_8799.n212 a_n8964_8799.n173 46.0096
R559 a_n8964_8799.n190 a_n8964_8799.n189 46.0096
R560 a_n8964_8799.n260 a_n8964_8799.n221 46.0096
R561 a_n8964_8799.n238 a_n8964_8799.n237 46.0096
R562 a_n8964_8799.n309 a_n8964_8799.n270 46.0096
R563 a_n8964_8799.n287 a_n8964_8799.n286 46.0096
R564 a_n8964_8799.n42 a_n8964_8799.n41 46.0096
R565 a_n8964_8799.n66 a_n8964_8799.n27 46.0096
R566 a_n8964_8799.n90 a_n8964_8799.n89 46.0096
R567 a_n8964_8799.n114 a_n8964_8799.n75 46.0096
R568 a_n8964_8799.n139 a_n8964_8799.n138 46.0096
R569 a_n8964_8799.n163 a_n8964_8799.n124 46.0096
R570 a_n8964_8799.n25 a_n8964_8799.n13 34.1553
R571 a_n8964_8799.n337 a_n8964_8799.n331 33.4185
R572 a_n8964_8799.n216 a_n8964_8799.n173 27.0217
R573 a_n8964_8799.n189 a_n8964_8799.n188 27.0217
R574 a_n8964_8799.n264 a_n8964_8799.n221 27.0217
R575 a_n8964_8799.n237 a_n8964_8799.n236 27.0217
R576 a_n8964_8799.n313 a_n8964_8799.n270 27.0217
R577 a_n8964_8799.n286 a_n8964_8799.n285 27.0217
R578 a_n8964_8799.n41 a_n8964_8799.n40 27.0217
R579 a_n8964_8799.n70 a_n8964_8799.n27 27.0217
R580 a_n8964_8799.n89 a_n8964_8799.n88 27.0217
R581 a_n8964_8799.n118 a_n8964_8799.n75 27.0217
R582 a_n8964_8799.n138 a_n8964_8799.n137 27.0217
R583 a_n8964_8799.n167 a_n8964_8799.n124 27.0217
R584 a_n8964_8799.n209 a_n8964_8799.n176 25.5611
R585 a_n8964_8799.n196 a_n8964_8799.n195 25.5611
R586 a_n8964_8799.n257 a_n8964_8799.n224 25.5611
R587 a_n8964_8799.n244 a_n8964_8799.n243 25.5611
R588 a_n8964_8799.n306 a_n8964_8799.n273 25.5611
R589 a_n8964_8799.n293 a_n8964_8799.n292 25.5611
R590 a_n8964_8799.n48 a_n8964_8799.n47 25.5611
R591 a_n8964_8799.n60 a_n8964_8799.n29 25.5611
R592 a_n8964_8799.n96 a_n8964_8799.n95 25.5611
R593 a_n8964_8799.n108 a_n8964_8799.n77 25.5611
R594 a_n8964_8799.n145 a_n8964_8799.n144 25.5611
R595 a_n8964_8799.n157 a_n8964_8799.n126 25.5611
R596 a_n8964_8799.n203 a_n8964_8799.n202 24.1005
R597 a_n8964_8799.n202 a_n8964_8799.n179 24.1005
R598 a_n8964_8799.n251 a_n8964_8799.n250 24.1005
R599 a_n8964_8799.n250 a_n8964_8799.n227 24.1005
R600 a_n8964_8799.n300 a_n8964_8799.n299 24.1005
R601 a_n8964_8799.n299 a_n8964_8799.n276 24.1005
R602 a_n8964_8799.n54 a_n8964_8799.n53 24.1005
R603 a_n8964_8799.n54 a_n8964_8799.n31 24.1005
R604 a_n8964_8799.n102 a_n8964_8799.n101 24.1005
R605 a_n8964_8799.n102 a_n8964_8799.n79 24.1005
R606 a_n8964_8799.n151 a_n8964_8799.n150 24.1005
R607 a_n8964_8799.n151 a_n8964_8799.n128 24.1005
R608 a_n8964_8799.n210 a_n8964_8799.n209 22.6399
R609 a_n8964_8799.n195 a_n8964_8799.n182 22.6399
R610 a_n8964_8799.n258 a_n8964_8799.n257 22.6399
R611 a_n8964_8799.n243 a_n8964_8799.n230 22.6399
R612 a_n8964_8799.n307 a_n8964_8799.n306 22.6399
R613 a_n8964_8799.n292 a_n8964_8799.n279 22.6399
R614 a_n8964_8799.n47 a_n8964_8799.n46 22.6399
R615 a_n8964_8799.n64 a_n8964_8799.n29 22.6399
R616 a_n8964_8799.n95 a_n8964_8799.n94 22.6399
R617 a_n8964_8799.n112 a_n8964_8799.n77 22.6399
R618 a_n8964_8799.n144 a_n8964_8799.n143 22.6399
R619 a_n8964_8799.n161 a_n8964_8799.n126 22.6399
R620 a_n8964_8799.n217 a_n8964_8799.n216 21.1793
R621 a_n8964_8799.n188 a_n8964_8799.n185 21.1793
R622 a_n8964_8799.n265 a_n8964_8799.n264 21.1793
R623 a_n8964_8799.n236 a_n8964_8799.n233 21.1793
R624 a_n8964_8799.n314 a_n8964_8799.n313 21.1793
R625 a_n8964_8799.n285 a_n8964_8799.n282 21.1793
R626 a_n8964_8799.n40 a_n8964_8799.n37 21.1793
R627 a_n8964_8799.n71 a_n8964_8799.n70 21.1793
R628 a_n8964_8799.n88 a_n8964_8799.n85 21.1793
R629 a_n8964_8799.n119 a_n8964_8799.n118 21.1793
R630 a_n8964_8799.n137 a_n8964_8799.n134 21.1793
R631 a_n8964_8799.n168 a_n8964_8799.n167 21.1793
R632 a_n8964_8799.n186 a_n8964_8799.n185 20.9576
R633 a_n8964_8799.n234 a_n8964_8799.n233 20.9576
R634 a_n8964_8799.n283 a_n8964_8799.n282 20.9576
R635 a_n8964_8799.n38 a_n8964_8799.n37 20.9576
R636 a_n8964_8799.n86 a_n8964_8799.n85 20.9576
R637 a_n8964_8799.n135 a_n8964_8799.n134 20.9576
R638 a_n8964_8799.n25 a_n8964_8799.n24 20.7339
R639 a_n8964_8799.n325 a_n8964_8799.n319 12.3339
R640 a_n8964_8799.n319 a_n8964_8799.n25 11.4887
R641 a_n8964_8799.n268 a_n8964_8799.n219 9.07815
R642 a_n8964_8799.n122 a_n8964_8799.n73 9.07815
R643 a_n8964_8799.n318 a_n8964_8799.n171 7.2142
R644 a_n8964_8799.n318 a_n8964_8799.n317 6.79277
R645 a_n8964_8799.n268 a_n8964_8799.n267 4.9702
R646 a_n8964_8799.n317 a_n8964_8799.n316 4.9702
R647 a_n8964_8799.n122 a_n8964_8799.n121 4.9702
R648 a_n8964_8799.n171 a_n8964_8799.n170 4.9702
R649 a_n8964_8799.n317 a_n8964_8799.n268 4.10845
R650 a_n8964_8799.n171 a_n8964_8799.n122 4.10845
R651 a_n8964_8799.n23 a_n8964_8799.t12 3.61217
R652 a_n8964_8799.n23 a_n8964_8799.t11 3.61217
R653 a_n8964_8799.n21 a_n8964_8799.t16 3.61217
R654 a_n8964_8799.n21 a_n8964_8799.t9 3.61217
R655 a_n8964_8799.n19 a_n8964_8799.t6 3.61217
R656 a_n8964_8799.n19 a_n8964_8799.t18 3.61217
R657 a_n8964_8799.n17 a_n8964_8799.t17 3.61217
R658 a_n8964_8799.n17 a_n8964_8799.t3 3.61217
R659 a_n8964_8799.n15 a_n8964_8799.t10 3.61217
R660 a_n8964_8799.n15 a_n8964_8799.t47 3.61217
R661 a_n8964_8799.n14 a_n8964_8799.t7 3.61217
R662 a_n8964_8799.n14 a_n8964_8799.t8 3.61217
R663 a_n8964_8799.n3 a_n8964_8799.t5 3.61217
R664 a_n8964_8799.n3 a_n8964_8799.t44 3.61217
R665 a_n8964_8799.n4 a_n8964_8799.t4 3.61217
R666 a_n8964_8799.n4 a_n8964_8799.t46 3.61217
R667 a_n8964_8799.n6 a_n8964_8799.t2 3.61217
R668 a_n8964_8799.n6 a_n8964_8799.t13 3.61217
R669 a_n8964_8799.n8 a_n8964_8799.t1 3.61217
R670 a_n8964_8799.n8 a_n8964_8799.t14 3.61217
R671 a_n8964_8799.n10 a_n8964_8799.t43 3.61217
R672 a_n8964_8799.n10 a_n8964_8799.t15 3.61217
R673 a_n8964_8799.n12 a_n8964_8799.t45 3.61217
R674 a_n8964_8799.n12 a_n8964_8799.t0 3.61217
R675 a_n8964_8799.n319 a_n8964_8799.n318 3.4105
R676 a_n8964_8799.n332 a_n8964_8799.t34 2.82907
R677 a_n8964_8799.n332 a_n8964_8799.t32 2.82907
R678 a_n8964_8799.n333 a_n8964_8799.t23 2.82907
R679 a_n8964_8799.n333 a_n8964_8799.t29 2.82907
R680 a_n8964_8799.n335 a_n8964_8799.t41 2.82907
R681 a_n8964_8799.n335 a_n8964_8799.t24 2.82907
R682 a_n8964_8799.n1 a_n8964_8799.t31 2.82907
R683 a_n8964_8799.n1 a_n8964_8799.t30 2.82907
R684 a_n8964_8799.n0 a_n8964_8799.t26 2.82907
R685 a_n8964_8799.n0 a_n8964_8799.t25 2.82907
R686 a_n8964_8799.n330 a_n8964_8799.t37 2.82907
R687 a_n8964_8799.n330 a_n8964_8799.t39 2.82907
R688 a_n8964_8799.n328 a_n8964_8799.t35 2.82907
R689 a_n8964_8799.n328 a_n8964_8799.t19 2.82907
R690 a_n8964_8799.n326 a_n8964_8799.t40 2.82907
R691 a_n8964_8799.n326 a_n8964_8799.t33 2.82907
R692 a_n8964_8799.n323 a_n8964_8799.t20 2.82907
R693 a_n8964_8799.n323 a_n8964_8799.t38 2.82907
R694 a_n8964_8799.n321 a_n8964_8799.t21 2.82907
R695 a_n8964_8799.n321 a_n8964_8799.t22 2.82907
R696 a_n8964_8799.n320 a_n8964_8799.t27 2.82907
R697 a_n8964_8799.n320 a_n8964_8799.t28 2.82907
R698 a_n8964_8799.n339 a_n8964_8799.t36 2.82907
R699 a_n8964_8799.t42 a_n8964_8799.n339 2.82907
R700 a_n8964_8799.n212 a_n8964_8799.n211 2.19141
R701 a_n8964_8799.n191 a_n8964_8799.n190 2.19141
R702 a_n8964_8799.n260 a_n8964_8799.n259 2.19141
R703 a_n8964_8799.n239 a_n8964_8799.n238 2.19141
R704 a_n8964_8799.n309 a_n8964_8799.n308 2.19141
R705 a_n8964_8799.n288 a_n8964_8799.n287 2.19141
R706 a_n8964_8799.n42 a_n8964_8799.n35 2.19141
R707 a_n8964_8799.n66 a_n8964_8799.n65 2.19141
R708 a_n8964_8799.n90 a_n8964_8799.n83 2.19141
R709 a_n8964_8799.n114 a_n8964_8799.n113 2.19141
R710 a_n8964_8799.n139 a_n8964_8799.n132 2.19141
R711 a_n8964_8799.n163 a_n8964_8799.n162 2.19141
R712 a_n8964_8799.n205 a_n8964_8799.n204 0.730803
R713 a_n8964_8799.n198 a_n8964_8799.n197 0.730803
R714 a_n8964_8799.n253 a_n8964_8799.n252 0.730803
R715 a_n8964_8799.n246 a_n8964_8799.n245 0.730803
R716 a_n8964_8799.n302 a_n8964_8799.n301 0.730803
R717 a_n8964_8799.n295 a_n8964_8799.n294 0.730803
R718 a_n8964_8799.n52 a_n8964_8799.n33 0.730803
R719 a_n8964_8799.n59 a_n8964_8799.n58 0.730803
R720 a_n8964_8799.n100 a_n8964_8799.n81 0.730803
R721 a_n8964_8799.n107 a_n8964_8799.n106 0.730803
R722 a_n8964_8799.n149 a_n8964_8799.n130 0.730803
R723 a_n8964_8799.n156 a_n8964_8799.n155 0.730803
R724 a_n8964_8799.n324 a_n8964_8799.n322 0.444466
R725 a_n8964_8799.n329 a_n8964_8799.n327 0.444466
R726 a_n8964_8799.n331 a_n8964_8799.n329 0.444466
R727 a_n8964_8799.n338 a_n8964_8799.n2 0.444466
R728 a_n8964_8799.n336 a_n8964_8799.n334 0.444466
R729 a_n8964_8799.n18 a_n8964_8799.n16 0.358259
R730 a_n8964_8799.n20 a_n8964_8799.n18 0.358259
R731 a_n8964_8799.n22 a_n8964_8799.n20 0.358259
R732 a_n8964_8799.n24 a_n8964_8799.n22 0.358259
R733 a_n8964_8799.n13 a_n8964_8799.n11 0.358259
R734 a_n8964_8799.n11 a_n8964_8799.n9 0.358259
R735 a_n8964_8799.n9 a_n8964_8799.n7 0.358259
R736 a_n8964_8799.n7 a_n8964_8799.n5 0.358259
R737 a_n8964_8799.n325 a_n8964_8799.n324 0.222483
R738 a_n8964_8799.n327 a_n8964_8799.n325 0.222483
R739 a_n8964_8799.n338 a_n8964_8799.n337 0.222483
R740 a_n8964_8799.n337 a_n8964_8799.n336 0.222483
R741 a_n8964_8799.n219 a_n8964_8799.n172 0.189894
R742 a_n8964_8799.n215 a_n8964_8799.n172 0.189894
R743 a_n8964_8799.n215 a_n8964_8799.n214 0.189894
R744 a_n8964_8799.n214 a_n8964_8799.n213 0.189894
R745 a_n8964_8799.n213 a_n8964_8799.n174 0.189894
R746 a_n8964_8799.n175 a_n8964_8799.n174 0.189894
R747 a_n8964_8799.n208 a_n8964_8799.n175 0.189894
R748 a_n8964_8799.n208 a_n8964_8799.n207 0.189894
R749 a_n8964_8799.n207 a_n8964_8799.n206 0.189894
R750 a_n8964_8799.n206 a_n8964_8799.n177 0.189894
R751 a_n8964_8799.n178 a_n8964_8799.n177 0.189894
R752 a_n8964_8799.n201 a_n8964_8799.n178 0.189894
R753 a_n8964_8799.n201 a_n8964_8799.n200 0.189894
R754 a_n8964_8799.n200 a_n8964_8799.n199 0.189894
R755 a_n8964_8799.n199 a_n8964_8799.n180 0.189894
R756 a_n8964_8799.n181 a_n8964_8799.n180 0.189894
R757 a_n8964_8799.n194 a_n8964_8799.n181 0.189894
R758 a_n8964_8799.n194 a_n8964_8799.n193 0.189894
R759 a_n8964_8799.n193 a_n8964_8799.n192 0.189894
R760 a_n8964_8799.n192 a_n8964_8799.n183 0.189894
R761 a_n8964_8799.n184 a_n8964_8799.n183 0.189894
R762 a_n8964_8799.n187 a_n8964_8799.n184 0.189894
R763 a_n8964_8799.n267 a_n8964_8799.n220 0.189894
R764 a_n8964_8799.n263 a_n8964_8799.n220 0.189894
R765 a_n8964_8799.n263 a_n8964_8799.n262 0.189894
R766 a_n8964_8799.n262 a_n8964_8799.n261 0.189894
R767 a_n8964_8799.n261 a_n8964_8799.n222 0.189894
R768 a_n8964_8799.n223 a_n8964_8799.n222 0.189894
R769 a_n8964_8799.n256 a_n8964_8799.n223 0.189894
R770 a_n8964_8799.n256 a_n8964_8799.n255 0.189894
R771 a_n8964_8799.n255 a_n8964_8799.n254 0.189894
R772 a_n8964_8799.n254 a_n8964_8799.n225 0.189894
R773 a_n8964_8799.n226 a_n8964_8799.n225 0.189894
R774 a_n8964_8799.n249 a_n8964_8799.n226 0.189894
R775 a_n8964_8799.n249 a_n8964_8799.n248 0.189894
R776 a_n8964_8799.n248 a_n8964_8799.n247 0.189894
R777 a_n8964_8799.n247 a_n8964_8799.n228 0.189894
R778 a_n8964_8799.n229 a_n8964_8799.n228 0.189894
R779 a_n8964_8799.n242 a_n8964_8799.n229 0.189894
R780 a_n8964_8799.n242 a_n8964_8799.n241 0.189894
R781 a_n8964_8799.n241 a_n8964_8799.n240 0.189894
R782 a_n8964_8799.n240 a_n8964_8799.n231 0.189894
R783 a_n8964_8799.n232 a_n8964_8799.n231 0.189894
R784 a_n8964_8799.n235 a_n8964_8799.n232 0.189894
R785 a_n8964_8799.n316 a_n8964_8799.n269 0.189894
R786 a_n8964_8799.n312 a_n8964_8799.n269 0.189894
R787 a_n8964_8799.n312 a_n8964_8799.n311 0.189894
R788 a_n8964_8799.n311 a_n8964_8799.n310 0.189894
R789 a_n8964_8799.n310 a_n8964_8799.n271 0.189894
R790 a_n8964_8799.n272 a_n8964_8799.n271 0.189894
R791 a_n8964_8799.n305 a_n8964_8799.n272 0.189894
R792 a_n8964_8799.n305 a_n8964_8799.n304 0.189894
R793 a_n8964_8799.n304 a_n8964_8799.n303 0.189894
R794 a_n8964_8799.n303 a_n8964_8799.n274 0.189894
R795 a_n8964_8799.n275 a_n8964_8799.n274 0.189894
R796 a_n8964_8799.n298 a_n8964_8799.n275 0.189894
R797 a_n8964_8799.n298 a_n8964_8799.n297 0.189894
R798 a_n8964_8799.n297 a_n8964_8799.n296 0.189894
R799 a_n8964_8799.n296 a_n8964_8799.n277 0.189894
R800 a_n8964_8799.n278 a_n8964_8799.n277 0.189894
R801 a_n8964_8799.n291 a_n8964_8799.n278 0.189894
R802 a_n8964_8799.n291 a_n8964_8799.n290 0.189894
R803 a_n8964_8799.n290 a_n8964_8799.n289 0.189894
R804 a_n8964_8799.n289 a_n8964_8799.n280 0.189894
R805 a_n8964_8799.n281 a_n8964_8799.n280 0.189894
R806 a_n8964_8799.n284 a_n8964_8799.n281 0.189894
R807 a_n8964_8799.n39 a_n8964_8799.n36 0.189894
R808 a_n8964_8799.n43 a_n8964_8799.n36 0.189894
R809 a_n8964_8799.n44 a_n8964_8799.n43 0.189894
R810 a_n8964_8799.n45 a_n8964_8799.n44 0.189894
R811 a_n8964_8799.n45 a_n8964_8799.n34 0.189894
R812 a_n8964_8799.n49 a_n8964_8799.n34 0.189894
R813 a_n8964_8799.n50 a_n8964_8799.n49 0.189894
R814 a_n8964_8799.n51 a_n8964_8799.n50 0.189894
R815 a_n8964_8799.n51 a_n8964_8799.n32 0.189894
R816 a_n8964_8799.n55 a_n8964_8799.n32 0.189894
R817 a_n8964_8799.n56 a_n8964_8799.n55 0.189894
R818 a_n8964_8799.n57 a_n8964_8799.n56 0.189894
R819 a_n8964_8799.n57 a_n8964_8799.n30 0.189894
R820 a_n8964_8799.n61 a_n8964_8799.n30 0.189894
R821 a_n8964_8799.n62 a_n8964_8799.n61 0.189894
R822 a_n8964_8799.n63 a_n8964_8799.n62 0.189894
R823 a_n8964_8799.n63 a_n8964_8799.n28 0.189894
R824 a_n8964_8799.n67 a_n8964_8799.n28 0.189894
R825 a_n8964_8799.n68 a_n8964_8799.n67 0.189894
R826 a_n8964_8799.n69 a_n8964_8799.n68 0.189894
R827 a_n8964_8799.n69 a_n8964_8799.n26 0.189894
R828 a_n8964_8799.n73 a_n8964_8799.n26 0.189894
R829 a_n8964_8799.n87 a_n8964_8799.n84 0.189894
R830 a_n8964_8799.n91 a_n8964_8799.n84 0.189894
R831 a_n8964_8799.n92 a_n8964_8799.n91 0.189894
R832 a_n8964_8799.n93 a_n8964_8799.n92 0.189894
R833 a_n8964_8799.n93 a_n8964_8799.n82 0.189894
R834 a_n8964_8799.n97 a_n8964_8799.n82 0.189894
R835 a_n8964_8799.n98 a_n8964_8799.n97 0.189894
R836 a_n8964_8799.n99 a_n8964_8799.n98 0.189894
R837 a_n8964_8799.n99 a_n8964_8799.n80 0.189894
R838 a_n8964_8799.n103 a_n8964_8799.n80 0.189894
R839 a_n8964_8799.n104 a_n8964_8799.n103 0.189894
R840 a_n8964_8799.n105 a_n8964_8799.n104 0.189894
R841 a_n8964_8799.n105 a_n8964_8799.n78 0.189894
R842 a_n8964_8799.n109 a_n8964_8799.n78 0.189894
R843 a_n8964_8799.n110 a_n8964_8799.n109 0.189894
R844 a_n8964_8799.n111 a_n8964_8799.n110 0.189894
R845 a_n8964_8799.n111 a_n8964_8799.n76 0.189894
R846 a_n8964_8799.n115 a_n8964_8799.n76 0.189894
R847 a_n8964_8799.n116 a_n8964_8799.n115 0.189894
R848 a_n8964_8799.n117 a_n8964_8799.n116 0.189894
R849 a_n8964_8799.n117 a_n8964_8799.n74 0.189894
R850 a_n8964_8799.n121 a_n8964_8799.n74 0.189894
R851 a_n8964_8799.n136 a_n8964_8799.n133 0.189894
R852 a_n8964_8799.n140 a_n8964_8799.n133 0.189894
R853 a_n8964_8799.n141 a_n8964_8799.n140 0.189894
R854 a_n8964_8799.n142 a_n8964_8799.n141 0.189894
R855 a_n8964_8799.n142 a_n8964_8799.n131 0.189894
R856 a_n8964_8799.n146 a_n8964_8799.n131 0.189894
R857 a_n8964_8799.n147 a_n8964_8799.n146 0.189894
R858 a_n8964_8799.n148 a_n8964_8799.n147 0.189894
R859 a_n8964_8799.n148 a_n8964_8799.n129 0.189894
R860 a_n8964_8799.n152 a_n8964_8799.n129 0.189894
R861 a_n8964_8799.n153 a_n8964_8799.n152 0.189894
R862 a_n8964_8799.n154 a_n8964_8799.n153 0.189894
R863 a_n8964_8799.n154 a_n8964_8799.n127 0.189894
R864 a_n8964_8799.n158 a_n8964_8799.n127 0.189894
R865 a_n8964_8799.n159 a_n8964_8799.n158 0.189894
R866 a_n8964_8799.n160 a_n8964_8799.n159 0.189894
R867 a_n8964_8799.n160 a_n8964_8799.n125 0.189894
R868 a_n8964_8799.n164 a_n8964_8799.n125 0.189894
R869 a_n8964_8799.n165 a_n8964_8799.n164 0.189894
R870 a_n8964_8799.n166 a_n8964_8799.n165 0.189894
R871 a_n8964_8799.n166 a_n8964_8799.n123 0.189894
R872 a_n8964_8799.n170 a_n8964_8799.n123 0.189894
R873 gnd.n7183 gnd.n447 1638.19
R874 gnd.n6487 gnd.n5135 939.716
R875 gnd.n7577 gnd.n107 795.207
R876 gnd.n7741 gnd.n103 795.207
R877 gnd.n4476 gnd.n4475 795.207
R878 gnd.n1688 gnd.n1687 795.207
R879 gnd.n4896 gnd.n1324 795.207
R880 gnd.n3349 gnd.n1322 795.207
R881 gnd.n2958 gnd.n1008 795.207
R882 gnd.n3021 gnd.n2959 795.207
R883 gnd.n7739 gnd.n109 775.989
R884 gnd.n178 gnd.n105 775.989
R885 gnd.n1986 gnd.n1984 775.989
R886 gnd.n1909 gnd.n1482 775.989
R887 gnd.n4898 gnd.n1319 775.989
R888 gnd.n3535 gnd.n1321 775.989
R889 gnd.n5057 gnd.n5056 775.989
R890 gnd.n5133 gnd.n1012 775.989
R891 gnd.n967 gnd.n953 766.379
R892 gnd.n6403 gnd.n6402 766.379
R893 gnd.n5618 gnd.n5517 766.379
R894 gnd.n5616 gnd.n5519 766.379
R895 gnd.n6488 gnd.n958 756.769
R896 gnd.n6389 gnd.n6388 756.769
R897 gnd.n5750 gnd.n5479 756.769
R898 gnd.n5736 gnd.n5468 756.769
R899 gnd.n3395 gnd.n1329 711.122
R900 gnd.n4738 gnd.n1455 711.122
R901 gnd.n3278 gnd.n2725 711.122
R902 gnd.n1798 gnd.n1457 711.122
R903 gnd.n6691 gnd.n739 703.915
R904 gnd.n7182 gnd.n448 703.915
R905 gnd.n7395 gnd.n7394 703.915
R906 gnd.n2859 gnd.n2856 703.915
R907 gnd.n6691 gnd.n6690 585
R908 gnd.n6692 gnd.n6691 585
R909 gnd.n6689 gnd.n741 585
R910 gnd.n741 gnd.n740 585
R911 gnd.n6688 gnd.n6687 585
R912 gnd.n6687 gnd.n6686 585
R913 gnd.n746 gnd.n745 585
R914 gnd.n6685 gnd.n746 585
R915 gnd.n6683 gnd.n6682 585
R916 gnd.n6684 gnd.n6683 585
R917 gnd.n6681 gnd.n748 585
R918 gnd.n748 gnd.n747 585
R919 gnd.n6680 gnd.n6679 585
R920 gnd.n6679 gnd.n6678 585
R921 gnd.n754 gnd.n753 585
R922 gnd.n6677 gnd.n754 585
R923 gnd.n6675 gnd.n6674 585
R924 gnd.n6676 gnd.n6675 585
R925 gnd.n6673 gnd.n756 585
R926 gnd.n756 gnd.n755 585
R927 gnd.n6672 gnd.n6671 585
R928 gnd.n6671 gnd.n6670 585
R929 gnd.n762 gnd.n761 585
R930 gnd.n6669 gnd.n762 585
R931 gnd.n6667 gnd.n6666 585
R932 gnd.n6668 gnd.n6667 585
R933 gnd.n6665 gnd.n764 585
R934 gnd.n764 gnd.n763 585
R935 gnd.n6664 gnd.n6663 585
R936 gnd.n6663 gnd.n6662 585
R937 gnd.n770 gnd.n769 585
R938 gnd.n6661 gnd.n770 585
R939 gnd.n6659 gnd.n6658 585
R940 gnd.n6660 gnd.n6659 585
R941 gnd.n6657 gnd.n772 585
R942 gnd.n772 gnd.n771 585
R943 gnd.n6656 gnd.n6655 585
R944 gnd.n6655 gnd.n6654 585
R945 gnd.n778 gnd.n777 585
R946 gnd.n6653 gnd.n778 585
R947 gnd.n6651 gnd.n6650 585
R948 gnd.n6652 gnd.n6651 585
R949 gnd.n6649 gnd.n780 585
R950 gnd.n780 gnd.n779 585
R951 gnd.n6648 gnd.n6647 585
R952 gnd.n6647 gnd.n6646 585
R953 gnd.n786 gnd.n785 585
R954 gnd.n6645 gnd.n786 585
R955 gnd.n6643 gnd.n6642 585
R956 gnd.n6644 gnd.n6643 585
R957 gnd.n6641 gnd.n788 585
R958 gnd.n788 gnd.n787 585
R959 gnd.n6640 gnd.n6639 585
R960 gnd.n6639 gnd.n6638 585
R961 gnd.n794 gnd.n793 585
R962 gnd.n6637 gnd.n794 585
R963 gnd.n6635 gnd.n6634 585
R964 gnd.n6636 gnd.n6635 585
R965 gnd.n6633 gnd.n796 585
R966 gnd.n796 gnd.n795 585
R967 gnd.n6632 gnd.n6631 585
R968 gnd.n6631 gnd.n6630 585
R969 gnd.n802 gnd.n801 585
R970 gnd.n6629 gnd.n802 585
R971 gnd.n6627 gnd.n6626 585
R972 gnd.n6628 gnd.n6627 585
R973 gnd.n6625 gnd.n804 585
R974 gnd.n804 gnd.n803 585
R975 gnd.n6624 gnd.n6623 585
R976 gnd.n6623 gnd.n6622 585
R977 gnd.n810 gnd.n809 585
R978 gnd.n6621 gnd.n810 585
R979 gnd.n6619 gnd.n6618 585
R980 gnd.n6620 gnd.n6619 585
R981 gnd.n6617 gnd.n812 585
R982 gnd.n812 gnd.n811 585
R983 gnd.n6616 gnd.n6615 585
R984 gnd.n6615 gnd.n6614 585
R985 gnd.n818 gnd.n817 585
R986 gnd.n6613 gnd.n818 585
R987 gnd.n6611 gnd.n6610 585
R988 gnd.n6612 gnd.n6611 585
R989 gnd.n6609 gnd.n820 585
R990 gnd.n820 gnd.n819 585
R991 gnd.n6608 gnd.n6607 585
R992 gnd.n6607 gnd.n6606 585
R993 gnd.n826 gnd.n825 585
R994 gnd.n6605 gnd.n826 585
R995 gnd.n6603 gnd.n6602 585
R996 gnd.n6604 gnd.n6603 585
R997 gnd.n6601 gnd.n828 585
R998 gnd.n828 gnd.n827 585
R999 gnd.n6600 gnd.n6599 585
R1000 gnd.n6599 gnd.n6598 585
R1001 gnd.n834 gnd.n833 585
R1002 gnd.n6597 gnd.n834 585
R1003 gnd.n6595 gnd.n6594 585
R1004 gnd.n6596 gnd.n6595 585
R1005 gnd.n6593 gnd.n836 585
R1006 gnd.n836 gnd.n835 585
R1007 gnd.n6592 gnd.n6591 585
R1008 gnd.n6591 gnd.n6590 585
R1009 gnd.n842 gnd.n841 585
R1010 gnd.n6589 gnd.n842 585
R1011 gnd.n6587 gnd.n6586 585
R1012 gnd.n6588 gnd.n6587 585
R1013 gnd.n6585 gnd.n844 585
R1014 gnd.n844 gnd.n843 585
R1015 gnd.n6584 gnd.n6583 585
R1016 gnd.n6583 gnd.n6582 585
R1017 gnd.n850 gnd.n849 585
R1018 gnd.n6581 gnd.n850 585
R1019 gnd.n6579 gnd.n6578 585
R1020 gnd.n6580 gnd.n6579 585
R1021 gnd.n6577 gnd.n852 585
R1022 gnd.n852 gnd.n851 585
R1023 gnd.n6576 gnd.n6575 585
R1024 gnd.n6575 gnd.n6574 585
R1025 gnd.n858 gnd.n857 585
R1026 gnd.n6573 gnd.n858 585
R1027 gnd.n6571 gnd.n6570 585
R1028 gnd.n6572 gnd.n6571 585
R1029 gnd.n6569 gnd.n860 585
R1030 gnd.n860 gnd.n859 585
R1031 gnd.n6568 gnd.n6567 585
R1032 gnd.n6567 gnd.n6566 585
R1033 gnd.n866 gnd.n865 585
R1034 gnd.n6565 gnd.n866 585
R1035 gnd.n6563 gnd.n6562 585
R1036 gnd.n6564 gnd.n6563 585
R1037 gnd.n6561 gnd.n868 585
R1038 gnd.n868 gnd.n867 585
R1039 gnd.n6560 gnd.n6559 585
R1040 gnd.n6559 gnd.n6558 585
R1041 gnd.n874 gnd.n873 585
R1042 gnd.n6557 gnd.n874 585
R1043 gnd.n6555 gnd.n6554 585
R1044 gnd.n6556 gnd.n6555 585
R1045 gnd.n6553 gnd.n876 585
R1046 gnd.n876 gnd.n875 585
R1047 gnd.n6552 gnd.n6551 585
R1048 gnd.n6551 gnd.n6550 585
R1049 gnd.n882 gnd.n881 585
R1050 gnd.n6549 gnd.n882 585
R1051 gnd.n6547 gnd.n6546 585
R1052 gnd.n6548 gnd.n6547 585
R1053 gnd.n6545 gnd.n884 585
R1054 gnd.n884 gnd.n883 585
R1055 gnd.n6544 gnd.n6543 585
R1056 gnd.n6543 gnd.n6542 585
R1057 gnd.n890 gnd.n889 585
R1058 gnd.n6541 gnd.n890 585
R1059 gnd.n6539 gnd.n6538 585
R1060 gnd.n6540 gnd.n6539 585
R1061 gnd.n6537 gnd.n892 585
R1062 gnd.n892 gnd.n891 585
R1063 gnd.n6536 gnd.n6535 585
R1064 gnd.n6535 gnd.n6534 585
R1065 gnd.n898 gnd.n897 585
R1066 gnd.n6533 gnd.n898 585
R1067 gnd.n6531 gnd.n6530 585
R1068 gnd.n6532 gnd.n6531 585
R1069 gnd.n6529 gnd.n900 585
R1070 gnd.n900 gnd.n899 585
R1071 gnd.n6528 gnd.n6527 585
R1072 gnd.n6527 gnd.n6526 585
R1073 gnd.n906 gnd.n905 585
R1074 gnd.n6525 gnd.n906 585
R1075 gnd.n739 gnd.n738 585
R1076 gnd.n6693 gnd.n739 585
R1077 gnd.n6696 gnd.n6695 585
R1078 gnd.n6695 gnd.n6694 585
R1079 gnd.n736 gnd.n735 585
R1080 gnd.n735 gnd.n734 585
R1081 gnd.n6701 gnd.n6700 585
R1082 gnd.n6702 gnd.n6701 585
R1083 gnd.n733 gnd.n732 585
R1084 gnd.n6703 gnd.n733 585
R1085 gnd.n6706 gnd.n6705 585
R1086 gnd.n6705 gnd.n6704 585
R1087 gnd.n730 gnd.n729 585
R1088 gnd.n729 gnd.n728 585
R1089 gnd.n6711 gnd.n6710 585
R1090 gnd.n6712 gnd.n6711 585
R1091 gnd.n727 gnd.n726 585
R1092 gnd.n6713 gnd.n727 585
R1093 gnd.n6716 gnd.n6715 585
R1094 gnd.n6715 gnd.n6714 585
R1095 gnd.n724 gnd.n723 585
R1096 gnd.n723 gnd.n722 585
R1097 gnd.n6721 gnd.n6720 585
R1098 gnd.n6722 gnd.n6721 585
R1099 gnd.n721 gnd.n720 585
R1100 gnd.n6723 gnd.n721 585
R1101 gnd.n6726 gnd.n6725 585
R1102 gnd.n6725 gnd.n6724 585
R1103 gnd.n718 gnd.n717 585
R1104 gnd.n717 gnd.n716 585
R1105 gnd.n6731 gnd.n6730 585
R1106 gnd.n6732 gnd.n6731 585
R1107 gnd.n715 gnd.n714 585
R1108 gnd.n6733 gnd.n715 585
R1109 gnd.n6736 gnd.n6735 585
R1110 gnd.n6735 gnd.n6734 585
R1111 gnd.n712 gnd.n711 585
R1112 gnd.n711 gnd.n710 585
R1113 gnd.n6741 gnd.n6740 585
R1114 gnd.n6742 gnd.n6741 585
R1115 gnd.n709 gnd.n708 585
R1116 gnd.n6743 gnd.n709 585
R1117 gnd.n6746 gnd.n6745 585
R1118 gnd.n6745 gnd.n6744 585
R1119 gnd.n706 gnd.n705 585
R1120 gnd.n705 gnd.n704 585
R1121 gnd.n6751 gnd.n6750 585
R1122 gnd.n6752 gnd.n6751 585
R1123 gnd.n703 gnd.n702 585
R1124 gnd.n6753 gnd.n703 585
R1125 gnd.n6756 gnd.n6755 585
R1126 gnd.n6755 gnd.n6754 585
R1127 gnd.n700 gnd.n699 585
R1128 gnd.n699 gnd.n698 585
R1129 gnd.n6761 gnd.n6760 585
R1130 gnd.n6762 gnd.n6761 585
R1131 gnd.n697 gnd.n696 585
R1132 gnd.n6763 gnd.n697 585
R1133 gnd.n6766 gnd.n6765 585
R1134 gnd.n6765 gnd.n6764 585
R1135 gnd.n694 gnd.n693 585
R1136 gnd.n693 gnd.n692 585
R1137 gnd.n6771 gnd.n6770 585
R1138 gnd.n6772 gnd.n6771 585
R1139 gnd.n691 gnd.n690 585
R1140 gnd.n6773 gnd.n691 585
R1141 gnd.n6776 gnd.n6775 585
R1142 gnd.n6775 gnd.n6774 585
R1143 gnd.n688 gnd.n687 585
R1144 gnd.n687 gnd.n686 585
R1145 gnd.n6781 gnd.n6780 585
R1146 gnd.n6782 gnd.n6781 585
R1147 gnd.n685 gnd.n684 585
R1148 gnd.n6783 gnd.n685 585
R1149 gnd.n6786 gnd.n6785 585
R1150 gnd.n6785 gnd.n6784 585
R1151 gnd.n682 gnd.n681 585
R1152 gnd.n681 gnd.n680 585
R1153 gnd.n6791 gnd.n6790 585
R1154 gnd.n6792 gnd.n6791 585
R1155 gnd.n679 gnd.n678 585
R1156 gnd.n6793 gnd.n679 585
R1157 gnd.n6796 gnd.n6795 585
R1158 gnd.n6795 gnd.n6794 585
R1159 gnd.n676 gnd.n675 585
R1160 gnd.n675 gnd.n674 585
R1161 gnd.n6801 gnd.n6800 585
R1162 gnd.n6802 gnd.n6801 585
R1163 gnd.n673 gnd.n672 585
R1164 gnd.n6803 gnd.n673 585
R1165 gnd.n6806 gnd.n6805 585
R1166 gnd.n6805 gnd.n6804 585
R1167 gnd.n670 gnd.n669 585
R1168 gnd.n669 gnd.n668 585
R1169 gnd.n6811 gnd.n6810 585
R1170 gnd.n6812 gnd.n6811 585
R1171 gnd.n667 gnd.n666 585
R1172 gnd.n6813 gnd.n667 585
R1173 gnd.n6816 gnd.n6815 585
R1174 gnd.n6815 gnd.n6814 585
R1175 gnd.n664 gnd.n663 585
R1176 gnd.n663 gnd.n662 585
R1177 gnd.n6821 gnd.n6820 585
R1178 gnd.n6822 gnd.n6821 585
R1179 gnd.n661 gnd.n660 585
R1180 gnd.n6823 gnd.n661 585
R1181 gnd.n6826 gnd.n6825 585
R1182 gnd.n6825 gnd.n6824 585
R1183 gnd.n658 gnd.n657 585
R1184 gnd.n657 gnd.n656 585
R1185 gnd.n6831 gnd.n6830 585
R1186 gnd.n6832 gnd.n6831 585
R1187 gnd.n655 gnd.n654 585
R1188 gnd.n6833 gnd.n655 585
R1189 gnd.n6836 gnd.n6835 585
R1190 gnd.n6835 gnd.n6834 585
R1191 gnd.n652 gnd.n651 585
R1192 gnd.n651 gnd.n650 585
R1193 gnd.n6841 gnd.n6840 585
R1194 gnd.n6842 gnd.n6841 585
R1195 gnd.n649 gnd.n648 585
R1196 gnd.n6843 gnd.n649 585
R1197 gnd.n6846 gnd.n6845 585
R1198 gnd.n6845 gnd.n6844 585
R1199 gnd.n646 gnd.n645 585
R1200 gnd.n645 gnd.n644 585
R1201 gnd.n6851 gnd.n6850 585
R1202 gnd.n6852 gnd.n6851 585
R1203 gnd.n643 gnd.n642 585
R1204 gnd.n6853 gnd.n643 585
R1205 gnd.n6856 gnd.n6855 585
R1206 gnd.n6855 gnd.n6854 585
R1207 gnd.n640 gnd.n639 585
R1208 gnd.n639 gnd.n638 585
R1209 gnd.n6861 gnd.n6860 585
R1210 gnd.n6862 gnd.n6861 585
R1211 gnd.n637 gnd.n636 585
R1212 gnd.n6863 gnd.n637 585
R1213 gnd.n6866 gnd.n6865 585
R1214 gnd.n6865 gnd.n6864 585
R1215 gnd.n634 gnd.n633 585
R1216 gnd.n633 gnd.n632 585
R1217 gnd.n6871 gnd.n6870 585
R1218 gnd.n6872 gnd.n6871 585
R1219 gnd.n631 gnd.n630 585
R1220 gnd.n6873 gnd.n631 585
R1221 gnd.n6876 gnd.n6875 585
R1222 gnd.n6875 gnd.n6874 585
R1223 gnd.n628 gnd.n627 585
R1224 gnd.n627 gnd.n626 585
R1225 gnd.n6881 gnd.n6880 585
R1226 gnd.n6882 gnd.n6881 585
R1227 gnd.n625 gnd.n624 585
R1228 gnd.n6883 gnd.n625 585
R1229 gnd.n6886 gnd.n6885 585
R1230 gnd.n6885 gnd.n6884 585
R1231 gnd.n622 gnd.n621 585
R1232 gnd.n621 gnd.n620 585
R1233 gnd.n6891 gnd.n6890 585
R1234 gnd.n6892 gnd.n6891 585
R1235 gnd.n619 gnd.n618 585
R1236 gnd.n6893 gnd.n619 585
R1237 gnd.n6896 gnd.n6895 585
R1238 gnd.n6895 gnd.n6894 585
R1239 gnd.n616 gnd.n615 585
R1240 gnd.n615 gnd.n614 585
R1241 gnd.n6901 gnd.n6900 585
R1242 gnd.n6902 gnd.n6901 585
R1243 gnd.n613 gnd.n612 585
R1244 gnd.n6903 gnd.n613 585
R1245 gnd.n6906 gnd.n6905 585
R1246 gnd.n6905 gnd.n6904 585
R1247 gnd.n610 gnd.n609 585
R1248 gnd.n609 gnd.n608 585
R1249 gnd.n6911 gnd.n6910 585
R1250 gnd.n6912 gnd.n6911 585
R1251 gnd.n607 gnd.n606 585
R1252 gnd.n6913 gnd.n607 585
R1253 gnd.n6916 gnd.n6915 585
R1254 gnd.n6915 gnd.n6914 585
R1255 gnd.n604 gnd.n603 585
R1256 gnd.n603 gnd.n602 585
R1257 gnd.n6921 gnd.n6920 585
R1258 gnd.n6922 gnd.n6921 585
R1259 gnd.n601 gnd.n600 585
R1260 gnd.n6923 gnd.n601 585
R1261 gnd.n6926 gnd.n6925 585
R1262 gnd.n6925 gnd.n6924 585
R1263 gnd.n598 gnd.n597 585
R1264 gnd.n597 gnd.n596 585
R1265 gnd.n6931 gnd.n6930 585
R1266 gnd.n6932 gnd.n6931 585
R1267 gnd.n595 gnd.n594 585
R1268 gnd.n6933 gnd.n595 585
R1269 gnd.n6936 gnd.n6935 585
R1270 gnd.n6935 gnd.n6934 585
R1271 gnd.n592 gnd.n591 585
R1272 gnd.n591 gnd.n590 585
R1273 gnd.n6941 gnd.n6940 585
R1274 gnd.n6942 gnd.n6941 585
R1275 gnd.n589 gnd.n588 585
R1276 gnd.n6943 gnd.n589 585
R1277 gnd.n6946 gnd.n6945 585
R1278 gnd.n6945 gnd.n6944 585
R1279 gnd.n586 gnd.n585 585
R1280 gnd.n585 gnd.n584 585
R1281 gnd.n6951 gnd.n6950 585
R1282 gnd.n6952 gnd.n6951 585
R1283 gnd.n583 gnd.n582 585
R1284 gnd.n6953 gnd.n583 585
R1285 gnd.n6956 gnd.n6955 585
R1286 gnd.n6955 gnd.n6954 585
R1287 gnd.n580 gnd.n579 585
R1288 gnd.n579 gnd.n578 585
R1289 gnd.n6961 gnd.n6960 585
R1290 gnd.n6962 gnd.n6961 585
R1291 gnd.n577 gnd.n576 585
R1292 gnd.n6963 gnd.n577 585
R1293 gnd.n6966 gnd.n6965 585
R1294 gnd.n6965 gnd.n6964 585
R1295 gnd.n574 gnd.n573 585
R1296 gnd.n573 gnd.n572 585
R1297 gnd.n6971 gnd.n6970 585
R1298 gnd.n6972 gnd.n6971 585
R1299 gnd.n571 gnd.n570 585
R1300 gnd.n6973 gnd.n571 585
R1301 gnd.n6976 gnd.n6975 585
R1302 gnd.n6975 gnd.n6974 585
R1303 gnd.n568 gnd.n567 585
R1304 gnd.n567 gnd.n566 585
R1305 gnd.n6981 gnd.n6980 585
R1306 gnd.n6982 gnd.n6981 585
R1307 gnd.n565 gnd.n564 585
R1308 gnd.n6983 gnd.n565 585
R1309 gnd.n6986 gnd.n6985 585
R1310 gnd.n6985 gnd.n6984 585
R1311 gnd.n562 gnd.n561 585
R1312 gnd.n561 gnd.n560 585
R1313 gnd.n6991 gnd.n6990 585
R1314 gnd.n6992 gnd.n6991 585
R1315 gnd.n559 gnd.n558 585
R1316 gnd.n6993 gnd.n559 585
R1317 gnd.n6996 gnd.n6995 585
R1318 gnd.n6995 gnd.n6994 585
R1319 gnd.n556 gnd.n555 585
R1320 gnd.n555 gnd.n554 585
R1321 gnd.n7001 gnd.n7000 585
R1322 gnd.n7002 gnd.n7001 585
R1323 gnd.n553 gnd.n552 585
R1324 gnd.n7003 gnd.n553 585
R1325 gnd.n7006 gnd.n7005 585
R1326 gnd.n7005 gnd.n7004 585
R1327 gnd.n550 gnd.n549 585
R1328 gnd.n549 gnd.n548 585
R1329 gnd.n7011 gnd.n7010 585
R1330 gnd.n7012 gnd.n7011 585
R1331 gnd.n547 gnd.n546 585
R1332 gnd.n7013 gnd.n547 585
R1333 gnd.n7016 gnd.n7015 585
R1334 gnd.n7015 gnd.n7014 585
R1335 gnd.n544 gnd.n543 585
R1336 gnd.n543 gnd.n542 585
R1337 gnd.n7021 gnd.n7020 585
R1338 gnd.n7022 gnd.n7021 585
R1339 gnd.n541 gnd.n540 585
R1340 gnd.n7023 gnd.n541 585
R1341 gnd.n7026 gnd.n7025 585
R1342 gnd.n7025 gnd.n7024 585
R1343 gnd.n538 gnd.n537 585
R1344 gnd.n537 gnd.n536 585
R1345 gnd.n7031 gnd.n7030 585
R1346 gnd.n7032 gnd.n7031 585
R1347 gnd.n535 gnd.n534 585
R1348 gnd.n7033 gnd.n535 585
R1349 gnd.n7036 gnd.n7035 585
R1350 gnd.n7035 gnd.n7034 585
R1351 gnd.n532 gnd.n531 585
R1352 gnd.n531 gnd.n530 585
R1353 gnd.n7041 gnd.n7040 585
R1354 gnd.n7042 gnd.n7041 585
R1355 gnd.n529 gnd.n528 585
R1356 gnd.n7043 gnd.n529 585
R1357 gnd.n7046 gnd.n7045 585
R1358 gnd.n7045 gnd.n7044 585
R1359 gnd.n526 gnd.n525 585
R1360 gnd.n525 gnd.n524 585
R1361 gnd.n7051 gnd.n7050 585
R1362 gnd.n7052 gnd.n7051 585
R1363 gnd.n523 gnd.n522 585
R1364 gnd.n7053 gnd.n523 585
R1365 gnd.n7056 gnd.n7055 585
R1366 gnd.n7055 gnd.n7054 585
R1367 gnd.n520 gnd.n519 585
R1368 gnd.n519 gnd.n518 585
R1369 gnd.n7061 gnd.n7060 585
R1370 gnd.n7062 gnd.n7061 585
R1371 gnd.n517 gnd.n516 585
R1372 gnd.n7063 gnd.n517 585
R1373 gnd.n7066 gnd.n7065 585
R1374 gnd.n7065 gnd.n7064 585
R1375 gnd.n514 gnd.n513 585
R1376 gnd.n513 gnd.n512 585
R1377 gnd.n7071 gnd.n7070 585
R1378 gnd.n7072 gnd.n7071 585
R1379 gnd.n511 gnd.n510 585
R1380 gnd.n7073 gnd.n511 585
R1381 gnd.n7076 gnd.n7075 585
R1382 gnd.n7075 gnd.n7074 585
R1383 gnd.n508 gnd.n507 585
R1384 gnd.n507 gnd.n506 585
R1385 gnd.n7081 gnd.n7080 585
R1386 gnd.n7082 gnd.n7081 585
R1387 gnd.n505 gnd.n504 585
R1388 gnd.n7083 gnd.n505 585
R1389 gnd.n7086 gnd.n7085 585
R1390 gnd.n7085 gnd.n7084 585
R1391 gnd.n502 gnd.n501 585
R1392 gnd.n501 gnd.n500 585
R1393 gnd.n7091 gnd.n7090 585
R1394 gnd.n7092 gnd.n7091 585
R1395 gnd.n499 gnd.n498 585
R1396 gnd.n7093 gnd.n499 585
R1397 gnd.n7096 gnd.n7095 585
R1398 gnd.n7095 gnd.n7094 585
R1399 gnd.n496 gnd.n495 585
R1400 gnd.n495 gnd.n494 585
R1401 gnd.n7101 gnd.n7100 585
R1402 gnd.n7102 gnd.n7101 585
R1403 gnd.n493 gnd.n492 585
R1404 gnd.n7103 gnd.n493 585
R1405 gnd.n7106 gnd.n7105 585
R1406 gnd.n7105 gnd.n7104 585
R1407 gnd.n490 gnd.n489 585
R1408 gnd.n489 gnd.n488 585
R1409 gnd.n7111 gnd.n7110 585
R1410 gnd.n7112 gnd.n7111 585
R1411 gnd.n487 gnd.n486 585
R1412 gnd.n7113 gnd.n487 585
R1413 gnd.n7116 gnd.n7115 585
R1414 gnd.n7115 gnd.n7114 585
R1415 gnd.n484 gnd.n483 585
R1416 gnd.n483 gnd.n482 585
R1417 gnd.n7121 gnd.n7120 585
R1418 gnd.n7122 gnd.n7121 585
R1419 gnd.n481 gnd.n480 585
R1420 gnd.n7123 gnd.n481 585
R1421 gnd.n7126 gnd.n7125 585
R1422 gnd.n7125 gnd.n7124 585
R1423 gnd.n478 gnd.n477 585
R1424 gnd.n477 gnd.n476 585
R1425 gnd.n7131 gnd.n7130 585
R1426 gnd.n7132 gnd.n7131 585
R1427 gnd.n475 gnd.n474 585
R1428 gnd.n7133 gnd.n475 585
R1429 gnd.n7136 gnd.n7135 585
R1430 gnd.n7135 gnd.n7134 585
R1431 gnd.n472 gnd.n471 585
R1432 gnd.n471 gnd.n470 585
R1433 gnd.n7141 gnd.n7140 585
R1434 gnd.n7142 gnd.n7141 585
R1435 gnd.n469 gnd.n468 585
R1436 gnd.n7143 gnd.n469 585
R1437 gnd.n7146 gnd.n7145 585
R1438 gnd.n7145 gnd.n7144 585
R1439 gnd.n466 gnd.n465 585
R1440 gnd.n465 gnd.n464 585
R1441 gnd.n7151 gnd.n7150 585
R1442 gnd.n7152 gnd.n7151 585
R1443 gnd.n463 gnd.n462 585
R1444 gnd.n7153 gnd.n463 585
R1445 gnd.n7156 gnd.n7155 585
R1446 gnd.n7155 gnd.n7154 585
R1447 gnd.n460 gnd.n459 585
R1448 gnd.n459 gnd.n458 585
R1449 gnd.n7161 gnd.n7160 585
R1450 gnd.n7162 gnd.n7161 585
R1451 gnd.n457 gnd.n456 585
R1452 gnd.n7163 gnd.n457 585
R1453 gnd.n7166 gnd.n7165 585
R1454 gnd.n7165 gnd.n7164 585
R1455 gnd.n454 gnd.n453 585
R1456 gnd.n453 gnd.n452 585
R1457 gnd.n7172 gnd.n7171 585
R1458 gnd.n7173 gnd.n7172 585
R1459 gnd.n451 gnd.n450 585
R1460 gnd.n7174 gnd.n451 585
R1461 gnd.n7177 gnd.n7176 585
R1462 gnd.n7176 gnd.n7175 585
R1463 gnd.n7178 gnd.n448 585
R1464 gnd.n448 gnd.n447 585
R1465 gnd.n323 gnd.n322 585
R1466 gnd.n7385 gnd.n322 585
R1467 gnd.n7388 gnd.n7387 585
R1468 gnd.n7387 gnd.n7386 585
R1469 gnd.n326 gnd.n325 585
R1470 gnd.n7384 gnd.n326 585
R1471 gnd.n7382 gnd.n7381 585
R1472 gnd.n7383 gnd.n7382 585
R1473 gnd.n329 gnd.n328 585
R1474 gnd.n328 gnd.n327 585
R1475 gnd.n7377 gnd.n7376 585
R1476 gnd.n7376 gnd.n7375 585
R1477 gnd.n332 gnd.n331 585
R1478 gnd.n7374 gnd.n332 585
R1479 gnd.n7372 gnd.n7371 585
R1480 gnd.n7373 gnd.n7372 585
R1481 gnd.n335 gnd.n334 585
R1482 gnd.n334 gnd.n333 585
R1483 gnd.n7367 gnd.n7366 585
R1484 gnd.n7366 gnd.n7365 585
R1485 gnd.n338 gnd.n337 585
R1486 gnd.n7364 gnd.n338 585
R1487 gnd.n7362 gnd.n7361 585
R1488 gnd.n7363 gnd.n7362 585
R1489 gnd.n341 gnd.n340 585
R1490 gnd.n340 gnd.n339 585
R1491 gnd.n7357 gnd.n7356 585
R1492 gnd.n7356 gnd.n7355 585
R1493 gnd.n344 gnd.n343 585
R1494 gnd.n7354 gnd.n344 585
R1495 gnd.n7352 gnd.n7351 585
R1496 gnd.n7353 gnd.n7352 585
R1497 gnd.n347 gnd.n346 585
R1498 gnd.n346 gnd.n345 585
R1499 gnd.n7347 gnd.n7346 585
R1500 gnd.n7346 gnd.n7345 585
R1501 gnd.n350 gnd.n349 585
R1502 gnd.n7344 gnd.n350 585
R1503 gnd.n7342 gnd.n7341 585
R1504 gnd.n7343 gnd.n7342 585
R1505 gnd.n353 gnd.n352 585
R1506 gnd.n352 gnd.n351 585
R1507 gnd.n7337 gnd.n7336 585
R1508 gnd.n7336 gnd.n7335 585
R1509 gnd.n356 gnd.n355 585
R1510 gnd.n7334 gnd.n356 585
R1511 gnd.n7332 gnd.n7331 585
R1512 gnd.n7333 gnd.n7332 585
R1513 gnd.n359 gnd.n358 585
R1514 gnd.n358 gnd.n357 585
R1515 gnd.n7327 gnd.n7326 585
R1516 gnd.n7326 gnd.n7325 585
R1517 gnd.n362 gnd.n361 585
R1518 gnd.n7324 gnd.n362 585
R1519 gnd.n7322 gnd.n7321 585
R1520 gnd.n7323 gnd.n7322 585
R1521 gnd.n365 gnd.n364 585
R1522 gnd.n364 gnd.n363 585
R1523 gnd.n7317 gnd.n7316 585
R1524 gnd.n7316 gnd.n7315 585
R1525 gnd.n368 gnd.n367 585
R1526 gnd.n7314 gnd.n368 585
R1527 gnd.n7312 gnd.n7311 585
R1528 gnd.n7313 gnd.n7312 585
R1529 gnd.n371 gnd.n370 585
R1530 gnd.n370 gnd.n369 585
R1531 gnd.n7307 gnd.n7306 585
R1532 gnd.n7306 gnd.n7305 585
R1533 gnd.n374 gnd.n373 585
R1534 gnd.n7304 gnd.n374 585
R1535 gnd.n7302 gnd.n7301 585
R1536 gnd.n7303 gnd.n7302 585
R1537 gnd.n377 gnd.n376 585
R1538 gnd.n376 gnd.n375 585
R1539 gnd.n7297 gnd.n7296 585
R1540 gnd.n7296 gnd.n7295 585
R1541 gnd.n380 gnd.n379 585
R1542 gnd.n7294 gnd.n380 585
R1543 gnd.n7292 gnd.n7291 585
R1544 gnd.n7293 gnd.n7292 585
R1545 gnd.n383 gnd.n382 585
R1546 gnd.n382 gnd.n381 585
R1547 gnd.n7287 gnd.n7286 585
R1548 gnd.n7286 gnd.n7285 585
R1549 gnd.n386 gnd.n385 585
R1550 gnd.n7284 gnd.n386 585
R1551 gnd.n7282 gnd.n7281 585
R1552 gnd.n7283 gnd.n7282 585
R1553 gnd.n389 gnd.n388 585
R1554 gnd.n388 gnd.n387 585
R1555 gnd.n7277 gnd.n7276 585
R1556 gnd.n7276 gnd.n7275 585
R1557 gnd.n392 gnd.n391 585
R1558 gnd.n7274 gnd.n392 585
R1559 gnd.n7272 gnd.n7271 585
R1560 gnd.n7273 gnd.n7272 585
R1561 gnd.n395 gnd.n394 585
R1562 gnd.n394 gnd.n393 585
R1563 gnd.n7267 gnd.n7266 585
R1564 gnd.n7266 gnd.n7265 585
R1565 gnd.n398 gnd.n397 585
R1566 gnd.n7264 gnd.n398 585
R1567 gnd.n7262 gnd.n7261 585
R1568 gnd.n7263 gnd.n7262 585
R1569 gnd.n401 gnd.n400 585
R1570 gnd.n400 gnd.n399 585
R1571 gnd.n7257 gnd.n7256 585
R1572 gnd.n7256 gnd.n7255 585
R1573 gnd.n404 gnd.n403 585
R1574 gnd.n7254 gnd.n404 585
R1575 gnd.n7252 gnd.n7251 585
R1576 gnd.n7253 gnd.n7252 585
R1577 gnd.n407 gnd.n406 585
R1578 gnd.n406 gnd.n405 585
R1579 gnd.n7247 gnd.n7246 585
R1580 gnd.n7246 gnd.n7245 585
R1581 gnd.n410 gnd.n409 585
R1582 gnd.n7244 gnd.n410 585
R1583 gnd.n7242 gnd.n7241 585
R1584 gnd.n7243 gnd.n7242 585
R1585 gnd.n413 gnd.n412 585
R1586 gnd.n412 gnd.n411 585
R1587 gnd.n7237 gnd.n7236 585
R1588 gnd.n7236 gnd.n7235 585
R1589 gnd.n416 gnd.n415 585
R1590 gnd.n7234 gnd.n416 585
R1591 gnd.n7232 gnd.n7231 585
R1592 gnd.n7233 gnd.n7232 585
R1593 gnd.n419 gnd.n418 585
R1594 gnd.n418 gnd.n417 585
R1595 gnd.n7227 gnd.n7226 585
R1596 gnd.n7226 gnd.n7225 585
R1597 gnd.n422 gnd.n421 585
R1598 gnd.n7224 gnd.n422 585
R1599 gnd.n7222 gnd.n7221 585
R1600 gnd.n7223 gnd.n7222 585
R1601 gnd.n425 gnd.n424 585
R1602 gnd.n424 gnd.n423 585
R1603 gnd.n7217 gnd.n7216 585
R1604 gnd.n7216 gnd.n7215 585
R1605 gnd.n428 gnd.n427 585
R1606 gnd.n7214 gnd.n428 585
R1607 gnd.n7212 gnd.n7211 585
R1608 gnd.n7213 gnd.n7212 585
R1609 gnd.n431 gnd.n430 585
R1610 gnd.n430 gnd.n429 585
R1611 gnd.n7207 gnd.n7206 585
R1612 gnd.n7206 gnd.n7205 585
R1613 gnd.n434 gnd.n433 585
R1614 gnd.n7204 gnd.n434 585
R1615 gnd.n7202 gnd.n7201 585
R1616 gnd.n7203 gnd.n7202 585
R1617 gnd.n437 gnd.n436 585
R1618 gnd.n436 gnd.n435 585
R1619 gnd.n7197 gnd.n7196 585
R1620 gnd.n7196 gnd.n7195 585
R1621 gnd.n440 gnd.n439 585
R1622 gnd.n7194 gnd.n440 585
R1623 gnd.n7192 gnd.n7191 585
R1624 gnd.n7193 gnd.n7192 585
R1625 gnd.n443 gnd.n442 585
R1626 gnd.n442 gnd.n441 585
R1627 gnd.n7187 gnd.n7186 585
R1628 gnd.n7186 gnd.n7185 585
R1629 gnd.n446 gnd.n445 585
R1630 gnd.n7184 gnd.n446 585
R1631 gnd.n7182 gnd.n7181 585
R1632 gnd.n7183 gnd.n7182 585
R1633 gnd.n4896 gnd.n4895 585
R1634 gnd.n4897 gnd.n4896 585
R1635 gnd.n1310 gnd.n1309 585
R1636 gnd.n3528 gnd.n1310 585
R1637 gnd.n4905 gnd.n4904 585
R1638 gnd.n4904 gnd.n4903 585
R1639 gnd.n4906 gnd.n1304 585
R1640 gnd.n3223 gnd.n1304 585
R1641 gnd.n4908 gnd.n4907 585
R1642 gnd.n4909 gnd.n4908 585
R1643 gnd.n1288 gnd.n1287 585
R1644 gnd.n3214 gnd.n1288 585
R1645 gnd.n4917 gnd.n4916 585
R1646 gnd.n4916 gnd.n4915 585
R1647 gnd.n4918 gnd.n1282 585
R1648 gnd.n3210 gnd.n1282 585
R1649 gnd.n4920 gnd.n4919 585
R1650 gnd.n4921 gnd.n4920 585
R1651 gnd.n1267 gnd.n1266 585
R1652 gnd.n3237 gnd.n1267 585
R1653 gnd.n4929 gnd.n4928 585
R1654 gnd.n4928 gnd.n4927 585
R1655 gnd.n4930 gnd.n1261 585
R1656 gnd.n3202 gnd.n1261 585
R1657 gnd.n4932 gnd.n4931 585
R1658 gnd.n4933 gnd.n4932 585
R1659 gnd.n1246 gnd.n1245 585
R1660 gnd.n3194 gnd.n1246 585
R1661 gnd.n4941 gnd.n4940 585
R1662 gnd.n4940 gnd.n4939 585
R1663 gnd.n4942 gnd.n1240 585
R1664 gnd.n3185 gnd.n1240 585
R1665 gnd.n4944 gnd.n4943 585
R1666 gnd.n4945 gnd.n4944 585
R1667 gnd.n1225 gnd.n1224 585
R1668 gnd.n3177 gnd.n1225 585
R1669 gnd.n4953 gnd.n4952 585
R1670 gnd.n4952 gnd.n4951 585
R1671 gnd.n4954 gnd.n1219 585
R1672 gnd.n3169 gnd.n1219 585
R1673 gnd.n4956 gnd.n4955 585
R1674 gnd.n4957 gnd.n4956 585
R1675 gnd.n1205 gnd.n1204 585
R1676 gnd.n3161 gnd.n1205 585
R1677 gnd.n4965 gnd.n4964 585
R1678 gnd.n4964 gnd.n4963 585
R1679 gnd.n4966 gnd.n1199 585
R1680 gnd.n3153 gnd.n1199 585
R1681 gnd.n4968 gnd.n4967 585
R1682 gnd.n4969 gnd.n4968 585
R1683 gnd.n1187 gnd.n1186 585
R1684 gnd.n3145 gnd.n1187 585
R1685 gnd.n4978 gnd.n4977 585
R1686 gnd.n4977 gnd.n4976 585
R1687 gnd.n4979 gnd.n1181 585
R1688 gnd.n3136 gnd.n1181 585
R1689 gnd.n4981 gnd.n4980 585
R1690 gnd.n4982 gnd.n4981 585
R1691 gnd.n1168 gnd.n1167 585
R1692 gnd.n3127 gnd.n1168 585
R1693 gnd.n4990 gnd.n4989 585
R1694 gnd.n4989 gnd.n4988 585
R1695 gnd.n4991 gnd.n1162 585
R1696 gnd.n3119 gnd.n1162 585
R1697 gnd.n4993 gnd.n4992 585
R1698 gnd.n4994 gnd.n4993 585
R1699 gnd.n1147 gnd.n1146 585
R1700 gnd.n3111 gnd.n1147 585
R1701 gnd.n5002 gnd.n5001 585
R1702 gnd.n5001 gnd.n5000 585
R1703 gnd.n5003 gnd.n1141 585
R1704 gnd.n3103 gnd.n1141 585
R1705 gnd.n5005 gnd.n5004 585
R1706 gnd.n5006 gnd.n5005 585
R1707 gnd.n1126 gnd.n1125 585
R1708 gnd.n3095 gnd.n1126 585
R1709 gnd.n5014 gnd.n5013 585
R1710 gnd.n5013 gnd.n5012 585
R1711 gnd.n5015 gnd.n1120 585
R1712 gnd.n3087 gnd.n1120 585
R1713 gnd.n5017 gnd.n5016 585
R1714 gnd.n5018 gnd.n5017 585
R1715 gnd.n1104 gnd.n1103 585
R1716 gnd.n3079 gnd.n1104 585
R1717 gnd.n5026 gnd.n5025 585
R1718 gnd.n5025 gnd.n5024 585
R1719 gnd.n5027 gnd.n1098 585
R1720 gnd.n1105 gnd.n1098 585
R1721 gnd.n5029 gnd.n5028 585
R1722 gnd.n5030 gnd.n5029 585
R1723 gnd.n1085 gnd.n1084 585
R1724 gnd.n1088 gnd.n1085 585
R1725 gnd.n5038 gnd.n5037 585
R1726 gnd.n5037 gnd.n5036 585
R1727 gnd.n5039 gnd.n1079 585
R1728 gnd.n1079 gnd.n1077 585
R1729 gnd.n5041 gnd.n5040 585
R1730 gnd.n5042 gnd.n5041 585
R1731 gnd.n1080 gnd.n1078 585
R1732 gnd.n1078 gnd.n1065 585
R1733 gnd.n3026 gnd.n1066 585
R1734 gnd.n5048 gnd.n1066 585
R1735 gnd.n2962 gnd.n2960 585
R1736 gnd.n2960 gnd.n1063 585
R1737 gnd.n3031 gnd.n3030 585
R1738 gnd.n3038 gnd.n3031 585
R1739 gnd.n2961 gnd.n2959 585
R1740 gnd.n2959 gnd.n1009 585
R1741 gnd.n3022 gnd.n3021 585
R1742 gnd.n3020 gnd.n3019 585
R1743 gnd.n3018 gnd.n3017 585
R1744 gnd.n3016 gnd.n3015 585
R1745 gnd.n3014 gnd.n3013 585
R1746 gnd.n3012 gnd.n3011 585
R1747 gnd.n3010 gnd.n3009 585
R1748 gnd.n3008 gnd.n3007 585
R1749 gnd.n3006 gnd.n3005 585
R1750 gnd.n3004 gnd.n3003 585
R1751 gnd.n3002 gnd.n3001 585
R1752 gnd.n3000 gnd.n2999 585
R1753 gnd.n2998 gnd.n2997 585
R1754 gnd.n2996 gnd.n2995 585
R1755 gnd.n2994 gnd.n2993 585
R1756 gnd.n2992 gnd.n2991 585
R1757 gnd.n2990 gnd.n2989 585
R1758 gnd.n2981 gnd.n2978 585
R1759 gnd.n2985 gnd.n1008 585
R1760 gnd.n5135 gnd.n1008 585
R1761 gnd.n3350 gnd.n3349 585
R1762 gnd.n3347 gnd.n3341 585
R1763 gnd.n3357 gnd.n3338 585
R1764 gnd.n3358 gnd.n3336 585
R1765 gnd.n3335 gnd.n3328 585
R1766 gnd.n3365 gnd.n3327 585
R1767 gnd.n3366 gnd.n3326 585
R1768 gnd.n3324 gnd.n3316 585
R1769 gnd.n3373 gnd.n3315 585
R1770 gnd.n3374 gnd.n3313 585
R1771 gnd.n3312 gnd.n3305 585
R1772 gnd.n3381 gnd.n3304 585
R1773 gnd.n3382 gnd.n3303 585
R1774 gnd.n3301 gnd.n3294 585
R1775 gnd.n3389 gnd.n3293 585
R1776 gnd.n3390 gnd.n3291 585
R1777 gnd.n3290 gnd.n3286 585
R1778 gnd.n3288 gnd.n3287 585
R1779 gnd.n1326 gnd.n1324 585
R1780 gnd.n2666 gnd.n1324 585
R1781 gnd.n2703 gnd.n1322 585
R1782 gnd.n4897 gnd.n1322 585
R1783 gnd.n3527 gnd.n3526 585
R1784 gnd.n3528 gnd.n3527 585
R1785 gnd.n2702 gnd.n1313 585
R1786 gnd.n4903 gnd.n1313 585
R1787 gnd.n3225 gnd.n3224 585
R1788 gnd.n3224 gnd.n3223 585
R1789 gnd.n2801 gnd.n1302 585
R1790 gnd.n4909 gnd.n1302 585
R1791 gnd.n3229 gnd.n2800 585
R1792 gnd.n3214 gnd.n2800 585
R1793 gnd.n3230 gnd.n1291 585
R1794 gnd.n4915 gnd.n1291 585
R1795 gnd.n3231 gnd.n2799 585
R1796 gnd.n3210 gnd.n2799 585
R1797 gnd.n2796 gnd.n1280 585
R1798 gnd.n4921 gnd.n1280 585
R1799 gnd.n3236 gnd.n3235 585
R1800 gnd.n3237 gnd.n3236 585
R1801 gnd.n2795 gnd.n1270 585
R1802 gnd.n4927 gnd.n1270 585
R1803 gnd.n3201 gnd.n3200 585
R1804 gnd.n3202 gnd.n3201 585
R1805 gnd.n2809 gnd.n1260 585
R1806 gnd.n4933 gnd.n1260 585
R1807 gnd.n3196 gnd.n3195 585
R1808 gnd.n3195 gnd.n3194 585
R1809 gnd.n2811 gnd.n1249 585
R1810 gnd.n4939 gnd.n1249 585
R1811 gnd.n3184 gnd.n3183 585
R1812 gnd.n3185 gnd.n3184 585
R1813 gnd.n2815 gnd.n1238 585
R1814 gnd.n4945 gnd.n1238 585
R1815 gnd.n3179 gnd.n3178 585
R1816 gnd.n3178 gnd.n3177 585
R1817 gnd.n2817 gnd.n1228 585
R1818 gnd.n4951 gnd.n1228 585
R1819 gnd.n3168 gnd.n3167 585
R1820 gnd.n3169 gnd.n3168 585
R1821 gnd.n2823 gnd.n1218 585
R1822 gnd.n4957 gnd.n1218 585
R1823 gnd.n3163 gnd.n3162 585
R1824 gnd.n3162 gnd.n3161 585
R1825 gnd.n2825 gnd.n1208 585
R1826 gnd.n4963 gnd.n1208 585
R1827 gnd.n3152 gnd.n3151 585
R1828 gnd.n3153 gnd.n3152 585
R1829 gnd.n2829 gnd.n1197 585
R1830 gnd.n4969 gnd.n1197 585
R1831 gnd.n3147 gnd.n3146 585
R1832 gnd.n3146 gnd.n3145 585
R1833 gnd.n2831 gnd.n1190 585
R1834 gnd.n4976 gnd.n1190 585
R1835 gnd.n3135 gnd.n3134 585
R1836 gnd.n3136 gnd.n3135 585
R1837 gnd.n2838 gnd.n1180 585
R1838 gnd.n4982 gnd.n1180 585
R1839 gnd.n3129 gnd.n3128 585
R1840 gnd.n3128 gnd.n3127 585
R1841 gnd.n2840 gnd.n1171 585
R1842 gnd.n4988 gnd.n1171 585
R1843 gnd.n3118 gnd.n3117 585
R1844 gnd.n3119 gnd.n3118 585
R1845 gnd.n2844 gnd.n1160 585
R1846 gnd.n4994 gnd.n1160 585
R1847 gnd.n3113 gnd.n3112 585
R1848 gnd.n3112 gnd.n3111 585
R1849 gnd.n2846 gnd.n1150 585
R1850 gnd.n5000 gnd.n1150 585
R1851 gnd.n3102 gnd.n3101 585
R1852 gnd.n3103 gnd.n3102 585
R1853 gnd.n2944 gnd.n1140 585
R1854 gnd.n5006 gnd.n1140 585
R1855 gnd.n3097 gnd.n3096 585
R1856 gnd.n3096 gnd.n3095 585
R1857 gnd.n2946 gnd.n1129 585
R1858 gnd.n5012 gnd.n1129 585
R1859 gnd.n3086 gnd.n3085 585
R1860 gnd.n3087 gnd.n3086 585
R1861 gnd.n2950 gnd.n1118 585
R1862 gnd.n5018 gnd.n1118 585
R1863 gnd.n3081 gnd.n3080 585
R1864 gnd.n3080 gnd.n3079 585
R1865 gnd.n3058 gnd.n1107 585
R1866 gnd.n5024 gnd.n1107 585
R1867 gnd.n3057 gnd.n3056 585
R1868 gnd.n3056 gnd.n1105 585
R1869 gnd.n2952 gnd.n1097 585
R1870 gnd.n5030 gnd.n1097 585
R1871 gnd.n3052 gnd.n3051 585
R1872 gnd.n3051 gnd.n1088 585
R1873 gnd.n3050 gnd.n1087 585
R1874 gnd.n5036 gnd.n1087 585
R1875 gnd.n3049 gnd.n3048 585
R1876 gnd.n3048 gnd.n1077 585
R1877 gnd.n2954 gnd.n1076 585
R1878 gnd.n5042 gnd.n1076 585
R1879 gnd.n3044 gnd.n3043 585
R1880 gnd.n3043 gnd.n1065 585
R1881 gnd.n3042 gnd.n1064 585
R1882 gnd.n5048 gnd.n1064 585
R1883 gnd.n3041 gnd.n3040 585
R1884 gnd.n3040 gnd.n1063 585
R1885 gnd.n3039 gnd.n2956 585
R1886 gnd.n3039 gnd.n3038 585
R1887 gnd.n2983 gnd.n2958 585
R1888 gnd.n2958 gnd.n1009 585
R1889 gnd.n7644 gnd.n107 585
R1890 gnd.n7740 gnd.n107 585
R1891 gnd.n7645 gnd.n7575 585
R1892 gnd.n7575 gnd.n104 585
R1893 gnd.n7646 gnd.n187 585
R1894 gnd.n7660 gnd.n187 585
R1895 gnd.n198 gnd.n196 585
R1896 gnd.n196 gnd.n186 585
R1897 gnd.n7651 gnd.n7650 585
R1898 gnd.n7652 gnd.n7651 585
R1899 gnd.n197 gnd.n195 585
R1900 gnd.n195 gnd.n193 585
R1901 gnd.n7571 gnd.n7570 585
R1902 gnd.n7570 gnd.n7569 585
R1903 gnd.n201 gnd.n200 585
R1904 gnd.n211 gnd.n201 585
R1905 gnd.n7560 gnd.n7559 585
R1906 gnd.n7561 gnd.n7560 585
R1907 gnd.n213 gnd.n212 585
R1908 gnd.n212 gnd.n208 585
R1909 gnd.n7555 gnd.n7554 585
R1910 gnd.n7554 gnd.n7553 585
R1911 gnd.n216 gnd.n215 585
R1912 gnd.n218 gnd.n216 585
R1913 gnd.n7544 gnd.n7543 585
R1914 gnd.n7545 gnd.n7544 585
R1915 gnd.n228 gnd.n227 585
R1916 gnd.n7447 gnd.n227 585
R1917 gnd.n7539 gnd.n7538 585
R1918 gnd.n7538 gnd.n7537 585
R1919 gnd.n231 gnd.n230 585
R1920 gnd.n7454 gnd.n231 585
R1921 gnd.n7528 gnd.n7527 585
R1922 gnd.n7529 gnd.n7528 585
R1923 gnd.n243 gnd.n242 585
R1924 gnd.n7414 gnd.n242 585
R1925 gnd.n7523 gnd.n7522 585
R1926 gnd.n7522 gnd.n7521 585
R1927 gnd.n246 gnd.n245 585
R1928 gnd.n7410 gnd.n246 585
R1929 gnd.n7512 gnd.n7511 585
R1930 gnd.n7513 gnd.n7512 585
R1931 gnd.n259 gnd.n258 585
R1932 gnd.n7403 gnd.n258 585
R1933 gnd.n7507 gnd.n7506 585
R1934 gnd.n7506 gnd.n7505 585
R1935 gnd.n262 gnd.n261 585
R1936 gnd.n7471 gnd.n262 585
R1937 gnd.n7484 gnd.n7483 585
R1938 gnd.n7483 gnd.n7482 585
R1939 gnd.n7485 gnd.n293 585
R1940 gnd.n7477 gnd.n293 585
R1941 gnd.n4644 gnd.n290 585
R1942 gnd.n4645 gnd.n4644 585
R1943 gnd.n7490 gnd.n289 585
R1944 gnd.n4657 gnd.n289 585
R1945 gnd.n7491 gnd.n288 585
R1946 gnd.n4661 gnd.n288 585
R1947 gnd.n7492 gnd.n287 585
R1948 gnd.n1541 gnd.n287 585
R1949 gnd.n284 gnd.n282 585
R1950 gnd.n4634 gnd.n282 585
R1951 gnd.n7497 gnd.n7496 585
R1952 gnd.n7498 gnd.n7497 585
R1953 gnd.n283 gnd.n281 585
R1954 gnd.n4622 gnd.n281 585
R1955 gnd.n4686 gnd.n4685 585
R1956 gnd.n4685 gnd.n4684 585
R1957 gnd.n4689 gnd.n1517 585
R1958 gnd.n1528 gnd.n1517 585
R1959 gnd.n4690 gnd.n1516 585
R1960 gnd.n4676 gnd.n1516 585
R1961 gnd.n4691 gnd.n1515 585
R1962 gnd.n4609 gnd.n1515 585
R1963 gnd.n1571 gnd.n1513 585
R1964 gnd.n1572 gnd.n1571 585
R1965 gnd.n4695 gnd.n1512 585
R1966 gnd.n4596 gnd.n1512 585
R1967 gnd.n4696 gnd.n1511 585
R1968 gnd.n1581 gnd.n1511 585
R1969 gnd.n4697 gnd.n1510 585
R1970 gnd.n4586 gnd.n1510 585
R1971 gnd.n4566 gnd.n1508 585
R1972 gnd.n4567 gnd.n4566 585
R1973 gnd.n4701 gnd.n1507 585
R1974 gnd.n1589 gnd.n1507 585
R1975 gnd.n4702 gnd.n1506 585
R1976 gnd.n4557 gnd.n1506 585
R1977 gnd.n4703 gnd.n1505 585
R1978 gnd.n1608 gnd.n1505 585
R1979 gnd.n4546 gnd.n1503 585
R1980 gnd.n4547 gnd.n4546 585
R1981 gnd.n4707 gnd.n1502 585
R1982 gnd.n4534 gnd.n1502 585
R1983 gnd.n4708 gnd.n1501 585
R1984 gnd.n1616 gnd.n1501 585
R1985 gnd.n4709 gnd.n1500 585
R1986 gnd.n4525 gnd.n1500 585
R1987 gnd.n1497 gnd.n1495 585
R1988 gnd.n1635 gnd.n1495 585
R1989 gnd.n4714 gnd.n4713 585
R1990 gnd.n4715 gnd.n4714 585
R1991 gnd.n1496 gnd.n1494 585
R1992 gnd.n4484 gnd.n1494 585
R1993 gnd.n1689 gnd.n1481 585
R1994 gnd.n4721 gnd.n1481 585
R1995 gnd.n1690 gnd.n1688 585
R1996 gnd.n1688 gnd.n1477 585
R1997 gnd.n1687 gnd.n1684 585
R1998 gnd.n1683 gnd.n1682 585
R1999 gnd.n1705 gnd.n1704 585
R2000 gnd.n1707 gnd.n1681 585
R2001 gnd.n1710 gnd.n1709 585
R2002 gnd.n1674 gnd.n1673 585
R2003 gnd.n1724 gnd.n1723 585
R2004 gnd.n1726 gnd.n1672 585
R2005 gnd.n1729 gnd.n1728 585
R2006 gnd.n1665 gnd.n1664 585
R2007 gnd.n1743 gnd.n1742 585
R2008 gnd.n1745 gnd.n1663 585
R2009 gnd.n1748 gnd.n1747 585
R2010 gnd.n1656 gnd.n1655 585
R2011 gnd.n1762 gnd.n1761 585
R2012 gnd.n1764 gnd.n1654 585
R2013 gnd.n1767 gnd.n1766 585
R2014 gnd.n1647 gnd.n1644 585
R2015 gnd.n4475 gnd.n4474 585
R2016 gnd.n4475 gnd.n1468 585
R2017 gnd.n7615 gnd.n103 585
R2018 gnd.n7616 gnd.n7613 585
R2019 gnd.n7617 gnd.n7609 585
R2020 gnd.n7607 gnd.n7605 585
R2021 gnd.n7621 gnd.n7604 585
R2022 gnd.n7622 gnd.n7602 585
R2023 gnd.n7623 gnd.n7601 585
R2024 gnd.n7599 gnd.n7597 585
R2025 gnd.n7627 gnd.n7596 585
R2026 gnd.n7628 gnd.n7594 585
R2027 gnd.n7629 gnd.n7593 585
R2028 gnd.n7591 gnd.n7589 585
R2029 gnd.n7633 gnd.n7588 585
R2030 gnd.n7634 gnd.n7586 585
R2031 gnd.n7635 gnd.n7585 585
R2032 gnd.n7583 gnd.n7581 585
R2033 gnd.n7639 gnd.n7580 585
R2034 gnd.n7640 gnd.n7578 585
R2035 gnd.n7641 gnd.n7577 585
R2036 gnd.n7577 gnd.n117 585
R2037 gnd.n7742 gnd.n7741 585
R2038 gnd.n7741 gnd.n7740 585
R2039 gnd.n7743 gnd.n101 585
R2040 gnd.n104 gnd.n101 585
R2041 gnd.n7744 gnd.n100 585
R2042 gnd.n7660 gnd.n100 585
R2043 gnd.n185 gnd.n98 585
R2044 gnd.n186 gnd.n185 585
R2045 gnd.n7748 gnd.n97 585
R2046 gnd.n7652 gnd.n97 585
R2047 gnd.n7749 gnd.n96 585
R2048 gnd.n193 gnd.n96 585
R2049 gnd.n7750 gnd.n95 585
R2050 gnd.n7569 gnd.n95 585
R2051 gnd.n210 gnd.n93 585
R2052 gnd.n211 gnd.n210 585
R2053 gnd.n7754 gnd.n92 585
R2054 gnd.n7561 gnd.n92 585
R2055 gnd.n7755 gnd.n91 585
R2056 gnd.n208 gnd.n91 585
R2057 gnd.n7756 gnd.n90 585
R2058 gnd.n7553 gnd.n90 585
R2059 gnd.n217 gnd.n88 585
R2060 gnd.n218 gnd.n217 585
R2061 gnd.n7760 gnd.n87 585
R2062 gnd.n7545 gnd.n87 585
R2063 gnd.n7761 gnd.n86 585
R2064 gnd.n7447 gnd.n86 585
R2065 gnd.n7762 gnd.n85 585
R2066 gnd.n7537 gnd.n85 585
R2067 gnd.n7453 gnd.n83 585
R2068 gnd.n7454 gnd.n7453 585
R2069 gnd.n7766 gnd.n82 585
R2070 gnd.n7529 gnd.n82 585
R2071 gnd.n7767 gnd.n81 585
R2072 gnd.n7414 gnd.n81 585
R2073 gnd.n7768 gnd.n80 585
R2074 gnd.n7521 gnd.n80 585
R2075 gnd.n7409 gnd.n78 585
R2076 gnd.n7410 gnd.n7409 585
R2077 gnd.n7772 gnd.n77 585
R2078 gnd.n7513 gnd.n77 585
R2079 gnd.n7773 gnd.n76 585
R2080 gnd.n7403 gnd.n76 585
R2081 gnd.n7774 gnd.n75 585
R2082 gnd.n7505 gnd.n75 585
R2083 gnd.n305 gnd.n73 585
R2084 gnd.n7471 gnd.n305 585
R2085 gnd.n7778 gnd.n72 585
R2086 gnd.n7482 gnd.n72 585
R2087 gnd.n7779 gnd.n71 585
R2088 gnd.n7477 gnd.n71 585
R2089 gnd.n7780 gnd.n70 585
R2090 gnd.n4645 gnd.n70 585
R2091 gnd.n4643 gnd.n69 585
R2092 gnd.n4657 gnd.n4643 585
R2093 gnd.n4627 gnd.n1543 585
R2094 gnd.n4661 gnd.n1543 585
R2095 gnd.n1553 gnd.n1551 585
R2096 gnd.n1551 gnd.n1541 585
R2097 gnd.n4632 gnd.n4631 585
R2098 gnd.n4634 gnd.n4632 585
R2099 gnd.n1552 gnd.n279 585
R2100 gnd.n7498 gnd.n279 585
R2101 gnd.n4624 gnd.n4623 585
R2102 gnd.n4623 gnd.n4622 585
R2103 gnd.n1555 gnd.n1519 585
R2104 gnd.n4684 gnd.n1519 585
R2105 gnd.n4602 gnd.n4601 585
R2106 gnd.n4601 gnd.n1528 585
R2107 gnd.n1564 gnd.n1527 585
R2108 gnd.n4676 gnd.n1527 585
R2109 gnd.n4607 gnd.n4606 585
R2110 gnd.n4609 gnd.n4607 585
R2111 gnd.n1563 gnd.n1562 585
R2112 gnd.n1572 gnd.n1562 585
R2113 gnd.n4598 gnd.n4597 585
R2114 gnd.n4597 gnd.n4596 585
R2115 gnd.n1567 gnd.n1566 585
R2116 gnd.n1581 gnd.n1567 585
R2117 gnd.n1593 gnd.n1580 585
R2118 gnd.n4586 gnd.n1580 585
R2119 gnd.n4565 gnd.n4564 585
R2120 gnd.n4567 gnd.n4565 585
R2121 gnd.n1592 gnd.n1591 585
R2122 gnd.n1591 gnd.n1589 585
R2123 gnd.n4559 gnd.n4558 585
R2124 gnd.n4558 gnd.n4557 585
R2125 gnd.n1596 gnd.n1595 585
R2126 gnd.n1608 gnd.n1596 585
R2127 gnd.n1620 gnd.n1607 585
R2128 gnd.n4547 gnd.n1607 585
R2129 gnd.n4533 gnd.n4532 585
R2130 gnd.n4534 gnd.n4533 585
R2131 gnd.n1619 gnd.n1618 585
R2132 gnd.n1618 gnd.n1616 585
R2133 gnd.n4527 gnd.n4526 585
R2134 gnd.n4526 gnd.n4525 585
R2135 gnd.n1623 gnd.n1622 585
R2136 gnd.n1635 gnd.n1623 585
R2137 gnd.n1642 gnd.n1492 585
R2138 gnd.n4715 gnd.n1492 585
R2139 gnd.n4483 gnd.n4482 585
R2140 gnd.n4484 gnd.n4483 585
R2141 gnd.n1641 gnd.n1479 585
R2142 gnd.n4721 gnd.n1479 585
R2143 gnd.n4477 gnd.n4476 585
R2144 gnd.n4476 gnd.n1477 585
R2145 gnd.n953 gnd.n952 585
R2146 gnd.n956 gnd.n953 585
R2147 gnd.n6498 gnd.n6497 585
R2148 gnd.n6497 gnd.n6496 585
R2149 gnd.n6499 gnd.n947 585
R2150 gnd.n6395 gnd.n947 585
R2151 gnd.n6501 gnd.n6500 585
R2152 gnd.n6502 gnd.n6501 585
R2153 gnd.n948 gnd.n946 585
R2154 gnd.n946 gnd.n942 585
R2155 gnd.n928 gnd.n927 585
R2156 gnd.n931 gnd.n928 585
R2157 gnd.n6512 gnd.n6511 585
R2158 gnd.n6511 gnd.n6510 585
R2159 gnd.n6513 gnd.n922 585
R2160 gnd.n6116 gnd.n922 585
R2161 gnd.n6515 gnd.n6514 585
R2162 gnd.n6516 gnd.n6515 585
R2163 gnd.n923 gnd.n921 585
R2164 gnd.n6100 gnd.n921 585
R2165 gnd.n6091 gnd.n6090 585
R2166 gnd.n6090 gnd.n909 585
R2167 gnd.n6089 gnd.n5208 585
R2168 gnd.n6089 gnd.n907 585
R2169 gnd.n6088 gnd.n5210 585
R2170 gnd.n6088 gnd.n6087 585
R2171 gnd.n6078 gnd.n5209 585
R2172 gnd.n5221 gnd.n5209 585
R2173 gnd.n6077 gnd.n6076 585
R2174 gnd.n6076 gnd.n6075 585
R2175 gnd.n5218 gnd.n5216 585
R2176 gnd.n6062 gnd.n5218 585
R2177 gnd.n6053 gnd.n6052 585
R2178 gnd.n6052 gnd.n6051 585
R2179 gnd.n5233 gnd.n5232 585
R2180 gnd.n5241 gnd.n5233 585
R2181 gnd.n6030 gnd.n6029 585
R2182 gnd.n6031 gnd.n6030 585
R2183 gnd.n5244 gnd.n5243 585
R2184 gnd.n5252 gnd.n5243 585
R2185 gnd.n6004 gnd.n5264 585
R2186 gnd.n5264 gnd.n5251 585
R2187 gnd.n6006 gnd.n6005 585
R2188 gnd.n6007 gnd.n6006 585
R2189 gnd.n5265 gnd.n5263 585
R2190 gnd.n5263 gnd.n5259 585
R2191 gnd.n5993 gnd.n5992 585
R2192 gnd.n5992 gnd.n5991 585
R2193 gnd.n5270 gnd.n5269 585
R2194 gnd.n5280 gnd.n5270 585
R2195 gnd.n5982 gnd.n5981 585
R2196 gnd.n5981 gnd.n5980 585
R2197 gnd.n5277 gnd.n5276 585
R2198 gnd.n5968 gnd.n5277 585
R2199 gnd.n5942 gnd.n5346 585
R2200 gnd.n5346 gnd.n5287 585
R2201 gnd.n5944 gnd.n5943 585
R2202 gnd.n5945 gnd.n5944 585
R2203 gnd.n5347 gnd.n5345 585
R2204 gnd.n5355 gnd.n5345 585
R2205 gnd.n5920 gnd.n5367 585
R2206 gnd.n5367 gnd.n5354 585
R2207 gnd.n5922 gnd.n5921 585
R2208 gnd.n5923 gnd.n5922 585
R2209 gnd.n5368 gnd.n5366 585
R2210 gnd.n5366 gnd.n5362 585
R2211 gnd.n5908 gnd.n5907 585
R2212 gnd.n5907 gnd.n5906 585
R2213 gnd.n5373 gnd.n5372 585
R2214 gnd.n5382 gnd.n5373 585
R2215 gnd.n5897 gnd.n5896 585
R2216 gnd.n5896 gnd.n5895 585
R2217 gnd.n5380 gnd.n5379 585
R2218 gnd.n5883 gnd.n5380 585
R2219 gnd.n5855 gnd.n5854 585
R2220 gnd.n5854 gnd.n5389 585
R2221 gnd.n5856 gnd.n5400 585
R2222 gnd.n5847 gnd.n5400 585
R2223 gnd.n5858 gnd.n5857 585
R2224 gnd.n5859 gnd.n5858 585
R2225 gnd.n5401 gnd.n5399 585
R2226 gnd.n5415 gnd.n5399 585
R2227 gnd.n5839 gnd.n5838 585
R2228 gnd.n5838 gnd.n5837 585
R2229 gnd.n5412 gnd.n5411 585
R2230 gnd.n5822 gnd.n5412 585
R2231 gnd.n5809 gnd.n5432 585
R2232 gnd.n5432 gnd.n5422 585
R2233 gnd.n5811 gnd.n5810 585
R2234 gnd.n5812 gnd.n5811 585
R2235 gnd.n5433 gnd.n5431 585
R2236 gnd.n5441 gnd.n5431 585
R2237 gnd.n5785 gnd.n5453 585
R2238 gnd.n5453 gnd.n5440 585
R2239 gnd.n5787 gnd.n5786 585
R2240 gnd.n5788 gnd.n5787 585
R2241 gnd.n5454 gnd.n5452 585
R2242 gnd.n5452 gnd.n5448 585
R2243 gnd.n5773 gnd.n5772 585
R2244 gnd.n5772 gnd.n5771 585
R2245 gnd.n5459 gnd.n5458 585
R2246 gnd.n5463 gnd.n5459 585
R2247 gnd.n5757 gnd.n5756 585
R2248 gnd.n5758 gnd.n5757 585
R2249 gnd.n5474 gnd.n5473 585
R2250 gnd.n5473 gnd.n5469 585
R2251 gnd.n5747 gnd.n5746 585
R2252 gnd.n5748 gnd.n5747 585
R2253 gnd.n5483 gnd.n5482 585
R2254 gnd.n5482 gnd.n5480 585
R2255 gnd.n5741 gnd.n5740 585
R2256 gnd.n5740 gnd.n5739 585
R2257 gnd.n5487 gnd.n5486 585
R2258 gnd.n5495 gnd.n5487 585
R2259 gnd.n5648 gnd.n5647 585
R2260 gnd.n5649 gnd.n5648 585
R2261 gnd.n5497 gnd.n5496 585
R2262 gnd.n5496 gnd.n5494 585
R2263 gnd.n5643 gnd.n5642 585
R2264 gnd.n5642 gnd.n5641 585
R2265 gnd.n5500 gnd.n5499 585
R2266 gnd.n5501 gnd.n5500 585
R2267 gnd.n5632 gnd.n5631 585
R2268 gnd.n5633 gnd.n5632 585
R2269 gnd.n5509 gnd.n5508 585
R2270 gnd.n5508 gnd.n5507 585
R2271 gnd.n5627 gnd.n5626 585
R2272 gnd.n5626 gnd.n5625 585
R2273 gnd.n5512 gnd.n5511 585
R2274 gnd.n5513 gnd.n5512 585
R2275 gnd.n5616 gnd.n5615 585
R2276 gnd.n5617 gnd.n5616 585
R2277 gnd.n5612 gnd.n5519 585
R2278 gnd.n5611 gnd.n5610 585
R2279 gnd.n5608 gnd.n5521 585
R2280 gnd.n5608 gnd.n5518 585
R2281 gnd.n5607 gnd.n5606 585
R2282 gnd.n5605 gnd.n5604 585
R2283 gnd.n5603 gnd.n5526 585
R2284 gnd.n5601 gnd.n5600 585
R2285 gnd.n5599 gnd.n5527 585
R2286 gnd.n5598 gnd.n5597 585
R2287 gnd.n5595 gnd.n5532 585
R2288 gnd.n5593 gnd.n5592 585
R2289 gnd.n5591 gnd.n5533 585
R2290 gnd.n5590 gnd.n5589 585
R2291 gnd.n5587 gnd.n5538 585
R2292 gnd.n5585 gnd.n5584 585
R2293 gnd.n5583 gnd.n5539 585
R2294 gnd.n5582 gnd.n5581 585
R2295 gnd.n5579 gnd.n5544 585
R2296 gnd.n5577 gnd.n5576 585
R2297 gnd.n5575 gnd.n5545 585
R2298 gnd.n5574 gnd.n5573 585
R2299 gnd.n5571 gnd.n5550 585
R2300 gnd.n5569 gnd.n5568 585
R2301 gnd.n5566 gnd.n5551 585
R2302 gnd.n5565 gnd.n5564 585
R2303 gnd.n5562 gnd.n5560 585
R2304 gnd.n5558 gnd.n5517 585
R2305 gnd.n6404 gnd.n6403 585
R2306 gnd.n6406 gnd.n6405 585
R2307 gnd.n6408 gnd.n6407 585
R2308 gnd.n6410 gnd.n6409 585
R2309 gnd.n6412 gnd.n6411 585
R2310 gnd.n6414 gnd.n6413 585
R2311 gnd.n6416 gnd.n6415 585
R2312 gnd.n6418 gnd.n6417 585
R2313 gnd.n6420 gnd.n6419 585
R2314 gnd.n6422 gnd.n6421 585
R2315 gnd.n6424 gnd.n6423 585
R2316 gnd.n6426 gnd.n6425 585
R2317 gnd.n6428 gnd.n6427 585
R2318 gnd.n6430 gnd.n6429 585
R2319 gnd.n6432 gnd.n6431 585
R2320 gnd.n6434 gnd.n6433 585
R2321 gnd.n6436 gnd.n6435 585
R2322 gnd.n6438 gnd.n6437 585
R2323 gnd.n6440 gnd.n6439 585
R2324 gnd.n6442 gnd.n6441 585
R2325 gnd.n6444 gnd.n6443 585
R2326 gnd.n6446 gnd.n6445 585
R2327 gnd.n6448 gnd.n6447 585
R2328 gnd.n6450 gnd.n6449 585
R2329 gnd.n6452 gnd.n6451 585
R2330 gnd.n6453 gnd.n5162 585
R2331 gnd.n6454 gnd.n967 585
R2332 gnd.n6487 gnd.n967 585
R2333 gnd.n6402 gnd.n6401 585
R2334 gnd.n6402 gnd.n956 585
R2335 gnd.n5191 gnd.n954 585
R2336 gnd.n6496 gnd.n954 585
R2337 gnd.n6397 gnd.n6396 585
R2338 gnd.n6396 gnd.n6395 585
R2339 gnd.n5193 gnd.n944 585
R2340 gnd.n6502 gnd.n944 585
R2341 gnd.n6110 gnd.n6109 585
R2342 gnd.n6110 gnd.n942 585
R2343 gnd.n6112 gnd.n6111 585
R2344 gnd.n6111 gnd.n931 585
R2345 gnd.n6113 gnd.n929 585
R2346 gnd.n6510 gnd.n929 585
R2347 gnd.n6115 gnd.n6114 585
R2348 gnd.n6116 gnd.n6115 585
R2349 gnd.n5202 gnd.n919 585
R2350 gnd.n6516 gnd.n919 585
R2351 gnd.n6102 gnd.n6101 585
R2352 gnd.n6101 gnd.n6100 585
R2353 gnd.n5205 gnd.n5204 585
R2354 gnd.n5205 gnd.n909 585
R2355 gnd.n6043 gnd.n6042 585
R2356 gnd.n6042 gnd.n907 585
R2357 gnd.n6044 gnd.n5212 585
R2358 gnd.n6087 gnd.n5212 585
R2359 gnd.n6046 gnd.n6045 585
R2360 gnd.n6045 gnd.n5221 585
R2361 gnd.n6047 gnd.n5219 585
R2362 gnd.n6075 gnd.n5219 585
R2363 gnd.n6048 gnd.n5229 585
R2364 gnd.n6062 gnd.n5229 585
R2365 gnd.n6050 gnd.n6049 585
R2366 gnd.n6051 gnd.n6050 585
R2367 gnd.n5236 gnd.n5235 585
R2368 gnd.n5241 gnd.n5235 585
R2369 gnd.n6033 gnd.n6032 585
R2370 gnd.n6032 gnd.n6031 585
R2371 gnd.n5239 gnd.n5238 585
R2372 gnd.n5252 gnd.n5239 585
R2373 gnd.n5958 gnd.n5957 585
R2374 gnd.n5957 gnd.n5251 585
R2375 gnd.n5959 gnd.n5261 585
R2376 gnd.n6007 gnd.n5261 585
R2377 gnd.n5961 gnd.n5960 585
R2378 gnd.n5960 gnd.n5259 585
R2379 gnd.n5962 gnd.n5272 585
R2380 gnd.n5991 gnd.n5272 585
R2381 gnd.n5964 gnd.n5963 585
R2382 gnd.n5963 gnd.n5280 585
R2383 gnd.n5965 gnd.n5279 585
R2384 gnd.n5980 gnd.n5279 585
R2385 gnd.n5967 gnd.n5966 585
R2386 gnd.n5968 gnd.n5967 585
R2387 gnd.n5291 gnd.n5290 585
R2388 gnd.n5290 gnd.n5287 585
R2389 gnd.n5947 gnd.n5946 585
R2390 gnd.n5946 gnd.n5945 585
R2391 gnd.n5342 gnd.n5341 585
R2392 gnd.n5355 gnd.n5342 585
R2393 gnd.n5868 gnd.n5867 585
R2394 gnd.n5867 gnd.n5354 585
R2395 gnd.n5869 gnd.n5364 585
R2396 gnd.n5923 gnd.n5364 585
R2397 gnd.n5872 gnd.n5871 585
R2398 gnd.n5871 gnd.n5362 585
R2399 gnd.n5873 gnd.n5375 585
R2400 gnd.n5906 gnd.n5375 585
R2401 gnd.n5876 gnd.n5875 585
R2402 gnd.n5875 gnd.n5382 585
R2403 gnd.n5877 gnd.n5381 585
R2404 gnd.n5895 gnd.n5381 585
R2405 gnd.n5880 gnd.n5879 585
R2406 gnd.n5883 gnd.n5880 585
R2407 gnd.n5865 gnd.n5391 585
R2408 gnd.n5391 gnd.n5389 585
R2409 gnd.n5396 gnd.n5392 585
R2410 gnd.n5847 gnd.n5396 585
R2411 gnd.n5861 gnd.n5860 585
R2412 gnd.n5860 gnd.n5859 585
R2413 gnd.n5395 gnd.n5394 585
R2414 gnd.n5415 gnd.n5395 585
R2415 gnd.n5819 gnd.n5414 585
R2416 gnd.n5837 gnd.n5414 585
R2417 gnd.n5821 gnd.n5820 585
R2418 gnd.n5822 gnd.n5821 585
R2419 gnd.n5425 gnd.n5424 585
R2420 gnd.n5424 gnd.n5422 585
R2421 gnd.n5814 gnd.n5813 585
R2422 gnd.n5813 gnd.n5812 585
R2423 gnd.n5428 gnd.n5427 585
R2424 gnd.n5441 gnd.n5428 585
R2425 gnd.n5665 gnd.n5664 585
R2426 gnd.n5664 gnd.n5440 585
R2427 gnd.n5666 gnd.n5450 585
R2428 gnd.n5788 gnd.n5450 585
R2429 gnd.n5668 gnd.n5667 585
R2430 gnd.n5667 gnd.n5448 585
R2431 gnd.n5669 gnd.n5460 585
R2432 gnd.n5771 gnd.n5460 585
R2433 gnd.n5671 gnd.n5670 585
R2434 gnd.n5670 gnd.n5463 585
R2435 gnd.n5672 gnd.n5471 585
R2436 gnd.n5758 gnd.n5471 585
R2437 gnd.n5674 gnd.n5673 585
R2438 gnd.n5673 gnd.n5469 585
R2439 gnd.n5675 gnd.n5481 585
R2440 gnd.n5748 gnd.n5481 585
R2441 gnd.n5676 gnd.n5489 585
R2442 gnd.n5489 gnd.n5480 585
R2443 gnd.n5678 gnd.n5677 585
R2444 gnd.n5739 gnd.n5678 585
R2445 gnd.n5490 gnd.n5488 585
R2446 gnd.n5495 gnd.n5488 585
R2447 gnd.n5651 gnd.n5650 585
R2448 gnd.n5650 gnd.n5649 585
R2449 gnd.n5493 gnd.n5492 585
R2450 gnd.n5494 gnd.n5493 585
R2451 gnd.n5640 gnd.n5639 585
R2452 gnd.n5641 gnd.n5640 585
R2453 gnd.n5503 gnd.n5502 585
R2454 gnd.n5502 gnd.n5501 585
R2455 gnd.n5635 gnd.n5634 585
R2456 gnd.n5634 gnd.n5633 585
R2457 gnd.n5506 gnd.n5505 585
R2458 gnd.n5507 gnd.n5506 585
R2459 gnd.n5624 gnd.n5623 585
R2460 gnd.n5625 gnd.n5624 585
R2461 gnd.n5515 gnd.n5514 585
R2462 gnd.n5514 gnd.n5513 585
R2463 gnd.n5619 gnd.n5618 585
R2464 gnd.n5618 gnd.n5617 585
R2465 gnd.n6492 gnd.n958 585
R2466 gnd.n966 gnd.n958 585
R2467 gnd.n6494 gnd.n6493 585
R2468 gnd.n6495 gnd.n6494 585
R2469 gnd.n959 gnd.n957 585
R2470 gnd.n6394 gnd.n957 585
R2471 gnd.n941 gnd.n940 585
R2472 gnd.n945 gnd.n941 585
R2473 gnd.n6505 gnd.n6504 585
R2474 gnd.n6504 gnd.n6503 585
R2475 gnd.n6506 gnd.n933 585
R2476 gnd.n5195 gnd.n933 585
R2477 gnd.n6508 gnd.n6507 585
R2478 gnd.n6509 gnd.n6508 585
R2479 gnd.n934 gnd.n932 585
R2480 gnd.n6117 gnd.n932 585
R2481 gnd.n917 gnd.n916 585
R2482 gnd.n920 gnd.n917 585
R2483 gnd.n6519 gnd.n6518 585
R2484 gnd.n6518 gnd.n6517 585
R2485 gnd.n6520 gnd.n911 585
R2486 gnd.n6099 gnd.n911 585
R2487 gnd.n6522 gnd.n6521 585
R2488 gnd.n6523 gnd.n6522 585
R2489 gnd.n912 gnd.n910 585
R2490 gnd.n6086 gnd.n910 585
R2491 gnd.n6071 gnd.n5223 585
R2492 gnd.n5223 gnd.n5211 585
R2493 gnd.n6073 gnd.n6072 585
R2494 gnd.n6074 gnd.n6073 585
R2495 gnd.n5224 gnd.n5222 585
R2496 gnd.n6061 gnd.n5222 585
R2497 gnd.n6065 gnd.n6064 585
R2498 gnd.n6064 gnd.n6063 585
R2499 gnd.n5227 gnd.n5226 585
R2500 gnd.n5234 gnd.n5227 585
R2501 gnd.n6017 gnd.n6016 585
R2502 gnd.n6016 gnd.n5242 585
R2503 gnd.n6018 gnd.n5254 585
R2504 gnd.n5254 gnd.n5240 585
R2505 gnd.n6020 gnd.n6019 585
R2506 gnd.n6021 gnd.n6020 585
R2507 gnd.n5255 gnd.n5253 585
R2508 gnd.n5262 gnd.n5253 585
R2509 gnd.n6010 gnd.n6009 585
R2510 gnd.n6009 gnd.n6008 585
R2511 gnd.n5258 gnd.n5257 585
R2512 gnd.n5990 gnd.n5258 585
R2513 gnd.n5976 gnd.n5282 585
R2514 gnd.n5282 gnd.n5271 585
R2515 gnd.n5978 gnd.n5977 585
R2516 gnd.n5979 gnd.n5978 585
R2517 gnd.n5283 gnd.n5281 585
R2518 gnd.n5281 gnd.n5278 585
R2519 gnd.n5971 gnd.n5970 585
R2520 gnd.n5970 gnd.n5969 585
R2521 gnd.n5286 gnd.n5285 585
R2522 gnd.n5344 gnd.n5286 585
R2523 gnd.n5931 gnd.n5357 585
R2524 gnd.n5357 gnd.n5343 585
R2525 gnd.n5933 gnd.n5932 585
R2526 gnd.n5934 gnd.n5933 585
R2527 gnd.n5358 gnd.n5356 585
R2528 gnd.n5365 gnd.n5356 585
R2529 gnd.n5926 gnd.n5925 585
R2530 gnd.n5925 gnd.n5924 585
R2531 gnd.n5361 gnd.n5360 585
R2532 gnd.n5905 gnd.n5361 585
R2533 gnd.n5891 gnd.n5384 585
R2534 gnd.n5384 gnd.n5374 585
R2535 gnd.n5893 gnd.n5892 585
R2536 gnd.n5894 gnd.n5893 585
R2537 gnd.n5385 gnd.n5383 585
R2538 gnd.n5882 gnd.n5383 585
R2539 gnd.n5886 gnd.n5885 585
R2540 gnd.n5885 gnd.n5884 585
R2541 gnd.n5388 gnd.n5387 585
R2542 gnd.n5848 gnd.n5388 585
R2543 gnd.n5832 gnd.n5831 585
R2544 gnd.n5831 gnd.n5398 585
R2545 gnd.n5833 gnd.n5417 585
R2546 gnd.n5417 gnd.n5397 585
R2547 gnd.n5835 gnd.n5834 585
R2548 gnd.n5836 gnd.n5835 585
R2549 gnd.n5418 gnd.n5416 585
R2550 gnd.n5416 gnd.n5413 585
R2551 gnd.n5825 gnd.n5824 585
R2552 gnd.n5824 gnd.n5823 585
R2553 gnd.n5421 gnd.n5420 585
R2554 gnd.n5430 gnd.n5421 585
R2555 gnd.n5796 gnd.n5443 585
R2556 gnd.n5443 gnd.n5429 585
R2557 gnd.n5798 gnd.n5797 585
R2558 gnd.n5799 gnd.n5798 585
R2559 gnd.n5444 gnd.n5442 585
R2560 gnd.n5451 gnd.n5442 585
R2561 gnd.n5791 gnd.n5790 585
R2562 gnd.n5790 gnd.n5789 585
R2563 gnd.n5447 gnd.n5446 585
R2564 gnd.n5770 gnd.n5447 585
R2565 gnd.n5766 gnd.n5765 585
R2566 gnd.n5767 gnd.n5766 585
R2567 gnd.n5465 gnd.n5464 585
R2568 gnd.n5472 gnd.n5464 585
R2569 gnd.n5761 gnd.n5760 585
R2570 gnd.n5760 gnd.n5759 585
R2571 gnd.n5468 gnd.n5467 585
R2572 gnd.n5749 gnd.n5468 585
R2573 gnd.n5736 gnd.n5735 585
R2574 gnd.n5734 gnd.n5687 585
R2575 gnd.n5733 gnd.n5686 585
R2576 gnd.n5738 gnd.n5686 585
R2577 gnd.n5732 gnd.n5731 585
R2578 gnd.n5730 gnd.n5729 585
R2579 gnd.n5728 gnd.n5727 585
R2580 gnd.n5726 gnd.n5725 585
R2581 gnd.n5724 gnd.n5723 585
R2582 gnd.n5722 gnd.n5721 585
R2583 gnd.n5720 gnd.n5719 585
R2584 gnd.n5718 gnd.n5717 585
R2585 gnd.n5716 gnd.n5715 585
R2586 gnd.n5714 gnd.n5713 585
R2587 gnd.n5712 gnd.n5711 585
R2588 gnd.n5710 gnd.n5709 585
R2589 gnd.n5708 gnd.n5707 585
R2590 gnd.n5703 gnd.n5479 585
R2591 gnd.n6388 gnd.n5157 585
R2592 gnd.n6460 gnd.n6459 585
R2593 gnd.n6462 gnd.n6461 585
R2594 gnd.n6464 gnd.n6463 585
R2595 gnd.n6466 gnd.n6465 585
R2596 gnd.n6468 gnd.n6467 585
R2597 gnd.n6470 gnd.n6469 585
R2598 gnd.n6472 gnd.n6471 585
R2599 gnd.n6474 gnd.n6473 585
R2600 gnd.n6476 gnd.n6475 585
R2601 gnd.n6478 gnd.n6477 585
R2602 gnd.n6480 gnd.n6479 585
R2603 gnd.n6482 gnd.n6481 585
R2604 gnd.n6483 gnd.n5143 585
R2605 gnd.n6485 gnd.n6484 585
R2606 gnd.n965 gnd.n964 585
R2607 gnd.n6489 gnd.n6488 585
R2608 gnd.n6488 gnd.n6487 585
R2609 gnd.n6390 gnd.n6389 585
R2610 gnd.n6389 gnd.n966 585
R2611 gnd.n6391 gnd.n955 585
R2612 gnd.n6495 gnd.n955 585
R2613 gnd.n6393 gnd.n6392 585
R2614 gnd.n6394 gnd.n6393 585
R2615 gnd.n6384 gnd.n5194 585
R2616 gnd.n5194 gnd.n945 585
R2617 gnd.n6382 gnd.n943 585
R2618 gnd.n6503 gnd.n943 585
R2619 gnd.n5197 gnd.n5196 585
R2620 gnd.n5196 gnd.n5195 585
R2621 gnd.n6120 gnd.n930 585
R2622 gnd.n6509 gnd.n930 585
R2623 gnd.n6119 gnd.n6118 585
R2624 gnd.n6118 gnd.n6117 585
R2625 gnd.n5201 gnd.n5199 585
R2626 gnd.n5201 gnd.n920 585
R2627 gnd.n6096 gnd.n918 585
R2628 gnd.n6517 gnd.n918 585
R2629 gnd.n6098 gnd.n6097 585
R2630 gnd.n6099 gnd.n6098 585
R2631 gnd.n5206 gnd.n908 585
R2632 gnd.n6523 gnd.n908 585
R2633 gnd.n6085 gnd.n6084 585
R2634 gnd.n6086 gnd.n6085 585
R2635 gnd.n5214 gnd.n5213 585
R2636 gnd.n5213 gnd.n5211 585
R2637 gnd.n6058 gnd.n5220 585
R2638 gnd.n6074 gnd.n5220 585
R2639 gnd.n6060 gnd.n6059 585
R2640 gnd.n6061 gnd.n6060 585
R2641 gnd.n5230 gnd.n5228 585
R2642 gnd.n6063 gnd.n5228 585
R2643 gnd.n6024 gnd.n5248 585
R2644 gnd.n6024 gnd.n5234 585
R2645 gnd.n6026 gnd.n6025 585
R2646 gnd.n6025 gnd.n5242 585
R2647 gnd.n6023 gnd.n5247 585
R2648 gnd.n6023 gnd.n5240 585
R2649 gnd.n6022 gnd.n5250 585
R2650 gnd.n6022 gnd.n6021 585
R2651 gnd.n5999 gnd.n5249 585
R2652 gnd.n5262 gnd.n5249 585
R2653 gnd.n5998 gnd.n5260 585
R2654 gnd.n6008 gnd.n5260 585
R2655 gnd.n5989 gnd.n5267 585
R2656 gnd.n5990 gnd.n5989 585
R2657 gnd.n5988 gnd.n5987 585
R2658 gnd.n5988 gnd.n5271 585
R2659 gnd.n5986 gnd.n5273 585
R2660 gnd.n5979 gnd.n5273 585
R2661 gnd.n5288 gnd.n5274 585
R2662 gnd.n5288 gnd.n5278 585
R2663 gnd.n5939 gnd.n5289 585
R2664 gnd.n5969 gnd.n5289 585
R2665 gnd.n5938 gnd.n5937 585
R2666 gnd.n5937 gnd.n5344 585
R2667 gnd.n5936 gnd.n5351 585
R2668 gnd.n5936 gnd.n5343 585
R2669 gnd.n5935 gnd.n5353 585
R2670 gnd.n5935 gnd.n5934 585
R2671 gnd.n5914 gnd.n5352 585
R2672 gnd.n5365 gnd.n5352 585
R2673 gnd.n5913 gnd.n5363 585
R2674 gnd.n5924 gnd.n5363 585
R2675 gnd.n5904 gnd.n5370 585
R2676 gnd.n5905 gnd.n5904 585
R2677 gnd.n5903 gnd.n5902 585
R2678 gnd.n5903 gnd.n5374 585
R2679 gnd.n5901 gnd.n5376 585
R2680 gnd.n5894 gnd.n5376 585
R2681 gnd.n5881 gnd.n5377 585
R2682 gnd.n5882 gnd.n5881 585
R2683 gnd.n5851 gnd.n5390 585
R2684 gnd.n5884 gnd.n5390 585
R2685 gnd.n5850 gnd.n5849 585
R2686 gnd.n5849 gnd.n5848 585
R2687 gnd.n5846 gnd.n5407 585
R2688 gnd.n5846 gnd.n5398 585
R2689 gnd.n5845 gnd.n5844 585
R2690 gnd.n5845 gnd.n5397 585
R2691 gnd.n5409 gnd.n5408 585
R2692 gnd.n5836 gnd.n5408 585
R2693 gnd.n5805 gnd.n5804 585
R2694 gnd.n5804 gnd.n5413 585
R2695 gnd.n5806 gnd.n5423 585
R2696 gnd.n5823 gnd.n5423 585
R2697 gnd.n5803 gnd.n5802 585
R2698 gnd.n5802 gnd.n5430 585
R2699 gnd.n5801 gnd.n5437 585
R2700 gnd.n5801 gnd.n5429 585
R2701 gnd.n5800 gnd.n5439 585
R2702 gnd.n5800 gnd.n5799 585
R2703 gnd.n5779 gnd.n5438 585
R2704 gnd.n5451 gnd.n5438 585
R2705 gnd.n5778 gnd.n5449 585
R2706 gnd.n5789 gnd.n5449 585
R2707 gnd.n5769 gnd.n5456 585
R2708 gnd.n5770 gnd.n5769 585
R2709 gnd.n5768 gnd.n5462 585
R2710 gnd.n5768 gnd.n5767 585
R2711 gnd.n5753 gnd.n5461 585
R2712 gnd.n5472 gnd.n5461 585
R2713 gnd.n5752 gnd.n5470 585
R2714 gnd.n5759 gnd.n5470 585
R2715 gnd.n5751 gnd.n5750 585
R2716 gnd.n5750 gnd.n5749 585
R2717 gnd.n4899 gnd.n4898 585
R2718 gnd.n4898 gnd.n4897 585
R2719 gnd.n4900 gnd.n1314 585
R2720 gnd.n3528 gnd.n1314 585
R2721 gnd.n4902 gnd.n4901 585
R2722 gnd.n4903 gnd.n4902 585
R2723 gnd.n1299 gnd.n1298 585
R2724 gnd.n3223 gnd.n1299 585
R2725 gnd.n4911 gnd.n4910 585
R2726 gnd.n4910 gnd.n4909 585
R2727 gnd.n4912 gnd.n1293 585
R2728 gnd.n3214 gnd.n1293 585
R2729 gnd.n4914 gnd.n4913 585
R2730 gnd.n4915 gnd.n4914 585
R2731 gnd.n1277 gnd.n1276 585
R2732 gnd.n3210 gnd.n1277 585
R2733 gnd.n4923 gnd.n4922 585
R2734 gnd.n4922 gnd.n4921 585
R2735 gnd.n4924 gnd.n1271 585
R2736 gnd.n3237 gnd.n1271 585
R2737 gnd.n4926 gnd.n4925 585
R2738 gnd.n4927 gnd.n4926 585
R2739 gnd.n1257 gnd.n1256 585
R2740 gnd.n3202 gnd.n1257 585
R2741 gnd.n4935 gnd.n4934 585
R2742 gnd.n4934 gnd.n4933 585
R2743 gnd.n4936 gnd.n1251 585
R2744 gnd.n3194 gnd.n1251 585
R2745 gnd.n4938 gnd.n4937 585
R2746 gnd.n4939 gnd.n4938 585
R2747 gnd.n1235 gnd.n1234 585
R2748 gnd.n3185 gnd.n1235 585
R2749 gnd.n4947 gnd.n4946 585
R2750 gnd.n4946 gnd.n4945 585
R2751 gnd.n4948 gnd.n1229 585
R2752 gnd.n3177 gnd.n1229 585
R2753 gnd.n4950 gnd.n4949 585
R2754 gnd.n4951 gnd.n4950 585
R2755 gnd.n1215 gnd.n1214 585
R2756 gnd.n3169 gnd.n1215 585
R2757 gnd.n4959 gnd.n4958 585
R2758 gnd.n4958 gnd.n4957 585
R2759 gnd.n4960 gnd.n1210 585
R2760 gnd.n3161 gnd.n1210 585
R2761 gnd.n4962 gnd.n4961 585
R2762 gnd.n4963 gnd.n4962 585
R2763 gnd.n1211 gnd.n1194 585
R2764 gnd.n3153 gnd.n1194 585
R2765 gnd.n4971 gnd.n4970 585
R2766 gnd.n4970 gnd.n4969 585
R2767 gnd.n4972 gnd.n1191 585
R2768 gnd.n3145 gnd.n1191 585
R2769 gnd.n4975 gnd.n4974 585
R2770 gnd.n4976 gnd.n4975 585
R2771 gnd.n1192 gnd.n1177 585
R2772 gnd.n3136 gnd.n1177 585
R2773 gnd.n4984 gnd.n4983 585
R2774 gnd.n4983 gnd.n4982 585
R2775 gnd.n4985 gnd.n1173 585
R2776 gnd.n3127 gnd.n1173 585
R2777 gnd.n4987 gnd.n4986 585
R2778 gnd.n4988 gnd.n4987 585
R2779 gnd.n1157 gnd.n1156 585
R2780 gnd.n3119 gnd.n1157 585
R2781 gnd.n4996 gnd.n4995 585
R2782 gnd.n4995 gnd.n4994 585
R2783 gnd.n4997 gnd.n1151 585
R2784 gnd.n3111 gnd.n1151 585
R2785 gnd.n4999 gnd.n4998 585
R2786 gnd.n5000 gnd.n4999 585
R2787 gnd.n1137 gnd.n1136 585
R2788 gnd.n3103 gnd.n1137 585
R2789 gnd.n5008 gnd.n5007 585
R2790 gnd.n5007 gnd.n5006 585
R2791 gnd.n5009 gnd.n1131 585
R2792 gnd.n3095 gnd.n1131 585
R2793 gnd.n5011 gnd.n5010 585
R2794 gnd.n5012 gnd.n5011 585
R2795 gnd.n1115 gnd.n1114 585
R2796 gnd.n3087 gnd.n1115 585
R2797 gnd.n5020 gnd.n5019 585
R2798 gnd.n5019 gnd.n5018 585
R2799 gnd.n5021 gnd.n1109 585
R2800 gnd.n3079 gnd.n1109 585
R2801 gnd.n5023 gnd.n5022 585
R2802 gnd.n5024 gnd.n5023 585
R2803 gnd.n1095 gnd.n1094 585
R2804 gnd.n1105 gnd.n1095 585
R2805 gnd.n5032 gnd.n5031 585
R2806 gnd.n5031 gnd.n5030 585
R2807 gnd.n5033 gnd.n1089 585
R2808 gnd.n1089 gnd.n1088 585
R2809 gnd.n5035 gnd.n5034 585
R2810 gnd.n5036 gnd.n5035 585
R2811 gnd.n1074 gnd.n1073 585
R2812 gnd.n1077 gnd.n1074 585
R2813 gnd.n5044 gnd.n5043 585
R2814 gnd.n5043 gnd.n5042 585
R2815 gnd.n5045 gnd.n1068 585
R2816 gnd.n1068 gnd.n1065 585
R2817 gnd.n5047 gnd.n5046 585
R2818 gnd.n5048 gnd.n5047 585
R2819 gnd.n1069 gnd.n1067 585
R2820 gnd.n1067 gnd.n1063 585
R2821 gnd.n3037 gnd.n3036 585
R2822 gnd.n3038 gnd.n3037 585
R2823 gnd.n3032 gnd.n1012 585
R2824 gnd.n1012 gnd.n1009 585
R2825 gnd.n5133 gnd.n5132 585
R2826 gnd.n5131 gnd.n1011 585
R2827 gnd.n5130 gnd.n1010 585
R2828 gnd.n5135 gnd.n1010 585
R2829 gnd.n5129 gnd.n5128 585
R2830 gnd.n5127 gnd.n5126 585
R2831 gnd.n5125 gnd.n5124 585
R2832 gnd.n5123 gnd.n5122 585
R2833 gnd.n5121 gnd.n5120 585
R2834 gnd.n5119 gnd.n5118 585
R2835 gnd.n5117 gnd.n5116 585
R2836 gnd.n5115 gnd.n5114 585
R2837 gnd.n5113 gnd.n5112 585
R2838 gnd.n5111 gnd.n5110 585
R2839 gnd.n5109 gnd.n5108 585
R2840 gnd.n5107 gnd.n5106 585
R2841 gnd.n5105 gnd.n5104 585
R2842 gnd.n5103 gnd.n5102 585
R2843 gnd.n5101 gnd.n5100 585
R2844 gnd.n5098 gnd.n5097 585
R2845 gnd.n5096 gnd.n5095 585
R2846 gnd.n5094 gnd.n5093 585
R2847 gnd.n5092 gnd.n5091 585
R2848 gnd.n5090 gnd.n5089 585
R2849 gnd.n5088 gnd.n5087 585
R2850 gnd.n5086 gnd.n5085 585
R2851 gnd.n5084 gnd.n5083 585
R2852 gnd.n5082 gnd.n5081 585
R2853 gnd.n5080 gnd.n5079 585
R2854 gnd.n5078 gnd.n5077 585
R2855 gnd.n5076 gnd.n5075 585
R2856 gnd.n5074 gnd.n5073 585
R2857 gnd.n5072 gnd.n5071 585
R2858 gnd.n5070 gnd.n5069 585
R2859 gnd.n5068 gnd.n5067 585
R2860 gnd.n5066 gnd.n5065 585
R2861 gnd.n5064 gnd.n5063 585
R2862 gnd.n5062 gnd.n1051 585
R2863 gnd.n1055 gnd.n1052 585
R2864 gnd.n5058 gnd.n5057 585
R2865 gnd.n3535 gnd.n3534 585
R2866 gnd.n3537 gnd.n2696 585
R2867 gnd.n3539 gnd.n3538 585
R2868 gnd.n3540 gnd.n2689 585
R2869 gnd.n3542 gnd.n3541 585
R2870 gnd.n3544 gnd.n2687 585
R2871 gnd.n3546 gnd.n3545 585
R2872 gnd.n3547 gnd.n2682 585
R2873 gnd.n3549 gnd.n3548 585
R2874 gnd.n3551 gnd.n2680 585
R2875 gnd.n3553 gnd.n3552 585
R2876 gnd.n3554 gnd.n2675 585
R2877 gnd.n3556 gnd.n3555 585
R2878 gnd.n3558 gnd.n2673 585
R2879 gnd.n3560 gnd.n3559 585
R2880 gnd.n3561 gnd.n2668 585
R2881 gnd.n3563 gnd.n3562 585
R2882 gnd.n3565 gnd.n2667 585
R2883 gnd.n3566 gnd.n2610 585
R2884 gnd.n3569 gnd.n3568 585
R2885 gnd.n2611 gnd.n2603 585
R2886 gnd.n2639 gnd.n2604 585
R2887 gnd.n2641 gnd.n2640 585
R2888 gnd.n2643 gnd.n2642 585
R2889 gnd.n2645 gnd.n2644 585
R2890 gnd.n2647 gnd.n2646 585
R2891 gnd.n2649 gnd.n2648 585
R2892 gnd.n2651 gnd.n2650 585
R2893 gnd.n2653 gnd.n2652 585
R2894 gnd.n2655 gnd.n2654 585
R2895 gnd.n2657 gnd.n2656 585
R2896 gnd.n2659 gnd.n2658 585
R2897 gnd.n2661 gnd.n2660 585
R2898 gnd.n2662 gnd.n2621 585
R2899 gnd.n2664 gnd.n2663 585
R2900 gnd.n2622 gnd.n2620 585
R2901 gnd.n2623 gnd.n1319 585
R2902 gnd.n2666 gnd.n1319 585
R2903 gnd.n3531 gnd.n1321 585
R2904 gnd.n4897 gnd.n1321 585
R2905 gnd.n3530 gnd.n3529 585
R2906 gnd.n3529 gnd.n3528 585
R2907 gnd.n2700 gnd.n1312 585
R2908 gnd.n4903 gnd.n1312 585
R2909 gnd.n3222 gnd.n3221 585
R2910 gnd.n3223 gnd.n3222 585
R2911 gnd.n2802 gnd.n1301 585
R2912 gnd.n4909 gnd.n1301 585
R2913 gnd.n3216 gnd.n3215 585
R2914 gnd.n3215 gnd.n3214 585
R2915 gnd.n3213 gnd.n1290 585
R2916 gnd.n4915 gnd.n1290 585
R2917 gnd.n3212 gnd.n3211 585
R2918 gnd.n3211 gnd.n3210 585
R2919 gnd.n2804 gnd.n1279 585
R2920 gnd.n4921 gnd.n1279 585
R2921 gnd.n3206 gnd.n2794 585
R2922 gnd.n3237 gnd.n2794 585
R2923 gnd.n3205 gnd.n1269 585
R2924 gnd.n4927 gnd.n1269 585
R2925 gnd.n3204 gnd.n3203 585
R2926 gnd.n3203 gnd.n3202 585
R2927 gnd.n2806 gnd.n1259 585
R2928 gnd.n4933 gnd.n1259 585
R2929 gnd.n3193 gnd.n3192 585
R2930 gnd.n3194 gnd.n3193 585
R2931 gnd.n2812 gnd.n1248 585
R2932 gnd.n4939 gnd.n1248 585
R2933 gnd.n3187 gnd.n3186 585
R2934 gnd.n3186 gnd.n3185 585
R2935 gnd.n2814 gnd.n1237 585
R2936 gnd.n4945 gnd.n1237 585
R2937 gnd.n3176 gnd.n3175 585
R2938 gnd.n3177 gnd.n3176 585
R2939 gnd.n2819 gnd.n1227 585
R2940 gnd.n4951 gnd.n1227 585
R2941 gnd.n3171 gnd.n3170 585
R2942 gnd.n3170 gnd.n3169 585
R2943 gnd.n2821 gnd.n1217 585
R2944 gnd.n4957 gnd.n1217 585
R2945 gnd.n3160 gnd.n3159 585
R2946 gnd.n3161 gnd.n3160 585
R2947 gnd.n2826 gnd.n1207 585
R2948 gnd.n4963 gnd.n1207 585
R2949 gnd.n3155 gnd.n3154 585
R2950 gnd.n3154 gnd.n3153 585
R2951 gnd.n2828 gnd.n1196 585
R2952 gnd.n4969 gnd.n1196 585
R2953 gnd.n3144 gnd.n3143 585
R2954 gnd.n3145 gnd.n3144 585
R2955 gnd.n2833 gnd.n1189 585
R2956 gnd.n4976 gnd.n1189 585
R2957 gnd.n3138 gnd.n3137 585
R2958 gnd.n3137 gnd.n3136 585
R2959 gnd.n2836 gnd.n1179 585
R2960 gnd.n4982 gnd.n1179 585
R2961 gnd.n3126 gnd.n3125 585
R2962 gnd.n3127 gnd.n3126 585
R2963 gnd.n2841 gnd.n1170 585
R2964 gnd.n4988 gnd.n1170 585
R2965 gnd.n3121 gnd.n3120 585
R2966 gnd.n3120 gnd.n3119 585
R2967 gnd.n2843 gnd.n1159 585
R2968 gnd.n4994 gnd.n1159 585
R2969 gnd.n3110 gnd.n3109 585
R2970 gnd.n3111 gnd.n3110 585
R2971 gnd.n2848 gnd.n1149 585
R2972 gnd.n5000 gnd.n1149 585
R2973 gnd.n3105 gnd.n3104 585
R2974 gnd.n3104 gnd.n3103 585
R2975 gnd.n2850 gnd.n1139 585
R2976 gnd.n5006 gnd.n1139 585
R2977 gnd.n3094 gnd.n3093 585
R2978 gnd.n3095 gnd.n3094 585
R2979 gnd.n2947 gnd.n1128 585
R2980 gnd.n5012 gnd.n1128 585
R2981 gnd.n3089 gnd.n3088 585
R2982 gnd.n3088 gnd.n3087 585
R2983 gnd.n2949 gnd.n1117 585
R2984 gnd.n5018 gnd.n1117 585
R2985 gnd.n3078 gnd.n3077 585
R2986 gnd.n3079 gnd.n3078 585
R2987 gnd.n3059 gnd.n1106 585
R2988 gnd.n5024 gnd.n1106 585
R2989 gnd.n3073 gnd.n3072 585
R2990 gnd.n3072 gnd.n1105 585
R2991 gnd.n3071 gnd.n1096 585
R2992 gnd.n5030 gnd.n1096 585
R2993 gnd.n3070 gnd.n3069 585
R2994 gnd.n3069 gnd.n1088 585
R2995 gnd.n3061 gnd.n1086 585
R2996 gnd.n5036 gnd.n1086 585
R2997 gnd.n3065 gnd.n3064 585
R2998 gnd.n3064 gnd.n1077 585
R2999 gnd.n3063 gnd.n1075 585
R3000 gnd.n5042 gnd.n1075 585
R3001 gnd.n1062 gnd.n1060 585
R3002 gnd.n1065 gnd.n1062 585
R3003 gnd.n5050 gnd.n5049 585
R3004 gnd.n5049 gnd.n5048 585
R3005 gnd.n1061 gnd.n1058 585
R3006 gnd.n1063 gnd.n1061 585
R3007 gnd.n5054 gnd.n1057 585
R3008 gnd.n3038 gnd.n1057 585
R3009 gnd.n5056 gnd.n5055 585
R3010 gnd.n5056 gnd.n1009 585
R3011 gnd.n7739 gnd.n7738 585
R3012 gnd.n7740 gnd.n7739 585
R3013 gnd.n110 gnd.n108 585
R3014 gnd.n108 gnd.n104 585
R3015 gnd.n7659 gnd.n7658 585
R3016 gnd.n7660 gnd.n7659 585
R3017 gnd.n189 gnd.n188 585
R3018 gnd.n188 gnd.n186 585
R3019 gnd.n7654 gnd.n7653 585
R3020 gnd.n7653 gnd.n7652 585
R3021 gnd.n192 gnd.n191 585
R3022 gnd.n193 gnd.n192 585
R3023 gnd.n7568 gnd.n7567 585
R3024 gnd.n7569 gnd.n7568 585
R3025 gnd.n204 gnd.n203 585
R3026 gnd.n211 gnd.n203 585
R3027 gnd.n7563 gnd.n7562 585
R3028 gnd.n7562 gnd.n7561 585
R3029 gnd.n207 gnd.n206 585
R3030 gnd.n208 gnd.n207 585
R3031 gnd.n7552 gnd.n7551 585
R3032 gnd.n7553 gnd.n7552 585
R3033 gnd.n221 gnd.n220 585
R3034 gnd.n220 gnd.n218 585
R3035 gnd.n7547 gnd.n7546 585
R3036 gnd.n7546 gnd.n7545 585
R3037 gnd.n224 gnd.n223 585
R3038 gnd.n7447 gnd.n224 585
R3039 gnd.n7536 gnd.n7535 585
R3040 gnd.n7537 gnd.n7536 585
R3041 gnd.n235 gnd.n234 585
R3042 gnd.n7454 gnd.n234 585
R3043 gnd.n7531 gnd.n7530 585
R3044 gnd.n7530 gnd.n7529 585
R3045 gnd.n238 gnd.n237 585
R3046 gnd.n7414 gnd.n238 585
R3047 gnd.n7520 gnd.n7519 585
R3048 gnd.n7521 gnd.n7520 585
R3049 gnd.n251 gnd.n250 585
R3050 gnd.n7410 gnd.n250 585
R3051 gnd.n7515 gnd.n7514 585
R3052 gnd.n7514 gnd.n7513 585
R3053 gnd.n254 gnd.n253 585
R3054 gnd.n7403 gnd.n254 585
R3055 gnd.n7504 gnd.n7503 585
R3056 gnd.n7505 gnd.n7504 585
R3057 gnd.n266 gnd.n265 585
R3058 gnd.n7471 gnd.n265 585
R3059 gnd.n7481 gnd.n7480 585
R3060 gnd.n7482 gnd.n7481 585
R3061 gnd.n7479 gnd.n7478 585
R3062 gnd.n7478 gnd.n7477 585
R3063 gnd.n1546 gnd.n297 585
R3064 gnd.n4645 gnd.n297 585
R3065 gnd.n4658 gnd.n1547 585
R3066 gnd.n4658 gnd.n4657 585
R3067 gnd.n4660 gnd.n4659 585
R3068 gnd.n4661 gnd.n4660 585
R3069 gnd.n1545 gnd.n272 585
R3070 gnd.n1545 gnd.n1541 585
R3071 gnd.n276 gnd.n273 585
R3072 gnd.n4634 gnd.n276 585
R3073 gnd.n7500 gnd.n7499 585
R3074 gnd.n7499 gnd.n7498 585
R3075 gnd.n275 gnd.n274 585
R3076 gnd.n4622 gnd.n275 585
R3077 gnd.n4683 gnd.n4682 585
R3078 gnd.n4684 gnd.n4683 585
R3079 gnd.n1522 gnd.n1521 585
R3080 gnd.n1528 gnd.n1521 585
R3081 gnd.n4678 gnd.n4677 585
R3082 gnd.n4677 gnd.n4676 585
R3083 gnd.n1525 gnd.n1524 585
R3084 gnd.n4609 gnd.n1525 585
R3085 gnd.n4593 gnd.n1573 585
R3086 gnd.n1573 gnd.n1572 585
R3087 gnd.n4595 gnd.n4594 585
R3088 gnd.n4596 gnd.n4595 585
R3089 gnd.n1574 gnd.n1570 585
R3090 gnd.n1581 gnd.n1570 585
R3091 gnd.n4588 gnd.n4587 585
R3092 gnd.n4587 gnd.n4586 585
R3093 gnd.n1577 gnd.n1576 585
R3094 gnd.n4567 gnd.n1577 585
R3095 gnd.n4554 gnd.n1600 585
R3096 gnd.n1600 gnd.n1589 585
R3097 gnd.n4556 gnd.n4555 585
R3098 gnd.n4557 gnd.n4556 585
R3099 gnd.n1601 gnd.n1599 585
R3100 gnd.n1608 gnd.n1599 585
R3101 gnd.n4549 gnd.n4548 585
R3102 gnd.n4548 gnd.n4547 585
R3103 gnd.n1604 gnd.n1603 585
R3104 gnd.n4534 gnd.n1604 585
R3105 gnd.n4522 gnd.n4518 585
R3106 gnd.n4518 gnd.n1616 585
R3107 gnd.n4524 gnd.n4523 585
R3108 gnd.n4525 gnd.n4524 585
R3109 gnd.n1489 gnd.n1488 585
R3110 gnd.n1635 gnd.n1489 585
R3111 gnd.n4717 gnd.n4716 585
R3112 gnd.n4716 gnd.n4715 585
R3113 gnd.n4718 gnd.n1483 585
R3114 gnd.n4484 gnd.n1483 585
R3115 gnd.n4720 gnd.n4719 585
R3116 gnd.n4721 gnd.n4720 585
R3117 gnd.n1484 gnd.n1482 585
R3118 gnd.n1482 gnd.n1477 585
R3119 gnd.n1909 gnd.n1908 585
R3120 gnd.n1912 gnd.n1911 585
R3121 gnd.n1905 gnd.n1904 585
R3122 gnd.n1904 gnd.n1468 585
R3123 gnd.n1917 gnd.n1916 585
R3124 gnd.n1919 gnd.n1903 585
R3125 gnd.n1922 gnd.n1921 585
R3126 gnd.n1901 gnd.n1900 585
R3127 gnd.n1927 gnd.n1926 585
R3128 gnd.n1929 gnd.n1899 585
R3129 gnd.n1932 gnd.n1931 585
R3130 gnd.n1897 gnd.n1896 585
R3131 gnd.n1938 gnd.n1937 585
R3132 gnd.n1940 gnd.n1895 585
R3133 gnd.n1941 gnd.n1892 585
R3134 gnd.n1944 gnd.n1943 585
R3135 gnd.n1894 gnd.n1889 585
R3136 gnd.n2029 gnd.n2028 585
R3137 gnd.n2026 gnd.n1951 585
R3138 gnd.n2024 gnd.n2023 585
R3139 gnd.n2022 gnd.n1952 585
R3140 gnd.n2021 gnd.n2020 585
R3141 gnd.n2018 gnd.n1957 585
R3142 gnd.n2016 gnd.n2015 585
R3143 gnd.n2014 gnd.n1958 585
R3144 gnd.n2013 gnd.n2012 585
R3145 gnd.n2010 gnd.n1963 585
R3146 gnd.n2008 gnd.n2007 585
R3147 gnd.n2006 gnd.n1964 585
R3148 gnd.n2005 gnd.n2004 585
R3149 gnd.n2002 gnd.n1969 585
R3150 gnd.n2000 gnd.n1999 585
R3151 gnd.n1998 gnd.n1970 585
R3152 gnd.n1997 gnd.n1996 585
R3153 gnd.n1994 gnd.n1975 585
R3154 gnd.n1992 gnd.n1991 585
R3155 gnd.n1979 gnd.n1976 585
R3156 gnd.n1987 gnd.n1986 585
R3157 gnd.n179 gnd.n178 585
R3158 gnd.n7668 gnd.n174 585
R3159 gnd.n7670 gnd.n7669 585
R3160 gnd.n7672 gnd.n172 585
R3161 gnd.n7674 gnd.n7673 585
R3162 gnd.n7675 gnd.n167 585
R3163 gnd.n7677 gnd.n7676 585
R3164 gnd.n7679 gnd.n165 585
R3165 gnd.n7681 gnd.n7680 585
R3166 gnd.n7682 gnd.n160 585
R3167 gnd.n7684 gnd.n7683 585
R3168 gnd.n7686 gnd.n158 585
R3169 gnd.n7688 gnd.n7687 585
R3170 gnd.n7689 gnd.n153 585
R3171 gnd.n7691 gnd.n7690 585
R3172 gnd.n7693 gnd.n151 585
R3173 gnd.n7695 gnd.n7694 585
R3174 gnd.n7696 gnd.n146 585
R3175 gnd.n7698 gnd.n7697 585
R3176 gnd.n7700 gnd.n144 585
R3177 gnd.n7702 gnd.n7701 585
R3178 gnd.n7706 gnd.n139 585
R3179 gnd.n7708 gnd.n7707 585
R3180 gnd.n7710 gnd.n137 585
R3181 gnd.n7712 gnd.n7711 585
R3182 gnd.n7713 gnd.n132 585
R3183 gnd.n7715 gnd.n7714 585
R3184 gnd.n7717 gnd.n130 585
R3185 gnd.n7719 gnd.n7718 585
R3186 gnd.n7720 gnd.n125 585
R3187 gnd.n7722 gnd.n7721 585
R3188 gnd.n7724 gnd.n123 585
R3189 gnd.n7726 gnd.n7725 585
R3190 gnd.n7727 gnd.n118 585
R3191 gnd.n7729 gnd.n7728 585
R3192 gnd.n7731 gnd.n115 585
R3193 gnd.n7733 gnd.n7732 585
R3194 gnd.n7734 gnd.n113 585
R3195 gnd.n7735 gnd.n109 585
R3196 gnd.n117 gnd.n109 585
R3197 gnd.n7664 gnd.n105 585
R3198 gnd.n7740 gnd.n105 585
R3199 gnd.n7663 gnd.n7662 585
R3200 gnd.n7662 gnd.n104 585
R3201 gnd.n7661 gnd.n183 585
R3202 gnd.n7661 gnd.n7660 585
R3203 gnd.n7433 gnd.n184 585
R3204 gnd.n186 gnd.n184 585
R3205 gnd.n7434 gnd.n194 585
R3206 gnd.n7652 gnd.n194 585
R3207 gnd.n7436 gnd.n7435 585
R3208 gnd.n7435 gnd.n193 585
R3209 gnd.n7437 gnd.n202 585
R3210 gnd.n7569 gnd.n202 585
R3211 gnd.n7439 gnd.n7438 585
R3212 gnd.n7438 gnd.n211 585
R3213 gnd.n7440 gnd.n209 585
R3214 gnd.n7561 gnd.n209 585
R3215 gnd.n7442 gnd.n7441 585
R3216 gnd.n7441 gnd.n208 585
R3217 gnd.n7443 gnd.n219 585
R3218 gnd.n7553 gnd.n219 585
R3219 gnd.n7445 gnd.n7444 585
R3220 gnd.n7444 gnd.n218 585
R3221 gnd.n7446 gnd.n226 585
R3222 gnd.n7545 gnd.n226 585
R3223 gnd.n7449 gnd.n7448 585
R3224 gnd.n7448 gnd.n7447 585
R3225 gnd.n7450 gnd.n232 585
R3226 gnd.n7537 gnd.n232 585
R3227 gnd.n7452 gnd.n7451 585
R3228 gnd.n7454 gnd.n7452 585
R3229 gnd.n7399 gnd.n240 585
R3230 gnd.n7529 gnd.n240 585
R3231 gnd.n7416 gnd.n7415 585
R3232 gnd.n7415 gnd.n7414 585
R3233 gnd.n7413 gnd.n248 585
R3234 gnd.n7521 gnd.n248 585
R3235 gnd.n7412 gnd.n7411 585
R3236 gnd.n7411 gnd.n7410 585
R3237 gnd.n7401 gnd.n256 585
R3238 gnd.n7513 gnd.n256 585
R3239 gnd.n7405 gnd.n7404 585
R3240 gnd.n7404 gnd.n7403 585
R3241 gnd.n304 gnd.n263 585
R3242 gnd.n7505 gnd.n263 585
R3243 gnd.n7473 gnd.n7472 585
R3244 gnd.n7472 gnd.n7471 585
R3245 gnd.n7474 gnd.n295 585
R3246 gnd.n7482 gnd.n295 585
R3247 gnd.n7476 gnd.n7475 585
R3248 gnd.n7477 gnd.n7476 585
R3249 gnd.n299 gnd.n298 585
R3250 gnd.n4645 gnd.n298 585
R3251 gnd.n4642 gnd.n4641 585
R3252 gnd.n4657 gnd.n4642 585
R3253 gnd.n1548 gnd.n1542 585
R3254 gnd.n4661 gnd.n1542 585
R3255 gnd.n4637 gnd.n4636 585
R3256 gnd.n4636 gnd.n1541 585
R3257 gnd.n4635 gnd.n1550 585
R3258 gnd.n4635 gnd.n4634 585
R3259 gnd.n4619 gnd.n278 585
R3260 gnd.n7498 gnd.n278 585
R3261 gnd.n4621 gnd.n4620 585
R3262 gnd.n4622 gnd.n4621 585
R3263 gnd.n1556 gnd.n1518 585
R3264 gnd.n4684 gnd.n1518 585
R3265 gnd.n4614 gnd.n4613 585
R3266 gnd.n4613 gnd.n1528 585
R3267 gnd.n4612 gnd.n1526 585
R3268 gnd.n4676 gnd.n1526 585
R3269 gnd.n4611 gnd.n4610 585
R3270 gnd.n4610 gnd.n4609 585
R3271 gnd.n1560 gnd.n1558 585
R3272 gnd.n1572 gnd.n1560 585
R3273 gnd.n4502 gnd.n1568 585
R3274 gnd.n4596 gnd.n1568 585
R3275 gnd.n4504 gnd.n4503 585
R3276 gnd.n4503 gnd.n1581 585
R3277 gnd.n4505 gnd.n1579 585
R3278 gnd.n4586 gnd.n1579 585
R3279 gnd.n4506 gnd.n1590 585
R3280 gnd.n4567 gnd.n1590 585
R3281 gnd.n4508 gnd.n4507 585
R3282 gnd.n4507 gnd.n1589 585
R3283 gnd.n4509 gnd.n1597 585
R3284 gnd.n4557 gnd.n1597 585
R3285 gnd.n4511 gnd.n4510 585
R3286 gnd.n4510 gnd.n1608 585
R3287 gnd.n4512 gnd.n1606 585
R3288 gnd.n4547 gnd.n1606 585
R3289 gnd.n4513 gnd.n1617 585
R3290 gnd.n4534 gnd.n1617 585
R3291 gnd.n4514 gnd.n1637 585
R3292 gnd.n1637 gnd.n1616 585
R3293 gnd.n4516 gnd.n4515 585
R3294 gnd.n4525 gnd.n4516 585
R3295 gnd.n1638 gnd.n1636 585
R3296 gnd.n1636 gnd.n1635 585
R3297 gnd.n4487 gnd.n1491 585
R3298 gnd.n4715 gnd.n1491 585
R3299 gnd.n4486 gnd.n4485 585
R3300 gnd.n4485 gnd.n4484 585
R3301 gnd.n1640 gnd.n1478 585
R3302 gnd.n4721 gnd.n1478 585
R3303 gnd.n1984 gnd.n1983 585
R3304 gnd.n1984 gnd.n1477 585
R3305 gnd.n4297 gnd.n4296 585
R3306 gnd.n4298 gnd.n4297 585
R3307 gnd.n4208 gnd.n2038 585
R3308 gnd.n2046 gnd.n2038 585
R3309 gnd.n4207 gnd.n4206 585
R3310 gnd.n4206 gnd.n4205 585
R3311 gnd.n2041 gnd.n2040 585
R3312 gnd.n4117 gnd.n2041 585
R3313 gnd.n4188 gnd.n4187 585
R3314 gnd.n4189 gnd.n4188 585
R3315 gnd.n4186 gnd.n2057 585
R3316 gnd.n2057 gnd.n2053 585
R3317 gnd.n4185 gnd.n4184 585
R3318 gnd.n4184 gnd.n4183 585
R3319 gnd.n2059 gnd.n2058 585
R3320 gnd.n4125 gnd.n2059 585
R3321 gnd.n4164 gnd.n4163 585
R3322 gnd.n4165 gnd.n4164 585
R3323 gnd.n4162 gnd.n2071 585
R3324 gnd.n2071 gnd.n2068 585
R3325 gnd.n4161 gnd.n4160 585
R3326 gnd.n4160 gnd.n4159 585
R3327 gnd.n2073 gnd.n2072 585
R3328 gnd.n4133 gnd.n2073 585
R3329 gnd.n4146 gnd.n4145 585
R3330 gnd.n4147 gnd.n4146 585
R3331 gnd.n4144 gnd.n2085 585
R3332 gnd.n4139 gnd.n2085 585
R3333 gnd.n4143 gnd.n4142 585
R3334 gnd.n4142 gnd.n4141 585
R3335 gnd.n2087 gnd.n2086 585
R3336 gnd.n4111 gnd.n2087 585
R3337 gnd.n4093 gnd.n2102 585
R3338 gnd.n2109 gnd.n2102 585
R3339 gnd.n4095 gnd.n4094 585
R3340 gnd.n4096 gnd.n4095 585
R3341 gnd.n4092 gnd.n2101 585
R3342 gnd.n2101 gnd.n2099 585
R3343 gnd.n4091 gnd.n4090 585
R3344 gnd.n4090 gnd.n4089 585
R3345 gnd.n2104 gnd.n2103 585
R3346 gnd.n4059 gnd.n2104 585
R3347 gnd.n4072 gnd.n4071 585
R3348 gnd.n4073 gnd.n4072 585
R3349 gnd.n4070 gnd.n2119 585
R3350 gnd.n4065 gnd.n2119 585
R3351 gnd.n4069 gnd.n4068 585
R3352 gnd.n4068 gnd.n4067 585
R3353 gnd.n2121 gnd.n2120 585
R3354 gnd.n4051 gnd.n2121 585
R3355 gnd.n4037 gnd.n2137 585
R3356 gnd.n2137 gnd.n2136 585
R3357 gnd.n4039 gnd.n4038 585
R3358 gnd.n4040 gnd.n4039 585
R3359 gnd.n4036 gnd.n2135 585
R3360 gnd.n2135 gnd.n2131 585
R3361 gnd.n4035 gnd.n4034 585
R3362 gnd.n4034 gnd.n4033 585
R3363 gnd.n2139 gnd.n2138 585
R3364 gnd.n3968 gnd.n2139 585
R3365 gnd.n4007 gnd.n4006 585
R3366 gnd.n4008 gnd.n4007 585
R3367 gnd.n4005 gnd.n2151 585
R3368 gnd.n2151 gnd.n2148 585
R3369 gnd.n4004 gnd.n4003 585
R3370 gnd.n4003 gnd.n4002 585
R3371 gnd.n2153 gnd.n2152 585
R3372 gnd.n3976 gnd.n2153 585
R3373 gnd.n3989 gnd.n3988 585
R3374 gnd.n3990 gnd.n3989 585
R3375 gnd.n3987 gnd.n2166 585
R3376 gnd.n2166 gnd.n2163 585
R3377 gnd.n3986 gnd.n3985 585
R3378 gnd.n3985 gnd.n3984 585
R3379 gnd.n2168 gnd.n2167 585
R3380 gnd.n2182 gnd.n2168 585
R3381 gnd.n3957 gnd.n3956 585
R3382 gnd.n3958 gnd.n3957 585
R3383 gnd.n3955 gnd.n2175 585
R3384 gnd.n3950 gnd.n2175 585
R3385 gnd.n3954 gnd.n3953 585
R3386 gnd.n3953 gnd.n3952 585
R3387 gnd.n2177 gnd.n2176 585
R3388 gnd.n3938 gnd.n2177 585
R3389 gnd.n3910 gnd.n2201 585
R3390 gnd.n2201 gnd.n2189 585
R3391 gnd.n3912 gnd.n3911 585
R3392 gnd.n3913 gnd.n3912 585
R3393 gnd.n3909 gnd.n2200 585
R3394 gnd.n2200 gnd.n2197 585
R3395 gnd.n3908 gnd.n3907 585
R3396 gnd.n3907 gnd.n3906 585
R3397 gnd.n2203 gnd.n2202 585
R3398 gnd.n2244 gnd.n2203 585
R3399 gnd.n3895 gnd.n3894 585
R3400 gnd.n3896 gnd.n3895 585
R3401 gnd.n3893 gnd.n2215 585
R3402 gnd.n2215 gnd.n2211 585
R3403 gnd.n3892 gnd.n3891 585
R3404 gnd.n3891 gnd.n3890 585
R3405 gnd.n2217 gnd.n2216 585
R3406 gnd.n3863 gnd.n2217 585
R3407 gnd.n3877 gnd.n3876 585
R3408 gnd.n3878 gnd.n3877 585
R3409 gnd.n3875 gnd.n2229 585
R3410 gnd.n3869 gnd.n2229 585
R3411 gnd.n3874 gnd.n3873 585
R3412 gnd.n3873 gnd.n3872 585
R3413 gnd.n2231 gnd.n2230 585
R3414 gnd.n3851 gnd.n2231 585
R3415 gnd.n3842 gnd.n2264 585
R3416 gnd.n2264 gnd.n2256 585
R3417 gnd.n3844 gnd.n3843 585
R3418 gnd.n3845 gnd.n3844 585
R3419 gnd.n3841 gnd.n2263 585
R3420 gnd.n3804 gnd.n2263 585
R3421 gnd.n3840 gnd.n3839 585
R3422 gnd.n3839 gnd.n3838 585
R3423 gnd.n2266 gnd.n2265 585
R3424 gnd.n2469 gnd.n2266 585
R3425 gnd.n3825 gnd.n3824 585
R3426 gnd.n3826 gnd.n3825 585
R3427 gnd.n3823 gnd.n2278 585
R3428 gnd.n2278 gnd.n2275 585
R3429 gnd.n3822 gnd.n3821 585
R3430 gnd.n3821 gnd.n3820 585
R3431 gnd.n2280 gnd.n2279 585
R3432 gnd.n2477 gnd.n2280 585
R3433 gnd.n3794 gnd.n3793 585
R3434 gnd.n3795 gnd.n3794 585
R3435 gnd.n3792 gnd.n2291 585
R3436 gnd.n2296 gnd.n2291 585
R3437 gnd.n3791 gnd.n3790 585
R3438 gnd.n3790 gnd.n3789 585
R3439 gnd.n2293 gnd.n2292 585
R3440 gnd.n2484 gnd.n2293 585
R3441 gnd.n3775 gnd.n3774 585
R3442 gnd.n3776 gnd.n3775 585
R3443 gnd.n3773 gnd.n2305 585
R3444 gnd.n3768 gnd.n2305 585
R3445 gnd.n3772 gnd.n3771 585
R3446 gnd.n3771 gnd.n3770 585
R3447 gnd.n2307 gnd.n2306 585
R3448 gnd.n2319 gnd.n2307 585
R3449 gnd.n3744 gnd.n2329 585
R3450 gnd.n2492 gnd.n2329 585
R3451 gnd.n3746 gnd.n3745 585
R3452 gnd.n3747 gnd.n3746 585
R3453 gnd.n3743 gnd.n2328 585
R3454 gnd.n2328 gnd.n2325 585
R3455 gnd.n3742 gnd.n3741 585
R3456 gnd.n3741 gnd.n3740 585
R3457 gnd.n2331 gnd.n2330 585
R3458 gnd.n2501 gnd.n2331 585
R3459 gnd.n3729 gnd.n3728 585
R3460 gnd.n3730 gnd.n3729 585
R3461 gnd.n3727 gnd.n2341 585
R3462 gnd.n2505 gnd.n2341 585
R3463 gnd.n3726 gnd.n3725 585
R3464 gnd.n3725 gnd.n3724 585
R3465 gnd.n2343 gnd.n2342 585
R3466 gnd.n2511 gnd.n2343 585
R3467 gnd.n3711 gnd.n3710 585
R3468 gnd.n3712 gnd.n3711 585
R3469 gnd.n3709 gnd.n2354 585
R3470 gnd.n2354 gnd.n2352 585
R3471 gnd.n3708 gnd.n3707 585
R3472 gnd.n3707 gnd.n3706 585
R3473 gnd.n2356 gnd.n2355 585
R3474 gnd.n2519 gnd.n2356 585
R3475 gnd.n3693 gnd.n3692 585
R3476 gnd.n3694 gnd.n3693 585
R3477 gnd.n3691 gnd.n2367 585
R3478 gnd.n3686 gnd.n2367 585
R3479 gnd.n3690 gnd.n3689 585
R3480 gnd.n3689 gnd.n3688 585
R3481 gnd.n2369 gnd.n2368 585
R3482 gnd.n3674 gnd.n2369 585
R3483 gnd.n3659 gnd.n2390 585
R3484 gnd.n2390 gnd.n2379 585
R3485 gnd.n3661 gnd.n3660 585
R3486 gnd.n3662 gnd.n3661 585
R3487 gnd.n3658 gnd.n2389 585
R3488 gnd.n2389 gnd.n2386 585
R3489 gnd.n3657 gnd.n3656 585
R3490 gnd.n3656 gnd.n3655 585
R3491 gnd.n2392 gnd.n2391 585
R3492 gnd.n2533 gnd.n2392 585
R3493 gnd.n3644 gnd.n3643 585
R3494 gnd.n3645 gnd.n3644 585
R3495 gnd.n3642 gnd.n2404 585
R3496 gnd.n2404 gnd.n2400 585
R3497 gnd.n3640 gnd.n3639 585
R3498 gnd.n2426 gnd.n2425 585
R3499 gnd.n3636 gnd.n3635 585
R3500 gnd.n3637 gnd.n3636 585
R3501 gnd.n3634 gnd.n2461 585
R3502 gnd.n3633 gnd.n3632 585
R3503 gnd.n3631 gnd.n3630 585
R3504 gnd.n3629 gnd.n3628 585
R3505 gnd.n3627 gnd.n3626 585
R3506 gnd.n3625 gnd.n3624 585
R3507 gnd.n3623 gnd.n3622 585
R3508 gnd.n3621 gnd.n3620 585
R3509 gnd.n3619 gnd.n3618 585
R3510 gnd.n3617 gnd.n3616 585
R3511 gnd.n3615 gnd.n3614 585
R3512 gnd.n3613 gnd.n3612 585
R3513 gnd.n3611 gnd.n3610 585
R3514 gnd.n3609 gnd.n3608 585
R3515 gnd.n3607 gnd.n3606 585
R3516 gnd.n3605 gnd.n3604 585
R3517 gnd.n3603 gnd.n3602 585
R3518 gnd.n3601 gnd.n3600 585
R3519 gnd.n3599 gnd.n3598 585
R3520 gnd.n3597 gnd.n3596 585
R3521 gnd.n3595 gnd.n3594 585
R3522 gnd.n3593 gnd.n3592 585
R3523 gnd.n3591 gnd.n3590 585
R3524 gnd.n3589 gnd.n3588 585
R3525 gnd.n3587 gnd.n3586 585
R3526 gnd.n3585 gnd.n3584 585
R3527 gnd.n3583 gnd.n3582 585
R3528 gnd.n3581 gnd.n3580 585
R3529 gnd.n3579 gnd.n3578 585
R3530 gnd.n3577 gnd.n3576 585
R3531 gnd.n3575 gnd.n2602 585
R3532 gnd.n2601 gnd.n2600 585
R3533 gnd.n2599 gnd.n2598 585
R3534 gnd.n2596 gnd.n2595 585
R3535 gnd.n2594 gnd.n2593 585
R3536 gnd.n2592 gnd.n2591 585
R3537 gnd.n2590 gnd.n2589 585
R3538 gnd.n2588 gnd.n2587 585
R3539 gnd.n2586 gnd.n2585 585
R3540 gnd.n2584 gnd.n2583 585
R3541 gnd.n2582 gnd.n2581 585
R3542 gnd.n2580 gnd.n2579 585
R3543 gnd.n2578 gnd.n2577 585
R3544 gnd.n2576 gnd.n2575 585
R3545 gnd.n2574 gnd.n2573 585
R3546 gnd.n2572 gnd.n2571 585
R3547 gnd.n2570 gnd.n2569 585
R3548 gnd.n2568 gnd.n2567 585
R3549 gnd.n2566 gnd.n2565 585
R3550 gnd.n2564 gnd.n2563 585
R3551 gnd.n2562 gnd.n2561 585
R3552 gnd.n2560 gnd.n2559 585
R3553 gnd.n2558 gnd.n2557 585
R3554 gnd.n2556 gnd.n2555 585
R3555 gnd.n2554 gnd.n2553 585
R3556 gnd.n2552 gnd.n2551 585
R3557 gnd.n2550 gnd.n2549 585
R3558 gnd.n2548 gnd.n2547 585
R3559 gnd.n2546 gnd.n2545 585
R3560 gnd.n2544 gnd.n2543 585
R3561 gnd.n2542 gnd.n2541 585
R3562 gnd.n2540 gnd.n2539 585
R3563 gnd.n4301 gnd.n4300 585
R3564 gnd.n4303 gnd.n4302 585
R3565 gnd.n4305 gnd.n4304 585
R3566 gnd.n4307 gnd.n4306 585
R3567 gnd.n4309 gnd.n4308 585
R3568 gnd.n4311 gnd.n4310 585
R3569 gnd.n4313 gnd.n4312 585
R3570 gnd.n4315 gnd.n4314 585
R3571 gnd.n4317 gnd.n4316 585
R3572 gnd.n4319 gnd.n4318 585
R3573 gnd.n4321 gnd.n4320 585
R3574 gnd.n4323 gnd.n4322 585
R3575 gnd.n4325 gnd.n4324 585
R3576 gnd.n4327 gnd.n4326 585
R3577 gnd.n4329 gnd.n4328 585
R3578 gnd.n4331 gnd.n4330 585
R3579 gnd.n4333 gnd.n4332 585
R3580 gnd.n4335 gnd.n4334 585
R3581 gnd.n4337 gnd.n4336 585
R3582 gnd.n4339 gnd.n4338 585
R3583 gnd.n4341 gnd.n4340 585
R3584 gnd.n4343 gnd.n4342 585
R3585 gnd.n4345 gnd.n4344 585
R3586 gnd.n4347 gnd.n4346 585
R3587 gnd.n4349 gnd.n4348 585
R3588 gnd.n4351 gnd.n4350 585
R3589 gnd.n4353 gnd.n4352 585
R3590 gnd.n4355 gnd.n4354 585
R3591 gnd.n4357 gnd.n4356 585
R3592 gnd.n4360 gnd.n4359 585
R3593 gnd.n4362 gnd.n4361 585
R3594 gnd.n4364 gnd.n4363 585
R3595 gnd.n4366 gnd.n4365 585
R3596 gnd.n4230 gnd.n2031 585
R3597 gnd.n4232 gnd.n4231 585
R3598 gnd.n4234 gnd.n4233 585
R3599 gnd.n4236 gnd.n4235 585
R3600 gnd.n4239 gnd.n4238 585
R3601 gnd.n4241 gnd.n4240 585
R3602 gnd.n4243 gnd.n4242 585
R3603 gnd.n4245 gnd.n4244 585
R3604 gnd.n4247 gnd.n4246 585
R3605 gnd.n4249 gnd.n4248 585
R3606 gnd.n4251 gnd.n4250 585
R3607 gnd.n4253 gnd.n4252 585
R3608 gnd.n4255 gnd.n4254 585
R3609 gnd.n4257 gnd.n4256 585
R3610 gnd.n4259 gnd.n4258 585
R3611 gnd.n4261 gnd.n4260 585
R3612 gnd.n4263 gnd.n4262 585
R3613 gnd.n4265 gnd.n4264 585
R3614 gnd.n4267 gnd.n4266 585
R3615 gnd.n4269 gnd.n4268 585
R3616 gnd.n4271 gnd.n4270 585
R3617 gnd.n4273 gnd.n4272 585
R3618 gnd.n4275 gnd.n4274 585
R3619 gnd.n4277 gnd.n4276 585
R3620 gnd.n4279 gnd.n4278 585
R3621 gnd.n4281 gnd.n4280 585
R3622 gnd.n4283 gnd.n4282 585
R3623 gnd.n4285 gnd.n4284 585
R3624 gnd.n4287 gnd.n4286 585
R3625 gnd.n4289 gnd.n4288 585
R3626 gnd.n4291 gnd.n4290 585
R3627 gnd.n4293 gnd.n4292 585
R3628 gnd.n4294 gnd.n2039 585
R3629 gnd.n4299 gnd.n2034 585
R3630 gnd.n4299 gnd.n4298 585
R3631 gnd.n4115 gnd.n2035 585
R3632 gnd.n2046 gnd.n2035 585
R3633 gnd.n4116 gnd.n2043 585
R3634 gnd.n4205 gnd.n2043 585
R3635 gnd.n4119 gnd.n4118 585
R3636 gnd.n4118 gnd.n4117 585
R3637 gnd.n4120 gnd.n2055 585
R3638 gnd.n4189 gnd.n2055 585
R3639 gnd.n4122 gnd.n4121 585
R3640 gnd.n4121 gnd.n2053 585
R3641 gnd.n4123 gnd.n2061 585
R3642 gnd.n4183 gnd.n2061 585
R3643 gnd.n4127 gnd.n4126 585
R3644 gnd.n4126 gnd.n4125 585
R3645 gnd.n4128 gnd.n2069 585
R3646 gnd.n4165 gnd.n2069 585
R3647 gnd.n4130 gnd.n4129 585
R3648 gnd.n4129 gnd.n2068 585
R3649 gnd.n4131 gnd.n2074 585
R3650 gnd.n4159 gnd.n2074 585
R3651 gnd.n4135 gnd.n4134 585
R3652 gnd.n4134 gnd.n4133 585
R3653 gnd.n4136 gnd.n2082 585
R3654 gnd.n4147 gnd.n2082 585
R3655 gnd.n4138 gnd.n4137 585
R3656 gnd.n4139 gnd.n4138 585
R3657 gnd.n4114 gnd.n2088 585
R3658 gnd.n4141 gnd.n2088 585
R3659 gnd.n4113 gnd.n4112 585
R3660 gnd.n4112 gnd.n4111 585
R3661 gnd.n2090 gnd.n2089 585
R3662 gnd.n2109 gnd.n2090 585
R3663 gnd.n4055 gnd.n2100 585
R3664 gnd.n4096 gnd.n2100 585
R3665 gnd.n4057 gnd.n4056 585
R3666 gnd.n4056 gnd.n2099 585
R3667 gnd.n4058 gnd.n2106 585
R3668 gnd.n4089 gnd.n2106 585
R3669 gnd.n4061 gnd.n4060 585
R3670 gnd.n4060 gnd.n4059 585
R3671 gnd.n4062 gnd.n2117 585
R3672 gnd.n4073 gnd.n2117 585
R3673 gnd.n4064 gnd.n4063 585
R3674 gnd.n4065 gnd.n4064 585
R3675 gnd.n4054 gnd.n2122 585
R3676 gnd.n4067 gnd.n2122 585
R3677 gnd.n4053 gnd.n4052 585
R3678 gnd.n4052 gnd.n4051 585
R3679 gnd.n2124 gnd.n2123 585
R3680 gnd.n2136 gnd.n2124 585
R3681 gnd.n3962 gnd.n2133 585
R3682 gnd.n4040 gnd.n2133 585
R3683 gnd.n3964 gnd.n3963 585
R3684 gnd.n3963 gnd.n2131 585
R3685 gnd.n3965 gnd.n2141 585
R3686 gnd.n4033 gnd.n2141 585
R3687 gnd.n3970 gnd.n3969 585
R3688 gnd.n3969 gnd.n3968 585
R3689 gnd.n3971 gnd.n2149 585
R3690 gnd.n4008 gnd.n2149 585
R3691 gnd.n3973 gnd.n3972 585
R3692 gnd.n3972 gnd.n2148 585
R3693 gnd.n3974 gnd.n2155 585
R3694 gnd.n4002 gnd.n2155 585
R3695 gnd.n3978 gnd.n3977 585
R3696 gnd.n3977 gnd.n3976 585
R3697 gnd.n3979 gnd.n2164 585
R3698 gnd.n3990 gnd.n2164 585
R3699 gnd.n3980 gnd.n2171 585
R3700 gnd.n2171 gnd.n2163 585
R3701 gnd.n3982 gnd.n3981 585
R3702 gnd.n3984 gnd.n3982 585
R3703 gnd.n3961 gnd.n2170 585
R3704 gnd.n2182 gnd.n2170 585
R3705 gnd.n3960 gnd.n3959 585
R3706 gnd.n3959 gnd.n3958 585
R3707 gnd.n2173 gnd.n2172 585
R3708 gnd.n3950 gnd.n2173 585
R3709 gnd.n2235 gnd.n2179 585
R3710 gnd.n3952 gnd.n2179 585
R3711 gnd.n2236 gnd.n2190 585
R3712 gnd.n3938 gnd.n2190 585
R3713 gnd.n2238 gnd.n2237 585
R3714 gnd.n2237 gnd.n2189 585
R3715 gnd.n2239 gnd.n2198 585
R3716 gnd.n3913 gnd.n2198 585
R3717 gnd.n2241 gnd.n2240 585
R3718 gnd.n2240 gnd.n2197 585
R3719 gnd.n2242 gnd.n2205 585
R3720 gnd.n3906 gnd.n2205 585
R3721 gnd.n2246 gnd.n2245 585
R3722 gnd.n2245 gnd.n2244 585
R3723 gnd.n2247 gnd.n2212 585
R3724 gnd.n3896 gnd.n2212 585
R3725 gnd.n2249 gnd.n2248 585
R3726 gnd.n2248 gnd.n2211 585
R3727 gnd.n2250 gnd.n2219 585
R3728 gnd.n3890 gnd.n2219 585
R3729 gnd.n3865 gnd.n3864 585
R3730 gnd.n3864 gnd.n3863 585
R3731 gnd.n3866 gnd.n2228 585
R3732 gnd.n3878 gnd.n2228 585
R3733 gnd.n3868 gnd.n3867 585
R3734 gnd.n3869 gnd.n3868 585
R3735 gnd.n2234 gnd.n2233 585
R3736 gnd.n3872 gnd.n2233 585
R3737 gnd.n3850 gnd.n3849 585
R3738 gnd.n3851 gnd.n3850 585
R3739 gnd.n3848 gnd.n2258 585
R3740 gnd.n2258 gnd.n2256 585
R3741 gnd.n3847 gnd.n3846 585
R3742 gnd.n3846 gnd.n3845 585
R3743 gnd.n2260 gnd.n2259 585
R3744 gnd.n3804 gnd.n2260 585
R3745 gnd.n2467 gnd.n2269 585
R3746 gnd.n3838 gnd.n2269 585
R3747 gnd.n2471 gnd.n2470 585
R3748 gnd.n2470 gnd.n2469 585
R3749 gnd.n2472 gnd.n2276 585
R3750 gnd.n3826 gnd.n2276 585
R3751 gnd.n2474 gnd.n2473 585
R3752 gnd.n2473 gnd.n2275 585
R3753 gnd.n2475 gnd.n2282 585
R3754 gnd.n3820 gnd.n2282 585
R3755 gnd.n2479 gnd.n2478 585
R3756 gnd.n2478 gnd.n2477 585
R3757 gnd.n2480 gnd.n2289 585
R3758 gnd.n3795 gnd.n2289 585
R3759 gnd.n2482 gnd.n2481 585
R3760 gnd.n2481 gnd.n2296 585
R3761 gnd.n2483 gnd.n2295 585
R3762 gnd.n3789 gnd.n2295 585
R3763 gnd.n2486 gnd.n2485 585
R3764 gnd.n2485 gnd.n2484 585
R3765 gnd.n2487 gnd.n2303 585
R3766 gnd.n3776 gnd.n2303 585
R3767 gnd.n2488 gnd.n2311 585
R3768 gnd.n3768 gnd.n2311 585
R3769 gnd.n2489 gnd.n2310 585
R3770 gnd.n3770 gnd.n2310 585
R3771 gnd.n2491 gnd.n2490 585
R3772 gnd.n2491 gnd.n2319 585
R3773 gnd.n2494 gnd.n2493 585
R3774 gnd.n2493 gnd.n2492 585
R3775 gnd.n2495 gnd.n2326 585
R3776 gnd.n3747 gnd.n2326 585
R3777 gnd.n2497 gnd.n2496 585
R3778 gnd.n2496 gnd.n2325 585
R3779 gnd.n2498 gnd.n2333 585
R3780 gnd.n3740 gnd.n2333 585
R3781 gnd.n2503 gnd.n2502 585
R3782 gnd.n2502 gnd.n2501 585
R3783 gnd.n2504 gnd.n2339 585
R3784 gnd.n3730 gnd.n2339 585
R3785 gnd.n2507 gnd.n2506 585
R3786 gnd.n2506 gnd.n2505 585
R3787 gnd.n2508 gnd.n2345 585
R3788 gnd.n3724 gnd.n2345 585
R3789 gnd.n2513 gnd.n2512 585
R3790 gnd.n2512 gnd.n2511 585
R3791 gnd.n2514 gnd.n2353 585
R3792 gnd.n3712 gnd.n2353 585
R3793 gnd.n2516 gnd.n2515 585
R3794 gnd.n2515 gnd.n2352 585
R3795 gnd.n2517 gnd.n2358 585
R3796 gnd.n3706 gnd.n2358 585
R3797 gnd.n2521 gnd.n2520 585
R3798 gnd.n2520 gnd.n2519 585
R3799 gnd.n2522 gnd.n2366 585
R3800 gnd.n3694 gnd.n2366 585
R3801 gnd.n2523 gnd.n2372 585
R3802 gnd.n3686 gnd.n2372 585
R3803 gnd.n2524 gnd.n2371 585
R3804 gnd.n3688 gnd.n2371 585
R3805 gnd.n2525 gnd.n2380 585
R3806 gnd.n3674 gnd.n2380 585
R3807 gnd.n2527 gnd.n2526 585
R3808 gnd.n2526 gnd.n2379 585
R3809 gnd.n2528 gnd.n2387 585
R3810 gnd.n3662 gnd.n2387 585
R3811 gnd.n2530 gnd.n2529 585
R3812 gnd.n2529 gnd.n2386 585
R3813 gnd.n2531 gnd.n2394 585
R3814 gnd.n3655 gnd.n2394 585
R3815 gnd.n2535 gnd.n2534 585
R3816 gnd.n2534 gnd.n2533 585
R3817 gnd.n2536 gnd.n2401 585
R3818 gnd.n3645 gnd.n2401 585
R3819 gnd.n2538 gnd.n2537 585
R3820 gnd.n2538 gnd.n2400 585
R3821 gnd.n2860 gnd.n2859 585
R3822 gnd.n2859 gnd.n1108 585
R3823 gnd.n7394 gnd.n7392 585
R3824 gnd.n7394 gnd.n7393 585
R3825 gnd.n7396 gnd.n7395 585
R3826 gnd.n7395 gnd.n225 585
R3827 gnd.n7397 gnd.n317 585
R3828 gnd.n317 gnd.n233 585
R3829 gnd.n7456 gnd.n7398 585
R3830 gnd.n7456 gnd.n7455 585
R3831 gnd.n7457 gnd.n316 585
R3832 gnd.n7457 gnd.n241 585
R3833 gnd.n7459 gnd.n7458 585
R3834 gnd.n7458 gnd.n239 585
R3835 gnd.n7460 gnd.n311 585
R3836 gnd.n311 gnd.n249 585
R3837 gnd.n7462 gnd.n7461 585
R3838 gnd.n7462 gnd.n247 585
R3839 gnd.n7463 gnd.n310 585
R3840 gnd.n7463 gnd.n257 585
R3841 gnd.n7465 gnd.n7464 585
R3842 gnd.n7464 gnd.n255 585
R3843 gnd.n7466 gnd.n307 585
R3844 gnd.n307 gnd.n264 585
R3845 gnd.n7469 gnd.n7468 585
R3846 gnd.n7470 gnd.n7469 585
R3847 gnd.n308 gnd.n306 585
R3848 gnd.n306 gnd.n296 585
R3849 gnd.n4651 gnd.n4650 585
R3850 gnd.n4650 gnd.n294 585
R3851 gnd.n4652 gnd.n4647 585
R3852 gnd.n4647 gnd.n4646 585
R3853 gnd.n4655 gnd.n4654 585
R3854 gnd.n4656 gnd.n4655 585
R3855 gnd.n4648 gnd.n1540 585
R3856 gnd.n1544 gnd.n1540 585
R3857 gnd.n4664 gnd.n4663 585
R3858 gnd.n4663 gnd.n4662 585
R3859 gnd.n4665 gnd.n1538 585
R3860 gnd.n4633 gnd.n1538 585
R3861 gnd.n4668 gnd.n4667 585
R3862 gnd.n4668 gnd.n280 585
R3863 gnd.n4669 gnd.n1537 585
R3864 gnd.n4669 gnd.n277 585
R3865 gnd.n4671 gnd.n4670 585
R3866 gnd.n4670 gnd.n1520 585
R3867 gnd.n4672 gnd.n1531 585
R3868 gnd.n1531 gnd.n1530 585
R3869 gnd.n4674 gnd.n4673 585
R3870 gnd.n4675 gnd.n4674 585
R3871 gnd.n1532 gnd.n1529 585
R3872 gnd.n4608 gnd.n1529 585
R3873 gnd.n4579 gnd.n4578 585
R3874 gnd.n4579 gnd.n1561 585
R3875 gnd.n4581 gnd.n4580 585
R3876 gnd.n4580 gnd.n1569 585
R3877 gnd.n4582 gnd.n1584 585
R3878 gnd.n1584 gnd.n1583 585
R3879 gnd.n4584 gnd.n4583 585
R3880 gnd.n4585 gnd.n4584 585
R3881 gnd.n1585 gnd.n1582 585
R3882 gnd.n1582 gnd.n1578 585
R3883 gnd.n4570 gnd.n4569 585
R3884 gnd.n4569 gnd.n4568 585
R3885 gnd.n1588 gnd.n1587 585
R3886 gnd.n1598 gnd.n1588 585
R3887 gnd.n4542 gnd.n1611 585
R3888 gnd.n1611 gnd.n1610 585
R3889 gnd.n4544 gnd.n4543 585
R3890 gnd.n4545 gnd.n4544 585
R3891 gnd.n1612 gnd.n1609 585
R3892 gnd.n1609 gnd.n1605 585
R3893 gnd.n4537 gnd.n4536 585
R3894 gnd.n4536 gnd.n4535 585
R3895 gnd.n1615 gnd.n1614 585
R3896 gnd.n4517 gnd.n1615 585
R3897 gnd.n1633 gnd.n1632 585
R3898 gnd.n1634 gnd.n1633 585
R3899 gnd.n1625 gnd.n1624 585
R3900 gnd.n1624 gnd.n1493 585
R3901 gnd.n1628 gnd.n1627 585
R3902 gnd.n1627 gnd.n1490 585
R3903 gnd.n1475 gnd.n1474 585
R3904 gnd.n1480 gnd.n1475 585
R3905 gnd.n4724 gnd.n4723 585
R3906 gnd.n4723 gnd.n4722 585
R3907 gnd.n4725 gnd.n1469 585
R3908 gnd.n1476 gnd.n1469 585
R3909 gnd.n4727 gnd.n4726 585
R3910 gnd.n4728 gnd.n4727 585
R3911 gnd.n1466 gnd.n1465 585
R3912 gnd.n4729 gnd.n1466 585
R3913 gnd.n4732 gnd.n4731 585
R3914 gnd.n4731 gnd.n4730 585
R3915 gnd.n4733 gnd.n1460 585
R3916 gnd.n1460 gnd.n1458 585
R3917 gnd.n4735 gnd.n4734 585
R3918 gnd.n4736 gnd.n4735 585
R3919 gnd.n1461 gnd.n1459 585
R3920 gnd.n1459 gnd.n1456 585
R3921 gnd.n4448 gnd.n4447 585
R3922 gnd.n4449 gnd.n4448 585
R3923 gnd.n1804 gnd.n1803 585
R3924 gnd.n4438 gnd.n1803 585
R3925 gnd.n4442 gnd.n4441 585
R3926 gnd.n4441 gnd.n4440 585
R3927 gnd.n1807 gnd.n1806 585
R3928 gnd.n4426 gnd.n1807 585
R3929 gnd.n4424 gnd.n4423 585
R3930 gnd.n4425 gnd.n4424 585
R3931 gnd.n1817 gnd.n1816 585
R3932 gnd.n4415 gnd.n1816 585
R3933 gnd.n4419 gnd.n4418 585
R3934 gnd.n4418 gnd.n4417 585
R3935 gnd.n1820 gnd.n1819 585
R3936 gnd.n4406 gnd.n1820 585
R3937 gnd.n4404 gnd.n4403 585
R3938 gnd.n4405 gnd.n4404 585
R3939 gnd.n1830 gnd.n1829 585
R3940 gnd.n4395 gnd.n1829 585
R3941 gnd.n4399 gnd.n4398 585
R3942 gnd.n4398 gnd.n4397 585
R3943 gnd.n1833 gnd.n1832 585
R3944 gnd.n4386 gnd.n1833 585
R3945 gnd.n4384 gnd.n4383 585
R3946 gnd.n4385 gnd.n4384 585
R3947 gnd.n1843 gnd.n1842 585
R3948 gnd.n4375 gnd.n1842 585
R3949 gnd.n4379 gnd.n4378 585
R3950 gnd.n4378 gnd.n4377 585
R3951 gnd.n1846 gnd.n1845 585
R3952 gnd.n1871 gnd.n1846 585
R3953 gnd.n4200 gnd.n4199 585
R3954 gnd.n4199 gnd.n1852 585
R3955 gnd.n4201 gnd.n2048 585
R3956 gnd.n2048 gnd.n2047 585
R3957 gnd.n4203 gnd.n4202 585
R3958 gnd.n4204 gnd.n4203 585
R3959 gnd.n2049 gnd.n2045 585
R3960 gnd.n2056 gnd.n2045 585
R3961 gnd.n4193 gnd.n4192 585
R3962 gnd.n4192 gnd.n4191 585
R3963 gnd.n2052 gnd.n2051 585
R3964 gnd.n2060 gnd.n2052 585
R3965 gnd.n4155 gnd.n2076 585
R3966 gnd.n2076 gnd.n2070 585
R3967 gnd.n4157 gnd.n4156 585
R3968 gnd.n4158 gnd.n4157 585
R3969 gnd.n2077 gnd.n2075 585
R3970 gnd.n4132 gnd.n2075 585
R3971 gnd.n4150 gnd.n4149 585
R3972 gnd.n4149 gnd.n4148 585
R3973 gnd.n2080 gnd.n2079 585
R3974 gnd.n4140 gnd.n2080 585
R3975 gnd.n4083 gnd.n4082 585
R3976 gnd.n4082 gnd.n2091 585
R3977 gnd.n4084 gnd.n2111 585
R3978 gnd.n2111 gnd.n2110 585
R3979 gnd.n4086 gnd.n4085 585
R3980 gnd.n4087 gnd.n4086 585
R3981 gnd.n2112 gnd.n2107 585
R3982 gnd.n2107 gnd.n2105 585
R3983 gnd.n4076 gnd.n4075 585
R3984 gnd.n4075 gnd.n4074 585
R3985 gnd.n2115 gnd.n2114 585
R3986 gnd.n4066 gnd.n2115 585
R3987 gnd.n4049 gnd.n4048 585
R3988 gnd.n4050 gnd.n4049 585
R3989 gnd.n2127 gnd.n2126 585
R3990 gnd.n2134 gnd.n2126 585
R3991 gnd.n4044 gnd.n4043 585
R3992 gnd.n4043 gnd.n4042 585
R3993 gnd.n2130 gnd.n2129 585
R3994 gnd.n2140 gnd.n2130 585
R3995 gnd.n3998 gnd.n2157 585
R3996 gnd.n2157 gnd.n2150 585
R3997 gnd.n4000 gnd.n3999 585
R3998 gnd.n4001 gnd.n4000 585
R3999 gnd.n2158 gnd.n2156 585
R4000 gnd.n3975 gnd.n2156 585
R4001 gnd.n3993 gnd.n3992 585
R4002 gnd.n3992 gnd.n3991 585
R4003 gnd.n2161 gnd.n2160 585
R4004 gnd.n3983 gnd.n2161 585
R4005 gnd.n3946 gnd.n2184 585
R4006 gnd.n2184 gnd.n2183 585
R4007 gnd.n3948 gnd.n3947 585
R4008 gnd.n3949 gnd.n3948 585
R4009 gnd.n2185 gnd.n2181 585
R4010 gnd.n2181 gnd.n2178 585
R4011 gnd.n3941 gnd.n3940 585
R4012 gnd.n3940 gnd.n3939 585
R4013 gnd.n2188 gnd.n2187 585
R4014 gnd.n3914 gnd.n2188 585
R4015 gnd.n3904 gnd.n3903 585
R4016 gnd.n3905 gnd.n3904 585
R4017 gnd.n2207 gnd.n2206 585
R4018 gnd.n2243 gnd.n2206 585
R4019 gnd.n3899 gnd.n3898 585
R4020 gnd.n3898 gnd.n3897 585
R4021 gnd.n2210 gnd.n2209 585
R4022 gnd.n3889 gnd.n2210 585
R4023 gnd.n3861 gnd.n3860 585
R4024 gnd.n3862 gnd.n3861 585
R4025 gnd.n2252 gnd.n2251 585
R4026 gnd.n2251 gnd.n2227 585
R4027 gnd.n3856 gnd.n3855 585
R4028 gnd.n3855 gnd.n2232 585
R4029 gnd.n3854 gnd.n2254 585
R4030 gnd.n3854 gnd.n3853 585
R4031 gnd.n3834 gnd.n2255 585
R4032 gnd.n2261 gnd.n2255 585
R4033 gnd.n3836 gnd.n3835 585
R4034 gnd.n3837 gnd.n3836 585
R4035 gnd.n2271 gnd.n2270 585
R4036 gnd.n2468 gnd.n2270 585
R4037 gnd.n3829 gnd.n3828 585
R4038 gnd.n3828 gnd.n3827 585
R4039 gnd.n2274 gnd.n2273 585
R4040 gnd.n2281 gnd.n2274 585
R4041 gnd.n3784 gnd.n2298 585
R4042 gnd.n2298 gnd.n2290 585
R4043 gnd.n3786 gnd.n3785 585
R4044 gnd.n3787 gnd.n3786 585
R4045 gnd.n2299 gnd.n2297 585
R4046 gnd.n2297 gnd.n2294 585
R4047 gnd.n3779 gnd.n3778 585
R4048 gnd.n3778 gnd.n3777 585
R4049 gnd.n2302 gnd.n2301 585
R4050 gnd.n3769 gnd.n2302 585
R4051 gnd.n3756 gnd.n3755 585
R4052 gnd.n3757 gnd.n3756 585
R4053 gnd.n2321 gnd.n2320 585
R4054 gnd.n2327 gnd.n2320 585
R4055 gnd.n3751 gnd.n3750 585
R4056 gnd.n3750 gnd.n3749 585
R4057 gnd.n2324 gnd.n2323 585
R4058 gnd.n2332 gnd.n2324 585
R4059 gnd.n3720 gnd.n2347 585
R4060 gnd.n2347 gnd.n2340 585
R4061 gnd.n3722 gnd.n3721 585
R4062 gnd.n3723 gnd.n3722 585
R4063 gnd.n2348 gnd.n2346 585
R4064 gnd.n2510 gnd.n2346 585
R4065 gnd.n3715 gnd.n3714 585
R4066 gnd.n3714 gnd.n3713 585
R4067 gnd.n2351 gnd.n2350 585
R4068 gnd.n3705 gnd.n2351 585
R4069 gnd.n3682 gnd.n2374 585
R4070 gnd.n2518 gnd.n2374 585
R4071 gnd.n3684 gnd.n3683 585
R4072 gnd.n3685 gnd.n3684 585
R4073 gnd.n2375 gnd.n2373 585
R4074 gnd.n2373 gnd.n2370 585
R4075 gnd.n3677 gnd.n3676 585
R4076 gnd.n3676 gnd.n3675 585
R4077 gnd.n2378 gnd.n2377 585
R4078 gnd.n3663 gnd.n2378 585
R4079 gnd.n3653 gnd.n3652 585
R4080 gnd.n3654 gnd.n3653 585
R4081 gnd.n2396 gnd.n2395 585
R4082 gnd.n2532 gnd.n2395 585
R4083 gnd.n3648 gnd.n3647 585
R4084 gnd.n3647 gnd.n3646 585
R4085 gnd.n2399 gnd.n2398 585
R4086 gnd.n3471 gnd.n2399 585
R4087 gnd.n3464 gnd.n2749 585
R4088 gnd.n2749 gnd.n2427 585
R4089 gnd.n3466 gnd.n3465 585
R4090 gnd.n3467 gnd.n3466 585
R4091 gnd.n2750 gnd.n2748 585
R4092 gnd.n3455 gnd.n2748 585
R4093 gnd.n3459 gnd.n3458 585
R4094 gnd.n3458 gnd.n3457 585
R4095 gnd.n2753 gnd.n2752 585
R4096 gnd.n3453 gnd.n2753 585
R4097 gnd.n3450 gnd.n3449 585
R4098 gnd.n3451 gnd.n3450 585
R4099 gnd.n2755 gnd.n2754 585
R4100 gnd.n3441 gnd.n2754 585
R4101 gnd.n3445 gnd.n3444 585
R4102 gnd.n3444 gnd.n3443 585
R4103 gnd.n2758 gnd.n2757 585
R4104 gnd.n3436 gnd.n2758 585
R4105 gnd.n3433 gnd.n3432 585
R4106 gnd.n3434 gnd.n3433 585
R4107 gnd.n2763 gnd.n2762 585
R4108 gnd.n3424 gnd.n2762 585
R4109 gnd.n3428 gnd.n3427 585
R4110 gnd.n3427 gnd.n3426 585
R4111 gnd.n2766 gnd.n2765 585
R4112 gnd.n3422 gnd.n2766 585
R4113 gnd.n3419 gnd.n3418 585
R4114 gnd.n3420 gnd.n3419 585
R4115 gnd.n2771 gnd.n2770 585
R4116 gnd.n3410 gnd.n2770 585
R4117 gnd.n3414 gnd.n3413 585
R4118 gnd.n3413 gnd.n3412 585
R4119 gnd.n2774 gnd.n2773 585
R4120 gnd.n3408 gnd.n2774 585
R4121 gnd.n3405 gnd.n3404 585
R4122 gnd.n3406 gnd.n3405 585
R4123 gnd.n2777 gnd.n2776 585
R4124 gnd.n2776 gnd.n2775 585
R4125 gnd.n3400 gnd.n3399 585
R4126 gnd.n3399 gnd.n3398 585
R4127 gnd.n2780 gnd.n2779 585
R4128 gnd.n3264 gnd.n2780 585
R4129 gnd.n3262 gnd.n3261 585
R4130 gnd.n3263 gnd.n3262 585
R4131 gnd.n2782 gnd.n2781 585
R4132 gnd.n2781 gnd.n1323 585
R4133 gnd.n3257 gnd.n3256 585
R4134 gnd.n3256 gnd.n1320 585
R4135 gnd.n3255 gnd.n2784 585
R4136 gnd.n3255 gnd.n2701 585
R4137 gnd.n3254 gnd.n3253 585
R4138 gnd.n3254 gnd.n1311 585
R4139 gnd.n2786 gnd.n2785 585
R4140 gnd.n2785 gnd.n1303 585
R4141 gnd.n3249 gnd.n3248 585
R4142 gnd.n3248 gnd.n1300 585
R4143 gnd.n3247 gnd.n2788 585
R4144 gnd.n3247 gnd.n1292 585
R4145 gnd.n3246 gnd.n3245 585
R4146 gnd.n3246 gnd.n1289 585
R4147 gnd.n2790 gnd.n2789 585
R4148 gnd.n2789 gnd.n1281 585
R4149 gnd.n3241 gnd.n3240 585
R4150 gnd.n3240 gnd.n1278 585
R4151 gnd.n3239 gnd.n2792 585
R4152 gnd.n3239 gnd.n3238 585
R4153 gnd.n2898 gnd.n2793 585
R4154 gnd.n2793 gnd.n1268 585
R4155 gnd.n2900 gnd.n2899 585
R4156 gnd.n2900 gnd.n2808 585
R4157 gnd.n2902 gnd.n2901 585
R4158 gnd.n2901 gnd.n1258 585
R4159 gnd.n2903 gnd.n2891 585
R4160 gnd.n2891 gnd.n1250 585
R4161 gnd.n2905 gnd.n2904 585
R4162 gnd.n2905 gnd.n1247 585
R4163 gnd.n2906 gnd.n2890 585
R4164 gnd.n2906 gnd.n1239 585
R4165 gnd.n2908 gnd.n2907 585
R4166 gnd.n2907 gnd.n1236 585
R4167 gnd.n2909 gnd.n2885 585
R4168 gnd.n2885 gnd.n2818 585
R4169 gnd.n2911 gnd.n2910 585
R4170 gnd.n2911 gnd.n1226 585
R4171 gnd.n2912 gnd.n2884 585
R4172 gnd.n2912 gnd.n2822 585
R4173 gnd.n2914 gnd.n2913 585
R4174 gnd.n2913 gnd.n1216 585
R4175 gnd.n2915 gnd.n2882 585
R4176 gnd.n2882 gnd.n1209 585
R4177 gnd.n2917 gnd.n2916 585
R4178 gnd.n2917 gnd.n1206 585
R4179 gnd.n2919 gnd.n2918 585
R4180 gnd.n2918 gnd.n1198 585
R4181 gnd.n2921 gnd.n2920 585
R4182 gnd.n2921 gnd.n1195 585
R4183 gnd.n2923 gnd.n2922 585
R4184 gnd.n2922 gnd.n2832 585
R4185 gnd.n2925 gnd.n2924 585
R4186 gnd.n2925 gnd.n1188 585
R4187 gnd.n2927 gnd.n2926 585
R4188 gnd.n2927 gnd.n2837 585
R4189 gnd.n2928 gnd.n2881 585
R4190 gnd.n2928 gnd.n1178 585
R4191 gnd.n2930 gnd.n2929 585
R4192 gnd.n2929 gnd.n1172 585
R4193 gnd.n2876 gnd.n2875 585
R4194 gnd.n2875 gnd.n1169 585
R4195 gnd.n2936 gnd.n2935 585
R4196 gnd.n2936 gnd.n1161 585
R4197 gnd.n2937 gnd.n2874 585
R4198 gnd.n2937 gnd.n1158 585
R4199 gnd.n2939 gnd.n2938 585
R4200 gnd.n2938 gnd.n2847 585
R4201 gnd.n2940 gnd.n2852 585
R4202 gnd.n2852 gnd.n1148 585
R4203 gnd.n2942 gnd.n2941 585
R4204 gnd.n2943 gnd.n2942 585
R4205 gnd.n2853 gnd.n2851 585
R4206 gnd.n2851 gnd.n1138 585
R4207 gnd.n2868 gnd.n2867 585
R4208 gnd.n2867 gnd.n1130 585
R4209 gnd.n2866 gnd.n2855 585
R4210 gnd.n2866 gnd.n1127 585
R4211 gnd.n2865 gnd.n2864 585
R4212 gnd.n2865 gnd.n1119 585
R4213 gnd.n2857 gnd.n2856 585
R4214 gnd.n2856 gnd.n1116 585
R4215 gnd.n4739 gnd.n4738 585
R4216 gnd.n4738 gnd.n4737 585
R4217 gnd.n4740 gnd.n1454 585
R4218 gnd.n4450 gnd.n1454 585
R4219 gnd.n4436 gnd.n1452 585
R4220 gnd.n4437 gnd.n4436 585
R4221 gnd.n4744 gnd.n1451 585
R4222 gnd.n4439 gnd.n1451 585
R4223 gnd.n4745 gnd.n1450 585
R4224 gnd.n1808 gnd.n1450 585
R4225 gnd.n4746 gnd.n1449 585
R4226 gnd.n4427 gnd.n1449 585
R4227 gnd.n1814 gnd.n1447 585
R4228 gnd.n1815 gnd.n1814 585
R4229 gnd.n4750 gnd.n1446 585
R4230 gnd.n4416 gnd.n1446 585
R4231 gnd.n4751 gnd.n1445 585
R4232 gnd.n1821 gnd.n1445 585
R4233 gnd.n4752 gnd.n1444 585
R4234 gnd.n4407 gnd.n1444 585
R4235 gnd.n1827 gnd.n1442 585
R4236 gnd.n1828 gnd.n1827 585
R4237 gnd.n4756 gnd.n1441 585
R4238 gnd.n4396 gnd.n1441 585
R4239 gnd.n4757 gnd.n1440 585
R4240 gnd.n1834 gnd.n1440 585
R4241 gnd.n4758 gnd.n1439 585
R4242 gnd.n4387 gnd.n1439 585
R4243 gnd.n1840 gnd.n1437 585
R4244 gnd.n1841 gnd.n1840 585
R4245 gnd.n4762 gnd.n1436 585
R4246 gnd.n4376 gnd.n1436 585
R4247 gnd.n4763 gnd.n1435 585
R4248 gnd.n1870 gnd.n1435 585
R4249 gnd.n4764 gnd.n1434 585
R4250 gnd.n4367 gnd.n1434 585
R4251 gnd.n2036 gnd.n1432 585
R4252 gnd.n2037 gnd.n2036 585
R4253 gnd.n4768 gnd.n1431 585
R4254 gnd.n2044 gnd.n1431 585
R4255 gnd.n4769 gnd.n1430 585
R4256 gnd.n2042 gnd.n1430 585
R4257 gnd.n4770 gnd.n1429 585
R4258 gnd.n4190 gnd.n1429 585
R4259 gnd.n4181 gnd.n1427 585
R4260 gnd.n4182 gnd.n4181 585
R4261 gnd.n4774 gnd.n1426 585
R4262 gnd.n4124 gnd.n1426 585
R4263 gnd.n4775 gnd.n1425 585
R4264 gnd.n4166 gnd.n1425 585
R4265 gnd.n4776 gnd.n1424 585
R4266 gnd.n4159 gnd.n1424 585
R4267 gnd.n2083 gnd.n1422 585
R4268 gnd.n2084 gnd.n2083 585
R4269 gnd.n4780 gnd.n1421 585
R4270 gnd.n2081 gnd.n1421 585
R4271 gnd.n4781 gnd.n1420 585
R4272 gnd.n4110 gnd.n1420 585
R4273 gnd.n4782 gnd.n1419 585
R4274 gnd.n2108 gnd.n1419 585
R4275 gnd.n4097 gnd.n1417 585
R4276 gnd.n4098 gnd.n4097 585
R4277 gnd.n4786 gnd.n1416 585
R4278 gnd.n4088 gnd.n1416 585
R4279 gnd.n4787 gnd.n1415 585
R4280 gnd.n2118 gnd.n1415 585
R4281 gnd.n4788 gnd.n1414 585
R4282 gnd.n2116 gnd.n1414 585
R4283 gnd.n4016 gnd.n1412 585
R4284 gnd.n4017 gnd.n4016 585
R4285 gnd.n4792 gnd.n1411 585
R4286 gnd.n2125 gnd.n1411 585
R4287 gnd.n4793 gnd.n1410 585
R4288 gnd.n4041 gnd.n1410 585
R4289 gnd.n4794 gnd.n1409 585
R4290 gnd.n4032 gnd.n1409 585
R4291 gnd.n3966 gnd.n1407 585
R4292 gnd.n3967 gnd.n3966 585
R4293 gnd.n4798 gnd.n1406 585
R4294 gnd.n4009 gnd.n1406 585
R4295 gnd.n4799 gnd.n1405 585
R4296 gnd.n2154 gnd.n1405 585
R4297 gnd.n4800 gnd.n1404 585
R4298 gnd.n2165 gnd.n1404 585
R4299 gnd.n2162 gnd.n1402 585
R4300 gnd.n2163 gnd.n2162 585
R4301 gnd.n4804 gnd.n1401 585
R4302 gnd.n2169 gnd.n1401 585
R4303 gnd.n4805 gnd.n1400 585
R4304 gnd.n2174 gnd.n1400 585
R4305 gnd.n4806 gnd.n1399 585
R4306 gnd.n3951 gnd.n1399 585
R4307 gnd.n3936 gnd.n1397 585
R4308 gnd.n3937 gnd.n3936 585
R4309 gnd.n4810 gnd.n1396 585
R4310 gnd.n2199 gnd.n1396 585
R4311 gnd.n4811 gnd.n1395 585
R4312 gnd.n3915 gnd.n1395 585
R4313 gnd.n4812 gnd.n1394 585
R4314 gnd.n2204 gnd.n1394 585
R4315 gnd.n2213 gnd.n1392 585
R4316 gnd.n2214 gnd.n2213 585
R4317 gnd.n4816 gnd.n1391 585
R4318 gnd.n3888 gnd.n1391 585
R4319 gnd.n4817 gnd.n1390 585
R4320 gnd.n2218 gnd.n1390 585
R4321 gnd.n4818 gnd.n1389 585
R4322 gnd.n3879 gnd.n1389 585
R4323 gnd.n3870 gnd.n1387 585
R4324 gnd.n3871 gnd.n3870 585
R4325 gnd.n4822 gnd.n1386 585
R4326 gnd.n3852 gnd.n1386 585
R4327 gnd.n4823 gnd.n1385 585
R4328 gnd.n2262 gnd.n1385 585
R4329 gnd.n4824 gnd.n1384 585
R4330 gnd.n3805 gnd.n1384 585
R4331 gnd.n2267 gnd.n1382 585
R4332 gnd.n2268 gnd.n2267 585
R4333 gnd.n4828 gnd.n1381 585
R4334 gnd.n3826 gnd.n1381 585
R4335 gnd.n4829 gnd.n1380 585
R4336 gnd.n3819 gnd.n1380 585
R4337 gnd.n4830 gnd.n1379 585
R4338 gnd.n2476 gnd.n1379 585
R4339 gnd.n3796 gnd.n1377 585
R4340 gnd.n3797 gnd.n3796 585
R4341 gnd.n4834 gnd.n1376 585
R4342 gnd.n3788 gnd.n1376 585
R4343 gnd.n4835 gnd.n1375 585
R4344 gnd.n2304 gnd.n1375 585
R4345 gnd.n4836 gnd.n1374 585
R4346 gnd.n3767 gnd.n1374 585
R4347 gnd.n2308 gnd.n1372 585
R4348 gnd.n2309 gnd.n2308 585
R4349 gnd.n4840 gnd.n1371 585
R4350 gnd.n3758 gnd.n1371 585
R4351 gnd.n4841 gnd.n1370 585
R4352 gnd.n3748 gnd.n1370 585
R4353 gnd.n4842 gnd.n1369 585
R4354 gnd.n3739 gnd.n1369 585
R4355 gnd.n2499 gnd.n1367 585
R4356 gnd.n2500 gnd.n2499 585
R4357 gnd.n4846 gnd.n1366 585
R4358 gnd.n3731 gnd.n1366 585
R4359 gnd.n4847 gnd.n1365 585
R4360 gnd.n2344 gnd.n1365 585
R4361 gnd.n4848 gnd.n1364 585
R4362 gnd.n2509 gnd.n1364 585
R4363 gnd.n3703 gnd.n1362 585
R4364 gnd.n3704 gnd.n3703 585
R4365 gnd.n4852 gnd.n1361 585
R4366 gnd.n2357 gnd.n1361 585
R4367 gnd.n4853 gnd.n1360 585
R4368 gnd.n3694 gnd.n1360 585
R4369 gnd.n4854 gnd.n1359 585
R4370 gnd.n3687 gnd.n1359 585
R4371 gnd.n3672 gnd.n1357 585
R4372 gnd.n3673 gnd.n3672 585
R4373 gnd.n4858 gnd.n1356 585
R4374 gnd.n2388 gnd.n1356 585
R4375 gnd.n4859 gnd.n1355 585
R4376 gnd.n3664 gnd.n1355 585
R4377 gnd.n4860 gnd.n1354 585
R4378 gnd.n2393 gnd.n1354 585
R4379 gnd.n2402 gnd.n1352 585
R4380 gnd.n2403 gnd.n2402 585
R4381 gnd.n4864 gnd.n1351 585
R4382 gnd.n3472 gnd.n1351 585
R4383 gnd.n4865 gnd.n1350 585
R4384 gnd.n2460 gnd.n1350 585
R4385 gnd.n4866 gnd.n1349 585
R4386 gnd.n3468 gnd.n1349 585
R4387 gnd.n2746 gnd.n1347 585
R4388 gnd.n2747 gnd.n2746 585
R4389 gnd.n4870 gnd.n1346 585
R4390 gnd.n3456 gnd.n1346 585
R4391 gnd.n4871 gnd.n1345 585
R4392 gnd.n3454 gnd.n1345 585
R4393 gnd.n4872 gnd.n1344 585
R4394 gnd.n3452 gnd.n1344 585
R4395 gnd.n3439 gnd.n1342 585
R4396 gnd.n3440 gnd.n3439 585
R4397 gnd.n4876 gnd.n1341 585
R4398 gnd.n3442 gnd.n1341 585
R4399 gnd.n4877 gnd.n1340 585
R4400 gnd.n3437 gnd.n1340 585
R4401 gnd.n4878 gnd.n1339 585
R4402 gnd.n3435 gnd.n1339 585
R4403 gnd.n2760 gnd.n1337 585
R4404 gnd.n2761 gnd.n2760 585
R4405 gnd.n4882 gnd.n1336 585
R4406 gnd.n3425 gnd.n1336 585
R4407 gnd.n4883 gnd.n1335 585
R4408 gnd.n3423 gnd.n1335 585
R4409 gnd.n4884 gnd.n1334 585
R4410 gnd.n3421 gnd.n1334 585
R4411 gnd.n2768 gnd.n1332 585
R4412 gnd.n2769 gnd.n2768 585
R4413 gnd.n4888 gnd.n1331 585
R4414 gnd.n3411 gnd.n1331 585
R4415 gnd.n4889 gnd.n1330 585
R4416 gnd.n3409 gnd.n1330 585
R4417 gnd.n4890 gnd.n1329 585
R4418 gnd.n3407 gnd.n1329 585
R4419 gnd.n3395 gnd.n3394 585
R4420 gnd.n3393 gnd.n3281 585
R4421 gnd.n3283 gnd.n3280 585
R4422 gnd.n3397 gnd.n3280 585
R4423 gnd.n3386 gnd.n3296 585
R4424 gnd.n3385 gnd.n3297 585
R4425 gnd.n3299 gnd.n3298 585
R4426 gnd.n3378 gnd.n3307 585
R4427 gnd.n3377 gnd.n3308 585
R4428 gnd.n3318 gnd.n3309 585
R4429 gnd.n3370 gnd.n3319 585
R4430 gnd.n3369 gnd.n3320 585
R4431 gnd.n3322 gnd.n3321 585
R4432 gnd.n3362 gnd.n3330 585
R4433 gnd.n3361 gnd.n3331 585
R4434 gnd.n3343 gnd.n3332 585
R4435 gnd.n3354 gnd.n3344 585
R4436 gnd.n3353 gnd.n3346 585
R4437 gnd.n3345 gnd.n2707 585
R4438 gnd.n3521 gnd.n2708 585
R4439 gnd.n3520 gnd.n2709 585
R4440 gnd.n3519 gnd.n2710 585
R4441 gnd.n3274 gnd.n2711 585
R4442 gnd.n3515 gnd.n2713 585
R4443 gnd.n3514 gnd.n2714 585
R4444 gnd.n3513 gnd.n2715 585
R4445 gnd.n3510 gnd.n2720 585
R4446 gnd.n3509 gnd.n2721 585
R4447 gnd.n3508 gnd.n2722 585
R4448 gnd.n3278 gnd.n2723 585
R4449 gnd.n4453 gnd.n1457 585
R4450 gnd.n4737 gnd.n1457 585
R4451 gnd.n4452 gnd.n4451 585
R4452 gnd.n4451 gnd.n4450 585
R4453 gnd.n1802 gnd.n1801 585
R4454 gnd.n4437 gnd.n1802 585
R4455 gnd.n4435 gnd.n4434 585
R4456 gnd.n4439 gnd.n4435 585
R4457 gnd.n1810 gnd.n1809 585
R4458 gnd.n1809 gnd.n1808 585
R4459 gnd.n4429 gnd.n4428 585
R4460 gnd.n4428 gnd.n4427 585
R4461 gnd.n1813 gnd.n1812 585
R4462 gnd.n1815 gnd.n1813 585
R4463 gnd.n4414 gnd.n4413 585
R4464 gnd.n4416 gnd.n4414 585
R4465 gnd.n1823 gnd.n1822 585
R4466 gnd.n1822 gnd.n1821 585
R4467 gnd.n4409 gnd.n4408 585
R4468 gnd.n4408 gnd.n4407 585
R4469 gnd.n1826 gnd.n1825 585
R4470 gnd.n1828 gnd.n1826 585
R4471 gnd.n4394 gnd.n4393 585
R4472 gnd.n4396 gnd.n4394 585
R4473 gnd.n1836 gnd.n1835 585
R4474 gnd.n1835 gnd.n1834 585
R4475 gnd.n4389 gnd.n4388 585
R4476 gnd.n4388 gnd.n4387 585
R4477 gnd.n1839 gnd.n1838 585
R4478 gnd.n1841 gnd.n1839 585
R4479 gnd.n4374 gnd.n4373 585
R4480 gnd.n4376 gnd.n4374 585
R4481 gnd.n1848 gnd.n1847 585
R4482 gnd.n1870 gnd.n1847 585
R4483 gnd.n4369 gnd.n4368 585
R4484 gnd.n4368 gnd.n4367 585
R4485 gnd.n1851 gnd.n1850 585
R4486 gnd.n2037 gnd.n1851 585
R4487 gnd.n4174 gnd.n4173 585
R4488 gnd.n4173 gnd.n2044 585
R4489 gnd.n4175 gnd.n4172 585
R4490 gnd.n4172 gnd.n2042 585
R4491 gnd.n2064 gnd.n2054 585
R4492 gnd.n4190 gnd.n2054 585
R4493 gnd.n4180 gnd.n4179 585
R4494 gnd.n4182 gnd.n4180 585
R4495 gnd.n2063 gnd.n2062 585
R4496 gnd.n4124 gnd.n2062 585
R4497 gnd.n4168 gnd.n4167 585
R4498 gnd.n4167 gnd.n4166 585
R4499 gnd.n2067 gnd.n2066 585
R4500 gnd.n4159 gnd.n2067 585
R4501 gnd.n4104 gnd.n4103 585
R4502 gnd.n4103 gnd.n2084 585
R4503 gnd.n2095 gnd.n2093 585
R4504 gnd.n2093 gnd.n2081 585
R4505 gnd.n4109 gnd.n4108 585
R4506 gnd.n4110 gnd.n4109 585
R4507 gnd.n2094 gnd.n2092 585
R4508 gnd.n2108 gnd.n2092 585
R4509 gnd.n4100 gnd.n4099 585
R4510 gnd.n4099 gnd.n4098 585
R4511 gnd.n2098 gnd.n2097 585
R4512 gnd.n4088 gnd.n2098 585
R4513 gnd.n4021 gnd.n4020 585
R4514 gnd.n4020 gnd.n2118 585
R4515 gnd.n4024 gnd.n4019 585
R4516 gnd.n4019 gnd.n2116 585
R4517 gnd.n4025 gnd.n4018 585
R4518 gnd.n4018 gnd.n4017 585
R4519 gnd.n4026 gnd.n4015 585
R4520 gnd.n4015 gnd.n2125 585
R4521 gnd.n2144 gnd.n2132 585
R4522 gnd.n4041 gnd.n2132 585
R4523 gnd.n4031 gnd.n4030 585
R4524 gnd.n4032 gnd.n4031 585
R4525 gnd.n2143 gnd.n2142 585
R4526 gnd.n3967 gnd.n2142 585
R4527 gnd.n4011 gnd.n4010 585
R4528 gnd.n4010 gnd.n4009 585
R4529 gnd.n2147 gnd.n2146 585
R4530 gnd.n2154 gnd.n2147 585
R4531 gnd.n3925 gnd.n3924 585
R4532 gnd.n3924 gnd.n2165 585
R4533 gnd.n3928 gnd.n3923 585
R4534 gnd.n3923 gnd.n2163 585
R4535 gnd.n3929 gnd.n3922 585
R4536 gnd.n3922 gnd.n2169 585
R4537 gnd.n3930 gnd.n3921 585
R4538 gnd.n3921 gnd.n2174 585
R4539 gnd.n2193 gnd.n2180 585
R4540 gnd.n3951 gnd.n2180 585
R4541 gnd.n3935 gnd.n3934 585
R4542 gnd.n3937 gnd.n3935 585
R4543 gnd.n2192 gnd.n2191 585
R4544 gnd.n2199 gnd.n2191 585
R4545 gnd.n3917 gnd.n3916 585
R4546 gnd.n3916 gnd.n3915 585
R4547 gnd.n2196 gnd.n2195 585
R4548 gnd.n2204 gnd.n2196 585
R4549 gnd.n2223 gnd.n2221 585
R4550 gnd.n2221 gnd.n2214 585
R4551 gnd.n3887 gnd.n3886 585
R4552 gnd.n3888 gnd.n3887 585
R4553 gnd.n2222 gnd.n2220 585
R4554 gnd.n2220 gnd.n2218 585
R4555 gnd.n3881 gnd.n3880 585
R4556 gnd.n3880 gnd.n3879 585
R4557 gnd.n2226 gnd.n2225 585
R4558 gnd.n3871 gnd.n2226 585
R4559 gnd.n3808 gnd.n2257 585
R4560 gnd.n3852 gnd.n2257 585
R4561 gnd.n3811 gnd.n3807 585
R4562 gnd.n3807 gnd.n2262 585
R4563 gnd.n3812 gnd.n3806 585
R4564 gnd.n3806 gnd.n3805 585
R4565 gnd.n3813 gnd.n3803 585
R4566 gnd.n3803 gnd.n2268 585
R4567 gnd.n2285 gnd.n2277 585
R4568 gnd.n3826 gnd.n2277 585
R4569 gnd.n3818 gnd.n3817 585
R4570 gnd.n3819 gnd.n3818 585
R4571 gnd.n2284 gnd.n2283 585
R4572 gnd.n2476 gnd.n2283 585
R4573 gnd.n3799 gnd.n3798 585
R4574 gnd.n3798 gnd.n3797 585
R4575 gnd.n2288 gnd.n2287 585
R4576 gnd.n3788 gnd.n2288 585
R4577 gnd.n2315 gnd.n2313 585
R4578 gnd.n2313 gnd.n2304 585
R4579 gnd.n3766 gnd.n3765 585
R4580 gnd.n3767 gnd.n3766 585
R4581 gnd.n2314 gnd.n2312 585
R4582 gnd.n2312 gnd.n2309 585
R4583 gnd.n3760 gnd.n3759 585
R4584 gnd.n3759 gnd.n3758 585
R4585 gnd.n2318 gnd.n2317 585
R4586 gnd.n3748 gnd.n2318 585
R4587 gnd.n3738 gnd.n3737 585
R4588 gnd.n3739 gnd.n3738 585
R4589 gnd.n2335 gnd.n2334 585
R4590 gnd.n2500 gnd.n2334 585
R4591 gnd.n3733 gnd.n3732 585
R4592 gnd.n3732 gnd.n3731 585
R4593 gnd.n2338 gnd.n2337 585
R4594 gnd.n2344 gnd.n2338 585
R4595 gnd.n2362 gnd.n2360 585
R4596 gnd.n2509 gnd.n2360 585
R4597 gnd.n3702 gnd.n3701 585
R4598 gnd.n3704 gnd.n3702 585
R4599 gnd.n2361 gnd.n2359 585
R4600 gnd.n2359 gnd.n2357 585
R4601 gnd.n3696 gnd.n3695 585
R4602 gnd.n3695 gnd.n3694 585
R4603 gnd.n2365 gnd.n2364 585
R4604 gnd.n3687 gnd.n2365 585
R4605 gnd.n3671 gnd.n3670 585
R4606 gnd.n3673 gnd.n3671 585
R4607 gnd.n2382 gnd.n2381 585
R4608 gnd.n2388 gnd.n2381 585
R4609 gnd.n3666 gnd.n3665 585
R4610 gnd.n3665 gnd.n3664 585
R4611 gnd.n2385 gnd.n2384 585
R4612 gnd.n2393 gnd.n2385 585
R4613 gnd.n3475 gnd.n3474 585
R4614 gnd.n3474 gnd.n2403 585
R4615 gnd.n3478 gnd.n3473 585
R4616 gnd.n3473 gnd.n3472 585
R4617 gnd.n3479 gnd.n3470 585
R4618 gnd.n3470 gnd.n2460 585
R4619 gnd.n3480 gnd.n3469 585
R4620 gnd.n3469 gnd.n3468 585
R4621 gnd.n2745 gnd.n2743 585
R4622 gnd.n2747 gnd.n2745 585
R4623 gnd.n3484 gnd.n2742 585
R4624 gnd.n3456 gnd.n2742 585
R4625 gnd.n3485 gnd.n2741 585
R4626 gnd.n3454 gnd.n2741 585
R4627 gnd.n3486 gnd.n2740 585
R4628 gnd.n3452 gnd.n2740 585
R4629 gnd.n3438 gnd.n2738 585
R4630 gnd.n3440 gnd.n3438 585
R4631 gnd.n3490 gnd.n2737 585
R4632 gnd.n3442 gnd.n2737 585
R4633 gnd.n3491 gnd.n2736 585
R4634 gnd.n3437 gnd.n2736 585
R4635 gnd.n3492 gnd.n2735 585
R4636 gnd.n3435 gnd.n2735 585
R4637 gnd.n2759 gnd.n2733 585
R4638 gnd.n2761 gnd.n2759 585
R4639 gnd.n3496 gnd.n2732 585
R4640 gnd.n3425 gnd.n2732 585
R4641 gnd.n3497 gnd.n2731 585
R4642 gnd.n3423 gnd.n2731 585
R4643 gnd.n3498 gnd.n2730 585
R4644 gnd.n3421 gnd.n2730 585
R4645 gnd.n2767 gnd.n2728 585
R4646 gnd.n2769 gnd.n2767 585
R4647 gnd.n3502 gnd.n2727 585
R4648 gnd.n3411 gnd.n2727 585
R4649 gnd.n3503 gnd.n2726 585
R4650 gnd.n3409 gnd.n2726 585
R4651 gnd.n3504 gnd.n2725 585
R4652 gnd.n3407 gnd.n2725 585
R4653 gnd.n1799 gnd.n1798 585
R4654 gnd.n1798 gnd.n1467 585
R4655 gnd.n4457 gnd.n1797 585
R4656 gnd.n4458 gnd.n1795 585
R4657 gnd.n4459 gnd.n1794 585
R4658 gnd.n1792 gnd.n1787 585
R4659 gnd.n4463 gnd.n1786 585
R4660 gnd.n4464 gnd.n1784 585
R4661 gnd.n4465 gnd.n1783 585
R4662 gnd.n1781 gnd.n1779 585
R4663 gnd.n4469 gnd.n1778 585
R4664 gnd.n4470 gnd.n1776 585
R4665 gnd.n4471 gnd.n1775 585
R4666 gnd.n1773 gnd.n1650 585
R4667 gnd.n1772 gnd.n1771 585
R4668 gnd.n1756 gnd.n1652 585
R4669 gnd.n1758 gnd.n1757 585
R4670 gnd.n1754 gnd.n1659 585
R4671 gnd.n1753 gnd.n1752 585
R4672 gnd.n1737 gnd.n1661 585
R4673 gnd.n1739 gnd.n1738 585
R4674 gnd.n1735 gnd.n1668 585
R4675 gnd.n1734 gnd.n1733 585
R4676 gnd.n1718 gnd.n1670 585
R4677 gnd.n1720 gnd.n1719 585
R4678 gnd.n1716 gnd.n1677 585
R4679 gnd.n1715 gnd.n1714 585
R4680 gnd.n1699 gnd.n1679 585
R4681 gnd.n1701 gnd.n1700 585
R4682 gnd.n1697 gnd.n1455 585
R4683 gnd.n4297 gnd.n2039 482.89
R4684 gnd.n4300 gnd.n4299 482.89
R4685 gnd.n2539 gnd.n2538 482.89
R4686 gnd.n3639 gnd.n2404 482.89
R4687 gnd.n6693 gnd.n6692 457.279
R4688 gnd.n2465 gnd.t243 443.966
R4689 gnd.n2032 gnd.t256 443.966
R4690 gnd.n2462 gnd.t284 443.966
R4691 gnd.n4228 gnd.t209 443.966
R4692 gnd.n2716 gnd.t233 371.625
R4693 gnd.n7610 gnd.t259 371.625
R4694 gnd.n1645 gnd.t250 371.625
R4695 gnd.n3339 gnd.t272 371.625
R4696 gnd.n1948 gnd.t227 371.625
R4697 gnd.n1977 gnd.t213 371.625
R4698 gnd.n180 gnd.t278 371.625
R4699 gnd.n7703 gnd.t202 371.625
R4700 gnd.n1031 gnd.t186 371.625
R4701 gnd.n1053 gnd.t269 371.625
R4702 gnd.n2694 gnd.t275 371.625
R4703 gnd.n2605 gnd.t194 371.625
R4704 gnd.n2979 gnd.t220 371.625
R4705 gnd.n1789 gnd.t190 371.625
R4706 gnd.n5704 gnd.t265 323.425
R4707 gnd.n5158 gnd.t198 323.425
R4708 gnd.n6372 gnd.n6346 289.615
R4709 gnd.n6340 gnd.n6314 289.615
R4710 gnd.n6308 gnd.n6282 289.615
R4711 gnd.n6277 gnd.n6251 289.615
R4712 gnd.n6245 gnd.n6219 289.615
R4713 gnd.n6213 gnd.n6187 289.615
R4714 gnd.n6181 gnd.n6155 289.615
R4715 gnd.n6150 gnd.n6124 289.615
R4716 gnd.n5554 gnd.t223 279.217
R4717 gnd.n5184 gnd.t182 279.217
R4718 gnd.n2411 gnd.t264 260.649
R4719 gnd.n4220 gnd.t208 260.649
R4720 gnd.n3638 gnd.n3637 256.663
R4721 gnd.n3637 gnd.n2428 256.663
R4722 gnd.n3637 gnd.n2429 256.663
R4723 gnd.n3637 gnd.n2430 256.663
R4724 gnd.n3637 gnd.n2431 256.663
R4725 gnd.n3637 gnd.n2432 256.663
R4726 gnd.n3637 gnd.n2433 256.663
R4727 gnd.n3637 gnd.n2434 256.663
R4728 gnd.n3637 gnd.n2435 256.663
R4729 gnd.n3637 gnd.n2436 256.663
R4730 gnd.n3637 gnd.n2437 256.663
R4731 gnd.n3637 gnd.n2438 256.663
R4732 gnd.n3637 gnd.n2439 256.663
R4733 gnd.n3637 gnd.n2440 256.663
R4734 gnd.n3637 gnd.n2441 256.663
R4735 gnd.n3637 gnd.n2442 256.663
R4736 gnd.n3577 gnd.n3574 256.663
R4737 gnd.n3637 gnd.n2443 256.663
R4738 gnd.n3637 gnd.n2444 256.663
R4739 gnd.n3637 gnd.n2445 256.663
R4740 gnd.n3637 gnd.n2446 256.663
R4741 gnd.n3637 gnd.n2447 256.663
R4742 gnd.n3637 gnd.n2448 256.663
R4743 gnd.n3637 gnd.n2449 256.663
R4744 gnd.n3637 gnd.n2450 256.663
R4745 gnd.n3637 gnd.n2451 256.663
R4746 gnd.n3637 gnd.n2452 256.663
R4747 gnd.n3637 gnd.n2453 256.663
R4748 gnd.n3637 gnd.n2454 256.663
R4749 gnd.n3637 gnd.n2455 256.663
R4750 gnd.n3637 gnd.n2456 256.663
R4751 gnd.n3637 gnd.n2457 256.663
R4752 gnd.n3637 gnd.n2458 256.663
R4753 gnd.n3637 gnd.n2459 256.663
R4754 gnd.n4366 gnd.n1872 256.663
R4755 gnd.n4366 gnd.n1873 256.663
R4756 gnd.n4366 gnd.n1874 256.663
R4757 gnd.n4366 gnd.n1875 256.663
R4758 gnd.n4366 gnd.n1876 256.663
R4759 gnd.n4366 gnd.n1877 256.663
R4760 gnd.n4366 gnd.n1878 256.663
R4761 gnd.n4366 gnd.n1879 256.663
R4762 gnd.n4366 gnd.n1880 256.663
R4763 gnd.n4366 gnd.n1881 256.663
R4764 gnd.n4366 gnd.n1882 256.663
R4765 gnd.n4366 gnd.n1883 256.663
R4766 gnd.n4366 gnd.n1884 256.663
R4767 gnd.n4366 gnd.n1885 256.663
R4768 gnd.n4366 gnd.n1886 256.663
R4769 gnd.n4366 gnd.n1887 256.663
R4770 gnd.n2031 gnd.n1888 256.663
R4771 gnd.n4366 gnd.n1869 256.663
R4772 gnd.n4366 gnd.n1868 256.663
R4773 gnd.n4366 gnd.n1867 256.663
R4774 gnd.n4366 gnd.n1866 256.663
R4775 gnd.n4366 gnd.n1865 256.663
R4776 gnd.n4366 gnd.n1864 256.663
R4777 gnd.n4366 gnd.n1863 256.663
R4778 gnd.n4366 gnd.n1862 256.663
R4779 gnd.n4366 gnd.n1861 256.663
R4780 gnd.n4366 gnd.n1860 256.663
R4781 gnd.n4366 gnd.n1859 256.663
R4782 gnd.n4366 gnd.n1858 256.663
R4783 gnd.n4366 gnd.n1857 256.663
R4784 gnd.n4366 gnd.n1856 256.663
R4785 gnd.n4366 gnd.n1855 256.663
R4786 gnd.n4366 gnd.n1854 256.663
R4787 gnd.n4366 gnd.n1853 256.663
R4788 gnd.n5135 gnd.n999 242.672
R4789 gnd.n5135 gnd.n1000 242.672
R4790 gnd.n5135 gnd.n1001 242.672
R4791 gnd.n5135 gnd.n1002 242.672
R4792 gnd.n5135 gnd.n1003 242.672
R4793 gnd.n5135 gnd.n1004 242.672
R4794 gnd.n5135 gnd.n1005 242.672
R4795 gnd.n5135 gnd.n1006 242.672
R4796 gnd.n5135 gnd.n1007 242.672
R4797 gnd.n3348 gnd.n2666 242.672
R4798 gnd.n3337 gnd.n2666 242.672
R4799 gnd.n3334 gnd.n2666 242.672
R4800 gnd.n3325 gnd.n2666 242.672
R4801 gnd.n3314 gnd.n2666 242.672
R4802 gnd.n3311 gnd.n2666 242.672
R4803 gnd.n3302 gnd.n2666 242.672
R4804 gnd.n3292 gnd.n2666 242.672
R4805 gnd.n3289 gnd.n2666 242.672
R4806 gnd.n1686 gnd.n1468 242.672
R4807 gnd.n1706 gnd.n1468 242.672
R4808 gnd.n1708 gnd.n1468 242.672
R4809 gnd.n1725 gnd.n1468 242.672
R4810 gnd.n1727 gnd.n1468 242.672
R4811 gnd.n1744 gnd.n1468 242.672
R4812 gnd.n1746 gnd.n1468 242.672
R4813 gnd.n1763 gnd.n1468 242.672
R4814 gnd.n1765 gnd.n1468 242.672
R4815 gnd.n7612 gnd.n117 242.672
R4816 gnd.n7608 gnd.n117 242.672
R4817 gnd.n7603 gnd.n117 242.672
R4818 gnd.n7600 gnd.n117 242.672
R4819 gnd.n7595 gnd.n117 242.672
R4820 gnd.n7592 gnd.n117 242.672
R4821 gnd.n7587 gnd.n117 242.672
R4822 gnd.n7584 gnd.n117 242.672
R4823 gnd.n7579 gnd.n117 242.672
R4824 gnd.n5609 gnd.n5518 242.672
R4825 gnd.n5522 gnd.n5518 242.672
R4826 gnd.n5602 gnd.n5518 242.672
R4827 gnd.n5596 gnd.n5518 242.672
R4828 gnd.n5594 gnd.n5518 242.672
R4829 gnd.n5588 gnd.n5518 242.672
R4830 gnd.n5586 gnd.n5518 242.672
R4831 gnd.n5580 gnd.n5518 242.672
R4832 gnd.n5578 gnd.n5518 242.672
R4833 gnd.n5572 gnd.n5518 242.672
R4834 gnd.n5570 gnd.n5518 242.672
R4835 gnd.n5563 gnd.n5518 242.672
R4836 gnd.n5561 gnd.n5518 242.672
R4837 gnd.n6487 gnd.n980 242.672
R4838 gnd.n6487 gnd.n979 242.672
R4839 gnd.n6487 gnd.n978 242.672
R4840 gnd.n6487 gnd.n977 242.672
R4841 gnd.n6487 gnd.n976 242.672
R4842 gnd.n6487 gnd.n975 242.672
R4843 gnd.n6487 gnd.n974 242.672
R4844 gnd.n6487 gnd.n973 242.672
R4845 gnd.n6487 gnd.n972 242.672
R4846 gnd.n6487 gnd.n971 242.672
R4847 gnd.n6487 gnd.n970 242.672
R4848 gnd.n6487 gnd.n969 242.672
R4849 gnd.n6487 gnd.n968 242.672
R4850 gnd.n5738 gnd.n5737 242.672
R4851 gnd.n5738 gnd.n5679 242.672
R4852 gnd.n5738 gnd.n5680 242.672
R4853 gnd.n5738 gnd.n5681 242.672
R4854 gnd.n5738 gnd.n5682 242.672
R4855 gnd.n5738 gnd.n5683 242.672
R4856 gnd.n5738 gnd.n5684 242.672
R4857 gnd.n5738 gnd.n5685 242.672
R4858 gnd.n6487 gnd.n5136 242.672
R4859 gnd.n6487 gnd.n5137 242.672
R4860 gnd.n6487 gnd.n5138 242.672
R4861 gnd.n6487 gnd.n5139 242.672
R4862 gnd.n6487 gnd.n5140 242.672
R4863 gnd.n6487 gnd.n5141 242.672
R4864 gnd.n6487 gnd.n5142 242.672
R4865 gnd.n6487 gnd.n6486 242.672
R4866 gnd.n5135 gnd.n5134 242.672
R4867 gnd.n5135 gnd.n981 242.672
R4868 gnd.n5135 gnd.n982 242.672
R4869 gnd.n5135 gnd.n983 242.672
R4870 gnd.n5135 gnd.n984 242.672
R4871 gnd.n5135 gnd.n985 242.672
R4872 gnd.n5135 gnd.n986 242.672
R4873 gnd.n5135 gnd.n987 242.672
R4874 gnd.n5135 gnd.n988 242.672
R4875 gnd.n5135 gnd.n989 242.672
R4876 gnd.n5135 gnd.n990 242.672
R4877 gnd.n5135 gnd.n991 242.672
R4878 gnd.n5135 gnd.n992 242.672
R4879 gnd.n5135 gnd.n993 242.672
R4880 gnd.n5135 gnd.n994 242.672
R4881 gnd.n5135 gnd.n995 242.672
R4882 gnd.n5135 gnd.n996 242.672
R4883 gnd.n5135 gnd.n997 242.672
R4884 gnd.n5135 gnd.n998 242.672
R4885 gnd.n3536 gnd.n2666 242.672
R4886 gnd.n2697 gnd.n2666 242.672
R4887 gnd.n3543 gnd.n2666 242.672
R4888 gnd.n2688 gnd.n2666 242.672
R4889 gnd.n3550 gnd.n2666 242.672
R4890 gnd.n2681 gnd.n2666 242.672
R4891 gnd.n3557 gnd.n2666 242.672
R4892 gnd.n2674 gnd.n2666 242.672
R4893 gnd.n3564 gnd.n2666 242.672
R4894 gnd.n3567 gnd.n2666 242.672
R4895 gnd.n2666 gnd.n2612 242.672
R4896 gnd.n3573 gnd.n2607 242.672
R4897 gnd.n2666 gnd.n2613 242.672
R4898 gnd.n2666 gnd.n2614 242.672
R4899 gnd.n2666 gnd.n2615 242.672
R4900 gnd.n2666 gnd.n2616 242.672
R4901 gnd.n2666 gnd.n2617 242.672
R4902 gnd.n2666 gnd.n2618 242.672
R4903 gnd.n2666 gnd.n2619 242.672
R4904 gnd.n2666 gnd.n2665 242.672
R4905 gnd.n1910 gnd.n1468 242.672
R4906 gnd.n1918 gnd.n1468 242.672
R4907 gnd.n1920 gnd.n1468 242.672
R4908 gnd.n1928 gnd.n1468 242.672
R4909 gnd.n1930 gnd.n1468 242.672
R4910 gnd.n1939 gnd.n1468 242.672
R4911 gnd.n1942 gnd.n1468 242.672
R4912 gnd.n1893 gnd.n1468 242.672
R4913 gnd.n2030 gnd.n1890 242.672
R4914 gnd.n2027 gnd.n1468 242.672
R4915 gnd.n2025 gnd.n1468 242.672
R4916 gnd.n2019 gnd.n1468 242.672
R4917 gnd.n2017 gnd.n1468 242.672
R4918 gnd.n2011 gnd.n1468 242.672
R4919 gnd.n2009 gnd.n1468 242.672
R4920 gnd.n2003 gnd.n1468 242.672
R4921 gnd.n2001 gnd.n1468 242.672
R4922 gnd.n1995 gnd.n1468 242.672
R4923 gnd.n1993 gnd.n1468 242.672
R4924 gnd.n1985 gnd.n1468 242.672
R4925 gnd.n177 gnd.n117 242.672
R4926 gnd.n7671 gnd.n117 242.672
R4927 gnd.n173 gnd.n117 242.672
R4928 gnd.n7678 gnd.n117 242.672
R4929 gnd.n166 gnd.n117 242.672
R4930 gnd.n7685 gnd.n117 242.672
R4931 gnd.n159 gnd.n117 242.672
R4932 gnd.n7692 gnd.n117 242.672
R4933 gnd.n152 gnd.n117 242.672
R4934 gnd.n7699 gnd.n117 242.672
R4935 gnd.n145 gnd.n117 242.672
R4936 gnd.n7709 gnd.n117 242.672
R4937 gnd.n138 gnd.n117 242.672
R4938 gnd.n7716 gnd.n117 242.672
R4939 gnd.n131 gnd.n117 242.672
R4940 gnd.n7723 gnd.n117 242.672
R4941 gnd.n124 gnd.n117 242.672
R4942 gnd.n7730 gnd.n117 242.672
R4943 gnd.n117 gnd.n116 242.672
R4944 gnd.n3397 gnd.n3396 242.672
R4945 gnd.n3397 gnd.n3265 242.672
R4946 gnd.n3397 gnd.n3266 242.672
R4947 gnd.n3397 gnd.n3267 242.672
R4948 gnd.n3397 gnd.n3268 242.672
R4949 gnd.n3397 gnd.n3269 242.672
R4950 gnd.n3397 gnd.n3270 242.672
R4951 gnd.n3397 gnd.n3271 242.672
R4952 gnd.n3397 gnd.n3272 242.672
R4953 gnd.n3397 gnd.n3273 242.672
R4954 gnd.n3397 gnd.n3275 242.672
R4955 gnd.n3397 gnd.n3276 242.672
R4956 gnd.n3397 gnd.n3277 242.672
R4957 gnd.n3397 gnd.n3279 242.672
R4958 gnd.n1796 gnd.n1467 242.672
R4959 gnd.n1793 gnd.n1467 242.672
R4960 gnd.n1785 gnd.n1467 242.672
R4961 gnd.n1782 gnd.n1467 242.672
R4962 gnd.n1777 gnd.n1467 242.672
R4963 gnd.n1774 gnd.n1467 242.672
R4964 gnd.n1651 gnd.n1467 242.672
R4965 gnd.n1755 gnd.n1467 242.672
R4966 gnd.n1660 gnd.n1467 242.672
R4967 gnd.n1736 gnd.n1467 242.672
R4968 gnd.n1669 gnd.n1467 242.672
R4969 gnd.n1717 gnd.n1467 242.672
R4970 gnd.n1678 gnd.n1467 242.672
R4971 gnd.n1698 gnd.n1467 242.672
R4972 gnd.n113 gnd.n109 240.244
R4973 gnd.n7732 gnd.n7731 240.244
R4974 gnd.n7729 gnd.n118 240.244
R4975 gnd.n7725 gnd.n7724 240.244
R4976 gnd.n7722 gnd.n125 240.244
R4977 gnd.n7718 gnd.n7717 240.244
R4978 gnd.n7715 gnd.n132 240.244
R4979 gnd.n7711 gnd.n7710 240.244
R4980 gnd.n7708 gnd.n139 240.244
R4981 gnd.n7701 gnd.n7700 240.244
R4982 gnd.n7698 gnd.n146 240.244
R4983 gnd.n7694 gnd.n7693 240.244
R4984 gnd.n7691 gnd.n153 240.244
R4985 gnd.n7687 gnd.n7686 240.244
R4986 gnd.n7684 gnd.n160 240.244
R4987 gnd.n7680 gnd.n7679 240.244
R4988 gnd.n7677 gnd.n167 240.244
R4989 gnd.n7673 gnd.n7672 240.244
R4990 gnd.n7670 gnd.n174 240.244
R4991 gnd.n1984 gnd.n1478 240.244
R4992 gnd.n4485 gnd.n1478 240.244
R4993 gnd.n4485 gnd.n1491 240.244
R4994 gnd.n1636 gnd.n1491 240.244
R4995 gnd.n4516 gnd.n1636 240.244
R4996 gnd.n4516 gnd.n1637 240.244
R4997 gnd.n1637 gnd.n1617 240.244
R4998 gnd.n1617 gnd.n1606 240.244
R4999 gnd.n4510 gnd.n1606 240.244
R5000 gnd.n4510 gnd.n1597 240.244
R5001 gnd.n4507 gnd.n1597 240.244
R5002 gnd.n4507 gnd.n1590 240.244
R5003 gnd.n1590 gnd.n1579 240.244
R5004 gnd.n4503 gnd.n1579 240.244
R5005 gnd.n4503 gnd.n1568 240.244
R5006 gnd.n1568 gnd.n1560 240.244
R5007 gnd.n4610 gnd.n1560 240.244
R5008 gnd.n4610 gnd.n1526 240.244
R5009 gnd.n4613 gnd.n1526 240.244
R5010 gnd.n4613 gnd.n1518 240.244
R5011 gnd.n4621 gnd.n1518 240.244
R5012 gnd.n4621 gnd.n278 240.244
R5013 gnd.n4635 gnd.n278 240.244
R5014 gnd.n4636 gnd.n4635 240.244
R5015 gnd.n4636 gnd.n1542 240.244
R5016 gnd.n4642 gnd.n1542 240.244
R5017 gnd.n4642 gnd.n298 240.244
R5018 gnd.n7476 gnd.n298 240.244
R5019 gnd.n7476 gnd.n295 240.244
R5020 gnd.n7472 gnd.n295 240.244
R5021 gnd.n7472 gnd.n263 240.244
R5022 gnd.n7404 gnd.n263 240.244
R5023 gnd.n7404 gnd.n256 240.244
R5024 gnd.n7411 gnd.n256 240.244
R5025 gnd.n7411 gnd.n248 240.244
R5026 gnd.n7415 gnd.n248 240.244
R5027 gnd.n7415 gnd.n240 240.244
R5028 gnd.n7452 gnd.n240 240.244
R5029 gnd.n7452 gnd.n232 240.244
R5030 gnd.n7448 gnd.n232 240.244
R5031 gnd.n7448 gnd.n226 240.244
R5032 gnd.n7444 gnd.n226 240.244
R5033 gnd.n7444 gnd.n219 240.244
R5034 gnd.n7441 gnd.n219 240.244
R5035 gnd.n7441 gnd.n209 240.244
R5036 gnd.n7438 gnd.n209 240.244
R5037 gnd.n7438 gnd.n202 240.244
R5038 gnd.n7435 gnd.n202 240.244
R5039 gnd.n7435 gnd.n194 240.244
R5040 gnd.n194 gnd.n184 240.244
R5041 gnd.n7661 gnd.n184 240.244
R5042 gnd.n7662 gnd.n7661 240.244
R5043 gnd.n7662 gnd.n105 240.244
R5044 gnd.n1911 gnd.n1904 240.244
R5045 gnd.n1917 gnd.n1904 240.244
R5046 gnd.n1921 gnd.n1919 240.244
R5047 gnd.n1927 gnd.n1900 240.244
R5048 gnd.n1931 gnd.n1929 240.244
R5049 gnd.n1938 gnd.n1896 240.244
R5050 gnd.n1941 gnd.n1940 240.244
R5051 gnd.n1943 gnd.n1894 240.244
R5052 gnd.n2028 gnd.n2026 240.244
R5053 gnd.n2024 gnd.n1952 240.244
R5054 gnd.n2020 gnd.n2018 240.244
R5055 gnd.n2016 gnd.n1958 240.244
R5056 gnd.n2012 gnd.n2010 240.244
R5057 gnd.n2008 gnd.n1964 240.244
R5058 gnd.n2004 gnd.n2002 240.244
R5059 gnd.n2000 gnd.n1970 240.244
R5060 gnd.n1996 gnd.n1994 240.244
R5061 gnd.n1992 gnd.n1976 240.244
R5062 gnd.n4720 gnd.n1482 240.244
R5063 gnd.n4720 gnd.n1483 240.244
R5064 gnd.n4716 gnd.n1483 240.244
R5065 gnd.n4716 gnd.n1489 240.244
R5066 gnd.n4524 gnd.n1489 240.244
R5067 gnd.n4524 gnd.n4518 240.244
R5068 gnd.n4518 gnd.n1604 240.244
R5069 gnd.n4548 gnd.n1604 240.244
R5070 gnd.n4548 gnd.n1599 240.244
R5071 gnd.n4556 gnd.n1599 240.244
R5072 gnd.n4556 gnd.n1600 240.244
R5073 gnd.n1600 gnd.n1577 240.244
R5074 gnd.n4587 gnd.n1577 240.244
R5075 gnd.n4587 gnd.n1570 240.244
R5076 gnd.n4595 gnd.n1570 240.244
R5077 gnd.n4595 gnd.n1573 240.244
R5078 gnd.n1573 gnd.n1525 240.244
R5079 gnd.n4677 gnd.n1525 240.244
R5080 gnd.n4677 gnd.n1521 240.244
R5081 gnd.n4683 gnd.n1521 240.244
R5082 gnd.n4683 gnd.n275 240.244
R5083 gnd.n7499 gnd.n275 240.244
R5084 gnd.n7499 gnd.n276 240.244
R5085 gnd.n1545 gnd.n276 240.244
R5086 gnd.n4660 gnd.n1545 240.244
R5087 gnd.n4660 gnd.n4658 240.244
R5088 gnd.n4658 gnd.n297 240.244
R5089 gnd.n7478 gnd.n297 240.244
R5090 gnd.n7481 gnd.n7478 240.244
R5091 gnd.n7481 gnd.n265 240.244
R5092 gnd.n7504 gnd.n265 240.244
R5093 gnd.n7504 gnd.n254 240.244
R5094 gnd.n7514 gnd.n254 240.244
R5095 gnd.n7514 gnd.n250 240.244
R5096 gnd.n7520 gnd.n250 240.244
R5097 gnd.n7520 gnd.n238 240.244
R5098 gnd.n7530 gnd.n238 240.244
R5099 gnd.n7530 gnd.n234 240.244
R5100 gnd.n7536 gnd.n234 240.244
R5101 gnd.n7536 gnd.n224 240.244
R5102 gnd.n7546 gnd.n224 240.244
R5103 gnd.n7546 gnd.n220 240.244
R5104 gnd.n7552 gnd.n220 240.244
R5105 gnd.n7552 gnd.n207 240.244
R5106 gnd.n7562 gnd.n207 240.244
R5107 gnd.n7562 gnd.n203 240.244
R5108 gnd.n7568 gnd.n203 240.244
R5109 gnd.n7568 gnd.n192 240.244
R5110 gnd.n7653 gnd.n192 240.244
R5111 gnd.n7653 gnd.n188 240.244
R5112 gnd.n7659 gnd.n188 240.244
R5113 gnd.n7659 gnd.n108 240.244
R5114 gnd.n7739 gnd.n108 240.244
R5115 gnd.n2620 gnd.n1319 240.244
R5116 gnd.n2664 gnd.n2621 240.244
R5117 gnd.n2660 gnd.n2659 240.244
R5118 gnd.n2656 gnd.n2655 240.244
R5119 gnd.n2652 gnd.n2651 240.244
R5120 gnd.n2648 gnd.n2647 240.244
R5121 gnd.n2644 gnd.n2643 240.244
R5122 gnd.n2640 gnd.n2639 240.244
R5123 gnd.n3568 gnd.n2611 240.244
R5124 gnd.n3566 gnd.n3565 240.244
R5125 gnd.n3563 gnd.n2668 240.244
R5126 gnd.n3559 gnd.n3558 240.244
R5127 gnd.n3556 gnd.n2675 240.244
R5128 gnd.n3552 gnd.n3551 240.244
R5129 gnd.n3549 gnd.n2682 240.244
R5130 gnd.n3545 gnd.n3544 240.244
R5131 gnd.n3542 gnd.n2689 240.244
R5132 gnd.n3538 gnd.n3537 240.244
R5133 gnd.n5056 gnd.n1057 240.244
R5134 gnd.n1061 gnd.n1057 240.244
R5135 gnd.n5049 gnd.n1061 240.244
R5136 gnd.n5049 gnd.n1062 240.244
R5137 gnd.n1075 gnd.n1062 240.244
R5138 gnd.n3064 gnd.n1075 240.244
R5139 gnd.n3064 gnd.n1086 240.244
R5140 gnd.n3069 gnd.n1086 240.244
R5141 gnd.n3069 gnd.n1096 240.244
R5142 gnd.n3072 gnd.n1096 240.244
R5143 gnd.n3072 gnd.n1106 240.244
R5144 gnd.n3078 gnd.n1106 240.244
R5145 gnd.n3078 gnd.n1117 240.244
R5146 gnd.n3088 gnd.n1117 240.244
R5147 gnd.n3088 gnd.n1128 240.244
R5148 gnd.n3094 gnd.n1128 240.244
R5149 gnd.n3094 gnd.n1139 240.244
R5150 gnd.n3104 gnd.n1139 240.244
R5151 gnd.n3104 gnd.n1149 240.244
R5152 gnd.n3110 gnd.n1149 240.244
R5153 gnd.n3110 gnd.n1159 240.244
R5154 gnd.n3120 gnd.n1159 240.244
R5155 gnd.n3120 gnd.n1170 240.244
R5156 gnd.n3126 gnd.n1170 240.244
R5157 gnd.n3126 gnd.n1179 240.244
R5158 gnd.n3137 gnd.n1179 240.244
R5159 gnd.n3137 gnd.n1189 240.244
R5160 gnd.n3144 gnd.n1189 240.244
R5161 gnd.n3144 gnd.n1196 240.244
R5162 gnd.n3154 gnd.n1196 240.244
R5163 gnd.n3154 gnd.n1207 240.244
R5164 gnd.n3160 gnd.n1207 240.244
R5165 gnd.n3160 gnd.n1217 240.244
R5166 gnd.n3170 gnd.n1217 240.244
R5167 gnd.n3170 gnd.n1227 240.244
R5168 gnd.n3176 gnd.n1227 240.244
R5169 gnd.n3176 gnd.n1237 240.244
R5170 gnd.n3186 gnd.n1237 240.244
R5171 gnd.n3186 gnd.n1248 240.244
R5172 gnd.n3193 gnd.n1248 240.244
R5173 gnd.n3193 gnd.n1259 240.244
R5174 gnd.n3203 gnd.n1259 240.244
R5175 gnd.n3203 gnd.n1269 240.244
R5176 gnd.n2794 gnd.n1269 240.244
R5177 gnd.n2794 gnd.n1279 240.244
R5178 gnd.n3211 gnd.n1279 240.244
R5179 gnd.n3211 gnd.n1290 240.244
R5180 gnd.n3215 gnd.n1290 240.244
R5181 gnd.n3215 gnd.n1301 240.244
R5182 gnd.n3222 gnd.n1301 240.244
R5183 gnd.n3222 gnd.n1312 240.244
R5184 gnd.n3529 gnd.n1312 240.244
R5185 gnd.n3529 gnd.n1321 240.244
R5186 gnd.n1011 gnd.n1010 240.244
R5187 gnd.n5128 gnd.n1010 240.244
R5188 gnd.n5126 gnd.n5125 240.244
R5189 gnd.n5122 gnd.n5121 240.244
R5190 gnd.n5118 gnd.n5117 240.244
R5191 gnd.n5114 gnd.n5113 240.244
R5192 gnd.n5110 gnd.n5109 240.244
R5193 gnd.n5106 gnd.n5105 240.244
R5194 gnd.n5102 gnd.n5101 240.244
R5195 gnd.n5097 gnd.n5096 240.244
R5196 gnd.n5093 gnd.n5092 240.244
R5197 gnd.n5089 gnd.n5088 240.244
R5198 gnd.n5085 gnd.n5084 240.244
R5199 gnd.n5081 gnd.n5080 240.244
R5200 gnd.n5077 gnd.n5076 240.244
R5201 gnd.n5073 gnd.n5072 240.244
R5202 gnd.n5069 gnd.n5068 240.244
R5203 gnd.n5065 gnd.n5064 240.244
R5204 gnd.n1052 gnd.n1051 240.244
R5205 gnd.n3037 gnd.n1012 240.244
R5206 gnd.n3037 gnd.n1067 240.244
R5207 gnd.n5047 gnd.n1067 240.244
R5208 gnd.n5047 gnd.n1068 240.244
R5209 gnd.n5043 gnd.n1068 240.244
R5210 gnd.n5043 gnd.n1074 240.244
R5211 gnd.n5035 gnd.n1074 240.244
R5212 gnd.n5035 gnd.n1089 240.244
R5213 gnd.n5031 gnd.n1089 240.244
R5214 gnd.n5031 gnd.n1095 240.244
R5215 gnd.n5023 gnd.n1095 240.244
R5216 gnd.n5023 gnd.n1109 240.244
R5217 gnd.n5019 gnd.n1109 240.244
R5218 gnd.n5019 gnd.n1115 240.244
R5219 gnd.n5011 gnd.n1115 240.244
R5220 gnd.n5011 gnd.n1131 240.244
R5221 gnd.n5007 gnd.n1131 240.244
R5222 gnd.n5007 gnd.n1137 240.244
R5223 gnd.n4999 gnd.n1137 240.244
R5224 gnd.n4999 gnd.n1151 240.244
R5225 gnd.n4995 gnd.n1151 240.244
R5226 gnd.n4995 gnd.n1157 240.244
R5227 gnd.n4987 gnd.n1157 240.244
R5228 gnd.n4987 gnd.n1173 240.244
R5229 gnd.n4983 gnd.n1173 240.244
R5230 gnd.n4983 gnd.n1177 240.244
R5231 gnd.n4975 gnd.n1177 240.244
R5232 gnd.n4975 gnd.n1191 240.244
R5233 gnd.n4970 gnd.n1191 240.244
R5234 gnd.n4970 gnd.n1194 240.244
R5235 gnd.n4962 gnd.n1194 240.244
R5236 gnd.n4962 gnd.n1210 240.244
R5237 gnd.n4958 gnd.n1210 240.244
R5238 gnd.n4958 gnd.n1215 240.244
R5239 gnd.n4950 gnd.n1215 240.244
R5240 gnd.n4950 gnd.n1229 240.244
R5241 gnd.n4946 gnd.n1229 240.244
R5242 gnd.n4946 gnd.n1235 240.244
R5243 gnd.n4938 gnd.n1235 240.244
R5244 gnd.n4938 gnd.n1251 240.244
R5245 gnd.n4934 gnd.n1251 240.244
R5246 gnd.n4934 gnd.n1257 240.244
R5247 gnd.n4926 gnd.n1257 240.244
R5248 gnd.n4926 gnd.n1271 240.244
R5249 gnd.n4922 gnd.n1271 240.244
R5250 gnd.n4922 gnd.n1277 240.244
R5251 gnd.n4914 gnd.n1277 240.244
R5252 gnd.n4914 gnd.n1293 240.244
R5253 gnd.n4910 gnd.n1293 240.244
R5254 gnd.n4910 gnd.n1299 240.244
R5255 gnd.n4902 gnd.n1299 240.244
R5256 gnd.n4902 gnd.n1314 240.244
R5257 gnd.n4898 gnd.n1314 240.244
R5258 gnd.n6488 gnd.n965 240.244
R5259 gnd.n6485 gnd.n5143 240.244
R5260 gnd.n6481 gnd.n6480 240.244
R5261 gnd.n6477 gnd.n6476 240.244
R5262 gnd.n6473 gnd.n6472 240.244
R5263 gnd.n6469 gnd.n6468 240.244
R5264 gnd.n6465 gnd.n6464 240.244
R5265 gnd.n6461 gnd.n6460 240.244
R5266 gnd.n5750 gnd.n5470 240.244
R5267 gnd.n5470 gnd.n5461 240.244
R5268 gnd.n5768 gnd.n5461 240.244
R5269 gnd.n5769 gnd.n5768 240.244
R5270 gnd.n5769 gnd.n5449 240.244
R5271 gnd.n5449 gnd.n5438 240.244
R5272 gnd.n5800 gnd.n5438 240.244
R5273 gnd.n5801 gnd.n5800 240.244
R5274 gnd.n5802 gnd.n5801 240.244
R5275 gnd.n5802 gnd.n5423 240.244
R5276 gnd.n5804 gnd.n5423 240.244
R5277 gnd.n5804 gnd.n5408 240.244
R5278 gnd.n5845 gnd.n5408 240.244
R5279 gnd.n5846 gnd.n5845 240.244
R5280 gnd.n5849 gnd.n5846 240.244
R5281 gnd.n5849 gnd.n5390 240.244
R5282 gnd.n5881 gnd.n5390 240.244
R5283 gnd.n5881 gnd.n5376 240.244
R5284 gnd.n5903 gnd.n5376 240.244
R5285 gnd.n5904 gnd.n5903 240.244
R5286 gnd.n5904 gnd.n5363 240.244
R5287 gnd.n5363 gnd.n5352 240.244
R5288 gnd.n5935 gnd.n5352 240.244
R5289 gnd.n5936 gnd.n5935 240.244
R5290 gnd.n5937 gnd.n5936 240.244
R5291 gnd.n5937 gnd.n5289 240.244
R5292 gnd.n5289 gnd.n5288 240.244
R5293 gnd.n5288 gnd.n5273 240.244
R5294 gnd.n5988 gnd.n5273 240.244
R5295 gnd.n5989 gnd.n5988 240.244
R5296 gnd.n5989 gnd.n5260 240.244
R5297 gnd.n5260 gnd.n5249 240.244
R5298 gnd.n6022 gnd.n5249 240.244
R5299 gnd.n6023 gnd.n6022 240.244
R5300 gnd.n6025 gnd.n6023 240.244
R5301 gnd.n6025 gnd.n6024 240.244
R5302 gnd.n6024 gnd.n5228 240.244
R5303 gnd.n6060 gnd.n5228 240.244
R5304 gnd.n6060 gnd.n5220 240.244
R5305 gnd.n5220 gnd.n5213 240.244
R5306 gnd.n6085 gnd.n5213 240.244
R5307 gnd.n6085 gnd.n908 240.244
R5308 gnd.n6098 gnd.n908 240.244
R5309 gnd.n6098 gnd.n918 240.244
R5310 gnd.n5201 gnd.n918 240.244
R5311 gnd.n6118 gnd.n5201 240.244
R5312 gnd.n6118 gnd.n930 240.244
R5313 gnd.n5196 gnd.n930 240.244
R5314 gnd.n5196 gnd.n943 240.244
R5315 gnd.n5194 gnd.n943 240.244
R5316 gnd.n6393 gnd.n5194 240.244
R5317 gnd.n6393 gnd.n955 240.244
R5318 gnd.n6389 gnd.n955 240.244
R5319 gnd.n5687 gnd.n5686 240.244
R5320 gnd.n5731 gnd.n5686 240.244
R5321 gnd.n5729 gnd.n5728 240.244
R5322 gnd.n5725 gnd.n5724 240.244
R5323 gnd.n5721 gnd.n5720 240.244
R5324 gnd.n5717 gnd.n5716 240.244
R5325 gnd.n5713 gnd.n5712 240.244
R5326 gnd.n5709 gnd.n5708 240.244
R5327 gnd.n5760 gnd.n5468 240.244
R5328 gnd.n5760 gnd.n5464 240.244
R5329 gnd.n5766 gnd.n5464 240.244
R5330 gnd.n5766 gnd.n5447 240.244
R5331 gnd.n5790 gnd.n5447 240.244
R5332 gnd.n5790 gnd.n5442 240.244
R5333 gnd.n5798 gnd.n5442 240.244
R5334 gnd.n5798 gnd.n5443 240.244
R5335 gnd.n5443 gnd.n5421 240.244
R5336 gnd.n5824 gnd.n5421 240.244
R5337 gnd.n5824 gnd.n5416 240.244
R5338 gnd.n5835 gnd.n5416 240.244
R5339 gnd.n5835 gnd.n5417 240.244
R5340 gnd.n5831 gnd.n5417 240.244
R5341 gnd.n5831 gnd.n5388 240.244
R5342 gnd.n5885 gnd.n5388 240.244
R5343 gnd.n5885 gnd.n5383 240.244
R5344 gnd.n5893 gnd.n5383 240.244
R5345 gnd.n5893 gnd.n5384 240.244
R5346 gnd.n5384 gnd.n5361 240.244
R5347 gnd.n5925 gnd.n5361 240.244
R5348 gnd.n5925 gnd.n5356 240.244
R5349 gnd.n5933 gnd.n5356 240.244
R5350 gnd.n5933 gnd.n5357 240.244
R5351 gnd.n5357 gnd.n5286 240.244
R5352 gnd.n5970 gnd.n5286 240.244
R5353 gnd.n5970 gnd.n5281 240.244
R5354 gnd.n5978 gnd.n5281 240.244
R5355 gnd.n5978 gnd.n5282 240.244
R5356 gnd.n5282 gnd.n5258 240.244
R5357 gnd.n6009 gnd.n5258 240.244
R5358 gnd.n6009 gnd.n5253 240.244
R5359 gnd.n6020 gnd.n5253 240.244
R5360 gnd.n6020 gnd.n5254 240.244
R5361 gnd.n6016 gnd.n5254 240.244
R5362 gnd.n6016 gnd.n5227 240.244
R5363 gnd.n6064 gnd.n5227 240.244
R5364 gnd.n6064 gnd.n5222 240.244
R5365 gnd.n6073 gnd.n5222 240.244
R5366 gnd.n6073 gnd.n5223 240.244
R5367 gnd.n5223 gnd.n910 240.244
R5368 gnd.n6522 gnd.n910 240.244
R5369 gnd.n6522 gnd.n911 240.244
R5370 gnd.n6518 gnd.n911 240.244
R5371 gnd.n6518 gnd.n917 240.244
R5372 gnd.n932 gnd.n917 240.244
R5373 gnd.n6508 gnd.n932 240.244
R5374 gnd.n6508 gnd.n933 240.244
R5375 gnd.n6504 gnd.n933 240.244
R5376 gnd.n6504 gnd.n941 240.244
R5377 gnd.n957 gnd.n941 240.244
R5378 gnd.n6494 gnd.n957 240.244
R5379 gnd.n6494 gnd.n958 240.244
R5380 gnd.n5162 gnd.n967 240.244
R5381 gnd.n6451 gnd.n6450 240.244
R5382 gnd.n6447 gnd.n6446 240.244
R5383 gnd.n6443 gnd.n6442 240.244
R5384 gnd.n6439 gnd.n6438 240.244
R5385 gnd.n6435 gnd.n6434 240.244
R5386 gnd.n6431 gnd.n6430 240.244
R5387 gnd.n6427 gnd.n6426 240.244
R5388 gnd.n6423 gnd.n6422 240.244
R5389 gnd.n6419 gnd.n6418 240.244
R5390 gnd.n6415 gnd.n6414 240.244
R5391 gnd.n6411 gnd.n6410 240.244
R5392 gnd.n6407 gnd.n6406 240.244
R5393 gnd.n5618 gnd.n5514 240.244
R5394 gnd.n5624 gnd.n5514 240.244
R5395 gnd.n5624 gnd.n5506 240.244
R5396 gnd.n5634 gnd.n5506 240.244
R5397 gnd.n5634 gnd.n5502 240.244
R5398 gnd.n5640 gnd.n5502 240.244
R5399 gnd.n5640 gnd.n5493 240.244
R5400 gnd.n5650 gnd.n5493 240.244
R5401 gnd.n5650 gnd.n5488 240.244
R5402 gnd.n5678 gnd.n5488 240.244
R5403 gnd.n5678 gnd.n5489 240.244
R5404 gnd.n5489 gnd.n5481 240.244
R5405 gnd.n5673 gnd.n5481 240.244
R5406 gnd.n5673 gnd.n5471 240.244
R5407 gnd.n5670 gnd.n5471 240.244
R5408 gnd.n5670 gnd.n5460 240.244
R5409 gnd.n5667 gnd.n5460 240.244
R5410 gnd.n5667 gnd.n5450 240.244
R5411 gnd.n5664 gnd.n5450 240.244
R5412 gnd.n5664 gnd.n5428 240.244
R5413 gnd.n5813 gnd.n5428 240.244
R5414 gnd.n5813 gnd.n5424 240.244
R5415 gnd.n5821 gnd.n5424 240.244
R5416 gnd.n5821 gnd.n5414 240.244
R5417 gnd.n5414 gnd.n5395 240.244
R5418 gnd.n5860 gnd.n5395 240.244
R5419 gnd.n5860 gnd.n5396 240.244
R5420 gnd.n5396 gnd.n5391 240.244
R5421 gnd.n5880 gnd.n5391 240.244
R5422 gnd.n5880 gnd.n5381 240.244
R5423 gnd.n5875 gnd.n5381 240.244
R5424 gnd.n5875 gnd.n5375 240.244
R5425 gnd.n5871 gnd.n5375 240.244
R5426 gnd.n5871 gnd.n5364 240.244
R5427 gnd.n5867 gnd.n5364 240.244
R5428 gnd.n5867 gnd.n5342 240.244
R5429 gnd.n5946 gnd.n5342 240.244
R5430 gnd.n5946 gnd.n5290 240.244
R5431 gnd.n5967 gnd.n5290 240.244
R5432 gnd.n5967 gnd.n5279 240.244
R5433 gnd.n5963 gnd.n5279 240.244
R5434 gnd.n5963 gnd.n5272 240.244
R5435 gnd.n5960 gnd.n5272 240.244
R5436 gnd.n5960 gnd.n5261 240.244
R5437 gnd.n5957 gnd.n5261 240.244
R5438 gnd.n5957 gnd.n5239 240.244
R5439 gnd.n6032 gnd.n5239 240.244
R5440 gnd.n6032 gnd.n5235 240.244
R5441 gnd.n6050 gnd.n5235 240.244
R5442 gnd.n6050 gnd.n5229 240.244
R5443 gnd.n5229 gnd.n5219 240.244
R5444 gnd.n6045 gnd.n5219 240.244
R5445 gnd.n6045 gnd.n5212 240.244
R5446 gnd.n6042 gnd.n5212 240.244
R5447 gnd.n6042 gnd.n5205 240.244
R5448 gnd.n6101 gnd.n5205 240.244
R5449 gnd.n6101 gnd.n919 240.244
R5450 gnd.n6115 gnd.n919 240.244
R5451 gnd.n6115 gnd.n929 240.244
R5452 gnd.n6111 gnd.n929 240.244
R5453 gnd.n6111 gnd.n6110 240.244
R5454 gnd.n6110 gnd.n944 240.244
R5455 gnd.n6396 gnd.n944 240.244
R5456 gnd.n6396 gnd.n954 240.244
R5457 gnd.n6402 gnd.n954 240.244
R5458 gnd.n5610 gnd.n5608 240.244
R5459 gnd.n5608 gnd.n5607 240.244
R5460 gnd.n5604 gnd.n5603 240.244
R5461 gnd.n5601 gnd.n5527 240.244
R5462 gnd.n5597 gnd.n5595 240.244
R5463 gnd.n5593 gnd.n5533 240.244
R5464 gnd.n5589 gnd.n5587 240.244
R5465 gnd.n5585 gnd.n5539 240.244
R5466 gnd.n5581 gnd.n5579 240.244
R5467 gnd.n5577 gnd.n5545 240.244
R5468 gnd.n5573 gnd.n5571 240.244
R5469 gnd.n5569 gnd.n5551 240.244
R5470 gnd.n5564 gnd.n5562 240.244
R5471 gnd.n5616 gnd.n5512 240.244
R5472 gnd.n5626 gnd.n5512 240.244
R5473 gnd.n5626 gnd.n5508 240.244
R5474 gnd.n5632 gnd.n5508 240.244
R5475 gnd.n5632 gnd.n5500 240.244
R5476 gnd.n5642 gnd.n5500 240.244
R5477 gnd.n5642 gnd.n5496 240.244
R5478 gnd.n5648 gnd.n5496 240.244
R5479 gnd.n5648 gnd.n5487 240.244
R5480 gnd.n5740 gnd.n5487 240.244
R5481 gnd.n5740 gnd.n5482 240.244
R5482 gnd.n5747 gnd.n5482 240.244
R5483 gnd.n5747 gnd.n5473 240.244
R5484 gnd.n5757 gnd.n5473 240.244
R5485 gnd.n5757 gnd.n5459 240.244
R5486 gnd.n5772 gnd.n5459 240.244
R5487 gnd.n5772 gnd.n5452 240.244
R5488 gnd.n5787 gnd.n5452 240.244
R5489 gnd.n5787 gnd.n5453 240.244
R5490 gnd.n5453 gnd.n5431 240.244
R5491 gnd.n5811 gnd.n5431 240.244
R5492 gnd.n5811 gnd.n5432 240.244
R5493 gnd.n5432 gnd.n5412 240.244
R5494 gnd.n5838 gnd.n5412 240.244
R5495 gnd.n5838 gnd.n5399 240.244
R5496 gnd.n5858 gnd.n5399 240.244
R5497 gnd.n5858 gnd.n5400 240.244
R5498 gnd.n5854 gnd.n5400 240.244
R5499 gnd.n5854 gnd.n5380 240.244
R5500 gnd.n5896 gnd.n5380 240.244
R5501 gnd.n5896 gnd.n5373 240.244
R5502 gnd.n5907 gnd.n5373 240.244
R5503 gnd.n5907 gnd.n5366 240.244
R5504 gnd.n5922 gnd.n5366 240.244
R5505 gnd.n5922 gnd.n5367 240.244
R5506 gnd.n5367 gnd.n5345 240.244
R5507 gnd.n5944 gnd.n5345 240.244
R5508 gnd.n5944 gnd.n5346 240.244
R5509 gnd.n5346 gnd.n5277 240.244
R5510 gnd.n5981 gnd.n5277 240.244
R5511 gnd.n5981 gnd.n5270 240.244
R5512 gnd.n5992 gnd.n5270 240.244
R5513 gnd.n5992 gnd.n5263 240.244
R5514 gnd.n6006 gnd.n5263 240.244
R5515 gnd.n6006 gnd.n5264 240.244
R5516 gnd.n5264 gnd.n5243 240.244
R5517 gnd.n6030 gnd.n5243 240.244
R5518 gnd.n6030 gnd.n5233 240.244
R5519 gnd.n6052 gnd.n5233 240.244
R5520 gnd.n6052 gnd.n5218 240.244
R5521 gnd.n6076 gnd.n5218 240.244
R5522 gnd.n6076 gnd.n5209 240.244
R5523 gnd.n6088 gnd.n5209 240.244
R5524 gnd.n6089 gnd.n6088 240.244
R5525 gnd.n6090 gnd.n6089 240.244
R5526 gnd.n6090 gnd.n921 240.244
R5527 gnd.n6515 gnd.n921 240.244
R5528 gnd.n6515 gnd.n922 240.244
R5529 gnd.n6511 gnd.n922 240.244
R5530 gnd.n6511 gnd.n928 240.244
R5531 gnd.n946 gnd.n928 240.244
R5532 gnd.n6501 gnd.n946 240.244
R5533 gnd.n6501 gnd.n947 240.244
R5534 gnd.n6497 gnd.n947 240.244
R5535 gnd.n6497 gnd.n953 240.244
R5536 gnd.n7578 gnd.n7577 240.244
R5537 gnd.n7583 gnd.n7580 240.244
R5538 gnd.n7586 gnd.n7585 240.244
R5539 gnd.n7591 gnd.n7588 240.244
R5540 gnd.n7594 gnd.n7593 240.244
R5541 gnd.n7599 gnd.n7596 240.244
R5542 gnd.n7602 gnd.n7601 240.244
R5543 gnd.n7607 gnd.n7604 240.244
R5544 gnd.n7613 gnd.n7609 240.244
R5545 gnd.n4476 gnd.n1479 240.244
R5546 gnd.n4483 gnd.n1479 240.244
R5547 gnd.n4483 gnd.n1492 240.244
R5548 gnd.n1623 gnd.n1492 240.244
R5549 gnd.n4526 gnd.n1623 240.244
R5550 gnd.n4526 gnd.n1618 240.244
R5551 gnd.n4533 gnd.n1618 240.244
R5552 gnd.n4533 gnd.n1607 240.244
R5553 gnd.n1607 gnd.n1596 240.244
R5554 gnd.n4558 gnd.n1596 240.244
R5555 gnd.n4558 gnd.n1591 240.244
R5556 gnd.n4565 gnd.n1591 240.244
R5557 gnd.n4565 gnd.n1580 240.244
R5558 gnd.n1580 gnd.n1567 240.244
R5559 gnd.n4597 gnd.n1567 240.244
R5560 gnd.n4597 gnd.n1562 240.244
R5561 gnd.n4607 gnd.n1562 240.244
R5562 gnd.n4607 gnd.n1527 240.244
R5563 gnd.n4601 gnd.n1527 240.244
R5564 gnd.n4601 gnd.n1519 240.244
R5565 gnd.n4623 gnd.n1519 240.244
R5566 gnd.n4623 gnd.n279 240.244
R5567 gnd.n4632 gnd.n279 240.244
R5568 gnd.n4632 gnd.n1551 240.244
R5569 gnd.n1551 gnd.n1543 240.244
R5570 gnd.n4643 gnd.n1543 240.244
R5571 gnd.n4643 gnd.n70 240.244
R5572 gnd.n71 gnd.n70 240.244
R5573 gnd.n72 gnd.n71 240.244
R5574 gnd.n305 gnd.n72 240.244
R5575 gnd.n305 gnd.n75 240.244
R5576 gnd.n76 gnd.n75 240.244
R5577 gnd.n77 gnd.n76 240.244
R5578 gnd.n7409 gnd.n77 240.244
R5579 gnd.n7409 gnd.n80 240.244
R5580 gnd.n81 gnd.n80 240.244
R5581 gnd.n82 gnd.n81 240.244
R5582 gnd.n7453 gnd.n82 240.244
R5583 gnd.n7453 gnd.n85 240.244
R5584 gnd.n86 gnd.n85 240.244
R5585 gnd.n87 gnd.n86 240.244
R5586 gnd.n217 gnd.n87 240.244
R5587 gnd.n217 gnd.n90 240.244
R5588 gnd.n91 gnd.n90 240.244
R5589 gnd.n92 gnd.n91 240.244
R5590 gnd.n210 gnd.n92 240.244
R5591 gnd.n210 gnd.n95 240.244
R5592 gnd.n96 gnd.n95 240.244
R5593 gnd.n97 gnd.n96 240.244
R5594 gnd.n185 gnd.n97 240.244
R5595 gnd.n185 gnd.n100 240.244
R5596 gnd.n101 gnd.n100 240.244
R5597 gnd.n7741 gnd.n101 240.244
R5598 gnd.n1705 gnd.n1682 240.244
R5599 gnd.n1709 gnd.n1707 240.244
R5600 gnd.n1724 gnd.n1673 240.244
R5601 gnd.n1728 gnd.n1726 240.244
R5602 gnd.n1743 gnd.n1664 240.244
R5603 gnd.n1747 gnd.n1745 240.244
R5604 gnd.n1762 gnd.n1655 240.244
R5605 gnd.n1766 gnd.n1764 240.244
R5606 gnd.n4475 gnd.n1644 240.244
R5607 gnd.n1688 gnd.n1481 240.244
R5608 gnd.n1494 gnd.n1481 240.244
R5609 gnd.n4714 gnd.n1494 240.244
R5610 gnd.n4714 gnd.n1495 240.244
R5611 gnd.n1500 gnd.n1495 240.244
R5612 gnd.n1501 gnd.n1500 240.244
R5613 gnd.n1502 gnd.n1501 240.244
R5614 gnd.n4546 gnd.n1502 240.244
R5615 gnd.n4546 gnd.n1505 240.244
R5616 gnd.n1506 gnd.n1505 240.244
R5617 gnd.n1507 gnd.n1506 240.244
R5618 gnd.n4566 gnd.n1507 240.244
R5619 gnd.n4566 gnd.n1510 240.244
R5620 gnd.n1511 gnd.n1510 240.244
R5621 gnd.n1512 gnd.n1511 240.244
R5622 gnd.n1571 gnd.n1512 240.244
R5623 gnd.n1571 gnd.n1515 240.244
R5624 gnd.n1516 gnd.n1515 240.244
R5625 gnd.n1517 gnd.n1516 240.244
R5626 gnd.n4685 gnd.n1517 240.244
R5627 gnd.n4685 gnd.n281 240.244
R5628 gnd.n7497 gnd.n281 240.244
R5629 gnd.n7497 gnd.n282 240.244
R5630 gnd.n287 gnd.n282 240.244
R5631 gnd.n288 gnd.n287 240.244
R5632 gnd.n289 gnd.n288 240.244
R5633 gnd.n4644 gnd.n289 240.244
R5634 gnd.n4644 gnd.n293 240.244
R5635 gnd.n7483 gnd.n293 240.244
R5636 gnd.n7483 gnd.n262 240.244
R5637 gnd.n7506 gnd.n262 240.244
R5638 gnd.n7506 gnd.n258 240.244
R5639 gnd.n7512 gnd.n258 240.244
R5640 gnd.n7512 gnd.n246 240.244
R5641 gnd.n7522 gnd.n246 240.244
R5642 gnd.n7522 gnd.n242 240.244
R5643 gnd.n7528 gnd.n242 240.244
R5644 gnd.n7528 gnd.n231 240.244
R5645 gnd.n7538 gnd.n231 240.244
R5646 gnd.n7538 gnd.n227 240.244
R5647 gnd.n7544 gnd.n227 240.244
R5648 gnd.n7544 gnd.n216 240.244
R5649 gnd.n7554 gnd.n216 240.244
R5650 gnd.n7554 gnd.n212 240.244
R5651 gnd.n7560 gnd.n212 240.244
R5652 gnd.n7560 gnd.n201 240.244
R5653 gnd.n7570 gnd.n201 240.244
R5654 gnd.n7570 gnd.n195 240.244
R5655 gnd.n7651 gnd.n195 240.244
R5656 gnd.n7651 gnd.n196 240.244
R5657 gnd.n196 gnd.n187 240.244
R5658 gnd.n7575 gnd.n187 240.244
R5659 gnd.n7575 gnd.n107 240.244
R5660 gnd.n3288 gnd.n1324 240.244
R5661 gnd.n3291 gnd.n3290 240.244
R5662 gnd.n3301 gnd.n3293 240.244
R5663 gnd.n3304 gnd.n3303 240.244
R5664 gnd.n3313 gnd.n3312 240.244
R5665 gnd.n3324 gnd.n3315 240.244
R5666 gnd.n3327 gnd.n3326 240.244
R5667 gnd.n3336 gnd.n3335 240.244
R5668 gnd.n3347 gnd.n3338 240.244
R5669 gnd.n3039 gnd.n2958 240.244
R5670 gnd.n3040 gnd.n3039 240.244
R5671 gnd.n3040 gnd.n1064 240.244
R5672 gnd.n3043 gnd.n1064 240.244
R5673 gnd.n3043 gnd.n1076 240.244
R5674 gnd.n3048 gnd.n1076 240.244
R5675 gnd.n3048 gnd.n1087 240.244
R5676 gnd.n3051 gnd.n1087 240.244
R5677 gnd.n3051 gnd.n1097 240.244
R5678 gnd.n3056 gnd.n1097 240.244
R5679 gnd.n3056 gnd.n1107 240.244
R5680 gnd.n3080 gnd.n1107 240.244
R5681 gnd.n3080 gnd.n1118 240.244
R5682 gnd.n3086 gnd.n1118 240.244
R5683 gnd.n3086 gnd.n1129 240.244
R5684 gnd.n3096 gnd.n1129 240.244
R5685 gnd.n3096 gnd.n1140 240.244
R5686 gnd.n3102 gnd.n1140 240.244
R5687 gnd.n3102 gnd.n1150 240.244
R5688 gnd.n3112 gnd.n1150 240.244
R5689 gnd.n3112 gnd.n1160 240.244
R5690 gnd.n3118 gnd.n1160 240.244
R5691 gnd.n3118 gnd.n1171 240.244
R5692 gnd.n3128 gnd.n1171 240.244
R5693 gnd.n3128 gnd.n1180 240.244
R5694 gnd.n3135 gnd.n1180 240.244
R5695 gnd.n3135 gnd.n1190 240.244
R5696 gnd.n3146 gnd.n1190 240.244
R5697 gnd.n3146 gnd.n1197 240.244
R5698 gnd.n3152 gnd.n1197 240.244
R5699 gnd.n3152 gnd.n1208 240.244
R5700 gnd.n3162 gnd.n1208 240.244
R5701 gnd.n3162 gnd.n1218 240.244
R5702 gnd.n3168 gnd.n1218 240.244
R5703 gnd.n3168 gnd.n1228 240.244
R5704 gnd.n3178 gnd.n1228 240.244
R5705 gnd.n3178 gnd.n1238 240.244
R5706 gnd.n3184 gnd.n1238 240.244
R5707 gnd.n3184 gnd.n1249 240.244
R5708 gnd.n3195 gnd.n1249 240.244
R5709 gnd.n3195 gnd.n1260 240.244
R5710 gnd.n3201 gnd.n1260 240.244
R5711 gnd.n3201 gnd.n1270 240.244
R5712 gnd.n3236 gnd.n1270 240.244
R5713 gnd.n3236 gnd.n1280 240.244
R5714 gnd.n2799 gnd.n1280 240.244
R5715 gnd.n2799 gnd.n1291 240.244
R5716 gnd.n2800 gnd.n1291 240.244
R5717 gnd.n2800 gnd.n1302 240.244
R5718 gnd.n3224 gnd.n1302 240.244
R5719 gnd.n3224 gnd.n1313 240.244
R5720 gnd.n3527 gnd.n1313 240.244
R5721 gnd.n3527 gnd.n1322 240.244
R5722 gnd.n3019 gnd.n3018 240.244
R5723 gnd.n3015 gnd.n3014 240.244
R5724 gnd.n3011 gnd.n3010 240.244
R5725 gnd.n3007 gnd.n3006 240.244
R5726 gnd.n3003 gnd.n3002 240.244
R5727 gnd.n2999 gnd.n2998 240.244
R5728 gnd.n2995 gnd.n2994 240.244
R5729 gnd.n2991 gnd.n2990 240.244
R5730 gnd.n2978 gnd.n1008 240.244
R5731 gnd.n3031 gnd.n2959 240.244
R5732 gnd.n3031 gnd.n2960 240.244
R5733 gnd.n2960 gnd.n1066 240.244
R5734 gnd.n1078 gnd.n1066 240.244
R5735 gnd.n5041 gnd.n1078 240.244
R5736 gnd.n5041 gnd.n1079 240.244
R5737 gnd.n5037 gnd.n1079 240.244
R5738 gnd.n5037 gnd.n1085 240.244
R5739 gnd.n5029 gnd.n1085 240.244
R5740 gnd.n5029 gnd.n1098 240.244
R5741 gnd.n5025 gnd.n1098 240.244
R5742 gnd.n5025 gnd.n1104 240.244
R5743 gnd.n5017 gnd.n1104 240.244
R5744 gnd.n5017 gnd.n1120 240.244
R5745 gnd.n5013 gnd.n1120 240.244
R5746 gnd.n5013 gnd.n1126 240.244
R5747 gnd.n5005 gnd.n1126 240.244
R5748 gnd.n5005 gnd.n1141 240.244
R5749 gnd.n5001 gnd.n1141 240.244
R5750 gnd.n5001 gnd.n1147 240.244
R5751 gnd.n4993 gnd.n1147 240.244
R5752 gnd.n4993 gnd.n1162 240.244
R5753 gnd.n4989 gnd.n1162 240.244
R5754 gnd.n4989 gnd.n1168 240.244
R5755 gnd.n4981 gnd.n1168 240.244
R5756 gnd.n4981 gnd.n1181 240.244
R5757 gnd.n4977 gnd.n1181 240.244
R5758 gnd.n4977 gnd.n1187 240.244
R5759 gnd.n4968 gnd.n1187 240.244
R5760 gnd.n4968 gnd.n1199 240.244
R5761 gnd.n4964 gnd.n1199 240.244
R5762 gnd.n4964 gnd.n1205 240.244
R5763 gnd.n4956 gnd.n1205 240.244
R5764 gnd.n4956 gnd.n1219 240.244
R5765 gnd.n4952 gnd.n1219 240.244
R5766 gnd.n4952 gnd.n1225 240.244
R5767 gnd.n4944 gnd.n1225 240.244
R5768 gnd.n4944 gnd.n1240 240.244
R5769 gnd.n4940 gnd.n1240 240.244
R5770 gnd.n4940 gnd.n1246 240.244
R5771 gnd.n4932 gnd.n1246 240.244
R5772 gnd.n4932 gnd.n1261 240.244
R5773 gnd.n4928 gnd.n1261 240.244
R5774 gnd.n4928 gnd.n1267 240.244
R5775 gnd.n4920 gnd.n1267 240.244
R5776 gnd.n4920 gnd.n1282 240.244
R5777 gnd.n4916 gnd.n1282 240.244
R5778 gnd.n4916 gnd.n1288 240.244
R5779 gnd.n4908 gnd.n1288 240.244
R5780 gnd.n4908 gnd.n1304 240.244
R5781 gnd.n4904 gnd.n1304 240.244
R5782 gnd.n4904 gnd.n1310 240.244
R5783 gnd.n4896 gnd.n1310 240.244
R5784 gnd.n6695 gnd.n739 240.244
R5785 gnd.n6695 gnd.n735 240.244
R5786 gnd.n6701 gnd.n735 240.244
R5787 gnd.n6701 gnd.n733 240.244
R5788 gnd.n6705 gnd.n733 240.244
R5789 gnd.n6705 gnd.n729 240.244
R5790 gnd.n6711 gnd.n729 240.244
R5791 gnd.n6711 gnd.n727 240.244
R5792 gnd.n6715 gnd.n727 240.244
R5793 gnd.n6715 gnd.n723 240.244
R5794 gnd.n6721 gnd.n723 240.244
R5795 gnd.n6721 gnd.n721 240.244
R5796 gnd.n6725 gnd.n721 240.244
R5797 gnd.n6725 gnd.n717 240.244
R5798 gnd.n6731 gnd.n717 240.244
R5799 gnd.n6731 gnd.n715 240.244
R5800 gnd.n6735 gnd.n715 240.244
R5801 gnd.n6735 gnd.n711 240.244
R5802 gnd.n6741 gnd.n711 240.244
R5803 gnd.n6741 gnd.n709 240.244
R5804 gnd.n6745 gnd.n709 240.244
R5805 gnd.n6745 gnd.n705 240.244
R5806 gnd.n6751 gnd.n705 240.244
R5807 gnd.n6751 gnd.n703 240.244
R5808 gnd.n6755 gnd.n703 240.244
R5809 gnd.n6755 gnd.n699 240.244
R5810 gnd.n6761 gnd.n699 240.244
R5811 gnd.n6761 gnd.n697 240.244
R5812 gnd.n6765 gnd.n697 240.244
R5813 gnd.n6765 gnd.n693 240.244
R5814 gnd.n6771 gnd.n693 240.244
R5815 gnd.n6771 gnd.n691 240.244
R5816 gnd.n6775 gnd.n691 240.244
R5817 gnd.n6775 gnd.n687 240.244
R5818 gnd.n6781 gnd.n687 240.244
R5819 gnd.n6781 gnd.n685 240.244
R5820 gnd.n6785 gnd.n685 240.244
R5821 gnd.n6785 gnd.n681 240.244
R5822 gnd.n6791 gnd.n681 240.244
R5823 gnd.n6791 gnd.n679 240.244
R5824 gnd.n6795 gnd.n679 240.244
R5825 gnd.n6795 gnd.n675 240.244
R5826 gnd.n6801 gnd.n675 240.244
R5827 gnd.n6801 gnd.n673 240.244
R5828 gnd.n6805 gnd.n673 240.244
R5829 gnd.n6805 gnd.n669 240.244
R5830 gnd.n6811 gnd.n669 240.244
R5831 gnd.n6811 gnd.n667 240.244
R5832 gnd.n6815 gnd.n667 240.244
R5833 gnd.n6815 gnd.n663 240.244
R5834 gnd.n6821 gnd.n663 240.244
R5835 gnd.n6821 gnd.n661 240.244
R5836 gnd.n6825 gnd.n661 240.244
R5837 gnd.n6825 gnd.n657 240.244
R5838 gnd.n6831 gnd.n657 240.244
R5839 gnd.n6831 gnd.n655 240.244
R5840 gnd.n6835 gnd.n655 240.244
R5841 gnd.n6835 gnd.n651 240.244
R5842 gnd.n6841 gnd.n651 240.244
R5843 gnd.n6841 gnd.n649 240.244
R5844 gnd.n6845 gnd.n649 240.244
R5845 gnd.n6845 gnd.n645 240.244
R5846 gnd.n6851 gnd.n645 240.244
R5847 gnd.n6851 gnd.n643 240.244
R5848 gnd.n6855 gnd.n643 240.244
R5849 gnd.n6855 gnd.n639 240.244
R5850 gnd.n6861 gnd.n639 240.244
R5851 gnd.n6861 gnd.n637 240.244
R5852 gnd.n6865 gnd.n637 240.244
R5853 gnd.n6865 gnd.n633 240.244
R5854 gnd.n6871 gnd.n633 240.244
R5855 gnd.n6871 gnd.n631 240.244
R5856 gnd.n6875 gnd.n631 240.244
R5857 gnd.n6875 gnd.n627 240.244
R5858 gnd.n6881 gnd.n627 240.244
R5859 gnd.n6881 gnd.n625 240.244
R5860 gnd.n6885 gnd.n625 240.244
R5861 gnd.n6885 gnd.n621 240.244
R5862 gnd.n6891 gnd.n621 240.244
R5863 gnd.n6891 gnd.n619 240.244
R5864 gnd.n6895 gnd.n619 240.244
R5865 gnd.n6895 gnd.n615 240.244
R5866 gnd.n6901 gnd.n615 240.244
R5867 gnd.n6901 gnd.n613 240.244
R5868 gnd.n6905 gnd.n613 240.244
R5869 gnd.n6905 gnd.n609 240.244
R5870 gnd.n6911 gnd.n609 240.244
R5871 gnd.n6911 gnd.n607 240.244
R5872 gnd.n6915 gnd.n607 240.244
R5873 gnd.n6915 gnd.n603 240.244
R5874 gnd.n6921 gnd.n603 240.244
R5875 gnd.n6921 gnd.n601 240.244
R5876 gnd.n6925 gnd.n601 240.244
R5877 gnd.n6925 gnd.n597 240.244
R5878 gnd.n6931 gnd.n597 240.244
R5879 gnd.n6931 gnd.n595 240.244
R5880 gnd.n6935 gnd.n595 240.244
R5881 gnd.n6935 gnd.n591 240.244
R5882 gnd.n6941 gnd.n591 240.244
R5883 gnd.n6941 gnd.n589 240.244
R5884 gnd.n6945 gnd.n589 240.244
R5885 gnd.n6945 gnd.n585 240.244
R5886 gnd.n6951 gnd.n585 240.244
R5887 gnd.n6951 gnd.n583 240.244
R5888 gnd.n6955 gnd.n583 240.244
R5889 gnd.n6955 gnd.n579 240.244
R5890 gnd.n6961 gnd.n579 240.244
R5891 gnd.n6961 gnd.n577 240.244
R5892 gnd.n6965 gnd.n577 240.244
R5893 gnd.n6965 gnd.n573 240.244
R5894 gnd.n6971 gnd.n573 240.244
R5895 gnd.n6971 gnd.n571 240.244
R5896 gnd.n6975 gnd.n571 240.244
R5897 gnd.n6975 gnd.n567 240.244
R5898 gnd.n6981 gnd.n567 240.244
R5899 gnd.n6981 gnd.n565 240.244
R5900 gnd.n6985 gnd.n565 240.244
R5901 gnd.n6985 gnd.n561 240.244
R5902 gnd.n6991 gnd.n561 240.244
R5903 gnd.n6991 gnd.n559 240.244
R5904 gnd.n6995 gnd.n559 240.244
R5905 gnd.n6995 gnd.n555 240.244
R5906 gnd.n7001 gnd.n555 240.244
R5907 gnd.n7001 gnd.n553 240.244
R5908 gnd.n7005 gnd.n553 240.244
R5909 gnd.n7005 gnd.n549 240.244
R5910 gnd.n7011 gnd.n549 240.244
R5911 gnd.n7011 gnd.n547 240.244
R5912 gnd.n7015 gnd.n547 240.244
R5913 gnd.n7015 gnd.n543 240.244
R5914 gnd.n7021 gnd.n543 240.244
R5915 gnd.n7021 gnd.n541 240.244
R5916 gnd.n7025 gnd.n541 240.244
R5917 gnd.n7025 gnd.n537 240.244
R5918 gnd.n7031 gnd.n537 240.244
R5919 gnd.n7031 gnd.n535 240.244
R5920 gnd.n7035 gnd.n535 240.244
R5921 gnd.n7035 gnd.n531 240.244
R5922 gnd.n7041 gnd.n531 240.244
R5923 gnd.n7041 gnd.n529 240.244
R5924 gnd.n7045 gnd.n529 240.244
R5925 gnd.n7045 gnd.n525 240.244
R5926 gnd.n7051 gnd.n525 240.244
R5927 gnd.n7051 gnd.n523 240.244
R5928 gnd.n7055 gnd.n523 240.244
R5929 gnd.n7055 gnd.n519 240.244
R5930 gnd.n7061 gnd.n519 240.244
R5931 gnd.n7061 gnd.n517 240.244
R5932 gnd.n7065 gnd.n517 240.244
R5933 gnd.n7065 gnd.n513 240.244
R5934 gnd.n7071 gnd.n513 240.244
R5935 gnd.n7071 gnd.n511 240.244
R5936 gnd.n7075 gnd.n511 240.244
R5937 gnd.n7075 gnd.n507 240.244
R5938 gnd.n7081 gnd.n507 240.244
R5939 gnd.n7081 gnd.n505 240.244
R5940 gnd.n7085 gnd.n505 240.244
R5941 gnd.n7085 gnd.n501 240.244
R5942 gnd.n7091 gnd.n501 240.244
R5943 gnd.n7091 gnd.n499 240.244
R5944 gnd.n7095 gnd.n499 240.244
R5945 gnd.n7095 gnd.n495 240.244
R5946 gnd.n7101 gnd.n495 240.244
R5947 gnd.n7101 gnd.n493 240.244
R5948 gnd.n7105 gnd.n493 240.244
R5949 gnd.n7105 gnd.n489 240.244
R5950 gnd.n7111 gnd.n489 240.244
R5951 gnd.n7111 gnd.n487 240.244
R5952 gnd.n7115 gnd.n487 240.244
R5953 gnd.n7115 gnd.n483 240.244
R5954 gnd.n7121 gnd.n483 240.244
R5955 gnd.n7121 gnd.n481 240.244
R5956 gnd.n7125 gnd.n481 240.244
R5957 gnd.n7125 gnd.n477 240.244
R5958 gnd.n7131 gnd.n477 240.244
R5959 gnd.n7131 gnd.n475 240.244
R5960 gnd.n7135 gnd.n475 240.244
R5961 gnd.n7135 gnd.n471 240.244
R5962 gnd.n7141 gnd.n471 240.244
R5963 gnd.n7141 gnd.n469 240.244
R5964 gnd.n7145 gnd.n469 240.244
R5965 gnd.n7145 gnd.n465 240.244
R5966 gnd.n7151 gnd.n465 240.244
R5967 gnd.n7151 gnd.n463 240.244
R5968 gnd.n7155 gnd.n463 240.244
R5969 gnd.n7155 gnd.n459 240.244
R5970 gnd.n7161 gnd.n459 240.244
R5971 gnd.n7161 gnd.n457 240.244
R5972 gnd.n7165 gnd.n457 240.244
R5973 gnd.n7165 gnd.n453 240.244
R5974 gnd.n7172 gnd.n453 240.244
R5975 gnd.n7172 gnd.n451 240.244
R5976 gnd.n7176 gnd.n451 240.244
R5977 gnd.n7176 gnd.n448 240.244
R5978 gnd.n7182 gnd.n446 240.244
R5979 gnd.n7186 gnd.n446 240.244
R5980 gnd.n7186 gnd.n442 240.244
R5981 gnd.n7192 gnd.n442 240.244
R5982 gnd.n7192 gnd.n440 240.244
R5983 gnd.n7196 gnd.n440 240.244
R5984 gnd.n7196 gnd.n436 240.244
R5985 gnd.n7202 gnd.n436 240.244
R5986 gnd.n7202 gnd.n434 240.244
R5987 gnd.n7206 gnd.n434 240.244
R5988 gnd.n7206 gnd.n430 240.244
R5989 gnd.n7212 gnd.n430 240.244
R5990 gnd.n7212 gnd.n428 240.244
R5991 gnd.n7216 gnd.n428 240.244
R5992 gnd.n7216 gnd.n424 240.244
R5993 gnd.n7222 gnd.n424 240.244
R5994 gnd.n7222 gnd.n422 240.244
R5995 gnd.n7226 gnd.n422 240.244
R5996 gnd.n7226 gnd.n418 240.244
R5997 gnd.n7232 gnd.n418 240.244
R5998 gnd.n7232 gnd.n416 240.244
R5999 gnd.n7236 gnd.n416 240.244
R6000 gnd.n7236 gnd.n412 240.244
R6001 gnd.n7242 gnd.n412 240.244
R6002 gnd.n7242 gnd.n410 240.244
R6003 gnd.n7246 gnd.n410 240.244
R6004 gnd.n7246 gnd.n406 240.244
R6005 gnd.n7252 gnd.n406 240.244
R6006 gnd.n7252 gnd.n404 240.244
R6007 gnd.n7256 gnd.n404 240.244
R6008 gnd.n7256 gnd.n400 240.244
R6009 gnd.n7262 gnd.n400 240.244
R6010 gnd.n7262 gnd.n398 240.244
R6011 gnd.n7266 gnd.n398 240.244
R6012 gnd.n7266 gnd.n394 240.244
R6013 gnd.n7272 gnd.n394 240.244
R6014 gnd.n7272 gnd.n392 240.244
R6015 gnd.n7276 gnd.n392 240.244
R6016 gnd.n7276 gnd.n388 240.244
R6017 gnd.n7282 gnd.n388 240.244
R6018 gnd.n7282 gnd.n386 240.244
R6019 gnd.n7286 gnd.n386 240.244
R6020 gnd.n7286 gnd.n382 240.244
R6021 gnd.n7292 gnd.n382 240.244
R6022 gnd.n7292 gnd.n380 240.244
R6023 gnd.n7296 gnd.n380 240.244
R6024 gnd.n7296 gnd.n376 240.244
R6025 gnd.n7302 gnd.n376 240.244
R6026 gnd.n7302 gnd.n374 240.244
R6027 gnd.n7306 gnd.n374 240.244
R6028 gnd.n7306 gnd.n370 240.244
R6029 gnd.n7312 gnd.n370 240.244
R6030 gnd.n7312 gnd.n368 240.244
R6031 gnd.n7316 gnd.n368 240.244
R6032 gnd.n7316 gnd.n364 240.244
R6033 gnd.n7322 gnd.n364 240.244
R6034 gnd.n7322 gnd.n362 240.244
R6035 gnd.n7326 gnd.n362 240.244
R6036 gnd.n7326 gnd.n358 240.244
R6037 gnd.n7332 gnd.n358 240.244
R6038 gnd.n7332 gnd.n356 240.244
R6039 gnd.n7336 gnd.n356 240.244
R6040 gnd.n7336 gnd.n352 240.244
R6041 gnd.n7342 gnd.n352 240.244
R6042 gnd.n7342 gnd.n350 240.244
R6043 gnd.n7346 gnd.n350 240.244
R6044 gnd.n7346 gnd.n346 240.244
R6045 gnd.n7352 gnd.n346 240.244
R6046 gnd.n7352 gnd.n344 240.244
R6047 gnd.n7356 gnd.n344 240.244
R6048 gnd.n7356 gnd.n340 240.244
R6049 gnd.n7362 gnd.n340 240.244
R6050 gnd.n7362 gnd.n338 240.244
R6051 gnd.n7366 gnd.n338 240.244
R6052 gnd.n7366 gnd.n334 240.244
R6053 gnd.n7372 gnd.n334 240.244
R6054 gnd.n7372 gnd.n332 240.244
R6055 gnd.n7376 gnd.n332 240.244
R6056 gnd.n7376 gnd.n328 240.244
R6057 gnd.n7382 gnd.n328 240.244
R6058 gnd.n7382 gnd.n326 240.244
R6059 gnd.n7387 gnd.n326 240.244
R6060 gnd.n7387 gnd.n322 240.244
R6061 gnd.n7394 gnd.n322 240.244
R6062 gnd.n2865 gnd.n2856 240.244
R6063 gnd.n2866 gnd.n2865 240.244
R6064 gnd.n2867 gnd.n2866 240.244
R6065 gnd.n2867 gnd.n2851 240.244
R6066 gnd.n2942 gnd.n2851 240.244
R6067 gnd.n2942 gnd.n2852 240.244
R6068 gnd.n2938 gnd.n2852 240.244
R6069 gnd.n2938 gnd.n2937 240.244
R6070 gnd.n2937 gnd.n2936 240.244
R6071 gnd.n2936 gnd.n2875 240.244
R6072 gnd.n2929 gnd.n2875 240.244
R6073 gnd.n2929 gnd.n2928 240.244
R6074 gnd.n2928 gnd.n2927 240.244
R6075 gnd.n2927 gnd.n2925 240.244
R6076 gnd.n2925 gnd.n2922 240.244
R6077 gnd.n2922 gnd.n2921 240.244
R6078 gnd.n2921 gnd.n2918 240.244
R6079 gnd.n2918 gnd.n2917 240.244
R6080 gnd.n2917 gnd.n2882 240.244
R6081 gnd.n2913 gnd.n2882 240.244
R6082 gnd.n2913 gnd.n2912 240.244
R6083 gnd.n2912 gnd.n2911 240.244
R6084 gnd.n2911 gnd.n2885 240.244
R6085 gnd.n2907 gnd.n2885 240.244
R6086 gnd.n2907 gnd.n2906 240.244
R6087 gnd.n2906 gnd.n2905 240.244
R6088 gnd.n2905 gnd.n2891 240.244
R6089 gnd.n2901 gnd.n2891 240.244
R6090 gnd.n2901 gnd.n2900 240.244
R6091 gnd.n2900 gnd.n2793 240.244
R6092 gnd.n3239 gnd.n2793 240.244
R6093 gnd.n3240 gnd.n3239 240.244
R6094 gnd.n3240 gnd.n2789 240.244
R6095 gnd.n3246 gnd.n2789 240.244
R6096 gnd.n3247 gnd.n3246 240.244
R6097 gnd.n3248 gnd.n3247 240.244
R6098 gnd.n3248 gnd.n2785 240.244
R6099 gnd.n3254 gnd.n2785 240.244
R6100 gnd.n3255 gnd.n3254 240.244
R6101 gnd.n3256 gnd.n3255 240.244
R6102 gnd.n3256 gnd.n2781 240.244
R6103 gnd.n3262 gnd.n2781 240.244
R6104 gnd.n3262 gnd.n2780 240.244
R6105 gnd.n3399 gnd.n2780 240.244
R6106 gnd.n3399 gnd.n2776 240.244
R6107 gnd.n3405 gnd.n2776 240.244
R6108 gnd.n3405 gnd.n2774 240.244
R6109 gnd.n3413 gnd.n2774 240.244
R6110 gnd.n3413 gnd.n2770 240.244
R6111 gnd.n3419 gnd.n2770 240.244
R6112 gnd.n3419 gnd.n2766 240.244
R6113 gnd.n3427 gnd.n2766 240.244
R6114 gnd.n3427 gnd.n2762 240.244
R6115 gnd.n3433 gnd.n2762 240.244
R6116 gnd.n3433 gnd.n2758 240.244
R6117 gnd.n3444 gnd.n2758 240.244
R6118 gnd.n3444 gnd.n2754 240.244
R6119 gnd.n3450 gnd.n2754 240.244
R6120 gnd.n3450 gnd.n2753 240.244
R6121 gnd.n3458 gnd.n2753 240.244
R6122 gnd.n3458 gnd.n2748 240.244
R6123 gnd.n3466 gnd.n2748 240.244
R6124 gnd.n3466 gnd.n2749 240.244
R6125 gnd.n2749 gnd.n2399 240.244
R6126 gnd.n3647 gnd.n2399 240.244
R6127 gnd.n3647 gnd.n2395 240.244
R6128 gnd.n3653 gnd.n2395 240.244
R6129 gnd.n3653 gnd.n2378 240.244
R6130 gnd.n3676 gnd.n2378 240.244
R6131 gnd.n3676 gnd.n2373 240.244
R6132 gnd.n3684 gnd.n2373 240.244
R6133 gnd.n3684 gnd.n2374 240.244
R6134 gnd.n2374 gnd.n2351 240.244
R6135 gnd.n3714 gnd.n2351 240.244
R6136 gnd.n3714 gnd.n2346 240.244
R6137 gnd.n3722 gnd.n2346 240.244
R6138 gnd.n3722 gnd.n2347 240.244
R6139 gnd.n2347 gnd.n2324 240.244
R6140 gnd.n3750 gnd.n2324 240.244
R6141 gnd.n3750 gnd.n2320 240.244
R6142 gnd.n3756 gnd.n2320 240.244
R6143 gnd.n3756 gnd.n2302 240.244
R6144 gnd.n3778 gnd.n2302 240.244
R6145 gnd.n3778 gnd.n2297 240.244
R6146 gnd.n3786 gnd.n2297 240.244
R6147 gnd.n3786 gnd.n2298 240.244
R6148 gnd.n2298 gnd.n2274 240.244
R6149 gnd.n3828 gnd.n2274 240.244
R6150 gnd.n3828 gnd.n2270 240.244
R6151 gnd.n3836 gnd.n2270 240.244
R6152 gnd.n3836 gnd.n2255 240.244
R6153 gnd.n3854 gnd.n2255 240.244
R6154 gnd.n3855 gnd.n3854 240.244
R6155 gnd.n3855 gnd.n2251 240.244
R6156 gnd.n3861 gnd.n2251 240.244
R6157 gnd.n3861 gnd.n2210 240.244
R6158 gnd.n3898 gnd.n2210 240.244
R6159 gnd.n3898 gnd.n2206 240.244
R6160 gnd.n3904 gnd.n2206 240.244
R6161 gnd.n3904 gnd.n2188 240.244
R6162 gnd.n3940 gnd.n2188 240.244
R6163 gnd.n3940 gnd.n2181 240.244
R6164 gnd.n3948 gnd.n2181 240.244
R6165 gnd.n3948 gnd.n2184 240.244
R6166 gnd.n2184 gnd.n2161 240.244
R6167 gnd.n3992 gnd.n2161 240.244
R6168 gnd.n3992 gnd.n2156 240.244
R6169 gnd.n4000 gnd.n2156 240.244
R6170 gnd.n4000 gnd.n2157 240.244
R6171 gnd.n2157 gnd.n2130 240.244
R6172 gnd.n4043 gnd.n2130 240.244
R6173 gnd.n4043 gnd.n2126 240.244
R6174 gnd.n4049 gnd.n2126 240.244
R6175 gnd.n4049 gnd.n2115 240.244
R6176 gnd.n4075 gnd.n2115 240.244
R6177 gnd.n4075 gnd.n2107 240.244
R6178 gnd.n4086 gnd.n2107 240.244
R6179 gnd.n4086 gnd.n2111 240.244
R6180 gnd.n4082 gnd.n2111 240.244
R6181 gnd.n4082 gnd.n2080 240.244
R6182 gnd.n4149 gnd.n2080 240.244
R6183 gnd.n4149 gnd.n2075 240.244
R6184 gnd.n4157 gnd.n2075 240.244
R6185 gnd.n4157 gnd.n2076 240.244
R6186 gnd.n2076 gnd.n2052 240.244
R6187 gnd.n4192 gnd.n2052 240.244
R6188 gnd.n4192 gnd.n2045 240.244
R6189 gnd.n4203 gnd.n2045 240.244
R6190 gnd.n4203 gnd.n2048 240.244
R6191 gnd.n4199 gnd.n2048 240.244
R6192 gnd.n4199 gnd.n1846 240.244
R6193 gnd.n4378 gnd.n1846 240.244
R6194 gnd.n4378 gnd.n1842 240.244
R6195 gnd.n4384 gnd.n1842 240.244
R6196 gnd.n4384 gnd.n1833 240.244
R6197 gnd.n4398 gnd.n1833 240.244
R6198 gnd.n4398 gnd.n1829 240.244
R6199 gnd.n4404 gnd.n1829 240.244
R6200 gnd.n4404 gnd.n1820 240.244
R6201 gnd.n4418 gnd.n1820 240.244
R6202 gnd.n4418 gnd.n1816 240.244
R6203 gnd.n4424 gnd.n1816 240.244
R6204 gnd.n4424 gnd.n1807 240.244
R6205 gnd.n4441 gnd.n1807 240.244
R6206 gnd.n4441 gnd.n1803 240.244
R6207 gnd.n4448 gnd.n1803 240.244
R6208 gnd.n4448 gnd.n1459 240.244
R6209 gnd.n4735 gnd.n1459 240.244
R6210 gnd.n4735 gnd.n1460 240.244
R6211 gnd.n4731 gnd.n1460 240.244
R6212 gnd.n4731 gnd.n1466 240.244
R6213 gnd.n4727 gnd.n1466 240.244
R6214 gnd.n4727 gnd.n1469 240.244
R6215 gnd.n4723 gnd.n1469 240.244
R6216 gnd.n4723 gnd.n1475 240.244
R6217 gnd.n1627 gnd.n1475 240.244
R6218 gnd.n1627 gnd.n1624 240.244
R6219 gnd.n1633 gnd.n1624 240.244
R6220 gnd.n1633 gnd.n1615 240.244
R6221 gnd.n4536 gnd.n1615 240.244
R6222 gnd.n4536 gnd.n1609 240.244
R6223 gnd.n4544 gnd.n1609 240.244
R6224 gnd.n4544 gnd.n1611 240.244
R6225 gnd.n1611 gnd.n1588 240.244
R6226 gnd.n4569 gnd.n1588 240.244
R6227 gnd.n4569 gnd.n1582 240.244
R6228 gnd.n4584 gnd.n1582 240.244
R6229 gnd.n4584 gnd.n1584 240.244
R6230 gnd.n4580 gnd.n1584 240.244
R6231 gnd.n4580 gnd.n4579 240.244
R6232 gnd.n4579 gnd.n1529 240.244
R6233 gnd.n4674 gnd.n1529 240.244
R6234 gnd.n4674 gnd.n1531 240.244
R6235 gnd.n4670 gnd.n1531 240.244
R6236 gnd.n4670 gnd.n4669 240.244
R6237 gnd.n4669 gnd.n4668 240.244
R6238 gnd.n4668 gnd.n1538 240.244
R6239 gnd.n4663 gnd.n1538 240.244
R6240 gnd.n4663 gnd.n1540 240.244
R6241 gnd.n4655 gnd.n1540 240.244
R6242 gnd.n4655 gnd.n4647 240.244
R6243 gnd.n4650 gnd.n4647 240.244
R6244 gnd.n4650 gnd.n306 240.244
R6245 gnd.n7469 gnd.n306 240.244
R6246 gnd.n7469 gnd.n307 240.244
R6247 gnd.n7464 gnd.n307 240.244
R6248 gnd.n7464 gnd.n7463 240.244
R6249 gnd.n7463 gnd.n7462 240.244
R6250 gnd.n7462 gnd.n311 240.244
R6251 gnd.n7458 gnd.n311 240.244
R6252 gnd.n7458 gnd.n7457 240.244
R6253 gnd.n7457 gnd.n7456 240.244
R6254 gnd.n7456 gnd.n317 240.244
R6255 gnd.n7395 gnd.n317 240.244
R6256 gnd.n6691 gnd.n741 240.244
R6257 gnd.n6687 gnd.n741 240.244
R6258 gnd.n6687 gnd.n746 240.244
R6259 gnd.n6683 gnd.n746 240.244
R6260 gnd.n6683 gnd.n748 240.244
R6261 gnd.n6679 gnd.n748 240.244
R6262 gnd.n6679 gnd.n754 240.244
R6263 gnd.n6675 gnd.n754 240.244
R6264 gnd.n6675 gnd.n756 240.244
R6265 gnd.n6671 gnd.n756 240.244
R6266 gnd.n6671 gnd.n762 240.244
R6267 gnd.n6667 gnd.n762 240.244
R6268 gnd.n6667 gnd.n764 240.244
R6269 gnd.n6663 gnd.n764 240.244
R6270 gnd.n6663 gnd.n770 240.244
R6271 gnd.n6659 gnd.n770 240.244
R6272 gnd.n6659 gnd.n772 240.244
R6273 gnd.n6655 gnd.n772 240.244
R6274 gnd.n6655 gnd.n778 240.244
R6275 gnd.n6651 gnd.n778 240.244
R6276 gnd.n6651 gnd.n780 240.244
R6277 gnd.n6647 gnd.n780 240.244
R6278 gnd.n6647 gnd.n786 240.244
R6279 gnd.n6643 gnd.n786 240.244
R6280 gnd.n6643 gnd.n788 240.244
R6281 gnd.n6639 gnd.n788 240.244
R6282 gnd.n6639 gnd.n794 240.244
R6283 gnd.n6635 gnd.n794 240.244
R6284 gnd.n6635 gnd.n796 240.244
R6285 gnd.n6631 gnd.n796 240.244
R6286 gnd.n6631 gnd.n802 240.244
R6287 gnd.n6627 gnd.n802 240.244
R6288 gnd.n6627 gnd.n804 240.244
R6289 gnd.n6623 gnd.n804 240.244
R6290 gnd.n6623 gnd.n810 240.244
R6291 gnd.n6619 gnd.n810 240.244
R6292 gnd.n6619 gnd.n812 240.244
R6293 gnd.n6615 gnd.n812 240.244
R6294 gnd.n6615 gnd.n818 240.244
R6295 gnd.n6611 gnd.n818 240.244
R6296 gnd.n6611 gnd.n820 240.244
R6297 gnd.n6607 gnd.n820 240.244
R6298 gnd.n6607 gnd.n826 240.244
R6299 gnd.n6603 gnd.n826 240.244
R6300 gnd.n6603 gnd.n828 240.244
R6301 gnd.n6599 gnd.n828 240.244
R6302 gnd.n6599 gnd.n834 240.244
R6303 gnd.n6595 gnd.n834 240.244
R6304 gnd.n6595 gnd.n836 240.244
R6305 gnd.n6591 gnd.n836 240.244
R6306 gnd.n6591 gnd.n842 240.244
R6307 gnd.n6587 gnd.n842 240.244
R6308 gnd.n6587 gnd.n844 240.244
R6309 gnd.n6583 gnd.n844 240.244
R6310 gnd.n6583 gnd.n850 240.244
R6311 gnd.n6579 gnd.n850 240.244
R6312 gnd.n6579 gnd.n852 240.244
R6313 gnd.n6575 gnd.n852 240.244
R6314 gnd.n6575 gnd.n858 240.244
R6315 gnd.n6571 gnd.n858 240.244
R6316 gnd.n6571 gnd.n860 240.244
R6317 gnd.n6567 gnd.n860 240.244
R6318 gnd.n6567 gnd.n866 240.244
R6319 gnd.n6563 gnd.n866 240.244
R6320 gnd.n6563 gnd.n868 240.244
R6321 gnd.n6559 gnd.n868 240.244
R6322 gnd.n6559 gnd.n874 240.244
R6323 gnd.n6555 gnd.n874 240.244
R6324 gnd.n6555 gnd.n876 240.244
R6325 gnd.n6551 gnd.n876 240.244
R6326 gnd.n6551 gnd.n882 240.244
R6327 gnd.n6547 gnd.n882 240.244
R6328 gnd.n6547 gnd.n884 240.244
R6329 gnd.n6543 gnd.n884 240.244
R6330 gnd.n6543 gnd.n890 240.244
R6331 gnd.n6539 gnd.n890 240.244
R6332 gnd.n6539 gnd.n892 240.244
R6333 gnd.n6535 gnd.n892 240.244
R6334 gnd.n6535 gnd.n898 240.244
R6335 gnd.n6531 gnd.n898 240.244
R6336 gnd.n6531 gnd.n900 240.244
R6337 gnd.n6527 gnd.n900 240.244
R6338 gnd.n6527 gnd.n906 240.244
R6339 gnd.n2859 gnd.n906 240.244
R6340 gnd.n1330 gnd.n1329 240.244
R6341 gnd.n1331 gnd.n1330 240.244
R6342 gnd.n2768 gnd.n1331 240.244
R6343 gnd.n2768 gnd.n1334 240.244
R6344 gnd.n1335 gnd.n1334 240.244
R6345 gnd.n1336 gnd.n1335 240.244
R6346 gnd.n2760 gnd.n1336 240.244
R6347 gnd.n2760 gnd.n1339 240.244
R6348 gnd.n1340 gnd.n1339 240.244
R6349 gnd.n1341 gnd.n1340 240.244
R6350 gnd.n3439 gnd.n1341 240.244
R6351 gnd.n3439 gnd.n1344 240.244
R6352 gnd.n1345 gnd.n1344 240.244
R6353 gnd.n1346 gnd.n1345 240.244
R6354 gnd.n2746 gnd.n1346 240.244
R6355 gnd.n2746 gnd.n1349 240.244
R6356 gnd.n1350 gnd.n1349 240.244
R6357 gnd.n1351 gnd.n1350 240.244
R6358 gnd.n2402 gnd.n1351 240.244
R6359 gnd.n2402 gnd.n1354 240.244
R6360 gnd.n1355 gnd.n1354 240.244
R6361 gnd.n1356 gnd.n1355 240.244
R6362 gnd.n3672 gnd.n1356 240.244
R6363 gnd.n3672 gnd.n1359 240.244
R6364 gnd.n1360 gnd.n1359 240.244
R6365 gnd.n1361 gnd.n1360 240.244
R6366 gnd.n3703 gnd.n1361 240.244
R6367 gnd.n3703 gnd.n1364 240.244
R6368 gnd.n1365 gnd.n1364 240.244
R6369 gnd.n1366 gnd.n1365 240.244
R6370 gnd.n2499 gnd.n1366 240.244
R6371 gnd.n2499 gnd.n1369 240.244
R6372 gnd.n1370 gnd.n1369 240.244
R6373 gnd.n1371 gnd.n1370 240.244
R6374 gnd.n2308 gnd.n1371 240.244
R6375 gnd.n2308 gnd.n1374 240.244
R6376 gnd.n1375 gnd.n1374 240.244
R6377 gnd.n1376 gnd.n1375 240.244
R6378 gnd.n3796 gnd.n1376 240.244
R6379 gnd.n3796 gnd.n1379 240.244
R6380 gnd.n1380 gnd.n1379 240.244
R6381 gnd.n1381 gnd.n1380 240.244
R6382 gnd.n2267 gnd.n1381 240.244
R6383 gnd.n2267 gnd.n1384 240.244
R6384 gnd.n1385 gnd.n1384 240.244
R6385 gnd.n1386 gnd.n1385 240.244
R6386 gnd.n3870 gnd.n1386 240.244
R6387 gnd.n3870 gnd.n1389 240.244
R6388 gnd.n1390 gnd.n1389 240.244
R6389 gnd.n1391 gnd.n1390 240.244
R6390 gnd.n2213 gnd.n1391 240.244
R6391 gnd.n2213 gnd.n1394 240.244
R6392 gnd.n1395 gnd.n1394 240.244
R6393 gnd.n1396 gnd.n1395 240.244
R6394 gnd.n3936 gnd.n1396 240.244
R6395 gnd.n3936 gnd.n1399 240.244
R6396 gnd.n1400 gnd.n1399 240.244
R6397 gnd.n1401 gnd.n1400 240.244
R6398 gnd.n2162 gnd.n1401 240.244
R6399 gnd.n2162 gnd.n1404 240.244
R6400 gnd.n1405 gnd.n1404 240.244
R6401 gnd.n1406 gnd.n1405 240.244
R6402 gnd.n3966 gnd.n1406 240.244
R6403 gnd.n3966 gnd.n1409 240.244
R6404 gnd.n1410 gnd.n1409 240.244
R6405 gnd.n1411 gnd.n1410 240.244
R6406 gnd.n4016 gnd.n1411 240.244
R6407 gnd.n4016 gnd.n1414 240.244
R6408 gnd.n1415 gnd.n1414 240.244
R6409 gnd.n1416 gnd.n1415 240.244
R6410 gnd.n4097 gnd.n1416 240.244
R6411 gnd.n4097 gnd.n1419 240.244
R6412 gnd.n1420 gnd.n1419 240.244
R6413 gnd.n1421 gnd.n1420 240.244
R6414 gnd.n2083 gnd.n1421 240.244
R6415 gnd.n2083 gnd.n1424 240.244
R6416 gnd.n1425 gnd.n1424 240.244
R6417 gnd.n1426 gnd.n1425 240.244
R6418 gnd.n4181 gnd.n1426 240.244
R6419 gnd.n4181 gnd.n1429 240.244
R6420 gnd.n1430 gnd.n1429 240.244
R6421 gnd.n1431 gnd.n1430 240.244
R6422 gnd.n2036 gnd.n1431 240.244
R6423 gnd.n2036 gnd.n1434 240.244
R6424 gnd.n1435 gnd.n1434 240.244
R6425 gnd.n1436 gnd.n1435 240.244
R6426 gnd.n1840 gnd.n1436 240.244
R6427 gnd.n1840 gnd.n1439 240.244
R6428 gnd.n1440 gnd.n1439 240.244
R6429 gnd.n1441 gnd.n1440 240.244
R6430 gnd.n1827 gnd.n1441 240.244
R6431 gnd.n1827 gnd.n1444 240.244
R6432 gnd.n1445 gnd.n1444 240.244
R6433 gnd.n1446 gnd.n1445 240.244
R6434 gnd.n1814 gnd.n1446 240.244
R6435 gnd.n1814 gnd.n1449 240.244
R6436 gnd.n1450 gnd.n1449 240.244
R6437 gnd.n1451 gnd.n1450 240.244
R6438 gnd.n4436 gnd.n1451 240.244
R6439 gnd.n4436 gnd.n1454 240.244
R6440 gnd.n4738 gnd.n1454 240.244
R6441 gnd.n3281 gnd.n3280 240.244
R6442 gnd.n3296 gnd.n3280 240.244
R6443 gnd.n3298 gnd.n3297 240.244
R6444 gnd.n3308 gnd.n3307 240.244
R6445 gnd.n3319 gnd.n3318 240.244
R6446 gnd.n3321 gnd.n3320 240.244
R6447 gnd.n3331 gnd.n3330 240.244
R6448 gnd.n3344 gnd.n3343 240.244
R6449 gnd.n3346 gnd.n3345 240.244
R6450 gnd.n2709 gnd.n2708 240.244
R6451 gnd.n3274 gnd.n2710 240.244
R6452 gnd.n2714 gnd.n2713 240.244
R6453 gnd.n2720 gnd.n2715 240.244
R6454 gnd.n2722 gnd.n2721 240.244
R6455 gnd.n2726 gnd.n2725 240.244
R6456 gnd.n2727 gnd.n2726 240.244
R6457 gnd.n2767 gnd.n2727 240.244
R6458 gnd.n2767 gnd.n2730 240.244
R6459 gnd.n2731 gnd.n2730 240.244
R6460 gnd.n2732 gnd.n2731 240.244
R6461 gnd.n2759 gnd.n2732 240.244
R6462 gnd.n2759 gnd.n2735 240.244
R6463 gnd.n2736 gnd.n2735 240.244
R6464 gnd.n2737 gnd.n2736 240.244
R6465 gnd.n3438 gnd.n2737 240.244
R6466 gnd.n3438 gnd.n2740 240.244
R6467 gnd.n2741 gnd.n2740 240.244
R6468 gnd.n2742 gnd.n2741 240.244
R6469 gnd.n2745 gnd.n2742 240.244
R6470 gnd.n3469 gnd.n2745 240.244
R6471 gnd.n3470 gnd.n3469 240.244
R6472 gnd.n3473 gnd.n3470 240.244
R6473 gnd.n3474 gnd.n3473 240.244
R6474 gnd.n3474 gnd.n2385 240.244
R6475 gnd.n3665 gnd.n2385 240.244
R6476 gnd.n3665 gnd.n2381 240.244
R6477 gnd.n3671 gnd.n2381 240.244
R6478 gnd.n3671 gnd.n2365 240.244
R6479 gnd.n3695 gnd.n2365 240.244
R6480 gnd.n3695 gnd.n2359 240.244
R6481 gnd.n3702 gnd.n2359 240.244
R6482 gnd.n3702 gnd.n2360 240.244
R6483 gnd.n2360 gnd.n2338 240.244
R6484 gnd.n3732 gnd.n2338 240.244
R6485 gnd.n3732 gnd.n2334 240.244
R6486 gnd.n3738 gnd.n2334 240.244
R6487 gnd.n3738 gnd.n2318 240.244
R6488 gnd.n3759 gnd.n2318 240.244
R6489 gnd.n3759 gnd.n2312 240.244
R6490 gnd.n3766 gnd.n2312 240.244
R6491 gnd.n3766 gnd.n2313 240.244
R6492 gnd.n2313 gnd.n2288 240.244
R6493 gnd.n3798 gnd.n2288 240.244
R6494 gnd.n3798 gnd.n2283 240.244
R6495 gnd.n3818 gnd.n2283 240.244
R6496 gnd.n3818 gnd.n2277 240.244
R6497 gnd.n3803 gnd.n2277 240.244
R6498 gnd.n3806 gnd.n3803 240.244
R6499 gnd.n3807 gnd.n3806 240.244
R6500 gnd.n3807 gnd.n2257 240.244
R6501 gnd.n2257 gnd.n2226 240.244
R6502 gnd.n3880 gnd.n2226 240.244
R6503 gnd.n3880 gnd.n2220 240.244
R6504 gnd.n3887 gnd.n2220 240.244
R6505 gnd.n3887 gnd.n2221 240.244
R6506 gnd.n2221 gnd.n2196 240.244
R6507 gnd.n3916 gnd.n2196 240.244
R6508 gnd.n3916 gnd.n2191 240.244
R6509 gnd.n3935 gnd.n2191 240.244
R6510 gnd.n3935 gnd.n2180 240.244
R6511 gnd.n3921 gnd.n2180 240.244
R6512 gnd.n3922 gnd.n3921 240.244
R6513 gnd.n3923 gnd.n3922 240.244
R6514 gnd.n3924 gnd.n3923 240.244
R6515 gnd.n3924 gnd.n2147 240.244
R6516 gnd.n4010 gnd.n2147 240.244
R6517 gnd.n4010 gnd.n2142 240.244
R6518 gnd.n4031 gnd.n2142 240.244
R6519 gnd.n4031 gnd.n2132 240.244
R6520 gnd.n4015 gnd.n2132 240.244
R6521 gnd.n4018 gnd.n4015 240.244
R6522 gnd.n4019 gnd.n4018 240.244
R6523 gnd.n4020 gnd.n4019 240.244
R6524 gnd.n4020 gnd.n2098 240.244
R6525 gnd.n4099 gnd.n2098 240.244
R6526 gnd.n4099 gnd.n2092 240.244
R6527 gnd.n4109 gnd.n2092 240.244
R6528 gnd.n4109 gnd.n2093 240.244
R6529 gnd.n4103 gnd.n2093 240.244
R6530 gnd.n4103 gnd.n2067 240.244
R6531 gnd.n4167 gnd.n2067 240.244
R6532 gnd.n4167 gnd.n2062 240.244
R6533 gnd.n4180 gnd.n2062 240.244
R6534 gnd.n4180 gnd.n2054 240.244
R6535 gnd.n4172 gnd.n2054 240.244
R6536 gnd.n4173 gnd.n4172 240.244
R6537 gnd.n4173 gnd.n1851 240.244
R6538 gnd.n4368 gnd.n1851 240.244
R6539 gnd.n4368 gnd.n1847 240.244
R6540 gnd.n4374 gnd.n1847 240.244
R6541 gnd.n4374 gnd.n1839 240.244
R6542 gnd.n4388 gnd.n1839 240.244
R6543 gnd.n4388 gnd.n1835 240.244
R6544 gnd.n4394 gnd.n1835 240.244
R6545 gnd.n4394 gnd.n1826 240.244
R6546 gnd.n4408 gnd.n1826 240.244
R6547 gnd.n4408 gnd.n1822 240.244
R6548 gnd.n4414 gnd.n1822 240.244
R6549 gnd.n4414 gnd.n1813 240.244
R6550 gnd.n4428 gnd.n1813 240.244
R6551 gnd.n4428 gnd.n1809 240.244
R6552 gnd.n4435 gnd.n1809 240.244
R6553 gnd.n4435 gnd.n1802 240.244
R6554 gnd.n4451 gnd.n1802 240.244
R6555 gnd.n4451 gnd.n1457 240.244
R6556 gnd.n1700 gnd.n1699 240.244
R6557 gnd.n1716 gnd.n1715 240.244
R6558 gnd.n1719 gnd.n1718 240.244
R6559 gnd.n1735 gnd.n1734 240.244
R6560 gnd.n1738 gnd.n1737 240.244
R6561 gnd.n1754 gnd.n1753 240.244
R6562 gnd.n1757 gnd.n1756 240.244
R6563 gnd.n1773 gnd.n1772 240.244
R6564 gnd.n1776 gnd.n1775 240.244
R6565 gnd.n1781 gnd.n1778 240.244
R6566 gnd.n1784 gnd.n1783 240.244
R6567 gnd.n1792 gnd.n1786 240.244
R6568 gnd.n1795 gnd.n1794 240.244
R6569 gnd.n1798 gnd.n1797 240.244
R6570 gnd.n2411 gnd.n2410 240.132
R6571 gnd.n4220 gnd.n4219 240.132
R6572 gnd.n6694 gnd.n6693 225.874
R6573 gnd.n6694 gnd.n734 225.874
R6574 gnd.n6702 gnd.n734 225.874
R6575 gnd.n6703 gnd.n6702 225.874
R6576 gnd.n6704 gnd.n6703 225.874
R6577 gnd.n6704 gnd.n728 225.874
R6578 gnd.n6712 gnd.n728 225.874
R6579 gnd.n6713 gnd.n6712 225.874
R6580 gnd.n6714 gnd.n6713 225.874
R6581 gnd.n6714 gnd.n722 225.874
R6582 gnd.n6722 gnd.n722 225.874
R6583 gnd.n6723 gnd.n6722 225.874
R6584 gnd.n6724 gnd.n6723 225.874
R6585 gnd.n6724 gnd.n716 225.874
R6586 gnd.n6732 gnd.n716 225.874
R6587 gnd.n6733 gnd.n6732 225.874
R6588 gnd.n6734 gnd.n6733 225.874
R6589 gnd.n6734 gnd.n710 225.874
R6590 gnd.n6742 gnd.n710 225.874
R6591 gnd.n6743 gnd.n6742 225.874
R6592 gnd.n6744 gnd.n6743 225.874
R6593 gnd.n6744 gnd.n704 225.874
R6594 gnd.n6752 gnd.n704 225.874
R6595 gnd.n6753 gnd.n6752 225.874
R6596 gnd.n6754 gnd.n6753 225.874
R6597 gnd.n6754 gnd.n698 225.874
R6598 gnd.n6762 gnd.n698 225.874
R6599 gnd.n6763 gnd.n6762 225.874
R6600 gnd.n6764 gnd.n6763 225.874
R6601 gnd.n6764 gnd.n692 225.874
R6602 gnd.n6772 gnd.n692 225.874
R6603 gnd.n6773 gnd.n6772 225.874
R6604 gnd.n6774 gnd.n6773 225.874
R6605 gnd.n6774 gnd.n686 225.874
R6606 gnd.n6782 gnd.n686 225.874
R6607 gnd.n6783 gnd.n6782 225.874
R6608 gnd.n6784 gnd.n6783 225.874
R6609 gnd.n6784 gnd.n680 225.874
R6610 gnd.n6792 gnd.n680 225.874
R6611 gnd.n6793 gnd.n6792 225.874
R6612 gnd.n6794 gnd.n6793 225.874
R6613 gnd.n6794 gnd.n674 225.874
R6614 gnd.n6802 gnd.n674 225.874
R6615 gnd.n6803 gnd.n6802 225.874
R6616 gnd.n6804 gnd.n6803 225.874
R6617 gnd.n6804 gnd.n668 225.874
R6618 gnd.n6812 gnd.n668 225.874
R6619 gnd.n6813 gnd.n6812 225.874
R6620 gnd.n6814 gnd.n6813 225.874
R6621 gnd.n6814 gnd.n662 225.874
R6622 gnd.n6822 gnd.n662 225.874
R6623 gnd.n6823 gnd.n6822 225.874
R6624 gnd.n6824 gnd.n6823 225.874
R6625 gnd.n6824 gnd.n656 225.874
R6626 gnd.n6832 gnd.n656 225.874
R6627 gnd.n6833 gnd.n6832 225.874
R6628 gnd.n6834 gnd.n6833 225.874
R6629 gnd.n6834 gnd.n650 225.874
R6630 gnd.n6842 gnd.n650 225.874
R6631 gnd.n6843 gnd.n6842 225.874
R6632 gnd.n6844 gnd.n6843 225.874
R6633 gnd.n6844 gnd.n644 225.874
R6634 gnd.n6852 gnd.n644 225.874
R6635 gnd.n6853 gnd.n6852 225.874
R6636 gnd.n6854 gnd.n6853 225.874
R6637 gnd.n6854 gnd.n638 225.874
R6638 gnd.n6862 gnd.n638 225.874
R6639 gnd.n6863 gnd.n6862 225.874
R6640 gnd.n6864 gnd.n6863 225.874
R6641 gnd.n6864 gnd.n632 225.874
R6642 gnd.n6872 gnd.n632 225.874
R6643 gnd.n6873 gnd.n6872 225.874
R6644 gnd.n6874 gnd.n6873 225.874
R6645 gnd.n6874 gnd.n626 225.874
R6646 gnd.n6882 gnd.n626 225.874
R6647 gnd.n6883 gnd.n6882 225.874
R6648 gnd.n6884 gnd.n6883 225.874
R6649 gnd.n6884 gnd.n620 225.874
R6650 gnd.n6892 gnd.n620 225.874
R6651 gnd.n6893 gnd.n6892 225.874
R6652 gnd.n6894 gnd.n6893 225.874
R6653 gnd.n6894 gnd.n614 225.874
R6654 gnd.n6902 gnd.n614 225.874
R6655 gnd.n6903 gnd.n6902 225.874
R6656 gnd.n6904 gnd.n6903 225.874
R6657 gnd.n6904 gnd.n608 225.874
R6658 gnd.n6912 gnd.n608 225.874
R6659 gnd.n6913 gnd.n6912 225.874
R6660 gnd.n6914 gnd.n6913 225.874
R6661 gnd.n6914 gnd.n602 225.874
R6662 gnd.n6922 gnd.n602 225.874
R6663 gnd.n6923 gnd.n6922 225.874
R6664 gnd.n6924 gnd.n6923 225.874
R6665 gnd.n6924 gnd.n596 225.874
R6666 gnd.n6932 gnd.n596 225.874
R6667 gnd.n6933 gnd.n6932 225.874
R6668 gnd.n6934 gnd.n6933 225.874
R6669 gnd.n6934 gnd.n590 225.874
R6670 gnd.n6942 gnd.n590 225.874
R6671 gnd.n6943 gnd.n6942 225.874
R6672 gnd.n6944 gnd.n6943 225.874
R6673 gnd.n6944 gnd.n584 225.874
R6674 gnd.n6952 gnd.n584 225.874
R6675 gnd.n6953 gnd.n6952 225.874
R6676 gnd.n6954 gnd.n6953 225.874
R6677 gnd.n6954 gnd.n578 225.874
R6678 gnd.n6962 gnd.n578 225.874
R6679 gnd.n6963 gnd.n6962 225.874
R6680 gnd.n6964 gnd.n6963 225.874
R6681 gnd.n6964 gnd.n572 225.874
R6682 gnd.n6972 gnd.n572 225.874
R6683 gnd.n6973 gnd.n6972 225.874
R6684 gnd.n6974 gnd.n6973 225.874
R6685 gnd.n6974 gnd.n566 225.874
R6686 gnd.n6982 gnd.n566 225.874
R6687 gnd.n6983 gnd.n6982 225.874
R6688 gnd.n6984 gnd.n6983 225.874
R6689 gnd.n6984 gnd.n560 225.874
R6690 gnd.n6992 gnd.n560 225.874
R6691 gnd.n6993 gnd.n6992 225.874
R6692 gnd.n6994 gnd.n6993 225.874
R6693 gnd.n6994 gnd.n554 225.874
R6694 gnd.n7002 gnd.n554 225.874
R6695 gnd.n7003 gnd.n7002 225.874
R6696 gnd.n7004 gnd.n7003 225.874
R6697 gnd.n7004 gnd.n548 225.874
R6698 gnd.n7012 gnd.n548 225.874
R6699 gnd.n7013 gnd.n7012 225.874
R6700 gnd.n7014 gnd.n7013 225.874
R6701 gnd.n7014 gnd.n542 225.874
R6702 gnd.n7022 gnd.n542 225.874
R6703 gnd.n7023 gnd.n7022 225.874
R6704 gnd.n7024 gnd.n7023 225.874
R6705 gnd.n7024 gnd.n536 225.874
R6706 gnd.n7032 gnd.n536 225.874
R6707 gnd.n7033 gnd.n7032 225.874
R6708 gnd.n7034 gnd.n7033 225.874
R6709 gnd.n7034 gnd.n530 225.874
R6710 gnd.n7042 gnd.n530 225.874
R6711 gnd.n7043 gnd.n7042 225.874
R6712 gnd.n7044 gnd.n7043 225.874
R6713 gnd.n7044 gnd.n524 225.874
R6714 gnd.n7052 gnd.n524 225.874
R6715 gnd.n7053 gnd.n7052 225.874
R6716 gnd.n7054 gnd.n7053 225.874
R6717 gnd.n7054 gnd.n518 225.874
R6718 gnd.n7062 gnd.n518 225.874
R6719 gnd.n7063 gnd.n7062 225.874
R6720 gnd.n7064 gnd.n7063 225.874
R6721 gnd.n7064 gnd.n512 225.874
R6722 gnd.n7072 gnd.n512 225.874
R6723 gnd.n7073 gnd.n7072 225.874
R6724 gnd.n7074 gnd.n7073 225.874
R6725 gnd.n7074 gnd.n506 225.874
R6726 gnd.n7082 gnd.n506 225.874
R6727 gnd.n7083 gnd.n7082 225.874
R6728 gnd.n7084 gnd.n7083 225.874
R6729 gnd.n7084 gnd.n500 225.874
R6730 gnd.n7092 gnd.n500 225.874
R6731 gnd.n7093 gnd.n7092 225.874
R6732 gnd.n7094 gnd.n7093 225.874
R6733 gnd.n7094 gnd.n494 225.874
R6734 gnd.n7102 gnd.n494 225.874
R6735 gnd.n7103 gnd.n7102 225.874
R6736 gnd.n7104 gnd.n7103 225.874
R6737 gnd.n7104 gnd.n488 225.874
R6738 gnd.n7112 gnd.n488 225.874
R6739 gnd.n7113 gnd.n7112 225.874
R6740 gnd.n7114 gnd.n7113 225.874
R6741 gnd.n7114 gnd.n482 225.874
R6742 gnd.n7122 gnd.n482 225.874
R6743 gnd.n7123 gnd.n7122 225.874
R6744 gnd.n7124 gnd.n7123 225.874
R6745 gnd.n7124 gnd.n476 225.874
R6746 gnd.n7132 gnd.n476 225.874
R6747 gnd.n7133 gnd.n7132 225.874
R6748 gnd.n7134 gnd.n7133 225.874
R6749 gnd.n7134 gnd.n470 225.874
R6750 gnd.n7142 gnd.n470 225.874
R6751 gnd.n7143 gnd.n7142 225.874
R6752 gnd.n7144 gnd.n7143 225.874
R6753 gnd.n7144 gnd.n464 225.874
R6754 gnd.n7152 gnd.n464 225.874
R6755 gnd.n7153 gnd.n7152 225.874
R6756 gnd.n7154 gnd.n7153 225.874
R6757 gnd.n7154 gnd.n458 225.874
R6758 gnd.n7162 gnd.n458 225.874
R6759 gnd.n7163 gnd.n7162 225.874
R6760 gnd.n7164 gnd.n7163 225.874
R6761 gnd.n7164 gnd.n452 225.874
R6762 gnd.n7173 gnd.n452 225.874
R6763 gnd.n7174 gnd.n7173 225.874
R6764 gnd.n7175 gnd.n7174 225.874
R6765 gnd.n7175 gnd.n447 225.874
R6766 gnd.n5554 gnd.t226 224.174
R6767 gnd.n5184 gnd.t184 224.174
R6768 gnd.n1893 gnd.n1890 199.319
R6769 gnd.n2027 gnd.n1890 199.319
R6770 gnd.n2613 gnd.n2607 199.319
R6771 gnd.n2612 gnd.n2607 199.319
R6772 gnd.n2412 gnd.n2409 186.49
R6773 gnd.n4221 gnd.n4218 186.49
R6774 gnd.n6373 gnd.n6372 185
R6775 gnd.n6371 gnd.n6370 185
R6776 gnd.n6350 gnd.n6349 185
R6777 gnd.n6365 gnd.n6364 185
R6778 gnd.n6363 gnd.n6362 185
R6779 gnd.n6354 gnd.n6353 185
R6780 gnd.n6357 gnd.n6356 185
R6781 gnd.n6341 gnd.n6340 185
R6782 gnd.n6339 gnd.n6338 185
R6783 gnd.n6318 gnd.n6317 185
R6784 gnd.n6333 gnd.n6332 185
R6785 gnd.n6331 gnd.n6330 185
R6786 gnd.n6322 gnd.n6321 185
R6787 gnd.n6325 gnd.n6324 185
R6788 gnd.n6309 gnd.n6308 185
R6789 gnd.n6307 gnd.n6306 185
R6790 gnd.n6286 gnd.n6285 185
R6791 gnd.n6301 gnd.n6300 185
R6792 gnd.n6299 gnd.n6298 185
R6793 gnd.n6290 gnd.n6289 185
R6794 gnd.n6293 gnd.n6292 185
R6795 gnd.n6278 gnd.n6277 185
R6796 gnd.n6276 gnd.n6275 185
R6797 gnd.n6255 gnd.n6254 185
R6798 gnd.n6270 gnd.n6269 185
R6799 gnd.n6268 gnd.n6267 185
R6800 gnd.n6259 gnd.n6258 185
R6801 gnd.n6262 gnd.n6261 185
R6802 gnd.n6246 gnd.n6245 185
R6803 gnd.n6244 gnd.n6243 185
R6804 gnd.n6223 gnd.n6222 185
R6805 gnd.n6238 gnd.n6237 185
R6806 gnd.n6236 gnd.n6235 185
R6807 gnd.n6227 gnd.n6226 185
R6808 gnd.n6230 gnd.n6229 185
R6809 gnd.n6214 gnd.n6213 185
R6810 gnd.n6212 gnd.n6211 185
R6811 gnd.n6191 gnd.n6190 185
R6812 gnd.n6206 gnd.n6205 185
R6813 gnd.n6204 gnd.n6203 185
R6814 gnd.n6195 gnd.n6194 185
R6815 gnd.n6198 gnd.n6197 185
R6816 gnd.n6182 gnd.n6181 185
R6817 gnd.n6180 gnd.n6179 185
R6818 gnd.n6159 gnd.n6158 185
R6819 gnd.n6174 gnd.n6173 185
R6820 gnd.n6172 gnd.n6171 185
R6821 gnd.n6163 gnd.n6162 185
R6822 gnd.n6166 gnd.n6165 185
R6823 gnd.n6151 gnd.n6150 185
R6824 gnd.n6149 gnd.n6148 185
R6825 gnd.n6128 gnd.n6127 185
R6826 gnd.n6143 gnd.n6142 185
R6827 gnd.n6141 gnd.n6140 185
R6828 gnd.n6132 gnd.n6131 185
R6829 gnd.n6135 gnd.n6134 185
R6830 gnd.n5555 gnd.t225 178.987
R6831 gnd.n5185 gnd.t185 178.987
R6832 gnd.n1 gnd.t30 170.774
R6833 gnd.n9 gnd.t91 170.103
R6834 gnd.n8 gnd.t40 170.103
R6835 gnd.n7 gnd.t311 170.103
R6836 gnd.n6 gnd.t38 170.103
R6837 gnd.n5 gnd.t299 170.103
R6838 gnd.n4 gnd.t294 170.103
R6839 gnd.n3 gnd.t331 170.103
R6840 gnd.n2 gnd.t85 170.103
R6841 gnd.n1 gnd.t1 170.103
R6842 gnd.n4292 gnd.n4291 163.367
R6843 gnd.n4288 gnd.n4287 163.367
R6844 gnd.n4284 gnd.n4283 163.367
R6845 gnd.n4280 gnd.n4279 163.367
R6846 gnd.n4276 gnd.n4275 163.367
R6847 gnd.n4272 gnd.n4271 163.367
R6848 gnd.n4268 gnd.n4267 163.367
R6849 gnd.n4264 gnd.n4263 163.367
R6850 gnd.n4260 gnd.n4259 163.367
R6851 gnd.n4256 gnd.n4255 163.367
R6852 gnd.n4252 gnd.n4251 163.367
R6853 gnd.n4248 gnd.n4247 163.367
R6854 gnd.n4244 gnd.n4243 163.367
R6855 gnd.n4240 gnd.n4239 163.367
R6856 gnd.n4235 gnd.n4234 163.367
R6857 gnd.n4231 gnd.n4230 163.367
R6858 gnd.n4365 gnd.n4364 163.367
R6859 gnd.n4361 gnd.n4360 163.367
R6860 gnd.n4356 gnd.n4355 163.367
R6861 gnd.n4352 gnd.n4351 163.367
R6862 gnd.n4348 gnd.n4347 163.367
R6863 gnd.n4344 gnd.n4343 163.367
R6864 gnd.n4340 gnd.n4339 163.367
R6865 gnd.n4336 gnd.n4335 163.367
R6866 gnd.n4332 gnd.n4331 163.367
R6867 gnd.n4328 gnd.n4327 163.367
R6868 gnd.n4324 gnd.n4323 163.367
R6869 gnd.n4320 gnd.n4319 163.367
R6870 gnd.n4316 gnd.n4315 163.367
R6871 gnd.n4312 gnd.n4311 163.367
R6872 gnd.n4308 gnd.n4307 163.367
R6873 gnd.n4304 gnd.n4303 163.367
R6874 gnd.n2538 gnd.n2401 163.367
R6875 gnd.n2534 gnd.n2401 163.367
R6876 gnd.n2534 gnd.n2394 163.367
R6877 gnd.n2529 gnd.n2394 163.367
R6878 gnd.n2529 gnd.n2387 163.367
R6879 gnd.n2526 gnd.n2387 163.367
R6880 gnd.n2526 gnd.n2380 163.367
R6881 gnd.n2380 gnd.n2371 163.367
R6882 gnd.n2372 gnd.n2371 163.367
R6883 gnd.n2372 gnd.n2366 163.367
R6884 gnd.n2520 gnd.n2366 163.367
R6885 gnd.n2520 gnd.n2358 163.367
R6886 gnd.n2515 gnd.n2358 163.367
R6887 gnd.n2515 gnd.n2353 163.367
R6888 gnd.n2512 gnd.n2353 163.367
R6889 gnd.n2512 gnd.n2345 163.367
R6890 gnd.n2506 gnd.n2345 163.367
R6891 gnd.n2506 gnd.n2339 163.367
R6892 gnd.n2502 gnd.n2339 163.367
R6893 gnd.n2502 gnd.n2333 163.367
R6894 gnd.n2496 gnd.n2333 163.367
R6895 gnd.n2496 gnd.n2326 163.367
R6896 gnd.n2493 gnd.n2326 163.367
R6897 gnd.n2493 gnd.n2491 163.367
R6898 gnd.n2491 gnd.n2310 163.367
R6899 gnd.n2311 gnd.n2310 163.367
R6900 gnd.n2311 gnd.n2303 163.367
R6901 gnd.n2485 gnd.n2303 163.367
R6902 gnd.n2485 gnd.n2295 163.367
R6903 gnd.n2481 gnd.n2295 163.367
R6904 gnd.n2481 gnd.n2289 163.367
R6905 gnd.n2478 gnd.n2289 163.367
R6906 gnd.n2478 gnd.n2282 163.367
R6907 gnd.n2473 gnd.n2282 163.367
R6908 gnd.n2473 gnd.n2276 163.367
R6909 gnd.n2470 gnd.n2276 163.367
R6910 gnd.n2470 gnd.n2269 163.367
R6911 gnd.n2269 gnd.n2260 163.367
R6912 gnd.n3846 gnd.n2260 163.367
R6913 gnd.n3846 gnd.n2258 163.367
R6914 gnd.n3850 gnd.n2258 163.367
R6915 gnd.n3850 gnd.n2233 163.367
R6916 gnd.n3868 gnd.n2233 163.367
R6917 gnd.n3868 gnd.n2228 163.367
R6918 gnd.n3864 gnd.n2228 163.367
R6919 gnd.n3864 gnd.n2219 163.367
R6920 gnd.n2248 gnd.n2219 163.367
R6921 gnd.n2248 gnd.n2212 163.367
R6922 gnd.n2245 gnd.n2212 163.367
R6923 gnd.n2245 gnd.n2205 163.367
R6924 gnd.n2240 gnd.n2205 163.367
R6925 gnd.n2240 gnd.n2198 163.367
R6926 gnd.n2237 gnd.n2198 163.367
R6927 gnd.n2237 gnd.n2190 163.367
R6928 gnd.n2190 gnd.n2179 163.367
R6929 gnd.n2179 gnd.n2173 163.367
R6930 gnd.n3959 gnd.n2173 163.367
R6931 gnd.n3959 gnd.n2170 163.367
R6932 gnd.n3982 gnd.n2170 163.367
R6933 gnd.n3982 gnd.n2171 163.367
R6934 gnd.n2171 gnd.n2164 163.367
R6935 gnd.n3977 gnd.n2164 163.367
R6936 gnd.n3977 gnd.n2155 163.367
R6937 gnd.n3972 gnd.n2155 163.367
R6938 gnd.n3972 gnd.n2149 163.367
R6939 gnd.n3969 gnd.n2149 163.367
R6940 gnd.n3969 gnd.n2141 163.367
R6941 gnd.n3963 gnd.n2141 163.367
R6942 gnd.n3963 gnd.n2133 163.367
R6943 gnd.n2133 gnd.n2124 163.367
R6944 gnd.n4052 gnd.n2124 163.367
R6945 gnd.n4052 gnd.n2122 163.367
R6946 gnd.n4064 gnd.n2122 163.367
R6947 gnd.n4064 gnd.n2117 163.367
R6948 gnd.n4060 gnd.n2117 163.367
R6949 gnd.n4060 gnd.n2106 163.367
R6950 gnd.n4056 gnd.n2106 163.367
R6951 gnd.n4056 gnd.n2100 163.367
R6952 gnd.n2100 gnd.n2090 163.367
R6953 gnd.n4112 gnd.n2090 163.367
R6954 gnd.n4112 gnd.n2088 163.367
R6955 gnd.n4138 gnd.n2088 163.367
R6956 gnd.n4138 gnd.n2082 163.367
R6957 gnd.n4134 gnd.n2082 163.367
R6958 gnd.n4134 gnd.n2074 163.367
R6959 gnd.n4129 gnd.n2074 163.367
R6960 gnd.n4129 gnd.n2069 163.367
R6961 gnd.n4126 gnd.n2069 163.367
R6962 gnd.n4126 gnd.n2061 163.367
R6963 gnd.n4121 gnd.n2061 163.367
R6964 gnd.n4121 gnd.n2055 163.367
R6965 gnd.n4118 gnd.n2055 163.367
R6966 gnd.n4118 gnd.n2043 163.367
R6967 gnd.n2043 gnd.n2035 163.367
R6968 gnd.n4299 gnd.n2035 163.367
R6969 gnd.n3636 gnd.n2426 163.367
R6970 gnd.n3636 gnd.n2461 163.367
R6971 gnd.n3632 gnd.n3631 163.367
R6972 gnd.n3628 gnd.n3627 163.367
R6973 gnd.n3624 gnd.n3623 163.367
R6974 gnd.n3620 gnd.n3619 163.367
R6975 gnd.n3616 gnd.n3615 163.367
R6976 gnd.n3612 gnd.n3611 163.367
R6977 gnd.n3608 gnd.n3607 163.367
R6978 gnd.n3604 gnd.n3603 163.367
R6979 gnd.n3600 gnd.n3599 163.367
R6980 gnd.n3596 gnd.n3595 163.367
R6981 gnd.n3592 gnd.n3591 163.367
R6982 gnd.n3588 gnd.n3587 163.367
R6983 gnd.n3584 gnd.n3583 163.367
R6984 gnd.n3580 gnd.n3579 163.367
R6985 gnd.n3576 gnd.n3575 163.367
R6986 gnd.n2600 gnd.n2599 163.367
R6987 gnd.n2595 gnd.n2594 163.367
R6988 gnd.n2591 gnd.n2590 163.367
R6989 gnd.n2587 gnd.n2586 163.367
R6990 gnd.n2583 gnd.n2582 163.367
R6991 gnd.n2579 gnd.n2578 163.367
R6992 gnd.n2575 gnd.n2574 163.367
R6993 gnd.n2571 gnd.n2570 163.367
R6994 gnd.n2567 gnd.n2566 163.367
R6995 gnd.n2563 gnd.n2562 163.367
R6996 gnd.n2559 gnd.n2558 163.367
R6997 gnd.n2555 gnd.n2554 163.367
R6998 gnd.n2551 gnd.n2550 163.367
R6999 gnd.n2547 gnd.n2546 163.367
R7000 gnd.n2543 gnd.n2542 163.367
R7001 gnd.n3644 gnd.n2404 163.367
R7002 gnd.n3644 gnd.n2392 163.367
R7003 gnd.n3656 gnd.n2392 163.367
R7004 gnd.n3656 gnd.n2389 163.367
R7005 gnd.n3661 gnd.n2389 163.367
R7006 gnd.n3661 gnd.n2390 163.367
R7007 gnd.n2390 gnd.n2369 163.367
R7008 gnd.n3689 gnd.n2369 163.367
R7009 gnd.n3689 gnd.n2367 163.367
R7010 gnd.n3693 gnd.n2367 163.367
R7011 gnd.n3693 gnd.n2356 163.367
R7012 gnd.n3707 gnd.n2356 163.367
R7013 gnd.n3707 gnd.n2354 163.367
R7014 gnd.n3711 gnd.n2354 163.367
R7015 gnd.n3711 gnd.n2343 163.367
R7016 gnd.n3725 gnd.n2343 163.367
R7017 gnd.n3725 gnd.n2341 163.367
R7018 gnd.n3729 gnd.n2341 163.367
R7019 gnd.n3729 gnd.n2331 163.367
R7020 gnd.n3741 gnd.n2331 163.367
R7021 gnd.n3741 gnd.n2328 163.367
R7022 gnd.n3746 gnd.n2328 163.367
R7023 gnd.n3746 gnd.n2329 163.367
R7024 gnd.n2329 gnd.n2307 163.367
R7025 gnd.n3771 gnd.n2307 163.367
R7026 gnd.n3771 gnd.n2305 163.367
R7027 gnd.n3775 gnd.n2305 163.367
R7028 gnd.n3775 gnd.n2293 163.367
R7029 gnd.n3790 gnd.n2293 163.367
R7030 gnd.n3790 gnd.n2291 163.367
R7031 gnd.n3794 gnd.n2291 163.367
R7032 gnd.n3794 gnd.n2280 163.367
R7033 gnd.n3821 gnd.n2280 163.367
R7034 gnd.n3821 gnd.n2278 163.367
R7035 gnd.n3825 gnd.n2278 163.367
R7036 gnd.n3825 gnd.n2266 163.367
R7037 gnd.n3839 gnd.n2266 163.367
R7038 gnd.n3839 gnd.n2263 163.367
R7039 gnd.n3844 gnd.n2263 163.367
R7040 gnd.n3844 gnd.n2264 163.367
R7041 gnd.n2264 gnd.n2231 163.367
R7042 gnd.n3873 gnd.n2231 163.367
R7043 gnd.n3873 gnd.n2229 163.367
R7044 gnd.n3877 gnd.n2229 163.367
R7045 gnd.n3877 gnd.n2217 163.367
R7046 gnd.n3891 gnd.n2217 163.367
R7047 gnd.n3891 gnd.n2215 163.367
R7048 gnd.n3895 gnd.n2215 163.367
R7049 gnd.n3895 gnd.n2203 163.367
R7050 gnd.n3907 gnd.n2203 163.367
R7051 gnd.n3907 gnd.n2200 163.367
R7052 gnd.n3912 gnd.n2200 163.367
R7053 gnd.n3912 gnd.n2201 163.367
R7054 gnd.n2201 gnd.n2177 163.367
R7055 gnd.n3953 gnd.n2177 163.367
R7056 gnd.n3953 gnd.n2175 163.367
R7057 gnd.n3957 gnd.n2175 163.367
R7058 gnd.n3957 gnd.n2168 163.367
R7059 gnd.n3985 gnd.n2168 163.367
R7060 gnd.n3985 gnd.n2166 163.367
R7061 gnd.n3989 gnd.n2166 163.367
R7062 gnd.n3989 gnd.n2153 163.367
R7063 gnd.n4003 gnd.n2153 163.367
R7064 gnd.n4003 gnd.n2151 163.367
R7065 gnd.n4007 gnd.n2151 163.367
R7066 gnd.n4007 gnd.n2139 163.367
R7067 gnd.n4034 gnd.n2139 163.367
R7068 gnd.n4034 gnd.n2135 163.367
R7069 gnd.n4039 gnd.n2135 163.367
R7070 gnd.n4039 gnd.n2137 163.367
R7071 gnd.n2137 gnd.n2121 163.367
R7072 gnd.n4068 gnd.n2121 163.367
R7073 gnd.n4068 gnd.n2119 163.367
R7074 gnd.n4072 gnd.n2119 163.367
R7075 gnd.n4072 gnd.n2104 163.367
R7076 gnd.n4090 gnd.n2104 163.367
R7077 gnd.n4090 gnd.n2101 163.367
R7078 gnd.n4095 gnd.n2101 163.367
R7079 gnd.n4095 gnd.n2102 163.367
R7080 gnd.n2102 gnd.n2087 163.367
R7081 gnd.n4142 gnd.n2087 163.367
R7082 gnd.n4142 gnd.n2085 163.367
R7083 gnd.n4146 gnd.n2085 163.367
R7084 gnd.n4146 gnd.n2073 163.367
R7085 gnd.n4160 gnd.n2073 163.367
R7086 gnd.n4160 gnd.n2071 163.367
R7087 gnd.n4164 gnd.n2071 163.367
R7088 gnd.n4164 gnd.n2059 163.367
R7089 gnd.n4184 gnd.n2059 163.367
R7090 gnd.n4184 gnd.n2057 163.367
R7091 gnd.n4188 gnd.n2057 163.367
R7092 gnd.n4188 gnd.n2041 163.367
R7093 gnd.n4206 gnd.n2041 163.367
R7094 gnd.n4206 gnd.n2038 163.367
R7095 gnd.n4297 gnd.n2038 163.367
R7096 gnd.n7184 gnd.n7183 157.537
R7097 gnd.n7185 gnd.n7184 157.537
R7098 gnd.n7185 gnd.n441 157.537
R7099 gnd.n7193 gnd.n441 157.537
R7100 gnd.n7194 gnd.n7193 157.537
R7101 gnd.n7195 gnd.n7194 157.537
R7102 gnd.n7195 gnd.n435 157.537
R7103 gnd.n7203 gnd.n435 157.537
R7104 gnd.n7204 gnd.n7203 157.537
R7105 gnd.n7205 gnd.n7204 157.537
R7106 gnd.n7205 gnd.n429 157.537
R7107 gnd.n7213 gnd.n429 157.537
R7108 gnd.n7214 gnd.n7213 157.537
R7109 gnd.n7215 gnd.n7214 157.537
R7110 gnd.n7215 gnd.n423 157.537
R7111 gnd.n7223 gnd.n423 157.537
R7112 gnd.n7224 gnd.n7223 157.537
R7113 gnd.n7225 gnd.n7224 157.537
R7114 gnd.n7225 gnd.n417 157.537
R7115 gnd.n7233 gnd.n417 157.537
R7116 gnd.n7234 gnd.n7233 157.537
R7117 gnd.n7235 gnd.n7234 157.537
R7118 gnd.n7235 gnd.n411 157.537
R7119 gnd.n7243 gnd.n411 157.537
R7120 gnd.n7244 gnd.n7243 157.537
R7121 gnd.n7245 gnd.n7244 157.537
R7122 gnd.n7245 gnd.n405 157.537
R7123 gnd.n7253 gnd.n405 157.537
R7124 gnd.n7254 gnd.n7253 157.537
R7125 gnd.n7255 gnd.n7254 157.537
R7126 gnd.n7255 gnd.n399 157.537
R7127 gnd.n7263 gnd.n399 157.537
R7128 gnd.n7264 gnd.n7263 157.537
R7129 gnd.n7265 gnd.n7264 157.537
R7130 gnd.n7265 gnd.n393 157.537
R7131 gnd.n7273 gnd.n393 157.537
R7132 gnd.n7274 gnd.n7273 157.537
R7133 gnd.n7275 gnd.n7274 157.537
R7134 gnd.n7275 gnd.n387 157.537
R7135 gnd.n7283 gnd.n387 157.537
R7136 gnd.n7284 gnd.n7283 157.537
R7137 gnd.n7285 gnd.n7284 157.537
R7138 gnd.n7285 gnd.n381 157.537
R7139 gnd.n7293 gnd.n381 157.537
R7140 gnd.n7294 gnd.n7293 157.537
R7141 gnd.n7295 gnd.n7294 157.537
R7142 gnd.n7295 gnd.n375 157.537
R7143 gnd.n7303 gnd.n375 157.537
R7144 gnd.n7304 gnd.n7303 157.537
R7145 gnd.n7305 gnd.n7304 157.537
R7146 gnd.n7305 gnd.n369 157.537
R7147 gnd.n7313 gnd.n369 157.537
R7148 gnd.n7314 gnd.n7313 157.537
R7149 gnd.n7315 gnd.n7314 157.537
R7150 gnd.n7315 gnd.n363 157.537
R7151 gnd.n7323 gnd.n363 157.537
R7152 gnd.n7324 gnd.n7323 157.537
R7153 gnd.n7325 gnd.n7324 157.537
R7154 gnd.n7325 gnd.n357 157.537
R7155 gnd.n7333 gnd.n357 157.537
R7156 gnd.n7334 gnd.n7333 157.537
R7157 gnd.n7335 gnd.n7334 157.537
R7158 gnd.n7335 gnd.n351 157.537
R7159 gnd.n7343 gnd.n351 157.537
R7160 gnd.n7344 gnd.n7343 157.537
R7161 gnd.n7345 gnd.n7344 157.537
R7162 gnd.n7345 gnd.n345 157.537
R7163 gnd.n7353 gnd.n345 157.537
R7164 gnd.n7354 gnd.n7353 157.537
R7165 gnd.n7355 gnd.n7354 157.537
R7166 gnd.n7355 gnd.n339 157.537
R7167 gnd.n7363 gnd.n339 157.537
R7168 gnd.n7364 gnd.n7363 157.537
R7169 gnd.n7365 gnd.n7364 157.537
R7170 gnd.n7365 gnd.n333 157.537
R7171 gnd.n7373 gnd.n333 157.537
R7172 gnd.n7374 gnd.n7373 157.537
R7173 gnd.n7375 gnd.n7374 157.537
R7174 gnd.n7375 gnd.n327 157.537
R7175 gnd.n7383 gnd.n327 157.537
R7176 gnd.n7384 gnd.n7383 157.537
R7177 gnd.n7386 gnd.n7384 157.537
R7178 gnd.n7386 gnd.n7385 157.537
R7179 gnd.n4227 gnd.n4226 156.462
R7180 gnd.n6313 gnd.n6281 153.042
R7181 gnd.n6377 gnd.n6376 152.079
R7182 gnd.n6345 gnd.n6344 152.079
R7183 gnd.n6313 gnd.n6312 152.079
R7184 gnd.n2417 gnd.n2416 152
R7185 gnd.n2418 gnd.n2407 152
R7186 gnd.n2420 gnd.n2419 152
R7187 gnd.n2422 gnd.n2405 152
R7188 gnd.n2424 gnd.n2423 152
R7189 gnd.n4225 gnd.n4209 152
R7190 gnd.n4217 gnd.n4210 152
R7191 gnd.n4216 gnd.n4215 152
R7192 gnd.n4214 gnd.n4211 152
R7193 gnd.n4212 gnd.t206 150.546
R7194 gnd.t150 gnd.n6355 147.661
R7195 gnd.t319 gnd.n6323 147.661
R7196 gnd.t71 gnd.n6291 147.661
R7197 gnd.t83 gnd.n6260 147.661
R7198 gnd.t106 gnd.n6228 147.661
R7199 gnd.t111 gnd.n6196 147.661
R7200 gnd.t87 gnd.n6164 147.661
R7201 gnd.t307 gnd.n6133 147.661
R7202 gnd.n1888 gnd.n1869 143.351
R7203 gnd.n3574 gnd.n2442 143.351
R7204 gnd.n3574 gnd.n2443 143.351
R7205 gnd.n2031 gnd.n2030 138.177
R7206 gnd.n3577 gnd.n3573 138.177
R7207 gnd.n2414 gnd.t247 130.484
R7208 gnd.n2423 gnd.t262 126.766
R7209 gnd.n2421 gnd.t217 126.766
R7210 gnd.n2407 gnd.t253 126.766
R7211 gnd.n2415 gnd.t237 126.766
R7212 gnd.n4213 gnd.t179 126.766
R7213 gnd.n4215 gnd.t281 126.766
R7214 gnd.n4224 gnd.t240 126.766
R7215 gnd.n4226 gnd.t230 126.766
R7216 gnd.n6372 gnd.n6371 104.615
R7217 gnd.n6371 gnd.n6349 104.615
R7218 gnd.n6364 gnd.n6349 104.615
R7219 gnd.n6364 gnd.n6363 104.615
R7220 gnd.n6363 gnd.n6353 104.615
R7221 gnd.n6356 gnd.n6353 104.615
R7222 gnd.n6340 gnd.n6339 104.615
R7223 gnd.n6339 gnd.n6317 104.615
R7224 gnd.n6332 gnd.n6317 104.615
R7225 gnd.n6332 gnd.n6331 104.615
R7226 gnd.n6331 gnd.n6321 104.615
R7227 gnd.n6324 gnd.n6321 104.615
R7228 gnd.n6308 gnd.n6307 104.615
R7229 gnd.n6307 gnd.n6285 104.615
R7230 gnd.n6300 gnd.n6285 104.615
R7231 gnd.n6300 gnd.n6299 104.615
R7232 gnd.n6299 gnd.n6289 104.615
R7233 gnd.n6292 gnd.n6289 104.615
R7234 gnd.n6277 gnd.n6276 104.615
R7235 gnd.n6276 gnd.n6254 104.615
R7236 gnd.n6269 gnd.n6254 104.615
R7237 gnd.n6269 gnd.n6268 104.615
R7238 gnd.n6268 gnd.n6258 104.615
R7239 gnd.n6261 gnd.n6258 104.615
R7240 gnd.n6245 gnd.n6244 104.615
R7241 gnd.n6244 gnd.n6222 104.615
R7242 gnd.n6237 gnd.n6222 104.615
R7243 gnd.n6237 gnd.n6236 104.615
R7244 gnd.n6236 gnd.n6226 104.615
R7245 gnd.n6229 gnd.n6226 104.615
R7246 gnd.n6213 gnd.n6212 104.615
R7247 gnd.n6212 gnd.n6190 104.615
R7248 gnd.n6205 gnd.n6190 104.615
R7249 gnd.n6205 gnd.n6204 104.615
R7250 gnd.n6204 gnd.n6194 104.615
R7251 gnd.n6197 gnd.n6194 104.615
R7252 gnd.n6181 gnd.n6180 104.615
R7253 gnd.n6180 gnd.n6158 104.615
R7254 gnd.n6173 gnd.n6158 104.615
R7255 gnd.n6173 gnd.n6172 104.615
R7256 gnd.n6172 gnd.n6162 104.615
R7257 gnd.n6165 gnd.n6162 104.615
R7258 gnd.n6150 gnd.n6149 104.615
R7259 gnd.n6149 gnd.n6127 104.615
R7260 gnd.n6142 gnd.n6127 104.615
R7261 gnd.n6142 gnd.n6141 104.615
R7262 gnd.n6141 gnd.n6131 104.615
R7263 gnd.n6134 gnd.n6131 104.615
R7264 gnd.n5704 gnd.t268 100.632
R7265 gnd.n5158 gnd.t200 100.632
R7266 gnd.n7732 gnd.n116 99.6594
R7267 gnd.n7730 gnd.n7729 99.6594
R7268 gnd.n7725 gnd.n124 99.6594
R7269 gnd.n7723 gnd.n7722 99.6594
R7270 gnd.n7718 gnd.n131 99.6594
R7271 gnd.n7716 gnd.n7715 99.6594
R7272 gnd.n7711 gnd.n138 99.6594
R7273 gnd.n7709 gnd.n7708 99.6594
R7274 gnd.n7701 gnd.n145 99.6594
R7275 gnd.n7699 gnd.n7698 99.6594
R7276 gnd.n7694 gnd.n152 99.6594
R7277 gnd.n7692 gnd.n7691 99.6594
R7278 gnd.n7687 gnd.n159 99.6594
R7279 gnd.n7685 gnd.n7684 99.6594
R7280 gnd.n7680 gnd.n166 99.6594
R7281 gnd.n7678 gnd.n7677 99.6594
R7282 gnd.n7673 gnd.n173 99.6594
R7283 gnd.n7671 gnd.n7670 99.6594
R7284 gnd.n178 gnd.n177 99.6594
R7285 gnd.n1910 gnd.n1909 99.6594
R7286 gnd.n1918 gnd.n1917 99.6594
R7287 gnd.n1921 gnd.n1920 99.6594
R7288 gnd.n1928 gnd.n1927 99.6594
R7289 gnd.n1931 gnd.n1930 99.6594
R7290 gnd.n1939 gnd.n1938 99.6594
R7291 gnd.n1942 gnd.n1941 99.6594
R7292 gnd.n1894 gnd.n1893 99.6594
R7293 gnd.n2026 gnd.n2025 99.6594
R7294 gnd.n2019 gnd.n1952 99.6594
R7295 gnd.n2018 gnd.n2017 99.6594
R7296 gnd.n2011 gnd.n1958 99.6594
R7297 gnd.n2010 gnd.n2009 99.6594
R7298 gnd.n2003 gnd.n1964 99.6594
R7299 gnd.n2002 gnd.n2001 99.6594
R7300 gnd.n1995 gnd.n1970 99.6594
R7301 gnd.n1994 gnd.n1993 99.6594
R7302 gnd.n1985 gnd.n1976 99.6594
R7303 gnd.n2665 gnd.n2664 99.6594
R7304 gnd.n2660 gnd.n2619 99.6594
R7305 gnd.n2656 gnd.n2618 99.6594
R7306 gnd.n2652 gnd.n2617 99.6594
R7307 gnd.n2648 gnd.n2616 99.6594
R7308 gnd.n2644 gnd.n2615 99.6594
R7309 gnd.n2640 gnd.n2614 99.6594
R7310 gnd.n2612 gnd.n2611 99.6594
R7311 gnd.n3567 gnd.n3566 99.6594
R7312 gnd.n3564 gnd.n3563 99.6594
R7313 gnd.n3559 gnd.n2674 99.6594
R7314 gnd.n3557 gnd.n3556 99.6594
R7315 gnd.n3552 gnd.n2681 99.6594
R7316 gnd.n3550 gnd.n3549 99.6594
R7317 gnd.n3545 gnd.n2688 99.6594
R7318 gnd.n3543 gnd.n3542 99.6594
R7319 gnd.n3538 gnd.n2697 99.6594
R7320 gnd.n3536 gnd.n3535 99.6594
R7321 gnd.n5134 gnd.n5133 99.6594
R7322 gnd.n5128 gnd.n981 99.6594
R7323 gnd.n5125 gnd.n982 99.6594
R7324 gnd.n5121 gnd.n983 99.6594
R7325 gnd.n5117 gnd.n984 99.6594
R7326 gnd.n5113 gnd.n985 99.6594
R7327 gnd.n5109 gnd.n986 99.6594
R7328 gnd.n5105 gnd.n987 99.6594
R7329 gnd.n5101 gnd.n988 99.6594
R7330 gnd.n5096 gnd.n989 99.6594
R7331 gnd.n5092 gnd.n990 99.6594
R7332 gnd.n5088 gnd.n991 99.6594
R7333 gnd.n5084 gnd.n992 99.6594
R7334 gnd.n5080 gnd.n993 99.6594
R7335 gnd.n5076 gnd.n994 99.6594
R7336 gnd.n5072 gnd.n995 99.6594
R7337 gnd.n5068 gnd.n996 99.6594
R7338 gnd.n5064 gnd.n997 99.6594
R7339 gnd.n1052 gnd.n998 99.6594
R7340 gnd.n6486 gnd.n6485 99.6594
R7341 gnd.n6481 gnd.n5142 99.6594
R7342 gnd.n6477 gnd.n5141 99.6594
R7343 gnd.n6473 gnd.n5140 99.6594
R7344 gnd.n6469 gnd.n5139 99.6594
R7345 gnd.n6465 gnd.n5138 99.6594
R7346 gnd.n6461 gnd.n5137 99.6594
R7347 gnd.n6388 gnd.n5136 99.6594
R7348 gnd.n5737 gnd.n5736 99.6594
R7349 gnd.n5731 gnd.n5679 99.6594
R7350 gnd.n5728 gnd.n5680 99.6594
R7351 gnd.n5724 gnd.n5681 99.6594
R7352 gnd.n5720 gnd.n5682 99.6594
R7353 gnd.n5716 gnd.n5683 99.6594
R7354 gnd.n5712 gnd.n5684 99.6594
R7355 gnd.n5708 gnd.n5685 99.6594
R7356 gnd.n6451 gnd.n968 99.6594
R7357 gnd.n6447 gnd.n969 99.6594
R7358 gnd.n6443 gnd.n970 99.6594
R7359 gnd.n6439 gnd.n971 99.6594
R7360 gnd.n6435 gnd.n972 99.6594
R7361 gnd.n6431 gnd.n973 99.6594
R7362 gnd.n6427 gnd.n974 99.6594
R7363 gnd.n6423 gnd.n975 99.6594
R7364 gnd.n6419 gnd.n976 99.6594
R7365 gnd.n6415 gnd.n977 99.6594
R7366 gnd.n6411 gnd.n978 99.6594
R7367 gnd.n6407 gnd.n979 99.6594
R7368 gnd.n6403 gnd.n980 99.6594
R7369 gnd.n5609 gnd.n5519 99.6594
R7370 gnd.n5607 gnd.n5522 99.6594
R7371 gnd.n5603 gnd.n5602 99.6594
R7372 gnd.n5596 gnd.n5527 99.6594
R7373 gnd.n5595 gnd.n5594 99.6594
R7374 gnd.n5588 gnd.n5533 99.6594
R7375 gnd.n5587 gnd.n5586 99.6594
R7376 gnd.n5580 gnd.n5539 99.6594
R7377 gnd.n5579 gnd.n5578 99.6594
R7378 gnd.n5572 gnd.n5545 99.6594
R7379 gnd.n5571 gnd.n5570 99.6594
R7380 gnd.n5563 gnd.n5551 99.6594
R7381 gnd.n5562 gnd.n5561 99.6594
R7382 gnd.n7580 gnd.n7579 99.6594
R7383 gnd.n7585 gnd.n7584 99.6594
R7384 gnd.n7588 gnd.n7587 99.6594
R7385 gnd.n7593 gnd.n7592 99.6594
R7386 gnd.n7596 gnd.n7595 99.6594
R7387 gnd.n7601 gnd.n7600 99.6594
R7388 gnd.n7604 gnd.n7603 99.6594
R7389 gnd.n7609 gnd.n7608 99.6594
R7390 gnd.n7612 gnd.n103 99.6594
R7391 gnd.n1687 gnd.n1686 99.6594
R7392 gnd.n1706 gnd.n1705 99.6594
R7393 gnd.n1709 gnd.n1708 99.6594
R7394 gnd.n1725 gnd.n1724 99.6594
R7395 gnd.n1728 gnd.n1727 99.6594
R7396 gnd.n1744 gnd.n1743 99.6594
R7397 gnd.n1747 gnd.n1746 99.6594
R7398 gnd.n1763 gnd.n1762 99.6594
R7399 gnd.n1766 gnd.n1765 99.6594
R7400 gnd.n3290 gnd.n3289 99.6594
R7401 gnd.n3293 gnd.n3292 99.6594
R7402 gnd.n3303 gnd.n3302 99.6594
R7403 gnd.n3312 gnd.n3311 99.6594
R7404 gnd.n3315 gnd.n3314 99.6594
R7405 gnd.n3326 gnd.n3325 99.6594
R7406 gnd.n3335 gnd.n3334 99.6594
R7407 gnd.n3338 gnd.n3337 99.6594
R7408 gnd.n3349 gnd.n3348 99.6594
R7409 gnd.n3021 gnd.n999 99.6594
R7410 gnd.n3018 gnd.n1000 99.6594
R7411 gnd.n3014 gnd.n1001 99.6594
R7412 gnd.n3010 gnd.n1002 99.6594
R7413 gnd.n3006 gnd.n1003 99.6594
R7414 gnd.n3002 gnd.n1004 99.6594
R7415 gnd.n2998 gnd.n1005 99.6594
R7416 gnd.n2994 gnd.n1006 99.6594
R7417 gnd.n2990 gnd.n1007 99.6594
R7418 gnd.n3019 gnd.n999 99.6594
R7419 gnd.n3015 gnd.n1000 99.6594
R7420 gnd.n3011 gnd.n1001 99.6594
R7421 gnd.n3007 gnd.n1002 99.6594
R7422 gnd.n3003 gnd.n1003 99.6594
R7423 gnd.n2999 gnd.n1004 99.6594
R7424 gnd.n2995 gnd.n1005 99.6594
R7425 gnd.n2991 gnd.n1006 99.6594
R7426 gnd.n2978 gnd.n1007 99.6594
R7427 gnd.n3348 gnd.n3347 99.6594
R7428 gnd.n3337 gnd.n3336 99.6594
R7429 gnd.n3334 gnd.n3327 99.6594
R7430 gnd.n3325 gnd.n3324 99.6594
R7431 gnd.n3314 gnd.n3313 99.6594
R7432 gnd.n3311 gnd.n3304 99.6594
R7433 gnd.n3302 gnd.n3301 99.6594
R7434 gnd.n3292 gnd.n3291 99.6594
R7435 gnd.n3289 gnd.n3288 99.6594
R7436 gnd.n1686 gnd.n1682 99.6594
R7437 gnd.n1707 gnd.n1706 99.6594
R7438 gnd.n1708 gnd.n1673 99.6594
R7439 gnd.n1726 gnd.n1725 99.6594
R7440 gnd.n1727 gnd.n1664 99.6594
R7441 gnd.n1745 gnd.n1744 99.6594
R7442 gnd.n1746 gnd.n1655 99.6594
R7443 gnd.n1764 gnd.n1763 99.6594
R7444 gnd.n1765 gnd.n1644 99.6594
R7445 gnd.n7613 gnd.n7612 99.6594
R7446 gnd.n7608 gnd.n7607 99.6594
R7447 gnd.n7603 gnd.n7602 99.6594
R7448 gnd.n7600 gnd.n7599 99.6594
R7449 gnd.n7595 gnd.n7594 99.6594
R7450 gnd.n7592 gnd.n7591 99.6594
R7451 gnd.n7587 gnd.n7586 99.6594
R7452 gnd.n7584 gnd.n7583 99.6594
R7453 gnd.n7579 gnd.n7578 99.6594
R7454 gnd.n5610 gnd.n5609 99.6594
R7455 gnd.n5604 gnd.n5522 99.6594
R7456 gnd.n5602 gnd.n5601 99.6594
R7457 gnd.n5597 gnd.n5596 99.6594
R7458 gnd.n5594 gnd.n5593 99.6594
R7459 gnd.n5589 gnd.n5588 99.6594
R7460 gnd.n5586 gnd.n5585 99.6594
R7461 gnd.n5581 gnd.n5580 99.6594
R7462 gnd.n5578 gnd.n5577 99.6594
R7463 gnd.n5573 gnd.n5572 99.6594
R7464 gnd.n5570 gnd.n5569 99.6594
R7465 gnd.n5564 gnd.n5563 99.6594
R7466 gnd.n5561 gnd.n5517 99.6594
R7467 gnd.n6406 gnd.n980 99.6594
R7468 gnd.n6410 gnd.n979 99.6594
R7469 gnd.n6414 gnd.n978 99.6594
R7470 gnd.n6418 gnd.n977 99.6594
R7471 gnd.n6422 gnd.n976 99.6594
R7472 gnd.n6426 gnd.n975 99.6594
R7473 gnd.n6430 gnd.n974 99.6594
R7474 gnd.n6434 gnd.n973 99.6594
R7475 gnd.n6438 gnd.n972 99.6594
R7476 gnd.n6442 gnd.n971 99.6594
R7477 gnd.n6446 gnd.n970 99.6594
R7478 gnd.n6450 gnd.n969 99.6594
R7479 gnd.n5162 gnd.n968 99.6594
R7480 gnd.n5737 gnd.n5687 99.6594
R7481 gnd.n5729 gnd.n5679 99.6594
R7482 gnd.n5725 gnd.n5680 99.6594
R7483 gnd.n5721 gnd.n5681 99.6594
R7484 gnd.n5717 gnd.n5682 99.6594
R7485 gnd.n5713 gnd.n5683 99.6594
R7486 gnd.n5709 gnd.n5684 99.6594
R7487 gnd.n5685 gnd.n5479 99.6594
R7488 gnd.n6460 gnd.n5136 99.6594
R7489 gnd.n6464 gnd.n5137 99.6594
R7490 gnd.n6468 gnd.n5138 99.6594
R7491 gnd.n6472 gnd.n5139 99.6594
R7492 gnd.n6476 gnd.n5140 99.6594
R7493 gnd.n6480 gnd.n5141 99.6594
R7494 gnd.n5143 gnd.n5142 99.6594
R7495 gnd.n6486 gnd.n965 99.6594
R7496 gnd.n5134 gnd.n1011 99.6594
R7497 gnd.n5126 gnd.n981 99.6594
R7498 gnd.n5122 gnd.n982 99.6594
R7499 gnd.n5118 gnd.n983 99.6594
R7500 gnd.n5114 gnd.n984 99.6594
R7501 gnd.n5110 gnd.n985 99.6594
R7502 gnd.n5106 gnd.n986 99.6594
R7503 gnd.n5102 gnd.n987 99.6594
R7504 gnd.n5097 gnd.n988 99.6594
R7505 gnd.n5093 gnd.n989 99.6594
R7506 gnd.n5089 gnd.n990 99.6594
R7507 gnd.n5085 gnd.n991 99.6594
R7508 gnd.n5081 gnd.n992 99.6594
R7509 gnd.n5077 gnd.n993 99.6594
R7510 gnd.n5073 gnd.n994 99.6594
R7511 gnd.n5069 gnd.n995 99.6594
R7512 gnd.n5065 gnd.n996 99.6594
R7513 gnd.n1051 gnd.n997 99.6594
R7514 gnd.n5057 gnd.n998 99.6594
R7515 gnd.n3537 gnd.n3536 99.6594
R7516 gnd.n2697 gnd.n2689 99.6594
R7517 gnd.n3544 gnd.n3543 99.6594
R7518 gnd.n2688 gnd.n2682 99.6594
R7519 gnd.n3551 gnd.n3550 99.6594
R7520 gnd.n2681 gnd.n2675 99.6594
R7521 gnd.n3558 gnd.n3557 99.6594
R7522 gnd.n2674 gnd.n2668 99.6594
R7523 gnd.n3565 gnd.n3564 99.6594
R7524 gnd.n3568 gnd.n3567 99.6594
R7525 gnd.n2639 gnd.n2613 99.6594
R7526 gnd.n2643 gnd.n2614 99.6594
R7527 gnd.n2647 gnd.n2615 99.6594
R7528 gnd.n2651 gnd.n2616 99.6594
R7529 gnd.n2655 gnd.n2617 99.6594
R7530 gnd.n2659 gnd.n2618 99.6594
R7531 gnd.n2621 gnd.n2619 99.6594
R7532 gnd.n2665 gnd.n2620 99.6594
R7533 gnd.n1911 gnd.n1910 99.6594
R7534 gnd.n1919 gnd.n1918 99.6594
R7535 gnd.n1920 gnd.n1900 99.6594
R7536 gnd.n1929 gnd.n1928 99.6594
R7537 gnd.n1930 gnd.n1896 99.6594
R7538 gnd.n1940 gnd.n1939 99.6594
R7539 gnd.n1943 gnd.n1942 99.6594
R7540 gnd.n2028 gnd.n2027 99.6594
R7541 gnd.n2025 gnd.n2024 99.6594
R7542 gnd.n2020 gnd.n2019 99.6594
R7543 gnd.n2017 gnd.n2016 99.6594
R7544 gnd.n2012 gnd.n2011 99.6594
R7545 gnd.n2009 gnd.n2008 99.6594
R7546 gnd.n2004 gnd.n2003 99.6594
R7547 gnd.n2001 gnd.n2000 99.6594
R7548 gnd.n1996 gnd.n1995 99.6594
R7549 gnd.n1993 gnd.n1992 99.6594
R7550 gnd.n1986 gnd.n1985 99.6594
R7551 gnd.n177 gnd.n174 99.6594
R7552 gnd.n7672 gnd.n7671 99.6594
R7553 gnd.n173 gnd.n167 99.6594
R7554 gnd.n7679 gnd.n7678 99.6594
R7555 gnd.n166 gnd.n160 99.6594
R7556 gnd.n7686 gnd.n7685 99.6594
R7557 gnd.n159 gnd.n153 99.6594
R7558 gnd.n7693 gnd.n7692 99.6594
R7559 gnd.n152 gnd.n146 99.6594
R7560 gnd.n7700 gnd.n7699 99.6594
R7561 gnd.n145 gnd.n139 99.6594
R7562 gnd.n7710 gnd.n7709 99.6594
R7563 gnd.n138 gnd.n132 99.6594
R7564 gnd.n7717 gnd.n7716 99.6594
R7565 gnd.n131 gnd.n125 99.6594
R7566 gnd.n7724 gnd.n7723 99.6594
R7567 gnd.n124 gnd.n118 99.6594
R7568 gnd.n7731 gnd.n7730 99.6594
R7569 gnd.n116 gnd.n113 99.6594
R7570 gnd.n3396 gnd.n3395 99.6594
R7571 gnd.n3296 gnd.n3265 99.6594
R7572 gnd.n3298 gnd.n3266 99.6594
R7573 gnd.n3308 gnd.n3267 99.6594
R7574 gnd.n3319 gnd.n3268 99.6594
R7575 gnd.n3321 gnd.n3269 99.6594
R7576 gnd.n3331 gnd.n3270 99.6594
R7577 gnd.n3344 gnd.n3271 99.6594
R7578 gnd.n3345 gnd.n3272 99.6594
R7579 gnd.n3273 gnd.n2709 99.6594
R7580 gnd.n3275 gnd.n3274 99.6594
R7581 gnd.n3276 gnd.n2714 99.6594
R7582 gnd.n3277 gnd.n2720 99.6594
R7583 gnd.n3279 gnd.n2722 99.6594
R7584 gnd.n3396 gnd.n3281 99.6594
R7585 gnd.n3297 gnd.n3265 99.6594
R7586 gnd.n3307 gnd.n3266 99.6594
R7587 gnd.n3318 gnd.n3267 99.6594
R7588 gnd.n3320 gnd.n3268 99.6594
R7589 gnd.n3330 gnd.n3269 99.6594
R7590 gnd.n3343 gnd.n3270 99.6594
R7591 gnd.n3346 gnd.n3271 99.6594
R7592 gnd.n3272 gnd.n2708 99.6594
R7593 gnd.n3273 gnd.n2710 99.6594
R7594 gnd.n3275 gnd.n2713 99.6594
R7595 gnd.n3276 gnd.n2715 99.6594
R7596 gnd.n3277 gnd.n2721 99.6594
R7597 gnd.n3279 gnd.n3278 99.6594
R7598 gnd.n1700 gnd.n1698 99.6594
R7599 gnd.n1715 gnd.n1678 99.6594
R7600 gnd.n1719 gnd.n1717 99.6594
R7601 gnd.n1734 gnd.n1669 99.6594
R7602 gnd.n1738 gnd.n1736 99.6594
R7603 gnd.n1753 gnd.n1660 99.6594
R7604 gnd.n1757 gnd.n1755 99.6594
R7605 gnd.n1772 gnd.n1651 99.6594
R7606 gnd.n1775 gnd.n1774 99.6594
R7607 gnd.n1778 gnd.n1777 99.6594
R7608 gnd.n1783 gnd.n1782 99.6594
R7609 gnd.n1786 gnd.n1785 99.6594
R7610 gnd.n1794 gnd.n1793 99.6594
R7611 gnd.n1797 gnd.n1796 99.6594
R7612 gnd.n1796 gnd.n1795 99.6594
R7613 gnd.n1793 gnd.n1792 99.6594
R7614 gnd.n1785 gnd.n1784 99.6594
R7615 gnd.n1782 gnd.n1781 99.6594
R7616 gnd.n1777 gnd.n1776 99.6594
R7617 gnd.n1774 gnd.n1773 99.6594
R7618 gnd.n1756 gnd.n1651 99.6594
R7619 gnd.n1755 gnd.n1754 99.6594
R7620 gnd.n1737 gnd.n1660 99.6594
R7621 gnd.n1736 gnd.n1735 99.6594
R7622 gnd.n1718 gnd.n1669 99.6594
R7623 gnd.n1717 gnd.n1716 99.6594
R7624 gnd.n1699 gnd.n1678 99.6594
R7625 gnd.n1698 gnd.n1455 99.6594
R7626 gnd.n2716 gnd.t236 98.63
R7627 gnd.n7610 gnd.t260 98.63
R7628 gnd.n1645 gnd.t252 98.63
R7629 gnd.n3339 gnd.t273 98.63
R7630 gnd.n1948 gnd.t229 98.63
R7631 gnd.n1977 gnd.t216 98.63
R7632 gnd.n180 gnd.t279 98.63
R7633 gnd.n7703 gnd.t204 98.63
R7634 gnd.n1031 gnd.t189 98.63
R7635 gnd.n1053 gnd.t271 98.63
R7636 gnd.n2694 gnd.t276 98.63
R7637 gnd.n2605 gnd.t196 98.63
R7638 gnd.n2979 gnd.t222 98.63
R7639 gnd.n1789 gnd.t192 98.63
R7640 gnd.n7385 gnd.n106 94.5225
R7641 gnd.n2465 gnd.t246 92.8196
R7642 gnd.n2032 gnd.t257 92.8196
R7643 gnd.n2462 gnd.t286 92.8118
R7644 gnd.n4228 gnd.t211 92.8118
R7645 gnd.n2414 gnd.n2413 81.8399
R7646 gnd.n5705 gnd.t267 74.8376
R7647 gnd.n5159 gnd.t201 74.8376
R7648 gnd.n2466 gnd.t245 72.8438
R7649 gnd.n2033 gnd.t258 72.8438
R7650 gnd.n2415 gnd.n2408 72.8411
R7651 gnd.n2421 gnd.n2406 72.8411
R7652 gnd.n4224 gnd.n4223 72.8411
R7653 gnd.n2717 gnd.t235 72.836
R7654 gnd.n2463 gnd.t285 72.836
R7655 gnd.n4229 gnd.t212 72.836
R7656 gnd.n7611 gnd.t261 72.836
R7657 gnd.n1646 gnd.t251 72.836
R7658 gnd.n3340 gnd.t274 72.836
R7659 gnd.n1949 gnd.t228 72.836
R7660 gnd.n1978 gnd.t215 72.836
R7661 gnd.n181 gnd.t280 72.836
R7662 gnd.n7704 gnd.t205 72.836
R7663 gnd.n1032 gnd.t188 72.836
R7664 gnd.n1054 gnd.t270 72.836
R7665 gnd.n2695 gnd.t277 72.836
R7666 gnd.n2606 gnd.t197 72.836
R7667 gnd.n2980 gnd.t221 72.836
R7668 gnd.n1790 gnd.t193 72.836
R7669 gnd.n4292 gnd.n1853 71.676
R7670 gnd.n4288 gnd.n1854 71.676
R7671 gnd.n4284 gnd.n1855 71.676
R7672 gnd.n4280 gnd.n1856 71.676
R7673 gnd.n4276 gnd.n1857 71.676
R7674 gnd.n4272 gnd.n1858 71.676
R7675 gnd.n4268 gnd.n1859 71.676
R7676 gnd.n4264 gnd.n1860 71.676
R7677 gnd.n4260 gnd.n1861 71.676
R7678 gnd.n4256 gnd.n1862 71.676
R7679 gnd.n4252 gnd.n1863 71.676
R7680 gnd.n4248 gnd.n1864 71.676
R7681 gnd.n4244 gnd.n1865 71.676
R7682 gnd.n4240 gnd.n1866 71.676
R7683 gnd.n4235 gnd.n1867 71.676
R7684 gnd.n4231 gnd.n1868 71.676
R7685 gnd.n4365 gnd.n1888 71.676
R7686 gnd.n4361 gnd.n1887 71.676
R7687 gnd.n4356 gnd.n1886 71.676
R7688 gnd.n4352 gnd.n1885 71.676
R7689 gnd.n4348 gnd.n1884 71.676
R7690 gnd.n4344 gnd.n1883 71.676
R7691 gnd.n4340 gnd.n1882 71.676
R7692 gnd.n4336 gnd.n1881 71.676
R7693 gnd.n4332 gnd.n1880 71.676
R7694 gnd.n4328 gnd.n1879 71.676
R7695 gnd.n4324 gnd.n1878 71.676
R7696 gnd.n4320 gnd.n1877 71.676
R7697 gnd.n4316 gnd.n1876 71.676
R7698 gnd.n4312 gnd.n1875 71.676
R7699 gnd.n4308 gnd.n1874 71.676
R7700 gnd.n4304 gnd.n1873 71.676
R7701 gnd.n4300 gnd.n1872 71.676
R7702 gnd.n3639 gnd.n3638 71.676
R7703 gnd.n2461 gnd.n2428 71.676
R7704 gnd.n3631 gnd.n2429 71.676
R7705 gnd.n3627 gnd.n2430 71.676
R7706 gnd.n3623 gnd.n2431 71.676
R7707 gnd.n3619 gnd.n2432 71.676
R7708 gnd.n3615 gnd.n2433 71.676
R7709 gnd.n3611 gnd.n2434 71.676
R7710 gnd.n3607 gnd.n2435 71.676
R7711 gnd.n3603 gnd.n2436 71.676
R7712 gnd.n3599 gnd.n2437 71.676
R7713 gnd.n3595 gnd.n2438 71.676
R7714 gnd.n3591 gnd.n2439 71.676
R7715 gnd.n3587 gnd.n2440 71.676
R7716 gnd.n3583 gnd.n2441 71.676
R7717 gnd.n3579 gnd.n2442 71.676
R7718 gnd.n3575 gnd.n2444 71.676
R7719 gnd.n2599 gnd.n2445 71.676
R7720 gnd.n2594 gnd.n2446 71.676
R7721 gnd.n2590 gnd.n2447 71.676
R7722 gnd.n2586 gnd.n2448 71.676
R7723 gnd.n2582 gnd.n2449 71.676
R7724 gnd.n2578 gnd.n2450 71.676
R7725 gnd.n2574 gnd.n2451 71.676
R7726 gnd.n2570 gnd.n2452 71.676
R7727 gnd.n2566 gnd.n2453 71.676
R7728 gnd.n2562 gnd.n2454 71.676
R7729 gnd.n2558 gnd.n2455 71.676
R7730 gnd.n2554 gnd.n2456 71.676
R7731 gnd.n2550 gnd.n2457 71.676
R7732 gnd.n2546 gnd.n2458 71.676
R7733 gnd.n2542 gnd.n2459 71.676
R7734 gnd.n3638 gnd.n2426 71.676
R7735 gnd.n3632 gnd.n2428 71.676
R7736 gnd.n3628 gnd.n2429 71.676
R7737 gnd.n3624 gnd.n2430 71.676
R7738 gnd.n3620 gnd.n2431 71.676
R7739 gnd.n3616 gnd.n2432 71.676
R7740 gnd.n3612 gnd.n2433 71.676
R7741 gnd.n3608 gnd.n2434 71.676
R7742 gnd.n3604 gnd.n2435 71.676
R7743 gnd.n3600 gnd.n2436 71.676
R7744 gnd.n3596 gnd.n2437 71.676
R7745 gnd.n3592 gnd.n2438 71.676
R7746 gnd.n3588 gnd.n2439 71.676
R7747 gnd.n3584 gnd.n2440 71.676
R7748 gnd.n3580 gnd.n2441 71.676
R7749 gnd.n3576 gnd.n2443 71.676
R7750 gnd.n2600 gnd.n2444 71.676
R7751 gnd.n2595 gnd.n2445 71.676
R7752 gnd.n2591 gnd.n2446 71.676
R7753 gnd.n2587 gnd.n2447 71.676
R7754 gnd.n2583 gnd.n2448 71.676
R7755 gnd.n2579 gnd.n2449 71.676
R7756 gnd.n2575 gnd.n2450 71.676
R7757 gnd.n2571 gnd.n2451 71.676
R7758 gnd.n2567 gnd.n2452 71.676
R7759 gnd.n2563 gnd.n2453 71.676
R7760 gnd.n2559 gnd.n2454 71.676
R7761 gnd.n2555 gnd.n2455 71.676
R7762 gnd.n2551 gnd.n2456 71.676
R7763 gnd.n2547 gnd.n2457 71.676
R7764 gnd.n2543 gnd.n2458 71.676
R7765 gnd.n2539 gnd.n2459 71.676
R7766 gnd.n4303 gnd.n1872 71.676
R7767 gnd.n4307 gnd.n1873 71.676
R7768 gnd.n4311 gnd.n1874 71.676
R7769 gnd.n4315 gnd.n1875 71.676
R7770 gnd.n4319 gnd.n1876 71.676
R7771 gnd.n4323 gnd.n1877 71.676
R7772 gnd.n4327 gnd.n1878 71.676
R7773 gnd.n4331 gnd.n1879 71.676
R7774 gnd.n4335 gnd.n1880 71.676
R7775 gnd.n4339 gnd.n1881 71.676
R7776 gnd.n4343 gnd.n1882 71.676
R7777 gnd.n4347 gnd.n1883 71.676
R7778 gnd.n4351 gnd.n1884 71.676
R7779 gnd.n4355 gnd.n1885 71.676
R7780 gnd.n4360 gnd.n1886 71.676
R7781 gnd.n4364 gnd.n1887 71.676
R7782 gnd.n4230 gnd.n1869 71.676
R7783 gnd.n4234 gnd.n1868 71.676
R7784 gnd.n4239 gnd.n1867 71.676
R7785 gnd.n4243 gnd.n1866 71.676
R7786 gnd.n4247 gnd.n1865 71.676
R7787 gnd.n4251 gnd.n1864 71.676
R7788 gnd.n4255 gnd.n1863 71.676
R7789 gnd.n4259 gnd.n1862 71.676
R7790 gnd.n4263 gnd.n1861 71.676
R7791 gnd.n4267 gnd.n1860 71.676
R7792 gnd.n4271 gnd.n1859 71.676
R7793 gnd.n4275 gnd.n1858 71.676
R7794 gnd.n4279 gnd.n1857 71.676
R7795 gnd.n4283 gnd.n1856 71.676
R7796 gnd.n4287 gnd.n1855 71.676
R7797 gnd.n4291 gnd.n1854 71.676
R7798 gnd.n2039 gnd.n1853 71.676
R7799 gnd.n10 gnd.t292 69.1507
R7800 gnd.n18 gnd.t288 68.4792
R7801 gnd.n17 gnd.t6 68.4792
R7802 gnd.n16 gnd.t8 68.4792
R7803 gnd.n15 gnd.t126 68.4792
R7804 gnd.n14 gnd.t324 68.4792
R7805 gnd.n13 gnd.t317 68.4792
R7806 gnd.n12 gnd.t309 68.4792
R7807 gnd.n11 gnd.t63 68.4792
R7808 gnd.n10 gnd.t154 68.4792
R7809 gnd.n5617 gnd.n5518 64.369
R7810 gnd.n2597 gnd.n2466 59.5399
R7811 gnd.n4358 gnd.n2033 59.5399
R7812 gnd.n2464 gnd.n2463 59.5399
R7813 gnd.n4237 gnd.n4229 59.5399
R7814 gnd.n3641 gnd.n2424 59.1804
R7815 gnd.n6487 gnd.n966 57.3586
R7816 gnd.n5135 gnd.n1009 57.3586
R7817 gnd.n5324 gnd.t117 56.607
R7818 gnd.n52 gnd.t168 56.607
R7819 gnd.n5293 gnd.t145 56.407
R7820 gnd.n5308 gnd.t97 56.407
R7821 gnd.n21 gnd.t160 56.407
R7822 gnd.n36 gnd.t73 56.407
R7823 gnd.n5337 gnd.t169 55.8337
R7824 gnd.n5306 gnd.t20 55.8337
R7825 gnd.n5321 gnd.t141 55.8337
R7826 gnd.n65 gnd.t328 55.8337
R7827 gnd.n34 gnd.t102 55.8337
R7828 gnd.n49 gnd.t18 55.8337
R7829 gnd.n2412 gnd.n2411 54.358
R7830 gnd.n4221 gnd.n4220 54.358
R7831 gnd.n5324 gnd.n5323 53.0052
R7832 gnd.n5326 gnd.n5325 53.0052
R7833 gnd.n5328 gnd.n5327 53.0052
R7834 gnd.n5330 gnd.n5329 53.0052
R7835 gnd.n5332 gnd.n5331 53.0052
R7836 gnd.n5334 gnd.n5333 53.0052
R7837 gnd.n5336 gnd.n5335 53.0052
R7838 gnd.n5293 gnd.n5292 53.0052
R7839 gnd.n5295 gnd.n5294 53.0052
R7840 gnd.n5297 gnd.n5296 53.0052
R7841 gnd.n5299 gnd.n5298 53.0052
R7842 gnd.n5301 gnd.n5300 53.0052
R7843 gnd.n5303 gnd.n5302 53.0052
R7844 gnd.n5305 gnd.n5304 53.0052
R7845 gnd.n5308 gnd.n5307 53.0052
R7846 gnd.n5310 gnd.n5309 53.0052
R7847 gnd.n5312 gnd.n5311 53.0052
R7848 gnd.n5314 gnd.n5313 53.0052
R7849 gnd.n5316 gnd.n5315 53.0052
R7850 gnd.n5318 gnd.n5317 53.0052
R7851 gnd.n5320 gnd.n5319 53.0052
R7852 gnd.n64 gnd.n63 53.0052
R7853 gnd.n62 gnd.n61 53.0052
R7854 gnd.n60 gnd.n59 53.0052
R7855 gnd.n58 gnd.n57 53.0052
R7856 gnd.n56 gnd.n55 53.0052
R7857 gnd.n54 gnd.n53 53.0052
R7858 gnd.n52 gnd.n51 53.0052
R7859 gnd.n33 gnd.n32 53.0052
R7860 gnd.n31 gnd.n30 53.0052
R7861 gnd.n29 gnd.n28 53.0052
R7862 gnd.n27 gnd.n26 53.0052
R7863 gnd.n25 gnd.n24 53.0052
R7864 gnd.n23 gnd.n22 53.0052
R7865 gnd.n21 gnd.n20 53.0052
R7866 gnd.n48 gnd.n47 53.0052
R7867 gnd.n46 gnd.n45 53.0052
R7868 gnd.n44 gnd.n43 53.0052
R7869 gnd.n42 gnd.n41 53.0052
R7870 gnd.n40 gnd.n39 53.0052
R7871 gnd.n38 gnd.n37 53.0052
R7872 gnd.n36 gnd.n35 53.0052
R7873 gnd.n4212 gnd.n4211 52.4801
R7874 gnd.n6356 gnd.t150 52.3082
R7875 gnd.n6324 gnd.t319 52.3082
R7876 gnd.n6292 gnd.t71 52.3082
R7877 gnd.n6261 gnd.t83 52.3082
R7878 gnd.n6229 gnd.t106 52.3082
R7879 gnd.n6197 gnd.t111 52.3082
R7880 gnd.n6165 gnd.t87 52.3082
R7881 gnd.n6134 gnd.t307 52.3082
R7882 gnd.n6186 gnd.n6154 51.4173
R7883 gnd.n6250 gnd.n6249 50.455
R7884 gnd.n6218 gnd.n6217 50.455
R7885 gnd.n6186 gnd.n6185 50.455
R7886 gnd.n5555 gnd.n5554 45.1884
R7887 gnd.n5185 gnd.n5184 45.1884
R7888 gnd.n4295 gnd.n4227 44.3322
R7889 gnd.n2415 gnd.n2414 44.3189
R7890 gnd.n7740 gnd.n106 43.6564
R7891 gnd.n2718 gnd.n2717 42.4732
R7892 gnd.n1791 gnd.n1790 42.4732
R7893 gnd.n5567 gnd.n5555 42.2793
R7894 gnd.n5186 gnd.n5185 42.2793
R7895 gnd.n5707 gnd.n5705 42.2793
R7896 gnd.n6459 gnd.n5159 42.2793
R7897 gnd.n7616 gnd.n7611 42.2793
R7898 gnd.n1647 gnd.n1646 42.2793
R7899 gnd.n3341 gnd.n3340 42.2793
R7900 gnd.n1979 gnd.n1978 42.2793
R7901 gnd.n7668 gnd.n181 42.2793
R7902 gnd.n7705 gnd.n7704 42.2793
R7903 gnd.n5099 gnd.n1032 42.2793
R7904 gnd.n1055 gnd.n1054 42.2793
R7905 gnd.n2696 gnd.n2695 42.2793
R7906 gnd.n2981 gnd.n2980 42.2793
R7907 gnd.n2413 gnd.n2412 41.6274
R7908 gnd.n4222 gnd.n4221 41.6274
R7909 gnd.n2422 gnd.n2421 40.8975
R7910 gnd.n4225 gnd.n4224 40.8975
R7911 gnd.n6692 gnd.n740 38.7329
R7912 gnd.n6686 gnd.n740 38.7329
R7913 gnd.n6686 gnd.n6685 38.7329
R7914 gnd.n6685 gnd.n6684 38.7329
R7915 gnd.n6684 gnd.n747 38.7329
R7916 gnd.n6678 gnd.n747 38.7329
R7917 gnd.n6678 gnd.n6677 38.7329
R7918 gnd.n6677 gnd.n6676 38.7329
R7919 gnd.n6676 gnd.n755 38.7329
R7920 gnd.n6670 gnd.n755 38.7329
R7921 gnd.n6670 gnd.n6669 38.7329
R7922 gnd.n6669 gnd.n6668 38.7329
R7923 gnd.n6668 gnd.n763 38.7329
R7924 gnd.n6662 gnd.n763 38.7329
R7925 gnd.n6662 gnd.n6661 38.7329
R7926 gnd.n6661 gnd.n6660 38.7329
R7927 gnd.n6660 gnd.n771 38.7329
R7928 gnd.n6654 gnd.n771 38.7329
R7929 gnd.n6654 gnd.n6653 38.7329
R7930 gnd.n6653 gnd.n6652 38.7329
R7931 gnd.n6652 gnd.n779 38.7329
R7932 gnd.n6646 gnd.n779 38.7329
R7933 gnd.n6646 gnd.n6645 38.7329
R7934 gnd.n6645 gnd.n6644 38.7329
R7935 gnd.n6644 gnd.n787 38.7329
R7936 gnd.n6638 gnd.n787 38.7329
R7937 gnd.n6638 gnd.n6637 38.7329
R7938 gnd.n6637 gnd.n6636 38.7329
R7939 gnd.n6636 gnd.n795 38.7329
R7940 gnd.n6630 gnd.n795 38.7329
R7941 gnd.n6630 gnd.n6629 38.7329
R7942 gnd.n6629 gnd.n6628 38.7329
R7943 gnd.n6628 gnd.n803 38.7329
R7944 gnd.n6622 gnd.n803 38.7329
R7945 gnd.n6622 gnd.n6621 38.7329
R7946 gnd.n6621 gnd.n6620 38.7329
R7947 gnd.n6620 gnd.n811 38.7329
R7948 gnd.n6614 gnd.n811 38.7329
R7949 gnd.n6614 gnd.n6613 38.7329
R7950 gnd.n6613 gnd.n6612 38.7329
R7951 gnd.n6612 gnd.n819 38.7329
R7952 gnd.n6606 gnd.n819 38.7329
R7953 gnd.n6606 gnd.n6605 38.7329
R7954 gnd.n6605 gnd.n6604 38.7329
R7955 gnd.n6604 gnd.n827 38.7329
R7956 gnd.n6598 gnd.n827 38.7329
R7957 gnd.n6598 gnd.n6597 38.7329
R7958 gnd.n6597 gnd.n6596 38.7329
R7959 gnd.n6596 gnd.n835 38.7329
R7960 gnd.n6590 gnd.n835 38.7329
R7961 gnd.n6590 gnd.n6589 38.7329
R7962 gnd.n6589 gnd.n6588 38.7329
R7963 gnd.n6588 gnd.n843 38.7329
R7964 gnd.n6582 gnd.n843 38.7329
R7965 gnd.n6582 gnd.n6581 38.7329
R7966 gnd.n6581 gnd.n6580 38.7329
R7967 gnd.n6580 gnd.n851 38.7329
R7968 gnd.n6574 gnd.n851 38.7329
R7969 gnd.n6574 gnd.n6573 38.7329
R7970 gnd.n6573 gnd.n6572 38.7329
R7971 gnd.n6572 gnd.n859 38.7329
R7972 gnd.n6566 gnd.n859 38.7329
R7973 gnd.n6566 gnd.n6565 38.7329
R7974 gnd.n6565 gnd.n6564 38.7329
R7975 gnd.n6564 gnd.n867 38.7329
R7976 gnd.n6558 gnd.n867 38.7329
R7977 gnd.n6558 gnd.n6557 38.7329
R7978 gnd.n6557 gnd.n6556 38.7329
R7979 gnd.n6556 gnd.n875 38.7329
R7980 gnd.n6550 gnd.n875 38.7329
R7981 gnd.n6550 gnd.n6549 38.7329
R7982 gnd.n6549 gnd.n6548 38.7329
R7983 gnd.n6548 gnd.n883 38.7329
R7984 gnd.n6542 gnd.n883 38.7329
R7985 gnd.n6542 gnd.n6541 38.7329
R7986 gnd.n6541 gnd.n6540 38.7329
R7987 gnd.n6540 gnd.n891 38.7329
R7988 gnd.n6534 gnd.n891 38.7329
R7989 gnd.n6534 gnd.n6533 38.7329
R7990 gnd.n6533 gnd.n6532 38.7329
R7991 gnd.n6532 gnd.n899 38.7329
R7992 gnd.n6526 gnd.n899 38.7329
R7993 gnd.n6526 gnd.n6525 38.7329
R7994 gnd.n2030 gnd.n1949 36.9518
R7995 gnd.n3573 gnd.n2606 36.9518
R7996 gnd.n2421 gnd.n2420 35.055
R7997 gnd.n2416 gnd.n2415 35.055
R7998 gnd.n4214 gnd.n4213 35.055
R7999 gnd.n4224 gnd.n4210 35.055
R8000 gnd.n5617 gnd.n5513 31.8661
R8001 gnd.n5625 gnd.n5513 31.8661
R8002 gnd.n5633 gnd.n5507 31.8661
R8003 gnd.n5633 gnd.n5501 31.8661
R8004 gnd.n5641 gnd.n5501 31.8661
R8005 gnd.n5641 gnd.n5494 31.8661
R8006 gnd.n5649 gnd.n5494 31.8661
R8007 gnd.n5649 gnd.n5495 31.8661
R8008 gnd.n5748 gnd.n5480 31.8661
R8009 gnd.n3038 gnd.n1009 31.8661
R8010 gnd.n5048 gnd.n1063 31.8661
R8011 gnd.n5048 gnd.n1065 31.8661
R8012 gnd.n5042 gnd.n1065 31.8661
R8013 gnd.n5042 gnd.n1077 31.8661
R8014 gnd.n5036 gnd.n1088 31.8661
R8015 gnd.n5030 gnd.n1088 31.8661
R8016 gnd.n5024 gnd.n1105 31.8661
R8017 gnd.n3264 gnd.n3263 31.8661
R8018 gnd.n3398 gnd.n3264 31.8661
R8019 gnd.n3406 gnd.n2775 31.8661
R8020 gnd.n4736 gnd.n1458 31.8661
R8021 gnd.n4730 gnd.n4729 31.8661
R8022 gnd.n4729 gnd.n4728 31.8661
R8023 gnd.n7553 gnd.n218 31.8661
R8024 gnd.n7561 gnd.n208 31.8661
R8025 gnd.n7561 gnd.n211 31.8661
R8026 gnd.n7569 gnd.n193 31.8661
R8027 gnd.n7652 gnd.n193 31.8661
R8028 gnd.n7652 gnd.n186 31.8661
R8029 gnd.n7660 gnd.n186 31.8661
R8030 gnd.n7740 gnd.n104 31.8661
R8031 gnd.n4301 gnd.n2034 31.3761
R8032 gnd.n2540 gnd.n2537 31.3761
R8033 gnd.n3079 gnd.n1116 29.3168
R8034 gnd.n5018 gnd.n1119 29.3168
R8035 gnd.n5012 gnd.n1130 29.3168
R8036 gnd.n3095 gnd.n1138 29.3168
R8037 gnd.n3103 gnd.n1148 29.3168
R8038 gnd.n3111 gnd.n1158 29.3168
R8039 gnd.n4994 gnd.n1161 29.3168
R8040 gnd.n4988 gnd.n1172 29.3168
R8041 gnd.n3127 gnd.n1178 29.3168
R8042 gnd.n3136 gnd.n1188 29.3168
R8043 gnd.n3145 gnd.n1195 29.3168
R8044 gnd.n4969 gnd.n1198 29.3168
R8045 gnd.n4963 gnd.n1209 29.3168
R8046 gnd.n3161 gnd.n1216 29.3168
R8047 gnd.n3169 gnd.n1226 29.3168
R8048 gnd.n3177 gnd.n1236 29.3168
R8049 gnd.n4945 gnd.n1239 29.3168
R8050 gnd.n4939 gnd.n1250 29.3168
R8051 gnd.n3194 gnd.n1258 29.3168
R8052 gnd.n3202 gnd.n1268 29.3168
R8053 gnd.n3237 gnd.n1278 29.3168
R8054 gnd.n4921 gnd.n1281 29.3168
R8055 gnd.n4915 gnd.n1292 29.3168
R8056 gnd.n3214 gnd.n1300 29.3168
R8057 gnd.n4909 gnd.n1303 29.3168
R8058 gnd.n3223 gnd.n1311 29.3168
R8059 gnd.n3528 gnd.n1320 29.3168
R8060 gnd.n4897 gnd.n1323 29.3168
R8061 gnd.n1477 gnd.n1476 29.3168
R8062 gnd.n4722 gnd.n4721 29.3168
R8063 gnd.n4715 gnd.n1490 29.3168
R8064 gnd.n1635 gnd.n1493 29.3168
R8065 gnd.n4525 gnd.n1634 29.3168
R8066 gnd.n4517 gnd.n1616 29.3168
R8067 gnd.n4547 gnd.n1605 29.3168
R8068 gnd.n4545 gnd.n1608 29.3168
R8069 gnd.n1598 gnd.n1589 29.3168
R8070 gnd.n4586 gnd.n1578 29.3168
R8071 gnd.n4585 gnd.n1581 29.3168
R8072 gnd.n1572 gnd.n1569 29.3168
R8073 gnd.n4609 gnd.n1561 29.3168
R8074 gnd.n4675 gnd.n1528 29.3168
R8075 gnd.n4622 gnd.n1520 29.3168
R8076 gnd.n7498 gnd.n277 29.3168
R8077 gnd.n4633 gnd.n1541 29.3168
R8078 gnd.n4662 gnd.n4661 29.3168
R8079 gnd.n4656 gnd.n4645 29.3168
R8080 gnd.n7482 gnd.n294 29.3168
R8081 gnd.n7471 gnd.n296 29.3168
R8082 gnd.n7403 gnd.n264 29.3168
R8083 gnd.n7513 gnd.n255 29.3168
R8084 gnd.n7521 gnd.n247 29.3168
R8085 gnd.n7529 gnd.n239 29.3168
R8086 gnd.n7454 gnd.n241 29.3168
R8087 gnd.n7447 gnd.n233 29.3168
R8088 gnd.n7545 gnd.n225 29.3168
R8089 gnd.n2666 gnd.n1323 28.0422
R8090 gnd.n1476 gnd.n1468 28.0422
R8091 gnd.n5000 gnd.t31 27.0862
R8092 gnd.n7410 gnd.t11 27.0862
R8093 gnd.n4976 gnd.t15 26.4489
R8094 gnd.n4657 gnd.t60 26.4489
R8095 gnd.n4951 gnd.t98 25.8116
R8096 gnd.n4676 gnd.t3 25.8116
R8097 gnd.n2717 gnd.n2716 25.7944
R8098 gnd.n5705 gnd.n5704 25.7944
R8099 gnd.n5159 gnd.n5158 25.7944
R8100 gnd.n7611 gnd.n7610 25.7944
R8101 gnd.n1646 gnd.n1645 25.7944
R8102 gnd.n3340 gnd.n3339 25.7944
R8103 gnd.n1949 gnd.n1948 25.7944
R8104 gnd.n1978 gnd.n1977 25.7944
R8105 gnd.n181 gnd.n180 25.7944
R8106 gnd.n7704 gnd.n7703 25.7944
R8107 gnd.n1032 gnd.n1031 25.7944
R8108 gnd.n1054 gnd.n1053 25.7944
R8109 gnd.n2695 gnd.n2694 25.7944
R8110 gnd.n2606 gnd.n2605 25.7944
R8111 gnd.n2980 gnd.n2979 25.7944
R8112 gnd.n1790 gnd.n1789 25.7944
R8113 gnd.n1105 gnd.t58 25.1743
R8114 gnd.n2808 gnd.t76 25.1743
R8115 gnd.n4927 gnd.t51 25.1743
R8116 gnd.n4557 gnd.t127 25.1743
R8117 gnd.n4568 gnd.t131 25.1743
R8118 gnd.n7553 gnd.t121 25.1743
R8119 gnd.n5749 gnd.n5469 24.8557
R8120 gnd.n5472 gnd.n5463 24.8557
R8121 gnd.n5770 gnd.n5448 24.8557
R8122 gnd.n5789 gnd.n5788 24.8557
R8123 gnd.n5799 gnd.n5441 24.8557
R8124 gnd.n5812 gnd.n5429 24.8557
R8125 gnd.n5837 gnd.n5413 24.8557
R8126 gnd.n5836 gnd.n5415 24.8557
R8127 gnd.n5859 gnd.n5397 24.8557
R8128 gnd.n5848 gnd.n5389 24.8557
R8129 gnd.n5884 gnd.n5883 24.8557
R8130 gnd.n5894 gnd.n5382 24.8557
R8131 gnd.n5906 gnd.n5374 24.8557
R8132 gnd.n5905 gnd.n5362 24.8557
R8133 gnd.n5924 gnd.n5923 24.8557
R8134 gnd.n5945 gnd.n5343 24.8557
R8135 gnd.n5969 gnd.n5968 24.8557
R8136 gnd.n5980 gnd.n5278 24.8557
R8137 gnd.n5979 gnd.n5280 24.8557
R8138 gnd.n5991 gnd.n5271 24.8557
R8139 gnd.n6008 gnd.n6007 24.8557
R8140 gnd.n5262 gnd.n5251 24.8557
R8141 gnd.n6031 gnd.n5240 24.8557
R8142 gnd.n5242 gnd.n5241 24.8557
R8143 gnd.n6051 gnd.n5234 24.8557
R8144 gnd.n6063 gnd.n6062 24.8557
R8145 gnd.n6074 gnd.n5221 24.8557
R8146 gnd.n6087 gnd.n5211 24.8557
R8147 gnd.n6523 gnd.n909 24.8557
R8148 gnd.n6517 gnd.n6516 24.8557
R8149 gnd.n6116 gnd.n920 24.8557
R8150 gnd.n6509 gnd.n931 24.8557
R8151 gnd.n5195 gnd.n942 24.8557
R8152 gnd.n6503 gnd.n6502 24.8557
R8153 gnd.n6495 gnd.n956 24.8557
R8154 gnd.n2822 gnd.t94 24.537
R8155 gnd.n1530 gnd.t118 24.537
R8156 gnd.n2837 gnd.t53 23.8997
R8157 gnd.n3398 gnd.n3397 23.8997
R8158 gnd.n4730 gnd.n1467 23.8997
R8159 gnd.n4646 gnd.t27 23.8997
R8160 gnd.n5767 gnd.t306 23.2624
R8161 gnd.n2943 gnd.t21 23.2624
R8162 gnd.t23 gnd.n249 23.2624
R8163 gnd.n6525 gnd.n6524 23.2399
R8164 gnd.n5759 gnd.t266 22.6251
R8165 gnd.n3038 gnd.t187 22.6251
R8166 gnd.t203 gnd.n104 22.6251
R8167 gnd.t45 gnd.n1108 21.6691
R8168 gnd.n7393 gnd.t35 21.6691
R8169 gnd.n5739 gnd.t82 21.3504
R8170 gnd.t136 gnd.n907 20.7131
R8171 gnd.t312 gnd.n5252 20.0758
R8172 gnd.n2701 gnd.t195 20.0758
R8173 gnd.t214 gnd.n1480 20.0758
R8174 gnd.n2466 gnd.n2465 19.9763
R8175 gnd.n2033 gnd.n2032 19.9763
R8176 gnd.n2463 gnd.n2462 19.9763
R8177 gnd.n4229 gnd.n4228 19.9763
R8178 gnd.n2409 gnd.t239 19.8005
R8179 gnd.n2409 gnd.t249 19.8005
R8180 gnd.n2410 gnd.t219 19.8005
R8181 gnd.n2410 gnd.t255 19.8005
R8182 gnd.n4218 gnd.t242 19.8005
R8183 gnd.n4218 gnd.t232 19.8005
R8184 gnd.n4219 gnd.t181 19.8005
R8185 gnd.n4219 gnd.t283 19.8005
R8186 gnd.n2406 gnd.n2405 19.5087
R8187 gnd.n2419 gnd.n2406 19.5087
R8188 gnd.n2417 gnd.n2408 19.5087
R8189 gnd.n4223 gnd.n4217 19.5087
R8190 gnd.t65 gnd.n5287 19.4385
R8191 gnd.n3504 gnd.n3503 19.3944
R8192 gnd.n3503 gnd.n3502 19.3944
R8193 gnd.n3502 gnd.n2728 19.3944
R8194 gnd.n3498 gnd.n2728 19.3944
R8195 gnd.n3498 gnd.n3497 19.3944
R8196 gnd.n3497 gnd.n3496 19.3944
R8197 gnd.n3496 gnd.n2733 19.3944
R8198 gnd.n3492 gnd.n2733 19.3944
R8199 gnd.n3492 gnd.n3491 19.3944
R8200 gnd.n3491 gnd.n3490 19.3944
R8201 gnd.n3490 gnd.n2738 19.3944
R8202 gnd.n3486 gnd.n2738 19.3944
R8203 gnd.n3486 gnd.n3485 19.3944
R8204 gnd.n3485 gnd.n3484 19.3944
R8205 gnd.n3484 gnd.n2743 19.3944
R8206 gnd.n3480 gnd.n2743 19.3944
R8207 gnd.n3480 gnd.n3479 19.3944
R8208 gnd.n3479 gnd.n3478 19.3944
R8209 gnd.n3478 gnd.n3475 19.3944
R8210 gnd.n3475 gnd.n2384 19.3944
R8211 gnd.n3666 gnd.n2384 19.3944
R8212 gnd.n3666 gnd.n2382 19.3944
R8213 gnd.n3670 gnd.n2382 19.3944
R8214 gnd.n3670 gnd.n2364 19.3944
R8215 gnd.n3696 gnd.n2364 19.3944
R8216 gnd.n3696 gnd.n2361 19.3944
R8217 gnd.n3701 gnd.n2361 19.3944
R8218 gnd.n3701 gnd.n2362 19.3944
R8219 gnd.n2362 gnd.n2337 19.3944
R8220 gnd.n3733 gnd.n2337 19.3944
R8221 gnd.n3733 gnd.n2335 19.3944
R8222 gnd.n3737 gnd.n2335 19.3944
R8223 gnd.n3737 gnd.n2317 19.3944
R8224 gnd.n3760 gnd.n2317 19.3944
R8225 gnd.n3760 gnd.n2314 19.3944
R8226 gnd.n3765 gnd.n2314 19.3944
R8227 gnd.n3765 gnd.n2315 19.3944
R8228 gnd.n2315 gnd.n2287 19.3944
R8229 gnd.n3799 gnd.n2287 19.3944
R8230 gnd.n3799 gnd.n2284 19.3944
R8231 gnd.n3817 gnd.n2284 19.3944
R8232 gnd.n3817 gnd.n2285 19.3944
R8233 gnd.n3813 gnd.n2285 19.3944
R8234 gnd.n3813 gnd.n3812 19.3944
R8235 gnd.n3812 gnd.n3811 19.3944
R8236 gnd.n3811 gnd.n3808 19.3944
R8237 gnd.n3808 gnd.n2225 19.3944
R8238 gnd.n3881 gnd.n2225 19.3944
R8239 gnd.n3881 gnd.n2222 19.3944
R8240 gnd.n3886 gnd.n2222 19.3944
R8241 gnd.n3886 gnd.n2223 19.3944
R8242 gnd.n2223 gnd.n2195 19.3944
R8243 gnd.n3917 gnd.n2195 19.3944
R8244 gnd.n3917 gnd.n2192 19.3944
R8245 gnd.n3934 gnd.n2192 19.3944
R8246 gnd.n3934 gnd.n2193 19.3944
R8247 gnd.n3930 gnd.n2193 19.3944
R8248 gnd.n3930 gnd.n3929 19.3944
R8249 gnd.n3929 gnd.n3928 19.3944
R8250 gnd.n3928 gnd.n3925 19.3944
R8251 gnd.n3925 gnd.n2146 19.3944
R8252 gnd.n4011 gnd.n2146 19.3944
R8253 gnd.n4011 gnd.n2143 19.3944
R8254 gnd.n4030 gnd.n2143 19.3944
R8255 gnd.n4030 gnd.n2144 19.3944
R8256 gnd.n4026 gnd.n2144 19.3944
R8257 gnd.n4026 gnd.n4025 19.3944
R8258 gnd.n4025 gnd.n4024 19.3944
R8259 gnd.n4024 gnd.n4021 19.3944
R8260 gnd.n4021 gnd.n2097 19.3944
R8261 gnd.n4100 gnd.n2097 19.3944
R8262 gnd.n4100 gnd.n2094 19.3944
R8263 gnd.n4108 gnd.n2094 19.3944
R8264 gnd.n4108 gnd.n2095 19.3944
R8265 gnd.n4104 gnd.n2095 19.3944
R8266 gnd.n4104 gnd.n2066 19.3944
R8267 gnd.n4168 gnd.n2066 19.3944
R8268 gnd.n4168 gnd.n2063 19.3944
R8269 gnd.n4179 gnd.n2063 19.3944
R8270 gnd.n4179 gnd.n2064 19.3944
R8271 gnd.n4175 gnd.n2064 19.3944
R8272 gnd.n4175 gnd.n4174 19.3944
R8273 gnd.n4174 gnd.n1850 19.3944
R8274 gnd.n4369 gnd.n1850 19.3944
R8275 gnd.n4369 gnd.n1848 19.3944
R8276 gnd.n4373 gnd.n1848 19.3944
R8277 gnd.n4373 gnd.n1838 19.3944
R8278 gnd.n4389 gnd.n1838 19.3944
R8279 gnd.n4389 gnd.n1836 19.3944
R8280 gnd.n4393 gnd.n1836 19.3944
R8281 gnd.n4393 gnd.n1825 19.3944
R8282 gnd.n4409 gnd.n1825 19.3944
R8283 gnd.n4409 gnd.n1823 19.3944
R8284 gnd.n4413 gnd.n1823 19.3944
R8285 gnd.n4413 gnd.n1812 19.3944
R8286 gnd.n4429 gnd.n1812 19.3944
R8287 gnd.n4429 gnd.n1810 19.3944
R8288 gnd.n4434 gnd.n1810 19.3944
R8289 gnd.n4434 gnd.n1801 19.3944
R8290 gnd.n4452 gnd.n1801 19.3944
R8291 gnd.n4453 gnd.n4452 19.3944
R8292 gnd.n3510 gnd.n3509 19.3944
R8293 gnd.n3509 gnd.n3508 19.3944
R8294 gnd.n3508 gnd.n2723 19.3944
R8295 gnd.n3394 gnd.n3393 19.3944
R8296 gnd.n3393 gnd.n3283 19.3944
R8297 gnd.n3386 gnd.n3283 19.3944
R8298 gnd.n3386 gnd.n3385 19.3944
R8299 gnd.n3385 gnd.n3299 19.3944
R8300 gnd.n3378 gnd.n3299 19.3944
R8301 gnd.n3378 gnd.n3377 19.3944
R8302 gnd.n3377 gnd.n3309 19.3944
R8303 gnd.n3370 gnd.n3309 19.3944
R8304 gnd.n3370 gnd.n3369 19.3944
R8305 gnd.n3369 gnd.n3322 19.3944
R8306 gnd.n3362 gnd.n3322 19.3944
R8307 gnd.n3362 gnd.n3361 19.3944
R8308 gnd.n3361 gnd.n3332 19.3944
R8309 gnd.n3354 gnd.n3332 19.3944
R8310 gnd.n3354 gnd.n3353 19.3944
R8311 gnd.n3353 gnd.n2707 19.3944
R8312 gnd.n3521 gnd.n2707 19.3944
R8313 gnd.n3521 gnd.n3520 19.3944
R8314 gnd.n3520 gnd.n3519 19.3944
R8315 gnd.n3519 gnd.n2711 19.3944
R8316 gnd.n3515 gnd.n2711 19.3944
R8317 gnd.n3515 gnd.n3514 19.3944
R8318 gnd.n3514 gnd.n3513 19.3944
R8319 gnd.n5612 gnd.n5611 19.3944
R8320 gnd.n5611 gnd.n5521 19.3944
R8321 gnd.n5606 gnd.n5521 19.3944
R8322 gnd.n5606 gnd.n5605 19.3944
R8323 gnd.n5605 gnd.n5526 19.3944
R8324 gnd.n5600 gnd.n5526 19.3944
R8325 gnd.n5600 gnd.n5599 19.3944
R8326 gnd.n5599 gnd.n5598 19.3944
R8327 gnd.n5598 gnd.n5532 19.3944
R8328 gnd.n5592 gnd.n5532 19.3944
R8329 gnd.n5592 gnd.n5591 19.3944
R8330 gnd.n5591 gnd.n5590 19.3944
R8331 gnd.n5590 gnd.n5538 19.3944
R8332 gnd.n5584 gnd.n5538 19.3944
R8333 gnd.n5584 gnd.n5583 19.3944
R8334 gnd.n5583 gnd.n5582 19.3944
R8335 gnd.n5582 gnd.n5544 19.3944
R8336 gnd.n5576 gnd.n5544 19.3944
R8337 gnd.n5576 gnd.n5575 19.3944
R8338 gnd.n5575 gnd.n5574 19.3944
R8339 gnd.n5574 gnd.n5550 19.3944
R8340 gnd.n5568 gnd.n5550 19.3944
R8341 gnd.n5566 gnd.n5565 19.3944
R8342 gnd.n5565 gnd.n5560 19.3944
R8343 gnd.n5560 gnd.n5558 19.3944
R8344 gnd.n6409 gnd.n6408 19.3944
R8345 gnd.n6408 gnd.n6405 19.3944
R8346 gnd.n6405 gnd.n6404 19.3944
R8347 gnd.n6454 gnd.n6453 19.3944
R8348 gnd.n6453 gnd.n6452 19.3944
R8349 gnd.n6452 gnd.n6449 19.3944
R8350 gnd.n6449 gnd.n6448 19.3944
R8351 gnd.n6448 gnd.n6445 19.3944
R8352 gnd.n6445 gnd.n6444 19.3944
R8353 gnd.n6444 gnd.n6441 19.3944
R8354 gnd.n6441 gnd.n6440 19.3944
R8355 gnd.n6440 gnd.n6437 19.3944
R8356 gnd.n6437 gnd.n6436 19.3944
R8357 gnd.n6436 gnd.n6433 19.3944
R8358 gnd.n6433 gnd.n6432 19.3944
R8359 gnd.n6432 gnd.n6429 19.3944
R8360 gnd.n6429 gnd.n6428 19.3944
R8361 gnd.n6428 gnd.n6425 19.3944
R8362 gnd.n6425 gnd.n6424 19.3944
R8363 gnd.n6424 gnd.n6421 19.3944
R8364 gnd.n6421 gnd.n6420 19.3944
R8365 gnd.n6420 gnd.n6417 19.3944
R8366 gnd.n6417 gnd.n6416 19.3944
R8367 gnd.n6416 gnd.n6413 19.3944
R8368 gnd.n6413 gnd.n6412 19.3944
R8369 gnd.n5752 gnd.n5751 19.3944
R8370 gnd.n5753 gnd.n5752 19.3944
R8371 gnd.n5753 gnd.n5462 19.3944
R8372 gnd.n5462 gnd.n5456 19.3944
R8373 gnd.n5778 gnd.n5456 19.3944
R8374 gnd.n5779 gnd.n5778 19.3944
R8375 gnd.n5779 gnd.n5439 19.3944
R8376 gnd.n5439 gnd.n5437 19.3944
R8377 gnd.n5803 gnd.n5437 19.3944
R8378 gnd.n5806 gnd.n5803 19.3944
R8379 gnd.n5806 gnd.n5805 19.3944
R8380 gnd.n5805 gnd.n5409 19.3944
R8381 gnd.n5844 gnd.n5409 19.3944
R8382 gnd.n5844 gnd.n5407 19.3944
R8383 gnd.n5850 gnd.n5407 19.3944
R8384 gnd.n5851 gnd.n5850 19.3944
R8385 gnd.n5851 gnd.n5377 19.3944
R8386 gnd.n5901 gnd.n5377 19.3944
R8387 gnd.n5902 gnd.n5901 19.3944
R8388 gnd.n5902 gnd.n5370 19.3944
R8389 gnd.n5913 gnd.n5370 19.3944
R8390 gnd.n5914 gnd.n5913 19.3944
R8391 gnd.n5914 gnd.n5353 19.3944
R8392 gnd.n5353 gnd.n5351 19.3944
R8393 gnd.n5938 gnd.n5351 19.3944
R8394 gnd.n5939 gnd.n5938 19.3944
R8395 gnd.n5939 gnd.n5274 19.3944
R8396 gnd.n5986 gnd.n5274 19.3944
R8397 gnd.n5987 gnd.n5986 19.3944
R8398 gnd.n5987 gnd.n5267 19.3944
R8399 gnd.n5998 gnd.n5267 19.3944
R8400 gnd.n5999 gnd.n5998 19.3944
R8401 gnd.n5999 gnd.n5250 19.3944
R8402 gnd.n5250 gnd.n5247 19.3944
R8403 gnd.n6026 gnd.n5247 19.3944
R8404 gnd.n6026 gnd.n5248 19.3944
R8405 gnd.n5248 gnd.n5230 19.3944
R8406 gnd.n6059 gnd.n5230 19.3944
R8407 gnd.n6059 gnd.n6058 19.3944
R8408 gnd.n6058 gnd.n5214 19.3944
R8409 gnd.n6084 gnd.n5214 19.3944
R8410 gnd.n6084 gnd.n5206 19.3944
R8411 gnd.n6097 gnd.n5206 19.3944
R8412 gnd.n6097 gnd.n6096 19.3944
R8413 gnd.n6096 gnd.n5199 19.3944
R8414 gnd.n6119 gnd.n5199 19.3944
R8415 gnd.n6120 gnd.n6119 19.3944
R8416 gnd.n6120 gnd.n5197 19.3944
R8417 gnd.n6382 gnd.n5197 19.3944
R8418 gnd.n6384 gnd.n6382 19.3944
R8419 gnd.n6392 gnd.n6384 19.3944
R8420 gnd.n6392 gnd.n6391 19.3944
R8421 gnd.n6391 gnd.n6390 19.3944
R8422 gnd.n5735 gnd.n5734 19.3944
R8423 gnd.n5734 gnd.n5733 19.3944
R8424 gnd.n5733 gnd.n5732 19.3944
R8425 gnd.n5732 gnd.n5730 19.3944
R8426 gnd.n5730 gnd.n5727 19.3944
R8427 gnd.n5727 gnd.n5726 19.3944
R8428 gnd.n5726 gnd.n5723 19.3944
R8429 gnd.n5723 gnd.n5722 19.3944
R8430 gnd.n5722 gnd.n5719 19.3944
R8431 gnd.n5719 gnd.n5718 19.3944
R8432 gnd.n5718 gnd.n5715 19.3944
R8433 gnd.n5715 gnd.n5714 19.3944
R8434 gnd.n5714 gnd.n5711 19.3944
R8435 gnd.n5711 gnd.n5710 19.3944
R8436 gnd.n5761 gnd.n5467 19.3944
R8437 gnd.n5761 gnd.n5465 19.3944
R8438 gnd.n5765 gnd.n5465 19.3944
R8439 gnd.n5765 gnd.n5446 19.3944
R8440 gnd.n5791 gnd.n5446 19.3944
R8441 gnd.n5791 gnd.n5444 19.3944
R8442 gnd.n5797 gnd.n5444 19.3944
R8443 gnd.n5797 gnd.n5796 19.3944
R8444 gnd.n5796 gnd.n5420 19.3944
R8445 gnd.n5825 gnd.n5420 19.3944
R8446 gnd.n5825 gnd.n5418 19.3944
R8447 gnd.n5834 gnd.n5418 19.3944
R8448 gnd.n5834 gnd.n5833 19.3944
R8449 gnd.n5833 gnd.n5832 19.3944
R8450 gnd.n5832 gnd.n5387 19.3944
R8451 gnd.n5886 gnd.n5387 19.3944
R8452 gnd.n5886 gnd.n5385 19.3944
R8453 gnd.n5892 gnd.n5385 19.3944
R8454 gnd.n5892 gnd.n5891 19.3944
R8455 gnd.n5891 gnd.n5360 19.3944
R8456 gnd.n5926 gnd.n5360 19.3944
R8457 gnd.n5926 gnd.n5358 19.3944
R8458 gnd.n5932 gnd.n5358 19.3944
R8459 gnd.n5932 gnd.n5931 19.3944
R8460 gnd.n5931 gnd.n5285 19.3944
R8461 gnd.n5971 gnd.n5285 19.3944
R8462 gnd.n5971 gnd.n5283 19.3944
R8463 gnd.n5977 gnd.n5283 19.3944
R8464 gnd.n5977 gnd.n5976 19.3944
R8465 gnd.n5976 gnd.n5257 19.3944
R8466 gnd.n6010 gnd.n5257 19.3944
R8467 gnd.n6010 gnd.n5255 19.3944
R8468 gnd.n6019 gnd.n5255 19.3944
R8469 gnd.n6019 gnd.n6018 19.3944
R8470 gnd.n6018 gnd.n6017 19.3944
R8471 gnd.n6017 gnd.n5226 19.3944
R8472 gnd.n6065 gnd.n5226 19.3944
R8473 gnd.n6065 gnd.n5224 19.3944
R8474 gnd.n6072 gnd.n5224 19.3944
R8475 gnd.n6072 gnd.n6071 19.3944
R8476 gnd.n6071 gnd.n912 19.3944
R8477 gnd.n6521 gnd.n912 19.3944
R8478 gnd.n6521 gnd.n6520 19.3944
R8479 gnd.n6520 gnd.n6519 19.3944
R8480 gnd.n6519 gnd.n916 19.3944
R8481 gnd.n934 gnd.n916 19.3944
R8482 gnd.n6507 gnd.n934 19.3944
R8483 gnd.n6507 gnd.n6506 19.3944
R8484 gnd.n6506 gnd.n6505 19.3944
R8485 gnd.n6505 gnd.n940 19.3944
R8486 gnd.n959 gnd.n940 19.3944
R8487 gnd.n6493 gnd.n959 19.3944
R8488 gnd.n6493 gnd.n6492 19.3944
R8489 gnd.n6489 gnd.n964 19.3944
R8490 gnd.n6484 gnd.n964 19.3944
R8491 gnd.n6484 gnd.n6483 19.3944
R8492 gnd.n6483 gnd.n6482 19.3944
R8493 gnd.n6482 gnd.n6479 19.3944
R8494 gnd.n6479 gnd.n6478 19.3944
R8495 gnd.n6478 gnd.n6475 19.3944
R8496 gnd.n6475 gnd.n6474 19.3944
R8497 gnd.n6474 gnd.n6471 19.3944
R8498 gnd.n6471 gnd.n6470 19.3944
R8499 gnd.n6470 gnd.n6467 19.3944
R8500 gnd.n6467 gnd.n6466 19.3944
R8501 gnd.n6466 gnd.n6463 19.3944
R8502 gnd.n6463 gnd.n6462 19.3944
R8503 gnd.n5619 gnd.n5515 19.3944
R8504 gnd.n5623 gnd.n5515 19.3944
R8505 gnd.n5623 gnd.n5505 19.3944
R8506 gnd.n5635 gnd.n5505 19.3944
R8507 gnd.n5635 gnd.n5503 19.3944
R8508 gnd.n5639 gnd.n5503 19.3944
R8509 gnd.n5639 gnd.n5492 19.3944
R8510 gnd.n5651 gnd.n5492 19.3944
R8511 gnd.n5651 gnd.n5490 19.3944
R8512 gnd.n5677 gnd.n5490 19.3944
R8513 gnd.n5677 gnd.n5676 19.3944
R8514 gnd.n5676 gnd.n5675 19.3944
R8515 gnd.n5675 gnd.n5674 19.3944
R8516 gnd.n5674 gnd.n5672 19.3944
R8517 gnd.n5672 gnd.n5671 19.3944
R8518 gnd.n5671 gnd.n5669 19.3944
R8519 gnd.n5669 gnd.n5668 19.3944
R8520 gnd.n5668 gnd.n5666 19.3944
R8521 gnd.n5666 gnd.n5665 19.3944
R8522 gnd.n5665 gnd.n5427 19.3944
R8523 gnd.n5814 gnd.n5427 19.3944
R8524 gnd.n5814 gnd.n5425 19.3944
R8525 gnd.n5820 gnd.n5425 19.3944
R8526 gnd.n5820 gnd.n5819 19.3944
R8527 gnd.n5819 gnd.n5394 19.3944
R8528 gnd.n5861 gnd.n5394 19.3944
R8529 gnd.n5861 gnd.n5392 19.3944
R8530 gnd.n5865 gnd.n5392 19.3944
R8531 gnd.n5879 gnd.n5865 19.3944
R8532 gnd.n5877 gnd.n5876 19.3944
R8533 gnd.n5873 gnd.n5872 19.3944
R8534 gnd.n5869 gnd.n5868 19.3944
R8535 gnd.n5947 gnd.n5341 19.3944
R8536 gnd.n5947 gnd.n5291 19.3944
R8537 gnd.n5966 gnd.n5291 19.3944
R8538 gnd.n5966 gnd.n5965 19.3944
R8539 gnd.n5965 gnd.n5964 19.3944
R8540 gnd.n5964 gnd.n5962 19.3944
R8541 gnd.n5962 gnd.n5961 19.3944
R8542 gnd.n5961 gnd.n5959 19.3944
R8543 gnd.n5959 gnd.n5958 19.3944
R8544 gnd.n5958 gnd.n5238 19.3944
R8545 gnd.n6033 gnd.n5238 19.3944
R8546 gnd.n6033 gnd.n5236 19.3944
R8547 gnd.n6049 gnd.n5236 19.3944
R8548 gnd.n6049 gnd.n6048 19.3944
R8549 gnd.n6048 gnd.n6047 19.3944
R8550 gnd.n6047 gnd.n6046 19.3944
R8551 gnd.n6046 gnd.n6044 19.3944
R8552 gnd.n6044 gnd.n6043 19.3944
R8553 gnd.n6043 gnd.n5204 19.3944
R8554 gnd.n6102 gnd.n5204 19.3944
R8555 gnd.n6102 gnd.n5202 19.3944
R8556 gnd.n6114 gnd.n5202 19.3944
R8557 gnd.n6114 gnd.n6113 19.3944
R8558 gnd.n6113 gnd.n6112 19.3944
R8559 gnd.n6112 gnd.n6109 19.3944
R8560 gnd.n6109 gnd.n5193 19.3944
R8561 gnd.n6397 gnd.n5193 19.3944
R8562 gnd.n6397 gnd.n5191 19.3944
R8563 gnd.n6401 gnd.n5191 19.3944
R8564 gnd.n5615 gnd.n5511 19.3944
R8565 gnd.n5627 gnd.n5511 19.3944
R8566 gnd.n5627 gnd.n5509 19.3944
R8567 gnd.n5631 gnd.n5509 19.3944
R8568 gnd.n5631 gnd.n5499 19.3944
R8569 gnd.n5643 gnd.n5499 19.3944
R8570 gnd.n5643 gnd.n5497 19.3944
R8571 gnd.n5647 gnd.n5497 19.3944
R8572 gnd.n5647 gnd.n5486 19.3944
R8573 gnd.n5741 gnd.n5486 19.3944
R8574 gnd.n5741 gnd.n5483 19.3944
R8575 gnd.n5746 gnd.n5483 19.3944
R8576 gnd.n5746 gnd.n5474 19.3944
R8577 gnd.n5756 gnd.n5474 19.3944
R8578 gnd.n5756 gnd.n5458 19.3944
R8579 gnd.n5773 gnd.n5458 19.3944
R8580 gnd.n5773 gnd.n5454 19.3944
R8581 gnd.n5786 gnd.n5454 19.3944
R8582 gnd.n5786 gnd.n5785 19.3944
R8583 gnd.n5785 gnd.n5433 19.3944
R8584 gnd.n5810 gnd.n5433 19.3944
R8585 gnd.n5810 gnd.n5809 19.3944
R8586 gnd.n5809 gnd.n5411 19.3944
R8587 gnd.n5839 gnd.n5411 19.3944
R8588 gnd.n5839 gnd.n5401 19.3944
R8589 gnd.n5857 gnd.n5401 19.3944
R8590 gnd.n5857 gnd.n5856 19.3944
R8591 gnd.n5856 gnd.n5855 19.3944
R8592 gnd.n5855 gnd.n5379 19.3944
R8593 gnd.n5897 gnd.n5379 19.3944
R8594 gnd.n5897 gnd.n5372 19.3944
R8595 gnd.n5908 gnd.n5372 19.3944
R8596 gnd.n5908 gnd.n5368 19.3944
R8597 gnd.n5921 gnd.n5368 19.3944
R8598 gnd.n5921 gnd.n5920 19.3944
R8599 gnd.n5920 gnd.n5347 19.3944
R8600 gnd.n5943 gnd.n5347 19.3944
R8601 gnd.n5943 gnd.n5942 19.3944
R8602 gnd.n5942 gnd.n5276 19.3944
R8603 gnd.n5982 gnd.n5276 19.3944
R8604 gnd.n5982 gnd.n5269 19.3944
R8605 gnd.n5993 gnd.n5269 19.3944
R8606 gnd.n5993 gnd.n5265 19.3944
R8607 gnd.n6005 gnd.n5265 19.3944
R8608 gnd.n6005 gnd.n6004 19.3944
R8609 gnd.n6004 gnd.n5244 19.3944
R8610 gnd.n6029 gnd.n5244 19.3944
R8611 gnd.n6029 gnd.n5232 19.3944
R8612 gnd.n6053 gnd.n5232 19.3944
R8613 gnd.n6053 gnd.n5216 19.3944
R8614 gnd.n6077 gnd.n5216 19.3944
R8615 gnd.n6078 gnd.n6077 19.3944
R8616 gnd.n6078 gnd.n5210 19.3944
R8617 gnd.n5210 gnd.n5208 19.3944
R8618 gnd.n6091 gnd.n5208 19.3944
R8619 gnd.n6091 gnd.n923 19.3944
R8620 gnd.n6514 gnd.n923 19.3944
R8621 gnd.n6514 gnd.n6513 19.3944
R8622 gnd.n6513 gnd.n6512 19.3944
R8623 gnd.n6512 gnd.n927 19.3944
R8624 gnd.n948 gnd.n927 19.3944
R8625 gnd.n6500 gnd.n948 19.3944
R8626 gnd.n6500 gnd.n6499 19.3944
R8627 gnd.n6499 gnd.n6498 19.3944
R8628 gnd.n6498 gnd.n952 19.3944
R8629 gnd.n4477 gnd.n1641 19.3944
R8630 gnd.n4482 gnd.n1641 19.3944
R8631 gnd.n4482 gnd.n1642 19.3944
R8632 gnd.n1642 gnd.n1622 19.3944
R8633 gnd.n4527 gnd.n1622 19.3944
R8634 gnd.n4527 gnd.n1619 19.3944
R8635 gnd.n4532 gnd.n1619 19.3944
R8636 gnd.n4532 gnd.n1620 19.3944
R8637 gnd.n1620 gnd.n1595 19.3944
R8638 gnd.n4559 gnd.n1595 19.3944
R8639 gnd.n4559 gnd.n1592 19.3944
R8640 gnd.n4564 gnd.n1592 19.3944
R8641 gnd.n4564 gnd.n1593 19.3944
R8642 gnd.n1593 gnd.n1566 19.3944
R8643 gnd.n4598 gnd.n1566 19.3944
R8644 gnd.n4598 gnd.n1563 19.3944
R8645 gnd.n4606 gnd.n1563 19.3944
R8646 gnd.n4606 gnd.n1564 19.3944
R8647 gnd.n4602 gnd.n1564 19.3944
R8648 gnd.n4602 gnd.n1555 19.3944
R8649 gnd.n4624 gnd.n1555 19.3944
R8650 gnd.n4624 gnd.n1552 19.3944
R8651 gnd.n4631 gnd.n1552 19.3944
R8652 gnd.n4631 gnd.n1553 19.3944
R8653 gnd.n4627 gnd.n1553 19.3944
R8654 gnd.n4627 gnd.n69 19.3944
R8655 gnd.n7780 gnd.n69 19.3944
R8656 gnd.n7780 gnd.n7779 19.3944
R8657 gnd.n7779 gnd.n7778 19.3944
R8658 gnd.n7778 gnd.n73 19.3944
R8659 gnd.n7774 gnd.n73 19.3944
R8660 gnd.n7774 gnd.n7773 19.3944
R8661 gnd.n7773 gnd.n7772 19.3944
R8662 gnd.n7772 gnd.n78 19.3944
R8663 gnd.n7768 gnd.n78 19.3944
R8664 gnd.n7768 gnd.n7767 19.3944
R8665 gnd.n7767 gnd.n7766 19.3944
R8666 gnd.n7766 gnd.n83 19.3944
R8667 gnd.n7762 gnd.n83 19.3944
R8668 gnd.n7762 gnd.n7761 19.3944
R8669 gnd.n7761 gnd.n7760 19.3944
R8670 gnd.n7760 gnd.n88 19.3944
R8671 gnd.n7756 gnd.n88 19.3944
R8672 gnd.n7756 gnd.n7755 19.3944
R8673 gnd.n7755 gnd.n7754 19.3944
R8674 gnd.n7754 gnd.n93 19.3944
R8675 gnd.n7750 gnd.n93 19.3944
R8676 gnd.n7750 gnd.n7749 19.3944
R8677 gnd.n7749 gnd.n7748 19.3944
R8678 gnd.n7748 gnd.n98 19.3944
R8679 gnd.n7744 gnd.n98 19.3944
R8680 gnd.n7744 gnd.n7743 19.3944
R8681 gnd.n7743 gnd.n7742 19.3944
R8682 gnd.n7641 gnd.n7640 19.3944
R8683 gnd.n7640 gnd.n7639 19.3944
R8684 gnd.n7639 gnd.n7581 19.3944
R8685 gnd.n7635 gnd.n7581 19.3944
R8686 gnd.n7635 gnd.n7634 19.3944
R8687 gnd.n7634 gnd.n7633 19.3944
R8688 gnd.n7633 gnd.n7589 19.3944
R8689 gnd.n7629 gnd.n7589 19.3944
R8690 gnd.n7629 gnd.n7628 19.3944
R8691 gnd.n7628 gnd.n7627 19.3944
R8692 gnd.n7627 gnd.n7597 19.3944
R8693 gnd.n7623 gnd.n7597 19.3944
R8694 gnd.n7623 gnd.n7622 19.3944
R8695 gnd.n7622 gnd.n7621 19.3944
R8696 gnd.n7621 gnd.n7605 19.3944
R8697 gnd.n7617 gnd.n7605 19.3944
R8698 gnd.n1684 gnd.n1683 19.3944
R8699 gnd.n1704 gnd.n1683 19.3944
R8700 gnd.n1704 gnd.n1681 19.3944
R8701 gnd.n1710 gnd.n1681 19.3944
R8702 gnd.n1710 gnd.n1674 19.3944
R8703 gnd.n1723 gnd.n1674 19.3944
R8704 gnd.n1723 gnd.n1672 19.3944
R8705 gnd.n1729 gnd.n1672 19.3944
R8706 gnd.n1729 gnd.n1665 19.3944
R8707 gnd.n1742 gnd.n1665 19.3944
R8708 gnd.n1742 gnd.n1663 19.3944
R8709 gnd.n1748 gnd.n1663 19.3944
R8710 gnd.n1748 gnd.n1656 19.3944
R8711 gnd.n1761 gnd.n1656 19.3944
R8712 gnd.n1761 gnd.n1654 19.3944
R8713 gnd.n1767 gnd.n1654 19.3944
R8714 gnd.n1690 gnd.n1689 19.3944
R8715 gnd.n1689 gnd.n1496 19.3944
R8716 gnd.n4713 gnd.n1496 19.3944
R8717 gnd.n4713 gnd.n1497 19.3944
R8718 gnd.n4709 gnd.n1497 19.3944
R8719 gnd.n4709 gnd.n4708 19.3944
R8720 gnd.n4708 gnd.n4707 19.3944
R8721 gnd.n4707 gnd.n1503 19.3944
R8722 gnd.n4703 gnd.n1503 19.3944
R8723 gnd.n4703 gnd.n4702 19.3944
R8724 gnd.n4702 gnd.n4701 19.3944
R8725 gnd.n4701 gnd.n1508 19.3944
R8726 gnd.n4697 gnd.n1508 19.3944
R8727 gnd.n4697 gnd.n4696 19.3944
R8728 gnd.n4696 gnd.n4695 19.3944
R8729 gnd.n4695 gnd.n1513 19.3944
R8730 gnd.n4691 gnd.n1513 19.3944
R8731 gnd.n4691 gnd.n4690 19.3944
R8732 gnd.n4690 gnd.n4689 19.3944
R8733 gnd.n4689 gnd.n4686 19.3944
R8734 gnd.n4686 gnd.n283 19.3944
R8735 gnd.n7496 gnd.n283 19.3944
R8736 gnd.n7496 gnd.n284 19.3944
R8737 gnd.n7492 gnd.n284 19.3944
R8738 gnd.n7492 gnd.n7491 19.3944
R8739 gnd.n7491 gnd.n7490 19.3944
R8740 gnd.n7490 gnd.n290 19.3944
R8741 gnd.n7485 gnd.n290 19.3944
R8742 gnd.n7485 gnd.n7484 19.3944
R8743 gnd.n7484 gnd.n261 19.3944
R8744 gnd.n7507 gnd.n261 19.3944
R8745 gnd.n7507 gnd.n259 19.3944
R8746 gnd.n7511 gnd.n259 19.3944
R8747 gnd.n7511 gnd.n245 19.3944
R8748 gnd.n7523 gnd.n245 19.3944
R8749 gnd.n7523 gnd.n243 19.3944
R8750 gnd.n7527 gnd.n243 19.3944
R8751 gnd.n7527 gnd.n230 19.3944
R8752 gnd.n7539 gnd.n230 19.3944
R8753 gnd.n7539 gnd.n228 19.3944
R8754 gnd.n7543 gnd.n228 19.3944
R8755 gnd.n7543 gnd.n215 19.3944
R8756 gnd.n7555 gnd.n215 19.3944
R8757 gnd.n7555 gnd.n213 19.3944
R8758 gnd.n7559 gnd.n213 19.3944
R8759 gnd.n7559 gnd.n200 19.3944
R8760 gnd.n7571 gnd.n200 19.3944
R8761 gnd.n7571 gnd.n197 19.3944
R8762 gnd.n7650 gnd.n197 19.3944
R8763 gnd.n7650 gnd.n198 19.3944
R8764 gnd.n7646 gnd.n198 19.3944
R8765 gnd.n7646 gnd.n7645 19.3944
R8766 gnd.n7645 gnd.n7644 19.3944
R8767 gnd.n3287 gnd.n1326 19.3944
R8768 gnd.n3287 gnd.n3286 19.3944
R8769 gnd.n3390 gnd.n3286 19.3944
R8770 gnd.n3390 gnd.n3389 19.3944
R8771 gnd.n3389 gnd.n3294 19.3944
R8772 gnd.n3382 gnd.n3294 19.3944
R8773 gnd.n3382 gnd.n3381 19.3944
R8774 gnd.n3381 gnd.n3305 19.3944
R8775 gnd.n3374 gnd.n3305 19.3944
R8776 gnd.n3374 gnd.n3373 19.3944
R8777 gnd.n3373 gnd.n3316 19.3944
R8778 gnd.n3366 gnd.n3316 19.3944
R8779 gnd.n3366 gnd.n3365 19.3944
R8780 gnd.n3365 gnd.n3328 19.3944
R8781 gnd.n3358 gnd.n3328 19.3944
R8782 gnd.n3358 gnd.n3357 19.3944
R8783 gnd.n7181 gnd.n445 19.3944
R8784 gnd.n7187 gnd.n445 19.3944
R8785 gnd.n7187 gnd.n443 19.3944
R8786 gnd.n7191 gnd.n443 19.3944
R8787 gnd.n7191 gnd.n439 19.3944
R8788 gnd.n7197 gnd.n439 19.3944
R8789 gnd.n7197 gnd.n437 19.3944
R8790 gnd.n7201 gnd.n437 19.3944
R8791 gnd.n7201 gnd.n433 19.3944
R8792 gnd.n7207 gnd.n433 19.3944
R8793 gnd.n7207 gnd.n431 19.3944
R8794 gnd.n7211 gnd.n431 19.3944
R8795 gnd.n7211 gnd.n427 19.3944
R8796 gnd.n7217 gnd.n427 19.3944
R8797 gnd.n7217 gnd.n425 19.3944
R8798 gnd.n7221 gnd.n425 19.3944
R8799 gnd.n7221 gnd.n421 19.3944
R8800 gnd.n7227 gnd.n421 19.3944
R8801 gnd.n7227 gnd.n419 19.3944
R8802 gnd.n7231 gnd.n419 19.3944
R8803 gnd.n7231 gnd.n415 19.3944
R8804 gnd.n7237 gnd.n415 19.3944
R8805 gnd.n7237 gnd.n413 19.3944
R8806 gnd.n7241 gnd.n413 19.3944
R8807 gnd.n7241 gnd.n409 19.3944
R8808 gnd.n7247 gnd.n409 19.3944
R8809 gnd.n7247 gnd.n407 19.3944
R8810 gnd.n7251 gnd.n407 19.3944
R8811 gnd.n7251 gnd.n403 19.3944
R8812 gnd.n7257 gnd.n403 19.3944
R8813 gnd.n7257 gnd.n401 19.3944
R8814 gnd.n7261 gnd.n401 19.3944
R8815 gnd.n7261 gnd.n397 19.3944
R8816 gnd.n7267 gnd.n397 19.3944
R8817 gnd.n7267 gnd.n395 19.3944
R8818 gnd.n7271 gnd.n395 19.3944
R8819 gnd.n7271 gnd.n391 19.3944
R8820 gnd.n7277 gnd.n391 19.3944
R8821 gnd.n7277 gnd.n389 19.3944
R8822 gnd.n7281 gnd.n389 19.3944
R8823 gnd.n7281 gnd.n385 19.3944
R8824 gnd.n7287 gnd.n385 19.3944
R8825 gnd.n7287 gnd.n383 19.3944
R8826 gnd.n7291 gnd.n383 19.3944
R8827 gnd.n7291 gnd.n379 19.3944
R8828 gnd.n7297 gnd.n379 19.3944
R8829 gnd.n7297 gnd.n377 19.3944
R8830 gnd.n7301 gnd.n377 19.3944
R8831 gnd.n7301 gnd.n373 19.3944
R8832 gnd.n7307 gnd.n373 19.3944
R8833 gnd.n7307 gnd.n371 19.3944
R8834 gnd.n7311 gnd.n371 19.3944
R8835 gnd.n7311 gnd.n367 19.3944
R8836 gnd.n7317 gnd.n367 19.3944
R8837 gnd.n7317 gnd.n365 19.3944
R8838 gnd.n7321 gnd.n365 19.3944
R8839 gnd.n7321 gnd.n361 19.3944
R8840 gnd.n7327 gnd.n361 19.3944
R8841 gnd.n7327 gnd.n359 19.3944
R8842 gnd.n7331 gnd.n359 19.3944
R8843 gnd.n7331 gnd.n355 19.3944
R8844 gnd.n7337 gnd.n355 19.3944
R8845 gnd.n7337 gnd.n353 19.3944
R8846 gnd.n7341 gnd.n353 19.3944
R8847 gnd.n7341 gnd.n349 19.3944
R8848 gnd.n7347 gnd.n349 19.3944
R8849 gnd.n7347 gnd.n347 19.3944
R8850 gnd.n7351 gnd.n347 19.3944
R8851 gnd.n7351 gnd.n343 19.3944
R8852 gnd.n7357 gnd.n343 19.3944
R8853 gnd.n7357 gnd.n341 19.3944
R8854 gnd.n7361 gnd.n341 19.3944
R8855 gnd.n7361 gnd.n337 19.3944
R8856 gnd.n7367 gnd.n337 19.3944
R8857 gnd.n7367 gnd.n335 19.3944
R8858 gnd.n7371 gnd.n335 19.3944
R8859 gnd.n7371 gnd.n331 19.3944
R8860 gnd.n7377 gnd.n331 19.3944
R8861 gnd.n7377 gnd.n329 19.3944
R8862 gnd.n7381 gnd.n329 19.3944
R8863 gnd.n7381 gnd.n325 19.3944
R8864 gnd.n7388 gnd.n325 19.3944
R8865 gnd.n7388 gnd.n323 19.3944
R8866 gnd.n7392 gnd.n323 19.3944
R8867 gnd.n6696 gnd.n738 19.3944
R8868 gnd.n6696 gnd.n736 19.3944
R8869 gnd.n6700 gnd.n736 19.3944
R8870 gnd.n6700 gnd.n732 19.3944
R8871 gnd.n6706 gnd.n732 19.3944
R8872 gnd.n6706 gnd.n730 19.3944
R8873 gnd.n6710 gnd.n730 19.3944
R8874 gnd.n6710 gnd.n726 19.3944
R8875 gnd.n6716 gnd.n726 19.3944
R8876 gnd.n6716 gnd.n724 19.3944
R8877 gnd.n6720 gnd.n724 19.3944
R8878 gnd.n6720 gnd.n720 19.3944
R8879 gnd.n6726 gnd.n720 19.3944
R8880 gnd.n6726 gnd.n718 19.3944
R8881 gnd.n6730 gnd.n718 19.3944
R8882 gnd.n6730 gnd.n714 19.3944
R8883 gnd.n6736 gnd.n714 19.3944
R8884 gnd.n6736 gnd.n712 19.3944
R8885 gnd.n6740 gnd.n712 19.3944
R8886 gnd.n6740 gnd.n708 19.3944
R8887 gnd.n6746 gnd.n708 19.3944
R8888 gnd.n6746 gnd.n706 19.3944
R8889 gnd.n6750 gnd.n706 19.3944
R8890 gnd.n6750 gnd.n702 19.3944
R8891 gnd.n6756 gnd.n702 19.3944
R8892 gnd.n6756 gnd.n700 19.3944
R8893 gnd.n6760 gnd.n700 19.3944
R8894 gnd.n6760 gnd.n696 19.3944
R8895 gnd.n6766 gnd.n696 19.3944
R8896 gnd.n6766 gnd.n694 19.3944
R8897 gnd.n6770 gnd.n694 19.3944
R8898 gnd.n6770 gnd.n690 19.3944
R8899 gnd.n6776 gnd.n690 19.3944
R8900 gnd.n6776 gnd.n688 19.3944
R8901 gnd.n6780 gnd.n688 19.3944
R8902 gnd.n6780 gnd.n684 19.3944
R8903 gnd.n6786 gnd.n684 19.3944
R8904 gnd.n6786 gnd.n682 19.3944
R8905 gnd.n6790 gnd.n682 19.3944
R8906 gnd.n6790 gnd.n678 19.3944
R8907 gnd.n6796 gnd.n678 19.3944
R8908 gnd.n6796 gnd.n676 19.3944
R8909 gnd.n6800 gnd.n676 19.3944
R8910 gnd.n6800 gnd.n672 19.3944
R8911 gnd.n6806 gnd.n672 19.3944
R8912 gnd.n6806 gnd.n670 19.3944
R8913 gnd.n6810 gnd.n670 19.3944
R8914 gnd.n6810 gnd.n666 19.3944
R8915 gnd.n6816 gnd.n666 19.3944
R8916 gnd.n6816 gnd.n664 19.3944
R8917 gnd.n6820 gnd.n664 19.3944
R8918 gnd.n6820 gnd.n660 19.3944
R8919 gnd.n6826 gnd.n660 19.3944
R8920 gnd.n6826 gnd.n658 19.3944
R8921 gnd.n6830 gnd.n658 19.3944
R8922 gnd.n6830 gnd.n654 19.3944
R8923 gnd.n6836 gnd.n654 19.3944
R8924 gnd.n6836 gnd.n652 19.3944
R8925 gnd.n6840 gnd.n652 19.3944
R8926 gnd.n6840 gnd.n648 19.3944
R8927 gnd.n6846 gnd.n648 19.3944
R8928 gnd.n6846 gnd.n646 19.3944
R8929 gnd.n6850 gnd.n646 19.3944
R8930 gnd.n6850 gnd.n642 19.3944
R8931 gnd.n6856 gnd.n642 19.3944
R8932 gnd.n6856 gnd.n640 19.3944
R8933 gnd.n6860 gnd.n640 19.3944
R8934 gnd.n6860 gnd.n636 19.3944
R8935 gnd.n6866 gnd.n636 19.3944
R8936 gnd.n6866 gnd.n634 19.3944
R8937 gnd.n6870 gnd.n634 19.3944
R8938 gnd.n6870 gnd.n630 19.3944
R8939 gnd.n6876 gnd.n630 19.3944
R8940 gnd.n6876 gnd.n628 19.3944
R8941 gnd.n6880 gnd.n628 19.3944
R8942 gnd.n6880 gnd.n624 19.3944
R8943 gnd.n6886 gnd.n624 19.3944
R8944 gnd.n6886 gnd.n622 19.3944
R8945 gnd.n6890 gnd.n622 19.3944
R8946 gnd.n6890 gnd.n618 19.3944
R8947 gnd.n6896 gnd.n618 19.3944
R8948 gnd.n6896 gnd.n616 19.3944
R8949 gnd.n6900 gnd.n616 19.3944
R8950 gnd.n6900 gnd.n612 19.3944
R8951 gnd.n6906 gnd.n612 19.3944
R8952 gnd.n6906 gnd.n610 19.3944
R8953 gnd.n6910 gnd.n610 19.3944
R8954 gnd.n6910 gnd.n606 19.3944
R8955 gnd.n6916 gnd.n606 19.3944
R8956 gnd.n6916 gnd.n604 19.3944
R8957 gnd.n6920 gnd.n604 19.3944
R8958 gnd.n6920 gnd.n600 19.3944
R8959 gnd.n6926 gnd.n600 19.3944
R8960 gnd.n6926 gnd.n598 19.3944
R8961 gnd.n6930 gnd.n598 19.3944
R8962 gnd.n6930 gnd.n594 19.3944
R8963 gnd.n6936 gnd.n594 19.3944
R8964 gnd.n6936 gnd.n592 19.3944
R8965 gnd.n6940 gnd.n592 19.3944
R8966 gnd.n6940 gnd.n588 19.3944
R8967 gnd.n6946 gnd.n588 19.3944
R8968 gnd.n6946 gnd.n586 19.3944
R8969 gnd.n6950 gnd.n586 19.3944
R8970 gnd.n6950 gnd.n582 19.3944
R8971 gnd.n6956 gnd.n582 19.3944
R8972 gnd.n6956 gnd.n580 19.3944
R8973 gnd.n6960 gnd.n580 19.3944
R8974 gnd.n6960 gnd.n576 19.3944
R8975 gnd.n6966 gnd.n576 19.3944
R8976 gnd.n6966 gnd.n574 19.3944
R8977 gnd.n6970 gnd.n574 19.3944
R8978 gnd.n6970 gnd.n570 19.3944
R8979 gnd.n6976 gnd.n570 19.3944
R8980 gnd.n6976 gnd.n568 19.3944
R8981 gnd.n6980 gnd.n568 19.3944
R8982 gnd.n6980 gnd.n564 19.3944
R8983 gnd.n6986 gnd.n564 19.3944
R8984 gnd.n6986 gnd.n562 19.3944
R8985 gnd.n6990 gnd.n562 19.3944
R8986 gnd.n6990 gnd.n558 19.3944
R8987 gnd.n6996 gnd.n558 19.3944
R8988 gnd.n6996 gnd.n556 19.3944
R8989 gnd.n7000 gnd.n556 19.3944
R8990 gnd.n7000 gnd.n552 19.3944
R8991 gnd.n7006 gnd.n552 19.3944
R8992 gnd.n7006 gnd.n550 19.3944
R8993 gnd.n7010 gnd.n550 19.3944
R8994 gnd.n7010 gnd.n546 19.3944
R8995 gnd.n7016 gnd.n546 19.3944
R8996 gnd.n7016 gnd.n544 19.3944
R8997 gnd.n7020 gnd.n544 19.3944
R8998 gnd.n7020 gnd.n540 19.3944
R8999 gnd.n7026 gnd.n540 19.3944
R9000 gnd.n7026 gnd.n538 19.3944
R9001 gnd.n7030 gnd.n538 19.3944
R9002 gnd.n7030 gnd.n534 19.3944
R9003 gnd.n7036 gnd.n534 19.3944
R9004 gnd.n7036 gnd.n532 19.3944
R9005 gnd.n7040 gnd.n532 19.3944
R9006 gnd.n7040 gnd.n528 19.3944
R9007 gnd.n7046 gnd.n528 19.3944
R9008 gnd.n7046 gnd.n526 19.3944
R9009 gnd.n7050 gnd.n526 19.3944
R9010 gnd.n7050 gnd.n522 19.3944
R9011 gnd.n7056 gnd.n522 19.3944
R9012 gnd.n7056 gnd.n520 19.3944
R9013 gnd.n7060 gnd.n520 19.3944
R9014 gnd.n7060 gnd.n516 19.3944
R9015 gnd.n7066 gnd.n516 19.3944
R9016 gnd.n7066 gnd.n514 19.3944
R9017 gnd.n7070 gnd.n514 19.3944
R9018 gnd.n7070 gnd.n510 19.3944
R9019 gnd.n7076 gnd.n510 19.3944
R9020 gnd.n7076 gnd.n508 19.3944
R9021 gnd.n7080 gnd.n508 19.3944
R9022 gnd.n7080 gnd.n504 19.3944
R9023 gnd.n7086 gnd.n504 19.3944
R9024 gnd.n7086 gnd.n502 19.3944
R9025 gnd.n7090 gnd.n502 19.3944
R9026 gnd.n7090 gnd.n498 19.3944
R9027 gnd.n7096 gnd.n498 19.3944
R9028 gnd.n7096 gnd.n496 19.3944
R9029 gnd.n7100 gnd.n496 19.3944
R9030 gnd.n7100 gnd.n492 19.3944
R9031 gnd.n7106 gnd.n492 19.3944
R9032 gnd.n7106 gnd.n490 19.3944
R9033 gnd.n7110 gnd.n490 19.3944
R9034 gnd.n7110 gnd.n486 19.3944
R9035 gnd.n7116 gnd.n486 19.3944
R9036 gnd.n7116 gnd.n484 19.3944
R9037 gnd.n7120 gnd.n484 19.3944
R9038 gnd.n7120 gnd.n480 19.3944
R9039 gnd.n7126 gnd.n480 19.3944
R9040 gnd.n7126 gnd.n478 19.3944
R9041 gnd.n7130 gnd.n478 19.3944
R9042 gnd.n7130 gnd.n474 19.3944
R9043 gnd.n7136 gnd.n474 19.3944
R9044 gnd.n7136 gnd.n472 19.3944
R9045 gnd.n7140 gnd.n472 19.3944
R9046 gnd.n7140 gnd.n468 19.3944
R9047 gnd.n7146 gnd.n468 19.3944
R9048 gnd.n7146 gnd.n466 19.3944
R9049 gnd.n7150 gnd.n466 19.3944
R9050 gnd.n7150 gnd.n462 19.3944
R9051 gnd.n7156 gnd.n462 19.3944
R9052 gnd.n7156 gnd.n460 19.3944
R9053 gnd.n7160 gnd.n460 19.3944
R9054 gnd.n7160 gnd.n456 19.3944
R9055 gnd.n7166 gnd.n456 19.3944
R9056 gnd.n7166 gnd.n454 19.3944
R9057 gnd.n7171 gnd.n454 19.3944
R9058 gnd.n7171 gnd.n450 19.3944
R9059 gnd.n7177 gnd.n450 19.3944
R9060 gnd.n7178 gnd.n7177 19.3944
R9061 gnd.n1912 gnd.n1908 19.3944
R9062 gnd.n1912 gnd.n1905 19.3944
R9063 gnd.n1916 gnd.n1905 19.3944
R9064 gnd.n1916 gnd.n1903 19.3944
R9065 gnd.n1922 gnd.n1903 19.3944
R9066 gnd.n1922 gnd.n1901 19.3944
R9067 gnd.n1926 gnd.n1901 19.3944
R9068 gnd.n1926 gnd.n1899 19.3944
R9069 gnd.n1932 gnd.n1899 19.3944
R9070 gnd.n1932 gnd.n1897 19.3944
R9071 gnd.n1937 gnd.n1897 19.3944
R9072 gnd.n1937 gnd.n1895 19.3944
R9073 gnd.n1895 gnd.n1892 19.3944
R9074 gnd.n1944 gnd.n1892 19.3944
R9075 gnd.n1944 gnd.n1889 19.3944
R9076 gnd.n2029 gnd.n1951 19.3944
R9077 gnd.n2023 gnd.n1951 19.3944
R9078 gnd.n2023 gnd.n2022 19.3944
R9079 gnd.n2022 gnd.n2021 19.3944
R9080 gnd.n2021 gnd.n1957 19.3944
R9081 gnd.n2015 gnd.n1957 19.3944
R9082 gnd.n2015 gnd.n2014 19.3944
R9083 gnd.n2014 gnd.n2013 19.3944
R9084 gnd.n2013 gnd.n1963 19.3944
R9085 gnd.n2007 gnd.n1963 19.3944
R9086 gnd.n2007 gnd.n2006 19.3944
R9087 gnd.n2006 gnd.n2005 19.3944
R9088 gnd.n2005 gnd.n1969 19.3944
R9089 gnd.n1999 gnd.n1969 19.3944
R9090 gnd.n1999 gnd.n1998 19.3944
R9091 gnd.n1998 gnd.n1997 19.3944
R9092 gnd.n1997 gnd.n1975 19.3944
R9093 gnd.n1991 gnd.n1975 19.3944
R9094 gnd.n1983 gnd.n1640 19.3944
R9095 gnd.n4486 gnd.n1640 19.3944
R9096 gnd.n4487 gnd.n4486 19.3944
R9097 gnd.n4487 gnd.n1638 19.3944
R9098 gnd.n4515 gnd.n1638 19.3944
R9099 gnd.n4515 gnd.n4514 19.3944
R9100 gnd.n4514 gnd.n4513 19.3944
R9101 gnd.n4513 gnd.n4512 19.3944
R9102 gnd.n4512 gnd.n4511 19.3944
R9103 gnd.n4511 gnd.n4509 19.3944
R9104 gnd.n4509 gnd.n4508 19.3944
R9105 gnd.n4508 gnd.n4506 19.3944
R9106 gnd.n4506 gnd.n4505 19.3944
R9107 gnd.n4505 gnd.n4504 19.3944
R9108 gnd.n4504 gnd.n4502 19.3944
R9109 gnd.n4502 gnd.n1558 19.3944
R9110 gnd.n4611 gnd.n1558 19.3944
R9111 gnd.n4612 gnd.n4611 19.3944
R9112 gnd.n4614 gnd.n4612 19.3944
R9113 gnd.n4614 gnd.n1556 19.3944
R9114 gnd.n4620 gnd.n1556 19.3944
R9115 gnd.n4620 gnd.n4619 19.3944
R9116 gnd.n4619 gnd.n1550 19.3944
R9117 gnd.n4637 gnd.n1550 19.3944
R9118 gnd.n4637 gnd.n1548 19.3944
R9119 gnd.n4641 gnd.n1548 19.3944
R9120 gnd.n4641 gnd.n299 19.3944
R9121 gnd.n7475 gnd.n299 19.3944
R9122 gnd.n7475 gnd.n7474 19.3944
R9123 gnd.n7474 gnd.n7473 19.3944
R9124 gnd.n7473 gnd.n304 19.3944
R9125 gnd.n7405 gnd.n304 19.3944
R9126 gnd.n7405 gnd.n7401 19.3944
R9127 gnd.n7412 gnd.n7401 19.3944
R9128 gnd.n7413 gnd.n7412 19.3944
R9129 gnd.n7416 gnd.n7413 19.3944
R9130 gnd.n7416 gnd.n7399 19.3944
R9131 gnd.n7451 gnd.n7399 19.3944
R9132 gnd.n7451 gnd.n7450 19.3944
R9133 gnd.n7450 gnd.n7449 19.3944
R9134 gnd.n7449 gnd.n7446 19.3944
R9135 gnd.n7446 gnd.n7445 19.3944
R9136 gnd.n7445 gnd.n7443 19.3944
R9137 gnd.n7443 gnd.n7442 19.3944
R9138 gnd.n7442 gnd.n7440 19.3944
R9139 gnd.n7440 gnd.n7439 19.3944
R9140 gnd.n7439 gnd.n7437 19.3944
R9141 gnd.n7437 gnd.n7436 19.3944
R9142 gnd.n7436 gnd.n7434 19.3944
R9143 gnd.n7434 gnd.n7433 19.3944
R9144 gnd.n7433 gnd.n183 19.3944
R9145 gnd.n7663 gnd.n183 19.3944
R9146 gnd.n7664 gnd.n7663 19.3944
R9147 gnd.n7702 gnd.n144 19.3944
R9148 gnd.n7697 gnd.n144 19.3944
R9149 gnd.n7697 gnd.n7696 19.3944
R9150 gnd.n7696 gnd.n7695 19.3944
R9151 gnd.n7695 gnd.n151 19.3944
R9152 gnd.n7690 gnd.n151 19.3944
R9153 gnd.n7690 gnd.n7689 19.3944
R9154 gnd.n7689 gnd.n7688 19.3944
R9155 gnd.n7688 gnd.n158 19.3944
R9156 gnd.n7683 gnd.n158 19.3944
R9157 gnd.n7683 gnd.n7682 19.3944
R9158 gnd.n7682 gnd.n7681 19.3944
R9159 gnd.n7681 gnd.n165 19.3944
R9160 gnd.n7676 gnd.n165 19.3944
R9161 gnd.n7676 gnd.n7675 19.3944
R9162 gnd.n7675 gnd.n7674 19.3944
R9163 gnd.n7674 gnd.n172 19.3944
R9164 gnd.n7669 gnd.n172 19.3944
R9165 gnd.n7735 gnd.n7734 19.3944
R9166 gnd.n7734 gnd.n7733 19.3944
R9167 gnd.n7733 gnd.n115 19.3944
R9168 gnd.n7728 gnd.n115 19.3944
R9169 gnd.n7728 gnd.n7727 19.3944
R9170 gnd.n7727 gnd.n7726 19.3944
R9171 gnd.n7726 gnd.n123 19.3944
R9172 gnd.n7721 gnd.n123 19.3944
R9173 gnd.n7721 gnd.n7720 19.3944
R9174 gnd.n7720 gnd.n7719 19.3944
R9175 gnd.n7719 gnd.n130 19.3944
R9176 gnd.n7714 gnd.n130 19.3944
R9177 gnd.n7714 gnd.n7713 19.3944
R9178 gnd.n7713 gnd.n7712 19.3944
R9179 gnd.n7712 gnd.n137 19.3944
R9180 gnd.n7707 gnd.n137 19.3944
R9181 gnd.n7707 gnd.n7706 19.3944
R9182 gnd.n4719 gnd.n1484 19.3944
R9183 gnd.n4719 gnd.n4718 19.3944
R9184 gnd.n4718 gnd.n4717 19.3944
R9185 gnd.n4717 gnd.n1488 19.3944
R9186 gnd.n4523 gnd.n1488 19.3944
R9187 gnd.n4523 gnd.n4522 19.3944
R9188 gnd.n4522 gnd.n1603 19.3944
R9189 gnd.n4549 gnd.n1603 19.3944
R9190 gnd.n4549 gnd.n1601 19.3944
R9191 gnd.n4555 gnd.n1601 19.3944
R9192 gnd.n4555 gnd.n4554 19.3944
R9193 gnd.n4554 gnd.n1576 19.3944
R9194 gnd.n4588 gnd.n1576 19.3944
R9195 gnd.n4588 gnd.n1574 19.3944
R9196 gnd.n4594 gnd.n1574 19.3944
R9197 gnd.n4594 gnd.n4593 19.3944
R9198 gnd.n4593 gnd.n1524 19.3944
R9199 gnd.n4678 gnd.n1524 19.3944
R9200 gnd.n4678 gnd.n1522 19.3944
R9201 gnd.n4682 gnd.n1522 19.3944
R9202 gnd.n4682 gnd.n274 19.3944
R9203 gnd.n7500 gnd.n274 19.3944
R9204 gnd.n273 gnd.n272 19.3944
R9205 gnd.n4659 gnd.n272 19.3944
R9206 gnd.n1547 gnd.n1546 19.3944
R9207 gnd.n7480 gnd.n7479 19.3944
R9208 gnd.n7503 gnd.n266 19.3944
R9209 gnd.n7503 gnd.n253 19.3944
R9210 gnd.n7515 gnd.n253 19.3944
R9211 gnd.n7515 gnd.n251 19.3944
R9212 gnd.n7519 gnd.n251 19.3944
R9213 gnd.n7519 gnd.n237 19.3944
R9214 gnd.n7531 gnd.n237 19.3944
R9215 gnd.n7531 gnd.n235 19.3944
R9216 gnd.n7535 gnd.n235 19.3944
R9217 gnd.n7535 gnd.n223 19.3944
R9218 gnd.n7547 gnd.n223 19.3944
R9219 gnd.n7547 gnd.n221 19.3944
R9220 gnd.n7551 gnd.n221 19.3944
R9221 gnd.n7551 gnd.n206 19.3944
R9222 gnd.n7563 gnd.n206 19.3944
R9223 gnd.n7563 gnd.n204 19.3944
R9224 gnd.n7567 gnd.n204 19.3944
R9225 gnd.n7567 gnd.n191 19.3944
R9226 gnd.n7654 gnd.n191 19.3944
R9227 gnd.n7654 gnd.n189 19.3944
R9228 gnd.n7658 gnd.n189 19.3944
R9229 gnd.n7658 gnd.n110 19.3944
R9230 gnd.n7738 gnd.n110 19.3944
R9231 gnd.n2864 gnd.n2857 19.3944
R9232 gnd.n2864 gnd.n2855 19.3944
R9233 gnd.n2868 gnd.n2855 19.3944
R9234 gnd.n2868 gnd.n2853 19.3944
R9235 gnd.n2941 gnd.n2853 19.3944
R9236 gnd.n2941 gnd.n2940 19.3944
R9237 gnd.n2940 gnd.n2939 19.3944
R9238 gnd.n2939 gnd.n2874 19.3944
R9239 gnd.n2935 gnd.n2874 19.3944
R9240 gnd.n2930 gnd.n2876 19.3944
R9241 gnd.n2926 gnd.n2881 19.3944
R9242 gnd.n2924 gnd.n2923 19.3944
R9243 gnd.n2920 gnd.n2919 19.3944
R9244 gnd.n2916 gnd.n2915 19.3944
R9245 gnd.n2915 gnd.n2914 19.3944
R9246 gnd.n2914 gnd.n2884 19.3944
R9247 gnd.n2910 gnd.n2884 19.3944
R9248 gnd.n2910 gnd.n2909 19.3944
R9249 gnd.n2909 gnd.n2908 19.3944
R9250 gnd.n2908 gnd.n2890 19.3944
R9251 gnd.n2904 gnd.n2890 19.3944
R9252 gnd.n2904 gnd.n2903 19.3944
R9253 gnd.n2903 gnd.n2902 19.3944
R9254 gnd.n2902 gnd.n2899 19.3944
R9255 gnd.n2899 gnd.n2898 19.3944
R9256 gnd.n2898 gnd.n2792 19.3944
R9257 gnd.n3241 gnd.n2792 19.3944
R9258 gnd.n3241 gnd.n2790 19.3944
R9259 gnd.n3245 gnd.n2790 19.3944
R9260 gnd.n3245 gnd.n2788 19.3944
R9261 gnd.n3249 gnd.n2788 19.3944
R9262 gnd.n3249 gnd.n2786 19.3944
R9263 gnd.n3253 gnd.n2786 19.3944
R9264 gnd.n3253 gnd.n2784 19.3944
R9265 gnd.n3257 gnd.n2784 19.3944
R9266 gnd.n3257 gnd.n2782 19.3944
R9267 gnd.n3261 gnd.n2782 19.3944
R9268 gnd.n3261 gnd.n2779 19.3944
R9269 gnd.n3400 gnd.n2779 19.3944
R9270 gnd.n3400 gnd.n2777 19.3944
R9271 gnd.n3404 gnd.n2777 19.3944
R9272 gnd.n3404 gnd.n2773 19.3944
R9273 gnd.n3414 gnd.n2773 19.3944
R9274 gnd.n3414 gnd.n2771 19.3944
R9275 gnd.n3418 gnd.n2771 19.3944
R9276 gnd.n3418 gnd.n2765 19.3944
R9277 gnd.n3428 gnd.n2765 19.3944
R9278 gnd.n3428 gnd.n2763 19.3944
R9279 gnd.n3432 gnd.n2763 19.3944
R9280 gnd.n3432 gnd.n2757 19.3944
R9281 gnd.n3445 gnd.n2757 19.3944
R9282 gnd.n3445 gnd.n2755 19.3944
R9283 gnd.n3449 gnd.n2755 19.3944
R9284 gnd.n3449 gnd.n2752 19.3944
R9285 gnd.n3459 gnd.n2752 19.3944
R9286 gnd.n3459 gnd.n2750 19.3944
R9287 gnd.n3465 gnd.n2750 19.3944
R9288 gnd.n3465 gnd.n3464 19.3944
R9289 gnd.n3464 gnd.n2398 19.3944
R9290 gnd.n3648 gnd.n2398 19.3944
R9291 gnd.n3648 gnd.n2396 19.3944
R9292 gnd.n3652 gnd.n2396 19.3944
R9293 gnd.n3652 gnd.n2377 19.3944
R9294 gnd.n3677 gnd.n2377 19.3944
R9295 gnd.n3677 gnd.n2375 19.3944
R9296 gnd.n3683 gnd.n2375 19.3944
R9297 gnd.n3683 gnd.n3682 19.3944
R9298 gnd.n3682 gnd.n2350 19.3944
R9299 gnd.n3715 gnd.n2350 19.3944
R9300 gnd.n3715 gnd.n2348 19.3944
R9301 gnd.n3721 gnd.n2348 19.3944
R9302 gnd.n3721 gnd.n3720 19.3944
R9303 gnd.n3720 gnd.n2323 19.3944
R9304 gnd.n3751 gnd.n2323 19.3944
R9305 gnd.n3751 gnd.n2321 19.3944
R9306 gnd.n3755 gnd.n2321 19.3944
R9307 gnd.n3755 gnd.n2301 19.3944
R9308 gnd.n3779 gnd.n2301 19.3944
R9309 gnd.n3779 gnd.n2299 19.3944
R9310 gnd.n3785 gnd.n2299 19.3944
R9311 gnd.n3785 gnd.n3784 19.3944
R9312 gnd.n3784 gnd.n2273 19.3944
R9313 gnd.n3829 gnd.n2273 19.3944
R9314 gnd.n3829 gnd.n2271 19.3944
R9315 gnd.n3835 gnd.n2271 19.3944
R9316 gnd.n3835 gnd.n3834 19.3944
R9317 gnd.n3834 gnd.n2254 19.3944
R9318 gnd.n3856 gnd.n2254 19.3944
R9319 gnd.n3856 gnd.n2252 19.3944
R9320 gnd.n3860 gnd.n2252 19.3944
R9321 gnd.n3860 gnd.n2209 19.3944
R9322 gnd.n3899 gnd.n2209 19.3944
R9323 gnd.n3899 gnd.n2207 19.3944
R9324 gnd.n3903 gnd.n2207 19.3944
R9325 gnd.n3903 gnd.n2187 19.3944
R9326 gnd.n3941 gnd.n2187 19.3944
R9327 gnd.n3941 gnd.n2185 19.3944
R9328 gnd.n3947 gnd.n2185 19.3944
R9329 gnd.n3947 gnd.n3946 19.3944
R9330 gnd.n3946 gnd.n2160 19.3944
R9331 gnd.n3993 gnd.n2160 19.3944
R9332 gnd.n3993 gnd.n2158 19.3944
R9333 gnd.n3999 gnd.n2158 19.3944
R9334 gnd.n3999 gnd.n3998 19.3944
R9335 gnd.n3998 gnd.n2129 19.3944
R9336 gnd.n4044 gnd.n2129 19.3944
R9337 gnd.n4044 gnd.n2127 19.3944
R9338 gnd.n4048 gnd.n2127 19.3944
R9339 gnd.n4048 gnd.n2114 19.3944
R9340 gnd.n4076 gnd.n2114 19.3944
R9341 gnd.n4076 gnd.n2112 19.3944
R9342 gnd.n4085 gnd.n2112 19.3944
R9343 gnd.n4085 gnd.n4084 19.3944
R9344 gnd.n4084 gnd.n4083 19.3944
R9345 gnd.n4083 gnd.n2079 19.3944
R9346 gnd.n4150 gnd.n2079 19.3944
R9347 gnd.n4150 gnd.n2077 19.3944
R9348 gnd.n4156 gnd.n2077 19.3944
R9349 gnd.n4156 gnd.n4155 19.3944
R9350 gnd.n4155 gnd.n2051 19.3944
R9351 gnd.n4193 gnd.n2051 19.3944
R9352 gnd.n4193 gnd.n2049 19.3944
R9353 gnd.n4202 gnd.n2049 19.3944
R9354 gnd.n4202 gnd.n4201 19.3944
R9355 gnd.n4201 gnd.n4200 19.3944
R9356 gnd.n4200 gnd.n1845 19.3944
R9357 gnd.n4379 gnd.n1845 19.3944
R9358 gnd.n4379 gnd.n1843 19.3944
R9359 gnd.n4383 gnd.n1843 19.3944
R9360 gnd.n4383 gnd.n1832 19.3944
R9361 gnd.n4399 gnd.n1832 19.3944
R9362 gnd.n4399 gnd.n1830 19.3944
R9363 gnd.n4403 gnd.n1830 19.3944
R9364 gnd.n4403 gnd.n1819 19.3944
R9365 gnd.n4419 gnd.n1819 19.3944
R9366 gnd.n4419 gnd.n1817 19.3944
R9367 gnd.n4423 gnd.n1817 19.3944
R9368 gnd.n4423 gnd.n1806 19.3944
R9369 gnd.n4442 gnd.n1806 19.3944
R9370 gnd.n4442 gnd.n1804 19.3944
R9371 gnd.n4447 gnd.n1804 19.3944
R9372 gnd.n4447 gnd.n1461 19.3944
R9373 gnd.n4734 gnd.n1461 19.3944
R9374 gnd.n4734 gnd.n4733 19.3944
R9375 gnd.n4733 gnd.n4732 19.3944
R9376 gnd.n4732 gnd.n1465 19.3944
R9377 gnd.n4726 gnd.n1465 19.3944
R9378 gnd.n4726 gnd.n4725 19.3944
R9379 gnd.n4725 gnd.n4724 19.3944
R9380 gnd.n4724 gnd.n1474 19.3944
R9381 gnd.n1628 gnd.n1474 19.3944
R9382 gnd.n1628 gnd.n1625 19.3944
R9383 gnd.n1632 gnd.n1625 19.3944
R9384 gnd.n1632 gnd.n1614 19.3944
R9385 gnd.n4537 gnd.n1614 19.3944
R9386 gnd.n4537 gnd.n1612 19.3944
R9387 gnd.n4543 gnd.n1612 19.3944
R9388 gnd.n4543 gnd.n4542 19.3944
R9389 gnd.n4542 gnd.n1587 19.3944
R9390 gnd.n4570 gnd.n1587 19.3944
R9391 gnd.n4570 gnd.n1585 19.3944
R9392 gnd.n4583 gnd.n1585 19.3944
R9393 gnd.n4583 gnd.n4582 19.3944
R9394 gnd.n4582 gnd.n4581 19.3944
R9395 gnd.n4581 gnd.n4578 19.3944
R9396 gnd.n4578 gnd.n1532 19.3944
R9397 gnd.n4673 gnd.n1532 19.3944
R9398 gnd.n4673 gnd.n4672 19.3944
R9399 gnd.n4672 gnd.n4671 19.3944
R9400 gnd.n4671 gnd.n1537 19.3944
R9401 gnd.n4667 gnd.n1537 19.3944
R9402 gnd.n4665 gnd.n4664 19.3944
R9403 gnd.n4654 gnd.n4648 19.3944
R9404 gnd.n4652 gnd.n4651 19.3944
R9405 gnd.n7468 gnd.n308 19.3944
R9406 gnd.n7466 gnd.n7465 19.3944
R9407 gnd.n7465 gnd.n310 19.3944
R9408 gnd.n7461 gnd.n310 19.3944
R9409 gnd.n7461 gnd.n7460 19.3944
R9410 gnd.n7460 gnd.n7459 19.3944
R9411 gnd.n7459 gnd.n316 19.3944
R9412 gnd.n7398 gnd.n316 19.3944
R9413 gnd.n7398 gnd.n7397 19.3944
R9414 gnd.n7397 gnd.n7396 19.3944
R9415 gnd.n5132 gnd.n5131 19.3944
R9416 gnd.n5131 gnd.n5130 19.3944
R9417 gnd.n5130 gnd.n5129 19.3944
R9418 gnd.n5129 gnd.n5127 19.3944
R9419 gnd.n5127 gnd.n5124 19.3944
R9420 gnd.n5124 gnd.n5123 19.3944
R9421 gnd.n5123 gnd.n5120 19.3944
R9422 gnd.n5120 gnd.n5119 19.3944
R9423 gnd.n5119 gnd.n5116 19.3944
R9424 gnd.n5116 gnd.n5115 19.3944
R9425 gnd.n5115 gnd.n5112 19.3944
R9426 gnd.n5112 gnd.n5111 19.3944
R9427 gnd.n5111 gnd.n5108 19.3944
R9428 gnd.n5108 gnd.n5107 19.3944
R9429 gnd.n5107 gnd.n5104 19.3944
R9430 gnd.n5104 gnd.n5103 19.3944
R9431 gnd.n5103 gnd.n5100 19.3944
R9432 gnd.n5098 gnd.n5095 19.3944
R9433 gnd.n5095 gnd.n5094 19.3944
R9434 gnd.n5094 gnd.n5091 19.3944
R9435 gnd.n5091 gnd.n5090 19.3944
R9436 gnd.n5090 gnd.n5087 19.3944
R9437 gnd.n5087 gnd.n5086 19.3944
R9438 gnd.n5086 gnd.n5083 19.3944
R9439 gnd.n5083 gnd.n5082 19.3944
R9440 gnd.n5082 gnd.n5079 19.3944
R9441 gnd.n5079 gnd.n5078 19.3944
R9442 gnd.n5078 gnd.n5075 19.3944
R9443 gnd.n5075 gnd.n5074 19.3944
R9444 gnd.n5074 gnd.n5071 19.3944
R9445 gnd.n5071 gnd.n5070 19.3944
R9446 gnd.n5070 gnd.n5067 19.3944
R9447 gnd.n5067 gnd.n5066 19.3944
R9448 gnd.n5066 gnd.n5063 19.3944
R9449 gnd.n5063 gnd.n5062 19.3944
R9450 gnd.n5055 gnd.n5054 19.3944
R9451 gnd.n5054 gnd.n1058 19.3944
R9452 gnd.n5050 gnd.n1058 19.3944
R9453 gnd.n5050 gnd.n1060 19.3944
R9454 gnd.n3063 gnd.n1060 19.3944
R9455 gnd.n3065 gnd.n3063 19.3944
R9456 gnd.n3065 gnd.n3061 19.3944
R9457 gnd.n3070 gnd.n3061 19.3944
R9458 gnd.n3071 gnd.n3070 19.3944
R9459 gnd.n3073 gnd.n3071 19.3944
R9460 gnd.n3073 gnd.n3059 19.3944
R9461 gnd.n3077 gnd.n3059 19.3944
R9462 gnd.n3077 gnd.n2949 19.3944
R9463 gnd.n3089 gnd.n2949 19.3944
R9464 gnd.n3089 gnd.n2947 19.3944
R9465 gnd.n3093 gnd.n2947 19.3944
R9466 gnd.n3093 gnd.n2850 19.3944
R9467 gnd.n3105 gnd.n2850 19.3944
R9468 gnd.n3105 gnd.n2848 19.3944
R9469 gnd.n3109 gnd.n2848 19.3944
R9470 gnd.n3109 gnd.n2843 19.3944
R9471 gnd.n3121 gnd.n2843 19.3944
R9472 gnd.n3121 gnd.n2841 19.3944
R9473 gnd.n3125 gnd.n2841 19.3944
R9474 gnd.n3125 gnd.n2836 19.3944
R9475 gnd.n3138 gnd.n2836 19.3944
R9476 gnd.n3138 gnd.n2833 19.3944
R9477 gnd.n3143 gnd.n2833 19.3944
R9478 gnd.n3143 gnd.n2828 19.3944
R9479 gnd.n3155 gnd.n2828 19.3944
R9480 gnd.n3155 gnd.n2826 19.3944
R9481 gnd.n3159 gnd.n2826 19.3944
R9482 gnd.n3159 gnd.n2821 19.3944
R9483 gnd.n3171 gnd.n2821 19.3944
R9484 gnd.n3171 gnd.n2819 19.3944
R9485 gnd.n3175 gnd.n2819 19.3944
R9486 gnd.n3175 gnd.n2814 19.3944
R9487 gnd.n3187 gnd.n2814 19.3944
R9488 gnd.n3187 gnd.n2812 19.3944
R9489 gnd.n3192 gnd.n2812 19.3944
R9490 gnd.n3192 gnd.n2806 19.3944
R9491 gnd.n3204 gnd.n2806 19.3944
R9492 gnd.n3205 gnd.n3204 19.3944
R9493 gnd.n3206 gnd.n3205 19.3944
R9494 gnd.n3206 gnd.n2804 19.3944
R9495 gnd.n3212 gnd.n2804 19.3944
R9496 gnd.n3213 gnd.n3212 19.3944
R9497 gnd.n3216 gnd.n3213 19.3944
R9498 gnd.n3216 gnd.n2802 19.3944
R9499 gnd.n3221 gnd.n2802 19.3944
R9500 gnd.n3221 gnd.n2700 19.3944
R9501 gnd.n3530 gnd.n2700 19.3944
R9502 gnd.n3531 gnd.n3530 19.3944
R9503 gnd.n3569 gnd.n2603 19.3944
R9504 gnd.n3569 gnd.n2610 19.3944
R9505 gnd.n2667 gnd.n2610 19.3944
R9506 gnd.n3562 gnd.n2667 19.3944
R9507 gnd.n3562 gnd.n3561 19.3944
R9508 gnd.n3561 gnd.n3560 19.3944
R9509 gnd.n3560 gnd.n2673 19.3944
R9510 gnd.n3555 gnd.n2673 19.3944
R9511 gnd.n3555 gnd.n3554 19.3944
R9512 gnd.n3554 gnd.n3553 19.3944
R9513 gnd.n3553 gnd.n2680 19.3944
R9514 gnd.n3548 gnd.n2680 19.3944
R9515 gnd.n3548 gnd.n3547 19.3944
R9516 gnd.n3547 gnd.n3546 19.3944
R9517 gnd.n3546 gnd.n2687 19.3944
R9518 gnd.n3541 gnd.n2687 19.3944
R9519 gnd.n3541 gnd.n3540 19.3944
R9520 gnd.n3540 gnd.n3539 19.3944
R9521 gnd.n2623 gnd.n2622 19.3944
R9522 gnd.n2663 gnd.n2622 19.3944
R9523 gnd.n2663 gnd.n2662 19.3944
R9524 gnd.n2662 gnd.n2661 19.3944
R9525 gnd.n2661 gnd.n2658 19.3944
R9526 gnd.n2658 gnd.n2657 19.3944
R9527 gnd.n2657 gnd.n2654 19.3944
R9528 gnd.n2654 gnd.n2653 19.3944
R9529 gnd.n2653 gnd.n2650 19.3944
R9530 gnd.n2650 gnd.n2649 19.3944
R9531 gnd.n2649 gnd.n2646 19.3944
R9532 gnd.n2646 gnd.n2645 19.3944
R9533 gnd.n2645 gnd.n2642 19.3944
R9534 gnd.n2642 gnd.n2641 19.3944
R9535 gnd.n2641 gnd.n2604 19.3944
R9536 gnd.n3030 gnd.n2961 19.3944
R9537 gnd.n3030 gnd.n2962 19.3944
R9538 gnd.n3026 gnd.n2962 19.3944
R9539 gnd.n3026 gnd.n1080 19.3944
R9540 gnd.n5040 gnd.n1080 19.3944
R9541 gnd.n5040 gnd.n5039 19.3944
R9542 gnd.n5039 gnd.n5038 19.3944
R9543 gnd.n5038 gnd.n1084 19.3944
R9544 gnd.n5028 gnd.n1084 19.3944
R9545 gnd.n5028 gnd.n5027 19.3944
R9546 gnd.n5027 gnd.n5026 19.3944
R9547 gnd.n5026 gnd.n1103 19.3944
R9548 gnd.n5016 gnd.n1103 19.3944
R9549 gnd.n5016 gnd.n5015 19.3944
R9550 gnd.n5015 gnd.n5014 19.3944
R9551 gnd.n5014 gnd.n1125 19.3944
R9552 gnd.n5004 gnd.n1125 19.3944
R9553 gnd.n5004 gnd.n5003 19.3944
R9554 gnd.n5003 gnd.n5002 19.3944
R9555 gnd.n5002 gnd.n1146 19.3944
R9556 gnd.n4992 gnd.n1146 19.3944
R9557 gnd.n4992 gnd.n4991 19.3944
R9558 gnd.n4991 gnd.n4990 19.3944
R9559 gnd.n4990 gnd.n1167 19.3944
R9560 gnd.n4980 gnd.n1167 19.3944
R9561 gnd.n4980 gnd.n4979 19.3944
R9562 gnd.n4979 gnd.n4978 19.3944
R9563 gnd.n4978 gnd.n1186 19.3944
R9564 gnd.n4967 gnd.n1186 19.3944
R9565 gnd.n4967 gnd.n4966 19.3944
R9566 gnd.n4966 gnd.n4965 19.3944
R9567 gnd.n4965 gnd.n1204 19.3944
R9568 gnd.n4955 gnd.n1204 19.3944
R9569 gnd.n4955 gnd.n4954 19.3944
R9570 gnd.n4954 gnd.n4953 19.3944
R9571 gnd.n4953 gnd.n1224 19.3944
R9572 gnd.n4943 gnd.n1224 19.3944
R9573 gnd.n4943 gnd.n4942 19.3944
R9574 gnd.n4942 gnd.n4941 19.3944
R9575 gnd.n4941 gnd.n1245 19.3944
R9576 gnd.n4931 gnd.n1245 19.3944
R9577 gnd.n4931 gnd.n4930 19.3944
R9578 gnd.n4930 gnd.n4929 19.3944
R9579 gnd.n4929 gnd.n1266 19.3944
R9580 gnd.n4919 gnd.n1266 19.3944
R9581 gnd.n4919 gnd.n4918 19.3944
R9582 gnd.n4918 gnd.n4917 19.3944
R9583 gnd.n4917 gnd.n1287 19.3944
R9584 gnd.n4907 gnd.n1287 19.3944
R9585 gnd.n4907 gnd.n4906 19.3944
R9586 gnd.n4906 gnd.n4905 19.3944
R9587 gnd.n4905 gnd.n1309 19.3944
R9588 gnd.n4895 gnd.n1309 19.3944
R9589 gnd.n3022 gnd.n3020 19.3944
R9590 gnd.n3020 gnd.n3017 19.3944
R9591 gnd.n3017 gnd.n3016 19.3944
R9592 gnd.n3016 gnd.n3013 19.3944
R9593 gnd.n3013 gnd.n3012 19.3944
R9594 gnd.n3012 gnd.n3009 19.3944
R9595 gnd.n3009 gnd.n3008 19.3944
R9596 gnd.n3008 gnd.n3005 19.3944
R9597 gnd.n3005 gnd.n3004 19.3944
R9598 gnd.n3004 gnd.n3001 19.3944
R9599 gnd.n3001 gnd.n3000 19.3944
R9600 gnd.n3000 gnd.n2997 19.3944
R9601 gnd.n2997 gnd.n2996 19.3944
R9602 gnd.n2996 gnd.n2993 19.3944
R9603 gnd.n2993 gnd.n2992 19.3944
R9604 gnd.n2992 gnd.n2989 19.3944
R9605 gnd.n2983 gnd.n2956 19.3944
R9606 gnd.n3041 gnd.n2956 19.3944
R9607 gnd.n3042 gnd.n3041 19.3944
R9608 gnd.n3044 gnd.n3042 19.3944
R9609 gnd.n3044 gnd.n2954 19.3944
R9610 gnd.n3049 gnd.n2954 19.3944
R9611 gnd.n3050 gnd.n3049 19.3944
R9612 gnd.n3052 gnd.n3050 19.3944
R9613 gnd.n3052 gnd.n2952 19.3944
R9614 gnd.n3057 gnd.n2952 19.3944
R9615 gnd.n3058 gnd.n3057 19.3944
R9616 gnd.n3081 gnd.n3058 19.3944
R9617 gnd.n3081 gnd.n2950 19.3944
R9618 gnd.n3085 gnd.n2950 19.3944
R9619 gnd.n3085 gnd.n2946 19.3944
R9620 gnd.n3097 gnd.n2946 19.3944
R9621 gnd.n3097 gnd.n2944 19.3944
R9622 gnd.n3101 gnd.n2944 19.3944
R9623 gnd.n3101 gnd.n2846 19.3944
R9624 gnd.n3113 gnd.n2846 19.3944
R9625 gnd.n3113 gnd.n2844 19.3944
R9626 gnd.n3117 gnd.n2844 19.3944
R9627 gnd.n3117 gnd.n2840 19.3944
R9628 gnd.n3129 gnd.n2840 19.3944
R9629 gnd.n3129 gnd.n2838 19.3944
R9630 gnd.n3134 gnd.n2838 19.3944
R9631 gnd.n3134 gnd.n2831 19.3944
R9632 gnd.n3147 gnd.n2831 19.3944
R9633 gnd.n3147 gnd.n2829 19.3944
R9634 gnd.n3151 gnd.n2829 19.3944
R9635 gnd.n3151 gnd.n2825 19.3944
R9636 gnd.n3163 gnd.n2825 19.3944
R9637 gnd.n3163 gnd.n2823 19.3944
R9638 gnd.n3167 gnd.n2823 19.3944
R9639 gnd.n3167 gnd.n2817 19.3944
R9640 gnd.n3179 gnd.n2817 19.3944
R9641 gnd.n3179 gnd.n2815 19.3944
R9642 gnd.n3183 gnd.n2815 19.3944
R9643 gnd.n3183 gnd.n2811 19.3944
R9644 gnd.n3196 gnd.n2811 19.3944
R9645 gnd.n3196 gnd.n2809 19.3944
R9646 gnd.n3200 gnd.n2809 19.3944
R9647 gnd.n3200 gnd.n2795 19.3944
R9648 gnd.n3235 gnd.n2795 19.3944
R9649 gnd.n3235 gnd.n2796 19.3944
R9650 gnd.n3231 gnd.n2796 19.3944
R9651 gnd.n3231 gnd.n3230 19.3944
R9652 gnd.n3230 gnd.n3229 19.3944
R9653 gnd.n3229 gnd.n2801 19.3944
R9654 gnd.n3225 gnd.n2801 19.3944
R9655 gnd.n3225 gnd.n2702 19.3944
R9656 gnd.n3526 gnd.n2702 19.3944
R9657 gnd.n3526 gnd.n2703 19.3944
R9658 gnd.n3036 gnd.n3032 19.3944
R9659 gnd.n3036 gnd.n1069 19.3944
R9660 gnd.n5046 gnd.n1069 19.3944
R9661 gnd.n5046 gnd.n5045 19.3944
R9662 gnd.n5045 gnd.n5044 19.3944
R9663 gnd.n5044 gnd.n1073 19.3944
R9664 gnd.n5034 gnd.n1073 19.3944
R9665 gnd.n5034 gnd.n5033 19.3944
R9666 gnd.n5033 gnd.n5032 19.3944
R9667 gnd.n5032 gnd.n1094 19.3944
R9668 gnd.n5022 gnd.n1094 19.3944
R9669 gnd.n5022 gnd.n5021 19.3944
R9670 gnd.n5021 gnd.n5020 19.3944
R9671 gnd.n5020 gnd.n1114 19.3944
R9672 gnd.n5010 gnd.n1114 19.3944
R9673 gnd.n5010 gnd.n5009 19.3944
R9674 gnd.n5009 gnd.n5008 19.3944
R9675 gnd.n5008 gnd.n1136 19.3944
R9676 gnd.n4998 gnd.n1136 19.3944
R9677 gnd.n4998 gnd.n4997 19.3944
R9678 gnd.n4997 gnd.n4996 19.3944
R9679 gnd.n4996 gnd.n1156 19.3944
R9680 gnd.n4986 gnd.n4985 19.3944
R9681 gnd.n4985 gnd.n4984 19.3944
R9682 gnd.n4974 gnd.n1192 19.3944
R9683 gnd.n4972 gnd.n4971 19.3944
R9684 gnd.n4961 gnd.n1211 19.3944
R9685 gnd.n4961 gnd.n4960 19.3944
R9686 gnd.n4960 gnd.n4959 19.3944
R9687 gnd.n4959 gnd.n1214 19.3944
R9688 gnd.n4949 gnd.n1214 19.3944
R9689 gnd.n4949 gnd.n4948 19.3944
R9690 gnd.n4948 gnd.n4947 19.3944
R9691 gnd.n4947 gnd.n1234 19.3944
R9692 gnd.n4937 gnd.n1234 19.3944
R9693 gnd.n4937 gnd.n4936 19.3944
R9694 gnd.n4936 gnd.n4935 19.3944
R9695 gnd.n4935 gnd.n1256 19.3944
R9696 gnd.n4925 gnd.n1256 19.3944
R9697 gnd.n4925 gnd.n4924 19.3944
R9698 gnd.n4924 gnd.n4923 19.3944
R9699 gnd.n4923 gnd.n1276 19.3944
R9700 gnd.n4913 gnd.n1276 19.3944
R9701 gnd.n4913 gnd.n4912 19.3944
R9702 gnd.n4912 gnd.n4911 19.3944
R9703 gnd.n4911 gnd.n1298 19.3944
R9704 gnd.n4901 gnd.n1298 19.3944
R9705 gnd.n4901 gnd.n4900 19.3944
R9706 gnd.n4900 gnd.n4899 19.3944
R9707 gnd.n6690 gnd.n6689 19.3944
R9708 gnd.n6689 gnd.n6688 19.3944
R9709 gnd.n6688 gnd.n745 19.3944
R9710 gnd.n6682 gnd.n745 19.3944
R9711 gnd.n6682 gnd.n6681 19.3944
R9712 gnd.n6681 gnd.n6680 19.3944
R9713 gnd.n6680 gnd.n753 19.3944
R9714 gnd.n6674 gnd.n753 19.3944
R9715 gnd.n6674 gnd.n6673 19.3944
R9716 gnd.n6673 gnd.n6672 19.3944
R9717 gnd.n6672 gnd.n761 19.3944
R9718 gnd.n6666 gnd.n761 19.3944
R9719 gnd.n6666 gnd.n6665 19.3944
R9720 gnd.n6665 gnd.n6664 19.3944
R9721 gnd.n6664 gnd.n769 19.3944
R9722 gnd.n6658 gnd.n769 19.3944
R9723 gnd.n6658 gnd.n6657 19.3944
R9724 gnd.n6657 gnd.n6656 19.3944
R9725 gnd.n6656 gnd.n777 19.3944
R9726 gnd.n6650 gnd.n777 19.3944
R9727 gnd.n6650 gnd.n6649 19.3944
R9728 gnd.n6649 gnd.n6648 19.3944
R9729 gnd.n6648 gnd.n785 19.3944
R9730 gnd.n6642 gnd.n785 19.3944
R9731 gnd.n6642 gnd.n6641 19.3944
R9732 gnd.n6641 gnd.n6640 19.3944
R9733 gnd.n6640 gnd.n793 19.3944
R9734 gnd.n6634 gnd.n793 19.3944
R9735 gnd.n6634 gnd.n6633 19.3944
R9736 gnd.n6633 gnd.n6632 19.3944
R9737 gnd.n6632 gnd.n801 19.3944
R9738 gnd.n6626 gnd.n801 19.3944
R9739 gnd.n6626 gnd.n6625 19.3944
R9740 gnd.n6625 gnd.n6624 19.3944
R9741 gnd.n6624 gnd.n809 19.3944
R9742 gnd.n6618 gnd.n809 19.3944
R9743 gnd.n6618 gnd.n6617 19.3944
R9744 gnd.n6617 gnd.n6616 19.3944
R9745 gnd.n6616 gnd.n817 19.3944
R9746 gnd.n6610 gnd.n817 19.3944
R9747 gnd.n6610 gnd.n6609 19.3944
R9748 gnd.n6609 gnd.n6608 19.3944
R9749 gnd.n6608 gnd.n825 19.3944
R9750 gnd.n6602 gnd.n825 19.3944
R9751 gnd.n6602 gnd.n6601 19.3944
R9752 gnd.n6601 gnd.n6600 19.3944
R9753 gnd.n6600 gnd.n833 19.3944
R9754 gnd.n6594 gnd.n833 19.3944
R9755 gnd.n6594 gnd.n6593 19.3944
R9756 gnd.n6593 gnd.n6592 19.3944
R9757 gnd.n6592 gnd.n841 19.3944
R9758 gnd.n6586 gnd.n841 19.3944
R9759 gnd.n6586 gnd.n6585 19.3944
R9760 gnd.n6585 gnd.n6584 19.3944
R9761 gnd.n6584 gnd.n849 19.3944
R9762 gnd.n6578 gnd.n849 19.3944
R9763 gnd.n6578 gnd.n6577 19.3944
R9764 gnd.n6577 gnd.n6576 19.3944
R9765 gnd.n6576 gnd.n857 19.3944
R9766 gnd.n6570 gnd.n857 19.3944
R9767 gnd.n6570 gnd.n6569 19.3944
R9768 gnd.n6569 gnd.n6568 19.3944
R9769 gnd.n6568 gnd.n865 19.3944
R9770 gnd.n6562 gnd.n865 19.3944
R9771 gnd.n6562 gnd.n6561 19.3944
R9772 gnd.n6561 gnd.n6560 19.3944
R9773 gnd.n6560 gnd.n873 19.3944
R9774 gnd.n6554 gnd.n873 19.3944
R9775 gnd.n6554 gnd.n6553 19.3944
R9776 gnd.n6553 gnd.n6552 19.3944
R9777 gnd.n6552 gnd.n881 19.3944
R9778 gnd.n6546 gnd.n881 19.3944
R9779 gnd.n6546 gnd.n6545 19.3944
R9780 gnd.n6545 gnd.n6544 19.3944
R9781 gnd.n6544 gnd.n889 19.3944
R9782 gnd.n6538 gnd.n889 19.3944
R9783 gnd.n6538 gnd.n6537 19.3944
R9784 gnd.n6537 gnd.n6536 19.3944
R9785 gnd.n6536 gnd.n897 19.3944
R9786 gnd.n6530 gnd.n897 19.3944
R9787 gnd.n6530 gnd.n6529 19.3944
R9788 gnd.n6529 gnd.n6528 19.3944
R9789 gnd.n6528 gnd.n905 19.3944
R9790 gnd.n2860 gnd.n905 19.3944
R9791 gnd.n4890 gnd.n4889 19.3944
R9792 gnd.n4889 gnd.n4888 19.3944
R9793 gnd.n4888 gnd.n1332 19.3944
R9794 gnd.n4884 gnd.n1332 19.3944
R9795 gnd.n4884 gnd.n4883 19.3944
R9796 gnd.n4883 gnd.n4882 19.3944
R9797 gnd.n4882 gnd.n1337 19.3944
R9798 gnd.n4878 gnd.n1337 19.3944
R9799 gnd.n4878 gnd.n4877 19.3944
R9800 gnd.n4877 gnd.n4876 19.3944
R9801 gnd.n4876 gnd.n1342 19.3944
R9802 gnd.n4872 gnd.n1342 19.3944
R9803 gnd.n4872 gnd.n4871 19.3944
R9804 gnd.n4871 gnd.n4870 19.3944
R9805 gnd.n4870 gnd.n1347 19.3944
R9806 gnd.n4866 gnd.n1347 19.3944
R9807 gnd.n4866 gnd.n4865 19.3944
R9808 gnd.n4865 gnd.n4864 19.3944
R9809 gnd.n4864 gnd.n1352 19.3944
R9810 gnd.n4860 gnd.n1352 19.3944
R9811 gnd.n4860 gnd.n4859 19.3944
R9812 gnd.n4859 gnd.n4858 19.3944
R9813 gnd.n4858 gnd.n1357 19.3944
R9814 gnd.n4854 gnd.n1357 19.3944
R9815 gnd.n4854 gnd.n4853 19.3944
R9816 gnd.n4853 gnd.n4852 19.3944
R9817 gnd.n4852 gnd.n1362 19.3944
R9818 gnd.n4848 gnd.n1362 19.3944
R9819 gnd.n4848 gnd.n4847 19.3944
R9820 gnd.n4847 gnd.n4846 19.3944
R9821 gnd.n4846 gnd.n1367 19.3944
R9822 gnd.n4842 gnd.n1367 19.3944
R9823 gnd.n4842 gnd.n4841 19.3944
R9824 gnd.n4841 gnd.n4840 19.3944
R9825 gnd.n4840 gnd.n1372 19.3944
R9826 gnd.n4836 gnd.n1372 19.3944
R9827 gnd.n4836 gnd.n4835 19.3944
R9828 gnd.n4835 gnd.n4834 19.3944
R9829 gnd.n4834 gnd.n1377 19.3944
R9830 gnd.n4830 gnd.n1377 19.3944
R9831 gnd.n4830 gnd.n4829 19.3944
R9832 gnd.n4829 gnd.n4828 19.3944
R9833 gnd.n4828 gnd.n1382 19.3944
R9834 gnd.n4824 gnd.n1382 19.3944
R9835 gnd.n4824 gnd.n4823 19.3944
R9836 gnd.n4823 gnd.n4822 19.3944
R9837 gnd.n4822 gnd.n1387 19.3944
R9838 gnd.n4818 gnd.n1387 19.3944
R9839 gnd.n4818 gnd.n4817 19.3944
R9840 gnd.n4817 gnd.n4816 19.3944
R9841 gnd.n4816 gnd.n1392 19.3944
R9842 gnd.n4812 gnd.n1392 19.3944
R9843 gnd.n4812 gnd.n4811 19.3944
R9844 gnd.n4811 gnd.n4810 19.3944
R9845 gnd.n4810 gnd.n1397 19.3944
R9846 gnd.n4806 gnd.n1397 19.3944
R9847 gnd.n4806 gnd.n4805 19.3944
R9848 gnd.n4805 gnd.n4804 19.3944
R9849 gnd.n4804 gnd.n1402 19.3944
R9850 gnd.n4800 gnd.n1402 19.3944
R9851 gnd.n4800 gnd.n4799 19.3944
R9852 gnd.n4799 gnd.n4798 19.3944
R9853 gnd.n4798 gnd.n1407 19.3944
R9854 gnd.n4794 gnd.n1407 19.3944
R9855 gnd.n4794 gnd.n4793 19.3944
R9856 gnd.n4793 gnd.n4792 19.3944
R9857 gnd.n4792 gnd.n1412 19.3944
R9858 gnd.n4788 gnd.n1412 19.3944
R9859 gnd.n4788 gnd.n4787 19.3944
R9860 gnd.n4787 gnd.n4786 19.3944
R9861 gnd.n4786 gnd.n1417 19.3944
R9862 gnd.n4782 gnd.n1417 19.3944
R9863 gnd.n4782 gnd.n4781 19.3944
R9864 gnd.n4781 gnd.n4780 19.3944
R9865 gnd.n4780 gnd.n1422 19.3944
R9866 gnd.n4776 gnd.n1422 19.3944
R9867 gnd.n4776 gnd.n4775 19.3944
R9868 gnd.n4775 gnd.n4774 19.3944
R9869 gnd.n4774 gnd.n1427 19.3944
R9870 gnd.n4770 gnd.n1427 19.3944
R9871 gnd.n4770 gnd.n4769 19.3944
R9872 gnd.n4769 gnd.n4768 19.3944
R9873 gnd.n4768 gnd.n1432 19.3944
R9874 gnd.n4764 gnd.n1432 19.3944
R9875 gnd.n4764 gnd.n4763 19.3944
R9876 gnd.n4763 gnd.n4762 19.3944
R9877 gnd.n4762 gnd.n1437 19.3944
R9878 gnd.n4758 gnd.n1437 19.3944
R9879 gnd.n4758 gnd.n4757 19.3944
R9880 gnd.n4757 gnd.n4756 19.3944
R9881 gnd.n4756 gnd.n1442 19.3944
R9882 gnd.n4752 gnd.n1442 19.3944
R9883 gnd.n4752 gnd.n4751 19.3944
R9884 gnd.n4751 gnd.n4750 19.3944
R9885 gnd.n4750 gnd.n1447 19.3944
R9886 gnd.n4746 gnd.n1447 19.3944
R9887 gnd.n4746 gnd.n4745 19.3944
R9888 gnd.n4745 gnd.n4744 19.3944
R9889 gnd.n4744 gnd.n1452 19.3944
R9890 gnd.n4740 gnd.n1452 19.3944
R9891 gnd.n4740 gnd.n4739 19.3944
R9892 gnd.n4459 gnd.n4458 19.3944
R9893 gnd.n4458 gnd.n4457 19.3944
R9894 gnd.n4457 gnd.n1799 19.3944
R9895 gnd.n1701 gnd.n1697 19.3944
R9896 gnd.n1701 gnd.n1679 19.3944
R9897 gnd.n1714 gnd.n1679 19.3944
R9898 gnd.n1714 gnd.n1677 19.3944
R9899 gnd.n1720 gnd.n1677 19.3944
R9900 gnd.n1720 gnd.n1670 19.3944
R9901 gnd.n1733 gnd.n1670 19.3944
R9902 gnd.n1733 gnd.n1668 19.3944
R9903 gnd.n1739 gnd.n1668 19.3944
R9904 gnd.n1739 gnd.n1661 19.3944
R9905 gnd.n1752 gnd.n1661 19.3944
R9906 gnd.n1752 gnd.n1659 19.3944
R9907 gnd.n1758 gnd.n1659 19.3944
R9908 gnd.n1758 gnd.n1652 19.3944
R9909 gnd.n1771 gnd.n1652 19.3944
R9910 gnd.n1771 gnd.n1650 19.3944
R9911 gnd.n4471 gnd.n1650 19.3944
R9912 gnd.n4471 gnd.n4470 19.3944
R9913 gnd.n4470 gnd.n4469 19.3944
R9914 gnd.n4469 gnd.n1779 19.3944
R9915 gnd.n4465 gnd.n1779 19.3944
R9916 gnd.n4465 gnd.n4464 19.3944
R9917 gnd.n4464 gnd.n4463 19.3944
R9918 gnd.n4463 gnd.n1787 19.3944
R9919 gnd.n3642 gnd.n3641 19.2005
R9920 gnd.n4296 gnd.n4295 19.2005
R9921 gnd.n5895 gnd.t80 18.8012
R9922 gnd.n5934 gnd.t318 18.8012
R9923 gnd.n5738 gnd.n5480 18.4825
R9924 gnd.n2030 gnd.n1889 18.4247
R9925 gnd.n3573 gnd.n2604 18.4247
R9926 gnd.n7617 gnd.n7616 18.2308
R9927 gnd.n1767 gnd.n1647 18.2308
R9928 gnd.n3357 gnd.n3341 18.2308
R9929 gnd.n2989 gnd.n2981 18.2308
R9930 gnd.t79 gnd.n5422 18.1639
R9931 gnd.n5451 gnd.t88 17.5266
R9932 gnd.t19 gnd.n1077 17.5266
R9933 gnd.n7569 gnd.t17 17.5266
R9934 gnd.t66 gnd.n5398 16.8893
R9935 gnd.n3087 gnd.t13 16.8893
R9936 gnd.n7537 gnd.t42 16.8893
R9937 gnd.t224 gnd.n5507 16.2519
R9938 gnd.n5365 gnd.t137 16.2519
R9939 gnd.n3119 gnd.t47 16.2519
R9940 gnd.n7505 gnd.t49 16.2519
R9941 gnd.n3407 gnd.n3406 15.9333
R9942 gnd.n3408 gnd.n3407 15.9333
R9943 gnd.n3409 gnd.n3408 15.9333
R9944 gnd.n3412 gnd.n3409 15.9333
R9945 gnd.n3411 gnd.n3410 15.9333
R9946 gnd.n3410 gnd.n2769 15.9333
R9947 gnd.n3420 gnd.n2769 15.9333
R9948 gnd.n3421 gnd.n3420 15.9333
R9949 gnd.n3422 gnd.n3421 15.9333
R9950 gnd.n3423 gnd.n3422 15.9333
R9951 gnd.n3426 gnd.n3423 15.9333
R9952 gnd.n3426 gnd.n3425 15.9333
R9953 gnd.n3425 gnd.n3424 15.9333
R9954 gnd.n3434 gnd.n2761 15.9333
R9955 gnd.n3435 gnd.n3434 15.9333
R9956 gnd.n3436 gnd.n3435 15.9333
R9957 gnd.n3437 gnd.n3436 15.9333
R9958 gnd.n3443 gnd.n3437 15.9333
R9959 gnd.n3443 gnd.n3442 15.9333
R9960 gnd.n3442 gnd.n3441 15.9333
R9961 gnd.n3441 gnd.n3440 15.9333
R9962 gnd.n3452 gnd.n3451 15.9333
R9963 gnd.n3453 gnd.n3452 15.9333
R9964 gnd.n3454 gnd.n3453 15.9333
R9965 gnd.n3457 gnd.n3454 15.9333
R9966 gnd.n3457 gnd.n3456 15.9333
R9967 gnd.n3456 gnd.n3455 15.9333
R9968 gnd.n3455 gnd.n2747 15.9333
R9969 gnd.n3467 gnd.n2747 15.9333
R9970 gnd.n3468 gnd.n2427 15.9333
R9971 gnd.n3471 gnd.n2460 15.9333
R9972 gnd.n2532 gnd.n2403 15.9333
R9973 gnd.n3673 gnd.n2370 15.9333
R9974 gnd.n3705 gnd.n3704 15.9333
R9975 gnd.n2510 gnd.n2344 15.9333
R9976 gnd.n2500 gnd.n2340 15.9333
R9977 gnd.n3749 gnd.n3748 15.9333
R9978 gnd.n3827 gnd.n3826 15.9333
R9979 gnd.n3853 gnd.n3852 15.9333
R9980 gnd.n3879 gnd.n2227 15.9333
R9981 gnd.n3889 gnd.n3888 15.9333
R9982 gnd.n2243 gnd.n2214 15.9333
R9983 gnd.n3915 gnd.n3914 15.9333
R9984 gnd.n3937 gnd.n2178 15.9333
R9985 gnd.n3991 gnd.n2163 15.9333
R9986 gnd.n4074 gnd.n2116 15.9333
R9987 gnd.n4088 gnd.n4087 15.9333
R9988 gnd.n2108 gnd.n2091 15.9333
R9989 gnd.n4148 gnd.n2081 15.9333
R9990 gnd.n4159 gnd.n4158 15.9333
R9991 gnd.n4204 gnd.n2044 15.9333
R9992 gnd.n2037 gnd.n1852 15.9333
R9993 gnd.n4367 gnd.n1852 15.9333
R9994 gnd.n1871 gnd.n1870 15.9333
R9995 gnd.n4377 gnd.n4376 15.9333
R9996 gnd.n4376 gnd.n4375 15.9333
R9997 gnd.n4375 gnd.n1841 15.9333
R9998 gnd.n4385 gnd.n1841 15.9333
R9999 gnd.n4387 gnd.n4385 15.9333
R10000 gnd.n4387 gnd.n4386 15.9333
R10001 gnd.n4386 gnd.n1834 15.9333
R10002 gnd.n4397 gnd.n1834 15.9333
R10003 gnd.n4396 gnd.n4395 15.9333
R10004 gnd.n4395 gnd.n1828 15.9333
R10005 gnd.n4405 gnd.n1828 15.9333
R10006 gnd.n4407 gnd.n4405 15.9333
R10007 gnd.n4407 gnd.n4406 15.9333
R10008 gnd.n4406 gnd.n1821 15.9333
R10009 gnd.n4417 gnd.n1821 15.9333
R10010 gnd.n4417 gnd.n4416 15.9333
R10011 gnd.n4415 gnd.n1815 15.9333
R10012 gnd.n4425 gnd.n1815 15.9333
R10013 gnd.n4427 gnd.n4425 15.9333
R10014 gnd.n4427 gnd.n4426 15.9333
R10015 gnd.n4426 gnd.n1808 15.9333
R10016 gnd.n4440 gnd.n1808 15.9333
R10017 gnd.n4440 gnd.n4439 15.9333
R10018 gnd.n4439 gnd.n4438 15.9333
R10019 gnd.n4438 gnd.n4437 15.9333
R10020 gnd.n4450 gnd.n4449 15.9333
R10021 gnd.n4450 gnd.n1456 15.9333
R10022 gnd.n4737 gnd.n1456 15.9333
R10023 gnd.n4737 gnd.n4736 15.9333
R10024 gnd.n6357 gnd.n6355 15.6674
R10025 gnd.n6325 gnd.n6323 15.6674
R10026 gnd.n6293 gnd.n6291 15.6674
R10027 gnd.n6262 gnd.n6260 15.6674
R10028 gnd.n6230 gnd.n6228 15.6674
R10029 gnd.n6198 gnd.n6196 15.6674
R10030 gnd.n6166 gnd.n6164 15.6674
R10031 gnd.n6135 gnd.n6133 15.6674
R10032 gnd.n5625 gnd.t224 15.6146
R10033 gnd.n6395 gnd.t183 15.6146
R10034 gnd.n6496 gnd.t199 15.6146
R10035 gnd.n3153 gnd.t114 15.6146
R10036 gnd.n4634 gnd.t74 15.6146
R10037 gnd.n3739 gnd.n2325 15.296
R10038 gnd.n2319 gnd.n2309 15.296
R10039 gnd.n3777 gnd.t107 15.296
R10040 gnd.n3890 gnd.n2218 15.296
R10041 gnd.n2244 gnd.n2204 15.296
R10042 gnd.n4042 gnd.t108 15.296
R10043 gnd.n4051 gnd.n2125 15.296
R10044 gnd.n4073 gnd.n2118 15.296
R10045 gnd.t210 gnd.n4190 15.296
R10046 gnd.n4213 gnd.n4212 15.0827
R10047 gnd.n2413 gnd.n2408 15.0481
R10048 gnd.n4223 gnd.n4222 15.0481
R10049 gnd.n6061 gnd.t148 14.9773
R10050 gnd.n3185 gnd.t33 14.9773
R10051 gnd.t96 gnd.n1289 14.9773
R10052 gnd.n3637 gnd.n2427 14.9773
R10053 gnd.n4535 gnd.t72 14.9773
R10054 gnd.n4596 gnd.t56 14.9773
R10055 gnd.t263 gnd.n3471 14.6587
R10056 gnd.n3713 gnd.n2352 14.6587
R10057 gnd.n2477 gnd.n2290 14.6587
R10058 gnd.n4002 gnd.n4001 14.6587
R10059 gnd.n4140 gnd.n4139 14.6587
R10060 gnd.n4124 gnd.t207 14.6587
R10061 gnd.n4125 gnd.n2060 14.6587
R10062 gnd.t105 gnd.n6099 14.34
R10063 gnd.n6117 gnd.t89 14.34
R10064 gnd.n5036 gnd.t19 14.34
R10065 gnd.t33 gnd.n1247 14.34
R10066 gnd.n3210 gnd.t96 14.34
R10067 gnd.t72 gnd.n4534 14.34
R10068 gnd.n1583 gnd.t56 14.34
R10069 gnd.n211 gnd.t17 14.34
R10070 gnd.n3675 gnd.t238 14.0214
R10071 gnd.n3731 gnd.n3730 14.0214
R10072 gnd.n3776 gnd.n2304 14.0214
R10073 gnd.n3871 gnd.n3869 14.0214
R10074 gnd.n3913 gnd.n2199 14.0214
R10075 gnd.n4032 gnd.n2131 14.0214
R10076 gnd.n4098 gnd.n2099 14.0214
R10077 gnd.n4205 gnd.n2042 14.0214
R10078 gnd.t70 gnd.n5822 13.7027
R10079 gnd.t114 gnd.n1206 13.7027
R10080 gnd.n3805 gnd.t293 13.7027
R10081 gnd.t323 gnd.n2174 13.7027
R10082 gnd.t74 gnd.n280 13.7027
R10083 gnd.n117 gnd.n106 13.7027
R10084 gnd.n5707 gnd.n5703 13.5763
R10085 gnd.n6459 gnd.n5157 13.5763
R10086 gnd.n1991 gnd.n1979 13.5763
R10087 gnd.n7669 gnd.n7668 13.5763
R10088 gnd.n5062 gnd.n1055 13.5763
R10089 gnd.n3539 gnd.n2696 13.5763
R10090 gnd.n5739 gnd.n5738 13.384
R10091 gnd.n3654 gnd.n2386 13.384
R10092 gnd.n3724 gnd.n3723 13.384
R10093 gnd.n3789 gnd.n2294 13.384
R10094 gnd.t68 gnd.n3787 13.384
R10095 gnd.t69 gnd.n2150 13.384
R10096 gnd.n3968 gnd.n2140 13.384
R10097 gnd.n2110 gnd.n2109 13.384
R10098 gnd.n4189 gnd.n2056 13.384
R10099 gnd.n2424 gnd.n2405 13.1884
R10100 gnd.n2419 gnd.n2418 13.1884
R10101 gnd.n2418 gnd.n2417 13.1884
R10102 gnd.n4216 gnd.n4211 13.1884
R10103 gnd.n4217 gnd.n4216 13.1884
R10104 gnd.n2420 gnd.n2407 13.146
R10105 gnd.n2416 gnd.n2407 13.146
R10106 gnd.n4215 gnd.n4214 13.146
R10107 gnd.n4215 gnd.n4210 13.146
R10108 gnd.t47 gnd.n1169 13.0654
R10109 gnd.n2518 gnd.t84 13.0654
R10110 gnd.n4132 gnd.t7 13.0654
R10111 gnd.n7470 gnd.t49 13.0654
R10112 gnd.n6358 gnd.n6354 12.8005
R10113 gnd.n6326 gnd.n6322 12.8005
R10114 gnd.n6294 gnd.n6290 12.8005
R10115 gnd.n6263 gnd.n6259 12.8005
R10116 gnd.n6231 gnd.n6227 12.8005
R10117 gnd.n6199 gnd.n6195 12.8005
R10118 gnd.n6167 gnd.n6163 12.8005
R10119 gnd.n6136 gnd.n6132 12.8005
R10120 gnd.n3662 gnd.n2388 12.7467
R10121 gnd.n3694 gnd.t248 12.7467
R10122 gnd.n2511 gnd.n2509 12.7467
R10123 gnd.n2262 gnd.n2256 12.7467
R10124 gnd.n3952 gnd.n3951 12.7467
R10125 gnd.n4111 gnd.n4110 12.7467
R10126 gnd.t13 gnd.n1127 12.4281
R10127 gnd.t29 gnd.n2761 12.4281
R10128 gnd.n4416 gnd.t287 12.4281
R10129 gnd.n7455 gnd.t42 12.4281
R10130 gnd.n5710 gnd.n5707 12.4126
R10131 gnd.n6462 gnd.n6459 12.4126
R10132 gnd.n1987 gnd.n1979 12.4126
R10133 gnd.n7668 gnd.n179 12.4126
R10134 gnd.n5058 gnd.n1055 12.4126
R10135 gnd.n3534 gnd.n2696 12.4126
R10136 gnd.n3641 gnd.n3640 12.1761
R10137 gnd.n4295 gnd.n4294 12.1761
R10138 gnd.n3646 gnd.n3645 12.1094
R10139 gnd.t218 gnd.n2393 12.1094
R10140 gnd.n2501 gnd.n2332 12.1094
R10141 gnd.n3769 gnd.n3768 12.1094
R10142 gnd.n4040 gnd.n2134 12.1094
R10143 gnd.n4089 gnd.n2105 12.1094
R10144 gnd.n2047 gnd.n2046 12.1094
R10145 gnd.n6362 gnd.n6361 12.0247
R10146 gnd.n6330 gnd.n6329 12.0247
R10147 gnd.n6298 gnd.n6297 12.0247
R10148 gnd.n6267 gnd.n6266 12.0247
R10149 gnd.n6235 gnd.n6234 12.0247
R10150 gnd.n6203 gnd.n6202 12.0247
R10151 gnd.n6171 gnd.n6170 12.0247
R10152 gnd.n6140 gnd.n6139 12.0247
R10153 gnd.n3688 gnd.n3687 11.4721
R10154 gnd.n3706 gnd.n2357 11.4721
R10155 gnd.t138 gnd.n2281 11.4721
R10156 gnd.n3820 gnd.n3819 11.4721
R10157 gnd.n3838 gnd.n2268 11.4721
R10158 gnd.n2182 gnd.n2169 11.4721
R10159 gnd.n3976 gnd.n2165 11.4721
R10160 gnd.n3975 gnd.t25 11.4721
R10161 gnd.n4147 gnd.n2084 11.4721
R10162 gnd.n4166 gnd.n4165 11.4721
R10163 gnd.n6365 gnd.n6352 11.249
R10164 gnd.n6333 gnd.n6320 11.249
R10165 gnd.n6301 gnd.n6288 11.249
R10166 gnd.n6270 gnd.n6257 11.249
R10167 gnd.n6238 gnd.n6225 11.249
R10168 gnd.n6206 gnd.n6193 11.249
R10169 gnd.n6174 gnd.n6161 11.249
R10170 gnd.n6143 gnd.n6130 11.249
R10171 gnd.n5823 gnd.t70 11.1535
R10172 gnd.t0 gnd.n3467 11.1535
R10173 gnd.n2296 gnd.t308 11.1535
R10174 gnd.t37 gnd.n4008 11.1535
R10175 gnd.n4377 gnd.t5 11.1535
R10176 gnd.n3747 gnd.n2327 10.8348
R10177 gnd.n2492 gnd.n2327 10.8348
R10178 gnd.n3897 gnd.n2211 10.8348
R10179 gnd.n3897 gnd.n3896 10.8348
R10180 gnd.n4067 gnd.n4066 10.8348
R10181 gnd.n4066 gnd.n4065 10.8348
R10182 gnd.n4363 gnd.n4362 10.6151
R10183 gnd.n4362 gnd.n4359 10.6151
R10184 gnd.n4357 gnd.n4354 10.6151
R10185 gnd.n4354 gnd.n4353 10.6151
R10186 gnd.n4353 gnd.n4350 10.6151
R10187 gnd.n4350 gnd.n4349 10.6151
R10188 gnd.n4349 gnd.n4346 10.6151
R10189 gnd.n4346 gnd.n4345 10.6151
R10190 gnd.n4345 gnd.n4342 10.6151
R10191 gnd.n4342 gnd.n4341 10.6151
R10192 gnd.n4341 gnd.n4338 10.6151
R10193 gnd.n4338 gnd.n4337 10.6151
R10194 gnd.n4337 gnd.n4334 10.6151
R10195 gnd.n4334 gnd.n4333 10.6151
R10196 gnd.n4333 gnd.n4330 10.6151
R10197 gnd.n4330 gnd.n4329 10.6151
R10198 gnd.n4329 gnd.n4326 10.6151
R10199 gnd.n4326 gnd.n4325 10.6151
R10200 gnd.n4325 gnd.n4322 10.6151
R10201 gnd.n4322 gnd.n4321 10.6151
R10202 gnd.n4321 gnd.n4318 10.6151
R10203 gnd.n4318 gnd.n4317 10.6151
R10204 gnd.n4317 gnd.n4314 10.6151
R10205 gnd.n4314 gnd.n4313 10.6151
R10206 gnd.n4313 gnd.n4310 10.6151
R10207 gnd.n4310 gnd.n4309 10.6151
R10208 gnd.n4309 gnd.n4306 10.6151
R10209 gnd.n4306 gnd.n4305 10.6151
R10210 gnd.n4305 gnd.n4302 10.6151
R10211 gnd.n4302 gnd.n4301 10.6151
R10212 gnd.n2537 gnd.n2536 10.6151
R10213 gnd.n2536 gnd.n2535 10.6151
R10214 gnd.n2535 gnd.n2531 10.6151
R10215 gnd.n2531 gnd.n2530 10.6151
R10216 gnd.n2530 gnd.n2528 10.6151
R10217 gnd.n2528 gnd.n2527 10.6151
R10218 gnd.n2527 gnd.n2525 10.6151
R10219 gnd.n2525 gnd.n2524 10.6151
R10220 gnd.n2524 gnd.n2523 10.6151
R10221 gnd.n2523 gnd.n2522 10.6151
R10222 gnd.n2522 gnd.n2521 10.6151
R10223 gnd.n2521 gnd.n2517 10.6151
R10224 gnd.n2517 gnd.n2516 10.6151
R10225 gnd.n2516 gnd.n2514 10.6151
R10226 gnd.n2514 gnd.n2513 10.6151
R10227 gnd.n2513 gnd.n2508 10.6151
R10228 gnd.n2508 gnd.n2507 10.6151
R10229 gnd.n2507 gnd.n2504 10.6151
R10230 gnd.n2504 gnd.n2503 10.6151
R10231 gnd.n2503 gnd.n2498 10.6151
R10232 gnd.n2498 gnd.n2497 10.6151
R10233 gnd.n2497 gnd.n2495 10.6151
R10234 gnd.n2495 gnd.n2494 10.6151
R10235 gnd.n2494 gnd.n2490 10.6151
R10236 gnd.n2490 gnd.n2489 10.6151
R10237 gnd.n2489 gnd.n2488 10.6151
R10238 gnd.n2488 gnd.n2487 10.6151
R10239 gnd.n2487 gnd.n2486 10.6151
R10240 gnd.n2486 gnd.n2483 10.6151
R10241 gnd.n2483 gnd.n2482 10.6151
R10242 gnd.n2482 gnd.n2480 10.6151
R10243 gnd.n2480 gnd.n2479 10.6151
R10244 gnd.n2479 gnd.n2475 10.6151
R10245 gnd.n2475 gnd.n2474 10.6151
R10246 gnd.n2474 gnd.n2472 10.6151
R10247 gnd.n2472 gnd.n2471 10.6151
R10248 gnd.n2471 gnd.n2467 10.6151
R10249 gnd.n2467 gnd.n2259 10.6151
R10250 gnd.n3847 gnd.n2259 10.6151
R10251 gnd.n3848 gnd.n3847 10.6151
R10252 gnd.n3849 gnd.n3848 10.6151
R10253 gnd.n3849 gnd.n2234 10.6151
R10254 gnd.n3867 gnd.n2234 10.6151
R10255 gnd.n3867 gnd.n3866 10.6151
R10256 gnd.n3866 gnd.n3865 10.6151
R10257 gnd.n3865 gnd.n2250 10.6151
R10258 gnd.n2250 gnd.n2249 10.6151
R10259 gnd.n2249 gnd.n2247 10.6151
R10260 gnd.n2247 gnd.n2246 10.6151
R10261 gnd.n2246 gnd.n2242 10.6151
R10262 gnd.n2242 gnd.n2241 10.6151
R10263 gnd.n2241 gnd.n2239 10.6151
R10264 gnd.n2239 gnd.n2238 10.6151
R10265 gnd.n2238 gnd.n2236 10.6151
R10266 gnd.n2236 gnd.n2235 10.6151
R10267 gnd.n2235 gnd.n2172 10.6151
R10268 gnd.n3960 gnd.n2172 10.6151
R10269 gnd.n3961 gnd.n3960 10.6151
R10270 gnd.n3981 gnd.n3961 10.6151
R10271 gnd.n3981 gnd.n3980 10.6151
R10272 gnd.n3980 gnd.n3979 10.6151
R10273 gnd.n3979 gnd.n3978 10.6151
R10274 gnd.n3978 gnd.n3974 10.6151
R10275 gnd.n3974 gnd.n3973 10.6151
R10276 gnd.n3973 gnd.n3971 10.6151
R10277 gnd.n3971 gnd.n3970 10.6151
R10278 gnd.n3970 gnd.n3965 10.6151
R10279 gnd.n3965 gnd.n3964 10.6151
R10280 gnd.n3964 gnd.n3962 10.6151
R10281 gnd.n3962 gnd.n2123 10.6151
R10282 gnd.n4053 gnd.n2123 10.6151
R10283 gnd.n4054 gnd.n4053 10.6151
R10284 gnd.n4063 gnd.n4054 10.6151
R10285 gnd.n4063 gnd.n4062 10.6151
R10286 gnd.n4062 gnd.n4061 10.6151
R10287 gnd.n4061 gnd.n4058 10.6151
R10288 gnd.n4058 gnd.n4057 10.6151
R10289 gnd.n4057 gnd.n4055 10.6151
R10290 gnd.n4055 gnd.n2089 10.6151
R10291 gnd.n4113 gnd.n2089 10.6151
R10292 gnd.n4114 gnd.n4113 10.6151
R10293 gnd.n4137 gnd.n4114 10.6151
R10294 gnd.n4137 gnd.n4136 10.6151
R10295 gnd.n4136 gnd.n4135 10.6151
R10296 gnd.n4135 gnd.n4131 10.6151
R10297 gnd.n4131 gnd.n4130 10.6151
R10298 gnd.n4130 gnd.n4128 10.6151
R10299 gnd.n4128 gnd.n4127 10.6151
R10300 gnd.n4127 gnd.n4123 10.6151
R10301 gnd.n4123 gnd.n4122 10.6151
R10302 gnd.n4122 gnd.n4120 10.6151
R10303 gnd.n4120 gnd.n4119 10.6151
R10304 gnd.n4119 gnd.n4116 10.6151
R10305 gnd.n4116 gnd.n4115 10.6151
R10306 gnd.n4115 gnd.n2034 10.6151
R10307 gnd.n2602 gnd.n2601 10.6151
R10308 gnd.n2601 gnd.n2598 10.6151
R10309 gnd.n2596 gnd.n2593 10.6151
R10310 gnd.n2593 gnd.n2592 10.6151
R10311 gnd.n2592 gnd.n2589 10.6151
R10312 gnd.n2589 gnd.n2588 10.6151
R10313 gnd.n2588 gnd.n2585 10.6151
R10314 gnd.n2585 gnd.n2584 10.6151
R10315 gnd.n2584 gnd.n2581 10.6151
R10316 gnd.n2581 gnd.n2580 10.6151
R10317 gnd.n2580 gnd.n2577 10.6151
R10318 gnd.n2577 gnd.n2576 10.6151
R10319 gnd.n2576 gnd.n2573 10.6151
R10320 gnd.n2573 gnd.n2572 10.6151
R10321 gnd.n2572 gnd.n2569 10.6151
R10322 gnd.n2569 gnd.n2568 10.6151
R10323 gnd.n2568 gnd.n2565 10.6151
R10324 gnd.n2565 gnd.n2564 10.6151
R10325 gnd.n2564 gnd.n2561 10.6151
R10326 gnd.n2561 gnd.n2560 10.6151
R10327 gnd.n2560 gnd.n2557 10.6151
R10328 gnd.n2557 gnd.n2556 10.6151
R10329 gnd.n2556 gnd.n2553 10.6151
R10330 gnd.n2553 gnd.n2552 10.6151
R10331 gnd.n2552 gnd.n2549 10.6151
R10332 gnd.n2549 gnd.n2548 10.6151
R10333 gnd.n2548 gnd.n2545 10.6151
R10334 gnd.n2545 gnd.n2544 10.6151
R10335 gnd.n2544 gnd.n2541 10.6151
R10336 gnd.n2541 gnd.n2540 10.6151
R10337 gnd.n3640 gnd.n2425 10.6151
R10338 gnd.n3635 gnd.n2425 10.6151
R10339 gnd.n3635 gnd.n3634 10.6151
R10340 gnd.n3634 gnd.n3633 10.6151
R10341 gnd.n3633 gnd.n3630 10.6151
R10342 gnd.n3630 gnd.n3629 10.6151
R10343 gnd.n3629 gnd.n3626 10.6151
R10344 gnd.n3626 gnd.n3625 10.6151
R10345 gnd.n3625 gnd.n3622 10.6151
R10346 gnd.n3622 gnd.n3621 10.6151
R10347 gnd.n3621 gnd.n3618 10.6151
R10348 gnd.n3618 gnd.n3617 10.6151
R10349 gnd.n3617 gnd.n3614 10.6151
R10350 gnd.n3614 gnd.n3613 10.6151
R10351 gnd.n3613 gnd.n3610 10.6151
R10352 gnd.n3610 gnd.n3609 10.6151
R10353 gnd.n3609 gnd.n3606 10.6151
R10354 gnd.n3606 gnd.n3605 10.6151
R10355 gnd.n3605 gnd.n3602 10.6151
R10356 gnd.n3602 gnd.n3601 10.6151
R10357 gnd.n3601 gnd.n3598 10.6151
R10358 gnd.n3598 gnd.n3597 10.6151
R10359 gnd.n3597 gnd.n3594 10.6151
R10360 gnd.n3594 gnd.n3593 10.6151
R10361 gnd.n3593 gnd.n3590 10.6151
R10362 gnd.n3590 gnd.n3589 10.6151
R10363 gnd.n3589 gnd.n3586 10.6151
R10364 gnd.n3586 gnd.n3585 10.6151
R10365 gnd.n3582 gnd.n3581 10.6151
R10366 gnd.n3581 gnd.n3578 10.6151
R10367 gnd.n4294 gnd.n4293 10.6151
R10368 gnd.n4293 gnd.n4290 10.6151
R10369 gnd.n4290 gnd.n4289 10.6151
R10370 gnd.n4289 gnd.n4286 10.6151
R10371 gnd.n4286 gnd.n4285 10.6151
R10372 gnd.n4285 gnd.n4282 10.6151
R10373 gnd.n4282 gnd.n4281 10.6151
R10374 gnd.n4281 gnd.n4278 10.6151
R10375 gnd.n4278 gnd.n4277 10.6151
R10376 gnd.n4277 gnd.n4274 10.6151
R10377 gnd.n4274 gnd.n4273 10.6151
R10378 gnd.n4273 gnd.n4270 10.6151
R10379 gnd.n4270 gnd.n4269 10.6151
R10380 gnd.n4269 gnd.n4266 10.6151
R10381 gnd.n4266 gnd.n4265 10.6151
R10382 gnd.n4265 gnd.n4262 10.6151
R10383 gnd.n4262 gnd.n4261 10.6151
R10384 gnd.n4261 gnd.n4258 10.6151
R10385 gnd.n4258 gnd.n4257 10.6151
R10386 gnd.n4257 gnd.n4254 10.6151
R10387 gnd.n4254 gnd.n4253 10.6151
R10388 gnd.n4253 gnd.n4250 10.6151
R10389 gnd.n4250 gnd.n4249 10.6151
R10390 gnd.n4249 gnd.n4246 10.6151
R10391 gnd.n4246 gnd.n4245 10.6151
R10392 gnd.n4245 gnd.n4242 10.6151
R10393 gnd.n4242 gnd.n4241 10.6151
R10394 gnd.n4241 gnd.n4238 10.6151
R10395 gnd.n4236 gnd.n4233 10.6151
R10396 gnd.n4233 gnd.n4232 10.6151
R10397 gnd.n3643 gnd.n3642 10.6151
R10398 gnd.n3643 gnd.n2391 10.6151
R10399 gnd.n3657 gnd.n2391 10.6151
R10400 gnd.n3658 gnd.n3657 10.6151
R10401 gnd.n3660 gnd.n3658 10.6151
R10402 gnd.n3660 gnd.n3659 10.6151
R10403 gnd.n3659 gnd.n2368 10.6151
R10404 gnd.n3690 gnd.n2368 10.6151
R10405 gnd.n3691 gnd.n3690 10.6151
R10406 gnd.n3692 gnd.n3691 10.6151
R10407 gnd.n3692 gnd.n2355 10.6151
R10408 gnd.n3708 gnd.n2355 10.6151
R10409 gnd.n3709 gnd.n3708 10.6151
R10410 gnd.n3710 gnd.n3709 10.6151
R10411 gnd.n3710 gnd.n2342 10.6151
R10412 gnd.n3726 gnd.n2342 10.6151
R10413 gnd.n3727 gnd.n3726 10.6151
R10414 gnd.n3728 gnd.n3727 10.6151
R10415 gnd.n3728 gnd.n2330 10.6151
R10416 gnd.n3742 gnd.n2330 10.6151
R10417 gnd.n3743 gnd.n3742 10.6151
R10418 gnd.n3745 gnd.n3743 10.6151
R10419 gnd.n3745 gnd.n3744 10.6151
R10420 gnd.n3744 gnd.n2306 10.6151
R10421 gnd.n3772 gnd.n2306 10.6151
R10422 gnd.n3773 gnd.n3772 10.6151
R10423 gnd.n3774 gnd.n3773 10.6151
R10424 gnd.n3774 gnd.n2292 10.6151
R10425 gnd.n3791 gnd.n2292 10.6151
R10426 gnd.n3792 gnd.n3791 10.6151
R10427 gnd.n3793 gnd.n3792 10.6151
R10428 gnd.n3793 gnd.n2279 10.6151
R10429 gnd.n3822 gnd.n2279 10.6151
R10430 gnd.n3823 gnd.n3822 10.6151
R10431 gnd.n3824 gnd.n3823 10.6151
R10432 gnd.n3824 gnd.n2265 10.6151
R10433 gnd.n3840 gnd.n2265 10.6151
R10434 gnd.n3841 gnd.n3840 10.6151
R10435 gnd.n3843 gnd.n3841 10.6151
R10436 gnd.n3843 gnd.n3842 10.6151
R10437 gnd.n3842 gnd.n2230 10.6151
R10438 gnd.n3874 gnd.n2230 10.6151
R10439 gnd.n3875 gnd.n3874 10.6151
R10440 gnd.n3876 gnd.n3875 10.6151
R10441 gnd.n3876 gnd.n2216 10.6151
R10442 gnd.n3892 gnd.n2216 10.6151
R10443 gnd.n3893 gnd.n3892 10.6151
R10444 gnd.n3894 gnd.n3893 10.6151
R10445 gnd.n3894 gnd.n2202 10.6151
R10446 gnd.n3908 gnd.n2202 10.6151
R10447 gnd.n3909 gnd.n3908 10.6151
R10448 gnd.n3911 gnd.n3909 10.6151
R10449 gnd.n3911 gnd.n3910 10.6151
R10450 gnd.n3910 gnd.n2176 10.6151
R10451 gnd.n3954 gnd.n2176 10.6151
R10452 gnd.n3955 gnd.n3954 10.6151
R10453 gnd.n3956 gnd.n3955 10.6151
R10454 gnd.n3956 gnd.n2167 10.6151
R10455 gnd.n3986 gnd.n2167 10.6151
R10456 gnd.n3987 gnd.n3986 10.6151
R10457 gnd.n3988 gnd.n3987 10.6151
R10458 gnd.n3988 gnd.n2152 10.6151
R10459 gnd.n4004 gnd.n2152 10.6151
R10460 gnd.n4005 gnd.n4004 10.6151
R10461 gnd.n4006 gnd.n4005 10.6151
R10462 gnd.n4006 gnd.n2138 10.6151
R10463 gnd.n4035 gnd.n2138 10.6151
R10464 gnd.n4036 gnd.n4035 10.6151
R10465 gnd.n4038 gnd.n4036 10.6151
R10466 gnd.n4038 gnd.n4037 10.6151
R10467 gnd.n4037 gnd.n2120 10.6151
R10468 gnd.n4069 gnd.n2120 10.6151
R10469 gnd.n4070 gnd.n4069 10.6151
R10470 gnd.n4071 gnd.n4070 10.6151
R10471 gnd.n4071 gnd.n2103 10.6151
R10472 gnd.n4091 gnd.n2103 10.6151
R10473 gnd.n4092 gnd.n4091 10.6151
R10474 gnd.n4094 gnd.n4092 10.6151
R10475 gnd.n4094 gnd.n4093 10.6151
R10476 gnd.n4093 gnd.n2086 10.6151
R10477 gnd.n4143 gnd.n2086 10.6151
R10478 gnd.n4144 gnd.n4143 10.6151
R10479 gnd.n4145 gnd.n4144 10.6151
R10480 gnd.n4145 gnd.n2072 10.6151
R10481 gnd.n4161 gnd.n2072 10.6151
R10482 gnd.n4162 gnd.n4161 10.6151
R10483 gnd.n4163 gnd.n4162 10.6151
R10484 gnd.n4163 gnd.n2058 10.6151
R10485 gnd.n4185 gnd.n2058 10.6151
R10486 gnd.n4186 gnd.n4185 10.6151
R10487 gnd.n4187 gnd.n4186 10.6151
R10488 gnd.n4187 gnd.n2040 10.6151
R10489 gnd.n4207 gnd.n2040 10.6151
R10490 gnd.n4208 gnd.n4207 10.6151
R10491 gnd.n4296 gnd.n4208 10.6151
R10492 gnd.n5495 gnd.t82 10.5161
R10493 gnd.n6100 gnd.t105 10.5161
R10494 gnd.n6510 gnd.t89 10.5161
R10495 gnd.n3758 gnd.t330 10.5161
R10496 gnd.n4017 gnd.t125 10.5161
R10497 gnd.n6366 gnd.n6350 10.4732
R10498 gnd.n6334 gnd.n6318 10.4732
R10499 gnd.n6302 gnd.n6286 10.4732
R10500 gnd.n6271 gnd.n6255 10.4732
R10501 gnd.n6239 gnd.n6223 10.4732
R10502 gnd.n6207 gnd.n6191 10.4732
R10503 gnd.n6175 gnd.n6159 10.4732
R10504 gnd.n6144 gnd.n6128 10.4732
R10505 gnd.n3687 gnd.n3686 10.1975
R10506 gnd.n3819 gnd.n2275 10.1975
R10507 gnd.n2469 gnd.n2268 10.1975
R10508 gnd.n3984 gnd.n2169 10.1975
R10509 gnd.n3990 gnd.n2165 10.1975
R10510 gnd.n4166 gnd.n2068 10.1975
R10511 gnd.t231 gnd.n1871 10.1975
R10512 gnd.n6075 gnd.t148 9.87883
R10513 gnd.n7783 gnd.n66 9.73455
R10514 gnd.n6370 gnd.n6369 9.69747
R10515 gnd.n6338 gnd.n6337 9.69747
R10516 gnd.n6306 gnd.n6305 9.69747
R10517 gnd.n6275 gnd.n6274 9.69747
R10518 gnd.n6243 gnd.n6242 9.69747
R10519 gnd.n6211 gnd.n6210 9.69747
R10520 gnd.n6179 gnd.n6178 9.69747
R10521 gnd.n6148 gnd.n6147 9.69747
R10522 gnd.n3646 gnd.n2400 9.56018
R10523 gnd.n3740 gnd.n2332 9.56018
R10524 gnd.n3770 gnd.n3769 9.56018
R10525 gnd.n2468 gnd.t173 9.56018
R10526 gnd.n3863 gnd.n3862 9.56018
R10527 gnd.n3906 gnd.n3905 9.56018
R10528 gnd.n3983 gnd.t172 9.56018
R10529 gnd.n2136 gnd.n2134 9.56018
R10530 gnd.n4059 gnd.n2105 9.56018
R10531 gnd.n4893 gnd.n1326 9.45751
R10532 gnd.n1692 gnd.n1684 9.45599
R10533 gnd.n6376 gnd.n6375 9.45567
R10534 gnd.n6344 gnd.n6343 9.45567
R10535 gnd.n6312 gnd.n6311 9.45567
R10536 gnd.n6281 gnd.n6280 9.45567
R10537 gnd.n6249 gnd.n6248 9.45567
R10538 gnd.n6217 gnd.n6216 9.45567
R10539 gnd.n6185 gnd.n6184 9.45567
R10540 gnd.n6154 gnd.n6153 9.45567
R10541 gnd.n5339 gnd.n5338 9.39724
R10542 gnd.n6375 gnd.n6374 9.3005
R10543 gnd.n6348 gnd.n6347 9.3005
R10544 gnd.n6369 gnd.n6368 9.3005
R10545 gnd.n6367 gnd.n6366 9.3005
R10546 gnd.n6352 gnd.n6351 9.3005
R10547 gnd.n6361 gnd.n6360 9.3005
R10548 gnd.n6359 gnd.n6358 9.3005
R10549 gnd.n6343 gnd.n6342 9.3005
R10550 gnd.n6316 gnd.n6315 9.3005
R10551 gnd.n6337 gnd.n6336 9.3005
R10552 gnd.n6335 gnd.n6334 9.3005
R10553 gnd.n6320 gnd.n6319 9.3005
R10554 gnd.n6329 gnd.n6328 9.3005
R10555 gnd.n6327 gnd.n6326 9.3005
R10556 gnd.n6311 gnd.n6310 9.3005
R10557 gnd.n6284 gnd.n6283 9.3005
R10558 gnd.n6305 gnd.n6304 9.3005
R10559 gnd.n6303 gnd.n6302 9.3005
R10560 gnd.n6288 gnd.n6287 9.3005
R10561 gnd.n6297 gnd.n6296 9.3005
R10562 gnd.n6295 gnd.n6294 9.3005
R10563 gnd.n6280 gnd.n6279 9.3005
R10564 gnd.n6253 gnd.n6252 9.3005
R10565 gnd.n6274 gnd.n6273 9.3005
R10566 gnd.n6272 gnd.n6271 9.3005
R10567 gnd.n6257 gnd.n6256 9.3005
R10568 gnd.n6266 gnd.n6265 9.3005
R10569 gnd.n6264 gnd.n6263 9.3005
R10570 gnd.n6248 gnd.n6247 9.3005
R10571 gnd.n6221 gnd.n6220 9.3005
R10572 gnd.n6242 gnd.n6241 9.3005
R10573 gnd.n6240 gnd.n6239 9.3005
R10574 gnd.n6225 gnd.n6224 9.3005
R10575 gnd.n6234 gnd.n6233 9.3005
R10576 gnd.n6232 gnd.n6231 9.3005
R10577 gnd.n6216 gnd.n6215 9.3005
R10578 gnd.n6189 gnd.n6188 9.3005
R10579 gnd.n6210 gnd.n6209 9.3005
R10580 gnd.n6208 gnd.n6207 9.3005
R10581 gnd.n6193 gnd.n6192 9.3005
R10582 gnd.n6202 gnd.n6201 9.3005
R10583 gnd.n6200 gnd.n6199 9.3005
R10584 gnd.n6184 gnd.n6183 9.3005
R10585 gnd.n6157 gnd.n6156 9.3005
R10586 gnd.n6178 gnd.n6177 9.3005
R10587 gnd.n6176 gnd.n6175 9.3005
R10588 gnd.n6161 gnd.n6160 9.3005
R10589 gnd.n6170 gnd.n6169 9.3005
R10590 gnd.n6168 gnd.n6167 9.3005
R10591 gnd.n6153 gnd.n6152 9.3005
R10592 gnd.n6126 gnd.n6125 9.3005
R10593 gnd.n6147 gnd.n6146 9.3005
R10594 gnd.n6145 gnd.n6144 9.3005
R10595 gnd.n6130 gnd.n6129 9.3005
R10596 gnd.n6139 gnd.n6138 9.3005
R10597 gnd.n6137 gnd.n6136 9.3005
R10598 gnd.n964 gnd.n963 9.3005
R10599 gnd.n6484 gnd.n5144 9.3005
R10600 gnd.n6483 gnd.n5145 9.3005
R10601 gnd.n6482 gnd.n5146 9.3005
R10602 gnd.n6479 gnd.n5147 9.3005
R10603 gnd.n6478 gnd.n5148 9.3005
R10604 gnd.n6475 gnd.n5149 9.3005
R10605 gnd.n6474 gnd.n5150 9.3005
R10606 gnd.n6471 gnd.n5151 9.3005
R10607 gnd.n6470 gnd.n5152 9.3005
R10608 gnd.n6467 gnd.n5153 9.3005
R10609 gnd.n6466 gnd.n5154 9.3005
R10610 gnd.n6463 gnd.n5155 9.3005
R10611 gnd.n6462 gnd.n5156 9.3005
R10612 gnd.n6459 gnd.n6458 9.3005
R10613 gnd.n6457 gnd.n5157 9.3005
R10614 gnd.n6490 gnd.n6489 9.3005
R10615 gnd.n5762 gnd.n5761 9.3005
R10616 gnd.n5763 gnd.n5465 9.3005
R10617 gnd.n5765 gnd.n5764 9.3005
R10618 gnd.n5446 gnd.n5445 9.3005
R10619 gnd.n5792 gnd.n5791 9.3005
R10620 gnd.n5793 gnd.n5444 9.3005
R10621 gnd.n5797 gnd.n5794 9.3005
R10622 gnd.n5796 gnd.n5795 9.3005
R10623 gnd.n5420 gnd.n5419 9.3005
R10624 gnd.n5826 gnd.n5825 9.3005
R10625 gnd.n5827 gnd.n5418 9.3005
R10626 gnd.n5834 gnd.n5828 9.3005
R10627 gnd.n5833 gnd.n5829 9.3005
R10628 gnd.n5832 gnd.n5830 9.3005
R10629 gnd.n5387 gnd.n5386 9.3005
R10630 gnd.n5887 gnd.n5886 9.3005
R10631 gnd.n5888 gnd.n5385 9.3005
R10632 gnd.n5892 gnd.n5889 9.3005
R10633 gnd.n5891 gnd.n5890 9.3005
R10634 gnd.n5360 gnd.n5359 9.3005
R10635 gnd.n5927 gnd.n5926 9.3005
R10636 gnd.n5928 gnd.n5358 9.3005
R10637 gnd.n5932 gnd.n5929 9.3005
R10638 gnd.n5931 gnd.n5930 9.3005
R10639 gnd.n5285 gnd.n5284 9.3005
R10640 gnd.n5972 gnd.n5971 9.3005
R10641 gnd.n5973 gnd.n5283 9.3005
R10642 gnd.n5977 gnd.n5974 9.3005
R10643 gnd.n5976 gnd.n5975 9.3005
R10644 gnd.n5257 gnd.n5256 9.3005
R10645 gnd.n6011 gnd.n6010 9.3005
R10646 gnd.n6012 gnd.n5255 9.3005
R10647 gnd.n6019 gnd.n6013 9.3005
R10648 gnd.n6018 gnd.n6014 9.3005
R10649 gnd.n6017 gnd.n6015 9.3005
R10650 gnd.n5226 gnd.n5225 9.3005
R10651 gnd.n6066 gnd.n6065 9.3005
R10652 gnd.n6067 gnd.n5224 9.3005
R10653 gnd.n6072 gnd.n6068 9.3005
R10654 gnd.n6071 gnd.n6070 9.3005
R10655 gnd.n6069 gnd.n912 9.3005
R10656 gnd.n6521 gnd.n913 9.3005
R10657 gnd.n6520 gnd.n914 9.3005
R10658 gnd.n6519 gnd.n915 9.3005
R10659 gnd.n935 gnd.n916 9.3005
R10660 gnd.n936 gnd.n934 9.3005
R10661 gnd.n6507 gnd.n937 9.3005
R10662 gnd.n6506 gnd.n938 9.3005
R10663 gnd.n6505 gnd.n939 9.3005
R10664 gnd.n960 gnd.n940 9.3005
R10665 gnd.n961 gnd.n959 9.3005
R10666 gnd.n6493 gnd.n962 9.3005
R10667 gnd.n6492 gnd.n6491 9.3005
R10668 gnd.n5467 gnd.n5466 9.3005
R10669 gnd.n5707 gnd.n5706 9.3005
R10670 gnd.n5710 gnd.n5702 9.3005
R10671 gnd.n5711 gnd.n5701 9.3005
R10672 gnd.n5714 gnd.n5700 9.3005
R10673 gnd.n5715 gnd.n5699 9.3005
R10674 gnd.n5718 gnd.n5698 9.3005
R10675 gnd.n5719 gnd.n5697 9.3005
R10676 gnd.n5722 gnd.n5696 9.3005
R10677 gnd.n5723 gnd.n5695 9.3005
R10678 gnd.n5726 gnd.n5694 9.3005
R10679 gnd.n5727 gnd.n5693 9.3005
R10680 gnd.n5730 gnd.n5692 9.3005
R10681 gnd.n5732 gnd.n5691 9.3005
R10682 gnd.n5733 gnd.n5690 9.3005
R10683 gnd.n5734 gnd.n5689 9.3005
R10684 gnd.n5735 gnd.n5688 9.3005
R10685 gnd.n5703 gnd.n5484 9.3005
R10686 gnd.n5752 gnd.n5475 9.3005
R10687 gnd.n5754 gnd.n5753 9.3005
R10688 gnd.n5462 gnd.n5457 9.3005
R10689 gnd.n5775 gnd.n5456 9.3005
R10690 gnd.n5778 gnd.n5777 9.3005
R10691 gnd.n5780 gnd.n5779 9.3005
R10692 gnd.n5783 gnd.n5439 9.3005
R10693 gnd.n5781 gnd.n5437 9.3005
R10694 gnd.n5803 gnd.n5435 9.3005
R10695 gnd.n5807 gnd.n5806 9.3005
R10696 gnd.n5805 gnd.n5410 9.3005
R10697 gnd.n5841 gnd.n5409 9.3005
R10698 gnd.n5844 gnd.n5843 9.3005
R10699 gnd.n5407 gnd.n5406 9.3005
R10700 gnd.n5850 gnd.n5404 9.3005
R10701 gnd.n5852 gnd.n5851 9.3005
R10702 gnd.n5378 gnd.n5377 9.3005
R10703 gnd.n5901 gnd.n5900 9.3005
R10704 gnd.n5902 gnd.n5371 9.3005
R10705 gnd.n5910 gnd.n5370 9.3005
R10706 gnd.n5913 gnd.n5912 9.3005
R10707 gnd.n5915 gnd.n5914 9.3005
R10708 gnd.n5918 gnd.n5353 9.3005
R10709 gnd.n5916 gnd.n5351 9.3005
R10710 gnd.n5938 gnd.n5349 9.3005
R10711 gnd.n5940 gnd.n5939 9.3005
R10712 gnd.n5275 gnd.n5274 9.3005
R10713 gnd.n5986 gnd.n5985 9.3005
R10714 gnd.n5987 gnd.n5268 9.3005
R10715 gnd.n5995 gnd.n5267 9.3005
R10716 gnd.n5998 gnd.n5997 9.3005
R10717 gnd.n6000 gnd.n5999 9.3005
R10718 gnd.n6002 gnd.n5250 9.3005
R10719 gnd.n5247 gnd.n5245 9.3005
R10720 gnd.n6027 gnd.n6026 9.3005
R10721 gnd.n5248 gnd.n5231 9.3005
R10722 gnd.n6055 gnd.n5230 9.3005
R10723 gnd.n6059 gnd.n6057 9.3005
R10724 gnd.n6058 gnd.n5215 9.3005
R10725 gnd.n6080 gnd.n5214 9.3005
R10726 gnd.n6084 gnd.n6083 9.3005
R10727 gnd.n5207 gnd.n5206 9.3005
R10728 gnd.n6097 gnd.n6093 9.3005
R10729 gnd.n6096 gnd.n6095 9.3005
R10730 gnd.n5199 gnd.n5198 9.3005
R10731 gnd.n6119 gnd.n5200 9.3005
R10732 gnd.n6121 gnd.n6120 9.3005
R10733 gnd.n6123 gnd.n5197 9.3005
R10734 gnd.n6382 gnd.n6381 9.3005
R10735 gnd.n6384 gnd.n6383 9.3005
R10736 gnd.n6392 gnd.n6385 9.3005
R10737 gnd.n6391 gnd.n6387 9.3005
R10738 gnd.n6390 gnd.n5160 9.3005
R10739 gnd.n5751 gnd.n5478 9.3005
R10740 gnd.n6453 gnd.n5161 9.3005
R10741 gnd.n6452 gnd.n5163 9.3005
R10742 gnd.n6449 gnd.n5164 9.3005
R10743 gnd.n6448 gnd.n5165 9.3005
R10744 gnd.n6445 gnd.n5166 9.3005
R10745 gnd.n6444 gnd.n5167 9.3005
R10746 gnd.n6441 gnd.n5168 9.3005
R10747 gnd.n6440 gnd.n5169 9.3005
R10748 gnd.n6437 gnd.n5170 9.3005
R10749 gnd.n6436 gnd.n5171 9.3005
R10750 gnd.n6433 gnd.n5172 9.3005
R10751 gnd.n6432 gnd.n5173 9.3005
R10752 gnd.n6429 gnd.n5174 9.3005
R10753 gnd.n6428 gnd.n5175 9.3005
R10754 gnd.n6425 gnd.n5176 9.3005
R10755 gnd.n6424 gnd.n5177 9.3005
R10756 gnd.n6421 gnd.n5178 9.3005
R10757 gnd.n6420 gnd.n5179 9.3005
R10758 gnd.n6417 gnd.n5180 9.3005
R10759 gnd.n6416 gnd.n5181 9.3005
R10760 gnd.n6413 gnd.n5182 9.3005
R10761 gnd.n6412 gnd.n5183 9.3005
R10762 gnd.n6409 gnd.n5187 9.3005
R10763 gnd.n6408 gnd.n5188 9.3005
R10764 gnd.n6405 gnd.n5189 9.3005
R10765 gnd.n6404 gnd.n5190 9.3005
R10766 gnd.n6455 gnd.n6454 9.3005
R10767 gnd.n5948 gnd.n5947 9.3005
R10768 gnd.n5949 gnd.n5291 9.3005
R10769 gnd.n5966 gnd.n5950 9.3005
R10770 gnd.n5965 gnd.n5951 9.3005
R10771 gnd.n5964 gnd.n5952 9.3005
R10772 gnd.n5962 gnd.n5953 9.3005
R10773 gnd.n5961 gnd.n5954 9.3005
R10774 gnd.n5959 gnd.n5955 9.3005
R10775 gnd.n5958 gnd.n5956 9.3005
R10776 gnd.n5238 gnd.n5237 9.3005
R10777 gnd.n6034 gnd.n6033 9.3005
R10778 gnd.n6035 gnd.n5236 9.3005
R10779 gnd.n6049 gnd.n6036 9.3005
R10780 gnd.n6048 gnd.n6037 9.3005
R10781 gnd.n6047 gnd.n6038 9.3005
R10782 gnd.n6046 gnd.n6039 9.3005
R10783 gnd.n6044 gnd.n6040 9.3005
R10784 gnd.n6043 gnd.n6041 9.3005
R10785 gnd.n5204 gnd.n5203 9.3005
R10786 gnd.n6103 gnd.n6102 9.3005
R10787 gnd.n6104 gnd.n5202 9.3005
R10788 gnd.n6114 gnd.n6105 9.3005
R10789 gnd.n6113 gnd.n6106 9.3005
R10790 gnd.n6112 gnd.n6107 9.3005
R10791 gnd.n6109 gnd.n6108 9.3005
R10792 gnd.n5193 gnd.n5192 9.3005
R10793 gnd.n6398 gnd.n6397 9.3005
R10794 gnd.n6399 gnd.n5191 9.3005
R10795 gnd.n6401 gnd.n6400 9.3005
R10796 gnd.n5621 gnd.n5515 9.3005
R10797 gnd.n5623 gnd.n5622 9.3005
R10798 gnd.n5505 gnd.n5504 9.3005
R10799 gnd.n5636 gnd.n5635 9.3005
R10800 gnd.n5637 gnd.n5503 9.3005
R10801 gnd.n5639 gnd.n5638 9.3005
R10802 gnd.n5492 gnd.n5491 9.3005
R10803 gnd.n5652 gnd.n5651 9.3005
R10804 gnd.n5653 gnd.n5490 9.3005
R10805 gnd.n5677 gnd.n5654 9.3005
R10806 gnd.n5676 gnd.n5655 9.3005
R10807 gnd.n5675 gnd.n5656 9.3005
R10808 gnd.n5674 gnd.n5657 9.3005
R10809 gnd.n5672 gnd.n5658 9.3005
R10810 gnd.n5671 gnd.n5659 9.3005
R10811 gnd.n5669 gnd.n5660 9.3005
R10812 gnd.n5668 gnd.n5661 9.3005
R10813 gnd.n5666 gnd.n5662 9.3005
R10814 gnd.n5665 gnd.n5663 9.3005
R10815 gnd.n5427 gnd.n5426 9.3005
R10816 gnd.n5815 gnd.n5814 9.3005
R10817 gnd.n5816 gnd.n5425 9.3005
R10818 gnd.n5820 gnd.n5817 9.3005
R10819 gnd.n5819 gnd.n5818 9.3005
R10820 gnd.n5394 gnd.n5393 9.3005
R10821 gnd.n5862 gnd.n5861 9.3005
R10822 gnd.n5863 gnd.n5392 9.3005
R10823 gnd.n5865 gnd.n5864 9.3005
R10824 gnd.n5620 gnd.n5619 9.3005
R10825 gnd.n5560 gnd.n5559 9.3005
R10826 gnd.n5565 gnd.n5557 9.3005
R10827 gnd.n5566 gnd.n5556 9.3005
R10828 gnd.n5568 gnd.n5553 9.3005
R10829 gnd.n5552 gnd.n5550 9.3005
R10830 gnd.n5574 gnd.n5549 9.3005
R10831 gnd.n5575 gnd.n5548 9.3005
R10832 gnd.n5576 gnd.n5547 9.3005
R10833 gnd.n5546 gnd.n5544 9.3005
R10834 gnd.n5582 gnd.n5543 9.3005
R10835 gnd.n5583 gnd.n5542 9.3005
R10836 gnd.n5584 gnd.n5541 9.3005
R10837 gnd.n5540 gnd.n5538 9.3005
R10838 gnd.n5590 gnd.n5537 9.3005
R10839 gnd.n5591 gnd.n5536 9.3005
R10840 gnd.n5592 gnd.n5535 9.3005
R10841 gnd.n5534 gnd.n5532 9.3005
R10842 gnd.n5598 gnd.n5531 9.3005
R10843 gnd.n5599 gnd.n5530 9.3005
R10844 gnd.n5600 gnd.n5529 9.3005
R10845 gnd.n5528 gnd.n5526 9.3005
R10846 gnd.n5605 gnd.n5525 9.3005
R10847 gnd.n5606 gnd.n5524 9.3005
R10848 gnd.n5523 gnd.n5521 9.3005
R10849 gnd.n5611 gnd.n5520 9.3005
R10850 gnd.n5613 gnd.n5612 9.3005
R10851 gnd.n5558 gnd.n5516 9.3005
R10852 gnd.n5511 gnd.n5510 9.3005
R10853 gnd.n5628 gnd.n5627 9.3005
R10854 gnd.n5629 gnd.n5509 9.3005
R10855 gnd.n5631 gnd.n5630 9.3005
R10856 gnd.n5499 gnd.n5498 9.3005
R10857 gnd.n5644 gnd.n5643 9.3005
R10858 gnd.n5645 gnd.n5497 9.3005
R10859 gnd.n5647 gnd.n5646 9.3005
R10860 gnd.n5486 gnd.n5485 9.3005
R10861 gnd.n5742 gnd.n5741 9.3005
R10862 gnd.n5744 gnd.n5483 9.3005
R10863 gnd.n5746 gnd.n5745 9.3005
R10864 gnd.n5477 gnd.n5474 9.3005
R10865 gnd.n5756 gnd.n5755 9.3005
R10866 gnd.n5476 gnd.n5458 9.3005
R10867 gnd.n5774 gnd.n5773 9.3005
R10868 gnd.n5776 gnd.n5454 9.3005
R10869 gnd.n5786 gnd.n5455 9.3005
R10870 gnd.n5785 gnd.n5784 9.3005
R10871 gnd.n5782 gnd.n5433 9.3005
R10872 gnd.n5810 gnd.n5434 9.3005
R10873 gnd.n5809 gnd.n5808 9.3005
R10874 gnd.n5436 gnd.n5411 9.3005
R10875 gnd.n5840 gnd.n5839 9.3005
R10876 gnd.n5842 gnd.n5401 9.3005
R10877 gnd.n5857 gnd.n5402 9.3005
R10878 gnd.n5856 gnd.n5403 9.3005
R10879 gnd.n5855 gnd.n5853 9.3005
R10880 gnd.n5405 gnd.n5379 9.3005
R10881 gnd.n5898 gnd.n5897 9.3005
R10882 gnd.n5899 gnd.n5372 9.3005
R10883 gnd.n5909 gnd.n5908 9.3005
R10884 gnd.n5911 gnd.n5368 9.3005
R10885 gnd.n5921 gnd.n5369 9.3005
R10886 gnd.n5920 gnd.n5919 9.3005
R10887 gnd.n5917 gnd.n5347 9.3005
R10888 gnd.n5943 gnd.n5348 9.3005
R10889 gnd.n5942 gnd.n5941 9.3005
R10890 gnd.n5350 gnd.n5276 9.3005
R10891 gnd.n5983 gnd.n5982 9.3005
R10892 gnd.n5984 gnd.n5269 9.3005
R10893 gnd.n5994 gnd.n5993 9.3005
R10894 gnd.n5996 gnd.n5265 9.3005
R10895 gnd.n6005 gnd.n5266 9.3005
R10896 gnd.n6004 gnd.n6003 9.3005
R10897 gnd.n6001 gnd.n5244 9.3005
R10898 gnd.n6029 gnd.n6028 9.3005
R10899 gnd.n5246 gnd.n5232 9.3005
R10900 gnd.n6054 gnd.n6053 9.3005
R10901 gnd.n6056 gnd.n5216 9.3005
R10902 gnd.n6077 gnd.n5217 9.3005
R10903 gnd.n6079 gnd.n6078 9.3005
R10904 gnd.n6081 gnd.n5210 9.3005
R10905 gnd.n6082 gnd.n5208 9.3005
R10906 gnd.n6092 gnd.n6091 9.3005
R10907 gnd.n6094 gnd.n923 9.3005
R10908 gnd.n6514 gnd.n924 9.3005
R10909 gnd.n6513 gnd.n925 9.3005
R10910 gnd.n6512 gnd.n926 9.3005
R10911 gnd.n6122 gnd.n927 9.3005
R10912 gnd.n6380 gnd.n948 9.3005
R10913 gnd.n6500 gnd.n949 9.3005
R10914 gnd.n6499 gnd.n950 9.3005
R10915 gnd.n6498 gnd.n951 9.3005
R10916 gnd.n6386 gnd.n952 9.3005
R10917 gnd.n5615 gnd.n5614 9.3005
R10918 gnd.n738 gnd.n737 9.3005
R10919 gnd.n6697 gnd.n6696 9.3005
R10920 gnd.n6698 gnd.n736 9.3005
R10921 gnd.n6700 gnd.n6699 9.3005
R10922 gnd.n732 gnd.n731 9.3005
R10923 gnd.n6707 gnd.n6706 9.3005
R10924 gnd.n6708 gnd.n730 9.3005
R10925 gnd.n6710 gnd.n6709 9.3005
R10926 gnd.n726 gnd.n725 9.3005
R10927 gnd.n6717 gnd.n6716 9.3005
R10928 gnd.n6718 gnd.n724 9.3005
R10929 gnd.n6720 gnd.n6719 9.3005
R10930 gnd.n720 gnd.n719 9.3005
R10931 gnd.n6727 gnd.n6726 9.3005
R10932 gnd.n6728 gnd.n718 9.3005
R10933 gnd.n6730 gnd.n6729 9.3005
R10934 gnd.n714 gnd.n713 9.3005
R10935 gnd.n6737 gnd.n6736 9.3005
R10936 gnd.n6738 gnd.n712 9.3005
R10937 gnd.n6740 gnd.n6739 9.3005
R10938 gnd.n708 gnd.n707 9.3005
R10939 gnd.n6747 gnd.n6746 9.3005
R10940 gnd.n6748 gnd.n706 9.3005
R10941 gnd.n6750 gnd.n6749 9.3005
R10942 gnd.n702 gnd.n701 9.3005
R10943 gnd.n6757 gnd.n6756 9.3005
R10944 gnd.n6758 gnd.n700 9.3005
R10945 gnd.n6760 gnd.n6759 9.3005
R10946 gnd.n696 gnd.n695 9.3005
R10947 gnd.n6767 gnd.n6766 9.3005
R10948 gnd.n6768 gnd.n694 9.3005
R10949 gnd.n6770 gnd.n6769 9.3005
R10950 gnd.n690 gnd.n689 9.3005
R10951 gnd.n6777 gnd.n6776 9.3005
R10952 gnd.n6778 gnd.n688 9.3005
R10953 gnd.n6780 gnd.n6779 9.3005
R10954 gnd.n684 gnd.n683 9.3005
R10955 gnd.n6787 gnd.n6786 9.3005
R10956 gnd.n6788 gnd.n682 9.3005
R10957 gnd.n6790 gnd.n6789 9.3005
R10958 gnd.n678 gnd.n677 9.3005
R10959 gnd.n6797 gnd.n6796 9.3005
R10960 gnd.n6798 gnd.n676 9.3005
R10961 gnd.n6800 gnd.n6799 9.3005
R10962 gnd.n672 gnd.n671 9.3005
R10963 gnd.n6807 gnd.n6806 9.3005
R10964 gnd.n6808 gnd.n670 9.3005
R10965 gnd.n6810 gnd.n6809 9.3005
R10966 gnd.n666 gnd.n665 9.3005
R10967 gnd.n6817 gnd.n6816 9.3005
R10968 gnd.n6818 gnd.n664 9.3005
R10969 gnd.n6820 gnd.n6819 9.3005
R10970 gnd.n660 gnd.n659 9.3005
R10971 gnd.n6827 gnd.n6826 9.3005
R10972 gnd.n6828 gnd.n658 9.3005
R10973 gnd.n6830 gnd.n6829 9.3005
R10974 gnd.n654 gnd.n653 9.3005
R10975 gnd.n6837 gnd.n6836 9.3005
R10976 gnd.n6838 gnd.n652 9.3005
R10977 gnd.n6840 gnd.n6839 9.3005
R10978 gnd.n648 gnd.n647 9.3005
R10979 gnd.n6847 gnd.n6846 9.3005
R10980 gnd.n6848 gnd.n646 9.3005
R10981 gnd.n6850 gnd.n6849 9.3005
R10982 gnd.n642 gnd.n641 9.3005
R10983 gnd.n6857 gnd.n6856 9.3005
R10984 gnd.n6858 gnd.n640 9.3005
R10985 gnd.n6860 gnd.n6859 9.3005
R10986 gnd.n636 gnd.n635 9.3005
R10987 gnd.n6867 gnd.n6866 9.3005
R10988 gnd.n6868 gnd.n634 9.3005
R10989 gnd.n6870 gnd.n6869 9.3005
R10990 gnd.n630 gnd.n629 9.3005
R10991 gnd.n6877 gnd.n6876 9.3005
R10992 gnd.n6878 gnd.n628 9.3005
R10993 gnd.n6880 gnd.n6879 9.3005
R10994 gnd.n624 gnd.n623 9.3005
R10995 gnd.n6887 gnd.n6886 9.3005
R10996 gnd.n6888 gnd.n622 9.3005
R10997 gnd.n6890 gnd.n6889 9.3005
R10998 gnd.n618 gnd.n617 9.3005
R10999 gnd.n6897 gnd.n6896 9.3005
R11000 gnd.n6898 gnd.n616 9.3005
R11001 gnd.n6900 gnd.n6899 9.3005
R11002 gnd.n612 gnd.n611 9.3005
R11003 gnd.n6907 gnd.n6906 9.3005
R11004 gnd.n6908 gnd.n610 9.3005
R11005 gnd.n6910 gnd.n6909 9.3005
R11006 gnd.n606 gnd.n605 9.3005
R11007 gnd.n6917 gnd.n6916 9.3005
R11008 gnd.n6918 gnd.n604 9.3005
R11009 gnd.n6920 gnd.n6919 9.3005
R11010 gnd.n600 gnd.n599 9.3005
R11011 gnd.n6927 gnd.n6926 9.3005
R11012 gnd.n6928 gnd.n598 9.3005
R11013 gnd.n6930 gnd.n6929 9.3005
R11014 gnd.n594 gnd.n593 9.3005
R11015 gnd.n6937 gnd.n6936 9.3005
R11016 gnd.n6938 gnd.n592 9.3005
R11017 gnd.n6940 gnd.n6939 9.3005
R11018 gnd.n588 gnd.n587 9.3005
R11019 gnd.n6947 gnd.n6946 9.3005
R11020 gnd.n6948 gnd.n586 9.3005
R11021 gnd.n6950 gnd.n6949 9.3005
R11022 gnd.n582 gnd.n581 9.3005
R11023 gnd.n6957 gnd.n6956 9.3005
R11024 gnd.n6958 gnd.n580 9.3005
R11025 gnd.n6960 gnd.n6959 9.3005
R11026 gnd.n576 gnd.n575 9.3005
R11027 gnd.n6967 gnd.n6966 9.3005
R11028 gnd.n6968 gnd.n574 9.3005
R11029 gnd.n6970 gnd.n6969 9.3005
R11030 gnd.n570 gnd.n569 9.3005
R11031 gnd.n6977 gnd.n6976 9.3005
R11032 gnd.n6978 gnd.n568 9.3005
R11033 gnd.n6980 gnd.n6979 9.3005
R11034 gnd.n564 gnd.n563 9.3005
R11035 gnd.n6987 gnd.n6986 9.3005
R11036 gnd.n6988 gnd.n562 9.3005
R11037 gnd.n6990 gnd.n6989 9.3005
R11038 gnd.n558 gnd.n557 9.3005
R11039 gnd.n6997 gnd.n6996 9.3005
R11040 gnd.n6998 gnd.n556 9.3005
R11041 gnd.n7000 gnd.n6999 9.3005
R11042 gnd.n552 gnd.n551 9.3005
R11043 gnd.n7007 gnd.n7006 9.3005
R11044 gnd.n7008 gnd.n550 9.3005
R11045 gnd.n7010 gnd.n7009 9.3005
R11046 gnd.n546 gnd.n545 9.3005
R11047 gnd.n7017 gnd.n7016 9.3005
R11048 gnd.n7018 gnd.n544 9.3005
R11049 gnd.n7020 gnd.n7019 9.3005
R11050 gnd.n540 gnd.n539 9.3005
R11051 gnd.n7027 gnd.n7026 9.3005
R11052 gnd.n7028 gnd.n538 9.3005
R11053 gnd.n7030 gnd.n7029 9.3005
R11054 gnd.n534 gnd.n533 9.3005
R11055 gnd.n7037 gnd.n7036 9.3005
R11056 gnd.n7038 gnd.n532 9.3005
R11057 gnd.n7040 gnd.n7039 9.3005
R11058 gnd.n528 gnd.n527 9.3005
R11059 gnd.n7047 gnd.n7046 9.3005
R11060 gnd.n7048 gnd.n526 9.3005
R11061 gnd.n7050 gnd.n7049 9.3005
R11062 gnd.n522 gnd.n521 9.3005
R11063 gnd.n7057 gnd.n7056 9.3005
R11064 gnd.n7058 gnd.n520 9.3005
R11065 gnd.n7060 gnd.n7059 9.3005
R11066 gnd.n516 gnd.n515 9.3005
R11067 gnd.n7067 gnd.n7066 9.3005
R11068 gnd.n7068 gnd.n514 9.3005
R11069 gnd.n7070 gnd.n7069 9.3005
R11070 gnd.n510 gnd.n509 9.3005
R11071 gnd.n7077 gnd.n7076 9.3005
R11072 gnd.n7078 gnd.n508 9.3005
R11073 gnd.n7080 gnd.n7079 9.3005
R11074 gnd.n504 gnd.n503 9.3005
R11075 gnd.n7087 gnd.n7086 9.3005
R11076 gnd.n7088 gnd.n502 9.3005
R11077 gnd.n7090 gnd.n7089 9.3005
R11078 gnd.n498 gnd.n497 9.3005
R11079 gnd.n7097 gnd.n7096 9.3005
R11080 gnd.n7098 gnd.n496 9.3005
R11081 gnd.n7100 gnd.n7099 9.3005
R11082 gnd.n492 gnd.n491 9.3005
R11083 gnd.n7107 gnd.n7106 9.3005
R11084 gnd.n7108 gnd.n490 9.3005
R11085 gnd.n7110 gnd.n7109 9.3005
R11086 gnd.n486 gnd.n485 9.3005
R11087 gnd.n7117 gnd.n7116 9.3005
R11088 gnd.n7118 gnd.n484 9.3005
R11089 gnd.n7120 gnd.n7119 9.3005
R11090 gnd.n480 gnd.n479 9.3005
R11091 gnd.n7127 gnd.n7126 9.3005
R11092 gnd.n7128 gnd.n478 9.3005
R11093 gnd.n7130 gnd.n7129 9.3005
R11094 gnd.n474 gnd.n473 9.3005
R11095 gnd.n7137 gnd.n7136 9.3005
R11096 gnd.n7138 gnd.n472 9.3005
R11097 gnd.n7140 gnd.n7139 9.3005
R11098 gnd.n468 gnd.n467 9.3005
R11099 gnd.n7147 gnd.n7146 9.3005
R11100 gnd.n7148 gnd.n466 9.3005
R11101 gnd.n7150 gnd.n7149 9.3005
R11102 gnd.n462 gnd.n461 9.3005
R11103 gnd.n7157 gnd.n7156 9.3005
R11104 gnd.n7158 gnd.n460 9.3005
R11105 gnd.n7160 gnd.n7159 9.3005
R11106 gnd.n456 gnd.n455 9.3005
R11107 gnd.n7167 gnd.n7166 9.3005
R11108 gnd.n7168 gnd.n454 9.3005
R11109 gnd.n7171 gnd.n7170 9.3005
R11110 gnd.n7169 gnd.n450 9.3005
R11111 gnd.n7177 gnd.n449 9.3005
R11112 gnd.n7179 gnd.n7178 9.3005
R11113 gnd.n445 gnd.n444 9.3005
R11114 gnd.n7188 gnd.n7187 9.3005
R11115 gnd.n7189 gnd.n443 9.3005
R11116 gnd.n7191 gnd.n7190 9.3005
R11117 gnd.n439 gnd.n438 9.3005
R11118 gnd.n7198 gnd.n7197 9.3005
R11119 gnd.n7199 gnd.n437 9.3005
R11120 gnd.n7201 gnd.n7200 9.3005
R11121 gnd.n433 gnd.n432 9.3005
R11122 gnd.n7208 gnd.n7207 9.3005
R11123 gnd.n7209 gnd.n431 9.3005
R11124 gnd.n7211 gnd.n7210 9.3005
R11125 gnd.n427 gnd.n426 9.3005
R11126 gnd.n7218 gnd.n7217 9.3005
R11127 gnd.n7219 gnd.n425 9.3005
R11128 gnd.n7221 gnd.n7220 9.3005
R11129 gnd.n421 gnd.n420 9.3005
R11130 gnd.n7228 gnd.n7227 9.3005
R11131 gnd.n7229 gnd.n419 9.3005
R11132 gnd.n7231 gnd.n7230 9.3005
R11133 gnd.n415 gnd.n414 9.3005
R11134 gnd.n7238 gnd.n7237 9.3005
R11135 gnd.n7239 gnd.n413 9.3005
R11136 gnd.n7241 gnd.n7240 9.3005
R11137 gnd.n409 gnd.n408 9.3005
R11138 gnd.n7248 gnd.n7247 9.3005
R11139 gnd.n7249 gnd.n407 9.3005
R11140 gnd.n7251 gnd.n7250 9.3005
R11141 gnd.n403 gnd.n402 9.3005
R11142 gnd.n7258 gnd.n7257 9.3005
R11143 gnd.n7259 gnd.n401 9.3005
R11144 gnd.n7261 gnd.n7260 9.3005
R11145 gnd.n397 gnd.n396 9.3005
R11146 gnd.n7268 gnd.n7267 9.3005
R11147 gnd.n7269 gnd.n395 9.3005
R11148 gnd.n7271 gnd.n7270 9.3005
R11149 gnd.n391 gnd.n390 9.3005
R11150 gnd.n7278 gnd.n7277 9.3005
R11151 gnd.n7279 gnd.n389 9.3005
R11152 gnd.n7281 gnd.n7280 9.3005
R11153 gnd.n385 gnd.n384 9.3005
R11154 gnd.n7288 gnd.n7287 9.3005
R11155 gnd.n7289 gnd.n383 9.3005
R11156 gnd.n7291 gnd.n7290 9.3005
R11157 gnd.n379 gnd.n378 9.3005
R11158 gnd.n7298 gnd.n7297 9.3005
R11159 gnd.n7299 gnd.n377 9.3005
R11160 gnd.n7301 gnd.n7300 9.3005
R11161 gnd.n373 gnd.n372 9.3005
R11162 gnd.n7308 gnd.n7307 9.3005
R11163 gnd.n7309 gnd.n371 9.3005
R11164 gnd.n7311 gnd.n7310 9.3005
R11165 gnd.n367 gnd.n366 9.3005
R11166 gnd.n7318 gnd.n7317 9.3005
R11167 gnd.n7319 gnd.n365 9.3005
R11168 gnd.n7321 gnd.n7320 9.3005
R11169 gnd.n361 gnd.n360 9.3005
R11170 gnd.n7328 gnd.n7327 9.3005
R11171 gnd.n7329 gnd.n359 9.3005
R11172 gnd.n7331 gnd.n7330 9.3005
R11173 gnd.n355 gnd.n354 9.3005
R11174 gnd.n7338 gnd.n7337 9.3005
R11175 gnd.n7339 gnd.n353 9.3005
R11176 gnd.n7341 gnd.n7340 9.3005
R11177 gnd.n349 gnd.n348 9.3005
R11178 gnd.n7348 gnd.n7347 9.3005
R11179 gnd.n7349 gnd.n347 9.3005
R11180 gnd.n7351 gnd.n7350 9.3005
R11181 gnd.n343 gnd.n342 9.3005
R11182 gnd.n7358 gnd.n7357 9.3005
R11183 gnd.n7359 gnd.n341 9.3005
R11184 gnd.n7361 gnd.n7360 9.3005
R11185 gnd.n337 gnd.n336 9.3005
R11186 gnd.n7368 gnd.n7367 9.3005
R11187 gnd.n7369 gnd.n335 9.3005
R11188 gnd.n7371 gnd.n7370 9.3005
R11189 gnd.n331 gnd.n330 9.3005
R11190 gnd.n7378 gnd.n7377 9.3005
R11191 gnd.n7379 gnd.n329 9.3005
R11192 gnd.n7381 gnd.n7380 9.3005
R11193 gnd.n325 gnd.n324 9.3005
R11194 gnd.n7389 gnd.n7388 9.3005
R11195 gnd.n7390 gnd.n323 9.3005
R11196 gnd.n7392 gnd.n7391 9.3005
R11197 gnd.n7181 gnd.n7180 9.3005
R11198 gnd.n7734 gnd.n112 9.3005
R11199 gnd.n7733 gnd.n114 9.3005
R11200 gnd.n119 gnd.n115 9.3005
R11201 gnd.n7728 gnd.n120 9.3005
R11202 gnd.n7727 gnd.n121 9.3005
R11203 gnd.n7726 gnd.n122 9.3005
R11204 gnd.n126 gnd.n123 9.3005
R11205 gnd.n7721 gnd.n127 9.3005
R11206 gnd.n7720 gnd.n128 9.3005
R11207 gnd.n7719 gnd.n129 9.3005
R11208 gnd.n133 gnd.n130 9.3005
R11209 gnd.n7714 gnd.n134 9.3005
R11210 gnd.n7713 gnd.n135 9.3005
R11211 gnd.n7712 gnd.n136 9.3005
R11212 gnd.n140 gnd.n137 9.3005
R11213 gnd.n7707 gnd.n141 9.3005
R11214 gnd.n7706 gnd.n142 9.3005
R11215 gnd.n7702 gnd.n143 9.3005
R11216 gnd.n147 gnd.n144 9.3005
R11217 gnd.n7697 gnd.n148 9.3005
R11218 gnd.n7696 gnd.n149 9.3005
R11219 gnd.n7695 gnd.n150 9.3005
R11220 gnd.n154 gnd.n151 9.3005
R11221 gnd.n7690 gnd.n155 9.3005
R11222 gnd.n7689 gnd.n156 9.3005
R11223 gnd.n7688 gnd.n157 9.3005
R11224 gnd.n161 gnd.n158 9.3005
R11225 gnd.n7683 gnd.n162 9.3005
R11226 gnd.n7682 gnd.n163 9.3005
R11227 gnd.n7681 gnd.n164 9.3005
R11228 gnd.n168 gnd.n165 9.3005
R11229 gnd.n7676 gnd.n169 9.3005
R11230 gnd.n7675 gnd.n170 9.3005
R11231 gnd.n7674 gnd.n171 9.3005
R11232 gnd.n175 gnd.n172 9.3005
R11233 gnd.n7669 gnd.n176 9.3005
R11234 gnd.n7668 gnd.n7667 9.3005
R11235 gnd.n7666 gnd.n179 9.3005
R11236 gnd.n7736 gnd.n7735 9.3005
R11237 gnd.n1981 gnd.n1640 9.3005
R11238 gnd.n4486 gnd.n1639 9.3005
R11239 gnd.n4488 gnd.n4487 9.3005
R11240 gnd.n4489 gnd.n1638 9.3005
R11241 gnd.n4515 gnd.n4490 9.3005
R11242 gnd.n4514 gnd.n4491 9.3005
R11243 gnd.n4513 gnd.n4492 9.3005
R11244 gnd.n4512 gnd.n4493 9.3005
R11245 gnd.n4511 gnd.n4494 9.3005
R11246 gnd.n4509 gnd.n4495 9.3005
R11247 gnd.n4508 gnd.n4496 9.3005
R11248 gnd.n4506 gnd.n4497 9.3005
R11249 gnd.n4505 gnd.n4498 9.3005
R11250 gnd.n4504 gnd.n4499 9.3005
R11251 gnd.n4502 gnd.n4501 9.3005
R11252 gnd.n4500 gnd.n1558 9.3005
R11253 gnd.n4611 gnd.n1559 9.3005
R11254 gnd.n4612 gnd.n1557 9.3005
R11255 gnd.n4615 gnd.n4614 9.3005
R11256 gnd.n4616 gnd.n1556 9.3005
R11257 gnd.n4620 gnd.n4617 9.3005
R11258 gnd.n4619 gnd.n4618 9.3005
R11259 gnd.n1550 gnd.n1549 9.3005
R11260 gnd.n4638 gnd.n4637 9.3005
R11261 gnd.n4639 gnd.n1548 9.3005
R11262 gnd.n4641 gnd.n4640 9.3005
R11263 gnd.n300 gnd.n299 9.3005
R11264 gnd.n7475 gnd.n301 9.3005
R11265 gnd.n7474 gnd.n302 9.3005
R11266 gnd.n7473 gnd.n303 9.3005
R11267 gnd.n7402 gnd.n304 9.3005
R11268 gnd.n7406 gnd.n7405 9.3005
R11269 gnd.n7407 gnd.n7401 9.3005
R11270 gnd.n7412 gnd.n7408 9.3005
R11271 gnd.n7413 gnd.n7400 9.3005
R11272 gnd.n7417 gnd.n7416 9.3005
R11273 gnd.n7418 gnd.n7399 9.3005
R11274 gnd.n7451 gnd.n7419 9.3005
R11275 gnd.n7450 gnd.n7420 9.3005
R11276 gnd.n7449 gnd.n7421 9.3005
R11277 gnd.n7446 gnd.n7422 9.3005
R11278 gnd.n7445 gnd.n7423 9.3005
R11279 gnd.n7443 gnd.n7424 9.3005
R11280 gnd.n7442 gnd.n7425 9.3005
R11281 gnd.n7440 gnd.n7426 9.3005
R11282 gnd.n7439 gnd.n7427 9.3005
R11283 gnd.n7437 gnd.n7428 9.3005
R11284 gnd.n7436 gnd.n7429 9.3005
R11285 gnd.n7434 gnd.n7430 9.3005
R11286 gnd.n7433 gnd.n7432 9.3005
R11287 gnd.n7431 gnd.n183 9.3005
R11288 gnd.n7663 gnd.n182 9.3005
R11289 gnd.n7665 gnd.n7664 9.3005
R11290 gnd.n1983 gnd.n1982 9.3005
R11291 gnd.n1991 gnd.n1990 9.3005
R11292 gnd.n1980 gnd.n1975 9.3005
R11293 gnd.n1997 gnd.n1974 9.3005
R11294 gnd.n1998 gnd.n1973 9.3005
R11295 gnd.n1999 gnd.n1972 9.3005
R11296 gnd.n1971 gnd.n1969 9.3005
R11297 gnd.n2005 gnd.n1968 9.3005
R11298 gnd.n2006 gnd.n1967 9.3005
R11299 gnd.n2007 gnd.n1966 9.3005
R11300 gnd.n1965 gnd.n1963 9.3005
R11301 gnd.n2013 gnd.n1962 9.3005
R11302 gnd.n2014 gnd.n1961 9.3005
R11303 gnd.n2015 gnd.n1960 9.3005
R11304 gnd.n1959 gnd.n1957 9.3005
R11305 gnd.n2021 gnd.n1956 9.3005
R11306 gnd.n2022 gnd.n1955 9.3005
R11307 gnd.n2023 gnd.n1954 9.3005
R11308 gnd.n1953 gnd.n1951 9.3005
R11309 gnd.n2029 gnd.n1950 9.3005
R11310 gnd.n1946 gnd.n1889 9.3005
R11311 gnd.n1945 gnd.n1944 9.3005
R11312 gnd.n1892 gnd.n1891 9.3005
R11313 gnd.n1935 gnd.n1895 9.3005
R11314 gnd.n1937 gnd.n1936 9.3005
R11315 gnd.n1934 gnd.n1897 9.3005
R11316 gnd.n1933 gnd.n1932 9.3005
R11317 gnd.n1899 gnd.n1898 9.3005
R11318 gnd.n1926 gnd.n1925 9.3005
R11319 gnd.n1924 gnd.n1901 9.3005
R11320 gnd.n1923 gnd.n1922 9.3005
R11321 gnd.n1903 gnd.n1902 9.3005
R11322 gnd.n1916 gnd.n1915 9.3005
R11323 gnd.n1914 gnd.n1905 9.3005
R11324 gnd.n1913 gnd.n1912 9.3005
R11325 gnd.n1908 gnd.n1907 9.3005
R11326 gnd.n1989 gnd.n1979 9.3005
R11327 gnd.n1988 gnd.n1987 9.3005
R11328 gnd.n4719 gnd.n1485 9.3005
R11329 gnd.n4718 gnd.n1486 9.3005
R11330 gnd.n4717 gnd.n1487 9.3005
R11331 gnd.n4519 gnd.n1488 9.3005
R11332 gnd.n4523 gnd.n4520 9.3005
R11333 gnd.n4522 gnd.n4521 9.3005
R11334 gnd.n1603 gnd.n1602 9.3005
R11335 gnd.n4550 gnd.n4549 9.3005
R11336 gnd.n4551 gnd.n1601 9.3005
R11337 gnd.n4555 gnd.n4552 9.3005
R11338 gnd.n4554 gnd.n4553 9.3005
R11339 gnd.n1576 gnd.n1575 9.3005
R11340 gnd.n4589 gnd.n4588 9.3005
R11341 gnd.n4590 gnd.n1574 9.3005
R11342 gnd.n4594 gnd.n4591 9.3005
R11343 gnd.n4593 gnd.n4592 9.3005
R11344 gnd.n1524 gnd.n1523 9.3005
R11345 gnd.n4679 gnd.n4678 9.3005
R11346 gnd.n4680 gnd.n1522 9.3005
R11347 gnd.n4682 gnd.n4681 9.3005
R11348 gnd.n274 gnd.n267 9.3005
R11349 gnd.n253 gnd.n252 9.3005
R11350 gnd.n7516 gnd.n7515 9.3005
R11351 gnd.n7517 gnd.n251 9.3005
R11352 gnd.n7519 gnd.n7518 9.3005
R11353 gnd.n237 gnd.n236 9.3005
R11354 gnd.n7532 gnd.n7531 9.3005
R11355 gnd.n7533 gnd.n235 9.3005
R11356 gnd.n7535 gnd.n7534 9.3005
R11357 gnd.n223 gnd.n222 9.3005
R11358 gnd.n7548 gnd.n7547 9.3005
R11359 gnd.n7549 gnd.n221 9.3005
R11360 gnd.n7551 gnd.n7550 9.3005
R11361 gnd.n206 gnd.n205 9.3005
R11362 gnd.n7564 gnd.n7563 9.3005
R11363 gnd.n7565 gnd.n204 9.3005
R11364 gnd.n7567 gnd.n7566 9.3005
R11365 gnd.n191 gnd.n190 9.3005
R11366 gnd.n7655 gnd.n7654 9.3005
R11367 gnd.n7656 gnd.n189 9.3005
R11368 gnd.n7658 gnd.n7657 9.3005
R11369 gnd.n111 gnd.n110 9.3005
R11370 gnd.n7738 gnd.n7737 9.3005
R11371 gnd.n1906 gnd.n1484 9.3005
R11372 gnd.n7502 gnd.n272 9.3005
R11373 gnd.n7503 gnd.n7502 9.3005
R11374 gnd.n2915 gnd.n2877 9.3005
R11375 gnd.n2914 gnd.n2883 9.3005
R11376 gnd.n2886 gnd.n2884 9.3005
R11377 gnd.n2910 gnd.n2887 9.3005
R11378 gnd.n2909 gnd.n2888 9.3005
R11379 gnd.n2908 gnd.n2889 9.3005
R11380 gnd.n2892 gnd.n2890 9.3005
R11381 gnd.n2904 gnd.n2893 9.3005
R11382 gnd.n2903 gnd.n2894 9.3005
R11383 gnd.n2902 gnd.n2895 9.3005
R11384 gnd.n2899 gnd.n2896 9.3005
R11385 gnd.n2898 gnd.n2897 9.3005
R11386 gnd.n2792 gnd.n2791 9.3005
R11387 gnd.n3242 gnd.n3241 9.3005
R11388 gnd.n3243 gnd.n2790 9.3005
R11389 gnd.n3245 gnd.n3244 9.3005
R11390 gnd.n2788 gnd.n2787 9.3005
R11391 gnd.n3250 gnd.n3249 9.3005
R11392 gnd.n3251 gnd.n2786 9.3005
R11393 gnd.n3253 gnd.n3252 9.3005
R11394 gnd.n2784 gnd.n2783 9.3005
R11395 gnd.n3258 gnd.n3257 9.3005
R11396 gnd.n3259 gnd.n2782 9.3005
R11397 gnd.n3261 gnd.n3260 9.3005
R11398 gnd.n2779 gnd.n2778 9.3005
R11399 gnd.n3401 gnd.n3400 9.3005
R11400 gnd.n3402 gnd.n2777 9.3005
R11401 gnd.n3404 gnd.n3403 9.3005
R11402 gnd.n2773 gnd.n2772 9.3005
R11403 gnd.n3415 gnd.n3414 9.3005
R11404 gnd.n3416 gnd.n2771 9.3005
R11405 gnd.n3418 gnd.n3417 9.3005
R11406 gnd.n2765 gnd.n2764 9.3005
R11407 gnd.n3429 gnd.n3428 9.3005
R11408 gnd.n3430 gnd.n2763 9.3005
R11409 gnd.n3432 gnd.n3431 9.3005
R11410 gnd.n2757 gnd.n2756 9.3005
R11411 gnd.n3446 gnd.n3445 9.3005
R11412 gnd.n3447 gnd.n2755 9.3005
R11413 gnd.n3449 gnd.n3448 9.3005
R11414 gnd.n2752 gnd.n2751 9.3005
R11415 gnd.n3460 gnd.n3459 9.3005
R11416 gnd.n3461 gnd.n2750 9.3005
R11417 gnd.n3465 gnd.n3462 9.3005
R11418 gnd.n3464 gnd.n3463 9.3005
R11419 gnd.n2398 gnd.n2397 9.3005
R11420 gnd.n3649 gnd.n3648 9.3005
R11421 gnd.n3650 gnd.n2396 9.3005
R11422 gnd.n3652 gnd.n3651 9.3005
R11423 gnd.n2377 gnd.n2376 9.3005
R11424 gnd.n3678 gnd.n3677 9.3005
R11425 gnd.n3679 gnd.n2375 9.3005
R11426 gnd.n3683 gnd.n3680 9.3005
R11427 gnd.n3682 gnd.n3681 9.3005
R11428 gnd.n2350 gnd.n2349 9.3005
R11429 gnd.n3716 gnd.n3715 9.3005
R11430 gnd.n3717 gnd.n2348 9.3005
R11431 gnd.n3721 gnd.n3718 9.3005
R11432 gnd.n3720 gnd.n3719 9.3005
R11433 gnd.n2323 gnd.n2322 9.3005
R11434 gnd.n3752 gnd.n3751 9.3005
R11435 gnd.n3753 gnd.n2321 9.3005
R11436 gnd.n3755 gnd.n3754 9.3005
R11437 gnd.n2301 gnd.n2300 9.3005
R11438 gnd.n3780 gnd.n3779 9.3005
R11439 gnd.n3781 gnd.n2299 9.3005
R11440 gnd.n3785 gnd.n3782 9.3005
R11441 gnd.n3784 gnd.n3783 9.3005
R11442 gnd.n2273 gnd.n2272 9.3005
R11443 gnd.n3830 gnd.n3829 9.3005
R11444 gnd.n3831 gnd.n2271 9.3005
R11445 gnd.n3835 gnd.n3832 9.3005
R11446 gnd.n3834 gnd.n3833 9.3005
R11447 gnd.n2254 gnd.n2253 9.3005
R11448 gnd.n3857 gnd.n3856 9.3005
R11449 gnd.n3858 gnd.n2252 9.3005
R11450 gnd.n3860 gnd.n3859 9.3005
R11451 gnd.n2209 gnd.n2208 9.3005
R11452 gnd.n3900 gnd.n3899 9.3005
R11453 gnd.n3901 gnd.n2207 9.3005
R11454 gnd.n3903 gnd.n3902 9.3005
R11455 gnd.n2187 gnd.n2186 9.3005
R11456 gnd.n3942 gnd.n3941 9.3005
R11457 gnd.n3943 gnd.n2185 9.3005
R11458 gnd.n3947 gnd.n3944 9.3005
R11459 gnd.n3946 gnd.n3945 9.3005
R11460 gnd.n2160 gnd.n2159 9.3005
R11461 gnd.n3994 gnd.n3993 9.3005
R11462 gnd.n3995 gnd.n2158 9.3005
R11463 gnd.n3999 gnd.n3996 9.3005
R11464 gnd.n3998 gnd.n3997 9.3005
R11465 gnd.n2129 gnd.n2128 9.3005
R11466 gnd.n4045 gnd.n4044 9.3005
R11467 gnd.n4046 gnd.n2127 9.3005
R11468 gnd.n4048 gnd.n4047 9.3005
R11469 gnd.n2114 gnd.n2113 9.3005
R11470 gnd.n4077 gnd.n4076 9.3005
R11471 gnd.n4078 gnd.n2112 9.3005
R11472 gnd.n4085 gnd.n4079 9.3005
R11473 gnd.n4084 gnd.n4080 9.3005
R11474 gnd.n4083 gnd.n4081 9.3005
R11475 gnd.n2079 gnd.n2078 9.3005
R11476 gnd.n4151 gnd.n4150 9.3005
R11477 gnd.n4152 gnd.n2077 9.3005
R11478 gnd.n4156 gnd.n4153 9.3005
R11479 gnd.n4155 gnd.n4154 9.3005
R11480 gnd.n2051 gnd.n2050 9.3005
R11481 gnd.n4194 gnd.n4193 9.3005
R11482 gnd.n4195 gnd.n2049 9.3005
R11483 gnd.n4202 gnd.n4196 9.3005
R11484 gnd.n4201 gnd.n4197 9.3005
R11485 gnd.n4200 gnd.n4198 9.3005
R11486 gnd.n1845 gnd.n1844 9.3005
R11487 gnd.n4380 gnd.n4379 9.3005
R11488 gnd.n4381 gnd.n1843 9.3005
R11489 gnd.n4383 gnd.n4382 9.3005
R11490 gnd.n1832 gnd.n1831 9.3005
R11491 gnd.n4400 gnd.n4399 9.3005
R11492 gnd.n4401 gnd.n1830 9.3005
R11493 gnd.n4403 gnd.n4402 9.3005
R11494 gnd.n1819 gnd.n1818 9.3005
R11495 gnd.n4420 gnd.n4419 9.3005
R11496 gnd.n4421 gnd.n1817 9.3005
R11497 gnd.n4423 gnd.n4422 9.3005
R11498 gnd.n1806 gnd.n1805 9.3005
R11499 gnd.n4443 gnd.n4442 9.3005
R11500 gnd.n4444 gnd.n1804 9.3005
R11501 gnd.n4447 gnd.n4446 9.3005
R11502 gnd.n4445 gnd.n1461 9.3005
R11503 gnd.n4734 gnd.n1462 9.3005
R11504 gnd.n4733 gnd.n1463 9.3005
R11505 gnd.n4732 gnd.n1464 9.3005
R11506 gnd.n1470 gnd.n1465 9.3005
R11507 gnd.n4726 gnd.n1471 9.3005
R11508 gnd.n4725 gnd.n1472 9.3005
R11509 gnd.n4724 gnd.n1473 9.3005
R11510 gnd.n1626 gnd.n1474 9.3005
R11511 gnd.n1629 gnd.n1628 9.3005
R11512 gnd.n1630 gnd.n1625 9.3005
R11513 gnd.n1632 gnd.n1631 9.3005
R11514 gnd.n1614 gnd.n1613 9.3005
R11515 gnd.n4538 gnd.n4537 9.3005
R11516 gnd.n4539 gnd.n1612 9.3005
R11517 gnd.n4543 gnd.n4540 9.3005
R11518 gnd.n4542 gnd.n4541 9.3005
R11519 gnd.n1587 gnd.n1586 9.3005
R11520 gnd.n4571 gnd.n4570 9.3005
R11521 gnd.n4572 gnd.n1585 9.3005
R11522 gnd.n4583 gnd.n4573 9.3005
R11523 gnd.n4582 gnd.n4574 9.3005
R11524 gnd.n4581 gnd.n4575 9.3005
R11525 gnd.n4578 gnd.n4577 9.3005
R11526 gnd.n4576 gnd.n1532 9.3005
R11527 gnd.n4673 gnd.n1533 9.3005
R11528 gnd.n4672 gnd.n1534 9.3005
R11529 gnd.n4671 gnd.n1535 9.3005
R11530 gnd.n1537 gnd.n1536 9.3005
R11531 gnd.n7465 gnd.n309 9.3005
R11532 gnd.n312 gnd.n310 9.3005
R11533 gnd.n7461 gnd.n313 9.3005
R11534 gnd.n7460 gnd.n314 9.3005
R11535 gnd.n7459 gnd.n315 9.3005
R11536 gnd.n318 gnd.n316 9.3005
R11537 gnd.n7398 gnd.n319 9.3005
R11538 gnd.n7397 gnd.n320 9.3005
R11539 gnd.n7396 gnd.n321 9.3005
R11540 gnd.n2608 gnd.n2604 9.3005
R11541 gnd.n2641 gnd.n2638 9.3005
R11542 gnd.n2642 gnd.n2637 9.3005
R11543 gnd.n2645 gnd.n2636 9.3005
R11544 gnd.n2646 gnd.n2635 9.3005
R11545 gnd.n2649 gnd.n2634 9.3005
R11546 gnd.n2650 gnd.n2633 9.3005
R11547 gnd.n2653 gnd.n2632 9.3005
R11548 gnd.n2654 gnd.n2631 9.3005
R11549 gnd.n2657 gnd.n2630 9.3005
R11550 gnd.n2658 gnd.n2629 9.3005
R11551 gnd.n2661 gnd.n2628 9.3005
R11552 gnd.n2662 gnd.n2627 9.3005
R11553 gnd.n2663 gnd.n2626 9.3005
R11554 gnd.n2625 gnd.n2622 9.3005
R11555 gnd.n2624 gnd.n2623 9.3005
R11556 gnd.n3570 gnd.n3569 9.3005
R11557 gnd.n2610 gnd.n2609 9.3005
R11558 gnd.n2669 gnd.n2667 9.3005
R11559 gnd.n3562 gnd.n2670 9.3005
R11560 gnd.n3561 gnd.n2671 9.3005
R11561 gnd.n3560 gnd.n2672 9.3005
R11562 gnd.n2676 gnd.n2673 9.3005
R11563 gnd.n3555 gnd.n2677 9.3005
R11564 gnd.n3554 gnd.n2678 9.3005
R11565 gnd.n3553 gnd.n2679 9.3005
R11566 gnd.n2683 gnd.n2680 9.3005
R11567 gnd.n3548 gnd.n2684 9.3005
R11568 gnd.n3547 gnd.n2685 9.3005
R11569 gnd.n3546 gnd.n2686 9.3005
R11570 gnd.n2690 gnd.n2687 9.3005
R11571 gnd.n3541 gnd.n2691 9.3005
R11572 gnd.n3540 gnd.n2692 9.3005
R11573 gnd.n3539 gnd.n2693 9.3005
R11574 gnd.n2698 gnd.n2696 9.3005
R11575 gnd.n3534 gnd.n3533 9.3005
R11576 gnd.n3571 gnd.n2603 9.3005
R11577 gnd.n2982 gnd.n2956 9.3005
R11578 gnd.n3041 gnd.n2957 9.3005
R11579 gnd.n3042 gnd.n2955 9.3005
R11580 gnd.n3045 gnd.n3044 9.3005
R11581 gnd.n3046 gnd.n2954 9.3005
R11582 gnd.n3049 gnd.n3047 9.3005
R11583 gnd.n3050 gnd.n2953 9.3005
R11584 gnd.n3053 gnd.n3052 9.3005
R11585 gnd.n3054 gnd.n2952 9.3005
R11586 gnd.n3057 gnd.n3055 9.3005
R11587 gnd.n3058 gnd.n2951 9.3005
R11588 gnd.n3082 gnd.n3081 9.3005
R11589 gnd.n3083 gnd.n2950 9.3005
R11590 gnd.n3085 gnd.n3084 9.3005
R11591 gnd.n2946 gnd.n2945 9.3005
R11592 gnd.n3098 gnd.n3097 9.3005
R11593 gnd.n3099 gnd.n2944 9.3005
R11594 gnd.n3101 gnd.n3100 9.3005
R11595 gnd.n2846 gnd.n2845 9.3005
R11596 gnd.n3114 gnd.n3113 9.3005
R11597 gnd.n3115 gnd.n2844 9.3005
R11598 gnd.n3117 gnd.n3116 9.3005
R11599 gnd.n2840 gnd.n2839 9.3005
R11600 gnd.n3130 gnd.n3129 9.3005
R11601 gnd.n3131 gnd.n2838 9.3005
R11602 gnd.n3134 gnd.n3133 9.3005
R11603 gnd.n2984 gnd.n2983 9.3005
R11604 gnd.n2989 gnd.n2988 9.3005
R11605 gnd.n2992 gnd.n2977 9.3005
R11606 gnd.n2993 gnd.n2976 9.3005
R11607 gnd.n2996 gnd.n2975 9.3005
R11608 gnd.n2997 gnd.n2974 9.3005
R11609 gnd.n3000 gnd.n2973 9.3005
R11610 gnd.n3001 gnd.n2972 9.3005
R11611 gnd.n3004 gnd.n2971 9.3005
R11612 gnd.n3005 gnd.n2970 9.3005
R11613 gnd.n3008 gnd.n2969 9.3005
R11614 gnd.n3009 gnd.n2968 9.3005
R11615 gnd.n3012 gnd.n2967 9.3005
R11616 gnd.n3013 gnd.n2966 9.3005
R11617 gnd.n3016 gnd.n2965 9.3005
R11618 gnd.n3017 gnd.n2964 9.3005
R11619 gnd.n3020 gnd.n2963 9.3005
R11620 gnd.n3023 gnd.n3022 9.3005
R11621 gnd.n2987 gnd.n2981 9.3005
R11622 gnd.n2986 gnd.n2985 9.3005
R11623 gnd.n3030 gnd.n3029 9.3005
R11624 gnd.n3028 gnd.n2962 9.3005
R11625 gnd.n3027 gnd.n3026 9.3005
R11626 gnd.n3025 gnd.n1080 9.3005
R11627 gnd.n5040 gnd.n1081 9.3005
R11628 gnd.n5039 gnd.n1082 9.3005
R11629 gnd.n5038 gnd.n1083 9.3005
R11630 gnd.n1099 gnd.n1084 9.3005
R11631 gnd.n5028 gnd.n1100 9.3005
R11632 gnd.n5027 gnd.n1101 9.3005
R11633 gnd.n5026 gnd.n1102 9.3005
R11634 gnd.n1121 gnd.n1103 9.3005
R11635 gnd.n5016 gnd.n1122 9.3005
R11636 gnd.n5015 gnd.n1123 9.3005
R11637 gnd.n5014 gnd.n1124 9.3005
R11638 gnd.n1142 gnd.n1125 9.3005
R11639 gnd.n5004 gnd.n1143 9.3005
R11640 gnd.n5003 gnd.n1144 9.3005
R11641 gnd.n5002 gnd.n1145 9.3005
R11642 gnd.n1163 gnd.n1146 9.3005
R11643 gnd.n4992 gnd.n1164 9.3005
R11644 gnd.n4991 gnd.n1165 9.3005
R11645 gnd.n4990 gnd.n1166 9.3005
R11646 gnd.n1182 gnd.n1167 9.3005
R11647 gnd.n4980 gnd.n1183 9.3005
R11648 gnd.n4979 gnd.n1184 9.3005
R11649 gnd.n4978 gnd.n1185 9.3005
R11650 gnd.n1200 gnd.n1186 9.3005
R11651 gnd.n4967 gnd.n1201 9.3005
R11652 gnd.n4966 gnd.n1202 9.3005
R11653 gnd.n4965 gnd.n1203 9.3005
R11654 gnd.n1220 gnd.n1204 9.3005
R11655 gnd.n4955 gnd.n1221 9.3005
R11656 gnd.n4954 gnd.n1222 9.3005
R11657 gnd.n4953 gnd.n1223 9.3005
R11658 gnd.n1241 gnd.n1224 9.3005
R11659 gnd.n4943 gnd.n1242 9.3005
R11660 gnd.n4942 gnd.n1243 9.3005
R11661 gnd.n4941 gnd.n1244 9.3005
R11662 gnd.n1262 gnd.n1245 9.3005
R11663 gnd.n4931 gnd.n1263 9.3005
R11664 gnd.n4930 gnd.n1264 9.3005
R11665 gnd.n4929 gnd.n1265 9.3005
R11666 gnd.n1283 gnd.n1266 9.3005
R11667 gnd.n4919 gnd.n1284 9.3005
R11668 gnd.n4918 gnd.n1285 9.3005
R11669 gnd.n4917 gnd.n1286 9.3005
R11670 gnd.n1305 gnd.n1287 9.3005
R11671 gnd.n4907 gnd.n1306 9.3005
R11672 gnd.n4906 gnd.n1307 9.3005
R11673 gnd.n4905 gnd.n1308 9.3005
R11674 gnd.n1325 gnd.n1309 9.3005
R11675 gnd.n4895 gnd.n4894 9.3005
R11676 gnd.n3024 gnd.n2961 9.3005
R11677 gnd.n5054 gnd.n5053 9.3005
R11678 gnd.n5052 gnd.n1058 9.3005
R11679 gnd.n5051 gnd.n5050 9.3005
R11680 gnd.n1060 gnd.n1059 9.3005
R11681 gnd.n3063 gnd.n3062 9.3005
R11682 gnd.n3066 gnd.n3065 9.3005
R11683 gnd.n3067 gnd.n3061 9.3005
R11684 gnd.n3070 gnd.n3068 9.3005
R11685 gnd.n3071 gnd.n3060 9.3005
R11686 gnd.n3074 gnd.n3073 9.3005
R11687 gnd.n3075 gnd.n3059 9.3005
R11688 gnd.n3077 gnd.n3076 9.3005
R11689 gnd.n2949 gnd.n2948 9.3005
R11690 gnd.n3090 gnd.n3089 9.3005
R11691 gnd.n3091 gnd.n2947 9.3005
R11692 gnd.n3093 gnd.n3092 9.3005
R11693 gnd.n2850 gnd.n2849 9.3005
R11694 gnd.n3106 gnd.n3105 9.3005
R11695 gnd.n3107 gnd.n2848 9.3005
R11696 gnd.n3109 gnd.n3108 9.3005
R11697 gnd.n2843 gnd.n2842 9.3005
R11698 gnd.n3122 gnd.n3121 9.3005
R11699 gnd.n3123 gnd.n2841 9.3005
R11700 gnd.n3125 gnd.n3124 9.3005
R11701 gnd.n2836 gnd.n2835 9.3005
R11702 gnd.n3139 gnd.n3138 9.3005
R11703 gnd.n3141 gnd.n2833 9.3005
R11704 gnd.n3143 gnd.n3142 9.3005
R11705 gnd.n2828 gnd.n2827 9.3005
R11706 gnd.n3156 gnd.n3155 9.3005
R11707 gnd.n3157 gnd.n2826 9.3005
R11708 gnd.n3159 gnd.n3158 9.3005
R11709 gnd.n2821 gnd.n2820 9.3005
R11710 gnd.n3172 gnd.n3171 9.3005
R11711 gnd.n3173 gnd.n2819 9.3005
R11712 gnd.n3175 gnd.n3174 9.3005
R11713 gnd.n2814 gnd.n2813 9.3005
R11714 gnd.n3188 gnd.n3187 9.3005
R11715 gnd.n3189 gnd.n2812 9.3005
R11716 gnd.n3192 gnd.n3191 9.3005
R11717 gnd.n3190 gnd.n2806 9.3005
R11718 gnd.n3204 gnd.n2807 9.3005
R11719 gnd.n3205 gnd.n2805 9.3005
R11720 gnd.n3207 gnd.n3206 9.3005
R11721 gnd.n3208 gnd.n2804 9.3005
R11722 gnd.n3212 gnd.n3209 9.3005
R11723 gnd.n3213 gnd.n2803 9.3005
R11724 gnd.n3217 gnd.n3216 9.3005
R11725 gnd.n3218 gnd.n2802 9.3005
R11726 gnd.n3221 gnd.n3220 9.3005
R11727 gnd.n3219 gnd.n2700 9.3005
R11728 gnd.n3530 gnd.n2699 9.3005
R11729 gnd.n3532 gnd.n3531 9.3005
R11730 gnd.n5055 gnd.n1056 9.3005
R11731 gnd.n5062 gnd.n5061 9.3005
R11732 gnd.n5063 gnd.n1050 9.3005
R11733 gnd.n5066 gnd.n1049 9.3005
R11734 gnd.n5067 gnd.n1048 9.3005
R11735 gnd.n5070 gnd.n1047 9.3005
R11736 gnd.n5071 gnd.n1046 9.3005
R11737 gnd.n5074 gnd.n1045 9.3005
R11738 gnd.n5075 gnd.n1044 9.3005
R11739 gnd.n5078 gnd.n1043 9.3005
R11740 gnd.n5079 gnd.n1042 9.3005
R11741 gnd.n5082 gnd.n1041 9.3005
R11742 gnd.n5083 gnd.n1040 9.3005
R11743 gnd.n5086 gnd.n1039 9.3005
R11744 gnd.n5087 gnd.n1038 9.3005
R11745 gnd.n5090 gnd.n1037 9.3005
R11746 gnd.n5091 gnd.n1036 9.3005
R11747 gnd.n5094 gnd.n1035 9.3005
R11748 gnd.n5095 gnd.n1034 9.3005
R11749 gnd.n5098 gnd.n1033 9.3005
R11750 gnd.n5100 gnd.n1030 9.3005
R11751 gnd.n5103 gnd.n1029 9.3005
R11752 gnd.n5104 gnd.n1028 9.3005
R11753 gnd.n5107 gnd.n1027 9.3005
R11754 gnd.n5108 gnd.n1026 9.3005
R11755 gnd.n5111 gnd.n1025 9.3005
R11756 gnd.n5112 gnd.n1024 9.3005
R11757 gnd.n5115 gnd.n1023 9.3005
R11758 gnd.n5116 gnd.n1022 9.3005
R11759 gnd.n5119 gnd.n1021 9.3005
R11760 gnd.n5120 gnd.n1020 9.3005
R11761 gnd.n5123 gnd.n1019 9.3005
R11762 gnd.n5124 gnd.n1018 9.3005
R11763 gnd.n5127 gnd.n1017 9.3005
R11764 gnd.n5129 gnd.n1016 9.3005
R11765 gnd.n5130 gnd.n1015 9.3005
R11766 gnd.n5131 gnd.n1014 9.3005
R11767 gnd.n5132 gnd.n1013 9.3005
R11768 gnd.n5060 gnd.n1055 9.3005
R11769 gnd.n5059 gnd.n5058 9.3005
R11770 gnd.n3036 gnd.n3035 9.3005
R11771 gnd.n3034 gnd.n1069 9.3005
R11772 gnd.n5046 gnd.n1070 9.3005
R11773 gnd.n5045 gnd.n1071 9.3005
R11774 gnd.n5044 gnd.n1072 9.3005
R11775 gnd.n1090 gnd.n1073 9.3005
R11776 gnd.n5034 gnd.n1091 9.3005
R11777 gnd.n5033 gnd.n1092 9.3005
R11778 gnd.n5032 gnd.n1093 9.3005
R11779 gnd.n1110 gnd.n1094 9.3005
R11780 gnd.n5022 gnd.n1111 9.3005
R11781 gnd.n5021 gnd.n1112 9.3005
R11782 gnd.n5020 gnd.n1113 9.3005
R11783 gnd.n1132 gnd.n1114 9.3005
R11784 gnd.n5010 gnd.n1133 9.3005
R11785 gnd.n5009 gnd.n1134 9.3005
R11786 gnd.n5008 gnd.n1135 9.3005
R11787 gnd.n1152 gnd.n1136 9.3005
R11788 gnd.n4998 gnd.n1153 9.3005
R11789 gnd.n4997 gnd.n1154 9.3005
R11790 gnd.n4996 gnd.n1155 9.3005
R11791 gnd.n4960 gnd.n1212 9.3005
R11792 gnd.n4959 gnd.n1213 9.3005
R11793 gnd.n1230 gnd.n1214 9.3005
R11794 gnd.n4949 gnd.n1231 9.3005
R11795 gnd.n4948 gnd.n1232 9.3005
R11796 gnd.n4947 gnd.n1233 9.3005
R11797 gnd.n1252 gnd.n1234 9.3005
R11798 gnd.n4937 gnd.n1253 9.3005
R11799 gnd.n4936 gnd.n1254 9.3005
R11800 gnd.n4935 gnd.n1255 9.3005
R11801 gnd.n1272 gnd.n1256 9.3005
R11802 gnd.n4925 gnd.n1273 9.3005
R11803 gnd.n4924 gnd.n1274 9.3005
R11804 gnd.n4923 gnd.n1275 9.3005
R11805 gnd.n1294 gnd.n1276 9.3005
R11806 gnd.n4913 gnd.n1295 9.3005
R11807 gnd.n4912 gnd.n1296 9.3005
R11808 gnd.n4911 gnd.n1297 9.3005
R11809 gnd.n1315 gnd.n1298 9.3005
R11810 gnd.n4901 gnd.n1316 9.3005
R11811 gnd.n4900 gnd.n1317 9.3005
R11812 gnd.n4899 gnd.n1318 9.3005
R11813 gnd.n3033 gnd.n3032 9.3005
R11814 gnd.n4985 gnd.n1175 9.3005
R11815 gnd.n4961 gnd.n1175 9.3005
R11816 gnd.n2864 gnd.n2863 9.3005
R11817 gnd.n2855 gnd.n2854 9.3005
R11818 gnd.n2869 gnd.n2868 9.3005
R11819 gnd.n2870 gnd.n2853 9.3005
R11820 gnd.n2941 gnd.n2871 9.3005
R11821 gnd.n2940 gnd.n2872 9.3005
R11822 gnd.n2939 gnd.n2873 9.3005
R11823 gnd.n2932 gnd.n2874 9.3005
R11824 gnd.n2862 gnd.n2857 9.3005
R11825 gnd.n2858 gnd.n905 9.3005
R11826 gnd.n6528 gnd.n904 9.3005
R11827 gnd.n6529 gnd.n903 9.3005
R11828 gnd.n6530 gnd.n902 9.3005
R11829 gnd.n901 gnd.n897 9.3005
R11830 gnd.n6536 gnd.n896 9.3005
R11831 gnd.n6537 gnd.n895 9.3005
R11832 gnd.n6538 gnd.n894 9.3005
R11833 gnd.n893 gnd.n889 9.3005
R11834 gnd.n6544 gnd.n888 9.3005
R11835 gnd.n6545 gnd.n887 9.3005
R11836 gnd.n6546 gnd.n886 9.3005
R11837 gnd.n885 gnd.n881 9.3005
R11838 gnd.n6552 gnd.n880 9.3005
R11839 gnd.n6553 gnd.n879 9.3005
R11840 gnd.n6554 gnd.n878 9.3005
R11841 gnd.n877 gnd.n873 9.3005
R11842 gnd.n6560 gnd.n872 9.3005
R11843 gnd.n6561 gnd.n871 9.3005
R11844 gnd.n6562 gnd.n870 9.3005
R11845 gnd.n869 gnd.n865 9.3005
R11846 gnd.n6568 gnd.n864 9.3005
R11847 gnd.n6569 gnd.n863 9.3005
R11848 gnd.n6570 gnd.n862 9.3005
R11849 gnd.n861 gnd.n857 9.3005
R11850 gnd.n6576 gnd.n856 9.3005
R11851 gnd.n6577 gnd.n855 9.3005
R11852 gnd.n6578 gnd.n854 9.3005
R11853 gnd.n853 gnd.n849 9.3005
R11854 gnd.n6584 gnd.n848 9.3005
R11855 gnd.n6585 gnd.n847 9.3005
R11856 gnd.n6586 gnd.n846 9.3005
R11857 gnd.n845 gnd.n841 9.3005
R11858 gnd.n6592 gnd.n840 9.3005
R11859 gnd.n6593 gnd.n839 9.3005
R11860 gnd.n6594 gnd.n838 9.3005
R11861 gnd.n837 gnd.n833 9.3005
R11862 gnd.n6600 gnd.n832 9.3005
R11863 gnd.n6601 gnd.n831 9.3005
R11864 gnd.n6602 gnd.n830 9.3005
R11865 gnd.n829 gnd.n825 9.3005
R11866 gnd.n6608 gnd.n824 9.3005
R11867 gnd.n6609 gnd.n823 9.3005
R11868 gnd.n6610 gnd.n822 9.3005
R11869 gnd.n821 gnd.n817 9.3005
R11870 gnd.n6616 gnd.n816 9.3005
R11871 gnd.n6617 gnd.n815 9.3005
R11872 gnd.n6618 gnd.n814 9.3005
R11873 gnd.n813 gnd.n809 9.3005
R11874 gnd.n6624 gnd.n808 9.3005
R11875 gnd.n6625 gnd.n807 9.3005
R11876 gnd.n6626 gnd.n806 9.3005
R11877 gnd.n805 gnd.n801 9.3005
R11878 gnd.n6632 gnd.n800 9.3005
R11879 gnd.n6633 gnd.n799 9.3005
R11880 gnd.n6634 gnd.n798 9.3005
R11881 gnd.n797 gnd.n793 9.3005
R11882 gnd.n6640 gnd.n792 9.3005
R11883 gnd.n6641 gnd.n791 9.3005
R11884 gnd.n6642 gnd.n790 9.3005
R11885 gnd.n789 gnd.n785 9.3005
R11886 gnd.n6648 gnd.n784 9.3005
R11887 gnd.n6649 gnd.n783 9.3005
R11888 gnd.n6650 gnd.n782 9.3005
R11889 gnd.n781 gnd.n777 9.3005
R11890 gnd.n6656 gnd.n776 9.3005
R11891 gnd.n6657 gnd.n775 9.3005
R11892 gnd.n6658 gnd.n774 9.3005
R11893 gnd.n773 gnd.n769 9.3005
R11894 gnd.n6664 gnd.n768 9.3005
R11895 gnd.n6665 gnd.n767 9.3005
R11896 gnd.n6666 gnd.n766 9.3005
R11897 gnd.n765 gnd.n761 9.3005
R11898 gnd.n6672 gnd.n760 9.3005
R11899 gnd.n6673 gnd.n759 9.3005
R11900 gnd.n6674 gnd.n758 9.3005
R11901 gnd.n757 gnd.n753 9.3005
R11902 gnd.n6680 gnd.n752 9.3005
R11903 gnd.n6681 gnd.n751 9.3005
R11904 gnd.n6682 gnd.n750 9.3005
R11905 gnd.n749 gnd.n745 9.3005
R11906 gnd.n6688 gnd.n744 9.3005
R11907 gnd.n6689 gnd.n743 9.3005
R11908 gnd.n6690 gnd.n742 9.3005
R11909 gnd.n2861 gnd.n2860 9.3005
R11910 gnd.n1702 gnd.n1701 9.3005
R11911 gnd.n1680 gnd.n1679 9.3005
R11912 gnd.n1714 gnd.n1713 9.3005
R11913 gnd.n1677 gnd.n1675 9.3005
R11914 gnd.n1721 gnd.n1720 9.3005
R11915 gnd.n1671 gnd.n1670 9.3005
R11916 gnd.n1733 gnd.n1732 9.3005
R11917 gnd.n1668 gnd.n1666 9.3005
R11918 gnd.n1740 gnd.n1739 9.3005
R11919 gnd.n1662 gnd.n1661 9.3005
R11920 gnd.n1752 gnd.n1751 9.3005
R11921 gnd.n1659 gnd.n1657 9.3005
R11922 gnd.n1759 gnd.n1758 9.3005
R11923 gnd.n1653 gnd.n1652 9.3005
R11924 gnd.n1771 gnd.n1770 9.3005
R11925 gnd.n1650 gnd.n1648 9.3005
R11926 gnd.n4472 gnd.n4471 9.3005
R11927 gnd.n4470 gnd.n1649 9.3005
R11928 gnd.n1697 gnd.n1695 9.3005
R11929 gnd.n1768 gnd.n1767 9.3005
R11930 gnd.n1658 gnd.n1654 9.3005
R11931 gnd.n1761 gnd.n1760 9.3005
R11932 gnd.n1750 gnd.n1656 9.3005
R11933 gnd.n1749 gnd.n1748 9.3005
R11934 gnd.n1667 gnd.n1663 9.3005
R11935 gnd.n1742 gnd.n1741 9.3005
R11936 gnd.n1731 gnd.n1665 9.3005
R11937 gnd.n1730 gnd.n1729 9.3005
R11938 gnd.n1676 gnd.n1672 9.3005
R11939 gnd.n1723 gnd.n1722 9.3005
R11940 gnd.n1712 gnd.n1674 9.3005
R11941 gnd.n1711 gnd.n1710 9.3005
R11942 gnd.n1696 gnd.n1681 9.3005
R11943 gnd.n1704 gnd.n1703 9.3005
R11944 gnd.n1694 gnd.n1683 9.3005
R11945 gnd.n1769 gnd.n1647 9.3005
R11946 gnd.n4474 gnd.n4473 9.3005
R11947 gnd.n4469 gnd.n4468 9.3005
R11948 gnd.n4467 gnd.n1779 9.3005
R11949 gnd.n4466 gnd.n4465 9.3005
R11950 gnd.n4464 gnd.n1780 9.3005
R11951 gnd.n4463 gnd.n4462 9.3005
R11952 gnd.n4461 gnd.n1787 9.3005
R11953 gnd.n4460 gnd.n4459 9.3005
R11954 gnd.n4458 gnd.n1788 9.3005
R11955 gnd.n4457 gnd.n4456 9.3005
R11956 gnd.n4455 gnd.n1799 9.3005
R11957 gnd.n3503 gnd.n2724 9.3005
R11958 gnd.n3502 gnd.n3501 9.3005
R11959 gnd.n3500 gnd.n2728 9.3005
R11960 gnd.n3499 gnd.n3498 9.3005
R11961 gnd.n3497 gnd.n2729 9.3005
R11962 gnd.n3496 gnd.n3495 9.3005
R11963 gnd.n3494 gnd.n2733 9.3005
R11964 gnd.n3493 gnd.n3492 9.3005
R11965 gnd.n3491 gnd.n2734 9.3005
R11966 gnd.n3490 gnd.n3489 9.3005
R11967 gnd.n3488 gnd.n2738 9.3005
R11968 gnd.n3487 gnd.n3486 9.3005
R11969 gnd.n3485 gnd.n2739 9.3005
R11970 gnd.n3484 gnd.n3483 9.3005
R11971 gnd.n3482 gnd.n2743 9.3005
R11972 gnd.n3481 gnd.n3480 9.3005
R11973 gnd.n3479 gnd.n2744 9.3005
R11974 gnd.n3478 gnd.n3477 9.3005
R11975 gnd.n3476 gnd.n3475 9.3005
R11976 gnd.n2384 gnd.n2383 9.3005
R11977 gnd.n3667 gnd.n3666 9.3005
R11978 gnd.n3668 gnd.n2382 9.3005
R11979 gnd.n3670 gnd.n3669 9.3005
R11980 gnd.n2364 gnd.n2363 9.3005
R11981 gnd.n3697 gnd.n3696 9.3005
R11982 gnd.n3698 gnd.n2361 9.3005
R11983 gnd.n3701 gnd.n3700 9.3005
R11984 gnd.n3699 gnd.n2362 9.3005
R11985 gnd.n2337 gnd.n2336 9.3005
R11986 gnd.n3734 gnd.n3733 9.3005
R11987 gnd.n3735 gnd.n2335 9.3005
R11988 gnd.n3737 gnd.n3736 9.3005
R11989 gnd.n2317 gnd.n2316 9.3005
R11990 gnd.n3761 gnd.n3760 9.3005
R11991 gnd.n3762 gnd.n2314 9.3005
R11992 gnd.n3765 gnd.n3764 9.3005
R11993 gnd.n3763 gnd.n2315 9.3005
R11994 gnd.n2287 gnd.n2286 9.3005
R11995 gnd.n3800 gnd.n3799 9.3005
R11996 gnd.n3801 gnd.n2284 9.3005
R11997 gnd.n3817 gnd.n3816 9.3005
R11998 gnd.n3815 gnd.n2285 9.3005
R11999 gnd.n3814 gnd.n3813 9.3005
R12000 gnd.n3812 gnd.n3802 9.3005
R12001 gnd.n3811 gnd.n3810 9.3005
R12002 gnd.n3809 gnd.n3808 9.3005
R12003 gnd.n2225 gnd.n2224 9.3005
R12004 gnd.n3882 gnd.n3881 9.3005
R12005 gnd.n3883 gnd.n2222 9.3005
R12006 gnd.n3886 gnd.n3885 9.3005
R12007 gnd.n3884 gnd.n2223 9.3005
R12008 gnd.n2195 gnd.n2194 9.3005
R12009 gnd.n3918 gnd.n3917 9.3005
R12010 gnd.n3919 gnd.n2192 9.3005
R12011 gnd.n3934 gnd.n3933 9.3005
R12012 gnd.n3932 gnd.n2193 9.3005
R12013 gnd.n3931 gnd.n3930 9.3005
R12014 gnd.n3929 gnd.n3920 9.3005
R12015 gnd.n3928 gnd.n3927 9.3005
R12016 gnd.n3926 gnd.n3925 9.3005
R12017 gnd.n2146 gnd.n2145 9.3005
R12018 gnd.n4012 gnd.n4011 9.3005
R12019 gnd.n4013 gnd.n2143 9.3005
R12020 gnd.n4030 gnd.n4029 9.3005
R12021 gnd.n4028 gnd.n2144 9.3005
R12022 gnd.n4027 gnd.n4026 9.3005
R12023 gnd.n4025 gnd.n4014 9.3005
R12024 gnd.n4024 gnd.n4023 9.3005
R12025 gnd.n4022 gnd.n4021 9.3005
R12026 gnd.n2097 gnd.n2096 9.3005
R12027 gnd.n4101 gnd.n4100 9.3005
R12028 gnd.n4102 gnd.n2094 9.3005
R12029 gnd.n4108 gnd.n4107 9.3005
R12030 gnd.n4106 gnd.n2095 9.3005
R12031 gnd.n4105 gnd.n4104 9.3005
R12032 gnd.n2066 gnd.n2065 9.3005
R12033 gnd.n4169 gnd.n4168 9.3005
R12034 gnd.n4170 gnd.n2063 9.3005
R12035 gnd.n4179 gnd.n4178 9.3005
R12036 gnd.n4177 gnd.n2064 9.3005
R12037 gnd.n4176 gnd.n4175 9.3005
R12038 gnd.n4174 gnd.n4171 9.3005
R12039 gnd.n1850 gnd.n1849 9.3005
R12040 gnd.n4370 gnd.n4369 9.3005
R12041 gnd.n4371 gnd.n1848 9.3005
R12042 gnd.n4373 gnd.n4372 9.3005
R12043 gnd.n1838 gnd.n1837 9.3005
R12044 gnd.n4390 gnd.n4389 9.3005
R12045 gnd.n4391 gnd.n1836 9.3005
R12046 gnd.n4393 gnd.n4392 9.3005
R12047 gnd.n1825 gnd.n1824 9.3005
R12048 gnd.n4410 gnd.n4409 9.3005
R12049 gnd.n4411 gnd.n1823 9.3005
R12050 gnd.n4413 gnd.n4412 9.3005
R12051 gnd.n1812 gnd.n1811 9.3005
R12052 gnd.n4430 gnd.n4429 9.3005
R12053 gnd.n4431 gnd.n1810 9.3005
R12054 gnd.n4434 gnd.n4433 9.3005
R12055 gnd.n4432 gnd.n1801 9.3005
R12056 gnd.n4452 gnd.n1800 9.3005
R12057 gnd.n4454 gnd.n4453 9.3005
R12058 gnd.n3505 gnd.n3504 9.3005
R12059 gnd.n3508 gnd.n3507 9.3005
R12060 gnd.n3509 gnd.n2719 9.3005
R12061 gnd.n3511 gnd.n3510 9.3005
R12062 gnd.n3513 gnd.n3512 9.3005
R12063 gnd.n3514 gnd.n2712 9.3005
R12064 gnd.n3516 gnd.n3515 9.3005
R12065 gnd.n3517 gnd.n2711 9.3005
R12066 gnd.n3519 gnd.n3518 9.3005
R12067 gnd.n3520 gnd.n2705 9.3005
R12068 gnd.n3506 gnd.n2723 9.3005
R12069 gnd.n2831 gnd.n2830 9.3005
R12070 gnd.n3148 gnd.n3147 9.3005
R12071 gnd.n3149 gnd.n2829 9.3005
R12072 gnd.n3151 gnd.n3150 9.3005
R12073 gnd.n2825 gnd.n2824 9.3005
R12074 gnd.n3164 gnd.n3163 9.3005
R12075 gnd.n3165 gnd.n2823 9.3005
R12076 gnd.n3167 gnd.n3166 9.3005
R12077 gnd.n2817 gnd.n2816 9.3005
R12078 gnd.n3180 gnd.n3179 9.3005
R12079 gnd.n3181 gnd.n2815 9.3005
R12080 gnd.n3183 gnd.n3182 9.3005
R12081 gnd.n2811 gnd.n2810 9.3005
R12082 gnd.n3197 gnd.n3196 9.3005
R12083 gnd.n3198 gnd.n2809 9.3005
R12084 gnd.n3200 gnd.n3199 9.3005
R12085 gnd.n2797 gnd.n2795 9.3005
R12086 gnd.n3235 gnd.n3234 9.3005
R12087 gnd.n3233 gnd.n2796 9.3005
R12088 gnd.n3232 gnd.n3231 9.3005
R12089 gnd.n3230 gnd.n2798 9.3005
R12090 gnd.n3229 gnd.n3228 9.3005
R12091 gnd.n3227 gnd.n2801 9.3005
R12092 gnd.n3226 gnd.n3225 9.3005
R12093 gnd.n2704 gnd.n2702 9.3005
R12094 gnd.n3526 gnd.n3525 9.3005
R12095 gnd.n3524 gnd.n2703 9.3005
R12096 gnd.n3522 gnd.n3521 9.3005
R12097 gnd.n2707 gnd.n2706 9.3005
R12098 gnd.n3353 gnd.n3352 9.3005
R12099 gnd.n3355 gnd.n3354 9.3005
R12100 gnd.n3333 gnd.n3332 9.3005
R12101 gnd.n3361 gnd.n3360 9.3005
R12102 gnd.n3363 gnd.n3362 9.3005
R12103 gnd.n3323 gnd.n3322 9.3005
R12104 gnd.n3369 gnd.n3368 9.3005
R12105 gnd.n3371 gnd.n3370 9.3005
R12106 gnd.n3310 gnd.n3309 9.3005
R12107 gnd.n3377 gnd.n3376 9.3005
R12108 gnd.n3379 gnd.n3378 9.3005
R12109 gnd.n3300 gnd.n3299 9.3005
R12110 gnd.n3385 gnd.n3384 9.3005
R12111 gnd.n3387 gnd.n3386 9.3005
R12112 gnd.n3285 gnd.n3283 9.3005
R12113 gnd.n3393 gnd.n3392 9.3005
R12114 gnd.n3394 gnd.n3282 9.3005
R12115 gnd.n3287 gnd.n1327 9.3005
R12116 gnd.n3286 gnd.n3284 9.3005
R12117 gnd.n3391 gnd.n3390 9.3005
R12118 gnd.n3389 gnd.n3388 9.3005
R12119 gnd.n3295 gnd.n3294 9.3005
R12120 gnd.n3383 gnd.n3382 9.3005
R12121 gnd.n3381 gnd.n3380 9.3005
R12122 gnd.n3306 gnd.n3305 9.3005
R12123 gnd.n3375 gnd.n3374 9.3005
R12124 gnd.n3373 gnd.n3372 9.3005
R12125 gnd.n3317 gnd.n3316 9.3005
R12126 gnd.n3367 gnd.n3366 9.3005
R12127 gnd.n3365 gnd.n3364 9.3005
R12128 gnd.n3329 gnd.n3328 9.3005
R12129 gnd.n3359 gnd.n3358 9.3005
R12130 gnd.n3357 gnd.n3356 9.3005
R12131 gnd.n3342 gnd.n3341 9.3005
R12132 gnd.n3351 gnd.n3350 9.3005
R12133 gnd.n4889 gnd.n1328 9.3005
R12134 gnd.n4888 gnd.n4887 9.3005
R12135 gnd.n4886 gnd.n1332 9.3005
R12136 gnd.n4885 gnd.n4884 9.3005
R12137 gnd.n4883 gnd.n1333 9.3005
R12138 gnd.n4882 gnd.n4881 9.3005
R12139 gnd.n4880 gnd.n1337 9.3005
R12140 gnd.n4879 gnd.n4878 9.3005
R12141 gnd.n4877 gnd.n1338 9.3005
R12142 gnd.n4876 gnd.n4875 9.3005
R12143 gnd.n4874 gnd.n1342 9.3005
R12144 gnd.n4873 gnd.n4872 9.3005
R12145 gnd.n4871 gnd.n1343 9.3005
R12146 gnd.n4870 gnd.n4869 9.3005
R12147 gnd.n4868 gnd.n1347 9.3005
R12148 gnd.n4867 gnd.n4866 9.3005
R12149 gnd.n4865 gnd.n1348 9.3005
R12150 gnd.n4864 gnd.n4863 9.3005
R12151 gnd.n4862 gnd.n1352 9.3005
R12152 gnd.n4861 gnd.n4860 9.3005
R12153 gnd.n4859 gnd.n1353 9.3005
R12154 gnd.n4858 gnd.n4857 9.3005
R12155 gnd.n4856 gnd.n1357 9.3005
R12156 gnd.n4855 gnd.n4854 9.3005
R12157 gnd.n4853 gnd.n1358 9.3005
R12158 gnd.n4852 gnd.n4851 9.3005
R12159 gnd.n4850 gnd.n1362 9.3005
R12160 gnd.n4849 gnd.n4848 9.3005
R12161 gnd.n4847 gnd.n1363 9.3005
R12162 gnd.n4846 gnd.n4845 9.3005
R12163 gnd.n4844 gnd.n1367 9.3005
R12164 gnd.n4843 gnd.n4842 9.3005
R12165 gnd.n4841 gnd.n1368 9.3005
R12166 gnd.n4840 gnd.n4839 9.3005
R12167 gnd.n4838 gnd.n1372 9.3005
R12168 gnd.n4837 gnd.n4836 9.3005
R12169 gnd.n4835 gnd.n1373 9.3005
R12170 gnd.n4834 gnd.n4833 9.3005
R12171 gnd.n4832 gnd.n1377 9.3005
R12172 gnd.n4831 gnd.n4830 9.3005
R12173 gnd.n4829 gnd.n1378 9.3005
R12174 gnd.n4828 gnd.n4827 9.3005
R12175 gnd.n4826 gnd.n1382 9.3005
R12176 gnd.n4825 gnd.n4824 9.3005
R12177 gnd.n4823 gnd.n1383 9.3005
R12178 gnd.n4822 gnd.n4821 9.3005
R12179 gnd.n4820 gnd.n1387 9.3005
R12180 gnd.n4819 gnd.n4818 9.3005
R12181 gnd.n4817 gnd.n1388 9.3005
R12182 gnd.n4816 gnd.n4815 9.3005
R12183 gnd.n4814 gnd.n1392 9.3005
R12184 gnd.n4813 gnd.n4812 9.3005
R12185 gnd.n4811 gnd.n1393 9.3005
R12186 gnd.n4810 gnd.n4809 9.3005
R12187 gnd.n4808 gnd.n1397 9.3005
R12188 gnd.n4807 gnd.n4806 9.3005
R12189 gnd.n4805 gnd.n1398 9.3005
R12190 gnd.n4804 gnd.n4803 9.3005
R12191 gnd.n4802 gnd.n1402 9.3005
R12192 gnd.n4801 gnd.n4800 9.3005
R12193 gnd.n4799 gnd.n1403 9.3005
R12194 gnd.n4798 gnd.n4797 9.3005
R12195 gnd.n4796 gnd.n1407 9.3005
R12196 gnd.n4795 gnd.n4794 9.3005
R12197 gnd.n4793 gnd.n1408 9.3005
R12198 gnd.n4792 gnd.n4791 9.3005
R12199 gnd.n4790 gnd.n1412 9.3005
R12200 gnd.n4789 gnd.n4788 9.3005
R12201 gnd.n4787 gnd.n1413 9.3005
R12202 gnd.n4786 gnd.n4785 9.3005
R12203 gnd.n4784 gnd.n1417 9.3005
R12204 gnd.n4783 gnd.n4782 9.3005
R12205 gnd.n4781 gnd.n1418 9.3005
R12206 gnd.n4780 gnd.n4779 9.3005
R12207 gnd.n4778 gnd.n1422 9.3005
R12208 gnd.n4777 gnd.n4776 9.3005
R12209 gnd.n4775 gnd.n1423 9.3005
R12210 gnd.n4774 gnd.n4773 9.3005
R12211 gnd.n4772 gnd.n1427 9.3005
R12212 gnd.n4771 gnd.n4770 9.3005
R12213 gnd.n4769 gnd.n1428 9.3005
R12214 gnd.n4768 gnd.n4767 9.3005
R12215 gnd.n4766 gnd.n1432 9.3005
R12216 gnd.n4765 gnd.n4764 9.3005
R12217 gnd.n4763 gnd.n1433 9.3005
R12218 gnd.n4762 gnd.n4761 9.3005
R12219 gnd.n4760 gnd.n1437 9.3005
R12220 gnd.n4759 gnd.n4758 9.3005
R12221 gnd.n4757 gnd.n1438 9.3005
R12222 gnd.n4756 gnd.n4755 9.3005
R12223 gnd.n4754 gnd.n1442 9.3005
R12224 gnd.n4753 gnd.n4752 9.3005
R12225 gnd.n4751 gnd.n1443 9.3005
R12226 gnd.n4750 gnd.n4749 9.3005
R12227 gnd.n4748 gnd.n1447 9.3005
R12228 gnd.n4747 gnd.n4746 9.3005
R12229 gnd.n4745 gnd.n1448 9.3005
R12230 gnd.n4744 gnd.n4743 9.3005
R12231 gnd.n4742 gnd.n1452 9.3005
R12232 gnd.n4741 gnd.n4740 9.3005
R12233 gnd.n4739 gnd.n1453 9.3005
R12234 gnd.n4891 gnd.n4890 9.3005
R12235 gnd.n1689 gnd.n1685 9.3005
R12236 gnd.n1498 gnd.n1496 9.3005
R12237 gnd.n4713 gnd.n4712 9.3005
R12238 gnd.n4711 gnd.n1497 9.3005
R12239 gnd.n4710 gnd.n4709 9.3005
R12240 gnd.n4708 gnd.n1499 9.3005
R12241 gnd.n4707 gnd.n4706 9.3005
R12242 gnd.n4705 gnd.n1503 9.3005
R12243 gnd.n4704 gnd.n4703 9.3005
R12244 gnd.n4702 gnd.n1504 9.3005
R12245 gnd.n4701 gnd.n4700 9.3005
R12246 gnd.n4699 gnd.n1508 9.3005
R12247 gnd.n4698 gnd.n4697 9.3005
R12248 gnd.n4696 gnd.n1509 9.3005
R12249 gnd.n4695 gnd.n4694 9.3005
R12250 gnd.n4693 gnd.n1513 9.3005
R12251 gnd.n4692 gnd.n4691 9.3005
R12252 gnd.n4690 gnd.n1514 9.3005
R12253 gnd.n4689 gnd.n4688 9.3005
R12254 gnd.n4687 gnd.n4686 9.3005
R12255 gnd.n285 gnd.n283 9.3005
R12256 gnd.n7496 gnd.n7495 9.3005
R12257 gnd.n7494 gnd.n284 9.3005
R12258 gnd.n7493 gnd.n7492 9.3005
R12259 gnd.n7491 gnd.n286 9.3005
R12260 gnd.n7490 gnd.n7489 9.3005
R12261 gnd.n7487 gnd.n290 9.3005
R12262 gnd.n7486 gnd.n7485 9.3005
R12263 gnd.n7484 gnd.n292 9.3005
R12264 gnd.n261 gnd.n260 9.3005
R12265 gnd.n7508 gnd.n7507 9.3005
R12266 gnd.n7509 gnd.n259 9.3005
R12267 gnd.n7511 gnd.n7510 9.3005
R12268 gnd.n245 gnd.n244 9.3005
R12269 gnd.n7524 gnd.n7523 9.3005
R12270 gnd.n7525 gnd.n243 9.3005
R12271 gnd.n7527 gnd.n7526 9.3005
R12272 gnd.n230 gnd.n229 9.3005
R12273 gnd.n7540 gnd.n7539 9.3005
R12274 gnd.n7541 gnd.n228 9.3005
R12275 gnd.n7543 gnd.n7542 9.3005
R12276 gnd.n215 gnd.n214 9.3005
R12277 gnd.n7556 gnd.n7555 9.3005
R12278 gnd.n7557 gnd.n213 9.3005
R12279 gnd.n7559 gnd.n7558 9.3005
R12280 gnd.n200 gnd.n199 9.3005
R12281 gnd.n7572 gnd.n7571 9.3005
R12282 gnd.n7573 gnd.n197 9.3005
R12283 gnd.n7650 gnd.n7649 9.3005
R12284 gnd.n7648 gnd.n198 9.3005
R12285 gnd.n7647 gnd.n7646 9.3005
R12286 gnd.n7645 gnd.n7574 9.3005
R12287 gnd.n7644 gnd.n7643 9.3005
R12288 gnd.n1691 gnd.n1690 9.3005
R12289 gnd.n7640 gnd.n7576 9.3005
R12290 gnd.n7639 gnd.n7638 9.3005
R12291 gnd.n7637 gnd.n7581 9.3005
R12292 gnd.n7636 gnd.n7635 9.3005
R12293 gnd.n7634 gnd.n7582 9.3005
R12294 gnd.n7633 gnd.n7632 9.3005
R12295 gnd.n7631 gnd.n7589 9.3005
R12296 gnd.n7630 gnd.n7629 9.3005
R12297 gnd.n7628 gnd.n7590 9.3005
R12298 gnd.n7627 gnd.n7626 9.3005
R12299 gnd.n7625 gnd.n7597 9.3005
R12300 gnd.n7624 gnd.n7623 9.3005
R12301 gnd.n7622 gnd.n7598 9.3005
R12302 gnd.n7621 gnd.n7620 9.3005
R12303 gnd.n7619 gnd.n7605 9.3005
R12304 gnd.n7618 gnd.n7617 9.3005
R12305 gnd.n7616 gnd.n7606 9.3005
R12306 gnd.n7615 gnd.n7614 9.3005
R12307 gnd.n7642 gnd.n7641 9.3005
R12308 gnd.n4479 gnd.n1641 9.3005
R12309 gnd.n4482 gnd.n4481 9.3005
R12310 gnd.n4480 gnd.n1642 9.3005
R12311 gnd.n1622 gnd.n1621 9.3005
R12312 gnd.n4528 gnd.n4527 9.3005
R12313 gnd.n4529 gnd.n1619 9.3005
R12314 gnd.n4532 gnd.n4531 9.3005
R12315 gnd.n4530 gnd.n1620 9.3005
R12316 gnd.n1595 gnd.n1594 9.3005
R12317 gnd.n4560 gnd.n4559 9.3005
R12318 gnd.n4561 gnd.n1592 9.3005
R12319 gnd.n4564 gnd.n4563 9.3005
R12320 gnd.n4562 gnd.n1593 9.3005
R12321 gnd.n1566 gnd.n1565 9.3005
R12322 gnd.n4599 gnd.n4598 9.3005
R12323 gnd.n4600 gnd.n1563 9.3005
R12324 gnd.n4606 gnd.n4605 9.3005
R12325 gnd.n4604 gnd.n1564 9.3005
R12326 gnd.n4603 gnd.n4602 9.3005
R12327 gnd.n1555 gnd.n1554 9.3005
R12328 gnd.n4625 gnd.n4624 9.3005
R12329 gnd.n4626 gnd.n1552 9.3005
R12330 gnd.n4631 gnd.n4630 9.3005
R12331 gnd.n4629 gnd.n1553 9.3005
R12332 gnd.n4628 gnd.n4627 9.3005
R12333 gnd.n69 gnd.n67 9.3005
R12334 gnd.n7781 gnd.n7780 9.3005
R12335 gnd.n7779 gnd.n68 9.3005
R12336 gnd.n7778 gnd.n7777 9.3005
R12337 gnd.n7776 gnd.n73 9.3005
R12338 gnd.n7775 gnd.n7774 9.3005
R12339 gnd.n7773 gnd.n74 9.3005
R12340 gnd.n7772 gnd.n7771 9.3005
R12341 gnd.n7770 gnd.n78 9.3005
R12342 gnd.n7769 gnd.n7768 9.3005
R12343 gnd.n7767 gnd.n79 9.3005
R12344 gnd.n7766 gnd.n7765 9.3005
R12345 gnd.n7764 gnd.n83 9.3005
R12346 gnd.n7763 gnd.n7762 9.3005
R12347 gnd.n7761 gnd.n84 9.3005
R12348 gnd.n7760 gnd.n7759 9.3005
R12349 gnd.n7758 gnd.n88 9.3005
R12350 gnd.n7757 gnd.n7756 9.3005
R12351 gnd.n7755 gnd.n89 9.3005
R12352 gnd.n7754 gnd.n7753 9.3005
R12353 gnd.n7752 gnd.n93 9.3005
R12354 gnd.n7751 gnd.n7750 9.3005
R12355 gnd.n7749 gnd.n94 9.3005
R12356 gnd.n7748 gnd.n7747 9.3005
R12357 gnd.n7746 gnd.n98 9.3005
R12358 gnd.n7745 gnd.n7744 9.3005
R12359 gnd.n7743 gnd.n99 9.3005
R12360 gnd.n7742 gnd.n102 9.3005
R12361 gnd.n4478 gnd.n4477 9.3005
R12362 gnd.t147 gnd.n5259 9.24152
R12363 gnd.t183 gnd.n945 9.24152
R12364 gnd.n6394 gnd.t199 9.24152
R12365 gnd.t187 gnd.n1063 9.24152
R12366 gnd.n4903 gnd.t195 9.24152
R12367 gnd.n4484 gnd.t214 9.24152
R12368 gnd.n7660 gnd.t203 9.24152
R12369 gnd.t110 gnd.t147 8.92286
R12370 gnd.n3664 gnd.t254 8.92286
R12371 gnd.n2388 gnd.n2379 8.92286
R12372 gnd.t2 gnd.n2357 8.92286
R12373 gnd.n3797 gnd.n3795 8.92286
R12374 gnd.n3845 gnd.n2262 8.92286
R12375 gnd.n3951 gnd.n3950 8.92286
R12376 gnd.n4009 gnd.n2148 8.92286
R12377 gnd.t175 gnd.n2084 8.92286
R12378 gnd.n4183 gnd.n4182 8.92286
R12379 gnd.n4298 gnd.t241 8.92286
R12380 gnd.n6373 gnd.n6348 8.92171
R12381 gnd.n6341 gnd.n6316 8.92171
R12382 gnd.n6309 gnd.n6284 8.92171
R12383 gnd.n6278 gnd.n6253 8.92171
R12384 gnd.n6246 gnd.n6221 8.92171
R12385 gnd.n6214 gnd.n6189 8.92171
R12386 gnd.n6182 gnd.n6157 8.92171
R12387 gnd.n6151 gnd.n6126 8.92171
R12388 gnd.n4227 gnd.n4209 8.72777
R12389 gnd.t137 gnd.n5354 8.60421
R12390 gnd.n3412 gnd.t234 8.60421
R12391 gnd.n3451 gnd.t291 8.60421
R12392 gnd.n4397 gnd.t90 8.60421
R12393 gnd.n4449 gnd.t191 8.60421
R12394 gnd.n5322 gnd.n5306 8.43467
R12395 gnd.n50 gnd.n34 8.43467
R12396 gnd.n3132 gnd.n0 8.41456
R12397 gnd.n7783 gnd.n7782 8.41456
R12398 gnd.n2484 gnd.n2294 8.28555
R12399 gnd.n3872 gnd.n2232 8.28555
R12400 gnd.n3939 gnd.n2189 8.28555
R12401 gnd.n4033 gnd.n2140 8.28555
R12402 gnd.n6374 gnd.n6346 8.14595
R12403 gnd.n6342 gnd.n6314 8.14595
R12404 gnd.n6310 gnd.n6282 8.14595
R12405 gnd.n6279 gnd.n6251 8.14595
R12406 gnd.n6247 gnd.n6219 8.14595
R12407 gnd.n6215 gnd.n6187 8.14595
R12408 gnd.n6183 gnd.n6155 8.14595
R12409 gnd.n6152 gnd.n6124 8.14595
R12410 gnd.n6379 gnd.n6378 7.97301
R12411 gnd.n5847 gnd.t66 7.9669
R12412 gnd.n3397 gnd.n2775 7.9669
R12413 gnd.n1467 gnd.n1458 7.9669
R12414 gnd.n7616 gnd.n7615 7.75808
R12415 gnd.n4474 gnd.n1647 7.75808
R12416 gnd.n3350 gnd.n3341 7.75808
R12417 gnd.n2985 gnd.n2981 7.75808
R12418 gnd.n3655 gnd.n2393 7.64824
R12419 gnd.n2484 gnd.n2304 7.64824
R12420 gnd.t109 gnd.n2261 7.64824
R12421 gnd.n3851 gnd.t10 7.64824
R12422 gnd.n3872 gnd.n3871 7.64824
R12423 gnd.n2199 gnd.n2189 7.64824
R12424 gnd.t174 gnd.n3938 7.64824
R12425 gnd.n3949 gnd.t171 7.64824
R12426 gnd.n4033 gnd.n4032 7.64824
R12427 gnd.t88 gnd.n5440 7.32958
R12428 gnd.t234 gnd.n3411 7.32958
R12429 gnd.n3440 gnd.t291 7.32958
R12430 gnd.n3655 gnd.t153 7.32958
R12431 gnd.n4117 gnd.t39 7.32958
R12432 gnd.t90 gnd.n4396 7.32958
R12433 gnd.n4437 gnd.t191 7.32958
R12434 gnd.n2423 gnd.n2422 7.30353
R12435 gnd.n4226 gnd.n4225 7.30353
R12436 gnd.n5749 gnd.n5748 7.01093
R12437 gnd.n5759 gnd.n5469 7.01093
R12438 gnd.n5758 gnd.n5472 7.01093
R12439 gnd.n5767 gnd.n5463 7.01093
R12440 gnd.n5771 gnd.n5770 7.01093
R12441 gnd.n5789 gnd.n5448 7.01093
R12442 gnd.n5788 gnd.n5451 7.01093
R12443 gnd.n5799 gnd.n5440 7.01093
R12444 gnd.n5441 gnd.n5429 7.01093
R12445 gnd.n5812 gnd.n5430 7.01093
R12446 gnd.n5823 gnd.n5422 7.01093
R12447 gnd.n5822 gnd.n5413 7.01093
R12448 gnd.n5415 gnd.n5397 7.01093
R12449 gnd.n5859 gnd.n5398 7.01093
R12450 gnd.n5848 gnd.n5847 7.01093
R12451 gnd.n5884 gnd.n5389 7.01093
R12452 gnd.n5895 gnd.n5894 7.01093
R12453 gnd.n5382 gnd.n5374 7.01093
R12454 gnd.n5924 gnd.n5362 7.01093
R12455 gnd.n5923 gnd.n5365 7.01093
R12456 gnd.n5934 gnd.n5354 7.01093
R12457 gnd.n5355 gnd.n5343 7.01093
R12458 gnd.n5945 gnd.n5344 7.01093
R12459 gnd.n5969 gnd.n5287 7.01093
R12460 gnd.n5968 gnd.n5278 7.01093
R12461 gnd.n5280 gnd.n5271 7.01093
R12462 gnd.n5991 gnd.n5990 7.01093
R12463 gnd.n6008 gnd.n5259 7.01093
R12464 gnd.n6007 gnd.n5262 7.01093
R12465 gnd.n6021 gnd.n5251 7.01093
R12466 gnd.n5252 gnd.n5240 7.01093
R12467 gnd.n6031 gnd.n5242 7.01093
R12468 gnd.n6062 gnd.n6061 7.01093
R12469 gnd.n6075 gnd.n6074 7.01093
R12470 gnd.n5221 gnd.n5211 7.01093
R12471 gnd.n6087 gnd.n6086 7.01093
R12472 gnd.n6099 gnd.n909 7.01093
R12473 gnd.n6516 gnd.n920 7.01093
R12474 gnd.n6117 gnd.n6116 7.01093
R12475 gnd.n6510 gnd.n6509 7.01093
R12476 gnd.n5195 gnd.n931 7.01093
R12477 gnd.n6503 gnd.n942 7.01093
R12478 gnd.n6502 gnd.n945 7.01093
R12479 gnd.n6395 gnd.n6394 7.01093
R12480 gnd.n6496 gnd.n6495 7.01093
R12481 gnd.n966 gnd.n956 7.01093
R12482 gnd.n3675 gnd.n2379 7.01093
R12483 gnd.n3713 gnd.n3712 7.01093
R12484 gnd.n2509 gnd.t144 7.01093
R12485 gnd.n3795 gnd.n2290 7.01093
R12486 gnd.n3804 gnd.t109 7.01093
R12487 gnd.n3845 gnd.n2261 7.01093
R12488 gnd.n3950 gnd.n3949 7.01093
R12489 gnd.n3958 gnd.t171 7.01093
R12490 gnd.n4001 gnd.n2148 7.01093
R12491 gnd.n4110 gnd.t104 7.01093
R12492 gnd.n4141 gnd.n4140 7.01093
R12493 gnd.n4183 gnd.n2060 7.01093
R12494 gnd.n5430 gnd.t79 6.69227
R12495 gnd.n5990 gnd.t110 6.69227
R12496 gnd.n6517 gnd.t300 6.69227
R12497 gnd.n5030 gnd.t58 6.69227
R12498 gnd.n3723 gnd.t62 6.69227
R12499 gnd.n2110 gnd.t310 6.69227
R12500 gnd.t121 gnd.n208 6.69227
R12501 gnd.n4359 gnd.n4358 6.5566
R12502 gnd.n2598 gnd.n2597 6.5566
R12503 gnd.n3582 gnd.n2464 6.5566
R12504 gnd.n4237 gnd.n4236 6.5566
R12505 gnd.n3472 gnd.n2400 6.37362
R12506 gnd.t254 gnd.t244 6.37362
R12507 gnd.n3770 gnd.n2309 6.37362
R12508 gnd.n3826 gnd.t173 6.37362
R12509 gnd.n3863 gnd.n2218 6.37362
R12510 gnd.n3906 gnd.n2204 6.37362
R12511 gnd.t172 gnd.n2163 6.37362
R12512 gnd.n2136 gnd.n2125 6.37362
R12513 gnd.n4182 gnd.t180 6.37362
R12514 gnd.t180 gnd.n2053 6.37362
R12515 gnd.n4298 gnd.n2037 6.37362
R12516 gnd.n3510 gnd.n2718 6.20656
R12517 gnd.n7705 gnd.n7702 6.20656
R12518 gnd.n5099 gnd.n5098 6.20656
R12519 gnd.n4459 gnd.n1791 6.20656
R12520 gnd.n5883 gnd.t86 6.05496
R12521 gnd.n5882 gnd.t80 6.05496
R12522 gnd.t318 gnd.n5355 6.05496
R12523 gnd.t81 gnd.n5234 6.05496
R12524 gnd.n5024 gnd.n1108 6.05496
R12525 gnd.n5006 gnd.t21 6.05496
R12526 gnd.t166 gnd.t316 6.05496
R12527 gnd.t151 gnd.t298 6.05496
R12528 gnd.n7414 gnd.t23 6.05496
R12529 gnd.n7393 gnd.n218 6.05496
R12530 gnd.n6376 gnd.n6346 5.81868
R12531 gnd.n6344 gnd.n6314 5.81868
R12532 gnd.n6312 gnd.n6282 5.81868
R12533 gnd.n6281 gnd.n6251 5.81868
R12534 gnd.n6249 gnd.n6219 5.81868
R12535 gnd.n6217 gnd.n6187 5.81868
R12536 gnd.n6185 gnd.n6155 5.81868
R12537 gnd.n6154 gnd.n6124 5.81868
R12538 gnd.n3686 gnd.n3685 5.73631
R12539 gnd.n2519 gnd.n2518 5.73631
R12540 gnd.n3827 gnd.n2275 5.73631
R12541 gnd.n2469 gnd.n2468 5.73631
R12542 gnd.t10 gnd.n2232 5.73631
R12543 gnd.n3939 gnd.t174 5.73631
R12544 gnd.n3984 gnd.n3983 5.73631
R12545 gnd.n3991 gnd.n3990 5.73631
R12546 gnd.n4133 gnd.n4132 5.73631
R12547 gnd.n4158 gnd.n2068 5.73631
R12548 gnd.n4363 gnd.n2031 5.62001
R12549 gnd.n3577 gnd.n2602 5.62001
R12550 gnd.n3578 gnd.n3577 5.62001
R12551 gnd.n4232 gnd.n2031 5.62001
R12552 gnd.n5567 gnd.n5566 5.4308
R12553 gnd.n6409 gnd.n5186 5.4308
R12554 gnd.n5344 gnd.t65 5.41765
R12555 gnd.t103 gnd.n5979 5.41765
R12556 gnd.n6063 gnd.t149 5.41765
R12557 gnd.n4982 gnd.t53 5.41765
R12558 gnd.t330 gnd.n3757 5.41765
R12559 gnd.n4050 gnd.t125 5.41765
R12560 gnd.n7477 gnd.t27 5.41765
R12561 gnd.n3731 gnd.t64 5.09899
R12562 gnd.n3748 gnd.n3747 5.09899
R12563 gnd.n3888 gnd.n2211 5.09899
R12564 gnd.n3896 gnd.n2214 5.09899
R12565 gnd.n4065 gnd.n2116 5.09899
R12566 gnd.n4098 gnd.t9 5.09899
R12567 gnd.n6374 gnd.n6373 5.04292
R12568 gnd.n6342 gnd.n6341 5.04292
R12569 gnd.n6310 gnd.n6309 5.04292
R12570 gnd.n6279 gnd.n6278 5.04292
R12571 gnd.n6247 gnd.n6246 5.04292
R12572 gnd.n6215 gnd.n6214 5.04292
R12573 gnd.n6183 gnd.n6182 5.04292
R12574 gnd.n6152 gnd.n6151 5.04292
R12575 gnd.n5338 gnd.n5337 4.82753
R12576 gnd.n66 gnd.n65 4.82753
R12577 gnd.t313 gnd.n5905 4.78034
R12578 gnd.n6021 gnd.t312 4.78034
R12579 gnd.n4957 gnd.t94 4.78034
R12580 gnd.n3468 gnd.t0 4.78034
R12581 gnd.n4366 gnd.t231 4.78034
R12582 gnd.n1870 gnd.t5 4.78034
R12583 gnd.n4684 gnd.t118 4.78034
R12584 gnd.n5879 gnd.n5878 4.74817
R12585 gnd.n5874 gnd.n5873 4.74817
R12586 gnd.n5870 gnd.n5869 4.74817
R12587 gnd.n5866 gnd.n5341 4.74817
R12588 gnd.n5878 gnd.n5877 4.74817
R12589 gnd.n5876 gnd.n5874 4.74817
R12590 gnd.n5872 gnd.n5870 4.74817
R12591 gnd.n5868 gnd.n5866 4.74817
R12592 gnd.n7501 gnd.n7500 4.74817
R12593 gnd.n1547 gnd.n271 4.74817
R12594 gnd.n7479 gnd.n270 4.74817
R12595 gnd.n269 gnd.n266 4.74817
R12596 gnd.n7501 gnd.n273 4.74817
R12597 gnd.n4659 gnd.n271 4.74817
R12598 gnd.n1546 gnd.n270 4.74817
R12599 gnd.n7480 gnd.n269 4.74817
R12600 gnd.n2935 gnd.n2934 4.74817
R12601 gnd.n2931 gnd.n2881 4.74817
R12602 gnd.n2924 gnd.n2880 4.74817
R12603 gnd.n2920 gnd.n2879 4.74817
R12604 gnd.n2916 gnd.n2878 4.74817
R12605 gnd.n4666 gnd.n4665 4.74817
R12606 gnd.n4648 gnd.n1539 4.74817
R12607 gnd.n4653 gnd.n4652 4.74817
R12608 gnd.n4649 gnd.n308 4.74817
R12609 gnd.n7467 gnd.n7466 4.74817
R12610 gnd.n4667 gnd.n4666 4.74817
R12611 gnd.n4664 gnd.n1539 4.74817
R12612 gnd.n4654 gnd.n4653 4.74817
R12613 gnd.n4651 gnd.n4649 4.74817
R12614 gnd.n7468 gnd.n7467 4.74817
R12615 gnd.n1174 gnd.n1156 4.74817
R12616 gnd.n1192 gnd.n1176 4.74817
R12617 gnd.n4973 gnd.n4972 4.74817
R12618 gnd.n1211 gnd.n1193 4.74817
R12619 gnd.n4986 gnd.n1174 4.74817
R12620 gnd.n4984 gnd.n1176 4.74817
R12621 gnd.n4974 gnd.n4973 4.74817
R12622 gnd.n4971 gnd.n1193 4.74817
R12623 gnd.n2934 gnd.n2876 4.74817
R12624 gnd.n2931 gnd.n2930 4.74817
R12625 gnd.n2926 gnd.n2880 4.74817
R12626 gnd.n2923 gnd.n2879 4.74817
R12627 gnd.n2919 gnd.n2878 4.74817
R12628 gnd.n5322 gnd.n5321 4.7074
R12629 gnd.n50 gnd.n49 4.7074
R12630 gnd.n5338 gnd.n5322 4.65959
R12631 gnd.n66 gnd.n50 4.65959
R12632 gnd.n2030 gnd.n1947 4.6132
R12633 gnd.n3573 gnd.n3572 4.6132
R12634 gnd.n3688 gnd.n2370 4.46168
R12635 gnd.n3706 gnd.n3705 4.46168
R12636 gnd.n2476 gnd.t138 4.46168
R12637 gnd.n3820 gnd.n2281 4.46168
R12638 gnd.n3838 gnd.n3837 4.46168
R12639 gnd.n2183 gnd.n2182 4.46168
R12640 gnd.n3976 gnd.n3975 4.46168
R12641 gnd.t25 gnd.n2154 4.46168
R12642 gnd.n4148 gnd.n4147 4.46168
R12643 gnd.n4165 gnd.n2070 4.46168
R12644 gnd.t282 gnd.n2042 4.46168
R12645 gnd.n4222 gnd.n4209 4.46111
R12646 gnd.n6359 gnd.n6355 4.38594
R12647 gnd.n6327 gnd.n6323 4.38594
R12648 gnd.n6295 gnd.n6291 4.38594
R12649 gnd.n6264 gnd.n6260 4.38594
R12650 gnd.n6232 gnd.n6228 4.38594
R12651 gnd.n6200 gnd.n6196 4.38594
R12652 gnd.n6168 gnd.n6164 4.38594
R12653 gnd.n6137 gnd.n6133 4.38594
R12654 gnd.n6370 gnd.n6348 4.26717
R12655 gnd.n6338 gnd.n6316 4.26717
R12656 gnd.n6306 gnd.n6284 4.26717
R12657 gnd.n6275 gnd.n6253 4.26717
R12658 gnd.n6243 gnd.n6221 4.26717
R12659 gnd.n6211 gnd.n6189 4.26717
R12660 gnd.n6179 gnd.n6157 4.26717
R12661 gnd.n6148 gnd.n6126 4.26717
R12662 gnd.t301 gnd.n5836 4.14303
R12663 gnd.n6086 gnd.t136 4.14303
R12664 gnd.n3079 gnd.t45 4.14303
R12665 gnd.n4933 gnd.t76 4.14303
R12666 gnd.n3238 gnd.t51 4.14303
R12667 gnd.n1610 gnd.t127 4.14303
R12668 gnd.t131 gnd.n4567 4.14303
R12669 gnd.n7545 gnd.t35 4.14303
R12670 gnd.n6378 gnd.n6377 4.08274
R12671 gnd.n4358 gnd.n4357 4.05904
R12672 gnd.n2597 gnd.n2596 4.05904
R12673 gnd.n3585 gnd.n2464 4.05904
R12674 gnd.n4238 gnd.n4237 4.05904
R12675 gnd.n19 gnd.n9 3.99943
R12676 gnd.n3263 gnd.n2666 3.82437
R12677 gnd.n3645 gnd.n2403 3.82437
R12678 gnd.n2501 gnd.n2500 3.82437
R12679 gnd.n2492 gnd.t139 3.82437
R12680 gnd.n3768 gnd.n3767 3.82437
R12681 gnd.n3879 gnd.n3878 3.82437
R12682 gnd.n3862 gnd.t166 3.82437
R12683 gnd.n3905 gnd.t151 3.82437
R12684 gnd.n3915 gnd.n2197 3.82437
R12685 gnd.n4041 gnd.n4040 3.82437
R12686 gnd.n4067 gnd.t67 3.82437
R12687 gnd.n4089 gnd.n4088 3.82437
R12688 gnd.n2046 gnd.n2044 3.82437
R12689 gnd.n4728 gnd.n1468 3.82437
R12690 gnd.n6378 gnd.n6250 3.70378
R12691 gnd.n5340 gnd.n5339 3.65935
R12692 gnd.n19 gnd.n18 3.60163
R12693 gnd.n6524 gnd.n907 3.50571
R12694 gnd.n6524 gnd.n6523 3.50571
R12695 gnd.n2818 gnd.t98 3.50571
R12696 gnd.n3424 gnd.t29 3.50571
R12697 gnd.t287 gnd.n4415 3.50571
R12698 gnd.n4608 gnd.t3 3.50571
R12699 gnd.n6369 gnd.n6350 3.49141
R12700 gnd.n6337 gnd.n6318 3.49141
R12701 gnd.n6305 gnd.n6286 3.49141
R12702 gnd.n6274 gnd.n6255 3.49141
R12703 gnd.n6242 gnd.n6223 3.49141
R12704 gnd.n6210 gnd.n6191 3.49141
R12705 gnd.n6178 gnd.n6159 3.49141
R12706 gnd.n6147 gnd.n6128 3.49141
R12707 gnd.n3663 gnd.n3662 3.18706
R12708 gnd.n3685 gnd.t248 3.18706
R12709 gnd.n2511 gnd.n2510 3.18706
R12710 gnd.n3740 gnd.t26 3.18706
R12711 gnd.t26 gnd.n3739 3.18706
R12712 gnd.n3787 gnd.n2296 3.18706
R12713 gnd.n3853 gnd.n2256 3.18706
R12714 gnd.n3952 gnd.n2178 3.18706
R12715 gnd.n4008 gnd.n2150 3.18706
R12716 gnd.t152 gnd.n2118 3.18706
R12717 gnd.n4059 gnd.t152 3.18706
R12718 gnd.n4111 gnd.n2091 3.18706
R12719 gnd.n4191 gnd.n2053 3.18706
R12720 gnd.n4117 gnd.t282 3.18706
R12721 gnd.n5837 gnd.t301 2.8684
R12722 gnd.n2832 gnd.t15 2.8684
R12723 gnd.n3694 gnd.t84 2.8684
R12724 gnd.n4159 gnd.t7 2.8684
R12725 gnd.t60 gnd.n1544 2.8684
R12726 gnd.n5323 gnd.t170 2.82907
R12727 gnd.n5323 gnd.t290 2.82907
R12728 gnd.n5325 gnd.t129 2.82907
R12729 gnd.n5325 gnd.t297 2.82907
R12730 gnd.n5327 gnd.t133 2.82907
R12731 gnd.n5327 gnd.t116 2.82907
R12732 gnd.n5329 gnd.t322 2.82907
R12733 gnd.n5329 gnd.t165 2.82907
R12734 gnd.n5331 gnd.t32 2.82907
R12735 gnd.n5331 gnd.t78 2.82907
R12736 gnd.n5333 gnd.t135 2.82907
R12737 gnd.n5333 gnd.t130 2.82907
R12738 gnd.n5335 gnd.t164 2.82907
R12739 gnd.n5335 gnd.t305 2.82907
R12740 gnd.n5292 gnd.t92 2.82907
R12741 gnd.n5292 gnd.t52 2.82907
R12742 gnd.n5294 gnd.t99 2.82907
R12743 gnd.n5294 gnd.t34 2.82907
R12744 gnd.n5296 gnd.t115 2.82907
R12745 gnd.n5296 gnd.t95 2.82907
R12746 gnd.n5298 gnd.t54 2.82907
R12747 gnd.n5298 gnd.t142 2.82907
R12748 gnd.n5300 gnd.t93 2.82907
R12749 gnd.n5300 gnd.t48 2.82907
R12750 gnd.n5302 gnd.t167 2.82907
R12751 gnd.n5302 gnd.t100 2.82907
R12752 gnd.n5304 gnd.t124 2.82907
R12753 gnd.n5304 gnd.t120 2.82907
R12754 gnd.n5307 gnd.t77 2.82907
R12755 gnd.n5307 gnd.t155 2.82907
R12756 gnd.n5309 gnd.t176 2.82907
R12757 gnd.n5309 gnd.t140 2.82907
R12758 gnd.n5311 gnd.t123 2.82907
R12759 gnd.n5311 gnd.t113 2.82907
R12760 gnd.n5313 gnd.t156 2.82907
R12761 gnd.n5313 gnd.t16 2.82907
R12762 gnd.n5315 gnd.t162 2.82907
R12763 gnd.n5315 gnd.t320 2.82907
R12764 gnd.n5317 gnd.t14 2.82907
R12765 gnd.n5317 gnd.t22 2.82907
R12766 gnd.n5319 gnd.t59 2.82907
R12767 gnd.n5319 gnd.t46 2.82907
R12768 gnd.n63 gnd.t36 2.82907
R12769 gnd.n63 gnd.t122 2.82907
R12770 gnd.n61 gnd.t326 2.82907
R12771 gnd.n61 gnd.t296 2.82907
R12772 gnd.n59 gnd.t321 2.82907
R12773 gnd.n59 gnd.t289 2.82907
R12774 gnd.n57 gnd.t295 2.82907
R12775 gnd.n57 gnd.t143 2.82907
R12776 gnd.n55 gnd.t163 2.82907
R12777 gnd.n55 gnd.t327 2.82907
R12778 gnd.n53 gnd.t315 2.82907
R12779 gnd.n53 gnd.t325 2.82907
R12780 gnd.n51 gnd.t329 2.82907
R12781 gnd.n51 gnd.t132 2.82907
R12782 gnd.n32 gnd.t146 2.82907
R12783 gnd.n32 gnd.t304 2.82907
R12784 gnd.n30 gnd.t24 2.82907
R12785 gnd.n30 gnd.t101 2.82907
R12786 gnd.n28 gnd.t159 2.82907
R12787 gnd.n28 gnd.t12 2.82907
R12788 gnd.n26 gnd.t61 2.82907
R12789 gnd.n26 gnd.t28 2.82907
R12790 gnd.n24 gnd.t314 2.82907
R12791 gnd.n24 gnd.t112 2.82907
R12792 gnd.n22 gnd.t177 2.82907
R12793 gnd.n22 gnd.t4 2.82907
R12794 gnd.n20 gnd.t178 2.82907
R12795 gnd.n20 gnd.t134 2.82907
R12796 gnd.n47 gnd.t158 2.82907
R12797 gnd.n47 gnd.t303 2.82907
R12798 gnd.n45 gnd.t41 2.82907
R12799 gnd.n45 gnd.t43 2.82907
R12800 gnd.n43 gnd.t50 2.82907
R12801 gnd.n43 gnd.t44 2.82907
R12802 gnd.n41 gnd.t161 2.82907
R12803 gnd.n41 gnd.t55 2.82907
R12804 gnd.n39 gnd.t119 2.82907
R12805 gnd.n39 gnd.t75 2.82907
R12806 gnd.n37 gnd.t57 2.82907
R12807 gnd.n37 gnd.t302 2.82907
R12808 gnd.n35 gnd.t128 2.82907
R12809 gnd.n35 gnd.t157 2.82907
R12810 gnd.n6366 gnd.n6365 2.71565
R12811 gnd.n6334 gnd.n6333 2.71565
R12812 gnd.n6302 gnd.n6301 2.71565
R12813 gnd.n6271 gnd.n6270 2.71565
R12814 gnd.n6239 gnd.n6238 2.71565
R12815 gnd.n6207 gnd.n6206 2.71565
R12816 gnd.n6175 gnd.n6174 2.71565
R12817 gnd.n6144 gnd.n6143 2.71565
R12818 gnd.n5018 gnd.n1116 2.54975
R12819 gnd.n3087 gnd.n1119 2.54975
R12820 gnd.n5012 gnd.n1127 2.54975
R12821 gnd.n3095 gnd.n1130 2.54975
R12822 gnd.n5006 gnd.n1138 2.54975
R12823 gnd.n3103 gnd.n2943 2.54975
R12824 gnd.n5000 gnd.n1148 2.54975
R12825 gnd.n3111 gnd.n2847 2.54975
R12826 gnd.n4994 gnd.n1158 2.54975
R12827 gnd.n3119 gnd.n1161 2.54975
R12828 gnd.n4988 gnd.n1169 2.54975
R12829 gnd.n3127 gnd.n1172 2.54975
R12830 gnd.n4982 gnd.n1178 2.54975
R12831 gnd.n3136 gnd.n2837 2.54975
R12832 gnd.n4976 gnd.n1188 2.54975
R12833 gnd.n3145 gnd.n2832 2.54975
R12834 gnd.n4969 gnd.n1195 2.54975
R12835 gnd.n3153 gnd.n1198 2.54975
R12836 gnd.n4963 gnd.n1206 2.54975
R12837 gnd.n3161 gnd.n1209 2.54975
R12838 gnd.n4957 gnd.n1216 2.54975
R12839 gnd.n3169 gnd.n2822 2.54975
R12840 gnd.n4951 gnd.n1226 2.54975
R12841 gnd.n3177 gnd.n2818 2.54975
R12842 gnd.n4945 gnd.n1236 2.54975
R12843 gnd.n3185 gnd.n1239 2.54975
R12844 gnd.n4939 gnd.n1247 2.54975
R12845 gnd.n3194 gnd.n1250 2.54975
R12846 gnd.n4933 gnd.n1258 2.54975
R12847 gnd.n3202 gnd.n2808 2.54975
R12848 gnd.n4927 gnd.n1268 2.54975
R12849 gnd.n3238 gnd.n3237 2.54975
R12850 gnd.n4921 gnd.n1278 2.54975
R12851 gnd.n3210 gnd.n1281 2.54975
R12852 gnd.n4915 gnd.n1289 2.54975
R12853 gnd.n3214 gnd.n1292 2.54975
R12854 gnd.n4909 gnd.n1300 2.54975
R12855 gnd.n3223 gnd.n1303 2.54975
R12856 gnd.n4903 gnd.n1311 2.54975
R12857 gnd.n3528 gnd.n2701 2.54975
R12858 gnd.n4897 gnd.n1320 2.54975
R12859 gnd.n3664 gnd.n2386 2.54975
R12860 gnd.n3724 gnd.n2344 2.54975
R12861 gnd.n2505 gnd.t64 2.54975
R12862 gnd.n3789 gnd.n3788 2.54975
R12863 gnd.n3788 gnd.t68 2.54975
R12864 gnd.n3852 gnd.n3851 2.54975
R12865 gnd.n3938 gnd.n3937 2.54975
R12866 gnd.n3967 gnd.t69 2.54975
R12867 gnd.n3968 gnd.n3967 2.54975
R12868 gnd.t9 gnd.n4096 2.54975
R12869 gnd.n2109 gnd.n2108 2.54975
R12870 gnd.n4190 gnd.n4189 2.54975
R12871 gnd.n4722 gnd.n1477 2.54975
R12872 gnd.n4721 gnd.n1480 2.54975
R12873 gnd.n4484 gnd.n1490 2.54975
R12874 gnd.n4715 gnd.n1493 2.54975
R12875 gnd.n1635 gnd.n1634 2.54975
R12876 gnd.n4525 gnd.n4517 2.54975
R12877 gnd.n4535 gnd.n1616 2.54975
R12878 gnd.n4534 gnd.n1605 2.54975
R12879 gnd.n4547 gnd.n4545 2.54975
R12880 gnd.n1610 gnd.n1608 2.54975
R12881 gnd.n4557 gnd.n1598 2.54975
R12882 gnd.n4568 gnd.n1589 2.54975
R12883 gnd.n4567 gnd.n1578 2.54975
R12884 gnd.n4586 gnd.n4585 2.54975
R12885 gnd.n1583 gnd.n1581 2.54975
R12886 gnd.n4596 gnd.n1569 2.54975
R12887 gnd.n1572 gnd.n1561 2.54975
R12888 gnd.n4609 gnd.n4608 2.54975
R12889 gnd.n4676 gnd.n4675 2.54975
R12890 gnd.n1530 gnd.n1528 2.54975
R12891 gnd.n4684 gnd.n1520 2.54975
R12892 gnd.n4622 gnd.n277 2.54975
R12893 gnd.n7498 gnd.n280 2.54975
R12894 gnd.n4634 gnd.n4633 2.54975
R12895 gnd.n4662 gnd.n1541 2.54975
R12896 gnd.n4661 gnd.n1544 2.54975
R12897 gnd.n4657 gnd.n4656 2.54975
R12898 gnd.n4646 gnd.n4645 2.54975
R12899 gnd.n7477 gnd.n294 2.54975
R12900 gnd.n7482 gnd.n296 2.54975
R12901 gnd.n7471 gnd.n7470 2.54975
R12902 gnd.n7505 gnd.n264 2.54975
R12903 gnd.n7403 gnd.n255 2.54975
R12904 gnd.n7513 gnd.n257 2.54975
R12905 gnd.n7410 gnd.n247 2.54975
R12906 gnd.n7521 gnd.n249 2.54975
R12907 gnd.n7414 gnd.n239 2.54975
R12908 gnd.n7529 gnd.n241 2.54975
R12909 gnd.n7455 gnd.n7454 2.54975
R12910 gnd.n7537 gnd.n233 2.54975
R12911 gnd.n7447 gnd.n225 2.54975
R12912 gnd.n5878 gnd.n5340 2.27742
R12913 gnd.n5874 gnd.n5340 2.27742
R12914 gnd.n5870 gnd.n5340 2.27742
R12915 gnd.n5866 gnd.n5340 2.27742
R12916 gnd.n7502 gnd.n7501 2.27742
R12917 gnd.n7502 gnd.n271 2.27742
R12918 gnd.n7502 gnd.n270 2.27742
R12919 gnd.n7502 gnd.n269 2.27742
R12920 gnd.n4666 gnd.n268 2.27742
R12921 gnd.n1539 gnd.n268 2.27742
R12922 gnd.n4653 gnd.n268 2.27742
R12923 gnd.n4649 gnd.n268 2.27742
R12924 gnd.n7467 gnd.n268 2.27742
R12925 gnd.n1175 gnd.n1174 2.27742
R12926 gnd.n1176 gnd.n1175 2.27742
R12927 gnd.n4973 gnd.n1175 2.27742
R12928 gnd.n1193 gnd.n1175 2.27742
R12929 gnd.n2934 gnd.n2933 2.27742
R12930 gnd.n2933 gnd.n2931 2.27742
R12931 gnd.n2933 gnd.n2880 2.27742
R12932 gnd.n2933 gnd.n2879 2.27742
R12933 gnd.n2933 gnd.n2878 2.27742
R12934 gnd.t266 gnd.n5758 2.23109
R12935 gnd.n5906 gnd.t313 2.23109
R12936 gnd.n2847 gnd.t31 2.23109
R12937 gnd.n3837 gnd.t293 2.23109
R12938 gnd.n3878 gnd.t316 2.23109
R12939 gnd.t298 gnd.n2197 2.23109
R12940 gnd.n2183 gnd.t323 2.23109
R12941 gnd.t11 gnd.n257 2.23109
R12942 gnd.n6362 gnd.n6352 1.93989
R12943 gnd.n6330 gnd.n6320 1.93989
R12944 gnd.n6298 gnd.n6288 1.93989
R12945 gnd.n6267 gnd.n6257 1.93989
R12946 gnd.n6235 gnd.n6225 1.93989
R12947 gnd.n6203 gnd.n6193 1.93989
R12948 gnd.n6171 gnd.n6161 1.93989
R12949 gnd.n6140 gnd.n6130 1.93989
R12950 gnd.n2533 gnd.n2532 1.91244
R12951 gnd.n2533 gnd.t218 1.91244
R12952 gnd.n3712 gnd.t144 1.91244
R12953 gnd.n3730 gnd.n2340 1.91244
R12954 gnd.n3777 gnd.n3776 1.91244
R12955 gnd.n3869 gnd.n2227 1.91244
R12956 gnd.n3914 gnd.n3913 1.91244
R12957 gnd.n4042 gnd.n2131 1.91244
R12958 gnd.n4087 gnd.n2099 1.91244
R12959 gnd.n4141 gnd.t104 1.91244
R12960 gnd.n4205 gnd.n4204 1.91244
R12961 gnd.n5771 gnd.t306 1.59378
R12962 gnd.n5980 gnd.t103 1.59378
R12963 gnd.n6051 gnd.t149 1.59378
R12964 gnd.n2505 gnd.t62 1.59378
R12965 gnd.n3797 gnd.t308 1.59378
R12966 gnd.n4009 gnd.t37 1.59378
R12967 gnd.n4096 gnd.t310 1.59378
R12968 gnd.n3472 gnd.t263 1.27512
R12969 gnd.n3674 gnd.n3673 1.27512
R12970 gnd.n2519 gnd.t2 1.27512
R12971 gnd.n3704 gnd.n2352 1.27512
R12972 gnd.n3758 gnd.t139 1.27512
R12973 gnd.n2477 gnd.n2476 1.27512
R12974 gnd.n3805 gnd.n3804 1.27512
R12975 gnd.n3958 gnd.n2174 1.27512
R12976 gnd.n4002 gnd.n2154 1.27512
R12977 gnd.n4017 gnd.t67 1.27512
R12978 gnd.n4139 gnd.n2081 1.27512
R12979 gnd.n4133 gnd.t175 1.27512
R12980 gnd.t207 gnd.n2070 1.27512
R12981 gnd.n4125 gnd.n4124 1.27512
R12982 gnd.n5568 gnd.n5567 1.16414
R12983 gnd.n6412 gnd.n5186 1.16414
R12984 gnd.n6361 gnd.n6354 1.16414
R12985 gnd.n6329 gnd.n6322 1.16414
R12986 gnd.n6297 gnd.n6290 1.16414
R12987 gnd.n6266 gnd.n6259 1.16414
R12988 gnd.n6234 gnd.n6227 1.16414
R12989 gnd.n6202 gnd.n6195 1.16414
R12990 gnd.n6170 gnd.n6163 1.16414
R12991 gnd.n6139 gnd.n6132 1.16414
R12992 gnd.n2030 gnd.n2029 0.970197
R12993 gnd.n3573 gnd.n2603 0.970197
R12994 gnd.n6345 gnd.n6313 0.962709
R12995 gnd.n6377 gnd.n6345 0.962709
R12996 gnd.n6218 gnd.n6186 0.962709
R12997 gnd.n6250 gnd.n6218 0.962709
R12998 gnd.t86 gnd.n5882 0.956468
R12999 gnd.n5241 gnd.t81 0.956468
R13000 gnd.n3637 gnd.n2460 0.956468
R13001 gnd.t153 gnd.n3654 0.956468
R13002 gnd.t39 gnd.n2056 0.956468
R13003 gnd.n4367 gnd.n4366 0.956468
R13004 gnd.n5332 gnd.n5330 0.773756
R13005 gnd.n60 gnd.n58 0.773756
R13006 gnd.n5337 gnd.n5336 0.773756
R13007 gnd.n5336 gnd.n5334 0.773756
R13008 gnd.n5334 gnd.n5332 0.773756
R13009 gnd.n5330 gnd.n5328 0.773756
R13010 gnd.n5328 gnd.n5326 0.773756
R13011 gnd.n5326 gnd.n5324 0.773756
R13012 gnd.n54 gnd.n52 0.773756
R13013 gnd.n56 gnd.n54 0.773756
R13014 gnd.n58 gnd.n56 0.773756
R13015 gnd.n62 gnd.n60 0.773756
R13016 gnd.n64 gnd.n62 0.773756
R13017 gnd.n65 gnd.n64 0.773756
R13018 gnd.n2 gnd.n1 0.672012
R13019 gnd.n3 gnd.n2 0.672012
R13020 gnd.n4 gnd.n3 0.672012
R13021 gnd.n5 gnd.n4 0.672012
R13022 gnd.n6 gnd.n5 0.672012
R13023 gnd.n7 gnd.n6 0.672012
R13024 gnd.n8 gnd.n7 0.672012
R13025 gnd.n9 gnd.n8 0.672012
R13026 gnd.n11 gnd.n10 0.672012
R13027 gnd.n12 gnd.n11 0.672012
R13028 gnd.n13 gnd.n12 0.672012
R13029 gnd.n14 gnd.n13 0.672012
R13030 gnd.n15 gnd.n14 0.672012
R13031 gnd.n16 gnd.n15 0.672012
R13032 gnd.n17 gnd.n16 0.672012
R13033 gnd.n18 gnd.n17 0.672012
R13034 gnd gnd.n0 0.665707
R13035 gnd.t244 gnd.n3663 0.637812
R13036 gnd.t238 gnd.n3674 0.637812
R13037 gnd.n3749 gnd.n2325 0.637812
R13038 gnd.n3757 gnd.n2319 0.637812
R13039 gnd.n3767 gnd.t107 0.637812
R13040 gnd.n3890 gnd.n3889 0.637812
R13041 gnd.n2244 gnd.n2243 0.637812
R13042 gnd.t108 gnd.n4041 0.637812
R13043 gnd.n4051 gnd.n4050 0.637812
R13044 gnd.n4074 gnd.n4073 0.637812
R13045 gnd.n4191 gnd.t210 0.637812
R13046 gnd.n2047 gnd.t241 0.637812
R13047 gnd.n5306 gnd.n5305 0.573776
R13048 gnd.n5305 gnd.n5303 0.573776
R13049 gnd.n5303 gnd.n5301 0.573776
R13050 gnd.n5301 gnd.n5299 0.573776
R13051 gnd.n5299 gnd.n5297 0.573776
R13052 gnd.n5297 gnd.n5295 0.573776
R13053 gnd.n5295 gnd.n5293 0.573776
R13054 gnd.n5321 gnd.n5320 0.573776
R13055 gnd.n5320 gnd.n5318 0.573776
R13056 gnd.n5318 gnd.n5316 0.573776
R13057 gnd.n5316 gnd.n5314 0.573776
R13058 gnd.n5314 gnd.n5312 0.573776
R13059 gnd.n5312 gnd.n5310 0.573776
R13060 gnd.n5310 gnd.n5308 0.573776
R13061 gnd.n23 gnd.n21 0.573776
R13062 gnd.n25 gnd.n23 0.573776
R13063 gnd.n27 gnd.n25 0.573776
R13064 gnd.n29 gnd.n27 0.573776
R13065 gnd.n31 gnd.n29 0.573776
R13066 gnd.n33 gnd.n31 0.573776
R13067 gnd.n34 gnd.n33 0.573776
R13068 gnd.n38 gnd.n36 0.573776
R13069 gnd.n40 gnd.n38 0.573776
R13070 gnd.n42 gnd.n40 0.573776
R13071 gnd.n44 gnd.n42 0.573776
R13072 gnd.n46 gnd.n44 0.573776
R13073 gnd.n48 gnd.n46 0.573776
R13074 gnd.n49 gnd.n48 0.573776
R13075 gnd.n7784 gnd.n7783 0.553847
R13076 gnd.n7502 gnd.n268 0.548625
R13077 gnd.n2933 gnd.n1175 0.548625
R13078 gnd.n2986 gnd.n2984 0.505073
R13079 gnd.n3024 gnd.n3023 0.505073
R13080 gnd.n7643 gnd.n7642 0.505073
R13081 gnd.n7614 gnd.n102 0.505073
R13082 gnd.n7737 gnd.n7736 0.492878
R13083 gnd.n7666 gnd.n7665 0.492878
R13084 gnd.n1988 gnd.n1982 0.492878
R13085 gnd.n1907 gnd.n1906 0.492878
R13086 gnd.n2624 gnd.n1318 0.492878
R13087 gnd.n3533 gnd.n3532 0.492878
R13088 gnd.n5059 gnd.n1056 0.492878
R13089 gnd.n3033 gnd.n1013 0.492878
R13090 gnd.n6400 gnd.n5190 0.486781
R13091 gnd.n1693 gnd.n1453 0.486781
R13092 gnd.n5620 gnd.n5516 0.48678
R13093 gnd.n4892 gnd.n4891 0.485256
R13094 gnd.n6491 gnd.n6490 0.480683
R13095 gnd.n5688 gnd.n5466 0.480683
R13096 gnd.n4455 gnd.n4454 0.451719
R13097 gnd.n3506 gnd.n3505 0.451719
R13098 gnd.n742 gnd.n737 0.447146
R13099 gnd.n7180 gnd.n7179 0.447146
R13100 gnd.n7391 gnd.n321 0.447146
R13101 gnd.n2862 gnd.n2861 0.447146
R13102 gnd.n4894 gnd.n4893 0.406268
R13103 gnd.n1692 gnd.n1691 0.404992
R13104 gnd.n3513 gnd.n2718 0.388379
R13105 gnd.n6358 gnd.n6357 0.388379
R13106 gnd.n6326 gnd.n6325 0.388379
R13107 gnd.n6294 gnd.n6293 0.388379
R13108 gnd.n6263 gnd.n6262 0.388379
R13109 gnd.n6231 gnd.n6230 0.388379
R13110 gnd.n6199 gnd.n6198 0.388379
R13111 gnd.n6167 gnd.n6166 0.388379
R13112 gnd.n6136 gnd.n6135 0.388379
R13113 gnd.n7706 gnd.n7705 0.388379
R13114 gnd.n5100 gnd.n5099 0.388379
R13115 gnd.n1791 gnd.n1787 0.388379
R13116 gnd.n7784 gnd.n19 0.374463
R13117 gnd gnd.n7784 0.367492
R13118 gnd.n6100 gnd.t300 0.319156
R13119 gnd.n5614 gnd.n5613 0.311721
R13120 gnd.n3524 gnd.n3523 0.27489
R13121 gnd.n4478 gnd.n1643 0.27489
R13122 gnd.n6457 gnd.n6456 0.268793
R13123 gnd.n6456 gnd.n6455 0.241354
R13124 gnd.n1947 gnd.n1946 0.229039
R13125 gnd.n1950 gnd.n1947 0.229039
R13126 gnd.n3572 gnd.n2608 0.229039
R13127 gnd.n3572 gnd.n3571 0.229039
R13128 gnd.n5743 gnd.n5484 0.206293
R13129 gnd.n5339 gnd.n0 0.169152
R13130 gnd.n6375 gnd.n6347 0.155672
R13131 gnd.n6368 gnd.n6347 0.155672
R13132 gnd.n6368 gnd.n6367 0.155672
R13133 gnd.n6367 gnd.n6351 0.155672
R13134 gnd.n6360 gnd.n6351 0.155672
R13135 gnd.n6360 gnd.n6359 0.155672
R13136 gnd.n6343 gnd.n6315 0.155672
R13137 gnd.n6336 gnd.n6315 0.155672
R13138 gnd.n6336 gnd.n6335 0.155672
R13139 gnd.n6335 gnd.n6319 0.155672
R13140 gnd.n6328 gnd.n6319 0.155672
R13141 gnd.n6328 gnd.n6327 0.155672
R13142 gnd.n6311 gnd.n6283 0.155672
R13143 gnd.n6304 gnd.n6283 0.155672
R13144 gnd.n6304 gnd.n6303 0.155672
R13145 gnd.n6303 gnd.n6287 0.155672
R13146 gnd.n6296 gnd.n6287 0.155672
R13147 gnd.n6296 gnd.n6295 0.155672
R13148 gnd.n6280 gnd.n6252 0.155672
R13149 gnd.n6273 gnd.n6252 0.155672
R13150 gnd.n6273 gnd.n6272 0.155672
R13151 gnd.n6272 gnd.n6256 0.155672
R13152 gnd.n6265 gnd.n6256 0.155672
R13153 gnd.n6265 gnd.n6264 0.155672
R13154 gnd.n6248 gnd.n6220 0.155672
R13155 gnd.n6241 gnd.n6220 0.155672
R13156 gnd.n6241 gnd.n6240 0.155672
R13157 gnd.n6240 gnd.n6224 0.155672
R13158 gnd.n6233 gnd.n6224 0.155672
R13159 gnd.n6233 gnd.n6232 0.155672
R13160 gnd.n6216 gnd.n6188 0.155672
R13161 gnd.n6209 gnd.n6188 0.155672
R13162 gnd.n6209 gnd.n6208 0.155672
R13163 gnd.n6208 gnd.n6192 0.155672
R13164 gnd.n6201 gnd.n6192 0.155672
R13165 gnd.n6201 gnd.n6200 0.155672
R13166 gnd.n6184 gnd.n6156 0.155672
R13167 gnd.n6177 gnd.n6156 0.155672
R13168 gnd.n6177 gnd.n6176 0.155672
R13169 gnd.n6176 gnd.n6160 0.155672
R13170 gnd.n6169 gnd.n6160 0.155672
R13171 gnd.n6169 gnd.n6168 0.155672
R13172 gnd.n6153 gnd.n6125 0.155672
R13173 gnd.n6146 gnd.n6125 0.155672
R13174 gnd.n6146 gnd.n6145 0.155672
R13175 gnd.n6145 gnd.n6129 0.155672
R13176 gnd.n6138 gnd.n6129 0.155672
R13177 gnd.n6138 gnd.n6137 0.155672
R13178 gnd.n6490 gnd.n963 0.152939
R13179 gnd.n5144 gnd.n963 0.152939
R13180 gnd.n5145 gnd.n5144 0.152939
R13181 gnd.n5146 gnd.n5145 0.152939
R13182 gnd.n5147 gnd.n5146 0.152939
R13183 gnd.n5148 gnd.n5147 0.152939
R13184 gnd.n5149 gnd.n5148 0.152939
R13185 gnd.n5150 gnd.n5149 0.152939
R13186 gnd.n5151 gnd.n5150 0.152939
R13187 gnd.n5152 gnd.n5151 0.152939
R13188 gnd.n5153 gnd.n5152 0.152939
R13189 gnd.n5154 gnd.n5153 0.152939
R13190 gnd.n5155 gnd.n5154 0.152939
R13191 gnd.n5156 gnd.n5155 0.152939
R13192 gnd.n6458 gnd.n5156 0.152939
R13193 gnd.n6458 gnd.n6457 0.152939
R13194 gnd.n5762 gnd.n5466 0.152939
R13195 gnd.n5763 gnd.n5762 0.152939
R13196 gnd.n5764 gnd.n5763 0.152939
R13197 gnd.n5764 gnd.n5445 0.152939
R13198 gnd.n5792 gnd.n5445 0.152939
R13199 gnd.n5793 gnd.n5792 0.152939
R13200 gnd.n5794 gnd.n5793 0.152939
R13201 gnd.n5795 gnd.n5794 0.152939
R13202 gnd.n5795 gnd.n5419 0.152939
R13203 gnd.n5826 gnd.n5419 0.152939
R13204 gnd.n5827 gnd.n5826 0.152939
R13205 gnd.n5828 gnd.n5827 0.152939
R13206 gnd.n5829 gnd.n5828 0.152939
R13207 gnd.n5830 gnd.n5829 0.152939
R13208 gnd.n5830 gnd.n5386 0.152939
R13209 gnd.n5887 gnd.n5386 0.152939
R13210 gnd.n5888 gnd.n5887 0.152939
R13211 gnd.n5889 gnd.n5888 0.152939
R13212 gnd.n5890 gnd.n5889 0.152939
R13213 gnd.n5890 gnd.n5359 0.152939
R13214 gnd.n5927 gnd.n5359 0.152939
R13215 gnd.n5928 gnd.n5927 0.152939
R13216 gnd.n5929 gnd.n5928 0.152939
R13217 gnd.n5930 gnd.n5929 0.152939
R13218 gnd.n5930 gnd.n5284 0.152939
R13219 gnd.n5972 gnd.n5284 0.152939
R13220 gnd.n5973 gnd.n5972 0.152939
R13221 gnd.n5974 gnd.n5973 0.152939
R13222 gnd.n5975 gnd.n5974 0.152939
R13223 gnd.n5975 gnd.n5256 0.152939
R13224 gnd.n6011 gnd.n5256 0.152939
R13225 gnd.n6012 gnd.n6011 0.152939
R13226 gnd.n6013 gnd.n6012 0.152939
R13227 gnd.n6014 gnd.n6013 0.152939
R13228 gnd.n6015 gnd.n6014 0.152939
R13229 gnd.n6015 gnd.n5225 0.152939
R13230 gnd.n6066 gnd.n5225 0.152939
R13231 gnd.n6067 gnd.n6066 0.152939
R13232 gnd.n6068 gnd.n6067 0.152939
R13233 gnd.n6070 gnd.n6068 0.152939
R13234 gnd.n6070 gnd.n6069 0.152939
R13235 gnd.n6069 gnd.n913 0.152939
R13236 gnd.n914 gnd.n913 0.152939
R13237 gnd.n915 gnd.n914 0.152939
R13238 gnd.n935 gnd.n915 0.152939
R13239 gnd.n936 gnd.n935 0.152939
R13240 gnd.n937 gnd.n936 0.152939
R13241 gnd.n938 gnd.n937 0.152939
R13242 gnd.n939 gnd.n938 0.152939
R13243 gnd.n960 gnd.n939 0.152939
R13244 gnd.n961 gnd.n960 0.152939
R13245 gnd.n962 gnd.n961 0.152939
R13246 gnd.n6491 gnd.n962 0.152939
R13247 gnd.n5689 gnd.n5688 0.152939
R13248 gnd.n5690 gnd.n5689 0.152939
R13249 gnd.n5691 gnd.n5690 0.152939
R13250 gnd.n5692 gnd.n5691 0.152939
R13251 gnd.n5693 gnd.n5692 0.152939
R13252 gnd.n5694 gnd.n5693 0.152939
R13253 gnd.n5695 gnd.n5694 0.152939
R13254 gnd.n5696 gnd.n5695 0.152939
R13255 gnd.n5697 gnd.n5696 0.152939
R13256 gnd.n5698 gnd.n5697 0.152939
R13257 gnd.n5699 gnd.n5698 0.152939
R13258 gnd.n5700 gnd.n5699 0.152939
R13259 gnd.n5701 gnd.n5700 0.152939
R13260 gnd.n5702 gnd.n5701 0.152939
R13261 gnd.n5706 gnd.n5702 0.152939
R13262 gnd.n5706 gnd.n5484 0.152939
R13263 gnd.n6455 gnd.n5161 0.152939
R13264 gnd.n5163 gnd.n5161 0.152939
R13265 gnd.n5164 gnd.n5163 0.152939
R13266 gnd.n5165 gnd.n5164 0.152939
R13267 gnd.n5166 gnd.n5165 0.152939
R13268 gnd.n5167 gnd.n5166 0.152939
R13269 gnd.n5168 gnd.n5167 0.152939
R13270 gnd.n5169 gnd.n5168 0.152939
R13271 gnd.n5170 gnd.n5169 0.152939
R13272 gnd.n5171 gnd.n5170 0.152939
R13273 gnd.n5172 gnd.n5171 0.152939
R13274 gnd.n5173 gnd.n5172 0.152939
R13275 gnd.n5174 gnd.n5173 0.152939
R13276 gnd.n5175 gnd.n5174 0.152939
R13277 gnd.n5176 gnd.n5175 0.152939
R13278 gnd.n5177 gnd.n5176 0.152939
R13279 gnd.n5178 gnd.n5177 0.152939
R13280 gnd.n5179 gnd.n5178 0.152939
R13281 gnd.n5180 gnd.n5179 0.152939
R13282 gnd.n5181 gnd.n5180 0.152939
R13283 gnd.n5182 gnd.n5181 0.152939
R13284 gnd.n5183 gnd.n5182 0.152939
R13285 gnd.n5187 gnd.n5183 0.152939
R13286 gnd.n5188 gnd.n5187 0.152939
R13287 gnd.n5189 gnd.n5188 0.152939
R13288 gnd.n5190 gnd.n5189 0.152939
R13289 gnd.n5949 gnd.n5948 0.152939
R13290 gnd.n5950 gnd.n5949 0.152939
R13291 gnd.n5951 gnd.n5950 0.152939
R13292 gnd.n5952 gnd.n5951 0.152939
R13293 gnd.n5953 gnd.n5952 0.152939
R13294 gnd.n5954 gnd.n5953 0.152939
R13295 gnd.n5955 gnd.n5954 0.152939
R13296 gnd.n5956 gnd.n5955 0.152939
R13297 gnd.n5956 gnd.n5237 0.152939
R13298 gnd.n6034 gnd.n5237 0.152939
R13299 gnd.n6035 gnd.n6034 0.152939
R13300 gnd.n6036 gnd.n6035 0.152939
R13301 gnd.n6037 gnd.n6036 0.152939
R13302 gnd.n6038 gnd.n6037 0.152939
R13303 gnd.n6039 gnd.n6038 0.152939
R13304 gnd.n6040 gnd.n6039 0.152939
R13305 gnd.n6041 gnd.n6040 0.152939
R13306 gnd.n6041 gnd.n5203 0.152939
R13307 gnd.n6103 gnd.n5203 0.152939
R13308 gnd.n6104 gnd.n6103 0.152939
R13309 gnd.n6105 gnd.n6104 0.152939
R13310 gnd.n6106 gnd.n6105 0.152939
R13311 gnd.n6107 gnd.n6106 0.152939
R13312 gnd.n6108 gnd.n6107 0.152939
R13313 gnd.n6108 gnd.n5192 0.152939
R13314 gnd.n6398 gnd.n5192 0.152939
R13315 gnd.n6399 gnd.n6398 0.152939
R13316 gnd.n6400 gnd.n6399 0.152939
R13317 gnd.n5621 gnd.n5620 0.152939
R13318 gnd.n5622 gnd.n5621 0.152939
R13319 gnd.n5622 gnd.n5504 0.152939
R13320 gnd.n5636 gnd.n5504 0.152939
R13321 gnd.n5637 gnd.n5636 0.152939
R13322 gnd.n5638 gnd.n5637 0.152939
R13323 gnd.n5638 gnd.n5491 0.152939
R13324 gnd.n5652 gnd.n5491 0.152939
R13325 gnd.n5653 gnd.n5652 0.152939
R13326 gnd.n5654 gnd.n5653 0.152939
R13327 gnd.n5655 gnd.n5654 0.152939
R13328 gnd.n5656 gnd.n5655 0.152939
R13329 gnd.n5657 gnd.n5656 0.152939
R13330 gnd.n5658 gnd.n5657 0.152939
R13331 gnd.n5659 gnd.n5658 0.152939
R13332 gnd.n5660 gnd.n5659 0.152939
R13333 gnd.n5661 gnd.n5660 0.152939
R13334 gnd.n5662 gnd.n5661 0.152939
R13335 gnd.n5663 gnd.n5662 0.152939
R13336 gnd.n5663 gnd.n5426 0.152939
R13337 gnd.n5815 gnd.n5426 0.152939
R13338 gnd.n5816 gnd.n5815 0.152939
R13339 gnd.n5817 gnd.n5816 0.152939
R13340 gnd.n5818 gnd.n5817 0.152939
R13341 gnd.n5818 gnd.n5393 0.152939
R13342 gnd.n5862 gnd.n5393 0.152939
R13343 gnd.n5863 gnd.n5862 0.152939
R13344 gnd.n5864 gnd.n5863 0.152939
R13345 gnd.n5613 gnd.n5520 0.152939
R13346 gnd.n5523 gnd.n5520 0.152939
R13347 gnd.n5524 gnd.n5523 0.152939
R13348 gnd.n5525 gnd.n5524 0.152939
R13349 gnd.n5528 gnd.n5525 0.152939
R13350 gnd.n5529 gnd.n5528 0.152939
R13351 gnd.n5530 gnd.n5529 0.152939
R13352 gnd.n5531 gnd.n5530 0.152939
R13353 gnd.n5534 gnd.n5531 0.152939
R13354 gnd.n5535 gnd.n5534 0.152939
R13355 gnd.n5536 gnd.n5535 0.152939
R13356 gnd.n5537 gnd.n5536 0.152939
R13357 gnd.n5540 gnd.n5537 0.152939
R13358 gnd.n5541 gnd.n5540 0.152939
R13359 gnd.n5542 gnd.n5541 0.152939
R13360 gnd.n5543 gnd.n5542 0.152939
R13361 gnd.n5546 gnd.n5543 0.152939
R13362 gnd.n5547 gnd.n5546 0.152939
R13363 gnd.n5548 gnd.n5547 0.152939
R13364 gnd.n5549 gnd.n5548 0.152939
R13365 gnd.n5552 gnd.n5549 0.152939
R13366 gnd.n5553 gnd.n5552 0.152939
R13367 gnd.n5556 gnd.n5553 0.152939
R13368 gnd.n5557 gnd.n5556 0.152939
R13369 gnd.n5559 gnd.n5557 0.152939
R13370 gnd.n5559 gnd.n5516 0.152939
R13371 gnd.n6697 gnd.n737 0.152939
R13372 gnd.n6698 gnd.n6697 0.152939
R13373 gnd.n6699 gnd.n6698 0.152939
R13374 gnd.n6699 gnd.n731 0.152939
R13375 gnd.n6707 gnd.n731 0.152939
R13376 gnd.n6708 gnd.n6707 0.152939
R13377 gnd.n6709 gnd.n6708 0.152939
R13378 gnd.n6709 gnd.n725 0.152939
R13379 gnd.n6717 gnd.n725 0.152939
R13380 gnd.n6718 gnd.n6717 0.152939
R13381 gnd.n6719 gnd.n6718 0.152939
R13382 gnd.n6719 gnd.n719 0.152939
R13383 gnd.n6727 gnd.n719 0.152939
R13384 gnd.n6728 gnd.n6727 0.152939
R13385 gnd.n6729 gnd.n6728 0.152939
R13386 gnd.n6729 gnd.n713 0.152939
R13387 gnd.n6737 gnd.n713 0.152939
R13388 gnd.n6738 gnd.n6737 0.152939
R13389 gnd.n6739 gnd.n6738 0.152939
R13390 gnd.n6739 gnd.n707 0.152939
R13391 gnd.n6747 gnd.n707 0.152939
R13392 gnd.n6748 gnd.n6747 0.152939
R13393 gnd.n6749 gnd.n6748 0.152939
R13394 gnd.n6749 gnd.n701 0.152939
R13395 gnd.n6757 gnd.n701 0.152939
R13396 gnd.n6758 gnd.n6757 0.152939
R13397 gnd.n6759 gnd.n6758 0.152939
R13398 gnd.n6759 gnd.n695 0.152939
R13399 gnd.n6767 gnd.n695 0.152939
R13400 gnd.n6768 gnd.n6767 0.152939
R13401 gnd.n6769 gnd.n6768 0.152939
R13402 gnd.n6769 gnd.n689 0.152939
R13403 gnd.n6777 gnd.n689 0.152939
R13404 gnd.n6778 gnd.n6777 0.152939
R13405 gnd.n6779 gnd.n6778 0.152939
R13406 gnd.n6779 gnd.n683 0.152939
R13407 gnd.n6787 gnd.n683 0.152939
R13408 gnd.n6788 gnd.n6787 0.152939
R13409 gnd.n6789 gnd.n6788 0.152939
R13410 gnd.n6789 gnd.n677 0.152939
R13411 gnd.n6797 gnd.n677 0.152939
R13412 gnd.n6798 gnd.n6797 0.152939
R13413 gnd.n6799 gnd.n6798 0.152939
R13414 gnd.n6799 gnd.n671 0.152939
R13415 gnd.n6807 gnd.n671 0.152939
R13416 gnd.n6808 gnd.n6807 0.152939
R13417 gnd.n6809 gnd.n6808 0.152939
R13418 gnd.n6809 gnd.n665 0.152939
R13419 gnd.n6817 gnd.n665 0.152939
R13420 gnd.n6818 gnd.n6817 0.152939
R13421 gnd.n6819 gnd.n6818 0.152939
R13422 gnd.n6819 gnd.n659 0.152939
R13423 gnd.n6827 gnd.n659 0.152939
R13424 gnd.n6828 gnd.n6827 0.152939
R13425 gnd.n6829 gnd.n6828 0.152939
R13426 gnd.n6829 gnd.n653 0.152939
R13427 gnd.n6837 gnd.n653 0.152939
R13428 gnd.n6838 gnd.n6837 0.152939
R13429 gnd.n6839 gnd.n6838 0.152939
R13430 gnd.n6839 gnd.n647 0.152939
R13431 gnd.n6847 gnd.n647 0.152939
R13432 gnd.n6848 gnd.n6847 0.152939
R13433 gnd.n6849 gnd.n6848 0.152939
R13434 gnd.n6849 gnd.n641 0.152939
R13435 gnd.n6857 gnd.n641 0.152939
R13436 gnd.n6858 gnd.n6857 0.152939
R13437 gnd.n6859 gnd.n6858 0.152939
R13438 gnd.n6859 gnd.n635 0.152939
R13439 gnd.n6867 gnd.n635 0.152939
R13440 gnd.n6868 gnd.n6867 0.152939
R13441 gnd.n6869 gnd.n6868 0.152939
R13442 gnd.n6869 gnd.n629 0.152939
R13443 gnd.n6877 gnd.n629 0.152939
R13444 gnd.n6878 gnd.n6877 0.152939
R13445 gnd.n6879 gnd.n6878 0.152939
R13446 gnd.n6879 gnd.n623 0.152939
R13447 gnd.n6887 gnd.n623 0.152939
R13448 gnd.n6888 gnd.n6887 0.152939
R13449 gnd.n6889 gnd.n6888 0.152939
R13450 gnd.n6889 gnd.n617 0.152939
R13451 gnd.n6897 gnd.n617 0.152939
R13452 gnd.n6898 gnd.n6897 0.152939
R13453 gnd.n6899 gnd.n6898 0.152939
R13454 gnd.n6899 gnd.n611 0.152939
R13455 gnd.n6907 gnd.n611 0.152939
R13456 gnd.n6908 gnd.n6907 0.152939
R13457 gnd.n6909 gnd.n6908 0.152939
R13458 gnd.n6909 gnd.n605 0.152939
R13459 gnd.n6917 gnd.n605 0.152939
R13460 gnd.n6918 gnd.n6917 0.152939
R13461 gnd.n6919 gnd.n6918 0.152939
R13462 gnd.n6919 gnd.n599 0.152939
R13463 gnd.n6927 gnd.n599 0.152939
R13464 gnd.n6928 gnd.n6927 0.152939
R13465 gnd.n6929 gnd.n6928 0.152939
R13466 gnd.n6929 gnd.n593 0.152939
R13467 gnd.n6937 gnd.n593 0.152939
R13468 gnd.n6938 gnd.n6937 0.152939
R13469 gnd.n6939 gnd.n6938 0.152939
R13470 gnd.n6939 gnd.n587 0.152939
R13471 gnd.n6947 gnd.n587 0.152939
R13472 gnd.n6948 gnd.n6947 0.152939
R13473 gnd.n6949 gnd.n6948 0.152939
R13474 gnd.n6949 gnd.n581 0.152939
R13475 gnd.n6957 gnd.n581 0.152939
R13476 gnd.n6958 gnd.n6957 0.152939
R13477 gnd.n6959 gnd.n6958 0.152939
R13478 gnd.n6959 gnd.n575 0.152939
R13479 gnd.n6967 gnd.n575 0.152939
R13480 gnd.n6968 gnd.n6967 0.152939
R13481 gnd.n6969 gnd.n6968 0.152939
R13482 gnd.n6969 gnd.n569 0.152939
R13483 gnd.n6977 gnd.n569 0.152939
R13484 gnd.n6978 gnd.n6977 0.152939
R13485 gnd.n6979 gnd.n6978 0.152939
R13486 gnd.n6979 gnd.n563 0.152939
R13487 gnd.n6987 gnd.n563 0.152939
R13488 gnd.n6988 gnd.n6987 0.152939
R13489 gnd.n6989 gnd.n6988 0.152939
R13490 gnd.n6989 gnd.n557 0.152939
R13491 gnd.n6997 gnd.n557 0.152939
R13492 gnd.n6998 gnd.n6997 0.152939
R13493 gnd.n6999 gnd.n6998 0.152939
R13494 gnd.n6999 gnd.n551 0.152939
R13495 gnd.n7007 gnd.n551 0.152939
R13496 gnd.n7008 gnd.n7007 0.152939
R13497 gnd.n7009 gnd.n7008 0.152939
R13498 gnd.n7009 gnd.n545 0.152939
R13499 gnd.n7017 gnd.n545 0.152939
R13500 gnd.n7018 gnd.n7017 0.152939
R13501 gnd.n7019 gnd.n7018 0.152939
R13502 gnd.n7019 gnd.n539 0.152939
R13503 gnd.n7027 gnd.n539 0.152939
R13504 gnd.n7028 gnd.n7027 0.152939
R13505 gnd.n7029 gnd.n7028 0.152939
R13506 gnd.n7029 gnd.n533 0.152939
R13507 gnd.n7037 gnd.n533 0.152939
R13508 gnd.n7038 gnd.n7037 0.152939
R13509 gnd.n7039 gnd.n7038 0.152939
R13510 gnd.n7039 gnd.n527 0.152939
R13511 gnd.n7047 gnd.n527 0.152939
R13512 gnd.n7048 gnd.n7047 0.152939
R13513 gnd.n7049 gnd.n7048 0.152939
R13514 gnd.n7049 gnd.n521 0.152939
R13515 gnd.n7057 gnd.n521 0.152939
R13516 gnd.n7058 gnd.n7057 0.152939
R13517 gnd.n7059 gnd.n7058 0.152939
R13518 gnd.n7059 gnd.n515 0.152939
R13519 gnd.n7067 gnd.n515 0.152939
R13520 gnd.n7068 gnd.n7067 0.152939
R13521 gnd.n7069 gnd.n7068 0.152939
R13522 gnd.n7069 gnd.n509 0.152939
R13523 gnd.n7077 gnd.n509 0.152939
R13524 gnd.n7078 gnd.n7077 0.152939
R13525 gnd.n7079 gnd.n7078 0.152939
R13526 gnd.n7079 gnd.n503 0.152939
R13527 gnd.n7087 gnd.n503 0.152939
R13528 gnd.n7088 gnd.n7087 0.152939
R13529 gnd.n7089 gnd.n7088 0.152939
R13530 gnd.n7089 gnd.n497 0.152939
R13531 gnd.n7097 gnd.n497 0.152939
R13532 gnd.n7098 gnd.n7097 0.152939
R13533 gnd.n7099 gnd.n7098 0.152939
R13534 gnd.n7099 gnd.n491 0.152939
R13535 gnd.n7107 gnd.n491 0.152939
R13536 gnd.n7108 gnd.n7107 0.152939
R13537 gnd.n7109 gnd.n7108 0.152939
R13538 gnd.n7109 gnd.n485 0.152939
R13539 gnd.n7117 gnd.n485 0.152939
R13540 gnd.n7118 gnd.n7117 0.152939
R13541 gnd.n7119 gnd.n7118 0.152939
R13542 gnd.n7119 gnd.n479 0.152939
R13543 gnd.n7127 gnd.n479 0.152939
R13544 gnd.n7128 gnd.n7127 0.152939
R13545 gnd.n7129 gnd.n7128 0.152939
R13546 gnd.n7129 gnd.n473 0.152939
R13547 gnd.n7137 gnd.n473 0.152939
R13548 gnd.n7138 gnd.n7137 0.152939
R13549 gnd.n7139 gnd.n7138 0.152939
R13550 gnd.n7139 gnd.n467 0.152939
R13551 gnd.n7147 gnd.n467 0.152939
R13552 gnd.n7148 gnd.n7147 0.152939
R13553 gnd.n7149 gnd.n7148 0.152939
R13554 gnd.n7149 gnd.n461 0.152939
R13555 gnd.n7157 gnd.n461 0.152939
R13556 gnd.n7158 gnd.n7157 0.152939
R13557 gnd.n7159 gnd.n7158 0.152939
R13558 gnd.n7159 gnd.n455 0.152939
R13559 gnd.n7167 gnd.n455 0.152939
R13560 gnd.n7168 gnd.n7167 0.152939
R13561 gnd.n7170 gnd.n7168 0.152939
R13562 gnd.n7170 gnd.n7169 0.152939
R13563 gnd.n7169 gnd.n449 0.152939
R13564 gnd.n7179 gnd.n449 0.152939
R13565 gnd.n7180 gnd.n444 0.152939
R13566 gnd.n7188 gnd.n444 0.152939
R13567 gnd.n7189 gnd.n7188 0.152939
R13568 gnd.n7190 gnd.n7189 0.152939
R13569 gnd.n7190 gnd.n438 0.152939
R13570 gnd.n7198 gnd.n438 0.152939
R13571 gnd.n7199 gnd.n7198 0.152939
R13572 gnd.n7200 gnd.n7199 0.152939
R13573 gnd.n7200 gnd.n432 0.152939
R13574 gnd.n7208 gnd.n432 0.152939
R13575 gnd.n7209 gnd.n7208 0.152939
R13576 gnd.n7210 gnd.n7209 0.152939
R13577 gnd.n7210 gnd.n426 0.152939
R13578 gnd.n7218 gnd.n426 0.152939
R13579 gnd.n7219 gnd.n7218 0.152939
R13580 gnd.n7220 gnd.n7219 0.152939
R13581 gnd.n7220 gnd.n420 0.152939
R13582 gnd.n7228 gnd.n420 0.152939
R13583 gnd.n7229 gnd.n7228 0.152939
R13584 gnd.n7230 gnd.n7229 0.152939
R13585 gnd.n7230 gnd.n414 0.152939
R13586 gnd.n7238 gnd.n414 0.152939
R13587 gnd.n7239 gnd.n7238 0.152939
R13588 gnd.n7240 gnd.n7239 0.152939
R13589 gnd.n7240 gnd.n408 0.152939
R13590 gnd.n7248 gnd.n408 0.152939
R13591 gnd.n7249 gnd.n7248 0.152939
R13592 gnd.n7250 gnd.n7249 0.152939
R13593 gnd.n7250 gnd.n402 0.152939
R13594 gnd.n7258 gnd.n402 0.152939
R13595 gnd.n7259 gnd.n7258 0.152939
R13596 gnd.n7260 gnd.n7259 0.152939
R13597 gnd.n7260 gnd.n396 0.152939
R13598 gnd.n7268 gnd.n396 0.152939
R13599 gnd.n7269 gnd.n7268 0.152939
R13600 gnd.n7270 gnd.n7269 0.152939
R13601 gnd.n7270 gnd.n390 0.152939
R13602 gnd.n7278 gnd.n390 0.152939
R13603 gnd.n7279 gnd.n7278 0.152939
R13604 gnd.n7280 gnd.n7279 0.152939
R13605 gnd.n7280 gnd.n384 0.152939
R13606 gnd.n7288 gnd.n384 0.152939
R13607 gnd.n7289 gnd.n7288 0.152939
R13608 gnd.n7290 gnd.n7289 0.152939
R13609 gnd.n7290 gnd.n378 0.152939
R13610 gnd.n7298 gnd.n378 0.152939
R13611 gnd.n7299 gnd.n7298 0.152939
R13612 gnd.n7300 gnd.n7299 0.152939
R13613 gnd.n7300 gnd.n372 0.152939
R13614 gnd.n7308 gnd.n372 0.152939
R13615 gnd.n7309 gnd.n7308 0.152939
R13616 gnd.n7310 gnd.n7309 0.152939
R13617 gnd.n7310 gnd.n366 0.152939
R13618 gnd.n7318 gnd.n366 0.152939
R13619 gnd.n7319 gnd.n7318 0.152939
R13620 gnd.n7320 gnd.n7319 0.152939
R13621 gnd.n7320 gnd.n360 0.152939
R13622 gnd.n7328 gnd.n360 0.152939
R13623 gnd.n7329 gnd.n7328 0.152939
R13624 gnd.n7330 gnd.n7329 0.152939
R13625 gnd.n7330 gnd.n354 0.152939
R13626 gnd.n7338 gnd.n354 0.152939
R13627 gnd.n7339 gnd.n7338 0.152939
R13628 gnd.n7340 gnd.n7339 0.152939
R13629 gnd.n7340 gnd.n348 0.152939
R13630 gnd.n7348 gnd.n348 0.152939
R13631 gnd.n7349 gnd.n7348 0.152939
R13632 gnd.n7350 gnd.n7349 0.152939
R13633 gnd.n7350 gnd.n342 0.152939
R13634 gnd.n7358 gnd.n342 0.152939
R13635 gnd.n7359 gnd.n7358 0.152939
R13636 gnd.n7360 gnd.n7359 0.152939
R13637 gnd.n7360 gnd.n336 0.152939
R13638 gnd.n7368 gnd.n336 0.152939
R13639 gnd.n7369 gnd.n7368 0.152939
R13640 gnd.n7370 gnd.n7369 0.152939
R13641 gnd.n7370 gnd.n330 0.152939
R13642 gnd.n7378 gnd.n330 0.152939
R13643 gnd.n7379 gnd.n7378 0.152939
R13644 gnd.n7380 gnd.n7379 0.152939
R13645 gnd.n7380 gnd.n324 0.152939
R13646 gnd.n7389 gnd.n324 0.152939
R13647 gnd.n7390 gnd.n7389 0.152939
R13648 gnd.n7391 gnd.n7390 0.152939
R13649 gnd.n312 gnd.n309 0.152939
R13650 gnd.n313 gnd.n312 0.152939
R13651 gnd.n314 gnd.n313 0.152939
R13652 gnd.n315 gnd.n314 0.152939
R13653 gnd.n318 gnd.n315 0.152939
R13654 gnd.n319 gnd.n318 0.152939
R13655 gnd.n320 gnd.n319 0.152939
R13656 gnd.n321 gnd.n320 0.152939
R13657 gnd.n7516 gnd.n252 0.152939
R13658 gnd.n7517 gnd.n7516 0.152939
R13659 gnd.n7518 gnd.n7517 0.152939
R13660 gnd.n7518 gnd.n236 0.152939
R13661 gnd.n7532 gnd.n236 0.152939
R13662 gnd.n7533 gnd.n7532 0.152939
R13663 gnd.n7534 gnd.n7533 0.152939
R13664 gnd.n7534 gnd.n222 0.152939
R13665 gnd.n7548 gnd.n222 0.152939
R13666 gnd.n7549 gnd.n7548 0.152939
R13667 gnd.n7550 gnd.n7549 0.152939
R13668 gnd.n7550 gnd.n205 0.152939
R13669 gnd.n7564 gnd.n205 0.152939
R13670 gnd.n7565 gnd.n7564 0.152939
R13671 gnd.n7566 gnd.n7565 0.152939
R13672 gnd.n7566 gnd.n190 0.152939
R13673 gnd.n7655 gnd.n190 0.152939
R13674 gnd.n7656 gnd.n7655 0.152939
R13675 gnd.n7657 gnd.n7656 0.152939
R13676 gnd.n7657 gnd.n111 0.152939
R13677 gnd.n7737 gnd.n111 0.152939
R13678 gnd.n7736 gnd.n112 0.152939
R13679 gnd.n114 gnd.n112 0.152939
R13680 gnd.n119 gnd.n114 0.152939
R13681 gnd.n120 gnd.n119 0.152939
R13682 gnd.n121 gnd.n120 0.152939
R13683 gnd.n122 gnd.n121 0.152939
R13684 gnd.n126 gnd.n122 0.152939
R13685 gnd.n127 gnd.n126 0.152939
R13686 gnd.n128 gnd.n127 0.152939
R13687 gnd.n129 gnd.n128 0.152939
R13688 gnd.n133 gnd.n129 0.152939
R13689 gnd.n134 gnd.n133 0.152939
R13690 gnd.n135 gnd.n134 0.152939
R13691 gnd.n136 gnd.n135 0.152939
R13692 gnd.n140 gnd.n136 0.152939
R13693 gnd.n141 gnd.n140 0.152939
R13694 gnd.n142 gnd.n141 0.152939
R13695 gnd.n143 gnd.n142 0.152939
R13696 gnd.n147 gnd.n143 0.152939
R13697 gnd.n148 gnd.n147 0.152939
R13698 gnd.n149 gnd.n148 0.152939
R13699 gnd.n150 gnd.n149 0.152939
R13700 gnd.n154 gnd.n150 0.152939
R13701 gnd.n155 gnd.n154 0.152939
R13702 gnd.n156 gnd.n155 0.152939
R13703 gnd.n157 gnd.n156 0.152939
R13704 gnd.n161 gnd.n157 0.152939
R13705 gnd.n162 gnd.n161 0.152939
R13706 gnd.n163 gnd.n162 0.152939
R13707 gnd.n164 gnd.n163 0.152939
R13708 gnd.n168 gnd.n164 0.152939
R13709 gnd.n169 gnd.n168 0.152939
R13710 gnd.n170 gnd.n169 0.152939
R13711 gnd.n171 gnd.n170 0.152939
R13712 gnd.n175 gnd.n171 0.152939
R13713 gnd.n176 gnd.n175 0.152939
R13714 gnd.n7667 gnd.n176 0.152939
R13715 gnd.n7667 gnd.n7666 0.152939
R13716 gnd.n1982 gnd.n1981 0.152939
R13717 gnd.n1981 gnd.n1639 0.152939
R13718 gnd.n4488 gnd.n1639 0.152939
R13719 gnd.n4489 gnd.n4488 0.152939
R13720 gnd.n4490 gnd.n4489 0.152939
R13721 gnd.n4491 gnd.n4490 0.152939
R13722 gnd.n4492 gnd.n4491 0.152939
R13723 gnd.n4493 gnd.n4492 0.152939
R13724 gnd.n4494 gnd.n4493 0.152939
R13725 gnd.n4495 gnd.n4494 0.152939
R13726 gnd.n4496 gnd.n4495 0.152939
R13727 gnd.n4497 gnd.n4496 0.152939
R13728 gnd.n4498 gnd.n4497 0.152939
R13729 gnd.n4499 gnd.n4498 0.152939
R13730 gnd.n4501 gnd.n4499 0.152939
R13731 gnd.n4501 gnd.n4500 0.152939
R13732 gnd.n4500 gnd.n1559 0.152939
R13733 gnd.n1559 gnd.n1557 0.152939
R13734 gnd.n4615 gnd.n1557 0.152939
R13735 gnd.n4616 gnd.n4615 0.152939
R13736 gnd.n4617 gnd.n4616 0.152939
R13737 gnd.n4618 gnd.n4617 0.152939
R13738 gnd.n4618 gnd.n1549 0.152939
R13739 gnd.n4638 gnd.n1549 0.152939
R13740 gnd.n4639 gnd.n4638 0.152939
R13741 gnd.n4640 gnd.n4639 0.152939
R13742 gnd.n301 gnd.n300 0.152939
R13743 gnd.n302 gnd.n301 0.152939
R13744 gnd.n303 gnd.n302 0.152939
R13745 gnd.n7402 gnd.n303 0.152939
R13746 gnd.n7406 gnd.n7402 0.152939
R13747 gnd.n7407 gnd.n7406 0.152939
R13748 gnd.n7408 gnd.n7407 0.152939
R13749 gnd.n7408 gnd.n7400 0.152939
R13750 gnd.n7417 gnd.n7400 0.152939
R13751 gnd.n7418 gnd.n7417 0.152939
R13752 gnd.n7419 gnd.n7418 0.152939
R13753 gnd.n7420 gnd.n7419 0.152939
R13754 gnd.n7421 gnd.n7420 0.152939
R13755 gnd.n7422 gnd.n7421 0.152939
R13756 gnd.n7423 gnd.n7422 0.152939
R13757 gnd.n7424 gnd.n7423 0.152939
R13758 gnd.n7425 gnd.n7424 0.152939
R13759 gnd.n7426 gnd.n7425 0.152939
R13760 gnd.n7427 gnd.n7426 0.152939
R13761 gnd.n7428 gnd.n7427 0.152939
R13762 gnd.n7429 gnd.n7428 0.152939
R13763 gnd.n7430 gnd.n7429 0.152939
R13764 gnd.n7432 gnd.n7430 0.152939
R13765 gnd.n7432 gnd.n7431 0.152939
R13766 gnd.n7431 gnd.n182 0.152939
R13767 gnd.n7665 gnd.n182 0.152939
R13768 gnd.n1913 gnd.n1907 0.152939
R13769 gnd.n1914 gnd.n1913 0.152939
R13770 gnd.n1915 gnd.n1914 0.152939
R13771 gnd.n1915 gnd.n1902 0.152939
R13772 gnd.n1923 gnd.n1902 0.152939
R13773 gnd.n1924 gnd.n1923 0.152939
R13774 gnd.n1925 gnd.n1924 0.152939
R13775 gnd.n1925 gnd.n1898 0.152939
R13776 gnd.n1933 gnd.n1898 0.152939
R13777 gnd.n1934 gnd.n1933 0.152939
R13778 gnd.n1936 gnd.n1934 0.152939
R13779 gnd.n1936 gnd.n1935 0.152939
R13780 gnd.n1935 gnd.n1891 0.152939
R13781 gnd.n1945 gnd.n1891 0.152939
R13782 gnd.n1946 gnd.n1945 0.152939
R13783 gnd.n1953 gnd.n1950 0.152939
R13784 gnd.n1954 gnd.n1953 0.152939
R13785 gnd.n1955 gnd.n1954 0.152939
R13786 gnd.n1956 gnd.n1955 0.152939
R13787 gnd.n1959 gnd.n1956 0.152939
R13788 gnd.n1960 gnd.n1959 0.152939
R13789 gnd.n1961 gnd.n1960 0.152939
R13790 gnd.n1962 gnd.n1961 0.152939
R13791 gnd.n1965 gnd.n1962 0.152939
R13792 gnd.n1966 gnd.n1965 0.152939
R13793 gnd.n1967 gnd.n1966 0.152939
R13794 gnd.n1968 gnd.n1967 0.152939
R13795 gnd.n1971 gnd.n1968 0.152939
R13796 gnd.n1972 gnd.n1971 0.152939
R13797 gnd.n1973 gnd.n1972 0.152939
R13798 gnd.n1974 gnd.n1973 0.152939
R13799 gnd.n1980 gnd.n1974 0.152939
R13800 gnd.n1990 gnd.n1980 0.152939
R13801 gnd.n1990 gnd.n1989 0.152939
R13802 gnd.n1989 gnd.n1988 0.152939
R13803 gnd.n1906 gnd.n1485 0.152939
R13804 gnd.n1486 gnd.n1485 0.152939
R13805 gnd.n1487 gnd.n1486 0.152939
R13806 gnd.n4519 gnd.n1487 0.152939
R13807 gnd.n4520 gnd.n4519 0.152939
R13808 gnd.n4521 gnd.n4520 0.152939
R13809 gnd.n4521 gnd.n1602 0.152939
R13810 gnd.n4550 gnd.n1602 0.152939
R13811 gnd.n4551 gnd.n4550 0.152939
R13812 gnd.n4552 gnd.n4551 0.152939
R13813 gnd.n4553 gnd.n4552 0.152939
R13814 gnd.n4553 gnd.n1575 0.152939
R13815 gnd.n4589 gnd.n1575 0.152939
R13816 gnd.n4590 gnd.n4589 0.152939
R13817 gnd.n4591 gnd.n4590 0.152939
R13818 gnd.n4592 gnd.n4591 0.152939
R13819 gnd.n4592 gnd.n1523 0.152939
R13820 gnd.n4679 gnd.n1523 0.152939
R13821 gnd.n4680 gnd.n4679 0.152939
R13822 gnd.n4681 gnd.n4680 0.152939
R13823 gnd.n4681 gnd.n267 0.152939
R13824 gnd.n2883 gnd.n2877 0.152939
R13825 gnd.n2886 gnd.n2883 0.152939
R13826 gnd.n2887 gnd.n2886 0.152939
R13827 gnd.n2888 gnd.n2887 0.152939
R13828 gnd.n2889 gnd.n2888 0.152939
R13829 gnd.n2892 gnd.n2889 0.152939
R13830 gnd.n2893 gnd.n2892 0.152939
R13831 gnd.n2894 gnd.n2893 0.152939
R13832 gnd.n2895 gnd.n2894 0.152939
R13833 gnd.n2896 gnd.n2895 0.152939
R13834 gnd.n2897 gnd.n2896 0.152939
R13835 gnd.n2897 gnd.n2791 0.152939
R13836 gnd.n3242 gnd.n2791 0.152939
R13837 gnd.n3243 gnd.n3242 0.152939
R13838 gnd.n3244 gnd.n3243 0.152939
R13839 gnd.n3244 gnd.n2787 0.152939
R13840 gnd.n3250 gnd.n2787 0.152939
R13841 gnd.n3251 gnd.n3250 0.152939
R13842 gnd.n3252 gnd.n3251 0.152939
R13843 gnd.n3252 gnd.n2783 0.152939
R13844 gnd.n3258 gnd.n2783 0.152939
R13845 gnd.n3259 gnd.n3258 0.152939
R13846 gnd.n3260 gnd.n3259 0.152939
R13847 gnd.n3260 gnd.n2778 0.152939
R13848 gnd.n3401 gnd.n2778 0.152939
R13849 gnd.n3402 gnd.n3401 0.152939
R13850 gnd.n3403 gnd.n3402 0.152939
R13851 gnd.n3403 gnd.n2772 0.152939
R13852 gnd.n3415 gnd.n2772 0.152939
R13853 gnd.n3416 gnd.n3415 0.152939
R13854 gnd.n3417 gnd.n3416 0.152939
R13855 gnd.n3417 gnd.n2764 0.152939
R13856 gnd.n3429 gnd.n2764 0.152939
R13857 gnd.n3430 gnd.n3429 0.152939
R13858 gnd.n3431 gnd.n3430 0.152939
R13859 gnd.n3431 gnd.n2756 0.152939
R13860 gnd.n3446 gnd.n2756 0.152939
R13861 gnd.n3447 gnd.n3446 0.152939
R13862 gnd.n3448 gnd.n3447 0.152939
R13863 gnd.n3448 gnd.n2751 0.152939
R13864 gnd.n3460 gnd.n2751 0.152939
R13865 gnd.n3461 gnd.n3460 0.152939
R13866 gnd.n3462 gnd.n3461 0.152939
R13867 gnd.n3463 gnd.n3462 0.152939
R13868 gnd.n3463 gnd.n2397 0.152939
R13869 gnd.n3649 gnd.n2397 0.152939
R13870 gnd.n3650 gnd.n3649 0.152939
R13871 gnd.n3651 gnd.n3650 0.152939
R13872 gnd.n3651 gnd.n2376 0.152939
R13873 gnd.n3678 gnd.n2376 0.152939
R13874 gnd.n3679 gnd.n3678 0.152939
R13875 gnd.n3680 gnd.n3679 0.152939
R13876 gnd.n3681 gnd.n3680 0.152939
R13877 gnd.n3681 gnd.n2349 0.152939
R13878 gnd.n3716 gnd.n2349 0.152939
R13879 gnd.n3717 gnd.n3716 0.152939
R13880 gnd.n3718 gnd.n3717 0.152939
R13881 gnd.n3719 gnd.n3718 0.152939
R13882 gnd.n3719 gnd.n2322 0.152939
R13883 gnd.n3752 gnd.n2322 0.152939
R13884 gnd.n3753 gnd.n3752 0.152939
R13885 gnd.n3754 gnd.n3753 0.152939
R13886 gnd.n3754 gnd.n2300 0.152939
R13887 gnd.n3780 gnd.n2300 0.152939
R13888 gnd.n3781 gnd.n3780 0.152939
R13889 gnd.n3782 gnd.n3781 0.152939
R13890 gnd.n3783 gnd.n3782 0.152939
R13891 gnd.n3783 gnd.n2272 0.152939
R13892 gnd.n3830 gnd.n2272 0.152939
R13893 gnd.n3831 gnd.n3830 0.152939
R13894 gnd.n3832 gnd.n3831 0.152939
R13895 gnd.n3833 gnd.n3832 0.152939
R13896 gnd.n3833 gnd.n2253 0.152939
R13897 gnd.n3857 gnd.n2253 0.152939
R13898 gnd.n3858 gnd.n3857 0.152939
R13899 gnd.n3859 gnd.n3858 0.152939
R13900 gnd.n3859 gnd.n2208 0.152939
R13901 gnd.n3900 gnd.n2208 0.152939
R13902 gnd.n3901 gnd.n3900 0.152939
R13903 gnd.n3902 gnd.n3901 0.152939
R13904 gnd.n3902 gnd.n2186 0.152939
R13905 gnd.n3942 gnd.n2186 0.152939
R13906 gnd.n3943 gnd.n3942 0.152939
R13907 gnd.n3944 gnd.n3943 0.152939
R13908 gnd.n3945 gnd.n3944 0.152939
R13909 gnd.n3945 gnd.n2159 0.152939
R13910 gnd.n3994 gnd.n2159 0.152939
R13911 gnd.n3995 gnd.n3994 0.152939
R13912 gnd.n3996 gnd.n3995 0.152939
R13913 gnd.n3997 gnd.n3996 0.152939
R13914 gnd.n3997 gnd.n2128 0.152939
R13915 gnd.n4045 gnd.n2128 0.152939
R13916 gnd.n4046 gnd.n4045 0.152939
R13917 gnd.n4047 gnd.n4046 0.152939
R13918 gnd.n4047 gnd.n2113 0.152939
R13919 gnd.n4077 gnd.n2113 0.152939
R13920 gnd.n4078 gnd.n4077 0.152939
R13921 gnd.n4079 gnd.n4078 0.152939
R13922 gnd.n4080 gnd.n4079 0.152939
R13923 gnd.n4081 gnd.n4080 0.152939
R13924 gnd.n4081 gnd.n2078 0.152939
R13925 gnd.n4151 gnd.n2078 0.152939
R13926 gnd.n4152 gnd.n4151 0.152939
R13927 gnd.n4153 gnd.n4152 0.152939
R13928 gnd.n4154 gnd.n4153 0.152939
R13929 gnd.n4154 gnd.n2050 0.152939
R13930 gnd.n4194 gnd.n2050 0.152939
R13931 gnd.n4195 gnd.n4194 0.152939
R13932 gnd.n4196 gnd.n4195 0.152939
R13933 gnd.n4197 gnd.n4196 0.152939
R13934 gnd.n4198 gnd.n4197 0.152939
R13935 gnd.n4198 gnd.n1844 0.152939
R13936 gnd.n4380 gnd.n1844 0.152939
R13937 gnd.n4381 gnd.n4380 0.152939
R13938 gnd.n4382 gnd.n4381 0.152939
R13939 gnd.n4382 gnd.n1831 0.152939
R13940 gnd.n4400 gnd.n1831 0.152939
R13941 gnd.n4401 gnd.n4400 0.152939
R13942 gnd.n4402 gnd.n4401 0.152939
R13943 gnd.n4402 gnd.n1818 0.152939
R13944 gnd.n4420 gnd.n1818 0.152939
R13945 gnd.n4421 gnd.n4420 0.152939
R13946 gnd.n4422 gnd.n4421 0.152939
R13947 gnd.n4422 gnd.n1805 0.152939
R13948 gnd.n4443 gnd.n1805 0.152939
R13949 gnd.n4444 gnd.n4443 0.152939
R13950 gnd.n4446 gnd.n4444 0.152939
R13951 gnd.n4446 gnd.n4445 0.152939
R13952 gnd.n4445 gnd.n1462 0.152939
R13953 gnd.n1463 gnd.n1462 0.152939
R13954 gnd.n1464 gnd.n1463 0.152939
R13955 gnd.n1470 gnd.n1464 0.152939
R13956 gnd.n1471 gnd.n1470 0.152939
R13957 gnd.n1472 gnd.n1471 0.152939
R13958 gnd.n1473 gnd.n1472 0.152939
R13959 gnd.n1626 gnd.n1473 0.152939
R13960 gnd.n1629 gnd.n1626 0.152939
R13961 gnd.n1630 gnd.n1629 0.152939
R13962 gnd.n1631 gnd.n1630 0.152939
R13963 gnd.n1631 gnd.n1613 0.152939
R13964 gnd.n4538 gnd.n1613 0.152939
R13965 gnd.n4539 gnd.n4538 0.152939
R13966 gnd.n4540 gnd.n4539 0.152939
R13967 gnd.n4541 gnd.n4540 0.152939
R13968 gnd.n4541 gnd.n1586 0.152939
R13969 gnd.n4571 gnd.n1586 0.152939
R13970 gnd.n4572 gnd.n4571 0.152939
R13971 gnd.n4573 gnd.n4572 0.152939
R13972 gnd.n4574 gnd.n4573 0.152939
R13973 gnd.n4575 gnd.n4574 0.152939
R13974 gnd.n4577 gnd.n4575 0.152939
R13975 gnd.n4577 gnd.n4576 0.152939
R13976 gnd.n4576 gnd.n1533 0.152939
R13977 gnd.n1534 gnd.n1533 0.152939
R13978 gnd.n1535 gnd.n1534 0.152939
R13979 gnd.n1536 gnd.n1535 0.152939
R13980 gnd.n1213 gnd.n1212 0.152939
R13981 gnd.n1230 gnd.n1213 0.152939
R13982 gnd.n1231 gnd.n1230 0.152939
R13983 gnd.n1232 gnd.n1231 0.152939
R13984 gnd.n1233 gnd.n1232 0.152939
R13985 gnd.n1252 gnd.n1233 0.152939
R13986 gnd.n1253 gnd.n1252 0.152939
R13987 gnd.n1254 gnd.n1253 0.152939
R13988 gnd.n1255 gnd.n1254 0.152939
R13989 gnd.n1272 gnd.n1255 0.152939
R13990 gnd.n1273 gnd.n1272 0.152939
R13991 gnd.n1274 gnd.n1273 0.152939
R13992 gnd.n1275 gnd.n1274 0.152939
R13993 gnd.n1294 gnd.n1275 0.152939
R13994 gnd.n1295 gnd.n1294 0.152939
R13995 gnd.n1296 gnd.n1295 0.152939
R13996 gnd.n1297 gnd.n1296 0.152939
R13997 gnd.n1315 gnd.n1297 0.152939
R13998 gnd.n1316 gnd.n1315 0.152939
R13999 gnd.n1317 gnd.n1316 0.152939
R14000 gnd.n1318 gnd.n1317 0.152939
R14001 gnd.n2625 gnd.n2624 0.152939
R14002 gnd.n2626 gnd.n2625 0.152939
R14003 gnd.n2627 gnd.n2626 0.152939
R14004 gnd.n2628 gnd.n2627 0.152939
R14005 gnd.n2629 gnd.n2628 0.152939
R14006 gnd.n2630 gnd.n2629 0.152939
R14007 gnd.n2631 gnd.n2630 0.152939
R14008 gnd.n2632 gnd.n2631 0.152939
R14009 gnd.n2633 gnd.n2632 0.152939
R14010 gnd.n2634 gnd.n2633 0.152939
R14011 gnd.n2635 gnd.n2634 0.152939
R14012 gnd.n2636 gnd.n2635 0.152939
R14013 gnd.n2637 gnd.n2636 0.152939
R14014 gnd.n2638 gnd.n2637 0.152939
R14015 gnd.n2638 gnd.n2608 0.152939
R14016 gnd.n3571 gnd.n3570 0.152939
R14017 gnd.n3570 gnd.n2609 0.152939
R14018 gnd.n2669 gnd.n2609 0.152939
R14019 gnd.n2670 gnd.n2669 0.152939
R14020 gnd.n2671 gnd.n2670 0.152939
R14021 gnd.n2672 gnd.n2671 0.152939
R14022 gnd.n2676 gnd.n2672 0.152939
R14023 gnd.n2677 gnd.n2676 0.152939
R14024 gnd.n2678 gnd.n2677 0.152939
R14025 gnd.n2679 gnd.n2678 0.152939
R14026 gnd.n2683 gnd.n2679 0.152939
R14027 gnd.n2684 gnd.n2683 0.152939
R14028 gnd.n2685 gnd.n2684 0.152939
R14029 gnd.n2686 gnd.n2685 0.152939
R14030 gnd.n2690 gnd.n2686 0.152939
R14031 gnd.n2691 gnd.n2690 0.152939
R14032 gnd.n2692 gnd.n2691 0.152939
R14033 gnd.n2693 gnd.n2692 0.152939
R14034 gnd.n2698 gnd.n2693 0.152939
R14035 gnd.n3533 gnd.n2698 0.152939
R14036 gnd.n2984 gnd.n2982 0.152939
R14037 gnd.n2982 gnd.n2957 0.152939
R14038 gnd.n2957 gnd.n2955 0.152939
R14039 gnd.n3045 gnd.n2955 0.152939
R14040 gnd.n3046 gnd.n3045 0.152939
R14041 gnd.n3047 gnd.n3046 0.152939
R14042 gnd.n3047 gnd.n2953 0.152939
R14043 gnd.n3053 gnd.n2953 0.152939
R14044 gnd.n3054 gnd.n3053 0.152939
R14045 gnd.n3055 gnd.n3054 0.152939
R14046 gnd.n3055 gnd.n2951 0.152939
R14047 gnd.n3082 gnd.n2951 0.152939
R14048 gnd.n3083 gnd.n3082 0.152939
R14049 gnd.n3084 gnd.n3083 0.152939
R14050 gnd.n3084 gnd.n2945 0.152939
R14051 gnd.n3098 gnd.n2945 0.152939
R14052 gnd.n3099 gnd.n3098 0.152939
R14053 gnd.n3100 gnd.n3099 0.152939
R14054 gnd.n3100 gnd.n2845 0.152939
R14055 gnd.n3114 gnd.n2845 0.152939
R14056 gnd.n3115 gnd.n3114 0.152939
R14057 gnd.n3116 gnd.n3115 0.152939
R14058 gnd.n3116 gnd.n2839 0.152939
R14059 gnd.n3130 gnd.n2839 0.152939
R14060 gnd.n3131 gnd.n3130 0.152939
R14061 gnd.n3133 gnd.n3131 0.152939
R14062 gnd.n3023 gnd.n2963 0.152939
R14063 gnd.n2964 gnd.n2963 0.152939
R14064 gnd.n2965 gnd.n2964 0.152939
R14065 gnd.n2966 gnd.n2965 0.152939
R14066 gnd.n2967 gnd.n2966 0.152939
R14067 gnd.n2968 gnd.n2967 0.152939
R14068 gnd.n2969 gnd.n2968 0.152939
R14069 gnd.n2970 gnd.n2969 0.152939
R14070 gnd.n2971 gnd.n2970 0.152939
R14071 gnd.n2972 gnd.n2971 0.152939
R14072 gnd.n2973 gnd.n2972 0.152939
R14073 gnd.n2974 gnd.n2973 0.152939
R14074 gnd.n2975 gnd.n2974 0.152939
R14075 gnd.n2976 gnd.n2975 0.152939
R14076 gnd.n2977 gnd.n2976 0.152939
R14077 gnd.n2988 gnd.n2977 0.152939
R14078 gnd.n2988 gnd.n2987 0.152939
R14079 gnd.n2987 gnd.n2986 0.152939
R14080 gnd.n3029 gnd.n3024 0.152939
R14081 gnd.n3029 gnd.n3028 0.152939
R14082 gnd.n3028 gnd.n3027 0.152939
R14083 gnd.n3027 gnd.n3025 0.152939
R14084 gnd.n3025 gnd.n1081 0.152939
R14085 gnd.n1082 gnd.n1081 0.152939
R14086 gnd.n1083 gnd.n1082 0.152939
R14087 gnd.n1099 gnd.n1083 0.152939
R14088 gnd.n1100 gnd.n1099 0.152939
R14089 gnd.n1101 gnd.n1100 0.152939
R14090 gnd.n1102 gnd.n1101 0.152939
R14091 gnd.n1121 gnd.n1102 0.152939
R14092 gnd.n1122 gnd.n1121 0.152939
R14093 gnd.n1123 gnd.n1122 0.152939
R14094 gnd.n1124 gnd.n1123 0.152939
R14095 gnd.n1142 gnd.n1124 0.152939
R14096 gnd.n1143 gnd.n1142 0.152939
R14097 gnd.n1144 gnd.n1143 0.152939
R14098 gnd.n1145 gnd.n1144 0.152939
R14099 gnd.n1163 gnd.n1145 0.152939
R14100 gnd.n1164 gnd.n1163 0.152939
R14101 gnd.n1165 gnd.n1164 0.152939
R14102 gnd.n1166 gnd.n1165 0.152939
R14103 gnd.n1182 gnd.n1166 0.152939
R14104 gnd.n1183 gnd.n1182 0.152939
R14105 gnd.n1184 gnd.n1183 0.152939
R14106 gnd.n1200 gnd.n1185 0.152939
R14107 gnd.n1201 gnd.n1200 0.152939
R14108 gnd.n1202 gnd.n1201 0.152939
R14109 gnd.n1203 gnd.n1202 0.152939
R14110 gnd.n1220 gnd.n1203 0.152939
R14111 gnd.n1221 gnd.n1220 0.152939
R14112 gnd.n1222 gnd.n1221 0.152939
R14113 gnd.n1223 gnd.n1222 0.152939
R14114 gnd.n1241 gnd.n1223 0.152939
R14115 gnd.n1242 gnd.n1241 0.152939
R14116 gnd.n1243 gnd.n1242 0.152939
R14117 gnd.n1244 gnd.n1243 0.152939
R14118 gnd.n1262 gnd.n1244 0.152939
R14119 gnd.n1263 gnd.n1262 0.152939
R14120 gnd.n1264 gnd.n1263 0.152939
R14121 gnd.n1265 gnd.n1264 0.152939
R14122 gnd.n1283 gnd.n1265 0.152939
R14123 gnd.n1284 gnd.n1283 0.152939
R14124 gnd.n1285 gnd.n1284 0.152939
R14125 gnd.n1286 gnd.n1285 0.152939
R14126 gnd.n1305 gnd.n1286 0.152939
R14127 gnd.n1306 gnd.n1305 0.152939
R14128 gnd.n1307 gnd.n1306 0.152939
R14129 gnd.n1308 gnd.n1307 0.152939
R14130 gnd.n1325 gnd.n1308 0.152939
R14131 gnd.n4894 gnd.n1325 0.152939
R14132 gnd.n5053 gnd.n1056 0.152939
R14133 gnd.n5053 gnd.n5052 0.152939
R14134 gnd.n5052 gnd.n5051 0.152939
R14135 gnd.n5051 gnd.n1059 0.152939
R14136 gnd.n3062 gnd.n1059 0.152939
R14137 gnd.n3066 gnd.n3062 0.152939
R14138 gnd.n3067 gnd.n3066 0.152939
R14139 gnd.n3068 gnd.n3067 0.152939
R14140 gnd.n3068 gnd.n3060 0.152939
R14141 gnd.n3074 gnd.n3060 0.152939
R14142 gnd.n3075 gnd.n3074 0.152939
R14143 gnd.n3076 gnd.n3075 0.152939
R14144 gnd.n3076 gnd.n2948 0.152939
R14145 gnd.n3090 gnd.n2948 0.152939
R14146 gnd.n3091 gnd.n3090 0.152939
R14147 gnd.n3092 gnd.n3091 0.152939
R14148 gnd.n3092 gnd.n2849 0.152939
R14149 gnd.n3106 gnd.n2849 0.152939
R14150 gnd.n3107 gnd.n3106 0.152939
R14151 gnd.n3108 gnd.n3107 0.152939
R14152 gnd.n3108 gnd.n2842 0.152939
R14153 gnd.n3122 gnd.n2842 0.152939
R14154 gnd.n3123 gnd.n3122 0.152939
R14155 gnd.n3124 gnd.n3123 0.152939
R14156 gnd.n3124 gnd.n2835 0.152939
R14157 gnd.n3139 gnd.n2835 0.152939
R14158 gnd.n3142 gnd.n3141 0.152939
R14159 gnd.n3142 gnd.n2827 0.152939
R14160 gnd.n3156 gnd.n2827 0.152939
R14161 gnd.n3157 gnd.n3156 0.152939
R14162 gnd.n3158 gnd.n3157 0.152939
R14163 gnd.n3158 gnd.n2820 0.152939
R14164 gnd.n3172 gnd.n2820 0.152939
R14165 gnd.n3173 gnd.n3172 0.152939
R14166 gnd.n3174 gnd.n3173 0.152939
R14167 gnd.n3174 gnd.n2813 0.152939
R14168 gnd.n3188 gnd.n2813 0.152939
R14169 gnd.n3189 gnd.n3188 0.152939
R14170 gnd.n3191 gnd.n3189 0.152939
R14171 gnd.n3191 gnd.n3190 0.152939
R14172 gnd.n3190 gnd.n2807 0.152939
R14173 gnd.n2807 gnd.n2805 0.152939
R14174 gnd.n3207 gnd.n2805 0.152939
R14175 gnd.n3208 gnd.n3207 0.152939
R14176 gnd.n3209 gnd.n3208 0.152939
R14177 gnd.n3209 gnd.n2803 0.152939
R14178 gnd.n3217 gnd.n2803 0.152939
R14179 gnd.n3218 gnd.n3217 0.152939
R14180 gnd.n3220 gnd.n3218 0.152939
R14181 gnd.n3220 gnd.n3219 0.152939
R14182 gnd.n3219 gnd.n2699 0.152939
R14183 gnd.n3532 gnd.n2699 0.152939
R14184 gnd.n1014 gnd.n1013 0.152939
R14185 gnd.n1015 gnd.n1014 0.152939
R14186 gnd.n1016 gnd.n1015 0.152939
R14187 gnd.n1017 gnd.n1016 0.152939
R14188 gnd.n1018 gnd.n1017 0.152939
R14189 gnd.n1019 gnd.n1018 0.152939
R14190 gnd.n1020 gnd.n1019 0.152939
R14191 gnd.n1021 gnd.n1020 0.152939
R14192 gnd.n1022 gnd.n1021 0.152939
R14193 gnd.n1023 gnd.n1022 0.152939
R14194 gnd.n1024 gnd.n1023 0.152939
R14195 gnd.n1025 gnd.n1024 0.152939
R14196 gnd.n1026 gnd.n1025 0.152939
R14197 gnd.n1027 gnd.n1026 0.152939
R14198 gnd.n1028 gnd.n1027 0.152939
R14199 gnd.n1029 gnd.n1028 0.152939
R14200 gnd.n1030 gnd.n1029 0.152939
R14201 gnd.n1033 gnd.n1030 0.152939
R14202 gnd.n1034 gnd.n1033 0.152939
R14203 gnd.n1035 gnd.n1034 0.152939
R14204 gnd.n1036 gnd.n1035 0.152939
R14205 gnd.n1037 gnd.n1036 0.152939
R14206 gnd.n1038 gnd.n1037 0.152939
R14207 gnd.n1039 gnd.n1038 0.152939
R14208 gnd.n1040 gnd.n1039 0.152939
R14209 gnd.n1041 gnd.n1040 0.152939
R14210 gnd.n1042 gnd.n1041 0.152939
R14211 gnd.n1043 gnd.n1042 0.152939
R14212 gnd.n1044 gnd.n1043 0.152939
R14213 gnd.n1045 gnd.n1044 0.152939
R14214 gnd.n1046 gnd.n1045 0.152939
R14215 gnd.n1047 gnd.n1046 0.152939
R14216 gnd.n1048 gnd.n1047 0.152939
R14217 gnd.n1049 gnd.n1048 0.152939
R14218 gnd.n1050 gnd.n1049 0.152939
R14219 gnd.n5061 gnd.n1050 0.152939
R14220 gnd.n5061 gnd.n5060 0.152939
R14221 gnd.n5060 gnd.n5059 0.152939
R14222 gnd.n3035 gnd.n3033 0.152939
R14223 gnd.n3035 gnd.n3034 0.152939
R14224 gnd.n3034 gnd.n1070 0.152939
R14225 gnd.n1071 gnd.n1070 0.152939
R14226 gnd.n1072 gnd.n1071 0.152939
R14227 gnd.n1090 gnd.n1072 0.152939
R14228 gnd.n1091 gnd.n1090 0.152939
R14229 gnd.n1092 gnd.n1091 0.152939
R14230 gnd.n1093 gnd.n1092 0.152939
R14231 gnd.n1110 gnd.n1093 0.152939
R14232 gnd.n1111 gnd.n1110 0.152939
R14233 gnd.n1112 gnd.n1111 0.152939
R14234 gnd.n1113 gnd.n1112 0.152939
R14235 gnd.n1132 gnd.n1113 0.152939
R14236 gnd.n1133 gnd.n1132 0.152939
R14237 gnd.n1134 gnd.n1133 0.152939
R14238 gnd.n1135 gnd.n1134 0.152939
R14239 gnd.n1152 gnd.n1135 0.152939
R14240 gnd.n1153 gnd.n1152 0.152939
R14241 gnd.n1154 gnd.n1153 0.152939
R14242 gnd.n1155 gnd.n1154 0.152939
R14243 gnd.n2863 gnd.n2862 0.152939
R14244 gnd.n2863 gnd.n2854 0.152939
R14245 gnd.n2869 gnd.n2854 0.152939
R14246 gnd.n2870 gnd.n2869 0.152939
R14247 gnd.n2871 gnd.n2870 0.152939
R14248 gnd.n2872 gnd.n2871 0.152939
R14249 gnd.n2873 gnd.n2872 0.152939
R14250 gnd.n2932 gnd.n2873 0.152939
R14251 gnd.n743 gnd.n742 0.152939
R14252 gnd.n744 gnd.n743 0.152939
R14253 gnd.n749 gnd.n744 0.152939
R14254 gnd.n750 gnd.n749 0.152939
R14255 gnd.n751 gnd.n750 0.152939
R14256 gnd.n752 gnd.n751 0.152939
R14257 gnd.n757 gnd.n752 0.152939
R14258 gnd.n758 gnd.n757 0.152939
R14259 gnd.n759 gnd.n758 0.152939
R14260 gnd.n760 gnd.n759 0.152939
R14261 gnd.n765 gnd.n760 0.152939
R14262 gnd.n766 gnd.n765 0.152939
R14263 gnd.n767 gnd.n766 0.152939
R14264 gnd.n768 gnd.n767 0.152939
R14265 gnd.n773 gnd.n768 0.152939
R14266 gnd.n774 gnd.n773 0.152939
R14267 gnd.n775 gnd.n774 0.152939
R14268 gnd.n776 gnd.n775 0.152939
R14269 gnd.n781 gnd.n776 0.152939
R14270 gnd.n782 gnd.n781 0.152939
R14271 gnd.n783 gnd.n782 0.152939
R14272 gnd.n784 gnd.n783 0.152939
R14273 gnd.n789 gnd.n784 0.152939
R14274 gnd.n790 gnd.n789 0.152939
R14275 gnd.n791 gnd.n790 0.152939
R14276 gnd.n792 gnd.n791 0.152939
R14277 gnd.n797 gnd.n792 0.152939
R14278 gnd.n798 gnd.n797 0.152939
R14279 gnd.n799 gnd.n798 0.152939
R14280 gnd.n800 gnd.n799 0.152939
R14281 gnd.n805 gnd.n800 0.152939
R14282 gnd.n806 gnd.n805 0.152939
R14283 gnd.n807 gnd.n806 0.152939
R14284 gnd.n808 gnd.n807 0.152939
R14285 gnd.n813 gnd.n808 0.152939
R14286 gnd.n814 gnd.n813 0.152939
R14287 gnd.n815 gnd.n814 0.152939
R14288 gnd.n816 gnd.n815 0.152939
R14289 gnd.n821 gnd.n816 0.152939
R14290 gnd.n822 gnd.n821 0.152939
R14291 gnd.n823 gnd.n822 0.152939
R14292 gnd.n824 gnd.n823 0.152939
R14293 gnd.n829 gnd.n824 0.152939
R14294 gnd.n830 gnd.n829 0.152939
R14295 gnd.n831 gnd.n830 0.152939
R14296 gnd.n832 gnd.n831 0.152939
R14297 gnd.n837 gnd.n832 0.152939
R14298 gnd.n838 gnd.n837 0.152939
R14299 gnd.n839 gnd.n838 0.152939
R14300 gnd.n840 gnd.n839 0.152939
R14301 gnd.n845 gnd.n840 0.152939
R14302 gnd.n846 gnd.n845 0.152939
R14303 gnd.n847 gnd.n846 0.152939
R14304 gnd.n848 gnd.n847 0.152939
R14305 gnd.n853 gnd.n848 0.152939
R14306 gnd.n854 gnd.n853 0.152939
R14307 gnd.n855 gnd.n854 0.152939
R14308 gnd.n856 gnd.n855 0.152939
R14309 gnd.n861 gnd.n856 0.152939
R14310 gnd.n862 gnd.n861 0.152939
R14311 gnd.n863 gnd.n862 0.152939
R14312 gnd.n864 gnd.n863 0.152939
R14313 gnd.n869 gnd.n864 0.152939
R14314 gnd.n870 gnd.n869 0.152939
R14315 gnd.n871 gnd.n870 0.152939
R14316 gnd.n872 gnd.n871 0.152939
R14317 gnd.n877 gnd.n872 0.152939
R14318 gnd.n878 gnd.n877 0.152939
R14319 gnd.n879 gnd.n878 0.152939
R14320 gnd.n880 gnd.n879 0.152939
R14321 gnd.n885 gnd.n880 0.152939
R14322 gnd.n886 gnd.n885 0.152939
R14323 gnd.n887 gnd.n886 0.152939
R14324 gnd.n888 gnd.n887 0.152939
R14325 gnd.n893 gnd.n888 0.152939
R14326 gnd.n894 gnd.n893 0.152939
R14327 gnd.n895 gnd.n894 0.152939
R14328 gnd.n896 gnd.n895 0.152939
R14329 gnd.n901 gnd.n896 0.152939
R14330 gnd.n902 gnd.n901 0.152939
R14331 gnd.n903 gnd.n902 0.152939
R14332 gnd.n904 gnd.n903 0.152939
R14333 gnd.n2858 gnd.n904 0.152939
R14334 gnd.n2861 gnd.n2858 0.152939
R14335 gnd.n4468 gnd.n4467 0.152939
R14336 gnd.n4467 gnd.n4466 0.152939
R14337 gnd.n4466 gnd.n1780 0.152939
R14338 gnd.n4462 gnd.n1780 0.152939
R14339 gnd.n4462 gnd.n4461 0.152939
R14340 gnd.n4461 gnd.n4460 0.152939
R14341 gnd.n4460 gnd.n1788 0.152939
R14342 gnd.n4456 gnd.n1788 0.152939
R14343 gnd.n4456 gnd.n4455 0.152939
R14344 gnd.n3505 gnd.n2724 0.152939
R14345 gnd.n3501 gnd.n2724 0.152939
R14346 gnd.n3501 gnd.n3500 0.152939
R14347 gnd.n3500 gnd.n3499 0.152939
R14348 gnd.n3499 gnd.n2729 0.152939
R14349 gnd.n3495 gnd.n2729 0.152939
R14350 gnd.n3495 gnd.n3494 0.152939
R14351 gnd.n3494 gnd.n3493 0.152939
R14352 gnd.n3493 gnd.n2734 0.152939
R14353 gnd.n3489 gnd.n2734 0.152939
R14354 gnd.n3489 gnd.n3488 0.152939
R14355 gnd.n3488 gnd.n3487 0.152939
R14356 gnd.n3487 gnd.n2739 0.152939
R14357 gnd.n3483 gnd.n2739 0.152939
R14358 gnd.n3483 gnd.n3482 0.152939
R14359 gnd.n3482 gnd.n3481 0.152939
R14360 gnd.n3481 gnd.n2744 0.152939
R14361 gnd.n3477 gnd.n2744 0.152939
R14362 gnd.n3477 gnd.n3476 0.152939
R14363 gnd.n3476 gnd.n2383 0.152939
R14364 gnd.n3667 gnd.n2383 0.152939
R14365 gnd.n3668 gnd.n3667 0.152939
R14366 gnd.n3669 gnd.n3668 0.152939
R14367 gnd.n3669 gnd.n2363 0.152939
R14368 gnd.n3697 gnd.n2363 0.152939
R14369 gnd.n3698 gnd.n3697 0.152939
R14370 gnd.n3700 gnd.n3698 0.152939
R14371 gnd.n3700 gnd.n3699 0.152939
R14372 gnd.n3699 gnd.n2336 0.152939
R14373 gnd.n3734 gnd.n2336 0.152939
R14374 gnd.n3735 gnd.n3734 0.152939
R14375 gnd.n3736 gnd.n3735 0.152939
R14376 gnd.n3736 gnd.n2316 0.152939
R14377 gnd.n3761 gnd.n2316 0.152939
R14378 gnd.n3762 gnd.n3761 0.152939
R14379 gnd.n3764 gnd.n3762 0.152939
R14380 gnd.n3764 gnd.n3763 0.152939
R14381 gnd.n3763 gnd.n2286 0.152939
R14382 gnd.n3800 gnd.n2286 0.152939
R14383 gnd.n3801 gnd.n3800 0.152939
R14384 gnd.n3816 gnd.n3801 0.152939
R14385 gnd.n3816 gnd.n3815 0.152939
R14386 gnd.n3815 gnd.n3814 0.152939
R14387 gnd.n3814 gnd.n3802 0.152939
R14388 gnd.n3810 gnd.n3802 0.152939
R14389 gnd.n3810 gnd.n3809 0.152939
R14390 gnd.n3809 gnd.n2224 0.152939
R14391 gnd.n3882 gnd.n2224 0.152939
R14392 gnd.n3883 gnd.n3882 0.152939
R14393 gnd.n3885 gnd.n3883 0.152939
R14394 gnd.n3885 gnd.n3884 0.152939
R14395 gnd.n3884 gnd.n2194 0.152939
R14396 gnd.n3918 gnd.n2194 0.152939
R14397 gnd.n3919 gnd.n3918 0.152939
R14398 gnd.n3933 gnd.n3919 0.152939
R14399 gnd.n3933 gnd.n3932 0.152939
R14400 gnd.n3932 gnd.n3931 0.152939
R14401 gnd.n3931 gnd.n3920 0.152939
R14402 gnd.n3927 gnd.n3920 0.152939
R14403 gnd.n3927 gnd.n3926 0.152939
R14404 gnd.n3926 gnd.n2145 0.152939
R14405 gnd.n4012 gnd.n2145 0.152939
R14406 gnd.n4013 gnd.n4012 0.152939
R14407 gnd.n4029 gnd.n4013 0.152939
R14408 gnd.n4029 gnd.n4028 0.152939
R14409 gnd.n4028 gnd.n4027 0.152939
R14410 gnd.n4027 gnd.n4014 0.152939
R14411 gnd.n4023 gnd.n4014 0.152939
R14412 gnd.n4023 gnd.n4022 0.152939
R14413 gnd.n4022 gnd.n2096 0.152939
R14414 gnd.n4101 gnd.n2096 0.152939
R14415 gnd.n4102 gnd.n4101 0.152939
R14416 gnd.n4107 gnd.n4102 0.152939
R14417 gnd.n4107 gnd.n4106 0.152939
R14418 gnd.n4106 gnd.n4105 0.152939
R14419 gnd.n4105 gnd.n2065 0.152939
R14420 gnd.n4169 gnd.n2065 0.152939
R14421 gnd.n4170 gnd.n4169 0.152939
R14422 gnd.n4178 gnd.n4170 0.152939
R14423 gnd.n4178 gnd.n4177 0.152939
R14424 gnd.n4177 gnd.n4176 0.152939
R14425 gnd.n4176 gnd.n4171 0.152939
R14426 gnd.n4171 gnd.n1849 0.152939
R14427 gnd.n4370 gnd.n1849 0.152939
R14428 gnd.n4371 gnd.n4370 0.152939
R14429 gnd.n4372 gnd.n4371 0.152939
R14430 gnd.n4372 gnd.n1837 0.152939
R14431 gnd.n4390 gnd.n1837 0.152939
R14432 gnd.n4391 gnd.n4390 0.152939
R14433 gnd.n4392 gnd.n4391 0.152939
R14434 gnd.n4392 gnd.n1824 0.152939
R14435 gnd.n4410 gnd.n1824 0.152939
R14436 gnd.n4411 gnd.n4410 0.152939
R14437 gnd.n4412 gnd.n4411 0.152939
R14438 gnd.n4412 gnd.n1811 0.152939
R14439 gnd.n4430 gnd.n1811 0.152939
R14440 gnd.n4431 gnd.n4430 0.152939
R14441 gnd.n4433 gnd.n4431 0.152939
R14442 gnd.n4433 gnd.n4432 0.152939
R14443 gnd.n4432 gnd.n1800 0.152939
R14444 gnd.n4454 gnd.n1800 0.152939
R14445 gnd.n3518 gnd.n2705 0.152939
R14446 gnd.n3518 gnd.n3517 0.152939
R14447 gnd.n3517 gnd.n3516 0.152939
R14448 gnd.n3516 gnd.n2712 0.152939
R14449 gnd.n3512 gnd.n2712 0.152939
R14450 gnd.n3512 gnd.n3511 0.152939
R14451 gnd.n3511 gnd.n2719 0.152939
R14452 gnd.n3507 gnd.n2719 0.152939
R14453 gnd.n3507 gnd.n3506 0.152939
R14454 gnd.n3148 gnd.n2830 0.152939
R14455 gnd.n3149 gnd.n3148 0.152939
R14456 gnd.n3150 gnd.n3149 0.152939
R14457 gnd.n3150 gnd.n2824 0.152939
R14458 gnd.n3164 gnd.n2824 0.152939
R14459 gnd.n3165 gnd.n3164 0.152939
R14460 gnd.n3166 gnd.n3165 0.152939
R14461 gnd.n3166 gnd.n2816 0.152939
R14462 gnd.n3180 gnd.n2816 0.152939
R14463 gnd.n3181 gnd.n3180 0.152939
R14464 gnd.n3182 gnd.n3181 0.152939
R14465 gnd.n3182 gnd.n2810 0.152939
R14466 gnd.n3197 gnd.n2810 0.152939
R14467 gnd.n3198 gnd.n3197 0.152939
R14468 gnd.n3199 gnd.n3198 0.152939
R14469 gnd.n3199 gnd.n2797 0.152939
R14470 gnd.n3234 gnd.n2797 0.152939
R14471 gnd.n3234 gnd.n3233 0.152939
R14472 gnd.n3233 gnd.n3232 0.152939
R14473 gnd.n3232 gnd.n2798 0.152939
R14474 gnd.n3228 gnd.n2798 0.152939
R14475 gnd.n3228 gnd.n3227 0.152939
R14476 gnd.n3227 gnd.n3226 0.152939
R14477 gnd.n3226 gnd.n2704 0.152939
R14478 gnd.n3525 gnd.n2704 0.152939
R14479 gnd.n3525 gnd.n3524 0.152939
R14480 gnd.n4891 gnd.n1328 0.152939
R14481 gnd.n4887 gnd.n1328 0.152939
R14482 gnd.n4887 gnd.n4886 0.152939
R14483 gnd.n4886 gnd.n4885 0.152939
R14484 gnd.n4885 gnd.n1333 0.152939
R14485 gnd.n4881 gnd.n1333 0.152939
R14486 gnd.n4881 gnd.n4880 0.152939
R14487 gnd.n4880 gnd.n4879 0.152939
R14488 gnd.n4879 gnd.n1338 0.152939
R14489 gnd.n4875 gnd.n1338 0.152939
R14490 gnd.n4875 gnd.n4874 0.152939
R14491 gnd.n4874 gnd.n4873 0.152939
R14492 gnd.n4873 gnd.n1343 0.152939
R14493 gnd.n4869 gnd.n1343 0.152939
R14494 gnd.n4869 gnd.n4868 0.152939
R14495 gnd.n4868 gnd.n4867 0.152939
R14496 gnd.n4867 gnd.n1348 0.152939
R14497 gnd.n4863 gnd.n1348 0.152939
R14498 gnd.n4863 gnd.n4862 0.152939
R14499 gnd.n4862 gnd.n4861 0.152939
R14500 gnd.n4861 gnd.n1353 0.152939
R14501 gnd.n4857 gnd.n1353 0.152939
R14502 gnd.n4857 gnd.n4856 0.152939
R14503 gnd.n4856 gnd.n4855 0.152939
R14504 gnd.n4855 gnd.n1358 0.152939
R14505 gnd.n4851 gnd.n1358 0.152939
R14506 gnd.n4851 gnd.n4850 0.152939
R14507 gnd.n4850 gnd.n4849 0.152939
R14508 gnd.n4849 gnd.n1363 0.152939
R14509 gnd.n4845 gnd.n1363 0.152939
R14510 gnd.n4845 gnd.n4844 0.152939
R14511 gnd.n4844 gnd.n4843 0.152939
R14512 gnd.n4843 gnd.n1368 0.152939
R14513 gnd.n4839 gnd.n1368 0.152939
R14514 gnd.n4839 gnd.n4838 0.152939
R14515 gnd.n4838 gnd.n4837 0.152939
R14516 gnd.n4837 gnd.n1373 0.152939
R14517 gnd.n4833 gnd.n1373 0.152939
R14518 gnd.n4833 gnd.n4832 0.152939
R14519 gnd.n4832 gnd.n4831 0.152939
R14520 gnd.n4831 gnd.n1378 0.152939
R14521 gnd.n4827 gnd.n1378 0.152939
R14522 gnd.n4827 gnd.n4826 0.152939
R14523 gnd.n4826 gnd.n4825 0.152939
R14524 gnd.n4825 gnd.n1383 0.152939
R14525 gnd.n4821 gnd.n1383 0.152939
R14526 gnd.n4821 gnd.n4820 0.152939
R14527 gnd.n4820 gnd.n4819 0.152939
R14528 gnd.n4819 gnd.n1388 0.152939
R14529 gnd.n4815 gnd.n1388 0.152939
R14530 gnd.n4815 gnd.n4814 0.152939
R14531 gnd.n4814 gnd.n4813 0.152939
R14532 gnd.n4813 gnd.n1393 0.152939
R14533 gnd.n4809 gnd.n1393 0.152939
R14534 gnd.n4809 gnd.n4808 0.152939
R14535 gnd.n4808 gnd.n4807 0.152939
R14536 gnd.n4807 gnd.n1398 0.152939
R14537 gnd.n4803 gnd.n1398 0.152939
R14538 gnd.n4803 gnd.n4802 0.152939
R14539 gnd.n4802 gnd.n4801 0.152939
R14540 gnd.n4801 gnd.n1403 0.152939
R14541 gnd.n4797 gnd.n1403 0.152939
R14542 gnd.n4797 gnd.n4796 0.152939
R14543 gnd.n4796 gnd.n4795 0.152939
R14544 gnd.n4795 gnd.n1408 0.152939
R14545 gnd.n4791 gnd.n1408 0.152939
R14546 gnd.n4791 gnd.n4790 0.152939
R14547 gnd.n4790 gnd.n4789 0.152939
R14548 gnd.n4789 gnd.n1413 0.152939
R14549 gnd.n4785 gnd.n1413 0.152939
R14550 gnd.n4785 gnd.n4784 0.152939
R14551 gnd.n4784 gnd.n4783 0.152939
R14552 gnd.n4783 gnd.n1418 0.152939
R14553 gnd.n4779 gnd.n1418 0.152939
R14554 gnd.n4779 gnd.n4778 0.152939
R14555 gnd.n4778 gnd.n4777 0.152939
R14556 gnd.n4777 gnd.n1423 0.152939
R14557 gnd.n4773 gnd.n1423 0.152939
R14558 gnd.n4773 gnd.n4772 0.152939
R14559 gnd.n4772 gnd.n4771 0.152939
R14560 gnd.n4771 gnd.n1428 0.152939
R14561 gnd.n4767 gnd.n1428 0.152939
R14562 gnd.n4767 gnd.n4766 0.152939
R14563 gnd.n4766 gnd.n4765 0.152939
R14564 gnd.n4765 gnd.n1433 0.152939
R14565 gnd.n4761 gnd.n1433 0.152939
R14566 gnd.n4761 gnd.n4760 0.152939
R14567 gnd.n4760 gnd.n4759 0.152939
R14568 gnd.n4759 gnd.n1438 0.152939
R14569 gnd.n4755 gnd.n1438 0.152939
R14570 gnd.n4755 gnd.n4754 0.152939
R14571 gnd.n4754 gnd.n4753 0.152939
R14572 gnd.n4753 gnd.n1443 0.152939
R14573 gnd.n4749 gnd.n1443 0.152939
R14574 gnd.n4749 gnd.n4748 0.152939
R14575 gnd.n4748 gnd.n4747 0.152939
R14576 gnd.n4747 gnd.n1448 0.152939
R14577 gnd.n4743 gnd.n1448 0.152939
R14578 gnd.n4743 gnd.n4742 0.152939
R14579 gnd.n4742 gnd.n4741 0.152939
R14580 gnd.n4741 gnd.n1453 0.152939
R14581 gnd.n1691 gnd.n1685 0.152939
R14582 gnd.n1685 gnd.n1498 0.152939
R14583 gnd.n4712 gnd.n1498 0.152939
R14584 gnd.n4712 gnd.n4711 0.152939
R14585 gnd.n4711 gnd.n4710 0.152939
R14586 gnd.n4710 gnd.n1499 0.152939
R14587 gnd.n4706 gnd.n1499 0.152939
R14588 gnd.n4706 gnd.n4705 0.152939
R14589 gnd.n4705 gnd.n4704 0.152939
R14590 gnd.n4704 gnd.n1504 0.152939
R14591 gnd.n4700 gnd.n1504 0.152939
R14592 gnd.n4700 gnd.n4699 0.152939
R14593 gnd.n4699 gnd.n4698 0.152939
R14594 gnd.n4698 gnd.n1509 0.152939
R14595 gnd.n4694 gnd.n1509 0.152939
R14596 gnd.n4694 gnd.n4693 0.152939
R14597 gnd.n4693 gnd.n4692 0.152939
R14598 gnd.n4692 gnd.n1514 0.152939
R14599 gnd.n4688 gnd.n1514 0.152939
R14600 gnd.n4688 gnd.n4687 0.152939
R14601 gnd.n4687 gnd.n285 0.152939
R14602 gnd.n7495 gnd.n285 0.152939
R14603 gnd.n7495 gnd.n7494 0.152939
R14604 gnd.n7494 gnd.n7493 0.152939
R14605 gnd.n7493 gnd.n286 0.152939
R14606 gnd.n7489 gnd.n286 0.152939
R14607 gnd.n7487 gnd.n7486 0.152939
R14608 gnd.n7486 gnd.n292 0.152939
R14609 gnd.n292 gnd.n260 0.152939
R14610 gnd.n7508 gnd.n260 0.152939
R14611 gnd.n7509 gnd.n7508 0.152939
R14612 gnd.n7510 gnd.n7509 0.152939
R14613 gnd.n7510 gnd.n244 0.152939
R14614 gnd.n7524 gnd.n244 0.152939
R14615 gnd.n7525 gnd.n7524 0.152939
R14616 gnd.n7526 gnd.n7525 0.152939
R14617 gnd.n7526 gnd.n229 0.152939
R14618 gnd.n7540 gnd.n229 0.152939
R14619 gnd.n7541 gnd.n7540 0.152939
R14620 gnd.n7542 gnd.n7541 0.152939
R14621 gnd.n7542 gnd.n214 0.152939
R14622 gnd.n7556 gnd.n214 0.152939
R14623 gnd.n7557 gnd.n7556 0.152939
R14624 gnd.n7558 gnd.n7557 0.152939
R14625 gnd.n7558 gnd.n199 0.152939
R14626 gnd.n7572 gnd.n199 0.152939
R14627 gnd.n7573 gnd.n7572 0.152939
R14628 gnd.n7649 gnd.n7573 0.152939
R14629 gnd.n7649 gnd.n7648 0.152939
R14630 gnd.n7648 gnd.n7647 0.152939
R14631 gnd.n7647 gnd.n7574 0.152939
R14632 gnd.n7643 gnd.n7574 0.152939
R14633 gnd.n7642 gnd.n7576 0.152939
R14634 gnd.n7638 gnd.n7576 0.152939
R14635 gnd.n7638 gnd.n7637 0.152939
R14636 gnd.n7637 gnd.n7636 0.152939
R14637 gnd.n7636 gnd.n7582 0.152939
R14638 gnd.n7632 gnd.n7582 0.152939
R14639 gnd.n7632 gnd.n7631 0.152939
R14640 gnd.n7631 gnd.n7630 0.152939
R14641 gnd.n7630 gnd.n7590 0.152939
R14642 gnd.n7626 gnd.n7590 0.152939
R14643 gnd.n7626 gnd.n7625 0.152939
R14644 gnd.n7625 gnd.n7624 0.152939
R14645 gnd.n7624 gnd.n7598 0.152939
R14646 gnd.n7620 gnd.n7598 0.152939
R14647 gnd.n7620 gnd.n7619 0.152939
R14648 gnd.n7619 gnd.n7618 0.152939
R14649 gnd.n7618 gnd.n7606 0.152939
R14650 gnd.n7614 gnd.n7606 0.152939
R14651 gnd.n4479 gnd.n4478 0.152939
R14652 gnd.n4481 gnd.n4479 0.152939
R14653 gnd.n4481 gnd.n4480 0.152939
R14654 gnd.n4480 gnd.n1621 0.152939
R14655 gnd.n4528 gnd.n1621 0.152939
R14656 gnd.n4529 gnd.n4528 0.152939
R14657 gnd.n4531 gnd.n4529 0.152939
R14658 gnd.n4531 gnd.n4530 0.152939
R14659 gnd.n4530 gnd.n1594 0.152939
R14660 gnd.n4560 gnd.n1594 0.152939
R14661 gnd.n4561 gnd.n4560 0.152939
R14662 gnd.n4563 gnd.n4561 0.152939
R14663 gnd.n4563 gnd.n4562 0.152939
R14664 gnd.n4562 gnd.n1565 0.152939
R14665 gnd.n4599 gnd.n1565 0.152939
R14666 gnd.n4600 gnd.n4599 0.152939
R14667 gnd.n4605 gnd.n4600 0.152939
R14668 gnd.n4605 gnd.n4604 0.152939
R14669 gnd.n4604 gnd.n4603 0.152939
R14670 gnd.n4603 gnd.n1554 0.152939
R14671 gnd.n4625 gnd.n1554 0.152939
R14672 gnd.n4626 gnd.n4625 0.152939
R14673 gnd.n4630 gnd.n4626 0.152939
R14674 gnd.n4630 gnd.n4629 0.152939
R14675 gnd.n4629 gnd.n4628 0.152939
R14676 gnd.n4628 gnd.n67 0.152939
R14677 gnd.n7781 gnd.n68 0.152939
R14678 gnd.n7777 gnd.n68 0.152939
R14679 gnd.n7777 gnd.n7776 0.152939
R14680 gnd.n7776 gnd.n7775 0.152939
R14681 gnd.n7775 gnd.n74 0.152939
R14682 gnd.n7771 gnd.n74 0.152939
R14683 gnd.n7771 gnd.n7770 0.152939
R14684 gnd.n7770 gnd.n7769 0.152939
R14685 gnd.n7769 gnd.n79 0.152939
R14686 gnd.n7765 gnd.n79 0.152939
R14687 gnd.n7765 gnd.n7764 0.152939
R14688 gnd.n7764 gnd.n7763 0.152939
R14689 gnd.n7763 gnd.n84 0.152939
R14690 gnd.n7759 gnd.n84 0.152939
R14691 gnd.n7759 gnd.n7758 0.152939
R14692 gnd.n7758 gnd.n7757 0.152939
R14693 gnd.n7757 gnd.n89 0.152939
R14694 gnd.n7753 gnd.n89 0.152939
R14695 gnd.n7753 gnd.n7752 0.152939
R14696 gnd.n7752 gnd.n7751 0.152939
R14697 gnd.n7751 gnd.n94 0.152939
R14698 gnd.n7747 gnd.n94 0.152939
R14699 gnd.n7747 gnd.n7746 0.152939
R14700 gnd.n7746 gnd.n7745 0.152939
R14701 gnd.n7745 gnd.n99 0.152939
R14702 gnd.n102 gnd.n99 0.152939
R14703 gnd.n4468 gnd.n1643 0.151415
R14704 gnd.n3523 gnd.n2705 0.151415
R14705 gnd.n309 gnd.n268 0.0889146
R14706 gnd.n2933 gnd.n2932 0.0889146
R14707 gnd.n5948 gnd.n5340 0.0767195
R14708 gnd.n5864 gnd.n5340 0.0767195
R14709 gnd.n7502 gnd.n252 0.0767195
R14710 gnd.n4640 gnd.n291 0.0767195
R14711 gnd.n300 gnd.n291 0.0767195
R14712 gnd.n7502 gnd.n267 0.0767195
R14713 gnd.n1212 gnd.n1175 0.0767195
R14714 gnd.n2834 gnd.n1184 0.0767195
R14715 gnd.n2834 gnd.n1185 0.0767195
R14716 gnd.n3140 gnd.n3139 0.0767195
R14717 gnd.n3141 gnd.n3140 0.0767195
R14718 gnd.n1175 gnd.n1155 0.0767195
R14719 gnd.n7489 gnd.n7488 0.0767195
R14720 gnd.n7488 gnd.n7487 0.0767195
R14721 gnd.n7782 gnd.n67 0.0767195
R14722 gnd.n7782 gnd.n7781 0.0767195
R14723 gnd.n3133 gnd.n3132 0.0695946
R14724 gnd.n3132 gnd.n2830 0.0695946
R14725 gnd.n2933 gnd.n2877 0.0645244
R14726 gnd.n1536 gnd.n268 0.0645244
R14727 gnd.n4893 gnd.n4892 0.063
R14728 gnd.n1693 gnd.n1692 0.063
R14729 gnd.n6456 gnd.n5160 0.0477147
R14730 gnd.n5614 gnd.n5510 0.0442063
R14731 gnd.n5628 gnd.n5510 0.0442063
R14732 gnd.n5629 gnd.n5628 0.0442063
R14733 gnd.n5630 gnd.n5629 0.0442063
R14734 gnd.n5630 gnd.n5498 0.0442063
R14735 gnd.n5644 gnd.n5498 0.0442063
R14736 gnd.n5645 gnd.n5644 0.0442063
R14737 gnd.n5646 gnd.n5645 0.0442063
R14738 gnd.n5646 gnd.n5485 0.0442063
R14739 gnd.n5742 gnd.n5485 0.0442063
R14740 gnd.n5745 gnd.n5744 0.0344674
R14741 gnd.n4472 gnd.n1649 0.0343753
R14742 gnd.n3522 gnd.n2706 0.0343753
R14743 gnd.n5478 gnd.n5477 0.0269946
R14744 gnd.n5755 gnd.n5475 0.0269946
R14745 gnd.n5754 gnd.n5476 0.0269946
R14746 gnd.n5774 gnd.n5457 0.0269946
R14747 gnd.n5776 gnd.n5775 0.0269946
R14748 gnd.n5777 gnd.n5455 0.0269946
R14749 gnd.n5784 gnd.n5780 0.0269946
R14750 gnd.n5783 gnd.n5782 0.0269946
R14751 gnd.n5781 gnd.n5434 0.0269946
R14752 gnd.n5808 gnd.n5435 0.0269946
R14753 gnd.n5807 gnd.n5436 0.0269946
R14754 gnd.n5840 gnd.n5410 0.0269946
R14755 gnd.n5842 gnd.n5841 0.0269946
R14756 gnd.n5843 gnd.n5402 0.0269946
R14757 gnd.n5406 gnd.n5403 0.0269946
R14758 gnd.n5853 gnd.n5404 0.0269946
R14759 gnd.n5852 gnd.n5405 0.0269946
R14760 gnd.n5898 gnd.n5378 0.0269946
R14761 gnd.n5900 gnd.n5899 0.0269946
R14762 gnd.n5909 gnd.n5371 0.0269946
R14763 gnd.n5911 gnd.n5910 0.0269946
R14764 gnd.n5912 gnd.n5369 0.0269946
R14765 gnd.n5919 gnd.n5915 0.0269946
R14766 gnd.n5918 gnd.n5917 0.0269946
R14767 gnd.n5916 gnd.n5348 0.0269946
R14768 gnd.n5941 gnd.n5349 0.0269946
R14769 gnd.n5940 gnd.n5350 0.0269946
R14770 gnd.n5983 gnd.n5275 0.0269946
R14771 gnd.n5985 gnd.n5984 0.0269946
R14772 gnd.n5994 gnd.n5268 0.0269946
R14773 gnd.n5996 gnd.n5995 0.0269946
R14774 gnd.n5997 gnd.n5266 0.0269946
R14775 gnd.n6003 gnd.n6000 0.0269946
R14776 gnd.n6002 gnd.n6001 0.0269946
R14777 gnd.n6028 gnd.n5245 0.0269946
R14778 gnd.n6027 gnd.n5246 0.0269946
R14779 gnd.n6054 gnd.n5231 0.0269946
R14780 gnd.n6056 gnd.n6055 0.0269946
R14781 gnd.n6057 gnd.n5217 0.0269946
R14782 gnd.n6079 gnd.n5215 0.0269946
R14783 gnd.n6081 gnd.n6080 0.0269946
R14784 gnd.n6083 gnd.n6082 0.0269946
R14785 gnd.n6092 gnd.n5207 0.0269946
R14786 gnd.n6094 gnd.n6093 0.0269946
R14787 gnd.n6095 gnd.n924 0.0269946
R14788 gnd.n5198 gnd.n925 0.0269946
R14789 gnd.n5200 gnd.n926 0.0269946
R14790 gnd.n6122 gnd.n6121 0.0269946
R14791 gnd.n6381 gnd.n949 0.0269946
R14792 gnd.n6383 gnd.n950 0.0269946
R14793 gnd.n6385 gnd.n951 0.0269946
R14794 gnd.n6387 gnd.n6386 0.0269946
R14795 gnd.n1694 gnd.n1693 0.0245515
R14796 gnd.n4892 gnd.n1327 0.0245515
R14797 gnd.n5744 gnd.n5743 0.0202011
R14798 gnd.n1695 gnd.n1694 0.0174377
R14799 gnd.n1703 gnd.n1695 0.0174377
R14800 gnd.n1703 gnd.n1702 0.0174377
R14801 gnd.n1702 gnd.n1696 0.0174377
R14802 gnd.n1696 gnd.n1680 0.0174377
R14803 gnd.n1711 gnd.n1680 0.0174377
R14804 gnd.n1713 gnd.n1711 0.0174377
R14805 gnd.n1713 gnd.n1712 0.0174377
R14806 gnd.n1712 gnd.n1675 0.0174377
R14807 gnd.n1722 gnd.n1675 0.0174377
R14808 gnd.n1722 gnd.n1721 0.0174377
R14809 gnd.n1721 gnd.n1676 0.0174377
R14810 gnd.n1676 gnd.n1671 0.0174377
R14811 gnd.n1730 gnd.n1671 0.0174377
R14812 gnd.n1732 gnd.n1730 0.0174377
R14813 gnd.n1732 gnd.n1731 0.0174377
R14814 gnd.n1731 gnd.n1666 0.0174377
R14815 gnd.n1741 gnd.n1666 0.0174377
R14816 gnd.n1741 gnd.n1740 0.0174377
R14817 gnd.n1740 gnd.n1667 0.0174377
R14818 gnd.n1667 gnd.n1662 0.0174377
R14819 gnd.n1749 gnd.n1662 0.0174377
R14820 gnd.n1751 gnd.n1749 0.0174377
R14821 gnd.n1751 gnd.n1750 0.0174377
R14822 gnd.n1750 gnd.n1657 0.0174377
R14823 gnd.n1760 gnd.n1657 0.0174377
R14824 gnd.n1760 gnd.n1759 0.0174377
R14825 gnd.n1759 gnd.n1658 0.0174377
R14826 gnd.n1658 gnd.n1653 0.0174377
R14827 gnd.n1768 gnd.n1653 0.0174377
R14828 gnd.n1770 gnd.n1768 0.0174377
R14829 gnd.n1770 gnd.n1769 0.0174377
R14830 gnd.n1769 gnd.n1648 0.0174377
R14831 gnd.n4473 gnd.n1648 0.0174377
R14832 gnd.n4473 gnd.n4472 0.0174377
R14833 gnd.n3282 gnd.n1327 0.0174377
R14834 gnd.n3284 gnd.n3282 0.0174377
R14835 gnd.n3392 gnd.n3284 0.0174377
R14836 gnd.n3392 gnd.n3391 0.0174377
R14837 gnd.n3391 gnd.n3285 0.0174377
R14838 gnd.n3388 gnd.n3285 0.0174377
R14839 gnd.n3388 gnd.n3387 0.0174377
R14840 gnd.n3387 gnd.n3295 0.0174377
R14841 gnd.n3384 gnd.n3295 0.0174377
R14842 gnd.n3384 gnd.n3383 0.0174377
R14843 gnd.n3383 gnd.n3300 0.0174377
R14844 gnd.n3380 gnd.n3300 0.0174377
R14845 gnd.n3380 gnd.n3379 0.0174377
R14846 gnd.n3379 gnd.n3306 0.0174377
R14847 gnd.n3376 gnd.n3306 0.0174377
R14848 gnd.n3376 gnd.n3375 0.0174377
R14849 gnd.n3375 gnd.n3310 0.0174377
R14850 gnd.n3372 gnd.n3310 0.0174377
R14851 gnd.n3372 gnd.n3371 0.0174377
R14852 gnd.n3371 gnd.n3317 0.0174377
R14853 gnd.n3368 gnd.n3317 0.0174377
R14854 gnd.n3368 gnd.n3367 0.0174377
R14855 gnd.n3367 gnd.n3323 0.0174377
R14856 gnd.n3364 gnd.n3323 0.0174377
R14857 gnd.n3364 gnd.n3363 0.0174377
R14858 gnd.n3363 gnd.n3329 0.0174377
R14859 gnd.n3360 gnd.n3329 0.0174377
R14860 gnd.n3360 gnd.n3359 0.0174377
R14861 gnd.n3359 gnd.n3333 0.0174377
R14862 gnd.n3356 gnd.n3333 0.0174377
R14863 gnd.n3356 gnd.n3355 0.0174377
R14864 gnd.n3355 gnd.n3342 0.0174377
R14865 gnd.n3352 gnd.n3342 0.0174377
R14866 gnd.n3352 gnd.n3351 0.0174377
R14867 gnd.n3351 gnd.n2706 0.0174377
R14868 gnd.n5743 gnd.n5742 0.0148637
R14869 gnd.n6379 gnd.n6123 0.0144266
R14870 gnd.n6380 gnd.n6379 0.0130679
R14871 gnd.n5745 gnd.n5478 0.00797283
R14872 gnd.n5477 gnd.n5475 0.00797283
R14873 gnd.n5755 gnd.n5754 0.00797283
R14874 gnd.n5476 gnd.n5457 0.00797283
R14875 gnd.n5775 gnd.n5774 0.00797283
R14876 gnd.n5777 gnd.n5776 0.00797283
R14877 gnd.n5780 gnd.n5455 0.00797283
R14878 gnd.n5784 gnd.n5783 0.00797283
R14879 gnd.n5782 gnd.n5781 0.00797283
R14880 gnd.n5435 gnd.n5434 0.00797283
R14881 gnd.n5808 gnd.n5807 0.00797283
R14882 gnd.n5436 gnd.n5410 0.00797283
R14883 gnd.n5841 gnd.n5840 0.00797283
R14884 gnd.n5843 gnd.n5842 0.00797283
R14885 gnd.n5406 gnd.n5402 0.00797283
R14886 gnd.n5404 gnd.n5403 0.00797283
R14887 gnd.n5853 gnd.n5852 0.00797283
R14888 gnd.n5405 gnd.n5378 0.00797283
R14889 gnd.n5900 gnd.n5898 0.00797283
R14890 gnd.n5899 gnd.n5371 0.00797283
R14891 gnd.n5910 gnd.n5909 0.00797283
R14892 gnd.n5912 gnd.n5911 0.00797283
R14893 gnd.n5915 gnd.n5369 0.00797283
R14894 gnd.n5919 gnd.n5918 0.00797283
R14895 gnd.n5917 gnd.n5916 0.00797283
R14896 gnd.n5349 gnd.n5348 0.00797283
R14897 gnd.n5941 gnd.n5940 0.00797283
R14898 gnd.n5350 gnd.n5275 0.00797283
R14899 gnd.n5985 gnd.n5983 0.00797283
R14900 gnd.n5984 gnd.n5268 0.00797283
R14901 gnd.n5995 gnd.n5994 0.00797283
R14902 gnd.n5997 gnd.n5996 0.00797283
R14903 gnd.n6000 gnd.n5266 0.00797283
R14904 gnd.n6003 gnd.n6002 0.00797283
R14905 gnd.n6001 gnd.n5245 0.00797283
R14906 gnd.n6028 gnd.n6027 0.00797283
R14907 gnd.n5246 gnd.n5231 0.00797283
R14908 gnd.n6055 gnd.n6054 0.00797283
R14909 gnd.n6057 gnd.n6056 0.00797283
R14910 gnd.n5217 gnd.n5215 0.00797283
R14911 gnd.n6080 gnd.n6079 0.00797283
R14912 gnd.n6083 gnd.n6081 0.00797283
R14913 gnd.n6082 gnd.n5207 0.00797283
R14914 gnd.n6093 gnd.n6092 0.00797283
R14915 gnd.n6095 gnd.n6094 0.00797283
R14916 gnd.n5198 gnd.n924 0.00797283
R14917 gnd.n5200 gnd.n925 0.00797283
R14918 gnd.n6121 gnd.n926 0.00797283
R14919 gnd.n6123 gnd.n6122 0.00797283
R14920 gnd.n6381 gnd.n6380 0.00797283
R14921 gnd.n6383 gnd.n949 0.00797283
R14922 gnd.n6385 gnd.n950 0.00797283
R14923 gnd.n6387 gnd.n951 0.00797283
R14924 gnd.n6386 gnd.n5160 0.00797283
R14925 gnd.n7488 gnd.n291 0.00507153
R14926 gnd.n3140 gnd.n2834 0.00507153
R14927 gnd.n1649 gnd.n1643 0.000838753
R14928 gnd.n3523 gnd.n3522 0.000838753
R14929 a_n2982_13878.n139 a_n2982_13878.t94 512.366
R14930 a_n2982_13878.n138 a_n2982_13878.t83 512.366
R14931 a_n2982_13878.n137 a_n2982_13878.t72 512.366
R14932 a_n2982_13878.n141 a_n2982_13878.t102 512.366
R14933 a_n2982_13878.n140 a_n2982_13878.t91 512.366
R14934 a_n2982_13878.n136 a_n2982_13878.t90 512.366
R14935 a_n2982_13878.n143 a_n2982_13878.t98 512.366
R14936 a_n2982_13878.n142 a_n2982_13878.t81 512.366
R14937 a_n2982_13878.n135 a_n2982_13878.t82 512.366
R14938 a_n2982_13878.n145 a_n2982_13878.t85 512.366
R14939 a_n2982_13878.n144 a_n2982_13878.t95 512.366
R14940 a_n2982_13878.n134 a_n2982_13878.t111 512.366
R14941 a_n2982_13878.n35 a_n2982_13878.t110 538.698
R14942 a_n2982_13878.n108 a_n2982_13878.t87 512.366
R14943 a_n2982_13878.n107 a_n2982_13878.t92 512.366
R14944 a_n2982_13878.n99 a_n2982_13878.t80 512.366
R14945 a_n2982_13878.n106 a_n2982_13878.t97 512.366
R14946 a_n2982_13878.n105 a_n2982_13878.t106 512.366
R14947 a_n2982_13878.n100 a_n2982_13878.t107 512.366
R14948 a_n2982_13878.n104 a_n2982_13878.t74 512.366
R14949 a_n2982_13878.n103 a_n2982_13878.t89 512.366
R14950 a_n2982_13878.n101 a_n2982_13878.t77 512.366
R14951 a_n2982_13878.n102 a_n2982_13878.t84 512.366
R14952 a_n2982_13878.n29 a_n2982_13878.t41 538.698
R14953 a_n2982_13878.n127 a_n2982_13878.t47 512.366
R14954 a_n2982_13878.n126 a_n2982_13878.t11 512.366
R14955 a_n2982_13878.n97 a_n2982_13878.t9 512.366
R14956 a_n2982_13878.n125 a_n2982_13878.t23 512.366
R14957 a_n2982_13878.n124 a_n2982_13878.t13 512.366
R14958 a_n2982_13878.n98 a_n2982_13878.t35 512.366
R14959 a_n2982_13878.n123 a_n2982_13878.t45 512.366
R14960 a_n2982_13878.n122 a_n2982_13878.t17 512.366
R14961 a_n2982_13878.n83 a_n2982_13878.t43 512.366
R14962 a_n2982_13878.n109 a_n2982_13878.t33 512.366
R14963 a_n2982_13878.n18 a_n2982_13878.t27 538.698
R14964 a_n2982_13878.n153 a_n2982_13878.t29 512.366
R14965 a_n2982_13878.n92 a_n2982_13878.t49 512.366
R14966 a_n2982_13878.n154 a_n2982_13878.t37 512.366
R14967 a_n2982_13878.n91 a_n2982_13878.t7 512.366
R14968 a_n2982_13878.n155 a_n2982_13878.t15 512.366
R14969 a_n2982_13878.n156 a_n2982_13878.t25 512.366
R14970 a_n2982_13878.n90 a_n2982_13878.t19 512.366
R14971 a_n2982_13878.n157 a_n2982_13878.t39 512.366
R14972 a_n2982_13878.n89 a_n2982_13878.t31 512.366
R14973 a_n2982_13878.n158 a_n2982_13878.t51 512.366
R14974 a_n2982_13878.n24 a_n2982_13878.t109 538.698
R14975 a_n2982_13878.n147 a_n2982_13878.t78 512.366
R14976 a_n2982_13878.n96 a_n2982_13878.t79 512.366
R14977 a_n2982_13878.n148 a_n2982_13878.t104 512.366
R14978 a_n2982_13878.n95 a_n2982_13878.t105 512.366
R14979 a_n2982_13878.n149 a_n2982_13878.t76 512.366
R14980 a_n2982_13878.n150 a_n2982_13878.t100 512.366
R14981 a_n2982_13878.n94 a_n2982_13878.t101 512.366
R14982 a_n2982_13878.n151 a_n2982_13878.t73 512.366
R14983 a_n2982_13878.n93 a_n2982_13878.t86 512.366
R14984 a_n2982_13878.n152 a_n2982_13878.t96 512.366
R14985 a_n2982_13878.n5 a_n2982_13878.n82 70.1674
R14986 a_n2982_13878.n7 a_n2982_13878.n80 70.1674
R14987 a_n2982_13878.n9 a_n2982_13878.n78 70.1674
R14988 a_n2982_13878.n11 a_n2982_13878.n76 70.1674
R14989 a_n2982_13878.n52 a_n2982_13878.n30 70.5844
R14990 a_n2982_13878.n37 a_n2982_13878.n36 44.7878
R14991 a_n2982_13878.n37 a_n2982_13878.n109 14.1664
R14992 a_n2982_13878.n30 a_n2982_13878.n50 70.1674
R14993 a_n2982_13878.n50 a_n2982_13878.n101 20.9683
R14994 a_n2982_13878.n49 a_n2982_13878.n31 74.73
R14995 a_n2982_13878.n103 a_n2982_13878.n49 11.843
R14996 a_n2982_13878.n48 a_n2982_13878.n31 80.4688
R14997 a_n2982_13878.n48 a_n2982_13878.n104 0.365327
R14998 a_n2982_13878.n32 a_n2982_13878.n47 75.0448
R14999 a_n2982_13878.n46 a_n2982_13878.n32 70.1674
R15000 a_n2982_13878.n106 a_n2982_13878.n46 20.9683
R15001 a_n2982_13878.n34 a_n2982_13878.n45 70.3058
R15002 a_n2982_13878.n45 a_n2982_13878.n99 20.6913
R15003 a_n2982_13878.n44 a_n2982_13878.n34 75.3623
R15004 a_n2982_13878.n107 a_n2982_13878.n44 10.5784
R15005 a_n2982_13878.n33 a_n2982_13878.n35 44.7878
R15006 a_n2982_13878.n58 a_n2982_13878.n36 44.5605
R15007 a_n2982_13878.n122 a_n2982_13878.n58 21.3688
R15008 a_n2982_13878.n57 a_n2982_13878.n25 80.4688
R15009 a_n2982_13878.n57 a_n2982_13878.n123 0.365327
R15010 a_n2982_13878.n26 a_n2982_13878.n56 75.0448
R15011 a_n2982_13878.n55 a_n2982_13878.n26 70.1674
R15012 a_n2982_13878.n125 a_n2982_13878.n55 20.9683
R15013 a_n2982_13878.n28 a_n2982_13878.n54 70.3058
R15014 a_n2982_13878.n54 a_n2982_13878.n97 20.6913
R15015 a_n2982_13878.n53 a_n2982_13878.n28 75.3623
R15016 a_n2982_13878.n126 a_n2982_13878.n53 10.5784
R15017 a_n2982_13878.n27 a_n2982_13878.n29 44.7878
R15018 a_n2982_13878.n14 a_n2982_13878.n74 70.5844
R15019 a_n2982_13878.n20 a_n2982_13878.n66 70.5844
R15020 a_n2982_13878.n65 a_n2982_13878.n20 70.1674
R15021 a_n2982_13878.n65 a_n2982_13878.n93 20.9683
R15022 a_n2982_13878.n19 a_n2982_13878.n64 74.73
R15023 a_n2982_13878.n151 a_n2982_13878.n64 11.843
R15024 a_n2982_13878.n63 a_n2982_13878.n19 80.4688
R15025 a_n2982_13878.n63 a_n2982_13878.n94 0.365327
R15026 a_n2982_13878.n21 a_n2982_13878.n62 75.0448
R15027 a_n2982_13878.n61 a_n2982_13878.n21 70.1674
R15028 a_n2982_13878.n61 a_n2982_13878.n95 20.9683
R15029 a_n2982_13878.n22 a_n2982_13878.n60 70.3058
R15030 a_n2982_13878.n148 a_n2982_13878.n60 20.6913
R15031 a_n2982_13878.n59 a_n2982_13878.n22 75.3623
R15032 a_n2982_13878.n59 a_n2982_13878.n96 10.5784
R15033 a_n2982_13878.n24 a_n2982_13878.n23 44.7878
R15034 a_n2982_13878.n73 a_n2982_13878.n14 70.1674
R15035 a_n2982_13878.n73 a_n2982_13878.n89 20.9683
R15036 a_n2982_13878.n13 a_n2982_13878.n72 74.73
R15037 a_n2982_13878.n157 a_n2982_13878.n72 11.843
R15038 a_n2982_13878.n71 a_n2982_13878.n13 80.4688
R15039 a_n2982_13878.n71 a_n2982_13878.n90 0.365327
R15040 a_n2982_13878.n15 a_n2982_13878.n70 75.0448
R15041 a_n2982_13878.n69 a_n2982_13878.n15 70.1674
R15042 a_n2982_13878.n69 a_n2982_13878.n91 20.9683
R15043 a_n2982_13878.n16 a_n2982_13878.n68 70.3058
R15044 a_n2982_13878.n154 a_n2982_13878.n68 20.6913
R15045 a_n2982_13878.n67 a_n2982_13878.n16 75.3623
R15046 a_n2982_13878.n67 a_n2982_13878.n92 10.5784
R15047 a_n2982_13878.n18 a_n2982_13878.n17 44.7878
R15048 a_n2982_13878.n76 a_n2982_13878.n134 20.9683
R15049 a_n2982_13878.n75 a_n2982_13878.n12 75.0448
R15050 a_n2982_13878.n144 a_n2982_13878.n75 11.2134
R15051 a_n2982_13878.n12 a_n2982_13878.n145 161.3
R15052 a_n2982_13878.n78 a_n2982_13878.n135 20.9683
R15053 a_n2982_13878.n77 a_n2982_13878.n10 75.0448
R15054 a_n2982_13878.n142 a_n2982_13878.n77 11.2134
R15055 a_n2982_13878.n10 a_n2982_13878.n143 161.3
R15056 a_n2982_13878.n80 a_n2982_13878.n136 20.9683
R15057 a_n2982_13878.n79 a_n2982_13878.n8 75.0448
R15058 a_n2982_13878.n140 a_n2982_13878.n79 11.2134
R15059 a_n2982_13878.n8 a_n2982_13878.n141 161.3
R15060 a_n2982_13878.n82 a_n2982_13878.n137 20.9683
R15061 a_n2982_13878.n81 a_n2982_13878.n6 75.0448
R15062 a_n2982_13878.n138 a_n2982_13878.n81 11.2134
R15063 a_n2982_13878.n6 a_n2982_13878.n139 161.3
R15064 a_n2982_13878.n3 a_n2982_13878.n119 81.3764
R15065 a_n2982_13878.n4 a_n2982_13878.n113 81.3764
R15066 a_n2982_13878.n0 a_n2982_13878.n110 81.3764
R15067 a_n2982_13878.n3 a_n2982_13878.n120 80.9324
R15068 a_n2982_13878.n2 a_n2982_13878.n121 80.9324
R15069 a_n2982_13878.n2 a_n2982_13878.n118 80.9324
R15070 a_n2982_13878.n2 a_n2982_13878.n117 80.9324
R15071 a_n2982_13878.n1 a_n2982_13878.n116 80.9324
R15072 a_n2982_13878.n4 a_n2982_13878.n114 80.9324
R15073 a_n2982_13878.n0 a_n2982_13878.n115 80.9324
R15074 a_n2982_13878.n0 a_n2982_13878.n112 80.9324
R15075 a_n2982_13878.n0 a_n2982_13878.n111 80.9324
R15076 a_n2982_13878.n41 a_n2982_13878.t28 74.6477
R15077 a_n2982_13878.n40 a_n2982_13878.t22 74.6477
R15078 a_n2982_13878.n39 a_n2982_13878.t42 74.2899
R15079 a_n2982_13878.t6 a_n2982_13878.n43 74.2898
R15080 a_n2982_13878.n43 a_n2982_13878.n88 70.6783
R15081 a_n2982_13878.n42 a_n2982_13878.n87 70.6783
R15082 a_n2982_13878.n42 a_n2982_13878.n86 70.6783
R15083 a_n2982_13878.n41 a_n2982_13878.n85 70.6783
R15084 a_n2982_13878.n41 a_n2982_13878.n84 70.6783
R15085 a_n2982_13878.n40 a_n2982_13878.n128 70.6783
R15086 a_n2982_13878.n40 a_n2982_13878.n129 70.6783
R15087 a_n2982_13878.n38 a_n2982_13878.n130 70.6783
R15088 a_n2982_13878.n38 a_n2982_13878.n131 70.6783
R15089 a_n2982_13878.n39 a_n2982_13878.n132 70.6783
R15090 a_n2982_13878.n139 a_n2982_13878.n138 48.2005
R15091 a_n2982_13878.t99 a_n2982_13878.n82 533.335
R15092 a_n2982_13878.n141 a_n2982_13878.n140 48.2005
R15093 a_n2982_13878.t108 a_n2982_13878.n80 533.335
R15094 a_n2982_13878.n143 a_n2982_13878.n142 48.2005
R15095 a_n2982_13878.t93 a_n2982_13878.n78 533.335
R15096 a_n2982_13878.n145 a_n2982_13878.n144 48.2005
R15097 a_n2982_13878.t88 a_n2982_13878.n76 533.335
R15098 a_n2982_13878.n108 a_n2982_13878.n107 48.2005
R15099 a_n2982_13878.n46 a_n2982_13878.n105 20.9683
R15100 a_n2982_13878.n104 a_n2982_13878.n100 48.2005
R15101 a_n2982_13878.n102 a_n2982_13878.n50 20.9683
R15102 a_n2982_13878.n127 a_n2982_13878.n126 48.2005
R15103 a_n2982_13878.n55 a_n2982_13878.n124 20.9683
R15104 a_n2982_13878.n123 a_n2982_13878.n98 48.2005
R15105 a_n2982_13878.n109 a_n2982_13878.n83 48.2005
R15106 a_n2982_13878.n153 a_n2982_13878.n92 48.2005
R15107 a_n2982_13878.n155 a_n2982_13878.n69 20.9683
R15108 a_n2982_13878.n156 a_n2982_13878.n90 48.2005
R15109 a_n2982_13878.n158 a_n2982_13878.n73 20.9683
R15110 a_n2982_13878.n147 a_n2982_13878.n96 48.2005
R15111 a_n2982_13878.n149 a_n2982_13878.n61 20.9683
R15112 a_n2982_13878.n150 a_n2982_13878.n94 48.2005
R15113 a_n2982_13878.n152 a_n2982_13878.n65 20.9683
R15114 a_n2982_13878.n106 a_n2982_13878.n45 21.4216
R15115 a_n2982_13878.n125 a_n2982_13878.n54 21.4216
R15116 a_n2982_13878.n91 a_n2982_13878.n68 21.4216
R15117 a_n2982_13878.n95 a_n2982_13878.n60 21.4216
R15118 a_n2982_13878.n52 a_n2982_13878.t103 532.5
R15119 a_n2982_13878.n37 a_n2982_13878.t21 538.699
R15120 a_n2982_13878.t5 a_n2982_13878.n74 532.5
R15121 a_n2982_13878.t75 a_n2982_13878.n66 532.5
R15122 a_n2982_13878.n1 a_n2982_13878.n0 32.6799
R15123 a_n2982_13878.n49 a_n2982_13878.n101 34.4824
R15124 a_n2982_13878.n58 a_n2982_13878.n83 20.5623
R15125 a_n2982_13878.n89 a_n2982_13878.n72 34.4824
R15126 a_n2982_13878.n93 a_n2982_13878.n64 34.4824
R15127 a_n2982_13878.n81 a_n2982_13878.n137 35.3134
R15128 a_n2982_13878.n79 a_n2982_13878.n136 35.3134
R15129 a_n2982_13878.n77 a_n2982_13878.n135 35.3134
R15130 a_n2982_13878.n75 a_n2982_13878.n134 35.3134
R15131 a_n2982_13878.n105 a_n2982_13878.n47 35.3134
R15132 a_n2982_13878.n47 a_n2982_13878.n100 11.2134
R15133 a_n2982_13878.n124 a_n2982_13878.n56 35.3134
R15134 a_n2982_13878.n56 a_n2982_13878.n98 11.2134
R15135 a_n2982_13878.n70 a_n2982_13878.n155 35.3134
R15136 a_n2982_13878.n156 a_n2982_13878.n70 11.2134
R15137 a_n2982_13878.n62 a_n2982_13878.n149 35.3134
R15138 a_n2982_13878.n150 a_n2982_13878.n62 11.2134
R15139 a_n2982_13878.n36 a_n2982_13878.n2 23.891
R15140 a_n2982_13878.n44 a_n2982_13878.n99 36.139
R15141 a_n2982_13878.n53 a_n2982_13878.n97 36.139
R15142 a_n2982_13878.n154 a_n2982_13878.n67 36.139
R15143 a_n2982_13878.n148 a_n2982_13878.n59 36.139
R15144 a_n2982_13878.n23 a_n2982_13878.n146 13.9285
R15145 a_n2982_13878.n30 a_n2982_13878.n51 13.724
R15146 a_n2982_13878.n133 a_n2982_13878.n27 12.4191
R15147 a_n2982_13878.n146 a_n2982_13878.n12 11.2486
R15148 a_n2982_13878.n5 a_n2982_13878.n51 11.2486
R15149 a_n2982_13878.n43 a_n2982_13878.n159 10.5745
R15150 a_n2982_13878.n159 a_n2982_13878.n14 8.58383
R15151 a_n2982_13878.n133 a_n2982_13878.n39 6.7311
R15152 a_n2982_13878.n159 a_n2982_13878.n51 5.3452
R15153 a_n2982_13878.n36 a_n2982_13878.n33 3.94368
R15154 a_n2982_13878.n17 a_n2982_13878.n20 3.94368
R15155 a_n2982_13878.n88 a_n2982_13878.t32 3.61217
R15156 a_n2982_13878.n88 a_n2982_13878.t52 3.61217
R15157 a_n2982_13878.n87 a_n2982_13878.t20 3.61217
R15158 a_n2982_13878.n87 a_n2982_13878.t40 3.61217
R15159 a_n2982_13878.n86 a_n2982_13878.t16 3.61217
R15160 a_n2982_13878.n86 a_n2982_13878.t26 3.61217
R15161 a_n2982_13878.n85 a_n2982_13878.t38 3.61217
R15162 a_n2982_13878.n85 a_n2982_13878.t8 3.61217
R15163 a_n2982_13878.n84 a_n2982_13878.t30 3.61217
R15164 a_n2982_13878.n84 a_n2982_13878.t50 3.61217
R15165 a_n2982_13878.n128 a_n2982_13878.t44 3.61217
R15166 a_n2982_13878.n128 a_n2982_13878.t34 3.61217
R15167 a_n2982_13878.n129 a_n2982_13878.t46 3.61217
R15168 a_n2982_13878.n129 a_n2982_13878.t18 3.61217
R15169 a_n2982_13878.n130 a_n2982_13878.t14 3.61217
R15170 a_n2982_13878.n130 a_n2982_13878.t36 3.61217
R15171 a_n2982_13878.n131 a_n2982_13878.t10 3.61217
R15172 a_n2982_13878.n131 a_n2982_13878.t24 3.61217
R15173 a_n2982_13878.n132 a_n2982_13878.t48 3.61217
R15174 a_n2982_13878.n132 a_n2982_13878.t12 3.61217
R15175 a_n2982_13878.n119 a_n2982_13878.t2 2.82907
R15176 a_n2982_13878.n119 a_n2982_13878.t66 2.82907
R15177 a_n2982_13878.n120 a_n2982_13878.t70 2.82907
R15178 a_n2982_13878.n120 a_n2982_13878.t60 2.82907
R15179 a_n2982_13878.n121 a_n2982_13878.t55 2.82907
R15180 a_n2982_13878.n121 a_n2982_13878.t61 2.82907
R15181 a_n2982_13878.n118 a_n2982_13878.t62 2.82907
R15182 a_n2982_13878.n118 a_n2982_13878.t58 2.82907
R15183 a_n2982_13878.n117 a_n2982_13878.t53 2.82907
R15184 a_n2982_13878.n117 a_n2982_13878.t4 2.82907
R15185 a_n2982_13878.n116 a_n2982_13878.t0 2.82907
R15186 a_n2982_13878.n116 a_n2982_13878.t63 2.82907
R15187 a_n2982_13878.n113 a_n2982_13878.t57 2.82907
R15188 a_n2982_13878.n113 a_n2982_13878.t67 2.82907
R15189 a_n2982_13878.n114 a_n2982_13878.t65 2.82907
R15190 a_n2982_13878.n114 a_n2982_13878.t1 2.82907
R15191 a_n2982_13878.n115 a_n2982_13878.t59 2.82907
R15192 a_n2982_13878.n115 a_n2982_13878.t54 2.82907
R15193 a_n2982_13878.n112 a_n2982_13878.t3 2.82907
R15194 a_n2982_13878.n112 a_n2982_13878.t56 2.82907
R15195 a_n2982_13878.n111 a_n2982_13878.t69 2.82907
R15196 a_n2982_13878.n111 a_n2982_13878.t71 2.82907
R15197 a_n2982_13878.n110 a_n2982_13878.t64 2.82907
R15198 a_n2982_13878.n110 a_n2982_13878.t68 2.82907
R15199 a_n2982_13878.n35 a_n2982_13878.n108 14.1668
R15200 a_n2982_13878.n102 a_n2982_13878.n52 22.3251
R15201 a_n2982_13878.n29 a_n2982_13878.n127 14.1668
R15202 a_n2982_13878.n153 a_n2982_13878.n18 14.1668
R15203 a_n2982_13878.n74 a_n2982_13878.n158 22.3251
R15204 a_n2982_13878.n147 a_n2982_13878.n24 14.1668
R15205 a_n2982_13878.n66 a_n2982_13878.n152 22.3251
R15206 a_n2982_13878.n146 a_n2982_13878.n133 1.30542
R15207 a_n2982_13878.n9 a_n2982_13878.n8 1.04595
R15208 a_n2982_13878.n48 a_n2982_13878.n103 47.835
R15209 a_n2982_13878.n57 a_n2982_13878.n122 47.835
R15210 a_n2982_13878.n157 a_n2982_13878.n71 47.835
R15211 a_n2982_13878.n151 a_n2982_13878.n63 47.835
R15212 a_n2982_13878.n0 a_n2982_13878.n4 1.3324
R15213 a_n2982_13878.n31 a_n2982_13878.n30 1.13686
R15214 a_n2982_13878.n20 a_n2982_13878.n19 1.13686
R15215 a_n2982_13878.n14 a_n2982_13878.n13 1.13686
R15216 a_n2982_13878.n36 a_n2982_13878.n25 1.09898
R15217 a_n2982_13878.n42 a_n2982_13878.n41 1.07378
R15218 a_n2982_13878.n39 a_n2982_13878.n38 1.07378
R15219 a_n2982_13878.n2 a_n2982_13878.n3 0.888431
R15220 a_n2982_13878.n2 a_n2982_13878.n1 0.888431
R15221 a_n2982_13878.n34 a_n2982_13878.n33 0.758076
R15222 a_n2982_13878.n34 a_n2982_13878.n32 0.758076
R15223 a_n2982_13878.n32 a_n2982_13878.n31 0.758076
R15224 a_n2982_13878.n28 a_n2982_13878.n27 0.758076
R15225 a_n2982_13878.n28 a_n2982_13878.n26 0.758076
R15226 a_n2982_13878.n26 a_n2982_13878.n25 0.758076
R15227 a_n2982_13878.n22 a_n2982_13878.n23 0.758076
R15228 a_n2982_13878.n21 a_n2982_13878.n22 0.758076
R15229 a_n2982_13878.n19 a_n2982_13878.n21 0.758076
R15230 a_n2982_13878.n16 a_n2982_13878.n17 0.758076
R15231 a_n2982_13878.n15 a_n2982_13878.n16 0.758076
R15232 a_n2982_13878.n13 a_n2982_13878.n15 0.758076
R15233 a_n2982_13878.n12 a_n2982_13878.n11 0.758076
R15234 a_n2982_13878.n10 a_n2982_13878.n9 0.758076
R15235 a_n2982_13878.n8 a_n2982_13878.n7 0.758076
R15236 a_n2982_13878.n6 a_n2982_13878.n5 0.758076
R15237 a_n2982_13878.n43 a_n2982_13878.n42 0.716017
R15238 a_n2982_13878.n38 a_n2982_13878.n40 0.716017
R15239 a_n2982_13878.n11 a_n2982_13878.n10 0.67853
R15240 a_n2982_13878.n7 a_n2982_13878.n6 0.67853
R15241 vdd.n315 vdd.n279 756.745
R15242 vdd.n260 vdd.n224 756.745
R15243 vdd.n217 vdd.n181 756.745
R15244 vdd.n162 vdd.n126 756.745
R15245 vdd.n120 vdd.n84 756.745
R15246 vdd.n65 vdd.n29 756.745
R15247 vdd.n2139 vdd.n2103 756.745
R15248 vdd.n2194 vdd.n2158 756.745
R15249 vdd.n2041 vdd.n2005 756.745
R15250 vdd.n2096 vdd.n2060 756.745
R15251 vdd.n1944 vdd.n1908 756.745
R15252 vdd.n1999 vdd.n1963 756.745
R15253 vdd.n1286 vdd.t200 640.208
R15254 vdd.n981 vdd.t245 640.208
R15255 vdd.n1290 vdd.t235 640.208
R15256 vdd.n972 vdd.t269 640.208
R15257 vdd.n867 vdd.t222 640.208
R15258 vdd.n2740 vdd.t263 640.208
R15259 vdd.n804 vdd.t211 640.208
R15260 vdd.n2737 vdd.t252 640.208
R15261 vdd.n768 vdd.t196 640.208
R15262 vdd.n1042 vdd.t259 640.208
R15263 vdd.n1603 vdd.t241 592.009
R15264 vdd.n1759 vdd.t256 592.009
R15265 vdd.n1795 vdd.t266 592.009
R15266 vdd.n2279 vdd.t226 592.009
R15267 vdd.n1219 vdd.t204 592.009
R15268 vdd.n1179 vdd.t208 592.009
R15269 vdd.n405 vdd.t238 592.009
R15270 vdd.n419 vdd.t214 592.009
R15271 vdd.n431 vdd.t229 592.009
R15272 vdd.n723 vdd.t232 592.009
R15273 vdd.n686 vdd.t249 592.009
R15274 vdd.n3285 vdd.t218 592.009
R15275 vdd.n316 vdd.n315 585
R15276 vdd.n314 vdd.n281 585
R15277 vdd.n313 vdd.n312 585
R15278 vdd.n284 vdd.n282 585
R15279 vdd.n307 vdd.n306 585
R15280 vdd.n305 vdd.n304 585
R15281 vdd.n288 vdd.n287 585
R15282 vdd.n299 vdd.n298 585
R15283 vdd.n297 vdd.n296 585
R15284 vdd.n292 vdd.n291 585
R15285 vdd.n261 vdd.n260 585
R15286 vdd.n259 vdd.n226 585
R15287 vdd.n258 vdd.n257 585
R15288 vdd.n229 vdd.n227 585
R15289 vdd.n252 vdd.n251 585
R15290 vdd.n250 vdd.n249 585
R15291 vdd.n233 vdd.n232 585
R15292 vdd.n244 vdd.n243 585
R15293 vdd.n242 vdd.n241 585
R15294 vdd.n237 vdd.n236 585
R15295 vdd.n218 vdd.n217 585
R15296 vdd.n216 vdd.n183 585
R15297 vdd.n215 vdd.n214 585
R15298 vdd.n186 vdd.n184 585
R15299 vdd.n209 vdd.n208 585
R15300 vdd.n207 vdd.n206 585
R15301 vdd.n190 vdd.n189 585
R15302 vdd.n201 vdd.n200 585
R15303 vdd.n199 vdd.n198 585
R15304 vdd.n194 vdd.n193 585
R15305 vdd.n163 vdd.n162 585
R15306 vdd.n161 vdd.n128 585
R15307 vdd.n160 vdd.n159 585
R15308 vdd.n131 vdd.n129 585
R15309 vdd.n154 vdd.n153 585
R15310 vdd.n152 vdd.n151 585
R15311 vdd.n135 vdd.n134 585
R15312 vdd.n146 vdd.n145 585
R15313 vdd.n144 vdd.n143 585
R15314 vdd.n139 vdd.n138 585
R15315 vdd.n121 vdd.n120 585
R15316 vdd.n119 vdd.n86 585
R15317 vdd.n118 vdd.n117 585
R15318 vdd.n89 vdd.n87 585
R15319 vdd.n112 vdd.n111 585
R15320 vdd.n110 vdd.n109 585
R15321 vdd.n93 vdd.n92 585
R15322 vdd.n104 vdd.n103 585
R15323 vdd.n102 vdd.n101 585
R15324 vdd.n97 vdd.n96 585
R15325 vdd.n66 vdd.n65 585
R15326 vdd.n64 vdd.n31 585
R15327 vdd.n63 vdd.n62 585
R15328 vdd.n34 vdd.n32 585
R15329 vdd.n57 vdd.n56 585
R15330 vdd.n55 vdd.n54 585
R15331 vdd.n38 vdd.n37 585
R15332 vdd.n49 vdd.n48 585
R15333 vdd.n47 vdd.n46 585
R15334 vdd.n42 vdd.n41 585
R15335 vdd.n2140 vdd.n2139 585
R15336 vdd.n2138 vdd.n2105 585
R15337 vdd.n2137 vdd.n2136 585
R15338 vdd.n2108 vdd.n2106 585
R15339 vdd.n2131 vdd.n2130 585
R15340 vdd.n2129 vdd.n2128 585
R15341 vdd.n2112 vdd.n2111 585
R15342 vdd.n2123 vdd.n2122 585
R15343 vdd.n2121 vdd.n2120 585
R15344 vdd.n2116 vdd.n2115 585
R15345 vdd.n2195 vdd.n2194 585
R15346 vdd.n2193 vdd.n2160 585
R15347 vdd.n2192 vdd.n2191 585
R15348 vdd.n2163 vdd.n2161 585
R15349 vdd.n2186 vdd.n2185 585
R15350 vdd.n2184 vdd.n2183 585
R15351 vdd.n2167 vdd.n2166 585
R15352 vdd.n2178 vdd.n2177 585
R15353 vdd.n2176 vdd.n2175 585
R15354 vdd.n2171 vdd.n2170 585
R15355 vdd.n2042 vdd.n2041 585
R15356 vdd.n2040 vdd.n2007 585
R15357 vdd.n2039 vdd.n2038 585
R15358 vdd.n2010 vdd.n2008 585
R15359 vdd.n2033 vdd.n2032 585
R15360 vdd.n2031 vdd.n2030 585
R15361 vdd.n2014 vdd.n2013 585
R15362 vdd.n2025 vdd.n2024 585
R15363 vdd.n2023 vdd.n2022 585
R15364 vdd.n2018 vdd.n2017 585
R15365 vdd.n2097 vdd.n2096 585
R15366 vdd.n2095 vdd.n2062 585
R15367 vdd.n2094 vdd.n2093 585
R15368 vdd.n2065 vdd.n2063 585
R15369 vdd.n2088 vdd.n2087 585
R15370 vdd.n2086 vdd.n2085 585
R15371 vdd.n2069 vdd.n2068 585
R15372 vdd.n2080 vdd.n2079 585
R15373 vdd.n2078 vdd.n2077 585
R15374 vdd.n2073 vdd.n2072 585
R15375 vdd.n1945 vdd.n1944 585
R15376 vdd.n1943 vdd.n1910 585
R15377 vdd.n1942 vdd.n1941 585
R15378 vdd.n1913 vdd.n1911 585
R15379 vdd.n1936 vdd.n1935 585
R15380 vdd.n1934 vdd.n1933 585
R15381 vdd.n1917 vdd.n1916 585
R15382 vdd.n1928 vdd.n1927 585
R15383 vdd.n1926 vdd.n1925 585
R15384 vdd.n1921 vdd.n1920 585
R15385 vdd.n2000 vdd.n1999 585
R15386 vdd.n1998 vdd.n1965 585
R15387 vdd.n1997 vdd.n1996 585
R15388 vdd.n1968 vdd.n1966 585
R15389 vdd.n1991 vdd.n1990 585
R15390 vdd.n1989 vdd.n1988 585
R15391 vdd.n1972 vdd.n1971 585
R15392 vdd.n1983 vdd.n1982 585
R15393 vdd.n1981 vdd.n1980 585
R15394 vdd.n1976 vdd.n1975 585
R15395 vdd.n445 vdd.n370 462.44
R15396 vdd.n3523 vdd.n372 462.44
R15397 vdd.n3418 vdd.n657 462.44
R15398 vdd.n3416 vdd.n660 462.44
R15399 vdd.n2274 vdd.n1502 462.44
R15400 vdd.n2277 vdd.n2276 462.44
R15401 vdd.n1830 vdd.n1600 462.44
R15402 vdd.n1827 vdd.n1598 462.44
R15403 vdd.n293 vdd.t88 329.043
R15404 vdd.n238 vdd.t177 329.043
R15405 vdd.n195 vdd.t71 329.043
R15406 vdd.n140 vdd.t169 329.043
R15407 vdd.n98 vdd.t137 329.043
R15408 vdd.n43 vdd.t122 329.043
R15409 vdd.n2117 vdd.t107 329.043
R15410 vdd.n2172 vdd.t135 329.043
R15411 vdd.n2019 vdd.t90 329.043
R15412 vdd.n2074 vdd.t124 329.043
R15413 vdd.n1922 vdd.t126 329.043
R15414 vdd.n1977 vdd.t139 329.043
R15415 vdd.n1603 vdd.t244 319.788
R15416 vdd.n1759 vdd.t258 319.788
R15417 vdd.n1795 vdd.t268 319.788
R15418 vdd.n2279 vdd.t227 319.788
R15419 vdd.n1219 vdd.t206 319.788
R15420 vdd.n1179 vdd.t209 319.788
R15421 vdd.n405 vdd.t239 319.788
R15422 vdd.n419 vdd.t216 319.788
R15423 vdd.n431 vdd.t230 319.788
R15424 vdd.n723 vdd.t234 319.788
R15425 vdd.n686 vdd.t251 319.788
R15426 vdd.n3285 vdd.t221 319.788
R15427 vdd.n1604 vdd.t243 303.69
R15428 vdd.n1760 vdd.t257 303.69
R15429 vdd.n1796 vdd.t267 303.69
R15430 vdd.n2280 vdd.t228 303.69
R15431 vdd.n1220 vdd.t207 303.69
R15432 vdd.n1180 vdd.t210 303.69
R15433 vdd.n406 vdd.t240 303.69
R15434 vdd.n420 vdd.t217 303.69
R15435 vdd.n432 vdd.t231 303.69
R15436 vdd.n724 vdd.t233 303.69
R15437 vdd.n687 vdd.t250 303.69
R15438 vdd.n3286 vdd.t220 303.69
R15439 vdd.n3007 vdd.n931 279.512
R15440 vdd.n3247 vdd.n778 279.512
R15441 vdd.n3184 vdd.n775 279.512
R15442 vdd.n2939 vdd.n2938 279.512
R15443 vdd.n2700 vdd.n969 279.512
R15444 vdd.n2631 vdd.n2630 279.512
R15445 vdd.n1326 vdd.n1325 279.512
R15446 vdd.n2425 vdd.n1109 279.512
R15447 vdd.n3163 vdd.n776 279.512
R15448 vdd.n3250 vdd.n3249 279.512
R15449 vdd.n2812 vdd.n2735 279.512
R15450 vdd.n2743 vdd.n927 279.512
R15451 vdd.n2628 vdd.n979 279.512
R15452 vdd.n977 vdd.n951 279.512
R15453 vdd.n1451 vdd.n1146 279.512
R15454 vdd.n1251 vdd.n1104 279.512
R15455 vdd.n2423 vdd.n1112 254.619
R15456 vdd.n756 vdd.n658 254.619
R15457 vdd.n3165 vdd.n776 185
R15458 vdd.n3248 vdd.n776 185
R15459 vdd.n3167 vdd.n3166 185
R15460 vdd.n3166 vdd.n774 185
R15461 vdd.n3168 vdd.n810 185
R15462 vdd.n3178 vdd.n810 185
R15463 vdd.n3169 vdd.n819 185
R15464 vdd.n819 vdd.n817 185
R15465 vdd.n3171 vdd.n3170 185
R15466 vdd.n3172 vdd.n3171 185
R15467 vdd.n3124 vdd.n818 185
R15468 vdd.n818 vdd.n814 185
R15469 vdd.n3123 vdd.n3122 185
R15470 vdd.n3122 vdd.n3121 185
R15471 vdd.n821 vdd.n820 185
R15472 vdd.n822 vdd.n821 185
R15473 vdd.n3114 vdd.n3113 185
R15474 vdd.n3115 vdd.n3114 185
R15475 vdd.n3112 vdd.n830 185
R15476 vdd.n835 vdd.n830 185
R15477 vdd.n3111 vdd.n3110 185
R15478 vdd.n3110 vdd.n3109 185
R15479 vdd.n832 vdd.n831 185
R15480 vdd.n841 vdd.n832 185
R15481 vdd.n3102 vdd.n3101 185
R15482 vdd.n3103 vdd.n3102 185
R15483 vdd.n3100 vdd.n842 185
R15484 vdd.n848 vdd.n842 185
R15485 vdd.n3099 vdd.n3098 185
R15486 vdd.n3098 vdd.n3097 185
R15487 vdd.n844 vdd.n843 185
R15488 vdd.n845 vdd.n844 185
R15489 vdd.n3090 vdd.n3089 185
R15490 vdd.n3091 vdd.n3090 185
R15491 vdd.n3088 vdd.n855 185
R15492 vdd.n855 vdd.n852 185
R15493 vdd.n3087 vdd.n3086 185
R15494 vdd.n3086 vdd.n3085 185
R15495 vdd.n857 vdd.n856 185
R15496 vdd.n858 vdd.n857 185
R15497 vdd.n3078 vdd.n3077 185
R15498 vdd.n3079 vdd.n3078 185
R15499 vdd.n3076 vdd.n866 185
R15500 vdd.n872 vdd.n866 185
R15501 vdd.n3075 vdd.n3074 185
R15502 vdd.n3074 vdd.n3073 185
R15503 vdd.n3064 vdd.n869 185
R15504 vdd.n879 vdd.n869 185
R15505 vdd.n3066 vdd.n3065 185
R15506 vdd.n3067 vdd.n3066 185
R15507 vdd.n3063 vdd.n880 185
R15508 vdd.n880 vdd.n876 185
R15509 vdd.n3062 vdd.n3061 185
R15510 vdd.n3061 vdd.n3060 185
R15511 vdd.n882 vdd.n881 185
R15512 vdd.n883 vdd.n882 185
R15513 vdd.n3053 vdd.n3052 185
R15514 vdd.n3054 vdd.n3053 185
R15515 vdd.n3051 vdd.n891 185
R15516 vdd.n896 vdd.n891 185
R15517 vdd.n3050 vdd.n3049 185
R15518 vdd.n3049 vdd.n3048 185
R15519 vdd.n893 vdd.n892 185
R15520 vdd.n902 vdd.n893 185
R15521 vdd.n3041 vdd.n3040 185
R15522 vdd.n3042 vdd.n3041 185
R15523 vdd.n3039 vdd.n903 185
R15524 vdd.n2915 vdd.n903 185
R15525 vdd.n3038 vdd.n3037 185
R15526 vdd.n3037 vdd.n3036 185
R15527 vdd.n905 vdd.n904 185
R15528 vdd.n2921 vdd.n905 185
R15529 vdd.n3029 vdd.n3028 185
R15530 vdd.n3030 vdd.n3029 185
R15531 vdd.n3027 vdd.n914 185
R15532 vdd.n914 vdd.n911 185
R15533 vdd.n3026 vdd.n3025 185
R15534 vdd.n3025 vdd.n3024 185
R15535 vdd.n916 vdd.n915 185
R15536 vdd.n917 vdd.n916 185
R15537 vdd.n3017 vdd.n3016 185
R15538 vdd.n3018 vdd.n3017 185
R15539 vdd.n3015 vdd.n925 185
R15540 vdd.n2933 vdd.n925 185
R15541 vdd.n3014 vdd.n3013 185
R15542 vdd.n3013 vdd.n3012 185
R15543 vdd.n927 vdd.n926 185
R15544 vdd.n928 vdd.n927 185
R15545 vdd.n2744 vdd.n2743 185
R15546 vdd.n2746 vdd.n2745 185
R15547 vdd.n2748 vdd.n2747 185
R15548 vdd.n2750 vdd.n2749 185
R15549 vdd.n2752 vdd.n2751 185
R15550 vdd.n2754 vdd.n2753 185
R15551 vdd.n2756 vdd.n2755 185
R15552 vdd.n2758 vdd.n2757 185
R15553 vdd.n2760 vdd.n2759 185
R15554 vdd.n2762 vdd.n2761 185
R15555 vdd.n2764 vdd.n2763 185
R15556 vdd.n2766 vdd.n2765 185
R15557 vdd.n2768 vdd.n2767 185
R15558 vdd.n2770 vdd.n2769 185
R15559 vdd.n2772 vdd.n2771 185
R15560 vdd.n2774 vdd.n2773 185
R15561 vdd.n2776 vdd.n2775 185
R15562 vdd.n2778 vdd.n2777 185
R15563 vdd.n2780 vdd.n2779 185
R15564 vdd.n2782 vdd.n2781 185
R15565 vdd.n2784 vdd.n2783 185
R15566 vdd.n2786 vdd.n2785 185
R15567 vdd.n2788 vdd.n2787 185
R15568 vdd.n2790 vdd.n2789 185
R15569 vdd.n2792 vdd.n2791 185
R15570 vdd.n2794 vdd.n2793 185
R15571 vdd.n2796 vdd.n2795 185
R15572 vdd.n2798 vdd.n2797 185
R15573 vdd.n2800 vdd.n2799 185
R15574 vdd.n2802 vdd.n2801 185
R15575 vdd.n2804 vdd.n2803 185
R15576 vdd.n2806 vdd.n2805 185
R15577 vdd.n2808 vdd.n2807 185
R15578 vdd.n2810 vdd.n2809 185
R15579 vdd.n2811 vdd.n2735 185
R15580 vdd.n3005 vdd.n2735 185
R15581 vdd.n3251 vdd.n3250 185
R15582 vdd.n3252 vdd.n767 185
R15583 vdd.n3254 vdd.n3253 185
R15584 vdd.n3256 vdd.n765 185
R15585 vdd.n3258 vdd.n3257 185
R15586 vdd.n3259 vdd.n764 185
R15587 vdd.n3261 vdd.n3260 185
R15588 vdd.n3263 vdd.n762 185
R15589 vdd.n3265 vdd.n3264 185
R15590 vdd.n3266 vdd.n761 185
R15591 vdd.n3268 vdd.n3267 185
R15592 vdd.n3270 vdd.n759 185
R15593 vdd.n3272 vdd.n3271 185
R15594 vdd.n3273 vdd.n758 185
R15595 vdd.n3275 vdd.n3274 185
R15596 vdd.n3277 vdd.n757 185
R15597 vdd.n3278 vdd.n754 185
R15598 vdd.n3281 vdd.n3280 185
R15599 vdd.n755 vdd.n753 185
R15600 vdd.n3137 vdd.n3136 185
R15601 vdd.n3139 vdd.n3138 185
R15602 vdd.n3141 vdd.n3133 185
R15603 vdd.n3143 vdd.n3142 185
R15604 vdd.n3144 vdd.n3132 185
R15605 vdd.n3146 vdd.n3145 185
R15606 vdd.n3148 vdd.n3130 185
R15607 vdd.n3150 vdd.n3149 185
R15608 vdd.n3151 vdd.n3129 185
R15609 vdd.n3153 vdd.n3152 185
R15610 vdd.n3155 vdd.n3127 185
R15611 vdd.n3157 vdd.n3156 185
R15612 vdd.n3158 vdd.n3126 185
R15613 vdd.n3160 vdd.n3159 185
R15614 vdd.n3162 vdd.n3125 185
R15615 vdd.n3164 vdd.n3163 185
R15616 vdd.n3163 vdd.n756 185
R15617 vdd.n3249 vdd.n771 185
R15618 vdd.n3249 vdd.n3248 185
R15619 vdd.n2866 vdd.n773 185
R15620 vdd.n774 vdd.n773 185
R15621 vdd.n2867 vdd.n809 185
R15622 vdd.n3178 vdd.n809 185
R15623 vdd.n2869 vdd.n2868 185
R15624 vdd.n2868 vdd.n817 185
R15625 vdd.n2870 vdd.n816 185
R15626 vdd.n3172 vdd.n816 185
R15627 vdd.n2872 vdd.n2871 185
R15628 vdd.n2871 vdd.n814 185
R15629 vdd.n2873 vdd.n824 185
R15630 vdd.n3121 vdd.n824 185
R15631 vdd.n2875 vdd.n2874 185
R15632 vdd.n2874 vdd.n822 185
R15633 vdd.n2876 vdd.n829 185
R15634 vdd.n3115 vdd.n829 185
R15635 vdd.n2878 vdd.n2877 185
R15636 vdd.n2877 vdd.n835 185
R15637 vdd.n2879 vdd.n834 185
R15638 vdd.n3109 vdd.n834 185
R15639 vdd.n2881 vdd.n2880 185
R15640 vdd.n2880 vdd.n841 185
R15641 vdd.n2882 vdd.n840 185
R15642 vdd.n3103 vdd.n840 185
R15643 vdd.n2884 vdd.n2883 185
R15644 vdd.n2883 vdd.n848 185
R15645 vdd.n2885 vdd.n847 185
R15646 vdd.n3097 vdd.n847 185
R15647 vdd.n2887 vdd.n2886 185
R15648 vdd.n2886 vdd.n845 185
R15649 vdd.n2888 vdd.n854 185
R15650 vdd.n3091 vdd.n854 185
R15651 vdd.n2890 vdd.n2889 185
R15652 vdd.n2889 vdd.n852 185
R15653 vdd.n2891 vdd.n860 185
R15654 vdd.n3085 vdd.n860 185
R15655 vdd.n2893 vdd.n2892 185
R15656 vdd.n2892 vdd.n858 185
R15657 vdd.n2894 vdd.n865 185
R15658 vdd.n3079 vdd.n865 185
R15659 vdd.n2896 vdd.n2895 185
R15660 vdd.n2895 vdd.n872 185
R15661 vdd.n2897 vdd.n871 185
R15662 vdd.n3073 vdd.n871 185
R15663 vdd.n2899 vdd.n2898 185
R15664 vdd.n2898 vdd.n879 185
R15665 vdd.n2900 vdd.n878 185
R15666 vdd.n3067 vdd.n878 185
R15667 vdd.n2902 vdd.n2901 185
R15668 vdd.n2901 vdd.n876 185
R15669 vdd.n2903 vdd.n885 185
R15670 vdd.n3060 vdd.n885 185
R15671 vdd.n2905 vdd.n2904 185
R15672 vdd.n2904 vdd.n883 185
R15673 vdd.n2906 vdd.n890 185
R15674 vdd.n3054 vdd.n890 185
R15675 vdd.n2908 vdd.n2907 185
R15676 vdd.n2907 vdd.n896 185
R15677 vdd.n2909 vdd.n895 185
R15678 vdd.n3048 vdd.n895 185
R15679 vdd.n2911 vdd.n2910 185
R15680 vdd.n2910 vdd.n902 185
R15681 vdd.n2912 vdd.n901 185
R15682 vdd.n3042 vdd.n901 185
R15683 vdd.n2914 vdd.n2913 185
R15684 vdd.n2915 vdd.n2914 185
R15685 vdd.n2815 vdd.n907 185
R15686 vdd.n3036 vdd.n907 185
R15687 vdd.n2923 vdd.n2922 185
R15688 vdd.n2922 vdd.n2921 185
R15689 vdd.n2924 vdd.n913 185
R15690 vdd.n3030 vdd.n913 185
R15691 vdd.n2926 vdd.n2925 185
R15692 vdd.n2925 vdd.n911 185
R15693 vdd.n2927 vdd.n919 185
R15694 vdd.n3024 vdd.n919 185
R15695 vdd.n2929 vdd.n2928 185
R15696 vdd.n2928 vdd.n917 185
R15697 vdd.n2930 vdd.n924 185
R15698 vdd.n3018 vdd.n924 185
R15699 vdd.n2932 vdd.n2931 185
R15700 vdd.n2933 vdd.n2932 185
R15701 vdd.n2814 vdd.n930 185
R15702 vdd.n3012 vdd.n930 185
R15703 vdd.n2813 vdd.n2812 185
R15704 vdd.n2812 vdd.n928 185
R15705 vdd.n2274 vdd.n2273 185
R15706 vdd.n2275 vdd.n2274 185
R15707 vdd.n1503 vdd.n1501 185
R15708 vdd.n1501 vdd.n1500 185
R15709 vdd.n2269 vdd.n2268 185
R15710 vdd.n2268 vdd.n2267 185
R15711 vdd.n1506 vdd.n1505 185
R15712 vdd.n1507 vdd.n1506 185
R15713 vdd.n2256 vdd.n2255 185
R15714 vdd.n2257 vdd.n2256 185
R15715 vdd.n1515 vdd.n1514 185
R15716 vdd.n2248 vdd.n1514 185
R15717 vdd.n2251 vdd.n2250 185
R15718 vdd.n2250 vdd.n2249 185
R15719 vdd.n1518 vdd.n1517 185
R15720 vdd.n1524 vdd.n1518 185
R15721 vdd.n2239 vdd.n2238 185
R15722 vdd.n2240 vdd.n2239 185
R15723 vdd.n1526 vdd.n1525 185
R15724 vdd.n2231 vdd.n1525 185
R15725 vdd.n2234 vdd.n2233 185
R15726 vdd.n2233 vdd.n2232 185
R15727 vdd.n1529 vdd.n1528 185
R15728 vdd.n1530 vdd.n1529 185
R15729 vdd.n2222 vdd.n2221 185
R15730 vdd.n2223 vdd.n2222 185
R15731 vdd.n1538 vdd.n1537 185
R15732 vdd.n1537 vdd.n1536 185
R15733 vdd.n2217 vdd.n2216 185
R15734 vdd.n2216 vdd.n2215 185
R15735 vdd.n1541 vdd.n1540 185
R15736 vdd.n1547 vdd.n1541 185
R15737 vdd.n2206 vdd.n2205 185
R15738 vdd.n2207 vdd.n2206 185
R15739 vdd.n1549 vdd.n1548 185
R15740 vdd.n1903 vdd.n1548 185
R15741 vdd.n1906 vdd.n1905 185
R15742 vdd.n1905 vdd.n1904 185
R15743 vdd.n1552 vdd.n1551 185
R15744 vdd.n1559 vdd.n1552 185
R15745 vdd.n1894 vdd.n1893 185
R15746 vdd.n1895 vdd.n1894 185
R15747 vdd.n1561 vdd.n1560 185
R15748 vdd.n1560 vdd.n1558 185
R15749 vdd.n1889 vdd.n1888 185
R15750 vdd.n1888 vdd.n1887 185
R15751 vdd.n1564 vdd.n1563 185
R15752 vdd.n1565 vdd.n1564 185
R15753 vdd.n1878 vdd.n1877 185
R15754 vdd.n1879 vdd.n1878 185
R15755 vdd.n1572 vdd.n1571 185
R15756 vdd.n1870 vdd.n1571 185
R15757 vdd.n1873 vdd.n1872 185
R15758 vdd.n1872 vdd.n1871 185
R15759 vdd.n1575 vdd.n1574 185
R15760 vdd.n1581 vdd.n1575 185
R15761 vdd.n1861 vdd.n1860 185
R15762 vdd.n1862 vdd.n1861 185
R15763 vdd.n1583 vdd.n1582 185
R15764 vdd.n1853 vdd.n1582 185
R15765 vdd.n1856 vdd.n1855 185
R15766 vdd.n1855 vdd.n1854 185
R15767 vdd.n1586 vdd.n1585 185
R15768 vdd.n1587 vdd.n1586 185
R15769 vdd.n1844 vdd.n1843 185
R15770 vdd.n1845 vdd.n1844 185
R15771 vdd.n1595 vdd.n1594 185
R15772 vdd.n1594 vdd.n1593 185
R15773 vdd.n1839 vdd.n1838 185
R15774 vdd.n1838 vdd.n1837 185
R15775 vdd.n1598 vdd.n1597 185
R15776 vdd.n1599 vdd.n1598 185
R15777 vdd.n1827 vdd.n1826 185
R15778 vdd.n1825 vdd.n1638 185
R15779 vdd.n1640 vdd.n1637 185
R15780 vdd.n1829 vdd.n1637 185
R15781 vdd.n1821 vdd.n1642 185
R15782 vdd.n1820 vdd.n1643 185
R15783 vdd.n1819 vdd.n1644 185
R15784 vdd.n1647 vdd.n1645 185
R15785 vdd.n1815 vdd.n1648 185
R15786 vdd.n1814 vdd.n1649 185
R15787 vdd.n1813 vdd.n1650 185
R15788 vdd.n1653 vdd.n1651 185
R15789 vdd.n1809 vdd.n1654 185
R15790 vdd.n1808 vdd.n1655 185
R15791 vdd.n1807 vdd.n1656 185
R15792 vdd.n1659 vdd.n1657 185
R15793 vdd.n1803 vdd.n1660 185
R15794 vdd.n1802 vdd.n1661 185
R15795 vdd.n1801 vdd.n1662 185
R15796 vdd.n1793 vdd.n1663 185
R15797 vdd.n1797 vdd.n1794 185
R15798 vdd.n1792 vdd.n1665 185
R15799 vdd.n1791 vdd.n1666 185
R15800 vdd.n1669 vdd.n1667 185
R15801 vdd.n1787 vdd.n1670 185
R15802 vdd.n1786 vdd.n1671 185
R15803 vdd.n1785 vdd.n1672 185
R15804 vdd.n1675 vdd.n1673 185
R15805 vdd.n1781 vdd.n1676 185
R15806 vdd.n1780 vdd.n1677 185
R15807 vdd.n1779 vdd.n1678 185
R15808 vdd.n1681 vdd.n1679 185
R15809 vdd.n1775 vdd.n1682 185
R15810 vdd.n1774 vdd.n1683 185
R15811 vdd.n1773 vdd.n1684 185
R15812 vdd.n1687 vdd.n1685 185
R15813 vdd.n1769 vdd.n1688 185
R15814 vdd.n1768 vdd.n1689 185
R15815 vdd.n1767 vdd.n1690 185
R15816 vdd.n1693 vdd.n1691 185
R15817 vdd.n1763 vdd.n1694 185
R15818 vdd.n1762 vdd.n1695 185
R15819 vdd.n1761 vdd.n1758 185
R15820 vdd.n1698 vdd.n1696 185
R15821 vdd.n1754 vdd.n1699 185
R15822 vdd.n1753 vdd.n1700 185
R15823 vdd.n1752 vdd.n1701 185
R15824 vdd.n1704 vdd.n1702 185
R15825 vdd.n1748 vdd.n1705 185
R15826 vdd.n1747 vdd.n1706 185
R15827 vdd.n1746 vdd.n1707 185
R15828 vdd.n1710 vdd.n1708 185
R15829 vdd.n1742 vdd.n1711 185
R15830 vdd.n1741 vdd.n1712 185
R15831 vdd.n1740 vdd.n1713 185
R15832 vdd.n1716 vdd.n1714 185
R15833 vdd.n1736 vdd.n1717 185
R15834 vdd.n1735 vdd.n1718 185
R15835 vdd.n1734 vdd.n1719 185
R15836 vdd.n1722 vdd.n1720 185
R15837 vdd.n1730 vdd.n1723 185
R15838 vdd.n1729 vdd.n1724 185
R15839 vdd.n1728 vdd.n1725 185
R15840 vdd.n1726 vdd.n1606 185
R15841 vdd.n1831 vdd.n1830 185
R15842 vdd.n1830 vdd.n1829 185
R15843 vdd.n2278 vdd.n2277 185
R15844 vdd.n2282 vdd.n1496 185
R15845 vdd.n1495 vdd.n1489 185
R15846 vdd.n1493 vdd.n1492 185
R15847 vdd.n1491 vdd.n1250 185
R15848 vdd.n2286 vdd.n1247 185
R15849 vdd.n2288 vdd.n2287 185
R15850 vdd.n2290 vdd.n1245 185
R15851 vdd.n2292 vdd.n2291 185
R15852 vdd.n2293 vdd.n1240 185
R15853 vdd.n2295 vdd.n2294 185
R15854 vdd.n2297 vdd.n1238 185
R15855 vdd.n2299 vdd.n2298 185
R15856 vdd.n2300 vdd.n1233 185
R15857 vdd.n2302 vdd.n2301 185
R15858 vdd.n2304 vdd.n1231 185
R15859 vdd.n2306 vdd.n2305 185
R15860 vdd.n2307 vdd.n1227 185
R15861 vdd.n2309 vdd.n2308 185
R15862 vdd.n2311 vdd.n1224 185
R15863 vdd.n2313 vdd.n2312 185
R15864 vdd.n1225 vdd.n1218 185
R15865 vdd.n2317 vdd.n1222 185
R15866 vdd.n2318 vdd.n1214 185
R15867 vdd.n2320 vdd.n2319 185
R15868 vdd.n2322 vdd.n1212 185
R15869 vdd.n2324 vdd.n2323 185
R15870 vdd.n2325 vdd.n1207 185
R15871 vdd.n2327 vdd.n2326 185
R15872 vdd.n2329 vdd.n1205 185
R15873 vdd.n2331 vdd.n2330 185
R15874 vdd.n2332 vdd.n1200 185
R15875 vdd.n2334 vdd.n2333 185
R15876 vdd.n2336 vdd.n1198 185
R15877 vdd.n2338 vdd.n2337 185
R15878 vdd.n2339 vdd.n1193 185
R15879 vdd.n2341 vdd.n2340 185
R15880 vdd.n2343 vdd.n1191 185
R15881 vdd.n2345 vdd.n2344 185
R15882 vdd.n2346 vdd.n1187 185
R15883 vdd.n2348 vdd.n2347 185
R15884 vdd.n2350 vdd.n1184 185
R15885 vdd.n2352 vdd.n2351 185
R15886 vdd.n1185 vdd.n1178 185
R15887 vdd.n2356 vdd.n1182 185
R15888 vdd.n2357 vdd.n1174 185
R15889 vdd.n2359 vdd.n2358 185
R15890 vdd.n2361 vdd.n1172 185
R15891 vdd.n2363 vdd.n2362 185
R15892 vdd.n2364 vdd.n1167 185
R15893 vdd.n2366 vdd.n2365 185
R15894 vdd.n2368 vdd.n1165 185
R15895 vdd.n2370 vdd.n2369 185
R15896 vdd.n2371 vdd.n1160 185
R15897 vdd.n2373 vdd.n2372 185
R15898 vdd.n2375 vdd.n1158 185
R15899 vdd.n2377 vdd.n2376 185
R15900 vdd.n2378 vdd.n1156 185
R15901 vdd.n2380 vdd.n2379 185
R15902 vdd.n2383 vdd.n2382 185
R15903 vdd.n2385 vdd.n2384 185
R15904 vdd.n2387 vdd.n1154 185
R15905 vdd.n2389 vdd.n2388 185
R15906 vdd.n1502 vdd.n1153 185
R15907 vdd.n2276 vdd.n1499 185
R15908 vdd.n2276 vdd.n2275 185
R15909 vdd.n1510 vdd.n1498 185
R15910 vdd.n1500 vdd.n1498 185
R15911 vdd.n2266 vdd.n2265 185
R15912 vdd.n2267 vdd.n2266 185
R15913 vdd.n1509 vdd.n1508 185
R15914 vdd.n1508 vdd.n1507 185
R15915 vdd.n2259 vdd.n2258 185
R15916 vdd.n2258 vdd.n2257 185
R15917 vdd.n1513 vdd.n1512 185
R15918 vdd.n2248 vdd.n1513 185
R15919 vdd.n2247 vdd.n2246 185
R15920 vdd.n2249 vdd.n2247 185
R15921 vdd.n1520 vdd.n1519 185
R15922 vdd.n1524 vdd.n1519 185
R15923 vdd.n2242 vdd.n2241 185
R15924 vdd.n2241 vdd.n2240 185
R15925 vdd.n1523 vdd.n1522 185
R15926 vdd.n2231 vdd.n1523 185
R15927 vdd.n2230 vdd.n2229 185
R15928 vdd.n2232 vdd.n2230 185
R15929 vdd.n1532 vdd.n1531 185
R15930 vdd.n1531 vdd.n1530 185
R15931 vdd.n2225 vdd.n2224 185
R15932 vdd.n2224 vdd.n2223 185
R15933 vdd.n1535 vdd.n1534 185
R15934 vdd.n1536 vdd.n1535 185
R15935 vdd.n2214 vdd.n2213 185
R15936 vdd.n2215 vdd.n2214 185
R15937 vdd.n1543 vdd.n1542 185
R15938 vdd.n1547 vdd.n1542 185
R15939 vdd.n2209 vdd.n2208 185
R15940 vdd.n2208 vdd.n2207 185
R15941 vdd.n1546 vdd.n1545 185
R15942 vdd.n1903 vdd.n1546 185
R15943 vdd.n1902 vdd.n1901 185
R15944 vdd.n1904 vdd.n1902 185
R15945 vdd.n1554 vdd.n1553 185
R15946 vdd.n1559 vdd.n1553 185
R15947 vdd.n1897 vdd.n1896 185
R15948 vdd.n1896 vdd.n1895 185
R15949 vdd.n1557 vdd.n1556 185
R15950 vdd.n1558 vdd.n1557 185
R15951 vdd.n1886 vdd.n1885 185
R15952 vdd.n1887 vdd.n1886 185
R15953 vdd.n1567 vdd.n1566 185
R15954 vdd.n1566 vdd.n1565 185
R15955 vdd.n1881 vdd.n1880 185
R15956 vdd.n1880 vdd.n1879 185
R15957 vdd.n1570 vdd.n1569 185
R15958 vdd.n1870 vdd.n1570 185
R15959 vdd.n1869 vdd.n1868 185
R15960 vdd.n1871 vdd.n1869 185
R15961 vdd.n1577 vdd.n1576 185
R15962 vdd.n1581 vdd.n1576 185
R15963 vdd.n1864 vdd.n1863 185
R15964 vdd.n1863 vdd.n1862 185
R15965 vdd.n1580 vdd.n1579 185
R15966 vdd.n1853 vdd.n1580 185
R15967 vdd.n1852 vdd.n1851 185
R15968 vdd.n1854 vdd.n1852 185
R15969 vdd.n1589 vdd.n1588 185
R15970 vdd.n1588 vdd.n1587 185
R15971 vdd.n1847 vdd.n1846 185
R15972 vdd.n1846 vdd.n1845 185
R15973 vdd.n1592 vdd.n1591 185
R15974 vdd.n1593 vdd.n1592 185
R15975 vdd.n1836 vdd.n1835 185
R15976 vdd.n1837 vdd.n1836 185
R15977 vdd.n1601 vdd.n1600 185
R15978 vdd.n1600 vdd.n1599 185
R15979 vdd.n971 vdd.n969 185
R15980 vdd.n2629 vdd.n969 185
R15981 vdd.n2551 vdd.n989 185
R15982 vdd.n989 vdd.n976 185
R15983 vdd.n2553 vdd.n2552 185
R15984 vdd.n2554 vdd.n2553 185
R15985 vdd.n2550 vdd.n988 185
R15986 vdd.n1370 vdd.n988 185
R15987 vdd.n2549 vdd.n2548 185
R15988 vdd.n2548 vdd.n2547 185
R15989 vdd.n991 vdd.n990 185
R15990 vdd.n992 vdd.n991 185
R15991 vdd.n2538 vdd.n2537 185
R15992 vdd.n2539 vdd.n2538 185
R15993 vdd.n2536 vdd.n1002 185
R15994 vdd.n1002 vdd.n999 185
R15995 vdd.n2535 vdd.n2534 185
R15996 vdd.n2534 vdd.n2533 185
R15997 vdd.n1004 vdd.n1003 185
R15998 vdd.n1396 vdd.n1004 185
R15999 vdd.n2526 vdd.n2525 185
R16000 vdd.n2527 vdd.n2526 185
R16001 vdd.n2524 vdd.n1012 185
R16002 vdd.n1017 vdd.n1012 185
R16003 vdd.n2523 vdd.n2522 185
R16004 vdd.n2522 vdd.n2521 185
R16005 vdd.n1014 vdd.n1013 185
R16006 vdd.n1023 vdd.n1014 185
R16007 vdd.n2514 vdd.n2513 185
R16008 vdd.n2515 vdd.n2514 185
R16009 vdd.n2512 vdd.n1024 185
R16010 vdd.n1408 vdd.n1024 185
R16011 vdd.n2511 vdd.n2510 185
R16012 vdd.n2510 vdd.n2509 185
R16013 vdd.n1026 vdd.n1025 185
R16014 vdd.n1027 vdd.n1026 185
R16015 vdd.n2502 vdd.n2501 185
R16016 vdd.n2503 vdd.n2502 185
R16017 vdd.n2500 vdd.n1036 185
R16018 vdd.n1036 vdd.n1033 185
R16019 vdd.n2499 vdd.n2498 185
R16020 vdd.n2498 vdd.n2497 185
R16021 vdd.n1038 vdd.n1037 185
R16022 vdd.n1047 vdd.n1038 185
R16023 vdd.n2489 vdd.n2488 185
R16024 vdd.n2490 vdd.n2489 185
R16025 vdd.n2487 vdd.n1048 185
R16026 vdd.n1054 vdd.n1048 185
R16027 vdd.n2486 vdd.n2485 185
R16028 vdd.n2485 vdd.n2484 185
R16029 vdd.n1050 vdd.n1049 185
R16030 vdd.n1051 vdd.n1050 185
R16031 vdd.n2477 vdd.n2476 185
R16032 vdd.n2478 vdd.n2477 185
R16033 vdd.n2475 vdd.n1061 185
R16034 vdd.n1061 vdd.n1058 185
R16035 vdd.n2474 vdd.n2473 185
R16036 vdd.n2473 vdd.n2472 185
R16037 vdd.n1063 vdd.n1062 185
R16038 vdd.n1064 vdd.n1063 185
R16039 vdd.n2465 vdd.n2464 185
R16040 vdd.n2466 vdd.n2465 185
R16041 vdd.n2463 vdd.n1072 185
R16042 vdd.n1077 vdd.n1072 185
R16043 vdd.n2462 vdd.n2461 185
R16044 vdd.n2461 vdd.n2460 185
R16045 vdd.n1074 vdd.n1073 185
R16046 vdd.n1083 vdd.n1074 185
R16047 vdd.n2453 vdd.n2452 185
R16048 vdd.n2454 vdd.n2453 185
R16049 vdd.n2451 vdd.n1084 185
R16050 vdd.n1090 vdd.n1084 185
R16051 vdd.n2450 vdd.n2449 185
R16052 vdd.n2449 vdd.n2448 185
R16053 vdd.n1086 vdd.n1085 185
R16054 vdd.n1087 vdd.n1086 185
R16055 vdd.n2441 vdd.n2440 185
R16056 vdd.n2442 vdd.n2441 185
R16057 vdd.n2439 vdd.n1097 185
R16058 vdd.n1097 vdd.n1094 185
R16059 vdd.n2438 vdd.n2437 185
R16060 vdd.n2437 vdd.n2436 185
R16061 vdd.n1099 vdd.n1098 185
R16062 vdd.n1108 vdd.n1099 185
R16063 vdd.n2429 vdd.n2428 185
R16064 vdd.n2430 vdd.n2429 185
R16065 vdd.n2427 vdd.n1109 185
R16066 vdd.n1109 vdd.n1105 185
R16067 vdd.n2426 vdd.n2425 185
R16068 vdd.n1111 vdd.n1110 185
R16069 vdd.n2422 vdd.n2421 185
R16070 vdd.n2423 vdd.n2422 185
R16071 vdd.n2420 vdd.n1147 185
R16072 vdd.n2419 vdd.n2418 185
R16073 vdd.n2417 vdd.n2416 185
R16074 vdd.n2415 vdd.n2414 185
R16075 vdd.n2413 vdd.n2412 185
R16076 vdd.n2411 vdd.n2410 185
R16077 vdd.n2409 vdd.n2408 185
R16078 vdd.n2407 vdd.n2406 185
R16079 vdd.n2405 vdd.n2404 185
R16080 vdd.n2403 vdd.n2402 185
R16081 vdd.n2401 vdd.n2400 185
R16082 vdd.n2399 vdd.n2398 185
R16083 vdd.n2397 vdd.n2396 185
R16084 vdd.n2395 vdd.n2394 185
R16085 vdd.n2393 vdd.n2392 185
R16086 vdd.n1292 vdd.n1148 185
R16087 vdd.n1294 vdd.n1293 185
R16088 vdd.n1296 vdd.n1295 185
R16089 vdd.n1298 vdd.n1297 185
R16090 vdd.n1300 vdd.n1299 185
R16091 vdd.n1302 vdd.n1301 185
R16092 vdd.n1304 vdd.n1303 185
R16093 vdd.n1306 vdd.n1305 185
R16094 vdd.n1308 vdd.n1307 185
R16095 vdd.n1310 vdd.n1309 185
R16096 vdd.n1312 vdd.n1311 185
R16097 vdd.n1314 vdd.n1313 185
R16098 vdd.n1316 vdd.n1315 185
R16099 vdd.n1318 vdd.n1317 185
R16100 vdd.n1321 vdd.n1320 185
R16101 vdd.n1323 vdd.n1322 185
R16102 vdd.n1325 vdd.n1324 185
R16103 vdd.n2632 vdd.n2631 185
R16104 vdd.n2634 vdd.n2633 185
R16105 vdd.n2636 vdd.n2635 185
R16106 vdd.n2639 vdd.n2638 185
R16107 vdd.n2641 vdd.n2640 185
R16108 vdd.n2643 vdd.n2642 185
R16109 vdd.n2645 vdd.n2644 185
R16110 vdd.n2647 vdd.n2646 185
R16111 vdd.n2649 vdd.n2648 185
R16112 vdd.n2651 vdd.n2650 185
R16113 vdd.n2653 vdd.n2652 185
R16114 vdd.n2655 vdd.n2654 185
R16115 vdd.n2657 vdd.n2656 185
R16116 vdd.n2659 vdd.n2658 185
R16117 vdd.n2661 vdd.n2660 185
R16118 vdd.n2663 vdd.n2662 185
R16119 vdd.n2665 vdd.n2664 185
R16120 vdd.n2667 vdd.n2666 185
R16121 vdd.n2669 vdd.n2668 185
R16122 vdd.n2671 vdd.n2670 185
R16123 vdd.n2673 vdd.n2672 185
R16124 vdd.n2675 vdd.n2674 185
R16125 vdd.n2677 vdd.n2676 185
R16126 vdd.n2679 vdd.n2678 185
R16127 vdd.n2681 vdd.n2680 185
R16128 vdd.n2683 vdd.n2682 185
R16129 vdd.n2685 vdd.n2684 185
R16130 vdd.n2687 vdd.n2686 185
R16131 vdd.n2689 vdd.n2688 185
R16132 vdd.n2691 vdd.n2690 185
R16133 vdd.n2693 vdd.n2692 185
R16134 vdd.n2695 vdd.n2694 185
R16135 vdd.n2697 vdd.n2696 185
R16136 vdd.n2698 vdd.n970 185
R16137 vdd.n2700 vdd.n2699 185
R16138 vdd.n2701 vdd.n2700 185
R16139 vdd.n2630 vdd.n974 185
R16140 vdd.n2630 vdd.n2629 185
R16141 vdd.n1368 vdd.n975 185
R16142 vdd.n976 vdd.n975 185
R16143 vdd.n1369 vdd.n986 185
R16144 vdd.n2554 vdd.n986 185
R16145 vdd.n1372 vdd.n1371 185
R16146 vdd.n1371 vdd.n1370 185
R16147 vdd.n1373 vdd.n993 185
R16148 vdd.n2547 vdd.n993 185
R16149 vdd.n1375 vdd.n1374 185
R16150 vdd.n1374 vdd.n992 185
R16151 vdd.n1376 vdd.n1000 185
R16152 vdd.n2539 vdd.n1000 185
R16153 vdd.n1378 vdd.n1377 185
R16154 vdd.n1377 vdd.n999 185
R16155 vdd.n1379 vdd.n1005 185
R16156 vdd.n2533 vdd.n1005 185
R16157 vdd.n1398 vdd.n1397 185
R16158 vdd.n1397 vdd.n1396 185
R16159 vdd.n1399 vdd.n1010 185
R16160 vdd.n2527 vdd.n1010 185
R16161 vdd.n1401 vdd.n1400 185
R16162 vdd.n1400 vdd.n1017 185
R16163 vdd.n1402 vdd.n1015 185
R16164 vdd.n2521 vdd.n1015 185
R16165 vdd.n1404 vdd.n1403 185
R16166 vdd.n1403 vdd.n1023 185
R16167 vdd.n1405 vdd.n1021 185
R16168 vdd.n2515 vdd.n1021 185
R16169 vdd.n1407 vdd.n1406 185
R16170 vdd.n1408 vdd.n1407 185
R16171 vdd.n1367 vdd.n1028 185
R16172 vdd.n2509 vdd.n1028 185
R16173 vdd.n1366 vdd.n1365 185
R16174 vdd.n1365 vdd.n1027 185
R16175 vdd.n1364 vdd.n1034 185
R16176 vdd.n2503 vdd.n1034 185
R16177 vdd.n1363 vdd.n1362 185
R16178 vdd.n1362 vdd.n1033 185
R16179 vdd.n1361 vdd.n1039 185
R16180 vdd.n2497 vdd.n1039 185
R16181 vdd.n1360 vdd.n1359 185
R16182 vdd.n1359 vdd.n1047 185
R16183 vdd.n1358 vdd.n1045 185
R16184 vdd.n2490 vdd.n1045 185
R16185 vdd.n1357 vdd.n1356 185
R16186 vdd.n1356 vdd.n1054 185
R16187 vdd.n1355 vdd.n1052 185
R16188 vdd.n2484 vdd.n1052 185
R16189 vdd.n1354 vdd.n1353 185
R16190 vdd.n1353 vdd.n1051 185
R16191 vdd.n1352 vdd.n1059 185
R16192 vdd.n2478 vdd.n1059 185
R16193 vdd.n1351 vdd.n1350 185
R16194 vdd.n1350 vdd.n1058 185
R16195 vdd.n1349 vdd.n1065 185
R16196 vdd.n2472 vdd.n1065 185
R16197 vdd.n1348 vdd.n1347 185
R16198 vdd.n1347 vdd.n1064 185
R16199 vdd.n1346 vdd.n1070 185
R16200 vdd.n2466 vdd.n1070 185
R16201 vdd.n1345 vdd.n1344 185
R16202 vdd.n1344 vdd.n1077 185
R16203 vdd.n1343 vdd.n1075 185
R16204 vdd.n2460 vdd.n1075 185
R16205 vdd.n1342 vdd.n1341 185
R16206 vdd.n1341 vdd.n1083 185
R16207 vdd.n1340 vdd.n1081 185
R16208 vdd.n2454 vdd.n1081 185
R16209 vdd.n1339 vdd.n1338 185
R16210 vdd.n1338 vdd.n1090 185
R16211 vdd.n1337 vdd.n1088 185
R16212 vdd.n2448 vdd.n1088 185
R16213 vdd.n1336 vdd.n1335 185
R16214 vdd.n1335 vdd.n1087 185
R16215 vdd.n1334 vdd.n1095 185
R16216 vdd.n2442 vdd.n1095 185
R16217 vdd.n1333 vdd.n1332 185
R16218 vdd.n1332 vdd.n1094 185
R16219 vdd.n1331 vdd.n1100 185
R16220 vdd.n2436 vdd.n1100 185
R16221 vdd.n1330 vdd.n1329 185
R16222 vdd.n1329 vdd.n1108 185
R16223 vdd.n1328 vdd.n1106 185
R16224 vdd.n2430 vdd.n1106 185
R16225 vdd.n1327 vdd.n1326 185
R16226 vdd.n1326 vdd.n1105 185
R16227 vdd.n370 vdd.n369 185
R16228 vdd.n3526 vdd.n370 185
R16229 vdd.n3529 vdd.n3528 185
R16230 vdd.n3528 vdd.n3527 185
R16231 vdd.n3530 vdd.n364 185
R16232 vdd.n364 vdd.n363 185
R16233 vdd.n3532 vdd.n3531 185
R16234 vdd.n3533 vdd.n3532 185
R16235 vdd.n359 vdd.n358 185
R16236 vdd.n3534 vdd.n359 185
R16237 vdd.n3537 vdd.n3536 185
R16238 vdd.n3536 vdd.n3535 185
R16239 vdd.n3538 vdd.n353 185
R16240 vdd.n3508 vdd.n353 185
R16241 vdd.n3540 vdd.n3539 185
R16242 vdd.n3541 vdd.n3540 185
R16243 vdd.n348 vdd.n347 185
R16244 vdd.n3542 vdd.n348 185
R16245 vdd.n3545 vdd.n3544 185
R16246 vdd.n3544 vdd.n3543 185
R16247 vdd.n3546 vdd.n342 185
R16248 vdd.n349 vdd.n342 185
R16249 vdd.n3548 vdd.n3547 185
R16250 vdd.n3549 vdd.n3548 185
R16251 vdd.n338 vdd.n337 185
R16252 vdd.n3550 vdd.n338 185
R16253 vdd.n3553 vdd.n3552 185
R16254 vdd.n3552 vdd.n3551 185
R16255 vdd.n3554 vdd.n333 185
R16256 vdd.n333 vdd.n332 185
R16257 vdd.n3556 vdd.n3555 185
R16258 vdd.n3557 vdd.n3556 185
R16259 vdd.n327 vdd.n325 185
R16260 vdd.n3558 vdd.n327 185
R16261 vdd.n3561 vdd.n3560 185
R16262 vdd.n3560 vdd.n3559 185
R16263 vdd.n326 vdd.n324 185
R16264 vdd.n328 vdd.n326 185
R16265 vdd.n3484 vdd.n3483 185
R16266 vdd.n3485 vdd.n3484 185
R16267 vdd.n615 vdd.n614 185
R16268 vdd.n614 vdd.n613 185
R16269 vdd.n3479 vdd.n3478 185
R16270 vdd.n3478 vdd.n3477 185
R16271 vdd.n618 vdd.n617 185
R16272 vdd.n624 vdd.n618 185
R16273 vdd.n3465 vdd.n3464 185
R16274 vdd.n3466 vdd.n3465 185
R16275 vdd.n626 vdd.n625 185
R16276 vdd.n3457 vdd.n625 185
R16277 vdd.n3460 vdd.n3459 185
R16278 vdd.n3459 vdd.n3458 185
R16279 vdd.n629 vdd.n628 185
R16280 vdd.n636 vdd.n629 185
R16281 vdd.n3448 vdd.n3447 185
R16282 vdd.n3449 vdd.n3448 185
R16283 vdd.n638 vdd.n637 185
R16284 vdd.n637 vdd.n635 185
R16285 vdd.n3443 vdd.n3442 185
R16286 vdd.n3442 vdd.n3441 185
R16287 vdd.n641 vdd.n640 185
R16288 vdd.n642 vdd.n641 185
R16289 vdd.n3432 vdd.n3431 185
R16290 vdd.n3433 vdd.n3432 185
R16291 vdd.n650 vdd.n649 185
R16292 vdd.n649 vdd.n648 185
R16293 vdd.n3427 vdd.n3426 185
R16294 vdd.n3426 vdd.n3425 185
R16295 vdd.n653 vdd.n652 185
R16296 vdd.n659 vdd.n653 185
R16297 vdd.n3416 vdd.n3415 185
R16298 vdd.n3417 vdd.n3416 185
R16299 vdd.n3412 vdd.n660 185
R16300 vdd.n3411 vdd.n3410 185
R16301 vdd.n3408 vdd.n662 185
R16302 vdd.n3408 vdd.n658 185
R16303 vdd.n3407 vdd.n3406 185
R16304 vdd.n3405 vdd.n3404 185
R16305 vdd.n3403 vdd.n3402 185
R16306 vdd.n3401 vdd.n3400 185
R16307 vdd.n3399 vdd.n668 185
R16308 vdd.n3397 vdd.n3396 185
R16309 vdd.n3395 vdd.n669 185
R16310 vdd.n3394 vdd.n3393 185
R16311 vdd.n3391 vdd.n674 185
R16312 vdd.n3389 vdd.n3388 185
R16313 vdd.n3387 vdd.n675 185
R16314 vdd.n3386 vdd.n3385 185
R16315 vdd.n3383 vdd.n680 185
R16316 vdd.n3381 vdd.n3380 185
R16317 vdd.n3379 vdd.n681 185
R16318 vdd.n3378 vdd.n3377 185
R16319 vdd.n3375 vdd.n688 185
R16320 vdd.n3373 vdd.n3372 185
R16321 vdd.n3371 vdd.n689 185
R16322 vdd.n3370 vdd.n3369 185
R16323 vdd.n3367 vdd.n694 185
R16324 vdd.n3365 vdd.n3364 185
R16325 vdd.n3363 vdd.n695 185
R16326 vdd.n3362 vdd.n3361 185
R16327 vdd.n3359 vdd.n700 185
R16328 vdd.n3357 vdd.n3356 185
R16329 vdd.n3355 vdd.n701 185
R16330 vdd.n3354 vdd.n3353 185
R16331 vdd.n3351 vdd.n706 185
R16332 vdd.n3349 vdd.n3348 185
R16333 vdd.n3347 vdd.n707 185
R16334 vdd.n3346 vdd.n3345 185
R16335 vdd.n3343 vdd.n712 185
R16336 vdd.n3341 vdd.n3340 185
R16337 vdd.n3339 vdd.n713 185
R16338 vdd.n3338 vdd.n3337 185
R16339 vdd.n3335 vdd.n718 185
R16340 vdd.n3333 vdd.n3332 185
R16341 vdd.n3331 vdd.n719 185
R16342 vdd.n728 vdd.n722 185
R16343 vdd.n3327 vdd.n3326 185
R16344 vdd.n3324 vdd.n726 185
R16345 vdd.n3323 vdd.n3322 185
R16346 vdd.n3321 vdd.n3320 185
R16347 vdd.n3319 vdd.n732 185
R16348 vdd.n3317 vdd.n3316 185
R16349 vdd.n3315 vdd.n733 185
R16350 vdd.n3314 vdd.n3313 185
R16351 vdd.n3311 vdd.n738 185
R16352 vdd.n3309 vdd.n3308 185
R16353 vdd.n3307 vdd.n739 185
R16354 vdd.n3306 vdd.n3305 185
R16355 vdd.n3303 vdd.n744 185
R16356 vdd.n3301 vdd.n3300 185
R16357 vdd.n3299 vdd.n745 185
R16358 vdd.n3298 vdd.n3297 185
R16359 vdd.n3295 vdd.n3294 185
R16360 vdd.n3293 vdd.n3292 185
R16361 vdd.n3291 vdd.n3290 185
R16362 vdd.n3289 vdd.n3288 185
R16363 vdd.n3284 vdd.n657 185
R16364 vdd.n658 vdd.n657 185
R16365 vdd.n3523 vdd.n3522 185
R16366 vdd.n599 vdd.n404 185
R16367 vdd.n598 vdd.n597 185
R16368 vdd.n596 vdd.n595 185
R16369 vdd.n594 vdd.n409 185
R16370 vdd.n590 vdd.n589 185
R16371 vdd.n588 vdd.n587 185
R16372 vdd.n586 vdd.n585 185
R16373 vdd.n584 vdd.n411 185
R16374 vdd.n580 vdd.n579 185
R16375 vdd.n578 vdd.n577 185
R16376 vdd.n576 vdd.n575 185
R16377 vdd.n574 vdd.n413 185
R16378 vdd.n570 vdd.n569 185
R16379 vdd.n568 vdd.n567 185
R16380 vdd.n566 vdd.n565 185
R16381 vdd.n564 vdd.n415 185
R16382 vdd.n560 vdd.n559 185
R16383 vdd.n558 vdd.n557 185
R16384 vdd.n556 vdd.n555 185
R16385 vdd.n554 vdd.n417 185
R16386 vdd.n550 vdd.n549 185
R16387 vdd.n548 vdd.n547 185
R16388 vdd.n546 vdd.n545 185
R16389 vdd.n544 vdd.n421 185
R16390 vdd.n540 vdd.n539 185
R16391 vdd.n538 vdd.n537 185
R16392 vdd.n536 vdd.n535 185
R16393 vdd.n534 vdd.n423 185
R16394 vdd.n530 vdd.n529 185
R16395 vdd.n528 vdd.n527 185
R16396 vdd.n526 vdd.n525 185
R16397 vdd.n524 vdd.n425 185
R16398 vdd.n520 vdd.n519 185
R16399 vdd.n518 vdd.n517 185
R16400 vdd.n516 vdd.n515 185
R16401 vdd.n514 vdd.n427 185
R16402 vdd.n510 vdd.n509 185
R16403 vdd.n508 vdd.n507 185
R16404 vdd.n506 vdd.n505 185
R16405 vdd.n504 vdd.n429 185
R16406 vdd.n500 vdd.n499 185
R16407 vdd.n498 vdd.n497 185
R16408 vdd.n496 vdd.n495 185
R16409 vdd.n494 vdd.n433 185
R16410 vdd.n490 vdd.n489 185
R16411 vdd.n488 vdd.n487 185
R16412 vdd.n486 vdd.n485 185
R16413 vdd.n484 vdd.n435 185
R16414 vdd.n480 vdd.n479 185
R16415 vdd.n478 vdd.n477 185
R16416 vdd.n476 vdd.n475 185
R16417 vdd.n474 vdd.n437 185
R16418 vdd.n470 vdd.n469 185
R16419 vdd.n468 vdd.n467 185
R16420 vdd.n466 vdd.n465 185
R16421 vdd.n464 vdd.n439 185
R16422 vdd.n460 vdd.n459 185
R16423 vdd.n458 vdd.n457 185
R16424 vdd.n456 vdd.n455 185
R16425 vdd.n454 vdd.n441 185
R16426 vdd.n450 vdd.n449 185
R16427 vdd.n448 vdd.n447 185
R16428 vdd.n446 vdd.n445 185
R16429 vdd.n3519 vdd.n372 185
R16430 vdd.n3526 vdd.n372 185
R16431 vdd.n3518 vdd.n371 185
R16432 vdd.n3527 vdd.n371 185
R16433 vdd.n3517 vdd.n3516 185
R16434 vdd.n3516 vdd.n363 185
R16435 vdd.n602 vdd.n362 185
R16436 vdd.n3533 vdd.n362 185
R16437 vdd.n3512 vdd.n361 185
R16438 vdd.n3534 vdd.n361 185
R16439 vdd.n3511 vdd.n360 185
R16440 vdd.n3535 vdd.n360 185
R16441 vdd.n3510 vdd.n3509 185
R16442 vdd.n3509 vdd.n3508 185
R16443 vdd.n604 vdd.n352 185
R16444 vdd.n3541 vdd.n352 185
R16445 vdd.n3504 vdd.n351 185
R16446 vdd.n3542 vdd.n351 185
R16447 vdd.n3503 vdd.n350 185
R16448 vdd.n3543 vdd.n350 185
R16449 vdd.n3502 vdd.n3501 185
R16450 vdd.n3501 vdd.n349 185
R16451 vdd.n606 vdd.n341 185
R16452 vdd.n3549 vdd.n341 185
R16453 vdd.n3497 vdd.n340 185
R16454 vdd.n3550 vdd.n340 185
R16455 vdd.n3496 vdd.n339 185
R16456 vdd.n3551 vdd.n339 185
R16457 vdd.n3495 vdd.n3494 185
R16458 vdd.n3494 vdd.n332 185
R16459 vdd.n608 vdd.n331 185
R16460 vdd.n3557 vdd.n331 185
R16461 vdd.n3490 vdd.n330 185
R16462 vdd.n3558 vdd.n330 185
R16463 vdd.n3489 vdd.n329 185
R16464 vdd.n3559 vdd.n329 185
R16465 vdd.n3488 vdd.n3487 185
R16466 vdd.n3487 vdd.n328 185
R16467 vdd.n3486 vdd.n610 185
R16468 vdd.n3486 vdd.n3485 185
R16469 vdd.n3474 vdd.n612 185
R16470 vdd.n613 vdd.n612 185
R16471 vdd.n3476 vdd.n3475 185
R16472 vdd.n3477 vdd.n3476 185
R16473 vdd.n620 vdd.n619 185
R16474 vdd.n624 vdd.n619 185
R16475 vdd.n3468 vdd.n3467 185
R16476 vdd.n3467 vdd.n3466 185
R16477 vdd.n623 vdd.n622 185
R16478 vdd.n3457 vdd.n623 185
R16479 vdd.n3456 vdd.n3455 185
R16480 vdd.n3458 vdd.n3456 185
R16481 vdd.n631 vdd.n630 185
R16482 vdd.n636 vdd.n630 185
R16483 vdd.n3451 vdd.n3450 185
R16484 vdd.n3450 vdd.n3449 185
R16485 vdd.n634 vdd.n633 185
R16486 vdd.n635 vdd.n634 185
R16487 vdd.n3440 vdd.n3439 185
R16488 vdd.n3441 vdd.n3440 185
R16489 vdd.n644 vdd.n643 185
R16490 vdd.n643 vdd.n642 185
R16491 vdd.n3435 vdd.n3434 185
R16492 vdd.n3434 vdd.n3433 185
R16493 vdd.n647 vdd.n646 185
R16494 vdd.n648 vdd.n647 185
R16495 vdd.n3424 vdd.n3423 185
R16496 vdd.n3425 vdd.n3424 185
R16497 vdd.n655 vdd.n654 185
R16498 vdd.n659 vdd.n654 185
R16499 vdd.n3419 vdd.n3418 185
R16500 vdd.n3418 vdd.n3417 185
R16501 vdd.n3008 vdd.n3007 185
R16502 vdd.n933 vdd.n932 185
R16503 vdd.n3004 vdd.n3003 185
R16504 vdd.n3005 vdd.n3004 185
R16505 vdd.n3002 vdd.n2736 185
R16506 vdd.n3001 vdd.n3000 185
R16507 vdd.n2999 vdd.n2998 185
R16508 vdd.n2997 vdd.n2996 185
R16509 vdd.n2995 vdd.n2994 185
R16510 vdd.n2993 vdd.n2992 185
R16511 vdd.n2991 vdd.n2990 185
R16512 vdd.n2989 vdd.n2988 185
R16513 vdd.n2987 vdd.n2986 185
R16514 vdd.n2985 vdd.n2984 185
R16515 vdd.n2983 vdd.n2982 185
R16516 vdd.n2981 vdd.n2980 185
R16517 vdd.n2979 vdd.n2978 185
R16518 vdd.n2977 vdd.n2976 185
R16519 vdd.n2975 vdd.n2974 185
R16520 vdd.n2973 vdd.n2972 185
R16521 vdd.n2971 vdd.n2970 185
R16522 vdd.n2969 vdd.n2968 185
R16523 vdd.n2967 vdd.n2966 185
R16524 vdd.n2965 vdd.n2964 185
R16525 vdd.n2963 vdd.n2962 185
R16526 vdd.n2961 vdd.n2960 185
R16527 vdd.n2959 vdd.n2958 185
R16528 vdd.n2957 vdd.n2956 185
R16529 vdd.n2955 vdd.n2954 185
R16530 vdd.n2953 vdd.n2952 185
R16531 vdd.n2951 vdd.n2950 185
R16532 vdd.n2949 vdd.n2948 185
R16533 vdd.n2947 vdd.n2946 185
R16534 vdd.n2944 vdd.n2943 185
R16535 vdd.n2942 vdd.n2941 185
R16536 vdd.n2940 vdd.n2939 185
R16537 vdd.n3185 vdd.n3184 185
R16538 vdd.n3186 vdd.n803 185
R16539 vdd.n3188 vdd.n3187 185
R16540 vdd.n3190 vdd.n801 185
R16541 vdd.n3192 vdd.n3191 185
R16542 vdd.n3193 vdd.n800 185
R16543 vdd.n3195 vdd.n3194 185
R16544 vdd.n3197 vdd.n798 185
R16545 vdd.n3199 vdd.n3198 185
R16546 vdd.n3200 vdd.n797 185
R16547 vdd.n3202 vdd.n3201 185
R16548 vdd.n3204 vdd.n795 185
R16549 vdd.n3206 vdd.n3205 185
R16550 vdd.n3207 vdd.n794 185
R16551 vdd.n3209 vdd.n3208 185
R16552 vdd.n3211 vdd.n792 185
R16553 vdd.n3213 vdd.n3212 185
R16554 vdd.n3215 vdd.n791 185
R16555 vdd.n3217 vdd.n3216 185
R16556 vdd.n3219 vdd.n789 185
R16557 vdd.n3221 vdd.n3220 185
R16558 vdd.n3222 vdd.n788 185
R16559 vdd.n3224 vdd.n3223 185
R16560 vdd.n3226 vdd.n786 185
R16561 vdd.n3228 vdd.n3227 185
R16562 vdd.n3229 vdd.n785 185
R16563 vdd.n3231 vdd.n3230 185
R16564 vdd.n3233 vdd.n783 185
R16565 vdd.n3235 vdd.n3234 185
R16566 vdd.n3236 vdd.n782 185
R16567 vdd.n3238 vdd.n3237 185
R16568 vdd.n3240 vdd.n781 185
R16569 vdd.n3241 vdd.n780 185
R16570 vdd.n3244 vdd.n3243 185
R16571 vdd.n3245 vdd.n778 185
R16572 vdd.n778 vdd.n756 185
R16573 vdd.n3182 vdd.n775 185
R16574 vdd.n3248 vdd.n775 185
R16575 vdd.n3181 vdd.n3180 185
R16576 vdd.n3180 vdd.n774 185
R16577 vdd.n3179 vdd.n807 185
R16578 vdd.n3179 vdd.n3178 185
R16579 vdd.n2822 vdd.n808 185
R16580 vdd.n817 vdd.n808 185
R16581 vdd.n2823 vdd.n815 185
R16582 vdd.n3172 vdd.n815 185
R16583 vdd.n2825 vdd.n2824 185
R16584 vdd.n2824 vdd.n814 185
R16585 vdd.n2826 vdd.n823 185
R16586 vdd.n3121 vdd.n823 185
R16587 vdd.n2828 vdd.n2827 185
R16588 vdd.n2827 vdd.n822 185
R16589 vdd.n2829 vdd.n828 185
R16590 vdd.n3115 vdd.n828 185
R16591 vdd.n2831 vdd.n2830 185
R16592 vdd.n2830 vdd.n835 185
R16593 vdd.n2832 vdd.n833 185
R16594 vdd.n3109 vdd.n833 185
R16595 vdd.n2834 vdd.n2833 185
R16596 vdd.n2833 vdd.n841 185
R16597 vdd.n2835 vdd.n839 185
R16598 vdd.n3103 vdd.n839 185
R16599 vdd.n2837 vdd.n2836 185
R16600 vdd.n2836 vdd.n848 185
R16601 vdd.n2838 vdd.n846 185
R16602 vdd.n3097 vdd.n846 185
R16603 vdd.n2840 vdd.n2839 185
R16604 vdd.n2839 vdd.n845 185
R16605 vdd.n2841 vdd.n853 185
R16606 vdd.n3091 vdd.n853 185
R16607 vdd.n2843 vdd.n2842 185
R16608 vdd.n2842 vdd.n852 185
R16609 vdd.n2844 vdd.n859 185
R16610 vdd.n3085 vdd.n859 185
R16611 vdd.n2846 vdd.n2845 185
R16612 vdd.n2845 vdd.n858 185
R16613 vdd.n2847 vdd.n864 185
R16614 vdd.n3079 vdd.n864 185
R16615 vdd.n2849 vdd.n2848 185
R16616 vdd.n2848 vdd.n872 185
R16617 vdd.n2850 vdd.n870 185
R16618 vdd.n3073 vdd.n870 185
R16619 vdd.n2852 vdd.n2851 185
R16620 vdd.n2851 vdd.n879 185
R16621 vdd.n2853 vdd.n877 185
R16622 vdd.n3067 vdd.n877 185
R16623 vdd.n2855 vdd.n2854 185
R16624 vdd.n2854 vdd.n876 185
R16625 vdd.n2856 vdd.n884 185
R16626 vdd.n3060 vdd.n884 185
R16627 vdd.n2858 vdd.n2857 185
R16628 vdd.n2857 vdd.n883 185
R16629 vdd.n2859 vdd.n889 185
R16630 vdd.n3054 vdd.n889 185
R16631 vdd.n2861 vdd.n2860 185
R16632 vdd.n2860 vdd.n896 185
R16633 vdd.n2862 vdd.n894 185
R16634 vdd.n3048 vdd.n894 185
R16635 vdd.n2864 vdd.n2863 185
R16636 vdd.n2863 vdd.n902 185
R16637 vdd.n2865 vdd.n900 185
R16638 vdd.n3042 vdd.n900 185
R16639 vdd.n2917 vdd.n2916 185
R16640 vdd.n2916 vdd.n2915 185
R16641 vdd.n2918 vdd.n906 185
R16642 vdd.n3036 vdd.n906 185
R16643 vdd.n2920 vdd.n2919 185
R16644 vdd.n2921 vdd.n2920 185
R16645 vdd.n2821 vdd.n912 185
R16646 vdd.n3030 vdd.n912 185
R16647 vdd.n2820 vdd.n2819 185
R16648 vdd.n2819 vdd.n911 185
R16649 vdd.n2818 vdd.n918 185
R16650 vdd.n3024 vdd.n918 185
R16651 vdd.n2817 vdd.n2816 185
R16652 vdd.n2816 vdd.n917 185
R16653 vdd.n2739 vdd.n923 185
R16654 vdd.n3018 vdd.n923 185
R16655 vdd.n2935 vdd.n2934 185
R16656 vdd.n2934 vdd.n2933 185
R16657 vdd.n2936 vdd.n929 185
R16658 vdd.n3012 vdd.n929 185
R16659 vdd.n2938 vdd.n2937 185
R16660 vdd.n2938 vdd.n928 185
R16661 vdd.n3009 vdd.n931 185
R16662 vdd.n931 vdd.n928 185
R16663 vdd.n3011 vdd.n3010 185
R16664 vdd.n3012 vdd.n3011 185
R16665 vdd.n922 vdd.n921 185
R16666 vdd.n2933 vdd.n922 185
R16667 vdd.n3020 vdd.n3019 185
R16668 vdd.n3019 vdd.n3018 185
R16669 vdd.n3021 vdd.n920 185
R16670 vdd.n920 vdd.n917 185
R16671 vdd.n3023 vdd.n3022 185
R16672 vdd.n3024 vdd.n3023 185
R16673 vdd.n910 vdd.n909 185
R16674 vdd.n911 vdd.n910 185
R16675 vdd.n3032 vdd.n3031 185
R16676 vdd.n3031 vdd.n3030 185
R16677 vdd.n3033 vdd.n908 185
R16678 vdd.n2921 vdd.n908 185
R16679 vdd.n3035 vdd.n3034 185
R16680 vdd.n3036 vdd.n3035 185
R16681 vdd.n899 vdd.n898 185
R16682 vdd.n2915 vdd.n899 185
R16683 vdd.n3044 vdd.n3043 185
R16684 vdd.n3043 vdd.n3042 185
R16685 vdd.n3045 vdd.n897 185
R16686 vdd.n902 vdd.n897 185
R16687 vdd.n3047 vdd.n3046 185
R16688 vdd.n3048 vdd.n3047 185
R16689 vdd.n888 vdd.n887 185
R16690 vdd.n896 vdd.n888 185
R16691 vdd.n3056 vdd.n3055 185
R16692 vdd.n3055 vdd.n3054 185
R16693 vdd.n3057 vdd.n886 185
R16694 vdd.n886 vdd.n883 185
R16695 vdd.n3059 vdd.n3058 185
R16696 vdd.n3060 vdd.n3059 185
R16697 vdd.n875 vdd.n874 185
R16698 vdd.n876 vdd.n875 185
R16699 vdd.n3069 vdd.n3068 185
R16700 vdd.n3068 vdd.n3067 185
R16701 vdd.n3070 vdd.n873 185
R16702 vdd.n879 vdd.n873 185
R16703 vdd.n3072 vdd.n3071 185
R16704 vdd.n3073 vdd.n3072 185
R16705 vdd.n863 vdd.n862 185
R16706 vdd.n872 vdd.n863 185
R16707 vdd.n3081 vdd.n3080 185
R16708 vdd.n3080 vdd.n3079 185
R16709 vdd.n3082 vdd.n861 185
R16710 vdd.n861 vdd.n858 185
R16711 vdd.n3084 vdd.n3083 185
R16712 vdd.n3085 vdd.n3084 185
R16713 vdd.n851 vdd.n850 185
R16714 vdd.n852 vdd.n851 185
R16715 vdd.n3093 vdd.n3092 185
R16716 vdd.n3092 vdd.n3091 185
R16717 vdd.n3094 vdd.n849 185
R16718 vdd.n849 vdd.n845 185
R16719 vdd.n3096 vdd.n3095 185
R16720 vdd.n3097 vdd.n3096 185
R16721 vdd.n838 vdd.n837 185
R16722 vdd.n848 vdd.n838 185
R16723 vdd.n3105 vdd.n3104 185
R16724 vdd.n3104 vdd.n3103 185
R16725 vdd.n3106 vdd.n836 185
R16726 vdd.n841 vdd.n836 185
R16727 vdd.n3108 vdd.n3107 185
R16728 vdd.n3109 vdd.n3108 185
R16729 vdd.n827 vdd.n826 185
R16730 vdd.n835 vdd.n827 185
R16731 vdd.n3117 vdd.n3116 185
R16732 vdd.n3116 vdd.n3115 185
R16733 vdd.n3118 vdd.n825 185
R16734 vdd.n825 vdd.n822 185
R16735 vdd.n3120 vdd.n3119 185
R16736 vdd.n3121 vdd.n3120 185
R16737 vdd.n813 vdd.n812 185
R16738 vdd.n814 vdd.n813 185
R16739 vdd.n3174 vdd.n3173 185
R16740 vdd.n3173 vdd.n3172 185
R16741 vdd.n3175 vdd.n811 185
R16742 vdd.n817 vdd.n811 185
R16743 vdd.n3177 vdd.n3176 185
R16744 vdd.n3178 vdd.n3177 185
R16745 vdd.n779 vdd.n777 185
R16746 vdd.n777 vdd.n774 185
R16747 vdd.n3247 vdd.n3246 185
R16748 vdd.n3248 vdd.n3247 185
R16749 vdd.n2628 vdd.n2627 185
R16750 vdd.n2629 vdd.n2628 185
R16751 vdd.n980 vdd.n978 185
R16752 vdd.n978 vdd.n976 185
R16753 vdd.n2543 vdd.n987 185
R16754 vdd.n2554 vdd.n987 185
R16755 vdd.n2544 vdd.n996 185
R16756 vdd.n1370 vdd.n996 185
R16757 vdd.n2546 vdd.n2545 185
R16758 vdd.n2547 vdd.n2546 185
R16759 vdd.n2542 vdd.n995 185
R16760 vdd.n995 vdd.n992 185
R16761 vdd.n2541 vdd.n2540 185
R16762 vdd.n2540 vdd.n2539 185
R16763 vdd.n998 vdd.n997 185
R16764 vdd.n999 vdd.n998 185
R16765 vdd.n2532 vdd.n2531 185
R16766 vdd.n2533 vdd.n2532 185
R16767 vdd.n2530 vdd.n1007 185
R16768 vdd.n1396 vdd.n1007 185
R16769 vdd.n2529 vdd.n2528 185
R16770 vdd.n2528 vdd.n2527 185
R16771 vdd.n1009 vdd.n1008 185
R16772 vdd.n1017 vdd.n1009 185
R16773 vdd.n2520 vdd.n2519 185
R16774 vdd.n2521 vdd.n2520 185
R16775 vdd.n2518 vdd.n1018 185
R16776 vdd.n1023 vdd.n1018 185
R16777 vdd.n2517 vdd.n2516 185
R16778 vdd.n2516 vdd.n2515 185
R16779 vdd.n1020 vdd.n1019 185
R16780 vdd.n1408 vdd.n1020 185
R16781 vdd.n2508 vdd.n2507 185
R16782 vdd.n2509 vdd.n2508 185
R16783 vdd.n2506 vdd.n1030 185
R16784 vdd.n1030 vdd.n1027 185
R16785 vdd.n2505 vdd.n2504 185
R16786 vdd.n2504 vdd.n2503 185
R16787 vdd.n1032 vdd.n1031 185
R16788 vdd.n1033 vdd.n1032 185
R16789 vdd.n2496 vdd.n2495 185
R16790 vdd.n2497 vdd.n2496 185
R16791 vdd.n2493 vdd.n1041 185
R16792 vdd.n1047 vdd.n1041 185
R16793 vdd.n2492 vdd.n2491 185
R16794 vdd.n2491 vdd.n2490 185
R16795 vdd.n1044 vdd.n1043 185
R16796 vdd.n1054 vdd.n1044 185
R16797 vdd.n2483 vdd.n2482 185
R16798 vdd.n2484 vdd.n2483 185
R16799 vdd.n2481 vdd.n1055 185
R16800 vdd.n1055 vdd.n1051 185
R16801 vdd.n2480 vdd.n2479 185
R16802 vdd.n2479 vdd.n2478 185
R16803 vdd.n1057 vdd.n1056 185
R16804 vdd.n1058 vdd.n1057 185
R16805 vdd.n2471 vdd.n2470 185
R16806 vdd.n2472 vdd.n2471 185
R16807 vdd.n2469 vdd.n1067 185
R16808 vdd.n1067 vdd.n1064 185
R16809 vdd.n2468 vdd.n2467 185
R16810 vdd.n2467 vdd.n2466 185
R16811 vdd.n1069 vdd.n1068 185
R16812 vdd.n1077 vdd.n1069 185
R16813 vdd.n2459 vdd.n2458 185
R16814 vdd.n2460 vdd.n2459 185
R16815 vdd.n2457 vdd.n1078 185
R16816 vdd.n1083 vdd.n1078 185
R16817 vdd.n2456 vdd.n2455 185
R16818 vdd.n2455 vdd.n2454 185
R16819 vdd.n1080 vdd.n1079 185
R16820 vdd.n1090 vdd.n1080 185
R16821 vdd.n2447 vdd.n2446 185
R16822 vdd.n2448 vdd.n2447 185
R16823 vdd.n2445 vdd.n1091 185
R16824 vdd.n1091 vdd.n1087 185
R16825 vdd.n2444 vdd.n2443 185
R16826 vdd.n2443 vdd.n2442 185
R16827 vdd.n1093 vdd.n1092 185
R16828 vdd.n1094 vdd.n1093 185
R16829 vdd.n2435 vdd.n2434 185
R16830 vdd.n2436 vdd.n2435 185
R16831 vdd.n2433 vdd.n1102 185
R16832 vdd.n1108 vdd.n1102 185
R16833 vdd.n2432 vdd.n2431 185
R16834 vdd.n2431 vdd.n2430 185
R16835 vdd.n1104 vdd.n1103 185
R16836 vdd.n1105 vdd.n1104 185
R16837 vdd.n2559 vdd.n951 185
R16838 vdd.n2701 vdd.n951 185
R16839 vdd.n2561 vdd.n2560 185
R16840 vdd.n2563 vdd.n2562 185
R16841 vdd.n2565 vdd.n2564 185
R16842 vdd.n2567 vdd.n2566 185
R16843 vdd.n2569 vdd.n2568 185
R16844 vdd.n2571 vdd.n2570 185
R16845 vdd.n2573 vdd.n2572 185
R16846 vdd.n2575 vdd.n2574 185
R16847 vdd.n2577 vdd.n2576 185
R16848 vdd.n2579 vdd.n2578 185
R16849 vdd.n2581 vdd.n2580 185
R16850 vdd.n2583 vdd.n2582 185
R16851 vdd.n2585 vdd.n2584 185
R16852 vdd.n2587 vdd.n2586 185
R16853 vdd.n2589 vdd.n2588 185
R16854 vdd.n2591 vdd.n2590 185
R16855 vdd.n2593 vdd.n2592 185
R16856 vdd.n2595 vdd.n2594 185
R16857 vdd.n2597 vdd.n2596 185
R16858 vdd.n2599 vdd.n2598 185
R16859 vdd.n2601 vdd.n2600 185
R16860 vdd.n2603 vdd.n2602 185
R16861 vdd.n2605 vdd.n2604 185
R16862 vdd.n2607 vdd.n2606 185
R16863 vdd.n2609 vdd.n2608 185
R16864 vdd.n2611 vdd.n2610 185
R16865 vdd.n2613 vdd.n2612 185
R16866 vdd.n2615 vdd.n2614 185
R16867 vdd.n2617 vdd.n2616 185
R16868 vdd.n2619 vdd.n2618 185
R16869 vdd.n2621 vdd.n2620 185
R16870 vdd.n2623 vdd.n2622 185
R16871 vdd.n2625 vdd.n2624 185
R16872 vdd.n2626 vdd.n979 185
R16873 vdd.n2558 vdd.n977 185
R16874 vdd.n2629 vdd.n977 185
R16875 vdd.n2557 vdd.n2556 185
R16876 vdd.n2556 vdd.n976 185
R16877 vdd.n2555 vdd.n984 185
R16878 vdd.n2555 vdd.n2554 185
R16879 vdd.n1386 vdd.n985 185
R16880 vdd.n1370 vdd.n985 185
R16881 vdd.n1387 vdd.n994 185
R16882 vdd.n2547 vdd.n994 185
R16883 vdd.n1389 vdd.n1388 185
R16884 vdd.n1388 vdd.n992 185
R16885 vdd.n1390 vdd.n1001 185
R16886 vdd.n2539 vdd.n1001 185
R16887 vdd.n1392 vdd.n1391 185
R16888 vdd.n1391 vdd.n999 185
R16889 vdd.n1393 vdd.n1006 185
R16890 vdd.n2533 vdd.n1006 185
R16891 vdd.n1395 vdd.n1394 185
R16892 vdd.n1396 vdd.n1395 185
R16893 vdd.n1385 vdd.n1011 185
R16894 vdd.n2527 vdd.n1011 185
R16895 vdd.n1384 vdd.n1383 185
R16896 vdd.n1383 vdd.n1017 185
R16897 vdd.n1382 vdd.n1016 185
R16898 vdd.n2521 vdd.n1016 185
R16899 vdd.n1381 vdd.n1380 185
R16900 vdd.n1380 vdd.n1023 185
R16901 vdd.n1289 vdd.n1022 185
R16902 vdd.n2515 vdd.n1022 185
R16903 vdd.n1410 vdd.n1409 185
R16904 vdd.n1409 vdd.n1408 185
R16905 vdd.n1411 vdd.n1029 185
R16906 vdd.n2509 vdd.n1029 185
R16907 vdd.n1413 vdd.n1412 185
R16908 vdd.n1412 vdd.n1027 185
R16909 vdd.n1414 vdd.n1035 185
R16910 vdd.n2503 vdd.n1035 185
R16911 vdd.n1416 vdd.n1415 185
R16912 vdd.n1415 vdd.n1033 185
R16913 vdd.n1417 vdd.n1040 185
R16914 vdd.n2497 vdd.n1040 185
R16915 vdd.n1419 vdd.n1418 185
R16916 vdd.n1418 vdd.n1047 185
R16917 vdd.n1420 vdd.n1046 185
R16918 vdd.n2490 vdd.n1046 185
R16919 vdd.n1422 vdd.n1421 185
R16920 vdd.n1421 vdd.n1054 185
R16921 vdd.n1423 vdd.n1053 185
R16922 vdd.n2484 vdd.n1053 185
R16923 vdd.n1425 vdd.n1424 185
R16924 vdd.n1424 vdd.n1051 185
R16925 vdd.n1426 vdd.n1060 185
R16926 vdd.n2478 vdd.n1060 185
R16927 vdd.n1428 vdd.n1427 185
R16928 vdd.n1427 vdd.n1058 185
R16929 vdd.n1429 vdd.n1066 185
R16930 vdd.n2472 vdd.n1066 185
R16931 vdd.n1431 vdd.n1430 185
R16932 vdd.n1430 vdd.n1064 185
R16933 vdd.n1432 vdd.n1071 185
R16934 vdd.n2466 vdd.n1071 185
R16935 vdd.n1434 vdd.n1433 185
R16936 vdd.n1433 vdd.n1077 185
R16937 vdd.n1435 vdd.n1076 185
R16938 vdd.n2460 vdd.n1076 185
R16939 vdd.n1437 vdd.n1436 185
R16940 vdd.n1436 vdd.n1083 185
R16941 vdd.n1438 vdd.n1082 185
R16942 vdd.n2454 vdd.n1082 185
R16943 vdd.n1440 vdd.n1439 185
R16944 vdd.n1439 vdd.n1090 185
R16945 vdd.n1441 vdd.n1089 185
R16946 vdd.n2448 vdd.n1089 185
R16947 vdd.n1443 vdd.n1442 185
R16948 vdd.n1442 vdd.n1087 185
R16949 vdd.n1444 vdd.n1096 185
R16950 vdd.n2442 vdd.n1096 185
R16951 vdd.n1446 vdd.n1445 185
R16952 vdd.n1445 vdd.n1094 185
R16953 vdd.n1447 vdd.n1101 185
R16954 vdd.n2436 vdd.n1101 185
R16955 vdd.n1449 vdd.n1448 185
R16956 vdd.n1448 vdd.n1108 185
R16957 vdd.n1450 vdd.n1107 185
R16958 vdd.n2430 vdd.n1107 185
R16959 vdd.n1452 vdd.n1451 185
R16960 vdd.n1451 vdd.n1105 185
R16961 vdd.n1252 vdd.n1251 185
R16962 vdd.n1254 vdd.n1253 185
R16963 vdd.n1256 vdd.n1255 185
R16964 vdd.n1258 vdd.n1257 185
R16965 vdd.n1260 vdd.n1259 185
R16966 vdd.n1262 vdd.n1261 185
R16967 vdd.n1264 vdd.n1263 185
R16968 vdd.n1266 vdd.n1265 185
R16969 vdd.n1268 vdd.n1267 185
R16970 vdd.n1270 vdd.n1269 185
R16971 vdd.n1272 vdd.n1271 185
R16972 vdd.n1274 vdd.n1273 185
R16973 vdd.n1276 vdd.n1275 185
R16974 vdd.n1278 vdd.n1277 185
R16975 vdd.n1280 vdd.n1279 185
R16976 vdd.n1282 vdd.n1281 185
R16977 vdd.n1284 vdd.n1283 185
R16978 vdd.n1486 vdd.n1285 185
R16979 vdd.n1485 vdd.n1484 185
R16980 vdd.n1483 vdd.n1482 185
R16981 vdd.n1481 vdd.n1480 185
R16982 vdd.n1479 vdd.n1478 185
R16983 vdd.n1477 vdd.n1476 185
R16984 vdd.n1475 vdd.n1474 185
R16985 vdd.n1473 vdd.n1472 185
R16986 vdd.n1471 vdd.n1470 185
R16987 vdd.n1469 vdd.n1468 185
R16988 vdd.n1467 vdd.n1466 185
R16989 vdd.n1465 vdd.n1464 185
R16990 vdd.n1463 vdd.n1462 185
R16991 vdd.n1461 vdd.n1460 185
R16992 vdd.n1459 vdd.n1458 185
R16993 vdd.n1457 vdd.n1456 185
R16994 vdd.n1455 vdd.n1454 185
R16995 vdd.n1453 vdd.n1146 185
R16996 vdd.n2423 vdd.n1146 185
R16997 vdd.n315 vdd.n314 171.744
R16998 vdd.n314 vdd.n313 171.744
R16999 vdd.n313 vdd.n282 171.744
R17000 vdd.n306 vdd.n282 171.744
R17001 vdd.n306 vdd.n305 171.744
R17002 vdd.n305 vdd.n287 171.744
R17003 vdd.n298 vdd.n287 171.744
R17004 vdd.n298 vdd.n297 171.744
R17005 vdd.n297 vdd.n291 171.744
R17006 vdd.n260 vdd.n259 171.744
R17007 vdd.n259 vdd.n258 171.744
R17008 vdd.n258 vdd.n227 171.744
R17009 vdd.n251 vdd.n227 171.744
R17010 vdd.n251 vdd.n250 171.744
R17011 vdd.n250 vdd.n232 171.744
R17012 vdd.n243 vdd.n232 171.744
R17013 vdd.n243 vdd.n242 171.744
R17014 vdd.n242 vdd.n236 171.744
R17015 vdd.n217 vdd.n216 171.744
R17016 vdd.n216 vdd.n215 171.744
R17017 vdd.n215 vdd.n184 171.744
R17018 vdd.n208 vdd.n184 171.744
R17019 vdd.n208 vdd.n207 171.744
R17020 vdd.n207 vdd.n189 171.744
R17021 vdd.n200 vdd.n189 171.744
R17022 vdd.n200 vdd.n199 171.744
R17023 vdd.n199 vdd.n193 171.744
R17024 vdd.n162 vdd.n161 171.744
R17025 vdd.n161 vdd.n160 171.744
R17026 vdd.n160 vdd.n129 171.744
R17027 vdd.n153 vdd.n129 171.744
R17028 vdd.n153 vdd.n152 171.744
R17029 vdd.n152 vdd.n134 171.744
R17030 vdd.n145 vdd.n134 171.744
R17031 vdd.n145 vdd.n144 171.744
R17032 vdd.n144 vdd.n138 171.744
R17033 vdd.n120 vdd.n119 171.744
R17034 vdd.n119 vdd.n118 171.744
R17035 vdd.n118 vdd.n87 171.744
R17036 vdd.n111 vdd.n87 171.744
R17037 vdd.n111 vdd.n110 171.744
R17038 vdd.n110 vdd.n92 171.744
R17039 vdd.n103 vdd.n92 171.744
R17040 vdd.n103 vdd.n102 171.744
R17041 vdd.n102 vdd.n96 171.744
R17042 vdd.n65 vdd.n64 171.744
R17043 vdd.n64 vdd.n63 171.744
R17044 vdd.n63 vdd.n32 171.744
R17045 vdd.n56 vdd.n32 171.744
R17046 vdd.n56 vdd.n55 171.744
R17047 vdd.n55 vdd.n37 171.744
R17048 vdd.n48 vdd.n37 171.744
R17049 vdd.n48 vdd.n47 171.744
R17050 vdd.n47 vdd.n41 171.744
R17051 vdd.n2139 vdd.n2138 171.744
R17052 vdd.n2138 vdd.n2137 171.744
R17053 vdd.n2137 vdd.n2106 171.744
R17054 vdd.n2130 vdd.n2106 171.744
R17055 vdd.n2130 vdd.n2129 171.744
R17056 vdd.n2129 vdd.n2111 171.744
R17057 vdd.n2122 vdd.n2111 171.744
R17058 vdd.n2122 vdd.n2121 171.744
R17059 vdd.n2121 vdd.n2115 171.744
R17060 vdd.n2194 vdd.n2193 171.744
R17061 vdd.n2193 vdd.n2192 171.744
R17062 vdd.n2192 vdd.n2161 171.744
R17063 vdd.n2185 vdd.n2161 171.744
R17064 vdd.n2185 vdd.n2184 171.744
R17065 vdd.n2184 vdd.n2166 171.744
R17066 vdd.n2177 vdd.n2166 171.744
R17067 vdd.n2177 vdd.n2176 171.744
R17068 vdd.n2176 vdd.n2170 171.744
R17069 vdd.n2041 vdd.n2040 171.744
R17070 vdd.n2040 vdd.n2039 171.744
R17071 vdd.n2039 vdd.n2008 171.744
R17072 vdd.n2032 vdd.n2008 171.744
R17073 vdd.n2032 vdd.n2031 171.744
R17074 vdd.n2031 vdd.n2013 171.744
R17075 vdd.n2024 vdd.n2013 171.744
R17076 vdd.n2024 vdd.n2023 171.744
R17077 vdd.n2023 vdd.n2017 171.744
R17078 vdd.n2096 vdd.n2095 171.744
R17079 vdd.n2095 vdd.n2094 171.744
R17080 vdd.n2094 vdd.n2063 171.744
R17081 vdd.n2087 vdd.n2063 171.744
R17082 vdd.n2087 vdd.n2086 171.744
R17083 vdd.n2086 vdd.n2068 171.744
R17084 vdd.n2079 vdd.n2068 171.744
R17085 vdd.n2079 vdd.n2078 171.744
R17086 vdd.n2078 vdd.n2072 171.744
R17087 vdd.n1944 vdd.n1943 171.744
R17088 vdd.n1943 vdd.n1942 171.744
R17089 vdd.n1942 vdd.n1911 171.744
R17090 vdd.n1935 vdd.n1911 171.744
R17091 vdd.n1935 vdd.n1934 171.744
R17092 vdd.n1934 vdd.n1916 171.744
R17093 vdd.n1927 vdd.n1916 171.744
R17094 vdd.n1927 vdd.n1926 171.744
R17095 vdd.n1926 vdd.n1920 171.744
R17096 vdd.n1999 vdd.n1998 171.744
R17097 vdd.n1998 vdd.n1997 171.744
R17098 vdd.n1997 vdd.n1966 171.744
R17099 vdd.n1990 vdd.n1966 171.744
R17100 vdd.n1990 vdd.n1989 171.744
R17101 vdd.n1989 vdd.n1971 171.744
R17102 vdd.n1982 vdd.n1971 171.744
R17103 vdd.n1982 vdd.n1981 171.744
R17104 vdd.n1981 vdd.n1975 171.744
R17105 vdd.n449 vdd.n448 146.341
R17106 vdd.n455 vdd.n454 146.341
R17107 vdd.n459 vdd.n458 146.341
R17108 vdd.n465 vdd.n464 146.341
R17109 vdd.n469 vdd.n468 146.341
R17110 vdd.n475 vdd.n474 146.341
R17111 vdd.n479 vdd.n478 146.341
R17112 vdd.n485 vdd.n484 146.341
R17113 vdd.n489 vdd.n488 146.341
R17114 vdd.n495 vdd.n494 146.341
R17115 vdd.n499 vdd.n498 146.341
R17116 vdd.n505 vdd.n504 146.341
R17117 vdd.n509 vdd.n508 146.341
R17118 vdd.n515 vdd.n514 146.341
R17119 vdd.n519 vdd.n518 146.341
R17120 vdd.n525 vdd.n524 146.341
R17121 vdd.n529 vdd.n528 146.341
R17122 vdd.n535 vdd.n534 146.341
R17123 vdd.n539 vdd.n538 146.341
R17124 vdd.n545 vdd.n544 146.341
R17125 vdd.n549 vdd.n548 146.341
R17126 vdd.n555 vdd.n554 146.341
R17127 vdd.n559 vdd.n558 146.341
R17128 vdd.n565 vdd.n564 146.341
R17129 vdd.n569 vdd.n568 146.341
R17130 vdd.n575 vdd.n574 146.341
R17131 vdd.n579 vdd.n578 146.341
R17132 vdd.n585 vdd.n584 146.341
R17133 vdd.n589 vdd.n588 146.341
R17134 vdd.n595 vdd.n594 146.341
R17135 vdd.n597 vdd.n404 146.341
R17136 vdd.n3418 vdd.n654 146.341
R17137 vdd.n3424 vdd.n654 146.341
R17138 vdd.n3424 vdd.n647 146.341
R17139 vdd.n3434 vdd.n647 146.341
R17140 vdd.n3434 vdd.n643 146.341
R17141 vdd.n3440 vdd.n643 146.341
R17142 vdd.n3440 vdd.n634 146.341
R17143 vdd.n3450 vdd.n634 146.341
R17144 vdd.n3450 vdd.n630 146.341
R17145 vdd.n3456 vdd.n630 146.341
R17146 vdd.n3456 vdd.n623 146.341
R17147 vdd.n3467 vdd.n623 146.341
R17148 vdd.n3467 vdd.n619 146.341
R17149 vdd.n3476 vdd.n619 146.341
R17150 vdd.n3476 vdd.n612 146.341
R17151 vdd.n3486 vdd.n612 146.341
R17152 vdd.n3487 vdd.n3486 146.341
R17153 vdd.n3487 vdd.n329 146.341
R17154 vdd.n330 vdd.n329 146.341
R17155 vdd.n331 vdd.n330 146.341
R17156 vdd.n3494 vdd.n331 146.341
R17157 vdd.n3494 vdd.n339 146.341
R17158 vdd.n340 vdd.n339 146.341
R17159 vdd.n341 vdd.n340 146.341
R17160 vdd.n3501 vdd.n341 146.341
R17161 vdd.n3501 vdd.n350 146.341
R17162 vdd.n351 vdd.n350 146.341
R17163 vdd.n352 vdd.n351 146.341
R17164 vdd.n3509 vdd.n352 146.341
R17165 vdd.n3509 vdd.n360 146.341
R17166 vdd.n361 vdd.n360 146.341
R17167 vdd.n362 vdd.n361 146.341
R17168 vdd.n3516 vdd.n362 146.341
R17169 vdd.n3516 vdd.n371 146.341
R17170 vdd.n372 vdd.n371 146.341
R17171 vdd.n3410 vdd.n3408 146.341
R17172 vdd.n3408 vdd.n3407 146.341
R17173 vdd.n3404 vdd.n3403 146.341
R17174 vdd.n3400 vdd.n3399 146.341
R17175 vdd.n3397 vdd.n669 146.341
R17176 vdd.n3393 vdd.n3391 146.341
R17177 vdd.n3389 vdd.n675 146.341
R17178 vdd.n3385 vdd.n3383 146.341
R17179 vdd.n3381 vdd.n681 146.341
R17180 vdd.n3377 vdd.n3375 146.341
R17181 vdd.n3373 vdd.n689 146.341
R17182 vdd.n3369 vdd.n3367 146.341
R17183 vdd.n3365 vdd.n695 146.341
R17184 vdd.n3361 vdd.n3359 146.341
R17185 vdd.n3357 vdd.n701 146.341
R17186 vdd.n3353 vdd.n3351 146.341
R17187 vdd.n3349 vdd.n707 146.341
R17188 vdd.n3345 vdd.n3343 146.341
R17189 vdd.n3341 vdd.n713 146.341
R17190 vdd.n3337 vdd.n3335 146.341
R17191 vdd.n3333 vdd.n719 146.341
R17192 vdd.n3326 vdd.n728 146.341
R17193 vdd.n3324 vdd.n3323 146.341
R17194 vdd.n3320 vdd.n3319 146.341
R17195 vdd.n3317 vdd.n733 146.341
R17196 vdd.n3313 vdd.n3311 146.341
R17197 vdd.n3309 vdd.n739 146.341
R17198 vdd.n3305 vdd.n3303 146.341
R17199 vdd.n3301 vdd.n745 146.341
R17200 vdd.n3297 vdd.n3295 146.341
R17201 vdd.n3292 vdd.n3291 146.341
R17202 vdd.n3288 vdd.n657 146.341
R17203 vdd.n3416 vdd.n653 146.341
R17204 vdd.n3426 vdd.n653 146.341
R17205 vdd.n3426 vdd.n649 146.341
R17206 vdd.n3432 vdd.n649 146.341
R17207 vdd.n3432 vdd.n641 146.341
R17208 vdd.n3442 vdd.n641 146.341
R17209 vdd.n3442 vdd.n637 146.341
R17210 vdd.n3448 vdd.n637 146.341
R17211 vdd.n3448 vdd.n629 146.341
R17212 vdd.n3459 vdd.n629 146.341
R17213 vdd.n3459 vdd.n625 146.341
R17214 vdd.n3465 vdd.n625 146.341
R17215 vdd.n3465 vdd.n618 146.341
R17216 vdd.n3478 vdd.n618 146.341
R17217 vdd.n3478 vdd.n614 146.341
R17218 vdd.n3484 vdd.n614 146.341
R17219 vdd.n3484 vdd.n326 146.341
R17220 vdd.n3560 vdd.n326 146.341
R17221 vdd.n3560 vdd.n327 146.341
R17222 vdd.n3556 vdd.n327 146.341
R17223 vdd.n3556 vdd.n333 146.341
R17224 vdd.n3552 vdd.n333 146.341
R17225 vdd.n3552 vdd.n338 146.341
R17226 vdd.n3548 vdd.n338 146.341
R17227 vdd.n3548 vdd.n342 146.341
R17228 vdd.n3544 vdd.n342 146.341
R17229 vdd.n3544 vdd.n348 146.341
R17230 vdd.n3540 vdd.n348 146.341
R17231 vdd.n3540 vdd.n353 146.341
R17232 vdd.n3536 vdd.n353 146.341
R17233 vdd.n3536 vdd.n359 146.341
R17234 vdd.n3532 vdd.n359 146.341
R17235 vdd.n3532 vdd.n364 146.341
R17236 vdd.n3528 vdd.n364 146.341
R17237 vdd.n3528 vdd.n370 146.341
R17238 vdd.n2388 vdd.n2387 146.341
R17239 vdd.n2385 vdd.n2382 146.341
R17240 vdd.n2380 vdd.n1156 146.341
R17241 vdd.n2376 vdd.n2375 146.341
R17242 vdd.n2373 vdd.n1160 146.341
R17243 vdd.n2369 vdd.n2368 146.341
R17244 vdd.n2366 vdd.n1167 146.341
R17245 vdd.n2362 vdd.n2361 146.341
R17246 vdd.n2359 vdd.n1174 146.341
R17247 vdd.n1185 vdd.n1182 146.341
R17248 vdd.n2351 vdd.n2350 146.341
R17249 vdd.n2348 vdd.n1187 146.341
R17250 vdd.n2344 vdd.n2343 146.341
R17251 vdd.n2341 vdd.n1193 146.341
R17252 vdd.n2337 vdd.n2336 146.341
R17253 vdd.n2334 vdd.n1200 146.341
R17254 vdd.n2330 vdd.n2329 146.341
R17255 vdd.n2327 vdd.n1207 146.341
R17256 vdd.n2323 vdd.n2322 146.341
R17257 vdd.n2320 vdd.n1214 146.341
R17258 vdd.n1225 vdd.n1222 146.341
R17259 vdd.n2312 vdd.n2311 146.341
R17260 vdd.n2309 vdd.n1227 146.341
R17261 vdd.n2305 vdd.n2304 146.341
R17262 vdd.n2302 vdd.n1233 146.341
R17263 vdd.n2298 vdd.n2297 146.341
R17264 vdd.n2295 vdd.n1240 146.341
R17265 vdd.n2291 vdd.n2290 146.341
R17266 vdd.n2288 vdd.n1247 146.341
R17267 vdd.n1493 vdd.n1491 146.341
R17268 vdd.n1496 vdd.n1495 146.341
R17269 vdd.n1836 vdd.n1600 146.341
R17270 vdd.n1836 vdd.n1592 146.341
R17271 vdd.n1846 vdd.n1592 146.341
R17272 vdd.n1846 vdd.n1588 146.341
R17273 vdd.n1852 vdd.n1588 146.341
R17274 vdd.n1852 vdd.n1580 146.341
R17275 vdd.n1863 vdd.n1580 146.341
R17276 vdd.n1863 vdd.n1576 146.341
R17277 vdd.n1869 vdd.n1576 146.341
R17278 vdd.n1869 vdd.n1570 146.341
R17279 vdd.n1880 vdd.n1570 146.341
R17280 vdd.n1880 vdd.n1566 146.341
R17281 vdd.n1886 vdd.n1566 146.341
R17282 vdd.n1886 vdd.n1557 146.341
R17283 vdd.n1896 vdd.n1557 146.341
R17284 vdd.n1896 vdd.n1553 146.341
R17285 vdd.n1902 vdd.n1553 146.341
R17286 vdd.n1902 vdd.n1546 146.341
R17287 vdd.n2208 vdd.n1546 146.341
R17288 vdd.n2208 vdd.n1542 146.341
R17289 vdd.n2214 vdd.n1542 146.341
R17290 vdd.n2214 vdd.n1535 146.341
R17291 vdd.n2224 vdd.n1535 146.341
R17292 vdd.n2224 vdd.n1531 146.341
R17293 vdd.n2230 vdd.n1531 146.341
R17294 vdd.n2230 vdd.n1523 146.341
R17295 vdd.n2241 vdd.n1523 146.341
R17296 vdd.n2241 vdd.n1519 146.341
R17297 vdd.n2247 vdd.n1519 146.341
R17298 vdd.n2247 vdd.n1513 146.341
R17299 vdd.n2258 vdd.n1513 146.341
R17300 vdd.n2258 vdd.n1508 146.341
R17301 vdd.n2266 vdd.n1508 146.341
R17302 vdd.n2266 vdd.n1498 146.341
R17303 vdd.n2276 vdd.n1498 146.341
R17304 vdd.n1638 vdd.n1637 146.341
R17305 vdd.n1642 vdd.n1637 146.341
R17306 vdd.n1644 vdd.n1643 146.341
R17307 vdd.n1648 vdd.n1647 146.341
R17308 vdd.n1650 vdd.n1649 146.341
R17309 vdd.n1654 vdd.n1653 146.341
R17310 vdd.n1656 vdd.n1655 146.341
R17311 vdd.n1660 vdd.n1659 146.341
R17312 vdd.n1662 vdd.n1661 146.341
R17313 vdd.n1794 vdd.n1793 146.341
R17314 vdd.n1666 vdd.n1665 146.341
R17315 vdd.n1670 vdd.n1669 146.341
R17316 vdd.n1672 vdd.n1671 146.341
R17317 vdd.n1676 vdd.n1675 146.341
R17318 vdd.n1678 vdd.n1677 146.341
R17319 vdd.n1682 vdd.n1681 146.341
R17320 vdd.n1684 vdd.n1683 146.341
R17321 vdd.n1688 vdd.n1687 146.341
R17322 vdd.n1690 vdd.n1689 146.341
R17323 vdd.n1694 vdd.n1693 146.341
R17324 vdd.n1758 vdd.n1695 146.341
R17325 vdd.n1699 vdd.n1698 146.341
R17326 vdd.n1701 vdd.n1700 146.341
R17327 vdd.n1705 vdd.n1704 146.341
R17328 vdd.n1707 vdd.n1706 146.341
R17329 vdd.n1711 vdd.n1710 146.341
R17330 vdd.n1713 vdd.n1712 146.341
R17331 vdd.n1717 vdd.n1716 146.341
R17332 vdd.n1719 vdd.n1718 146.341
R17333 vdd.n1723 vdd.n1722 146.341
R17334 vdd.n1725 vdd.n1724 146.341
R17335 vdd.n1830 vdd.n1606 146.341
R17336 vdd.n1838 vdd.n1598 146.341
R17337 vdd.n1838 vdd.n1594 146.341
R17338 vdd.n1844 vdd.n1594 146.341
R17339 vdd.n1844 vdd.n1586 146.341
R17340 vdd.n1855 vdd.n1586 146.341
R17341 vdd.n1855 vdd.n1582 146.341
R17342 vdd.n1861 vdd.n1582 146.341
R17343 vdd.n1861 vdd.n1575 146.341
R17344 vdd.n1872 vdd.n1575 146.341
R17345 vdd.n1872 vdd.n1571 146.341
R17346 vdd.n1878 vdd.n1571 146.341
R17347 vdd.n1878 vdd.n1564 146.341
R17348 vdd.n1888 vdd.n1564 146.341
R17349 vdd.n1888 vdd.n1560 146.341
R17350 vdd.n1894 vdd.n1560 146.341
R17351 vdd.n1894 vdd.n1552 146.341
R17352 vdd.n1905 vdd.n1552 146.341
R17353 vdd.n1905 vdd.n1548 146.341
R17354 vdd.n2206 vdd.n1548 146.341
R17355 vdd.n2206 vdd.n1541 146.341
R17356 vdd.n2216 vdd.n1541 146.341
R17357 vdd.n2216 vdd.n1537 146.341
R17358 vdd.n2222 vdd.n1537 146.341
R17359 vdd.n2222 vdd.n1529 146.341
R17360 vdd.n2233 vdd.n1529 146.341
R17361 vdd.n2233 vdd.n1525 146.341
R17362 vdd.n2239 vdd.n1525 146.341
R17363 vdd.n2239 vdd.n1518 146.341
R17364 vdd.n2250 vdd.n1518 146.341
R17365 vdd.n2250 vdd.n1514 146.341
R17366 vdd.n2256 vdd.n1514 146.341
R17367 vdd.n2256 vdd.n1506 146.341
R17368 vdd.n2268 vdd.n1506 146.341
R17369 vdd.n2268 vdd.n1501 146.341
R17370 vdd.n2274 vdd.n1501 146.341
R17371 vdd.n1286 vdd.t203 127.284
R17372 vdd.n981 vdd.t247 127.284
R17373 vdd.n1290 vdd.t237 127.284
R17374 vdd.n972 vdd.t270 127.284
R17375 vdd.n867 vdd.t224 127.284
R17376 vdd.n867 vdd.t225 127.284
R17377 vdd.n2740 vdd.t265 127.284
R17378 vdd.n804 vdd.t212 127.284
R17379 vdd.n2737 vdd.t255 127.284
R17380 vdd.n768 vdd.t198 127.284
R17381 vdd.n1042 vdd.t261 127.284
R17382 vdd.n1042 vdd.t262 127.284
R17383 vdd.n22 vdd.n20 117.314
R17384 vdd.n17 vdd.n15 117.314
R17385 vdd.n27 vdd.n26 116.927
R17386 vdd.n24 vdd.n23 116.927
R17387 vdd.n22 vdd.n21 116.927
R17388 vdd.n17 vdd.n16 116.927
R17389 vdd.n19 vdd.n18 116.927
R17390 vdd.n27 vdd.n25 116.927
R17391 vdd.n1287 vdd.t202 111.188
R17392 vdd.n982 vdd.t248 111.188
R17393 vdd.n1291 vdd.t236 111.188
R17394 vdd.n973 vdd.t271 111.188
R17395 vdd.n2741 vdd.t264 111.188
R17396 vdd.n805 vdd.t213 111.188
R17397 vdd.n2738 vdd.t254 111.188
R17398 vdd.n769 vdd.t199 111.188
R17399 vdd.n3011 vdd.n931 99.5127
R17400 vdd.n3011 vdd.n922 99.5127
R17401 vdd.n3019 vdd.n922 99.5127
R17402 vdd.n3019 vdd.n920 99.5127
R17403 vdd.n3023 vdd.n920 99.5127
R17404 vdd.n3023 vdd.n910 99.5127
R17405 vdd.n3031 vdd.n910 99.5127
R17406 vdd.n3031 vdd.n908 99.5127
R17407 vdd.n3035 vdd.n908 99.5127
R17408 vdd.n3035 vdd.n899 99.5127
R17409 vdd.n3043 vdd.n899 99.5127
R17410 vdd.n3043 vdd.n897 99.5127
R17411 vdd.n3047 vdd.n897 99.5127
R17412 vdd.n3047 vdd.n888 99.5127
R17413 vdd.n3055 vdd.n888 99.5127
R17414 vdd.n3055 vdd.n886 99.5127
R17415 vdd.n3059 vdd.n886 99.5127
R17416 vdd.n3059 vdd.n875 99.5127
R17417 vdd.n3068 vdd.n875 99.5127
R17418 vdd.n3068 vdd.n873 99.5127
R17419 vdd.n3072 vdd.n873 99.5127
R17420 vdd.n3072 vdd.n863 99.5127
R17421 vdd.n3080 vdd.n863 99.5127
R17422 vdd.n3080 vdd.n861 99.5127
R17423 vdd.n3084 vdd.n861 99.5127
R17424 vdd.n3084 vdd.n851 99.5127
R17425 vdd.n3092 vdd.n851 99.5127
R17426 vdd.n3092 vdd.n849 99.5127
R17427 vdd.n3096 vdd.n849 99.5127
R17428 vdd.n3096 vdd.n838 99.5127
R17429 vdd.n3104 vdd.n838 99.5127
R17430 vdd.n3104 vdd.n836 99.5127
R17431 vdd.n3108 vdd.n836 99.5127
R17432 vdd.n3108 vdd.n827 99.5127
R17433 vdd.n3116 vdd.n827 99.5127
R17434 vdd.n3116 vdd.n825 99.5127
R17435 vdd.n3120 vdd.n825 99.5127
R17436 vdd.n3120 vdd.n813 99.5127
R17437 vdd.n3173 vdd.n813 99.5127
R17438 vdd.n3173 vdd.n811 99.5127
R17439 vdd.n3177 vdd.n811 99.5127
R17440 vdd.n3177 vdd.n777 99.5127
R17441 vdd.n3247 vdd.n777 99.5127
R17442 vdd.n3243 vdd.n778 99.5127
R17443 vdd.n3241 vdd.n3240 99.5127
R17444 vdd.n3238 vdd.n782 99.5127
R17445 vdd.n3234 vdd.n3233 99.5127
R17446 vdd.n3231 vdd.n785 99.5127
R17447 vdd.n3227 vdd.n3226 99.5127
R17448 vdd.n3224 vdd.n788 99.5127
R17449 vdd.n3220 vdd.n3219 99.5127
R17450 vdd.n3217 vdd.n791 99.5127
R17451 vdd.n3212 vdd.n3211 99.5127
R17452 vdd.n3209 vdd.n794 99.5127
R17453 vdd.n3205 vdd.n3204 99.5127
R17454 vdd.n3202 vdd.n797 99.5127
R17455 vdd.n3198 vdd.n3197 99.5127
R17456 vdd.n3195 vdd.n800 99.5127
R17457 vdd.n3191 vdd.n3190 99.5127
R17458 vdd.n3188 vdd.n803 99.5127
R17459 vdd.n2938 vdd.n929 99.5127
R17460 vdd.n2934 vdd.n929 99.5127
R17461 vdd.n2934 vdd.n923 99.5127
R17462 vdd.n2816 vdd.n923 99.5127
R17463 vdd.n2816 vdd.n918 99.5127
R17464 vdd.n2819 vdd.n918 99.5127
R17465 vdd.n2819 vdd.n912 99.5127
R17466 vdd.n2920 vdd.n912 99.5127
R17467 vdd.n2920 vdd.n906 99.5127
R17468 vdd.n2916 vdd.n906 99.5127
R17469 vdd.n2916 vdd.n900 99.5127
R17470 vdd.n2863 vdd.n900 99.5127
R17471 vdd.n2863 vdd.n894 99.5127
R17472 vdd.n2860 vdd.n894 99.5127
R17473 vdd.n2860 vdd.n889 99.5127
R17474 vdd.n2857 vdd.n889 99.5127
R17475 vdd.n2857 vdd.n884 99.5127
R17476 vdd.n2854 vdd.n884 99.5127
R17477 vdd.n2854 vdd.n877 99.5127
R17478 vdd.n2851 vdd.n877 99.5127
R17479 vdd.n2851 vdd.n870 99.5127
R17480 vdd.n2848 vdd.n870 99.5127
R17481 vdd.n2848 vdd.n864 99.5127
R17482 vdd.n2845 vdd.n864 99.5127
R17483 vdd.n2845 vdd.n859 99.5127
R17484 vdd.n2842 vdd.n859 99.5127
R17485 vdd.n2842 vdd.n853 99.5127
R17486 vdd.n2839 vdd.n853 99.5127
R17487 vdd.n2839 vdd.n846 99.5127
R17488 vdd.n2836 vdd.n846 99.5127
R17489 vdd.n2836 vdd.n839 99.5127
R17490 vdd.n2833 vdd.n839 99.5127
R17491 vdd.n2833 vdd.n833 99.5127
R17492 vdd.n2830 vdd.n833 99.5127
R17493 vdd.n2830 vdd.n828 99.5127
R17494 vdd.n2827 vdd.n828 99.5127
R17495 vdd.n2827 vdd.n823 99.5127
R17496 vdd.n2824 vdd.n823 99.5127
R17497 vdd.n2824 vdd.n815 99.5127
R17498 vdd.n815 vdd.n808 99.5127
R17499 vdd.n3179 vdd.n808 99.5127
R17500 vdd.n3180 vdd.n3179 99.5127
R17501 vdd.n3180 vdd.n775 99.5127
R17502 vdd.n3004 vdd.n933 99.5127
R17503 vdd.n3004 vdd.n2736 99.5127
R17504 vdd.n3000 vdd.n2999 99.5127
R17505 vdd.n2996 vdd.n2995 99.5127
R17506 vdd.n2992 vdd.n2991 99.5127
R17507 vdd.n2988 vdd.n2987 99.5127
R17508 vdd.n2984 vdd.n2983 99.5127
R17509 vdd.n2980 vdd.n2979 99.5127
R17510 vdd.n2976 vdd.n2975 99.5127
R17511 vdd.n2972 vdd.n2971 99.5127
R17512 vdd.n2968 vdd.n2967 99.5127
R17513 vdd.n2964 vdd.n2963 99.5127
R17514 vdd.n2960 vdd.n2959 99.5127
R17515 vdd.n2956 vdd.n2955 99.5127
R17516 vdd.n2952 vdd.n2951 99.5127
R17517 vdd.n2948 vdd.n2947 99.5127
R17518 vdd.n2943 vdd.n2942 99.5127
R17519 vdd.n2700 vdd.n970 99.5127
R17520 vdd.n2696 vdd.n2695 99.5127
R17521 vdd.n2692 vdd.n2691 99.5127
R17522 vdd.n2688 vdd.n2687 99.5127
R17523 vdd.n2684 vdd.n2683 99.5127
R17524 vdd.n2680 vdd.n2679 99.5127
R17525 vdd.n2676 vdd.n2675 99.5127
R17526 vdd.n2672 vdd.n2671 99.5127
R17527 vdd.n2668 vdd.n2667 99.5127
R17528 vdd.n2664 vdd.n2663 99.5127
R17529 vdd.n2660 vdd.n2659 99.5127
R17530 vdd.n2656 vdd.n2655 99.5127
R17531 vdd.n2652 vdd.n2651 99.5127
R17532 vdd.n2648 vdd.n2647 99.5127
R17533 vdd.n2644 vdd.n2643 99.5127
R17534 vdd.n2640 vdd.n2639 99.5127
R17535 vdd.n2635 vdd.n2634 99.5127
R17536 vdd.n1326 vdd.n1106 99.5127
R17537 vdd.n1329 vdd.n1106 99.5127
R17538 vdd.n1329 vdd.n1100 99.5127
R17539 vdd.n1332 vdd.n1100 99.5127
R17540 vdd.n1332 vdd.n1095 99.5127
R17541 vdd.n1335 vdd.n1095 99.5127
R17542 vdd.n1335 vdd.n1088 99.5127
R17543 vdd.n1338 vdd.n1088 99.5127
R17544 vdd.n1338 vdd.n1081 99.5127
R17545 vdd.n1341 vdd.n1081 99.5127
R17546 vdd.n1341 vdd.n1075 99.5127
R17547 vdd.n1344 vdd.n1075 99.5127
R17548 vdd.n1344 vdd.n1070 99.5127
R17549 vdd.n1347 vdd.n1070 99.5127
R17550 vdd.n1347 vdd.n1065 99.5127
R17551 vdd.n1350 vdd.n1065 99.5127
R17552 vdd.n1350 vdd.n1059 99.5127
R17553 vdd.n1353 vdd.n1059 99.5127
R17554 vdd.n1353 vdd.n1052 99.5127
R17555 vdd.n1356 vdd.n1052 99.5127
R17556 vdd.n1356 vdd.n1045 99.5127
R17557 vdd.n1359 vdd.n1045 99.5127
R17558 vdd.n1359 vdd.n1039 99.5127
R17559 vdd.n1362 vdd.n1039 99.5127
R17560 vdd.n1362 vdd.n1034 99.5127
R17561 vdd.n1365 vdd.n1034 99.5127
R17562 vdd.n1365 vdd.n1028 99.5127
R17563 vdd.n1407 vdd.n1028 99.5127
R17564 vdd.n1407 vdd.n1021 99.5127
R17565 vdd.n1403 vdd.n1021 99.5127
R17566 vdd.n1403 vdd.n1015 99.5127
R17567 vdd.n1400 vdd.n1015 99.5127
R17568 vdd.n1400 vdd.n1010 99.5127
R17569 vdd.n1397 vdd.n1010 99.5127
R17570 vdd.n1397 vdd.n1005 99.5127
R17571 vdd.n1377 vdd.n1005 99.5127
R17572 vdd.n1377 vdd.n1000 99.5127
R17573 vdd.n1374 vdd.n1000 99.5127
R17574 vdd.n1374 vdd.n993 99.5127
R17575 vdd.n1371 vdd.n993 99.5127
R17576 vdd.n1371 vdd.n986 99.5127
R17577 vdd.n986 vdd.n975 99.5127
R17578 vdd.n2630 vdd.n975 99.5127
R17579 vdd.n2422 vdd.n1111 99.5127
R17580 vdd.n2422 vdd.n1147 99.5127
R17581 vdd.n2418 vdd.n2417 99.5127
R17582 vdd.n2414 vdd.n2413 99.5127
R17583 vdd.n2410 vdd.n2409 99.5127
R17584 vdd.n2406 vdd.n2405 99.5127
R17585 vdd.n2402 vdd.n2401 99.5127
R17586 vdd.n2398 vdd.n2397 99.5127
R17587 vdd.n2394 vdd.n2393 99.5127
R17588 vdd.n1293 vdd.n1292 99.5127
R17589 vdd.n1297 vdd.n1296 99.5127
R17590 vdd.n1301 vdd.n1300 99.5127
R17591 vdd.n1305 vdd.n1304 99.5127
R17592 vdd.n1309 vdd.n1308 99.5127
R17593 vdd.n1313 vdd.n1312 99.5127
R17594 vdd.n1317 vdd.n1316 99.5127
R17595 vdd.n1322 vdd.n1321 99.5127
R17596 vdd.n2429 vdd.n1109 99.5127
R17597 vdd.n2429 vdd.n1099 99.5127
R17598 vdd.n2437 vdd.n1099 99.5127
R17599 vdd.n2437 vdd.n1097 99.5127
R17600 vdd.n2441 vdd.n1097 99.5127
R17601 vdd.n2441 vdd.n1086 99.5127
R17602 vdd.n2449 vdd.n1086 99.5127
R17603 vdd.n2449 vdd.n1084 99.5127
R17604 vdd.n2453 vdd.n1084 99.5127
R17605 vdd.n2453 vdd.n1074 99.5127
R17606 vdd.n2461 vdd.n1074 99.5127
R17607 vdd.n2461 vdd.n1072 99.5127
R17608 vdd.n2465 vdd.n1072 99.5127
R17609 vdd.n2465 vdd.n1063 99.5127
R17610 vdd.n2473 vdd.n1063 99.5127
R17611 vdd.n2473 vdd.n1061 99.5127
R17612 vdd.n2477 vdd.n1061 99.5127
R17613 vdd.n2477 vdd.n1050 99.5127
R17614 vdd.n2485 vdd.n1050 99.5127
R17615 vdd.n2485 vdd.n1048 99.5127
R17616 vdd.n2489 vdd.n1048 99.5127
R17617 vdd.n2489 vdd.n1038 99.5127
R17618 vdd.n2498 vdd.n1038 99.5127
R17619 vdd.n2498 vdd.n1036 99.5127
R17620 vdd.n2502 vdd.n1036 99.5127
R17621 vdd.n2502 vdd.n1026 99.5127
R17622 vdd.n2510 vdd.n1026 99.5127
R17623 vdd.n2510 vdd.n1024 99.5127
R17624 vdd.n2514 vdd.n1024 99.5127
R17625 vdd.n2514 vdd.n1014 99.5127
R17626 vdd.n2522 vdd.n1014 99.5127
R17627 vdd.n2522 vdd.n1012 99.5127
R17628 vdd.n2526 vdd.n1012 99.5127
R17629 vdd.n2526 vdd.n1004 99.5127
R17630 vdd.n2534 vdd.n1004 99.5127
R17631 vdd.n2534 vdd.n1002 99.5127
R17632 vdd.n2538 vdd.n1002 99.5127
R17633 vdd.n2538 vdd.n991 99.5127
R17634 vdd.n2548 vdd.n991 99.5127
R17635 vdd.n2548 vdd.n988 99.5127
R17636 vdd.n2553 vdd.n988 99.5127
R17637 vdd.n2553 vdd.n989 99.5127
R17638 vdd.n989 vdd.n969 99.5127
R17639 vdd.n3163 vdd.n3162 99.5127
R17640 vdd.n3160 vdd.n3126 99.5127
R17641 vdd.n3156 vdd.n3155 99.5127
R17642 vdd.n3153 vdd.n3129 99.5127
R17643 vdd.n3149 vdd.n3148 99.5127
R17644 vdd.n3146 vdd.n3132 99.5127
R17645 vdd.n3142 vdd.n3141 99.5127
R17646 vdd.n3139 vdd.n3136 99.5127
R17647 vdd.n3280 vdd.n755 99.5127
R17648 vdd.n3278 vdd.n3277 99.5127
R17649 vdd.n3275 vdd.n758 99.5127
R17650 vdd.n3271 vdd.n3270 99.5127
R17651 vdd.n3268 vdd.n761 99.5127
R17652 vdd.n3264 vdd.n3263 99.5127
R17653 vdd.n3261 vdd.n764 99.5127
R17654 vdd.n3257 vdd.n3256 99.5127
R17655 vdd.n3254 vdd.n767 99.5127
R17656 vdd.n2812 vdd.n930 99.5127
R17657 vdd.n2932 vdd.n930 99.5127
R17658 vdd.n2932 vdd.n924 99.5127
R17659 vdd.n2928 vdd.n924 99.5127
R17660 vdd.n2928 vdd.n919 99.5127
R17661 vdd.n2925 vdd.n919 99.5127
R17662 vdd.n2925 vdd.n913 99.5127
R17663 vdd.n2922 vdd.n913 99.5127
R17664 vdd.n2922 vdd.n907 99.5127
R17665 vdd.n2914 vdd.n907 99.5127
R17666 vdd.n2914 vdd.n901 99.5127
R17667 vdd.n2910 vdd.n901 99.5127
R17668 vdd.n2910 vdd.n895 99.5127
R17669 vdd.n2907 vdd.n895 99.5127
R17670 vdd.n2907 vdd.n890 99.5127
R17671 vdd.n2904 vdd.n890 99.5127
R17672 vdd.n2904 vdd.n885 99.5127
R17673 vdd.n2901 vdd.n885 99.5127
R17674 vdd.n2901 vdd.n878 99.5127
R17675 vdd.n2898 vdd.n878 99.5127
R17676 vdd.n2898 vdd.n871 99.5127
R17677 vdd.n2895 vdd.n871 99.5127
R17678 vdd.n2895 vdd.n865 99.5127
R17679 vdd.n2892 vdd.n865 99.5127
R17680 vdd.n2892 vdd.n860 99.5127
R17681 vdd.n2889 vdd.n860 99.5127
R17682 vdd.n2889 vdd.n854 99.5127
R17683 vdd.n2886 vdd.n854 99.5127
R17684 vdd.n2886 vdd.n847 99.5127
R17685 vdd.n2883 vdd.n847 99.5127
R17686 vdd.n2883 vdd.n840 99.5127
R17687 vdd.n2880 vdd.n840 99.5127
R17688 vdd.n2880 vdd.n834 99.5127
R17689 vdd.n2877 vdd.n834 99.5127
R17690 vdd.n2877 vdd.n829 99.5127
R17691 vdd.n2874 vdd.n829 99.5127
R17692 vdd.n2874 vdd.n824 99.5127
R17693 vdd.n2871 vdd.n824 99.5127
R17694 vdd.n2871 vdd.n816 99.5127
R17695 vdd.n2868 vdd.n816 99.5127
R17696 vdd.n2868 vdd.n809 99.5127
R17697 vdd.n809 vdd.n773 99.5127
R17698 vdd.n3249 vdd.n773 99.5127
R17699 vdd.n2747 vdd.n2746 99.5127
R17700 vdd.n2751 vdd.n2750 99.5127
R17701 vdd.n2755 vdd.n2754 99.5127
R17702 vdd.n2759 vdd.n2758 99.5127
R17703 vdd.n2763 vdd.n2762 99.5127
R17704 vdd.n2767 vdd.n2766 99.5127
R17705 vdd.n2771 vdd.n2770 99.5127
R17706 vdd.n2775 vdd.n2774 99.5127
R17707 vdd.n2779 vdd.n2778 99.5127
R17708 vdd.n2783 vdd.n2782 99.5127
R17709 vdd.n2787 vdd.n2786 99.5127
R17710 vdd.n2791 vdd.n2790 99.5127
R17711 vdd.n2795 vdd.n2794 99.5127
R17712 vdd.n2799 vdd.n2798 99.5127
R17713 vdd.n2803 vdd.n2802 99.5127
R17714 vdd.n2807 vdd.n2806 99.5127
R17715 vdd.n2809 vdd.n2735 99.5127
R17716 vdd.n3013 vdd.n927 99.5127
R17717 vdd.n3013 vdd.n925 99.5127
R17718 vdd.n3017 vdd.n925 99.5127
R17719 vdd.n3017 vdd.n916 99.5127
R17720 vdd.n3025 vdd.n916 99.5127
R17721 vdd.n3025 vdd.n914 99.5127
R17722 vdd.n3029 vdd.n914 99.5127
R17723 vdd.n3029 vdd.n905 99.5127
R17724 vdd.n3037 vdd.n905 99.5127
R17725 vdd.n3037 vdd.n903 99.5127
R17726 vdd.n3041 vdd.n903 99.5127
R17727 vdd.n3041 vdd.n893 99.5127
R17728 vdd.n3049 vdd.n893 99.5127
R17729 vdd.n3049 vdd.n891 99.5127
R17730 vdd.n3053 vdd.n891 99.5127
R17731 vdd.n3053 vdd.n882 99.5127
R17732 vdd.n3061 vdd.n882 99.5127
R17733 vdd.n3061 vdd.n880 99.5127
R17734 vdd.n3066 vdd.n880 99.5127
R17735 vdd.n3066 vdd.n869 99.5127
R17736 vdd.n3074 vdd.n869 99.5127
R17737 vdd.n3074 vdd.n866 99.5127
R17738 vdd.n3078 vdd.n866 99.5127
R17739 vdd.n3078 vdd.n857 99.5127
R17740 vdd.n3086 vdd.n857 99.5127
R17741 vdd.n3086 vdd.n855 99.5127
R17742 vdd.n3090 vdd.n855 99.5127
R17743 vdd.n3090 vdd.n844 99.5127
R17744 vdd.n3098 vdd.n844 99.5127
R17745 vdd.n3098 vdd.n842 99.5127
R17746 vdd.n3102 vdd.n842 99.5127
R17747 vdd.n3102 vdd.n832 99.5127
R17748 vdd.n3110 vdd.n832 99.5127
R17749 vdd.n3110 vdd.n830 99.5127
R17750 vdd.n3114 vdd.n830 99.5127
R17751 vdd.n3114 vdd.n821 99.5127
R17752 vdd.n3122 vdd.n821 99.5127
R17753 vdd.n3122 vdd.n818 99.5127
R17754 vdd.n3171 vdd.n818 99.5127
R17755 vdd.n3171 vdd.n819 99.5127
R17756 vdd.n819 vdd.n810 99.5127
R17757 vdd.n3166 vdd.n810 99.5127
R17758 vdd.n3166 vdd.n776 99.5127
R17759 vdd.n2624 vdd.n2623 99.5127
R17760 vdd.n2620 vdd.n2619 99.5127
R17761 vdd.n2616 vdd.n2615 99.5127
R17762 vdd.n2612 vdd.n2611 99.5127
R17763 vdd.n2608 vdd.n2607 99.5127
R17764 vdd.n2604 vdd.n2603 99.5127
R17765 vdd.n2600 vdd.n2599 99.5127
R17766 vdd.n2596 vdd.n2595 99.5127
R17767 vdd.n2592 vdd.n2591 99.5127
R17768 vdd.n2588 vdd.n2587 99.5127
R17769 vdd.n2584 vdd.n2583 99.5127
R17770 vdd.n2580 vdd.n2579 99.5127
R17771 vdd.n2576 vdd.n2575 99.5127
R17772 vdd.n2572 vdd.n2571 99.5127
R17773 vdd.n2568 vdd.n2567 99.5127
R17774 vdd.n2564 vdd.n2563 99.5127
R17775 vdd.n2560 vdd.n951 99.5127
R17776 vdd.n1451 vdd.n1107 99.5127
R17777 vdd.n1448 vdd.n1107 99.5127
R17778 vdd.n1448 vdd.n1101 99.5127
R17779 vdd.n1445 vdd.n1101 99.5127
R17780 vdd.n1445 vdd.n1096 99.5127
R17781 vdd.n1442 vdd.n1096 99.5127
R17782 vdd.n1442 vdd.n1089 99.5127
R17783 vdd.n1439 vdd.n1089 99.5127
R17784 vdd.n1439 vdd.n1082 99.5127
R17785 vdd.n1436 vdd.n1082 99.5127
R17786 vdd.n1436 vdd.n1076 99.5127
R17787 vdd.n1433 vdd.n1076 99.5127
R17788 vdd.n1433 vdd.n1071 99.5127
R17789 vdd.n1430 vdd.n1071 99.5127
R17790 vdd.n1430 vdd.n1066 99.5127
R17791 vdd.n1427 vdd.n1066 99.5127
R17792 vdd.n1427 vdd.n1060 99.5127
R17793 vdd.n1424 vdd.n1060 99.5127
R17794 vdd.n1424 vdd.n1053 99.5127
R17795 vdd.n1421 vdd.n1053 99.5127
R17796 vdd.n1421 vdd.n1046 99.5127
R17797 vdd.n1418 vdd.n1046 99.5127
R17798 vdd.n1418 vdd.n1040 99.5127
R17799 vdd.n1415 vdd.n1040 99.5127
R17800 vdd.n1415 vdd.n1035 99.5127
R17801 vdd.n1412 vdd.n1035 99.5127
R17802 vdd.n1412 vdd.n1029 99.5127
R17803 vdd.n1409 vdd.n1029 99.5127
R17804 vdd.n1409 vdd.n1022 99.5127
R17805 vdd.n1380 vdd.n1022 99.5127
R17806 vdd.n1380 vdd.n1016 99.5127
R17807 vdd.n1383 vdd.n1016 99.5127
R17808 vdd.n1383 vdd.n1011 99.5127
R17809 vdd.n1395 vdd.n1011 99.5127
R17810 vdd.n1395 vdd.n1006 99.5127
R17811 vdd.n1391 vdd.n1006 99.5127
R17812 vdd.n1391 vdd.n1001 99.5127
R17813 vdd.n1388 vdd.n1001 99.5127
R17814 vdd.n1388 vdd.n994 99.5127
R17815 vdd.n994 vdd.n985 99.5127
R17816 vdd.n2555 vdd.n985 99.5127
R17817 vdd.n2556 vdd.n2555 99.5127
R17818 vdd.n2556 vdd.n977 99.5127
R17819 vdd.n1255 vdd.n1254 99.5127
R17820 vdd.n1259 vdd.n1258 99.5127
R17821 vdd.n1263 vdd.n1262 99.5127
R17822 vdd.n1267 vdd.n1266 99.5127
R17823 vdd.n1271 vdd.n1270 99.5127
R17824 vdd.n1275 vdd.n1274 99.5127
R17825 vdd.n1279 vdd.n1278 99.5127
R17826 vdd.n1283 vdd.n1282 99.5127
R17827 vdd.n1484 vdd.n1285 99.5127
R17828 vdd.n1482 vdd.n1481 99.5127
R17829 vdd.n1478 vdd.n1477 99.5127
R17830 vdd.n1474 vdd.n1473 99.5127
R17831 vdd.n1470 vdd.n1469 99.5127
R17832 vdd.n1466 vdd.n1465 99.5127
R17833 vdd.n1462 vdd.n1461 99.5127
R17834 vdd.n1458 vdd.n1457 99.5127
R17835 vdd.n1454 vdd.n1146 99.5127
R17836 vdd.n2431 vdd.n1104 99.5127
R17837 vdd.n2431 vdd.n1102 99.5127
R17838 vdd.n2435 vdd.n1102 99.5127
R17839 vdd.n2435 vdd.n1093 99.5127
R17840 vdd.n2443 vdd.n1093 99.5127
R17841 vdd.n2443 vdd.n1091 99.5127
R17842 vdd.n2447 vdd.n1091 99.5127
R17843 vdd.n2447 vdd.n1080 99.5127
R17844 vdd.n2455 vdd.n1080 99.5127
R17845 vdd.n2455 vdd.n1078 99.5127
R17846 vdd.n2459 vdd.n1078 99.5127
R17847 vdd.n2459 vdd.n1069 99.5127
R17848 vdd.n2467 vdd.n1069 99.5127
R17849 vdd.n2467 vdd.n1067 99.5127
R17850 vdd.n2471 vdd.n1067 99.5127
R17851 vdd.n2471 vdd.n1057 99.5127
R17852 vdd.n2479 vdd.n1057 99.5127
R17853 vdd.n2479 vdd.n1055 99.5127
R17854 vdd.n2483 vdd.n1055 99.5127
R17855 vdd.n2483 vdd.n1044 99.5127
R17856 vdd.n2491 vdd.n1044 99.5127
R17857 vdd.n2491 vdd.n1041 99.5127
R17858 vdd.n2496 vdd.n1041 99.5127
R17859 vdd.n2496 vdd.n1032 99.5127
R17860 vdd.n2504 vdd.n1032 99.5127
R17861 vdd.n2504 vdd.n1030 99.5127
R17862 vdd.n2508 vdd.n1030 99.5127
R17863 vdd.n2508 vdd.n1020 99.5127
R17864 vdd.n2516 vdd.n1020 99.5127
R17865 vdd.n2516 vdd.n1018 99.5127
R17866 vdd.n2520 vdd.n1018 99.5127
R17867 vdd.n2520 vdd.n1009 99.5127
R17868 vdd.n2528 vdd.n1009 99.5127
R17869 vdd.n2528 vdd.n1007 99.5127
R17870 vdd.n2532 vdd.n1007 99.5127
R17871 vdd.n2532 vdd.n998 99.5127
R17872 vdd.n2540 vdd.n998 99.5127
R17873 vdd.n2540 vdd.n995 99.5127
R17874 vdd.n2546 vdd.n995 99.5127
R17875 vdd.n2546 vdd.n996 99.5127
R17876 vdd.n996 vdd.n987 99.5127
R17877 vdd.n987 vdd.n978 99.5127
R17878 vdd.n2628 vdd.n978 99.5127
R17879 vdd.n9 vdd.n7 98.9633
R17880 vdd.n2 vdd.n0 98.9633
R17881 vdd.n9 vdd.n8 98.6055
R17882 vdd.n11 vdd.n10 98.6055
R17883 vdd.n13 vdd.n12 98.6055
R17884 vdd.n6 vdd.n5 98.6055
R17885 vdd.n4 vdd.n3 98.6055
R17886 vdd.n2 vdd.n1 98.6055
R17887 vdd.t88 vdd.n291 85.8723
R17888 vdd.t177 vdd.n236 85.8723
R17889 vdd.t71 vdd.n193 85.8723
R17890 vdd.t169 vdd.n138 85.8723
R17891 vdd.t137 vdd.n96 85.8723
R17892 vdd.t122 vdd.n41 85.8723
R17893 vdd.t107 vdd.n2115 85.8723
R17894 vdd.t135 vdd.n2170 85.8723
R17895 vdd.t90 vdd.n2017 85.8723
R17896 vdd.t124 vdd.n2072 85.8723
R17897 vdd.t126 vdd.n1920 85.8723
R17898 vdd.t139 vdd.n1975 85.8723
R17899 vdd.n868 vdd.n867 78.546
R17900 vdd.n2494 vdd.n1042 78.546
R17901 vdd.n278 vdd.n277 75.1835
R17902 vdd.n276 vdd.n275 75.1835
R17903 vdd.n274 vdd.n273 75.1835
R17904 vdd.n272 vdd.n271 75.1835
R17905 vdd.n270 vdd.n269 75.1835
R17906 vdd.n268 vdd.n267 75.1835
R17907 vdd.n266 vdd.n265 75.1835
R17908 vdd.n180 vdd.n179 75.1835
R17909 vdd.n178 vdd.n177 75.1835
R17910 vdd.n176 vdd.n175 75.1835
R17911 vdd.n174 vdd.n173 75.1835
R17912 vdd.n172 vdd.n171 75.1835
R17913 vdd.n170 vdd.n169 75.1835
R17914 vdd.n168 vdd.n167 75.1835
R17915 vdd.n83 vdd.n82 75.1835
R17916 vdd.n81 vdd.n80 75.1835
R17917 vdd.n79 vdd.n78 75.1835
R17918 vdd.n77 vdd.n76 75.1835
R17919 vdd.n75 vdd.n74 75.1835
R17920 vdd.n73 vdd.n72 75.1835
R17921 vdd.n71 vdd.n70 75.1835
R17922 vdd.n2145 vdd.n2144 75.1835
R17923 vdd.n2147 vdd.n2146 75.1835
R17924 vdd.n2149 vdd.n2148 75.1835
R17925 vdd.n2151 vdd.n2150 75.1835
R17926 vdd.n2153 vdd.n2152 75.1835
R17927 vdd.n2155 vdd.n2154 75.1835
R17928 vdd.n2157 vdd.n2156 75.1835
R17929 vdd.n2047 vdd.n2046 75.1835
R17930 vdd.n2049 vdd.n2048 75.1835
R17931 vdd.n2051 vdd.n2050 75.1835
R17932 vdd.n2053 vdd.n2052 75.1835
R17933 vdd.n2055 vdd.n2054 75.1835
R17934 vdd.n2057 vdd.n2056 75.1835
R17935 vdd.n2059 vdd.n2058 75.1835
R17936 vdd.n1950 vdd.n1949 75.1835
R17937 vdd.n1952 vdd.n1951 75.1835
R17938 vdd.n1954 vdd.n1953 75.1835
R17939 vdd.n1956 vdd.n1955 75.1835
R17940 vdd.n1958 vdd.n1957 75.1835
R17941 vdd.n1960 vdd.n1959 75.1835
R17942 vdd.n1962 vdd.n1961 75.1835
R17943 vdd.n3005 vdd.n2718 72.8958
R17944 vdd.n3005 vdd.n2719 72.8958
R17945 vdd.n3005 vdd.n2720 72.8958
R17946 vdd.n3005 vdd.n2721 72.8958
R17947 vdd.n3005 vdd.n2722 72.8958
R17948 vdd.n3005 vdd.n2723 72.8958
R17949 vdd.n3005 vdd.n2724 72.8958
R17950 vdd.n3005 vdd.n2725 72.8958
R17951 vdd.n3005 vdd.n2726 72.8958
R17952 vdd.n3005 vdd.n2727 72.8958
R17953 vdd.n3005 vdd.n2728 72.8958
R17954 vdd.n3005 vdd.n2729 72.8958
R17955 vdd.n3005 vdd.n2730 72.8958
R17956 vdd.n3005 vdd.n2731 72.8958
R17957 vdd.n3005 vdd.n2732 72.8958
R17958 vdd.n3005 vdd.n2733 72.8958
R17959 vdd.n3005 vdd.n2734 72.8958
R17960 vdd.n772 vdd.n756 72.8958
R17961 vdd.n3255 vdd.n756 72.8958
R17962 vdd.n766 vdd.n756 72.8958
R17963 vdd.n3262 vdd.n756 72.8958
R17964 vdd.n763 vdd.n756 72.8958
R17965 vdd.n3269 vdd.n756 72.8958
R17966 vdd.n760 vdd.n756 72.8958
R17967 vdd.n3276 vdd.n756 72.8958
R17968 vdd.n3279 vdd.n756 72.8958
R17969 vdd.n3135 vdd.n756 72.8958
R17970 vdd.n3140 vdd.n756 72.8958
R17971 vdd.n3134 vdd.n756 72.8958
R17972 vdd.n3147 vdd.n756 72.8958
R17973 vdd.n3131 vdd.n756 72.8958
R17974 vdd.n3154 vdd.n756 72.8958
R17975 vdd.n3128 vdd.n756 72.8958
R17976 vdd.n3161 vdd.n756 72.8958
R17977 vdd.n2424 vdd.n2423 72.8958
R17978 vdd.n2423 vdd.n1113 72.8958
R17979 vdd.n2423 vdd.n1114 72.8958
R17980 vdd.n2423 vdd.n1115 72.8958
R17981 vdd.n2423 vdd.n1116 72.8958
R17982 vdd.n2423 vdd.n1117 72.8958
R17983 vdd.n2423 vdd.n1118 72.8958
R17984 vdd.n2423 vdd.n1119 72.8958
R17985 vdd.n2423 vdd.n1120 72.8958
R17986 vdd.n2423 vdd.n1121 72.8958
R17987 vdd.n2423 vdd.n1122 72.8958
R17988 vdd.n2423 vdd.n1123 72.8958
R17989 vdd.n2423 vdd.n1124 72.8958
R17990 vdd.n2423 vdd.n1125 72.8958
R17991 vdd.n2423 vdd.n1126 72.8958
R17992 vdd.n2423 vdd.n1127 72.8958
R17993 vdd.n2423 vdd.n1128 72.8958
R17994 vdd.n2701 vdd.n952 72.8958
R17995 vdd.n2701 vdd.n953 72.8958
R17996 vdd.n2701 vdd.n954 72.8958
R17997 vdd.n2701 vdd.n955 72.8958
R17998 vdd.n2701 vdd.n956 72.8958
R17999 vdd.n2701 vdd.n957 72.8958
R18000 vdd.n2701 vdd.n958 72.8958
R18001 vdd.n2701 vdd.n959 72.8958
R18002 vdd.n2701 vdd.n960 72.8958
R18003 vdd.n2701 vdd.n961 72.8958
R18004 vdd.n2701 vdd.n962 72.8958
R18005 vdd.n2701 vdd.n963 72.8958
R18006 vdd.n2701 vdd.n964 72.8958
R18007 vdd.n2701 vdd.n965 72.8958
R18008 vdd.n2701 vdd.n966 72.8958
R18009 vdd.n2701 vdd.n967 72.8958
R18010 vdd.n2701 vdd.n968 72.8958
R18011 vdd.n3006 vdd.n3005 72.8958
R18012 vdd.n3005 vdd.n2702 72.8958
R18013 vdd.n3005 vdd.n2703 72.8958
R18014 vdd.n3005 vdd.n2704 72.8958
R18015 vdd.n3005 vdd.n2705 72.8958
R18016 vdd.n3005 vdd.n2706 72.8958
R18017 vdd.n3005 vdd.n2707 72.8958
R18018 vdd.n3005 vdd.n2708 72.8958
R18019 vdd.n3005 vdd.n2709 72.8958
R18020 vdd.n3005 vdd.n2710 72.8958
R18021 vdd.n3005 vdd.n2711 72.8958
R18022 vdd.n3005 vdd.n2712 72.8958
R18023 vdd.n3005 vdd.n2713 72.8958
R18024 vdd.n3005 vdd.n2714 72.8958
R18025 vdd.n3005 vdd.n2715 72.8958
R18026 vdd.n3005 vdd.n2716 72.8958
R18027 vdd.n3005 vdd.n2717 72.8958
R18028 vdd.n3183 vdd.n756 72.8958
R18029 vdd.n3189 vdd.n756 72.8958
R18030 vdd.n802 vdd.n756 72.8958
R18031 vdd.n3196 vdd.n756 72.8958
R18032 vdd.n799 vdd.n756 72.8958
R18033 vdd.n3203 vdd.n756 72.8958
R18034 vdd.n796 vdd.n756 72.8958
R18035 vdd.n3210 vdd.n756 72.8958
R18036 vdd.n793 vdd.n756 72.8958
R18037 vdd.n3218 vdd.n756 72.8958
R18038 vdd.n790 vdd.n756 72.8958
R18039 vdd.n3225 vdd.n756 72.8958
R18040 vdd.n787 vdd.n756 72.8958
R18041 vdd.n3232 vdd.n756 72.8958
R18042 vdd.n784 vdd.n756 72.8958
R18043 vdd.n3239 vdd.n756 72.8958
R18044 vdd.n3242 vdd.n756 72.8958
R18045 vdd.n2701 vdd.n950 72.8958
R18046 vdd.n2701 vdd.n949 72.8958
R18047 vdd.n2701 vdd.n948 72.8958
R18048 vdd.n2701 vdd.n947 72.8958
R18049 vdd.n2701 vdd.n946 72.8958
R18050 vdd.n2701 vdd.n945 72.8958
R18051 vdd.n2701 vdd.n944 72.8958
R18052 vdd.n2701 vdd.n943 72.8958
R18053 vdd.n2701 vdd.n942 72.8958
R18054 vdd.n2701 vdd.n941 72.8958
R18055 vdd.n2701 vdd.n940 72.8958
R18056 vdd.n2701 vdd.n939 72.8958
R18057 vdd.n2701 vdd.n938 72.8958
R18058 vdd.n2701 vdd.n937 72.8958
R18059 vdd.n2701 vdd.n936 72.8958
R18060 vdd.n2701 vdd.n935 72.8958
R18061 vdd.n2701 vdd.n934 72.8958
R18062 vdd.n2423 vdd.n1129 72.8958
R18063 vdd.n2423 vdd.n1130 72.8958
R18064 vdd.n2423 vdd.n1131 72.8958
R18065 vdd.n2423 vdd.n1132 72.8958
R18066 vdd.n2423 vdd.n1133 72.8958
R18067 vdd.n2423 vdd.n1134 72.8958
R18068 vdd.n2423 vdd.n1135 72.8958
R18069 vdd.n2423 vdd.n1136 72.8958
R18070 vdd.n2423 vdd.n1137 72.8958
R18071 vdd.n2423 vdd.n1138 72.8958
R18072 vdd.n2423 vdd.n1139 72.8958
R18073 vdd.n2423 vdd.n1140 72.8958
R18074 vdd.n2423 vdd.n1141 72.8958
R18075 vdd.n2423 vdd.n1142 72.8958
R18076 vdd.n2423 vdd.n1143 72.8958
R18077 vdd.n2423 vdd.n1144 72.8958
R18078 vdd.n2423 vdd.n1145 72.8958
R18079 vdd.n1829 vdd.n1828 66.2847
R18080 vdd.n1829 vdd.n1607 66.2847
R18081 vdd.n1829 vdd.n1608 66.2847
R18082 vdd.n1829 vdd.n1609 66.2847
R18083 vdd.n1829 vdd.n1610 66.2847
R18084 vdd.n1829 vdd.n1611 66.2847
R18085 vdd.n1829 vdd.n1612 66.2847
R18086 vdd.n1829 vdd.n1613 66.2847
R18087 vdd.n1829 vdd.n1614 66.2847
R18088 vdd.n1829 vdd.n1615 66.2847
R18089 vdd.n1829 vdd.n1616 66.2847
R18090 vdd.n1829 vdd.n1617 66.2847
R18091 vdd.n1829 vdd.n1618 66.2847
R18092 vdd.n1829 vdd.n1619 66.2847
R18093 vdd.n1829 vdd.n1620 66.2847
R18094 vdd.n1829 vdd.n1621 66.2847
R18095 vdd.n1829 vdd.n1622 66.2847
R18096 vdd.n1829 vdd.n1623 66.2847
R18097 vdd.n1829 vdd.n1624 66.2847
R18098 vdd.n1829 vdd.n1625 66.2847
R18099 vdd.n1829 vdd.n1626 66.2847
R18100 vdd.n1829 vdd.n1627 66.2847
R18101 vdd.n1829 vdd.n1628 66.2847
R18102 vdd.n1829 vdd.n1629 66.2847
R18103 vdd.n1829 vdd.n1630 66.2847
R18104 vdd.n1829 vdd.n1631 66.2847
R18105 vdd.n1829 vdd.n1632 66.2847
R18106 vdd.n1829 vdd.n1633 66.2847
R18107 vdd.n1829 vdd.n1634 66.2847
R18108 vdd.n1829 vdd.n1635 66.2847
R18109 vdd.n1829 vdd.n1636 66.2847
R18110 vdd.n1497 vdd.n1112 66.2847
R18111 vdd.n1494 vdd.n1112 66.2847
R18112 vdd.n1490 vdd.n1112 66.2847
R18113 vdd.n2289 vdd.n1112 66.2847
R18114 vdd.n1246 vdd.n1112 66.2847
R18115 vdd.n2296 vdd.n1112 66.2847
R18116 vdd.n1239 vdd.n1112 66.2847
R18117 vdd.n2303 vdd.n1112 66.2847
R18118 vdd.n1232 vdd.n1112 66.2847
R18119 vdd.n2310 vdd.n1112 66.2847
R18120 vdd.n1226 vdd.n1112 66.2847
R18121 vdd.n1221 vdd.n1112 66.2847
R18122 vdd.n2321 vdd.n1112 66.2847
R18123 vdd.n1213 vdd.n1112 66.2847
R18124 vdd.n2328 vdd.n1112 66.2847
R18125 vdd.n1206 vdd.n1112 66.2847
R18126 vdd.n2335 vdd.n1112 66.2847
R18127 vdd.n1199 vdd.n1112 66.2847
R18128 vdd.n2342 vdd.n1112 66.2847
R18129 vdd.n1192 vdd.n1112 66.2847
R18130 vdd.n2349 vdd.n1112 66.2847
R18131 vdd.n1186 vdd.n1112 66.2847
R18132 vdd.n1181 vdd.n1112 66.2847
R18133 vdd.n2360 vdd.n1112 66.2847
R18134 vdd.n1173 vdd.n1112 66.2847
R18135 vdd.n2367 vdd.n1112 66.2847
R18136 vdd.n1166 vdd.n1112 66.2847
R18137 vdd.n2374 vdd.n1112 66.2847
R18138 vdd.n1159 vdd.n1112 66.2847
R18139 vdd.n2381 vdd.n1112 66.2847
R18140 vdd.n2386 vdd.n1112 66.2847
R18141 vdd.n1155 vdd.n1112 66.2847
R18142 vdd.n3409 vdd.n658 66.2847
R18143 vdd.n663 vdd.n658 66.2847
R18144 vdd.n666 vdd.n658 66.2847
R18145 vdd.n3398 vdd.n658 66.2847
R18146 vdd.n3392 vdd.n658 66.2847
R18147 vdd.n3390 vdd.n658 66.2847
R18148 vdd.n3384 vdd.n658 66.2847
R18149 vdd.n3382 vdd.n658 66.2847
R18150 vdd.n3376 vdd.n658 66.2847
R18151 vdd.n3374 vdd.n658 66.2847
R18152 vdd.n3368 vdd.n658 66.2847
R18153 vdd.n3366 vdd.n658 66.2847
R18154 vdd.n3360 vdd.n658 66.2847
R18155 vdd.n3358 vdd.n658 66.2847
R18156 vdd.n3352 vdd.n658 66.2847
R18157 vdd.n3350 vdd.n658 66.2847
R18158 vdd.n3344 vdd.n658 66.2847
R18159 vdd.n3342 vdd.n658 66.2847
R18160 vdd.n3336 vdd.n658 66.2847
R18161 vdd.n3334 vdd.n658 66.2847
R18162 vdd.n727 vdd.n658 66.2847
R18163 vdd.n3325 vdd.n658 66.2847
R18164 vdd.n729 vdd.n658 66.2847
R18165 vdd.n3318 vdd.n658 66.2847
R18166 vdd.n3312 vdd.n658 66.2847
R18167 vdd.n3310 vdd.n658 66.2847
R18168 vdd.n3304 vdd.n658 66.2847
R18169 vdd.n3302 vdd.n658 66.2847
R18170 vdd.n3296 vdd.n658 66.2847
R18171 vdd.n750 vdd.n658 66.2847
R18172 vdd.n752 vdd.n658 66.2847
R18173 vdd.n3525 vdd.n3524 66.2847
R18174 vdd.n3525 vdd.n403 66.2847
R18175 vdd.n3525 vdd.n402 66.2847
R18176 vdd.n3525 vdd.n401 66.2847
R18177 vdd.n3525 vdd.n400 66.2847
R18178 vdd.n3525 vdd.n399 66.2847
R18179 vdd.n3525 vdd.n398 66.2847
R18180 vdd.n3525 vdd.n397 66.2847
R18181 vdd.n3525 vdd.n396 66.2847
R18182 vdd.n3525 vdd.n395 66.2847
R18183 vdd.n3525 vdd.n394 66.2847
R18184 vdd.n3525 vdd.n393 66.2847
R18185 vdd.n3525 vdd.n392 66.2847
R18186 vdd.n3525 vdd.n391 66.2847
R18187 vdd.n3525 vdd.n390 66.2847
R18188 vdd.n3525 vdd.n389 66.2847
R18189 vdd.n3525 vdd.n388 66.2847
R18190 vdd.n3525 vdd.n387 66.2847
R18191 vdd.n3525 vdd.n386 66.2847
R18192 vdd.n3525 vdd.n385 66.2847
R18193 vdd.n3525 vdd.n384 66.2847
R18194 vdd.n3525 vdd.n383 66.2847
R18195 vdd.n3525 vdd.n382 66.2847
R18196 vdd.n3525 vdd.n381 66.2847
R18197 vdd.n3525 vdd.n380 66.2847
R18198 vdd.n3525 vdd.n379 66.2847
R18199 vdd.n3525 vdd.n378 66.2847
R18200 vdd.n3525 vdd.n377 66.2847
R18201 vdd.n3525 vdd.n376 66.2847
R18202 vdd.n3525 vdd.n375 66.2847
R18203 vdd.n3525 vdd.n374 66.2847
R18204 vdd.n3525 vdd.n373 66.2847
R18205 vdd.n448 vdd.n373 52.4337
R18206 vdd.n454 vdd.n374 52.4337
R18207 vdd.n458 vdd.n375 52.4337
R18208 vdd.n464 vdd.n376 52.4337
R18209 vdd.n468 vdd.n377 52.4337
R18210 vdd.n474 vdd.n378 52.4337
R18211 vdd.n478 vdd.n379 52.4337
R18212 vdd.n484 vdd.n380 52.4337
R18213 vdd.n488 vdd.n381 52.4337
R18214 vdd.n494 vdd.n382 52.4337
R18215 vdd.n498 vdd.n383 52.4337
R18216 vdd.n504 vdd.n384 52.4337
R18217 vdd.n508 vdd.n385 52.4337
R18218 vdd.n514 vdd.n386 52.4337
R18219 vdd.n518 vdd.n387 52.4337
R18220 vdd.n524 vdd.n388 52.4337
R18221 vdd.n528 vdd.n389 52.4337
R18222 vdd.n534 vdd.n390 52.4337
R18223 vdd.n538 vdd.n391 52.4337
R18224 vdd.n544 vdd.n392 52.4337
R18225 vdd.n548 vdd.n393 52.4337
R18226 vdd.n554 vdd.n394 52.4337
R18227 vdd.n558 vdd.n395 52.4337
R18228 vdd.n564 vdd.n396 52.4337
R18229 vdd.n568 vdd.n397 52.4337
R18230 vdd.n574 vdd.n398 52.4337
R18231 vdd.n578 vdd.n399 52.4337
R18232 vdd.n584 vdd.n400 52.4337
R18233 vdd.n588 vdd.n401 52.4337
R18234 vdd.n594 vdd.n402 52.4337
R18235 vdd.n597 vdd.n403 52.4337
R18236 vdd.n3524 vdd.n3523 52.4337
R18237 vdd.n3409 vdd.n660 52.4337
R18238 vdd.n3407 vdd.n663 52.4337
R18239 vdd.n3403 vdd.n666 52.4337
R18240 vdd.n3399 vdd.n3398 52.4337
R18241 vdd.n3392 vdd.n669 52.4337
R18242 vdd.n3391 vdd.n3390 52.4337
R18243 vdd.n3384 vdd.n675 52.4337
R18244 vdd.n3383 vdd.n3382 52.4337
R18245 vdd.n3376 vdd.n681 52.4337
R18246 vdd.n3375 vdd.n3374 52.4337
R18247 vdd.n3368 vdd.n689 52.4337
R18248 vdd.n3367 vdd.n3366 52.4337
R18249 vdd.n3360 vdd.n695 52.4337
R18250 vdd.n3359 vdd.n3358 52.4337
R18251 vdd.n3352 vdd.n701 52.4337
R18252 vdd.n3351 vdd.n3350 52.4337
R18253 vdd.n3344 vdd.n707 52.4337
R18254 vdd.n3343 vdd.n3342 52.4337
R18255 vdd.n3336 vdd.n713 52.4337
R18256 vdd.n3335 vdd.n3334 52.4337
R18257 vdd.n727 vdd.n719 52.4337
R18258 vdd.n3326 vdd.n3325 52.4337
R18259 vdd.n3323 vdd.n729 52.4337
R18260 vdd.n3319 vdd.n3318 52.4337
R18261 vdd.n3312 vdd.n733 52.4337
R18262 vdd.n3311 vdd.n3310 52.4337
R18263 vdd.n3304 vdd.n739 52.4337
R18264 vdd.n3303 vdd.n3302 52.4337
R18265 vdd.n3296 vdd.n745 52.4337
R18266 vdd.n3295 vdd.n750 52.4337
R18267 vdd.n3291 vdd.n752 52.4337
R18268 vdd.n2388 vdd.n1155 52.4337
R18269 vdd.n2386 vdd.n2385 52.4337
R18270 vdd.n2381 vdd.n2380 52.4337
R18271 vdd.n2376 vdd.n1159 52.4337
R18272 vdd.n2374 vdd.n2373 52.4337
R18273 vdd.n2369 vdd.n1166 52.4337
R18274 vdd.n2367 vdd.n2366 52.4337
R18275 vdd.n2362 vdd.n1173 52.4337
R18276 vdd.n2360 vdd.n2359 52.4337
R18277 vdd.n1182 vdd.n1181 52.4337
R18278 vdd.n2351 vdd.n1186 52.4337
R18279 vdd.n2349 vdd.n2348 52.4337
R18280 vdd.n2344 vdd.n1192 52.4337
R18281 vdd.n2342 vdd.n2341 52.4337
R18282 vdd.n2337 vdd.n1199 52.4337
R18283 vdd.n2335 vdd.n2334 52.4337
R18284 vdd.n2330 vdd.n1206 52.4337
R18285 vdd.n2328 vdd.n2327 52.4337
R18286 vdd.n2323 vdd.n1213 52.4337
R18287 vdd.n2321 vdd.n2320 52.4337
R18288 vdd.n1222 vdd.n1221 52.4337
R18289 vdd.n2312 vdd.n1226 52.4337
R18290 vdd.n2310 vdd.n2309 52.4337
R18291 vdd.n2305 vdd.n1232 52.4337
R18292 vdd.n2303 vdd.n2302 52.4337
R18293 vdd.n2298 vdd.n1239 52.4337
R18294 vdd.n2296 vdd.n2295 52.4337
R18295 vdd.n2291 vdd.n1246 52.4337
R18296 vdd.n2289 vdd.n2288 52.4337
R18297 vdd.n1491 vdd.n1490 52.4337
R18298 vdd.n1495 vdd.n1494 52.4337
R18299 vdd.n2277 vdd.n1497 52.4337
R18300 vdd.n1828 vdd.n1827 52.4337
R18301 vdd.n1642 vdd.n1607 52.4337
R18302 vdd.n1644 vdd.n1608 52.4337
R18303 vdd.n1648 vdd.n1609 52.4337
R18304 vdd.n1650 vdd.n1610 52.4337
R18305 vdd.n1654 vdd.n1611 52.4337
R18306 vdd.n1656 vdd.n1612 52.4337
R18307 vdd.n1660 vdd.n1613 52.4337
R18308 vdd.n1662 vdd.n1614 52.4337
R18309 vdd.n1794 vdd.n1615 52.4337
R18310 vdd.n1666 vdd.n1616 52.4337
R18311 vdd.n1670 vdd.n1617 52.4337
R18312 vdd.n1672 vdd.n1618 52.4337
R18313 vdd.n1676 vdd.n1619 52.4337
R18314 vdd.n1678 vdd.n1620 52.4337
R18315 vdd.n1682 vdd.n1621 52.4337
R18316 vdd.n1684 vdd.n1622 52.4337
R18317 vdd.n1688 vdd.n1623 52.4337
R18318 vdd.n1690 vdd.n1624 52.4337
R18319 vdd.n1694 vdd.n1625 52.4337
R18320 vdd.n1758 vdd.n1626 52.4337
R18321 vdd.n1699 vdd.n1627 52.4337
R18322 vdd.n1701 vdd.n1628 52.4337
R18323 vdd.n1705 vdd.n1629 52.4337
R18324 vdd.n1707 vdd.n1630 52.4337
R18325 vdd.n1711 vdd.n1631 52.4337
R18326 vdd.n1713 vdd.n1632 52.4337
R18327 vdd.n1717 vdd.n1633 52.4337
R18328 vdd.n1719 vdd.n1634 52.4337
R18329 vdd.n1723 vdd.n1635 52.4337
R18330 vdd.n1725 vdd.n1636 52.4337
R18331 vdd.n1828 vdd.n1638 52.4337
R18332 vdd.n1643 vdd.n1607 52.4337
R18333 vdd.n1647 vdd.n1608 52.4337
R18334 vdd.n1649 vdd.n1609 52.4337
R18335 vdd.n1653 vdd.n1610 52.4337
R18336 vdd.n1655 vdd.n1611 52.4337
R18337 vdd.n1659 vdd.n1612 52.4337
R18338 vdd.n1661 vdd.n1613 52.4337
R18339 vdd.n1793 vdd.n1614 52.4337
R18340 vdd.n1665 vdd.n1615 52.4337
R18341 vdd.n1669 vdd.n1616 52.4337
R18342 vdd.n1671 vdd.n1617 52.4337
R18343 vdd.n1675 vdd.n1618 52.4337
R18344 vdd.n1677 vdd.n1619 52.4337
R18345 vdd.n1681 vdd.n1620 52.4337
R18346 vdd.n1683 vdd.n1621 52.4337
R18347 vdd.n1687 vdd.n1622 52.4337
R18348 vdd.n1689 vdd.n1623 52.4337
R18349 vdd.n1693 vdd.n1624 52.4337
R18350 vdd.n1695 vdd.n1625 52.4337
R18351 vdd.n1698 vdd.n1626 52.4337
R18352 vdd.n1700 vdd.n1627 52.4337
R18353 vdd.n1704 vdd.n1628 52.4337
R18354 vdd.n1706 vdd.n1629 52.4337
R18355 vdd.n1710 vdd.n1630 52.4337
R18356 vdd.n1712 vdd.n1631 52.4337
R18357 vdd.n1716 vdd.n1632 52.4337
R18358 vdd.n1718 vdd.n1633 52.4337
R18359 vdd.n1722 vdd.n1634 52.4337
R18360 vdd.n1724 vdd.n1635 52.4337
R18361 vdd.n1636 vdd.n1606 52.4337
R18362 vdd.n1497 vdd.n1496 52.4337
R18363 vdd.n1494 vdd.n1493 52.4337
R18364 vdd.n1490 vdd.n1247 52.4337
R18365 vdd.n2290 vdd.n2289 52.4337
R18366 vdd.n1246 vdd.n1240 52.4337
R18367 vdd.n2297 vdd.n2296 52.4337
R18368 vdd.n1239 vdd.n1233 52.4337
R18369 vdd.n2304 vdd.n2303 52.4337
R18370 vdd.n1232 vdd.n1227 52.4337
R18371 vdd.n2311 vdd.n2310 52.4337
R18372 vdd.n1226 vdd.n1225 52.4337
R18373 vdd.n1221 vdd.n1214 52.4337
R18374 vdd.n2322 vdd.n2321 52.4337
R18375 vdd.n1213 vdd.n1207 52.4337
R18376 vdd.n2329 vdd.n2328 52.4337
R18377 vdd.n1206 vdd.n1200 52.4337
R18378 vdd.n2336 vdd.n2335 52.4337
R18379 vdd.n1199 vdd.n1193 52.4337
R18380 vdd.n2343 vdd.n2342 52.4337
R18381 vdd.n1192 vdd.n1187 52.4337
R18382 vdd.n2350 vdd.n2349 52.4337
R18383 vdd.n1186 vdd.n1185 52.4337
R18384 vdd.n1181 vdd.n1174 52.4337
R18385 vdd.n2361 vdd.n2360 52.4337
R18386 vdd.n1173 vdd.n1167 52.4337
R18387 vdd.n2368 vdd.n2367 52.4337
R18388 vdd.n1166 vdd.n1160 52.4337
R18389 vdd.n2375 vdd.n2374 52.4337
R18390 vdd.n1159 vdd.n1156 52.4337
R18391 vdd.n2382 vdd.n2381 52.4337
R18392 vdd.n2387 vdd.n2386 52.4337
R18393 vdd.n1502 vdd.n1155 52.4337
R18394 vdd.n3410 vdd.n3409 52.4337
R18395 vdd.n3404 vdd.n663 52.4337
R18396 vdd.n3400 vdd.n666 52.4337
R18397 vdd.n3398 vdd.n3397 52.4337
R18398 vdd.n3393 vdd.n3392 52.4337
R18399 vdd.n3390 vdd.n3389 52.4337
R18400 vdd.n3385 vdd.n3384 52.4337
R18401 vdd.n3382 vdd.n3381 52.4337
R18402 vdd.n3377 vdd.n3376 52.4337
R18403 vdd.n3374 vdd.n3373 52.4337
R18404 vdd.n3369 vdd.n3368 52.4337
R18405 vdd.n3366 vdd.n3365 52.4337
R18406 vdd.n3361 vdd.n3360 52.4337
R18407 vdd.n3358 vdd.n3357 52.4337
R18408 vdd.n3353 vdd.n3352 52.4337
R18409 vdd.n3350 vdd.n3349 52.4337
R18410 vdd.n3345 vdd.n3344 52.4337
R18411 vdd.n3342 vdd.n3341 52.4337
R18412 vdd.n3337 vdd.n3336 52.4337
R18413 vdd.n3334 vdd.n3333 52.4337
R18414 vdd.n728 vdd.n727 52.4337
R18415 vdd.n3325 vdd.n3324 52.4337
R18416 vdd.n3320 vdd.n729 52.4337
R18417 vdd.n3318 vdd.n3317 52.4337
R18418 vdd.n3313 vdd.n3312 52.4337
R18419 vdd.n3310 vdd.n3309 52.4337
R18420 vdd.n3305 vdd.n3304 52.4337
R18421 vdd.n3302 vdd.n3301 52.4337
R18422 vdd.n3297 vdd.n3296 52.4337
R18423 vdd.n3292 vdd.n750 52.4337
R18424 vdd.n3288 vdd.n752 52.4337
R18425 vdd.n3524 vdd.n404 52.4337
R18426 vdd.n595 vdd.n403 52.4337
R18427 vdd.n589 vdd.n402 52.4337
R18428 vdd.n585 vdd.n401 52.4337
R18429 vdd.n579 vdd.n400 52.4337
R18430 vdd.n575 vdd.n399 52.4337
R18431 vdd.n569 vdd.n398 52.4337
R18432 vdd.n565 vdd.n397 52.4337
R18433 vdd.n559 vdd.n396 52.4337
R18434 vdd.n555 vdd.n395 52.4337
R18435 vdd.n549 vdd.n394 52.4337
R18436 vdd.n545 vdd.n393 52.4337
R18437 vdd.n539 vdd.n392 52.4337
R18438 vdd.n535 vdd.n391 52.4337
R18439 vdd.n529 vdd.n390 52.4337
R18440 vdd.n525 vdd.n389 52.4337
R18441 vdd.n519 vdd.n388 52.4337
R18442 vdd.n515 vdd.n387 52.4337
R18443 vdd.n509 vdd.n386 52.4337
R18444 vdd.n505 vdd.n385 52.4337
R18445 vdd.n499 vdd.n384 52.4337
R18446 vdd.n495 vdd.n383 52.4337
R18447 vdd.n489 vdd.n382 52.4337
R18448 vdd.n485 vdd.n381 52.4337
R18449 vdd.n479 vdd.n380 52.4337
R18450 vdd.n475 vdd.n379 52.4337
R18451 vdd.n469 vdd.n378 52.4337
R18452 vdd.n465 vdd.n377 52.4337
R18453 vdd.n459 vdd.n376 52.4337
R18454 vdd.n455 vdd.n375 52.4337
R18455 vdd.n449 vdd.n374 52.4337
R18456 vdd.n445 vdd.n373 52.4337
R18457 vdd.t17 vdd.t30 51.4683
R18458 vdd.n266 vdd.n264 42.0461
R18459 vdd.n168 vdd.n166 42.0461
R18460 vdd.n71 vdd.n69 42.0461
R18461 vdd.n2145 vdd.n2143 42.0461
R18462 vdd.n2047 vdd.n2045 42.0461
R18463 vdd.n1950 vdd.n1948 42.0461
R18464 vdd.n320 vdd.n319 41.6884
R18465 vdd.n222 vdd.n221 41.6884
R18466 vdd.n125 vdd.n124 41.6884
R18467 vdd.n2199 vdd.n2198 41.6884
R18468 vdd.n2101 vdd.n2100 41.6884
R18469 vdd.n2004 vdd.n2003 41.6884
R18470 vdd.n1605 vdd.n1604 41.1157
R18471 vdd.n1761 vdd.n1760 41.1157
R18472 vdd.n1797 vdd.n1796 41.1157
R18473 vdd.n407 vdd.n406 41.1157
R18474 vdd.n547 vdd.n420 41.1157
R18475 vdd.n433 vdd.n432 41.1157
R18476 vdd.n3242 vdd.n3241 39.2114
R18477 vdd.n3239 vdd.n3238 39.2114
R18478 vdd.n3234 vdd.n784 39.2114
R18479 vdd.n3232 vdd.n3231 39.2114
R18480 vdd.n3227 vdd.n787 39.2114
R18481 vdd.n3225 vdd.n3224 39.2114
R18482 vdd.n3220 vdd.n790 39.2114
R18483 vdd.n3218 vdd.n3217 39.2114
R18484 vdd.n3212 vdd.n793 39.2114
R18485 vdd.n3210 vdd.n3209 39.2114
R18486 vdd.n3205 vdd.n796 39.2114
R18487 vdd.n3203 vdd.n3202 39.2114
R18488 vdd.n3198 vdd.n799 39.2114
R18489 vdd.n3196 vdd.n3195 39.2114
R18490 vdd.n3191 vdd.n802 39.2114
R18491 vdd.n3189 vdd.n3188 39.2114
R18492 vdd.n3184 vdd.n3183 39.2114
R18493 vdd.n3007 vdd.n3006 39.2114
R18494 vdd.n2736 vdd.n2702 39.2114
R18495 vdd.n2999 vdd.n2703 39.2114
R18496 vdd.n2995 vdd.n2704 39.2114
R18497 vdd.n2991 vdd.n2705 39.2114
R18498 vdd.n2987 vdd.n2706 39.2114
R18499 vdd.n2983 vdd.n2707 39.2114
R18500 vdd.n2979 vdd.n2708 39.2114
R18501 vdd.n2975 vdd.n2709 39.2114
R18502 vdd.n2971 vdd.n2710 39.2114
R18503 vdd.n2967 vdd.n2711 39.2114
R18504 vdd.n2963 vdd.n2712 39.2114
R18505 vdd.n2959 vdd.n2713 39.2114
R18506 vdd.n2955 vdd.n2714 39.2114
R18507 vdd.n2951 vdd.n2715 39.2114
R18508 vdd.n2947 vdd.n2716 39.2114
R18509 vdd.n2942 vdd.n2717 39.2114
R18510 vdd.n2696 vdd.n968 39.2114
R18511 vdd.n2692 vdd.n967 39.2114
R18512 vdd.n2688 vdd.n966 39.2114
R18513 vdd.n2684 vdd.n965 39.2114
R18514 vdd.n2680 vdd.n964 39.2114
R18515 vdd.n2676 vdd.n963 39.2114
R18516 vdd.n2672 vdd.n962 39.2114
R18517 vdd.n2668 vdd.n961 39.2114
R18518 vdd.n2664 vdd.n960 39.2114
R18519 vdd.n2660 vdd.n959 39.2114
R18520 vdd.n2656 vdd.n958 39.2114
R18521 vdd.n2652 vdd.n957 39.2114
R18522 vdd.n2648 vdd.n956 39.2114
R18523 vdd.n2644 vdd.n955 39.2114
R18524 vdd.n2640 vdd.n954 39.2114
R18525 vdd.n2635 vdd.n953 39.2114
R18526 vdd.n2631 vdd.n952 39.2114
R18527 vdd.n2425 vdd.n2424 39.2114
R18528 vdd.n1147 vdd.n1113 39.2114
R18529 vdd.n2417 vdd.n1114 39.2114
R18530 vdd.n2413 vdd.n1115 39.2114
R18531 vdd.n2409 vdd.n1116 39.2114
R18532 vdd.n2405 vdd.n1117 39.2114
R18533 vdd.n2401 vdd.n1118 39.2114
R18534 vdd.n2397 vdd.n1119 39.2114
R18535 vdd.n2393 vdd.n1120 39.2114
R18536 vdd.n1293 vdd.n1121 39.2114
R18537 vdd.n1297 vdd.n1122 39.2114
R18538 vdd.n1301 vdd.n1123 39.2114
R18539 vdd.n1305 vdd.n1124 39.2114
R18540 vdd.n1309 vdd.n1125 39.2114
R18541 vdd.n1313 vdd.n1126 39.2114
R18542 vdd.n1317 vdd.n1127 39.2114
R18543 vdd.n1322 vdd.n1128 39.2114
R18544 vdd.n3161 vdd.n3160 39.2114
R18545 vdd.n3156 vdd.n3128 39.2114
R18546 vdd.n3154 vdd.n3153 39.2114
R18547 vdd.n3149 vdd.n3131 39.2114
R18548 vdd.n3147 vdd.n3146 39.2114
R18549 vdd.n3142 vdd.n3134 39.2114
R18550 vdd.n3140 vdd.n3139 39.2114
R18551 vdd.n3135 vdd.n755 39.2114
R18552 vdd.n3279 vdd.n3278 39.2114
R18553 vdd.n3276 vdd.n3275 39.2114
R18554 vdd.n3271 vdd.n760 39.2114
R18555 vdd.n3269 vdd.n3268 39.2114
R18556 vdd.n3264 vdd.n763 39.2114
R18557 vdd.n3262 vdd.n3261 39.2114
R18558 vdd.n3257 vdd.n766 39.2114
R18559 vdd.n3255 vdd.n3254 39.2114
R18560 vdd.n3250 vdd.n772 39.2114
R18561 vdd.n2743 vdd.n2718 39.2114
R18562 vdd.n2747 vdd.n2719 39.2114
R18563 vdd.n2751 vdd.n2720 39.2114
R18564 vdd.n2755 vdd.n2721 39.2114
R18565 vdd.n2759 vdd.n2722 39.2114
R18566 vdd.n2763 vdd.n2723 39.2114
R18567 vdd.n2767 vdd.n2724 39.2114
R18568 vdd.n2771 vdd.n2725 39.2114
R18569 vdd.n2775 vdd.n2726 39.2114
R18570 vdd.n2779 vdd.n2727 39.2114
R18571 vdd.n2783 vdd.n2728 39.2114
R18572 vdd.n2787 vdd.n2729 39.2114
R18573 vdd.n2791 vdd.n2730 39.2114
R18574 vdd.n2795 vdd.n2731 39.2114
R18575 vdd.n2799 vdd.n2732 39.2114
R18576 vdd.n2803 vdd.n2733 39.2114
R18577 vdd.n2807 vdd.n2734 39.2114
R18578 vdd.n2746 vdd.n2718 39.2114
R18579 vdd.n2750 vdd.n2719 39.2114
R18580 vdd.n2754 vdd.n2720 39.2114
R18581 vdd.n2758 vdd.n2721 39.2114
R18582 vdd.n2762 vdd.n2722 39.2114
R18583 vdd.n2766 vdd.n2723 39.2114
R18584 vdd.n2770 vdd.n2724 39.2114
R18585 vdd.n2774 vdd.n2725 39.2114
R18586 vdd.n2778 vdd.n2726 39.2114
R18587 vdd.n2782 vdd.n2727 39.2114
R18588 vdd.n2786 vdd.n2728 39.2114
R18589 vdd.n2790 vdd.n2729 39.2114
R18590 vdd.n2794 vdd.n2730 39.2114
R18591 vdd.n2798 vdd.n2731 39.2114
R18592 vdd.n2802 vdd.n2732 39.2114
R18593 vdd.n2806 vdd.n2733 39.2114
R18594 vdd.n2809 vdd.n2734 39.2114
R18595 vdd.n772 vdd.n767 39.2114
R18596 vdd.n3256 vdd.n3255 39.2114
R18597 vdd.n766 vdd.n764 39.2114
R18598 vdd.n3263 vdd.n3262 39.2114
R18599 vdd.n763 vdd.n761 39.2114
R18600 vdd.n3270 vdd.n3269 39.2114
R18601 vdd.n760 vdd.n758 39.2114
R18602 vdd.n3277 vdd.n3276 39.2114
R18603 vdd.n3280 vdd.n3279 39.2114
R18604 vdd.n3136 vdd.n3135 39.2114
R18605 vdd.n3141 vdd.n3140 39.2114
R18606 vdd.n3134 vdd.n3132 39.2114
R18607 vdd.n3148 vdd.n3147 39.2114
R18608 vdd.n3131 vdd.n3129 39.2114
R18609 vdd.n3155 vdd.n3154 39.2114
R18610 vdd.n3128 vdd.n3126 39.2114
R18611 vdd.n3162 vdd.n3161 39.2114
R18612 vdd.n2424 vdd.n1111 39.2114
R18613 vdd.n2418 vdd.n1113 39.2114
R18614 vdd.n2414 vdd.n1114 39.2114
R18615 vdd.n2410 vdd.n1115 39.2114
R18616 vdd.n2406 vdd.n1116 39.2114
R18617 vdd.n2402 vdd.n1117 39.2114
R18618 vdd.n2398 vdd.n1118 39.2114
R18619 vdd.n2394 vdd.n1119 39.2114
R18620 vdd.n1292 vdd.n1120 39.2114
R18621 vdd.n1296 vdd.n1121 39.2114
R18622 vdd.n1300 vdd.n1122 39.2114
R18623 vdd.n1304 vdd.n1123 39.2114
R18624 vdd.n1308 vdd.n1124 39.2114
R18625 vdd.n1312 vdd.n1125 39.2114
R18626 vdd.n1316 vdd.n1126 39.2114
R18627 vdd.n1321 vdd.n1127 39.2114
R18628 vdd.n1325 vdd.n1128 39.2114
R18629 vdd.n2634 vdd.n952 39.2114
R18630 vdd.n2639 vdd.n953 39.2114
R18631 vdd.n2643 vdd.n954 39.2114
R18632 vdd.n2647 vdd.n955 39.2114
R18633 vdd.n2651 vdd.n956 39.2114
R18634 vdd.n2655 vdd.n957 39.2114
R18635 vdd.n2659 vdd.n958 39.2114
R18636 vdd.n2663 vdd.n959 39.2114
R18637 vdd.n2667 vdd.n960 39.2114
R18638 vdd.n2671 vdd.n961 39.2114
R18639 vdd.n2675 vdd.n962 39.2114
R18640 vdd.n2679 vdd.n963 39.2114
R18641 vdd.n2683 vdd.n964 39.2114
R18642 vdd.n2687 vdd.n965 39.2114
R18643 vdd.n2691 vdd.n966 39.2114
R18644 vdd.n2695 vdd.n967 39.2114
R18645 vdd.n970 vdd.n968 39.2114
R18646 vdd.n3006 vdd.n933 39.2114
R18647 vdd.n3000 vdd.n2702 39.2114
R18648 vdd.n2996 vdd.n2703 39.2114
R18649 vdd.n2992 vdd.n2704 39.2114
R18650 vdd.n2988 vdd.n2705 39.2114
R18651 vdd.n2984 vdd.n2706 39.2114
R18652 vdd.n2980 vdd.n2707 39.2114
R18653 vdd.n2976 vdd.n2708 39.2114
R18654 vdd.n2972 vdd.n2709 39.2114
R18655 vdd.n2968 vdd.n2710 39.2114
R18656 vdd.n2964 vdd.n2711 39.2114
R18657 vdd.n2960 vdd.n2712 39.2114
R18658 vdd.n2956 vdd.n2713 39.2114
R18659 vdd.n2952 vdd.n2714 39.2114
R18660 vdd.n2948 vdd.n2715 39.2114
R18661 vdd.n2943 vdd.n2716 39.2114
R18662 vdd.n2939 vdd.n2717 39.2114
R18663 vdd.n3183 vdd.n803 39.2114
R18664 vdd.n3190 vdd.n3189 39.2114
R18665 vdd.n802 vdd.n800 39.2114
R18666 vdd.n3197 vdd.n3196 39.2114
R18667 vdd.n799 vdd.n797 39.2114
R18668 vdd.n3204 vdd.n3203 39.2114
R18669 vdd.n796 vdd.n794 39.2114
R18670 vdd.n3211 vdd.n3210 39.2114
R18671 vdd.n793 vdd.n791 39.2114
R18672 vdd.n3219 vdd.n3218 39.2114
R18673 vdd.n790 vdd.n788 39.2114
R18674 vdd.n3226 vdd.n3225 39.2114
R18675 vdd.n787 vdd.n785 39.2114
R18676 vdd.n3233 vdd.n3232 39.2114
R18677 vdd.n784 vdd.n782 39.2114
R18678 vdd.n3240 vdd.n3239 39.2114
R18679 vdd.n3243 vdd.n3242 39.2114
R18680 vdd.n979 vdd.n934 39.2114
R18681 vdd.n2623 vdd.n935 39.2114
R18682 vdd.n2619 vdd.n936 39.2114
R18683 vdd.n2615 vdd.n937 39.2114
R18684 vdd.n2611 vdd.n938 39.2114
R18685 vdd.n2607 vdd.n939 39.2114
R18686 vdd.n2603 vdd.n940 39.2114
R18687 vdd.n2599 vdd.n941 39.2114
R18688 vdd.n2595 vdd.n942 39.2114
R18689 vdd.n2591 vdd.n943 39.2114
R18690 vdd.n2587 vdd.n944 39.2114
R18691 vdd.n2583 vdd.n945 39.2114
R18692 vdd.n2579 vdd.n946 39.2114
R18693 vdd.n2575 vdd.n947 39.2114
R18694 vdd.n2571 vdd.n948 39.2114
R18695 vdd.n2567 vdd.n949 39.2114
R18696 vdd.n2563 vdd.n950 39.2114
R18697 vdd.n1251 vdd.n1129 39.2114
R18698 vdd.n1255 vdd.n1130 39.2114
R18699 vdd.n1259 vdd.n1131 39.2114
R18700 vdd.n1263 vdd.n1132 39.2114
R18701 vdd.n1267 vdd.n1133 39.2114
R18702 vdd.n1271 vdd.n1134 39.2114
R18703 vdd.n1275 vdd.n1135 39.2114
R18704 vdd.n1279 vdd.n1136 39.2114
R18705 vdd.n1283 vdd.n1137 39.2114
R18706 vdd.n1484 vdd.n1138 39.2114
R18707 vdd.n1481 vdd.n1139 39.2114
R18708 vdd.n1477 vdd.n1140 39.2114
R18709 vdd.n1473 vdd.n1141 39.2114
R18710 vdd.n1469 vdd.n1142 39.2114
R18711 vdd.n1465 vdd.n1143 39.2114
R18712 vdd.n1461 vdd.n1144 39.2114
R18713 vdd.n1457 vdd.n1145 39.2114
R18714 vdd.n2560 vdd.n950 39.2114
R18715 vdd.n2564 vdd.n949 39.2114
R18716 vdd.n2568 vdd.n948 39.2114
R18717 vdd.n2572 vdd.n947 39.2114
R18718 vdd.n2576 vdd.n946 39.2114
R18719 vdd.n2580 vdd.n945 39.2114
R18720 vdd.n2584 vdd.n944 39.2114
R18721 vdd.n2588 vdd.n943 39.2114
R18722 vdd.n2592 vdd.n942 39.2114
R18723 vdd.n2596 vdd.n941 39.2114
R18724 vdd.n2600 vdd.n940 39.2114
R18725 vdd.n2604 vdd.n939 39.2114
R18726 vdd.n2608 vdd.n938 39.2114
R18727 vdd.n2612 vdd.n937 39.2114
R18728 vdd.n2616 vdd.n936 39.2114
R18729 vdd.n2620 vdd.n935 39.2114
R18730 vdd.n2624 vdd.n934 39.2114
R18731 vdd.n1254 vdd.n1129 39.2114
R18732 vdd.n1258 vdd.n1130 39.2114
R18733 vdd.n1262 vdd.n1131 39.2114
R18734 vdd.n1266 vdd.n1132 39.2114
R18735 vdd.n1270 vdd.n1133 39.2114
R18736 vdd.n1274 vdd.n1134 39.2114
R18737 vdd.n1278 vdd.n1135 39.2114
R18738 vdd.n1282 vdd.n1136 39.2114
R18739 vdd.n1285 vdd.n1137 39.2114
R18740 vdd.n1482 vdd.n1138 39.2114
R18741 vdd.n1478 vdd.n1139 39.2114
R18742 vdd.n1474 vdd.n1140 39.2114
R18743 vdd.n1470 vdd.n1141 39.2114
R18744 vdd.n1466 vdd.n1142 39.2114
R18745 vdd.n1462 vdd.n1143 39.2114
R18746 vdd.n1458 vdd.n1144 39.2114
R18747 vdd.n1454 vdd.n1145 39.2114
R18748 vdd.n2281 vdd.n2280 37.2369
R18749 vdd.n2317 vdd.n1220 37.2369
R18750 vdd.n2356 vdd.n1180 37.2369
R18751 vdd.n3331 vdd.n724 37.2369
R18752 vdd.n688 vdd.n687 37.2369
R18753 vdd.n3287 vdd.n3286 37.2369
R18754 vdd.n1288 vdd.n1287 30.449
R18755 vdd.n983 vdd.n982 30.449
R18756 vdd.n1319 vdd.n1291 30.449
R18757 vdd.n2637 vdd.n973 30.449
R18758 vdd.n2742 vdd.n2741 30.449
R18759 vdd.n806 vdd.n805 30.449
R18760 vdd.n2945 vdd.n2738 30.449
R18761 vdd.n770 vdd.n769 30.449
R18762 vdd.n2427 vdd.n2426 29.8151
R18763 vdd.n2699 vdd.n971 29.8151
R18764 vdd.n2632 vdd.n974 29.8151
R18765 vdd.n1327 vdd.n1324 29.8151
R18766 vdd.n2940 vdd.n2937 29.8151
R18767 vdd.n3185 vdd.n3182 29.8151
R18768 vdd.n3009 vdd.n3008 29.8151
R18769 vdd.n3246 vdd.n3245 29.8151
R18770 vdd.n3165 vdd.n3164 29.8151
R18771 vdd.n3251 vdd.n771 29.8151
R18772 vdd.n2813 vdd.n2811 29.8151
R18773 vdd.n2744 vdd.n926 29.8151
R18774 vdd.n1252 vdd.n1103 29.8151
R18775 vdd.n2627 vdd.n2626 29.8151
R18776 vdd.n2559 vdd.n2558 29.8151
R18777 vdd.n1453 vdd.n1452 29.8151
R18778 vdd.n1835 vdd.n1601 19.3944
R18779 vdd.n1835 vdd.n1591 19.3944
R18780 vdd.n1847 vdd.n1591 19.3944
R18781 vdd.n1847 vdd.n1589 19.3944
R18782 vdd.n1851 vdd.n1589 19.3944
R18783 vdd.n1851 vdd.n1579 19.3944
R18784 vdd.n1864 vdd.n1579 19.3944
R18785 vdd.n1864 vdd.n1577 19.3944
R18786 vdd.n1868 vdd.n1577 19.3944
R18787 vdd.n1868 vdd.n1569 19.3944
R18788 vdd.n1881 vdd.n1569 19.3944
R18789 vdd.n1881 vdd.n1567 19.3944
R18790 vdd.n1885 vdd.n1567 19.3944
R18791 vdd.n1885 vdd.n1556 19.3944
R18792 vdd.n1897 vdd.n1556 19.3944
R18793 vdd.n1897 vdd.n1554 19.3944
R18794 vdd.n1901 vdd.n1554 19.3944
R18795 vdd.n1901 vdd.n1545 19.3944
R18796 vdd.n2209 vdd.n1545 19.3944
R18797 vdd.n2209 vdd.n1543 19.3944
R18798 vdd.n2213 vdd.n1543 19.3944
R18799 vdd.n2213 vdd.n1534 19.3944
R18800 vdd.n2225 vdd.n1534 19.3944
R18801 vdd.n2225 vdd.n1532 19.3944
R18802 vdd.n2229 vdd.n1532 19.3944
R18803 vdd.n2229 vdd.n1522 19.3944
R18804 vdd.n2242 vdd.n1522 19.3944
R18805 vdd.n2242 vdd.n1520 19.3944
R18806 vdd.n2246 vdd.n1520 19.3944
R18807 vdd.n2246 vdd.n1512 19.3944
R18808 vdd.n2259 vdd.n1512 19.3944
R18809 vdd.n2259 vdd.n1509 19.3944
R18810 vdd.n2265 vdd.n1509 19.3944
R18811 vdd.n2265 vdd.n1510 19.3944
R18812 vdd.n1510 vdd.n1499 19.3944
R18813 vdd.n1754 vdd.n1696 19.3944
R18814 vdd.n1754 vdd.n1753 19.3944
R18815 vdd.n1753 vdd.n1752 19.3944
R18816 vdd.n1752 vdd.n1702 19.3944
R18817 vdd.n1748 vdd.n1702 19.3944
R18818 vdd.n1748 vdd.n1747 19.3944
R18819 vdd.n1747 vdd.n1746 19.3944
R18820 vdd.n1746 vdd.n1708 19.3944
R18821 vdd.n1742 vdd.n1708 19.3944
R18822 vdd.n1742 vdd.n1741 19.3944
R18823 vdd.n1741 vdd.n1740 19.3944
R18824 vdd.n1740 vdd.n1714 19.3944
R18825 vdd.n1736 vdd.n1714 19.3944
R18826 vdd.n1736 vdd.n1735 19.3944
R18827 vdd.n1735 vdd.n1734 19.3944
R18828 vdd.n1734 vdd.n1720 19.3944
R18829 vdd.n1730 vdd.n1720 19.3944
R18830 vdd.n1730 vdd.n1729 19.3944
R18831 vdd.n1729 vdd.n1728 19.3944
R18832 vdd.n1728 vdd.n1726 19.3944
R18833 vdd.n1792 vdd.n1791 19.3944
R18834 vdd.n1791 vdd.n1667 19.3944
R18835 vdd.n1787 vdd.n1667 19.3944
R18836 vdd.n1787 vdd.n1786 19.3944
R18837 vdd.n1786 vdd.n1785 19.3944
R18838 vdd.n1785 vdd.n1673 19.3944
R18839 vdd.n1781 vdd.n1673 19.3944
R18840 vdd.n1781 vdd.n1780 19.3944
R18841 vdd.n1780 vdd.n1779 19.3944
R18842 vdd.n1779 vdd.n1679 19.3944
R18843 vdd.n1775 vdd.n1679 19.3944
R18844 vdd.n1775 vdd.n1774 19.3944
R18845 vdd.n1774 vdd.n1773 19.3944
R18846 vdd.n1773 vdd.n1685 19.3944
R18847 vdd.n1769 vdd.n1685 19.3944
R18848 vdd.n1769 vdd.n1768 19.3944
R18849 vdd.n1768 vdd.n1767 19.3944
R18850 vdd.n1767 vdd.n1691 19.3944
R18851 vdd.n1763 vdd.n1691 19.3944
R18852 vdd.n1763 vdd.n1762 19.3944
R18853 vdd.n1826 vdd.n1825 19.3944
R18854 vdd.n1825 vdd.n1640 19.3944
R18855 vdd.n1821 vdd.n1640 19.3944
R18856 vdd.n1821 vdd.n1820 19.3944
R18857 vdd.n1820 vdd.n1819 19.3944
R18858 vdd.n1819 vdd.n1645 19.3944
R18859 vdd.n1815 vdd.n1645 19.3944
R18860 vdd.n1815 vdd.n1814 19.3944
R18861 vdd.n1814 vdd.n1813 19.3944
R18862 vdd.n1813 vdd.n1651 19.3944
R18863 vdd.n1809 vdd.n1651 19.3944
R18864 vdd.n1809 vdd.n1808 19.3944
R18865 vdd.n1808 vdd.n1807 19.3944
R18866 vdd.n1807 vdd.n1657 19.3944
R18867 vdd.n1803 vdd.n1657 19.3944
R18868 vdd.n1803 vdd.n1802 19.3944
R18869 vdd.n1802 vdd.n1801 19.3944
R18870 vdd.n1801 vdd.n1663 19.3944
R18871 vdd.n2313 vdd.n1218 19.3944
R18872 vdd.n2313 vdd.n1224 19.3944
R18873 vdd.n2308 vdd.n1224 19.3944
R18874 vdd.n2308 vdd.n2307 19.3944
R18875 vdd.n2307 vdd.n2306 19.3944
R18876 vdd.n2306 vdd.n1231 19.3944
R18877 vdd.n2301 vdd.n1231 19.3944
R18878 vdd.n2301 vdd.n2300 19.3944
R18879 vdd.n2300 vdd.n2299 19.3944
R18880 vdd.n2299 vdd.n1238 19.3944
R18881 vdd.n2294 vdd.n1238 19.3944
R18882 vdd.n2294 vdd.n2293 19.3944
R18883 vdd.n2293 vdd.n2292 19.3944
R18884 vdd.n2292 vdd.n1245 19.3944
R18885 vdd.n2287 vdd.n1245 19.3944
R18886 vdd.n2287 vdd.n2286 19.3944
R18887 vdd.n1492 vdd.n1250 19.3944
R18888 vdd.n2282 vdd.n1489 19.3944
R18889 vdd.n2352 vdd.n1178 19.3944
R18890 vdd.n2352 vdd.n1184 19.3944
R18891 vdd.n2347 vdd.n1184 19.3944
R18892 vdd.n2347 vdd.n2346 19.3944
R18893 vdd.n2346 vdd.n2345 19.3944
R18894 vdd.n2345 vdd.n1191 19.3944
R18895 vdd.n2340 vdd.n1191 19.3944
R18896 vdd.n2340 vdd.n2339 19.3944
R18897 vdd.n2339 vdd.n2338 19.3944
R18898 vdd.n2338 vdd.n1198 19.3944
R18899 vdd.n2333 vdd.n1198 19.3944
R18900 vdd.n2333 vdd.n2332 19.3944
R18901 vdd.n2332 vdd.n2331 19.3944
R18902 vdd.n2331 vdd.n1205 19.3944
R18903 vdd.n2326 vdd.n1205 19.3944
R18904 vdd.n2326 vdd.n2325 19.3944
R18905 vdd.n2325 vdd.n2324 19.3944
R18906 vdd.n2324 vdd.n1212 19.3944
R18907 vdd.n2319 vdd.n1212 19.3944
R18908 vdd.n2319 vdd.n2318 19.3944
R18909 vdd.n2389 vdd.n1153 19.3944
R18910 vdd.n2389 vdd.n1154 19.3944
R18911 vdd.n2384 vdd.n2383 19.3944
R18912 vdd.n2379 vdd.n2378 19.3944
R18913 vdd.n2378 vdd.n2377 19.3944
R18914 vdd.n2377 vdd.n1158 19.3944
R18915 vdd.n2372 vdd.n1158 19.3944
R18916 vdd.n2372 vdd.n2371 19.3944
R18917 vdd.n2371 vdd.n2370 19.3944
R18918 vdd.n2370 vdd.n1165 19.3944
R18919 vdd.n2365 vdd.n1165 19.3944
R18920 vdd.n2365 vdd.n2364 19.3944
R18921 vdd.n2364 vdd.n2363 19.3944
R18922 vdd.n2363 vdd.n1172 19.3944
R18923 vdd.n2358 vdd.n1172 19.3944
R18924 vdd.n2358 vdd.n2357 19.3944
R18925 vdd.n1839 vdd.n1597 19.3944
R18926 vdd.n1839 vdd.n1595 19.3944
R18927 vdd.n1843 vdd.n1595 19.3944
R18928 vdd.n1843 vdd.n1585 19.3944
R18929 vdd.n1856 vdd.n1585 19.3944
R18930 vdd.n1856 vdd.n1583 19.3944
R18931 vdd.n1860 vdd.n1583 19.3944
R18932 vdd.n1860 vdd.n1574 19.3944
R18933 vdd.n1873 vdd.n1574 19.3944
R18934 vdd.n1873 vdd.n1572 19.3944
R18935 vdd.n1877 vdd.n1572 19.3944
R18936 vdd.n1877 vdd.n1563 19.3944
R18937 vdd.n1889 vdd.n1563 19.3944
R18938 vdd.n1889 vdd.n1561 19.3944
R18939 vdd.n1893 vdd.n1561 19.3944
R18940 vdd.n1893 vdd.n1551 19.3944
R18941 vdd.n1906 vdd.n1551 19.3944
R18942 vdd.n1906 vdd.n1549 19.3944
R18943 vdd.n2205 vdd.n1549 19.3944
R18944 vdd.n2205 vdd.n1540 19.3944
R18945 vdd.n2217 vdd.n1540 19.3944
R18946 vdd.n2217 vdd.n1538 19.3944
R18947 vdd.n2221 vdd.n1538 19.3944
R18948 vdd.n2221 vdd.n1528 19.3944
R18949 vdd.n2234 vdd.n1528 19.3944
R18950 vdd.n2234 vdd.n1526 19.3944
R18951 vdd.n2238 vdd.n1526 19.3944
R18952 vdd.n2238 vdd.n1517 19.3944
R18953 vdd.n2251 vdd.n1517 19.3944
R18954 vdd.n2251 vdd.n1515 19.3944
R18955 vdd.n2255 vdd.n1515 19.3944
R18956 vdd.n2255 vdd.n1505 19.3944
R18957 vdd.n2269 vdd.n1505 19.3944
R18958 vdd.n2269 vdd.n1503 19.3944
R18959 vdd.n2273 vdd.n1503 19.3944
R18960 vdd.n3419 vdd.n655 19.3944
R18961 vdd.n3423 vdd.n655 19.3944
R18962 vdd.n3423 vdd.n646 19.3944
R18963 vdd.n3435 vdd.n646 19.3944
R18964 vdd.n3435 vdd.n644 19.3944
R18965 vdd.n3439 vdd.n644 19.3944
R18966 vdd.n3439 vdd.n633 19.3944
R18967 vdd.n3451 vdd.n633 19.3944
R18968 vdd.n3451 vdd.n631 19.3944
R18969 vdd.n3455 vdd.n631 19.3944
R18970 vdd.n3455 vdd.n622 19.3944
R18971 vdd.n3468 vdd.n622 19.3944
R18972 vdd.n3468 vdd.n620 19.3944
R18973 vdd.n3475 vdd.n620 19.3944
R18974 vdd.n3475 vdd.n3474 19.3944
R18975 vdd.n3474 vdd.n610 19.3944
R18976 vdd.n3488 vdd.n610 19.3944
R18977 vdd.n3489 vdd.n3488 19.3944
R18978 vdd.n3490 vdd.n3489 19.3944
R18979 vdd.n3490 vdd.n608 19.3944
R18980 vdd.n3495 vdd.n608 19.3944
R18981 vdd.n3496 vdd.n3495 19.3944
R18982 vdd.n3497 vdd.n3496 19.3944
R18983 vdd.n3497 vdd.n606 19.3944
R18984 vdd.n3502 vdd.n606 19.3944
R18985 vdd.n3503 vdd.n3502 19.3944
R18986 vdd.n3504 vdd.n3503 19.3944
R18987 vdd.n3504 vdd.n604 19.3944
R18988 vdd.n3510 vdd.n604 19.3944
R18989 vdd.n3511 vdd.n3510 19.3944
R18990 vdd.n3512 vdd.n3511 19.3944
R18991 vdd.n3512 vdd.n602 19.3944
R18992 vdd.n3517 vdd.n602 19.3944
R18993 vdd.n3518 vdd.n3517 19.3944
R18994 vdd.n3519 vdd.n3518 19.3944
R18995 vdd.n550 vdd.n417 19.3944
R18996 vdd.n556 vdd.n417 19.3944
R18997 vdd.n557 vdd.n556 19.3944
R18998 vdd.n560 vdd.n557 19.3944
R18999 vdd.n560 vdd.n415 19.3944
R19000 vdd.n566 vdd.n415 19.3944
R19001 vdd.n567 vdd.n566 19.3944
R19002 vdd.n570 vdd.n567 19.3944
R19003 vdd.n570 vdd.n413 19.3944
R19004 vdd.n576 vdd.n413 19.3944
R19005 vdd.n577 vdd.n576 19.3944
R19006 vdd.n580 vdd.n577 19.3944
R19007 vdd.n580 vdd.n411 19.3944
R19008 vdd.n586 vdd.n411 19.3944
R19009 vdd.n587 vdd.n586 19.3944
R19010 vdd.n590 vdd.n587 19.3944
R19011 vdd.n590 vdd.n409 19.3944
R19012 vdd.n596 vdd.n409 19.3944
R19013 vdd.n598 vdd.n596 19.3944
R19014 vdd.n599 vdd.n598 19.3944
R19015 vdd.n497 vdd.n496 19.3944
R19016 vdd.n500 vdd.n497 19.3944
R19017 vdd.n500 vdd.n429 19.3944
R19018 vdd.n506 vdd.n429 19.3944
R19019 vdd.n507 vdd.n506 19.3944
R19020 vdd.n510 vdd.n507 19.3944
R19021 vdd.n510 vdd.n427 19.3944
R19022 vdd.n516 vdd.n427 19.3944
R19023 vdd.n517 vdd.n516 19.3944
R19024 vdd.n520 vdd.n517 19.3944
R19025 vdd.n520 vdd.n425 19.3944
R19026 vdd.n526 vdd.n425 19.3944
R19027 vdd.n527 vdd.n526 19.3944
R19028 vdd.n530 vdd.n527 19.3944
R19029 vdd.n530 vdd.n423 19.3944
R19030 vdd.n536 vdd.n423 19.3944
R19031 vdd.n537 vdd.n536 19.3944
R19032 vdd.n540 vdd.n537 19.3944
R19033 vdd.n540 vdd.n421 19.3944
R19034 vdd.n546 vdd.n421 19.3944
R19035 vdd.n447 vdd.n446 19.3944
R19036 vdd.n450 vdd.n447 19.3944
R19037 vdd.n450 vdd.n441 19.3944
R19038 vdd.n456 vdd.n441 19.3944
R19039 vdd.n457 vdd.n456 19.3944
R19040 vdd.n460 vdd.n457 19.3944
R19041 vdd.n460 vdd.n439 19.3944
R19042 vdd.n466 vdd.n439 19.3944
R19043 vdd.n467 vdd.n466 19.3944
R19044 vdd.n470 vdd.n467 19.3944
R19045 vdd.n470 vdd.n437 19.3944
R19046 vdd.n476 vdd.n437 19.3944
R19047 vdd.n477 vdd.n476 19.3944
R19048 vdd.n480 vdd.n477 19.3944
R19049 vdd.n480 vdd.n435 19.3944
R19050 vdd.n486 vdd.n435 19.3944
R19051 vdd.n487 vdd.n486 19.3944
R19052 vdd.n490 vdd.n487 19.3944
R19053 vdd.n3415 vdd.n652 19.3944
R19054 vdd.n3427 vdd.n652 19.3944
R19055 vdd.n3427 vdd.n650 19.3944
R19056 vdd.n3431 vdd.n650 19.3944
R19057 vdd.n3431 vdd.n640 19.3944
R19058 vdd.n3443 vdd.n640 19.3944
R19059 vdd.n3443 vdd.n638 19.3944
R19060 vdd.n3447 vdd.n638 19.3944
R19061 vdd.n3447 vdd.n628 19.3944
R19062 vdd.n3460 vdd.n628 19.3944
R19063 vdd.n3460 vdd.n626 19.3944
R19064 vdd.n3464 vdd.n626 19.3944
R19065 vdd.n3464 vdd.n617 19.3944
R19066 vdd.n3479 vdd.n617 19.3944
R19067 vdd.n3479 vdd.n615 19.3944
R19068 vdd.n3483 vdd.n615 19.3944
R19069 vdd.n3483 vdd.n324 19.3944
R19070 vdd.n3561 vdd.n324 19.3944
R19071 vdd.n3561 vdd.n325 19.3944
R19072 vdd.n3555 vdd.n325 19.3944
R19073 vdd.n3555 vdd.n3554 19.3944
R19074 vdd.n3554 vdd.n3553 19.3944
R19075 vdd.n3553 vdd.n337 19.3944
R19076 vdd.n3547 vdd.n337 19.3944
R19077 vdd.n3547 vdd.n3546 19.3944
R19078 vdd.n3546 vdd.n3545 19.3944
R19079 vdd.n3545 vdd.n347 19.3944
R19080 vdd.n3539 vdd.n347 19.3944
R19081 vdd.n3539 vdd.n3538 19.3944
R19082 vdd.n3538 vdd.n3537 19.3944
R19083 vdd.n3537 vdd.n358 19.3944
R19084 vdd.n3531 vdd.n358 19.3944
R19085 vdd.n3531 vdd.n3530 19.3944
R19086 vdd.n3530 vdd.n3529 19.3944
R19087 vdd.n3529 vdd.n369 19.3944
R19088 vdd.n3372 vdd.n3371 19.3944
R19089 vdd.n3371 vdd.n3370 19.3944
R19090 vdd.n3370 vdd.n694 19.3944
R19091 vdd.n3364 vdd.n694 19.3944
R19092 vdd.n3364 vdd.n3363 19.3944
R19093 vdd.n3363 vdd.n3362 19.3944
R19094 vdd.n3362 vdd.n700 19.3944
R19095 vdd.n3356 vdd.n700 19.3944
R19096 vdd.n3356 vdd.n3355 19.3944
R19097 vdd.n3355 vdd.n3354 19.3944
R19098 vdd.n3354 vdd.n706 19.3944
R19099 vdd.n3348 vdd.n706 19.3944
R19100 vdd.n3348 vdd.n3347 19.3944
R19101 vdd.n3347 vdd.n3346 19.3944
R19102 vdd.n3346 vdd.n712 19.3944
R19103 vdd.n3340 vdd.n712 19.3944
R19104 vdd.n3340 vdd.n3339 19.3944
R19105 vdd.n3339 vdd.n3338 19.3944
R19106 vdd.n3338 vdd.n718 19.3944
R19107 vdd.n3332 vdd.n718 19.3944
R19108 vdd.n3412 vdd.n3411 19.3944
R19109 vdd.n3411 vdd.n662 19.3944
R19110 vdd.n3406 vdd.n3405 19.3944
R19111 vdd.n3402 vdd.n3401 19.3944
R19112 vdd.n3401 vdd.n668 19.3944
R19113 vdd.n3396 vdd.n668 19.3944
R19114 vdd.n3396 vdd.n3395 19.3944
R19115 vdd.n3395 vdd.n3394 19.3944
R19116 vdd.n3394 vdd.n674 19.3944
R19117 vdd.n3388 vdd.n674 19.3944
R19118 vdd.n3388 vdd.n3387 19.3944
R19119 vdd.n3387 vdd.n3386 19.3944
R19120 vdd.n3386 vdd.n680 19.3944
R19121 vdd.n3380 vdd.n680 19.3944
R19122 vdd.n3380 vdd.n3379 19.3944
R19123 vdd.n3379 vdd.n3378 19.3944
R19124 vdd.n3327 vdd.n722 19.3944
R19125 vdd.n3327 vdd.n726 19.3944
R19126 vdd.n3322 vdd.n726 19.3944
R19127 vdd.n3322 vdd.n3321 19.3944
R19128 vdd.n3321 vdd.n732 19.3944
R19129 vdd.n3316 vdd.n732 19.3944
R19130 vdd.n3316 vdd.n3315 19.3944
R19131 vdd.n3315 vdd.n3314 19.3944
R19132 vdd.n3314 vdd.n738 19.3944
R19133 vdd.n3308 vdd.n738 19.3944
R19134 vdd.n3308 vdd.n3307 19.3944
R19135 vdd.n3307 vdd.n3306 19.3944
R19136 vdd.n3306 vdd.n744 19.3944
R19137 vdd.n3300 vdd.n744 19.3944
R19138 vdd.n3300 vdd.n3299 19.3944
R19139 vdd.n3299 vdd.n3298 19.3944
R19140 vdd.n3294 vdd.n3293 19.3944
R19141 vdd.n3290 vdd.n3289 19.3944
R19142 vdd.n1761 vdd.n1696 19.0066
R19143 vdd.n2317 vdd.n1218 19.0066
R19144 vdd.n550 vdd.n547 19.0066
R19145 vdd.n3331 vdd.n722 19.0066
R19146 vdd.n1829 vdd.n1599 18.5924
R19147 vdd.n2275 vdd.n1112 18.5924
R19148 vdd.n3417 vdd.n658 18.5924
R19149 vdd.n3526 vdd.n3525 18.5924
R19150 vdd.n1287 vdd.n1286 16.0975
R19151 vdd.n982 vdd.n981 16.0975
R19152 vdd.n1604 vdd.n1603 16.0975
R19153 vdd.n1760 vdd.n1759 16.0975
R19154 vdd.n1796 vdd.n1795 16.0975
R19155 vdd.n2280 vdd.n2279 16.0975
R19156 vdd.n1220 vdd.n1219 16.0975
R19157 vdd.n1180 vdd.n1179 16.0975
R19158 vdd.n1291 vdd.n1290 16.0975
R19159 vdd.n973 vdd.n972 16.0975
R19160 vdd.n2741 vdd.n2740 16.0975
R19161 vdd.n406 vdd.n405 16.0975
R19162 vdd.n420 vdd.n419 16.0975
R19163 vdd.n432 vdd.n431 16.0975
R19164 vdd.n724 vdd.n723 16.0975
R19165 vdd.n687 vdd.n686 16.0975
R19166 vdd.n805 vdd.n804 16.0975
R19167 vdd.n2738 vdd.n2737 16.0975
R19168 vdd.n3286 vdd.n3285 16.0975
R19169 vdd.n769 vdd.n768 16.0975
R19170 vdd.t30 vdd.n2701 15.4182
R19171 vdd.n3005 vdd.t17 15.4182
R19172 vdd.n28 vdd.n27 14.8356
R19173 vdd.n316 vdd.n281 13.1884
R19174 vdd.n261 vdd.n226 13.1884
R19175 vdd.n218 vdd.n183 13.1884
R19176 vdd.n163 vdd.n128 13.1884
R19177 vdd.n121 vdd.n86 13.1884
R19178 vdd.n66 vdd.n31 13.1884
R19179 vdd.n2140 vdd.n2105 13.1884
R19180 vdd.n2195 vdd.n2160 13.1884
R19181 vdd.n2042 vdd.n2007 13.1884
R19182 vdd.n2097 vdd.n2062 13.1884
R19183 vdd.n1945 vdd.n1910 13.1884
R19184 vdd.n2000 vdd.n1965 13.1884
R19185 vdd.n2423 vdd.n1105 13.1509
R19186 vdd.n3248 vdd.n756 13.1509
R19187 vdd.n1797 vdd.n1792 12.9944
R19188 vdd.n1797 vdd.n1663 12.9944
R19189 vdd.n2356 vdd.n1178 12.9944
R19190 vdd.n2357 vdd.n2356 12.9944
R19191 vdd.n496 vdd.n433 12.9944
R19192 vdd.n490 vdd.n433 12.9944
R19193 vdd.n3372 vdd.n688 12.9944
R19194 vdd.n3378 vdd.n688 12.9944
R19195 vdd.n317 vdd.n279 12.8005
R19196 vdd.n312 vdd.n283 12.8005
R19197 vdd.n262 vdd.n224 12.8005
R19198 vdd.n257 vdd.n228 12.8005
R19199 vdd.n219 vdd.n181 12.8005
R19200 vdd.n214 vdd.n185 12.8005
R19201 vdd.n164 vdd.n126 12.8005
R19202 vdd.n159 vdd.n130 12.8005
R19203 vdd.n122 vdd.n84 12.8005
R19204 vdd.n117 vdd.n88 12.8005
R19205 vdd.n67 vdd.n29 12.8005
R19206 vdd.n62 vdd.n33 12.8005
R19207 vdd.n2141 vdd.n2103 12.8005
R19208 vdd.n2136 vdd.n2107 12.8005
R19209 vdd.n2196 vdd.n2158 12.8005
R19210 vdd.n2191 vdd.n2162 12.8005
R19211 vdd.n2043 vdd.n2005 12.8005
R19212 vdd.n2038 vdd.n2009 12.8005
R19213 vdd.n2098 vdd.n2060 12.8005
R19214 vdd.n2093 vdd.n2064 12.8005
R19215 vdd.n1946 vdd.n1908 12.8005
R19216 vdd.n1941 vdd.n1912 12.8005
R19217 vdd.n2001 vdd.n1963 12.8005
R19218 vdd.n1996 vdd.n1967 12.8005
R19219 vdd.n311 vdd.n284 12.0247
R19220 vdd.n256 vdd.n229 12.0247
R19221 vdd.n213 vdd.n186 12.0247
R19222 vdd.n158 vdd.n131 12.0247
R19223 vdd.n116 vdd.n89 12.0247
R19224 vdd.n61 vdd.n34 12.0247
R19225 vdd.n2135 vdd.n2108 12.0247
R19226 vdd.n2190 vdd.n2163 12.0247
R19227 vdd.n2037 vdd.n2010 12.0247
R19228 vdd.n2092 vdd.n2065 12.0247
R19229 vdd.n1940 vdd.n1913 12.0247
R19230 vdd.n1995 vdd.n1968 12.0247
R19231 vdd.n1837 vdd.n1599 11.337
R19232 vdd.n1845 vdd.n1593 11.337
R19233 vdd.n1845 vdd.n1587 11.337
R19234 vdd.n1854 vdd.n1587 11.337
R19235 vdd.n1862 vdd.n1581 11.337
R19236 vdd.n1871 vdd.n1870 11.337
R19237 vdd.n1887 vdd.n1565 11.337
R19238 vdd.n1895 vdd.n1558 11.337
R19239 vdd.n1904 vdd.n1903 11.337
R19240 vdd.n2207 vdd.n1547 11.337
R19241 vdd.n2223 vdd.n1536 11.337
R19242 vdd.n2232 vdd.n1530 11.337
R19243 vdd.n2240 vdd.n1524 11.337
R19244 vdd.n2249 vdd.n2248 11.337
R19245 vdd.n2257 vdd.n1507 11.337
R19246 vdd.n2267 vdd.n1507 11.337
R19247 vdd.n2275 vdd.n1500 11.337
R19248 vdd.n3417 vdd.n659 11.337
R19249 vdd.n3425 vdd.n648 11.337
R19250 vdd.n3433 vdd.n648 11.337
R19251 vdd.n3441 vdd.n642 11.337
R19252 vdd.n3449 vdd.n635 11.337
R19253 vdd.n3458 vdd.n3457 11.337
R19254 vdd.n3466 vdd.n624 11.337
R19255 vdd.n3485 vdd.n613 11.337
R19256 vdd.n3559 vdd.n328 11.337
R19257 vdd.n3557 vdd.n332 11.337
R19258 vdd.n3551 vdd.n3550 11.337
R19259 vdd.n3543 vdd.n349 11.337
R19260 vdd.n3542 vdd.n3541 11.337
R19261 vdd.n3535 vdd.n3534 11.337
R19262 vdd.n3534 vdd.n3533 11.337
R19263 vdd.n3533 vdd.n363 11.337
R19264 vdd.n3527 vdd.n3526 11.337
R19265 vdd.n308 vdd.n307 11.249
R19266 vdd.n253 vdd.n252 11.249
R19267 vdd.n210 vdd.n209 11.249
R19268 vdd.n155 vdd.n154 11.249
R19269 vdd.n113 vdd.n112 11.249
R19270 vdd.n58 vdd.n57 11.249
R19271 vdd.n2132 vdd.n2131 11.249
R19272 vdd.n2187 vdd.n2186 11.249
R19273 vdd.n2034 vdd.n2033 11.249
R19274 vdd.n2089 vdd.n2088 11.249
R19275 vdd.n1937 vdd.n1936 11.249
R19276 vdd.n1992 vdd.n1991 11.249
R19277 vdd.n2257 vdd.t89 10.7702
R19278 vdd.n3433 vdd.t121 10.7702
R19279 vdd.n293 vdd.n292 10.7238
R19280 vdd.n238 vdd.n237 10.7238
R19281 vdd.n195 vdd.n194 10.7238
R19282 vdd.n140 vdd.n139 10.7238
R19283 vdd.n98 vdd.n97 10.7238
R19284 vdd.n43 vdd.n42 10.7238
R19285 vdd.n2117 vdd.n2116 10.7238
R19286 vdd.n2172 vdd.n2171 10.7238
R19287 vdd.n2019 vdd.n2018 10.7238
R19288 vdd.n2074 vdd.n2073 10.7238
R19289 vdd.n1922 vdd.n1921 10.7238
R19290 vdd.n1977 vdd.n1976 10.7238
R19291 vdd.n2428 vdd.n2427 10.6151
R19292 vdd.n2428 vdd.n1098 10.6151
R19293 vdd.n2438 vdd.n1098 10.6151
R19294 vdd.n2439 vdd.n2438 10.6151
R19295 vdd.n2440 vdd.n2439 10.6151
R19296 vdd.n2440 vdd.n1085 10.6151
R19297 vdd.n2450 vdd.n1085 10.6151
R19298 vdd.n2451 vdd.n2450 10.6151
R19299 vdd.n2452 vdd.n2451 10.6151
R19300 vdd.n2452 vdd.n1073 10.6151
R19301 vdd.n2462 vdd.n1073 10.6151
R19302 vdd.n2463 vdd.n2462 10.6151
R19303 vdd.n2464 vdd.n2463 10.6151
R19304 vdd.n2464 vdd.n1062 10.6151
R19305 vdd.n2474 vdd.n1062 10.6151
R19306 vdd.n2475 vdd.n2474 10.6151
R19307 vdd.n2476 vdd.n2475 10.6151
R19308 vdd.n2476 vdd.n1049 10.6151
R19309 vdd.n2486 vdd.n1049 10.6151
R19310 vdd.n2487 vdd.n2486 10.6151
R19311 vdd.n2488 vdd.n2487 10.6151
R19312 vdd.n2488 vdd.n1037 10.6151
R19313 vdd.n2499 vdd.n1037 10.6151
R19314 vdd.n2500 vdd.n2499 10.6151
R19315 vdd.n2501 vdd.n2500 10.6151
R19316 vdd.n2501 vdd.n1025 10.6151
R19317 vdd.n2511 vdd.n1025 10.6151
R19318 vdd.n2512 vdd.n2511 10.6151
R19319 vdd.n2513 vdd.n2512 10.6151
R19320 vdd.n2513 vdd.n1013 10.6151
R19321 vdd.n2523 vdd.n1013 10.6151
R19322 vdd.n2524 vdd.n2523 10.6151
R19323 vdd.n2525 vdd.n2524 10.6151
R19324 vdd.n2525 vdd.n1003 10.6151
R19325 vdd.n2535 vdd.n1003 10.6151
R19326 vdd.n2536 vdd.n2535 10.6151
R19327 vdd.n2537 vdd.n2536 10.6151
R19328 vdd.n2537 vdd.n990 10.6151
R19329 vdd.n2549 vdd.n990 10.6151
R19330 vdd.n2550 vdd.n2549 10.6151
R19331 vdd.n2552 vdd.n2550 10.6151
R19332 vdd.n2552 vdd.n2551 10.6151
R19333 vdd.n2551 vdd.n971 10.6151
R19334 vdd.n2699 vdd.n2698 10.6151
R19335 vdd.n2698 vdd.n2697 10.6151
R19336 vdd.n2697 vdd.n2694 10.6151
R19337 vdd.n2694 vdd.n2693 10.6151
R19338 vdd.n2693 vdd.n2690 10.6151
R19339 vdd.n2690 vdd.n2689 10.6151
R19340 vdd.n2689 vdd.n2686 10.6151
R19341 vdd.n2686 vdd.n2685 10.6151
R19342 vdd.n2685 vdd.n2682 10.6151
R19343 vdd.n2682 vdd.n2681 10.6151
R19344 vdd.n2681 vdd.n2678 10.6151
R19345 vdd.n2678 vdd.n2677 10.6151
R19346 vdd.n2677 vdd.n2674 10.6151
R19347 vdd.n2674 vdd.n2673 10.6151
R19348 vdd.n2673 vdd.n2670 10.6151
R19349 vdd.n2670 vdd.n2669 10.6151
R19350 vdd.n2669 vdd.n2666 10.6151
R19351 vdd.n2666 vdd.n2665 10.6151
R19352 vdd.n2665 vdd.n2662 10.6151
R19353 vdd.n2662 vdd.n2661 10.6151
R19354 vdd.n2661 vdd.n2658 10.6151
R19355 vdd.n2658 vdd.n2657 10.6151
R19356 vdd.n2657 vdd.n2654 10.6151
R19357 vdd.n2654 vdd.n2653 10.6151
R19358 vdd.n2653 vdd.n2650 10.6151
R19359 vdd.n2650 vdd.n2649 10.6151
R19360 vdd.n2649 vdd.n2646 10.6151
R19361 vdd.n2646 vdd.n2645 10.6151
R19362 vdd.n2645 vdd.n2642 10.6151
R19363 vdd.n2642 vdd.n2641 10.6151
R19364 vdd.n2641 vdd.n2638 10.6151
R19365 vdd.n2636 vdd.n2633 10.6151
R19366 vdd.n2633 vdd.n2632 10.6151
R19367 vdd.n1328 vdd.n1327 10.6151
R19368 vdd.n1330 vdd.n1328 10.6151
R19369 vdd.n1331 vdd.n1330 10.6151
R19370 vdd.n1333 vdd.n1331 10.6151
R19371 vdd.n1334 vdd.n1333 10.6151
R19372 vdd.n1336 vdd.n1334 10.6151
R19373 vdd.n1337 vdd.n1336 10.6151
R19374 vdd.n1339 vdd.n1337 10.6151
R19375 vdd.n1340 vdd.n1339 10.6151
R19376 vdd.n1342 vdd.n1340 10.6151
R19377 vdd.n1343 vdd.n1342 10.6151
R19378 vdd.n1345 vdd.n1343 10.6151
R19379 vdd.n1346 vdd.n1345 10.6151
R19380 vdd.n1348 vdd.n1346 10.6151
R19381 vdd.n1349 vdd.n1348 10.6151
R19382 vdd.n1351 vdd.n1349 10.6151
R19383 vdd.n1352 vdd.n1351 10.6151
R19384 vdd.n1354 vdd.n1352 10.6151
R19385 vdd.n1355 vdd.n1354 10.6151
R19386 vdd.n1357 vdd.n1355 10.6151
R19387 vdd.n1358 vdd.n1357 10.6151
R19388 vdd.n1360 vdd.n1358 10.6151
R19389 vdd.n1361 vdd.n1360 10.6151
R19390 vdd.n1363 vdd.n1361 10.6151
R19391 vdd.n1364 vdd.n1363 10.6151
R19392 vdd.n1366 vdd.n1364 10.6151
R19393 vdd.n1367 vdd.n1366 10.6151
R19394 vdd.n1406 vdd.n1367 10.6151
R19395 vdd.n1406 vdd.n1405 10.6151
R19396 vdd.n1405 vdd.n1404 10.6151
R19397 vdd.n1404 vdd.n1402 10.6151
R19398 vdd.n1402 vdd.n1401 10.6151
R19399 vdd.n1401 vdd.n1399 10.6151
R19400 vdd.n1399 vdd.n1398 10.6151
R19401 vdd.n1398 vdd.n1379 10.6151
R19402 vdd.n1379 vdd.n1378 10.6151
R19403 vdd.n1378 vdd.n1376 10.6151
R19404 vdd.n1376 vdd.n1375 10.6151
R19405 vdd.n1375 vdd.n1373 10.6151
R19406 vdd.n1373 vdd.n1372 10.6151
R19407 vdd.n1372 vdd.n1369 10.6151
R19408 vdd.n1369 vdd.n1368 10.6151
R19409 vdd.n1368 vdd.n974 10.6151
R19410 vdd.n2426 vdd.n1110 10.6151
R19411 vdd.n2421 vdd.n1110 10.6151
R19412 vdd.n2421 vdd.n2420 10.6151
R19413 vdd.n2420 vdd.n2419 10.6151
R19414 vdd.n2419 vdd.n2416 10.6151
R19415 vdd.n2416 vdd.n2415 10.6151
R19416 vdd.n2415 vdd.n2412 10.6151
R19417 vdd.n2412 vdd.n2411 10.6151
R19418 vdd.n2411 vdd.n2408 10.6151
R19419 vdd.n2408 vdd.n2407 10.6151
R19420 vdd.n2407 vdd.n2404 10.6151
R19421 vdd.n2404 vdd.n2403 10.6151
R19422 vdd.n2403 vdd.n2400 10.6151
R19423 vdd.n2400 vdd.n2399 10.6151
R19424 vdd.n2399 vdd.n2396 10.6151
R19425 vdd.n2396 vdd.n2395 10.6151
R19426 vdd.n2395 vdd.n2392 10.6151
R19427 vdd.n2392 vdd.n1148 10.6151
R19428 vdd.n1294 vdd.n1148 10.6151
R19429 vdd.n1295 vdd.n1294 10.6151
R19430 vdd.n1298 vdd.n1295 10.6151
R19431 vdd.n1299 vdd.n1298 10.6151
R19432 vdd.n1302 vdd.n1299 10.6151
R19433 vdd.n1303 vdd.n1302 10.6151
R19434 vdd.n1306 vdd.n1303 10.6151
R19435 vdd.n1307 vdd.n1306 10.6151
R19436 vdd.n1310 vdd.n1307 10.6151
R19437 vdd.n1311 vdd.n1310 10.6151
R19438 vdd.n1314 vdd.n1311 10.6151
R19439 vdd.n1315 vdd.n1314 10.6151
R19440 vdd.n1318 vdd.n1315 10.6151
R19441 vdd.n1323 vdd.n1320 10.6151
R19442 vdd.n1324 vdd.n1323 10.6151
R19443 vdd.n2937 vdd.n2936 10.6151
R19444 vdd.n2936 vdd.n2935 10.6151
R19445 vdd.n2935 vdd.n2739 10.6151
R19446 vdd.n2817 vdd.n2739 10.6151
R19447 vdd.n2818 vdd.n2817 10.6151
R19448 vdd.n2820 vdd.n2818 10.6151
R19449 vdd.n2821 vdd.n2820 10.6151
R19450 vdd.n2919 vdd.n2821 10.6151
R19451 vdd.n2919 vdd.n2918 10.6151
R19452 vdd.n2918 vdd.n2917 10.6151
R19453 vdd.n2917 vdd.n2865 10.6151
R19454 vdd.n2865 vdd.n2864 10.6151
R19455 vdd.n2864 vdd.n2862 10.6151
R19456 vdd.n2862 vdd.n2861 10.6151
R19457 vdd.n2861 vdd.n2859 10.6151
R19458 vdd.n2859 vdd.n2858 10.6151
R19459 vdd.n2858 vdd.n2856 10.6151
R19460 vdd.n2856 vdd.n2855 10.6151
R19461 vdd.n2855 vdd.n2853 10.6151
R19462 vdd.n2853 vdd.n2852 10.6151
R19463 vdd.n2852 vdd.n2850 10.6151
R19464 vdd.n2850 vdd.n2849 10.6151
R19465 vdd.n2849 vdd.n2847 10.6151
R19466 vdd.n2847 vdd.n2846 10.6151
R19467 vdd.n2846 vdd.n2844 10.6151
R19468 vdd.n2844 vdd.n2843 10.6151
R19469 vdd.n2843 vdd.n2841 10.6151
R19470 vdd.n2841 vdd.n2840 10.6151
R19471 vdd.n2840 vdd.n2838 10.6151
R19472 vdd.n2838 vdd.n2837 10.6151
R19473 vdd.n2837 vdd.n2835 10.6151
R19474 vdd.n2835 vdd.n2834 10.6151
R19475 vdd.n2834 vdd.n2832 10.6151
R19476 vdd.n2832 vdd.n2831 10.6151
R19477 vdd.n2831 vdd.n2829 10.6151
R19478 vdd.n2829 vdd.n2828 10.6151
R19479 vdd.n2828 vdd.n2826 10.6151
R19480 vdd.n2826 vdd.n2825 10.6151
R19481 vdd.n2825 vdd.n2823 10.6151
R19482 vdd.n2823 vdd.n2822 10.6151
R19483 vdd.n2822 vdd.n807 10.6151
R19484 vdd.n3181 vdd.n807 10.6151
R19485 vdd.n3182 vdd.n3181 10.6151
R19486 vdd.n3008 vdd.n932 10.6151
R19487 vdd.n3003 vdd.n932 10.6151
R19488 vdd.n3003 vdd.n3002 10.6151
R19489 vdd.n3002 vdd.n3001 10.6151
R19490 vdd.n3001 vdd.n2998 10.6151
R19491 vdd.n2998 vdd.n2997 10.6151
R19492 vdd.n2997 vdd.n2994 10.6151
R19493 vdd.n2994 vdd.n2993 10.6151
R19494 vdd.n2993 vdd.n2990 10.6151
R19495 vdd.n2990 vdd.n2989 10.6151
R19496 vdd.n2989 vdd.n2986 10.6151
R19497 vdd.n2986 vdd.n2985 10.6151
R19498 vdd.n2985 vdd.n2982 10.6151
R19499 vdd.n2982 vdd.n2981 10.6151
R19500 vdd.n2981 vdd.n2978 10.6151
R19501 vdd.n2978 vdd.n2977 10.6151
R19502 vdd.n2977 vdd.n2974 10.6151
R19503 vdd.n2974 vdd.n2973 10.6151
R19504 vdd.n2973 vdd.n2970 10.6151
R19505 vdd.n2970 vdd.n2969 10.6151
R19506 vdd.n2969 vdd.n2966 10.6151
R19507 vdd.n2966 vdd.n2965 10.6151
R19508 vdd.n2965 vdd.n2962 10.6151
R19509 vdd.n2962 vdd.n2961 10.6151
R19510 vdd.n2961 vdd.n2958 10.6151
R19511 vdd.n2958 vdd.n2957 10.6151
R19512 vdd.n2957 vdd.n2954 10.6151
R19513 vdd.n2954 vdd.n2953 10.6151
R19514 vdd.n2953 vdd.n2950 10.6151
R19515 vdd.n2950 vdd.n2949 10.6151
R19516 vdd.n2949 vdd.n2946 10.6151
R19517 vdd.n2944 vdd.n2941 10.6151
R19518 vdd.n2941 vdd.n2940 10.6151
R19519 vdd.n3010 vdd.n3009 10.6151
R19520 vdd.n3010 vdd.n921 10.6151
R19521 vdd.n3020 vdd.n921 10.6151
R19522 vdd.n3021 vdd.n3020 10.6151
R19523 vdd.n3022 vdd.n3021 10.6151
R19524 vdd.n3022 vdd.n909 10.6151
R19525 vdd.n3032 vdd.n909 10.6151
R19526 vdd.n3033 vdd.n3032 10.6151
R19527 vdd.n3034 vdd.n3033 10.6151
R19528 vdd.n3034 vdd.n898 10.6151
R19529 vdd.n3044 vdd.n898 10.6151
R19530 vdd.n3045 vdd.n3044 10.6151
R19531 vdd.n3046 vdd.n3045 10.6151
R19532 vdd.n3046 vdd.n887 10.6151
R19533 vdd.n3056 vdd.n887 10.6151
R19534 vdd.n3057 vdd.n3056 10.6151
R19535 vdd.n3058 vdd.n3057 10.6151
R19536 vdd.n3058 vdd.n874 10.6151
R19537 vdd.n3069 vdd.n874 10.6151
R19538 vdd.n3070 vdd.n3069 10.6151
R19539 vdd.n3071 vdd.n3070 10.6151
R19540 vdd.n3071 vdd.n862 10.6151
R19541 vdd.n3081 vdd.n862 10.6151
R19542 vdd.n3082 vdd.n3081 10.6151
R19543 vdd.n3083 vdd.n3082 10.6151
R19544 vdd.n3083 vdd.n850 10.6151
R19545 vdd.n3093 vdd.n850 10.6151
R19546 vdd.n3094 vdd.n3093 10.6151
R19547 vdd.n3095 vdd.n3094 10.6151
R19548 vdd.n3095 vdd.n837 10.6151
R19549 vdd.n3105 vdd.n837 10.6151
R19550 vdd.n3106 vdd.n3105 10.6151
R19551 vdd.n3107 vdd.n3106 10.6151
R19552 vdd.n3107 vdd.n826 10.6151
R19553 vdd.n3117 vdd.n826 10.6151
R19554 vdd.n3118 vdd.n3117 10.6151
R19555 vdd.n3119 vdd.n3118 10.6151
R19556 vdd.n3119 vdd.n812 10.6151
R19557 vdd.n3174 vdd.n812 10.6151
R19558 vdd.n3175 vdd.n3174 10.6151
R19559 vdd.n3176 vdd.n3175 10.6151
R19560 vdd.n3176 vdd.n779 10.6151
R19561 vdd.n3246 vdd.n779 10.6151
R19562 vdd.n3245 vdd.n3244 10.6151
R19563 vdd.n3244 vdd.n780 10.6151
R19564 vdd.n781 vdd.n780 10.6151
R19565 vdd.n3237 vdd.n781 10.6151
R19566 vdd.n3237 vdd.n3236 10.6151
R19567 vdd.n3236 vdd.n3235 10.6151
R19568 vdd.n3235 vdd.n783 10.6151
R19569 vdd.n3230 vdd.n783 10.6151
R19570 vdd.n3230 vdd.n3229 10.6151
R19571 vdd.n3229 vdd.n3228 10.6151
R19572 vdd.n3228 vdd.n786 10.6151
R19573 vdd.n3223 vdd.n786 10.6151
R19574 vdd.n3223 vdd.n3222 10.6151
R19575 vdd.n3222 vdd.n3221 10.6151
R19576 vdd.n3221 vdd.n789 10.6151
R19577 vdd.n3216 vdd.n789 10.6151
R19578 vdd.n3216 vdd.n3215 10.6151
R19579 vdd.n3215 vdd.n3213 10.6151
R19580 vdd.n3213 vdd.n792 10.6151
R19581 vdd.n3208 vdd.n792 10.6151
R19582 vdd.n3208 vdd.n3207 10.6151
R19583 vdd.n3207 vdd.n3206 10.6151
R19584 vdd.n3206 vdd.n795 10.6151
R19585 vdd.n3201 vdd.n795 10.6151
R19586 vdd.n3201 vdd.n3200 10.6151
R19587 vdd.n3200 vdd.n3199 10.6151
R19588 vdd.n3199 vdd.n798 10.6151
R19589 vdd.n3194 vdd.n798 10.6151
R19590 vdd.n3194 vdd.n3193 10.6151
R19591 vdd.n3193 vdd.n3192 10.6151
R19592 vdd.n3192 vdd.n801 10.6151
R19593 vdd.n3187 vdd.n3186 10.6151
R19594 vdd.n3186 vdd.n3185 10.6151
R19595 vdd.n3164 vdd.n3125 10.6151
R19596 vdd.n3159 vdd.n3125 10.6151
R19597 vdd.n3159 vdd.n3158 10.6151
R19598 vdd.n3158 vdd.n3157 10.6151
R19599 vdd.n3157 vdd.n3127 10.6151
R19600 vdd.n3152 vdd.n3127 10.6151
R19601 vdd.n3152 vdd.n3151 10.6151
R19602 vdd.n3151 vdd.n3150 10.6151
R19603 vdd.n3150 vdd.n3130 10.6151
R19604 vdd.n3145 vdd.n3130 10.6151
R19605 vdd.n3145 vdd.n3144 10.6151
R19606 vdd.n3144 vdd.n3143 10.6151
R19607 vdd.n3143 vdd.n3133 10.6151
R19608 vdd.n3138 vdd.n3133 10.6151
R19609 vdd.n3138 vdd.n3137 10.6151
R19610 vdd.n3137 vdd.n753 10.6151
R19611 vdd.n3281 vdd.n753 10.6151
R19612 vdd.n3281 vdd.n754 10.6151
R19613 vdd.n757 vdd.n754 10.6151
R19614 vdd.n3274 vdd.n757 10.6151
R19615 vdd.n3274 vdd.n3273 10.6151
R19616 vdd.n3273 vdd.n3272 10.6151
R19617 vdd.n3272 vdd.n759 10.6151
R19618 vdd.n3267 vdd.n759 10.6151
R19619 vdd.n3267 vdd.n3266 10.6151
R19620 vdd.n3266 vdd.n3265 10.6151
R19621 vdd.n3265 vdd.n762 10.6151
R19622 vdd.n3260 vdd.n762 10.6151
R19623 vdd.n3260 vdd.n3259 10.6151
R19624 vdd.n3259 vdd.n3258 10.6151
R19625 vdd.n3258 vdd.n765 10.6151
R19626 vdd.n3253 vdd.n3252 10.6151
R19627 vdd.n3252 vdd.n3251 10.6151
R19628 vdd.n2814 vdd.n2813 10.6151
R19629 vdd.n2931 vdd.n2814 10.6151
R19630 vdd.n2931 vdd.n2930 10.6151
R19631 vdd.n2930 vdd.n2929 10.6151
R19632 vdd.n2929 vdd.n2927 10.6151
R19633 vdd.n2927 vdd.n2926 10.6151
R19634 vdd.n2926 vdd.n2924 10.6151
R19635 vdd.n2924 vdd.n2923 10.6151
R19636 vdd.n2923 vdd.n2815 10.6151
R19637 vdd.n2913 vdd.n2815 10.6151
R19638 vdd.n2913 vdd.n2912 10.6151
R19639 vdd.n2912 vdd.n2911 10.6151
R19640 vdd.n2911 vdd.n2909 10.6151
R19641 vdd.n2909 vdd.n2908 10.6151
R19642 vdd.n2908 vdd.n2906 10.6151
R19643 vdd.n2906 vdd.n2905 10.6151
R19644 vdd.n2905 vdd.n2903 10.6151
R19645 vdd.n2903 vdd.n2902 10.6151
R19646 vdd.n2902 vdd.n2900 10.6151
R19647 vdd.n2900 vdd.n2899 10.6151
R19648 vdd.n2899 vdd.n2897 10.6151
R19649 vdd.n2897 vdd.n2896 10.6151
R19650 vdd.n2896 vdd.n2894 10.6151
R19651 vdd.n2894 vdd.n2893 10.6151
R19652 vdd.n2893 vdd.n2891 10.6151
R19653 vdd.n2891 vdd.n2890 10.6151
R19654 vdd.n2890 vdd.n2888 10.6151
R19655 vdd.n2888 vdd.n2887 10.6151
R19656 vdd.n2887 vdd.n2885 10.6151
R19657 vdd.n2885 vdd.n2884 10.6151
R19658 vdd.n2884 vdd.n2882 10.6151
R19659 vdd.n2882 vdd.n2881 10.6151
R19660 vdd.n2881 vdd.n2879 10.6151
R19661 vdd.n2879 vdd.n2878 10.6151
R19662 vdd.n2878 vdd.n2876 10.6151
R19663 vdd.n2876 vdd.n2875 10.6151
R19664 vdd.n2875 vdd.n2873 10.6151
R19665 vdd.n2873 vdd.n2872 10.6151
R19666 vdd.n2872 vdd.n2870 10.6151
R19667 vdd.n2870 vdd.n2869 10.6151
R19668 vdd.n2869 vdd.n2867 10.6151
R19669 vdd.n2867 vdd.n2866 10.6151
R19670 vdd.n2866 vdd.n771 10.6151
R19671 vdd.n2745 vdd.n2744 10.6151
R19672 vdd.n2748 vdd.n2745 10.6151
R19673 vdd.n2749 vdd.n2748 10.6151
R19674 vdd.n2752 vdd.n2749 10.6151
R19675 vdd.n2753 vdd.n2752 10.6151
R19676 vdd.n2756 vdd.n2753 10.6151
R19677 vdd.n2757 vdd.n2756 10.6151
R19678 vdd.n2760 vdd.n2757 10.6151
R19679 vdd.n2761 vdd.n2760 10.6151
R19680 vdd.n2764 vdd.n2761 10.6151
R19681 vdd.n2765 vdd.n2764 10.6151
R19682 vdd.n2768 vdd.n2765 10.6151
R19683 vdd.n2769 vdd.n2768 10.6151
R19684 vdd.n2772 vdd.n2769 10.6151
R19685 vdd.n2773 vdd.n2772 10.6151
R19686 vdd.n2776 vdd.n2773 10.6151
R19687 vdd.n2777 vdd.n2776 10.6151
R19688 vdd.n2780 vdd.n2777 10.6151
R19689 vdd.n2781 vdd.n2780 10.6151
R19690 vdd.n2784 vdd.n2781 10.6151
R19691 vdd.n2785 vdd.n2784 10.6151
R19692 vdd.n2788 vdd.n2785 10.6151
R19693 vdd.n2789 vdd.n2788 10.6151
R19694 vdd.n2792 vdd.n2789 10.6151
R19695 vdd.n2793 vdd.n2792 10.6151
R19696 vdd.n2796 vdd.n2793 10.6151
R19697 vdd.n2797 vdd.n2796 10.6151
R19698 vdd.n2800 vdd.n2797 10.6151
R19699 vdd.n2801 vdd.n2800 10.6151
R19700 vdd.n2804 vdd.n2801 10.6151
R19701 vdd.n2805 vdd.n2804 10.6151
R19702 vdd.n2810 vdd.n2808 10.6151
R19703 vdd.n2811 vdd.n2810 10.6151
R19704 vdd.n3014 vdd.n926 10.6151
R19705 vdd.n3015 vdd.n3014 10.6151
R19706 vdd.n3016 vdd.n3015 10.6151
R19707 vdd.n3016 vdd.n915 10.6151
R19708 vdd.n3026 vdd.n915 10.6151
R19709 vdd.n3027 vdd.n3026 10.6151
R19710 vdd.n3028 vdd.n3027 10.6151
R19711 vdd.n3028 vdd.n904 10.6151
R19712 vdd.n3038 vdd.n904 10.6151
R19713 vdd.n3039 vdd.n3038 10.6151
R19714 vdd.n3040 vdd.n3039 10.6151
R19715 vdd.n3040 vdd.n892 10.6151
R19716 vdd.n3050 vdd.n892 10.6151
R19717 vdd.n3051 vdd.n3050 10.6151
R19718 vdd.n3052 vdd.n3051 10.6151
R19719 vdd.n3052 vdd.n881 10.6151
R19720 vdd.n3062 vdd.n881 10.6151
R19721 vdd.n3063 vdd.n3062 10.6151
R19722 vdd.n3065 vdd.n3063 10.6151
R19723 vdd.n3065 vdd.n3064 10.6151
R19724 vdd.n3076 vdd.n3075 10.6151
R19725 vdd.n3077 vdd.n3076 10.6151
R19726 vdd.n3077 vdd.n856 10.6151
R19727 vdd.n3087 vdd.n856 10.6151
R19728 vdd.n3088 vdd.n3087 10.6151
R19729 vdd.n3089 vdd.n3088 10.6151
R19730 vdd.n3089 vdd.n843 10.6151
R19731 vdd.n3099 vdd.n843 10.6151
R19732 vdd.n3100 vdd.n3099 10.6151
R19733 vdd.n3101 vdd.n3100 10.6151
R19734 vdd.n3101 vdd.n831 10.6151
R19735 vdd.n3111 vdd.n831 10.6151
R19736 vdd.n3112 vdd.n3111 10.6151
R19737 vdd.n3113 vdd.n3112 10.6151
R19738 vdd.n3113 vdd.n820 10.6151
R19739 vdd.n3123 vdd.n820 10.6151
R19740 vdd.n3124 vdd.n3123 10.6151
R19741 vdd.n3170 vdd.n3124 10.6151
R19742 vdd.n3170 vdd.n3169 10.6151
R19743 vdd.n3169 vdd.n3168 10.6151
R19744 vdd.n3168 vdd.n3167 10.6151
R19745 vdd.n3167 vdd.n3165 10.6151
R19746 vdd.n2432 vdd.n1103 10.6151
R19747 vdd.n2433 vdd.n2432 10.6151
R19748 vdd.n2434 vdd.n2433 10.6151
R19749 vdd.n2434 vdd.n1092 10.6151
R19750 vdd.n2444 vdd.n1092 10.6151
R19751 vdd.n2445 vdd.n2444 10.6151
R19752 vdd.n2446 vdd.n2445 10.6151
R19753 vdd.n2446 vdd.n1079 10.6151
R19754 vdd.n2456 vdd.n1079 10.6151
R19755 vdd.n2457 vdd.n2456 10.6151
R19756 vdd.n2458 vdd.n2457 10.6151
R19757 vdd.n2458 vdd.n1068 10.6151
R19758 vdd.n2468 vdd.n1068 10.6151
R19759 vdd.n2469 vdd.n2468 10.6151
R19760 vdd.n2470 vdd.n2469 10.6151
R19761 vdd.n2470 vdd.n1056 10.6151
R19762 vdd.n2480 vdd.n1056 10.6151
R19763 vdd.n2481 vdd.n2480 10.6151
R19764 vdd.n2482 vdd.n2481 10.6151
R19765 vdd.n2482 vdd.n1043 10.6151
R19766 vdd.n2492 vdd.n1043 10.6151
R19767 vdd.n2493 vdd.n2492 10.6151
R19768 vdd.n2495 vdd.n1031 10.6151
R19769 vdd.n2505 vdd.n1031 10.6151
R19770 vdd.n2506 vdd.n2505 10.6151
R19771 vdd.n2507 vdd.n2506 10.6151
R19772 vdd.n2507 vdd.n1019 10.6151
R19773 vdd.n2517 vdd.n1019 10.6151
R19774 vdd.n2518 vdd.n2517 10.6151
R19775 vdd.n2519 vdd.n2518 10.6151
R19776 vdd.n2519 vdd.n1008 10.6151
R19777 vdd.n2529 vdd.n1008 10.6151
R19778 vdd.n2530 vdd.n2529 10.6151
R19779 vdd.n2531 vdd.n2530 10.6151
R19780 vdd.n2531 vdd.n997 10.6151
R19781 vdd.n2541 vdd.n997 10.6151
R19782 vdd.n2542 vdd.n2541 10.6151
R19783 vdd.n2545 vdd.n2542 10.6151
R19784 vdd.n2545 vdd.n2544 10.6151
R19785 vdd.n2544 vdd.n2543 10.6151
R19786 vdd.n2543 vdd.n980 10.6151
R19787 vdd.n2627 vdd.n980 10.6151
R19788 vdd.n2626 vdd.n2625 10.6151
R19789 vdd.n2625 vdd.n2622 10.6151
R19790 vdd.n2622 vdd.n2621 10.6151
R19791 vdd.n2621 vdd.n2618 10.6151
R19792 vdd.n2618 vdd.n2617 10.6151
R19793 vdd.n2617 vdd.n2614 10.6151
R19794 vdd.n2614 vdd.n2613 10.6151
R19795 vdd.n2613 vdd.n2610 10.6151
R19796 vdd.n2610 vdd.n2609 10.6151
R19797 vdd.n2609 vdd.n2606 10.6151
R19798 vdd.n2606 vdd.n2605 10.6151
R19799 vdd.n2605 vdd.n2602 10.6151
R19800 vdd.n2602 vdd.n2601 10.6151
R19801 vdd.n2601 vdd.n2598 10.6151
R19802 vdd.n2598 vdd.n2597 10.6151
R19803 vdd.n2597 vdd.n2594 10.6151
R19804 vdd.n2594 vdd.n2593 10.6151
R19805 vdd.n2593 vdd.n2590 10.6151
R19806 vdd.n2590 vdd.n2589 10.6151
R19807 vdd.n2589 vdd.n2586 10.6151
R19808 vdd.n2586 vdd.n2585 10.6151
R19809 vdd.n2585 vdd.n2582 10.6151
R19810 vdd.n2582 vdd.n2581 10.6151
R19811 vdd.n2581 vdd.n2578 10.6151
R19812 vdd.n2578 vdd.n2577 10.6151
R19813 vdd.n2577 vdd.n2574 10.6151
R19814 vdd.n2574 vdd.n2573 10.6151
R19815 vdd.n2573 vdd.n2570 10.6151
R19816 vdd.n2570 vdd.n2569 10.6151
R19817 vdd.n2569 vdd.n2566 10.6151
R19818 vdd.n2566 vdd.n2565 10.6151
R19819 vdd.n2562 vdd.n2561 10.6151
R19820 vdd.n2561 vdd.n2559 10.6151
R19821 vdd.n1452 vdd.n1450 10.6151
R19822 vdd.n1450 vdd.n1449 10.6151
R19823 vdd.n1449 vdd.n1447 10.6151
R19824 vdd.n1447 vdd.n1446 10.6151
R19825 vdd.n1446 vdd.n1444 10.6151
R19826 vdd.n1444 vdd.n1443 10.6151
R19827 vdd.n1443 vdd.n1441 10.6151
R19828 vdd.n1441 vdd.n1440 10.6151
R19829 vdd.n1440 vdd.n1438 10.6151
R19830 vdd.n1438 vdd.n1437 10.6151
R19831 vdd.n1437 vdd.n1435 10.6151
R19832 vdd.n1435 vdd.n1434 10.6151
R19833 vdd.n1434 vdd.n1432 10.6151
R19834 vdd.n1432 vdd.n1431 10.6151
R19835 vdd.n1431 vdd.n1429 10.6151
R19836 vdd.n1429 vdd.n1428 10.6151
R19837 vdd.n1428 vdd.n1426 10.6151
R19838 vdd.n1426 vdd.n1425 10.6151
R19839 vdd.n1425 vdd.n1423 10.6151
R19840 vdd.n1423 vdd.n1422 10.6151
R19841 vdd.n1422 vdd.n1420 10.6151
R19842 vdd.n1420 vdd.n1419 10.6151
R19843 vdd.n1419 vdd.n1417 10.6151
R19844 vdd.n1417 vdd.n1416 10.6151
R19845 vdd.n1416 vdd.n1414 10.6151
R19846 vdd.n1414 vdd.n1413 10.6151
R19847 vdd.n1413 vdd.n1411 10.6151
R19848 vdd.n1411 vdd.n1410 10.6151
R19849 vdd.n1410 vdd.n1289 10.6151
R19850 vdd.n1381 vdd.n1289 10.6151
R19851 vdd.n1382 vdd.n1381 10.6151
R19852 vdd.n1384 vdd.n1382 10.6151
R19853 vdd.n1385 vdd.n1384 10.6151
R19854 vdd.n1394 vdd.n1385 10.6151
R19855 vdd.n1394 vdd.n1393 10.6151
R19856 vdd.n1393 vdd.n1392 10.6151
R19857 vdd.n1392 vdd.n1390 10.6151
R19858 vdd.n1390 vdd.n1389 10.6151
R19859 vdd.n1389 vdd.n1387 10.6151
R19860 vdd.n1387 vdd.n1386 10.6151
R19861 vdd.n1386 vdd.n984 10.6151
R19862 vdd.n2557 vdd.n984 10.6151
R19863 vdd.n2558 vdd.n2557 10.6151
R19864 vdd.n1253 vdd.n1252 10.6151
R19865 vdd.n1256 vdd.n1253 10.6151
R19866 vdd.n1257 vdd.n1256 10.6151
R19867 vdd.n1260 vdd.n1257 10.6151
R19868 vdd.n1261 vdd.n1260 10.6151
R19869 vdd.n1264 vdd.n1261 10.6151
R19870 vdd.n1265 vdd.n1264 10.6151
R19871 vdd.n1268 vdd.n1265 10.6151
R19872 vdd.n1269 vdd.n1268 10.6151
R19873 vdd.n1272 vdd.n1269 10.6151
R19874 vdd.n1273 vdd.n1272 10.6151
R19875 vdd.n1276 vdd.n1273 10.6151
R19876 vdd.n1277 vdd.n1276 10.6151
R19877 vdd.n1280 vdd.n1277 10.6151
R19878 vdd.n1281 vdd.n1280 10.6151
R19879 vdd.n1284 vdd.n1281 10.6151
R19880 vdd.n1486 vdd.n1284 10.6151
R19881 vdd.n1486 vdd.n1485 10.6151
R19882 vdd.n1485 vdd.n1483 10.6151
R19883 vdd.n1483 vdd.n1480 10.6151
R19884 vdd.n1480 vdd.n1479 10.6151
R19885 vdd.n1479 vdd.n1476 10.6151
R19886 vdd.n1476 vdd.n1475 10.6151
R19887 vdd.n1475 vdd.n1472 10.6151
R19888 vdd.n1472 vdd.n1471 10.6151
R19889 vdd.n1471 vdd.n1468 10.6151
R19890 vdd.n1468 vdd.n1467 10.6151
R19891 vdd.n1467 vdd.n1464 10.6151
R19892 vdd.n1464 vdd.n1463 10.6151
R19893 vdd.n1463 vdd.n1460 10.6151
R19894 vdd.n1460 vdd.n1459 10.6151
R19895 vdd.n1456 vdd.n1455 10.6151
R19896 vdd.n1455 vdd.n1453 10.6151
R19897 vdd.t64 vdd.n2231 10.5435
R19898 vdd.n636 vdd.t75 10.5435
R19899 vdd.n304 vdd.n286 10.4732
R19900 vdd.n249 vdd.n231 10.4732
R19901 vdd.n206 vdd.n188 10.4732
R19902 vdd.n151 vdd.n133 10.4732
R19903 vdd.n109 vdd.n91 10.4732
R19904 vdd.n54 vdd.n36 10.4732
R19905 vdd.n2128 vdd.n2110 10.4732
R19906 vdd.n2183 vdd.n2165 10.4732
R19907 vdd.n2030 vdd.n2012 10.4732
R19908 vdd.n2085 vdd.n2067 10.4732
R19909 vdd.n1933 vdd.n1915 10.4732
R19910 vdd.n1988 vdd.n1970 10.4732
R19911 vdd.n2215 vdd.t58 10.3167
R19912 vdd.n3477 vdd.t119 10.3167
R19913 vdd.t128 vdd.n1559 10.09
R19914 vdd.n2267 vdd.t205 10.09
R19915 vdd.n3425 vdd.t219 10.09
R19916 vdd.n3558 vdd.t102 10.09
R19917 vdd.n2392 vdd.n2391 9.98956
R19918 vdd.n3215 vdd.n3214 9.98956
R19919 vdd.n3282 vdd.n3281 9.98956
R19920 vdd.n2284 vdd.n1486 9.98956
R19921 vdd.n1879 vdd.t144 9.86327
R19922 vdd.n3549 vdd.t93 9.86327
R19923 vdd.n2629 vdd.t48 9.7499
R19924 vdd.t35 vdd.n928 9.7499
R19925 vdd.n303 vdd.n288 9.69747
R19926 vdd.n248 vdd.n233 9.69747
R19927 vdd.n205 vdd.n190 9.69747
R19928 vdd.n150 vdd.n135 9.69747
R19929 vdd.n108 vdd.n93 9.69747
R19930 vdd.n53 vdd.n38 9.69747
R19931 vdd.n2127 vdd.n2112 9.69747
R19932 vdd.n2182 vdd.n2167 9.69747
R19933 vdd.n2029 vdd.n2014 9.69747
R19934 vdd.n2084 vdd.n2069 9.69747
R19935 vdd.n1932 vdd.n1917 9.69747
R19936 vdd.n1987 vdd.n1972 9.69747
R19937 vdd.t123 vdd.n1853 9.63654
R19938 vdd.n3508 vdd.t70 9.63654
R19939 vdd.n319 vdd.n318 9.45567
R19940 vdd.n264 vdd.n263 9.45567
R19941 vdd.n221 vdd.n220 9.45567
R19942 vdd.n166 vdd.n165 9.45567
R19943 vdd.n124 vdd.n123 9.45567
R19944 vdd.n69 vdd.n68 9.45567
R19945 vdd.n2143 vdd.n2142 9.45567
R19946 vdd.n2198 vdd.n2197 9.45567
R19947 vdd.n2045 vdd.n2044 9.45567
R19948 vdd.n2100 vdd.n2099 9.45567
R19949 vdd.n1948 vdd.n1947 9.45567
R19950 vdd.n2003 vdd.n2002 9.45567
R19951 vdd.n2354 vdd.n1178 9.3005
R19952 vdd.n2353 vdd.n2352 9.3005
R19953 vdd.n1184 vdd.n1183 9.3005
R19954 vdd.n2347 vdd.n1188 9.3005
R19955 vdd.n2346 vdd.n1189 9.3005
R19956 vdd.n2345 vdd.n1190 9.3005
R19957 vdd.n1194 vdd.n1191 9.3005
R19958 vdd.n2340 vdd.n1195 9.3005
R19959 vdd.n2339 vdd.n1196 9.3005
R19960 vdd.n2338 vdd.n1197 9.3005
R19961 vdd.n1201 vdd.n1198 9.3005
R19962 vdd.n2333 vdd.n1202 9.3005
R19963 vdd.n2332 vdd.n1203 9.3005
R19964 vdd.n2331 vdd.n1204 9.3005
R19965 vdd.n1208 vdd.n1205 9.3005
R19966 vdd.n2326 vdd.n1209 9.3005
R19967 vdd.n2325 vdd.n1210 9.3005
R19968 vdd.n2324 vdd.n1211 9.3005
R19969 vdd.n1215 vdd.n1212 9.3005
R19970 vdd.n2319 vdd.n1216 9.3005
R19971 vdd.n2318 vdd.n1217 9.3005
R19972 vdd.n2317 vdd.n2316 9.3005
R19973 vdd.n2315 vdd.n1218 9.3005
R19974 vdd.n2314 vdd.n2313 9.3005
R19975 vdd.n1224 vdd.n1223 9.3005
R19976 vdd.n2308 vdd.n1228 9.3005
R19977 vdd.n2307 vdd.n1229 9.3005
R19978 vdd.n2306 vdd.n1230 9.3005
R19979 vdd.n1234 vdd.n1231 9.3005
R19980 vdd.n2301 vdd.n1235 9.3005
R19981 vdd.n2300 vdd.n1236 9.3005
R19982 vdd.n2299 vdd.n1237 9.3005
R19983 vdd.n1241 vdd.n1238 9.3005
R19984 vdd.n2294 vdd.n1242 9.3005
R19985 vdd.n2293 vdd.n1243 9.3005
R19986 vdd.n2292 vdd.n1244 9.3005
R19987 vdd.n1248 vdd.n1245 9.3005
R19988 vdd.n2287 vdd.n1249 9.3005
R19989 vdd.n2356 vdd.n2355 9.3005
R19990 vdd.n2378 vdd.n1149 9.3005
R19991 vdd.n2377 vdd.n1157 9.3005
R19992 vdd.n1161 vdd.n1158 9.3005
R19993 vdd.n2372 vdd.n1162 9.3005
R19994 vdd.n2371 vdd.n1163 9.3005
R19995 vdd.n2370 vdd.n1164 9.3005
R19996 vdd.n1168 vdd.n1165 9.3005
R19997 vdd.n2365 vdd.n1169 9.3005
R19998 vdd.n2364 vdd.n1170 9.3005
R19999 vdd.n2363 vdd.n1171 9.3005
R20000 vdd.n1175 vdd.n1172 9.3005
R20001 vdd.n2358 vdd.n1176 9.3005
R20002 vdd.n2357 vdd.n1177 9.3005
R20003 vdd.n2390 vdd.n2389 9.3005
R20004 vdd.n1153 vdd.n1152 9.3005
R20005 vdd.n2203 vdd.n1549 9.3005
R20006 vdd.n2205 vdd.n2204 9.3005
R20007 vdd.n1540 vdd.n1539 9.3005
R20008 vdd.n2218 vdd.n2217 9.3005
R20009 vdd.n2219 vdd.n1538 9.3005
R20010 vdd.n2221 vdd.n2220 9.3005
R20011 vdd.n1528 vdd.n1527 9.3005
R20012 vdd.n2235 vdd.n2234 9.3005
R20013 vdd.n2236 vdd.n1526 9.3005
R20014 vdd.n2238 vdd.n2237 9.3005
R20015 vdd.n1517 vdd.n1516 9.3005
R20016 vdd.n2252 vdd.n2251 9.3005
R20017 vdd.n2253 vdd.n1515 9.3005
R20018 vdd.n2255 vdd.n2254 9.3005
R20019 vdd.n1505 vdd.n1504 9.3005
R20020 vdd.n2270 vdd.n2269 9.3005
R20021 vdd.n2271 vdd.n1503 9.3005
R20022 vdd.n2273 vdd.n2272 9.3005
R20023 vdd.n295 vdd.n294 9.3005
R20024 vdd.n290 vdd.n289 9.3005
R20025 vdd.n301 vdd.n300 9.3005
R20026 vdd.n303 vdd.n302 9.3005
R20027 vdd.n286 vdd.n285 9.3005
R20028 vdd.n309 vdd.n308 9.3005
R20029 vdd.n311 vdd.n310 9.3005
R20030 vdd.n283 vdd.n280 9.3005
R20031 vdd.n318 vdd.n317 9.3005
R20032 vdd.n240 vdd.n239 9.3005
R20033 vdd.n235 vdd.n234 9.3005
R20034 vdd.n246 vdd.n245 9.3005
R20035 vdd.n248 vdd.n247 9.3005
R20036 vdd.n231 vdd.n230 9.3005
R20037 vdd.n254 vdd.n253 9.3005
R20038 vdd.n256 vdd.n255 9.3005
R20039 vdd.n228 vdd.n225 9.3005
R20040 vdd.n263 vdd.n262 9.3005
R20041 vdd.n197 vdd.n196 9.3005
R20042 vdd.n192 vdd.n191 9.3005
R20043 vdd.n203 vdd.n202 9.3005
R20044 vdd.n205 vdd.n204 9.3005
R20045 vdd.n188 vdd.n187 9.3005
R20046 vdd.n211 vdd.n210 9.3005
R20047 vdd.n213 vdd.n212 9.3005
R20048 vdd.n185 vdd.n182 9.3005
R20049 vdd.n220 vdd.n219 9.3005
R20050 vdd.n142 vdd.n141 9.3005
R20051 vdd.n137 vdd.n136 9.3005
R20052 vdd.n148 vdd.n147 9.3005
R20053 vdd.n150 vdd.n149 9.3005
R20054 vdd.n133 vdd.n132 9.3005
R20055 vdd.n156 vdd.n155 9.3005
R20056 vdd.n158 vdd.n157 9.3005
R20057 vdd.n130 vdd.n127 9.3005
R20058 vdd.n165 vdd.n164 9.3005
R20059 vdd.n100 vdd.n99 9.3005
R20060 vdd.n95 vdd.n94 9.3005
R20061 vdd.n106 vdd.n105 9.3005
R20062 vdd.n108 vdd.n107 9.3005
R20063 vdd.n91 vdd.n90 9.3005
R20064 vdd.n114 vdd.n113 9.3005
R20065 vdd.n116 vdd.n115 9.3005
R20066 vdd.n88 vdd.n85 9.3005
R20067 vdd.n123 vdd.n122 9.3005
R20068 vdd.n45 vdd.n44 9.3005
R20069 vdd.n40 vdd.n39 9.3005
R20070 vdd.n51 vdd.n50 9.3005
R20071 vdd.n53 vdd.n52 9.3005
R20072 vdd.n36 vdd.n35 9.3005
R20073 vdd.n59 vdd.n58 9.3005
R20074 vdd.n61 vdd.n60 9.3005
R20075 vdd.n33 vdd.n30 9.3005
R20076 vdd.n68 vdd.n67 9.3005
R20077 vdd.n3331 vdd.n3330 9.3005
R20078 vdd.n3332 vdd.n721 9.3005
R20079 vdd.n720 vdd.n718 9.3005
R20080 vdd.n3338 vdd.n717 9.3005
R20081 vdd.n3339 vdd.n716 9.3005
R20082 vdd.n3340 vdd.n715 9.3005
R20083 vdd.n714 vdd.n712 9.3005
R20084 vdd.n3346 vdd.n711 9.3005
R20085 vdd.n3347 vdd.n710 9.3005
R20086 vdd.n3348 vdd.n709 9.3005
R20087 vdd.n708 vdd.n706 9.3005
R20088 vdd.n3354 vdd.n705 9.3005
R20089 vdd.n3355 vdd.n704 9.3005
R20090 vdd.n3356 vdd.n703 9.3005
R20091 vdd.n702 vdd.n700 9.3005
R20092 vdd.n3362 vdd.n699 9.3005
R20093 vdd.n3363 vdd.n698 9.3005
R20094 vdd.n3364 vdd.n697 9.3005
R20095 vdd.n696 vdd.n694 9.3005
R20096 vdd.n3370 vdd.n693 9.3005
R20097 vdd.n3371 vdd.n692 9.3005
R20098 vdd.n3372 vdd.n691 9.3005
R20099 vdd.n690 vdd.n688 9.3005
R20100 vdd.n3378 vdd.n685 9.3005
R20101 vdd.n3379 vdd.n684 9.3005
R20102 vdd.n3380 vdd.n683 9.3005
R20103 vdd.n682 vdd.n680 9.3005
R20104 vdd.n3386 vdd.n679 9.3005
R20105 vdd.n3387 vdd.n678 9.3005
R20106 vdd.n3388 vdd.n677 9.3005
R20107 vdd.n676 vdd.n674 9.3005
R20108 vdd.n3394 vdd.n673 9.3005
R20109 vdd.n3395 vdd.n672 9.3005
R20110 vdd.n3396 vdd.n671 9.3005
R20111 vdd.n670 vdd.n668 9.3005
R20112 vdd.n3401 vdd.n667 9.3005
R20113 vdd.n3411 vdd.n661 9.3005
R20114 vdd.n3413 vdd.n3412 9.3005
R20115 vdd.n652 vdd.n651 9.3005
R20116 vdd.n3428 vdd.n3427 9.3005
R20117 vdd.n3429 vdd.n650 9.3005
R20118 vdd.n3431 vdd.n3430 9.3005
R20119 vdd.n640 vdd.n639 9.3005
R20120 vdd.n3444 vdd.n3443 9.3005
R20121 vdd.n3445 vdd.n638 9.3005
R20122 vdd.n3447 vdd.n3446 9.3005
R20123 vdd.n628 vdd.n627 9.3005
R20124 vdd.n3461 vdd.n3460 9.3005
R20125 vdd.n3462 vdd.n626 9.3005
R20126 vdd.n3464 vdd.n3463 9.3005
R20127 vdd.n617 vdd.n616 9.3005
R20128 vdd.n3480 vdd.n3479 9.3005
R20129 vdd.n3481 vdd.n615 9.3005
R20130 vdd.n3483 vdd.n3482 9.3005
R20131 vdd.n324 vdd.n322 9.3005
R20132 vdd.n3415 vdd.n3414 9.3005
R20133 vdd.n3562 vdd.n3561 9.3005
R20134 vdd.n325 vdd.n323 9.3005
R20135 vdd.n3555 vdd.n334 9.3005
R20136 vdd.n3554 vdd.n335 9.3005
R20137 vdd.n3553 vdd.n336 9.3005
R20138 vdd.n343 vdd.n337 9.3005
R20139 vdd.n3547 vdd.n344 9.3005
R20140 vdd.n3546 vdd.n345 9.3005
R20141 vdd.n3545 vdd.n346 9.3005
R20142 vdd.n354 vdd.n347 9.3005
R20143 vdd.n3539 vdd.n355 9.3005
R20144 vdd.n3538 vdd.n356 9.3005
R20145 vdd.n3537 vdd.n357 9.3005
R20146 vdd.n365 vdd.n358 9.3005
R20147 vdd.n3531 vdd.n366 9.3005
R20148 vdd.n3530 vdd.n367 9.3005
R20149 vdd.n3529 vdd.n368 9.3005
R20150 vdd.n443 vdd.n369 9.3005
R20151 vdd.n447 vdd.n442 9.3005
R20152 vdd.n451 vdd.n450 9.3005
R20153 vdd.n452 vdd.n441 9.3005
R20154 vdd.n456 vdd.n453 9.3005
R20155 vdd.n457 vdd.n440 9.3005
R20156 vdd.n461 vdd.n460 9.3005
R20157 vdd.n462 vdd.n439 9.3005
R20158 vdd.n466 vdd.n463 9.3005
R20159 vdd.n467 vdd.n438 9.3005
R20160 vdd.n471 vdd.n470 9.3005
R20161 vdd.n472 vdd.n437 9.3005
R20162 vdd.n476 vdd.n473 9.3005
R20163 vdd.n477 vdd.n436 9.3005
R20164 vdd.n481 vdd.n480 9.3005
R20165 vdd.n482 vdd.n435 9.3005
R20166 vdd.n486 vdd.n483 9.3005
R20167 vdd.n487 vdd.n434 9.3005
R20168 vdd.n491 vdd.n490 9.3005
R20169 vdd.n492 vdd.n433 9.3005
R20170 vdd.n496 vdd.n493 9.3005
R20171 vdd.n497 vdd.n430 9.3005
R20172 vdd.n501 vdd.n500 9.3005
R20173 vdd.n502 vdd.n429 9.3005
R20174 vdd.n506 vdd.n503 9.3005
R20175 vdd.n507 vdd.n428 9.3005
R20176 vdd.n511 vdd.n510 9.3005
R20177 vdd.n512 vdd.n427 9.3005
R20178 vdd.n516 vdd.n513 9.3005
R20179 vdd.n517 vdd.n426 9.3005
R20180 vdd.n521 vdd.n520 9.3005
R20181 vdd.n522 vdd.n425 9.3005
R20182 vdd.n526 vdd.n523 9.3005
R20183 vdd.n527 vdd.n424 9.3005
R20184 vdd.n531 vdd.n530 9.3005
R20185 vdd.n532 vdd.n423 9.3005
R20186 vdd.n536 vdd.n533 9.3005
R20187 vdd.n537 vdd.n422 9.3005
R20188 vdd.n541 vdd.n540 9.3005
R20189 vdd.n542 vdd.n421 9.3005
R20190 vdd.n546 vdd.n543 9.3005
R20191 vdd.n547 vdd.n418 9.3005
R20192 vdd.n551 vdd.n550 9.3005
R20193 vdd.n552 vdd.n417 9.3005
R20194 vdd.n556 vdd.n553 9.3005
R20195 vdd.n557 vdd.n416 9.3005
R20196 vdd.n561 vdd.n560 9.3005
R20197 vdd.n562 vdd.n415 9.3005
R20198 vdd.n566 vdd.n563 9.3005
R20199 vdd.n567 vdd.n414 9.3005
R20200 vdd.n571 vdd.n570 9.3005
R20201 vdd.n572 vdd.n413 9.3005
R20202 vdd.n576 vdd.n573 9.3005
R20203 vdd.n577 vdd.n412 9.3005
R20204 vdd.n581 vdd.n580 9.3005
R20205 vdd.n582 vdd.n411 9.3005
R20206 vdd.n586 vdd.n583 9.3005
R20207 vdd.n587 vdd.n410 9.3005
R20208 vdd.n591 vdd.n590 9.3005
R20209 vdd.n592 vdd.n409 9.3005
R20210 vdd.n596 vdd.n593 9.3005
R20211 vdd.n598 vdd.n408 9.3005
R20212 vdd.n600 vdd.n599 9.3005
R20213 vdd.n3522 vdd.n3521 9.3005
R20214 vdd.n446 vdd.n444 9.3005
R20215 vdd.n3421 vdd.n655 9.3005
R20216 vdd.n3423 vdd.n3422 9.3005
R20217 vdd.n646 vdd.n645 9.3005
R20218 vdd.n3436 vdd.n3435 9.3005
R20219 vdd.n3437 vdd.n644 9.3005
R20220 vdd.n3439 vdd.n3438 9.3005
R20221 vdd.n633 vdd.n632 9.3005
R20222 vdd.n3452 vdd.n3451 9.3005
R20223 vdd.n3453 vdd.n631 9.3005
R20224 vdd.n3455 vdd.n3454 9.3005
R20225 vdd.n622 vdd.n621 9.3005
R20226 vdd.n3469 vdd.n3468 9.3005
R20227 vdd.n3470 vdd.n620 9.3005
R20228 vdd.n3475 vdd.n3471 9.3005
R20229 vdd.n3474 vdd.n3473 9.3005
R20230 vdd.n3472 vdd.n610 9.3005
R20231 vdd.n3488 vdd.n611 9.3005
R20232 vdd.n3489 vdd.n609 9.3005
R20233 vdd.n3491 vdd.n3490 9.3005
R20234 vdd.n3492 vdd.n608 9.3005
R20235 vdd.n3495 vdd.n3493 9.3005
R20236 vdd.n3496 vdd.n607 9.3005
R20237 vdd.n3498 vdd.n3497 9.3005
R20238 vdd.n3499 vdd.n606 9.3005
R20239 vdd.n3502 vdd.n3500 9.3005
R20240 vdd.n3503 vdd.n605 9.3005
R20241 vdd.n3505 vdd.n3504 9.3005
R20242 vdd.n3506 vdd.n604 9.3005
R20243 vdd.n3510 vdd.n3507 9.3005
R20244 vdd.n3511 vdd.n603 9.3005
R20245 vdd.n3513 vdd.n3512 9.3005
R20246 vdd.n3514 vdd.n602 9.3005
R20247 vdd.n3517 vdd.n3515 9.3005
R20248 vdd.n3518 vdd.n601 9.3005
R20249 vdd.n3520 vdd.n3519 9.3005
R20250 vdd.n3420 vdd.n3419 9.3005
R20251 vdd.n3284 vdd.n656 9.3005
R20252 vdd.n3289 vdd.n3283 9.3005
R20253 vdd.n3299 vdd.n748 9.3005
R20254 vdd.n3300 vdd.n747 9.3005
R20255 vdd.n746 vdd.n744 9.3005
R20256 vdd.n3306 vdd.n743 9.3005
R20257 vdd.n3307 vdd.n742 9.3005
R20258 vdd.n3308 vdd.n741 9.3005
R20259 vdd.n740 vdd.n738 9.3005
R20260 vdd.n3314 vdd.n737 9.3005
R20261 vdd.n3315 vdd.n736 9.3005
R20262 vdd.n3316 vdd.n735 9.3005
R20263 vdd.n734 vdd.n732 9.3005
R20264 vdd.n3321 vdd.n731 9.3005
R20265 vdd.n3322 vdd.n730 9.3005
R20266 vdd.n726 vdd.n725 9.3005
R20267 vdd.n3328 vdd.n3327 9.3005
R20268 vdd.n3329 vdd.n722 9.3005
R20269 vdd.n2283 vdd.n2282 9.3005
R20270 vdd.n2278 vdd.n1488 9.3005
R20271 vdd.n1835 vdd.n1834 9.3005
R20272 vdd.n1591 vdd.n1590 9.3005
R20273 vdd.n1848 vdd.n1847 9.3005
R20274 vdd.n1849 vdd.n1589 9.3005
R20275 vdd.n1851 vdd.n1850 9.3005
R20276 vdd.n1579 vdd.n1578 9.3005
R20277 vdd.n1865 vdd.n1864 9.3005
R20278 vdd.n1866 vdd.n1577 9.3005
R20279 vdd.n1868 vdd.n1867 9.3005
R20280 vdd.n1569 vdd.n1568 9.3005
R20281 vdd.n1882 vdd.n1881 9.3005
R20282 vdd.n1883 vdd.n1567 9.3005
R20283 vdd.n1885 vdd.n1884 9.3005
R20284 vdd.n1556 vdd.n1555 9.3005
R20285 vdd.n1898 vdd.n1897 9.3005
R20286 vdd.n1899 vdd.n1554 9.3005
R20287 vdd.n1901 vdd.n1900 9.3005
R20288 vdd.n1545 vdd.n1544 9.3005
R20289 vdd.n2210 vdd.n2209 9.3005
R20290 vdd.n2211 vdd.n1543 9.3005
R20291 vdd.n2213 vdd.n2212 9.3005
R20292 vdd.n1534 vdd.n1533 9.3005
R20293 vdd.n2226 vdd.n2225 9.3005
R20294 vdd.n2227 vdd.n1532 9.3005
R20295 vdd.n2229 vdd.n2228 9.3005
R20296 vdd.n1522 vdd.n1521 9.3005
R20297 vdd.n2243 vdd.n2242 9.3005
R20298 vdd.n2244 vdd.n1520 9.3005
R20299 vdd.n2246 vdd.n2245 9.3005
R20300 vdd.n1512 vdd.n1511 9.3005
R20301 vdd.n2260 vdd.n2259 9.3005
R20302 vdd.n2261 vdd.n1509 9.3005
R20303 vdd.n2265 vdd.n2264 9.3005
R20304 vdd.n2263 vdd.n1510 9.3005
R20305 vdd.n2262 vdd.n1499 9.3005
R20306 vdd.n1833 vdd.n1601 9.3005
R20307 vdd.n1726 vdd.n1602 9.3005
R20308 vdd.n1728 vdd.n1727 9.3005
R20309 vdd.n1729 vdd.n1721 9.3005
R20310 vdd.n1731 vdd.n1730 9.3005
R20311 vdd.n1732 vdd.n1720 9.3005
R20312 vdd.n1734 vdd.n1733 9.3005
R20313 vdd.n1735 vdd.n1715 9.3005
R20314 vdd.n1737 vdd.n1736 9.3005
R20315 vdd.n1738 vdd.n1714 9.3005
R20316 vdd.n1740 vdd.n1739 9.3005
R20317 vdd.n1741 vdd.n1709 9.3005
R20318 vdd.n1743 vdd.n1742 9.3005
R20319 vdd.n1744 vdd.n1708 9.3005
R20320 vdd.n1746 vdd.n1745 9.3005
R20321 vdd.n1747 vdd.n1703 9.3005
R20322 vdd.n1749 vdd.n1748 9.3005
R20323 vdd.n1750 vdd.n1702 9.3005
R20324 vdd.n1752 vdd.n1751 9.3005
R20325 vdd.n1753 vdd.n1697 9.3005
R20326 vdd.n1755 vdd.n1754 9.3005
R20327 vdd.n1756 vdd.n1696 9.3005
R20328 vdd.n1761 vdd.n1757 9.3005
R20329 vdd.n1762 vdd.n1692 9.3005
R20330 vdd.n1764 vdd.n1763 9.3005
R20331 vdd.n1765 vdd.n1691 9.3005
R20332 vdd.n1767 vdd.n1766 9.3005
R20333 vdd.n1768 vdd.n1686 9.3005
R20334 vdd.n1770 vdd.n1769 9.3005
R20335 vdd.n1771 vdd.n1685 9.3005
R20336 vdd.n1773 vdd.n1772 9.3005
R20337 vdd.n1774 vdd.n1680 9.3005
R20338 vdd.n1776 vdd.n1775 9.3005
R20339 vdd.n1777 vdd.n1679 9.3005
R20340 vdd.n1779 vdd.n1778 9.3005
R20341 vdd.n1780 vdd.n1674 9.3005
R20342 vdd.n1782 vdd.n1781 9.3005
R20343 vdd.n1783 vdd.n1673 9.3005
R20344 vdd.n1785 vdd.n1784 9.3005
R20345 vdd.n1786 vdd.n1668 9.3005
R20346 vdd.n1788 vdd.n1787 9.3005
R20347 vdd.n1789 vdd.n1667 9.3005
R20348 vdd.n1791 vdd.n1790 9.3005
R20349 vdd.n1792 vdd.n1664 9.3005
R20350 vdd.n1798 vdd.n1797 9.3005
R20351 vdd.n1799 vdd.n1663 9.3005
R20352 vdd.n1801 vdd.n1800 9.3005
R20353 vdd.n1802 vdd.n1658 9.3005
R20354 vdd.n1804 vdd.n1803 9.3005
R20355 vdd.n1805 vdd.n1657 9.3005
R20356 vdd.n1807 vdd.n1806 9.3005
R20357 vdd.n1808 vdd.n1652 9.3005
R20358 vdd.n1810 vdd.n1809 9.3005
R20359 vdd.n1811 vdd.n1651 9.3005
R20360 vdd.n1813 vdd.n1812 9.3005
R20361 vdd.n1814 vdd.n1646 9.3005
R20362 vdd.n1816 vdd.n1815 9.3005
R20363 vdd.n1817 vdd.n1645 9.3005
R20364 vdd.n1819 vdd.n1818 9.3005
R20365 vdd.n1820 vdd.n1641 9.3005
R20366 vdd.n1822 vdd.n1821 9.3005
R20367 vdd.n1823 vdd.n1640 9.3005
R20368 vdd.n1825 vdd.n1824 9.3005
R20369 vdd.n1826 vdd.n1639 9.3005
R20370 vdd.n1832 vdd.n1831 9.3005
R20371 vdd.n1840 vdd.n1839 9.3005
R20372 vdd.n1841 vdd.n1595 9.3005
R20373 vdd.n1843 vdd.n1842 9.3005
R20374 vdd.n1585 vdd.n1584 9.3005
R20375 vdd.n1857 vdd.n1856 9.3005
R20376 vdd.n1858 vdd.n1583 9.3005
R20377 vdd.n1860 vdd.n1859 9.3005
R20378 vdd.n1574 vdd.n1573 9.3005
R20379 vdd.n1874 vdd.n1873 9.3005
R20380 vdd.n1875 vdd.n1572 9.3005
R20381 vdd.n1877 vdd.n1876 9.3005
R20382 vdd.n1563 vdd.n1562 9.3005
R20383 vdd.n1890 vdd.n1889 9.3005
R20384 vdd.n1891 vdd.n1561 9.3005
R20385 vdd.n1893 vdd.n1892 9.3005
R20386 vdd.n1551 vdd.n1550 9.3005
R20387 vdd.n1907 vdd.n1906 9.3005
R20388 vdd.n1597 vdd.n1596 9.3005
R20389 vdd.n2119 vdd.n2118 9.3005
R20390 vdd.n2114 vdd.n2113 9.3005
R20391 vdd.n2125 vdd.n2124 9.3005
R20392 vdd.n2127 vdd.n2126 9.3005
R20393 vdd.n2110 vdd.n2109 9.3005
R20394 vdd.n2133 vdd.n2132 9.3005
R20395 vdd.n2135 vdd.n2134 9.3005
R20396 vdd.n2107 vdd.n2104 9.3005
R20397 vdd.n2142 vdd.n2141 9.3005
R20398 vdd.n2174 vdd.n2173 9.3005
R20399 vdd.n2169 vdd.n2168 9.3005
R20400 vdd.n2180 vdd.n2179 9.3005
R20401 vdd.n2182 vdd.n2181 9.3005
R20402 vdd.n2165 vdd.n2164 9.3005
R20403 vdd.n2188 vdd.n2187 9.3005
R20404 vdd.n2190 vdd.n2189 9.3005
R20405 vdd.n2162 vdd.n2159 9.3005
R20406 vdd.n2197 vdd.n2196 9.3005
R20407 vdd.n2021 vdd.n2020 9.3005
R20408 vdd.n2016 vdd.n2015 9.3005
R20409 vdd.n2027 vdd.n2026 9.3005
R20410 vdd.n2029 vdd.n2028 9.3005
R20411 vdd.n2012 vdd.n2011 9.3005
R20412 vdd.n2035 vdd.n2034 9.3005
R20413 vdd.n2037 vdd.n2036 9.3005
R20414 vdd.n2009 vdd.n2006 9.3005
R20415 vdd.n2044 vdd.n2043 9.3005
R20416 vdd.n2076 vdd.n2075 9.3005
R20417 vdd.n2071 vdd.n2070 9.3005
R20418 vdd.n2082 vdd.n2081 9.3005
R20419 vdd.n2084 vdd.n2083 9.3005
R20420 vdd.n2067 vdd.n2066 9.3005
R20421 vdd.n2090 vdd.n2089 9.3005
R20422 vdd.n2092 vdd.n2091 9.3005
R20423 vdd.n2064 vdd.n2061 9.3005
R20424 vdd.n2099 vdd.n2098 9.3005
R20425 vdd.n1924 vdd.n1923 9.3005
R20426 vdd.n1919 vdd.n1918 9.3005
R20427 vdd.n1930 vdd.n1929 9.3005
R20428 vdd.n1932 vdd.n1931 9.3005
R20429 vdd.n1915 vdd.n1914 9.3005
R20430 vdd.n1938 vdd.n1937 9.3005
R20431 vdd.n1940 vdd.n1939 9.3005
R20432 vdd.n1912 vdd.n1909 9.3005
R20433 vdd.n1947 vdd.n1946 9.3005
R20434 vdd.n1979 vdd.n1978 9.3005
R20435 vdd.n1974 vdd.n1973 9.3005
R20436 vdd.n1985 vdd.n1984 9.3005
R20437 vdd.n1987 vdd.n1986 9.3005
R20438 vdd.n1970 vdd.n1969 9.3005
R20439 vdd.n1993 vdd.n1992 9.3005
R20440 vdd.n1995 vdd.n1994 9.3005
R20441 vdd.n1967 vdd.n1964 9.3005
R20442 vdd.n2002 vdd.n2001 9.3005
R20443 vdd.n1853 vdd.t91 9.18308
R20444 vdd.n3508 vdd.t167 9.18308
R20445 vdd.n1879 vdd.t97 8.95635
R20446 vdd.t68 vdd.n3549 8.95635
R20447 vdd.n300 vdd.n299 8.92171
R20448 vdd.n245 vdd.n244 8.92171
R20449 vdd.n202 vdd.n201 8.92171
R20450 vdd.n147 vdd.n146 8.92171
R20451 vdd.n105 vdd.n104 8.92171
R20452 vdd.n50 vdd.n49 8.92171
R20453 vdd.n2124 vdd.n2123 8.92171
R20454 vdd.n2179 vdd.n2178 8.92171
R20455 vdd.n2026 vdd.n2025 8.92171
R20456 vdd.n2081 vdd.n2080 8.92171
R20457 vdd.n1929 vdd.n1928 8.92171
R20458 vdd.n1984 vdd.n1983 8.92171
R20459 vdd.n223 vdd.n125 8.81535
R20460 vdd.n2102 vdd.n2004 8.81535
R20461 vdd.n1559 vdd.t105 8.72962
R20462 vdd.t60 vdd.n3558 8.72962
R20463 vdd.n2215 vdd.t81 8.50289
R20464 vdd.n3477 vdd.t66 8.50289
R20465 vdd.n28 vdd.n14 8.42249
R20466 vdd.n2231 vdd.t132 8.27616
R20467 vdd.t72 vdd.n636 8.27616
R20468 vdd.n3564 vdd.n3563 8.16225
R20469 vdd.n2202 vdd.n2201 8.16225
R20470 vdd.n296 vdd.n290 8.14595
R20471 vdd.n241 vdd.n235 8.14595
R20472 vdd.n198 vdd.n192 8.14595
R20473 vdd.n143 vdd.n137 8.14595
R20474 vdd.n101 vdd.n95 8.14595
R20475 vdd.n46 vdd.n40 8.14595
R20476 vdd.n2120 vdd.n2114 8.14595
R20477 vdd.n2175 vdd.n2169 8.14595
R20478 vdd.n2022 vdd.n2016 8.14595
R20479 vdd.n2077 vdd.n2071 8.14595
R20480 vdd.n1925 vdd.n1919 8.14595
R20481 vdd.n1980 vdd.n1974 8.14595
R20482 vdd.t242 vdd.n1593 7.8227
R20483 vdd.t215 vdd.n363 7.8227
R20484 vdd.n2430 vdd.n1105 7.70933
R20485 vdd.n2430 vdd.n1108 7.70933
R20486 vdd.n2436 vdd.n1094 7.70933
R20487 vdd.n2442 vdd.n1094 7.70933
R20488 vdd.n2442 vdd.n1087 7.70933
R20489 vdd.n2448 vdd.n1087 7.70933
R20490 vdd.n2448 vdd.n1090 7.70933
R20491 vdd.n2454 vdd.n1083 7.70933
R20492 vdd.n2460 vdd.n1077 7.70933
R20493 vdd.n2466 vdd.n1064 7.70933
R20494 vdd.n2472 vdd.n1064 7.70933
R20495 vdd.n2478 vdd.n1058 7.70933
R20496 vdd.n2484 vdd.n1051 7.70933
R20497 vdd.n2484 vdd.n1054 7.70933
R20498 vdd.n2490 vdd.n1047 7.70933
R20499 vdd.n2497 vdd.n1033 7.70933
R20500 vdd.n2503 vdd.n1033 7.70933
R20501 vdd.n2509 vdd.n1027 7.70933
R20502 vdd.n2515 vdd.n1023 7.70933
R20503 vdd.n2521 vdd.n1017 7.70933
R20504 vdd.n2539 vdd.n999 7.70933
R20505 vdd.n2539 vdd.n992 7.70933
R20506 vdd.n2547 vdd.n992 7.70933
R20507 vdd.n2629 vdd.n976 7.70933
R20508 vdd.n3012 vdd.n928 7.70933
R20509 vdd.n3024 vdd.n917 7.70933
R20510 vdd.n3024 vdd.n911 7.70933
R20511 vdd.n3030 vdd.n911 7.70933
R20512 vdd.n3042 vdd.n902 7.70933
R20513 vdd.n3048 vdd.n896 7.70933
R20514 vdd.n3060 vdd.n883 7.70933
R20515 vdd.n3067 vdd.n876 7.70933
R20516 vdd.n3067 vdd.n879 7.70933
R20517 vdd.n3073 vdd.n872 7.70933
R20518 vdd.n3079 vdd.n858 7.70933
R20519 vdd.n3085 vdd.n858 7.70933
R20520 vdd.n3091 vdd.n852 7.70933
R20521 vdd.n3097 vdd.n845 7.70933
R20522 vdd.n3097 vdd.n848 7.70933
R20523 vdd.n3103 vdd.n841 7.70933
R20524 vdd.n3109 vdd.n835 7.70933
R20525 vdd.n3115 vdd.n822 7.70933
R20526 vdd.n3121 vdd.n822 7.70933
R20527 vdd.n3121 vdd.n814 7.70933
R20528 vdd.n3172 vdd.n814 7.70933
R20529 vdd.n3172 vdd.n817 7.70933
R20530 vdd.n3178 vdd.n774 7.70933
R20531 vdd.n3248 vdd.n774 7.70933
R20532 vdd.n295 vdd.n292 7.3702
R20533 vdd.n240 vdd.n237 7.3702
R20534 vdd.n197 vdd.n194 7.3702
R20535 vdd.n142 vdd.n139 7.3702
R20536 vdd.n100 vdd.n97 7.3702
R20537 vdd.n45 vdd.n42 7.3702
R20538 vdd.n2119 vdd.n2116 7.3702
R20539 vdd.n2174 vdd.n2171 7.3702
R20540 vdd.n2021 vdd.n2018 7.3702
R20541 vdd.n2076 vdd.n2073 7.3702
R20542 vdd.n1924 vdd.n1921 7.3702
R20543 vdd.n1979 vdd.n1976 7.3702
R20544 vdd.n1077 vdd.t53 7.36923
R20545 vdd.n3103 vdd.t32 7.36923
R20546 vdd.n2454 vdd.t7 7.1425
R20547 vdd.n1396 vdd.t1 7.1425
R20548 vdd.n3036 vdd.t6 7.1425
R20549 vdd.n835 vdd.t16 7.1425
R20550 vdd.n1762 vdd.n1761 6.98232
R20551 vdd.n2318 vdd.n2317 6.98232
R20552 vdd.n547 vdd.n546 6.98232
R20553 vdd.n3332 vdd.n3331 6.98232
R20554 vdd.n2249 vdd.t130 6.91577
R20555 vdd.n3441 vdd.t95 6.91577
R20556 vdd.n1396 vdd.t2 6.80241
R20557 vdd.n3036 vdd.t46 6.80241
R20558 vdd.t86 vdd.n1530 6.68904
R20559 vdd.n3457 vdd.t146 6.68904
R20560 vdd.n2207 vdd.t62 6.46231
R20561 vdd.n2478 vdd.t14 6.46231
R20562 vdd.t19 vdd.n1027 6.46231
R20563 vdd.n3060 vdd.t24 6.46231
R20564 vdd.t38 vdd.n852 6.46231
R20565 vdd.n3485 vdd.t109 6.46231
R20566 vdd.n2554 vdd.t50 6.34895
R20567 vdd.n2933 vdd.t4 6.34895
R20568 vdd.n3564 vdd.n321 6.32949
R20569 vdd.n2201 vdd.n2200 6.32949
R20570 vdd.n3075 vdd.n868 6.2444
R20571 vdd.n2494 vdd.n2493 6.2444
R20572 vdd.t56 vdd.n1558 6.23558
R20573 vdd.t150 vdd.n332 6.23558
R20574 vdd.n1871 vdd.t116 6.00885
R20575 vdd.n3543 vdd.t114 6.00885
R20576 vdd.n2515 vdd.t43 5.89549
R20577 vdd.n896 vdd.t20 5.89549
R20578 vdd.n296 vdd.n295 5.81868
R20579 vdd.n241 vdd.n240 5.81868
R20580 vdd.n198 vdd.n197 5.81868
R20581 vdd.n143 vdd.n142 5.81868
R20582 vdd.n101 vdd.n100 5.81868
R20583 vdd.n46 vdd.n45 5.81868
R20584 vdd.n2120 vdd.n2119 5.81868
R20585 vdd.n2175 vdd.n2174 5.81868
R20586 vdd.n2022 vdd.n2021 5.81868
R20587 vdd.n2077 vdd.n2076 5.81868
R20588 vdd.n1925 vdd.n1924 5.81868
R20589 vdd.n1980 vdd.n1979 5.81868
R20590 vdd.n2637 vdd.n2636 5.77611
R20591 vdd.n1320 vdd.n1319 5.77611
R20592 vdd.n2945 vdd.n2944 5.77611
R20593 vdd.n3187 vdd.n806 5.77611
R20594 vdd.n3253 vdd.n770 5.77611
R20595 vdd.n2808 vdd.n2742 5.77611
R20596 vdd.n2562 vdd.n983 5.77611
R20597 vdd.n1456 vdd.n1288 5.77611
R20598 vdd.n1831 vdd.n1605 5.62474
R20599 vdd.n2281 vdd.n2278 5.62474
R20600 vdd.n3522 vdd.n407 5.62474
R20601 vdd.n3287 vdd.n3284 5.62474
R20602 vdd.n2490 vdd.t34 5.55539
R20603 vdd.n872 vdd.t10 5.55539
R20604 vdd.n1581 vdd.t116 5.32866
R20605 vdd.t114 vdd.n3542 5.32866
R20606 vdd.n1887 vdd.t56 5.10193
R20607 vdd.n3551 vdd.t150 5.10193
R20608 vdd.n299 vdd.n290 5.04292
R20609 vdd.n244 vdd.n235 5.04292
R20610 vdd.n201 vdd.n192 5.04292
R20611 vdd.n146 vdd.n137 5.04292
R20612 vdd.n104 vdd.n95 5.04292
R20613 vdd.n49 vdd.n40 5.04292
R20614 vdd.n2123 vdd.n2114 5.04292
R20615 vdd.n2178 vdd.n2169 5.04292
R20616 vdd.n2025 vdd.n2016 5.04292
R20617 vdd.n2080 vdd.n2071 5.04292
R20618 vdd.n1928 vdd.n1919 5.04292
R20619 vdd.n1983 vdd.n1974 5.04292
R20620 vdd.n1903 vdd.t62 4.8752
R20621 vdd.t13 vdd.t26 4.8752
R20622 vdd.t54 vdd.t0 4.8752
R20623 vdd.t109 vdd.n328 4.8752
R20624 vdd.n2638 vdd.n2637 4.83952
R20625 vdd.n1319 vdd.n1318 4.83952
R20626 vdd.n2946 vdd.n2945 4.83952
R20627 vdd.n806 vdd.n801 4.83952
R20628 vdd.n770 vdd.n765 4.83952
R20629 vdd.n2805 vdd.n2742 4.83952
R20630 vdd.n2565 vdd.n983 4.83952
R20631 vdd.n1459 vdd.n1288 4.83952
R20632 vdd.n1370 vdd.t22 4.76184
R20633 vdd.n3018 vdd.t8 4.76184
R20634 vdd.n2286 vdd.n2285 4.74817
R20635 vdd.n1492 vdd.n1487 4.74817
R20636 vdd.n1154 vdd.n1151 4.74817
R20637 vdd.n2379 vdd.n1150 4.74817
R20638 vdd.n2384 vdd.n1151 4.74817
R20639 vdd.n2383 vdd.n1150 4.74817
R20640 vdd.n664 vdd.n662 4.74817
R20641 vdd.n3402 vdd.n665 4.74817
R20642 vdd.n3405 vdd.n665 4.74817
R20643 vdd.n3406 vdd.n664 4.74817
R20644 vdd.n3294 vdd.n749 4.74817
R20645 vdd.n3290 vdd.n751 4.74817
R20646 vdd.n3293 vdd.n751 4.74817
R20647 vdd.n3298 vdd.n749 4.74817
R20648 vdd.n2285 vdd.n1250 4.74817
R20649 vdd.n1489 vdd.n1487 4.74817
R20650 vdd.n321 vdd.n320 4.7074
R20651 vdd.n223 vdd.n222 4.7074
R20652 vdd.n2200 vdd.n2199 4.7074
R20653 vdd.n2102 vdd.n2101 4.7074
R20654 vdd.n2223 vdd.t86 4.64847
R20655 vdd.t15 vdd.n1058 4.64847
R20656 vdd.n2509 vdd.t52 4.64847
R20657 vdd.t41 vdd.n883 4.64847
R20658 vdd.n3091 vdd.t37 4.64847
R20659 vdd.n3466 vdd.t146 4.64847
R20660 vdd.n1047 vdd.t260 4.53511
R20661 vdd.n3073 vdd.t223 4.53511
R20662 vdd.n1524 vdd.t130 4.42174
R20663 vdd.n2436 vdd.t201 4.42174
R20664 vdd.n1370 vdd.t246 4.42174
R20665 vdd.n3018 vdd.t253 4.42174
R20666 vdd.n817 vdd.t197 4.42174
R20667 vdd.t95 vdd.n635 4.42174
R20668 vdd.n3064 vdd.n868 4.37123
R20669 vdd.n2495 vdd.n2494 4.37123
R20670 vdd.n2533 vdd.t39 4.30838
R20671 vdd.n2921 vdd.t28 4.30838
R20672 vdd.n300 vdd.n288 4.26717
R20673 vdd.n245 vdd.n233 4.26717
R20674 vdd.n202 vdd.n190 4.26717
R20675 vdd.n147 vdd.n135 4.26717
R20676 vdd.n105 vdd.n93 4.26717
R20677 vdd.n50 vdd.n38 4.26717
R20678 vdd.n2124 vdd.n2112 4.26717
R20679 vdd.n2179 vdd.n2167 4.26717
R20680 vdd.n2026 vdd.n2014 4.26717
R20681 vdd.n2081 vdd.n2069 4.26717
R20682 vdd.n1929 vdd.n1917 4.26717
R20683 vdd.n1984 vdd.n1972 4.26717
R20684 vdd.n321 vdd.n223 4.10845
R20685 vdd.n2200 vdd.n2102 4.10845
R20686 vdd.n277 vdd.t143 4.06363
R20687 vdd.n277 vdd.t178 4.06363
R20688 vdd.n275 vdd.t69 4.06363
R20689 vdd.n275 vdd.t112 4.06363
R20690 vdd.n273 vdd.t113 4.06363
R20691 vdd.n273 vdd.t158 4.06363
R20692 vdd.n271 vdd.t160 4.06363
R20693 vdd.n271 vdd.t61 4.06363
R20694 vdd.n269 vdd.t85 4.06363
R20695 vdd.n269 vdd.t138 4.06363
R20696 vdd.n267 vdd.t161 4.06363
R20697 vdd.n267 vdd.t174 4.06363
R20698 vdd.n265 vdd.t179 4.06363
R20699 vdd.n265 vdd.t78 4.06363
R20700 vdd.n179 vdd.t136 4.06363
R20701 vdd.n179 vdd.t168 4.06363
R20702 vdd.n177 vdd.t182 4.06363
R20703 vdd.n177 vdd.t94 4.06363
R20704 vdd.n175 vdd.t103 4.06363
R20705 vdd.n175 vdd.t151 4.06363
R20706 vdd.n173 vdd.t152 4.06363
R20707 vdd.n173 vdd.t175 4.06363
R20708 vdd.n171 vdd.t67 4.06363
R20709 vdd.n171 vdd.t120 4.06363
R20710 vdd.n169 vdd.t155 4.06363
R20711 vdd.n169 vdd.t162 4.06363
R20712 vdd.n167 vdd.t170 4.06363
R20713 vdd.n167 vdd.t73 4.06363
R20714 vdd.n82 vdd.t115 4.06363
R20715 vdd.n82 vdd.t180 4.06363
R20716 vdd.n80 vdd.t100 4.06363
R20717 vdd.n80 vdd.t165 4.06363
R20718 vdd.n78 vdd.t125 4.06363
R20719 vdd.n78 vdd.t153 4.06363
R20720 vdd.n76 vdd.t110 4.06363
R20721 vdd.n76 vdd.t172 4.06363
R20722 vdd.n74 vdd.t77 4.06363
R20723 vdd.n74 vdd.t159 4.06363
R20724 vdd.n72 vdd.t76 4.06363
R20725 vdd.n72 vdd.t147 4.06363
R20726 vdd.n70 vdd.t96 4.06363
R20727 vdd.n70 vdd.t163 4.06363
R20728 vdd.n2144 vdd.t142 4.06363
R20729 vdd.n2144 vdd.t141 4.06363
R20730 vdd.n2146 vdd.t104 4.06363
R20731 vdd.n2146 vdd.t84 4.06363
R20732 vdd.n2148 vdd.t80 4.06363
R20733 vdd.n2148 vdd.t140 4.06363
R20734 vdd.n2150 vdd.t118 4.06363
R20735 vdd.n2150 vdd.t83 4.06363
R20736 vdd.n2152 vdd.t74 4.06363
R20737 vdd.n2152 vdd.t157 4.06363
R20738 vdd.n2154 vdd.t156 4.06363
R20739 vdd.n2154 vdd.t98 4.06363
R20740 vdd.n2156 vdd.t108 4.06363
R20741 vdd.n2156 vdd.t181 4.06363
R20742 vdd.n2046 vdd.t133 4.06363
R20743 vdd.n2046 vdd.t131 4.06363
R20744 vdd.n2048 vdd.t87 4.06363
R20745 vdd.n2048 vdd.t65 4.06363
R20746 vdd.n2050 vdd.t59 4.06363
R20747 vdd.n2050 vdd.t127 4.06363
R20748 vdd.n2052 vdd.t106 4.06363
R20749 vdd.n2052 vdd.t63 4.06363
R20750 vdd.n2054 vdd.t57 4.06363
R20751 vdd.n2054 vdd.t149 4.06363
R20752 vdd.n2056 vdd.t145 4.06363
R20753 vdd.n2056 vdd.t101 4.06363
R20754 vdd.n2058 vdd.t92 4.06363
R20755 vdd.n2058 vdd.t171 4.06363
R20756 vdd.n1949 vdd.t164 4.06363
R20757 vdd.n1949 vdd.t183 4.06363
R20758 vdd.n1951 vdd.t148 4.06363
R20759 vdd.n1951 vdd.t79 4.06363
R20760 vdd.n1953 vdd.t134 4.06363
R20761 vdd.n1953 vdd.t82 4.06363
R20762 vdd.n1955 vdd.t173 4.06363
R20763 vdd.n1955 vdd.t111 4.06363
R20764 vdd.n1957 vdd.t154 4.06363
R20765 vdd.n1957 vdd.t129 4.06363
R20766 vdd.n1959 vdd.t166 4.06363
R20767 vdd.n1959 vdd.t99 4.06363
R20768 vdd.n1961 vdd.t176 4.06363
R20769 vdd.n1961 vdd.t117 4.06363
R20770 vdd.n1083 vdd.t45 3.96828
R20771 vdd.n2527 vdd.t25 3.96828
R20772 vdd.n2915 vdd.t42 3.96828
R20773 vdd.n3109 vdd.t33 3.96828
R20774 vdd.n26 vdd.t191 3.9605
R20775 vdd.n26 vdd.t194 3.9605
R20776 vdd.n23 vdd.t187 3.9605
R20777 vdd.n23 vdd.t275 3.9605
R20778 vdd.n21 vdd.t273 3.9605
R20779 vdd.n21 vdd.t185 3.9605
R20780 vdd.n20 vdd.t189 3.9605
R20781 vdd.n20 vdd.t186 3.9605
R20782 vdd.n15 vdd.t272 3.9605
R20783 vdd.n15 vdd.t190 3.9605
R20784 vdd.n16 vdd.t195 3.9605
R20785 vdd.n16 vdd.t192 3.9605
R20786 vdd.n18 vdd.t274 3.9605
R20787 vdd.n18 vdd.t188 3.9605
R20788 vdd.n25 vdd.t193 3.9605
R20789 vdd.n25 vdd.t184 3.9605
R20790 vdd.n2460 vdd.t45 3.74155
R20791 vdd.n1017 vdd.t25 3.74155
R20792 vdd.n3042 vdd.t42 3.74155
R20793 vdd.n841 vdd.t33 3.74155
R20794 vdd.n7 vdd.t55 3.61217
R20795 vdd.n7 vdd.t21 3.61217
R20796 vdd.n8 vdd.t29 3.61217
R20797 vdd.n8 vdd.t47 3.61217
R20798 vdd.n10 vdd.t5 3.61217
R20799 vdd.n10 vdd.t9 3.61217
R20800 vdd.n12 vdd.t18 3.61217
R20801 vdd.n12 vdd.t36 3.61217
R20802 vdd.n5 vdd.t49 3.61217
R20803 vdd.n5 vdd.t31 3.61217
R20804 vdd.n3 vdd.t23 3.61217
R20805 vdd.n3 vdd.t51 3.61217
R20806 vdd.n1 vdd.t3 3.61217
R20807 vdd.n1 vdd.t40 3.61217
R20808 vdd.n0 vdd.t44 3.61217
R20809 vdd.n0 vdd.t27 3.61217
R20810 vdd.n1837 vdd.t242 3.51482
R20811 vdd.n3527 vdd.t215 3.51482
R20812 vdd.n304 vdd.n303 3.49141
R20813 vdd.n249 vdd.n248 3.49141
R20814 vdd.n206 vdd.n205 3.49141
R20815 vdd.n151 vdd.n150 3.49141
R20816 vdd.n109 vdd.n108 3.49141
R20817 vdd.n54 vdd.n53 3.49141
R20818 vdd.n2128 vdd.n2127 3.49141
R20819 vdd.n2183 vdd.n2182 3.49141
R20820 vdd.n2030 vdd.n2029 3.49141
R20821 vdd.n2085 vdd.n2084 3.49141
R20822 vdd.n1933 vdd.n1932 3.49141
R20823 vdd.n1988 vdd.n1987 3.49141
R20824 vdd.t39 vdd.n999 3.40145
R20825 vdd.n2701 vdd.t48 3.40145
R20826 vdd.n3005 vdd.t35 3.40145
R20827 vdd.n3030 vdd.t28 3.40145
R20828 vdd.n1108 vdd.t201 3.28809
R20829 vdd.n2554 vdd.t246 3.28809
R20830 vdd.n2933 vdd.t253 3.28809
R20831 vdd.n3178 vdd.t197 3.28809
R20832 vdd.n2240 vdd.t132 3.06136
R20833 vdd.n2472 vdd.t15 3.06136
R20834 vdd.n1408 vdd.t52 3.06136
R20835 vdd.n3054 vdd.t41 3.06136
R20836 vdd.t37 vdd.n845 3.06136
R20837 vdd.n3449 vdd.t72 3.06136
R20838 vdd.n2547 vdd.t22 2.94799
R20839 vdd.t8 vdd.n917 2.94799
R20840 vdd.t81 vdd.n1536 2.83463
R20841 vdd.n624 vdd.t66 2.83463
R20842 vdd.n307 vdd.n286 2.71565
R20843 vdd.n252 vdd.n231 2.71565
R20844 vdd.n209 vdd.n188 2.71565
R20845 vdd.n154 vdd.n133 2.71565
R20846 vdd.n112 vdd.n91 2.71565
R20847 vdd.n57 vdd.n36 2.71565
R20848 vdd.n2131 vdd.n2110 2.71565
R20849 vdd.n2186 vdd.n2165 2.71565
R20850 vdd.n2033 vdd.n2012 2.71565
R20851 vdd.n2088 vdd.n2067 2.71565
R20852 vdd.n1936 vdd.n1915 2.71565
R20853 vdd.n1991 vdd.n1970 2.71565
R20854 vdd.n1904 vdd.t105 2.6079
R20855 vdd.n3559 vdd.t60 2.6079
R20856 vdd.n2521 vdd.t26 2.49453
R20857 vdd.n902 vdd.t54 2.49453
R20858 vdd.n294 vdd.n293 2.4129
R20859 vdd.n239 vdd.n238 2.4129
R20860 vdd.n196 vdd.n195 2.4129
R20861 vdd.n141 vdd.n140 2.4129
R20862 vdd.n99 vdd.n98 2.4129
R20863 vdd.n44 vdd.n43 2.4129
R20864 vdd.n2118 vdd.n2117 2.4129
R20865 vdd.n2173 vdd.n2172 2.4129
R20866 vdd.n2020 vdd.n2019 2.4129
R20867 vdd.n2075 vdd.n2074 2.4129
R20868 vdd.n1923 vdd.n1922 2.4129
R20869 vdd.n1978 vdd.n1977 2.4129
R20870 vdd.t97 vdd.n1565 2.38117
R20871 vdd.n3550 vdd.t68 2.38117
R20872 vdd.n2391 vdd.n1151 2.27742
R20873 vdd.n2391 vdd.n1150 2.27742
R20874 vdd.n3214 vdd.n665 2.27742
R20875 vdd.n3214 vdd.n664 2.27742
R20876 vdd.n3282 vdd.n751 2.27742
R20877 vdd.n3282 vdd.n749 2.27742
R20878 vdd.n2285 vdd.n2284 2.27742
R20879 vdd.n2284 vdd.n1487 2.27742
R20880 vdd.n1862 vdd.t91 2.15444
R20881 vdd.n1054 vdd.t34 2.15444
R20882 vdd.n2497 vdd.t12 2.15444
R20883 vdd.n879 vdd.t11 2.15444
R20884 vdd.n3079 vdd.t10 2.15444
R20885 vdd.n3541 vdd.t167 2.15444
R20886 vdd.n308 vdd.n284 1.93989
R20887 vdd.n253 vdd.n229 1.93989
R20888 vdd.n210 vdd.n186 1.93989
R20889 vdd.n155 vdd.n131 1.93989
R20890 vdd.n113 vdd.n89 1.93989
R20891 vdd.n58 vdd.n34 1.93989
R20892 vdd.n2132 vdd.n2108 1.93989
R20893 vdd.n2187 vdd.n2163 1.93989
R20894 vdd.n2034 vdd.n2010 1.93989
R20895 vdd.n2089 vdd.n2065 1.93989
R20896 vdd.n1937 vdd.n1913 1.93989
R20897 vdd.n1992 vdd.n1968 1.93989
R20898 vdd.n1408 vdd.t43 1.81434
R20899 vdd.n3054 vdd.t20 1.81434
R20900 vdd.n1854 vdd.t123 1.70098
R20901 vdd.n3535 vdd.t70 1.70098
R20902 vdd.n1870 vdd.t144 1.47425
R20903 vdd.n349 vdd.t93 1.47425
R20904 vdd.t50 vdd.n976 1.36088
R20905 vdd.n3012 vdd.t4 1.36088
R20906 vdd.n1895 vdd.t128 1.24752
R20907 vdd.t205 vdd.n1500 1.24752
R20908 vdd.t14 vdd.n1051 1.24752
R20909 vdd.n2503 vdd.t19 1.24752
R20910 vdd.t24 vdd.n876 1.24752
R20911 vdd.n3085 vdd.t38 1.24752
R20912 vdd.n659 vdd.t219 1.24752
R20913 vdd.t102 vdd.n3557 1.24752
R20914 vdd.n2201 vdd.n28 1.16438
R20915 vdd.n319 vdd.n279 1.16414
R20916 vdd.n312 vdd.n311 1.16414
R20917 vdd.n264 vdd.n224 1.16414
R20918 vdd.n257 vdd.n256 1.16414
R20919 vdd.n221 vdd.n181 1.16414
R20920 vdd.n214 vdd.n213 1.16414
R20921 vdd.n166 vdd.n126 1.16414
R20922 vdd.n159 vdd.n158 1.16414
R20923 vdd.n124 vdd.n84 1.16414
R20924 vdd.n117 vdd.n116 1.16414
R20925 vdd.n69 vdd.n29 1.16414
R20926 vdd.n62 vdd.n61 1.16414
R20927 vdd.n2143 vdd.n2103 1.16414
R20928 vdd.n2136 vdd.n2135 1.16414
R20929 vdd.n2198 vdd.n2158 1.16414
R20930 vdd.n2191 vdd.n2190 1.16414
R20931 vdd.n2045 vdd.n2005 1.16414
R20932 vdd.n2038 vdd.n2037 1.16414
R20933 vdd.n2100 vdd.n2060 1.16414
R20934 vdd.n2093 vdd.n2092 1.16414
R20935 vdd.n1948 vdd.n1908 1.16414
R20936 vdd.n1941 vdd.n1940 1.16414
R20937 vdd.n2003 vdd.n1963 1.16414
R20938 vdd.n1996 vdd.n1995 1.16414
R20939 vdd vdd.n3564 1.15654
R20940 vdd.n1547 vdd.t58 1.02079
R20941 vdd.t260 vdd.t12 1.02079
R20942 vdd.t11 vdd.t223 1.02079
R20943 vdd.t119 vdd.n613 1.02079
R20944 vdd.n1726 vdd.n1605 0.970197
R20945 vdd.n2282 vdd.n2281 0.970197
R20946 vdd.n599 vdd.n407 0.970197
R20947 vdd.n3289 vdd.n3287 0.970197
R20948 vdd.n2527 vdd.t2 0.907421
R20949 vdd.n2915 vdd.t46 0.907421
R20950 vdd.n2232 vdd.t64 0.794056
R20951 vdd.n3458 vdd.t75 0.794056
R20952 vdd.n2248 vdd.t89 0.567326
R20953 vdd.n1090 vdd.t7 0.567326
R20954 vdd.n2533 vdd.t1 0.567326
R20955 vdd.n2921 vdd.t6 0.567326
R20956 vdd.n3115 vdd.t16 0.567326
R20957 vdd.t121 vdd.n642 0.567326
R20958 vdd.n2272 vdd.n1152 0.482207
R20959 vdd.n3414 vdd.n3413 0.482207
R20960 vdd.n444 vdd.n443 0.482207
R20961 vdd.n3521 vdd.n3520 0.482207
R20962 vdd.n3420 vdd.n656 0.482207
R20963 vdd.n2262 vdd.n1488 0.482207
R20964 vdd.n1833 vdd.n1832 0.482207
R20965 vdd.n1639 vdd.n1596 0.482207
R20966 vdd.n4 vdd.n2 0.459552
R20967 vdd.n11 vdd.n9 0.459552
R20968 vdd.n317 vdd.n316 0.388379
R20969 vdd.n283 vdd.n281 0.388379
R20970 vdd.n262 vdd.n261 0.388379
R20971 vdd.n228 vdd.n226 0.388379
R20972 vdd.n219 vdd.n218 0.388379
R20973 vdd.n185 vdd.n183 0.388379
R20974 vdd.n164 vdd.n163 0.388379
R20975 vdd.n130 vdd.n128 0.388379
R20976 vdd.n122 vdd.n121 0.388379
R20977 vdd.n88 vdd.n86 0.388379
R20978 vdd.n67 vdd.n66 0.388379
R20979 vdd.n33 vdd.n31 0.388379
R20980 vdd.n2141 vdd.n2140 0.388379
R20981 vdd.n2107 vdd.n2105 0.388379
R20982 vdd.n2196 vdd.n2195 0.388379
R20983 vdd.n2162 vdd.n2160 0.388379
R20984 vdd.n2043 vdd.n2042 0.388379
R20985 vdd.n2009 vdd.n2007 0.388379
R20986 vdd.n2098 vdd.n2097 0.388379
R20987 vdd.n2064 vdd.n2062 0.388379
R20988 vdd.n1946 vdd.n1945 0.388379
R20989 vdd.n1912 vdd.n1910 0.388379
R20990 vdd.n2001 vdd.n2000 0.388379
R20991 vdd.n1967 vdd.n1965 0.388379
R20992 vdd.n19 vdd.n17 0.387128
R20993 vdd.n24 vdd.n22 0.387128
R20994 vdd.n6 vdd.n4 0.358259
R20995 vdd.n13 vdd.n11 0.358259
R20996 vdd.n268 vdd.n266 0.358259
R20997 vdd.n270 vdd.n268 0.358259
R20998 vdd.n272 vdd.n270 0.358259
R20999 vdd.n274 vdd.n272 0.358259
R21000 vdd.n276 vdd.n274 0.358259
R21001 vdd.n278 vdd.n276 0.358259
R21002 vdd.n320 vdd.n278 0.358259
R21003 vdd.n170 vdd.n168 0.358259
R21004 vdd.n172 vdd.n170 0.358259
R21005 vdd.n174 vdd.n172 0.358259
R21006 vdd.n176 vdd.n174 0.358259
R21007 vdd.n178 vdd.n176 0.358259
R21008 vdd.n180 vdd.n178 0.358259
R21009 vdd.n222 vdd.n180 0.358259
R21010 vdd.n73 vdd.n71 0.358259
R21011 vdd.n75 vdd.n73 0.358259
R21012 vdd.n77 vdd.n75 0.358259
R21013 vdd.n79 vdd.n77 0.358259
R21014 vdd.n81 vdd.n79 0.358259
R21015 vdd.n83 vdd.n81 0.358259
R21016 vdd.n125 vdd.n83 0.358259
R21017 vdd.n2199 vdd.n2157 0.358259
R21018 vdd.n2157 vdd.n2155 0.358259
R21019 vdd.n2155 vdd.n2153 0.358259
R21020 vdd.n2153 vdd.n2151 0.358259
R21021 vdd.n2151 vdd.n2149 0.358259
R21022 vdd.n2149 vdd.n2147 0.358259
R21023 vdd.n2147 vdd.n2145 0.358259
R21024 vdd.n2101 vdd.n2059 0.358259
R21025 vdd.n2059 vdd.n2057 0.358259
R21026 vdd.n2057 vdd.n2055 0.358259
R21027 vdd.n2055 vdd.n2053 0.358259
R21028 vdd.n2053 vdd.n2051 0.358259
R21029 vdd.n2051 vdd.n2049 0.358259
R21030 vdd.n2049 vdd.n2047 0.358259
R21031 vdd.n2004 vdd.n1962 0.358259
R21032 vdd.n1962 vdd.n1960 0.358259
R21033 vdd.n1960 vdd.n1958 0.358259
R21034 vdd.n1958 vdd.n1956 0.358259
R21035 vdd.n1956 vdd.n1954 0.358259
R21036 vdd.n1954 vdd.n1952 0.358259
R21037 vdd.n1952 vdd.n1950 0.358259
R21038 vdd.n2466 vdd.t53 0.340595
R21039 vdd.n1023 vdd.t13 0.340595
R21040 vdd.n3048 vdd.t0 0.340595
R21041 vdd.n848 vdd.t32 0.340595
R21042 vdd.n14 vdd.n6 0.334552
R21043 vdd.n14 vdd.n13 0.334552
R21044 vdd.n27 vdd.n19 0.21707
R21045 vdd.n27 vdd.n24 0.21707
R21046 vdd.n318 vdd.n280 0.155672
R21047 vdd.n310 vdd.n280 0.155672
R21048 vdd.n310 vdd.n309 0.155672
R21049 vdd.n309 vdd.n285 0.155672
R21050 vdd.n302 vdd.n285 0.155672
R21051 vdd.n302 vdd.n301 0.155672
R21052 vdd.n301 vdd.n289 0.155672
R21053 vdd.n294 vdd.n289 0.155672
R21054 vdd.n263 vdd.n225 0.155672
R21055 vdd.n255 vdd.n225 0.155672
R21056 vdd.n255 vdd.n254 0.155672
R21057 vdd.n254 vdd.n230 0.155672
R21058 vdd.n247 vdd.n230 0.155672
R21059 vdd.n247 vdd.n246 0.155672
R21060 vdd.n246 vdd.n234 0.155672
R21061 vdd.n239 vdd.n234 0.155672
R21062 vdd.n220 vdd.n182 0.155672
R21063 vdd.n212 vdd.n182 0.155672
R21064 vdd.n212 vdd.n211 0.155672
R21065 vdd.n211 vdd.n187 0.155672
R21066 vdd.n204 vdd.n187 0.155672
R21067 vdd.n204 vdd.n203 0.155672
R21068 vdd.n203 vdd.n191 0.155672
R21069 vdd.n196 vdd.n191 0.155672
R21070 vdd.n165 vdd.n127 0.155672
R21071 vdd.n157 vdd.n127 0.155672
R21072 vdd.n157 vdd.n156 0.155672
R21073 vdd.n156 vdd.n132 0.155672
R21074 vdd.n149 vdd.n132 0.155672
R21075 vdd.n149 vdd.n148 0.155672
R21076 vdd.n148 vdd.n136 0.155672
R21077 vdd.n141 vdd.n136 0.155672
R21078 vdd.n123 vdd.n85 0.155672
R21079 vdd.n115 vdd.n85 0.155672
R21080 vdd.n115 vdd.n114 0.155672
R21081 vdd.n114 vdd.n90 0.155672
R21082 vdd.n107 vdd.n90 0.155672
R21083 vdd.n107 vdd.n106 0.155672
R21084 vdd.n106 vdd.n94 0.155672
R21085 vdd.n99 vdd.n94 0.155672
R21086 vdd.n68 vdd.n30 0.155672
R21087 vdd.n60 vdd.n30 0.155672
R21088 vdd.n60 vdd.n59 0.155672
R21089 vdd.n59 vdd.n35 0.155672
R21090 vdd.n52 vdd.n35 0.155672
R21091 vdd.n52 vdd.n51 0.155672
R21092 vdd.n51 vdd.n39 0.155672
R21093 vdd.n44 vdd.n39 0.155672
R21094 vdd.n2142 vdd.n2104 0.155672
R21095 vdd.n2134 vdd.n2104 0.155672
R21096 vdd.n2134 vdd.n2133 0.155672
R21097 vdd.n2133 vdd.n2109 0.155672
R21098 vdd.n2126 vdd.n2109 0.155672
R21099 vdd.n2126 vdd.n2125 0.155672
R21100 vdd.n2125 vdd.n2113 0.155672
R21101 vdd.n2118 vdd.n2113 0.155672
R21102 vdd.n2197 vdd.n2159 0.155672
R21103 vdd.n2189 vdd.n2159 0.155672
R21104 vdd.n2189 vdd.n2188 0.155672
R21105 vdd.n2188 vdd.n2164 0.155672
R21106 vdd.n2181 vdd.n2164 0.155672
R21107 vdd.n2181 vdd.n2180 0.155672
R21108 vdd.n2180 vdd.n2168 0.155672
R21109 vdd.n2173 vdd.n2168 0.155672
R21110 vdd.n2044 vdd.n2006 0.155672
R21111 vdd.n2036 vdd.n2006 0.155672
R21112 vdd.n2036 vdd.n2035 0.155672
R21113 vdd.n2035 vdd.n2011 0.155672
R21114 vdd.n2028 vdd.n2011 0.155672
R21115 vdd.n2028 vdd.n2027 0.155672
R21116 vdd.n2027 vdd.n2015 0.155672
R21117 vdd.n2020 vdd.n2015 0.155672
R21118 vdd.n2099 vdd.n2061 0.155672
R21119 vdd.n2091 vdd.n2061 0.155672
R21120 vdd.n2091 vdd.n2090 0.155672
R21121 vdd.n2090 vdd.n2066 0.155672
R21122 vdd.n2083 vdd.n2066 0.155672
R21123 vdd.n2083 vdd.n2082 0.155672
R21124 vdd.n2082 vdd.n2070 0.155672
R21125 vdd.n2075 vdd.n2070 0.155672
R21126 vdd.n1947 vdd.n1909 0.155672
R21127 vdd.n1939 vdd.n1909 0.155672
R21128 vdd.n1939 vdd.n1938 0.155672
R21129 vdd.n1938 vdd.n1914 0.155672
R21130 vdd.n1931 vdd.n1914 0.155672
R21131 vdd.n1931 vdd.n1930 0.155672
R21132 vdd.n1930 vdd.n1918 0.155672
R21133 vdd.n1923 vdd.n1918 0.155672
R21134 vdd.n2002 vdd.n1964 0.155672
R21135 vdd.n1994 vdd.n1964 0.155672
R21136 vdd.n1994 vdd.n1993 0.155672
R21137 vdd.n1993 vdd.n1969 0.155672
R21138 vdd.n1986 vdd.n1969 0.155672
R21139 vdd.n1986 vdd.n1985 0.155672
R21140 vdd.n1985 vdd.n1973 0.155672
R21141 vdd.n1978 vdd.n1973 0.155672
R21142 vdd.n1157 vdd.n1149 0.152939
R21143 vdd.n1161 vdd.n1157 0.152939
R21144 vdd.n1162 vdd.n1161 0.152939
R21145 vdd.n1163 vdd.n1162 0.152939
R21146 vdd.n1164 vdd.n1163 0.152939
R21147 vdd.n1168 vdd.n1164 0.152939
R21148 vdd.n1169 vdd.n1168 0.152939
R21149 vdd.n1170 vdd.n1169 0.152939
R21150 vdd.n1171 vdd.n1170 0.152939
R21151 vdd.n1175 vdd.n1171 0.152939
R21152 vdd.n1176 vdd.n1175 0.152939
R21153 vdd.n1177 vdd.n1176 0.152939
R21154 vdd.n2355 vdd.n1177 0.152939
R21155 vdd.n2355 vdd.n2354 0.152939
R21156 vdd.n2354 vdd.n2353 0.152939
R21157 vdd.n2353 vdd.n1183 0.152939
R21158 vdd.n1188 vdd.n1183 0.152939
R21159 vdd.n1189 vdd.n1188 0.152939
R21160 vdd.n1190 vdd.n1189 0.152939
R21161 vdd.n1194 vdd.n1190 0.152939
R21162 vdd.n1195 vdd.n1194 0.152939
R21163 vdd.n1196 vdd.n1195 0.152939
R21164 vdd.n1197 vdd.n1196 0.152939
R21165 vdd.n1201 vdd.n1197 0.152939
R21166 vdd.n1202 vdd.n1201 0.152939
R21167 vdd.n1203 vdd.n1202 0.152939
R21168 vdd.n1204 vdd.n1203 0.152939
R21169 vdd.n1208 vdd.n1204 0.152939
R21170 vdd.n1209 vdd.n1208 0.152939
R21171 vdd.n1210 vdd.n1209 0.152939
R21172 vdd.n1211 vdd.n1210 0.152939
R21173 vdd.n1215 vdd.n1211 0.152939
R21174 vdd.n1216 vdd.n1215 0.152939
R21175 vdd.n1217 vdd.n1216 0.152939
R21176 vdd.n2316 vdd.n1217 0.152939
R21177 vdd.n2316 vdd.n2315 0.152939
R21178 vdd.n2315 vdd.n2314 0.152939
R21179 vdd.n2314 vdd.n1223 0.152939
R21180 vdd.n1228 vdd.n1223 0.152939
R21181 vdd.n1229 vdd.n1228 0.152939
R21182 vdd.n1230 vdd.n1229 0.152939
R21183 vdd.n1234 vdd.n1230 0.152939
R21184 vdd.n1235 vdd.n1234 0.152939
R21185 vdd.n1236 vdd.n1235 0.152939
R21186 vdd.n1237 vdd.n1236 0.152939
R21187 vdd.n1241 vdd.n1237 0.152939
R21188 vdd.n1242 vdd.n1241 0.152939
R21189 vdd.n1243 vdd.n1242 0.152939
R21190 vdd.n1244 vdd.n1243 0.152939
R21191 vdd.n1248 vdd.n1244 0.152939
R21192 vdd.n1249 vdd.n1248 0.152939
R21193 vdd.n2390 vdd.n1152 0.152939
R21194 vdd.n2204 vdd.n2203 0.152939
R21195 vdd.n2204 vdd.n1539 0.152939
R21196 vdd.n2218 vdd.n1539 0.152939
R21197 vdd.n2219 vdd.n2218 0.152939
R21198 vdd.n2220 vdd.n2219 0.152939
R21199 vdd.n2220 vdd.n1527 0.152939
R21200 vdd.n2235 vdd.n1527 0.152939
R21201 vdd.n2236 vdd.n2235 0.152939
R21202 vdd.n2237 vdd.n2236 0.152939
R21203 vdd.n2237 vdd.n1516 0.152939
R21204 vdd.n2252 vdd.n1516 0.152939
R21205 vdd.n2253 vdd.n2252 0.152939
R21206 vdd.n2254 vdd.n2253 0.152939
R21207 vdd.n2254 vdd.n1504 0.152939
R21208 vdd.n2270 vdd.n1504 0.152939
R21209 vdd.n2271 vdd.n2270 0.152939
R21210 vdd.n2272 vdd.n2271 0.152939
R21211 vdd.n670 vdd.n667 0.152939
R21212 vdd.n671 vdd.n670 0.152939
R21213 vdd.n672 vdd.n671 0.152939
R21214 vdd.n673 vdd.n672 0.152939
R21215 vdd.n676 vdd.n673 0.152939
R21216 vdd.n677 vdd.n676 0.152939
R21217 vdd.n678 vdd.n677 0.152939
R21218 vdd.n679 vdd.n678 0.152939
R21219 vdd.n682 vdd.n679 0.152939
R21220 vdd.n683 vdd.n682 0.152939
R21221 vdd.n684 vdd.n683 0.152939
R21222 vdd.n685 vdd.n684 0.152939
R21223 vdd.n690 vdd.n685 0.152939
R21224 vdd.n691 vdd.n690 0.152939
R21225 vdd.n692 vdd.n691 0.152939
R21226 vdd.n693 vdd.n692 0.152939
R21227 vdd.n696 vdd.n693 0.152939
R21228 vdd.n697 vdd.n696 0.152939
R21229 vdd.n698 vdd.n697 0.152939
R21230 vdd.n699 vdd.n698 0.152939
R21231 vdd.n702 vdd.n699 0.152939
R21232 vdd.n703 vdd.n702 0.152939
R21233 vdd.n704 vdd.n703 0.152939
R21234 vdd.n705 vdd.n704 0.152939
R21235 vdd.n708 vdd.n705 0.152939
R21236 vdd.n709 vdd.n708 0.152939
R21237 vdd.n710 vdd.n709 0.152939
R21238 vdd.n711 vdd.n710 0.152939
R21239 vdd.n714 vdd.n711 0.152939
R21240 vdd.n715 vdd.n714 0.152939
R21241 vdd.n716 vdd.n715 0.152939
R21242 vdd.n717 vdd.n716 0.152939
R21243 vdd.n720 vdd.n717 0.152939
R21244 vdd.n721 vdd.n720 0.152939
R21245 vdd.n3330 vdd.n721 0.152939
R21246 vdd.n3330 vdd.n3329 0.152939
R21247 vdd.n3329 vdd.n3328 0.152939
R21248 vdd.n3328 vdd.n725 0.152939
R21249 vdd.n730 vdd.n725 0.152939
R21250 vdd.n731 vdd.n730 0.152939
R21251 vdd.n734 vdd.n731 0.152939
R21252 vdd.n735 vdd.n734 0.152939
R21253 vdd.n736 vdd.n735 0.152939
R21254 vdd.n737 vdd.n736 0.152939
R21255 vdd.n740 vdd.n737 0.152939
R21256 vdd.n741 vdd.n740 0.152939
R21257 vdd.n742 vdd.n741 0.152939
R21258 vdd.n743 vdd.n742 0.152939
R21259 vdd.n746 vdd.n743 0.152939
R21260 vdd.n747 vdd.n746 0.152939
R21261 vdd.n748 vdd.n747 0.152939
R21262 vdd.n3413 vdd.n661 0.152939
R21263 vdd.n3414 vdd.n651 0.152939
R21264 vdd.n3428 vdd.n651 0.152939
R21265 vdd.n3429 vdd.n3428 0.152939
R21266 vdd.n3430 vdd.n3429 0.152939
R21267 vdd.n3430 vdd.n639 0.152939
R21268 vdd.n3444 vdd.n639 0.152939
R21269 vdd.n3445 vdd.n3444 0.152939
R21270 vdd.n3446 vdd.n3445 0.152939
R21271 vdd.n3446 vdd.n627 0.152939
R21272 vdd.n3461 vdd.n627 0.152939
R21273 vdd.n3462 vdd.n3461 0.152939
R21274 vdd.n3463 vdd.n3462 0.152939
R21275 vdd.n3463 vdd.n616 0.152939
R21276 vdd.n3480 vdd.n616 0.152939
R21277 vdd.n3481 vdd.n3480 0.152939
R21278 vdd.n3482 vdd.n3481 0.152939
R21279 vdd.n3482 vdd.n322 0.152939
R21280 vdd.n3562 vdd.n323 0.152939
R21281 vdd.n334 vdd.n323 0.152939
R21282 vdd.n335 vdd.n334 0.152939
R21283 vdd.n336 vdd.n335 0.152939
R21284 vdd.n343 vdd.n336 0.152939
R21285 vdd.n344 vdd.n343 0.152939
R21286 vdd.n345 vdd.n344 0.152939
R21287 vdd.n346 vdd.n345 0.152939
R21288 vdd.n354 vdd.n346 0.152939
R21289 vdd.n355 vdd.n354 0.152939
R21290 vdd.n356 vdd.n355 0.152939
R21291 vdd.n357 vdd.n356 0.152939
R21292 vdd.n365 vdd.n357 0.152939
R21293 vdd.n366 vdd.n365 0.152939
R21294 vdd.n367 vdd.n366 0.152939
R21295 vdd.n368 vdd.n367 0.152939
R21296 vdd.n443 vdd.n368 0.152939
R21297 vdd.n444 vdd.n442 0.152939
R21298 vdd.n451 vdd.n442 0.152939
R21299 vdd.n452 vdd.n451 0.152939
R21300 vdd.n453 vdd.n452 0.152939
R21301 vdd.n453 vdd.n440 0.152939
R21302 vdd.n461 vdd.n440 0.152939
R21303 vdd.n462 vdd.n461 0.152939
R21304 vdd.n463 vdd.n462 0.152939
R21305 vdd.n463 vdd.n438 0.152939
R21306 vdd.n471 vdd.n438 0.152939
R21307 vdd.n472 vdd.n471 0.152939
R21308 vdd.n473 vdd.n472 0.152939
R21309 vdd.n473 vdd.n436 0.152939
R21310 vdd.n481 vdd.n436 0.152939
R21311 vdd.n482 vdd.n481 0.152939
R21312 vdd.n483 vdd.n482 0.152939
R21313 vdd.n483 vdd.n434 0.152939
R21314 vdd.n491 vdd.n434 0.152939
R21315 vdd.n492 vdd.n491 0.152939
R21316 vdd.n493 vdd.n492 0.152939
R21317 vdd.n493 vdd.n430 0.152939
R21318 vdd.n501 vdd.n430 0.152939
R21319 vdd.n502 vdd.n501 0.152939
R21320 vdd.n503 vdd.n502 0.152939
R21321 vdd.n503 vdd.n428 0.152939
R21322 vdd.n511 vdd.n428 0.152939
R21323 vdd.n512 vdd.n511 0.152939
R21324 vdd.n513 vdd.n512 0.152939
R21325 vdd.n513 vdd.n426 0.152939
R21326 vdd.n521 vdd.n426 0.152939
R21327 vdd.n522 vdd.n521 0.152939
R21328 vdd.n523 vdd.n522 0.152939
R21329 vdd.n523 vdd.n424 0.152939
R21330 vdd.n531 vdd.n424 0.152939
R21331 vdd.n532 vdd.n531 0.152939
R21332 vdd.n533 vdd.n532 0.152939
R21333 vdd.n533 vdd.n422 0.152939
R21334 vdd.n541 vdd.n422 0.152939
R21335 vdd.n542 vdd.n541 0.152939
R21336 vdd.n543 vdd.n542 0.152939
R21337 vdd.n543 vdd.n418 0.152939
R21338 vdd.n551 vdd.n418 0.152939
R21339 vdd.n552 vdd.n551 0.152939
R21340 vdd.n553 vdd.n552 0.152939
R21341 vdd.n553 vdd.n416 0.152939
R21342 vdd.n561 vdd.n416 0.152939
R21343 vdd.n562 vdd.n561 0.152939
R21344 vdd.n563 vdd.n562 0.152939
R21345 vdd.n563 vdd.n414 0.152939
R21346 vdd.n571 vdd.n414 0.152939
R21347 vdd.n572 vdd.n571 0.152939
R21348 vdd.n573 vdd.n572 0.152939
R21349 vdd.n573 vdd.n412 0.152939
R21350 vdd.n581 vdd.n412 0.152939
R21351 vdd.n582 vdd.n581 0.152939
R21352 vdd.n583 vdd.n582 0.152939
R21353 vdd.n583 vdd.n410 0.152939
R21354 vdd.n591 vdd.n410 0.152939
R21355 vdd.n592 vdd.n591 0.152939
R21356 vdd.n593 vdd.n592 0.152939
R21357 vdd.n593 vdd.n408 0.152939
R21358 vdd.n600 vdd.n408 0.152939
R21359 vdd.n3521 vdd.n600 0.152939
R21360 vdd.n3421 vdd.n3420 0.152939
R21361 vdd.n3422 vdd.n3421 0.152939
R21362 vdd.n3422 vdd.n645 0.152939
R21363 vdd.n3436 vdd.n645 0.152939
R21364 vdd.n3437 vdd.n3436 0.152939
R21365 vdd.n3438 vdd.n3437 0.152939
R21366 vdd.n3438 vdd.n632 0.152939
R21367 vdd.n3452 vdd.n632 0.152939
R21368 vdd.n3453 vdd.n3452 0.152939
R21369 vdd.n3454 vdd.n3453 0.152939
R21370 vdd.n3454 vdd.n621 0.152939
R21371 vdd.n3469 vdd.n621 0.152939
R21372 vdd.n3470 vdd.n3469 0.152939
R21373 vdd.n3471 vdd.n3470 0.152939
R21374 vdd.n3473 vdd.n3471 0.152939
R21375 vdd.n3473 vdd.n3472 0.152939
R21376 vdd.n3472 vdd.n611 0.152939
R21377 vdd.n611 vdd.n609 0.152939
R21378 vdd.n3491 vdd.n609 0.152939
R21379 vdd.n3492 vdd.n3491 0.152939
R21380 vdd.n3493 vdd.n3492 0.152939
R21381 vdd.n3493 vdd.n607 0.152939
R21382 vdd.n3498 vdd.n607 0.152939
R21383 vdd.n3499 vdd.n3498 0.152939
R21384 vdd.n3500 vdd.n3499 0.152939
R21385 vdd.n3500 vdd.n605 0.152939
R21386 vdd.n3505 vdd.n605 0.152939
R21387 vdd.n3506 vdd.n3505 0.152939
R21388 vdd.n3507 vdd.n3506 0.152939
R21389 vdd.n3507 vdd.n603 0.152939
R21390 vdd.n3513 vdd.n603 0.152939
R21391 vdd.n3514 vdd.n3513 0.152939
R21392 vdd.n3515 vdd.n3514 0.152939
R21393 vdd.n3515 vdd.n601 0.152939
R21394 vdd.n3520 vdd.n601 0.152939
R21395 vdd.n3283 vdd.n656 0.152939
R21396 vdd.n2283 vdd.n1488 0.152939
R21397 vdd.n1834 vdd.n1833 0.152939
R21398 vdd.n1834 vdd.n1590 0.152939
R21399 vdd.n1848 vdd.n1590 0.152939
R21400 vdd.n1849 vdd.n1848 0.152939
R21401 vdd.n1850 vdd.n1849 0.152939
R21402 vdd.n1850 vdd.n1578 0.152939
R21403 vdd.n1865 vdd.n1578 0.152939
R21404 vdd.n1866 vdd.n1865 0.152939
R21405 vdd.n1867 vdd.n1866 0.152939
R21406 vdd.n1867 vdd.n1568 0.152939
R21407 vdd.n1882 vdd.n1568 0.152939
R21408 vdd.n1883 vdd.n1882 0.152939
R21409 vdd.n1884 vdd.n1883 0.152939
R21410 vdd.n1884 vdd.n1555 0.152939
R21411 vdd.n1898 vdd.n1555 0.152939
R21412 vdd.n1899 vdd.n1898 0.152939
R21413 vdd.n1900 vdd.n1899 0.152939
R21414 vdd.n1900 vdd.n1544 0.152939
R21415 vdd.n2210 vdd.n1544 0.152939
R21416 vdd.n2211 vdd.n2210 0.152939
R21417 vdd.n2212 vdd.n2211 0.152939
R21418 vdd.n2212 vdd.n1533 0.152939
R21419 vdd.n2226 vdd.n1533 0.152939
R21420 vdd.n2227 vdd.n2226 0.152939
R21421 vdd.n2228 vdd.n2227 0.152939
R21422 vdd.n2228 vdd.n1521 0.152939
R21423 vdd.n2243 vdd.n1521 0.152939
R21424 vdd.n2244 vdd.n2243 0.152939
R21425 vdd.n2245 vdd.n2244 0.152939
R21426 vdd.n2245 vdd.n1511 0.152939
R21427 vdd.n2260 vdd.n1511 0.152939
R21428 vdd.n2261 vdd.n2260 0.152939
R21429 vdd.n2264 vdd.n2261 0.152939
R21430 vdd.n2264 vdd.n2263 0.152939
R21431 vdd.n2263 vdd.n2262 0.152939
R21432 vdd.n1824 vdd.n1639 0.152939
R21433 vdd.n1824 vdd.n1823 0.152939
R21434 vdd.n1823 vdd.n1822 0.152939
R21435 vdd.n1822 vdd.n1641 0.152939
R21436 vdd.n1818 vdd.n1641 0.152939
R21437 vdd.n1818 vdd.n1817 0.152939
R21438 vdd.n1817 vdd.n1816 0.152939
R21439 vdd.n1816 vdd.n1646 0.152939
R21440 vdd.n1812 vdd.n1646 0.152939
R21441 vdd.n1812 vdd.n1811 0.152939
R21442 vdd.n1811 vdd.n1810 0.152939
R21443 vdd.n1810 vdd.n1652 0.152939
R21444 vdd.n1806 vdd.n1652 0.152939
R21445 vdd.n1806 vdd.n1805 0.152939
R21446 vdd.n1805 vdd.n1804 0.152939
R21447 vdd.n1804 vdd.n1658 0.152939
R21448 vdd.n1800 vdd.n1658 0.152939
R21449 vdd.n1800 vdd.n1799 0.152939
R21450 vdd.n1799 vdd.n1798 0.152939
R21451 vdd.n1798 vdd.n1664 0.152939
R21452 vdd.n1790 vdd.n1664 0.152939
R21453 vdd.n1790 vdd.n1789 0.152939
R21454 vdd.n1789 vdd.n1788 0.152939
R21455 vdd.n1788 vdd.n1668 0.152939
R21456 vdd.n1784 vdd.n1668 0.152939
R21457 vdd.n1784 vdd.n1783 0.152939
R21458 vdd.n1783 vdd.n1782 0.152939
R21459 vdd.n1782 vdd.n1674 0.152939
R21460 vdd.n1778 vdd.n1674 0.152939
R21461 vdd.n1778 vdd.n1777 0.152939
R21462 vdd.n1777 vdd.n1776 0.152939
R21463 vdd.n1776 vdd.n1680 0.152939
R21464 vdd.n1772 vdd.n1680 0.152939
R21465 vdd.n1772 vdd.n1771 0.152939
R21466 vdd.n1771 vdd.n1770 0.152939
R21467 vdd.n1770 vdd.n1686 0.152939
R21468 vdd.n1766 vdd.n1686 0.152939
R21469 vdd.n1766 vdd.n1765 0.152939
R21470 vdd.n1765 vdd.n1764 0.152939
R21471 vdd.n1764 vdd.n1692 0.152939
R21472 vdd.n1757 vdd.n1692 0.152939
R21473 vdd.n1757 vdd.n1756 0.152939
R21474 vdd.n1756 vdd.n1755 0.152939
R21475 vdd.n1755 vdd.n1697 0.152939
R21476 vdd.n1751 vdd.n1697 0.152939
R21477 vdd.n1751 vdd.n1750 0.152939
R21478 vdd.n1750 vdd.n1749 0.152939
R21479 vdd.n1749 vdd.n1703 0.152939
R21480 vdd.n1745 vdd.n1703 0.152939
R21481 vdd.n1745 vdd.n1744 0.152939
R21482 vdd.n1744 vdd.n1743 0.152939
R21483 vdd.n1743 vdd.n1709 0.152939
R21484 vdd.n1739 vdd.n1709 0.152939
R21485 vdd.n1739 vdd.n1738 0.152939
R21486 vdd.n1738 vdd.n1737 0.152939
R21487 vdd.n1737 vdd.n1715 0.152939
R21488 vdd.n1733 vdd.n1715 0.152939
R21489 vdd.n1733 vdd.n1732 0.152939
R21490 vdd.n1732 vdd.n1731 0.152939
R21491 vdd.n1731 vdd.n1721 0.152939
R21492 vdd.n1727 vdd.n1721 0.152939
R21493 vdd.n1727 vdd.n1602 0.152939
R21494 vdd.n1832 vdd.n1602 0.152939
R21495 vdd.n1840 vdd.n1596 0.152939
R21496 vdd.n1841 vdd.n1840 0.152939
R21497 vdd.n1842 vdd.n1841 0.152939
R21498 vdd.n1842 vdd.n1584 0.152939
R21499 vdd.n1857 vdd.n1584 0.152939
R21500 vdd.n1858 vdd.n1857 0.152939
R21501 vdd.n1859 vdd.n1858 0.152939
R21502 vdd.n1859 vdd.n1573 0.152939
R21503 vdd.n1874 vdd.n1573 0.152939
R21504 vdd.n1875 vdd.n1874 0.152939
R21505 vdd.n1876 vdd.n1875 0.152939
R21506 vdd.n1876 vdd.n1562 0.152939
R21507 vdd.n1890 vdd.n1562 0.152939
R21508 vdd.n1891 vdd.n1890 0.152939
R21509 vdd.n1892 vdd.n1891 0.152939
R21510 vdd.n1892 vdd.n1550 0.152939
R21511 vdd.n1907 vdd.n1550 0.152939
R21512 vdd.n2391 vdd.n2390 0.110256
R21513 vdd.n3214 vdd.n661 0.110256
R21514 vdd.n3283 vdd.n3282 0.110256
R21515 vdd.n2284 vdd.n2283 0.110256
R21516 vdd.n2203 vdd.n2202 0.0695946
R21517 vdd.n3563 vdd.n322 0.0695946
R21518 vdd.n3563 vdd.n3562 0.0695946
R21519 vdd.n2202 vdd.n1907 0.0695946
R21520 vdd.n2391 vdd.n1149 0.0431829
R21521 vdd.n2284 vdd.n1249 0.0431829
R21522 vdd.n3214 vdd.n667 0.0431829
R21523 vdd.n3282 vdd.n748 0.0431829
R21524 vdd vdd.n28 0.00833333
R21525 a_n2804_13878.n29 a_n2804_13878.n28 98.9632
R21526 a_n2804_13878.n2 a_n2804_13878.n0 98.7517
R21527 a_n2804_13878.n22 a_n2804_13878.n21 98.6055
R21528 a_n2804_13878.n24 a_n2804_13878.n23 98.6055
R21529 a_n2804_13878.n26 a_n2804_13878.n25 98.6055
R21530 a_n2804_13878.n28 a_n2804_13878.n27 98.6055
R21531 a_n2804_13878.n10 a_n2804_13878.n9 98.6055
R21532 a_n2804_13878.n8 a_n2804_13878.n7 98.6055
R21533 a_n2804_13878.n6 a_n2804_13878.n5 98.6055
R21534 a_n2804_13878.n4 a_n2804_13878.n3 98.6055
R21535 a_n2804_13878.n2 a_n2804_13878.n1 98.6055
R21536 a_n2804_13878.n20 a_n2804_13878.n19 98.6054
R21537 a_n2804_13878.n12 a_n2804_13878.t25 74.6477
R21538 a_n2804_13878.n17 a_n2804_13878.t26 74.2899
R21539 a_n2804_13878.n14 a_n2804_13878.t27 74.2899
R21540 a_n2804_13878.n13 a_n2804_13878.t24 74.2899
R21541 a_n2804_13878.n16 a_n2804_13878.n15 70.6783
R21542 a_n2804_13878.n12 a_n2804_13878.n11 70.6783
R21543 a_n2804_13878.n18 a_n2804_13878.n10 15.7159
R21544 a_n2804_13878.n20 a_n2804_13878.n18 12.6495
R21545 a_n2804_13878.n18 a_n2804_13878.n17 8.38735
R21546 a_n2804_13878.n19 a_n2804_13878.t7 3.61217
R21547 a_n2804_13878.n19 a_n2804_13878.t16 3.61217
R21548 a_n2804_13878.n21 a_n2804_13878.t20 3.61217
R21549 a_n2804_13878.n21 a_n2804_13878.t6 3.61217
R21550 a_n2804_13878.n23 a_n2804_13878.t10 3.61217
R21551 a_n2804_13878.n23 a_n2804_13878.t11 3.61217
R21552 a_n2804_13878.n25 a_n2804_13878.t21 3.61217
R21553 a_n2804_13878.n25 a_n2804_13878.t22 3.61217
R21554 a_n2804_13878.n27 a_n2804_13878.t0 3.61217
R21555 a_n2804_13878.n27 a_n2804_13878.t12 3.61217
R21556 a_n2804_13878.n15 a_n2804_13878.t30 3.61217
R21557 a_n2804_13878.n15 a_n2804_13878.t31 3.61217
R21558 a_n2804_13878.n11 a_n2804_13878.t28 3.61217
R21559 a_n2804_13878.n11 a_n2804_13878.t29 3.61217
R21560 a_n2804_13878.n9 a_n2804_13878.t13 3.61217
R21561 a_n2804_13878.n9 a_n2804_13878.t1 3.61217
R21562 a_n2804_13878.n7 a_n2804_13878.t18 3.61217
R21563 a_n2804_13878.n7 a_n2804_13878.t3 3.61217
R21564 a_n2804_13878.n5 a_n2804_13878.t2 3.61217
R21565 a_n2804_13878.n5 a_n2804_13878.t5 3.61217
R21566 a_n2804_13878.n3 a_n2804_13878.t15 3.61217
R21567 a_n2804_13878.n3 a_n2804_13878.t8 3.61217
R21568 a_n2804_13878.n1 a_n2804_13878.t19 3.61217
R21569 a_n2804_13878.n1 a_n2804_13878.t9 3.61217
R21570 a_n2804_13878.n0 a_n2804_13878.t4 3.61217
R21571 a_n2804_13878.n0 a_n2804_13878.t14 3.61217
R21572 a_n2804_13878.n29 a_n2804_13878.t17 3.61217
R21573 a_n2804_13878.t23 a_n2804_13878.n29 3.61217
R21574 a_n2804_13878.n13 a_n2804_13878.n12 0.358259
R21575 a_n2804_13878.n16 a_n2804_13878.n14 0.358259
R21576 a_n2804_13878.n17 a_n2804_13878.n16 0.358259
R21577 a_n2804_13878.n28 a_n2804_13878.n26 0.358259
R21578 a_n2804_13878.n26 a_n2804_13878.n24 0.358259
R21579 a_n2804_13878.n24 a_n2804_13878.n22 0.358259
R21580 a_n2804_13878.n22 a_n2804_13878.n20 0.358259
R21581 a_n2804_13878.n4 a_n2804_13878.n2 0.146627
R21582 a_n2804_13878.n6 a_n2804_13878.n4 0.146627
R21583 a_n2804_13878.n8 a_n2804_13878.n6 0.146627
R21584 a_n2804_13878.n10 a_n2804_13878.n8 0.146627
R21585 a_n2804_13878.n14 a_n2804_13878.n13 0.101793
R21586 CSoutput.n19 CSoutput.t164 184.661
R21587 CSoutput.n78 CSoutput.n77 165.8
R21588 CSoutput.n76 CSoutput.n0 165.8
R21589 CSoutput.n75 CSoutput.n74 165.8
R21590 CSoutput.n73 CSoutput.n72 165.8
R21591 CSoutput.n71 CSoutput.n2 165.8
R21592 CSoutput.n69 CSoutput.n68 165.8
R21593 CSoutput.n67 CSoutput.n3 165.8
R21594 CSoutput.n66 CSoutput.n65 165.8
R21595 CSoutput.n63 CSoutput.n4 165.8
R21596 CSoutput.n61 CSoutput.n60 165.8
R21597 CSoutput.n59 CSoutput.n5 165.8
R21598 CSoutput.n58 CSoutput.n57 165.8
R21599 CSoutput.n55 CSoutput.n6 165.8
R21600 CSoutput.n54 CSoutput.n53 165.8
R21601 CSoutput.n52 CSoutput.n51 165.8
R21602 CSoutput.n50 CSoutput.n8 165.8
R21603 CSoutput.n48 CSoutput.n47 165.8
R21604 CSoutput.n46 CSoutput.n9 165.8
R21605 CSoutput.n45 CSoutput.n44 165.8
R21606 CSoutput.n42 CSoutput.n10 165.8
R21607 CSoutput.n41 CSoutput.n40 165.8
R21608 CSoutput.n39 CSoutput.n38 165.8
R21609 CSoutput.n37 CSoutput.n12 165.8
R21610 CSoutput.n35 CSoutput.n34 165.8
R21611 CSoutput.n33 CSoutput.n13 165.8
R21612 CSoutput.n32 CSoutput.n31 165.8
R21613 CSoutput.n29 CSoutput.n14 165.8
R21614 CSoutput.n28 CSoutput.n27 165.8
R21615 CSoutput.n26 CSoutput.n25 165.8
R21616 CSoutput.n24 CSoutput.n16 165.8
R21617 CSoutput.n22 CSoutput.n21 165.8
R21618 CSoutput.n20 CSoutput.n17 165.8
R21619 CSoutput.n77 CSoutput.t165 162.194
R21620 CSoutput.n18 CSoutput.t166 120.501
R21621 CSoutput.n23 CSoutput.t174 120.501
R21622 CSoutput.n15 CSoutput.t170 120.501
R21623 CSoutput.n30 CSoutput.t167 120.501
R21624 CSoutput.n36 CSoutput.t177 120.501
R21625 CSoutput.n11 CSoutput.t180 120.501
R21626 CSoutput.n43 CSoutput.t169 120.501
R21627 CSoutput.n49 CSoutput.t181 120.501
R21628 CSoutput.n7 CSoutput.t160 120.501
R21629 CSoutput.n56 CSoutput.t176 120.501
R21630 CSoutput.n62 CSoutput.t168 120.501
R21631 CSoutput.n64 CSoutput.t162 120.501
R21632 CSoutput.n70 CSoutput.t179 120.501
R21633 CSoutput.n1 CSoutput.t173 120.501
R21634 CSoutput.n310 CSoutput.n308 103.469
R21635 CSoutput.n294 CSoutput.n292 103.469
R21636 CSoutput.n279 CSoutput.n277 103.469
R21637 CSoutput.n112 CSoutput.n110 103.469
R21638 CSoutput.n96 CSoutput.n94 103.469
R21639 CSoutput.n81 CSoutput.n79 103.469
R21640 CSoutput.n320 CSoutput.n319 103.111
R21641 CSoutput.n318 CSoutput.n317 103.111
R21642 CSoutput.n316 CSoutput.n315 103.111
R21643 CSoutput.n314 CSoutput.n313 103.111
R21644 CSoutput.n312 CSoutput.n311 103.111
R21645 CSoutput.n310 CSoutput.n309 103.111
R21646 CSoutput.n306 CSoutput.n305 103.111
R21647 CSoutput.n304 CSoutput.n303 103.111
R21648 CSoutput.n302 CSoutput.n301 103.111
R21649 CSoutput.n300 CSoutput.n299 103.111
R21650 CSoutput.n298 CSoutput.n297 103.111
R21651 CSoutput.n296 CSoutput.n295 103.111
R21652 CSoutput.n294 CSoutput.n293 103.111
R21653 CSoutput.n291 CSoutput.n290 103.111
R21654 CSoutput.n289 CSoutput.n288 103.111
R21655 CSoutput.n287 CSoutput.n286 103.111
R21656 CSoutput.n285 CSoutput.n284 103.111
R21657 CSoutput.n283 CSoutput.n282 103.111
R21658 CSoutput.n281 CSoutput.n280 103.111
R21659 CSoutput.n279 CSoutput.n278 103.111
R21660 CSoutput.n112 CSoutput.n111 103.111
R21661 CSoutput.n114 CSoutput.n113 103.111
R21662 CSoutput.n116 CSoutput.n115 103.111
R21663 CSoutput.n118 CSoutput.n117 103.111
R21664 CSoutput.n120 CSoutput.n119 103.111
R21665 CSoutput.n122 CSoutput.n121 103.111
R21666 CSoutput.n124 CSoutput.n123 103.111
R21667 CSoutput.n96 CSoutput.n95 103.111
R21668 CSoutput.n98 CSoutput.n97 103.111
R21669 CSoutput.n100 CSoutput.n99 103.111
R21670 CSoutput.n102 CSoutput.n101 103.111
R21671 CSoutput.n104 CSoutput.n103 103.111
R21672 CSoutput.n106 CSoutput.n105 103.111
R21673 CSoutput.n108 CSoutput.n107 103.111
R21674 CSoutput.n81 CSoutput.n80 103.111
R21675 CSoutput.n83 CSoutput.n82 103.111
R21676 CSoutput.n85 CSoutput.n84 103.111
R21677 CSoutput.n87 CSoutput.n86 103.111
R21678 CSoutput.n89 CSoutput.n88 103.111
R21679 CSoutput.n91 CSoutput.n90 103.111
R21680 CSoutput.n93 CSoutput.n92 103.111
R21681 CSoutput.n322 CSoutput.n321 103.111
R21682 CSoutput.n342 CSoutput.n340 81.5057
R21683 CSoutput.n327 CSoutput.n325 81.5057
R21684 CSoutput.n374 CSoutput.n372 81.5057
R21685 CSoutput.n359 CSoutput.n357 81.5057
R21686 CSoutput.n354 CSoutput.n353 80.9324
R21687 CSoutput.n352 CSoutput.n351 80.9324
R21688 CSoutput.n350 CSoutput.n349 80.9324
R21689 CSoutput.n348 CSoutput.n347 80.9324
R21690 CSoutput.n346 CSoutput.n345 80.9324
R21691 CSoutput.n344 CSoutput.n343 80.9324
R21692 CSoutput.n342 CSoutput.n341 80.9324
R21693 CSoutput.n339 CSoutput.n338 80.9324
R21694 CSoutput.n337 CSoutput.n336 80.9324
R21695 CSoutput.n335 CSoutput.n334 80.9324
R21696 CSoutput.n333 CSoutput.n332 80.9324
R21697 CSoutput.n331 CSoutput.n330 80.9324
R21698 CSoutput.n329 CSoutput.n328 80.9324
R21699 CSoutput.n327 CSoutput.n326 80.9324
R21700 CSoutput.n374 CSoutput.n373 80.9324
R21701 CSoutput.n376 CSoutput.n375 80.9324
R21702 CSoutput.n378 CSoutput.n377 80.9324
R21703 CSoutput.n380 CSoutput.n379 80.9324
R21704 CSoutput.n382 CSoutput.n381 80.9324
R21705 CSoutput.n384 CSoutput.n383 80.9324
R21706 CSoutput.n386 CSoutput.n385 80.9324
R21707 CSoutput.n359 CSoutput.n358 80.9324
R21708 CSoutput.n361 CSoutput.n360 80.9324
R21709 CSoutput.n363 CSoutput.n362 80.9324
R21710 CSoutput.n365 CSoutput.n364 80.9324
R21711 CSoutput.n367 CSoutput.n366 80.9324
R21712 CSoutput.n369 CSoutput.n368 80.9324
R21713 CSoutput.n371 CSoutput.n370 80.9324
R21714 CSoutput.n25 CSoutput.n24 48.1486
R21715 CSoutput.n69 CSoutput.n3 48.1486
R21716 CSoutput.n38 CSoutput.n37 48.1486
R21717 CSoutput.n42 CSoutput.n41 48.1486
R21718 CSoutput.n51 CSoutput.n50 48.1486
R21719 CSoutput.n55 CSoutput.n54 48.1486
R21720 CSoutput.n22 CSoutput.n17 46.462
R21721 CSoutput.n72 CSoutput.n71 46.462
R21722 CSoutput.n20 CSoutput.n19 44.9055
R21723 CSoutput.n29 CSoutput.n28 43.7635
R21724 CSoutput.n65 CSoutput.n63 43.7635
R21725 CSoutput.n35 CSoutput.n13 41.7396
R21726 CSoutput.n57 CSoutput.n5 41.7396
R21727 CSoutput.n44 CSoutput.n9 37.0171
R21728 CSoutput.n48 CSoutput.n9 37.0171
R21729 CSoutput.n76 CSoutput.n75 34.9932
R21730 CSoutput.n31 CSoutput.n13 32.2947
R21731 CSoutput.n61 CSoutput.n5 32.2947
R21732 CSoutput.n30 CSoutput.n29 29.6014
R21733 CSoutput.n63 CSoutput.n62 29.6014
R21734 CSoutput.n19 CSoutput.n18 28.4085
R21735 CSoutput.n18 CSoutput.n17 25.1176
R21736 CSoutput.n72 CSoutput.n1 25.1176
R21737 CSoutput.n43 CSoutput.n42 22.0922
R21738 CSoutput.n50 CSoutput.n49 22.0922
R21739 CSoutput.n77 CSoutput.n76 21.8586
R21740 CSoutput.n37 CSoutput.n36 18.9681
R21741 CSoutput.n56 CSoutput.n55 18.9681
R21742 CSoutput.n25 CSoutput.n15 17.6292
R21743 CSoutput.n64 CSoutput.n3 17.6292
R21744 CSoutput.n24 CSoutput.n23 15.844
R21745 CSoutput.n70 CSoutput.n69 15.844
R21746 CSoutput.n38 CSoutput.n11 14.5051
R21747 CSoutput.n54 CSoutput.n7 14.5051
R21748 CSoutput.n389 CSoutput.n78 11.6139
R21749 CSoutput.n41 CSoutput.n11 11.3811
R21750 CSoutput.n51 CSoutput.n7 11.3811
R21751 CSoutput.n23 CSoutput.n22 10.0422
R21752 CSoutput.n71 CSoutput.n70 10.0422
R21753 CSoutput.n307 CSoutput.n291 9.25285
R21754 CSoutput.n109 CSoutput.n93 9.25285
R21755 CSoutput.n355 CSoutput.n339 8.97993
R21756 CSoutput.n387 CSoutput.n371 8.97993
R21757 CSoutput.n356 CSoutput.n324 8.71993
R21758 CSoutput.n28 CSoutput.n15 8.25698
R21759 CSoutput.n65 CSoutput.n64 8.25698
R21760 CSoutput.n356 CSoutput.n355 7.89345
R21761 CSoutput.n388 CSoutput.n387 7.89345
R21762 CSoutput.n324 CSoutput.n323 7.12641
R21763 CSoutput.n126 CSoutput.n125 7.12641
R21764 CSoutput.n36 CSoutput.n35 6.91809
R21765 CSoutput.n57 CSoutput.n56 6.91809
R21766 CSoutput.n355 CSoutput.n354 5.25266
R21767 CSoutput.n387 CSoutput.n386 5.25266
R21768 CSoutput.n323 CSoutput.n322 5.1449
R21769 CSoutput.n307 CSoutput.n306 5.1449
R21770 CSoutput.n125 CSoutput.n124 5.1449
R21771 CSoutput.n109 CSoutput.n108 5.1449
R21772 CSoutput.n389 CSoutput.n126 5.12749
R21773 CSoutput.n217 CSoutput.n170 4.5005
R21774 CSoutput.n186 CSoutput.n170 4.5005
R21775 CSoutput.n181 CSoutput.n165 4.5005
R21776 CSoutput.n181 CSoutput.n167 4.5005
R21777 CSoutput.n181 CSoutput.n164 4.5005
R21778 CSoutput.n181 CSoutput.n168 4.5005
R21779 CSoutput.n181 CSoutput.n163 4.5005
R21780 CSoutput.n181 CSoutput.t175 4.5005
R21781 CSoutput.n181 CSoutput.n162 4.5005
R21782 CSoutput.n181 CSoutput.n169 4.5005
R21783 CSoutput.n181 CSoutput.n170 4.5005
R21784 CSoutput.n179 CSoutput.n165 4.5005
R21785 CSoutput.n179 CSoutput.n167 4.5005
R21786 CSoutput.n179 CSoutput.n164 4.5005
R21787 CSoutput.n179 CSoutput.n168 4.5005
R21788 CSoutput.n179 CSoutput.n163 4.5005
R21789 CSoutput.n179 CSoutput.t175 4.5005
R21790 CSoutput.n179 CSoutput.n162 4.5005
R21791 CSoutput.n179 CSoutput.n169 4.5005
R21792 CSoutput.n179 CSoutput.n170 4.5005
R21793 CSoutput.n178 CSoutput.n165 4.5005
R21794 CSoutput.n178 CSoutput.n167 4.5005
R21795 CSoutput.n178 CSoutput.n164 4.5005
R21796 CSoutput.n178 CSoutput.n168 4.5005
R21797 CSoutput.n178 CSoutput.n163 4.5005
R21798 CSoutput.n178 CSoutput.t175 4.5005
R21799 CSoutput.n178 CSoutput.n162 4.5005
R21800 CSoutput.n178 CSoutput.n169 4.5005
R21801 CSoutput.n178 CSoutput.n170 4.5005
R21802 CSoutput.n263 CSoutput.n165 4.5005
R21803 CSoutput.n263 CSoutput.n167 4.5005
R21804 CSoutput.n263 CSoutput.n164 4.5005
R21805 CSoutput.n263 CSoutput.n168 4.5005
R21806 CSoutput.n263 CSoutput.n163 4.5005
R21807 CSoutput.n263 CSoutput.t175 4.5005
R21808 CSoutput.n263 CSoutput.n162 4.5005
R21809 CSoutput.n263 CSoutput.n169 4.5005
R21810 CSoutput.n263 CSoutput.n170 4.5005
R21811 CSoutput.n261 CSoutput.n165 4.5005
R21812 CSoutput.n261 CSoutput.n167 4.5005
R21813 CSoutput.n261 CSoutput.n164 4.5005
R21814 CSoutput.n261 CSoutput.n168 4.5005
R21815 CSoutput.n261 CSoutput.n163 4.5005
R21816 CSoutput.n261 CSoutput.t175 4.5005
R21817 CSoutput.n261 CSoutput.n162 4.5005
R21818 CSoutput.n261 CSoutput.n169 4.5005
R21819 CSoutput.n259 CSoutput.n165 4.5005
R21820 CSoutput.n259 CSoutput.n167 4.5005
R21821 CSoutput.n259 CSoutput.n164 4.5005
R21822 CSoutput.n259 CSoutput.n168 4.5005
R21823 CSoutput.n259 CSoutput.n163 4.5005
R21824 CSoutput.n259 CSoutput.t175 4.5005
R21825 CSoutput.n259 CSoutput.n162 4.5005
R21826 CSoutput.n259 CSoutput.n169 4.5005
R21827 CSoutput.n189 CSoutput.n165 4.5005
R21828 CSoutput.n189 CSoutput.n167 4.5005
R21829 CSoutput.n189 CSoutput.n164 4.5005
R21830 CSoutput.n189 CSoutput.n168 4.5005
R21831 CSoutput.n189 CSoutput.n163 4.5005
R21832 CSoutput.n189 CSoutput.t175 4.5005
R21833 CSoutput.n189 CSoutput.n162 4.5005
R21834 CSoutput.n189 CSoutput.n169 4.5005
R21835 CSoutput.n189 CSoutput.n170 4.5005
R21836 CSoutput.n188 CSoutput.n165 4.5005
R21837 CSoutput.n188 CSoutput.n167 4.5005
R21838 CSoutput.n188 CSoutput.n164 4.5005
R21839 CSoutput.n188 CSoutput.n168 4.5005
R21840 CSoutput.n188 CSoutput.n163 4.5005
R21841 CSoutput.n188 CSoutput.t175 4.5005
R21842 CSoutput.n188 CSoutput.n162 4.5005
R21843 CSoutput.n188 CSoutput.n169 4.5005
R21844 CSoutput.n188 CSoutput.n170 4.5005
R21845 CSoutput.n192 CSoutput.n165 4.5005
R21846 CSoutput.n192 CSoutput.n167 4.5005
R21847 CSoutput.n192 CSoutput.n164 4.5005
R21848 CSoutput.n192 CSoutput.n168 4.5005
R21849 CSoutput.n192 CSoutput.n163 4.5005
R21850 CSoutput.n192 CSoutput.t175 4.5005
R21851 CSoutput.n192 CSoutput.n162 4.5005
R21852 CSoutput.n192 CSoutput.n169 4.5005
R21853 CSoutput.n192 CSoutput.n170 4.5005
R21854 CSoutput.n191 CSoutput.n165 4.5005
R21855 CSoutput.n191 CSoutput.n167 4.5005
R21856 CSoutput.n191 CSoutput.n164 4.5005
R21857 CSoutput.n191 CSoutput.n168 4.5005
R21858 CSoutput.n191 CSoutput.n163 4.5005
R21859 CSoutput.n191 CSoutput.t175 4.5005
R21860 CSoutput.n191 CSoutput.n162 4.5005
R21861 CSoutput.n191 CSoutput.n169 4.5005
R21862 CSoutput.n191 CSoutput.n170 4.5005
R21863 CSoutput.n174 CSoutput.n165 4.5005
R21864 CSoutput.n174 CSoutput.n167 4.5005
R21865 CSoutput.n174 CSoutput.n164 4.5005
R21866 CSoutput.n174 CSoutput.n168 4.5005
R21867 CSoutput.n174 CSoutput.n163 4.5005
R21868 CSoutput.n174 CSoutput.t175 4.5005
R21869 CSoutput.n174 CSoutput.n162 4.5005
R21870 CSoutput.n174 CSoutput.n169 4.5005
R21871 CSoutput.n174 CSoutput.n170 4.5005
R21872 CSoutput.n266 CSoutput.n165 4.5005
R21873 CSoutput.n266 CSoutput.n167 4.5005
R21874 CSoutput.n266 CSoutput.n164 4.5005
R21875 CSoutput.n266 CSoutput.n168 4.5005
R21876 CSoutput.n266 CSoutput.n163 4.5005
R21877 CSoutput.n266 CSoutput.t175 4.5005
R21878 CSoutput.n266 CSoutput.n162 4.5005
R21879 CSoutput.n266 CSoutput.n169 4.5005
R21880 CSoutput.n266 CSoutput.n170 4.5005
R21881 CSoutput.n253 CSoutput.n224 4.5005
R21882 CSoutput.n253 CSoutput.n230 4.5005
R21883 CSoutput.n211 CSoutput.n200 4.5005
R21884 CSoutput.n211 CSoutput.n202 4.5005
R21885 CSoutput.n211 CSoutput.n199 4.5005
R21886 CSoutput.n211 CSoutput.n203 4.5005
R21887 CSoutput.n211 CSoutput.n198 4.5005
R21888 CSoutput.n211 CSoutput.t171 4.5005
R21889 CSoutput.n211 CSoutput.n197 4.5005
R21890 CSoutput.n211 CSoutput.n204 4.5005
R21891 CSoutput.n253 CSoutput.n211 4.5005
R21892 CSoutput.n232 CSoutput.n200 4.5005
R21893 CSoutput.n232 CSoutput.n202 4.5005
R21894 CSoutput.n232 CSoutput.n199 4.5005
R21895 CSoutput.n232 CSoutput.n203 4.5005
R21896 CSoutput.n232 CSoutput.n198 4.5005
R21897 CSoutput.n232 CSoutput.t171 4.5005
R21898 CSoutput.n232 CSoutput.n197 4.5005
R21899 CSoutput.n232 CSoutput.n204 4.5005
R21900 CSoutput.n253 CSoutput.n232 4.5005
R21901 CSoutput.n210 CSoutput.n200 4.5005
R21902 CSoutput.n210 CSoutput.n202 4.5005
R21903 CSoutput.n210 CSoutput.n199 4.5005
R21904 CSoutput.n210 CSoutput.n203 4.5005
R21905 CSoutput.n210 CSoutput.n198 4.5005
R21906 CSoutput.n210 CSoutput.t171 4.5005
R21907 CSoutput.n210 CSoutput.n197 4.5005
R21908 CSoutput.n210 CSoutput.n204 4.5005
R21909 CSoutput.n253 CSoutput.n210 4.5005
R21910 CSoutput.n234 CSoutput.n200 4.5005
R21911 CSoutput.n234 CSoutput.n202 4.5005
R21912 CSoutput.n234 CSoutput.n199 4.5005
R21913 CSoutput.n234 CSoutput.n203 4.5005
R21914 CSoutput.n234 CSoutput.n198 4.5005
R21915 CSoutput.n234 CSoutput.t171 4.5005
R21916 CSoutput.n234 CSoutput.n197 4.5005
R21917 CSoutput.n234 CSoutput.n204 4.5005
R21918 CSoutput.n253 CSoutput.n234 4.5005
R21919 CSoutput.n200 CSoutput.n195 4.5005
R21920 CSoutput.n202 CSoutput.n195 4.5005
R21921 CSoutput.n199 CSoutput.n195 4.5005
R21922 CSoutput.n203 CSoutput.n195 4.5005
R21923 CSoutput.n198 CSoutput.n195 4.5005
R21924 CSoutput.t171 CSoutput.n195 4.5005
R21925 CSoutput.n197 CSoutput.n195 4.5005
R21926 CSoutput.n204 CSoutput.n195 4.5005
R21927 CSoutput.n256 CSoutput.n200 4.5005
R21928 CSoutput.n256 CSoutput.n202 4.5005
R21929 CSoutput.n256 CSoutput.n199 4.5005
R21930 CSoutput.n256 CSoutput.n203 4.5005
R21931 CSoutput.n256 CSoutput.n198 4.5005
R21932 CSoutput.n256 CSoutput.t171 4.5005
R21933 CSoutput.n256 CSoutput.n197 4.5005
R21934 CSoutput.n256 CSoutput.n204 4.5005
R21935 CSoutput.n254 CSoutput.n200 4.5005
R21936 CSoutput.n254 CSoutput.n202 4.5005
R21937 CSoutput.n254 CSoutput.n199 4.5005
R21938 CSoutput.n254 CSoutput.n203 4.5005
R21939 CSoutput.n254 CSoutput.n198 4.5005
R21940 CSoutput.n254 CSoutput.t171 4.5005
R21941 CSoutput.n254 CSoutput.n197 4.5005
R21942 CSoutput.n254 CSoutput.n204 4.5005
R21943 CSoutput.n254 CSoutput.n253 4.5005
R21944 CSoutput.n236 CSoutput.n200 4.5005
R21945 CSoutput.n236 CSoutput.n202 4.5005
R21946 CSoutput.n236 CSoutput.n199 4.5005
R21947 CSoutput.n236 CSoutput.n203 4.5005
R21948 CSoutput.n236 CSoutput.n198 4.5005
R21949 CSoutput.n236 CSoutput.t171 4.5005
R21950 CSoutput.n236 CSoutput.n197 4.5005
R21951 CSoutput.n236 CSoutput.n204 4.5005
R21952 CSoutput.n253 CSoutput.n236 4.5005
R21953 CSoutput.n208 CSoutput.n200 4.5005
R21954 CSoutput.n208 CSoutput.n202 4.5005
R21955 CSoutput.n208 CSoutput.n199 4.5005
R21956 CSoutput.n208 CSoutput.n203 4.5005
R21957 CSoutput.n208 CSoutput.n198 4.5005
R21958 CSoutput.n208 CSoutput.t171 4.5005
R21959 CSoutput.n208 CSoutput.n197 4.5005
R21960 CSoutput.n208 CSoutput.n204 4.5005
R21961 CSoutput.n253 CSoutput.n208 4.5005
R21962 CSoutput.n238 CSoutput.n200 4.5005
R21963 CSoutput.n238 CSoutput.n202 4.5005
R21964 CSoutput.n238 CSoutput.n199 4.5005
R21965 CSoutput.n238 CSoutput.n203 4.5005
R21966 CSoutput.n238 CSoutput.n198 4.5005
R21967 CSoutput.n238 CSoutput.t171 4.5005
R21968 CSoutput.n238 CSoutput.n197 4.5005
R21969 CSoutput.n238 CSoutput.n204 4.5005
R21970 CSoutput.n253 CSoutput.n238 4.5005
R21971 CSoutput.n207 CSoutput.n200 4.5005
R21972 CSoutput.n207 CSoutput.n202 4.5005
R21973 CSoutput.n207 CSoutput.n199 4.5005
R21974 CSoutput.n207 CSoutput.n203 4.5005
R21975 CSoutput.n207 CSoutput.n198 4.5005
R21976 CSoutput.n207 CSoutput.t171 4.5005
R21977 CSoutput.n207 CSoutput.n197 4.5005
R21978 CSoutput.n207 CSoutput.n204 4.5005
R21979 CSoutput.n253 CSoutput.n207 4.5005
R21980 CSoutput.n252 CSoutput.n200 4.5005
R21981 CSoutput.n252 CSoutput.n202 4.5005
R21982 CSoutput.n252 CSoutput.n199 4.5005
R21983 CSoutput.n252 CSoutput.n203 4.5005
R21984 CSoutput.n252 CSoutput.n198 4.5005
R21985 CSoutput.n252 CSoutput.t171 4.5005
R21986 CSoutput.n252 CSoutput.n197 4.5005
R21987 CSoutput.n252 CSoutput.n204 4.5005
R21988 CSoutput.n253 CSoutput.n252 4.5005
R21989 CSoutput.n251 CSoutput.n136 4.5005
R21990 CSoutput.n152 CSoutput.n136 4.5005
R21991 CSoutput.n147 CSoutput.n131 4.5005
R21992 CSoutput.n147 CSoutput.n133 4.5005
R21993 CSoutput.n147 CSoutput.n130 4.5005
R21994 CSoutput.n147 CSoutput.n134 4.5005
R21995 CSoutput.n147 CSoutput.n129 4.5005
R21996 CSoutput.n147 CSoutput.t161 4.5005
R21997 CSoutput.n147 CSoutput.n128 4.5005
R21998 CSoutput.n147 CSoutput.n135 4.5005
R21999 CSoutput.n147 CSoutput.n136 4.5005
R22000 CSoutput.n145 CSoutput.n131 4.5005
R22001 CSoutput.n145 CSoutput.n133 4.5005
R22002 CSoutput.n145 CSoutput.n130 4.5005
R22003 CSoutput.n145 CSoutput.n134 4.5005
R22004 CSoutput.n145 CSoutput.n129 4.5005
R22005 CSoutput.n145 CSoutput.t161 4.5005
R22006 CSoutput.n145 CSoutput.n128 4.5005
R22007 CSoutput.n145 CSoutput.n135 4.5005
R22008 CSoutput.n145 CSoutput.n136 4.5005
R22009 CSoutput.n144 CSoutput.n131 4.5005
R22010 CSoutput.n144 CSoutput.n133 4.5005
R22011 CSoutput.n144 CSoutput.n130 4.5005
R22012 CSoutput.n144 CSoutput.n134 4.5005
R22013 CSoutput.n144 CSoutput.n129 4.5005
R22014 CSoutput.n144 CSoutput.t161 4.5005
R22015 CSoutput.n144 CSoutput.n128 4.5005
R22016 CSoutput.n144 CSoutput.n135 4.5005
R22017 CSoutput.n144 CSoutput.n136 4.5005
R22018 CSoutput.n273 CSoutput.n131 4.5005
R22019 CSoutput.n273 CSoutput.n133 4.5005
R22020 CSoutput.n273 CSoutput.n130 4.5005
R22021 CSoutput.n273 CSoutput.n134 4.5005
R22022 CSoutput.n273 CSoutput.n129 4.5005
R22023 CSoutput.n273 CSoutput.t161 4.5005
R22024 CSoutput.n273 CSoutput.n128 4.5005
R22025 CSoutput.n273 CSoutput.n135 4.5005
R22026 CSoutput.n273 CSoutput.n136 4.5005
R22027 CSoutput.n271 CSoutput.n131 4.5005
R22028 CSoutput.n271 CSoutput.n133 4.5005
R22029 CSoutput.n271 CSoutput.n130 4.5005
R22030 CSoutput.n271 CSoutput.n134 4.5005
R22031 CSoutput.n271 CSoutput.n129 4.5005
R22032 CSoutput.n271 CSoutput.t161 4.5005
R22033 CSoutput.n271 CSoutput.n128 4.5005
R22034 CSoutput.n271 CSoutput.n135 4.5005
R22035 CSoutput.n269 CSoutput.n131 4.5005
R22036 CSoutput.n269 CSoutput.n133 4.5005
R22037 CSoutput.n269 CSoutput.n130 4.5005
R22038 CSoutput.n269 CSoutput.n134 4.5005
R22039 CSoutput.n269 CSoutput.n129 4.5005
R22040 CSoutput.n269 CSoutput.t161 4.5005
R22041 CSoutput.n269 CSoutput.n128 4.5005
R22042 CSoutput.n269 CSoutput.n135 4.5005
R22043 CSoutput.n155 CSoutput.n131 4.5005
R22044 CSoutput.n155 CSoutput.n133 4.5005
R22045 CSoutput.n155 CSoutput.n130 4.5005
R22046 CSoutput.n155 CSoutput.n134 4.5005
R22047 CSoutput.n155 CSoutput.n129 4.5005
R22048 CSoutput.n155 CSoutput.t161 4.5005
R22049 CSoutput.n155 CSoutput.n128 4.5005
R22050 CSoutput.n155 CSoutput.n135 4.5005
R22051 CSoutput.n155 CSoutput.n136 4.5005
R22052 CSoutput.n154 CSoutput.n131 4.5005
R22053 CSoutput.n154 CSoutput.n133 4.5005
R22054 CSoutput.n154 CSoutput.n130 4.5005
R22055 CSoutput.n154 CSoutput.n134 4.5005
R22056 CSoutput.n154 CSoutput.n129 4.5005
R22057 CSoutput.n154 CSoutput.t161 4.5005
R22058 CSoutput.n154 CSoutput.n128 4.5005
R22059 CSoutput.n154 CSoutput.n135 4.5005
R22060 CSoutput.n154 CSoutput.n136 4.5005
R22061 CSoutput.n158 CSoutput.n131 4.5005
R22062 CSoutput.n158 CSoutput.n133 4.5005
R22063 CSoutput.n158 CSoutput.n130 4.5005
R22064 CSoutput.n158 CSoutput.n134 4.5005
R22065 CSoutput.n158 CSoutput.n129 4.5005
R22066 CSoutput.n158 CSoutput.t161 4.5005
R22067 CSoutput.n158 CSoutput.n128 4.5005
R22068 CSoutput.n158 CSoutput.n135 4.5005
R22069 CSoutput.n158 CSoutput.n136 4.5005
R22070 CSoutput.n157 CSoutput.n131 4.5005
R22071 CSoutput.n157 CSoutput.n133 4.5005
R22072 CSoutput.n157 CSoutput.n130 4.5005
R22073 CSoutput.n157 CSoutput.n134 4.5005
R22074 CSoutput.n157 CSoutput.n129 4.5005
R22075 CSoutput.n157 CSoutput.t161 4.5005
R22076 CSoutput.n157 CSoutput.n128 4.5005
R22077 CSoutput.n157 CSoutput.n135 4.5005
R22078 CSoutput.n157 CSoutput.n136 4.5005
R22079 CSoutput.n140 CSoutput.n131 4.5005
R22080 CSoutput.n140 CSoutput.n133 4.5005
R22081 CSoutput.n140 CSoutput.n130 4.5005
R22082 CSoutput.n140 CSoutput.n134 4.5005
R22083 CSoutput.n140 CSoutput.n129 4.5005
R22084 CSoutput.n140 CSoutput.t161 4.5005
R22085 CSoutput.n140 CSoutput.n128 4.5005
R22086 CSoutput.n140 CSoutput.n135 4.5005
R22087 CSoutput.n140 CSoutput.n136 4.5005
R22088 CSoutput.n276 CSoutput.n131 4.5005
R22089 CSoutput.n276 CSoutput.n133 4.5005
R22090 CSoutput.n276 CSoutput.n130 4.5005
R22091 CSoutput.n276 CSoutput.n134 4.5005
R22092 CSoutput.n276 CSoutput.n129 4.5005
R22093 CSoutput.n276 CSoutput.t161 4.5005
R22094 CSoutput.n276 CSoutput.n128 4.5005
R22095 CSoutput.n276 CSoutput.n135 4.5005
R22096 CSoutput.n276 CSoutput.n136 4.5005
R22097 CSoutput.n323 CSoutput.n307 4.10845
R22098 CSoutput.n125 CSoutput.n109 4.10845
R22099 CSoutput.n321 CSoutput.t99 4.06363
R22100 CSoutput.n321 CSoutput.t29 4.06363
R22101 CSoutput.n319 CSoutput.t45 4.06363
R22102 CSoutput.n319 CSoutput.t69 4.06363
R22103 CSoutput.n317 CSoutput.t81 4.06363
R22104 CSoutput.n317 CSoutput.t16 4.06363
R22105 CSoutput.n315 CSoutput.t12 4.06363
R22106 CSoutput.n315 CSoutput.t47 4.06363
R22107 CSoutput.n313 CSoutput.t63 4.06363
R22108 CSoutput.n313 CSoutput.t83 4.06363
R22109 CSoutput.n311 CSoutput.t96 4.06363
R22110 CSoutput.n311 CSoutput.t26 4.06363
R22111 CSoutput.n309 CSoutput.t32 4.06363
R22112 CSoutput.n309 CSoutput.t84 4.06363
R22113 CSoutput.n308 CSoutput.t98 4.06363
R22114 CSoutput.n308 CSoutput.t100 4.06363
R22115 CSoutput.n305 CSoutput.t90 4.06363
R22116 CSoutput.n305 CSoutput.t17 4.06363
R22117 CSoutput.n303 CSoutput.t33 4.06363
R22118 CSoutput.n303 CSoutput.t61 4.06363
R22119 CSoutput.n301 CSoutput.t74 4.06363
R22120 CSoutput.n301 CSoutput.t104 4.06363
R22121 CSoutput.n299 CSoutput.t97 4.06363
R22122 CSoutput.n299 CSoutput.t38 4.06363
R22123 CSoutput.n297 CSoutput.t51 4.06363
R22124 CSoutput.n297 CSoutput.t75 4.06363
R22125 CSoutput.n295 CSoutput.t85 4.06363
R22126 CSoutput.n295 CSoutput.t15 4.06363
R22127 CSoutput.n293 CSoutput.t18 4.06363
R22128 CSoutput.n293 CSoutput.t78 4.06363
R22129 CSoutput.n292 CSoutput.t91 4.06363
R22130 CSoutput.n292 CSoutput.t92 4.06363
R22131 CSoutput.n290 CSoutput.t101 4.06363
R22132 CSoutput.n290 CSoutput.t62 4.06363
R22133 CSoutput.n288 CSoutput.t88 4.06363
R22134 CSoutput.n288 CSoutput.t48 4.06363
R22135 CSoutput.n286 CSoutput.t76 4.06363
R22136 CSoutput.n286 CSoutput.t36 4.06363
R22137 CSoutput.n284 CSoutput.t94 4.06363
R22138 CSoutput.n284 CSoutput.t55 4.06363
R22139 CSoutput.n282 CSoutput.t82 4.06363
R22140 CSoutput.n282 CSoutput.t43 4.06363
R22141 CSoutput.n280 CSoutput.t71 4.06363
R22142 CSoutput.n280 CSoutput.t25 4.06363
R22143 CSoutput.n278 CSoutput.t86 4.06363
R22144 CSoutput.n278 CSoutput.t20 4.06363
R22145 CSoutput.n277 CSoutput.t52 4.06363
R22146 CSoutput.n277 CSoutput.t34 4.06363
R22147 CSoutput.n110 CSoutput.t66 4.06363
R22148 CSoutput.n110 CSoutput.t41 4.06363
R22149 CSoutput.n111 CSoutput.t24 4.06363
R22150 CSoutput.n111 CSoutput.t68 4.06363
R22151 CSoutput.n113 CSoutput.t65 4.06363
R22152 CSoutput.n113 CSoutput.t39 4.06363
R22153 CSoutput.n115 CSoutput.t23 4.06363
R22154 CSoutput.n115 CSoutput.t22 4.06363
R22155 CSoutput.n117 CSoutput.t80 4.06363
R22156 CSoutput.n117 CSoutput.t50 4.06363
R22157 CSoutput.n119 CSoutput.t46 4.06363
R22158 CSoutput.n119 CSoutput.t19 4.06363
R22159 CSoutput.n121 CSoutput.t103 4.06363
R22160 CSoutput.n121 CSoutput.t79 4.06363
R22161 CSoutput.n123 CSoutput.t67 4.06363
R22162 CSoutput.n123 CSoutput.t42 4.06363
R22163 CSoutput.n94 CSoutput.t57 4.06363
R22164 CSoutput.n94 CSoutput.t30 4.06363
R22165 CSoutput.n95 CSoutput.t14 4.06363
R22166 CSoutput.n95 CSoutput.t59 4.06363
R22167 CSoutput.n97 CSoutput.t54 4.06363
R22168 CSoutput.n97 CSoutput.t27 4.06363
R22169 CSoutput.n99 CSoutput.t13 4.06363
R22170 CSoutput.n99 CSoutput.t11 4.06363
R22171 CSoutput.n101 CSoutput.t73 4.06363
R22172 CSoutput.n101 CSoutput.t40 4.06363
R22173 CSoutput.n103 CSoutput.t37 4.06363
R22174 CSoutput.n103 CSoutput.t10 4.06363
R22175 CSoutput.n105 CSoutput.t93 4.06363
R22176 CSoutput.n105 CSoutput.t70 4.06363
R22177 CSoutput.n107 CSoutput.t58 4.06363
R22178 CSoutput.n107 CSoutput.t31 4.06363
R22179 CSoutput.n79 CSoutput.t105 4.06363
R22180 CSoutput.n79 CSoutput.t53 4.06363
R22181 CSoutput.n80 CSoutput.t21 4.06363
R22182 CSoutput.n80 CSoutput.t87 4.06363
R22183 CSoutput.n82 CSoutput.t28 4.06363
R22184 CSoutput.n82 CSoutput.t72 4.06363
R22185 CSoutput.n84 CSoutput.t44 4.06363
R22186 CSoutput.n84 CSoutput.t60 4.06363
R22187 CSoutput.n86 CSoutput.t56 4.06363
R22188 CSoutput.n86 CSoutput.t95 4.06363
R22189 CSoutput.n88 CSoutput.t35 4.06363
R22190 CSoutput.n88 CSoutput.t77 4.06363
R22191 CSoutput.n90 CSoutput.t49 4.06363
R22192 CSoutput.n90 CSoutput.t89 4.06363
R22193 CSoutput.n92 CSoutput.t64 4.06363
R22194 CSoutput.n92 CSoutput.t102 4.06363
R22195 CSoutput.n44 CSoutput.n43 3.79402
R22196 CSoutput.n49 CSoutput.n48 3.79402
R22197 CSoutput.n389 CSoutput.n388 3.57343
R22198 CSoutput.n388 CSoutput.n356 3.3798
R22199 CSoutput.n324 CSoutput.n126 2.99158
R22200 CSoutput.n353 CSoutput.t157 2.82907
R22201 CSoutput.n353 CSoutput.t128 2.82907
R22202 CSoutput.n351 CSoutput.t127 2.82907
R22203 CSoutput.n351 CSoutput.t142 2.82907
R22204 CSoutput.n349 CSoutput.t1 2.82907
R22205 CSoutput.n349 CSoutput.t7 2.82907
R22206 CSoutput.n347 CSoutput.t8 2.82907
R22207 CSoutput.n347 CSoutput.t147 2.82907
R22208 CSoutput.n345 CSoutput.t129 2.82907
R22209 CSoutput.n345 CSoutput.t117 2.82907
R22210 CSoutput.n343 CSoutput.t0 2.82907
R22211 CSoutput.n343 CSoutput.t158 2.82907
R22212 CSoutput.n341 CSoutput.t137 2.82907
R22213 CSoutput.n341 CSoutput.t153 2.82907
R22214 CSoutput.n340 CSoutput.t148 2.82907
R22215 CSoutput.n340 CSoutput.t154 2.82907
R22216 CSoutput.n338 CSoutput.t156 2.82907
R22217 CSoutput.n338 CSoutput.t4 2.82907
R22218 CSoutput.n336 CSoutput.t107 2.82907
R22219 CSoutput.n336 CSoutput.t146 2.82907
R22220 CSoutput.n334 CSoutput.t108 2.82907
R22221 CSoutput.n334 CSoutput.t106 2.82907
R22222 CSoutput.n332 CSoutput.t114 2.82907
R22223 CSoutput.n332 CSoutput.t111 2.82907
R22224 CSoutput.n330 CSoutput.t119 2.82907
R22225 CSoutput.n330 CSoutput.t149 2.82907
R22226 CSoutput.n328 CSoutput.t155 2.82907
R22227 CSoutput.n328 CSoutput.t132 2.82907
R22228 CSoutput.n326 CSoutput.t145 2.82907
R22229 CSoutput.n326 CSoutput.t115 2.82907
R22230 CSoutput.n325 CSoutput.t118 2.82907
R22231 CSoutput.n325 CSoutput.t136 2.82907
R22232 CSoutput.n372 CSoutput.t112 2.82907
R22233 CSoutput.n372 CSoutput.t141 2.82907
R22234 CSoutput.n373 CSoutput.t9 2.82907
R22235 CSoutput.n373 CSoutput.t121 2.82907
R22236 CSoutput.n375 CSoutput.t123 2.82907
R22237 CSoutput.n375 CSoutput.t125 2.82907
R22238 CSoutput.n377 CSoutput.t140 2.82907
R22239 CSoutput.n377 CSoutput.t131 2.82907
R22240 CSoutput.n379 CSoutput.t110 2.82907
R22241 CSoutput.n379 CSoutput.t113 2.82907
R22242 CSoutput.n381 CSoutput.t126 2.82907
R22243 CSoutput.n381 CSoutput.t122 2.82907
R22244 CSoutput.n383 CSoutput.t133 2.82907
R22245 CSoutput.n383 CSoutput.t151 2.82907
R22246 CSoutput.n385 CSoutput.t5 2.82907
R22247 CSoutput.n385 CSoutput.t135 2.82907
R22248 CSoutput.n357 CSoutput.t143 2.82907
R22249 CSoutput.n357 CSoutput.t124 2.82907
R22250 CSoutput.n358 CSoutput.t138 2.82907
R22251 CSoutput.n358 CSoutput.t120 2.82907
R22252 CSoutput.n360 CSoutput.t130 2.82907
R22253 CSoutput.n360 CSoutput.t152 2.82907
R22254 CSoutput.n362 CSoutput.t3 2.82907
R22255 CSoutput.n362 CSoutput.t134 2.82907
R22256 CSoutput.n364 CSoutput.t159 2.82907
R22257 CSoutput.n364 CSoutput.t144 2.82907
R22258 CSoutput.n366 CSoutput.t6 2.82907
R22259 CSoutput.n366 CSoutput.t150 2.82907
R22260 CSoutput.n368 CSoutput.t109 2.82907
R22261 CSoutput.n368 CSoutput.t2 2.82907
R22262 CSoutput.n370 CSoutput.t139 2.82907
R22263 CSoutput.n370 CSoutput.t116 2.82907
R22264 CSoutput.n75 CSoutput.n1 2.45513
R22265 CSoutput.n217 CSoutput.n215 2.251
R22266 CSoutput.n217 CSoutput.n214 2.251
R22267 CSoutput.n217 CSoutput.n213 2.251
R22268 CSoutput.n217 CSoutput.n212 2.251
R22269 CSoutput.n186 CSoutput.n185 2.251
R22270 CSoutput.n186 CSoutput.n184 2.251
R22271 CSoutput.n186 CSoutput.n183 2.251
R22272 CSoutput.n186 CSoutput.n182 2.251
R22273 CSoutput.n259 CSoutput.n258 2.251
R22274 CSoutput.n224 CSoutput.n222 2.251
R22275 CSoutput.n224 CSoutput.n221 2.251
R22276 CSoutput.n224 CSoutput.n220 2.251
R22277 CSoutput.n242 CSoutput.n224 2.251
R22278 CSoutput.n230 CSoutput.n229 2.251
R22279 CSoutput.n230 CSoutput.n228 2.251
R22280 CSoutput.n230 CSoutput.n227 2.251
R22281 CSoutput.n230 CSoutput.n226 2.251
R22282 CSoutput.n256 CSoutput.n196 2.251
R22283 CSoutput.n251 CSoutput.n249 2.251
R22284 CSoutput.n251 CSoutput.n248 2.251
R22285 CSoutput.n251 CSoutput.n247 2.251
R22286 CSoutput.n251 CSoutput.n246 2.251
R22287 CSoutput.n152 CSoutput.n151 2.251
R22288 CSoutput.n152 CSoutput.n150 2.251
R22289 CSoutput.n152 CSoutput.n149 2.251
R22290 CSoutput.n152 CSoutput.n148 2.251
R22291 CSoutput.n269 CSoutput.n268 2.251
R22292 CSoutput.n186 CSoutput.n166 2.2505
R22293 CSoutput.n181 CSoutput.n166 2.2505
R22294 CSoutput.n179 CSoutput.n166 2.2505
R22295 CSoutput.n178 CSoutput.n166 2.2505
R22296 CSoutput.n263 CSoutput.n166 2.2505
R22297 CSoutput.n261 CSoutput.n166 2.2505
R22298 CSoutput.n259 CSoutput.n166 2.2505
R22299 CSoutput.n189 CSoutput.n166 2.2505
R22300 CSoutput.n188 CSoutput.n166 2.2505
R22301 CSoutput.n192 CSoutput.n166 2.2505
R22302 CSoutput.n191 CSoutput.n166 2.2505
R22303 CSoutput.n174 CSoutput.n166 2.2505
R22304 CSoutput.n266 CSoutput.n166 2.2505
R22305 CSoutput.n266 CSoutput.n265 2.2505
R22306 CSoutput.n230 CSoutput.n201 2.2505
R22307 CSoutput.n211 CSoutput.n201 2.2505
R22308 CSoutput.n232 CSoutput.n201 2.2505
R22309 CSoutput.n210 CSoutput.n201 2.2505
R22310 CSoutput.n234 CSoutput.n201 2.2505
R22311 CSoutput.n201 CSoutput.n195 2.2505
R22312 CSoutput.n256 CSoutput.n201 2.2505
R22313 CSoutput.n254 CSoutput.n201 2.2505
R22314 CSoutput.n236 CSoutput.n201 2.2505
R22315 CSoutput.n208 CSoutput.n201 2.2505
R22316 CSoutput.n238 CSoutput.n201 2.2505
R22317 CSoutput.n207 CSoutput.n201 2.2505
R22318 CSoutput.n252 CSoutput.n201 2.2505
R22319 CSoutput.n252 CSoutput.n205 2.2505
R22320 CSoutput.n152 CSoutput.n132 2.2505
R22321 CSoutput.n147 CSoutput.n132 2.2505
R22322 CSoutput.n145 CSoutput.n132 2.2505
R22323 CSoutput.n144 CSoutput.n132 2.2505
R22324 CSoutput.n273 CSoutput.n132 2.2505
R22325 CSoutput.n271 CSoutput.n132 2.2505
R22326 CSoutput.n269 CSoutput.n132 2.2505
R22327 CSoutput.n155 CSoutput.n132 2.2505
R22328 CSoutput.n154 CSoutput.n132 2.2505
R22329 CSoutput.n158 CSoutput.n132 2.2505
R22330 CSoutput.n157 CSoutput.n132 2.2505
R22331 CSoutput.n140 CSoutput.n132 2.2505
R22332 CSoutput.n276 CSoutput.n132 2.2505
R22333 CSoutput.n276 CSoutput.n275 2.2505
R22334 CSoutput.n194 CSoutput.n187 2.25024
R22335 CSoutput.n194 CSoutput.n180 2.25024
R22336 CSoutput.n262 CSoutput.n194 2.25024
R22337 CSoutput.n194 CSoutput.n190 2.25024
R22338 CSoutput.n194 CSoutput.n193 2.25024
R22339 CSoutput.n194 CSoutput.n161 2.25024
R22340 CSoutput.n244 CSoutput.n241 2.25024
R22341 CSoutput.n244 CSoutput.n240 2.25024
R22342 CSoutput.n244 CSoutput.n239 2.25024
R22343 CSoutput.n244 CSoutput.n206 2.25024
R22344 CSoutput.n244 CSoutput.n243 2.25024
R22345 CSoutput.n245 CSoutput.n244 2.25024
R22346 CSoutput.n160 CSoutput.n153 2.25024
R22347 CSoutput.n160 CSoutput.n146 2.25024
R22348 CSoutput.n272 CSoutput.n160 2.25024
R22349 CSoutput.n160 CSoutput.n156 2.25024
R22350 CSoutput.n160 CSoutput.n159 2.25024
R22351 CSoutput.n160 CSoutput.n127 2.25024
R22352 CSoutput.n261 CSoutput.n171 1.50111
R22353 CSoutput.n209 CSoutput.n195 1.50111
R22354 CSoutput.n271 CSoutput.n137 1.50111
R22355 CSoutput.n217 CSoutput.n216 1.501
R22356 CSoutput.n224 CSoutput.n223 1.501
R22357 CSoutput.n251 CSoutput.n250 1.501
R22358 CSoutput.n265 CSoutput.n176 1.12536
R22359 CSoutput.n265 CSoutput.n177 1.12536
R22360 CSoutput.n265 CSoutput.n264 1.12536
R22361 CSoutput.n225 CSoutput.n205 1.12536
R22362 CSoutput.n231 CSoutput.n205 1.12536
R22363 CSoutput.n233 CSoutput.n205 1.12536
R22364 CSoutput.n275 CSoutput.n142 1.12536
R22365 CSoutput.n275 CSoutput.n143 1.12536
R22366 CSoutput.n275 CSoutput.n274 1.12536
R22367 CSoutput.n265 CSoutput.n172 1.12536
R22368 CSoutput.n265 CSoutput.n173 1.12536
R22369 CSoutput.n265 CSoutput.n175 1.12536
R22370 CSoutput.n255 CSoutput.n205 1.12536
R22371 CSoutput.n235 CSoutput.n205 1.12536
R22372 CSoutput.n237 CSoutput.n205 1.12536
R22373 CSoutput.n275 CSoutput.n138 1.12536
R22374 CSoutput.n275 CSoutput.n139 1.12536
R22375 CSoutput.n275 CSoutput.n141 1.12536
R22376 CSoutput.n31 CSoutput.n30 0.669944
R22377 CSoutput.n62 CSoutput.n61 0.669944
R22378 CSoutput.n344 CSoutput.n342 0.573776
R22379 CSoutput.n346 CSoutput.n344 0.573776
R22380 CSoutput.n348 CSoutput.n346 0.573776
R22381 CSoutput.n350 CSoutput.n348 0.573776
R22382 CSoutput.n352 CSoutput.n350 0.573776
R22383 CSoutput.n354 CSoutput.n352 0.573776
R22384 CSoutput.n329 CSoutput.n327 0.573776
R22385 CSoutput.n331 CSoutput.n329 0.573776
R22386 CSoutput.n333 CSoutput.n331 0.573776
R22387 CSoutput.n335 CSoutput.n333 0.573776
R22388 CSoutput.n337 CSoutput.n335 0.573776
R22389 CSoutput.n339 CSoutput.n337 0.573776
R22390 CSoutput.n386 CSoutput.n384 0.573776
R22391 CSoutput.n384 CSoutput.n382 0.573776
R22392 CSoutput.n382 CSoutput.n380 0.573776
R22393 CSoutput.n380 CSoutput.n378 0.573776
R22394 CSoutput.n378 CSoutput.n376 0.573776
R22395 CSoutput.n376 CSoutput.n374 0.573776
R22396 CSoutput.n371 CSoutput.n369 0.573776
R22397 CSoutput.n369 CSoutput.n367 0.573776
R22398 CSoutput.n367 CSoutput.n365 0.573776
R22399 CSoutput.n365 CSoutput.n363 0.573776
R22400 CSoutput.n363 CSoutput.n361 0.573776
R22401 CSoutput.n361 CSoutput.n359 0.573776
R22402 CSoutput.n389 CSoutput.n276 0.53442
R22403 CSoutput.n312 CSoutput.n310 0.358259
R22404 CSoutput.n314 CSoutput.n312 0.358259
R22405 CSoutput.n316 CSoutput.n314 0.358259
R22406 CSoutput.n318 CSoutput.n316 0.358259
R22407 CSoutput.n320 CSoutput.n318 0.358259
R22408 CSoutput.n322 CSoutput.n320 0.358259
R22409 CSoutput.n296 CSoutput.n294 0.358259
R22410 CSoutput.n298 CSoutput.n296 0.358259
R22411 CSoutput.n300 CSoutput.n298 0.358259
R22412 CSoutput.n302 CSoutput.n300 0.358259
R22413 CSoutput.n304 CSoutput.n302 0.358259
R22414 CSoutput.n306 CSoutput.n304 0.358259
R22415 CSoutput.n281 CSoutput.n279 0.358259
R22416 CSoutput.n283 CSoutput.n281 0.358259
R22417 CSoutput.n285 CSoutput.n283 0.358259
R22418 CSoutput.n287 CSoutput.n285 0.358259
R22419 CSoutput.n289 CSoutput.n287 0.358259
R22420 CSoutput.n291 CSoutput.n289 0.358259
R22421 CSoutput.n124 CSoutput.n122 0.358259
R22422 CSoutput.n122 CSoutput.n120 0.358259
R22423 CSoutput.n120 CSoutput.n118 0.358259
R22424 CSoutput.n118 CSoutput.n116 0.358259
R22425 CSoutput.n116 CSoutput.n114 0.358259
R22426 CSoutput.n114 CSoutput.n112 0.358259
R22427 CSoutput.n108 CSoutput.n106 0.358259
R22428 CSoutput.n106 CSoutput.n104 0.358259
R22429 CSoutput.n104 CSoutput.n102 0.358259
R22430 CSoutput.n102 CSoutput.n100 0.358259
R22431 CSoutput.n100 CSoutput.n98 0.358259
R22432 CSoutput.n98 CSoutput.n96 0.358259
R22433 CSoutput.n93 CSoutput.n91 0.358259
R22434 CSoutput.n91 CSoutput.n89 0.358259
R22435 CSoutput.n89 CSoutput.n87 0.358259
R22436 CSoutput.n87 CSoutput.n85 0.358259
R22437 CSoutput.n85 CSoutput.n83 0.358259
R22438 CSoutput.n83 CSoutput.n81 0.358259
R22439 CSoutput.n21 CSoutput.n20 0.169105
R22440 CSoutput.n21 CSoutput.n16 0.169105
R22441 CSoutput.n26 CSoutput.n16 0.169105
R22442 CSoutput.n27 CSoutput.n26 0.169105
R22443 CSoutput.n27 CSoutput.n14 0.169105
R22444 CSoutput.n32 CSoutput.n14 0.169105
R22445 CSoutput.n33 CSoutput.n32 0.169105
R22446 CSoutput.n34 CSoutput.n33 0.169105
R22447 CSoutput.n34 CSoutput.n12 0.169105
R22448 CSoutput.n39 CSoutput.n12 0.169105
R22449 CSoutput.n40 CSoutput.n39 0.169105
R22450 CSoutput.n40 CSoutput.n10 0.169105
R22451 CSoutput.n45 CSoutput.n10 0.169105
R22452 CSoutput.n46 CSoutput.n45 0.169105
R22453 CSoutput.n47 CSoutput.n46 0.169105
R22454 CSoutput.n47 CSoutput.n8 0.169105
R22455 CSoutput.n52 CSoutput.n8 0.169105
R22456 CSoutput.n53 CSoutput.n52 0.169105
R22457 CSoutput.n53 CSoutput.n6 0.169105
R22458 CSoutput.n58 CSoutput.n6 0.169105
R22459 CSoutput.n59 CSoutput.n58 0.169105
R22460 CSoutput.n60 CSoutput.n59 0.169105
R22461 CSoutput.n60 CSoutput.n4 0.169105
R22462 CSoutput.n66 CSoutput.n4 0.169105
R22463 CSoutput.n67 CSoutput.n66 0.169105
R22464 CSoutput.n68 CSoutput.n67 0.169105
R22465 CSoutput.n68 CSoutput.n2 0.169105
R22466 CSoutput.n73 CSoutput.n2 0.169105
R22467 CSoutput.n74 CSoutput.n73 0.169105
R22468 CSoutput.n74 CSoutput.n0 0.169105
R22469 CSoutput.n78 CSoutput.n0 0.169105
R22470 CSoutput.n219 CSoutput.n218 0.0910737
R22471 CSoutput.n270 CSoutput.n267 0.0723685
R22472 CSoutput.n224 CSoutput.n219 0.0522944
R22473 CSoutput.n267 CSoutput.n266 0.0499135
R22474 CSoutput.n218 CSoutput.n217 0.0499135
R22475 CSoutput.n252 CSoutput.n251 0.0464294
R22476 CSoutput.n260 CSoutput.n257 0.0391444
R22477 CSoutput.n219 CSoutput.t178 0.023435
R22478 CSoutput.n267 CSoutput.t172 0.02262
R22479 CSoutput.n218 CSoutput.t163 0.02262
R22480 CSoutput CSoutput.n389 0.0052
R22481 CSoutput.n189 CSoutput.n172 0.00365111
R22482 CSoutput.n192 CSoutput.n173 0.00365111
R22483 CSoutput.n175 CSoutput.n174 0.00365111
R22484 CSoutput.n217 CSoutput.n176 0.00365111
R22485 CSoutput.n181 CSoutput.n177 0.00365111
R22486 CSoutput.n264 CSoutput.n178 0.00365111
R22487 CSoutput.n255 CSoutput.n254 0.00365111
R22488 CSoutput.n235 CSoutput.n208 0.00365111
R22489 CSoutput.n237 CSoutput.n207 0.00365111
R22490 CSoutput.n225 CSoutput.n224 0.00365111
R22491 CSoutput.n231 CSoutput.n211 0.00365111
R22492 CSoutput.n233 CSoutput.n210 0.00365111
R22493 CSoutput.n155 CSoutput.n138 0.00365111
R22494 CSoutput.n158 CSoutput.n139 0.00365111
R22495 CSoutput.n141 CSoutput.n140 0.00365111
R22496 CSoutput.n251 CSoutput.n142 0.00365111
R22497 CSoutput.n147 CSoutput.n143 0.00365111
R22498 CSoutput.n274 CSoutput.n144 0.00365111
R22499 CSoutput.n186 CSoutput.n176 0.00340054
R22500 CSoutput.n179 CSoutput.n177 0.00340054
R22501 CSoutput.n264 CSoutput.n263 0.00340054
R22502 CSoutput.n259 CSoutput.n172 0.00340054
R22503 CSoutput.n188 CSoutput.n173 0.00340054
R22504 CSoutput.n191 CSoutput.n175 0.00340054
R22505 CSoutput.n230 CSoutput.n225 0.00340054
R22506 CSoutput.n232 CSoutput.n231 0.00340054
R22507 CSoutput.n234 CSoutput.n233 0.00340054
R22508 CSoutput.n256 CSoutput.n255 0.00340054
R22509 CSoutput.n236 CSoutput.n235 0.00340054
R22510 CSoutput.n238 CSoutput.n237 0.00340054
R22511 CSoutput.n152 CSoutput.n142 0.00340054
R22512 CSoutput.n145 CSoutput.n143 0.00340054
R22513 CSoutput.n274 CSoutput.n273 0.00340054
R22514 CSoutput.n269 CSoutput.n138 0.00340054
R22515 CSoutput.n154 CSoutput.n139 0.00340054
R22516 CSoutput.n157 CSoutput.n141 0.00340054
R22517 CSoutput.n187 CSoutput.n181 0.00252698
R22518 CSoutput.n180 CSoutput.n178 0.00252698
R22519 CSoutput.n262 CSoutput.n261 0.00252698
R22520 CSoutput.n190 CSoutput.n188 0.00252698
R22521 CSoutput.n193 CSoutput.n191 0.00252698
R22522 CSoutput.n266 CSoutput.n161 0.00252698
R22523 CSoutput.n187 CSoutput.n186 0.00252698
R22524 CSoutput.n180 CSoutput.n179 0.00252698
R22525 CSoutput.n263 CSoutput.n262 0.00252698
R22526 CSoutput.n190 CSoutput.n189 0.00252698
R22527 CSoutput.n193 CSoutput.n192 0.00252698
R22528 CSoutput.n174 CSoutput.n161 0.00252698
R22529 CSoutput.n241 CSoutput.n211 0.00252698
R22530 CSoutput.n240 CSoutput.n210 0.00252698
R22531 CSoutput.n239 CSoutput.n195 0.00252698
R22532 CSoutput.n236 CSoutput.n206 0.00252698
R22533 CSoutput.n243 CSoutput.n238 0.00252698
R22534 CSoutput.n252 CSoutput.n245 0.00252698
R22535 CSoutput.n241 CSoutput.n230 0.00252698
R22536 CSoutput.n240 CSoutput.n232 0.00252698
R22537 CSoutput.n239 CSoutput.n234 0.00252698
R22538 CSoutput.n254 CSoutput.n206 0.00252698
R22539 CSoutput.n243 CSoutput.n208 0.00252698
R22540 CSoutput.n245 CSoutput.n207 0.00252698
R22541 CSoutput.n153 CSoutput.n147 0.00252698
R22542 CSoutput.n146 CSoutput.n144 0.00252698
R22543 CSoutput.n272 CSoutput.n271 0.00252698
R22544 CSoutput.n156 CSoutput.n154 0.00252698
R22545 CSoutput.n159 CSoutput.n157 0.00252698
R22546 CSoutput.n276 CSoutput.n127 0.00252698
R22547 CSoutput.n153 CSoutput.n152 0.00252698
R22548 CSoutput.n146 CSoutput.n145 0.00252698
R22549 CSoutput.n273 CSoutput.n272 0.00252698
R22550 CSoutput.n156 CSoutput.n155 0.00252698
R22551 CSoutput.n159 CSoutput.n158 0.00252698
R22552 CSoutput.n140 CSoutput.n127 0.00252698
R22553 CSoutput.n261 CSoutput.n260 0.0020275
R22554 CSoutput.n260 CSoutput.n259 0.0020275
R22555 CSoutput.n257 CSoutput.n195 0.0020275
R22556 CSoutput.n257 CSoutput.n256 0.0020275
R22557 CSoutput.n271 CSoutput.n270 0.0020275
R22558 CSoutput.n270 CSoutput.n269 0.0020275
R22559 CSoutput.n171 CSoutput.n170 0.00166668
R22560 CSoutput.n253 CSoutput.n209 0.00166668
R22561 CSoutput.n137 CSoutput.n136 0.00166668
R22562 CSoutput.n275 CSoutput.n137 0.00133328
R22563 CSoutput.n209 CSoutput.n205 0.00133328
R22564 CSoutput.n265 CSoutput.n171 0.00133328
R22565 CSoutput.n268 CSoutput.n160 0.001
R22566 CSoutput.n246 CSoutput.n160 0.001
R22567 CSoutput.n148 CSoutput.n128 0.001
R22568 CSoutput.n247 CSoutput.n128 0.001
R22569 CSoutput.n149 CSoutput.n129 0.001
R22570 CSoutput.n248 CSoutput.n129 0.001
R22571 CSoutput.n150 CSoutput.n130 0.001
R22572 CSoutput.n249 CSoutput.n130 0.001
R22573 CSoutput.n151 CSoutput.n131 0.001
R22574 CSoutput.n250 CSoutput.n131 0.001
R22575 CSoutput.n244 CSoutput.n196 0.001
R22576 CSoutput.n244 CSoutput.n242 0.001
R22577 CSoutput.n226 CSoutput.n197 0.001
R22578 CSoutput.n220 CSoutput.n197 0.001
R22579 CSoutput.n227 CSoutput.n198 0.001
R22580 CSoutput.n221 CSoutput.n198 0.001
R22581 CSoutput.n228 CSoutput.n199 0.001
R22582 CSoutput.n222 CSoutput.n199 0.001
R22583 CSoutput.n229 CSoutput.n200 0.001
R22584 CSoutput.n223 CSoutput.n200 0.001
R22585 CSoutput.n258 CSoutput.n194 0.001
R22586 CSoutput.n212 CSoutput.n194 0.001
R22587 CSoutput.n182 CSoutput.n162 0.001
R22588 CSoutput.n213 CSoutput.n162 0.001
R22589 CSoutput.n183 CSoutput.n163 0.001
R22590 CSoutput.n214 CSoutput.n163 0.001
R22591 CSoutput.n184 CSoutput.n164 0.001
R22592 CSoutput.n215 CSoutput.n164 0.001
R22593 CSoutput.n185 CSoutput.n165 0.001
R22594 CSoutput.n216 CSoutput.n165 0.001
R22595 CSoutput.n216 CSoutput.n166 0.001
R22596 CSoutput.n215 CSoutput.n167 0.001
R22597 CSoutput.n214 CSoutput.n168 0.001
R22598 CSoutput.n213 CSoutput.t175 0.001
R22599 CSoutput.n212 CSoutput.n169 0.001
R22600 CSoutput.n185 CSoutput.n167 0.001
R22601 CSoutput.n184 CSoutput.n168 0.001
R22602 CSoutput.n183 CSoutput.t175 0.001
R22603 CSoutput.n182 CSoutput.n169 0.001
R22604 CSoutput.n258 CSoutput.n170 0.001
R22605 CSoutput.n223 CSoutput.n201 0.001
R22606 CSoutput.n222 CSoutput.n202 0.001
R22607 CSoutput.n221 CSoutput.n203 0.001
R22608 CSoutput.n220 CSoutput.t171 0.001
R22609 CSoutput.n242 CSoutput.n204 0.001
R22610 CSoutput.n229 CSoutput.n202 0.001
R22611 CSoutput.n228 CSoutput.n203 0.001
R22612 CSoutput.n227 CSoutput.t171 0.001
R22613 CSoutput.n226 CSoutput.n204 0.001
R22614 CSoutput.n253 CSoutput.n196 0.001
R22615 CSoutput.n250 CSoutput.n132 0.001
R22616 CSoutput.n249 CSoutput.n133 0.001
R22617 CSoutput.n248 CSoutput.n134 0.001
R22618 CSoutput.n247 CSoutput.t161 0.001
R22619 CSoutput.n246 CSoutput.n135 0.001
R22620 CSoutput.n151 CSoutput.n133 0.001
R22621 CSoutput.n150 CSoutput.n134 0.001
R22622 CSoutput.n149 CSoutput.t161 0.001
R22623 CSoutput.n148 CSoutput.n135 0.001
R22624 CSoutput.n268 CSoutput.n136 0.001
R22625 minus.n53 minus.t28 323.478
R22626 minus.n11 minus.t8 323.478
R22627 minus.n82 minus.t13 297.12
R22628 minus.n80 minus.t15 297.12
R22629 minus.n44 minus.t5 297.12
R22630 minus.n74 minus.t6 297.12
R22631 minus.n46 minus.t26 297.12
R22632 minus.n68 minus.t21 297.12
R22633 minus.n48 minus.t23 297.12
R22634 minus.n62 minus.t16 297.12
R22635 minus.n50 minus.t17 297.12
R22636 minus.n56 minus.t9 297.12
R22637 minus.n52 minus.t27 297.12
R22638 minus.n10 minus.t7 297.12
R22639 minus.n14 minus.t11 297.12
R22640 minus.n16 minus.t10 297.12
R22641 minus.n20 minus.t12 297.12
R22642 minus.n22 minus.t20 297.12
R22643 minus.n26 minus.t18 297.12
R22644 minus.n28 minus.t25 297.12
R22645 minus.n32 minus.t24 297.12
R22646 minus.n34 minus.t14 297.12
R22647 minus.n38 minus.t22 297.12
R22648 minus.n40 minus.t19 297.12
R22649 minus.n88 minus.t2 243.255
R22650 minus.n87 minus.n85 224.169
R22651 minus.n87 minus.n86 223.454
R22652 minus.n55 minus.n54 161.3
R22653 minus.n56 minus.n51 161.3
R22654 minus.n58 minus.n57 161.3
R22655 minus.n59 minus.n50 161.3
R22656 minus.n61 minus.n60 161.3
R22657 minus.n62 minus.n49 161.3
R22658 minus.n64 minus.n63 161.3
R22659 minus.n65 minus.n48 161.3
R22660 minus.n67 minus.n66 161.3
R22661 minus.n68 minus.n47 161.3
R22662 minus.n70 minus.n69 161.3
R22663 minus.n71 minus.n46 161.3
R22664 minus.n73 minus.n72 161.3
R22665 minus.n74 minus.n45 161.3
R22666 minus.n76 minus.n75 161.3
R22667 minus.n77 minus.n44 161.3
R22668 minus.n79 minus.n78 161.3
R22669 minus.n80 minus.n43 161.3
R22670 minus.n81 minus.n42 161.3
R22671 minus.n83 minus.n82 161.3
R22672 minus.n41 minus.n40 161.3
R22673 minus.n39 minus.n0 161.3
R22674 minus.n38 minus.n37 161.3
R22675 minus.n36 minus.n1 161.3
R22676 minus.n35 minus.n34 161.3
R22677 minus.n33 minus.n2 161.3
R22678 minus.n32 minus.n31 161.3
R22679 minus.n30 minus.n3 161.3
R22680 minus.n29 minus.n28 161.3
R22681 minus.n27 minus.n4 161.3
R22682 minus.n26 minus.n25 161.3
R22683 minus.n24 minus.n5 161.3
R22684 minus.n23 minus.n22 161.3
R22685 minus.n21 minus.n6 161.3
R22686 minus.n20 minus.n19 161.3
R22687 minus.n18 minus.n7 161.3
R22688 minus.n17 minus.n16 161.3
R22689 minus.n15 minus.n8 161.3
R22690 minus.n14 minus.n13 161.3
R22691 minus.n12 minus.n9 161.3
R22692 minus.n82 minus.n81 46.0096
R22693 minus.n40 minus.n39 46.0096
R22694 minus.n12 minus.n11 45.0871
R22695 minus.n54 minus.n53 45.0871
R22696 minus.n80 minus.n79 41.6278
R22697 minus.n55 minus.n52 41.6278
R22698 minus.n10 minus.n9 41.6278
R22699 minus.n38 minus.n1 41.6278
R22700 minus.n75 minus.n44 37.246
R22701 minus.n57 minus.n56 37.246
R22702 minus.n15 minus.n14 37.246
R22703 minus.n34 minus.n33 37.246
R22704 minus.n84 minus.n83 33.3925
R22705 minus.n74 minus.n73 32.8641
R22706 minus.n61 minus.n50 32.8641
R22707 minus.n16 minus.n7 32.8641
R22708 minus.n32 minus.n3 32.8641
R22709 minus.n69 minus.n46 28.4823
R22710 minus.n63 minus.n62 28.4823
R22711 minus.n21 minus.n20 28.4823
R22712 minus.n28 minus.n27 28.4823
R22713 minus.n68 minus.n67 24.1005
R22714 minus.n67 minus.n48 24.1005
R22715 minus.n22 minus.n5 24.1005
R22716 minus.n26 minus.n5 24.1005
R22717 minus.n86 minus.t4 19.8005
R22718 minus.n86 minus.t3 19.8005
R22719 minus.n85 minus.t1 19.8005
R22720 minus.n85 minus.t0 19.8005
R22721 minus.n69 minus.n68 19.7187
R22722 minus.n63 minus.n48 19.7187
R22723 minus.n22 minus.n21 19.7187
R22724 minus.n27 minus.n26 19.7187
R22725 minus.n73 minus.n46 15.3369
R22726 minus.n62 minus.n61 15.3369
R22727 minus.n20 minus.n7 15.3369
R22728 minus.n28 minus.n3 15.3369
R22729 minus.n53 minus.n52 14.1472
R22730 minus.n11 minus.n10 14.1472
R22731 minus.n84 minus.n41 12.0933
R22732 minus minus.n89 11.7006
R22733 minus.n75 minus.n74 10.955
R22734 minus.n57 minus.n50 10.955
R22735 minus.n16 minus.n15 10.955
R22736 minus.n33 minus.n32 10.955
R22737 minus.n79 minus.n44 6.57323
R22738 minus.n56 minus.n55 6.57323
R22739 minus.n14 minus.n9 6.57323
R22740 minus.n34 minus.n1 6.57323
R22741 minus.n89 minus.n88 4.80222
R22742 minus.n81 minus.n80 2.19141
R22743 minus.n39 minus.n38 2.19141
R22744 minus.n89 minus.n84 0.972091
R22745 minus.n88 minus.n87 0.716017
R22746 minus.n83 minus.n42 0.189894
R22747 minus.n43 minus.n42 0.189894
R22748 minus.n78 minus.n43 0.189894
R22749 minus.n78 minus.n77 0.189894
R22750 minus.n77 minus.n76 0.189894
R22751 minus.n76 minus.n45 0.189894
R22752 minus.n72 minus.n45 0.189894
R22753 minus.n72 minus.n71 0.189894
R22754 minus.n71 minus.n70 0.189894
R22755 minus.n70 minus.n47 0.189894
R22756 minus.n66 minus.n47 0.189894
R22757 minus.n66 minus.n65 0.189894
R22758 minus.n65 minus.n64 0.189894
R22759 minus.n64 minus.n49 0.189894
R22760 minus.n60 minus.n49 0.189894
R22761 minus.n60 minus.n59 0.189894
R22762 minus.n59 minus.n58 0.189894
R22763 minus.n58 minus.n51 0.189894
R22764 minus.n54 minus.n51 0.189894
R22765 minus.n13 minus.n12 0.189894
R22766 minus.n13 minus.n8 0.189894
R22767 minus.n17 minus.n8 0.189894
R22768 minus.n18 minus.n17 0.189894
R22769 minus.n19 minus.n18 0.189894
R22770 minus.n19 minus.n6 0.189894
R22771 minus.n23 minus.n6 0.189894
R22772 minus.n24 minus.n23 0.189894
R22773 minus.n25 minus.n24 0.189894
R22774 minus.n25 minus.n4 0.189894
R22775 minus.n29 minus.n4 0.189894
R22776 minus.n30 minus.n29 0.189894
R22777 minus.n31 minus.n30 0.189894
R22778 minus.n31 minus.n2 0.189894
R22779 minus.n35 minus.n2 0.189894
R22780 minus.n36 minus.n35 0.189894
R22781 minus.n37 minus.n36 0.189894
R22782 minus.n37 minus.n0 0.189894
R22783 minus.n41 minus.n0 0.189894
R22784 commonsourceibias.n35 commonsourceibias.t16 223.028
R22785 commonsourceibias.n128 commonsourceibias.t85 223.028
R22786 commonsourceibias.n217 commonsourceibias.t75 223.028
R22787 commonsourceibias.n364 commonsourceibias.t54 223.028
R22788 commonsourceibias.n305 commonsourceibias.t91 223.028
R22789 commonsourceibias.n499 commonsourceibias.t78 223.028
R22790 commonsourceibias.n99 commonsourceibias.t60 207.983
R22791 commonsourceibias.n192 commonsourceibias.t92 207.983
R22792 commonsourceibias.n281 commonsourceibias.t81 207.983
R22793 commonsourceibias.n430 commonsourceibias.t8 207.983
R22794 commonsourceibias.n476 commonsourceibias.t110 207.983
R22795 commonsourceibias.n565 commonsourceibias.t97 207.983
R22796 commonsourceibias.n97 commonsourceibias.t14 168.701
R22797 commonsourceibias.n91 commonsourceibias.t38 168.701
R22798 commonsourceibias.n17 commonsourceibias.t4 168.701
R22799 commonsourceibias.n83 commonsourceibias.t28 168.701
R22800 commonsourceibias.n77 commonsourceibias.t62 168.701
R22801 commonsourceibias.n22 commonsourceibias.t18 168.701
R22802 commonsourceibias.n69 commonsourceibias.t26 168.701
R22803 commonsourceibias.n63 commonsourceibias.t6 168.701
R22804 commonsourceibias.n25 commonsourceibias.t32 168.701
R22805 commonsourceibias.n27 commonsourceibias.t42 168.701
R22806 commonsourceibias.n29 commonsourceibias.t20 168.701
R22807 commonsourceibias.n46 commonsourceibias.t30 168.701
R22808 commonsourceibias.n40 commonsourceibias.t56 168.701
R22809 commonsourceibias.n34 commonsourceibias.t12 168.701
R22810 commonsourceibias.n190 commonsourceibias.t106 168.701
R22811 commonsourceibias.n184 commonsourceibias.t119 168.701
R22812 commonsourceibias.n5 commonsourceibias.t84 168.701
R22813 commonsourceibias.n176 commonsourceibias.t100 168.701
R22814 commonsourceibias.n170 commonsourceibias.t114 168.701
R22815 commonsourceibias.n10 commonsourceibias.t80 168.701
R22816 commonsourceibias.n162 commonsourceibias.t76 168.701
R22817 commonsourceibias.n156 commonsourceibias.t105 168.701
R22818 commonsourceibias.n118 commonsourceibias.t121 168.701
R22819 commonsourceibias.n120 commonsourceibias.t71 168.701
R22820 commonsourceibias.n122 commonsourceibias.t99 168.701
R22821 commonsourceibias.n139 commonsourceibias.t95 168.701
R22822 commonsourceibias.n133 commonsourceibias.t109 168.701
R22823 commonsourceibias.n127 commonsourceibias.t89 168.701
R22824 commonsourceibias.n216 commonsourceibias.t77 168.701
R22825 commonsourceibias.n222 commonsourceibias.t96 168.701
R22826 commonsourceibias.n228 commonsourceibias.t82 168.701
R22827 commonsourceibias.n211 commonsourceibias.t86 168.701
R22828 commonsourceibias.n209 commonsourceibias.t127 168.701
R22829 commonsourceibias.n207 commonsourceibias.t108 168.701
R22830 commonsourceibias.n245 commonsourceibias.t93 168.701
R22831 commonsourceibias.n251 commonsourceibias.t67 168.701
R22832 commonsourceibias.n204 commonsourceibias.t70 168.701
R22833 commonsourceibias.n259 commonsourceibias.t101 168.701
R22834 commonsourceibias.n265 commonsourceibias.t87 168.701
R22835 commonsourceibias.n199 commonsourceibias.t74 168.701
R22836 commonsourceibias.n273 commonsourceibias.t107 168.701
R22837 commonsourceibias.n279 commonsourceibias.t94 168.701
R22838 commonsourceibias.n363 commonsourceibias.t52 168.701
R22839 commonsourceibias.n369 commonsourceibias.t2 168.701
R22840 commonsourceibias.n375 commonsourceibias.t48 168.701
R22841 commonsourceibias.n358 commonsourceibias.t40 168.701
R22842 commonsourceibias.n356 commonsourceibias.t58 168.701
R22843 commonsourceibias.n354 commonsourceibias.t50 168.701
R22844 commonsourceibias.n392 commonsourceibias.t24 168.701
R22845 commonsourceibias.n398 commonsourceibias.t44 168.701
R22846 commonsourceibias.n400 commonsourceibias.t36 168.701
R22847 commonsourceibias.n407 commonsourceibias.t10 168.701
R22848 commonsourceibias.n413 commonsourceibias.t46 168.701
R22849 commonsourceibias.n415 commonsourceibias.t22 168.701
R22850 commonsourceibias.n422 commonsourceibias.t0 168.701
R22851 commonsourceibias.n428 commonsourceibias.t34 168.701
R22852 commonsourceibias.n474 commonsourceibias.t123 168.701
R22853 commonsourceibias.n468 commonsourceibias.t68 168.701
R22854 commonsourceibias.n461 commonsourceibias.t102 168.701
R22855 commonsourceibias.n459 commonsourceibias.t117 168.701
R22856 commonsourceibias.n453 commonsourceibias.t64 168.701
R22857 commonsourceibias.n446 commonsourceibias.t72 168.701
R22858 commonsourceibias.n444 commonsourceibias.t90 168.701
R22859 commonsourceibias.n304 commonsourceibias.t83 168.701
R22860 commonsourceibias.n310 commonsourceibias.t126 168.701
R22861 commonsourceibias.n316 commonsourceibias.t113 168.701
R22862 commonsourceibias.n299 commonsourceibias.t116 168.701
R22863 commonsourceibias.n297 commonsourceibias.t66 168.701
R22864 commonsourceibias.n295 commonsourceibias.t69 168.701
R22865 commonsourceibias.n333 commonsourceibias.t122 168.701
R22866 commonsourceibias.n498 commonsourceibias.t73 168.701
R22867 commonsourceibias.n504 commonsourceibias.t115 168.701
R22868 commonsourceibias.n510 commonsourceibias.t98 168.701
R22869 commonsourceibias.n493 commonsourceibias.t103 168.701
R22870 commonsourceibias.n491 commonsourceibias.t120 168.701
R22871 commonsourceibias.n489 commonsourceibias.t125 168.701
R22872 commonsourceibias.n527 commonsourceibias.t111 168.701
R22873 commonsourceibias.n533 commonsourceibias.t79 168.701
R22874 commonsourceibias.n535 commonsourceibias.t65 168.701
R22875 commonsourceibias.n542 commonsourceibias.t118 168.701
R22876 commonsourceibias.n548 commonsourceibias.t104 168.701
R22877 commonsourceibias.n550 commonsourceibias.t88 168.701
R22878 commonsourceibias.n557 commonsourceibias.t124 168.701
R22879 commonsourceibias.n563 commonsourceibias.t112 168.701
R22880 commonsourceibias.n36 commonsourceibias.n33 161.3
R22881 commonsourceibias.n38 commonsourceibias.n37 161.3
R22882 commonsourceibias.n39 commonsourceibias.n32 161.3
R22883 commonsourceibias.n42 commonsourceibias.n41 161.3
R22884 commonsourceibias.n43 commonsourceibias.n31 161.3
R22885 commonsourceibias.n45 commonsourceibias.n44 161.3
R22886 commonsourceibias.n47 commonsourceibias.n30 161.3
R22887 commonsourceibias.n49 commonsourceibias.n48 161.3
R22888 commonsourceibias.n51 commonsourceibias.n50 161.3
R22889 commonsourceibias.n52 commonsourceibias.n28 161.3
R22890 commonsourceibias.n54 commonsourceibias.n53 161.3
R22891 commonsourceibias.n56 commonsourceibias.n55 161.3
R22892 commonsourceibias.n57 commonsourceibias.n26 161.3
R22893 commonsourceibias.n59 commonsourceibias.n58 161.3
R22894 commonsourceibias.n61 commonsourceibias.n60 161.3
R22895 commonsourceibias.n62 commonsourceibias.n24 161.3
R22896 commonsourceibias.n65 commonsourceibias.n64 161.3
R22897 commonsourceibias.n66 commonsourceibias.n23 161.3
R22898 commonsourceibias.n68 commonsourceibias.n67 161.3
R22899 commonsourceibias.n70 commonsourceibias.n21 161.3
R22900 commonsourceibias.n72 commonsourceibias.n71 161.3
R22901 commonsourceibias.n73 commonsourceibias.n20 161.3
R22902 commonsourceibias.n75 commonsourceibias.n74 161.3
R22903 commonsourceibias.n76 commonsourceibias.n19 161.3
R22904 commonsourceibias.n79 commonsourceibias.n78 161.3
R22905 commonsourceibias.n80 commonsourceibias.n18 161.3
R22906 commonsourceibias.n82 commonsourceibias.n81 161.3
R22907 commonsourceibias.n84 commonsourceibias.n16 161.3
R22908 commonsourceibias.n86 commonsourceibias.n85 161.3
R22909 commonsourceibias.n87 commonsourceibias.n15 161.3
R22910 commonsourceibias.n89 commonsourceibias.n88 161.3
R22911 commonsourceibias.n90 commonsourceibias.n14 161.3
R22912 commonsourceibias.n93 commonsourceibias.n92 161.3
R22913 commonsourceibias.n94 commonsourceibias.n13 161.3
R22914 commonsourceibias.n96 commonsourceibias.n95 161.3
R22915 commonsourceibias.n98 commonsourceibias.n12 161.3
R22916 commonsourceibias.n129 commonsourceibias.n126 161.3
R22917 commonsourceibias.n131 commonsourceibias.n130 161.3
R22918 commonsourceibias.n132 commonsourceibias.n125 161.3
R22919 commonsourceibias.n135 commonsourceibias.n134 161.3
R22920 commonsourceibias.n136 commonsourceibias.n124 161.3
R22921 commonsourceibias.n138 commonsourceibias.n137 161.3
R22922 commonsourceibias.n140 commonsourceibias.n123 161.3
R22923 commonsourceibias.n142 commonsourceibias.n141 161.3
R22924 commonsourceibias.n144 commonsourceibias.n143 161.3
R22925 commonsourceibias.n145 commonsourceibias.n121 161.3
R22926 commonsourceibias.n147 commonsourceibias.n146 161.3
R22927 commonsourceibias.n149 commonsourceibias.n148 161.3
R22928 commonsourceibias.n150 commonsourceibias.n119 161.3
R22929 commonsourceibias.n152 commonsourceibias.n151 161.3
R22930 commonsourceibias.n154 commonsourceibias.n153 161.3
R22931 commonsourceibias.n155 commonsourceibias.n117 161.3
R22932 commonsourceibias.n158 commonsourceibias.n157 161.3
R22933 commonsourceibias.n159 commonsourceibias.n11 161.3
R22934 commonsourceibias.n161 commonsourceibias.n160 161.3
R22935 commonsourceibias.n163 commonsourceibias.n9 161.3
R22936 commonsourceibias.n165 commonsourceibias.n164 161.3
R22937 commonsourceibias.n166 commonsourceibias.n8 161.3
R22938 commonsourceibias.n168 commonsourceibias.n167 161.3
R22939 commonsourceibias.n169 commonsourceibias.n7 161.3
R22940 commonsourceibias.n172 commonsourceibias.n171 161.3
R22941 commonsourceibias.n173 commonsourceibias.n6 161.3
R22942 commonsourceibias.n175 commonsourceibias.n174 161.3
R22943 commonsourceibias.n177 commonsourceibias.n4 161.3
R22944 commonsourceibias.n179 commonsourceibias.n178 161.3
R22945 commonsourceibias.n180 commonsourceibias.n3 161.3
R22946 commonsourceibias.n182 commonsourceibias.n181 161.3
R22947 commonsourceibias.n183 commonsourceibias.n2 161.3
R22948 commonsourceibias.n186 commonsourceibias.n185 161.3
R22949 commonsourceibias.n187 commonsourceibias.n1 161.3
R22950 commonsourceibias.n189 commonsourceibias.n188 161.3
R22951 commonsourceibias.n191 commonsourceibias.n0 161.3
R22952 commonsourceibias.n280 commonsourceibias.n194 161.3
R22953 commonsourceibias.n278 commonsourceibias.n277 161.3
R22954 commonsourceibias.n276 commonsourceibias.n195 161.3
R22955 commonsourceibias.n275 commonsourceibias.n274 161.3
R22956 commonsourceibias.n272 commonsourceibias.n196 161.3
R22957 commonsourceibias.n271 commonsourceibias.n270 161.3
R22958 commonsourceibias.n269 commonsourceibias.n197 161.3
R22959 commonsourceibias.n268 commonsourceibias.n267 161.3
R22960 commonsourceibias.n266 commonsourceibias.n198 161.3
R22961 commonsourceibias.n264 commonsourceibias.n263 161.3
R22962 commonsourceibias.n262 commonsourceibias.n200 161.3
R22963 commonsourceibias.n261 commonsourceibias.n260 161.3
R22964 commonsourceibias.n258 commonsourceibias.n201 161.3
R22965 commonsourceibias.n257 commonsourceibias.n256 161.3
R22966 commonsourceibias.n255 commonsourceibias.n202 161.3
R22967 commonsourceibias.n254 commonsourceibias.n253 161.3
R22968 commonsourceibias.n252 commonsourceibias.n203 161.3
R22969 commonsourceibias.n250 commonsourceibias.n249 161.3
R22970 commonsourceibias.n248 commonsourceibias.n205 161.3
R22971 commonsourceibias.n247 commonsourceibias.n246 161.3
R22972 commonsourceibias.n244 commonsourceibias.n206 161.3
R22973 commonsourceibias.n243 commonsourceibias.n242 161.3
R22974 commonsourceibias.n241 commonsourceibias.n240 161.3
R22975 commonsourceibias.n239 commonsourceibias.n208 161.3
R22976 commonsourceibias.n238 commonsourceibias.n237 161.3
R22977 commonsourceibias.n236 commonsourceibias.n235 161.3
R22978 commonsourceibias.n234 commonsourceibias.n210 161.3
R22979 commonsourceibias.n233 commonsourceibias.n232 161.3
R22980 commonsourceibias.n231 commonsourceibias.n230 161.3
R22981 commonsourceibias.n229 commonsourceibias.n212 161.3
R22982 commonsourceibias.n227 commonsourceibias.n226 161.3
R22983 commonsourceibias.n225 commonsourceibias.n213 161.3
R22984 commonsourceibias.n224 commonsourceibias.n223 161.3
R22985 commonsourceibias.n221 commonsourceibias.n214 161.3
R22986 commonsourceibias.n220 commonsourceibias.n219 161.3
R22987 commonsourceibias.n218 commonsourceibias.n215 161.3
R22988 commonsourceibias.n429 commonsourceibias.n343 161.3
R22989 commonsourceibias.n427 commonsourceibias.n426 161.3
R22990 commonsourceibias.n425 commonsourceibias.n344 161.3
R22991 commonsourceibias.n424 commonsourceibias.n423 161.3
R22992 commonsourceibias.n421 commonsourceibias.n345 161.3
R22993 commonsourceibias.n420 commonsourceibias.n419 161.3
R22994 commonsourceibias.n418 commonsourceibias.n346 161.3
R22995 commonsourceibias.n417 commonsourceibias.n416 161.3
R22996 commonsourceibias.n414 commonsourceibias.n347 161.3
R22997 commonsourceibias.n412 commonsourceibias.n411 161.3
R22998 commonsourceibias.n410 commonsourceibias.n348 161.3
R22999 commonsourceibias.n409 commonsourceibias.n408 161.3
R23000 commonsourceibias.n406 commonsourceibias.n349 161.3
R23001 commonsourceibias.n405 commonsourceibias.n404 161.3
R23002 commonsourceibias.n403 commonsourceibias.n350 161.3
R23003 commonsourceibias.n402 commonsourceibias.n401 161.3
R23004 commonsourceibias.n399 commonsourceibias.n351 161.3
R23005 commonsourceibias.n397 commonsourceibias.n396 161.3
R23006 commonsourceibias.n395 commonsourceibias.n352 161.3
R23007 commonsourceibias.n394 commonsourceibias.n393 161.3
R23008 commonsourceibias.n391 commonsourceibias.n353 161.3
R23009 commonsourceibias.n390 commonsourceibias.n389 161.3
R23010 commonsourceibias.n388 commonsourceibias.n387 161.3
R23011 commonsourceibias.n386 commonsourceibias.n355 161.3
R23012 commonsourceibias.n385 commonsourceibias.n384 161.3
R23013 commonsourceibias.n383 commonsourceibias.n382 161.3
R23014 commonsourceibias.n381 commonsourceibias.n357 161.3
R23015 commonsourceibias.n380 commonsourceibias.n379 161.3
R23016 commonsourceibias.n378 commonsourceibias.n377 161.3
R23017 commonsourceibias.n376 commonsourceibias.n359 161.3
R23018 commonsourceibias.n374 commonsourceibias.n373 161.3
R23019 commonsourceibias.n372 commonsourceibias.n360 161.3
R23020 commonsourceibias.n371 commonsourceibias.n370 161.3
R23021 commonsourceibias.n368 commonsourceibias.n361 161.3
R23022 commonsourceibias.n367 commonsourceibias.n366 161.3
R23023 commonsourceibias.n365 commonsourceibias.n362 161.3
R23024 commonsourceibias.n335 commonsourceibias.n334 161.3
R23025 commonsourceibias.n332 commonsourceibias.n294 161.3
R23026 commonsourceibias.n331 commonsourceibias.n330 161.3
R23027 commonsourceibias.n329 commonsourceibias.n328 161.3
R23028 commonsourceibias.n327 commonsourceibias.n296 161.3
R23029 commonsourceibias.n326 commonsourceibias.n325 161.3
R23030 commonsourceibias.n324 commonsourceibias.n323 161.3
R23031 commonsourceibias.n322 commonsourceibias.n298 161.3
R23032 commonsourceibias.n321 commonsourceibias.n320 161.3
R23033 commonsourceibias.n319 commonsourceibias.n318 161.3
R23034 commonsourceibias.n317 commonsourceibias.n300 161.3
R23035 commonsourceibias.n315 commonsourceibias.n314 161.3
R23036 commonsourceibias.n313 commonsourceibias.n301 161.3
R23037 commonsourceibias.n312 commonsourceibias.n311 161.3
R23038 commonsourceibias.n309 commonsourceibias.n302 161.3
R23039 commonsourceibias.n308 commonsourceibias.n307 161.3
R23040 commonsourceibias.n306 commonsourceibias.n303 161.3
R23041 commonsourceibias.n441 commonsourceibias.n293 161.3
R23042 commonsourceibias.n475 commonsourceibias.n284 161.3
R23043 commonsourceibias.n473 commonsourceibias.n472 161.3
R23044 commonsourceibias.n471 commonsourceibias.n285 161.3
R23045 commonsourceibias.n470 commonsourceibias.n469 161.3
R23046 commonsourceibias.n467 commonsourceibias.n286 161.3
R23047 commonsourceibias.n466 commonsourceibias.n465 161.3
R23048 commonsourceibias.n464 commonsourceibias.n287 161.3
R23049 commonsourceibias.n463 commonsourceibias.n462 161.3
R23050 commonsourceibias.n460 commonsourceibias.n288 161.3
R23051 commonsourceibias.n458 commonsourceibias.n457 161.3
R23052 commonsourceibias.n456 commonsourceibias.n289 161.3
R23053 commonsourceibias.n455 commonsourceibias.n454 161.3
R23054 commonsourceibias.n452 commonsourceibias.n290 161.3
R23055 commonsourceibias.n451 commonsourceibias.n450 161.3
R23056 commonsourceibias.n449 commonsourceibias.n291 161.3
R23057 commonsourceibias.n448 commonsourceibias.n447 161.3
R23058 commonsourceibias.n445 commonsourceibias.n292 161.3
R23059 commonsourceibias.n443 commonsourceibias.n442 161.3
R23060 commonsourceibias.n564 commonsourceibias.n478 161.3
R23061 commonsourceibias.n562 commonsourceibias.n561 161.3
R23062 commonsourceibias.n560 commonsourceibias.n479 161.3
R23063 commonsourceibias.n559 commonsourceibias.n558 161.3
R23064 commonsourceibias.n556 commonsourceibias.n480 161.3
R23065 commonsourceibias.n555 commonsourceibias.n554 161.3
R23066 commonsourceibias.n553 commonsourceibias.n481 161.3
R23067 commonsourceibias.n552 commonsourceibias.n551 161.3
R23068 commonsourceibias.n549 commonsourceibias.n482 161.3
R23069 commonsourceibias.n547 commonsourceibias.n546 161.3
R23070 commonsourceibias.n545 commonsourceibias.n483 161.3
R23071 commonsourceibias.n544 commonsourceibias.n543 161.3
R23072 commonsourceibias.n541 commonsourceibias.n484 161.3
R23073 commonsourceibias.n540 commonsourceibias.n539 161.3
R23074 commonsourceibias.n538 commonsourceibias.n485 161.3
R23075 commonsourceibias.n537 commonsourceibias.n536 161.3
R23076 commonsourceibias.n534 commonsourceibias.n486 161.3
R23077 commonsourceibias.n532 commonsourceibias.n531 161.3
R23078 commonsourceibias.n530 commonsourceibias.n487 161.3
R23079 commonsourceibias.n529 commonsourceibias.n528 161.3
R23080 commonsourceibias.n526 commonsourceibias.n488 161.3
R23081 commonsourceibias.n525 commonsourceibias.n524 161.3
R23082 commonsourceibias.n523 commonsourceibias.n522 161.3
R23083 commonsourceibias.n521 commonsourceibias.n490 161.3
R23084 commonsourceibias.n520 commonsourceibias.n519 161.3
R23085 commonsourceibias.n518 commonsourceibias.n517 161.3
R23086 commonsourceibias.n516 commonsourceibias.n492 161.3
R23087 commonsourceibias.n515 commonsourceibias.n514 161.3
R23088 commonsourceibias.n513 commonsourceibias.n512 161.3
R23089 commonsourceibias.n511 commonsourceibias.n494 161.3
R23090 commonsourceibias.n509 commonsourceibias.n508 161.3
R23091 commonsourceibias.n507 commonsourceibias.n495 161.3
R23092 commonsourceibias.n506 commonsourceibias.n505 161.3
R23093 commonsourceibias.n503 commonsourceibias.n496 161.3
R23094 commonsourceibias.n502 commonsourceibias.n501 161.3
R23095 commonsourceibias.n500 commonsourceibias.n497 161.3
R23096 commonsourceibias.n111 commonsourceibias.n109 81.5057
R23097 commonsourceibias.n338 commonsourceibias.n336 81.5057
R23098 commonsourceibias.n111 commonsourceibias.n110 80.9324
R23099 commonsourceibias.n113 commonsourceibias.n112 80.9324
R23100 commonsourceibias.n115 commonsourceibias.n114 80.9324
R23101 commonsourceibias.n108 commonsourceibias.n107 80.9324
R23102 commonsourceibias.n106 commonsourceibias.n105 80.9324
R23103 commonsourceibias.n104 commonsourceibias.n103 80.9324
R23104 commonsourceibias.n102 commonsourceibias.n101 80.9324
R23105 commonsourceibias.n433 commonsourceibias.n432 80.9324
R23106 commonsourceibias.n435 commonsourceibias.n434 80.9324
R23107 commonsourceibias.n437 commonsourceibias.n436 80.9324
R23108 commonsourceibias.n439 commonsourceibias.n438 80.9324
R23109 commonsourceibias.n342 commonsourceibias.n341 80.9324
R23110 commonsourceibias.n340 commonsourceibias.n339 80.9324
R23111 commonsourceibias.n338 commonsourceibias.n337 80.9324
R23112 commonsourceibias.n100 commonsourceibias.n99 80.6037
R23113 commonsourceibias.n193 commonsourceibias.n192 80.6037
R23114 commonsourceibias.n282 commonsourceibias.n281 80.6037
R23115 commonsourceibias.n431 commonsourceibias.n430 80.6037
R23116 commonsourceibias.n477 commonsourceibias.n476 80.6037
R23117 commonsourceibias.n566 commonsourceibias.n565 80.6037
R23118 commonsourceibias.n85 commonsourceibias.n84 56.5617
R23119 commonsourceibias.n71 commonsourceibias.n70 56.5617
R23120 commonsourceibias.n62 commonsourceibias.n61 56.5617
R23121 commonsourceibias.n48 commonsourceibias.n47 56.5617
R23122 commonsourceibias.n178 commonsourceibias.n177 56.5617
R23123 commonsourceibias.n164 commonsourceibias.n163 56.5617
R23124 commonsourceibias.n155 commonsourceibias.n154 56.5617
R23125 commonsourceibias.n141 commonsourceibias.n140 56.5617
R23126 commonsourceibias.n230 commonsourceibias.n229 56.5617
R23127 commonsourceibias.n244 commonsourceibias.n243 56.5617
R23128 commonsourceibias.n253 commonsourceibias.n252 56.5617
R23129 commonsourceibias.n267 commonsourceibias.n266 56.5617
R23130 commonsourceibias.n377 commonsourceibias.n376 56.5617
R23131 commonsourceibias.n391 commonsourceibias.n390 56.5617
R23132 commonsourceibias.n401 commonsourceibias.n399 56.5617
R23133 commonsourceibias.n416 commonsourceibias.n414 56.5617
R23134 commonsourceibias.n462 commonsourceibias.n460 56.5617
R23135 commonsourceibias.n447 commonsourceibias.n445 56.5617
R23136 commonsourceibias.n318 commonsourceibias.n317 56.5617
R23137 commonsourceibias.n332 commonsourceibias.n331 56.5617
R23138 commonsourceibias.n512 commonsourceibias.n511 56.5617
R23139 commonsourceibias.n526 commonsourceibias.n525 56.5617
R23140 commonsourceibias.n536 commonsourceibias.n534 56.5617
R23141 commonsourceibias.n551 commonsourceibias.n549 56.5617
R23142 commonsourceibias.n76 commonsourceibias.n75 56.0773
R23143 commonsourceibias.n57 commonsourceibias.n56 56.0773
R23144 commonsourceibias.n169 commonsourceibias.n168 56.0773
R23145 commonsourceibias.n150 commonsourceibias.n149 56.0773
R23146 commonsourceibias.n239 commonsourceibias.n238 56.0773
R23147 commonsourceibias.n258 commonsourceibias.n257 56.0773
R23148 commonsourceibias.n386 commonsourceibias.n385 56.0773
R23149 commonsourceibias.n406 commonsourceibias.n405 56.0773
R23150 commonsourceibias.n452 commonsourceibias.n451 56.0773
R23151 commonsourceibias.n327 commonsourceibias.n326 56.0773
R23152 commonsourceibias.n521 commonsourceibias.n520 56.0773
R23153 commonsourceibias.n541 commonsourceibias.n540 56.0773
R23154 commonsourceibias.n99 commonsourceibias.n98 55.3321
R23155 commonsourceibias.n192 commonsourceibias.n191 55.3321
R23156 commonsourceibias.n281 commonsourceibias.n280 55.3321
R23157 commonsourceibias.n430 commonsourceibias.n429 55.3321
R23158 commonsourceibias.n476 commonsourceibias.n475 55.3321
R23159 commonsourceibias.n565 commonsourceibias.n564 55.3321
R23160 commonsourceibias.n90 commonsourceibias.n89 55.1086
R23161 commonsourceibias.n41 commonsourceibias.n31 55.1086
R23162 commonsourceibias.n183 commonsourceibias.n182 55.1086
R23163 commonsourceibias.n134 commonsourceibias.n124 55.1086
R23164 commonsourceibias.n223 commonsourceibias.n213 55.1086
R23165 commonsourceibias.n272 commonsourceibias.n271 55.1086
R23166 commonsourceibias.n370 commonsourceibias.n360 55.1086
R23167 commonsourceibias.n421 commonsourceibias.n420 55.1086
R23168 commonsourceibias.n467 commonsourceibias.n466 55.1086
R23169 commonsourceibias.n311 commonsourceibias.n301 55.1086
R23170 commonsourceibias.n505 commonsourceibias.n495 55.1086
R23171 commonsourceibias.n556 commonsourceibias.n555 55.1086
R23172 commonsourceibias.n35 commonsourceibias.n34 47.4592
R23173 commonsourceibias.n128 commonsourceibias.n127 47.4592
R23174 commonsourceibias.n217 commonsourceibias.n216 47.4592
R23175 commonsourceibias.n364 commonsourceibias.n363 47.4592
R23176 commonsourceibias.n305 commonsourceibias.n304 47.4592
R23177 commonsourceibias.n499 commonsourceibias.n498 47.4592
R23178 commonsourceibias.n218 commonsourceibias.n217 44.0436
R23179 commonsourceibias.n365 commonsourceibias.n364 44.0436
R23180 commonsourceibias.n306 commonsourceibias.n305 44.0436
R23181 commonsourceibias.n500 commonsourceibias.n499 44.0436
R23182 commonsourceibias.n36 commonsourceibias.n35 44.0436
R23183 commonsourceibias.n129 commonsourceibias.n128 44.0436
R23184 commonsourceibias.n92 commonsourceibias.n13 42.5146
R23185 commonsourceibias.n39 commonsourceibias.n38 42.5146
R23186 commonsourceibias.n185 commonsourceibias.n1 42.5146
R23187 commonsourceibias.n132 commonsourceibias.n131 42.5146
R23188 commonsourceibias.n221 commonsourceibias.n220 42.5146
R23189 commonsourceibias.n274 commonsourceibias.n195 42.5146
R23190 commonsourceibias.n368 commonsourceibias.n367 42.5146
R23191 commonsourceibias.n423 commonsourceibias.n344 42.5146
R23192 commonsourceibias.n469 commonsourceibias.n285 42.5146
R23193 commonsourceibias.n309 commonsourceibias.n308 42.5146
R23194 commonsourceibias.n503 commonsourceibias.n502 42.5146
R23195 commonsourceibias.n558 commonsourceibias.n479 42.5146
R23196 commonsourceibias.n78 commonsourceibias.n18 41.5458
R23197 commonsourceibias.n53 commonsourceibias.n52 41.5458
R23198 commonsourceibias.n171 commonsourceibias.n6 41.5458
R23199 commonsourceibias.n146 commonsourceibias.n145 41.5458
R23200 commonsourceibias.n235 commonsourceibias.n234 41.5458
R23201 commonsourceibias.n260 commonsourceibias.n200 41.5458
R23202 commonsourceibias.n382 commonsourceibias.n381 41.5458
R23203 commonsourceibias.n408 commonsourceibias.n348 41.5458
R23204 commonsourceibias.n454 commonsourceibias.n289 41.5458
R23205 commonsourceibias.n323 commonsourceibias.n322 41.5458
R23206 commonsourceibias.n517 commonsourceibias.n516 41.5458
R23207 commonsourceibias.n543 commonsourceibias.n483 41.5458
R23208 commonsourceibias.n68 commonsourceibias.n23 40.577
R23209 commonsourceibias.n64 commonsourceibias.n23 40.577
R23210 commonsourceibias.n161 commonsourceibias.n11 40.577
R23211 commonsourceibias.n157 commonsourceibias.n11 40.577
R23212 commonsourceibias.n246 commonsourceibias.n205 40.577
R23213 commonsourceibias.n250 commonsourceibias.n205 40.577
R23214 commonsourceibias.n393 commonsourceibias.n352 40.577
R23215 commonsourceibias.n397 commonsourceibias.n352 40.577
R23216 commonsourceibias.n443 commonsourceibias.n293 40.577
R23217 commonsourceibias.n334 commonsourceibias.n293 40.577
R23218 commonsourceibias.n528 commonsourceibias.n487 40.577
R23219 commonsourceibias.n532 commonsourceibias.n487 40.577
R23220 commonsourceibias.n82 commonsourceibias.n18 39.6083
R23221 commonsourceibias.n52 commonsourceibias.n51 39.6083
R23222 commonsourceibias.n175 commonsourceibias.n6 39.6083
R23223 commonsourceibias.n145 commonsourceibias.n144 39.6083
R23224 commonsourceibias.n234 commonsourceibias.n233 39.6083
R23225 commonsourceibias.n264 commonsourceibias.n200 39.6083
R23226 commonsourceibias.n381 commonsourceibias.n380 39.6083
R23227 commonsourceibias.n412 commonsourceibias.n348 39.6083
R23228 commonsourceibias.n458 commonsourceibias.n289 39.6083
R23229 commonsourceibias.n322 commonsourceibias.n321 39.6083
R23230 commonsourceibias.n516 commonsourceibias.n515 39.6083
R23231 commonsourceibias.n547 commonsourceibias.n483 39.6083
R23232 commonsourceibias.n96 commonsourceibias.n13 38.6395
R23233 commonsourceibias.n38 commonsourceibias.n33 38.6395
R23234 commonsourceibias.n189 commonsourceibias.n1 38.6395
R23235 commonsourceibias.n131 commonsourceibias.n126 38.6395
R23236 commonsourceibias.n220 commonsourceibias.n215 38.6395
R23237 commonsourceibias.n278 commonsourceibias.n195 38.6395
R23238 commonsourceibias.n367 commonsourceibias.n362 38.6395
R23239 commonsourceibias.n427 commonsourceibias.n344 38.6395
R23240 commonsourceibias.n473 commonsourceibias.n285 38.6395
R23241 commonsourceibias.n308 commonsourceibias.n303 38.6395
R23242 commonsourceibias.n502 commonsourceibias.n497 38.6395
R23243 commonsourceibias.n562 commonsourceibias.n479 38.6395
R23244 commonsourceibias.n89 commonsourceibias.n15 26.0455
R23245 commonsourceibias.n45 commonsourceibias.n31 26.0455
R23246 commonsourceibias.n182 commonsourceibias.n3 26.0455
R23247 commonsourceibias.n138 commonsourceibias.n124 26.0455
R23248 commonsourceibias.n227 commonsourceibias.n213 26.0455
R23249 commonsourceibias.n271 commonsourceibias.n197 26.0455
R23250 commonsourceibias.n374 commonsourceibias.n360 26.0455
R23251 commonsourceibias.n420 commonsourceibias.n346 26.0455
R23252 commonsourceibias.n466 commonsourceibias.n287 26.0455
R23253 commonsourceibias.n315 commonsourceibias.n301 26.0455
R23254 commonsourceibias.n509 commonsourceibias.n495 26.0455
R23255 commonsourceibias.n555 commonsourceibias.n481 26.0455
R23256 commonsourceibias.n75 commonsourceibias.n20 25.0767
R23257 commonsourceibias.n58 commonsourceibias.n57 25.0767
R23258 commonsourceibias.n168 commonsourceibias.n8 25.0767
R23259 commonsourceibias.n151 commonsourceibias.n150 25.0767
R23260 commonsourceibias.n240 commonsourceibias.n239 25.0767
R23261 commonsourceibias.n257 commonsourceibias.n202 25.0767
R23262 commonsourceibias.n387 commonsourceibias.n386 25.0767
R23263 commonsourceibias.n405 commonsourceibias.n350 25.0767
R23264 commonsourceibias.n451 commonsourceibias.n291 25.0767
R23265 commonsourceibias.n328 commonsourceibias.n327 25.0767
R23266 commonsourceibias.n522 commonsourceibias.n521 25.0767
R23267 commonsourceibias.n540 commonsourceibias.n485 25.0767
R23268 commonsourceibias.n71 commonsourceibias.n22 24.3464
R23269 commonsourceibias.n61 commonsourceibias.n25 24.3464
R23270 commonsourceibias.n164 commonsourceibias.n10 24.3464
R23271 commonsourceibias.n154 commonsourceibias.n118 24.3464
R23272 commonsourceibias.n243 commonsourceibias.n207 24.3464
R23273 commonsourceibias.n253 commonsourceibias.n204 24.3464
R23274 commonsourceibias.n390 commonsourceibias.n354 24.3464
R23275 commonsourceibias.n401 commonsourceibias.n400 24.3464
R23276 commonsourceibias.n447 commonsourceibias.n446 24.3464
R23277 commonsourceibias.n331 commonsourceibias.n295 24.3464
R23278 commonsourceibias.n525 commonsourceibias.n489 24.3464
R23279 commonsourceibias.n536 commonsourceibias.n535 24.3464
R23280 commonsourceibias.n85 commonsourceibias.n17 23.8546
R23281 commonsourceibias.n47 commonsourceibias.n46 23.8546
R23282 commonsourceibias.n178 commonsourceibias.n5 23.8546
R23283 commonsourceibias.n140 commonsourceibias.n139 23.8546
R23284 commonsourceibias.n229 commonsourceibias.n228 23.8546
R23285 commonsourceibias.n267 commonsourceibias.n199 23.8546
R23286 commonsourceibias.n376 commonsourceibias.n375 23.8546
R23287 commonsourceibias.n416 commonsourceibias.n415 23.8546
R23288 commonsourceibias.n462 commonsourceibias.n461 23.8546
R23289 commonsourceibias.n317 commonsourceibias.n316 23.8546
R23290 commonsourceibias.n511 commonsourceibias.n510 23.8546
R23291 commonsourceibias.n551 commonsourceibias.n550 23.8546
R23292 commonsourceibias.n98 commonsourceibias.n97 17.4607
R23293 commonsourceibias.n191 commonsourceibias.n190 17.4607
R23294 commonsourceibias.n280 commonsourceibias.n279 17.4607
R23295 commonsourceibias.n429 commonsourceibias.n428 17.4607
R23296 commonsourceibias.n475 commonsourceibias.n474 17.4607
R23297 commonsourceibias.n564 commonsourceibias.n563 17.4607
R23298 commonsourceibias.n84 commonsourceibias.n83 16.9689
R23299 commonsourceibias.n48 commonsourceibias.n29 16.9689
R23300 commonsourceibias.n177 commonsourceibias.n176 16.9689
R23301 commonsourceibias.n141 commonsourceibias.n122 16.9689
R23302 commonsourceibias.n230 commonsourceibias.n211 16.9689
R23303 commonsourceibias.n266 commonsourceibias.n265 16.9689
R23304 commonsourceibias.n377 commonsourceibias.n358 16.9689
R23305 commonsourceibias.n414 commonsourceibias.n413 16.9689
R23306 commonsourceibias.n460 commonsourceibias.n459 16.9689
R23307 commonsourceibias.n318 commonsourceibias.n299 16.9689
R23308 commonsourceibias.n512 commonsourceibias.n493 16.9689
R23309 commonsourceibias.n549 commonsourceibias.n548 16.9689
R23310 commonsourceibias.n70 commonsourceibias.n69 16.477
R23311 commonsourceibias.n63 commonsourceibias.n62 16.477
R23312 commonsourceibias.n163 commonsourceibias.n162 16.477
R23313 commonsourceibias.n156 commonsourceibias.n155 16.477
R23314 commonsourceibias.n245 commonsourceibias.n244 16.477
R23315 commonsourceibias.n252 commonsourceibias.n251 16.477
R23316 commonsourceibias.n392 commonsourceibias.n391 16.477
R23317 commonsourceibias.n399 commonsourceibias.n398 16.477
R23318 commonsourceibias.n445 commonsourceibias.n444 16.477
R23319 commonsourceibias.n333 commonsourceibias.n332 16.477
R23320 commonsourceibias.n527 commonsourceibias.n526 16.477
R23321 commonsourceibias.n534 commonsourceibias.n533 16.477
R23322 commonsourceibias.n77 commonsourceibias.n76 15.9852
R23323 commonsourceibias.n56 commonsourceibias.n27 15.9852
R23324 commonsourceibias.n170 commonsourceibias.n169 15.9852
R23325 commonsourceibias.n149 commonsourceibias.n120 15.9852
R23326 commonsourceibias.n238 commonsourceibias.n209 15.9852
R23327 commonsourceibias.n259 commonsourceibias.n258 15.9852
R23328 commonsourceibias.n385 commonsourceibias.n356 15.9852
R23329 commonsourceibias.n407 commonsourceibias.n406 15.9852
R23330 commonsourceibias.n453 commonsourceibias.n452 15.9852
R23331 commonsourceibias.n326 commonsourceibias.n297 15.9852
R23332 commonsourceibias.n520 commonsourceibias.n491 15.9852
R23333 commonsourceibias.n542 commonsourceibias.n541 15.9852
R23334 commonsourceibias.n91 commonsourceibias.n90 15.4934
R23335 commonsourceibias.n41 commonsourceibias.n40 15.4934
R23336 commonsourceibias.n184 commonsourceibias.n183 15.4934
R23337 commonsourceibias.n134 commonsourceibias.n133 15.4934
R23338 commonsourceibias.n223 commonsourceibias.n222 15.4934
R23339 commonsourceibias.n273 commonsourceibias.n272 15.4934
R23340 commonsourceibias.n370 commonsourceibias.n369 15.4934
R23341 commonsourceibias.n422 commonsourceibias.n421 15.4934
R23342 commonsourceibias.n468 commonsourceibias.n467 15.4934
R23343 commonsourceibias.n311 commonsourceibias.n310 15.4934
R23344 commonsourceibias.n505 commonsourceibias.n504 15.4934
R23345 commonsourceibias.n557 commonsourceibias.n556 15.4934
R23346 commonsourceibias.n102 commonsourceibias.n100 13.2663
R23347 commonsourceibias.n433 commonsourceibias.n431 13.2663
R23348 commonsourceibias.n568 commonsourceibias.n283 12.2777
R23349 commonsourceibias.n568 commonsourceibias.n567 10.3347
R23350 commonsourceibias.n159 commonsourceibias.n116 9.50363
R23351 commonsourceibias.n441 commonsourceibias.n440 9.50363
R23352 commonsourceibias.n92 commonsourceibias.n91 9.09948
R23353 commonsourceibias.n40 commonsourceibias.n39 9.09948
R23354 commonsourceibias.n185 commonsourceibias.n184 9.09948
R23355 commonsourceibias.n133 commonsourceibias.n132 9.09948
R23356 commonsourceibias.n222 commonsourceibias.n221 9.09948
R23357 commonsourceibias.n274 commonsourceibias.n273 9.09948
R23358 commonsourceibias.n369 commonsourceibias.n368 9.09948
R23359 commonsourceibias.n423 commonsourceibias.n422 9.09948
R23360 commonsourceibias.n469 commonsourceibias.n468 9.09948
R23361 commonsourceibias.n310 commonsourceibias.n309 9.09948
R23362 commonsourceibias.n504 commonsourceibias.n503 9.09948
R23363 commonsourceibias.n558 commonsourceibias.n557 9.09948
R23364 commonsourceibias.n283 commonsourceibias.n193 8.79261
R23365 commonsourceibias.n567 commonsourceibias.n477 8.79261
R23366 commonsourceibias.n78 commonsourceibias.n77 8.60764
R23367 commonsourceibias.n53 commonsourceibias.n27 8.60764
R23368 commonsourceibias.n171 commonsourceibias.n170 8.60764
R23369 commonsourceibias.n146 commonsourceibias.n120 8.60764
R23370 commonsourceibias.n235 commonsourceibias.n209 8.60764
R23371 commonsourceibias.n260 commonsourceibias.n259 8.60764
R23372 commonsourceibias.n382 commonsourceibias.n356 8.60764
R23373 commonsourceibias.n408 commonsourceibias.n407 8.60764
R23374 commonsourceibias.n454 commonsourceibias.n453 8.60764
R23375 commonsourceibias.n323 commonsourceibias.n297 8.60764
R23376 commonsourceibias.n517 commonsourceibias.n491 8.60764
R23377 commonsourceibias.n543 commonsourceibias.n542 8.60764
R23378 commonsourceibias.n69 commonsourceibias.n68 8.11581
R23379 commonsourceibias.n64 commonsourceibias.n63 8.11581
R23380 commonsourceibias.n162 commonsourceibias.n161 8.11581
R23381 commonsourceibias.n157 commonsourceibias.n156 8.11581
R23382 commonsourceibias.n246 commonsourceibias.n245 8.11581
R23383 commonsourceibias.n251 commonsourceibias.n250 8.11581
R23384 commonsourceibias.n393 commonsourceibias.n392 8.11581
R23385 commonsourceibias.n398 commonsourceibias.n397 8.11581
R23386 commonsourceibias.n444 commonsourceibias.n443 8.11581
R23387 commonsourceibias.n334 commonsourceibias.n333 8.11581
R23388 commonsourceibias.n528 commonsourceibias.n527 8.11581
R23389 commonsourceibias.n533 commonsourceibias.n532 8.11581
R23390 commonsourceibias.n83 commonsourceibias.n82 7.62397
R23391 commonsourceibias.n51 commonsourceibias.n29 7.62397
R23392 commonsourceibias.n176 commonsourceibias.n175 7.62397
R23393 commonsourceibias.n144 commonsourceibias.n122 7.62397
R23394 commonsourceibias.n233 commonsourceibias.n211 7.62397
R23395 commonsourceibias.n265 commonsourceibias.n264 7.62397
R23396 commonsourceibias.n380 commonsourceibias.n358 7.62397
R23397 commonsourceibias.n413 commonsourceibias.n412 7.62397
R23398 commonsourceibias.n459 commonsourceibias.n458 7.62397
R23399 commonsourceibias.n321 commonsourceibias.n299 7.62397
R23400 commonsourceibias.n515 commonsourceibias.n493 7.62397
R23401 commonsourceibias.n548 commonsourceibias.n547 7.62397
R23402 commonsourceibias.n97 commonsourceibias.n96 7.13213
R23403 commonsourceibias.n34 commonsourceibias.n33 7.13213
R23404 commonsourceibias.n190 commonsourceibias.n189 7.13213
R23405 commonsourceibias.n127 commonsourceibias.n126 7.13213
R23406 commonsourceibias.n216 commonsourceibias.n215 7.13213
R23407 commonsourceibias.n279 commonsourceibias.n278 7.13213
R23408 commonsourceibias.n363 commonsourceibias.n362 7.13213
R23409 commonsourceibias.n428 commonsourceibias.n427 7.13213
R23410 commonsourceibias.n474 commonsourceibias.n473 7.13213
R23411 commonsourceibias.n304 commonsourceibias.n303 7.13213
R23412 commonsourceibias.n498 commonsourceibias.n497 7.13213
R23413 commonsourceibias.n563 commonsourceibias.n562 7.13213
R23414 commonsourceibias.n283 commonsourceibias.n282 5.06534
R23415 commonsourceibias.n567 commonsourceibias.n566 5.06534
R23416 commonsourceibias commonsourceibias.n568 4.04308
R23417 commonsourceibias.n109 commonsourceibias.t13 2.82907
R23418 commonsourceibias.n109 commonsourceibias.t17 2.82907
R23419 commonsourceibias.n110 commonsourceibias.t31 2.82907
R23420 commonsourceibias.n110 commonsourceibias.t57 2.82907
R23421 commonsourceibias.n112 commonsourceibias.t43 2.82907
R23422 commonsourceibias.n112 commonsourceibias.t21 2.82907
R23423 commonsourceibias.n114 commonsourceibias.t7 2.82907
R23424 commonsourceibias.n114 commonsourceibias.t33 2.82907
R23425 commonsourceibias.n107 commonsourceibias.t19 2.82907
R23426 commonsourceibias.n107 commonsourceibias.t27 2.82907
R23427 commonsourceibias.n105 commonsourceibias.t29 2.82907
R23428 commonsourceibias.n105 commonsourceibias.t63 2.82907
R23429 commonsourceibias.n103 commonsourceibias.t39 2.82907
R23430 commonsourceibias.n103 commonsourceibias.t5 2.82907
R23431 commonsourceibias.n101 commonsourceibias.t61 2.82907
R23432 commonsourceibias.n101 commonsourceibias.t15 2.82907
R23433 commonsourceibias.n432 commonsourceibias.t35 2.82907
R23434 commonsourceibias.n432 commonsourceibias.t9 2.82907
R23435 commonsourceibias.n434 commonsourceibias.t23 2.82907
R23436 commonsourceibias.n434 commonsourceibias.t1 2.82907
R23437 commonsourceibias.n436 commonsourceibias.t11 2.82907
R23438 commonsourceibias.n436 commonsourceibias.t47 2.82907
R23439 commonsourceibias.n438 commonsourceibias.t45 2.82907
R23440 commonsourceibias.n438 commonsourceibias.t37 2.82907
R23441 commonsourceibias.n341 commonsourceibias.t51 2.82907
R23442 commonsourceibias.n341 commonsourceibias.t25 2.82907
R23443 commonsourceibias.n339 commonsourceibias.t41 2.82907
R23444 commonsourceibias.n339 commonsourceibias.t59 2.82907
R23445 commonsourceibias.n337 commonsourceibias.t3 2.82907
R23446 commonsourceibias.n337 commonsourceibias.t49 2.82907
R23447 commonsourceibias.n336 commonsourceibias.t55 2.82907
R23448 commonsourceibias.n336 commonsourceibias.t53 2.82907
R23449 commonsourceibias.n17 commonsourceibias.n15 0.738255
R23450 commonsourceibias.n46 commonsourceibias.n45 0.738255
R23451 commonsourceibias.n5 commonsourceibias.n3 0.738255
R23452 commonsourceibias.n139 commonsourceibias.n138 0.738255
R23453 commonsourceibias.n228 commonsourceibias.n227 0.738255
R23454 commonsourceibias.n199 commonsourceibias.n197 0.738255
R23455 commonsourceibias.n375 commonsourceibias.n374 0.738255
R23456 commonsourceibias.n415 commonsourceibias.n346 0.738255
R23457 commonsourceibias.n461 commonsourceibias.n287 0.738255
R23458 commonsourceibias.n316 commonsourceibias.n315 0.738255
R23459 commonsourceibias.n510 commonsourceibias.n509 0.738255
R23460 commonsourceibias.n550 commonsourceibias.n481 0.738255
R23461 commonsourceibias.n104 commonsourceibias.n102 0.573776
R23462 commonsourceibias.n106 commonsourceibias.n104 0.573776
R23463 commonsourceibias.n108 commonsourceibias.n106 0.573776
R23464 commonsourceibias.n115 commonsourceibias.n113 0.573776
R23465 commonsourceibias.n113 commonsourceibias.n111 0.573776
R23466 commonsourceibias.n340 commonsourceibias.n338 0.573776
R23467 commonsourceibias.n342 commonsourceibias.n340 0.573776
R23468 commonsourceibias.n439 commonsourceibias.n437 0.573776
R23469 commonsourceibias.n437 commonsourceibias.n435 0.573776
R23470 commonsourceibias.n435 commonsourceibias.n433 0.573776
R23471 commonsourceibias.n116 commonsourceibias.n108 0.287138
R23472 commonsourceibias.n116 commonsourceibias.n115 0.287138
R23473 commonsourceibias.n440 commonsourceibias.n342 0.287138
R23474 commonsourceibias.n440 commonsourceibias.n439 0.287138
R23475 commonsourceibias.n100 commonsourceibias.n12 0.285035
R23476 commonsourceibias.n193 commonsourceibias.n0 0.285035
R23477 commonsourceibias.n282 commonsourceibias.n194 0.285035
R23478 commonsourceibias.n431 commonsourceibias.n343 0.285035
R23479 commonsourceibias.n477 commonsourceibias.n284 0.285035
R23480 commonsourceibias.n566 commonsourceibias.n478 0.285035
R23481 commonsourceibias.n22 commonsourceibias.n20 0.246418
R23482 commonsourceibias.n58 commonsourceibias.n25 0.246418
R23483 commonsourceibias.n10 commonsourceibias.n8 0.246418
R23484 commonsourceibias.n151 commonsourceibias.n118 0.246418
R23485 commonsourceibias.n240 commonsourceibias.n207 0.246418
R23486 commonsourceibias.n204 commonsourceibias.n202 0.246418
R23487 commonsourceibias.n387 commonsourceibias.n354 0.246418
R23488 commonsourceibias.n400 commonsourceibias.n350 0.246418
R23489 commonsourceibias.n446 commonsourceibias.n291 0.246418
R23490 commonsourceibias.n328 commonsourceibias.n295 0.246418
R23491 commonsourceibias.n522 commonsourceibias.n489 0.246418
R23492 commonsourceibias.n535 commonsourceibias.n485 0.246418
R23493 commonsourceibias.n95 commonsourceibias.n12 0.189894
R23494 commonsourceibias.n95 commonsourceibias.n94 0.189894
R23495 commonsourceibias.n94 commonsourceibias.n93 0.189894
R23496 commonsourceibias.n93 commonsourceibias.n14 0.189894
R23497 commonsourceibias.n88 commonsourceibias.n14 0.189894
R23498 commonsourceibias.n88 commonsourceibias.n87 0.189894
R23499 commonsourceibias.n87 commonsourceibias.n86 0.189894
R23500 commonsourceibias.n86 commonsourceibias.n16 0.189894
R23501 commonsourceibias.n81 commonsourceibias.n16 0.189894
R23502 commonsourceibias.n81 commonsourceibias.n80 0.189894
R23503 commonsourceibias.n80 commonsourceibias.n79 0.189894
R23504 commonsourceibias.n79 commonsourceibias.n19 0.189894
R23505 commonsourceibias.n74 commonsourceibias.n19 0.189894
R23506 commonsourceibias.n74 commonsourceibias.n73 0.189894
R23507 commonsourceibias.n73 commonsourceibias.n72 0.189894
R23508 commonsourceibias.n72 commonsourceibias.n21 0.189894
R23509 commonsourceibias.n67 commonsourceibias.n21 0.189894
R23510 commonsourceibias.n67 commonsourceibias.n66 0.189894
R23511 commonsourceibias.n66 commonsourceibias.n65 0.189894
R23512 commonsourceibias.n65 commonsourceibias.n24 0.189894
R23513 commonsourceibias.n60 commonsourceibias.n24 0.189894
R23514 commonsourceibias.n60 commonsourceibias.n59 0.189894
R23515 commonsourceibias.n59 commonsourceibias.n26 0.189894
R23516 commonsourceibias.n55 commonsourceibias.n26 0.189894
R23517 commonsourceibias.n55 commonsourceibias.n54 0.189894
R23518 commonsourceibias.n54 commonsourceibias.n28 0.189894
R23519 commonsourceibias.n50 commonsourceibias.n28 0.189894
R23520 commonsourceibias.n50 commonsourceibias.n49 0.189894
R23521 commonsourceibias.n49 commonsourceibias.n30 0.189894
R23522 commonsourceibias.n44 commonsourceibias.n30 0.189894
R23523 commonsourceibias.n44 commonsourceibias.n43 0.189894
R23524 commonsourceibias.n43 commonsourceibias.n42 0.189894
R23525 commonsourceibias.n42 commonsourceibias.n32 0.189894
R23526 commonsourceibias.n37 commonsourceibias.n32 0.189894
R23527 commonsourceibias.n37 commonsourceibias.n36 0.189894
R23528 commonsourceibias.n158 commonsourceibias.n117 0.189894
R23529 commonsourceibias.n153 commonsourceibias.n117 0.189894
R23530 commonsourceibias.n153 commonsourceibias.n152 0.189894
R23531 commonsourceibias.n152 commonsourceibias.n119 0.189894
R23532 commonsourceibias.n148 commonsourceibias.n119 0.189894
R23533 commonsourceibias.n148 commonsourceibias.n147 0.189894
R23534 commonsourceibias.n147 commonsourceibias.n121 0.189894
R23535 commonsourceibias.n143 commonsourceibias.n121 0.189894
R23536 commonsourceibias.n143 commonsourceibias.n142 0.189894
R23537 commonsourceibias.n142 commonsourceibias.n123 0.189894
R23538 commonsourceibias.n137 commonsourceibias.n123 0.189894
R23539 commonsourceibias.n137 commonsourceibias.n136 0.189894
R23540 commonsourceibias.n136 commonsourceibias.n135 0.189894
R23541 commonsourceibias.n135 commonsourceibias.n125 0.189894
R23542 commonsourceibias.n130 commonsourceibias.n125 0.189894
R23543 commonsourceibias.n130 commonsourceibias.n129 0.189894
R23544 commonsourceibias.n188 commonsourceibias.n0 0.189894
R23545 commonsourceibias.n188 commonsourceibias.n187 0.189894
R23546 commonsourceibias.n187 commonsourceibias.n186 0.189894
R23547 commonsourceibias.n186 commonsourceibias.n2 0.189894
R23548 commonsourceibias.n181 commonsourceibias.n2 0.189894
R23549 commonsourceibias.n181 commonsourceibias.n180 0.189894
R23550 commonsourceibias.n180 commonsourceibias.n179 0.189894
R23551 commonsourceibias.n179 commonsourceibias.n4 0.189894
R23552 commonsourceibias.n174 commonsourceibias.n4 0.189894
R23553 commonsourceibias.n174 commonsourceibias.n173 0.189894
R23554 commonsourceibias.n173 commonsourceibias.n172 0.189894
R23555 commonsourceibias.n172 commonsourceibias.n7 0.189894
R23556 commonsourceibias.n167 commonsourceibias.n7 0.189894
R23557 commonsourceibias.n167 commonsourceibias.n166 0.189894
R23558 commonsourceibias.n166 commonsourceibias.n165 0.189894
R23559 commonsourceibias.n165 commonsourceibias.n9 0.189894
R23560 commonsourceibias.n160 commonsourceibias.n9 0.189894
R23561 commonsourceibias.n277 commonsourceibias.n194 0.189894
R23562 commonsourceibias.n277 commonsourceibias.n276 0.189894
R23563 commonsourceibias.n276 commonsourceibias.n275 0.189894
R23564 commonsourceibias.n275 commonsourceibias.n196 0.189894
R23565 commonsourceibias.n270 commonsourceibias.n196 0.189894
R23566 commonsourceibias.n270 commonsourceibias.n269 0.189894
R23567 commonsourceibias.n269 commonsourceibias.n268 0.189894
R23568 commonsourceibias.n268 commonsourceibias.n198 0.189894
R23569 commonsourceibias.n263 commonsourceibias.n198 0.189894
R23570 commonsourceibias.n263 commonsourceibias.n262 0.189894
R23571 commonsourceibias.n262 commonsourceibias.n261 0.189894
R23572 commonsourceibias.n261 commonsourceibias.n201 0.189894
R23573 commonsourceibias.n256 commonsourceibias.n201 0.189894
R23574 commonsourceibias.n256 commonsourceibias.n255 0.189894
R23575 commonsourceibias.n255 commonsourceibias.n254 0.189894
R23576 commonsourceibias.n254 commonsourceibias.n203 0.189894
R23577 commonsourceibias.n249 commonsourceibias.n203 0.189894
R23578 commonsourceibias.n249 commonsourceibias.n248 0.189894
R23579 commonsourceibias.n248 commonsourceibias.n247 0.189894
R23580 commonsourceibias.n247 commonsourceibias.n206 0.189894
R23581 commonsourceibias.n242 commonsourceibias.n206 0.189894
R23582 commonsourceibias.n242 commonsourceibias.n241 0.189894
R23583 commonsourceibias.n241 commonsourceibias.n208 0.189894
R23584 commonsourceibias.n237 commonsourceibias.n208 0.189894
R23585 commonsourceibias.n237 commonsourceibias.n236 0.189894
R23586 commonsourceibias.n236 commonsourceibias.n210 0.189894
R23587 commonsourceibias.n232 commonsourceibias.n210 0.189894
R23588 commonsourceibias.n232 commonsourceibias.n231 0.189894
R23589 commonsourceibias.n231 commonsourceibias.n212 0.189894
R23590 commonsourceibias.n226 commonsourceibias.n212 0.189894
R23591 commonsourceibias.n226 commonsourceibias.n225 0.189894
R23592 commonsourceibias.n225 commonsourceibias.n224 0.189894
R23593 commonsourceibias.n224 commonsourceibias.n214 0.189894
R23594 commonsourceibias.n219 commonsourceibias.n214 0.189894
R23595 commonsourceibias.n219 commonsourceibias.n218 0.189894
R23596 commonsourceibias.n366 commonsourceibias.n365 0.189894
R23597 commonsourceibias.n366 commonsourceibias.n361 0.189894
R23598 commonsourceibias.n371 commonsourceibias.n361 0.189894
R23599 commonsourceibias.n372 commonsourceibias.n371 0.189894
R23600 commonsourceibias.n373 commonsourceibias.n372 0.189894
R23601 commonsourceibias.n373 commonsourceibias.n359 0.189894
R23602 commonsourceibias.n378 commonsourceibias.n359 0.189894
R23603 commonsourceibias.n379 commonsourceibias.n378 0.189894
R23604 commonsourceibias.n379 commonsourceibias.n357 0.189894
R23605 commonsourceibias.n383 commonsourceibias.n357 0.189894
R23606 commonsourceibias.n384 commonsourceibias.n383 0.189894
R23607 commonsourceibias.n384 commonsourceibias.n355 0.189894
R23608 commonsourceibias.n388 commonsourceibias.n355 0.189894
R23609 commonsourceibias.n389 commonsourceibias.n388 0.189894
R23610 commonsourceibias.n389 commonsourceibias.n353 0.189894
R23611 commonsourceibias.n394 commonsourceibias.n353 0.189894
R23612 commonsourceibias.n395 commonsourceibias.n394 0.189894
R23613 commonsourceibias.n396 commonsourceibias.n395 0.189894
R23614 commonsourceibias.n396 commonsourceibias.n351 0.189894
R23615 commonsourceibias.n402 commonsourceibias.n351 0.189894
R23616 commonsourceibias.n403 commonsourceibias.n402 0.189894
R23617 commonsourceibias.n404 commonsourceibias.n403 0.189894
R23618 commonsourceibias.n404 commonsourceibias.n349 0.189894
R23619 commonsourceibias.n409 commonsourceibias.n349 0.189894
R23620 commonsourceibias.n410 commonsourceibias.n409 0.189894
R23621 commonsourceibias.n411 commonsourceibias.n410 0.189894
R23622 commonsourceibias.n411 commonsourceibias.n347 0.189894
R23623 commonsourceibias.n417 commonsourceibias.n347 0.189894
R23624 commonsourceibias.n418 commonsourceibias.n417 0.189894
R23625 commonsourceibias.n419 commonsourceibias.n418 0.189894
R23626 commonsourceibias.n419 commonsourceibias.n345 0.189894
R23627 commonsourceibias.n424 commonsourceibias.n345 0.189894
R23628 commonsourceibias.n425 commonsourceibias.n424 0.189894
R23629 commonsourceibias.n426 commonsourceibias.n425 0.189894
R23630 commonsourceibias.n426 commonsourceibias.n343 0.189894
R23631 commonsourceibias.n307 commonsourceibias.n306 0.189894
R23632 commonsourceibias.n307 commonsourceibias.n302 0.189894
R23633 commonsourceibias.n312 commonsourceibias.n302 0.189894
R23634 commonsourceibias.n313 commonsourceibias.n312 0.189894
R23635 commonsourceibias.n314 commonsourceibias.n313 0.189894
R23636 commonsourceibias.n314 commonsourceibias.n300 0.189894
R23637 commonsourceibias.n319 commonsourceibias.n300 0.189894
R23638 commonsourceibias.n320 commonsourceibias.n319 0.189894
R23639 commonsourceibias.n320 commonsourceibias.n298 0.189894
R23640 commonsourceibias.n324 commonsourceibias.n298 0.189894
R23641 commonsourceibias.n325 commonsourceibias.n324 0.189894
R23642 commonsourceibias.n325 commonsourceibias.n296 0.189894
R23643 commonsourceibias.n329 commonsourceibias.n296 0.189894
R23644 commonsourceibias.n330 commonsourceibias.n329 0.189894
R23645 commonsourceibias.n330 commonsourceibias.n294 0.189894
R23646 commonsourceibias.n335 commonsourceibias.n294 0.189894
R23647 commonsourceibias.n442 commonsourceibias.n292 0.189894
R23648 commonsourceibias.n448 commonsourceibias.n292 0.189894
R23649 commonsourceibias.n449 commonsourceibias.n448 0.189894
R23650 commonsourceibias.n450 commonsourceibias.n449 0.189894
R23651 commonsourceibias.n450 commonsourceibias.n290 0.189894
R23652 commonsourceibias.n455 commonsourceibias.n290 0.189894
R23653 commonsourceibias.n456 commonsourceibias.n455 0.189894
R23654 commonsourceibias.n457 commonsourceibias.n456 0.189894
R23655 commonsourceibias.n457 commonsourceibias.n288 0.189894
R23656 commonsourceibias.n463 commonsourceibias.n288 0.189894
R23657 commonsourceibias.n464 commonsourceibias.n463 0.189894
R23658 commonsourceibias.n465 commonsourceibias.n464 0.189894
R23659 commonsourceibias.n465 commonsourceibias.n286 0.189894
R23660 commonsourceibias.n470 commonsourceibias.n286 0.189894
R23661 commonsourceibias.n471 commonsourceibias.n470 0.189894
R23662 commonsourceibias.n472 commonsourceibias.n471 0.189894
R23663 commonsourceibias.n472 commonsourceibias.n284 0.189894
R23664 commonsourceibias.n501 commonsourceibias.n500 0.189894
R23665 commonsourceibias.n501 commonsourceibias.n496 0.189894
R23666 commonsourceibias.n506 commonsourceibias.n496 0.189894
R23667 commonsourceibias.n507 commonsourceibias.n506 0.189894
R23668 commonsourceibias.n508 commonsourceibias.n507 0.189894
R23669 commonsourceibias.n508 commonsourceibias.n494 0.189894
R23670 commonsourceibias.n513 commonsourceibias.n494 0.189894
R23671 commonsourceibias.n514 commonsourceibias.n513 0.189894
R23672 commonsourceibias.n514 commonsourceibias.n492 0.189894
R23673 commonsourceibias.n518 commonsourceibias.n492 0.189894
R23674 commonsourceibias.n519 commonsourceibias.n518 0.189894
R23675 commonsourceibias.n519 commonsourceibias.n490 0.189894
R23676 commonsourceibias.n523 commonsourceibias.n490 0.189894
R23677 commonsourceibias.n524 commonsourceibias.n523 0.189894
R23678 commonsourceibias.n524 commonsourceibias.n488 0.189894
R23679 commonsourceibias.n529 commonsourceibias.n488 0.189894
R23680 commonsourceibias.n530 commonsourceibias.n529 0.189894
R23681 commonsourceibias.n531 commonsourceibias.n530 0.189894
R23682 commonsourceibias.n531 commonsourceibias.n486 0.189894
R23683 commonsourceibias.n537 commonsourceibias.n486 0.189894
R23684 commonsourceibias.n538 commonsourceibias.n537 0.189894
R23685 commonsourceibias.n539 commonsourceibias.n538 0.189894
R23686 commonsourceibias.n539 commonsourceibias.n484 0.189894
R23687 commonsourceibias.n544 commonsourceibias.n484 0.189894
R23688 commonsourceibias.n545 commonsourceibias.n544 0.189894
R23689 commonsourceibias.n546 commonsourceibias.n545 0.189894
R23690 commonsourceibias.n546 commonsourceibias.n482 0.189894
R23691 commonsourceibias.n552 commonsourceibias.n482 0.189894
R23692 commonsourceibias.n553 commonsourceibias.n552 0.189894
R23693 commonsourceibias.n554 commonsourceibias.n553 0.189894
R23694 commonsourceibias.n554 commonsourceibias.n480 0.189894
R23695 commonsourceibias.n559 commonsourceibias.n480 0.189894
R23696 commonsourceibias.n560 commonsourceibias.n559 0.189894
R23697 commonsourceibias.n561 commonsourceibias.n560 0.189894
R23698 commonsourceibias.n561 commonsourceibias.n478 0.189894
R23699 commonsourceibias.n159 commonsourceibias.n158 0.170955
R23700 commonsourceibias.n160 commonsourceibias.n159 0.170955
R23701 commonsourceibias.n441 commonsourceibias.n335 0.170955
R23702 commonsourceibias.n442 commonsourceibias.n441 0.170955
R23703 diffpairibias.n0 diffpairibias.t27 436.822
R23704 diffpairibias.n27 diffpairibias.t24 435.479
R23705 diffpairibias.n26 diffpairibias.t21 435.479
R23706 diffpairibias.n25 diffpairibias.t22 435.479
R23707 diffpairibias.n24 diffpairibias.t26 435.479
R23708 diffpairibias.n23 diffpairibias.t20 435.479
R23709 diffpairibias.n0 diffpairibias.t23 435.479
R23710 diffpairibias.n1 diffpairibias.t28 435.479
R23711 diffpairibias.n2 diffpairibias.t25 435.479
R23712 diffpairibias.n3 diffpairibias.t29 435.479
R23713 diffpairibias.n13 diffpairibias.t14 377.536
R23714 diffpairibias.n13 diffpairibias.t0 376.193
R23715 diffpairibias.n14 diffpairibias.t10 376.193
R23716 diffpairibias.n15 diffpairibias.t12 376.193
R23717 diffpairibias.n16 diffpairibias.t6 376.193
R23718 diffpairibias.n17 diffpairibias.t2 376.193
R23719 diffpairibias.n18 diffpairibias.t16 376.193
R23720 diffpairibias.n19 diffpairibias.t4 376.193
R23721 diffpairibias.n20 diffpairibias.t18 376.193
R23722 diffpairibias.n21 diffpairibias.t8 376.193
R23723 diffpairibias.n4 diffpairibias.t15 113.368
R23724 diffpairibias.n4 diffpairibias.t1 112.698
R23725 diffpairibias.n5 diffpairibias.t11 112.698
R23726 diffpairibias.n6 diffpairibias.t13 112.698
R23727 diffpairibias.n7 diffpairibias.t7 112.698
R23728 diffpairibias.n8 diffpairibias.t3 112.698
R23729 diffpairibias.n9 diffpairibias.t17 112.698
R23730 diffpairibias.n10 diffpairibias.t5 112.698
R23731 diffpairibias.n11 diffpairibias.t19 112.698
R23732 diffpairibias.n12 diffpairibias.t9 112.698
R23733 diffpairibias.n22 diffpairibias.n21 4.77242
R23734 diffpairibias.n22 diffpairibias.n12 4.30807
R23735 diffpairibias.n23 diffpairibias.n22 4.13945
R23736 diffpairibias.n21 diffpairibias.n20 1.34352
R23737 diffpairibias.n20 diffpairibias.n19 1.34352
R23738 diffpairibias.n19 diffpairibias.n18 1.34352
R23739 diffpairibias.n18 diffpairibias.n17 1.34352
R23740 diffpairibias.n17 diffpairibias.n16 1.34352
R23741 diffpairibias.n16 diffpairibias.n15 1.34352
R23742 diffpairibias.n15 diffpairibias.n14 1.34352
R23743 diffpairibias.n14 diffpairibias.n13 1.34352
R23744 diffpairibias.n3 diffpairibias.n2 1.34352
R23745 diffpairibias.n2 diffpairibias.n1 1.34352
R23746 diffpairibias.n1 diffpairibias.n0 1.34352
R23747 diffpairibias.n24 diffpairibias.n23 1.34352
R23748 diffpairibias.n25 diffpairibias.n24 1.34352
R23749 diffpairibias.n26 diffpairibias.n25 1.34352
R23750 diffpairibias.n27 diffpairibias.n26 1.34352
R23751 diffpairibias.n28 diffpairibias.n27 0.862419
R23752 diffpairibias diffpairibias.n28 0.684875
R23753 diffpairibias.n12 diffpairibias.n11 0.672012
R23754 diffpairibias.n11 diffpairibias.n10 0.672012
R23755 diffpairibias.n10 diffpairibias.n9 0.672012
R23756 diffpairibias.n9 diffpairibias.n8 0.672012
R23757 diffpairibias.n8 diffpairibias.n7 0.672012
R23758 diffpairibias.n7 diffpairibias.n6 0.672012
R23759 diffpairibias.n6 diffpairibias.n5 0.672012
R23760 diffpairibias.n5 diffpairibias.n4 0.672012
R23761 diffpairibias.n28 diffpairibias.n3 0.190907
R23762 output.n41 output.n15 289.615
R23763 output.n72 output.n46 289.615
R23764 output.n104 output.n78 289.615
R23765 output.n136 output.n110 289.615
R23766 output.n77 output.n45 197.26
R23767 output.n77 output.n76 196.298
R23768 output.n109 output.n108 196.298
R23769 output.n141 output.n140 196.298
R23770 output.n42 output.n41 185
R23771 output.n40 output.n39 185
R23772 output.n19 output.n18 185
R23773 output.n34 output.n33 185
R23774 output.n32 output.n31 185
R23775 output.n23 output.n22 185
R23776 output.n26 output.n25 185
R23777 output.n73 output.n72 185
R23778 output.n71 output.n70 185
R23779 output.n50 output.n49 185
R23780 output.n65 output.n64 185
R23781 output.n63 output.n62 185
R23782 output.n54 output.n53 185
R23783 output.n57 output.n56 185
R23784 output.n105 output.n104 185
R23785 output.n103 output.n102 185
R23786 output.n82 output.n81 185
R23787 output.n97 output.n96 185
R23788 output.n95 output.n94 185
R23789 output.n86 output.n85 185
R23790 output.n89 output.n88 185
R23791 output.n137 output.n136 185
R23792 output.n135 output.n134 185
R23793 output.n114 output.n113 185
R23794 output.n129 output.n128 185
R23795 output.n127 output.n126 185
R23796 output.n118 output.n117 185
R23797 output.n121 output.n120 185
R23798 output.t2 output.n24 147.661
R23799 output.t19 output.n55 147.661
R23800 output.t0 output.n87 147.661
R23801 output.t1 output.n119 147.661
R23802 output.n41 output.n40 104.615
R23803 output.n40 output.n18 104.615
R23804 output.n33 output.n18 104.615
R23805 output.n33 output.n32 104.615
R23806 output.n32 output.n22 104.615
R23807 output.n25 output.n22 104.615
R23808 output.n72 output.n71 104.615
R23809 output.n71 output.n49 104.615
R23810 output.n64 output.n49 104.615
R23811 output.n64 output.n63 104.615
R23812 output.n63 output.n53 104.615
R23813 output.n56 output.n53 104.615
R23814 output.n104 output.n103 104.615
R23815 output.n103 output.n81 104.615
R23816 output.n96 output.n81 104.615
R23817 output.n96 output.n95 104.615
R23818 output.n95 output.n85 104.615
R23819 output.n88 output.n85 104.615
R23820 output.n136 output.n135 104.615
R23821 output.n135 output.n113 104.615
R23822 output.n128 output.n113 104.615
R23823 output.n128 output.n127 104.615
R23824 output.n127 output.n117 104.615
R23825 output.n120 output.n117 104.615
R23826 output.n1 output.t15 77.056
R23827 output.n14 output.t16 76.6694
R23828 output.n1 output.n0 72.7095
R23829 output.n3 output.n2 72.7095
R23830 output.n5 output.n4 72.7095
R23831 output.n7 output.n6 72.7095
R23832 output.n9 output.n8 72.7095
R23833 output.n11 output.n10 72.7095
R23834 output.n13 output.n12 72.7095
R23835 output.n25 output.t2 52.3082
R23836 output.n56 output.t19 52.3082
R23837 output.n88 output.t0 52.3082
R23838 output.n120 output.t1 52.3082
R23839 output.n26 output.n24 15.6674
R23840 output.n57 output.n55 15.6674
R23841 output.n89 output.n87 15.6674
R23842 output.n121 output.n119 15.6674
R23843 output.n27 output.n23 12.8005
R23844 output.n58 output.n54 12.8005
R23845 output.n90 output.n86 12.8005
R23846 output.n122 output.n118 12.8005
R23847 output.n31 output.n30 12.0247
R23848 output.n62 output.n61 12.0247
R23849 output.n94 output.n93 12.0247
R23850 output.n126 output.n125 12.0247
R23851 output.n34 output.n21 11.249
R23852 output.n65 output.n52 11.249
R23853 output.n97 output.n84 11.249
R23854 output.n129 output.n116 11.249
R23855 output.n35 output.n19 10.4732
R23856 output.n66 output.n50 10.4732
R23857 output.n98 output.n82 10.4732
R23858 output.n130 output.n114 10.4732
R23859 output.n39 output.n38 9.69747
R23860 output.n70 output.n69 9.69747
R23861 output.n102 output.n101 9.69747
R23862 output.n134 output.n133 9.69747
R23863 output.n45 output.n44 9.45567
R23864 output.n76 output.n75 9.45567
R23865 output.n108 output.n107 9.45567
R23866 output.n140 output.n139 9.45567
R23867 output.n44 output.n43 9.3005
R23868 output.n17 output.n16 9.3005
R23869 output.n38 output.n37 9.3005
R23870 output.n36 output.n35 9.3005
R23871 output.n21 output.n20 9.3005
R23872 output.n30 output.n29 9.3005
R23873 output.n28 output.n27 9.3005
R23874 output.n75 output.n74 9.3005
R23875 output.n48 output.n47 9.3005
R23876 output.n69 output.n68 9.3005
R23877 output.n67 output.n66 9.3005
R23878 output.n52 output.n51 9.3005
R23879 output.n61 output.n60 9.3005
R23880 output.n59 output.n58 9.3005
R23881 output.n107 output.n106 9.3005
R23882 output.n80 output.n79 9.3005
R23883 output.n101 output.n100 9.3005
R23884 output.n99 output.n98 9.3005
R23885 output.n84 output.n83 9.3005
R23886 output.n93 output.n92 9.3005
R23887 output.n91 output.n90 9.3005
R23888 output.n139 output.n138 9.3005
R23889 output.n112 output.n111 9.3005
R23890 output.n133 output.n132 9.3005
R23891 output.n131 output.n130 9.3005
R23892 output.n116 output.n115 9.3005
R23893 output.n125 output.n124 9.3005
R23894 output.n123 output.n122 9.3005
R23895 output.n42 output.n17 8.92171
R23896 output.n73 output.n48 8.92171
R23897 output.n105 output.n80 8.92171
R23898 output.n137 output.n112 8.92171
R23899 output output.n141 8.15037
R23900 output.n43 output.n15 8.14595
R23901 output.n74 output.n46 8.14595
R23902 output.n106 output.n78 8.14595
R23903 output.n138 output.n110 8.14595
R23904 output.n45 output.n15 5.81868
R23905 output.n76 output.n46 5.81868
R23906 output.n108 output.n78 5.81868
R23907 output.n140 output.n110 5.81868
R23908 output.n43 output.n42 5.04292
R23909 output.n74 output.n73 5.04292
R23910 output.n106 output.n105 5.04292
R23911 output.n138 output.n137 5.04292
R23912 output.n28 output.n24 4.38594
R23913 output.n59 output.n55 4.38594
R23914 output.n91 output.n87 4.38594
R23915 output.n123 output.n119 4.38594
R23916 output.n39 output.n17 4.26717
R23917 output.n70 output.n48 4.26717
R23918 output.n102 output.n80 4.26717
R23919 output.n134 output.n112 4.26717
R23920 output.n0 output.t5 3.9605
R23921 output.n0 output.t9 3.9605
R23922 output.n2 output.t12 3.9605
R23923 output.n2 output.t17 3.9605
R23924 output.n4 output.t18 3.9605
R23925 output.n4 output.t7 3.9605
R23926 output.n6 output.t11 3.9605
R23927 output.n6 output.t3 3.9605
R23928 output.n8 output.t6 3.9605
R23929 output.n8 output.t4 3.9605
R23930 output.n10 output.t10 3.9605
R23931 output.n10 output.t13 3.9605
R23932 output.n12 output.t14 3.9605
R23933 output.n12 output.t8 3.9605
R23934 output.n38 output.n19 3.49141
R23935 output.n69 output.n50 3.49141
R23936 output.n101 output.n82 3.49141
R23937 output.n133 output.n114 3.49141
R23938 output.n35 output.n34 2.71565
R23939 output.n66 output.n65 2.71565
R23940 output.n98 output.n97 2.71565
R23941 output.n130 output.n129 2.71565
R23942 output.n31 output.n21 1.93989
R23943 output.n62 output.n52 1.93989
R23944 output.n94 output.n84 1.93989
R23945 output.n126 output.n116 1.93989
R23946 output.n30 output.n23 1.16414
R23947 output.n61 output.n54 1.16414
R23948 output.n93 output.n86 1.16414
R23949 output.n125 output.n118 1.16414
R23950 output.n141 output.n109 0.962709
R23951 output.n109 output.n77 0.962709
R23952 output.n27 output.n26 0.388379
R23953 output.n58 output.n57 0.388379
R23954 output.n90 output.n89 0.388379
R23955 output.n122 output.n121 0.388379
R23956 output.n14 output.n13 0.387128
R23957 output.n13 output.n11 0.387128
R23958 output.n11 output.n9 0.387128
R23959 output.n9 output.n7 0.387128
R23960 output.n7 output.n5 0.387128
R23961 output.n5 output.n3 0.387128
R23962 output.n3 output.n1 0.387128
R23963 output.n44 output.n16 0.155672
R23964 output.n37 output.n16 0.155672
R23965 output.n37 output.n36 0.155672
R23966 output.n36 output.n20 0.155672
R23967 output.n29 output.n20 0.155672
R23968 output.n29 output.n28 0.155672
R23969 output.n75 output.n47 0.155672
R23970 output.n68 output.n47 0.155672
R23971 output.n68 output.n67 0.155672
R23972 output.n67 output.n51 0.155672
R23973 output.n60 output.n51 0.155672
R23974 output.n60 output.n59 0.155672
R23975 output.n107 output.n79 0.155672
R23976 output.n100 output.n79 0.155672
R23977 output.n100 output.n99 0.155672
R23978 output.n99 output.n83 0.155672
R23979 output.n92 output.n83 0.155672
R23980 output.n92 output.n91 0.155672
R23981 output.n139 output.n111 0.155672
R23982 output.n132 output.n111 0.155672
R23983 output.n132 output.n131 0.155672
R23984 output.n131 output.n115 0.155672
R23985 output.n124 output.n115 0.155672
R23986 output.n124 output.n123 0.155672
R23987 output output.n14 0.126227
R23988 a_n2982_8322.n12 a_n2982_8322.t27 74.6477
R23989 a_n2982_8322.n1 a_n2982_8322.t6 74.6477
R23990 a_n2982_8322.n28 a_n2982_8322.t21 74.6474
R23991 a_n2982_8322.n20 a_n2982_8322.t1 74.2899
R23992 a_n2982_8322.n13 a_n2982_8322.t25 74.2899
R23993 a_n2982_8322.n14 a_n2982_8322.t28 74.2899
R23994 a_n2982_8322.n17 a_n2982_8322.t29 74.2899
R23995 a_n2982_8322.n10 a_n2982_8322.t0 74.2899
R23996 a_n2982_8322.n28 a_n2982_8322.n27 70.6783
R23997 a_n2982_8322.n26 a_n2982_8322.n25 70.6783
R23998 a_n2982_8322.n24 a_n2982_8322.n23 70.6783
R23999 a_n2982_8322.n22 a_n2982_8322.n21 70.6783
R24000 a_n2982_8322.n12 a_n2982_8322.n11 70.6783
R24001 a_n2982_8322.n16 a_n2982_8322.n15 70.6783
R24002 a_n2982_8322.n1 a_n2982_8322.n0 70.6783
R24003 a_n2982_8322.n3 a_n2982_8322.n2 70.6783
R24004 a_n2982_8322.n5 a_n2982_8322.n4 70.6783
R24005 a_n2982_8322.n7 a_n2982_8322.n6 70.6783
R24006 a_n2982_8322.n9 a_n2982_8322.n8 70.6783
R24007 a_n2982_8322.n30 a_n2982_8322.n29 70.6782
R24008 a_n2982_8322.n18 a_n2982_8322.n10 24.9022
R24009 a_n2982_8322.n19 a_n2982_8322.t32 9.79689
R24010 a_n2982_8322.n18 a_n2982_8322.n17 8.38735
R24011 a_n2982_8322.n20 a_n2982_8322.n19 6.90998
R24012 a_n2982_8322.n19 a_n2982_8322.n18 5.3452
R24013 a_n2982_8322.n27 a_n2982_8322.t14 3.61217
R24014 a_n2982_8322.n27 a_n2982_8322.t10 3.61217
R24015 a_n2982_8322.n25 a_n2982_8322.t20 3.61217
R24016 a_n2982_8322.n25 a_n2982_8322.t8 3.61217
R24017 a_n2982_8322.n23 a_n2982_8322.t5 3.61217
R24018 a_n2982_8322.n23 a_n2982_8322.t4 3.61217
R24019 a_n2982_8322.n21 a_n2982_8322.t18 3.61217
R24020 a_n2982_8322.n21 a_n2982_8322.t17 3.61217
R24021 a_n2982_8322.n11 a_n2982_8322.t31 3.61217
R24022 a_n2982_8322.n11 a_n2982_8322.t30 3.61217
R24023 a_n2982_8322.n15 a_n2982_8322.t26 3.61217
R24024 a_n2982_8322.n15 a_n2982_8322.t24 3.61217
R24025 a_n2982_8322.n0 a_n2982_8322.t19 3.61217
R24026 a_n2982_8322.n0 a_n2982_8322.t15 3.61217
R24027 a_n2982_8322.n2 a_n2982_8322.t22 3.61217
R24028 a_n2982_8322.n2 a_n2982_8322.t12 3.61217
R24029 a_n2982_8322.n4 a_n2982_8322.t3 3.61217
R24030 a_n2982_8322.n4 a_n2982_8322.t2 3.61217
R24031 a_n2982_8322.n6 a_n2982_8322.t16 3.61217
R24032 a_n2982_8322.n6 a_n2982_8322.t9 3.61217
R24033 a_n2982_8322.n8 a_n2982_8322.t13 3.61217
R24034 a_n2982_8322.n8 a_n2982_8322.t11 3.61217
R24035 a_n2982_8322.n30 a_n2982_8322.t7 3.61217
R24036 a_n2982_8322.t23 a_n2982_8322.n30 3.61217
R24037 a_n2982_8322.n17 a_n2982_8322.n16 0.358259
R24038 a_n2982_8322.n16 a_n2982_8322.n14 0.358259
R24039 a_n2982_8322.n13 a_n2982_8322.n12 0.358259
R24040 a_n2982_8322.n10 a_n2982_8322.n9 0.358259
R24041 a_n2982_8322.n9 a_n2982_8322.n7 0.358259
R24042 a_n2982_8322.n7 a_n2982_8322.n5 0.358259
R24043 a_n2982_8322.n5 a_n2982_8322.n3 0.358259
R24044 a_n2982_8322.n3 a_n2982_8322.n1 0.358259
R24045 a_n2982_8322.n22 a_n2982_8322.n20 0.358259
R24046 a_n2982_8322.n24 a_n2982_8322.n22 0.358259
R24047 a_n2982_8322.n26 a_n2982_8322.n24 0.358259
R24048 a_n2982_8322.n29 a_n2982_8322.n26 0.358259
R24049 a_n2982_8322.n29 a_n2982_8322.n28 0.358259
R24050 a_n2982_8322.n14 a_n2982_8322.n13 0.101793
R24051 a_n2982_8322.t34 a_n2982_8322.t37 0.0788333
R24052 a_n2982_8322.t33 a_n2982_8322.t35 0.0788333
R24053 a_n2982_8322.t32 a_n2982_8322.t36 0.0788333
R24054 a_n2982_8322.t33 a_n2982_8322.t34 0.0318333
R24055 a_n2982_8322.t32 a_n2982_8322.t35 0.0318333
R24056 a_n2982_8322.t37 a_n2982_8322.t35 0.0318333
R24057 a_n2982_8322.t36 a_n2982_8322.t33 0.0318333
R24058 outputibias.n27 outputibias.n1 289.615
R24059 outputibias.n58 outputibias.n32 289.615
R24060 outputibias.n90 outputibias.n64 289.615
R24061 outputibias.n122 outputibias.n96 289.615
R24062 outputibias.n28 outputibias.n27 185
R24063 outputibias.n26 outputibias.n25 185
R24064 outputibias.n5 outputibias.n4 185
R24065 outputibias.n20 outputibias.n19 185
R24066 outputibias.n18 outputibias.n17 185
R24067 outputibias.n9 outputibias.n8 185
R24068 outputibias.n12 outputibias.n11 185
R24069 outputibias.n59 outputibias.n58 185
R24070 outputibias.n57 outputibias.n56 185
R24071 outputibias.n36 outputibias.n35 185
R24072 outputibias.n51 outputibias.n50 185
R24073 outputibias.n49 outputibias.n48 185
R24074 outputibias.n40 outputibias.n39 185
R24075 outputibias.n43 outputibias.n42 185
R24076 outputibias.n91 outputibias.n90 185
R24077 outputibias.n89 outputibias.n88 185
R24078 outputibias.n68 outputibias.n67 185
R24079 outputibias.n83 outputibias.n82 185
R24080 outputibias.n81 outputibias.n80 185
R24081 outputibias.n72 outputibias.n71 185
R24082 outputibias.n75 outputibias.n74 185
R24083 outputibias.n123 outputibias.n122 185
R24084 outputibias.n121 outputibias.n120 185
R24085 outputibias.n100 outputibias.n99 185
R24086 outputibias.n115 outputibias.n114 185
R24087 outputibias.n113 outputibias.n112 185
R24088 outputibias.n104 outputibias.n103 185
R24089 outputibias.n107 outputibias.n106 185
R24090 outputibias.n0 outputibias.t8 178.945
R24091 outputibias.n133 outputibias.t11 177.018
R24092 outputibias.n132 outputibias.t9 177.018
R24093 outputibias.n0 outputibias.t10 177.018
R24094 outputibias.t5 outputibias.n10 147.661
R24095 outputibias.t7 outputibias.n41 147.661
R24096 outputibias.t1 outputibias.n73 147.661
R24097 outputibias.t3 outputibias.n105 147.661
R24098 outputibias.n128 outputibias.t4 132.363
R24099 outputibias.n128 outputibias.t6 130.436
R24100 outputibias.n129 outputibias.t0 130.436
R24101 outputibias.n130 outputibias.t2 130.436
R24102 outputibias.n27 outputibias.n26 104.615
R24103 outputibias.n26 outputibias.n4 104.615
R24104 outputibias.n19 outputibias.n4 104.615
R24105 outputibias.n19 outputibias.n18 104.615
R24106 outputibias.n18 outputibias.n8 104.615
R24107 outputibias.n11 outputibias.n8 104.615
R24108 outputibias.n58 outputibias.n57 104.615
R24109 outputibias.n57 outputibias.n35 104.615
R24110 outputibias.n50 outputibias.n35 104.615
R24111 outputibias.n50 outputibias.n49 104.615
R24112 outputibias.n49 outputibias.n39 104.615
R24113 outputibias.n42 outputibias.n39 104.615
R24114 outputibias.n90 outputibias.n89 104.615
R24115 outputibias.n89 outputibias.n67 104.615
R24116 outputibias.n82 outputibias.n67 104.615
R24117 outputibias.n82 outputibias.n81 104.615
R24118 outputibias.n81 outputibias.n71 104.615
R24119 outputibias.n74 outputibias.n71 104.615
R24120 outputibias.n122 outputibias.n121 104.615
R24121 outputibias.n121 outputibias.n99 104.615
R24122 outputibias.n114 outputibias.n99 104.615
R24123 outputibias.n114 outputibias.n113 104.615
R24124 outputibias.n113 outputibias.n103 104.615
R24125 outputibias.n106 outputibias.n103 104.615
R24126 outputibias.n63 outputibias.n31 95.6354
R24127 outputibias.n63 outputibias.n62 94.6732
R24128 outputibias.n95 outputibias.n94 94.6732
R24129 outputibias.n127 outputibias.n126 94.6732
R24130 outputibias.n11 outputibias.t5 52.3082
R24131 outputibias.n42 outputibias.t7 52.3082
R24132 outputibias.n74 outputibias.t1 52.3082
R24133 outputibias.n106 outputibias.t3 52.3082
R24134 outputibias.n12 outputibias.n10 15.6674
R24135 outputibias.n43 outputibias.n41 15.6674
R24136 outputibias.n75 outputibias.n73 15.6674
R24137 outputibias.n107 outputibias.n105 15.6674
R24138 outputibias.n13 outputibias.n9 12.8005
R24139 outputibias.n44 outputibias.n40 12.8005
R24140 outputibias.n76 outputibias.n72 12.8005
R24141 outputibias.n108 outputibias.n104 12.8005
R24142 outputibias.n17 outputibias.n16 12.0247
R24143 outputibias.n48 outputibias.n47 12.0247
R24144 outputibias.n80 outputibias.n79 12.0247
R24145 outputibias.n112 outputibias.n111 12.0247
R24146 outputibias.n20 outputibias.n7 11.249
R24147 outputibias.n51 outputibias.n38 11.249
R24148 outputibias.n83 outputibias.n70 11.249
R24149 outputibias.n115 outputibias.n102 11.249
R24150 outputibias.n21 outputibias.n5 10.4732
R24151 outputibias.n52 outputibias.n36 10.4732
R24152 outputibias.n84 outputibias.n68 10.4732
R24153 outputibias.n116 outputibias.n100 10.4732
R24154 outputibias.n25 outputibias.n24 9.69747
R24155 outputibias.n56 outputibias.n55 9.69747
R24156 outputibias.n88 outputibias.n87 9.69747
R24157 outputibias.n120 outputibias.n119 9.69747
R24158 outputibias.n31 outputibias.n30 9.45567
R24159 outputibias.n62 outputibias.n61 9.45567
R24160 outputibias.n94 outputibias.n93 9.45567
R24161 outputibias.n126 outputibias.n125 9.45567
R24162 outputibias.n30 outputibias.n29 9.3005
R24163 outputibias.n3 outputibias.n2 9.3005
R24164 outputibias.n24 outputibias.n23 9.3005
R24165 outputibias.n22 outputibias.n21 9.3005
R24166 outputibias.n7 outputibias.n6 9.3005
R24167 outputibias.n16 outputibias.n15 9.3005
R24168 outputibias.n14 outputibias.n13 9.3005
R24169 outputibias.n61 outputibias.n60 9.3005
R24170 outputibias.n34 outputibias.n33 9.3005
R24171 outputibias.n55 outputibias.n54 9.3005
R24172 outputibias.n53 outputibias.n52 9.3005
R24173 outputibias.n38 outputibias.n37 9.3005
R24174 outputibias.n47 outputibias.n46 9.3005
R24175 outputibias.n45 outputibias.n44 9.3005
R24176 outputibias.n93 outputibias.n92 9.3005
R24177 outputibias.n66 outputibias.n65 9.3005
R24178 outputibias.n87 outputibias.n86 9.3005
R24179 outputibias.n85 outputibias.n84 9.3005
R24180 outputibias.n70 outputibias.n69 9.3005
R24181 outputibias.n79 outputibias.n78 9.3005
R24182 outputibias.n77 outputibias.n76 9.3005
R24183 outputibias.n125 outputibias.n124 9.3005
R24184 outputibias.n98 outputibias.n97 9.3005
R24185 outputibias.n119 outputibias.n118 9.3005
R24186 outputibias.n117 outputibias.n116 9.3005
R24187 outputibias.n102 outputibias.n101 9.3005
R24188 outputibias.n111 outputibias.n110 9.3005
R24189 outputibias.n109 outputibias.n108 9.3005
R24190 outputibias.n28 outputibias.n3 8.92171
R24191 outputibias.n59 outputibias.n34 8.92171
R24192 outputibias.n91 outputibias.n66 8.92171
R24193 outputibias.n123 outputibias.n98 8.92171
R24194 outputibias.n29 outputibias.n1 8.14595
R24195 outputibias.n60 outputibias.n32 8.14595
R24196 outputibias.n92 outputibias.n64 8.14595
R24197 outputibias.n124 outputibias.n96 8.14595
R24198 outputibias.n31 outputibias.n1 5.81868
R24199 outputibias.n62 outputibias.n32 5.81868
R24200 outputibias.n94 outputibias.n64 5.81868
R24201 outputibias.n126 outputibias.n96 5.81868
R24202 outputibias.n131 outputibias.n130 5.20947
R24203 outputibias.n29 outputibias.n28 5.04292
R24204 outputibias.n60 outputibias.n59 5.04292
R24205 outputibias.n92 outputibias.n91 5.04292
R24206 outputibias.n124 outputibias.n123 5.04292
R24207 outputibias.n131 outputibias.n127 4.42209
R24208 outputibias.n14 outputibias.n10 4.38594
R24209 outputibias.n45 outputibias.n41 4.38594
R24210 outputibias.n77 outputibias.n73 4.38594
R24211 outputibias.n109 outputibias.n105 4.38594
R24212 outputibias.n132 outputibias.n131 4.28454
R24213 outputibias.n25 outputibias.n3 4.26717
R24214 outputibias.n56 outputibias.n34 4.26717
R24215 outputibias.n88 outputibias.n66 4.26717
R24216 outputibias.n120 outputibias.n98 4.26717
R24217 outputibias.n24 outputibias.n5 3.49141
R24218 outputibias.n55 outputibias.n36 3.49141
R24219 outputibias.n87 outputibias.n68 3.49141
R24220 outputibias.n119 outputibias.n100 3.49141
R24221 outputibias.n21 outputibias.n20 2.71565
R24222 outputibias.n52 outputibias.n51 2.71565
R24223 outputibias.n84 outputibias.n83 2.71565
R24224 outputibias.n116 outputibias.n115 2.71565
R24225 outputibias.n17 outputibias.n7 1.93989
R24226 outputibias.n48 outputibias.n38 1.93989
R24227 outputibias.n80 outputibias.n70 1.93989
R24228 outputibias.n112 outputibias.n102 1.93989
R24229 outputibias.n130 outputibias.n129 1.9266
R24230 outputibias.n129 outputibias.n128 1.9266
R24231 outputibias.n133 outputibias.n132 1.92658
R24232 outputibias.n134 outputibias.n133 1.29913
R24233 outputibias.n16 outputibias.n9 1.16414
R24234 outputibias.n47 outputibias.n40 1.16414
R24235 outputibias.n79 outputibias.n72 1.16414
R24236 outputibias.n111 outputibias.n104 1.16414
R24237 outputibias.n127 outputibias.n95 0.962709
R24238 outputibias.n95 outputibias.n63 0.962709
R24239 outputibias.n13 outputibias.n12 0.388379
R24240 outputibias.n44 outputibias.n43 0.388379
R24241 outputibias.n76 outputibias.n75 0.388379
R24242 outputibias.n108 outputibias.n107 0.388379
R24243 outputibias.n134 outputibias.n0 0.337251
R24244 outputibias outputibias.n134 0.302375
R24245 outputibias.n30 outputibias.n2 0.155672
R24246 outputibias.n23 outputibias.n2 0.155672
R24247 outputibias.n23 outputibias.n22 0.155672
R24248 outputibias.n22 outputibias.n6 0.155672
R24249 outputibias.n15 outputibias.n6 0.155672
R24250 outputibias.n15 outputibias.n14 0.155672
R24251 outputibias.n61 outputibias.n33 0.155672
R24252 outputibias.n54 outputibias.n33 0.155672
R24253 outputibias.n54 outputibias.n53 0.155672
R24254 outputibias.n53 outputibias.n37 0.155672
R24255 outputibias.n46 outputibias.n37 0.155672
R24256 outputibias.n46 outputibias.n45 0.155672
R24257 outputibias.n93 outputibias.n65 0.155672
R24258 outputibias.n86 outputibias.n65 0.155672
R24259 outputibias.n86 outputibias.n85 0.155672
R24260 outputibias.n85 outputibias.n69 0.155672
R24261 outputibias.n78 outputibias.n69 0.155672
R24262 outputibias.n78 outputibias.n77 0.155672
R24263 outputibias.n125 outputibias.n97 0.155672
R24264 outputibias.n118 outputibias.n97 0.155672
R24265 outputibias.n118 outputibias.n117 0.155672
R24266 outputibias.n117 outputibias.n101 0.155672
R24267 outputibias.n110 outputibias.n101 0.155672
R24268 outputibias.n110 outputibias.n109 0.155672
C0 output outputibias 2.34152f
C1 vdd output 7.23429f
C2 CSoutput output 6.13571f
C3 CSoutput outputibias 0.032386f
C4 vdd CSoutput 0.117223p
C5 minus diffpairibias 4.33e-19
C6 commonsourceibias output 0.006808f
C7 vdd plus 0.095585f
C8 CSoutput minus 2.89653f
C9 plus diffpairibias 4.56e-19
C10 commonsourceibias outputibias 0.003832f
C11 CSoutput plus 0.892085f
C12 vdd commonsourceibias 0.004218f
C13 commonsourceibias diffpairibias 0.052527f
C14 minus plus 9.92364f
C15 CSoutput commonsourceibias 37.4715f
C16 minus commonsourceibias 0.337549f
C17 plus commonsourceibias 0.283677f
C18 diffpairibias gnd 59.99123f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.150736p
C22 plus gnd 36.888f
C23 minus gnd 30.042679f
C24 CSoutput gnd 0.102106p
C25 vdd gnd 0.512126p
C26 outputibias.t10 gnd 0.11477f
C27 outputibias.t8 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t5 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t7 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t1 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t3 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t2 gnd 0.108319f
C161 outputibias.t0 gnd 0.108319f
C162 outputibias.t6 gnd 0.108319f
C163 outputibias.t4 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t9 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t11 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 a_n2982_8322.t7 gnd 0.100113f
C174 a_n2982_8322.t35 gnd 20.7695f
C175 a_n2982_8322.t37 gnd 20.6238f
C176 a_n2982_8322.t34 gnd 20.6238f
C177 a_n2982_8322.t33 gnd 20.7695f
C178 a_n2982_8322.t36 gnd 20.6238f
C179 a_n2982_8322.t32 gnd 29.446598f
C180 a_n2982_8322.t6 gnd 0.937411f
C181 a_n2982_8322.t19 gnd 0.100113f
C182 a_n2982_8322.t15 gnd 0.100113f
C183 a_n2982_8322.n0 gnd 0.705199f
C184 a_n2982_8322.n1 gnd 0.787956f
C185 a_n2982_8322.t22 gnd 0.100113f
C186 a_n2982_8322.t12 gnd 0.100113f
C187 a_n2982_8322.n2 gnd 0.705199f
C188 a_n2982_8322.n3 gnd 0.40035f
C189 a_n2982_8322.t3 gnd 0.100113f
C190 a_n2982_8322.t2 gnd 0.100113f
C191 a_n2982_8322.n4 gnd 0.705199f
C192 a_n2982_8322.n5 gnd 0.40035f
C193 a_n2982_8322.t16 gnd 0.100113f
C194 a_n2982_8322.t9 gnd 0.100113f
C195 a_n2982_8322.n6 gnd 0.705199f
C196 a_n2982_8322.n7 gnd 0.40035f
C197 a_n2982_8322.t13 gnd 0.100113f
C198 a_n2982_8322.t11 gnd 0.100113f
C199 a_n2982_8322.n8 gnd 0.705199f
C200 a_n2982_8322.n9 gnd 0.40035f
C201 a_n2982_8322.t0 gnd 0.935545f
C202 a_n2982_8322.n10 gnd 1.87053f
C203 a_n2982_8322.t27 gnd 0.937411f
C204 a_n2982_8322.t31 gnd 0.100113f
C205 a_n2982_8322.t30 gnd 0.100113f
C206 a_n2982_8322.n11 gnd 0.705199f
C207 a_n2982_8322.n12 gnd 0.787956f
C208 a_n2982_8322.t25 gnd 0.935545f
C209 a_n2982_8322.n13 gnd 0.39651f
C210 a_n2982_8322.t28 gnd 0.935545f
C211 a_n2982_8322.n14 gnd 0.39651f
C212 a_n2982_8322.t26 gnd 0.100113f
C213 a_n2982_8322.t24 gnd 0.100113f
C214 a_n2982_8322.n15 gnd 0.705199f
C215 a_n2982_8322.n16 gnd 0.40035f
C216 a_n2982_8322.t29 gnd 0.935545f
C217 a_n2982_8322.n17 gnd 1.47073f
C218 a_n2982_8322.n18 gnd 2.35026f
C219 a_n2982_8322.n19 gnd 3.52538f
C220 a_n2982_8322.t1 gnd 0.935545f
C221 a_n2982_8322.n20 gnd 1.11095f
C222 a_n2982_8322.t18 gnd 0.100113f
C223 a_n2982_8322.t17 gnd 0.100113f
C224 a_n2982_8322.n21 gnd 0.705199f
C225 a_n2982_8322.n22 gnd 0.40035f
C226 a_n2982_8322.t5 gnd 0.100113f
C227 a_n2982_8322.t4 gnd 0.100113f
C228 a_n2982_8322.n23 gnd 0.705199f
C229 a_n2982_8322.n24 gnd 0.40035f
C230 a_n2982_8322.t20 gnd 0.100113f
C231 a_n2982_8322.t8 gnd 0.100113f
C232 a_n2982_8322.n25 gnd 0.705199f
C233 a_n2982_8322.n26 gnd 0.40035f
C234 a_n2982_8322.t21 gnd 0.937409f
C235 a_n2982_8322.t14 gnd 0.100113f
C236 a_n2982_8322.t10 gnd 0.100113f
C237 a_n2982_8322.n27 gnd 0.705199f
C238 a_n2982_8322.n28 gnd 0.787958f
C239 a_n2982_8322.n29 gnd 0.400348f
C240 a_n2982_8322.n30 gnd 0.705201f
C241 a_n2982_8322.t23 gnd 0.100113f
C242 output.t15 gnd 0.464308f
C243 output.t5 gnd 0.044422f
C244 output.t9 gnd 0.044422f
C245 output.n0 gnd 0.364624f
C246 output.n1 gnd 0.614102f
C247 output.t12 gnd 0.044422f
C248 output.t17 gnd 0.044422f
C249 output.n2 gnd 0.364624f
C250 output.n3 gnd 0.350265f
C251 output.t18 gnd 0.044422f
C252 output.t7 gnd 0.044422f
C253 output.n4 gnd 0.364624f
C254 output.n5 gnd 0.350265f
C255 output.t11 gnd 0.044422f
C256 output.t3 gnd 0.044422f
C257 output.n6 gnd 0.364624f
C258 output.n7 gnd 0.350265f
C259 output.t6 gnd 0.044422f
C260 output.t4 gnd 0.044422f
C261 output.n8 gnd 0.364624f
C262 output.n9 gnd 0.350265f
C263 output.t10 gnd 0.044422f
C264 output.t13 gnd 0.044422f
C265 output.n10 gnd 0.364624f
C266 output.n11 gnd 0.350265f
C267 output.t14 gnd 0.044422f
C268 output.t8 gnd 0.044422f
C269 output.n12 gnd 0.364624f
C270 output.n13 gnd 0.350265f
C271 output.t16 gnd 0.462979f
C272 output.n14 gnd 0.28994f
C273 output.n15 gnd 0.015803f
C274 output.n16 gnd 0.011243f
C275 output.n17 gnd 0.006041f
C276 output.n18 gnd 0.01428f
C277 output.n19 gnd 0.006397f
C278 output.n20 gnd 0.011243f
C279 output.n21 gnd 0.006041f
C280 output.n22 gnd 0.01428f
C281 output.n23 gnd 0.006397f
C282 output.n24 gnd 0.048111f
C283 output.t2 gnd 0.023274f
C284 output.n25 gnd 0.01071f
C285 output.n26 gnd 0.008435f
C286 output.n27 gnd 0.006041f
C287 output.n28 gnd 0.267512f
C288 output.n29 gnd 0.011243f
C289 output.n30 gnd 0.006041f
C290 output.n31 gnd 0.006397f
C291 output.n32 gnd 0.01428f
C292 output.n33 gnd 0.01428f
C293 output.n34 gnd 0.006397f
C294 output.n35 gnd 0.006041f
C295 output.n36 gnd 0.011243f
C296 output.n37 gnd 0.011243f
C297 output.n38 gnd 0.006041f
C298 output.n39 gnd 0.006397f
C299 output.n40 gnd 0.01428f
C300 output.n41 gnd 0.030913f
C301 output.n42 gnd 0.006397f
C302 output.n43 gnd 0.006041f
C303 output.n44 gnd 0.025987f
C304 output.n45 gnd 0.097665f
C305 output.n46 gnd 0.015803f
C306 output.n47 gnd 0.011243f
C307 output.n48 gnd 0.006041f
C308 output.n49 gnd 0.01428f
C309 output.n50 gnd 0.006397f
C310 output.n51 gnd 0.011243f
C311 output.n52 gnd 0.006041f
C312 output.n53 gnd 0.01428f
C313 output.n54 gnd 0.006397f
C314 output.n55 gnd 0.048111f
C315 output.t19 gnd 0.023274f
C316 output.n56 gnd 0.01071f
C317 output.n57 gnd 0.008435f
C318 output.n58 gnd 0.006041f
C319 output.n59 gnd 0.267512f
C320 output.n60 gnd 0.011243f
C321 output.n61 gnd 0.006041f
C322 output.n62 gnd 0.006397f
C323 output.n63 gnd 0.01428f
C324 output.n64 gnd 0.01428f
C325 output.n65 gnd 0.006397f
C326 output.n66 gnd 0.006041f
C327 output.n67 gnd 0.011243f
C328 output.n68 gnd 0.011243f
C329 output.n69 gnd 0.006041f
C330 output.n70 gnd 0.006397f
C331 output.n71 gnd 0.01428f
C332 output.n72 gnd 0.030913f
C333 output.n73 gnd 0.006397f
C334 output.n74 gnd 0.006041f
C335 output.n75 gnd 0.025987f
C336 output.n76 gnd 0.09306f
C337 output.n77 gnd 1.65264f
C338 output.n78 gnd 0.015803f
C339 output.n79 gnd 0.011243f
C340 output.n80 gnd 0.006041f
C341 output.n81 gnd 0.01428f
C342 output.n82 gnd 0.006397f
C343 output.n83 gnd 0.011243f
C344 output.n84 gnd 0.006041f
C345 output.n85 gnd 0.01428f
C346 output.n86 gnd 0.006397f
C347 output.n87 gnd 0.048111f
C348 output.t0 gnd 0.023274f
C349 output.n88 gnd 0.01071f
C350 output.n89 gnd 0.008435f
C351 output.n90 gnd 0.006041f
C352 output.n91 gnd 0.267512f
C353 output.n92 gnd 0.011243f
C354 output.n93 gnd 0.006041f
C355 output.n94 gnd 0.006397f
C356 output.n95 gnd 0.01428f
C357 output.n96 gnd 0.01428f
C358 output.n97 gnd 0.006397f
C359 output.n98 gnd 0.006041f
C360 output.n99 gnd 0.011243f
C361 output.n100 gnd 0.011243f
C362 output.n101 gnd 0.006041f
C363 output.n102 gnd 0.006397f
C364 output.n103 gnd 0.01428f
C365 output.n104 gnd 0.030913f
C366 output.n105 gnd 0.006397f
C367 output.n106 gnd 0.006041f
C368 output.n107 gnd 0.025987f
C369 output.n108 gnd 0.09306f
C370 output.n109 gnd 0.713089f
C371 output.n110 gnd 0.015803f
C372 output.n111 gnd 0.011243f
C373 output.n112 gnd 0.006041f
C374 output.n113 gnd 0.01428f
C375 output.n114 gnd 0.006397f
C376 output.n115 gnd 0.011243f
C377 output.n116 gnd 0.006041f
C378 output.n117 gnd 0.01428f
C379 output.n118 gnd 0.006397f
C380 output.n119 gnd 0.048111f
C381 output.t1 gnd 0.023274f
C382 output.n120 gnd 0.01071f
C383 output.n121 gnd 0.008435f
C384 output.n122 gnd 0.006041f
C385 output.n123 gnd 0.267512f
C386 output.n124 gnd 0.011243f
C387 output.n125 gnd 0.006041f
C388 output.n126 gnd 0.006397f
C389 output.n127 gnd 0.01428f
C390 output.n128 gnd 0.01428f
C391 output.n129 gnd 0.006397f
C392 output.n130 gnd 0.006041f
C393 output.n131 gnd 0.011243f
C394 output.n132 gnd 0.011243f
C395 output.n133 gnd 0.006041f
C396 output.n134 gnd 0.006397f
C397 output.n135 gnd 0.01428f
C398 output.n136 gnd 0.030913f
C399 output.n137 gnd 0.006397f
C400 output.n138 gnd 0.006041f
C401 output.n139 gnd 0.025987f
C402 output.n140 gnd 0.09306f
C403 output.n141 gnd 1.67353f
C404 diffpairibias.t27 gnd 0.090128f
C405 diffpairibias.t23 gnd 0.08996f
C406 diffpairibias.n0 gnd 0.105991f
C407 diffpairibias.t28 gnd 0.08996f
C408 diffpairibias.n1 gnd 0.051736f
C409 diffpairibias.t25 gnd 0.08996f
C410 diffpairibias.n2 gnd 0.051736f
C411 diffpairibias.t29 gnd 0.08996f
C412 diffpairibias.n3 gnd 0.041084f
C413 diffpairibias.t15 gnd 0.086371f
C414 diffpairibias.t1 gnd 0.085993f
C415 diffpairibias.n4 gnd 0.13579f
C416 diffpairibias.t11 gnd 0.085993f
C417 diffpairibias.n5 gnd 0.072463f
C418 diffpairibias.t13 gnd 0.085993f
C419 diffpairibias.n6 gnd 0.072463f
C420 diffpairibias.t7 gnd 0.085993f
C421 diffpairibias.n7 gnd 0.072463f
C422 diffpairibias.t3 gnd 0.085993f
C423 diffpairibias.n8 gnd 0.072463f
C424 diffpairibias.t17 gnd 0.085993f
C425 diffpairibias.n9 gnd 0.072463f
C426 diffpairibias.t5 gnd 0.085993f
C427 diffpairibias.n10 gnd 0.072463f
C428 diffpairibias.t19 gnd 0.085993f
C429 diffpairibias.n11 gnd 0.072463f
C430 diffpairibias.t9 gnd 0.085993f
C431 diffpairibias.n12 gnd 0.102883f
C432 diffpairibias.t14 gnd 0.086899f
C433 diffpairibias.t0 gnd 0.086748f
C434 diffpairibias.n13 gnd 0.094648f
C435 diffpairibias.t10 gnd 0.086748f
C436 diffpairibias.n14 gnd 0.052262f
C437 diffpairibias.t12 gnd 0.086748f
C438 diffpairibias.n15 gnd 0.052262f
C439 diffpairibias.t6 gnd 0.086748f
C440 diffpairibias.n16 gnd 0.052262f
C441 diffpairibias.t2 gnd 0.086748f
C442 diffpairibias.n17 gnd 0.052262f
C443 diffpairibias.t16 gnd 0.086748f
C444 diffpairibias.n18 gnd 0.052262f
C445 diffpairibias.t4 gnd 0.086748f
C446 diffpairibias.n19 gnd 0.052262f
C447 diffpairibias.t18 gnd 0.086748f
C448 diffpairibias.n20 gnd 0.052262f
C449 diffpairibias.t8 gnd 0.086748f
C450 diffpairibias.n21 gnd 0.061849f
C451 diffpairibias.n22 gnd 0.233513f
C452 diffpairibias.t20 gnd 0.08996f
C453 diffpairibias.n23 gnd 0.051747f
C454 diffpairibias.t26 gnd 0.08996f
C455 diffpairibias.n24 gnd 0.051736f
C456 diffpairibias.t22 gnd 0.08996f
C457 diffpairibias.n25 gnd 0.051736f
C458 diffpairibias.t21 gnd 0.08996f
C459 diffpairibias.n26 gnd 0.051736f
C460 diffpairibias.t24 gnd 0.08996f
C461 diffpairibias.n27 gnd 0.04729f
C462 diffpairibias.n28 gnd 0.047711f
C463 commonsourceibias.n0 gnd 0.010571f
C464 commonsourceibias.t92 gnd 0.160069f
C465 commonsourceibias.t106 gnd 0.148006f
C466 commonsourceibias.n1 gnd 0.006439f
C467 commonsourceibias.n2 gnd 0.007922f
C468 commonsourceibias.t119 gnd 0.148006f
C469 commonsourceibias.n3 gnd 0.008036f
C470 commonsourceibias.n4 gnd 0.007922f
C471 commonsourceibias.t84 gnd 0.148006f
C472 commonsourceibias.n5 gnd 0.059054f
C473 commonsourceibias.t100 gnd 0.148006f
C474 commonsourceibias.n6 gnd 0.006408f
C475 commonsourceibias.n7 gnd 0.007922f
C476 commonsourceibias.t114 gnd 0.148006f
C477 commonsourceibias.n8 gnd 0.007648f
C478 commonsourceibias.n9 gnd 0.007922f
C479 commonsourceibias.t80 gnd 0.148006f
C480 commonsourceibias.n10 gnd 0.059054f
C481 commonsourceibias.t76 gnd 0.148006f
C482 commonsourceibias.n11 gnd 0.006398f
C483 commonsourceibias.n12 gnd 0.010571f
C484 commonsourceibias.t60 gnd 0.160069f
C485 commonsourceibias.t14 gnd 0.148006f
C486 commonsourceibias.n13 gnd 0.006439f
C487 commonsourceibias.n14 gnd 0.007922f
C488 commonsourceibias.t38 gnd 0.148006f
C489 commonsourceibias.n15 gnd 0.008036f
C490 commonsourceibias.n16 gnd 0.007922f
C491 commonsourceibias.t4 gnd 0.148006f
C492 commonsourceibias.n17 gnd 0.059054f
C493 commonsourceibias.t28 gnd 0.148006f
C494 commonsourceibias.n18 gnd 0.006408f
C495 commonsourceibias.n19 gnd 0.007922f
C496 commonsourceibias.t62 gnd 0.148006f
C497 commonsourceibias.n20 gnd 0.007648f
C498 commonsourceibias.n21 gnd 0.007922f
C499 commonsourceibias.t18 gnd 0.148006f
C500 commonsourceibias.n22 gnd 0.059054f
C501 commonsourceibias.t26 gnd 0.148006f
C502 commonsourceibias.n23 gnd 0.006398f
C503 commonsourceibias.n24 gnd 0.007922f
C504 commonsourceibias.t6 gnd 0.148006f
C505 commonsourceibias.t32 gnd 0.148006f
C506 commonsourceibias.n25 gnd 0.059054f
C507 commonsourceibias.n26 gnd 0.007922f
C508 commonsourceibias.t42 gnd 0.148006f
C509 commonsourceibias.n27 gnd 0.059054f
C510 commonsourceibias.n28 gnd 0.007922f
C511 commonsourceibias.t20 gnd 0.148006f
C512 commonsourceibias.n29 gnd 0.059054f
C513 commonsourceibias.n30 gnd 0.007922f
C514 commonsourceibias.t30 gnd 0.148006f
C515 commonsourceibias.n31 gnd 0.009005f
C516 commonsourceibias.n32 gnd 0.007922f
C517 commonsourceibias.t56 gnd 0.148006f
C518 commonsourceibias.n33 gnd 0.010649f
C519 commonsourceibias.t16 gnd 0.164876f
C520 commonsourceibias.t12 gnd 0.148006f
C521 commonsourceibias.n34 gnd 0.065802f
C522 commonsourceibias.n35 gnd 0.070497f
C523 commonsourceibias.n36 gnd 0.03372f
C524 commonsourceibias.n37 gnd 0.007922f
C525 commonsourceibias.n38 gnd 0.006439f
C526 commonsourceibias.n39 gnd 0.010916f
C527 commonsourceibias.n40 gnd 0.059054f
C528 commonsourceibias.n41 gnd 0.010963f
C529 commonsourceibias.n42 gnd 0.007922f
C530 commonsourceibias.n43 gnd 0.007922f
C531 commonsourceibias.n44 gnd 0.007922f
C532 commonsourceibias.n45 gnd 0.008036f
C533 commonsourceibias.n46 gnd 0.059054f
C534 commonsourceibias.n47 gnd 0.009764f
C535 commonsourceibias.n48 gnd 0.010802f
C536 commonsourceibias.n49 gnd 0.007922f
C537 commonsourceibias.n50 gnd 0.007922f
C538 commonsourceibias.n51 gnd 0.010731f
C539 commonsourceibias.n52 gnd 0.006408f
C540 commonsourceibias.n53 gnd 0.010864f
C541 commonsourceibias.n54 gnd 0.007922f
C542 commonsourceibias.n55 gnd 0.007922f
C543 commonsourceibias.n56 gnd 0.010931f
C544 commonsourceibias.n57 gnd 0.009425f
C545 commonsourceibias.n58 gnd 0.007648f
C546 commonsourceibias.n59 gnd 0.007922f
C547 commonsourceibias.n60 gnd 0.007922f
C548 commonsourceibias.n61 gnd 0.00969f
C549 commonsourceibias.n62 gnd 0.010876f
C550 commonsourceibias.n63 gnd 0.059054f
C551 commonsourceibias.n64 gnd 0.010803f
C552 commonsourceibias.n65 gnd 0.007922f
C553 commonsourceibias.n66 gnd 0.007922f
C554 commonsourceibias.n67 gnd 0.007922f
C555 commonsourceibias.n68 gnd 0.010803f
C556 commonsourceibias.n69 gnd 0.059054f
C557 commonsourceibias.n70 gnd 0.010876f
C558 commonsourceibias.n71 gnd 0.00969f
C559 commonsourceibias.n72 gnd 0.007922f
C560 commonsourceibias.n73 gnd 0.007922f
C561 commonsourceibias.n74 gnd 0.007922f
C562 commonsourceibias.n75 gnd 0.009425f
C563 commonsourceibias.n76 gnd 0.010931f
C564 commonsourceibias.n77 gnd 0.059054f
C565 commonsourceibias.n78 gnd 0.010864f
C566 commonsourceibias.n79 gnd 0.007922f
C567 commonsourceibias.n80 gnd 0.007922f
C568 commonsourceibias.n81 gnd 0.007922f
C569 commonsourceibias.n82 gnd 0.010731f
C570 commonsourceibias.n83 gnd 0.059054f
C571 commonsourceibias.n84 gnd 0.010802f
C572 commonsourceibias.n85 gnd 0.009764f
C573 commonsourceibias.n86 gnd 0.007922f
C574 commonsourceibias.n87 gnd 0.007922f
C575 commonsourceibias.n88 gnd 0.007922f
C576 commonsourceibias.n89 gnd 0.009005f
C577 commonsourceibias.n90 gnd 0.010963f
C578 commonsourceibias.n91 gnd 0.059054f
C579 commonsourceibias.n92 gnd 0.010916f
C580 commonsourceibias.n93 gnd 0.007922f
C581 commonsourceibias.n94 gnd 0.007922f
C582 commonsourceibias.n95 gnd 0.007922f
C583 commonsourceibias.n96 gnd 0.010649f
C584 commonsourceibias.n97 gnd 0.059054f
C585 commonsourceibias.n98 gnd 0.010674f
C586 commonsourceibias.n99 gnd 0.071211f
C587 commonsourceibias.n100 gnd 0.079625f
C588 commonsourceibias.t61 gnd 0.017095f
C589 commonsourceibias.t15 gnd 0.017095f
C590 commonsourceibias.n101 gnd 0.151055f
C591 commonsourceibias.n102 gnd 0.130846f
C592 commonsourceibias.t39 gnd 0.017095f
C593 commonsourceibias.t5 gnd 0.017095f
C594 commonsourceibias.n103 gnd 0.151055f
C595 commonsourceibias.n104 gnd 0.069385f
C596 commonsourceibias.t29 gnd 0.017095f
C597 commonsourceibias.t63 gnd 0.017095f
C598 commonsourceibias.n105 gnd 0.151055f
C599 commonsourceibias.n106 gnd 0.069385f
C600 commonsourceibias.t19 gnd 0.017095f
C601 commonsourceibias.t27 gnd 0.017095f
C602 commonsourceibias.n107 gnd 0.151055f
C603 commonsourceibias.n108 gnd 0.057968f
C604 commonsourceibias.t13 gnd 0.017095f
C605 commonsourceibias.t17 gnd 0.017095f
C606 commonsourceibias.n109 gnd 0.15156f
C607 commonsourceibias.t31 gnd 0.017095f
C608 commonsourceibias.t57 gnd 0.017095f
C609 commonsourceibias.n110 gnd 0.151055f
C610 commonsourceibias.n111 gnd 0.140755f
C611 commonsourceibias.t43 gnd 0.017095f
C612 commonsourceibias.t21 gnd 0.017095f
C613 commonsourceibias.n112 gnd 0.151055f
C614 commonsourceibias.n113 gnd 0.069385f
C615 commonsourceibias.t7 gnd 0.017095f
C616 commonsourceibias.t33 gnd 0.017095f
C617 commonsourceibias.n114 gnd 0.151055f
C618 commonsourceibias.n115 gnd 0.057968f
C619 commonsourceibias.n116 gnd 0.070193f
C620 commonsourceibias.n117 gnd 0.007922f
C621 commonsourceibias.t105 gnd 0.148006f
C622 commonsourceibias.t121 gnd 0.148006f
C623 commonsourceibias.n118 gnd 0.059054f
C624 commonsourceibias.n119 gnd 0.007922f
C625 commonsourceibias.t71 gnd 0.148006f
C626 commonsourceibias.n120 gnd 0.059054f
C627 commonsourceibias.n121 gnd 0.007922f
C628 commonsourceibias.t99 gnd 0.148006f
C629 commonsourceibias.n122 gnd 0.059054f
C630 commonsourceibias.n123 gnd 0.007922f
C631 commonsourceibias.t95 gnd 0.148006f
C632 commonsourceibias.n124 gnd 0.009005f
C633 commonsourceibias.n125 gnd 0.007922f
C634 commonsourceibias.t109 gnd 0.148006f
C635 commonsourceibias.n126 gnd 0.010649f
C636 commonsourceibias.t85 gnd 0.164876f
C637 commonsourceibias.t89 gnd 0.148006f
C638 commonsourceibias.n127 gnd 0.065802f
C639 commonsourceibias.n128 gnd 0.070497f
C640 commonsourceibias.n129 gnd 0.03372f
C641 commonsourceibias.n130 gnd 0.007922f
C642 commonsourceibias.n131 gnd 0.006439f
C643 commonsourceibias.n132 gnd 0.010916f
C644 commonsourceibias.n133 gnd 0.059054f
C645 commonsourceibias.n134 gnd 0.010963f
C646 commonsourceibias.n135 gnd 0.007922f
C647 commonsourceibias.n136 gnd 0.007922f
C648 commonsourceibias.n137 gnd 0.007922f
C649 commonsourceibias.n138 gnd 0.008036f
C650 commonsourceibias.n139 gnd 0.059054f
C651 commonsourceibias.n140 gnd 0.009764f
C652 commonsourceibias.n141 gnd 0.010802f
C653 commonsourceibias.n142 gnd 0.007922f
C654 commonsourceibias.n143 gnd 0.007922f
C655 commonsourceibias.n144 gnd 0.010731f
C656 commonsourceibias.n145 gnd 0.006408f
C657 commonsourceibias.n146 gnd 0.010864f
C658 commonsourceibias.n147 gnd 0.007922f
C659 commonsourceibias.n148 gnd 0.007922f
C660 commonsourceibias.n149 gnd 0.010931f
C661 commonsourceibias.n150 gnd 0.009425f
C662 commonsourceibias.n151 gnd 0.007648f
C663 commonsourceibias.n152 gnd 0.007922f
C664 commonsourceibias.n153 gnd 0.007922f
C665 commonsourceibias.n154 gnd 0.00969f
C666 commonsourceibias.n155 gnd 0.010876f
C667 commonsourceibias.n156 gnd 0.059054f
C668 commonsourceibias.n157 gnd 0.010803f
C669 commonsourceibias.n158 gnd 0.007884f
C670 commonsourceibias.n159 gnd 0.057266f
C671 commonsourceibias.n160 gnd 0.007884f
C672 commonsourceibias.n161 gnd 0.010803f
C673 commonsourceibias.n162 gnd 0.059054f
C674 commonsourceibias.n163 gnd 0.010876f
C675 commonsourceibias.n164 gnd 0.00969f
C676 commonsourceibias.n165 gnd 0.007922f
C677 commonsourceibias.n166 gnd 0.007922f
C678 commonsourceibias.n167 gnd 0.007922f
C679 commonsourceibias.n168 gnd 0.009425f
C680 commonsourceibias.n169 gnd 0.010931f
C681 commonsourceibias.n170 gnd 0.059054f
C682 commonsourceibias.n171 gnd 0.010864f
C683 commonsourceibias.n172 gnd 0.007922f
C684 commonsourceibias.n173 gnd 0.007922f
C685 commonsourceibias.n174 gnd 0.007922f
C686 commonsourceibias.n175 gnd 0.010731f
C687 commonsourceibias.n176 gnd 0.059054f
C688 commonsourceibias.n177 gnd 0.010802f
C689 commonsourceibias.n178 gnd 0.009764f
C690 commonsourceibias.n179 gnd 0.007922f
C691 commonsourceibias.n180 gnd 0.007922f
C692 commonsourceibias.n181 gnd 0.007922f
C693 commonsourceibias.n182 gnd 0.009005f
C694 commonsourceibias.n183 gnd 0.010963f
C695 commonsourceibias.n184 gnd 0.059054f
C696 commonsourceibias.n185 gnd 0.010916f
C697 commonsourceibias.n186 gnd 0.007922f
C698 commonsourceibias.n187 gnd 0.007922f
C699 commonsourceibias.n188 gnd 0.007922f
C700 commonsourceibias.n189 gnd 0.010649f
C701 commonsourceibias.n190 gnd 0.059054f
C702 commonsourceibias.n191 gnd 0.010674f
C703 commonsourceibias.n192 gnd 0.071211f
C704 commonsourceibias.n193 gnd 0.047027f
C705 commonsourceibias.n194 gnd 0.010571f
C706 commonsourceibias.t94 gnd 0.148006f
C707 commonsourceibias.n195 gnd 0.006439f
C708 commonsourceibias.n196 gnd 0.007922f
C709 commonsourceibias.t107 gnd 0.148006f
C710 commonsourceibias.n197 gnd 0.008036f
C711 commonsourceibias.n198 gnd 0.007922f
C712 commonsourceibias.t74 gnd 0.148006f
C713 commonsourceibias.n199 gnd 0.059054f
C714 commonsourceibias.t87 gnd 0.148006f
C715 commonsourceibias.n200 gnd 0.006408f
C716 commonsourceibias.n201 gnd 0.007922f
C717 commonsourceibias.t101 gnd 0.148006f
C718 commonsourceibias.n202 gnd 0.007648f
C719 commonsourceibias.n203 gnd 0.007922f
C720 commonsourceibias.t70 gnd 0.148006f
C721 commonsourceibias.n204 gnd 0.059054f
C722 commonsourceibias.t67 gnd 0.148006f
C723 commonsourceibias.n205 gnd 0.006398f
C724 commonsourceibias.n206 gnd 0.007922f
C725 commonsourceibias.t93 gnd 0.148006f
C726 commonsourceibias.t108 gnd 0.148006f
C727 commonsourceibias.n207 gnd 0.059054f
C728 commonsourceibias.n208 gnd 0.007922f
C729 commonsourceibias.t127 gnd 0.148006f
C730 commonsourceibias.n209 gnd 0.059054f
C731 commonsourceibias.n210 gnd 0.007922f
C732 commonsourceibias.t86 gnd 0.148006f
C733 commonsourceibias.n211 gnd 0.059054f
C734 commonsourceibias.n212 gnd 0.007922f
C735 commonsourceibias.t82 gnd 0.148006f
C736 commonsourceibias.n213 gnd 0.009005f
C737 commonsourceibias.n214 gnd 0.007922f
C738 commonsourceibias.t96 gnd 0.148006f
C739 commonsourceibias.n215 gnd 0.010649f
C740 commonsourceibias.t75 gnd 0.164876f
C741 commonsourceibias.t77 gnd 0.148006f
C742 commonsourceibias.n216 gnd 0.065802f
C743 commonsourceibias.n217 gnd 0.070497f
C744 commonsourceibias.n218 gnd 0.03372f
C745 commonsourceibias.n219 gnd 0.007922f
C746 commonsourceibias.n220 gnd 0.006439f
C747 commonsourceibias.n221 gnd 0.010916f
C748 commonsourceibias.n222 gnd 0.059054f
C749 commonsourceibias.n223 gnd 0.010963f
C750 commonsourceibias.n224 gnd 0.007922f
C751 commonsourceibias.n225 gnd 0.007922f
C752 commonsourceibias.n226 gnd 0.007922f
C753 commonsourceibias.n227 gnd 0.008036f
C754 commonsourceibias.n228 gnd 0.059054f
C755 commonsourceibias.n229 gnd 0.009764f
C756 commonsourceibias.n230 gnd 0.010802f
C757 commonsourceibias.n231 gnd 0.007922f
C758 commonsourceibias.n232 gnd 0.007922f
C759 commonsourceibias.n233 gnd 0.010731f
C760 commonsourceibias.n234 gnd 0.006408f
C761 commonsourceibias.n235 gnd 0.010864f
C762 commonsourceibias.n236 gnd 0.007922f
C763 commonsourceibias.n237 gnd 0.007922f
C764 commonsourceibias.n238 gnd 0.010931f
C765 commonsourceibias.n239 gnd 0.009425f
C766 commonsourceibias.n240 gnd 0.007648f
C767 commonsourceibias.n241 gnd 0.007922f
C768 commonsourceibias.n242 gnd 0.007922f
C769 commonsourceibias.n243 gnd 0.00969f
C770 commonsourceibias.n244 gnd 0.010876f
C771 commonsourceibias.n245 gnd 0.059054f
C772 commonsourceibias.n246 gnd 0.010803f
C773 commonsourceibias.n247 gnd 0.007922f
C774 commonsourceibias.n248 gnd 0.007922f
C775 commonsourceibias.n249 gnd 0.007922f
C776 commonsourceibias.n250 gnd 0.010803f
C777 commonsourceibias.n251 gnd 0.059054f
C778 commonsourceibias.n252 gnd 0.010876f
C779 commonsourceibias.n253 gnd 0.00969f
C780 commonsourceibias.n254 gnd 0.007922f
C781 commonsourceibias.n255 gnd 0.007922f
C782 commonsourceibias.n256 gnd 0.007922f
C783 commonsourceibias.n257 gnd 0.009425f
C784 commonsourceibias.n258 gnd 0.010931f
C785 commonsourceibias.n259 gnd 0.059054f
C786 commonsourceibias.n260 gnd 0.010864f
C787 commonsourceibias.n261 gnd 0.007922f
C788 commonsourceibias.n262 gnd 0.007922f
C789 commonsourceibias.n263 gnd 0.007922f
C790 commonsourceibias.n264 gnd 0.010731f
C791 commonsourceibias.n265 gnd 0.059054f
C792 commonsourceibias.n266 gnd 0.010802f
C793 commonsourceibias.n267 gnd 0.009764f
C794 commonsourceibias.n268 gnd 0.007922f
C795 commonsourceibias.n269 gnd 0.007922f
C796 commonsourceibias.n270 gnd 0.007922f
C797 commonsourceibias.n271 gnd 0.009005f
C798 commonsourceibias.n272 gnd 0.010963f
C799 commonsourceibias.n273 gnd 0.059054f
C800 commonsourceibias.n274 gnd 0.010916f
C801 commonsourceibias.n275 gnd 0.007922f
C802 commonsourceibias.n276 gnd 0.007922f
C803 commonsourceibias.n277 gnd 0.007922f
C804 commonsourceibias.n278 gnd 0.010649f
C805 commonsourceibias.n279 gnd 0.059054f
C806 commonsourceibias.n280 gnd 0.010674f
C807 commonsourceibias.t81 gnd 0.160069f
C808 commonsourceibias.n281 gnd 0.071211f
C809 commonsourceibias.n282 gnd 0.025411f
C810 commonsourceibias.n283 gnd 0.458519f
C811 commonsourceibias.n284 gnd 0.010571f
C812 commonsourceibias.t110 gnd 0.160069f
C813 commonsourceibias.t123 gnd 0.148006f
C814 commonsourceibias.n285 gnd 0.006439f
C815 commonsourceibias.n286 gnd 0.007922f
C816 commonsourceibias.t68 gnd 0.148006f
C817 commonsourceibias.n287 gnd 0.008036f
C818 commonsourceibias.n288 gnd 0.007922f
C819 commonsourceibias.t117 gnd 0.148006f
C820 commonsourceibias.n289 gnd 0.006408f
C821 commonsourceibias.n290 gnd 0.007922f
C822 commonsourceibias.t64 gnd 0.148006f
C823 commonsourceibias.n291 gnd 0.007648f
C824 commonsourceibias.n292 gnd 0.007922f
C825 commonsourceibias.t90 gnd 0.148006f
C826 commonsourceibias.n293 gnd 0.006398f
C827 commonsourceibias.n294 gnd 0.007922f
C828 commonsourceibias.t122 gnd 0.148006f
C829 commonsourceibias.t69 gnd 0.148006f
C830 commonsourceibias.n295 gnd 0.059054f
C831 commonsourceibias.n296 gnd 0.007922f
C832 commonsourceibias.t66 gnd 0.148006f
C833 commonsourceibias.n297 gnd 0.059054f
C834 commonsourceibias.n298 gnd 0.007922f
C835 commonsourceibias.t116 gnd 0.148006f
C836 commonsourceibias.n299 gnd 0.059054f
C837 commonsourceibias.n300 gnd 0.007922f
C838 commonsourceibias.t113 gnd 0.148006f
C839 commonsourceibias.n301 gnd 0.009005f
C840 commonsourceibias.n302 gnd 0.007922f
C841 commonsourceibias.t126 gnd 0.148006f
C842 commonsourceibias.n303 gnd 0.010649f
C843 commonsourceibias.t91 gnd 0.164876f
C844 commonsourceibias.t83 gnd 0.148006f
C845 commonsourceibias.n304 gnd 0.065802f
C846 commonsourceibias.n305 gnd 0.070497f
C847 commonsourceibias.n306 gnd 0.03372f
C848 commonsourceibias.n307 gnd 0.007922f
C849 commonsourceibias.n308 gnd 0.006439f
C850 commonsourceibias.n309 gnd 0.010916f
C851 commonsourceibias.n310 gnd 0.059054f
C852 commonsourceibias.n311 gnd 0.010963f
C853 commonsourceibias.n312 gnd 0.007922f
C854 commonsourceibias.n313 gnd 0.007922f
C855 commonsourceibias.n314 gnd 0.007922f
C856 commonsourceibias.n315 gnd 0.008036f
C857 commonsourceibias.n316 gnd 0.059054f
C858 commonsourceibias.n317 gnd 0.009764f
C859 commonsourceibias.n318 gnd 0.010802f
C860 commonsourceibias.n319 gnd 0.007922f
C861 commonsourceibias.n320 gnd 0.007922f
C862 commonsourceibias.n321 gnd 0.010731f
C863 commonsourceibias.n322 gnd 0.006408f
C864 commonsourceibias.n323 gnd 0.010864f
C865 commonsourceibias.n324 gnd 0.007922f
C866 commonsourceibias.n325 gnd 0.007922f
C867 commonsourceibias.n326 gnd 0.010931f
C868 commonsourceibias.n327 gnd 0.009425f
C869 commonsourceibias.n328 gnd 0.007648f
C870 commonsourceibias.n329 gnd 0.007922f
C871 commonsourceibias.n330 gnd 0.007922f
C872 commonsourceibias.n331 gnd 0.00969f
C873 commonsourceibias.n332 gnd 0.010876f
C874 commonsourceibias.n333 gnd 0.059054f
C875 commonsourceibias.n334 gnd 0.010803f
C876 commonsourceibias.n335 gnd 0.007884f
C877 commonsourceibias.t55 gnd 0.017095f
C878 commonsourceibias.t53 gnd 0.017095f
C879 commonsourceibias.n336 gnd 0.15156f
C880 commonsourceibias.t3 gnd 0.017095f
C881 commonsourceibias.t49 gnd 0.017095f
C882 commonsourceibias.n337 gnd 0.151055f
C883 commonsourceibias.n338 gnd 0.140755f
C884 commonsourceibias.t41 gnd 0.017095f
C885 commonsourceibias.t59 gnd 0.017095f
C886 commonsourceibias.n339 gnd 0.151055f
C887 commonsourceibias.n340 gnd 0.069385f
C888 commonsourceibias.t51 gnd 0.017095f
C889 commonsourceibias.t25 gnd 0.017095f
C890 commonsourceibias.n341 gnd 0.151055f
C891 commonsourceibias.n342 gnd 0.057968f
C892 commonsourceibias.n343 gnd 0.010571f
C893 commonsourceibias.t34 gnd 0.148006f
C894 commonsourceibias.n344 gnd 0.006439f
C895 commonsourceibias.n345 gnd 0.007922f
C896 commonsourceibias.t0 gnd 0.148006f
C897 commonsourceibias.n346 gnd 0.008036f
C898 commonsourceibias.n347 gnd 0.007922f
C899 commonsourceibias.t46 gnd 0.148006f
C900 commonsourceibias.n348 gnd 0.006408f
C901 commonsourceibias.n349 gnd 0.007922f
C902 commonsourceibias.t10 gnd 0.148006f
C903 commonsourceibias.n350 gnd 0.007648f
C904 commonsourceibias.n351 gnd 0.007922f
C905 commonsourceibias.t44 gnd 0.148006f
C906 commonsourceibias.n352 gnd 0.006398f
C907 commonsourceibias.n353 gnd 0.007922f
C908 commonsourceibias.t24 gnd 0.148006f
C909 commonsourceibias.t50 gnd 0.148006f
C910 commonsourceibias.n354 gnd 0.059054f
C911 commonsourceibias.n355 gnd 0.007922f
C912 commonsourceibias.t58 gnd 0.148006f
C913 commonsourceibias.n356 gnd 0.059054f
C914 commonsourceibias.n357 gnd 0.007922f
C915 commonsourceibias.t40 gnd 0.148006f
C916 commonsourceibias.n358 gnd 0.059054f
C917 commonsourceibias.n359 gnd 0.007922f
C918 commonsourceibias.t48 gnd 0.148006f
C919 commonsourceibias.n360 gnd 0.009005f
C920 commonsourceibias.n361 gnd 0.007922f
C921 commonsourceibias.t2 gnd 0.148006f
C922 commonsourceibias.n362 gnd 0.010649f
C923 commonsourceibias.t54 gnd 0.164876f
C924 commonsourceibias.t52 gnd 0.148006f
C925 commonsourceibias.n363 gnd 0.065802f
C926 commonsourceibias.n364 gnd 0.070497f
C927 commonsourceibias.n365 gnd 0.03372f
C928 commonsourceibias.n366 gnd 0.007922f
C929 commonsourceibias.n367 gnd 0.006439f
C930 commonsourceibias.n368 gnd 0.010916f
C931 commonsourceibias.n369 gnd 0.059054f
C932 commonsourceibias.n370 gnd 0.010963f
C933 commonsourceibias.n371 gnd 0.007922f
C934 commonsourceibias.n372 gnd 0.007922f
C935 commonsourceibias.n373 gnd 0.007922f
C936 commonsourceibias.n374 gnd 0.008036f
C937 commonsourceibias.n375 gnd 0.059054f
C938 commonsourceibias.n376 gnd 0.009764f
C939 commonsourceibias.n377 gnd 0.010802f
C940 commonsourceibias.n378 gnd 0.007922f
C941 commonsourceibias.n379 gnd 0.007922f
C942 commonsourceibias.n380 gnd 0.010731f
C943 commonsourceibias.n381 gnd 0.006408f
C944 commonsourceibias.n382 gnd 0.010864f
C945 commonsourceibias.n383 gnd 0.007922f
C946 commonsourceibias.n384 gnd 0.007922f
C947 commonsourceibias.n385 gnd 0.010931f
C948 commonsourceibias.n386 gnd 0.009425f
C949 commonsourceibias.n387 gnd 0.007648f
C950 commonsourceibias.n388 gnd 0.007922f
C951 commonsourceibias.n389 gnd 0.007922f
C952 commonsourceibias.n390 gnd 0.00969f
C953 commonsourceibias.n391 gnd 0.010876f
C954 commonsourceibias.n392 gnd 0.059054f
C955 commonsourceibias.n393 gnd 0.010803f
C956 commonsourceibias.n394 gnd 0.007922f
C957 commonsourceibias.n395 gnd 0.007922f
C958 commonsourceibias.n396 gnd 0.007922f
C959 commonsourceibias.n397 gnd 0.010803f
C960 commonsourceibias.n398 gnd 0.059054f
C961 commonsourceibias.n399 gnd 0.010876f
C962 commonsourceibias.t36 gnd 0.148006f
C963 commonsourceibias.n400 gnd 0.059054f
C964 commonsourceibias.n401 gnd 0.00969f
C965 commonsourceibias.n402 gnd 0.007922f
C966 commonsourceibias.n403 gnd 0.007922f
C967 commonsourceibias.n404 gnd 0.007922f
C968 commonsourceibias.n405 gnd 0.009425f
C969 commonsourceibias.n406 gnd 0.010931f
C970 commonsourceibias.n407 gnd 0.059054f
C971 commonsourceibias.n408 gnd 0.010864f
C972 commonsourceibias.n409 gnd 0.007922f
C973 commonsourceibias.n410 gnd 0.007922f
C974 commonsourceibias.n411 gnd 0.007922f
C975 commonsourceibias.n412 gnd 0.010731f
C976 commonsourceibias.n413 gnd 0.059054f
C977 commonsourceibias.n414 gnd 0.010802f
C978 commonsourceibias.t22 gnd 0.148006f
C979 commonsourceibias.n415 gnd 0.059054f
C980 commonsourceibias.n416 gnd 0.009764f
C981 commonsourceibias.n417 gnd 0.007922f
C982 commonsourceibias.n418 gnd 0.007922f
C983 commonsourceibias.n419 gnd 0.007922f
C984 commonsourceibias.n420 gnd 0.009005f
C985 commonsourceibias.n421 gnd 0.010963f
C986 commonsourceibias.n422 gnd 0.059054f
C987 commonsourceibias.n423 gnd 0.010916f
C988 commonsourceibias.n424 gnd 0.007922f
C989 commonsourceibias.n425 gnd 0.007922f
C990 commonsourceibias.n426 gnd 0.007922f
C991 commonsourceibias.n427 gnd 0.010649f
C992 commonsourceibias.n428 gnd 0.059054f
C993 commonsourceibias.n429 gnd 0.010674f
C994 commonsourceibias.t8 gnd 0.160069f
C995 commonsourceibias.n430 gnd 0.071211f
C996 commonsourceibias.n431 gnd 0.079625f
C997 commonsourceibias.t35 gnd 0.017095f
C998 commonsourceibias.t9 gnd 0.017095f
C999 commonsourceibias.n432 gnd 0.151055f
C1000 commonsourceibias.n433 gnd 0.130846f
C1001 commonsourceibias.t23 gnd 0.017095f
C1002 commonsourceibias.t1 gnd 0.017095f
C1003 commonsourceibias.n434 gnd 0.151055f
C1004 commonsourceibias.n435 gnd 0.069385f
C1005 commonsourceibias.t11 gnd 0.017095f
C1006 commonsourceibias.t47 gnd 0.017095f
C1007 commonsourceibias.n436 gnd 0.151055f
C1008 commonsourceibias.n437 gnd 0.069385f
C1009 commonsourceibias.t45 gnd 0.017095f
C1010 commonsourceibias.t37 gnd 0.017095f
C1011 commonsourceibias.n438 gnd 0.151055f
C1012 commonsourceibias.n439 gnd 0.057968f
C1013 commonsourceibias.n440 gnd 0.070193f
C1014 commonsourceibias.n441 gnd 0.057266f
C1015 commonsourceibias.n442 gnd 0.007884f
C1016 commonsourceibias.n443 gnd 0.010803f
C1017 commonsourceibias.n444 gnd 0.059054f
C1018 commonsourceibias.n445 gnd 0.010876f
C1019 commonsourceibias.t72 gnd 0.148006f
C1020 commonsourceibias.n446 gnd 0.059054f
C1021 commonsourceibias.n447 gnd 0.00969f
C1022 commonsourceibias.n448 gnd 0.007922f
C1023 commonsourceibias.n449 gnd 0.007922f
C1024 commonsourceibias.n450 gnd 0.007922f
C1025 commonsourceibias.n451 gnd 0.009425f
C1026 commonsourceibias.n452 gnd 0.010931f
C1027 commonsourceibias.n453 gnd 0.059054f
C1028 commonsourceibias.n454 gnd 0.010864f
C1029 commonsourceibias.n455 gnd 0.007922f
C1030 commonsourceibias.n456 gnd 0.007922f
C1031 commonsourceibias.n457 gnd 0.007922f
C1032 commonsourceibias.n458 gnd 0.010731f
C1033 commonsourceibias.n459 gnd 0.059054f
C1034 commonsourceibias.n460 gnd 0.010802f
C1035 commonsourceibias.t102 gnd 0.148006f
C1036 commonsourceibias.n461 gnd 0.059054f
C1037 commonsourceibias.n462 gnd 0.009764f
C1038 commonsourceibias.n463 gnd 0.007922f
C1039 commonsourceibias.n464 gnd 0.007922f
C1040 commonsourceibias.n465 gnd 0.007922f
C1041 commonsourceibias.n466 gnd 0.009005f
C1042 commonsourceibias.n467 gnd 0.010963f
C1043 commonsourceibias.n468 gnd 0.059054f
C1044 commonsourceibias.n469 gnd 0.010916f
C1045 commonsourceibias.n470 gnd 0.007922f
C1046 commonsourceibias.n471 gnd 0.007922f
C1047 commonsourceibias.n472 gnd 0.007922f
C1048 commonsourceibias.n473 gnd 0.010649f
C1049 commonsourceibias.n474 gnd 0.059054f
C1050 commonsourceibias.n475 gnd 0.010674f
C1051 commonsourceibias.n476 gnd 0.071211f
C1052 commonsourceibias.n477 gnd 0.047027f
C1053 commonsourceibias.n478 gnd 0.010571f
C1054 commonsourceibias.t112 gnd 0.148006f
C1055 commonsourceibias.n479 gnd 0.006439f
C1056 commonsourceibias.n480 gnd 0.007922f
C1057 commonsourceibias.t124 gnd 0.148006f
C1058 commonsourceibias.n481 gnd 0.008036f
C1059 commonsourceibias.n482 gnd 0.007922f
C1060 commonsourceibias.t104 gnd 0.148006f
C1061 commonsourceibias.n483 gnd 0.006408f
C1062 commonsourceibias.n484 gnd 0.007922f
C1063 commonsourceibias.t118 gnd 0.148006f
C1064 commonsourceibias.n485 gnd 0.007648f
C1065 commonsourceibias.n486 gnd 0.007922f
C1066 commonsourceibias.t79 gnd 0.148006f
C1067 commonsourceibias.n487 gnd 0.006398f
C1068 commonsourceibias.n488 gnd 0.007922f
C1069 commonsourceibias.t111 gnd 0.148006f
C1070 commonsourceibias.t125 gnd 0.148006f
C1071 commonsourceibias.n489 gnd 0.059054f
C1072 commonsourceibias.n490 gnd 0.007922f
C1073 commonsourceibias.t120 gnd 0.148006f
C1074 commonsourceibias.n491 gnd 0.059054f
C1075 commonsourceibias.n492 gnd 0.007922f
C1076 commonsourceibias.t103 gnd 0.148006f
C1077 commonsourceibias.n493 gnd 0.059054f
C1078 commonsourceibias.n494 gnd 0.007922f
C1079 commonsourceibias.t98 gnd 0.148006f
C1080 commonsourceibias.n495 gnd 0.009005f
C1081 commonsourceibias.n496 gnd 0.007922f
C1082 commonsourceibias.t115 gnd 0.148006f
C1083 commonsourceibias.n497 gnd 0.010649f
C1084 commonsourceibias.t78 gnd 0.164876f
C1085 commonsourceibias.t73 gnd 0.148006f
C1086 commonsourceibias.n498 gnd 0.065802f
C1087 commonsourceibias.n499 gnd 0.070497f
C1088 commonsourceibias.n500 gnd 0.03372f
C1089 commonsourceibias.n501 gnd 0.007922f
C1090 commonsourceibias.n502 gnd 0.006439f
C1091 commonsourceibias.n503 gnd 0.010916f
C1092 commonsourceibias.n504 gnd 0.059054f
C1093 commonsourceibias.n505 gnd 0.010963f
C1094 commonsourceibias.n506 gnd 0.007922f
C1095 commonsourceibias.n507 gnd 0.007922f
C1096 commonsourceibias.n508 gnd 0.007922f
C1097 commonsourceibias.n509 gnd 0.008036f
C1098 commonsourceibias.n510 gnd 0.059054f
C1099 commonsourceibias.n511 gnd 0.009764f
C1100 commonsourceibias.n512 gnd 0.010802f
C1101 commonsourceibias.n513 gnd 0.007922f
C1102 commonsourceibias.n514 gnd 0.007922f
C1103 commonsourceibias.n515 gnd 0.010731f
C1104 commonsourceibias.n516 gnd 0.006408f
C1105 commonsourceibias.n517 gnd 0.010864f
C1106 commonsourceibias.n518 gnd 0.007922f
C1107 commonsourceibias.n519 gnd 0.007922f
C1108 commonsourceibias.n520 gnd 0.010931f
C1109 commonsourceibias.n521 gnd 0.009425f
C1110 commonsourceibias.n522 gnd 0.007648f
C1111 commonsourceibias.n523 gnd 0.007922f
C1112 commonsourceibias.n524 gnd 0.007922f
C1113 commonsourceibias.n525 gnd 0.00969f
C1114 commonsourceibias.n526 gnd 0.010876f
C1115 commonsourceibias.n527 gnd 0.059054f
C1116 commonsourceibias.n528 gnd 0.010803f
C1117 commonsourceibias.n529 gnd 0.007922f
C1118 commonsourceibias.n530 gnd 0.007922f
C1119 commonsourceibias.n531 gnd 0.007922f
C1120 commonsourceibias.n532 gnd 0.010803f
C1121 commonsourceibias.n533 gnd 0.059054f
C1122 commonsourceibias.n534 gnd 0.010876f
C1123 commonsourceibias.t65 gnd 0.148006f
C1124 commonsourceibias.n535 gnd 0.059054f
C1125 commonsourceibias.n536 gnd 0.00969f
C1126 commonsourceibias.n537 gnd 0.007922f
C1127 commonsourceibias.n538 gnd 0.007922f
C1128 commonsourceibias.n539 gnd 0.007922f
C1129 commonsourceibias.n540 gnd 0.009425f
C1130 commonsourceibias.n541 gnd 0.010931f
C1131 commonsourceibias.n542 gnd 0.059054f
C1132 commonsourceibias.n543 gnd 0.010864f
C1133 commonsourceibias.n544 gnd 0.007922f
C1134 commonsourceibias.n545 gnd 0.007922f
C1135 commonsourceibias.n546 gnd 0.007922f
C1136 commonsourceibias.n547 gnd 0.010731f
C1137 commonsourceibias.n548 gnd 0.059054f
C1138 commonsourceibias.n549 gnd 0.010802f
C1139 commonsourceibias.t88 gnd 0.148006f
C1140 commonsourceibias.n550 gnd 0.059054f
C1141 commonsourceibias.n551 gnd 0.009764f
C1142 commonsourceibias.n552 gnd 0.007922f
C1143 commonsourceibias.n553 gnd 0.007922f
C1144 commonsourceibias.n554 gnd 0.007922f
C1145 commonsourceibias.n555 gnd 0.009005f
C1146 commonsourceibias.n556 gnd 0.010963f
C1147 commonsourceibias.n557 gnd 0.059054f
C1148 commonsourceibias.n558 gnd 0.010916f
C1149 commonsourceibias.n559 gnd 0.007922f
C1150 commonsourceibias.n560 gnd 0.007922f
C1151 commonsourceibias.n561 gnd 0.007922f
C1152 commonsourceibias.n562 gnd 0.010649f
C1153 commonsourceibias.n563 gnd 0.059054f
C1154 commonsourceibias.n564 gnd 0.010674f
C1155 commonsourceibias.t97 gnd 0.160069f
C1156 commonsourceibias.n565 gnd 0.071211f
C1157 commonsourceibias.n566 gnd 0.025411f
C1158 commonsourceibias.n567 gnd 0.219034f
C1159 commonsourceibias.n568 gnd 4.63083f
C1160 minus.n0 gnd 0.031797f
C1161 minus.n1 gnd 0.007215f
C1162 minus.n2 gnd 0.031797f
C1163 minus.n3 gnd 0.007215f
C1164 minus.n4 gnd 0.031797f
C1165 minus.n5 gnd 0.007215f
C1166 minus.n6 gnd 0.031797f
C1167 minus.n7 gnd 0.007215f
C1168 minus.n8 gnd 0.031797f
C1169 minus.n9 gnd 0.007215f
C1170 minus.t8 gnd 0.466068f
C1171 minus.t7 gnd 0.449743f
C1172 minus.n10 gnd 0.206297f
C1173 minus.n11 gnd 0.185158f
C1174 minus.n12 gnd 0.136889f
C1175 minus.n13 gnd 0.031797f
C1176 minus.t11 gnd 0.449743f
C1177 minus.n14 gnd 0.19979f
C1178 minus.n15 gnd 0.007215f
C1179 minus.t10 gnd 0.449743f
C1180 minus.n16 gnd 0.19979f
C1181 minus.n17 gnd 0.031797f
C1182 minus.n18 gnd 0.031797f
C1183 minus.n19 gnd 0.031797f
C1184 minus.t12 gnd 0.449743f
C1185 minus.n20 gnd 0.19979f
C1186 minus.n21 gnd 0.007215f
C1187 minus.t20 gnd 0.449743f
C1188 minus.n22 gnd 0.19979f
C1189 minus.n23 gnd 0.031797f
C1190 minus.n24 gnd 0.031797f
C1191 minus.n25 gnd 0.031797f
C1192 minus.t18 gnd 0.449743f
C1193 minus.n26 gnd 0.19979f
C1194 minus.n27 gnd 0.007215f
C1195 minus.t25 gnd 0.449743f
C1196 minus.n28 gnd 0.19979f
C1197 minus.n29 gnd 0.031797f
C1198 minus.n30 gnd 0.031797f
C1199 minus.n31 gnd 0.031797f
C1200 minus.t24 gnd 0.449743f
C1201 minus.n32 gnd 0.19979f
C1202 minus.n33 gnd 0.007215f
C1203 minus.t14 gnd 0.449743f
C1204 minus.n34 gnd 0.19979f
C1205 minus.n35 gnd 0.031797f
C1206 minus.n36 gnd 0.031797f
C1207 minus.n37 gnd 0.031797f
C1208 minus.t22 gnd 0.449743f
C1209 minus.n38 gnd 0.19979f
C1210 minus.n39 gnd 0.007215f
C1211 minus.t19 gnd 0.449743f
C1212 minus.n40 gnd 0.200084f
C1213 minus.n41 gnd 0.368244f
C1214 minus.n42 gnd 0.031797f
C1215 minus.t13 gnd 0.449743f
C1216 minus.t15 gnd 0.449743f
C1217 minus.n43 gnd 0.031797f
C1218 minus.t5 gnd 0.449743f
C1219 minus.n44 gnd 0.19979f
C1220 minus.n45 gnd 0.031797f
C1221 minus.t6 gnd 0.449743f
C1222 minus.t26 gnd 0.449743f
C1223 minus.n46 gnd 0.19979f
C1224 minus.n47 gnd 0.031797f
C1225 minus.t21 gnd 0.449743f
C1226 minus.t23 gnd 0.449743f
C1227 minus.n48 gnd 0.19979f
C1228 minus.n49 gnd 0.031797f
C1229 minus.t16 gnd 0.449743f
C1230 minus.t17 gnd 0.449743f
C1231 minus.n50 gnd 0.19979f
C1232 minus.n51 gnd 0.031797f
C1233 minus.t9 gnd 0.449743f
C1234 minus.t27 gnd 0.449743f
C1235 minus.n52 gnd 0.206297f
C1236 minus.t28 gnd 0.466068f
C1237 minus.n53 gnd 0.185158f
C1238 minus.n54 gnd 0.136889f
C1239 minus.n55 gnd 0.007215f
C1240 minus.n56 gnd 0.19979f
C1241 minus.n57 gnd 0.007215f
C1242 minus.n58 gnd 0.031797f
C1243 minus.n59 gnd 0.031797f
C1244 minus.n60 gnd 0.031797f
C1245 minus.n61 gnd 0.007215f
C1246 minus.n62 gnd 0.19979f
C1247 minus.n63 gnd 0.007215f
C1248 minus.n64 gnd 0.031797f
C1249 minus.n65 gnd 0.031797f
C1250 minus.n66 gnd 0.031797f
C1251 minus.n67 gnd 0.007215f
C1252 minus.n68 gnd 0.19979f
C1253 minus.n69 gnd 0.007215f
C1254 minus.n70 gnd 0.031797f
C1255 minus.n71 gnd 0.031797f
C1256 minus.n72 gnd 0.031797f
C1257 minus.n73 gnd 0.007215f
C1258 minus.n74 gnd 0.19979f
C1259 minus.n75 gnd 0.007215f
C1260 minus.n76 gnd 0.031797f
C1261 minus.n77 gnd 0.031797f
C1262 minus.n78 gnd 0.031797f
C1263 minus.n79 gnd 0.007215f
C1264 minus.n80 gnd 0.19979f
C1265 minus.n81 gnd 0.007215f
C1266 minus.n82 gnd 0.200084f
C1267 minus.n83 gnd 1.06524f
C1268 minus.n84 gnd 1.58719f
C1269 minus.t1 gnd 0.009802f
C1270 minus.t0 gnd 0.009802f
C1271 minus.n85 gnd 0.032232f
C1272 minus.t4 gnd 0.009802f
C1273 minus.t3 gnd 0.009802f
C1274 minus.n86 gnd 0.03179f
C1275 minus.n87 gnd 0.271314f
C1276 minus.t2 gnd 0.054558f
C1277 minus.n88 gnd 0.148054f
C1278 minus.n89 gnd 2.10933f
C1279 CSoutput.n0 gnd 0.044585f
C1280 CSoutput.t173 gnd 0.294918f
C1281 CSoutput.n1 gnd 0.13317f
C1282 CSoutput.n2 gnd 0.044585f
C1283 CSoutput.t179 gnd 0.294918f
C1284 CSoutput.n3 gnd 0.035337f
C1285 CSoutput.n4 gnd 0.044585f
C1286 CSoutput.t168 gnd 0.294918f
C1287 CSoutput.n5 gnd 0.030471f
C1288 CSoutput.n6 gnd 0.044585f
C1289 CSoutput.t176 gnd 0.294918f
C1290 CSoutput.t160 gnd 0.294918f
C1291 CSoutput.n7 gnd 0.131719f
C1292 CSoutput.n8 gnd 0.044585f
C1293 CSoutput.t181 gnd 0.294918f
C1294 CSoutput.n9 gnd 0.029053f
C1295 CSoutput.n10 gnd 0.044585f
C1296 CSoutput.t169 gnd 0.294918f
C1297 CSoutput.t180 gnd 0.294918f
C1298 CSoutput.n11 gnd 0.131719f
C1299 CSoutput.n12 gnd 0.044585f
C1300 CSoutput.t177 gnd 0.294918f
C1301 CSoutput.n13 gnd 0.030471f
C1302 CSoutput.n14 gnd 0.044585f
C1303 CSoutput.t167 gnd 0.294918f
C1304 CSoutput.t170 gnd 0.294918f
C1305 CSoutput.n15 gnd 0.131719f
C1306 CSoutput.n16 gnd 0.044585f
C1307 CSoutput.t174 gnd 0.294918f
C1308 CSoutput.n17 gnd 0.032545f
C1309 CSoutput.t164 gnd 0.352435f
C1310 CSoutput.t166 gnd 0.294918f
C1311 CSoutput.n18 gnd 0.168154f
C1312 CSoutput.n19 gnd 0.163167f
C1313 CSoutput.n20 gnd 0.189294f
C1314 CSoutput.n21 gnd 0.044585f
C1315 CSoutput.n22 gnd 0.037211f
C1316 CSoutput.n23 gnd 0.131719f
C1317 CSoutput.n24 gnd 0.03587f
C1318 CSoutput.n25 gnd 0.035337f
C1319 CSoutput.n26 gnd 0.044585f
C1320 CSoutput.n27 gnd 0.044585f
C1321 CSoutput.n28 gnd 0.036925f
C1322 CSoutput.n29 gnd 0.03135f
C1323 CSoutput.n30 gnd 0.134651f
C1324 CSoutput.n31 gnd 0.031782f
C1325 CSoutput.n32 gnd 0.044585f
C1326 CSoutput.n33 gnd 0.044585f
C1327 CSoutput.n34 gnd 0.044585f
C1328 CSoutput.n35 gnd 0.036532f
C1329 CSoutput.n36 gnd 0.131719f
C1330 CSoutput.n37 gnd 0.034937f
C1331 CSoutput.n38 gnd 0.03627f
C1332 CSoutput.n39 gnd 0.044585f
C1333 CSoutput.n40 gnd 0.044585f
C1334 CSoutput.n41 gnd 0.037203f
C1335 CSoutput.n42 gnd 0.034004f
C1336 CSoutput.n43 gnd 0.131719f
C1337 CSoutput.n44 gnd 0.034866f
C1338 CSoutput.n45 gnd 0.044585f
C1339 CSoutput.n46 gnd 0.044585f
C1340 CSoutput.n47 gnd 0.044585f
C1341 CSoutput.n48 gnd 0.034866f
C1342 CSoutput.n49 gnd 0.131719f
C1343 CSoutput.n50 gnd 0.034004f
C1344 CSoutput.n51 gnd 0.037203f
C1345 CSoutput.n52 gnd 0.044585f
C1346 CSoutput.n53 gnd 0.044585f
C1347 CSoutput.n54 gnd 0.03627f
C1348 CSoutput.n55 gnd 0.034937f
C1349 CSoutput.n56 gnd 0.131719f
C1350 CSoutput.n57 gnd 0.036532f
C1351 CSoutput.n58 gnd 0.044585f
C1352 CSoutput.n59 gnd 0.044585f
C1353 CSoutput.n60 gnd 0.044585f
C1354 CSoutput.n61 gnd 0.031782f
C1355 CSoutput.n62 gnd 0.134651f
C1356 CSoutput.n63 gnd 0.03135f
C1357 CSoutput.t162 gnd 0.294918f
C1358 CSoutput.n64 gnd 0.131719f
C1359 CSoutput.n65 gnd 0.036925f
C1360 CSoutput.n66 gnd 0.044585f
C1361 CSoutput.n67 gnd 0.044585f
C1362 CSoutput.n68 gnd 0.044585f
C1363 CSoutput.n69 gnd 0.03587f
C1364 CSoutput.n70 gnd 0.131719f
C1365 CSoutput.n71 gnd 0.037211f
C1366 CSoutput.n72 gnd 0.032545f
C1367 CSoutput.n73 gnd 0.044585f
C1368 CSoutput.n74 gnd 0.044585f
C1369 CSoutput.n75 gnd 0.033751f
C1370 CSoutput.n76 gnd 0.020045f
C1371 CSoutput.t165 gnd 0.331362f
C1372 CSoutput.n77 gnd 0.164607f
C1373 CSoutput.n78 gnd 0.704339f
C1374 CSoutput.t105 gnd 0.055613f
C1375 CSoutput.t53 gnd 0.055613f
C1376 CSoutput.n79 gnd 0.430575f
C1377 CSoutput.t21 gnd 0.055613f
C1378 CSoutput.t87 gnd 0.055613f
C1379 CSoutput.n80 gnd 0.429808f
C1380 CSoutput.n81 gnd 0.436254f
C1381 CSoutput.t28 gnd 0.055613f
C1382 CSoutput.t72 gnd 0.055613f
C1383 CSoutput.n82 gnd 0.429808f
C1384 CSoutput.n83 gnd 0.214968f
C1385 CSoutput.t44 gnd 0.055613f
C1386 CSoutput.t60 gnd 0.055613f
C1387 CSoutput.n84 gnd 0.429808f
C1388 CSoutput.n85 gnd 0.214968f
C1389 CSoutput.t56 gnd 0.055613f
C1390 CSoutput.t95 gnd 0.055613f
C1391 CSoutput.n86 gnd 0.429808f
C1392 CSoutput.n87 gnd 0.214968f
C1393 CSoutput.t35 gnd 0.055613f
C1394 CSoutput.t77 gnd 0.055613f
C1395 CSoutput.n88 gnd 0.429808f
C1396 CSoutput.n89 gnd 0.214968f
C1397 CSoutput.t49 gnd 0.055613f
C1398 CSoutput.t89 gnd 0.055613f
C1399 CSoutput.n90 gnd 0.429808f
C1400 CSoutput.n91 gnd 0.214968f
C1401 CSoutput.t64 gnd 0.055613f
C1402 CSoutput.t102 gnd 0.055613f
C1403 CSoutput.n92 gnd 0.429808f
C1404 CSoutput.n93 gnd 0.394201f
C1405 CSoutput.t57 gnd 0.055613f
C1406 CSoutput.t30 gnd 0.055613f
C1407 CSoutput.n94 gnd 0.430575f
C1408 CSoutput.t14 gnd 0.055613f
C1409 CSoutput.t59 gnd 0.055613f
C1410 CSoutput.n95 gnd 0.429808f
C1411 CSoutput.n96 gnd 0.436254f
C1412 CSoutput.t54 gnd 0.055613f
C1413 CSoutput.t27 gnd 0.055613f
C1414 CSoutput.n97 gnd 0.429808f
C1415 CSoutput.n98 gnd 0.214968f
C1416 CSoutput.t13 gnd 0.055613f
C1417 CSoutput.t11 gnd 0.055613f
C1418 CSoutput.n99 gnd 0.429808f
C1419 CSoutput.n100 gnd 0.214968f
C1420 CSoutput.t73 gnd 0.055613f
C1421 CSoutput.t40 gnd 0.055613f
C1422 CSoutput.n101 gnd 0.429808f
C1423 CSoutput.n102 gnd 0.214968f
C1424 CSoutput.t37 gnd 0.055613f
C1425 CSoutput.t10 gnd 0.055613f
C1426 CSoutput.n103 gnd 0.429808f
C1427 CSoutput.n104 gnd 0.214968f
C1428 CSoutput.t93 gnd 0.055613f
C1429 CSoutput.t70 gnd 0.055613f
C1430 CSoutput.n105 gnd 0.429808f
C1431 CSoutput.n106 gnd 0.214968f
C1432 CSoutput.t58 gnd 0.055613f
C1433 CSoutput.t31 gnd 0.055613f
C1434 CSoutput.n107 gnd 0.429808f
C1435 CSoutput.n108 gnd 0.320571f
C1436 CSoutput.n109 gnd 0.404238f
C1437 CSoutput.t66 gnd 0.055613f
C1438 CSoutput.t41 gnd 0.055613f
C1439 CSoutput.n110 gnd 0.430575f
C1440 CSoutput.t24 gnd 0.055613f
C1441 CSoutput.t68 gnd 0.055613f
C1442 CSoutput.n111 gnd 0.429808f
C1443 CSoutput.n112 gnd 0.436254f
C1444 CSoutput.t65 gnd 0.055613f
C1445 CSoutput.t39 gnd 0.055613f
C1446 CSoutput.n113 gnd 0.429808f
C1447 CSoutput.n114 gnd 0.214968f
C1448 CSoutput.t23 gnd 0.055613f
C1449 CSoutput.t22 gnd 0.055613f
C1450 CSoutput.n115 gnd 0.429808f
C1451 CSoutput.n116 gnd 0.214968f
C1452 CSoutput.t80 gnd 0.055613f
C1453 CSoutput.t50 gnd 0.055613f
C1454 CSoutput.n117 gnd 0.429808f
C1455 CSoutput.n118 gnd 0.214968f
C1456 CSoutput.t46 gnd 0.055613f
C1457 CSoutput.t19 gnd 0.055613f
C1458 CSoutput.n119 gnd 0.429808f
C1459 CSoutput.n120 gnd 0.214968f
C1460 CSoutput.t103 gnd 0.055613f
C1461 CSoutput.t79 gnd 0.055613f
C1462 CSoutput.n121 gnd 0.429808f
C1463 CSoutput.n122 gnd 0.214968f
C1464 CSoutput.t67 gnd 0.055613f
C1465 CSoutput.t42 gnd 0.055613f
C1466 CSoutput.n123 gnd 0.429808f
C1467 CSoutput.n124 gnd 0.320571f
C1468 CSoutput.n125 gnd 0.451834f
C1469 CSoutput.n126 gnd 8.9793f
C1470 CSoutput.n128 gnd 0.788695f
C1471 CSoutput.n129 gnd 0.591522f
C1472 CSoutput.n130 gnd 0.788695f
C1473 CSoutput.n131 gnd 0.788695f
C1474 CSoutput.n132 gnd 2.12341f
C1475 CSoutput.n133 gnd 0.788695f
C1476 CSoutput.n134 gnd 0.788695f
C1477 CSoutput.t161 gnd 0.985869f
C1478 CSoutput.n135 gnd 0.788695f
C1479 CSoutput.n136 gnd 0.788695f
C1480 CSoutput.n140 gnd 0.788695f
C1481 CSoutput.n144 gnd 0.788695f
C1482 CSoutput.n145 gnd 0.788695f
C1483 CSoutput.n147 gnd 0.788695f
C1484 CSoutput.n152 gnd 0.788695f
C1485 CSoutput.n154 gnd 0.788695f
C1486 CSoutput.n155 gnd 0.788695f
C1487 CSoutput.n157 gnd 0.788695f
C1488 CSoutput.n158 gnd 0.788695f
C1489 CSoutput.n160 gnd 0.788695f
C1490 CSoutput.t172 gnd 13.179f
C1491 CSoutput.n162 gnd 0.788695f
C1492 CSoutput.n163 gnd 0.591522f
C1493 CSoutput.n164 gnd 0.788695f
C1494 CSoutput.n165 gnd 0.788695f
C1495 CSoutput.n166 gnd 2.12341f
C1496 CSoutput.n167 gnd 0.788695f
C1497 CSoutput.n168 gnd 0.788695f
C1498 CSoutput.t175 gnd 0.985869f
C1499 CSoutput.n169 gnd 0.788695f
C1500 CSoutput.n170 gnd 0.788695f
C1501 CSoutput.n174 gnd 0.788695f
C1502 CSoutput.n178 gnd 0.788695f
C1503 CSoutput.n179 gnd 0.788695f
C1504 CSoutput.n181 gnd 0.788695f
C1505 CSoutput.n186 gnd 0.788695f
C1506 CSoutput.n188 gnd 0.788695f
C1507 CSoutput.n189 gnd 0.788695f
C1508 CSoutput.n191 gnd 0.788695f
C1509 CSoutput.n192 gnd 0.788695f
C1510 CSoutput.n194 gnd 0.788695f
C1511 CSoutput.n195 gnd 0.591522f
C1512 CSoutput.n197 gnd 0.788695f
C1513 CSoutput.n198 gnd 0.591522f
C1514 CSoutput.n199 gnd 0.788695f
C1515 CSoutput.n200 gnd 0.788695f
C1516 CSoutput.n201 gnd 2.12341f
C1517 CSoutput.n202 gnd 0.788695f
C1518 CSoutput.n203 gnd 0.788695f
C1519 CSoutput.t171 gnd 0.985869f
C1520 CSoutput.n204 gnd 0.788695f
C1521 CSoutput.n205 gnd 2.12341f
C1522 CSoutput.n207 gnd 0.788695f
C1523 CSoutput.n208 gnd 0.788695f
C1524 CSoutput.n210 gnd 0.788695f
C1525 CSoutput.n211 gnd 0.788695f
C1526 CSoutput.t178 gnd 12.9642f
C1527 CSoutput.t163 gnd 13.179f
C1528 CSoutput.n217 gnd 2.47425f
C1529 CSoutput.n218 gnd 10.0792f
C1530 CSoutput.n219 gnd 10.501f
C1531 CSoutput.n224 gnd 2.68028f
C1532 CSoutput.n230 gnd 0.788695f
C1533 CSoutput.n232 gnd 0.788695f
C1534 CSoutput.n234 gnd 0.788695f
C1535 CSoutput.n236 gnd 0.788695f
C1536 CSoutput.n238 gnd 0.788695f
C1537 CSoutput.n244 gnd 0.788695f
C1538 CSoutput.n251 gnd 1.44695f
C1539 CSoutput.n252 gnd 1.44695f
C1540 CSoutput.n253 gnd 0.788695f
C1541 CSoutput.n254 gnd 0.788695f
C1542 CSoutput.n256 gnd 0.591522f
C1543 CSoutput.n257 gnd 0.506585f
C1544 CSoutput.n259 gnd 0.591522f
C1545 CSoutput.n260 gnd 0.506585f
C1546 CSoutput.n261 gnd 0.591522f
C1547 CSoutput.n263 gnd 0.788695f
C1548 CSoutput.n265 gnd 2.12341f
C1549 CSoutput.n266 gnd 2.47425f
C1550 CSoutput.n267 gnd 9.27028f
C1551 CSoutput.n269 gnd 0.591522f
C1552 CSoutput.n270 gnd 1.52202f
C1553 CSoutput.n271 gnd 0.591522f
C1554 CSoutput.n273 gnd 0.788695f
C1555 CSoutput.n275 gnd 2.12341f
C1556 CSoutput.n276 gnd 4.62513f
C1557 CSoutput.t52 gnd 0.055613f
C1558 CSoutput.t34 gnd 0.055613f
C1559 CSoutput.n277 gnd 0.430575f
C1560 CSoutput.t86 gnd 0.055613f
C1561 CSoutput.t20 gnd 0.055613f
C1562 CSoutput.n278 gnd 0.429808f
C1563 CSoutput.n279 gnd 0.436254f
C1564 CSoutput.t71 gnd 0.055613f
C1565 CSoutput.t25 gnd 0.055613f
C1566 CSoutput.n280 gnd 0.429808f
C1567 CSoutput.n281 gnd 0.214968f
C1568 CSoutput.t82 gnd 0.055613f
C1569 CSoutput.t43 gnd 0.055613f
C1570 CSoutput.n282 gnd 0.429808f
C1571 CSoutput.n283 gnd 0.214968f
C1572 CSoutput.t94 gnd 0.055613f
C1573 CSoutput.t55 gnd 0.055613f
C1574 CSoutput.n284 gnd 0.429808f
C1575 CSoutput.n285 gnd 0.214968f
C1576 CSoutput.t76 gnd 0.055613f
C1577 CSoutput.t36 gnd 0.055613f
C1578 CSoutput.n286 gnd 0.429808f
C1579 CSoutput.n287 gnd 0.214968f
C1580 CSoutput.t88 gnd 0.055613f
C1581 CSoutput.t48 gnd 0.055613f
C1582 CSoutput.n288 gnd 0.429808f
C1583 CSoutput.n289 gnd 0.214968f
C1584 CSoutput.t101 gnd 0.055613f
C1585 CSoutput.t62 gnd 0.055613f
C1586 CSoutput.n290 gnd 0.429808f
C1587 CSoutput.n291 gnd 0.394201f
C1588 CSoutput.t91 gnd 0.055613f
C1589 CSoutput.t92 gnd 0.055613f
C1590 CSoutput.n292 gnd 0.430575f
C1591 CSoutput.t18 gnd 0.055613f
C1592 CSoutput.t78 gnd 0.055613f
C1593 CSoutput.n293 gnd 0.429808f
C1594 CSoutput.n294 gnd 0.436254f
C1595 CSoutput.t85 gnd 0.055613f
C1596 CSoutput.t15 gnd 0.055613f
C1597 CSoutput.n295 gnd 0.429808f
C1598 CSoutput.n296 gnd 0.214968f
C1599 CSoutput.t51 gnd 0.055613f
C1600 CSoutput.t75 gnd 0.055613f
C1601 CSoutput.n297 gnd 0.429808f
C1602 CSoutput.n298 gnd 0.214968f
C1603 CSoutput.t97 gnd 0.055613f
C1604 CSoutput.t38 gnd 0.055613f
C1605 CSoutput.n299 gnd 0.429808f
C1606 CSoutput.n300 gnd 0.214968f
C1607 CSoutput.t74 gnd 0.055613f
C1608 CSoutput.t104 gnd 0.055613f
C1609 CSoutput.n301 gnd 0.429808f
C1610 CSoutput.n302 gnd 0.214968f
C1611 CSoutput.t33 gnd 0.055613f
C1612 CSoutput.t61 gnd 0.055613f
C1613 CSoutput.n303 gnd 0.429808f
C1614 CSoutput.n304 gnd 0.214968f
C1615 CSoutput.t90 gnd 0.055613f
C1616 CSoutput.t17 gnd 0.055613f
C1617 CSoutput.n305 gnd 0.429808f
C1618 CSoutput.n306 gnd 0.320571f
C1619 CSoutput.n307 gnd 0.404238f
C1620 CSoutput.t98 gnd 0.055613f
C1621 CSoutput.t100 gnd 0.055613f
C1622 CSoutput.n308 gnd 0.430575f
C1623 CSoutput.t32 gnd 0.055613f
C1624 CSoutput.t84 gnd 0.055613f
C1625 CSoutput.n309 gnd 0.429808f
C1626 CSoutput.n310 gnd 0.436254f
C1627 CSoutput.t96 gnd 0.055613f
C1628 CSoutput.t26 gnd 0.055613f
C1629 CSoutput.n311 gnd 0.429808f
C1630 CSoutput.n312 gnd 0.214968f
C1631 CSoutput.t63 gnd 0.055613f
C1632 CSoutput.t83 gnd 0.055613f
C1633 CSoutput.n313 gnd 0.429808f
C1634 CSoutput.n314 gnd 0.214968f
C1635 CSoutput.t12 gnd 0.055613f
C1636 CSoutput.t47 gnd 0.055613f
C1637 CSoutput.n315 gnd 0.429808f
C1638 CSoutput.n316 gnd 0.214968f
C1639 CSoutput.t81 gnd 0.055613f
C1640 CSoutput.t16 gnd 0.055613f
C1641 CSoutput.n317 gnd 0.429808f
C1642 CSoutput.n318 gnd 0.214968f
C1643 CSoutput.t45 gnd 0.055613f
C1644 CSoutput.t69 gnd 0.055613f
C1645 CSoutput.n319 gnd 0.429808f
C1646 CSoutput.n320 gnd 0.214968f
C1647 CSoutput.t99 gnd 0.055613f
C1648 CSoutput.t29 gnd 0.055613f
C1649 CSoutput.n321 gnd 0.429806f
C1650 CSoutput.n322 gnd 0.320572f
C1651 CSoutput.n323 gnd 0.451834f
C1652 CSoutput.n324 gnd 12.5737f
C1653 CSoutput.t118 gnd 0.048662f
C1654 CSoutput.t136 gnd 0.048662f
C1655 CSoutput.n325 gnd 0.431429f
C1656 CSoutput.t145 gnd 0.048662f
C1657 CSoutput.t115 gnd 0.048662f
C1658 CSoutput.n326 gnd 0.42999f
C1659 CSoutput.n327 gnd 0.40067f
C1660 CSoutput.t155 gnd 0.048662f
C1661 CSoutput.t132 gnd 0.048662f
C1662 CSoutput.n328 gnd 0.42999f
C1663 CSoutput.n329 gnd 0.197512f
C1664 CSoutput.t119 gnd 0.048662f
C1665 CSoutput.t149 gnd 0.048662f
C1666 CSoutput.n330 gnd 0.42999f
C1667 CSoutput.n331 gnd 0.197512f
C1668 CSoutput.t114 gnd 0.048662f
C1669 CSoutput.t111 gnd 0.048662f
C1670 CSoutput.n332 gnd 0.42999f
C1671 CSoutput.n333 gnd 0.197512f
C1672 CSoutput.t108 gnd 0.048662f
C1673 CSoutput.t106 gnd 0.048662f
C1674 CSoutput.n334 gnd 0.42999f
C1675 CSoutput.n335 gnd 0.197512f
C1676 CSoutput.t107 gnd 0.048662f
C1677 CSoutput.t146 gnd 0.048662f
C1678 CSoutput.n336 gnd 0.42999f
C1679 CSoutput.n337 gnd 0.197512f
C1680 CSoutput.t156 gnd 0.048662f
C1681 CSoutput.t4 gnd 0.048662f
C1682 CSoutput.n338 gnd 0.42999f
C1683 CSoutput.n339 gnd 0.364251f
C1684 CSoutput.t148 gnd 0.048662f
C1685 CSoutput.t154 gnd 0.048662f
C1686 CSoutput.n340 gnd 0.431429f
C1687 CSoutput.t137 gnd 0.048662f
C1688 CSoutput.t153 gnd 0.048662f
C1689 CSoutput.n341 gnd 0.42999f
C1690 CSoutput.n342 gnd 0.40067f
C1691 CSoutput.t0 gnd 0.048662f
C1692 CSoutput.t158 gnd 0.048662f
C1693 CSoutput.n343 gnd 0.42999f
C1694 CSoutput.n344 gnd 0.197512f
C1695 CSoutput.t129 gnd 0.048662f
C1696 CSoutput.t117 gnd 0.048662f
C1697 CSoutput.n345 gnd 0.42999f
C1698 CSoutput.n346 gnd 0.197512f
C1699 CSoutput.t8 gnd 0.048662f
C1700 CSoutput.t147 gnd 0.048662f
C1701 CSoutput.n347 gnd 0.42999f
C1702 CSoutput.n348 gnd 0.197512f
C1703 CSoutput.t1 gnd 0.048662f
C1704 CSoutput.t7 gnd 0.048662f
C1705 CSoutput.n349 gnd 0.42999f
C1706 CSoutput.n350 gnd 0.197512f
C1707 CSoutput.t127 gnd 0.048662f
C1708 CSoutput.t142 gnd 0.048662f
C1709 CSoutput.n351 gnd 0.42999f
C1710 CSoutput.n352 gnd 0.197512f
C1711 CSoutput.t157 gnd 0.048662f
C1712 CSoutput.t128 gnd 0.048662f
C1713 CSoutput.n353 gnd 0.42999f
C1714 CSoutput.n354 gnd 0.299865f
C1715 CSoutput.n355 gnd 0.557172f
C1716 CSoutput.n356 gnd 12.877f
C1717 CSoutput.t143 gnd 0.048662f
C1718 CSoutput.t124 gnd 0.048662f
C1719 CSoutput.n357 gnd 0.431429f
C1720 CSoutput.t138 gnd 0.048662f
C1721 CSoutput.t120 gnd 0.048662f
C1722 CSoutput.n358 gnd 0.42999f
C1723 CSoutput.n359 gnd 0.40067f
C1724 CSoutput.t130 gnd 0.048662f
C1725 CSoutput.t152 gnd 0.048662f
C1726 CSoutput.n360 gnd 0.42999f
C1727 CSoutput.n361 gnd 0.197512f
C1728 CSoutput.t3 gnd 0.048662f
C1729 CSoutput.t134 gnd 0.048662f
C1730 CSoutput.n362 gnd 0.42999f
C1731 CSoutput.n363 gnd 0.197512f
C1732 CSoutput.t159 gnd 0.048662f
C1733 CSoutput.t144 gnd 0.048662f
C1734 CSoutput.n364 gnd 0.42999f
C1735 CSoutput.n365 gnd 0.197512f
C1736 CSoutput.t6 gnd 0.048662f
C1737 CSoutput.t150 gnd 0.048662f
C1738 CSoutput.n366 gnd 0.42999f
C1739 CSoutput.n367 gnd 0.197512f
C1740 CSoutput.t109 gnd 0.048662f
C1741 CSoutput.t2 gnd 0.048662f
C1742 CSoutput.n368 gnd 0.42999f
C1743 CSoutput.n369 gnd 0.197512f
C1744 CSoutput.t139 gnd 0.048662f
C1745 CSoutput.t116 gnd 0.048662f
C1746 CSoutput.n370 gnd 0.42999f
C1747 CSoutput.n371 gnd 0.364251f
C1748 CSoutput.t112 gnd 0.048662f
C1749 CSoutput.t141 gnd 0.048662f
C1750 CSoutput.n372 gnd 0.431429f
C1751 CSoutput.t9 gnd 0.048662f
C1752 CSoutput.t121 gnd 0.048662f
C1753 CSoutput.n373 gnd 0.42999f
C1754 CSoutput.n374 gnd 0.40067f
C1755 CSoutput.t123 gnd 0.048662f
C1756 CSoutput.t125 gnd 0.048662f
C1757 CSoutput.n375 gnd 0.42999f
C1758 CSoutput.n376 gnd 0.197512f
C1759 CSoutput.t140 gnd 0.048662f
C1760 CSoutput.t131 gnd 0.048662f
C1761 CSoutput.n377 gnd 0.42999f
C1762 CSoutput.n378 gnd 0.197512f
C1763 CSoutput.t110 gnd 0.048662f
C1764 CSoutput.t113 gnd 0.048662f
C1765 CSoutput.n379 gnd 0.42999f
C1766 CSoutput.n380 gnd 0.197512f
C1767 CSoutput.t126 gnd 0.048662f
C1768 CSoutput.t122 gnd 0.048662f
C1769 CSoutput.n381 gnd 0.42999f
C1770 CSoutput.n382 gnd 0.197512f
C1771 CSoutput.t133 gnd 0.048662f
C1772 CSoutput.t151 gnd 0.048662f
C1773 CSoutput.n383 gnd 0.42999f
C1774 CSoutput.n384 gnd 0.197512f
C1775 CSoutput.t5 gnd 0.048662f
C1776 CSoutput.t135 gnd 0.048662f
C1777 CSoutput.n385 gnd 0.42999f
C1778 CSoutput.n386 gnd 0.299865f
C1779 CSoutput.n387 gnd 0.557172f
C1780 CSoutput.n388 gnd 7.74668f
C1781 CSoutput.n389 gnd 14.2929f
C1782 a_n2804_13878.t17 gnd 0.194556f
C1783 a_n2804_13878.t4 gnd 0.194556f
C1784 a_n2804_13878.t14 gnd 0.194556f
C1785 a_n2804_13878.n0 gnd 1.53358f
C1786 a_n2804_13878.t19 gnd 0.194556f
C1787 a_n2804_13878.t9 gnd 0.194556f
C1788 a_n2804_13878.n1 gnd 1.53196f
C1789 a_n2804_13878.n2 gnd 2.14061f
C1790 a_n2804_13878.t15 gnd 0.194556f
C1791 a_n2804_13878.t8 gnd 0.194556f
C1792 a_n2804_13878.n3 gnd 1.53196f
C1793 a_n2804_13878.n4 gnd 1.04414f
C1794 a_n2804_13878.t2 gnd 0.194556f
C1795 a_n2804_13878.t5 gnd 0.194556f
C1796 a_n2804_13878.n5 gnd 1.53196f
C1797 a_n2804_13878.n6 gnd 1.04414f
C1798 a_n2804_13878.t18 gnd 0.194556f
C1799 a_n2804_13878.t3 gnd 0.194556f
C1800 a_n2804_13878.n7 gnd 1.53196f
C1801 a_n2804_13878.n8 gnd 1.04414f
C1802 a_n2804_13878.t13 gnd 0.194556f
C1803 a_n2804_13878.t1 gnd 0.194556f
C1804 a_n2804_13878.n9 gnd 1.53196f
C1805 a_n2804_13878.n10 gnd 4.90178f
C1806 a_n2804_13878.t25 gnd 1.82172f
C1807 a_n2804_13878.t28 gnd 0.194556f
C1808 a_n2804_13878.t29 gnd 0.194556f
C1809 a_n2804_13878.n11 gnd 1.37045f
C1810 a_n2804_13878.n12 gnd 1.53128f
C1811 a_n2804_13878.t24 gnd 1.81809f
C1812 a_n2804_13878.n13 gnd 0.770559f
C1813 a_n2804_13878.t27 gnd 1.81809f
C1814 a_n2804_13878.n14 gnd 0.770559f
C1815 a_n2804_13878.t30 gnd 0.194556f
C1816 a_n2804_13878.t31 gnd 0.194556f
C1817 a_n2804_13878.n15 gnd 1.37045f
C1818 a_n2804_13878.n16 gnd 0.778022f
C1819 a_n2804_13878.t26 gnd 1.81809f
C1820 a_n2804_13878.n17 gnd 2.85814f
C1821 a_n2804_13878.n18 gnd 3.74876f
C1822 a_n2804_13878.t7 gnd 0.194556f
C1823 a_n2804_13878.t16 gnd 0.194556f
C1824 a_n2804_13878.n19 gnd 1.53195f
C1825 a_n2804_13878.n20 gnd 2.50239f
C1826 a_n2804_13878.t20 gnd 0.194556f
C1827 a_n2804_13878.t6 gnd 0.194556f
C1828 a_n2804_13878.n21 gnd 1.53196f
C1829 a_n2804_13878.n22 gnd 0.678771f
C1830 a_n2804_13878.t10 gnd 0.194556f
C1831 a_n2804_13878.t11 gnd 0.194556f
C1832 a_n2804_13878.n23 gnd 1.53196f
C1833 a_n2804_13878.n24 gnd 0.678771f
C1834 a_n2804_13878.t21 gnd 0.194556f
C1835 a_n2804_13878.t22 gnd 0.194556f
C1836 a_n2804_13878.n25 gnd 1.53196f
C1837 a_n2804_13878.n26 gnd 0.678771f
C1838 a_n2804_13878.t0 gnd 0.194556f
C1839 a_n2804_13878.t12 gnd 0.194556f
C1840 a_n2804_13878.n27 gnd 1.53196f
C1841 a_n2804_13878.n28 gnd 1.37704f
C1842 a_n2804_13878.n29 gnd 1.5345f
C1843 a_n2804_13878.t23 gnd 0.194556f
C1844 vdd.t44 gnd 0.034706f
C1845 vdd.t27 gnd 0.034706f
C1846 vdd.n0 gnd 0.273732f
C1847 vdd.t3 gnd 0.034706f
C1848 vdd.t40 gnd 0.034706f
C1849 vdd.n1 gnd 0.27328f
C1850 vdd.n2 gnd 0.252016f
C1851 vdd.t23 gnd 0.034706f
C1852 vdd.t51 gnd 0.034706f
C1853 vdd.n3 gnd 0.27328f
C1854 vdd.n4 gnd 0.127454f
C1855 vdd.t49 gnd 0.034706f
C1856 vdd.t31 gnd 0.034706f
C1857 vdd.n5 gnd 0.27328f
C1858 vdd.n6 gnd 0.119592f
C1859 vdd.t55 gnd 0.034706f
C1860 vdd.t21 gnd 0.034706f
C1861 vdd.n7 gnd 0.273732f
C1862 vdd.t29 gnd 0.034706f
C1863 vdd.t47 gnd 0.034706f
C1864 vdd.n8 gnd 0.27328f
C1865 vdd.n9 gnd 0.252016f
C1866 vdd.t5 gnd 0.034706f
C1867 vdd.t9 gnd 0.034706f
C1868 vdd.n10 gnd 0.27328f
C1869 vdd.n11 gnd 0.127454f
C1870 vdd.t18 gnd 0.034706f
C1871 vdd.t36 gnd 0.034706f
C1872 vdd.n12 gnd 0.27328f
C1873 vdd.n13 gnd 0.119592f
C1874 vdd.n14 gnd 0.084549f
C1875 vdd.t272 gnd 0.019281f
C1876 vdd.t190 gnd 0.019281f
C1877 vdd.n15 gnd 0.177474f
C1878 vdd.t195 gnd 0.019281f
C1879 vdd.t192 gnd 0.019281f
C1880 vdd.n16 gnd 0.176955f
C1881 vdd.n17 gnd 0.307957f
C1882 vdd.t274 gnd 0.019281f
C1883 vdd.t188 gnd 0.019281f
C1884 vdd.n18 gnd 0.176955f
C1885 vdd.n19 gnd 0.127406f
C1886 vdd.t189 gnd 0.019281f
C1887 vdd.t186 gnd 0.019281f
C1888 vdd.n20 gnd 0.177474f
C1889 vdd.t273 gnd 0.019281f
C1890 vdd.t185 gnd 0.019281f
C1891 vdd.n21 gnd 0.176955f
C1892 vdd.n22 gnd 0.307957f
C1893 vdd.t187 gnd 0.019281f
C1894 vdd.t275 gnd 0.019281f
C1895 vdd.n23 gnd 0.176955f
C1896 vdd.n24 gnd 0.127406f
C1897 vdd.t193 gnd 0.019281f
C1898 vdd.t184 gnd 0.019281f
C1899 vdd.n25 gnd 0.176955f
C1900 vdd.t191 gnd 0.019281f
C1901 vdd.t194 gnd 0.019281f
C1902 vdd.n26 gnd 0.176955f
C1903 vdd.n27 gnd 20.5711f
C1904 vdd.n28 gnd 8.01923f
C1905 vdd.n29 gnd 0.005259f
C1906 vdd.n30 gnd 0.00488f
C1907 vdd.n31 gnd 0.002699f
C1908 vdd.n32 gnd 0.006198f
C1909 vdd.n33 gnd 0.002622f
C1910 vdd.n34 gnd 0.002776f
C1911 vdd.n35 gnd 0.00488f
C1912 vdd.n36 gnd 0.002622f
C1913 vdd.n37 gnd 0.006198f
C1914 vdd.n38 gnd 0.002776f
C1915 vdd.n39 gnd 0.00488f
C1916 vdd.n40 gnd 0.002622f
C1917 vdd.n41 gnd 0.004648f
C1918 vdd.n42 gnd 0.004662f
C1919 vdd.t122 gnd 0.013316f
C1920 vdd.n43 gnd 0.029628f
C1921 vdd.n44 gnd 0.154189f
C1922 vdd.n45 gnd 0.002622f
C1923 vdd.n46 gnd 0.002776f
C1924 vdd.n47 gnd 0.006198f
C1925 vdd.n48 gnd 0.006198f
C1926 vdd.n49 gnd 0.002776f
C1927 vdd.n50 gnd 0.002622f
C1928 vdd.n51 gnd 0.00488f
C1929 vdd.n52 gnd 0.00488f
C1930 vdd.n53 gnd 0.002622f
C1931 vdd.n54 gnd 0.002776f
C1932 vdd.n55 gnd 0.006198f
C1933 vdd.n56 gnd 0.006198f
C1934 vdd.n57 gnd 0.002776f
C1935 vdd.n58 gnd 0.002622f
C1936 vdd.n59 gnd 0.00488f
C1937 vdd.n60 gnd 0.00488f
C1938 vdd.n61 gnd 0.002622f
C1939 vdd.n62 gnd 0.002776f
C1940 vdd.n63 gnd 0.006198f
C1941 vdd.n64 gnd 0.006198f
C1942 vdd.n65 gnd 0.014653f
C1943 vdd.n66 gnd 0.002699f
C1944 vdd.n67 gnd 0.002622f
C1945 vdd.n68 gnd 0.012613f
C1946 vdd.n69 gnd 0.008806f
C1947 vdd.t96 gnd 0.03085f
C1948 vdd.t163 gnd 0.03085f
C1949 vdd.n70 gnd 0.212021f
C1950 vdd.n71 gnd 0.166722f
C1951 vdd.t76 gnd 0.03085f
C1952 vdd.t147 gnd 0.03085f
C1953 vdd.n72 gnd 0.212021f
C1954 vdd.n73 gnd 0.134544f
C1955 vdd.t77 gnd 0.03085f
C1956 vdd.t159 gnd 0.03085f
C1957 vdd.n74 gnd 0.212021f
C1958 vdd.n75 gnd 0.134544f
C1959 vdd.t110 gnd 0.03085f
C1960 vdd.t172 gnd 0.03085f
C1961 vdd.n76 gnd 0.212021f
C1962 vdd.n77 gnd 0.134544f
C1963 vdd.t125 gnd 0.03085f
C1964 vdd.t153 gnd 0.03085f
C1965 vdd.n78 gnd 0.212021f
C1966 vdd.n79 gnd 0.134544f
C1967 vdd.t100 gnd 0.03085f
C1968 vdd.t165 gnd 0.03085f
C1969 vdd.n80 gnd 0.212021f
C1970 vdd.n81 gnd 0.134544f
C1971 vdd.t115 gnd 0.03085f
C1972 vdd.t180 gnd 0.03085f
C1973 vdd.n82 gnd 0.212021f
C1974 vdd.n83 gnd 0.134544f
C1975 vdd.n84 gnd 0.005259f
C1976 vdd.n85 gnd 0.00488f
C1977 vdd.n86 gnd 0.002699f
C1978 vdd.n87 gnd 0.006198f
C1979 vdd.n88 gnd 0.002622f
C1980 vdd.n89 gnd 0.002776f
C1981 vdd.n90 gnd 0.00488f
C1982 vdd.n91 gnd 0.002622f
C1983 vdd.n92 gnd 0.006198f
C1984 vdd.n93 gnd 0.002776f
C1985 vdd.n94 gnd 0.00488f
C1986 vdd.n95 gnd 0.002622f
C1987 vdd.n96 gnd 0.004648f
C1988 vdd.n97 gnd 0.004662f
C1989 vdd.t137 gnd 0.013316f
C1990 vdd.n98 gnd 0.029628f
C1991 vdd.n99 gnd 0.154189f
C1992 vdd.n100 gnd 0.002622f
C1993 vdd.n101 gnd 0.002776f
C1994 vdd.n102 gnd 0.006198f
C1995 vdd.n103 gnd 0.006198f
C1996 vdd.n104 gnd 0.002776f
C1997 vdd.n105 gnd 0.002622f
C1998 vdd.n106 gnd 0.00488f
C1999 vdd.n107 gnd 0.00488f
C2000 vdd.n108 gnd 0.002622f
C2001 vdd.n109 gnd 0.002776f
C2002 vdd.n110 gnd 0.006198f
C2003 vdd.n111 gnd 0.006198f
C2004 vdd.n112 gnd 0.002776f
C2005 vdd.n113 gnd 0.002622f
C2006 vdd.n114 gnd 0.00488f
C2007 vdd.n115 gnd 0.00488f
C2008 vdd.n116 gnd 0.002622f
C2009 vdd.n117 gnd 0.002776f
C2010 vdd.n118 gnd 0.006198f
C2011 vdd.n119 gnd 0.006198f
C2012 vdd.n120 gnd 0.014653f
C2013 vdd.n121 gnd 0.002699f
C2014 vdd.n122 gnd 0.002622f
C2015 vdd.n123 gnd 0.012613f
C2016 vdd.n124 gnd 0.008529f
C2017 vdd.n125 gnd 0.100101f
C2018 vdd.n126 gnd 0.005259f
C2019 vdd.n127 gnd 0.00488f
C2020 vdd.n128 gnd 0.002699f
C2021 vdd.n129 gnd 0.006198f
C2022 vdd.n130 gnd 0.002622f
C2023 vdd.n131 gnd 0.002776f
C2024 vdd.n132 gnd 0.00488f
C2025 vdd.n133 gnd 0.002622f
C2026 vdd.n134 gnd 0.006198f
C2027 vdd.n135 gnd 0.002776f
C2028 vdd.n136 gnd 0.00488f
C2029 vdd.n137 gnd 0.002622f
C2030 vdd.n138 gnd 0.004648f
C2031 vdd.n139 gnd 0.004662f
C2032 vdd.t169 gnd 0.013316f
C2033 vdd.n140 gnd 0.029628f
C2034 vdd.n141 gnd 0.154189f
C2035 vdd.n142 gnd 0.002622f
C2036 vdd.n143 gnd 0.002776f
C2037 vdd.n144 gnd 0.006198f
C2038 vdd.n145 gnd 0.006198f
C2039 vdd.n146 gnd 0.002776f
C2040 vdd.n147 gnd 0.002622f
C2041 vdd.n148 gnd 0.00488f
C2042 vdd.n149 gnd 0.00488f
C2043 vdd.n150 gnd 0.002622f
C2044 vdd.n151 gnd 0.002776f
C2045 vdd.n152 gnd 0.006198f
C2046 vdd.n153 gnd 0.006198f
C2047 vdd.n154 gnd 0.002776f
C2048 vdd.n155 gnd 0.002622f
C2049 vdd.n156 gnd 0.00488f
C2050 vdd.n157 gnd 0.00488f
C2051 vdd.n158 gnd 0.002622f
C2052 vdd.n159 gnd 0.002776f
C2053 vdd.n160 gnd 0.006198f
C2054 vdd.n161 gnd 0.006198f
C2055 vdd.n162 gnd 0.014653f
C2056 vdd.n163 gnd 0.002699f
C2057 vdd.n164 gnd 0.002622f
C2058 vdd.n165 gnd 0.012613f
C2059 vdd.n166 gnd 0.008806f
C2060 vdd.t170 gnd 0.03085f
C2061 vdd.t73 gnd 0.03085f
C2062 vdd.n167 gnd 0.212021f
C2063 vdd.n168 gnd 0.166722f
C2064 vdd.t155 gnd 0.03085f
C2065 vdd.t162 gnd 0.03085f
C2066 vdd.n169 gnd 0.212021f
C2067 vdd.n170 gnd 0.134544f
C2068 vdd.t67 gnd 0.03085f
C2069 vdd.t120 gnd 0.03085f
C2070 vdd.n171 gnd 0.212021f
C2071 vdd.n172 gnd 0.134544f
C2072 vdd.t152 gnd 0.03085f
C2073 vdd.t175 gnd 0.03085f
C2074 vdd.n173 gnd 0.212021f
C2075 vdd.n174 gnd 0.134544f
C2076 vdd.t103 gnd 0.03085f
C2077 vdd.t151 gnd 0.03085f
C2078 vdd.n175 gnd 0.212021f
C2079 vdd.n176 gnd 0.134544f
C2080 vdd.t182 gnd 0.03085f
C2081 vdd.t94 gnd 0.03085f
C2082 vdd.n177 gnd 0.212021f
C2083 vdd.n178 gnd 0.134544f
C2084 vdd.t136 gnd 0.03085f
C2085 vdd.t168 gnd 0.03085f
C2086 vdd.n179 gnd 0.212021f
C2087 vdd.n180 gnd 0.134544f
C2088 vdd.n181 gnd 0.005259f
C2089 vdd.n182 gnd 0.00488f
C2090 vdd.n183 gnd 0.002699f
C2091 vdd.n184 gnd 0.006198f
C2092 vdd.n185 gnd 0.002622f
C2093 vdd.n186 gnd 0.002776f
C2094 vdd.n187 gnd 0.00488f
C2095 vdd.n188 gnd 0.002622f
C2096 vdd.n189 gnd 0.006198f
C2097 vdd.n190 gnd 0.002776f
C2098 vdd.n191 gnd 0.00488f
C2099 vdd.n192 gnd 0.002622f
C2100 vdd.n193 gnd 0.004648f
C2101 vdd.n194 gnd 0.004662f
C2102 vdd.t71 gnd 0.013316f
C2103 vdd.n195 gnd 0.029628f
C2104 vdd.n196 gnd 0.154189f
C2105 vdd.n197 gnd 0.002622f
C2106 vdd.n198 gnd 0.002776f
C2107 vdd.n199 gnd 0.006198f
C2108 vdd.n200 gnd 0.006198f
C2109 vdd.n201 gnd 0.002776f
C2110 vdd.n202 gnd 0.002622f
C2111 vdd.n203 gnd 0.00488f
C2112 vdd.n204 gnd 0.00488f
C2113 vdd.n205 gnd 0.002622f
C2114 vdd.n206 gnd 0.002776f
C2115 vdd.n207 gnd 0.006198f
C2116 vdd.n208 gnd 0.006198f
C2117 vdd.n209 gnd 0.002776f
C2118 vdd.n210 gnd 0.002622f
C2119 vdd.n211 gnd 0.00488f
C2120 vdd.n212 gnd 0.00488f
C2121 vdd.n213 gnd 0.002622f
C2122 vdd.n214 gnd 0.002776f
C2123 vdd.n215 gnd 0.006198f
C2124 vdd.n216 gnd 0.006198f
C2125 vdd.n217 gnd 0.014653f
C2126 vdd.n218 gnd 0.002699f
C2127 vdd.n219 gnd 0.002622f
C2128 vdd.n220 gnd 0.012613f
C2129 vdd.n221 gnd 0.008529f
C2130 vdd.n222 gnd 0.05955f
C2131 vdd.n223 gnd 0.214575f
C2132 vdd.n224 gnd 0.005259f
C2133 vdd.n225 gnd 0.00488f
C2134 vdd.n226 gnd 0.002699f
C2135 vdd.n227 gnd 0.006198f
C2136 vdd.n228 gnd 0.002622f
C2137 vdd.n229 gnd 0.002776f
C2138 vdd.n230 gnd 0.00488f
C2139 vdd.n231 gnd 0.002622f
C2140 vdd.n232 gnd 0.006198f
C2141 vdd.n233 gnd 0.002776f
C2142 vdd.n234 gnd 0.00488f
C2143 vdd.n235 gnd 0.002622f
C2144 vdd.n236 gnd 0.004648f
C2145 vdd.n237 gnd 0.004662f
C2146 vdd.t177 gnd 0.013316f
C2147 vdd.n238 gnd 0.029628f
C2148 vdd.n239 gnd 0.154189f
C2149 vdd.n240 gnd 0.002622f
C2150 vdd.n241 gnd 0.002776f
C2151 vdd.n242 gnd 0.006198f
C2152 vdd.n243 gnd 0.006198f
C2153 vdd.n244 gnd 0.002776f
C2154 vdd.n245 gnd 0.002622f
C2155 vdd.n246 gnd 0.00488f
C2156 vdd.n247 gnd 0.00488f
C2157 vdd.n248 gnd 0.002622f
C2158 vdd.n249 gnd 0.002776f
C2159 vdd.n250 gnd 0.006198f
C2160 vdd.n251 gnd 0.006198f
C2161 vdd.n252 gnd 0.002776f
C2162 vdd.n253 gnd 0.002622f
C2163 vdd.n254 gnd 0.00488f
C2164 vdd.n255 gnd 0.00488f
C2165 vdd.n256 gnd 0.002622f
C2166 vdd.n257 gnd 0.002776f
C2167 vdd.n258 gnd 0.006198f
C2168 vdd.n259 gnd 0.006198f
C2169 vdd.n260 gnd 0.014653f
C2170 vdd.n261 gnd 0.002699f
C2171 vdd.n262 gnd 0.002622f
C2172 vdd.n263 gnd 0.012613f
C2173 vdd.n264 gnd 0.008806f
C2174 vdd.t179 gnd 0.03085f
C2175 vdd.t78 gnd 0.03085f
C2176 vdd.n265 gnd 0.212021f
C2177 vdd.n266 gnd 0.166722f
C2178 vdd.t161 gnd 0.03085f
C2179 vdd.t174 gnd 0.03085f
C2180 vdd.n267 gnd 0.212021f
C2181 vdd.n268 gnd 0.134544f
C2182 vdd.t85 gnd 0.03085f
C2183 vdd.t138 gnd 0.03085f
C2184 vdd.n269 gnd 0.212021f
C2185 vdd.n270 gnd 0.134544f
C2186 vdd.t160 gnd 0.03085f
C2187 vdd.t61 gnd 0.03085f
C2188 vdd.n271 gnd 0.212021f
C2189 vdd.n272 gnd 0.134544f
C2190 vdd.t113 gnd 0.03085f
C2191 vdd.t158 gnd 0.03085f
C2192 vdd.n273 gnd 0.212021f
C2193 vdd.n274 gnd 0.134544f
C2194 vdd.t69 gnd 0.03085f
C2195 vdd.t112 gnd 0.03085f
C2196 vdd.n275 gnd 0.212021f
C2197 vdd.n276 gnd 0.134544f
C2198 vdd.t143 gnd 0.03085f
C2199 vdd.t178 gnd 0.03085f
C2200 vdd.n277 gnd 0.212021f
C2201 vdd.n278 gnd 0.134544f
C2202 vdd.n279 gnd 0.005259f
C2203 vdd.n280 gnd 0.00488f
C2204 vdd.n281 gnd 0.002699f
C2205 vdd.n282 gnd 0.006198f
C2206 vdd.n283 gnd 0.002622f
C2207 vdd.n284 gnd 0.002776f
C2208 vdd.n285 gnd 0.00488f
C2209 vdd.n286 gnd 0.002622f
C2210 vdd.n287 gnd 0.006198f
C2211 vdd.n288 gnd 0.002776f
C2212 vdd.n289 gnd 0.00488f
C2213 vdd.n290 gnd 0.002622f
C2214 vdd.n291 gnd 0.004648f
C2215 vdd.n292 gnd 0.004662f
C2216 vdd.t88 gnd 0.013316f
C2217 vdd.n293 gnd 0.029628f
C2218 vdd.n294 gnd 0.154189f
C2219 vdd.n295 gnd 0.002622f
C2220 vdd.n296 gnd 0.002776f
C2221 vdd.n297 gnd 0.006198f
C2222 vdd.n298 gnd 0.006198f
C2223 vdd.n299 gnd 0.002776f
C2224 vdd.n300 gnd 0.002622f
C2225 vdd.n301 gnd 0.00488f
C2226 vdd.n302 gnd 0.00488f
C2227 vdd.n303 gnd 0.002622f
C2228 vdd.n304 gnd 0.002776f
C2229 vdd.n305 gnd 0.006198f
C2230 vdd.n306 gnd 0.006198f
C2231 vdd.n307 gnd 0.002776f
C2232 vdd.n308 gnd 0.002622f
C2233 vdd.n309 gnd 0.00488f
C2234 vdd.n310 gnd 0.00488f
C2235 vdd.n311 gnd 0.002622f
C2236 vdd.n312 gnd 0.002776f
C2237 vdd.n313 gnd 0.006198f
C2238 vdd.n314 gnd 0.006198f
C2239 vdd.n315 gnd 0.014653f
C2240 vdd.n316 gnd 0.002699f
C2241 vdd.n317 gnd 0.002622f
C2242 vdd.n318 gnd 0.012613f
C2243 vdd.n319 gnd 0.008529f
C2244 vdd.n320 gnd 0.05955f
C2245 vdd.n321 gnd 0.240295f
C2246 vdd.n322 gnd 0.007364f
C2247 vdd.n323 gnd 0.009582f
C2248 vdd.n324 gnd 0.007712f
C2249 vdd.n325 gnd 0.007712f
C2250 vdd.n326 gnd 0.009582f
C2251 vdd.n327 gnd 0.009582f
C2252 vdd.n328 gnd 0.700161f
C2253 vdd.n329 gnd 0.009582f
C2254 vdd.n330 gnd 0.009582f
C2255 vdd.n331 gnd 0.009582f
C2256 vdd.n332 gnd 0.758916f
C2257 vdd.n333 gnd 0.009582f
C2258 vdd.n334 gnd 0.009582f
C2259 vdd.n335 gnd 0.009582f
C2260 vdd.n336 gnd 0.009582f
C2261 vdd.n337 gnd 0.007712f
C2262 vdd.n338 gnd 0.009582f
C2263 vdd.t150 gnd 0.489623f
C2264 vdd.n339 gnd 0.009582f
C2265 vdd.n340 gnd 0.009582f
C2266 vdd.n341 gnd 0.009582f
C2267 vdd.t93 gnd 0.489623f
C2268 vdd.n342 gnd 0.009582f
C2269 vdd.n343 gnd 0.009582f
C2270 vdd.n344 gnd 0.009582f
C2271 vdd.n345 gnd 0.009582f
C2272 vdd.n346 gnd 0.009582f
C2273 vdd.n347 gnd 0.007712f
C2274 vdd.n348 gnd 0.009582f
C2275 vdd.n349 gnd 0.553274f
C2276 vdd.n350 gnd 0.009582f
C2277 vdd.n351 gnd 0.009582f
C2278 vdd.n352 gnd 0.009582f
C2279 vdd.t167 gnd 0.489623f
C2280 vdd.n353 gnd 0.009582f
C2281 vdd.n354 gnd 0.009582f
C2282 vdd.n355 gnd 0.009582f
C2283 vdd.n356 gnd 0.009582f
C2284 vdd.n357 gnd 0.009582f
C2285 vdd.n358 gnd 0.007712f
C2286 vdd.n359 gnd 0.009582f
C2287 vdd.t70 gnd 0.489623f
C2288 vdd.n360 gnd 0.009582f
C2289 vdd.n361 gnd 0.009582f
C2290 vdd.n362 gnd 0.009582f
C2291 vdd.n363 gnd 0.827463f
C2292 vdd.n364 gnd 0.009582f
C2293 vdd.n365 gnd 0.009582f
C2294 vdd.n366 gnd 0.009582f
C2295 vdd.n367 gnd 0.009582f
C2296 vdd.n368 gnd 0.009582f
C2297 vdd.n369 gnd 0.006401f
C2298 vdd.n370 gnd 0.021821f
C2299 vdd.t215 gnd 0.489623f
C2300 vdd.n371 gnd 0.009582f
C2301 vdd.n372 gnd 0.021821f
C2302 vdd.n404 gnd 0.009582f
C2303 vdd.t240 gnd 0.117885f
C2304 vdd.t239 gnd 0.125987f
C2305 vdd.t238 gnd 0.153957f
C2306 vdd.n405 gnd 0.19735f
C2307 vdd.n406 gnd 0.166581f
C2308 vdd.n407 gnd 0.012648f
C2309 vdd.n408 gnd 0.009582f
C2310 vdd.n409 gnd 0.007712f
C2311 vdd.n410 gnd 0.009582f
C2312 vdd.n411 gnd 0.007712f
C2313 vdd.n412 gnd 0.009582f
C2314 vdd.n413 gnd 0.007712f
C2315 vdd.n414 gnd 0.009582f
C2316 vdd.n415 gnd 0.007712f
C2317 vdd.n416 gnd 0.009582f
C2318 vdd.n417 gnd 0.007712f
C2319 vdd.n418 gnd 0.009582f
C2320 vdd.t217 gnd 0.117885f
C2321 vdd.t216 gnd 0.125987f
C2322 vdd.t214 gnd 0.153957f
C2323 vdd.n419 gnd 0.19735f
C2324 vdd.n420 gnd 0.166581f
C2325 vdd.n421 gnd 0.007712f
C2326 vdd.n422 gnd 0.009582f
C2327 vdd.n423 gnd 0.007712f
C2328 vdd.n424 gnd 0.009582f
C2329 vdd.n425 gnd 0.007712f
C2330 vdd.n426 gnd 0.009582f
C2331 vdd.n427 gnd 0.007712f
C2332 vdd.n428 gnd 0.009582f
C2333 vdd.n429 gnd 0.007712f
C2334 vdd.n430 gnd 0.009582f
C2335 vdd.t231 gnd 0.117885f
C2336 vdd.t230 gnd 0.125987f
C2337 vdd.t229 gnd 0.153957f
C2338 vdd.n431 gnd 0.19735f
C2339 vdd.n432 gnd 0.166581f
C2340 vdd.n433 gnd 0.016505f
C2341 vdd.n434 gnd 0.009582f
C2342 vdd.n435 gnd 0.007712f
C2343 vdd.n436 gnd 0.009582f
C2344 vdd.n437 gnd 0.007712f
C2345 vdd.n438 gnd 0.009582f
C2346 vdd.n439 gnd 0.007712f
C2347 vdd.n440 gnd 0.009582f
C2348 vdd.n441 gnd 0.007712f
C2349 vdd.n442 gnd 0.009582f
C2350 vdd.n443 gnd 0.021821f
C2351 vdd.n444 gnd 0.02197f
C2352 vdd.n445 gnd 0.02197f
C2353 vdd.n446 gnd 0.006401f
C2354 vdd.n447 gnd 0.007712f
C2355 vdd.n448 gnd 0.009582f
C2356 vdd.n449 gnd 0.009582f
C2357 vdd.n450 gnd 0.007712f
C2358 vdd.n451 gnd 0.009582f
C2359 vdd.n452 gnd 0.009582f
C2360 vdd.n453 gnd 0.009582f
C2361 vdd.n454 gnd 0.009582f
C2362 vdd.n455 gnd 0.009582f
C2363 vdd.n456 gnd 0.007712f
C2364 vdd.n457 gnd 0.007712f
C2365 vdd.n458 gnd 0.009582f
C2366 vdd.n459 gnd 0.009582f
C2367 vdd.n460 gnd 0.007712f
C2368 vdd.n461 gnd 0.009582f
C2369 vdd.n462 gnd 0.009582f
C2370 vdd.n463 gnd 0.009582f
C2371 vdd.n464 gnd 0.009582f
C2372 vdd.n465 gnd 0.009582f
C2373 vdd.n466 gnd 0.007712f
C2374 vdd.n467 gnd 0.007712f
C2375 vdd.n468 gnd 0.009582f
C2376 vdd.n469 gnd 0.009582f
C2377 vdd.n470 gnd 0.007712f
C2378 vdd.n471 gnd 0.009582f
C2379 vdd.n472 gnd 0.009582f
C2380 vdd.n473 gnd 0.009582f
C2381 vdd.n474 gnd 0.009582f
C2382 vdd.n475 gnd 0.009582f
C2383 vdd.n476 gnd 0.007712f
C2384 vdd.n477 gnd 0.007712f
C2385 vdd.n478 gnd 0.009582f
C2386 vdd.n479 gnd 0.009582f
C2387 vdd.n480 gnd 0.007712f
C2388 vdd.n481 gnd 0.009582f
C2389 vdd.n482 gnd 0.009582f
C2390 vdd.n483 gnd 0.009582f
C2391 vdd.n484 gnd 0.009582f
C2392 vdd.n485 gnd 0.009582f
C2393 vdd.n486 gnd 0.007712f
C2394 vdd.n487 gnd 0.007712f
C2395 vdd.n488 gnd 0.009582f
C2396 vdd.n489 gnd 0.009582f
C2397 vdd.n490 gnd 0.00644f
C2398 vdd.n491 gnd 0.009582f
C2399 vdd.n492 gnd 0.009582f
C2400 vdd.n493 gnd 0.009582f
C2401 vdd.n494 gnd 0.009582f
C2402 vdd.n495 gnd 0.009582f
C2403 vdd.n496 gnd 0.00644f
C2404 vdd.n497 gnd 0.007712f
C2405 vdd.n498 gnd 0.009582f
C2406 vdd.n499 gnd 0.009582f
C2407 vdd.n500 gnd 0.007712f
C2408 vdd.n501 gnd 0.009582f
C2409 vdd.n502 gnd 0.009582f
C2410 vdd.n503 gnd 0.009582f
C2411 vdd.n504 gnd 0.009582f
C2412 vdd.n505 gnd 0.009582f
C2413 vdd.n506 gnd 0.007712f
C2414 vdd.n507 gnd 0.007712f
C2415 vdd.n508 gnd 0.009582f
C2416 vdd.n509 gnd 0.009582f
C2417 vdd.n510 gnd 0.007712f
C2418 vdd.n511 gnd 0.009582f
C2419 vdd.n512 gnd 0.009582f
C2420 vdd.n513 gnd 0.009582f
C2421 vdd.n514 gnd 0.009582f
C2422 vdd.n515 gnd 0.009582f
C2423 vdd.n516 gnd 0.007712f
C2424 vdd.n517 gnd 0.007712f
C2425 vdd.n518 gnd 0.009582f
C2426 vdd.n519 gnd 0.009582f
C2427 vdd.n520 gnd 0.007712f
C2428 vdd.n521 gnd 0.009582f
C2429 vdd.n522 gnd 0.009582f
C2430 vdd.n523 gnd 0.009582f
C2431 vdd.n524 gnd 0.009582f
C2432 vdd.n525 gnd 0.009582f
C2433 vdd.n526 gnd 0.007712f
C2434 vdd.n527 gnd 0.007712f
C2435 vdd.n528 gnd 0.009582f
C2436 vdd.n529 gnd 0.009582f
C2437 vdd.n530 gnd 0.007712f
C2438 vdd.n531 gnd 0.009582f
C2439 vdd.n532 gnd 0.009582f
C2440 vdd.n533 gnd 0.009582f
C2441 vdd.n534 gnd 0.009582f
C2442 vdd.n535 gnd 0.009582f
C2443 vdd.n536 gnd 0.007712f
C2444 vdd.n537 gnd 0.007712f
C2445 vdd.n538 gnd 0.009582f
C2446 vdd.n539 gnd 0.009582f
C2447 vdd.n540 gnd 0.007712f
C2448 vdd.n541 gnd 0.009582f
C2449 vdd.n542 gnd 0.009582f
C2450 vdd.n543 gnd 0.009582f
C2451 vdd.n544 gnd 0.009582f
C2452 vdd.n545 gnd 0.009582f
C2453 vdd.n546 gnd 0.005244f
C2454 vdd.n547 gnd 0.016505f
C2455 vdd.n548 gnd 0.009582f
C2456 vdd.n549 gnd 0.009582f
C2457 vdd.n550 gnd 0.007635f
C2458 vdd.n551 gnd 0.009582f
C2459 vdd.n552 gnd 0.009582f
C2460 vdd.n553 gnd 0.009582f
C2461 vdd.n554 gnd 0.009582f
C2462 vdd.n555 gnd 0.009582f
C2463 vdd.n556 gnd 0.007712f
C2464 vdd.n557 gnd 0.007712f
C2465 vdd.n558 gnd 0.009582f
C2466 vdd.n559 gnd 0.009582f
C2467 vdd.n560 gnd 0.007712f
C2468 vdd.n561 gnd 0.009582f
C2469 vdd.n562 gnd 0.009582f
C2470 vdd.n563 gnd 0.009582f
C2471 vdd.n564 gnd 0.009582f
C2472 vdd.n565 gnd 0.009582f
C2473 vdd.n566 gnd 0.007712f
C2474 vdd.n567 gnd 0.007712f
C2475 vdd.n568 gnd 0.009582f
C2476 vdd.n569 gnd 0.009582f
C2477 vdd.n570 gnd 0.007712f
C2478 vdd.n571 gnd 0.009582f
C2479 vdd.n572 gnd 0.009582f
C2480 vdd.n573 gnd 0.009582f
C2481 vdd.n574 gnd 0.009582f
C2482 vdd.n575 gnd 0.009582f
C2483 vdd.n576 gnd 0.007712f
C2484 vdd.n577 gnd 0.007712f
C2485 vdd.n578 gnd 0.009582f
C2486 vdd.n579 gnd 0.009582f
C2487 vdd.n580 gnd 0.007712f
C2488 vdd.n581 gnd 0.009582f
C2489 vdd.n582 gnd 0.009582f
C2490 vdd.n583 gnd 0.009582f
C2491 vdd.n584 gnd 0.009582f
C2492 vdd.n585 gnd 0.009582f
C2493 vdd.n586 gnd 0.007712f
C2494 vdd.n587 gnd 0.007712f
C2495 vdd.n588 gnd 0.009582f
C2496 vdd.n589 gnd 0.009582f
C2497 vdd.n590 gnd 0.007712f
C2498 vdd.n591 gnd 0.009582f
C2499 vdd.n592 gnd 0.009582f
C2500 vdd.n593 gnd 0.009582f
C2501 vdd.n594 gnd 0.009582f
C2502 vdd.n595 gnd 0.009582f
C2503 vdd.n596 gnd 0.007712f
C2504 vdd.n597 gnd 0.009582f
C2505 vdd.n598 gnd 0.007712f
C2506 vdd.n599 gnd 0.004049f
C2507 vdd.n600 gnd 0.009582f
C2508 vdd.n601 gnd 0.009582f
C2509 vdd.n602 gnd 0.007712f
C2510 vdd.n603 gnd 0.009582f
C2511 vdd.n604 gnd 0.007712f
C2512 vdd.n605 gnd 0.009582f
C2513 vdd.n606 gnd 0.007712f
C2514 vdd.n607 gnd 0.009582f
C2515 vdd.n608 gnd 0.007712f
C2516 vdd.n609 gnd 0.009582f
C2517 vdd.n610 gnd 0.007712f
C2518 vdd.n611 gnd 0.009582f
C2519 vdd.n612 gnd 0.009582f
C2520 vdd.n613 gnd 0.533689f
C2521 vdd.t109 gnd 0.489623f
C2522 vdd.n614 gnd 0.009582f
C2523 vdd.n615 gnd 0.007712f
C2524 vdd.n616 gnd 0.009582f
C2525 vdd.n617 gnd 0.007712f
C2526 vdd.n618 gnd 0.009582f
C2527 vdd.t66 gnd 0.489623f
C2528 vdd.n619 gnd 0.009582f
C2529 vdd.n620 gnd 0.007712f
C2530 vdd.n621 gnd 0.009582f
C2531 vdd.n622 gnd 0.007712f
C2532 vdd.n623 gnd 0.009582f
C2533 vdd.t146 gnd 0.489623f
C2534 vdd.n624 gnd 0.612029f
C2535 vdd.n625 gnd 0.009582f
C2536 vdd.n626 gnd 0.007712f
C2537 vdd.n627 gnd 0.009582f
C2538 vdd.n628 gnd 0.007712f
C2539 vdd.n629 gnd 0.009582f
C2540 vdd.t75 gnd 0.489623f
C2541 vdd.n630 gnd 0.009582f
C2542 vdd.n631 gnd 0.007712f
C2543 vdd.n632 gnd 0.009582f
C2544 vdd.n633 gnd 0.007712f
C2545 vdd.n634 gnd 0.009582f
C2546 vdd.n635 gnd 0.680576f
C2547 vdd.n636 gnd 0.812775f
C2548 vdd.t72 gnd 0.489623f
C2549 vdd.n637 gnd 0.009582f
C2550 vdd.n638 gnd 0.007712f
C2551 vdd.n639 gnd 0.009582f
C2552 vdd.n640 gnd 0.007712f
C2553 vdd.n641 gnd 0.009582f
C2554 vdd.n642 gnd 0.514104f
C2555 vdd.n643 gnd 0.009582f
C2556 vdd.n644 gnd 0.007712f
C2557 vdd.n645 gnd 0.009582f
C2558 vdd.n646 gnd 0.007712f
C2559 vdd.n647 gnd 0.009582f
C2560 vdd.n648 gnd 0.979246f
C2561 vdd.t121 gnd 0.489623f
C2562 vdd.n649 gnd 0.009582f
C2563 vdd.n650 gnd 0.007712f
C2564 vdd.n651 gnd 0.009582f
C2565 vdd.n652 gnd 0.007712f
C2566 vdd.n653 gnd 0.009582f
C2567 vdd.t219 gnd 0.489623f
C2568 vdd.n654 gnd 0.009582f
C2569 vdd.n655 gnd 0.007712f
C2570 vdd.n656 gnd 0.02197f
C2571 vdd.n657 gnd 0.02197f
C2572 vdd.n658 gnd 11.799901f
C2573 vdd.n659 gnd 0.543482f
C2574 vdd.n660 gnd 0.02197f
C2575 vdd.n661 gnd 0.008241f
C2576 vdd.n662 gnd 0.007712f
C2577 vdd.n667 gnd 0.006133f
C2578 vdd.n668 gnd 0.007712f
C2579 vdd.n669 gnd 0.009582f
C2580 vdd.n670 gnd 0.009582f
C2581 vdd.n671 gnd 0.009582f
C2582 vdd.n672 gnd 0.009582f
C2583 vdd.n673 gnd 0.009582f
C2584 vdd.n674 gnd 0.007712f
C2585 vdd.n675 gnd 0.009582f
C2586 vdd.n676 gnd 0.009582f
C2587 vdd.n677 gnd 0.009582f
C2588 vdd.n678 gnd 0.009582f
C2589 vdd.n679 gnd 0.009582f
C2590 vdd.n680 gnd 0.007712f
C2591 vdd.n681 gnd 0.009582f
C2592 vdd.n682 gnd 0.009582f
C2593 vdd.n683 gnd 0.009582f
C2594 vdd.n684 gnd 0.009582f
C2595 vdd.n685 gnd 0.009582f
C2596 vdd.t250 gnd 0.117885f
C2597 vdd.t251 gnd 0.125987f
C2598 vdd.t249 gnd 0.153957f
C2599 vdd.n686 gnd 0.19735f
C2600 vdd.n687 gnd 0.16581f
C2601 vdd.n688 gnd 0.015733f
C2602 vdd.n689 gnd 0.009582f
C2603 vdd.n690 gnd 0.009582f
C2604 vdd.n691 gnd 0.009582f
C2605 vdd.n692 gnd 0.009582f
C2606 vdd.n693 gnd 0.009582f
C2607 vdd.n694 gnd 0.007712f
C2608 vdd.n695 gnd 0.009582f
C2609 vdd.n696 gnd 0.009582f
C2610 vdd.n697 gnd 0.009582f
C2611 vdd.n698 gnd 0.009582f
C2612 vdd.n699 gnd 0.009582f
C2613 vdd.n700 gnd 0.007712f
C2614 vdd.n701 gnd 0.009582f
C2615 vdd.n702 gnd 0.009582f
C2616 vdd.n703 gnd 0.009582f
C2617 vdd.n704 gnd 0.009582f
C2618 vdd.n705 gnd 0.009582f
C2619 vdd.n706 gnd 0.007712f
C2620 vdd.n707 gnd 0.009582f
C2621 vdd.n708 gnd 0.009582f
C2622 vdd.n709 gnd 0.009582f
C2623 vdd.n710 gnd 0.009582f
C2624 vdd.n711 gnd 0.009582f
C2625 vdd.n712 gnd 0.007712f
C2626 vdd.n713 gnd 0.009582f
C2627 vdd.n714 gnd 0.009582f
C2628 vdd.n715 gnd 0.009582f
C2629 vdd.n716 gnd 0.009582f
C2630 vdd.n717 gnd 0.009582f
C2631 vdd.n718 gnd 0.007712f
C2632 vdd.n719 gnd 0.009582f
C2633 vdd.n720 gnd 0.009582f
C2634 vdd.n721 gnd 0.009582f
C2635 vdd.n722 gnd 0.007635f
C2636 vdd.t233 gnd 0.117885f
C2637 vdd.t234 gnd 0.125987f
C2638 vdd.t232 gnd 0.153957f
C2639 vdd.n723 gnd 0.19735f
C2640 vdd.n724 gnd 0.16581f
C2641 vdd.n725 gnd 0.009582f
C2642 vdd.n726 gnd 0.007712f
C2643 vdd.n728 gnd 0.009582f
C2644 vdd.n730 gnd 0.009582f
C2645 vdd.n731 gnd 0.009582f
C2646 vdd.n732 gnd 0.007712f
C2647 vdd.n733 gnd 0.009582f
C2648 vdd.n734 gnd 0.009582f
C2649 vdd.n735 gnd 0.009582f
C2650 vdd.n736 gnd 0.009582f
C2651 vdd.n737 gnd 0.009582f
C2652 vdd.n738 gnd 0.007712f
C2653 vdd.n739 gnd 0.009582f
C2654 vdd.n740 gnd 0.009582f
C2655 vdd.n741 gnd 0.009582f
C2656 vdd.n742 gnd 0.009582f
C2657 vdd.n743 gnd 0.009582f
C2658 vdd.n744 gnd 0.007712f
C2659 vdd.n745 gnd 0.009582f
C2660 vdd.n746 gnd 0.009582f
C2661 vdd.n747 gnd 0.009582f
C2662 vdd.n748 gnd 0.006133f
C2663 vdd.n753 gnd 0.006516f
C2664 vdd.n754 gnd 0.006516f
C2665 vdd.n755 gnd 0.006516f
C2666 vdd.n756 gnd 11.5649f
C2667 vdd.n757 gnd 0.006516f
C2668 vdd.n758 gnd 0.006516f
C2669 vdd.n759 gnd 0.006516f
C2670 vdd.n761 gnd 0.006516f
C2671 vdd.n762 gnd 0.006516f
C2672 vdd.n764 gnd 0.006516f
C2673 vdd.n765 gnd 0.004743f
C2674 vdd.n767 gnd 0.006516f
C2675 vdd.t199 gnd 0.263304f
C2676 vdd.t198 gnd 0.269524f
C2677 vdd.t196 gnd 0.171895f
C2678 vdd.n768 gnd 0.0929f
C2679 vdd.n769 gnd 0.052696f
C2680 vdd.n770 gnd 0.009312f
C2681 vdd.n771 gnd 0.014795f
C2682 vdd.n773 gnd 0.006516f
C2683 vdd.n774 gnd 0.665888f
C2684 vdd.n775 gnd 0.013951f
C2685 vdd.n776 gnd 0.013951f
C2686 vdd.n777 gnd 0.006516f
C2687 vdd.n778 gnd 0.014795f
C2688 vdd.n779 gnd 0.006516f
C2689 vdd.n780 gnd 0.006516f
C2690 vdd.n781 gnd 0.006516f
C2691 vdd.n782 gnd 0.006516f
C2692 vdd.n783 gnd 0.006516f
C2693 vdd.n785 gnd 0.006516f
C2694 vdd.n786 gnd 0.006516f
C2695 vdd.n788 gnd 0.006516f
C2696 vdd.n789 gnd 0.006516f
C2697 vdd.n791 gnd 0.006516f
C2698 vdd.n792 gnd 0.006516f
C2699 vdd.n794 gnd 0.006516f
C2700 vdd.n795 gnd 0.006516f
C2701 vdd.n797 gnd 0.006516f
C2702 vdd.n798 gnd 0.006516f
C2703 vdd.n800 gnd 0.006516f
C2704 vdd.n801 gnd 0.004743f
C2705 vdd.n803 gnd 0.006516f
C2706 vdd.t213 gnd 0.263304f
C2707 vdd.t212 gnd 0.269524f
C2708 vdd.t211 gnd 0.171895f
C2709 vdd.n804 gnd 0.0929f
C2710 vdd.n805 gnd 0.052696f
C2711 vdd.n806 gnd 0.009312f
C2712 vdd.n807 gnd 0.006516f
C2713 vdd.n808 gnd 0.006516f
C2714 vdd.t197 gnd 0.332944f
C2715 vdd.n809 gnd 0.006516f
C2716 vdd.n810 gnd 0.006516f
C2717 vdd.n811 gnd 0.006516f
C2718 vdd.n812 gnd 0.006516f
C2719 vdd.n813 gnd 0.006516f
C2720 vdd.n814 gnd 0.665888f
C2721 vdd.n815 gnd 0.006516f
C2722 vdd.n816 gnd 0.006516f
C2723 vdd.n817 gnd 0.523897f
C2724 vdd.n818 gnd 0.006516f
C2725 vdd.n819 gnd 0.006516f
C2726 vdd.n820 gnd 0.006516f
C2727 vdd.n821 gnd 0.006516f
C2728 vdd.n822 gnd 0.665888f
C2729 vdd.n823 gnd 0.006516f
C2730 vdd.n824 gnd 0.006516f
C2731 vdd.n825 gnd 0.006516f
C2732 vdd.n826 gnd 0.006516f
C2733 vdd.n827 gnd 0.006516f
C2734 vdd.t16 gnd 0.332944f
C2735 vdd.n828 gnd 0.006516f
C2736 vdd.n829 gnd 0.006516f
C2737 vdd.n830 gnd 0.006516f
C2738 vdd.n831 gnd 0.006516f
C2739 vdd.n832 gnd 0.006516f
C2740 vdd.t33 gnd 0.332944f
C2741 vdd.n833 gnd 0.006516f
C2742 vdd.n834 gnd 0.006516f
C2743 vdd.n835 gnd 0.641406f
C2744 vdd.n836 gnd 0.006516f
C2745 vdd.n837 gnd 0.006516f
C2746 vdd.n838 gnd 0.006516f
C2747 vdd.t32 gnd 0.332944f
C2748 vdd.n839 gnd 0.006516f
C2749 vdd.n840 gnd 0.006516f
C2750 vdd.n841 gnd 0.494519f
C2751 vdd.n842 gnd 0.006516f
C2752 vdd.n843 gnd 0.006516f
C2753 vdd.n844 gnd 0.006516f
C2754 vdd.n845 gnd 0.465142f
C2755 vdd.n846 gnd 0.006516f
C2756 vdd.n847 gnd 0.006516f
C2757 vdd.n848 gnd 0.347632f
C2758 vdd.n849 gnd 0.006516f
C2759 vdd.n850 gnd 0.006516f
C2760 vdd.n851 gnd 0.006516f
C2761 vdd.n852 gnd 0.612029f
C2762 vdd.n853 gnd 0.006516f
C2763 vdd.n854 gnd 0.006516f
C2764 vdd.t37 gnd 0.332944f
C2765 vdd.n855 gnd 0.006516f
C2766 vdd.n856 gnd 0.006516f
C2767 vdd.n857 gnd 0.006516f
C2768 vdd.n858 gnd 0.665888f
C2769 vdd.n859 gnd 0.006516f
C2770 vdd.n860 gnd 0.006516f
C2771 vdd.t38 gnd 0.332944f
C2772 vdd.n861 gnd 0.006516f
C2773 vdd.n862 gnd 0.006516f
C2774 vdd.n863 gnd 0.006516f
C2775 vdd.t10 gnd 0.332944f
C2776 vdd.n864 gnd 0.006516f
C2777 vdd.n865 gnd 0.006516f
C2778 vdd.n866 gnd 0.006516f
C2779 vdd.t224 gnd 0.269524f
C2780 vdd.t222 gnd 0.171895f
C2781 vdd.t225 gnd 0.269524f
C2782 vdd.n867 gnd 0.151484f
C2783 vdd.n868 gnd 0.018876f
C2784 vdd.n869 gnd 0.006516f
C2785 vdd.t223 gnd 0.239915f
C2786 vdd.n870 gnd 0.006516f
C2787 vdd.n871 gnd 0.006516f
C2788 vdd.n872 gnd 0.572859f
C2789 vdd.n873 gnd 0.006516f
C2790 vdd.n874 gnd 0.006516f
C2791 vdd.n875 gnd 0.006516f
C2792 vdd.n876 gnd 0.386802f
C2793 vdd.n877 gnd 0.006516f
C2794 vdd.n878 gnd 0.006516f
C2795 vdd.t11 gnd 0.137094f
C2796 vdd.n879 gnd 0.425972f
C2797 vdd.n880 gnd 0.006516f
C2798 vdd.n881 gnd 0.006516f
C2799 vdd.n882 gnd 0.006516f
C2800 vdd.n883 gnd 0.533689f
C2801 vdd.n884 gnd 0.006516f
C2802 vdd.n885 gnd 0.006516f
C2803 vdd.t24 gnd 0.332944f
C2804 vdd.n886 gnd 0.006516f
C2805 vdd.n887 gnd 0.006516f
C2806 vdd.n888 gnd 0.006516f
C2807 vdd.t20 gnd 0.332944f
C2808 vdd.n889 gnd 0.006516f
C2809 vdd.n890 gnd 0.006516f
C2810 vdd.t41 gnd 0.332944f
C2811 vdd.n891 gnd 0.006516f
C2812 vdd.n892 gnd 0.006516f
C2813 vdd.n893 gnd 0.006516f
C2814 vdd.t0 gnd 0.225227f
C2815 vdd.n894 gnd 0.006516f
C2816 vdd.n895 gnd 0.006516f
C2817 vdd.n896 gnd 0.587548f
C2818 vdd.n897 gnd 0.006516f
C2819 vdd.n898 gnd 0.006516f
C2820 vdd.n899 gnd 0.006516f
C2821 vdd.t42 gnd 0.332944f
C2822 vdd.n900 gnd 0.006516f
C2823 vdd.n901 gnd 0.006516f
C2824 vdd.t54 gnd 0.318255f
C2825 vdd.n902 gnd 0.440661f
C2826 vdd.n903 gnd 0.006516f
C2827 vdd.n904 gnd 0.006516f
C2828 vdd.n905 gnd 0.006516f
C2829 vdd.t6 gnd 0.332944f
C2830 vdd.n906 gnd 0.006516f
C2831 vdd.n907 gnd 0.006516f
C2832 vdd.t46 gnd 0.332944f
C2833 vdd.n908 gnd 0.006516f
C2834 vdd.n909 gnd 0.006516f
C2835 vdd.n910 gnd 0.006516f
C2836 vdd.n911 gnd 0.665888f
C2837 vdd.n912 gnd 0.006516f
C2838 vdd.n913 gnd 0.006516f
C2839 vdd.t28 gnd 0.332944f
C2840 vdd.n914 gnd 0.006516f
C2841 vdd.n915 gnd 0.006516f
C2842 vdd.n916 gnd 0.006516f
C2843 vdd.n917 gnd 0.460246f
C2844 vdd.n918 gnd 0.006516f
C2845 vdd.n919 gnd 0.006516f
C2846 vdd.n920 gnd 0.006516f
C2847 vdd.n921 gnd 0.006516f
C2848 vdd.n922 gnd 0.006516f
C2849 vdd.t253 gnd 0.332944f
C2850 vdd.n923 gnd 0.006516f
C2851 vdd.n924 gnd 0.006516f
C2852 vdd.t8 gnd 0.332944f
C2853 vdd.n925 gnd 0.006516f
C2854 vdd.n926 gnd 0.013951f
C2855 vdd.n927 gnd 0.013951f
C2856 vdd.n928 gnd 0.75402f
C2857 vdd.n929 gnd 0.006516f
C2858 vdd.n930 gnd 0.006516f
C2859 vdd.t4 gnd 0.332944f
C2860 vdd.n931 gnd 0.013951f
C2861 vdd.n932 gnd 0.006516f
C2862 vdd.n933 gnd 0.006516f
C2863 vdd.t48 gnd 0.567963f
C2864 vdd.n951 gnd 0.014795f
C2865 vdd.n969 gnd 0.013951f
C2866 vdd.n970 gnd 0.006516f
C2867 vdd.n971 gnd 0.013951f
C2868 vdd.t271 gnd 0.263304f
C2869 vdd.t270 gnd 0.269524f
C2870 vdd.t269 gnd 0.171895f
C2871 vdd.n972 gnd 0.0929f
C2872 vdd.n973 gnd 0.052696f
C2873 vdd.n974 gnd 0.014795f
C2874 vdd.n975 gnd 0.006516f
C2875 vdd.n976 gnd 0.391699f
C2876 vdd.n977 gnd 0.013951f
C2877 vdd.n978 gnd 0.006516f
C2878 vdd.n979 gnd 0.014795f
C2879 vdd.n980 gnd 0.006516f
C2880 vdd.t248 gnd 0.263304f
C2881 vdd.t247 gnd 0.269524f
C2882 vdd.t245 gnd 0.171895f
C2883 vdd.n981 gnd 0.0929f
C2884 vdd.n982 gnd 0.052696f
C2885 vdd.n983 gnd 0.009312f
C2886 vdd.n984 gnd 0.006516f
C2887 vdd.n985 gnd 0.006516f
C2888 vdd.t246 gnd 0.332944f
C2889 vdd.n986 gnd 0.006516f
C2890 vdd.t50 gnd 0.332944f
C2891 vdd.n987 gnd 0.006516f
C2892 vdd.n988 gnd 0.006516f
C2893 vdd.n989 gnd 0.006516f
C2894 vdd.n990 gnd 0.006516f
C2895 vdd.n991 gnd 0.006516f
C2896 vdd.n992 gnd 0.665888f
C2897 vdd.n993 gnd 0.006516f
C2898 vdd.n994 gnd 0.006516f
C2899 vdd.t22 gnd 0.332944f
C2900 vdd.n995 gnd 0.006516f
C2901 vdd.n996 gnd 0.006516f
C2902 vdd.n997 gnd 0.006516f
C2903 vdd.n998 gnd 0.006516f
C2904 vdd.n999 gnd 0.479831f
C2905 vdd.n1000 gnd 0.006516f
C2906 vdd.n1001 gnd 0.006516f
C2907 vdd.n1002 gnd 0.006516f
C2908 vdd.n1003 gnd 0.006516f
C2909 vdd.n1004 gnd 0.006516f
C2910 vdd.t1 gnd 0.332944f
C2911 vdd.n1005 gnd 0.006516f
C2912 vdd.n1006 gnd 0.006516f
C2913 vdd.t39 gnd 0.332944f
C2914 vdd.n1007 gnd 0.006516f
C2915 vdd.n1008 gnd 0.006516f
C2916 vdd.n1009 gnd 0.006516f
C2917 vdd.t25 gnd 0.332944f
C2918 vdd.n1010 gnd 0.006516f
C2919 vdd.n1011 gnd 0.006516f
C2920 vdd.t2 gnd 0.332944f
C2921 vdd.n1012 gnd 0.006516f
C2922 vdd.n1013 gnd 0.006516f
C2923 vdd.n1014 gnd 0.006516f
C2924 vdd.t26 gnd 0.318255f
C2925 vdd.n1015 gnd 0.006516f
C2926 vdd.n1016 gnd 0.006516f
C2927 vdd.n1017 gnd 0.494519f
C2928 vdd.n1018 gnd 0.006516f
C2929 vdd.n1019 gnd 0.006516f
C2930 vdd.n1020 gnd 0.006516f
C2931 vdd.t43 gnd 0.332944f
C2932 vdd.n1021 gnd 0.006516f
C2933 vdd.n1022 gnd 0.006516f
C2934 vdd.t13 gnd 0.225227f
C2935 vdd.n1023 gnd 0.347632f
C2936 vdd.n1024 gnd 0.006516f
C2937 vdd.n1025 gnd 0.006516f
C2938 vdd.n1026 gnd 0.006516f
C2939 vdd.n1027 gnd 0.612029f
C2940 vdd.n1028 gnd 0.006516f
C2941 vdd.n1029 gnd 0.006516f
C2942 vdd.t52 gnd 0.332944f
C2943 vdd.n1030 gnd 0.006516f
C2944 vdd.n1031 gnd 0.006516f
C2945 vdd.n1032 gnd 0.006516f
C2946 vdd.n1033 gnd 0.665888f
C2947 vdd.n1034 gnd 0.006516f
C2948 vdd.n1035 gnd 0.006516f
C2949 vdd.t19 gnd 0.332944f
C2950 vdd.n1036 gnd 0.006516f
C2951 vdd.n1037 gnd 0.006516f
C2952 vdd.n1038 gnd 0.006516f
C2953 vdd.t12 gnd 0.137094f
C2954 vdd.n1039 gnd 0.006516f
C2955 vdd.n1040 gnd 0.006516f
C2956 vdd.n1041 gnd 0.006516f
C2957 vdd.t261 gnd 0.269524f
C2958 vdd.t259 gnd 0.171895f
C2959 vdd.t262 gnd 0.269524f
C2960 vdd.n1042 gnd 0.151484f
C2961 vdd.n1043 gnd 0.006516f
C2962 vdd.n1044 gnd 0.006516f
C2963 vdd.t34 gnd 0.332944f
C2964 vdd.n1045 gnd 0.006516f
C2965 vdd.n1046 gnd 0.006516f
C2966 vdd.t260 gnd 0.239915f
C2967 vdd.n1047 gnd 0.528793f
C2968 vdd.n1048 gnd 0.006516f
C2969 vdd.n1049 gnd 0.006516f
C2970 vdd.n1050 gnd 0.006516f
C2971 vdd.n1051 gnd 0.386802f
C2972 vdd.n1052 gnd 0.006516f
C2973 vdd.n1053 gnd 0.006516f
C2974 vdd.n1054 gnd 0.425972f
C2975 vdd.n1055 gnd 0.006516f
C2976 vdd.n1056 gnd 0.006516f
C2977 vdd.n1057 gnd 0.006516f
C2978 vdd.n1058 gnd 0.533689f
C2979 vdd.n1059 gnd 0.006516f
C2980 vdd.n1060 gnd 0.006516f
C2981 vdd.t14 gnd 0.332944f
C2982 vdd.n1061 gnd 0.006516f
C2983 vdd.n1062 gnd 0.006516f
C2984 vdd.n1063 gnd 0.006516f
C2985 vdd.n1064 gnd 0.665888f
C2986 vdd.n1065 gnd 0.006516f
C2987 vdd.n1066 gnd 0.006516f
C2988 vdd.t15 gnd 0.332944f
C2989 vdd.n1067 gnd 0.006516f
C2990 vdd.n1068 gnd 0.006516f
C2991 vdd.n1069 gnd 0.006516f
C2992 vdd.t53 gnd 0.332944f
C2993 vdd.n1070 gnd 0.006516f
C2994 vdd.n1071 gnd 0.006516f
C2995 vdd.n1072 gnd 0.006516f
C2996 vdd.n1073 gnd 0.006516f
C2997 vdd.n1074 gnd 0.006516f
C2998 vdd.t45 gnd 0.332944f
C2999 vdd.n1075 gnd 0.006516f
C3000 vdd.n1076 gnd 0.006516f
C3001 vdd.n1077 gnd 0.651199f
C3002 vdd.n1078 gnd 0.006516f
C3003 vdd.n1079 gnd 0.006516f
C3004 vdd.n1080 gnd 0.006516f
C3005 vdd.t7 gnd 0.332944f
C3006 vdd.n1081 gnd 0.006516f
C3007 vdd.n1082 gnd 0.006516f
C3008 vdd.n1083 gnd 0.504312f
C3009 vdd.n1084 gnd 0.006516f
C3010 vdd.n1085 gnd 0.006516f
C3011 vdd.n1086 gnd 0.006516f
C3012 vdd.n1087 gnd 0.665888f
C3013 vdd.n1088 gnd 0.006516f
C3014 vdd.n1089 gnd 0.006516f
C3015 vdd.n1090 gnd 0.357425f
C3016 vdd.n1091 gnd 0.006516f
C3017 vdd.n1092 gnd 0.006516f
C3018 vdd.n1093 gnd 0.006516f
C3019 vdd.n1094 gnd 0.665888f
C3020 vdd.n1095 gnd 0.006516f
C3021 vdd.n1096 gnd 0.006516f
C3022 vdd.n1097 gnd 0.006516f
C3023 vdd.n1098 gnd 0.006516f
C3024 vdd.n1099 gnd 0.006516f
C3025 vdd.t201 gnd 0.332944f
C3026 vdd.n1100 gnd 0.006516f
C3027 vdd.n1101 gnd 0.006516f
C3028 vdd.n1102 gnd 0.006516f
C3029 vdd.n1103 gnd 0.013951f
C3030 vdd.n1104 gnd 0.013951f
C3031 vdd.n1105 gnd 0.900907f
C3032 vdd.n1106 gnd 0.006516f
C3033 vdd.n1107 gnd 0.006516f
C3034 vdd.n1108 gnd 0.474935f
C3035 vdd.n1109 gnd 0.013951f
C3036 vdd.n1110 gnd 0.006516f
C3037 vdd.n1111 gnd 0.006516f
C3038 vdd.n1112 gnd 11.799901f
C3039 vdd.n1146 gnd 0.014795f
C3040 vdd.n1147 gnd 0.006516f
C3041 vdd.n1148 gnd 0.006516f
C3042 vdd.n1149 gnd 0.006133f
C3043 vdd.n1152 gnd 0.02197f
C3044 vdd.n1153 gnd 0.006401f
C3045 vdd.n1154 gnd 0.007712f
C3046 vdd.n1156 gnd 0.009582f
C3047 vdd.n1157 gnd 0.009582f
C3048 vdd.n1158 gnd 0.007712f
C3049 vdd.n1160 gnd 0.009582f
C3050 vdd.n1161 gnd 0.009582f
C3051 vdd.n1162 gnd 0.009582f
C3052 vdd.n1163 gnd 0.009582f
C3053 vdd.n1164 gnd 0.009582f
C3054 vdd.n1165 gnd 0.007712f
C3055 vdd.n1167 gnd 0.009582f
C3056 vdd.n1168 gnd 0.009582f
C3057 vdd.n1169 gnd 0.009582f
C3058 vdd.n1170 gnd 0.009582f
C3059 vdd.n1171 gnd 0.009582f
C3060 vdd.n1172 gnd 0.007712f
C3061 vdd.n1174 gnd 0.009582f
C3062 vdd.n1175 gnd 0.009582f
C3063 vdd.n1176 gnd 0.009582f
C3064 vdd.n1177 gnd 0.009582f
C3065 vdd.n1178 gnd 0.00644f
C3066 vdd.t210 gnd 0.117885f
C3067 vdd.t209 gnd 0.125987f
C3068 vdd.t208 gnd 0.153957f
C3069 vdd.n1179 gnd 0.19735f
C3070 vdd.n1180 gnd 0.16581f
C3071 vdd.n1182 gnd 0.009582f
C3072 vdd.n1183 gnd 0.009582f
C3073 vdd.n1184 gnd 0.007712f
C3074 vdd.n1185 gnd 0.009582f
C3075 vdd.n1187 gnd 0.009582f
C3076 vdd.n1188 gnd 0.009582f
C3077 vdd.n1189 gnd 0.009582f
C3078 vdd.n1190 gnd 0.009582f
C3079 vdd.n1191 gnd 0.007712f
C3080 vdd.n1193 gnd 0.009582f
C3081 vdd.n1194 gnd 0.009582f
C3082 vdd.n1195 gnd 0.009582f
C3083 vdd.n1196 gnd 0.009582f
C3084 vdd.n1197 gnd 0.009582f
C3085 vdd.n1198 gnd 0.007712f
C3086 vdd.n1200 gnd 0.009582f
C3087 vdd.n1201 gnd 0.009582f
C3088 vdd.n1202 gnd 0.009582f
C3089 vdd.n1203 gnd 0.009582f
C3090 vdd.n1204 gnd 0.009582f
C3091 vdd.n1205 gnd 0.007712f
C3092 vdd.n1207 gnd 0.009582f
C3093 vdd.n1208 gnd 0.009582f
C3094 vdd.n1209 gnd 0.009582f
C3095 vdd.n1210 gnd 0.009582f
C3096 vdd.n1211 gnd 0.009582f
C3097 vdd.n1212 gnd 0.007712f
C3098 vdd.n1214 gnd 0.009582f
C3099 vdd.n1215 gnd 0.009582f
C3100 vdd.n1216 gnd 0.009582f
C3101 vdd.n1217 gnd 0.009582f
C3102 vdd.n1218 gnd 0.007635f
C3103 vdd.t207 gnd 0.117885f
C3104 vdd.t206 gnd 0.125987f
C3105 vdd.t204 gnd 0.153957f
C3106 vdd.n1219 gnd 0.19735f
C3107 vdd.n1220 gnd 0.16581f
C3108 vdd.n1222 gnd 0.009582f
C3109 vdd.n1223 gnd 0.009582f
C3110 vdd.n1224 gnd 0.007712f
C3111 vdd.n1225 gnd 0.009582f
C3112 vdd.n1227 gnd 0.009582f
C3113 vdd.n1228 gnd 0.009582f
C3114 vdd.n1229 gnd 0.009582f
C3115 vdd.n1230 gnd 0.009582f
C3116 vdd.n1231 gnd 0.007712f
C3117 vdd.n1233 gnd 0.009582f
C3118 vdd.n1234 gnd 0.009582f
C3119 vdd.n1235 gnd 0.009582f
C3120 vdd.n1236 gnd 0.009582f
C3121 vdd.n1237 gnd 0.009582f
C3122 vdd.n1238 gnd 0.007712f
C3123 vdd.n1240 gnd 0.009582f
C3124 vdd.n1241 gnd 0.009582f
C3125 vdd.n1242 gnd 0.009582f
C3126 vdd.n1243 gnd 0.009582f
C3127 vdd.n1244 gnd 0.009582f
C3128 vdd.n1245 gnd 0.007712f
C3129 vdd.n1247 gnd 0.009582f
C3130 vdd.n1248 gnd 0.009582f
C3131 vdd.n1249 gnd 0.006133f
C3132 vdd.n1250 gnd 0.007712f
C3133 vdd.n1251 gnd 0.014795f
C3134 vdd.n1252 gnd 0.014795f
C3135 vdd.n1253 gnd 0.006516f
C3136 vdd.n1254 gnd 0.006516f
C3137 vdd.n1255 gnd 0.006516f
C3138 vdd.n1256 gnd 0.006516f
C3139 vdd.n1257 gnd 0.006516f
C3140 vdd.n1258 gnd 0.006516f
C3141 vdd.n1259 gnd 0.006516f
C3142 vdd.n1260 gnd 0.006516f
C3143 vdd.n1261 gnd 0.006516f
C3144 vdd.n1262 gnd 0.006516f
C3145 vdd.n1263 gnd 0.006516f
C3146 vdd.n1264 gnd 0.006516f
C3147 vdd.n1265 gnd 0.006516f
C3148 vdd.n1266 gnd 0.006516f
C3149 vdd.n1267 gnd 0.006516f
C3150 vdd.n1268 gnd 0.006516f
C3151 vdd.n1269 gnd 0.006516f
C3152 vdd.n1270 gnd 0.006516f
C3153 vdd.n1271 gnd 0.006516f
C3154 vdd.n1272 gnd 0.006516f
C3155 vdd.n1273 gnd 0.006516f
C3156 vdd.n1274 gnd 0.006516f
C3157 vdd.n1275 gnd 0.006516f
C3158 vdd.n1276 gnd 0.006516f
C3159 vdd.n1277 gnd 0.006516f
C3160 vdd.n1278 gnd 0.006516f
C3161 vdd.n1279 gnd 0.006516f
C3162 vdd.n1280 gnd 0.006516f
C3163 vdd.n1281 gnd 0.006516f
C3164 vdd.n1282 gnd 0.006516f
C3165 vdd.n1283 gnd 0.006516f
C3166 vdd.n1284 gnd 0.006516f
C3167 vdd.n1285 gnd 0.006516f
C3168 vdd.t202 gnd 0.263304f
C3169 vdd.t203 gnd 0.269524f
C3170 vdd.t200 gnd 0.171895f
C3171 vdd.n1286 gnd 0.0929f
C3172 vdd.n1287 gnd 0.052696f
C3173 vdd.n1288 gnd 0.009312f
C3174 vdd.n1289 gnd 0.006516f
C3175 vdd.t236 gnd 0.263304f
C3176 vdd.t237 gnd 0.269524f
C3177 vdd.t235 gnd 0.171895f
C3178 vdd.n1290 gnd 0.0929f
C3179 vdd.n1291 gnd 0.052696f
C3180 vdd.n1292 gnd 0.006516f
C3181 vdd.n1293 gnd 0.006516f
C3182 vdd.n1294 gnd 0.006516f
C3183 vdd.n1295 gnd 0.006516f
C3184 vdd.n1296 gnd 0.006516f
C3185 vdd.n1297 gnd 0.006516f
C3186 vdd.n1298 gnd 0.006516f
C3187 vdd.n1299 gnd 0.006516f
C3188 vdd.n1300 gnd 0.006516f
C3189 vdd.n1301 gnd 0.006516f
C3190 vdd.n1302 gnd 0.006516f
C3191 vdd.n1303 gnd 0.006516f
C3192 vdd.n1304 gnd 0.006516f
C3193 vdd.n1305 gnd 0.006516f
C3194 vdd.n1306 gnd 0.006516f
C3195 vdd.n1307 gnd 0.006516f
C3196 vdd.n1308 gnd 0.006516f
C3197 vdd.n1309 gnd 0.006516f
C3198 vdd.n1310 gnd 0.006516f
C3199 vdd.n1311 gnd 0.006516f
C3200 vdd.n1312 gnd 0.006516f
C3201 vdd.n1313 gnd 0.006516f
C3202 vdd.n1314 gnd 0.006516f
C3203 vdd.n1315 gnd 0.006516f
C3204 vdd.n1316 gnd 0.006516f
C3205 vdd.n1317 gnd 0.006516f
C3206 vdd.n1318 gnd 0.004743f
C3207 vdd.n1319 gnd 0.009312f
C3208 vdd.n1320 gnd 0.005031f
C3209 vdd.n1321 gnd 0.006516f
C3210 vdd.n1322 gnd 0.006516f
C3211 vdd.n1323 gnd 0.006516f
C3212 vdd.n1324 gnd 0.014795f
C3213 vdd.n1325 gnd 0.014795f
C3214 vdd.n1326 gnd 0.013951f
C3215 vdd.n1327 gnd 0.013951f
C3216 vdd.n1328 gnd 0.006516f
C3217 vdd.n1329 gnd 0.006516f
C3218 vdd.n1330 gnd 0.006516f
C3219 vdd.n1331 gnd 0.006516f
C3220 vdd.n1332 gnd 0.006516f
C3221 vdd.n1333 gnd 0.006516f
C3222 vdd.n1334 gnd 0.006516f
C3223 vdd.n1335 gnd 0.006516f
C3224 vdd.n1336 gnd 0.006516f
C3225 vdd.n1337 gnd 0.006516f
C3226 vdd.n1338 gnd 0.006516f
C3227 vdd.n1339 gnd 0.006516f
C3228 vdd.n1340 gnd 0.006516f
C3229 vdd.n1341 gnd 0.006516f
C3230 vdd.n1342 gnd 0.006516f
C3231 vdd.n1343 gnd 0.006516f
C3232 vdd.n1344 gnd 0.006516f
C3233 vdd.n1345 gnd 0.006516f
C3234 vdd.n1346 gnd 0.006516f
C3235 vdd.n1347 gnd 0.006516f
C3236 vdd.n1348 gnd 0.006516f
C3237 vdd.n1349 gnd 0.006516f
C3238 vdd.n1350 gnd 0.006516f
C3239 vdd.n1351 gnd 0.006516f
C3240 vdd.n1352 gnd 0.006516f
C3241 vdd.n1353 gnd 0.006516f
C3242 vdd.n1354 gnd 0.006516f
C3243 vdd.n1355 gnd 0.006516f
C3244 vdd.n1356 gnd 0.006516f
C3245 vdd.n1357 gnd 0.006516f
C3246 vdd.n1358 gnd 0.006516f
C3247 vdd.n1359 gnd 0.006516f
C3248 vdd.n1360 gnd 0.006516f
C3249 vdd.n1361 gnd 0.006516f
C3250 vdd.n1362 gnd 0.006516f
C3251 vdd.n1363 gnd 0.006516f
C3252 vdd.n1364 gnd 0.006516f
C3253 vdd.n1365 gnd 0.006516f
C3254 vdd.n1366 gnd 0.006516f
C3255 vdd.n1367 gnd 0.006516f
C3256 vdd.n1368 gnd 0.006516f
C3257 vdd.n1369 gnd 0.006516f
C3258 vdd.n1370 gnd 0.396595f
C3259 vdd.n1371 gnd 0.006516f
C3260 vdd.n1372 gnd 0.006516f
C3261 vdd.n1373 gnd 0.006516f
C3262 vdd.n1374 gnd 0.006516f
C3263 vdd.n1375 gnd 0.006516f
C3264 vdd.n1376 gnd 0.006516f
C3265 vdd.n1377 gnd 0.006516f
C3266 vdd.n1378 gnd 0.006516f
C3267 vdd.n1379 gnd 0.006516f
C3268 vdd.n1380 gnd 0.006516f
C3269 vdd.n1381 gnd 0.006516f
C3270 vdd.n1382 gnd 0.006516f
C3271 vdd.n1383 gnd 0.006516f
C3272 vdd.n1384 gnd 0.006516f
C3273 vdd.n1385 gnd 0.006516f
C3274 vdd.n1386 gnd 0.006516f
C3275 vdd.n1387 gnd 0.006516f
C3276 vdd.n1388 gnd 0.006516f
C3277 vdd.n1389 gnd 0.006516f
C3278 vdd.n1390 gnd 0.006516f
C3279 vdd.n1391 gnd 0.006516f
C3280 vdd.n1392 gnd 0.006516f
C3281 vdd.n1393 gnd 0.006516f
C3282 vdd.n1394 gnd 0.006516f
C3283 vdd.n1395 gnd 0.006516f
C3284 vdd.n1396 gnd 0.602237f
C3285 vdd.n1397 gnd 0.006516f
C3286 vdd.n1398 gnd 0.006516f
C3287 vdd.n1399 gnd 0.006516f
C3288 vdd.n1400 gnd 0.006516f
C3289 vdd.n1401 gnd 0.006516f
C3290 vdd.n1402 gnd 0.006516f
C3291 vdd.n1403 gnd 0.006516f
C3292 vdd.n1404 gnd 0.006516f
C3293 vdd.n1405 gnd 0.006516f
C3294 vdd.n1406 gnd 0.006516f
C3295 vdd.n1407 gnd 0.006516f
C3296 vdd.n1408 gnd 0.210538f
C3297 vdd.n1409 gnd 0.006516f
C3298 vdd.n1410 gnd 0.006516f
C3299 vdd.n1411 gnd 0.006516f
C3300 vdd.n1412 gnd 0.006516f
C3301 vdd.n1413 gnd 0.006516f
C3302 vdd.n1414 gnd 0.006516f
C3303 vdd.n1415 gnd 0.006516f
C3304 vdd.n1416 gnd 0.006516f
C3305 vdd.n1417 gnd 0.006516f
C3306 vdd.n1418 gnd 0.006516f
C3307 vdd.n1419 gnd 0.006516f
C3308 vdd.n1420 gnd 0.006516f
C3309 vdd.n1421 gnd 0.006516f
C3310 vdd.n1422 gnd 0.006516f
C3311 vdd.n1423 gnd 0.006516f
C3312 vdd.n1424 gnd 0.006516f
C3313 vdd.n1425 gnd 0.006516f
C3314 vdd.n1426 gnd 0.006516f
C3315 vdd.n1427 gnd 0.006516f
C3316 vdd.n1428 gnd 0.006516f
C3317 vdd.n1429 gnd 0.006516f
C3318 vdd.n1430 gnd 0.006516f
C3319 vdd.n1431 gnd 0.006516f
C3320 vdd.n1432 gnd 0.006516f
C3321 vdd.n1433 gnd 0.006516f
C3322 vdd.n1434 gnd 0.006516f
C3323 vdd.n1435 gnd 0.006516f
C3324 vdd.n1436 gnd 0.006516f
C3325 vdd.n1437 gnd 0.006516f
C3326 vdd.n1438 gnd 0.006516f
C3327 vdd.n1439 gnd 0.006516f
C3328 vdd.n1440 gnd 0.006516f
C3329 vdd.n1441 gnd 0.006516f
C3330 vdd.n1442 gnd 0.006516f
C3331 vdd.n1443 gnd 0.006516f
C3332 vdd.n1444 gnd 0.006516f
C3333 vdd.n1445 gnd 0.006516f
C3334 vdd.n1446 gnd 0.006516f
C3335 vdd.n1447 gnd 0.006516f
C3336 vdd.n1448 gnd 0.006516f
C3337 vdd.n1449 gnd 0.006516f
C3338 vdd.n1450 gnd 0.006516f
C3339 vdd.n1451 gnd 0.013951f
C3340 vdd.n1452 gnd 0.013951f
C3341 vdd.n1453 gnd 0.014795f
C3342 vdd.n1454 gnd 0.006516f
C3343 vdd.n1455 gnd 0.006516f
C3344 vdd.n1456 gnd 0.005031f
C3345 vdd.n1457 gnd 0.006516f
C3346 vdd.n1458 gnd 0.006516f
C3347 vdd.n1459 gnd 0.004743f
C3348 vdd.n1460 gnd 0.006516f
C3349 vdd.n1461 gnd 0.006516f
C3350 vdd.n1462 gnd 0.006516f
C3351 vdd.n1463 gnd 0.006516f
C3352 vdd.n1464 gnd 0.006516f
C3353 vdd.n1465 gnd 0.006516f
C3354 vdd.n1466 gnd 0.006516f
C3355 vdd.n1467 gnd 0.006516f
C3356 vdd.n1468 gnd 0.006516f
C3357 vdd.n1469 gnd 0.006516f
C3358 vdd.n1470 gnd 0.006516f
C3359 vdd.n1471 gnd 0.006516f
C3360 vdd.n1472 gnd 0.006516f
C3361 vdd.n1473 gnd 0.006516f
C3362 vdd.n1474 gnd 0.006516f
C3363 vdd.n1475 gnd 0.006516f
C3364 vdd.n1476 gnd 0.006516f
C3365 vdd.n1477 gnd 0.006516f
C3366 vdd.n1478 gnd 0.006516f
C3367 vdd.n1479 gnd 0.006516f
C3368 vdd.n1480 gnd 0.006516f
C3369 vdd.n1481 gnd 0.006516f
C3370 vdd.n1482 gnd 0.006516f
C3371 vdd.n1483 gnd 0.006516f
C3372 vdd.n1484 gnd 0.006516f
C3373 vdd.n1485 gnd 0.006516f
C3374 vdd.n1486 gnd 0.043894f
C3375 vdd.n1488 gnd 0.02197f
C3376 vdd.n1489 gnd 0.007712f
C3377 vdd.n1491 gnd 0.009582f
C3378 vdd.n1492 gnd 0.007712f
C3379 vdd.n1493 gnd 0.009582f
C3380 vdd.n1495 gnd 0.009582f
C3381 vdd.n1496 gnd 0.009582f
C3382 vdd.n1498 gnd 0.009582f
C3383 vdd.n1499 gnd 0.006401f
C3384 vdd.n1500 gnd 0.543482f
C3385 vdd.n1501 gnd 0.009582f
C3386 vdd.n1502 gnd 0.02197f
C3387 vdd.n1503 gnd 0.007712f
C3388 vdd.n1504 gnd 0.009582f
C3389 vdd.n1505 gnd 0.007712f
C3390 vdd.n1506 gnd 0.009582f
C3391 vdd.n1507 gnd 0.979246f
C3392 vdd.n1508 gnd 0.009582f
C3393 vdd.n1509 gnd 0.007712f
C3394 vdd.n1510 gnd 0.007712f
C3395 vdd.n1511 gnd 0.009582f
C3396 vdd.n1512 gnd 0.007712f
C3397 vdd.n1513 gnd 0.009582f
C3398 vdd.t89 gnd 0.489623f
C3399 vdd.n1514 gnd 0.009582f
C3400 vdd.n1515 gnd 0.007712f
C3401 vdd.n1516 gnd 0.009582f
C3402 vdd.n1517 gnd 0.007712f
C3403 vdd.n1518 gnd 0.009582f
C3404 vdd.t130 gnd 0.489623f
C3405 vdd.n1519 gnd 0.009582f
C3406 vdd.n1520 gnd 0.007712f
C3407 vdd.n1521 gnd 0.009582f
C3408 vdd.n1522 gnd 0.007712f
C3409 vdd.n1523 gnd 0.009582f
C3410 vdd.t132 gnd 0.489623f
C3411 vdd.n1524 gnd 0.680576f
C3412 vdd.n1525 gnd 0.009582f
C3413 vdd.n1526 gnd 0.007712f
C3414 vdd.n1527 gnd 0.009582f
C3415 vdd.n1528 gnd 0.007712f
C3416 vdd.n1529 gnd 0.009582f
C3417 vdd.n1530 gnd 0.778501f
C3418 vdd.n1531 gnd 0.009582f
C3419 vdd.n1532 gnd 0.007712f
C3420 vdd.n1533 gnd 0.009582f
C3421 vdd.n1534 gnd 0.007712f
C3422 vdd.n1535 gnd 0.009582f
C3423 vdd.n1536 gnd 0.612029f
C3424 vdd.t86 gnd 0.489623f
C3425 vdd.n1537 gnd 0.009582f
C3426 vdd.n1538 gnd 0.007712f
C3427 vdd.n1539 gnd 0.009582f
C3428 vdd.n1540 gnd 0.007712f
C3429 vdd.n1541 gnd 0.009582f
C3430 vdd.t58 gnd 0.489623f
C3431 vdd.n1542 gnd 0.009582f
C3432 vdd.n1543 gnd 0.007712f
C3433 vdd.n1544 gnd 0.009582f
C3434 vdd.n1545 gnd 0.007712f
C3435 vdd.n1546 gnd 0.009582f
C3436 vdd.t62 gnd 0.489623f
C3437 vdd.n1547 gnd 0.533689f
C3438 vdd.n1548 gnd 0.009582f
C3439 vdd.n1549 gnd 0.007712f
C3440 vdd.n1550 gnd 0.009582f
C3441 vdd.n1551 gnd 0.007712f
C3442 vdd.n1552 gnd 0.009582f
C3443 vdd.t105 gnd 0.489623f
C3444 vdd.n1553 gnd 0.009582f
C3445 vdd.n1554 gnd 0.007712f
C3446 vdd.n1555 gnd 0.009582f
C3447 vdd.n1556 gnd 0.007712f
C3448 vdd.n1557 gnd 0.009582f
C3449 vdd.n1558 gnd 0.758916f
C3450 vdd.n1559 gnd 0.812775f
C3451 vdd.t128 gnd 0.489623f
C3452 vdd.n1560 gnd 0.009582f
C3453 vdd.n1561 gnd 0.007712f
C3454 vdd.n1562 gnd 0.009582f
C3455 vdd.n1563 gnd 0.007712f
C3456 vdd.n1564 gnd 0.009582f
C3457 vdd.n1565 gnd 0.592444f
C3458 vdd.n1566 gnd 0.009582f
C3459 vdd.n1567 gnd 0.007712f
C3460 vdd.n1568 gnd 0.009582f
C3461 vdd.n1569 gnd 0.007712f
C3462 vdd.n1570 gnd 0.009582f
C3463 vdd.t144 gnd 0.489623f
C3464 vdd.t97 gnd 0.489623f
C3465 vdd.n1571 gnd 0.009582f
C3466 vdd.n1572 gnd 0.007712f
C3467 vdd.n1573 gnd 0.009582f
C3468 vdd.n1574 gnd 0.007712f
C3469 vdd.n1575 gnd 0.009582f
C3470 vdd.t116 gnd 0.489623f
C3471 vdd.n1576 gnd 0.009582f
C3472 vdd.n1577 gnd 0.007712f
C3473 vdd.n1578 gnd 0.009582f
C3474 vdd.n1579 gnd 0.007712f
C3475 vdd.n1580 gnd 0.009582f
C3476 vdd.t91 gnd 0.489623f
C3477 vdd.n1581 gnd 0.719746f
C3478 vdd.n1582 gnd 0.009582f
C3479 vdd.n1583 gnd 0.007712f
C3480 vdd.n1584 gnd 0.009582f
C3481 vdd.n1585 gnd 0.007712f
C3482 vdd.n1586 gnd 0.009582f
C3483 vdd.n1587 gnd 0.979246f
C3484 vdd.n1588 gnd 0.009582f
C3485 vdd.n1589 gnd 0.007712f
C3486 vdd.n1590 gnd 0.009582f
C3487 vdd.n1591 gnd 0.007712f
C3488 vdd.n1592 gnd 0.009582f
C3489 vdd.n1593 gnd 0.827463f
C3490 vdd.n1594 gnd 0.009582f
C3491 vdd.n1595 gnd 0.007712f
C3492 vdd.n1596 gnd 0.021821f
C3493 vdd.n1597 gnd 0.006401f
C3494 vdd.n1598 gnd 0.021821f
C3495 vdd.n1599 gnd 1.29261f
C3496 vdd.n1600 gnd 0.021821f
C3497 vdd.n1601 gnd 0.006401f
C3498 vdd.n1602 gnd 0.009582f
C3499 vdd.t243 gnd 0.117885f
C3500 vdd.t244 gnd 0.125987f
C3501 vdd.t241 gnd 0.153957f
C3502 vdd.n1603 gnd 0.19735f
C3503 vdd.n1604 gnd 0.166581f
C3504 vdd.n1605 gnd 0.012648f
C3505 vdd.n1606 gnd 0.009582f
C3506 vdd.n1637 gnd 0.009582f
C3507 vdd.n1638 gnd 0.009582f
C3508 vdd.n1639 gnd 0.02197f
C3509 vdd.n1640 gnd 0.007712f
C3510 vdd.n1641 gnd 0.009582f
C3511 vdd.n1642 gnd 0.009582f
C3512 vdd.n1643 gnd 0.009582f
C3513 vdd.n1644 gnd 0.009582f
C3514 vdd.n1645 gnd 0.007712f
C3515 vdd.n1646 gnd 0.009582f
C3516 vdd.n1647 gnd 0.009582f
C3517 vdd.n1648 gnd 0.009582f
C3518 vdd.n1649 gnd 0.009582f
C3519 vdd.n1650 gnd 0.009582f
C3520 vdd.n1651 gnd 0.007712f
C3521 vdd.n1652 gnd 0.009582f
C3522 vdd.n1653 gnd 0.009582f
C3523 vdd.n1654 gnd 0.009582f
C3524 vdd.n1655 gnd 0.009582f
C3525 vdd.n1656 gnd 0.009582f
C3526 vdd.n1657 gnd 0.007712f
C3527 vdd.n1658 gnd 0.009582f
C3528 vdd.n1659 gnd 0.009582f
C3529 vdd.n1660 gnd 0.009582f
C3530 vdd.n1661 gnd 0.009582f
C3531 vdd.n1662 gnd 0.009582f
C3532 vdd.n1663 gnd 0.00644f
C3533 vdd.n1664 gnd 0.009582f
C3534 vdd.n1665 gnd 0.009582f
C3535 vdd.n1666 gnd 0.009582f
C3536 vdd.n1667 gnd 0.007712f
C3537 vdd.n1668 gnd 0.009582f
C3538 vdd.n1669 gnd 0.009582f
C3539 vdd.n1670 gnd 0.009582f
C3540 vdd.n1671 gnd 0.009582f
C3541 vdd.n1672 gnd 0.009582f
C3542 vdd.n1673 gnd 0.007712f
C3543 vdd.n1674 gnd 0.009582f
C3544 vdd.n1675 gnd 0.009582f
C3545 vdd.n1676 gnd 0.009582f
C3546 vdd.n1677 gnd 0.009582f
C3547 vdd.n1678 gnd 0.009582f
C3548 vdd.n1679 gnd 0.007712f
C3549 vdd.n1680 gnd 0.009582f
C3550 vdd.n1681 gnd 0.009582f
C3551 vdd.n1682 gnd 0.009582f
C3552 vdd.n1683 gnd 0.009582f
C3553 vdd.n1684 gnd 0.009582f
C3554 vdd.n1685 gnd 0.007712f
C3555 vdd.n1686 gnd 0.009582f
C3556 vdd.n1687 gnd 0.009582f
C3557 vdd.n1688 gnd 0.009582f
C3558 vdd.n1689 gnd 0.009582f
C3559 vdd.n1690 gnd 0.009582f
C3560 vdd.n1691 gnd 0.007712f
C3561 vdd.n1692 gnd 0.009582f
C3562 vdd.n1693 gnd 0.009582f
C3563 vdd.n1694 gnd 0.009582f
C3564 vdd.n1695 gnd 0.009582f
C3565 vdd.n1696 gnd 0.007635f
C3566 vdd.n1697 gnd 0.009582f
C3567 vdd.n1698 gnd 0.009582f
C3568 vdd.n1699 gnd 0.009582f
C3569 vdd.n1700 gnd 0.009582f
C3570 vdd.n1701 gnd 0.009582f
C3571 vdd.n1702 gnd 0.007712f
C3572 vdd.n1703 gnd 0.009582f
C3573 vdd.n1704 gnd 0.009582f
C3574 vdd.n1705 gnd 0.009582f
C3575 vdd.n1706 gnd 0.009582f
C3576 vdd.n1707 gnd 0.009582f
C3577 vdd.n1708 gnd 0.007712f
C3578 vdd.n1709 gnd 0.009582f
C3579 vdd.n1710 gnd 0.009582f
C3580 vdd.n1711 gnd 0.009582f
C3581 vdd.n1712 gnd 0.009582f
C3582 vdd.n1713 gnd 0.009582f
C3583 vdd.n1714 gnd 0.007712f
C3584 vdd.n1715 gnd 0.009582f
C3585 vdd.n1716 gnd 0.009582f
C3586 vdd.n1717 gnd 0.009582f
C3587 vdd.n1718 gnd 0.009582f
C3588 vdd.n1719 gnd 0.009582f
C3589 vdd.n1720 gnd 0.007712f
C3590 vdd.n1721 gnd 0.009582f
C3591 vdd.n1722 gnd 0.009582f
C3592 vdd.n1723 gnd 0.009582f
C3593 vdd.n1724 gnd 0.009582f
C3594 vdd.n1725 gnd 0.009582f
C3595 vdd.n1726 gnd 0.004049f
C3596 vdd.n1727 gnd 0.009582f
C3597 vdd.n1728 gnd 0.007712f
C3598 vdd.n1729 gnd 0.007712f
C3599 vdd.n1730 gnd 0.007712f
C3600 vdd.n1731 gnd 0.009582f
C3601 vdd.n1732 gnd 0.009582f
C3602 vdd.n1733 gnd 0.009582f
C3603 vdd.n1734 gnd 0.007712f
C3604 vdd.n1735 gnd 0.007712f
C3605 vdd.n1736 gnd 0.007712f
C3606 vdd.n1737 gnd 0.009582f
C3607 vdd.n1738 gnd 0.009582f
C3608 vdd.n1739 gnd 0.009582f
C3609 vdd.n1740 gnd 0.007712f
C3610 vdd.n1741 gnd 0.007712f
C3611 vdd.n1742 gnd 0.007712f
C3612 vdd.n1743 gnd 0.009582f
C3613 vdd.n1744 gnd 0.009582f
C3614 vdd.n1745 gnd 0.009582f
C3615 vdd.n1746 gnd 0.007712f
C3616 vdd.n1747 gnd 0.007712f
C3617 vdd.n1748 gnd 0.007712f
C3618 vdd.n1749 gnd 0.009582f
C3619 vdd.n1750 gnd 0.009582f
C3620 vdd.n1751 gnd 0.009582f
C3621 vdd.n1752 gnd 0.007712f
C3622 vdd.n1753 gnd 0.007712f
C3623 vdd.n1754 gnd 0.007712f
C3624 vdd.n1755 gnd 0.009582f
C3625 vdd.n1756 gnd 0.009582f
C3626 vdd.n1757 gnd 0.009582f
C3627 vdd.n1758 gnd 0.009582f
C3628 vdd.t257 gnd 0.117885f
C3629 vdd.t258 gnd 0.125987f
C3630 vdd.t256 gnd 0.153957f
C3631 vdd.n1759 gnd 0.19735f
C3632 vdd.n1760 gnd 0.166581f
C3633 vdd.n1761 gnd 0.016505f
C3634 vdd.n1762 gnd 0.005244f
C3635 vdd.n1763 gnd 0.007712f
C3636 vdd.n1764 gnd 0.009582f
C3637 vdd.n1765 gnd 0.009582f
C3638 vdd.n1766 gnd 0.009582f
C3639 vdd.n1767 gnd 0.007712f
C3640 vdd.n1768 gnd 0.007712f
C3641 vdd.n1769 gnd 0.007712f
C3642 vdd.n1770 gnd 0.009582f
C3643 vdd.n1771 gnd 0.009582f
C3644 vdd.n1772 gnd 0.009582f
C3645 vdd.n1773 gnd 0.007712f
C3646 vdd.n1774 gnd 0.007712f
C3647 vdd.n1775 gnd 0.007712f
C3648 vdd.n1776 gnd 0.009582f
C3649 vdd.n1777 gnd 0.009582f
C3650 vdd.n1778 gnd 0.009582f
C3651 vdd.n1779 gnd 0.007712f
C3652 vdd.n1780 gnd 0.007712f
C3653 vdd.n1781 gnd 0.007712f
C3654 vdd.n1782 gnd 0.009582f
C3655 vdd.n1783 gnd 0.009582f
C3656 vdd.n1784 gnd 0.009582f
C3657 vdd.n1785 gnd 0.007712f
C3658 vdd.n1786 gnd 0.007712f
C3659 vdd.n1787 gnd 0.007712f
C3660 vdd.n1788 gnd 0.009582f
C3661 vdd.n1789 gnd 0.009582f
C3662 vdd.n1790 gnd 0.009582f
C3663 vdd.n1791 gnd 0.007712f
C3664 vdd.n1792 gnd 0.00644f
C3665 vdd.n1793 gnd 0.009582f
C3666 vdd.n1794 gnd 0.009582f
C3667 vdd.t267 gnd 0.117885f
C3668 vdd.t268 gnd 0.125987f
C3669 vdd.t266 gnd 0.153957f
C3670 vdd.n1795 gnd 0.19735f
C3671 vdd.n1796 gnd 0.166581f
C3672 vdd.n1797 gnd 0.016505f
C3673 vdd.n1798 gnd 0.009582f
C3674 vdd.n1799 gnd 0.009582f
C3675 vdd.n1800 gnd 0.009582f
C3676 vdd.n1801 gnd 0.007712f
C3677 vdd.n1802 gnd 0.007712f
C3678 vdd.n1803 gnd 0.007712f
C3679 vdd.n1804 gnd 0.009582f
C3680 vdd.n1805 gnd 0.009582f
C3681 vdd.n1806 gnd 0.009582f
C3682 vdd.n1807 gnd 0.007712f
C3683 vdd.n1808 gnd 0.007712f
C3684 vdd.n1809 gnd 0.007712f
C3685 vdd.n1810 gnd 0.009582f
C3686 vdd.n1811 gnd 0.009582f
C3687 vdd.n1812 gnd 0.009582f
C3688 vdd.n1813 gnd 0.007712f
C3689 vdd.n1814 gnd 0.007712f
C3690 vdd.n1815 gnd 0.007712f
C3691 vdd.n1816 gnd 0.009582f
C3692 vdd.n1817 gnd 0.009582f
C3693 vdd.n1818 gnd 0.009582f
C3694 vdd.n1819 gnd 0.007712f
C3695 vdd.n1820 gnd 0.007712f
C3696 vdd.n1821 gnd 0.007712f
C3697 vdd.n1822 gnd 0.009582f
C3698 vdd.n1823 gnd 0.009582f
C3699 vdd.n1824 gnd 0.009582f
C3700 vdd.n1825 gnd 0.007712f
C3701 vdd.n1826 gnd 0.006401f
C3702 vdd.n1827 gnd 0.02197f
C3703 vdd.n1829 gnd 2.16413f
C3704 vdd.n1830 gnd 0.02197f
C3705 vdd.n1831 gnd 0.003663f
C3706 vdd.n1832 gnd 0.02197f
C3707 vdd.n1833 gnd 0.021821f
C3708 vdd.n1834 gnd 0.009582f
C3709 vdd.n1835 gnd 0.007712f
C3710 vdd.n1836 gnd 0.009582f
C3711 vdd.t242 gnd 0.489623f
C3712 vdd.n1837 gnd 0.641406f
C3713 vdd.n1838 gnd 0.009582f
C3714 vdd.n1839 gnd 0.007712f
C3715 vdd.n1840 gnd 0.009582f
C3716 vdd.n1841 gnd 0.009582f
C3717 vdd.n1842 gnd 0.009582f
C3718 vdd.n1843 gnd 0.007712f
C3719 vdd.n1844 gnd 0.009582f
C3720 vdd.n1845 gnd 0.979246f
C3721 vdd.n1846 gnd 0.009582f
C3722 vdd.n1847 gnd 0.007712f
C3723 vdd.n1848 gnd 0.009582f
C3724 vdd.n1849 gnd 0.009582f
C3725 vdd.n1850 gnd 0.009582f
C3726 vdd.n1851 gnd 0.007712f
C3727 vdd.n1852 gnd 0.009582f
C3728 vdd.n1853 gnd 0.812775f
C3729 vdd.t123 gnd 0.489623f
C3730 vdd.n1854 gnd 0.563067f
C3731 vdd.n1855 gnd 0.009582f
C3732 vdd.n1856 gnd 0.007712f
C3733 vdd.n1857 gnd 0.009582f
C3734 vdd.n1858 gnd 0.009582f
C3735 vdd.n1859 gnd 0.009582f
C3736 vdd.n1860 gnd 0.007712f
C3737 vdd.n1861 gnd 0.009582f
C3738 vdd.n1862 gnd 0.582652f
C3739 vdd.n1863 gnd 0.009582f
C3740 vdd.n1864 gnd 0.007712f
C3741 vdd.n1865 gnd 0.009582f
C3742 vdd.n1866 gnd 0.009582f
C3743 vdd.n1867 gnd 0.009582f
C3744 vdd.n1868 gnd 0.007712f
C3745 vdd.n1869 gnd 0.009582f
C3746 vdd.n1870 gnd 0.553274f
C3747 vdd.n1871 gnd 0.749124f
C3748 vdd.n1872 gnd 0.009582f
C3749 vdd.n1873 gnd 0.007712f
C3750 vdd.n1874 gnd 0.009582f
C3751 vdd.n1875 gnd 0.009582f
C3752 vdd.n1876 gnd 0.009582f
C3753 vdd.n1877 gnd 0.007712f
C3754 vdd.n1878 gnd 0.009582f
C3755 vdd.n1879 gnd 0.812775f
C3756 vdd.n1880 gnd 0.009582f
C3757 vdd.n1881 gnd 0.007712f
C3758 vdd.n1882 gnd 0.009582f
C3759 vdd.n1883 gnd 0.009582f
C3760 vdd.n1884 gnd 0.009582f
C3761 vdd.n1885 gnd 0.007712f
C3762 vdd.n1886 gnd 0.009582f
C3763 vdd.t56 gnd 0.489623f
C3764 vdd.n1887 gnd 0.709954f
C3765 vdd.n1888 gnd 0.009582f
C3766 vdd.n1889 gnd 0.007712f
C3767 vdd.n1890 gnd 0.009582f
C3768 vdd.n1891 gnd 0.009582f
C3769 vdd.n1892 gnd 0.009582f
C3770 vdd.n1893 gnd 0.007712f
C3771 vdd.n1894 gnd 0.009582f
C3772 vdd.n1895 gnd 0.543482f
C3773 vdd.n1896 gnd 0.009582f
C3774 vdd.n1897 gnd 0.007712f
C3775 vdd.n1898 gnd 0.009582f
C3776 vdd.n1899 gnd 0.009582f
C3777 vdd.n1900 gnd 0.009582f
C3778 vdd.n1901 gnd 0.007712f
C3779 vdd.n1902 gnd 0.009582f
C3780 vdd.n1903 gnd 0.700161f
C3781 vdd.n1904 gnd 0.602237f
C3782 vdd.n1905 gnd 0.009582f
C3783 vdd.n1906 gnd 0.007712f
C3784 vdd.n1907 gnd 0.007364f
C3785 vdd.n1908 gnd 0.005259f
C3786 vdd.n1909 gnd 0.00488f
C3787 vdd.n1910 gnd 0.002699f
C3788 vdd.n1911 gnd 0.006198f
C3789 vdd.n1912 gnd 0.002622f
C3790 vdd.n1913 gnd 0.002776f
C3791 vdd.n1914 gnd 0.00488f
C3792 vdd.n1915 gnd 0.002622f
C3793 vdd.n1916 gnd 0.006198f
C3794 vdd.n1917 gnd 0.002776f
C3795 vdd.n1918 gnd 0.00488f
C3796 vdd.n1919 gnd 0.002622f
C3797 vdd.n1920 gnd 0.004648f
C3798 vdd.n1921 gnd 0.004662f
C3799 vdd.t126 gnd 0.013316f
C3800 vdd.n1922 gnd 0.029628f
C3801 vdd.n1923 gnd 0.154189f
C3802 vdd.n1924 gnd 0.002622f
C3803 vdd.n1925 gnd 0.002776f
C3804 vdd.n1926 gnd 0.006198f
C3805 vdd.n1927 gnd 0.006198f
C3806 vdd.n1928 gnd 0.002776f
C3807 vdd.n1929 gnd 0.002622f
C3808 vdd.n1930 gnd 0.00488f
C3809 vdd.n1931 gnd 0.00488f
C3810 vdd.n1932 gnd 0.002622f
C3811 vdd.n1933 gnd 0.002776f
C3812 vdd.n1934 gnd 0.006198f
C3813 vdd.n1935 gnd 0.006198f
C3814 vdd.n1936 gnd 0.002776f
C3815 vdd.n1937 gnd 0.002622f
C3816 vdd.n1938 gnd 0.00488f
C3817 vdd.n1939 gnd 0.00488f
C3818 vdd.n1940 gnd 0.002622f
C3819 vdd.n1941 gnd 0.002776f
C3820 vdd.n1942 gnd 0.006198f
C3821 vdd.n1943 gnd 0.006198f
C3822 vdd.n1944 gnd 0.014653f
C3823 vdd.n1945 gnd 0.002699f
C3824 vdd.n1946 gnd 0.002622f
C3825 vdd.n1947 gnd 0.012613f
C3826 vdd.n1948 gnd 0.008806f
C3827 vdd.t164 gnd 0.03085f
C3828 vdd.t183 gnd 0.03085f
C3829 vdd.n1949 gnd 0.212021f
C3830 vdd.n1950 gnd 0.166722f
C3831 vdd.t148 gnd 0.03085f
C3832 vdd.t79 gnd 0.03085f
C3833 vdd.n1951 gnd 0.212021f
C3834 vdd.n1952 gnd 0.134544f
C3835 vdd.t134 gnd 0.03085f
C3836 vdd.t82 gnd 0.03085f
C3837 vdd.n1953 gnd 0.212021f
C3838 vdd.n1954 gnd 0.134544f
C3839 vdd.t173 gnd 0.03085f
C3840 vdd.t111 gnd 0.03085f
C3841 vdd.n1955 gnd 0.212021f
C3842 vdd.n1956 gnd 0.134544f
C3843 vdd.t154 gnd 0.03085f
C3844 vdd.t129 gnd 0.03085f
C3845 vdd.n1957 gnd 0.212021f
C3846 vdd.n1958 gnd 0.134544f
C3847 vdd.t166 gnd 0.03085f
C3848 vdd.t99 gnd 0.03085f
C3849 vdd.n1959 gnd 0.212021f
C3850 vdd.n1960 gnd 0.134544f
C3851 vdd.t176 gnd 0.03085f
C3852 vdd.t117 gnd 0.03085f
C3853 vdd.n1961 gnd 0.212021f
C3854 vdd.n1962 gnd 0.134544f
C3855 vdd.n1963 gnd 0.005259f
C3856 vdd.n1964 gnd 0.00488f
C3857 vdd.n1965 gnd 0.002699f
C3858 vdd.n1966 gnd 0.006198f
C3859 vdd.n1967 gnd 0.002622f
C3860 vdd.n1968 gnd 0.002776f
C3861 vdd.n1969 gnd 0.00488f
C3862 vdd.n1970 gnd 0.002622f
C3863 vdd.n1971 gnd 0.006198f
C3864 vdd.n1972 gnd 0.002776f
C3865 vdd.n1973 gnd 0.00488f
C3866 vdd.n1974 gnd 0.002622f
C3867 vdd.n1975 gnd 0.004648f
C3868 vdd.n1976 gnd 0.004662f
C3869 vdd.t139 gnd 0.013316f
C3870 vdd.n1977 gnd 0.029628f
C3871 vdd.n1978 gnd 0.154189f
C3872 vdd.n1979 gnd 0.002622f
C3873 vdd.n1980 gnd 0.002776f
C3874 vdd.n1981 gnd 0.006198f
C3875 vdd.n1982 gnd 0.006198f
C3876 vdd.n1983 gnd 0.002776f
C3877 vdd.n1984 gnd 0.002622f
C3878 vdd.n1985 gnd 0.00488f
C3879 vdd.n1986 gnd 0.00488f
C3880 vdd.n1987 gnd 0.002622f
C3881 vdd.n1988 gnd 0.002776f
C3882 vdd.n1989 gnd 0.006198f
C3883 vdd.n1990 gnd 0.006198f
C3884 vdd.n1991 gnd 0.002776f
C3885 vdd.n1992 gnd 0.002622f
C3886 vdd.n1993 gnd 0.00488f
C3887 vdd.n1994 gnd 0.00488f
C3888 vdd.n1995 gnd 0.002622f
C3889 vdd.n1996 gnd 0.002776f
C3890 vdd.n1997 gnd 0.006198f
C3891 vdd.n1998 gnd 0.006198f
C3892 vdd.n1999 gnd 0.014653f
C3893 vdd.n2000 gnd 0.002699f
C3894 vdd.n2001 gnd 0.002622f
C3895 vdd.n2002 gnd 0.012613f
C3896 vdd.n2003 gnd 0.008529f
C3897 vdd.n2004 gnd 0.100101f
C3898 vdd.n2005 gnd 0.005259f
C3899 vdd.n2006 gnd 0.00488f
C3900 vdd.n2007 gnd 0.002699f
C3901 vdd.n2008 gnd 0.006198f
C3902 vdd.n2009 gnd 0.002622f
C3903 vdd.n2010 gnd 0.002776f
C3904 vdd.n2011 gnd 0.00488f
C3905 vdd.n2012 gnd 0.002622f
C3906 vdd.n2013 gnd 0.006198f
C3907 vdd.n2014 gnd 0.002776f
C3908 vdd.n2015 gnd 0.00488f
C3909 vdd.n2016 gnd 0.002622f
C3910 vdd.n2017 gnd 0.004648f
C3911 vdd.n2018 gnd 0.004662f
C3912 vdd.t90 gnd 0.013316f
C3913 vdd.n2019 gnd 0.029628f
C3914 vdd.n2020 gnd 0.154189f
C3915 vdd.n2021 gnd 0.002622f
C3916 vdd.n2022 gnd 0.002776f
C3917 vdd.n2023 gnd 0.006198f
C3918 vdd.n2024 gnd 0.006198f
C3919 vdd.n2025 gnd 0.002776f
C3920 vdd.n2026 gnd 0.002622f
C3921 vdd.n2027 gnd 0.00488f
C3922 vdd.n2028 gnd 0.00488f
C3923 vdd.n2029 gnd 0.002622f
C3924 vdd.n2030 gnd 0.002776f
C3925 vdd.n2031 gnd 0.006198f
C3926 vdd.n2032 gnd 0.006198f
C3927 vdd.n2033 gnd 0.002776f
C3928 vdd.n2034 gnd 0.002622f
C3929 vdd.n2035 gnd 0.00488f
C3930 vdd.n2036 gnd 0.00488f
C3931 vdd.n2037 gnd 0.002622f
C3932 vdd.n2038 gnd 0.002776f
C3933 vdd.n2039 gnd 0.006198f
C3934 vdd.n2040 gnd 0.006198f
C3935 vdd.n2041 gnd 0.014653f
C3936 vdd.n2042 gnd 0.002699f
C3937 vdd.n2043 gnd 0.002622f
C3938 vdd.n2044 gnd 0.012613f
C3939 vdd.n2045 gnd 0.008806f
C3940 vdd.t133 gnd 0.03085f
C3941 vdd.t131 gnd 0.03085f
C3942 vdd.n2046 gnd 0.212021f
C3943 vdd.n2047 gnd 0.166722f
C3944 vdd.t87 gnd 0.03085f
C3945 vdd.t65 gnd 0.03085f
C3946 vdd.n2048 gnd 0.212021f
C3947 vdd.n2049 gnd 0.134544f
C3948 vdd.t59 gnd 0.03085f
C3949 vdd.t127 gnd 0.03085f
C3950 vdd.n2050 gnd 0.212021f
C3951 vdd.n2051 gnd 0.134544f
C3952 vdd.t106 gnd 0.03085f
C3953 vdd.t63 gnd 0.03085f
C3954 vdd.n2052 gnd 0.212021f
C3955 vdd.n2053 gnd 0.134544f
C3956 vdd.t57 gnd 0.03085f
C3957 vdd.t149 gnd 0.03085f
C3958 vdd.n2054 gnd 0.212021f
C3959 vdd.n2055 gnd 0.134544f
C3960 vdd.t145 gnd 0.03085f
C3961 vdd.t101 gnd 0.03085f
C3962 vdd.n2056 gnd 0.212021f
C3963 vdd.n2057 gnd 0.134544f
C3964 vdd.t92 gnd 0.03085f
C3965 vdd.t171 gnd 0.03085f
C3966 vdd.n2058 gnd 0.212021f
C3967 vdd.n2059 gnd 0.134544f
C3968 vdd.n2060 gnd 0.005259f
C3969 vdd.n2061 gnd 0.00488f
C3970 vdd.n2062 gnd 0.002699f
C3971 vdd.n2063 gnd 0.006198f
C3972 vdd.n2064 gnd 0.002622f
C3973 vdd.n2065 gnd 0.002776f
C3974 vdd.n2066 gnd 0.00488f
C3975 vdd.n2067 gnd 0.002622f
C3976 vdd.n2068 gnd 0.006198f
C3977 vdd.n2069 gnd 0.002776f
C3978 vdd.n2070 gnd 0.00488f
C3979 vdd.n2071 gnd 0.002622f
C3980 vdd.n2072 gnd 0.004648f
C3981 vdd.n2073 gnd 0.004662f
C3982 vdd.t124 gnd 0.013316f
C3983 vdd.n2074 gnd 0.029628f
C3984 vdd.n2075 gnd 0.154189f
C3985 vdd.n2076 gnd 0.002622f
C3986 vdd.n2077 gnd 0.002776f
C3987 vdd.n2078 gnd 0.006198f
C3988 vdd.n2079 gnd 0.006198f
C3989 vdd.n2080 gnd 0.002776f
C3990 vdd.n2081 gnd 0.002622f
C3991 vdd.n2082 gnd 0.00488f
C3992 vdd.n2083 gnd 0.00488f
C3993 vdd.n2084 gnd 0.002622f
C3994 vdd.n2085 gnd 0.002776f
C3995 vdd.n2086 gnd 0.006198f
C3996 vdd.n2087 gnd 0.006198f
C3997 vdd.n2088 gnd 0.002776f
C3998 vdd.n2089 gnd 0.002622f
C3999 vdd.n2090 gnd 0.00488f
C4000 vdd.n2091 gnd 0.00488f
C4001 vdd.n2092 gnd 0.002622f
C4002 vdd.n2093 gnd 0.002776f
C4003 vdd.n2094 gnd 0.006198f
C4004 vdd.n2095 gnd 0.006198f
C4005 vdd.n2096 gnd 0.014653f
C4006 vdd.n2097 gnd 0.002699f
C4007 vdd.n2098 gnd 0.002622f
C4008 vdd.n2099 gnd 0.012613f
C4009 vdd.n2100 gnd 0.008529f
C4010 vdd.n2101 gnd 0.05955f
C4011 vdd.n2102 gnd 0.214575f
C4012 vdd.n2103 gnd 0.005259f
C4013 vdd.n2104 gnd 0.00488f
C4014 vdd.n2105 gnd 0.002699f
C4015 vdd.n2106 gnd 0.006198f
C4016 vdd.n2107 gnd 0.002622f
C4017 vdd.n2108 gnd 0.002776f
C4018 vdd.n2109 gnd 0.00488f
C4019 vdd.n2110 gnd 0.002622f
C4020 vdd.n2111 gnd 0.006198f
C4021 vdd.n2112 gnd 0.002776f
C4022 vdd.n2113 gnd 0.00488f
C4023 vdd.n2114 gnd 0.002622f
C4024 vdd.n2115 gnd 0.004648f
C4025 vdd.n2116 gnd 0.004662f
C4026 vdd.t107 gnd 0.013316f
C4027 vdd.n2117 gnd 0.029628f
C4028 vdd.n2118 gnd 0.154189f
C4029 vdd.n2119 gnd 0.002622f
C4030 vdd.n2120 gnd 0.002776f
C4031 vdd.n2121 gnd 0.006198f
C4032 vdd.n2122 gnd 0.006198f
C4033 vdd.n2123 gnd 0.002776f
C4034 vdd.n2124 gnd 0.002622f
C4035 vdd.n2125 gnd 0.00488f
C4036 vdd.n2126 gnd 0.00488f
C4037 vdd.n2127 gnd 0.002622f
C4038 vdd.n2128 gnd 0.002776f
C4039 vdd.n2129 gnd 0.006198f
C4040 vdd.n2130 gnd 0.006198f
C4041 vdd.n2131 gnd 0.002776f
C4042 vdd.n2132 gnd 0.002622f
C4043 vdd.n2133 gnd 0.00488f
C4044 vdd.n2134 gnd 0.00488f
C4045 vdd.n2135 gnd 0.002622f
C4046 vdd.n2136 gnd 0.002776f
C4047 vdd.n2137 gnd 0.006198f
C4048 vdd.n2138 gnd 0.006198f
C4049 vdd.n2139 gnd 0.014653f
C4050 vdd.n2140 gnd 0.002699f
C4051 vdd.n2141 gnd 0.002622f
C4052 vdd.n2142 gnd 0.012613f
C4053 vdd.n2143 gnd 0.008806f
C4054 vdd.t142 gnd 0.03085f
C4055 vdd.t141 gnd 0.03085f
C4056 vdd.n2144 gnd 0.212021f
C4057 vdd.n2145 gnd 0.166722f
C4058 vdd.t104 gnd 0.03085f
C4059 vdd.t84 gnd 0.03085f
C4060 vdd.n2146 gnd 0.212021f
C4061 vdd.n2147 gnd 0.134544f
C4062 vdd.t80 gnd 0.03085f
C4063 vdd.t140 gnd 0.03085f
C4064 vdd.n2148 gnd 0.212021f
C4065 vdd.n2149 gnd 0.134544f
C4066 vdd.t118 gnd 0.03085f
C4067 vdd.t83 gnd 0.03085f
C4068 vdd.n2150 gnd 0.212021f
C4069 vdd.n2151 gnd 0.134544f
C4070 vdd.t74 gnd 0.03085f
C4071 vdd.t157 gnd 0.03085f
C4072 vdd.n2152 gnd 0.212021f
C4073 vdd.n2153 gnd 0.134544f
C4074 vdd.t156 gnd 0.03085f
C4075 vdd.t98 gnd 0.03085f
C4076 vdd.n2154 gnd 0.212021f
C4077 vdd.n2155 gnd 0.134544f
C4078 vdd.t108 gnd 0.03085f
C4079 vdd.t181 gnd 0.03085f
C4080 vdd.n2156 gnd 0.212021f
C4081 vdd.n2157 gnd 0.134544f
C4082 vdd.n2158 gnd 0.005259f
C4083 vdd.n2159 gnd 0.00488f
C4084 vdd.n2160 gnd 0.002699f
C4085 vdd.n2161 gnd 0.006198f
C4086 vdd.n2162 gnd 0.002622f
C4087 vdd.n2163 gnd 0.002776f
C4088 vdd.n2164 gnd 0.00488f
C4089 vdd.n2165 gnd 0.002622f
C4090 vdd.n2166 gnd 0.006198f
C4091 vdd.n2167 gnd 0.002776f
C4092 vdd.n2168 gnd 0.00488f
C4093 vdd.n2169 gnd 0.002622f
C4094 vdd.n2170 gnd 0.004648f
C4095 vdd.n2171 gnd 0.004662f
C4096 vdd.t135 gnd 0.013316f
C4097 vdd.n2172 gnd 0.029628f
C4098 vdd.n2173 gnd 0.154189f
C4099 vdd.n2174 gnd 0.002622f
C4100 vdd.n2175 gnd 0.002776f
C4101 vdd.n2176 gnd 0.006198f
C4102 vdd.n2177 gnd 0.006198f
C4103 vdd.n2178 gnd 0.002776f
C4104 vdd.n2179 gnd 0.002622f
C4105 vdd.n2180 gnd 0.00488f
C4106 vdd.n2181 gnd 0.00488f
C4107 vdd.n2182 gnd 0.002622f
C4108 vdd.n2183 gnd 0.002776f
C4109 vdd.n2184 gnd 0.006198f
C4110 vdd.n2185 gnd 0.006198f
C4111 vdd.n2186 gnd 0.002776f
C4112 vdd.n2187 gnd 0.002622f
C4113 vdd.n2188 gnd 0.00488f
C4114 vdd.n2189 gnd 0.00488f
C4115 vdd.n2190 gnd 0.002622f
C4116 vdd.n2191 gnd 0.002776f
C4117 vdd.n2192 gnd 0.006198f
C4118 vdd.n2193 gnd 0.006198f
C4119 vdd.n2194 gnd 0.014653f
C4120 vdd.n2195 gnd 0.002699f
C4121 vdd.n2196 gnd 0.002622f
C4122 vdd.n2197 gnd 0.012613f
C4123 vdd.n2198 gnd 0.008529f
C4124 vdd.n2199 gnd 0.05955f
C4125 vdd.n2200 gnd 0.240295f
C4126 vdd.n2201 gnd 2.63972f
C4127 vdd.n2202 gnd 0.565189f
C4128 vdd.n2203 gnd 0.007364f
C4129 vdd.n2204 gnd 0.009582f
C4130 vdd.n2205 gnd 0.007712f
C4131 vdd.n2206 gnd 0.009582f
C4132 vdd.n2207 gnd 0.768708f
C4133 vdd.n2208 gnd 0.009582f
C4134 vdd.n2209 gnd 0.007712f
C4135 vdd.n2210 gnd 0.009582f
C4136 vdd.n2211 gnd 0.009582f
C4137 vdd.n2212 gnd 0.009582f
C4138 vdd.n2213 gnd 0.007712f
C4139 vdd.n2214 gnd 0.009582f
C4140 vdd.t81 gnd 0.489623f
C4141 vdd.n2215 gnd 0.812775f
C4142 vdd.n2216 gnd 0.009582f
C4143 vdd.n2217 gnd 0.007712f
C4144 vdd.n2218 gnd 0.009582f
C4145 vdd.n2219 gnd 0.009582f
C4146 vdd.n2220 gnd 0.009582f
C4147 vdd.n2221 gnd 0.007712f
C4148 vdd.n2222 gnd 0.009582f
C4149 vdd.n2223 gnd 0.690369f
C4150 vdd.n2224 gnd 0.009582f
C4151 vdd.n2225 gnd 0.007712f
C4152 vdd.n2226 gnd 0.009582f
C4153 vdd.n2227 gnd 0.009582f
C4154 vdd.n2228 gnd 0.009582f
C4155 vdd.n2229 gnd 0.007712f
C4156 vdd.n2230 gnd 0.009582f
C4157 vdd.n2231 gnd 0.812775f
C4158 vdd.t64 gnd 0.489623f
C4159 vdd.n2232 gnd 0.523897f
C4160 vdd.n2233 gnd 0.009582f
C4161 vdd.n2234 gnd 0.007712f
C4162 vdd.n2235 gnd 0.009582f
C4163 vdd.n2236 gnd 0.009582f
C4164 vdd.n2237 gnd 0.009582f
C4165 vdd.n2238 gnd 0.007712f
C4166 vdd.n2239 gnd 0.009582f
C4167 vdd.n2240 gnd 0.621821f
C4168 vdd.n2241 gnd 0.009582f
C4169 vdd.n2242 gnd 0.007712f
C4170 vdd.n2243 gnd 0.009582f
C4171 vdd.n2244 gnd 0.009582f
C4172 vdd.n2245 gnd 0.009582f
C4173 vdd.n2246 gnd 0.007712f
C4174 vdd.n2247 gnd 0.009582f
C4175 vdd.n2248 gnd 0.514104f
C4176 vdd.n2249 gnd 0.788293f
C4177 vdd.n2250 gnd 0.009582f
C4178 vdd.n2251 gnd 0.007712f
C4179 vdd.n2252 gnd 0.009582f
C4180 vdd.n2253 gnd 0.009582f
C4181 vdd.n2254 gnd 0.009582f
C4182 vdd.n2255 gnd 0.007712f
C4183 vdd.n2256 gnd 0.009582f
C4184 vdd.n2257 gnd 0.954765f
C4185 vdd.n2258 gnd 0.009582f
C4186 vdd.n2259 gnd 0.007712f
C4187 vdd.n2260 gnd 0.009582f
C4188 vdd.n2261 gnd 0.009582f
C4189 vdd.n2262 gnd 0.021821f
C4190 vdd.n2263 gnd 0.009582f
C4191 vdd.n2264 gnd 0.009582f
C4192 vdd.n2265 gnd 0.007712f
C4193 vdd.n2266 gnd 0.009582f
C4194 vdd.t205 gnd 0.489623f
C4195 vdd.n2267 gnd 0.925388f
C4196 vdd.n2268 gnd 0.009582f
C4197 vdd.n2269 gnd 0.007712f
C4198 vdd.n2270 gnd 0.009582f
C4199 vdd.n2271 gnd 0.009582f
C4200 vdd.n2272 gnd 0.021821f
C4201 vdd.n2273 gnd 0.006401f
C4202 vdd.n2274 gnd 0.021821f
C4203 vdd.n2275 gnd 1.29261f
C4204 vdd.n2276 gnd 0.021821f
C4205 vdd.n2277 gnd 0.02197f
C4206 vdd.n2278 gnd 0.003663f
C4207 vdd.t228 gnd 0.117885f
C4208 vdd.t227 gnd 0.125987f
C4209 vdd.t226 gnd 0.153957f
C4210 vdd.n2279 gnd 0.19735f
C4211 vdd.n2280 gnd 0.16581f
C4212 vdd.n2281 gnd 0.011877f
C4213 vdd.n2282 gnd 0.004049f
C4214 vdd.n2283 gnd 0.008241f
C4215 vdd.n2284 gnd 1.01724f
C4216 vdd.n2286 gnd 0.007712f
C4217 vdd.n2287 gnd 0.007712f
C4218 vdd.n2288 gnd 0.009582f
C4219 vdd.n2290 gnd 0.009582f
C4220 vdd.n2291 gnd 0.009582f
C4221 vdd.n2292 gnd 0.007712f
C4222 vdd.n2293 gnd 0.007712f
C4223 vdd.n2294 gnd 0.007712f
C4224 vdd.n2295 gnd 0.009582f
C4225 vdd.n2297 gnd 0.009582f
C4226 vdd.n2298 gnd 0.009582f
C4227 vdd.n2299 gnd 0.007712f
C4228 vdd.n2300 gnd 0.007712f
C4229 vdd.n2301 gnd 0.007712f
C4230 vdd.n2302 gnd 0.009582f
C4231 vdd.n2304 gnd 0.009582f
C4232 vdd.n2305 gnd 0.009582f
C4233 vdd.n2306 gnd 0.007712f
C4234 vdd.n2307 gnd 0.007712f
C4235 vdd.n2308 gnd 0.007712f
C4236 vdd.n2309 gnd 0.009582f
C4237 vdd.n2311 gnd 0.009582f
C4238 vdd.n2312 gnd 0.009582f
C4239 vdd.n2313 gnd 0.007712f
C4240 vdd.n2314 gnd 0.009582f
C4241 vdd.n2315 gnd 0.009582f
C4242 vdd.n2316 gnd 0.009582f
C4243 vdd.n2317 gnd 0.015733f
C4244 vdd.n2318 gnd 0.005244f
C4245 vdd.n2319 gnd 0.007712f
C4246 vdd.n2320 gnd 0.009582f
C4247 vdd.n2322 gnd 0.009582f
C4248 vdd.n2323 gnd 0.009582f
C4249 vdd.n2324 gnd 0.007712f
C4250 vdd.n2325 gnd 0.007712f
C4251 vdd.n2326 gnd 0.007712f
C4252 vdd.n2327 gnd 0.009582f
C4253 vdd.n2329 gnd 0.009582f
C4254 vdd.n2330 gnd 0.009582f
C4255 vdd.n2331 gnd 0.007712f
C4256 vdd.n2332 gnd 0.007712f
C4257 vdd.n2333 gnd 0.007712f
C4258 vdd.n2334 gnd 0.009582f
C4259 vdd.n2336 gnd 0.009582f
C4260 vdd.n2337 gnd 0.009582f
C4261 vdd.n2338 gnd 0.007712f
C4262 vdd.n2339 gnd 0.007712f
C4263 vdd.n2340 gnd 0.007712f
C4264 vdd.n2341 gnd 0.009582f
C4265 vdd.n2343 gnd 0.009582f
C4266 vdd.n2344 gnd 0.009582f
C4267 vdd.n2345 gnd 0.007712f
C4268 vdd.n2346 gnd 0.007712f
C4269 vdd.n2347 gnd 0.007712f
C4270 vdd.n2348 gnd 0.009582f
C4271 vdd.n2350 gnd 0.009582f
C4272 vdd.n2351 gnd 0.009582f
C4273 vdd.n2352 gnd 0.007712f
C4274 vdd.n2353 gnd 0.009582f
C4275 vdd.n2354 gnd 0.009582f
C4276 vdd.n2355 gnd 0.009582f
C4277 vdd.n2356 gnd 0.015733f
C4278 vdd.n2357 gnd 0.00644f
C4279 vdd.n2358 gnd 0.007712f
C4280 vdd.n2359 gnd 0.009582f
C4281 vdd.n2361 gnd 0.009582f
C4282 vdd.n2362 gnd 0.009582f
C4283 vdd.n2363 gnd 0.007712f
C4284 vdd.n2364 gnd 0.007712f
C4285 vdd.n2365 gnd 0.007712f
C4286 vdd.n2366 gnd 0.009582f
C4287 vdd.n2368 gnd 0.009582f
C4288 vdd.n2369 gnd 0.009582f
C4289 vdd.n2370 gnd 0.007712f
C4290 vdd.n2371 gnd 0.007712f
C4291 vdd.n2372 gnd 0.007712f
C4292 vdd.n2373 gnd 0.009582f
C4293 vdd.n2375 gnd 0.009582f
C4294 vdd.n2376 gnd 0.009582f
C4295 vdd.n2377 gnd 0.007712f
C4296 vdd.n2378 gnd 0.007712f
C4297 vdd.n2379 gnd 0.007712f
C4298 vdd.n2380 gnd 0.009582f
C4299 vdd.n2382 gnd 0.009582f
C4300 vdd.n2383 gnd 0.007712f
C4301 vdd.n2384 gnd 0.007712f
C4302 vdd.n2385 gnd 0.009582f
C4303 vdd.n2387 gnd 0.009582f
C4304 vdd.n2388 gnd 0.009582f
C4305 vdd.n2389 gnd 0.007712f
C4306 vdd.n2390 gnd 0.008241f
C4307 vdd.n2391 gnd 1.01724f
C4308 vdd.n2392 gnd 0.043894f
C4309 vdd.n2393 gnd 0.006516f
C4310 vdd.n2394 gnd 0.006516f
C4311 vdd.n2395 gnd 0.006516f
C4312 vdd.n2396 gnd 0.006516f
C4313 vdd.n2397 gnd 0.006516f
C4314 vdd.n2398 gnd 0.006516f
C4315 vdd.n2399 gnd 0.006516f
C4316 vdd.n2400 gnd 0.006516f
C4317 vdd.n2401 gnd 0.006516f
C4318 vdd.n2402 gnd 0.006516f
C4319 vdd.n2403 gnd 0.006516f
C4320 vdd.n2404 gnd 0.006516f
C4321 vdd.n2405 gnd 0.006516f
C4322 vdd.n2406 gnd 0.006516f
C4323 vdd.n2407 gnd 0.006516f
C4324 vdd.n2408 gnd 0.006516f
C4325 vdd.n2409 gnd 0.006516f
C4326 vdd.n2410 gnd 0.006516f
C4327 vdd.n2411 gnd 0.006516f
C4328 vdd.n2412 gnd 0.006516f
C4329 vdd.n2413 gnd 0.006516f
C4330 vdd.n2414 gnd 0.006516f
C4331 vdd.n2415 gnd 0.006516f
C4332 vdd.n2416 gnd 0.006516f
C4333 vdd.n2417 gnd 0.006516f
C4334 vdd.n2418 gnd 0.006516f
C4335 vdd.n2419 gnd 0.006516f
C4336 vdd.n2420 gnd 0.006516f
C4337 vdd.n2421 gnd 0.006516f
C4338 vdd.n2422 gnd 0.006516f
C4339 vdd.n2423 gnd 11.5649f
C4340 vdd.n2425 gnd 0.014795f
C4341 vdd.n2426 gnd 0.014795f
C4342 vdd.n2427 gnd 0.013951f
C4343 vdd.n2428 gnd 0.006516f
C4344 vdd.n2429 gnd 0.006516f
C4345 vdd.n2430 gnd 0.665888f
C4346 vdd.n2431 gnd 0.006516f
C4347 vdd.n2432 gnd 0.006516f
C4348 vdd.n2433 gnd 0.006516f
C4349 vdd.n2434 gnd 0.006516f
C4350 vdd.n2435 gnd 0.006516f
C4351 vdd.n2436 gnd 0.523897f
C4352 vdd.n2437 gnd 0.006516f
C4353 vdd.n2438 gnd 0.006516f
C4354 vdd.n2439 gnd 0.006516f
C4355 vdd.n2440 gnd 0.006516f
C4356 vdd.n2441 gnd 0.006516f
C4357 vdd.n2442 gnd 0.665888f
C4358 vdd.n2443 gnd 0.006516f
C4359 vdd.n2444 gnd 0.006516f
C4360 vdd.n2445 gnd 0.006516f
C4361 vdd.n2446 gnd 0.006516f
C4362 vdd.n2447 gnd 0.006516f
C4363 vdd.n2448 gnd 0.665888f
C4364 vdd.n2449 gnd 0.006516f
C4365 vdd.n2450 gnd 0.006516f
C4366 vdd.n2451 gnd 0.006516f
C4367 vdd.n2452 gnd 0.006516f
C4368 vdd.n2453 gnd 0.006516f
C4369 vdd.n2454 gnd 0.641406f
C4370 vdd.n2455 gnd 0.006516f
C4371 vdd.n2456 gnd 0.006516f
C4372 vdd.n2457 gnd 0.006516f
C4373 vdd.n2458 gnd 0.006516f
C4374 vdd.n2459 gnd 0.006516f
C4375 vdd.n2460 gnd 0.494519f
C4376 vdd.n2461 gnd 0.006516f
C4377 vdd.n2462 gnd 0.006516f
C4378 vdd.n2463 gnd 0.006516f
C4379 vdd.n2464 gnd 0.006516f
C4380 vdd.n2465 gnd 0.006516f
C4381 vdd.n2466 gnd 0.347632f
C4382 vdd.n2467 gnd 0.006516f
C4383 vdd.n2468 gnd 0.006516f
C4384 vdd.n2469 gnd 0.006516f
C4385 vdd.n2470 gnd 0.006516f
C4386 vdd.n2471 gnd 0.006516f
C4387 vdd.n2472 gnd 0.465142f
C4388 vdd.n2473 gnd 0.006516f
C4389 vdd.n2474 gnd 0.006516f
C4390 vdd.n2475 gnd 0.006516f
C4391 vdd.n2476 gnd 0.006516f
C4392 vdd.n2477 gnd 0.006516f
C4393 vdd.n2478 gnd 0.612029f
C4394 vdd.n2479 gnd 0.006516f
C4395 vdd.n2480 gnd 0.006516f
C4396 vdd.n2481 gnd 0.006516f
C4397 vdd.n2482 gnd 0.006516f
C4398 vdd.n2483 gnd 0.006516f
C4399 vdd.n2484 gnd 0.665888f
C4400 vdd.n2485 gnd 0.006516f
C4401 vdd.n2486 gnd 0.006516f
C4402 vdd.n2487 gnd 0.006516f
C4403 vdd.n2488 gnd 0.006516f
C4404 vdd.n2489 gnd 0.006516f
C4405 vdd.n2490 gnd 0.572859f
C4406 vdd.n2491 gnd 0.006516f
C4407 vdd.n2492 gnd 0.006516f
C4408 vdd.n2493 gnd 0.005174f
C4409 vdd.n2494 gnd 0.018876f
C4410 vdd.n2495 gnd 0.004599f
C4411 vdd.n2496 gnd 0.006516f
C4412 vdd.n2497 gnd 0.425972f
C4413 vdd.n2498 gnd 0.006516f
C4414 vdd.n2499 gnd 0.006516f
C4415 vdd.n2500 gnd 0.006516f
C4416 vdd.n2501 gnd 0.006516f
C4417 vdd.n2502 gnd 0.006516f
C4418 vdd.n2503 gnd 0.386802f
C4419 vdd.n2504 gnd 0.006516f
C4420 vdd.n2505 gnd 0.006516f
C4421 vdd.n2506 gnd 0.006516f
C4422 vdd.n2507 gnd 0.006516f
C4423 vdd.n2508 gnd 0.006516f
C4424 vdd.n2509 gnd 0.533689f
C4425 vdd.n2510 gnd 0.006516f
C4426 vdd.n2511 gnd 0.006516f
C4427 vdd.n2512 gnd 0.006516f
C4428 vdd.n2513 gnd 0.006516f
C4429 vdd.n2514 gnd 0.006516f
C4430 vdd.n2515 gnd 0.587548f
C4431 vdd.n2516 gnd 0.006516f
C4432 vdd.n2517 gnd 0.006516f
C4433 vdd.n2518 gnd 0.006516f
C4434 vdd.n2519 gnd 0.006516f
C4435 vdd.n2520 gnd 0.006516f
C4436 vdd.n2521 gnd 0.440661f
C4437 vdd.n2522 gnd 0.006516f
C4438 vdd.n2523 gnd 0.006516f
C4439 vdd.n2524 gnd 0.006516f
C4440 vdd.n2525 gnd 0.006516f
C4441 vdd.n2526 gnd 0.006516f
C4442 vdd.n2527 gnd 0.210538f
C4443 vdd.n2528 gnd 0.006516f
C4444 vdd.n2529 gnd 0.006516f
C4445 vdd.n2530 gnd 0.006516f
C4446 vdd.n2531 gnd 0.006516f
C4447 vdd.n2532 gnd 0.006516f
C4448 vdd.n2533 gnd 0.210538f
C4449 vdd.n2534 gnd 0.006516f
C4450 vdd.n2535 gnd 0.006516f
C4451 vdd.n2536 gnd 0.006516f
C4452 vdd.n2537 gnd 0.006516f
C4453 vdd.n2538 gnd 0.006516f
C4454 vdd.n2539 gnd 0.665888f
C4455 vdd.n2540 gnd 0.006516f
C4456 vdd.n2541 gnd 0.006516f
C4457 vdd.n2542 gnd 0.006516f
C4458 vdd.n2543 gnd 0.006516f
C4459 vdd.n2544 gnd 0.006516f
C4460 vdd.n2545 gnd 0.006516f
C4461 vdd.n2546 gnd 0.006516f
C4462 vdd.n2547 gnd 0.460246f
C4463 vdd.n2548 gnd 0.006516f
C4464 vdd.n2549 gnd 0.006516f
C4465 vdd.n2550 gnd 0.006516f
C4466 vdd.n2551 gnd 0.006516f
C4467 vdd.n2552 gnd 0.006516f
C4468 vdd.n2553 gnd 0.006516f
C4469 vdd.n2554 gnd 0.41618f
C4470 vdd.n2555 gnd 0.006516f
C4471 vdd.n2556 gnd 0.006516f
C4472 vdd.n2557 gnd 0.006516f
C4473 vdd.n2558 gnd 0.014795f
C4474 vdd.n2559 gnd 0.013951f
C4475 vdd.n2560 gnd 0.006516f
C4476 vdd.n2561 gnd 0.006516f
C4477 vdd.n2562 gnd 0.005031f
C4478 vdd.n2563 gnd 0.006516f
C4479 vdd.n2564 gnd 0.006516f
C4480 vdd.n2565 gnd 0.004743f
C4481 vdd.n2566 gnd 0.006516f
C4482 vdd.n2567 gnd 0.006516f
C4483 vdd.n2568 gnd 0.006516f
C4484 vdd.n2569 gnd 0.006516f
C4485 vdd.n2570 gnd 0.006516f
C4486 vdd.n2571 gnd 0.006516f
C4487 vdd.n2572 gnd 0.006516f
C4488 vdd.n2573 gnd 0.006516f
C4489 vdd.n2574 gnd 0.006516f
C4490 vdd.n2575 gnd 0.006516f
C4491 vdd.n2576 gnd 0.006516f
C4492 vdd.n2577 gnd 0.006516f
C4493 vdd.n2578 gnd 0.006516f
C4494 vdd.n2579 gnd 0.006516f
C4495 vdd.n2580 gnd 0.006516f
C4496 vdd.n2581 gnd 0.006516f
C4497 vdd.n2582 gnd 0.006516f
C4498 vdd.n2583 gnd 0.006516f
C4499 vdd.n2584 gnd 0.006516f
C4500 vdd.n2585 gnd 0.006516f
C4501 vdd.n2586 gnd 0.006516f
C4502 vdd.n2587 gnd 0.006516f
C4503 vdd.n2588 gnd 0.006516f
C4504 vdd.n2589 gnd 0.006516f
C4505 vdd.n2590 gnd 0.006516f
C4506 vdd.n2591 gnd 0.006516f
C4507 vdd.n2592 gnd 0.006516f
C4508 vdd.n2593 gnd 0.006516f
C4509 vdd.n2594 gnd 0.006516f
C4510 vdd.n2595 gnd 0.006516f
C4511 vdd.n2596 gnd 0.006516f
C4512 vdd.n2597 gnd 0.006516f
C4513 vdd.n2598 gnd 0.006516f
C4514 vdd.n2599 gnd 0.006516f
C4515 vdd.n2600 gnd 0.006516f
C4516 vdd.n2601 gnd 0.006516f
C4517 vdd.n2602 gnd 0.006516f
C4518 vdd.n2603 gnd 0.006516f
C4519 vdd.n2604 gnd 0.006516f
C4520 vdd.n2605 gnd 0.006516f
C4521 vdd.n2606 gnd 0.006516f
C4522 vdd.n2607 gnd 0.006516f
C4523 vdd.n2608 gnd 0.006516f
C4524 vdd.n2609 gnd 0.006516f
C4525 vdd.n2610 gnd 0.006516f
C4526 vdd.n2611 gnd 0.006516f
C4527 vdd.n2612 gnd 0.006516f
C4528 vdd.n2613 gnd 0.006516f
C4529 vdd.n2614 gnd 0.006516f
C4530 vdd.n2615 gnd 0.006516f
C4531 vdd.n2616 gnd 0.006516f
C4532 vdd.n2617 gnd 0.006516f
C4533 vdd.n2618 gnd 0.006516f
C4534 vdd.n2619 gnd 0.006516f
C4535 vdd.n2620 gnd 0.006516f
C4536 vdd.n2621 gnd 0.006516f
C4537 vdd.n2622 gnd 0.006516f
C4538 vdd.n2623 gnd 0.006516f
C4539 vdd.n2624 gnd 0.006516f
C4540 vdd.n2625 gnd 0.006516f
C4541 vdd.n2626 gnd 0.014795f
C4542 vdd.n2627 gnd 0.013951f
C4543 vdd.n2628 gnd 0.013951f
C4544 vdd.n2629 gnd 0.75402f
C4545 vdd.n2630 gnd 0.013951f
C4546 vdd.n2631 gnd 0.014795f
C4547 vdd.n2632 gnd 0.013951f
C4548 vdd.n2633 gnd 0.006516f
C4549 vdd.n2634 gnd 0.006516f
C4550 vdd.n2635 gnd 0.006516f
C4551 vdd.n2636 gnd 0.005031f
C4552 vdd.n2637 gnd 0.009312f
C4553 vdd.n2638 gnd 0.004743f
C4554 vdd.n2639 gnd 0.006516f
C4555 vdd.n2640 gnd 0.006516f
C4556 vdd.n2641 gnd 0.006516f
C4557 vdd.n2642 gnd 0.006516f
C4558 vdd.n2643 gnd 0.006516f
C4559 vdd.n2644 gnd 0.006516f
C4560 vdd.n2645 gnd 0.006516f
C4561 vdd.n2646 gnd 0.006516f
C4562 vdd.n2647 gnd 0.006516f
C4563 vdd.n2648 gnd 0.006516f
C4564 vdd.n2649 gnd 0.006516f
C4565 vdd.n2650 gnd 0.006516f
C4566 vdd.n2651 gnd 0.006516f
C4567 vdd.n2652 gnd 0.006516f
C4568 vdd.n2653 gnd 0.006516f
C4569 vdd.n2654 gnd 0.006516f
C4570 vdd.n2655 gnd 0.006516f
C4571 vdd.n2656 gnd 0.006516f
C4572 vdd.n2657 gnd 0.006516f
C4573 vdd.n2658 gnd 0.006516f
C4574 vdd.n2659 gnd 0.006516f
C4575 vdd.n2660 gnd 0.006516f
C4576 vdd.n2661 gnd 0.006516f
C4577 vdd.n2662 gnd 0.006516f
C4578 vdd.n2663 gnd 0.006516f
C4579 vdd.n2664 gnd 0.006516f
C4580 vdd.n2665 gnd 0.006516f
C4581 vdd.n2666 gnd 0.006516f
C4582 vdd.n2667 gnd 0.006516f
C4583 vdd.n2668 gnd 0.006516f
C4584 vdd.n2669 gnd 0.006516f
C4585 vdd.n2670 gnd 0.006516f
C4586 vdd.n2671 gnd 0.006516f
C4587 vdd.n2672 gnd 0.006516f
C4588 vdd.n2673 gnd 0.006516f
C4589 vdd.n2674 gnd 0.006516f
C4590 vdd.n2675 gnd 0.006516f
C4591 vdd.n2676 gnd 0.006516f
C4592 vdd.n2677 gnd 0.006516f
C4593 vdd.n2678 gnd 0.006516f
C4594 vdd.n2679 gnd 0.006516f
C4595 vdd.n2680 gnd 0.006516f
C4596 vdd.n2681 gnd 0.006516f
C4597 vdd.n2682 gnd 0.006516f
C4598 vdd.n2683 gnd 0.006516f
C4599 vdd.n2684 gnd 0.006516f
C4600 vdd.n2685 gnd 0.006516f
C4601 vdd.n2686 gnd 0.006516f
C4602 vdd.n2687 gnd 0.006516f
C4603 vdd.n2688 gnd 0.006516f
C4604 vdd.n2689 gnd 0.006516f
C4605 vdd.n2690 gnd 0.006516f
C4606 vdd.n2691 gnd 0.006516f
C4607 vdd.n2692 gnd 0.006516f
C4608 vdd.n2693 gnd 0.006516f
C4609 vdd.n2694 gnd 0.006516f
C4610 vdd.n2695 gnd 0.006516f
C4611 vdd.n2696 gnd 0.006516f
C4612 vdd.n2697 gnd 0.006516f
C4613 vdd.n2698 gnd 0.006516f
C4614 vdd.n2699 gnd 0.014795f
C4615 vdd.n2700 gnd 0.014795f
C4616 vdd.n2701 gnd 0.812775f
C4617 vdd.t30 gnd 2.88878f
C4618 vdd.t17 gnd 2.88878f
C4619 vdd.n2735 gnd 0.014795f
C4620 vdd.t35 gnd 0.567963f
C4621 vdd.n2736 gnd 0.006516f
C4622 vdd.t254 gnd 0.263304f
C4623 vdd.t255 gnd 0.269524f
C4624 vdd.t252 gnd 0.171895f
C4625 vdd.n2737 gnd 0.0929f
C4626 vdd.n2738 gnd 0.052696f
C4627 vdd.n2739 gnd 0.006516f
C4628 vdd.t264 gnd 0.263304f
C4629 vdd.t265 gnd 0.269524f
C4630 vdd.t263 gnd 0.171895f
C4631 vdd.n2740 gnd 0.0929f
C4632 vdd.n2741 gnd 0.052696f
C4633 vdd.n2742 gnd 0.009312f
C4634 vdd.n2743 gnd 0.014795f
C4635 vdd.n2744 gnd 0.014795f
C4636 vdd.n2745 gnd 0.006516f
C4637 vdd.n2746 gnd 0.006516f
C4638 vdd.n2747 gnd 0.006516f
C4639 vdd.n2748 gnd 0.006516f
C4640 vdd.n2749 gnd 0.006516f
C4641 vdd.n2750 gnd 0.006516f
C4642 vdd.n2751 gnd 0.006516f
C4643 vdd.n2752 gnd 0.006516f
C4644 vdd.n2753 gnd 0.006516f
C4645 vdd.n2754 gnd 0.006516f
C4646 vdd.n2755 gnd 0.006516f
C4647 vdd.n2756 gnd 0.006516f
C4648 vdd.n2757 gnd 0.006516f
C4649 vdd.n2758 gnd 0.006516f
C4650 vdd.n2759 gnd 0.006516f
C4651 vdd.n2760 gnd 0.006516f
C4652 vdd.n2761 gnd 0.006516f
C4653 vdd.n2762 gnd 0.006516f
C4654 vdd.n2763 gnd 0.006516f
C4655 vdd.n2764 gnd 0.006516f
C4656 vdd.n2765 gnd 0.006516f
C4657 vdd.n2766 gnd 0.006516f
C4658 vdd.n2767 gnd 0.006516f
C4659 vdd.n2768 gnd 0.006516f
C4660 vdd.n2769 gnd 0.006516f
C4661 vdd.n2770 gnd 0.006516f
C4662 vdd.n2771 gnd 0.006516f
C4663 vdd.n2772 gnd 0.006516f
C4664 vdd.n2773 gnd 0.006516f
C4665 vdd.n2774 gnd 0.006516f
C4666 vdd.n2775 gnd 0.006516f
C4667 vdd.n2776 gnd 0.006516f
C4668 vdd.n2777 gnd 0.006516f
C4669 vdd.n2778 gnd 0.006516f
C4670 vdd.n2779 gnd 0.006516f
C4671 vdd.n2780 gnd 0.006516f
C4672 vdd.n2781 gnd 0.006516f
C4673 vdd.n2782 gnd 0.006516f
C4674 vdd.n2783 gnd 0.006516f
C4675 vdd.n2784 gnd 0.006516f
C4676 vdd.n2785 gnd 0.006516f
C4677 vdd.n2786 gnd 0.006516f
C4678 vdd.n2787 gnd 0.006516f
C4679 vdd.n2788 gnd 0.006516f
C4680 vdd.n2789 gnd 0.006516f
C4681 vdd.n2790 gnd 0.006516f
C4682 vdd.n2791 gnd 0.006516f
C4683 vdd.n2792 gnd 0.006516f
C4684 vdd.n2793 gnd 0.006516f
C4685 vdd.n2794 gnd 0.006516f
C4686 vdd.n2795 gnd 0.006516f
C4687 vdd.n2796 gnd 0.006516f
C4688 vdd.n2797 gnd 0.006516f
C4689 vdd.n2798 gnd 0.006516f
C4690 vdd.n2799 gnd 0.006516f
C4691 vdd.n2800 gnd 0.006516f
C4692 vdd.n2801 gnd 0.006516f
C4693 vdd.n2802 gnd 0.006516f
C4694 vdd.n2803 gnd 0.006516f
C4695 vdd.n2804 gnd 0.006516f
C4696 vdd.n2805 gnd 0.004743f
C4697 vdd.n2806 gnd 0.006516f
C4698 vdd.n2807 gnd 0.006516f
C4699 vdd.n2808 gnd 0.005031f
C4700 vdd.n2809 gnd 0.006516f
C4701 vdd.n2810 gnd 0.006516f
C4702 vdd.n2811 gnd 0.014795f
C4703 vdd.n2812 gnd 0.013951f
C4704 vdd.n2813 gnd 0.013951f
C4705 vdd.n2814 gnd 0.006516f
C4706 vdd.n2815 gnd 0.006516f
C4707 vdd.n2816 gnd 0.006516f
C4708 vdd.n2817 gnd 0.006516f
C4709 vdd.n2818 gnd 0.006516f
C4710 vdd.n2819 gnd 0.006516f
C4711 vdd.n2820 gnd 0.006516f
C4712 vdd.n2821 gnd 0.006516f
C4713 vdd.n2822 gnd 0.006516f
C4714 vdd.n2823 gnd 0.006516f
C4715 vdd.n2824 gnd 0.006516f
C4716 vdd.n2825 gnd 0.006516f
C4717 vdd.n2826 gnd 0.006516f
C4718 vdd.n2827 gnd 0.006516f
C4719 vdd.n2828 gnd 0.006516f
C4720 vdd.n2829 gnd 0.006516f
C4721 vdd.n2830 gnd 0.006516f
C4722 vdd.n2831 gnd 0.006516f
C4723 vdd.n2832 gnd 0.006516f
C4724 vdd.n2833 gnd 0.006516f
C4725 vdd.n2834 gnd 0.006516f
C4726 vdd.n2835 gnd 0.006516f
C4727 vdd.n2836 gnd 0.006516f
C4728 vdd.n2837 gnd 0.006516f
C4729 vdd.n2838 gnd 0.006516f
C4730 vdd.n2839 gnd 0.006516f
C4731 vdd.n2840 gnd 0.006516f
C4732 vdd.n2841 gnd 0.006516f
C4733 vdd.n2842 gnd 0.006516f
C4734 vdd.n2843 gnd 0.006516f
C4735 vdd.n2844 gnd 0.006516f
C4736 vdd.n2845 gnd 0.006516f
C4737 vdd.n2846 gnd 0.006516f
C4738 vdd.n2847 gnd 0.006516f
C4739 vdd.n2848 gnd 0.006516f
C4740 vdd.n2849 gnd 0.006516f
C4741 vdd.n2850 gnd 0.006516f
C4742 vdd.n2851 gnd 0.006516f
C4743 vdd.n2852 gnd 0.006516f
C4744 vdd.n2853 gnd 0.006516f
C4745 vdd.n2854 gnd 0.006516f
C4746 vdd.n2855 gnd 0.006516f
C4747 vdd.n2856 gnd 0.006516f
C4748 vdd.n2857 gnd 0.006516f
C4749 vdd.n2858 gnd 0.006516f
C4750 vdd.n2859 gnd 0.006516f
C4751 vdd.n2860 gnd 0.006516f
C4752 vdd.n2861 gnd 0.006516f
C4753 vdd.n2862 gnd 0.006516f
C4754 vdd.n2863 gnd 0.006516f
C4755 vdd.n2864 gnd 0.006516f
C4756 vdd.n2865 gnd 0.006516f
C4757 vdd.n2866 gnd 0.006516f
C4758 vdd.n2867 gnd 0.006516f
C4759 vdd.n2868 gnd 0.006516f
C4760 vdd.n2869 gnd 0.006516f
C4761 vdd.n2870 gnd 0.006516f
C4762 vdd.n2871 gnd 0.006516f
C4763 vdd.n2872 gnd 0.006516f
C4764 vdd.n2873 gnd 0.006516f
C4765 vdd.n2874 gnd 0.006516f
C4766 vdd.n2875 gnd 0.006516f
C4767 vdd.n2876 gnd 0.006516f
C4768 vdd.n2877 gnd 0.006516f
C4769 vdd.n2878 gnd 0.006516f
C4770 vdd.n2879 gnd 0.006516f
C4771 vdd.n2880 gnd 0.006516f
C4772 vdd.n2881 gnd 0.006516f
C4773 vdd.n2882 gnd 0.006516f
C4774 vdd.n2883 gnd 0.006516f
C4775 vdd.n2884 gnd 0.006516f
C4776 vdd.n2885 gnd 0.006516f
C4777 vdd.n2886 gnd 0.006516f
C4778 vdd.n2887 gnd 0.006516f
C4779 vdd.n2888 gnd 0.006516f
C4780 vdd.n2889 gnd 0.006516f
C4781 vdd.n2890 gnd 0.006516f
C4782 vdd.n2891 gnd 0.006516f
C4783 vdd.n2892 gnd 0.006516f
C4784 vdd.n2893 gnd 0.006516f
C4785 vdd.n2894 gnd 0.006516f
C4786 vdd.n2895 gnd 0.006516f
C4787 vdd.n2896 gnd 0.006516f
C4788 vdd.n2897 gnd 0.006516f
C4789 vdd.n2898 gnd 0.006516f
C4790 vdd.n2899 gnd 0.006516f
C4791 vdd.n2900 gnd 0.006516f
C4792 vdd.n2901 gnd 0.006516f
C4793 vdd.n2902 gnd 0.006516f
C4794 vdd.n2903 gnd 0.006516f
C4795 vdd.n2904 gnd 0.006516f
C4796 vdd.n2905 gnd 0.006516f
C4797 vdd.n2906 gnd 0.006516f
C4798 vdd.n2907 gnd 0.006516f
C4799 vdd.n2908 gnd 0.006516f
C4800 vdd.n2909 gnd 0.006516f
C4801 vdd.n2910 gnd 0.006516f
C4802 vdd.n2911 gnd 0.006516f
C4803 vdd.n2912 gnd 0.006516f
C4804 vdd.n2913 gnd 0.006516f
C4805 vdd.n2914 gnd 0.006516f
C4806 vdd.n2915 gnd 0.210538f
C4807 vdd.n2916 gnd 0.006516f
C4808 vdd.n2917 gnd 0.006516f
C4809 vdd.n2918 gnd 0.006516f
C4810 vdd.n2919 gnd 0.006516f
C4811 vdd.n2920 gnd 0.006516f
C4812 vdd.n2921 gnd 0.210538f
C4813 vdd.n2922 gnd 0.006516f
C4814 vdd.n2923 gnd 0.006516f
C4815 vdd.n2924 gnd 0.006516f
C4816 vdd.n2925 gnd 0.006516f
C4817 vdd.n2926 gnd 0.006516f
C4818 vdd.n2927 gnd 0.006516f
C4819 vdd.n2928 gnd 0.006516f
C4820 vdd.n2929 gnd 0.006516f
C4821 vdd.n2930 gnd 0.006516f
C4822 vdd.n2931 gnd 0.006516f
C4823 vdd.n2932 gnd 0.006516f
C4824 vdd.n2933 gnd 0.41618f
C4825 vdd.n2934 gnd 0.006516f
C4826 vdd.n2935 gnd 0.006516f
C4827 vdd.n2936 gnd 0.006516f
C4828 vdd.n2937 gnd 0.013951f
C4829 vdd.n2938 gnd 0.013951f
C4830 vdd.n2939 gnd 0.014795f
C4831 vdd.n2940 gnd 0.014795f
C4832 vdd.n2941 gnd 0.006516f
C4833 vdd.n2942 gnd 0.006516f
C4834 vdd.n2943 gnd 0.006516f
C4835 vdd.n2944 gnd 0.005031f
C4836 vdd.n2945 gnd 0.009312f
C4837 vdd.n2946 gnd 0.004743f
C4838 vdd.n2947 gnd 0.006516f
C4839 vdd.n2948 gnd 0.006516f
C4840 vdd.n2949 gnd 0.006516f
C4841 vdd.n2950 gnd 0.006516f
C4842 vdd.n2951 gnd 0.006516f
C4843 vdd.n2952 gnd 0.006516f
C4844 vdd.n2953 gnd 0.006516f
C4845 vdd.n2954 gnd 0.006516f
C4846 vdd.n2955 gnd 0.006516f
C4847 vdd.n2956 gnd 0.006516f
C4848 vdd.n2957 gnd 0.006516f
C4849 vdd.n2958 gnd 0.006516f
C4850 vdd.n2959 gnd 0.006516f
C4851 vdd.n2960 gnd 0.006516f
C4852 vdd.n2961 gnd 0.006516f
C4853 vdd.n2962 gnd 0.006516f
C4854 vdd.n2963 gnd 0.006516f
C4855 vdd.n2964 gnd 0.006516f
C4856 vdd.n2965 gnd 0.006516f
C4857 vdd.n2966 gnd 0.006516f
C4858 vdd.n2967 gnd 0.006516f
C4859 vdd.n2968 gnd 0.006516f
C4860 vdd.n2969 gnd 0.006516f
C4861 vdd.n2970 gnd 0.006516f
C4862 vdd.n2971 gnd 0.006516f
C4863 vdd.n2972 gnd 0.006516f
C4864 vdd.n2973 gnd 0.006516f
C4865 vdd.n2974 gnd 0.006516f
C4866 vdd.n2975 gnd 0.006516f
C4867 vdd.n2976 gnd 0.006516f
C4868 vdd.n2977 gnd 0.006516f
C4869 vdd.n2978 gnd 0.006516f
C4870 vdd.n2979 gnd 0.006516f
C4871 vdd.n2980 gnd 0.006516f
C4872 vdd.n2981 gnd 0.006516f
C4873 vdd.n2982 gnd 0.006516f
C4874 vdd.n2983 gnd 0.006516f
C4875 vdd.n2984 gnd 0.006516f
C4876 vdd.n2985 gnd 0.006516f
C4877 vdd.n2986 gnd 0.006516f
C4878 vdd.n2987 gnd 0.006516f
C4879 vdd.n2988 gnd 0.006516f
C4880 vdd.n2989 gnd 0.006516f
C4881 vdd.n2990 gnd 0.006516f
C4882 vdd.n2991 gnd 0.006516f
C4883 vdd.n2992 gnd 0.006516f
C4884 vdd.n2993 gnd 0.006516f
C4885 vdd.n2994 gnd 0.006516f
C4886 vdd.n2995 gnd 0.006516f
C4887 vdd.n2996 gnd 0.006516f
C4888 vdd.n2997 gnd 0.006516f
C4889 vdd.n2998 gnd 0.006516f
C4890 vdd.n2999 gnd 0.006516f
C4891 vdd.n3000 gnd 0.006516f
C4892 vdd.n3001 gnd 0.006516f
C4893 vdd.n3002 gnd 0.006516f
C4894 vdd.n3003 gnd 0.006516f
C4895 vdd.n3004 gnd 0.006516f
C4896 vdd.n3005 gnd 0.812775f
C4897 vdd.n3007 gnd 0.014795f
C4898 vdd.n3008 gnd 0.014795f
C4899 vdd.n3009 gnd 0.013951f
C4900 vdd.n3010 gnd 0.006516f
C4901 vdd.n3011 gnd 0.006516f
C4902 vdd.n3012 gnd 0.391699f
C4903 vdd.n3013 gnd 0.006516f
C4904 vdd.n3014 gnd 0.006516f
C4905 vdd.n3015 gnd 0.006516f
C4906 vdd.n3016 gnd 0.006516f
C4907 vdd.n3017 gnd 0.006516f
C4908 vdd.n3018 gnd 0.396595f
C4909 vdd.n3019 gnd 0.006516f
C4910 vdd.n3020 gnd 0.006516f
C4911 vdd.n3021 gnd 0.006516f
C4912 vdd.n3022 gnd 0.006516f
C4913 vdd.n3023 gnd 0.006516f
C4914 vdd.n3024 gnd 0.665888f
C4915 vdd.n3025 gnd 0.006516f
C4916 vdd.n3026 gnd 0.006516f
C4917 vdd.n3027 gnd 0.006516f
C4918 vdd.n3028 gnd 0.006516f
C4919 vdd.n3029 gnd 0.006516f
C4920 vdd.n3030 gnd 0.479831f
C4921 vdd.n3031 gnd 0.006516f
C4922 vdd.n3032 gnd 0.006516f
C4923 vdd.n3033 gnd 0.006516f
C4924 vdd.n3034 gnd 0.006516f
C4925 vdd.n3035 gnd 0.006516f
C4926 vdd.n3036 gnd 0.602237f
C4927 vdd.n3037 gnd 0.006516f
C4928 vdd.n3038 gnd 0.006516f
C4929 vdd.n3039 gnd 0.006516f
C4930 vdd.n3040 gnd 0.006516f
C4931 vdd.n3041 gnd 0.006516f
C4932 vdd.n3042 gnd 0.494519f
C4933 vdd.n3043 gnd 0.006516f
C4934 vdd.n3044 gnd 0.006516f
C4935 vdd.n3045 gnd 0.006516f
C4936 vdd.n3046 gnd 0.006516f
C4937 vdd.n3047 gnd 0.006516f
C4938 vdd.n3048 gnd 0.347632f
C4939 vdd.n3049 gnd 0.006516f
C4940 vdd.n3050 gnd 0.006516f
C4941 vdd.n3051 gnd 0.006516f
C4942 vdd.n3052 gnd 0.006516f
C4943 vdd.n3053 gnd 0.006516f
C4944 vdd.n3054 gnd 0.210538f
C4945 vdd.n3055 gnd 0.006516f
C4946 vdd.n3056 gnd 0.006516f
C4947 vdd.n3057 gnd 0.006516f
C4948 vdd.n3058 gnd 0.006516f
C4949 vdd.n3059 gnd 0.006516f
C4950 vdd.n3060 gnd 0.612029f
C4951 vdd.n3061 gnd 0.006516f
C4952 vdd.n3062 gnd 0.006516f
C4953 vdd.n3063 gnd 0.006516f
C4954 vdd.n3064 gnd 0.004599f
C4955 vdd.n3065 gnd 0.006516f
C4956 vdd.n3066 gnd 0.006516f
C4957 vdd.n3067 gnd 0.665888f
C4958 vdd.n3068 gnd 0.006516f
C4959 vdd.n3069 gnd 0.006516f
C4960 vdd.n3070 gnd 0.006516f
C4961 vdd.n3071 gnd 0.006516f
C4962 vdd.n3072 gnd 0.006516f
C4963 vdd.n3073 gnd 0.528793f
C4964 vdd.n3074 gnd 0.006516f
C4965 vdd.n3075 gnd 0.005174f
C4966 vdd.n3076 gnd 0.006516f
C4967 vdd.n3077 gnd 0.006516f
C4968 vdd.n3078 gnd 0.006516f
C4969 vdd.n3079 gnd 0.425972f
C4970 vdd.n3080 gnd 0.006516f
C4971 vdd.n3081 gnd 0.006516f
C4972 vdd.n3082 gnd 0.006516f
C4973 vdd.n3083 gnd 0.006516f
C4974 vdd.n3084 gnd 0.006516f
C4975 vdd.n3085 gnd 0.386802f
C4976 vdd.n3086 gnd 0.006516f
C4977 vdd.n3087 gnd 0.006516f
C4978 vdd.n3088 gnd 0.006516f
C4979 vdd.n3089 gnd 0.006516f
C4980 vdd.n3090 gnd 0.006516f
C4981 vdd.n3091 gnd 0.533689f
C4982 vdd.n3092 gnd 0.006516f
C4983 vdd.n3093 gnd 0.006516f
C4984 vdd.n3094 gnd 0.006516f
C4985 vdd.n3095 gnd 0.006516f
C4986 vdd.n3096 gnd 0.006516f
C4987 vdd.n3097 gnd 0.665888f
C4988 vdd.n3098 gnd 0.006516f
C4989 vdd.n3099 gnd 0.006516f
C4990 vdd.n3100 gnd 0.006516f
C4991 vdd.n3101 gnd 0.006516f
C4992 vdd.n3102 gnd 0.006516f
C4993 vdd.n3103 gnd 0.651199f
C4994 vdd.n3104 gnd 0.006516f
C4995 vdd.n3105 gnd 0.006516f
C4996 vdd.n3106 gnd 0.006516f
C4997 vdd.n3107 gnd 0.006516f
C4998 vdd.n3108 gnd 0.006516f
C4999 vdd.n3109 gnd 0.504312f
C5000 vdd.n3110 gnd 0.006516f
C5001 vdd.n3111 gnd 0.006516f
C5002 vdd.n3112 gnd 0.006516f
C5003 vdd.n3113 gnd 0.006516f
C5004 vdd.n3114 gnd 0.006516f
C5005 vdd.n3115 gnd 0.357425f
C5006 vdd.n3116 gnd 0.006516f
C5007 vdd.n3117 gnd 0.006516f
C5008 vdd.n3118 gnd 0.006516f
C5009 vdd.n3119 gnd 0.006516f
C5010 vdd.n3120 gnd 0.006516f
C5011 vdd.n3121 gnd 0.665888f
C5012 vdd.n3122 gnd 0.006516f
C5013 vdd.n3123 gnd 0.006516f
C5014 vdd.n3124 gnd 0.006516f
C5015 vdd.n3125 gnd 0.006516f
C5016 vdd.n3126 gnd 0.006516f
C5017 vdd.n3127 gnd 0.006516f
C5018 vdd.n3129 gnd 0.006516f
C5019 vdd.n3130 gnd 0.006516f
C5020 vdd.n3132 gnd 0.006516f
C5021 vdd.n3133 gnd 0.006516f
C5022 vdd.n3136 gnd 0.006516f
C5023 vdd.n3137 gnd 0.006516f
C5024 vdd.n3138 gnd 0.006516f
C5025 vdd.n3139 gnd 0.006516f
C5026 vdd.n3141 gnd 0.006516f
C5027 vdd.n3142 gnd 0.006516f
C5028 vdd.n3143 gnd 0.006516f
C5029 vdd.n3144 gnd 0.006516f
C5030 vdd.n3145 gnd 0.006516f
C5031 vdd.n3146 gnd 0.006516f
C5032 vdd.n3148 gnd 0.006516f
C5033 vdd.n3149 gnd 0.006516f
C5034 vdd.n3150 gnd 0.006516f
C5035 vdd.n3151 gnd 0.006516f
C5036 vdd.n3152 gnd 0.006516f
C5037 vdd.n3153 gnd 0.006516f
C5038 vdd.n3155 gnd 0.006516f
C5039 vdd.n3156 gnd 0.006516f
C5040 vdd.n3157 gnd 0.006516f
C5041 vdd.n3158 gnd 0.006516f
C5042 vdd.n3159 gnd 0.006516f
C5043 vdd.n3160 gnd 0.006516f
C5044 vdd.n3162 gnd 0.006516f
C5045 vdd.n3163 gnd 0.014795f
C5046 vdd.n3164 gnd 0.014795f
C5047 vdd.n3165 gnd 0.013951f
C5048 vdd.n3166 gnd 0.006516f
C5049 vdd.n3167 gnd 0.006516f
C5050 vdd.n3168 gnd 0.006516f
C5051 vdd.n3169 gnd 0.006516f
C5052 vdd.n3170 gnd 0.006516f
C5053 vdd.n3171 gnd 0.006516f
C5054 vdd.n3172 gnd 0.665888f
C5055 vdd.n3173 gnd 0.006516f
C5056 vdd.n3174 gnd 0.006516f
C5057 vdd.n3175 gnd 0.006516f
C5058 vdd.n3176 gnd 0.006516f
C5059 vdd.n3177 gnd 0.006516f
C5060 vdd.n3178 gnd 0.474935f
C5061 vdd.n3179 gnd 0.006516f
C5062 vdd.n3180 gnd 0.006516f
C5063 vdd.n3181 gnd 0.006516f
C5064 vdd.n3182 gnd 0.014795f
C5065 vdd.n3184 gnd 0.014795f
C5066 vdd.n3185 gnd 0.013951f
C5067 vdd.n3186 gnd 0.006516f
C5068 vdd.n3187 gnd 0.005031f
C5069 vdd.n3188 gnd 0.006516f
C5070 vdd.n3190 gnd 0.006516f
C5071 vdd.n3191 gnd 0.006516f
C5072 vdd.n3192 gnd 0.006516f
C5073 vdd.n3193 gnd 0.006516f
C5074 vdd.n3194 gnd 0.006516f
C5075 vdd.n3195 gnd 0.006516f
C5076 vdd.n3197 gnd 0.006516f
C5077 vdd.n3198 gnd 0.006516f
C5078 vdd.n3199 gnd 0.006516f
C5079 vdd.n3200 gnd 0.006516f
C5080 vdd.n3201 gnd 0.006516f
C5081 vdd.n3202 gnd 0.006516f
C5082 vdd.n3204 gnd 0.006516f
C5083 vdd.n3205 gnd 0.006516f
C5084 vdd.n3206 gnd 0.006516f
C5085 vdd.n3207 gnd 0.006516f
C5086 vdd.n3208 gnd 0.006516f
C5087 vdd.n3209 gnd 0.006516f
C5088 vdd.n3211 gnd 0.006516f
C5089 vdd.n3212 gnd 0.006516f
C5090 vdd.n3213 gnd 0.006516f
C5091 vdd.n3214 gnd 1.0209f
C5092 vdd.n3215 gnd 0.040234f
C5093 vdd.n3216 gnd 0.006516f
C5094 vdd.n3217 gnd 0.006516f
C5095 vdd.n3219 gnd 0.006516f
C5096 vdd.n3220 gnd 0.006516f
C5097 vdd.n3221 gnd 0.006516f
C5098 vdd.n3222 gnd 0.006516f
C5099 vdd.n3223 gnd 0.006516f
C5100 vdd.n3224 gnd 0.006516f
C5101 vdd.n3226 gnd 0.006516f
C5102 vdd.n3227 gnd 0.006516f
C5103 vdd.n3228 gnd 0.006516f
C5104 vdd.n3229 gnd 0.006516f
C5105 vdd.n3230 gnd 0.006516f
C5106 vdd.n3231 gnd 0.006516f
C5107 vdd.n3233 gnd 0.006516f
C5108 vdd.n3234 gnd 0.006516f
C5109 vdd.n3235 gnd 0.006516f
C5110 vdd.n3236 gnd 0.006516f
C5111 vdd.n3237 gnd 0.006516f
C5112 vdd.n3238 gnd 0.006516f
C5113 vdd.n3240 gnd 0.006516f
C5114 vdd.n3241 gnd 0.006516f
C5115 vdd.n3243 gnd 0.006516f
C5116 vdd.n3244 gnd 0.006516f
C5117 vdd.n3245 gnd 0.014795f
C5118 vdd.n3246 gnd 0.013951f
C5119 vdd.n3247 gnd 0.013951f
C5120 vdd.n3248 gnd 0.900907f
C5121 vdd.n3249 gnd 0.013951f
C5122 vdd.n3250 gnd 0.014795f
C5123 vdd.n3251 gnd 0.013951f
C5124 vdd.n3252 gnd 0.006516f
C5125 vdd.n3253 gnd 0.005031f
C5126 vdd.n3254 gnd 0.006516f
C5127 vdd.n3256 gnd 0.006516f
C5128 vdd.n3257 gnd 0.006516f
C5129 vdd.n3258 gnd 0.006516f
C5130 vdd.n3259 gnd 0.006516f
C5131 vdd.n3260 gnd 0.006516f
C5132 vdd.n3261 gnd 0.006516f
C5133 vdd.n3263 gnd 0.006516f
C5134 vdd.n3264 gnd 0.006516f
C5135 vdd.n3265 gnd 0.006516f
C5136 vdd.n3266 gnd 0.006516f
C5137 vdd.n3267 gnd 0.006516f
C5138 vdd.n3268 gnd 0.006516f
C5139 vdd.n3270 gnd 0.006516f
C5140 vdd.n3271 gnd 0.006516f
C5141 vdd.n3272 gnd 0.006516f
C5142 vdd.n3273 gnd 0.006516f
C5143 vdd.n3274 gnd 0.006516f
C5144 vdd.n3275 gnd 0.006516f
C5145 vdd.n3277 gnd 0.006516f
C5146 vdd.n3278 gnd 0.006516f
C5147 vdd.n3280 gnd 0.006516f
C5148 vdd.n3281 gnd 0.040234f
C5149 vdd.n3282 gnd 1.0209f
C5150 vdd.n3283 gnd 0.008241f
C5151 vdd.n3284 gnd 0.003663f
C5152 vdd.t220 gnd 0.117885f
C5153 vdd.t221 gnd 0.125987f
C5154 vdd.t218 gnd 0.153957f
C5155 vdd.n3285 gnd 0.19735f
C5156 vdd.n3286 gnd 0.16581f
C5157 vdd.n3287 gnd 0.011877f
C5158 vdd.n3288 gnd 0.009582f
C5159 vdd.n3289 gnd 0.004049f
C5160 vdd.n3290 gnd 0.007712f
C5161 vdd.n3291 gnd 0.009582f
C5162 vdd.n3292 gnd 0.009582f
C5163 vdd.n3293 gnd 0.007712f
C5164 vdd.n3294 gnd 0.007712f
C5165 vdd.n3295 gnd 0.009582f
C5166 vdd.n3297 gnd 0.009582f
C5167 vdd.n3298 gnd 0.007712f
C5168 vdd.n3299 gnd 0.007712f
C5169 vdd.n3300 gnd 0.007712f
C5170 vdd.n3301 gnd 0.009582f
C5171 vdd.n3303 gnd 0.009582f
C5172 vdd.n3305 gnd 0.009582f
C5173 vdd.n3306 gnd 0.007712f
C5174 vdd.n3307 gnd 0.007712f
C5175 vdd.n3308 gnd 0.007712f
C5176 vdd.n3309 gnd 0.009582f
C5177 vdd.n3311 gnd 0.009582f
C5178 vdd.n3313 gnd 0.009582f
C5179 vdd.n3314 gnd 0.007712f
C5180 vdd.n3315 gnd 0.007712f
C5181 vdd.n3316 gnd 0.007712f
C5182 vdd.n3317 gnd 0.009582f
C5183 vdd.n3319 gnd 0.009582f
C5184 vdd.n3320 gnd 0.009582f
C5185 vdd.n3321 gnd 0.007712f
C5186 vdd.n3322 gnd 0.007712f
C5187 vdd.n3323 gnd 0.009582f
C5188 vdd.n3324 gnd 0.009582f
C5189 vdd.n3326 gnd 0.009582f
C5190 vdd.n3327 gnd 0.007712f
C5191 vdd.n3328 gnd 0.009582f
C5192 vdd.n3329 gnd 0.009582f
C5193 vdd.n3330 gnd 0.009582f
C5194 vdd.n3331 gnd 0.015733f
C5195 vdd.n3332 gnd 0.005244f
C5196 vdd.n3333 gnd 0.009582f
C5197 vdd.n3335 gnd 0.009582f
C5198 vdd.n3337 gnd 0.009582f
C5199 vdd.n3338 gnd 0.007712f
C5200 vdd.n3339 gnd 0.007712f
C5201 vdd.n3340 gnd 0.007712f
C5202 vdd.n3341 gnd 0.009582f
C5203 vdd.n3343 gnd 0.009582f
C5204 vdd.n3345 gnd 0.009582f
C5205 vdd.n3346 gnd 0.007712f
C5206 vdd.n3347 gnd 0.007712f
C5207 vdd.n3348 gnd 0.007712f
C5208 vdd.n3349 gnd 0.009582f
C5209 vdd.n3351 gnd 0.009582f
C5210 vdd.n3353 gnd 0.009582f
C5211 vdd.n3354 gnd 0.007712f
C5212 vdd.n3355 gnd 0.007712f
C5213 vdd.n3356 gnd 0.007712f
C5214 vdd.n3357 gnd 0.009582f
C5215 vdd.n3359 gnd 0.009582f
C5216 vdd.n3361 gnd 0.009582f
C5217 vdd.n3362 gnd 0.007712f
C5218 vdd.n3363 gnd 0.007712f
C5219 vdd.n3364 gnd 0.007712f
C5220 vdd.n3365 gnd 0.009582f
C5221 vdd.n3367 gnd 0.009582f
C5222 vdd.n3369 gnd 0.009582f
C5223 vdd.n3370 gnd 0.007712f
C5224 vdd.n3371 gnd 0.007712f
C5225 vdd.n3372 gnd 0.00644f
C5226 vdd.n3373 gnd 0.009582f
C5227 vdd.n3375 gnd 0.009582f
C5228 vdd.n3377 gnd 0.009582f
C5229 vdd.n3378 gnd 0.00644f
C5230 vdd.n3379 gnd 0.007712f
C5231 vdd.n3380 gnd 0.007712f
C5232 vdd.n3381 gnd 0.009582f
C5233 vdd.n3383 gnd 0.009582f
C5234 vdd.n3385 gnd 0.009582f
C5235 vdd.n3386 gnd 0.007712f
C5236 vdd.n3387 gnd 0.007712f
C5237 vdd.n3388 gnd 0.007712f
C5238 vdd.n3389 gnd 0.009582f
C5239 vdd.n3391 gnd 0.009582f
C5240 vdd.n3393 gnd 0.009582f
C5241 vdd.n3394 gnd 0.007712f
C5242 vdd.n3395 gnd 0.007712f
C5243 vdd.n3396 gnd 0.007712f
C5244 vdd.n3397 gnd 0.009582f
C5245 vdd.n3399 gnd 0.009582f
C5246 vdd.n3400 gnd 0.009582f
C5247 vdd.n3401 gnd 0.007712f
C5248 vdd.n3402 gnd 0.007712f
C5249 vdd.n3403 gnd 0.009582f
C5250 vdd.n3404 gnd 0.009582f
C5251 vdd.n3405 gnd 0.007712f
C5252 vdd.n3406 gnd 0.007712f
C5253 vdd.n3407 gnd 0.009582f
C5254 vdd.n3408 gnd 0.009582f
C5255 vdd.n3410 gnd 0.009582f
C5256 vdd.n3411 gnd 0.007712f
C5257 vdd.n3412 gnd 0.006401f
C5258 vdd.n3413 gnd 0.02197f
C5259 vdd.n3414 gnd 0.021821f
C5260 vdd.n3415 gnd 0.006401f
C5261 vdd.n3416 gnd 0.021821f
C5262 vdd.n3417 gnd 1.29261f
C5263 vdd.n3418 gnd 0.021821f
C5264 vdd.n3419 gnd 0.006401f
C5265 vdd.n3420 gnd 0.021821f
C5266 vdd.n3421 gnd 0.009582f
C5267 vdd.n3422 gnd 0.009582f
C5268 vdd.n3423 gnd 0.007712f
C5269 vdd.n3424 gnd 0.009582f
C5270 vdd.n3425 gnd 0.925388f
C5271 vdd.n3426 gnd 0.009582f
C5272 vdd.n3427 gnd 0.007712f
C5273 vdd.n3428 gnd 0.009582f
C5274 vdd.n3429 gnd 0.009582f
C5275 vdd.n3430 gnd 0.009582f
C5276 vdd.n3431 gnd 0.007712f
C5277 vdd.n3432 gnd 0.009582f
C5278 vdd.n3433 gnd 0.954765f
C5279 vdd.n3434 gnd 0.009582f
C5280 vdd.n3435 gnd 0.007712f
C5281 vdd.n3436 gnd 0.009582f
C5282 vdd.n3437 gnd 0.009582f
C5283 vdd.n3438 gnd 0.009582f
C5284 vdd.n3439 gnd 0.007712f
C5285 vdd.n3440 gnd 0.009582f
C5286 vdd.t95 gnd 0.489623f
C5287 vdd.n3441 gnd 0.788293f
C5288 vdd.n3442 gnd 0.009582f
C5289 vdd.n3443 gnd 0.007712f
C5290 vdd.n3444 gnd 0.009582f
C5291 vdd.n3445 gnd 0.009582f
C5292 vdd.n3446 gnd 0.009582f
C5293 vdd.n3447 gnd 0.007712f
C5294 vdd.n3448 gnd 0.009582f
C5295 vdd.n3449 gnd 0.621821f
C5296 vdd.n3450 gnd 0.009582f
C5297 vdd.n3451 gnd 0.007712f
C5298 vdd.n3452 gnd 0.009582f
C5299 vdd.n3453 gnd 0.009582f
C5300 vdd.n3454 gnd 0.009582f
C5301 vdd.n3455 gnd 0.007712f
C5302 vdd.n3456 gnd 0.009582f
C5303 vdd.n3457 gnd 0.778501f
C5304 vdd.n3458 gnd 0.523897f
C5305 vdd.n3459 gnd 0.009582f
C5306 vdd.n3460 gnd 0.007712f
C5307 vdd.n3461 gnd 0.009582f
C5308 vdd.n3462 gnd 0.009582f
C5309 vdd.n3463 gnd 0.009582f
C5310 vdd.n3464 gnd 0.007712f
C5311 vdd.n3465 gnd 0.009582f
C5312 vdd.n3466 gnd 0.690369f
C5313 vdd.n3467 gnd 0.009582f
C5314 vdd.n3468 gnd 0.007712f
C5315 vdd.n3469 gnd 0.009582f
C5316 vdd.n3470 gnd 0.009582f
C5317 vdd.n3471 gnd 0.009582f
C5318 vdd.n3472 gnd 0.009582f
C5319 vdd.n3473 gnd 0.009582f
C5320 vdd.n3474 gnd 0.007712f
C5321 vdd.n3475 gnd 0.007712f
C5322 vdd.n3476 gnd 0.009582f
C5323 vdd.t119 gnd 0.489623f
C5324 vdd.n3477 gnd 0.812775f
C5325 vdd.n3478 gnd 0.009582f
C5326 vdd.n3479 gnd 0.007712f
C5327 vdd.n3480 gnd 0.009582f
C5328 vdd.n3481 gnd 0.009582f
C5329 vdd.n3482 gnd 0.009582f
C5330 vdd.n3483 gnd 0.007712f
C5331 vdd.n3484 gnd 0.009582f
C5332 vdd.n3485 gnd 0.768708f
C5333 vdd.n3486 gnd 0.009582f
C5334 vdd.n3487 gnd 0.009582f
C5335 vdd.n3488 gnd 0.007712f
C5336 vdd.n3489 gnd 0.007712f
C5337 vdd.n3490 gnd 0.007712f
C5338 vdd.n3491 gnd 0.009582f
C5339 vdd.n3492 gnd 0.009582f
C5340 vdd.n3493 gnd 0.009582f
C5341 vdd.n3494 gnd 0.009582f
C5342 vdd.n3495 gnd 0.007712f
C5343 vdd.n3496 gnd 0.007712f
C5344 vdd.n3497 gnd 0.007712f
C5345 vdd.n3498 gnd 0.009582f
C5346 vdd.n3499 gnd 0.009582f
C5347 vdd.n3500 gnd 0.009582f
C5348 vdd.n3501 gnd 0.009582f
C5349 vdd.n3502 gnd 0.007712f
C5350 vdd.n3503 gnd 0.007712f
C5351 vdd.n3504 gnd 0.007712f
C5352 vdd.n3505 gnd 0.009582f
C5353 vdd.n3506 gnd 0.009582f
C5354 vdd.n3507 gnd 0.009582f
C5355 vdd.n3508 gnd 0.812775f
C5356 vdd.n3509 gnd 0.009582f
C5357 vdd.n3510 gnd 0.007712f
C5358 vdd.n3511 gnd 0.007712f
C5359 vdd.n3512 gnd 0.007712f
C5360 vdd.n3513 gnd 0.009582f
C5361 vdd.n3514 gnd 0.009582f
C5362 vdd.n3515 gnd 0.009582f
C5363 vdd.n3516 gnd 0.009582f
C5364 vdd.n3517 gnd 0.007712f
C5365 vdd.n3518 gnd 0.007712f
C5366 vdd.n3519 gnd 0.006401f
C5367 vdd.n3520 gnd 0.021821f
C5368 vdd.n3521 gnd 0.02197f
C5369 vdd.n3522 gnd 0.003663f
C5370 vdd.n3523 gnd 0.02197f
C5371 vdd.n3525 gnd 2.16413f
C5372 vdd.n3526 gnd 1.29261f
C5373 vdd.n3527 gnd 0.641406f
C5374 vdd.n3528 gnd 0.009582f
C5375 vdd.n3529 gnd 0.007712f
C5376 vdd.n3530 gnd 0.007712f
C5377 vdd.n3531 gnd 0.007712f
C5378 vdd.n3532 gnd 0.009582f
C5379 vdd.n3533 gnd 0.979246f
C5380 vdd.n3534 gnd 0.979246f
C5381 vdd.n3535 gnd 0.563067f
C5382 vdd.n3536 gnd 0.009582f
C5383 vdd.n3537 gnd 0.007712f
C5384 vdd.n3538 gnd 0.007712f
C5385 vdd.n3539 gnd 0.007712f
C5386 vdd.n3540 gnd 0.009582f
C5387 vdd.n3541 gnd 0.582652f
C5388 vdd.n3542 gnd 0.719746f
C5389 vdd.t114 gnd 0.489623f
C5390 vdd.n3543 gnd 0.749124f
C5391 vdd.n3544 gnd 0.009582f
C5392 vdd.n3545 gnd 0.007712f
C5393 vdd.n3546 gnd 0.007712f
C5394 vdd.n3547 gnd 0.007712f
C5395 vdd.n3548 gnd 0.009582f
C5396 vdd.n3549 gnd 0.812775f
C5397 vdd.t68 gnd 0.489623f
C5398 vdd.n3550 gnd 0.592444f
C5399 vdd.n3551 gnd 0.709954f
C5400 vdd.n3552 gnd 0.009582f
C5401 vdd.n3553 gnd 0.007712f
C5402 vdd.n3554 gnd 0.007712f
C5403 vdd.n3555 gnd 0.007712f
C5404 vdd.n3556 gnd 0.009582f
C5405 vdd.n3557 gnd 0.543482f
C5406 vdd.t102 gnd 0.489623f
C5407 vdd.n3558 gnd 0.812775f
C5408 vdd.t60 gnd 0.489623f
C5409 vdd.n3559 gnd 0.602237f
C5410 vdd.n3560 gnd 0.009582f
C5411 vdd.n3561 gnd 0.007712f
C5412 vdd.n3562 gnd 0.007364f
C5413 vdd.n3563 gnd 0.565189f
C5414 vdd.n3564 gnd 2.62939f
C5415 a_n2982_13878.n0 gnd 3.88594f
C5416 a_n2982_13878.n1 gnd 2.85743f
C5417 a_n2982_13878.n2 gnd 3.82475f
C5418 a_n2982_13878.n3 gnd 0.806598f
C5419 a_n2982_13878.n4 gnd 0.8066f
C5420 a_n2982_13878.n5 gnd 0.916876f
C5421 a_n2982_13878.n6 gnd 0.201555f
C5422 a_n2982_13878.n7 gnd 0.148449f
C5423 a_n2982_13878.n8 gnd 0.233314f
C5424 a_n2982_13878.n9 gnd 0.180209f
C5425 a_n2982_13878.n10 gnd 0.201555f
C5426 a_n2982_13878.n11 gnd 0.148449f
C5427 a_n2982_13878.n12 gnd 0.969982f
C5428 a_n2982_13878.n13 gnd 0.212423f
C5429 a_n2982_13878.n14 gnd 0.747657f
C5430 a_n2982_13878.n15 gnd 0.212423f
C5431 a_n2982_13878.n16 gnd 0.212423f
C5432 a_n2982_13878.n17 gnd 0.483791f
C5433 a_n2982_13878.n18 gnd 0.278519f
C5434 a_n2982_13878.n19 gnd 0.212423f
C5435 a_n2982_13878.n20 gnd 0.536897f
C5436 a_n2982_13878.n21 gnd 0.212423f
C5437 a_n2982_13878.n22 gnd 0.212423f
C5438 a_n2982_13878.n23 gnd 0.945129f
C5439 a_n2982_13878.n24 gnd 0.278519f
C5440 a_n2982_13878.n25 gnd 0.106212f
C5441 a_n2982_13878.n26 gnd 0.212423f
C5442 a_n2982_13878.n27 gnd 0.85592f
C5443 a_n2982_13878.n28 gnd 0.212423f
C5444 a_n2982_13878.n29 gnd 0.278519f
C5445 a_n2982_13878.n30 gnd 0.985615f
C5446 a_n2982_13878.n31 gnd 0.212423f
C5447 a_n2982_13878.n32 gnd 0.212423f
C5448 a_n2982_13878.n33 gnd 0.483791f
C5449 a_n2982_13878.n34 gnd 0.212423f
C5450 a_n2982_13878.n35 gnd 0.278519f
C5451 a_n2982_13878.n36 gnd 3.26746f
C5452 a_n2982_13878.n37 gnd 0.278518f
C5453 a_n2982_13878.n38 gnd 1.17841f
C5454 a_n2982_13878.n39 gnd 2.1518f
C5455 a_n2982_13878.n40 gnd 1.74886f
C5456 a_n2982_13878.n41 gnd 1.74886f
C5457 a_n2982_13878.n42 gnd 1.17841f
C5458 a_n2982_13878.n43 gnd 2.35355f
C5459 a_n2982_13878.n44 gnd 0.008523f
C5460 a_n2982_13878.n45 gnd 4.11e-19
C5461 a_n2982_13878.n47 gnd 0.008224f
C5462 a_n2982_13878.n48 gnd 0.011959f
C5463 a_n2982_13878.n49 gnd 0.007912f
C5464 a_n2982_13878.n51 gnd 1.6691f
C5465 a_n2982_13878.n52 gnd 0.28176f
C5466 a_n2982_13878.n53 gnd 0.008523f
C5467 a_n2982_13878.n54 gnd 4.11e-19
C5468 a_n2982_13878.n56 gnd 0.008224f
C5469 a_n2982_13878.n57 gnd 0.011959f
C5470 a_n2982_13878.n58 gnd 0.004385f
C5471 a_n2982_13878.n59 gnd 0.008523f
C5472 a_n2982_13878.n60 gnd 4.11e-19
C5473 a_n2982_13878.n62 gnd 0.008224f
C5474 a_n2982_13878.n63 gnd 0.011959f
C5475 a_n2982_13878.n64 gnd 0.007912f
C5476 a_n2982_13878.n66 gnd 0.28176f
C5477 a_n2982_13878.n67 gnd 0.008523f
C5478 a_n2982_13878.n68 gnd 4.11e-19
C5479 a_n2982_13878.n70 gnd 0.008224f
C5480 a_n2982_13878.n71 gnd 0.011959f
C5481 a_n2982_13878.n72 gnd 0.007912f
C5482 a_n2982_13878.n74 gnd 0.28176f
C5483 a_n2982_13878.n75 gnd 0.008224f
C5484 a_n2982_13878.n76 gnd 0.280611f
C5485 a_n2982_13878.n77 gnd 0.008224f
C5486 a_n2982_13878.n78 gnd 0.280611f
C5487 a_n2982_13878.n79 gnd 0.008224f
C5488 a_n2982_13878.n80 gnd 0.280611f
C5489 a_n2982_13878.n81 gnd 0.008224f
C5490 a_n2982_13878.n82 gnd 0.280611f
C5491 a_n2982_13878.n83 gnd 0.301308f
C5492 a_n2982_13878.t28 gnd 1.37961f
C5493 a_n2982_13878.t30 gnd 0.147339f
C5494 a_n2982_13878.t50 gnd 0.147339f
C5495 a_n2982_13878.n84 gnd 1.03786f
C5496 a_n2982_13878.t38 gnd 0.147339f
C5497 a_n2982_13878.t8 gnd 0.147339f
C5498 a_n2982_13878.n85 gnd 1.03786f
C5499 a_n2982_13878.t16 gnd 0.147339f
C5500 a_n2982_13878.t26 gnd 0.147339f
C5501 a_n2982_13878.n86 gnd 1.03786f
C5502 a_n2982_13878.t20 gnd 0.147339f
C5503 a_n2982_13878.t40 gnd 0.147339f
C5504 a_n2982_13878.n87 gnd 1.03786f
C5505 a_n2982_13878.t32 gnd 0.147339f
C5506 a_n2982_13878.t52 gnd 0.147339f
C5507 a_n2982_13878.n88 gnd 1.03786f
C5508 a_n2982_13878.t31 gnd 0.68535f
C5509 a_n2982_13878.n89 gnd 0.301308f
C5510 a_n2982_13878.t51 gnd 0.68535f
C5511 a_n2982_13878.t19 gnd 0.68535f
C5512 a_n2982_13878.n90 gnd 0.292258f
C5513 a_n2982_13878.t7 gnd 0.68535f
C5514 a_n2982_13878.n91 gnd 0.303898f
C5515 a_n2982_13878.t15 gnd 0.68535f
C5516 a_n2982_13878.t49 gnd 0.68535f
C5517 a_n2982_13878.n92 gnd 0.297169f
C5518 a_n2982_13878.t27 gnd 0.699618f
C5519 a_n2982_13878.t86 gnd 0.68535f
C5520 a_n2982_13878.n93 gnd 0.301308f
C5521 a_n2982_13878.t96 gnd 0.68535f
C5522 a_n2982_13878.t101 gnd 0.68535f
C5523 a_n2982_13878.n94 gnd 0.292258f
C5524 a_n2982_13878.t105 gnd 0.68535f
C5525 a_n2982_13878.n95 gnd 0.303898f
C5526 a_n2982_13878.t76 gnd 0.68535f
C5527 a_n2982_13878.t79 gnd 0.68535f
C5528 a_n2982_13878.n96 gnd 0.297169f
C5529 a_n2982_13878.t109 gnd 0.699618f
C5530 a_n2982_13878.t41 gnd 0.699618f
C5531 a_n2982_13878.t47 gnd 0.68535f
C5532 a_n2982_13878.t11 gnd 0.68535f
C5533 a_n2982_13878.t9 gnd 0.68535f
C5534 a_n2982_13878.n97 gnd 0.301188f
C5535 a_n2982_13878.t23 gnd 0.68535f
C5536 a_n2982_13878.t13 gnd 0.68535f
C5537 a_n2982_13878.t35 gnd 0.68535f
C5538 a_n2982_13878.n98 gnd 0.297497f
C5539 a_n2982_13878.t45 gnd 0.68535f
C5540 a_n2982_13878.t17 gnd 0.68535f
C5541 a_n2982_13878.t43 gnd 0.68535f
C5542 a_n2982_13878.t33 gnd 0.68535f
C5543 a_n2982_13878.t21 gnd 0.699618f
C5544 a_n2982_13878.t110 gnd 0.699618f
C5545 a_n2982_13878.t87 gnd 0.68535f
C5546 a_n2982_13878.t92 gnd 0.68535f
C5547 a_n2982_13878.t80 gnd 0.68535f
C5548 a_n2982_13878.n99 gnd 0.301188f
C5549 a_n2982_13878.t97 gnd 0.68535f
C5550 a_n2982_13878.t106 gnd 0.68535f
C5551 a_n2982_13878.t107 gnd 0.68535f
C5552 a_n2982_13878.n100 gnd 0.297497f
C5553 a_n2982_13878.t74 gnd 0.68535f
C5554 a_n2982_13878.t89 gnd 0.68535f
C5555 a_n2982_13878.t77 gnd 0.68535f
C5556 a_n2982_13878.n101 gnd 0.301308f
C5557 a_n2982_13878.t84 gnd 0.68535f
C5558 a_n2982_13878.t103 gnd 0.696376f
C5559 a_n2982_13878.n102 gnd 0.303454f
C5560 a_n2982_13878.n103 gnd 0.297752f
C5561 a_n2982_13878.n104 gnd 0.292258f
C5562 a_n2982_13878.n105 gnd 0.301323f
C5563 a_n2982_13878.n106 gnd 0.303898f
C5564 a_n2982_13878.n107 gnd 0.297169f
C5565 a_n2982_13878.n108 gnd 0.303453f
C5566 a_n2982_13878.n109 gnd 0.303454f
C5567 a_n2982_13878.t64 gnd 0.114597f
C5568 a_n2982_13878.t68 gnd 0.114597f
C5569 a_n2982_13878.n110 gnd 1.01487f
C5570 a_n2982_13878.t69 gnd 0.114597f
C5571 a_n2982_13878.t71 gnd 0.114597f
C5572 a_n2982_13878.n111 gnd 1.01262f
C5573 a_n2982_13878.t3 gnd 0.114597f
C5574 a_n2982_13878.t56 gnd 0.114597f
C5575 a_n2982_13878.n112 gnd 1.01262f
C5576 a_n2982_13878.t57 gnd 0.114597f
C5577 a_n2982_13878.t67 gnd 0.114597f
C5578 a_n2982_13878.n113 gnd 1.01487f
C5579 a_n2982_13878.t65 gnd 0.114597f
C5580 a_n2982_13878.t1 gnd 0.114597f
C5581 a_n2982_13878.n114 gnd 1.01262f
C5582 a_n2982_13878.t59 gnd 0.114597f
C5583 a_n2982_13878.t54 gnd 0.114597f
C5584 a_n2982_13878.n115 gnd 1.01262f
C5585 a_n2982_13878.t0 gnd 0.114597f
C5586 a_n2982_13878.t63 gnd 0.114597f
C5587 a_n2982_13878.n116 gnd 1.01262f
C5588 a_n2982_13878.t53 gnd 0.114597f
C5589 a_n2982_13878.t4 gnd 0.114597f
C5590 a_n2982_13878.n117 gnd 1.01262f
C5591 a_n2982_13878.t62 gnd 0.114597f
C5592 a_n2982_13878.t58 gnd 0.114597f
C5593 a_n2982_13878.n118 gnd 1.01262f
C5594 a_n2982_13878.t2 gnd 0.114597f
C5595 a_n2982_13878.t66 gnd 0.114597f
C5596 a_n2982_13878.n119 gnd 1.01487f
C5597 a_n2982_13878.t70 gnd 0.114597f
C5598 a_n2982_13878.t60 gnd 0.114597f
C5599 a_n2982_13878.n120 gnd 1.01262f
C5600 a_n2982_13878.t55 gnd 0.114597f
C5601 a_n2982_13878.t61 gnd 0.114597f
C5602 a_n2982_13878.n121 gnd 1.01262f
C5603 a_n2982_13878.n122 gnd 0.30128f
C5604 a_n2982_13878.n123 gnd 0.292258f
C5605 a_n2982_13878.n124 gnd 0.301323f
C5606 a_n2982_13878.n125 gnd 0.303898f
C5607 a_n2982_13878.n126 gnd 0.297169f
C5608 a_n2982_13878.n127 gnd 0.303453f
C5609 a_n2982_13878.t22 gnd 1.37961f
C5610 a_n2982_13878.t44 gnd 0.147339f
C5611 a_n2982_13878.t34 gnd 0.147339f
C5612 a_n2982_13878.n128 gnd 1.03786f
C5613 a_n2982_13878.t46 gnd 0.147339f
C5614 a_n2982_13878.t18 gnd 0.147339f
C5615 a_n2982_13878.n129 gnd 1.03786f
C5616 a_n2982_13878.t14 gnd 0.147339f
C5617 a_n2982_13878.t36 gnd 0.147339f
C5618 a_n2982_13878.n130 gnd 1.03786f
C5619 a_n2982_13878.t10 gnd 0.147339f
C5620 a_n2982_13878.t24 gnd 0.147339f
C5621 a_n2982_13878.n131 gnd 1.03786f
C5622 a_n2982_13878.t48 gnd 0.147339f
C5623 a_n2982_13878.t12 gnd 0.147339f
C5624 a_n2982_13878.n132 gnd 1.03786f
C5625 a_n2982_13878.t42 gnd 1.37686f
C5626 a_n2982_13878.n133 gnd 1.00893f
C5627 a_n2982_13878.t85 gnd 0.68535f
C5628 a_n2982_13878.t95 gnd 0.68535f
C5629 a_n2982_13878.t111 gnd 0.68535f
C5630 a_n2982_13878.n134 gnd 0.301323f
C5631 a_n2982_13878.t98 gnd 0.68535f
C5632 a_n2982_13878.t81 gnd 0.68535f
C5633 a_n2982_13878.t82 gnd 0.68535f
C5634 a_n2982_13878.n135 gnd 0.301323f
C5635 a_n2982_13878.t102 gnd 0.68535f
C5636 a_n2982_13878.t91 gnd 0.68535f
C5637 a_n2982_13878.t90 gnd 0.68535f
C5638 a_n2982_13878.n136 gnd 0.301323f
C5639 a_n2982_13878.t94 gnd 0.68535f
C5640 a_n2982_13878.t83 gnd 0.68535f
C5641 a_n2982_13878.t72 gnd 0.68535f
C5642 a_n2982_13878.n137 gnd 0.301323f
C5643 a_n2982_13878.t99 gnd 0.696834f
C5644 a_n2982_13878.n138 gnd 0.297497f
C5645 a_n2982_13878.n139 gnd 0.292094f
C5646 a_n2982_13878.t108 gnd 0.696834f
C5647 a_n2982_13878.n140 gnd 0.297497f
C5648 a_n2982_13878.n141 gnd 0.292094f
C5649 a_n2982_13878.t93 gnd 0.696834f
C5650 a_n2982_13878.n142 gnd 0.297497f
C5651 a_n2982_13878.n143 gnd 0.292094f
C5652 a_n2982_13878.t88 gnd 0.696834f
C5653 a_n2982_13878.n144 gnd 0.297497f
C5654 a_n2982_13878.n145 gnd 0.292094f
C5655 a_n2982_13878.n146 gnd 1.34265f
C5656 a_n2982_13878.t78 gnd 0.68535f
C5657 a_n2982_13878.n147 gnd 0.303453f
C5658 a_n2982_13878.t104 gnd 0.68535f
C5659 a_n2982_13878.n148 gnd 0.301188f
C5660 a_n2982_13878.n149 gnd 0.301323f
C5661 a_n2982_13878.t100 gnd 0.68535f
C5662 a_n2982_13878.n150 gnd 0.297497f
C5663 a_n2982_13878.t73 gnd 0.68535f
C5664 a_n2982_13878.n151 gnd 0.297752f
C5665 a_n2982_13878.n152 gnd 0.303454f
C5666 a_n2982_13878.t75 gnd 0.696376f
C5667 a_n2982_13878.t29 gnd 0.68535f
C5668 a_n2982_13878.n153 gnd 0.303453f
C5669 a_n2982_13878.t37 gnd 0.68535f
C5670 a_n2982_13878.n154 gnd 0.301188f
C5671 a_n2982_13878.n155 gnd 0.301323f
C5672 a_n2982_13878.t25 gnd 0.68535f
C5673 a_n2982_13878.n156 gnd 0.297497f
C5674 a_n2982_13878.t39 gnd 0.68535f
C5675 a_n2982_13878.n157 gnd 0.297752f
C5676 a_n2982_13878.n158 gnd 0.303454f
C5677 a_n2982_13878.t5 gnd 0.696376f
C5678 a_n2982_13878.n159 gnd 1.32692f
C5679 a_n2982_13878.t6 gnd 1.37686f
C5680 a_n8964_8799.t36 gnd 0.114243f
C5681 a_n8964_8799.t26 gnd 0.114243f
C5682 a_n8964_8799.t25 gnd 0.114243f
C5683 a_n8964_8799.n0 gnd 1.01173f
C5684 a_n8964_8799.t31 gnd 0.114243f
C5685 a_n8964_8799.t30 gnd 0.114243f
C5686 a_n8964_8799.n1 gnd 1.00949f
C5687 a_n8964_8799.n2 gnd 0.804105f
C5688 a_n8964_8799.t5 gnd 0.146883f
C5689 a_n8964_8799.t44 gnd 0.146883f
C5690 a_n8964_8799.n3 gnd 1.15849f
C5691 a_n8964_8799.t4 gnd 0.146883f
C5692 a_n8964_8799.t46 gnd 0.146883f
C5693 a_n8964_8799.n4 gnd 1.15658f
C5694 a_n8964_8799.n5 gnd 1.03963f
C5695 a_n8964_8799.t2 gnd 0.146883f
C5696 a_n8964_8799.t13 gnd 0.146883f
C5697 a_n8964_8799.n6 gnd 1.15658f
C5698 a_n8964_8799.n7 gnd 0.51245f
C5699 a_n8964_8799.t1 gnd 0.146883f
C5700 a_n8964_8799.t14 gnd 0.146883f
C5701 a_n8964_8799.n8 gnd 1.15658f
C5702 a_n8964_8799.n9 gnd 0.51245f
C5703 a_n8964_8799.t43 gnd 0.146883f
C5704 a_n8964_8799.t15 gnd 0.146883f
C5705 a_n8964_8799.n10 gnd 1.15658f
C5706 a_n8964_8799.n11 gnd 0.51245f
C5707 a_n8964_8799.t45 gnd 0.146883f
C5708 a_n8964_8799.t0 gnd 0.146883f
C5709 a_n8964_8799.n12 gnd 1.15658f
C5710 a_n8964_8799.n13 gnd 3.78338f
C5711 a_n8964_8799.t7 gnd 0.146883f
C5712 a_n8964_8799.t8 gnd 0.146883f
C5713 a_n8964_8799.n14 gnd 1.15849f
C5714 a_n8964_8799.t10 gnd 0.146883f
C5715 a_n8964_8799.t47 gnd 0.146883f
C5716 a_n8964_8799.n15 gnd 1.15658f
C5717 a_n8964_8799.n16 gnd 1.03962f
C5718 a_n8964_8799.t17 gnd 0.146883f
C5719 a_n8964_8799.t3 gnd 0.146883f
C5720 a_n8964_8799.n17 gnd 1.15658f
C5721 a_n8964_8799.n18 gnd 0.51245f
C5722 a_n8964_8799.t6 gnd 0.146883f
C5723 a_n8964_8799.t18 gnd 0.146883f
C5724 a_n8964_8799.n19 gnd 1.15658f
C5725 a_n8964_8799.n20 gnd 0.51245f
C5726 a_n8964_8799.t16 gnd 0.146883f
C5727 a_n8964_8799.t9 gnd 0.146883f
C5728 a_n8964_8799.n21 gnd 1.15658f
C5729 a_n8964_8799.n22 gnd 0.51245f
C5730 a_n8964_8799.t12 gnd 0.146883f
C5731 a_n8964_8799.t11 gnd 0.146883f
C5732 a_n8964_8799.n23 gnd 1.15658f
C5733 a_n8964_8799.n24 gnd 2.52923f
C5734 a_n8964_8799.n25 gnd 7.77025f
C5735 a_n8964_8799.n26 gnd 0.052942f
C5736 a_n8964_8799.t85 gnd 0.609047f
C5737 a_n8964_8799.n27 gnd 0.272012f
C5738 a_n8964_8799.n28 gnd 0.052942f
C5739 a_n8964_8799.n29 gnd 0.012014f
C5740 a_n8964_8799.t114 gnd 0.609047f
C5741 a_n8964_8799.n30 gnd 0.052942f
C5742 a_n8964_8799.t130 gnd 0.609047f
C5743 a_n8964_8799.n31 gnd 0.271849f
C5744 a_n8964_8799.t131 gnd 0.609047f
C5745 a_n8964_8799.n32 gnd 0.052942f
C5746 a_n8964_8799.n33 gnd 0.012014f
C5747 a_n8964_8799.t73 gnd 0.609047f
C5748 a_n8964_8799.n34 gnd 0.052942f
C5749 a_n8964_8799.t74 gnd 0.609047f
C5750 a_n8964_8799.n35 gnd 0.266953f
C5751 a_n8964_8799.t107 gnd 0.609047f
C5752 a_n8964_8799.n36 gnd 0.052942f
C5753 a_n8964_8799.t111 gnd 0.609047f
C5754 a_n8964_8799.n37 gnd 0.271196f
C5755 a_n8964_8799.t86 gnd 0.620574f
C5756 a_n8964_8799.n38 gnd 0.255339f
C5757 a_n8964_8799.n39 gnd 0.173109f
C5758 a_n8964_8799.n40 gnd 0.012014f
C5759 a_n8964_8799.t50 gnd 0.609047f
C5760 a_n8964_8799.n41 gnd 0.272012f
C5761 a_n8964_8799.n42 gnd 0.012014f
C5762 a_n8964_8799.n43 gnd 0.052942f
C5763 a_n8964_8799.n44 gnd 0.052942f
C5764 a_n8964_8799.n45 gnd 0.052942f
C5765 a_n8964_8799.n46 gnd 0.271522f
C5766 a_n8964_8799.n47 gnd 0.012014f
C5767 a_n8964_8799.t134 gnd 0.609047f
C5768 a_n8964_8799.n48 gnd 0.272012f
C5769 a_n8964_8799.n49 gnd 0.052942f
C5770 a_n8964_8799.n50 gnd 0.052942f
C5771 a_n8964_8799.n51 gnd 0.052942f
C5772 a_n8964_8799.n52 gnd 0.266626f
C5773 a_n8964_8799.t103 gnd 0.609047f
C5774 a_n8964_8799.n53 gnd 0.271849f
C5775 a_n8964_8799.n54 gnd 0.012014f
C5776 a_n8964_8799.n55 gnd 0.052942f
C5777 a_n8964_8799.n56 gnd 0.052942f
C5778 a_n8964_8799.n57 gnd 0.052942f
C5779 a_n8964_8799.n58 gnd 0.266626f
C5780 a_n8964_8799.n59 gnd 0.012014f
C5781 a_n8964_8799.t88 gnd 0.609047f
C5782 a_n8964_8799.n60 gnd 0.272012f
C5783 a_n8964_8799.n61 gnd 0.052942f
C5784 a_n8964_8799.n62 gnd 0.052942f
C5785 a_n8964_8799.n63 gnd 0.052942f
C5786 a_n8964_8799.n64 gnd 0.271522f
C5787 a_n8964_8799.t129 gnd 0.609047f
C5788 a_n8964_8799.n65 gnd 0.266953f
C5789 a_n8964_8799.n66 gnd 0.012014f
C5790 a_n8964_8799.n67 gnd 0.052942f
C5791 a_n8964_8799.n68 gnd 0.052942f
C5792 a_n8964_8799.n69 gnd 0.052942f
C5793 a_n8964_8799.n70 gnd 0.012014f
C5794 a_n8964_8799.t87 gnd 0.609047f
C5795 a_n8964_8799.n71 gnd 0.271196f
C5796 a_n8964_8799.t112 gnd 0.609047f
C5797 a_n8964_8799.n72 gnd 0.266463f
C5798 a_n8964_8799.n73 gnd 0.305039f
C5799 a_n8964_8799.n74 gnd 0.052942f
C5800 a_n8964_8799.t94 gnd 0.609047f
C5801 a_n8964_8799.n75 gnd 0.272012f
C5802 a_n8964_8799.n76 gnd 0.052942f
C5803 a_n8964_8799.n77 gnd 0.012014f
C5804 a_n8964_8799.t126 gnd 0.609047f
C5805 a_n8964_8799.n78 gnd 0.052942f
C5806 a_n8964_8799.t140 gnd 0.609047f
C5807 a_n8964_8799.n79 gnd 0.271849f
C5808 a_n8964_8799.t142 gnd 0.609047f
C5809 a_n8964_8799.n80 gnd 0.052942f
C5810 a_n8964_8799.n81 gnd 0.012014f
C5811 a_n8964_8799.t80 gnd 0.609047f
C5812 a_n8964_8799.n82 gnd 0.052942f
C5813 a_n8964_8799.t83 gnd 0.609047f
C5814 a_n8964_8799.n83 gnd 0.266953f
C5815 a_n8964_8799.t116 gnd 0.609047f
C5816 a_n8964_8799.n84 gnd 0.052942f
C5817 a_n8964_8799.t122 gnd 0.609047f
C5818 a_n8964_8799.n85 gnd 0.271196f
C5819 a_n8964_8799.t95 gnd 0.620574f
C5820 a_n8964_8799.n86 gnd 0.255339f
C5821 a_n8964_8799.n87 gnd 0.173109f
C5822 a_n8964_8799.n88 gnd 0.012014f
C5823 a_n8964_8799.t60 gnd 0.609047f
C5824 a_n8964_8799.n89 gnd 0.272012f
C5825 a_n8964_8799.n90 gnd 0.012014f
C5826 a_n8964_8799.n91 gnd 0.052942f
C5827 a_n8964_8799.n92 gnd 0.052942f
C5828 a_n8964_8799.n93 gnd 0.052942f
C5829 a_n8964_8799.n94 gnd 0.271522f
C5830 a_n8964_8799.n95 gnd 0.012014f
C5831 a_n8964_8799.t143 gnd 0.609047f
C5832 a_n8964_8799.n96 gnd 0.272012f
C5833 a_n8964_8799.n97 gnd 0.052942f
C5834 a_n8964_8799.n98 gnd 0.052942f
C5835 a_n8964_8799.n99 gnd 0.052942f
C5836 a_n8964_8799.n100 gnd 0.266626f
C5837 a_n8964_8799.t113 gnd 0.609047f
C5838 a_n8964_8799.n101 gnd 0.271849f
C5839 a_n8964_8799.n102 gnd 0.012014f
C5840 a_n8964_8799.n103 gnd 0.052942f
C5841 a_n8964_8799.n104 gnd 0.052942f
C5842 a_n8964_8799.n105 gnd 0.052942f
C5843 a_n8964_8799.n106 gnd 0.266626f
C5844 a_n8964_8799.n107 gnd 0.012014f
C5845 a_n8964_8799.t99 gnd 0.609047f
C5846 a_n8964_8799.n108 gnd 0.272012f
C5847 a_n8964_8799.n109 gnd 0.052942f
C5848 a_n8964_8799.n110 gnd 0.052942f
C5849 a_n8964_8799.n111 gnd 0.052942f
C5850 a_n8964_8799.n112 gnd 0.271522f
C5851 a_n8964_8799.t139 gnd 0.609047f
C5852 a_n8964_8799.n113 gnd 0.266953f
C5853 a_n8964_8799.n114 gnd 0.012014f
C5854 a_n8964_8799.n115 gnd 0.052942f
C5855 a_n8964_8799.n116 gnd 0.052942f
C5856 a_n8964_8799.n117 gnd 0.052942f
C5857 a_n8964_8799.n118 gnd 0.012014f
C5858 a_n8964_8799.t96 gnd 0.609047f
C5859 a_n8964_8799.n119 gnd 0.271196f
C5860 a_n8964_8799.t123 gnd 0.609047f
C5861 a_n8964_8799.n120 gnd 0.266463f
C5862 a_n8964_8799.n121 gnd 0.137159f
C5863 a_n8964_8799.n122 gnd 0.917292f
C5864 a_n8964_8799.n123 gnd 0.052942f
C5865 a_n8964_8799.t66 gnd 0.609047f
C5866 a_n8964_8799.n124 gnd 0.272012f
C5867 a_n8964_8799.n125 gnd 0.052942f
C5868 a_n8964_8799.n126 gnd 0.012014f
C5869 a_n8964_8799.t81 gnd 0.609047f
C5870 a_n8964_8799.n127 gnd 0.052942f
C5871 a_n8964_8799.t109 gnd 0.609047f
C5872 a_n8964_8799.n128 gnd 0.271849f
C5873 a_n8964_8799.t93 gnd 0.609047f
C5874 a_n8964_8799.n129 gnd 0.052942f
C5875 a_n8964_8799.n130 gnd 0.012014f
C5876 a_n8964_8799.t97 gnd 0.609047f
C5877 a_n8964_8799.n131 gnd 0.052942f
C5878 a_n8964_8799.t64 gnd 0.609047f
C5879 a_n8964_8799.n132 gnd 0.266953f
C5880 a_n8964_8799.t118 gnd 0.609047f
C5881 a_n8964_8799.n133 gnd 0.052942f
C5882 a_n8964_8799.t51 gnd 0.609047f
C5883 a_n8964_8799.n134 gnd 0.271196f
C5884 a_n8964_8799.t89 gnd 0.620574f
C5885 a_n8964_8799.n135 gnd 0.255339f
C5886 a_n8964_8799.n136 gnd 0.173109f
C5887 a_n8964_8799.n137 gnd 0.012014f
C5888 a_n8964_8799.t104 gnd 0.609047f
C5889 a_n8964_8799.n138 gnd 0.272012f
C5890 a_n8964_8799.n139 gnd 0.012014f
C5891 a_n8964_8799.n140 gnd 0.052942f
C5892 a_n8964_8799.n141 gnd 0.052942f
C5893 a_n8964_8799.n142 gnd 0.052942f
C5894 a_n8964_8799.n143 gnd 0.271522f
C5895 a_n8964_8799.n144 gnd 0.012014f
C5896 a_n8964_8799.t76 gnd 0.609047f
C5897 a_n8964_8799.n145 gnd 0.272012f
C5898 a_n8964_8799.n146 gnd 0.052942f
C5899 a_n8964_8799.n147 gnd 0.052942f
C5900 a_n8964_8799.n148 gnd 0.052942f
C5901 a_n8964_8799.n149 gnd 0.266626f
C5902 a_n8964_8799.t58 gnd 0.609047f
C5903 a_n8964_8799.n150 gnd 0.271849f
C5904 a_n8964_8799.n151 gnd 0.012014f
C5905 a_n8964_8799.n152 gnd 0.052942f
C5906 a_n8964_8799.n153 gnd 0.052942f
C5907 a_n8964_8799.n154 gnd 0.052942f
C5908 a_n8964_8799.n155 gnd 0.266626f
C5909 a_n8964_8799.n156 gnd 0.012014f
C5910 a_n8964_8799.t125 gnd 0.609047f
C5911 a_n8964_8799.n157 gnd 0.272012f
C5912 a_n8964_8799.n158 gnd 0.052942f
C5913 a_n8964_8799.n159 gnd 0.052942f
C5914 a_n8964_8799.n160 gnd 0.052942f
C5915 a_n8964_8799.n161 gnd 0.271522f
C5916 a_n8964_8799.t132 gnd 0.609047f
C5917 a_n8964_8799.n162 gnd 0.266953f
C5918 a_n8964_8799.n163 gnd 0.012014f
C5919 a_n8964_8799.n164 gnd 0.052942f
C5920 a_n8964_8799.n165 gnd 0.052942f
C5921 a_n8964_8799.n166 gnd 0.052942f
C5922 a_n8964_8799.n167 gnd 0.012014f
C5923 a_n8964_8799.t48 gnd 0.609047f
C5924 a_n8964_8799.n168 gnd 0.271196f
C5925 a_n8964_8799.t100 gnd 0.609047f
C5926 a_n8964_8799.n169 gnd 0.266463f
C5927 a_n8964_8799.n170 gnd 0.137159f
C5928 a_n8964_8799.n171 gnd 1.93567f
C5929 a_n8964_8799.n172 gnd 0.052942f
C5930 a_n8964_8799.t55 gnd 0.609047f
C5931 a_n8964_8799.t53 gnd 0.609047f
C5932 a_n8964_8799.t121 gnd 0.609047f
C5933 a_n8964_8799.n173 gnd 0.272012f
C5934 a_n8964_8799.n174 gnd 0.052942f
C5935 a_n8964_8799.t69 gnd 0.609047f
C5936 a_n8964_8799.t57 gnd 0.609047f
C5937 a_n8964_8799.n175 gnd 0.052942f
C5938 a_n8964_8799.t127 gnd 0.609047f
C5939 a_n8964_8799.n176 gnd 0.272012f
C5940 a_n8964_8799.n177 gnd 0.052942f
C5941 a_n8964_8799.t90 gnd 0.609047f
C5942 a_n8964_8799.t70 gnd 0.609047f
C5943 a_n8964_8799.n178 gnd 0.052942f
C5944 a_n8964_8799.t141 gnd 0.609047f
C5945 a_n8964_8799.n179 gnd 0.271849f
C5946 a_n8964_8799.n180 gnd 0.052942f
C5947 a_n8964_8799.t106 gnd 0.609047f
C5948 a_n8964_8799.t72 gnd 0.609047f
C5949 a_n8964_8799.n181 gnd 0.052942f
C5950 a_n8964_8799.t137 gnd 0.609047f
C5951 a_n8964_8799.n182 gnd 0.271522f
C5952 a_n8964_8799.n183 gnd 0.052942f
C5953 a_n8964_8799.t108 gnd 0.609047f
C5954 a_n8964_8799.t84 gnd 0.609047f
C5955 a_n8964_8799.n184 gnd 0.052942f
C5956 a_n8964_8799.t54 gnd 0.609047f
C5957 a_n8964_8799.n185 gnd 0.271196f
C5958 a_n8964_8799.t124 gnd 0.620574f
C5959 a_n8964_8799.n186 gnd 0.255339f
C5960 a_n8964_8799.n187 gnd 0.17311f
C5961 a_n8964_8799.n188 gnd 0.012014f
C5962 a_n8964_8799.n189 gnd 0.272012f
C5963 a_n8964_8799.n190 gnd 0.012014f
C5964 a_n8964_8799.n191 gnd 0.266953f
C5965 a_n8964_8799.n192 gnd 0.052942f
C5966 a_n8964_8799.n193 gnd 0.052942f
C5967 a_n8964_8799.n194 gnd 0.052942f
C5968 a_n8964_8799.n195 gnd 0.012014f
C5969 a_n8964_8799.n196 gnd 0.272012f
C5970 a_n8964_8799.n197 gnd 0.012014f
C5971 a_n8964_8799.n198 gnd 0.266626f
C5972 a_n8964_8799.n199 gnd 0.052942f
C5973 a_n8964_8799.n200 gnd 0.052942f
C5974 a_n8964_8799.n201 gnd 0.052942f
C5975 a_n8964_8799.n202 gnd 0.012014f
C5976 a_n8964_8799.n203 gnd 0.271849f
C5977 a_n8964_8799.n204 gnd 0.266626f
C5978 a_n8964_8799.n205 gnd 0.012014f
C5979 a_n8964_8799.n206 gnd 0.052942f
C5980 a_n8964_8799.n207 gnd 0.052942f
C5981 a_n8964_8799.n208 gnd 0.052942f
C5982 a_n8964_8799.n209 gnd 0.012014f
C5983 a_n8964_8799.n210 gnd 0.271522f
C5984 a_n8964_8799.n211 gnd 0.266953f
C5985 a_n8964_8799.n212 gnd 0.012014f
C5986 a_n8964_8799.n213 gnd 0.052942f
C5987 a_n8964_8799.n214 gnd 0.052942f
C5988 a_n8964_8799.n215 gnd 0.052942f
C5989 a_n8964_8799.n216 gnd 0.012014f
C5990 a_n8964_8799.n217 gnd 0.271196f
C5991 a_n8964_8799.n218 gnd 0.266463f
C5992 a_n8964_8799.n219 gnd 0.305039f
C5993 a_n8964_8799.n220 gnd 0.052942f
C5994 a_n8964_8799.t62 gnd 0.609047f
C5995 a_n8964_8799.t61 gnd 0.609047f
C5996 a_n8964_8799.t135 gnd 0.609047f
C5997 a_n8964_8799.n221 gnd 0.272012f
C5998 a_n8964_8799.n222 gnd 0.052942f
C5999 a_n8964_8799.t75 gnd 0.609047f
C6000 a_n8964_8799.t68 gnd 0.609047f
C6001 a_n8964_8799.n223 gnd 0.052942f
C6002 a_n8964_8799.t138 gnd 0.609047f
C6003 a_n8964_8799.n224 gnd 0.272012f
C6004 a_n8964_8799.n225 gnd 0.052942f
C6005 a_n8964_8799.t102 gnd 0.609047f
C6006 a_n8964_8799.t78 gnd 0.609047f
C6007 a_n8964_8799.n226 gnd 0.052942f
C6008 a_n8964_8799.t56 gnd 0.609047f
C6009 a_n8964_8799.n227 gnd 0.271849f
C6010 a_n8964_8799.n228 gnd 0.052942f
C6011 a_n8964_8799.t115 gnd 0.609047f
C6012 a_n8964_8799.t79 gnd 0.609047f
C6013 a_n8964_8799.n229 gnd 0.052942f
C6014 a_n8964_8799.t49 gnd 0.609047f
C6015 a_n8964_8799.n230 gnd 0.271522f
C6016 a_n8964_8799.n231 gnd 0.052942f
C6017 a_n8964_8799.t120 gnd 0.609047f
C6018 a_n8964_8799.t92 gnd 0.609047f
C6019 a_n8964_8799.n232 gnd 0.052942f
C6020 a_n8964_8799.t63 gnd 0.609047f
C6021 a_n8964_8799.n233 gnd 0.271196f
C6022 a_n8964_8799.t136 gnd 0.620574f
C6023 a_n8964_8799.n234 gnd 0.255339f
C6024 a_n8964_8799.n235 gnd 0.17311f
C6025 a_n8964_8799.n236 gnd 0.012014f
C6026 a_n8964_8799.n237 gnd 0.272012f
C6027 a_n8964_8799.n238 gnd 0.012014f
C6028 a_n8964_8799.n239 gnd 0.266953f
C6029 a_n8964_8799.n240 gnd 0.052942f
C6030 a_n8964_8799.n241 gnd 0.052942f
C6031 a_n8964_8799.n242 gnd 0.052942f
C6032 a_n8964_8799.n243 gnd 0.012014f
C6033 a_n8964_8799.n244 gnd 0.272012f
C6034 a_n8964_8799.n245 gnd 0.012014f
C6035 a_n8964_8799.n246 gnd 0.266626f
C6036 a_n8964_8799.n247 gnd 0.052942f
C6037 a_n8964_8799.n248 gnd 0.052942f
C6038 a_n8964_8799.n249 gnd 0.052942f
C6039 a_n8964_8799.n250 gnd 0.012014f
C6040 a_n8964_8799.n251 gnd 0.271849f
C6041 a_n8964_8799.n252 gnd 0.266626f
C6042 a_n8964_8799.n253 gnd 0.012014f
C6043 a_n8964_8799.n254 gnd 0.052942f
C6044 a_n8964_8799.n255 gnd 0.052942f
C6045 a_n8964_8799.n256 gnd 0.052942f
C6046 a_n8964_8799.n257 gnd 0.012014f
C6047 a_n8964_8799.n258 gnd 0.271522f
C6048 a_n8964_8799.n259 gnd 0.266953f
C6049 a_n8964_8799.n260 gnd 0.012014f
C6050 a_n8964_8799.n261 gnd 0.052942f
C6051 a_n8964_8799.n262 gnd 0.052942f
C6052 a_n8964_8799.n263 gnd 0.052942f
C6053 a_n8964_8799.n264 gnd 0.012014f
C6054 a_n8964_8799.n265 gnd 0.271196f
C6055 a_n8964_8799.n266 gnd 0.266463f
C6056 a_n8964_8799.n267 gnd 0.137159f
C6057 a_n8964_8799.n268 gnd 0.917292f
C6058 a_n8964_8799.n269 gnd 0.052942f
C6059 a_n8964_8799.t101 gnd 0.609047f
C6060 a_n8964_8799.t119 gnd 0.609047f
C6061 a_n8964_8799.t67 gnd 0.609047f
C6062 a_n8964_8799.n270 gnd 0.272012f
C6063 a_n8964_8799.n271 gnd 0.052942f
C6064 a_n8964_8799.t133 gnd 0.609047f
C6065 a_n8964_8799.t82 gnd 0.609047f
C6066 a_n8964_8799.n272 gnd 0.052942f
C6067 a_n8964_8799.t128 gnd 0.609047f
C6068 a_n8964_8799.n273 gnd 0.272012f
C6069 a_n8964_8799.n274 gnd 0.052942f
C6070 a_n8964_8799.t71 gnd 0.609047f
C6071 a_n8964_8799.t110 gnd 0.609047f
C6072 a_n8964_8799.n275 gnd 0.052942f
C6073 a_n8964_8799.t59 gnd 0.609047f
C6074 a_n8964_8799.n276 gnd 0.271849f
C6075 a_n8964_8799.n277 gnd 0.052942f
C6076 a_n8964_8799.t98 gnd 0.609047f
C6077 a_n8964_8799.t77 gnd 0.609047f
C6078 a_n8964_8799.n278 gnd 0.052942f
C6079 a_n8964_8799.t117 gnd 0.609047f
C6080 a_n8964_8799.n279 gnd 0.271522f
C6081 a_n8964_8799.n280 gnd 0.052942f
C6082 a_n8964_8799.t65 gnd 0.609047f
C6083 a_n8964_8799.t105 gnd 0.609047f
C6084 a_n8964_8799.n281 gnd 0.052942f
C6085 a_n8964_8799.t52 gnd 0.609047f
C6086 a_n8964_8799.n282 gnd 0.271196f
C6087 a_n8964_8799.t91 gnd 0.620574f
C6088 a_n8964_8799.n283 gnd 0.255339f
C6089 a_n8964_8799.n284 gnd 0.17311f
C6090 a_n8964_8799.n285 gnd 0.012014f
C6091 a_n8964_8799.n286 gnd 0.272012f
C6092 a_n8964_8799.n287 gnd 0.012014f
C6093 a_n8964_8799.n288 gnd 0.266953f
C6094 a_n8964_8799.n289 gnd 0.052942f
C6095 a_n8964_8799.n290 gnd 0.052942f
C6096 a_n8964_8799.n291 gnd 0.052942f
C6097 a_n8964_8799.n292 gnd 0.012014f
C6098 a_n8964_8799.n293 gnd 0.272012f
C6099 a_n8964_8799.n294 gnd 0.012014f
C6100 a_n8964_8799.n295 gnd 0.266626f
C6101 a_n8964_8799.n296 gnd 0.052942f
C6102 a_n8964_8799.n297 gnd 0.052942f
C6103 a_n8964_8799.n298 gnd 0.052942f
C6104 a_n8964_8799.n299 gnd 0.012014f
C6105 a_n8964_8799.n300 gnd 0.271849f
C6106 a_n8964_8799.n301 gnd 0.266626f
C6107 a_n8964_8799.n302 gnd 0.012014f
C6108 a_n8964_8799.n303 gnd 0.052942f
C6109 a_n8964_8799.n304 gnd 0.052942f
C6110 a_n8964_8799.n305 gnd 0.052942f
C6111 a_n8964_8799.n306 gnd 0.012014f
C6112 a_n8964_8799.n307 gnd 0.271522f
C6113 a_n8964_8799.n308 gnd 0.266953f
C6114 a_n8964_8799.n309 gnd 0.012014f
C6115 a_n8964_8799.n310 gnd 0.052942f
C6116 a_n8964_8799.n311 gnd 0.052942f
C6117 a_n8964_8799.n312 gnd 0.052942f
C6118 a_n8964_8799.n313 gnd 0.012014f
C6119 a_n8964_8799.n314 gnd 0.271196f
C6120 a_n8964_8799.n315 gnd 0.266463f
C6121 a_n8964_8799.n316 gnd 0.137159f
C6122 a_n8964_8799.n317 gnd 1.40346f
C6123 a_n8964_8799.n318 gnd 17.687399f
C6124 a_n8964_8799.n319 gnd 4.45734f
C6125 a_n8964_8799.t27 gnd 0.114243f
C6126 a_n8964_8799.t28 gnd 0.114243f
C6127 a_n8964_8799.n320 gnd 1.01173f
C6128 a_n8964_8799.t21 gnd 0.114243f
C6129 a_n8964_8799.t22 gnd 0.114243f
C6130 a_n8964_8799.n321 gnd 1.00949f
C6131 a_n8964_8799.n322 gnd 0.804103f
C6132 a_n8964_8799.t20 gnd 0.114243f
C6133 a_n8964_8799.t38 gnd 0.114243f
C6134 a_n8964_8799.n323 gnd 1.00949f
C6135 a_n8964_8799.n324 gnd 0.335766f
C6136 a_n8964_8799.n325 gnd 0.479366f
C6137 a_n8964_8799.t40 gnd 0.114243f
C6138 a_n8964_8799.t33 gnd 0.114243f
C6139 a_n8964_8799.n326 gnd 1.00949f
C6140 a_n8964_8799.n327 gnd 0.335766f
C6141 a_n8964_8799.t35 gnd 0.114243f
C6142 a_n8964_8799.t19 gnd 0.114243f
C6143 a_n8964_8799.n328 gnd 1.00949f
C6144 a_n8964_8799.n329 gnd 0.394856f
C6145 a_n8964_8799.t37 gnd 0.114243f
C6146 a_n8964_8799.t39 gnd 0.114243f
C6147 a_n8964_8799.n330 gnd 1.00949f
C6148 a_n8964_8799.n331 gnd 2.90698f
C6149 a_n8964_8799.t34 gnd 0.114243f
C6150 a_n8964_8799.t32 gnd 0.114243f
C6151 a_n8964_8799.n332 gnd 1.01173f
C6152 a_n8964_8799.t23 gnd 0.114243f
C6153 a_n8964_8799.t29 gnd 0.114243f
C6154 a_n8964_8799.n333 gnd 1.00949f
C6155 a_n8964_8799.n334 gnd 0.804105f
C6156 a_n8964_8799.t41 gnd 0.114243f
C6157 a_n8964_8799.t24 gnd 0.114243f
C6158 a_n8964_8799.n335 gnd 1.00949f
C6159 a_n8964_8799.n336 gnd 0.335767f
C6160 a_n8964_8799.n337 gnd 2.44664f
C6161 a_n8964_8799.n338 gnd 0.33577f
C6162 a_n8964_8799.n339 gnd 1.00948f
C6163 a_n8964_8799.t42 gnd 0.114243f
C6164 a_n3827_n3924.n0 gnd 1.99733f
C6165 a_n3827_n3924.n1 gnd 2.17486f
C6166 a_n3827_n3924.n2 gnd 1.44807f
C6167 a_n3827_n3924.n3 gnd 1.31657f
C6168 a_n3827_n3924.n4 gnd 1.81285f
C6169 a_n3827_n3924.n5 gnd 0.914318f
C6170 a_n3827_n3924.n6 gnd 3.90473f
C6171 a_n3827_n3924.n7 gnd 0.886511f
C6172 a_n3827_n3924.n8 gnd 1.77302f
C6173 a_n3827_n3924.n9 gnd 2.49022f
C6174 a_n3827_n3924.n10 gnd 0.954549f
C6175 a_n3827_n3924.n11 gnd 0.724032f
C6176 a_n3827_n3924.n12 gnd 1.2733f
C6177 a_n3827_n3924.t6 gnd 1.26048f
C6178 a_n3827_n3924.t0 gnd 1.25868f
C6179 a_n3827_n3924.t13 gnd 1.25868f
C6180 a_n3827_n3924.t57 gnd 1.25868f
C6181 a_n3827_n3924.t49 gnd 1.25868f
C6182 a_n3827_n3924.t50 gnd 1.25868f
C6183 a_n3827_n3924.t7 gnd 1.25868f
C6184 a_n3827_n3924.t56 gnd 1.25868f
C6185 a_n3827_n3924.t8 gnd 1.25868f
C6186 a_n3827_n3924.t14 gnd 1.26084f
C6187 a_n3827_n3924.t26 gnd 1.01304f
C6188 a_n3827_n3924.t34 gnd 0.097472f
C6189 a_n3827_n3924.t47 gnd 0.097472f
C6190 a_n3827_n3924.n13 gnd 0.796068f
C6191 a_n3827_n3924.t36 gnd 0.097472f
C6192 a_n3827_n3924.t35 gnd 0.097472f
C6193 a_n3827_n3924.n14 gnd 0.796068f
C6194 a_n3827_n3924.t31 gnd 0.097472f
C6195 a_n3827_n3924.t43 gnd 0.097472f
C6196 a_n3827_n3924.n15 gnd 0.796068f
C6197 a_n3827_n3924.t28 gnd 0.097472f
C6198 a_n3827_n3924.t30 gnd 0.097472f
C6199 a_n3827_n3924.n16 gnd 0.796068f
C6200 a_n3827_n3924.t27 gnd 0.097472f
C6201 a_n3827_n3924.t48 gnd 0.097472f
C6202 a_n3827_n3924.n17 gnd 0.796068f
C6203 a_n3827_n3924.t29 gnd 1.01304f
C6204 a_n3827_n3924.t22 gnd 1.01304f
C6205 a_n3827_n3924.t52 gnd 0.097472f
C6206 a_n3827_n3924.t53 gnd 0.097472f
C6207 a_n3827_n3924.n18 gnd 0.796068f
C6208 a_n3827_n3924.t55 gnd 0.097472f
C6209 a_n3827_n3924.t4 gnd 0.097472f
C6210 a_n3827_n3924.n19 gnd 0.796068f
C6211 a_n3827_n3924.t12 gnd 0.097472f
C6212 a_n3827_n3924.t17 gnd 0.097472f
C6213 a_n3827_n3924.n20 gnd 0.796068f
C6214 a_n3827_n3924.t10 gnd 0.097472f
C6215 a_n3827_n3924.t23 gnd 0.097472f
C6216 a_n3827_n3924.n21 gnd 0.796068f
C6217 a_n3827_n3924.t2 gnd 0.097472f
C6218 a_n3827_n3924.t15 gnd 0.097472f
C6219 a_n3827_n3924.n22 gnd 0.796068f
C6220 a_n3827_n3924.t51 gnd 1.01304f
C6221 a_n3827_n3924.n23 gnd 0.914318f
C6222 a_n3827_n3924.t45 gnd 1.01304f
C6223 a_n3827_n3924.t32 gnd 0.097472f
C6224 a_n3827_n3924.t33 gnd 0.097472f
C6225 a_n3827_n3924.n24 gnd 0.796069f
C6226 a_n3827_n3924.t38 gnd 0.097472f
C6227 a_n3827_n3924.t37 gnd 0.097472f
C6228 a_n3827_n3924.n25 gnd 0.796069f
C6229 a_n3827_n3924.t41 gnd 0.097472f
C6230 a_n3827_n3924.t42 gnd 0.097472f
C6231 a_n3827_n3924.n26 gnd 0.796069f
C6232 a_n3827_n3924.t40 gnd 0.097472f
C6233 a_n3827_n3924.t44 gnd 0.097472f
C6234 a_n3827_n3924.n27 gnd 0.796069f
C6235 a_n3827_n3924.t46 gnd 0.097472f
C6236 a_n3827_n3924.t39 gnd 0.097472f
C6237 a_n3827_n3924.n28 gnd 0.796069f
C6238 a_n3827_n3924.t25 gnd 1.01304f
C6239 a_n3827_n3924.t24 gnd 1.01304f
C6240 a_n3827_n3924.t18 gnd 0.097472f
C6241 a_n3827_n3924.t3 gnd 0.097472f
C6242 a_n3827_n3924.n29 gnd 0.796069f
C6243 a_n3827_n3924.t19 gnd 0.097472f
C6244 a_n3827_n3924.t54 gnd 0.097472f
C6245 a_n3827_n3924.n30 gnd 0.796069f
C6246 a_n3827_n3924.t16 gnd 0.097472f
C6247 a_n3827_n3924.t11 gnd 0.097472f
C6248 a_n3827_n3924.n31 gnd 0.796069f
C6249 a_n3827_n3924.t5 gnd 0.097472f
C6250 a_n3827_n3924.t20 gnd 0.097472f
C6251 a_n3827_n3924.n32 gnd 0.796069f
C6252 a_n3827_n3924.t21 gnd 0.097472f
C6253 a_n3827_n3924.t9 gnd 0.097472f
C6254 a_n3827_n3924.n33 gnd 0.796069f
C6255 a_n3827_n3924.t1 gnd 1.01304f
C6256 plus.n0 gnd 0.023479f
C6257 plus.t21 gnd 0.332087f
C6258 plus.n1 gnd 0.023479f
C6259 plus.t22 gnd 0.332087f
C6260 plus.t16 gnd 0.332087f
C6261 plus.n2 gnd 0.147524f
C6262 plus.n3 gnd 0.023479f
C6263 plus.t17 gnd 0.332087f
C6264 plus.t11 gnd 0.332087f
C6265 plus.n4 gnd 0.147524f
C6266 plus.n5 gnd 0.023479f
C6267 plus.t5 gnd 0.332087f
C6268 plus.t6 gnd 0.332087f
C6269 plus.n6 gnd 0.147524f
C6270 plus.n7 gnd 0.023479f
C6271 plus.t23 gnd 0.332087f
C6272 plus.t24 gnd 0.332087f
C6273 plus.n8 gnd 0.147524f
C6274 plus.n9 gnd 0.023479f
C6275 plus.t18 gnd 0.332087f
C6276 plus.t13 gnd 0.332087f
C6277 plus.n10 gnd 0.152328f
C6278 plus.t15 gnd 0.344141f
C6279 plus.n11 gnd 0.136719f
C6280 plus.n12 gnd 0.101078f
C6281 plus.n13 gnd 0.005328f
C6282 plus.n14 gnd 0.147524f
C6283 plus.n15 gnd 0.005328f
C6284 plus.n16 gnd 0.023479f
C6285 plus.n17 gnd 0.023479f
C6286 plus.n18 gnd 0.023479f
C6287 plus.n19 gnd 0.005328f
C6288 plus.n20 gnd 0.147524f
C6289 plus.n21 gnd 0.005328f
C6290 plus.n22 gnd 0.023479f
C6291 plus.n23 gnd 0.023479f
C6292 plus.n24 gnd 0.023479f
C6293 plus.n25 gnd 0.005328f
C6294 plus.n26 gnd 0.147524f
C6295 plus.n27 gnd 0.005328f
C6296 plus.n28 gnd 0.023479f
C6297 plus.n29 gnd 0.023479f
C6298 plus.n30 gnd 0.023479f
C6299 plus.n31 gnd 0.005328f
C6300 plus.n32 gnd 0.147524f
C6301 plus.n33 gnd 0.005328f
C6302 plus.n34 gnd 0.023479f
C6303 plus.n35 gnd 0.023479f
C6304 plus.n36 gnd 0.023479f
C6305 plus.n37 gnd 0.005328f
C6306 plus.n38 gnd 0.147524f
C6307 plus.n39 gnd 0.005328f
C6308 plus.n40 gnd 0.147741f
C6309 plus.n41 gnd 0.265862f
C6310 plus.n42 gnd 0.023479f
C6311 plus.n43 gnd 0.005328f
C6312 plus.t10 gnd 0.332087f
C6313 plus.n44 gnd 0.023479f
C6314 plus.n45 gnd 0.005328f
C6315 plus.t12 gnd 0.332087f
C6316 plus.n46 gnd 0.023479f
C6317 plus.n47 gnd 0.005328f
C6318 plus.t7 gnd 0.332087f
C6319 plus.n48 gnd 0.023479f
C6320 plus.n49 gnd 0.005328f
C6321 plus.t27 gnd 0.332087f
C6322 plus.n50 gnd 0.023479f
C6323 plus.n51 gnd 0.005328f
C6324 plus.t26 gnd 0.332087f
C6325 plus.t20 gnd 0.344141f
C6326 plus.t19 gnd 0.332087f
C6327 plus.n52 gnd 0.152328f
C6328 plus.n53 gnd 0.136719f
C6329 plus.n54 gnd 0.101078f
C6330 plus.n55 gnd 0.023479f
C6331 plus.n56 gnd 0.147524f
C6332 plus.n57 gnd 0.005328f
C6333 plus.t25 gnd 0.332087f
C6334 plus.n58 gnd 0.147524f
C6335 plus.n59 gnd 0.023479f
C6336 plus.n60 gnd 0.023479f
C6337 plus.n61 gnd 0.023479f
C6338 plus.n62 gnd 0.147524f
C6339 plus.n63 gnd 0.005328f
C6340 plus.t9 gnd 0.332087f
C6341 plus.n64 gnd 0.147524f
C6342 plus.n65 gnd 0.023479f
C6343 plus.n66 gnd 0.023479f
C6344 plus.n67 gnd 0.023479f
C6345 plus.n68 gnd 0.147524f
C6346 plus.n69 gnd 0.005328f
C6347 plus.t14 gnd 0.332087f
C6348 plus.n70 gnd 0.147524f
C6349 plus.n71 gnd 0.023479f
C6350 plus.n72 gnd 0.023479f
C6351 plus.n73 gnd 0.023479f
C6352 plus.n74 gnd 0.147524f
C6353 plus.n75 gnd 0.005328f
C6354 plus.t28 gnd 0.332087f
C6355 plus.n76 gnd 0.147524f
C6356 plus.n77 gnd 0.023479f
C6357 plus.n78 gnd 0.023479f
C6358 plus.n79 gnd 0.023479f
C6359 plus.n80 gnd 0.147524f
C6360 plus.n81 gnd 0.005328f
C6361 plus.t8 gnd 0.332087f
C6362 plus.n82 gnd 0.147741f
C6363 plus.n83 gnd 0.777153f
C6364 plus.n84 gnd 1.16267f
C6365 plus.t2 gnd 0.040531f
C6366 plus.t3 gnd 0.007238f
C6367 plus.t1 gnd 0.007238f
C6368 plus.n85 gnd 0.023474f
C6369 plus.n86 gnd 0.182228f
C6370 plus.t4 gnd 0.007238f
C6371 plus.t0 gnd 0.007238f
C6372 plus.n87 gnd 0.023474f
C6373 plus.n88 gnd 0.136784f
C6374 plus.n89 gnd 2.9595f
.ends

