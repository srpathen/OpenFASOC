* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right.t15 minus.t0 source.t18 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X1 source.t2 plus.t0 drain_left.t15 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X2 drain_right.t14 minus.t1 source.t23 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X3 source.t29 minus.t2 drain_right.t13 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X4 source.t19 minus.t3 drain_right.t12 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X5 source.t9 plus.t1 drain_left.t14 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X6 a_n2210_n2088# a_n2210_n2088# a_n2210_n2088# a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.5
X7 source.t27 minus.t4 drain_right.t11 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X8 drain_right.t10 minus.t5 source.t25 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X9 drain_right.t9 minus.t6 source.t22 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X10 a_n2210_n2088# a_n2210_n2088# a_n2210_n2088# a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X11 drain_right.t8 minus.t7 source.t24 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X12 drain_left.t13 plus.t2 source.t6 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X13 source.t7 plus.t3 drain_left.t12 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X14 source.t26 minus.t8 drain_right.t7 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X15 source.t15 minus.t9 drain_right.t6 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X16 drain_left.t11 plus.t4 source.t10 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X17 source.t5 plus.t5 drain_left.t10 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X18 a_n2210_n2088# a_n2210_n2088# a_n2210_n2088# a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X19 source.t14 plus.t6 drain_left.t9 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X20 drain_right.t5 minus.t10 source.t17 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X21 source.t31 plus.t7 drain_left.t8 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X22 drain_left.t7 plus.t8 source.t3 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X23 a_n2210_n2088# a_n2210_n2088# a_n2210_n2088# a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.5
X24 drain_left.t6 plus.t9 source.t11 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X25 drain_right.t4 minus.t11 source.t20 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X26 source.t21 minus.t12 drain_right.t3 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.5
X27 source.t16 minus.t13 drain_right.t2 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X28 source.t4 plus.t10 drain_left.t5 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X29 source.t28 minus.t14 drain_right.t1 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X30 drain_left.t4 plus.t11 source.t8 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X31 drain_left.t3 plus.t12 source.t12 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
X32 source.t0 plus.t13 drain_left.t2 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X33 drain_left.t1 plus.t14 source.t13 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X34 drain_left.t0 plus.t15 source.t1 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.5
X35 drain_right.t0 minus.t15 source.t30 a_n2210_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.5
R0 minus.n5 minus.t10 388.748
R1 minus.n27 minus.t12 388.748
R2 minus.n6 minus.t3 367.767
R3 minus.n8 minus.t7 367.767
R4 minus.n12 minus.t13 367.767
R5 minus.n13 minus.t6 367.767
R6 minus.n1 minus.t8 367.767
R7 minus.n19 minus.t0 367.767
R8 minus.n20 minus.t9 367.767
R9 minus.n28 minus.t11 367.767
R10 minus.n30 minus.t2 367.767
R11 minus.n34 minus.t1 367.767
R12 minus.n35 minus.t14 367.767
R13 minus.n23 minus.t5 367.767
R14 minus.n41 minus.t4 367.767
R15 minus.n42 minus.t15 367.767
R16 minus.n21 minus.n20 161.3
R17 minus.n19 minus.n0 161.3
R18 minus.n18 minus.n17 161.3
R19 minus.n16 minus.n1 161.3
R20 minus.n15 minus.n14 161.3
R21 minus.n13 minus.n2 161.3
R22 minus.n12 minus.n11 161.3
R23 minus.n10 minus.n3 161.3
R24 minus.n9 minus.n8 161.3
R25 minus.n7 minus.n4 161.3
R26 minus.n43 minus.n42 161.3
R27 minus.n41 minus.n22 161.3
R28 minus.n40 minus.n39 161.3
R29 minus.n38 minus.n23 161.3
R30 minus.n37 minus.n36 161.3
R31 minus.n35 minus.n24 161.3
R32 minus.n34 minus.n33 161.3
R33 minus.n32 minus.n25 161.3
R34 minus.n31 minus.n30 161.3
R35 minus.n29 minus.n26 161.3
R36 minus.n5 minus.n4 70.4033
R37 minus.n27 minus.n26 70.4033
R38 minus.n13 minus.n12 48.2005
R39 minus.n20 minus.n19 48.2005
R40 minus.n35 minus.n34 48.2005
R41 minus.n42 minus.n41 48.2005
R42 minus.n8 minus.n7 37.246
R43 minus.n18 minus.n1 37.246
R44 minus.n30 minus.n29 37.246
R45 minus.n40 minus.n23 37.246
R46 minus.n8 minus.n3 35.7853
R47 minus.n14 minus.n1 35.7853
R48 minus.n30 minus.n25 35.7853
R49 minus.n36 minus.n23 35.7853
R50 minus.n44 minus.n21 33.0081
R51 minus.n6 minus.n5 20.9576
R52 minus.n28 minus.n27 20.9576
R53 minus.n12 minus.n3 12.4157
R54 minus.n14 minus.n13 12.4157
R55 minus.n34 minus.n25 12.4157
R56 minus.n36 minus.n35 12.4157
R57 minus.n7 minus.n6 10.955
R58 minus.n19 minus.n18 10.955
R59 minus.n29 minus.n28 10.955
R60 minus.n41 minus.n40 10.955
R61 minus.n44 minus.n43 6.56111
R62 minus.n21 minus.n0 0.189894
R63 minus.n17 minus.n0 0.189894
R64 minus.n17 minus.n16 0.189894
R65 minus.n16 minus.n15 0.189894
R66 minus.n15 minus.n2 0.189894
R67 minus.n11 minus.n2 0.189894
R68 minus.n11 minus.n10 0.189894
R69 minus.n10 minus.n9 0.189894
R70 minus.n9 minus.n4 0.189894
R71 minus.n31 minus.n26 0.189894
R72 minus.n32 minus.n31 0.189894
R73 minus.n33 minus.n32 0.189894
R74 minus.n33 minus.n24 0.189894
R75 minus.n37 minus.n24 0.189894
R76 minus.n38 minus.n37 0.189894
R77 minus.n39 minus.n38 0.189894
R78 minus.n39 minus.n22 0.189894
R79 minus.n43 minus.n22 0.189894
R80 minus minus.n44 0.188
R81 source.n274 source.n248 289.615
R82 source.n236 source.n210 289.615
R83 source.n204 source.n178 289.615
R84 source.n166 source.n140 289.615
R85 source.n26 source.n0 289.615
R86 source.n64 source.n38 289.615
R87 source.n96 source.n70 289.615
R88 source.n134 source.n108 289.615
R89 source.n259 source.n258 185
R90 source.n256 source.n255 185
R91 source.n265 source.n264 185
R92 source.n267 source.n266 185
R93 source.n252 source.n251 185
R94 source.n273 source.n272 185
R95 source.n275 source.n274 185
R96 source.n221 source.n220 185
R97 source.n218 source.n217 185
R98 source.n227 source.n226 185
R99 source.n229 source.n228 185
R100 source.n214 source.n213 185
R101 source.n235 source.n234 185
R102 source.n237 source.n236 185
R103 source.n189 source.n188 185
R104 source.n186 source.n185 185
R105 source.n195 source.n194 185
R106 source.n197 source.n196 185
R107 source.n182 source.n181 185
R108 source.n203 source.n202 185
R109 source.n205 source.n204 185
R110 source.n151 source.n150 185
R111 source.n148 source.n147 185
R112 source.n157 source.n156 185
R113 source.n159 source.n158 185
R114 source.n144 source.n143 185
R115 source.n165 source.n164 185
R116 source.n167 source.n166 185
R117 source.n27 source.n26 185
R118 source.n25 source.n24 185
R119 source.n4 source.n3 185
R120 source.n19 source.n18 185
R121 source.n17 source.n16 185
R122 source.n8 source.n7 185
R123 source.n11 source.n10 185
R124 source.n65 source.n64 185
R125 source.n63 source.n62 185
R126 source.n42 source.n41 185
R127 source.n57 source.n56 185
R128 source.n55 source.n54 185
R129 source.n46 source.n45 185
R130 source.n49 source.n48 185
R131 source.n97 source.n96 185
R132 source.n95 source.n94 185
R133 source.n74 source.n73 185
R134 source.n89 source.n88 185
R135 source.n87 source.n86 185
R136 source.n78 source.n77 185
R137 source.n81 source.n80 185
R138 source.n135 source.n134 185
R139 source.n133 source.n132 185
R140 source.n112 source.n111 185
R141 source.n127 source.n126 185
R142 source.n125 source.n124 185
R143 source.n116 source.n115 185
R144 source.n119 source.n118 185
R145 source.t30 source.n257 147.661
R146 source.t21 source.n219 147.661
R147 source.t10 source.n187 147.661
R148 source.t14 source.n149 147.661
R149 source.t12 source.n9 147.661
R150 source.t9 source.n47 147.661
R151 source.t17 source.n79 147.661
R152 source.t15 source.n117 147.661
R153 source.n258 source.n255 104.615
R154 source.n265 source.n255 104.615
R155 source.n266 source.n265 104.615
R156 source.n266 source.n251 104.615
R157 source.n273 source.n251 104.615
R158 source.n274 source.n273 104.615
R159 source.n220 source.n217 104.615
R160 source.n227 source.n217 104.615
R161 source.n228 source.n227 104.615
R162 source.n228 source.n213 104.615
R163 source.n235 source.n213 104.615
R164 source.n236 source.n235 104.615
R165 source.n188 source.n185 104.615
R166 source.n195 source.n185 104.615
R167 source.n196 source.n195 104.615
R168 source.n196 source.n181 104.615
R169 source.n203 source.n181 104.615
R170 source.n204 source.n203 104.615
R171 source.n150 source.n147 104.615
R172 source.n157 source.n147 104.615
R173 source.n158 source.n157 104.615
R174 source.n158 source.n143 104.615
R175 source.n165 source.n143 104.615
R176 source.n166 source.n165 104.615
R177 source.n26 source.n25 104.615
R178 source.n25 source.n3 104.615
R179 source.n18 source.n3 104.615
R180 source.n18 source.n17 104.615
R181 source.n17 source.n7 104.615
R182 source.n10 source.n7 104.615
R183 source.n64 source.n63 104.615
R184 source.n63 source.n41 104.615
R185 source.n56 source.n41 104.615
R186 source.n56 source.n55 104.615
R187 source.n55 source.n45 104.615
R188 source.n48 source.n45 104.615
R189 source.n96 source.n95 104.615
R190 source.n95 source.n73 104.615
R191 source.n88 source.n73 104.615
R192 source.n88 source.n87 104.615
R193 source.n87 source.n77 104.615
R194 source.n80 source.n77 104.615
R195 source.n134 source.n133 104.615
R196 source.n133 source.n111 104.615
R197 source.n126 source.n111 104.615
R198 source.n126 source.n125 104.615
R199 source.n125 source.n115 104.615
R200 source.n118 source.n115 104.615
R201 source.n258 source.t30 52.3082
R202 source.n220 source.t21 52.3082
R203 source.n188 source.t10 52.3082
R204 source.n150 source.t14 52.3082
R205 source.n10 source.t12 52.3082
R206 source.n48 source.t9 52.3082
R207 source.n80 source.t17 52.3082
R208 source.n118 source.t15 52.3082
R209 source.n33 source.n32 50.512
R210 source.n35 source.n34 50.512
R211 source.n37 source.n36 50.512
R212 source.n103 source.n102 50.512
R213 source.n105 source.n104 50.512
R214 source.n107 source.n106 50.512
R215 source.n247 source.n246 50.5119
R216 source.n245 source.n244 50.5119
R217 source.n243 source.n242 50.5119
R218 source.n177 source.n176 50.5119
R219 source.n175 source.n174 50.5119
R220 source.n173 source.n172 50.5119
R221 source.n279 source.n278 32.1853
R222 source.n241 source.n240 32.1853
R223 source.n209 source.n208 32.1853
R224 source.n171 source.n170 32.1853
R225 source.n31 source.n30 32.1853
R226 source.n69 source.n68 32.1853
R227 source.n101 source.n100 32.1853
R228 source.n139 source.n138 32.1853
R229 source.n171 source.n139 17.4578
R230 source.n259 source.n257 15.6674
R231 source.n221 source.n219 15.6674
R232 source.n189 source.n187 15.6674
R233 source.n151 source.n149 15.6674
R234 source.n11 source.n9 15.6674
R235 source.n49 source.n47 15.6674
R236 source.n81 source.n79 15.6674
R237 source.n119 source.n117 15.6674
R238 source.n260 source.n256 12.8005
R239 source.n222 source.n218 12.8005
R240 source.n190 source.n186 12.8005
R241 source.n152 source.n148 12.8005
R242 source.n12 source.n8 12.8005
R243 source.n50 source.n46 12.8005
R244 source.n82 source.n78 12.8005
R245 source.n120 source.n116 12.8005
R246 source.n264 source.n263 12.0247
R247 source.n226 source.n225 12.0247
R248 source.n194 source.n193 12.0247
R249 source.n156 source.n155 12.0247
R250 source.n16 source.n15 12.0247
R251 source.n54 source.n53 12.0247
R252 source.n86 source.n85 12.0247
R253 source.n124 source.n123 12.0247
R254 source.n280 source.n31 11.8371
R255 source.n267 source.n254 11.249
R256 source.n229 source.n216 11.249
R257 source.n197 source.n184 11.249
R258 source.n159 source.n146 11.249
R259 source.n19 source.n6 11.249
R260 source.n57 source.n44 11.249
R261 source.n89 source.n76 11.249
R262 source.n127 source.n114 11.249
R263 source.n268 source.n252 10.4732
R264 source.n230 source.n214 10.4732
R265 source.n198 source.n182 10.4732
R266 source.n160 source.n144 10.4732
R267 source.n20 source.n4 10.4732
R268 source.n58 source.n42 10.4732
R269 source.n90 source.n74 10.4732
R270 source.n128 source.n112 10.4732
R271 source.n272 source.n271 9.69747
R272 source.n234 source.n233 9.69747
R273 source.n202 source.n201 9.69747
R274 source.n164 source.n163 9.69747
R275 source.n24 source.n23 9.69747
R276 source.n62 source.n61 9.69747
R277 source.n94 source.n93 9.69747
R278 source.n132 source.n131 9.69747
R279 source.n278 source.n277 9.45567
R280 source.n240 source.n239 9.45567
R281 source.n208 source.n207 9.45567
R282 source.n170 source.n169 9.45567
R283 source.n30 source.n29 9.45567
R284 source.n68 source.n67 9.45567
R285 source.n100 source.n99 9.45567
R286 source.n138 source.n137 9.45567
R287 source.n277 source.n276 9.3005
R288 source.n250 source.n249 9.3005
R289 source.n271 source.n270 9.3005
R290 source.n269 source.n268 9.3005
R291 source.n254 source.n253 9.3005
R292 source.n263 source.n262 9.3005
R293 source.n261 source.n260 9.3005
R294 source.n239 source.n238 9.3005
R295 source.n212 source.n211 9.3005
R296 source.n233 source.n232 9.3005
R297 source.n231 source.n230 9.3005
R298 source.n216 source.n215 9.3005
R299 source.n225 source.n224 9.3005
R300 source.n223 source.n222 9.3005
R301 source.n207 source.n206 9.3005
R302 source.n180 source.n179 9.3005
R303 source.n201 source.n200 9.3005
R304 source.n199 source.n198 9.3005
R305 source.n184 source.n183 9.3005
R306 source.n193 source.n192 9.3005
R307 source.n191 source.n190 9.3005
R308 source.n169 source.n168 9.3005
R309 source.n142 source.n141 9.3005
R310 source.n163 source.n162 9.3005
R311 source.n161 source.n160 9.3005
R312 source.n146 source.n145 9.3005
R313 source.n155 source.n154 9.3005
R314 source.n153 source.n152 9.3005
R315 source.n29 source.n28 9.3005
R316 source.n2 source.n1 9.3005
R317 source.n23 source.n22 9.3005
R318 source.n21 source.n20 9.3005
R319 source.n6 source.n5 9.3005
R320 source.n15 source.n14 9.3005
R321 source.n13 source.n12 9.3005
R322 source.n67 source.n66 9.3005
R323 source.n40 source.n39 9.3005
R324 source.n61 source.n60 9.3005
R325 source.n59 source.n58 9.3005
R326 source.n44 source.n43 9.3005
R327 source.n53 source.n52 9.3005
R328 source.n51 source.n50 9.3005
R329 source.n99 source.n98 9.3005
R330 source.n72 source.n71 9.3005
R331 source.n93 source.n92 9.3005
R332 source.n91 source.n90 9.3005
R333 source.n76 source.n75 9.3005
R334 source.n85 source.n84 9.3005
R335 source.n83 source.n82 9.3005
R336 source.n137 source.n136 9.3005
R337 source.n110 source.n109 9.3005
R338 source.n131 source.n130 9.3005
R339 source.n129 source.n128 9.3005
R340 source.n114 source.n113 9.3005
R341 source.n123 source.n122 9.3005
R342 source.n121 source.n120 9.3005
R343 source.n275 source.n250 8.92171
R344 source.n237 source.n212 8.92171
R345 source.n205 source.n180 8.92171
R346 source.n167 source.n142 8.92171
R347 source.n27 source.n2 8.92171
R348 source.n65 source.n40 8.92171
R349 source.n97 source.n72 8.92171
R350 source.n135 source.n110 8.92171
R351 source.n276 source.n248 8.14595
R352 source.n238 source.n210 8.14595
R353 source.n206 source.n178 8.14595
R354 source.n168 source.n140 8.14595
R355 source.n28 source.n0 8.14595
R356 source.n66 source.n38 8.14595
R357 source.n98 source.n70 8.14595
R358 source.n136 source.n108 8.14595
R359 source.n278 source.n248 5.81868
R360 source.n240 source.n210 5.81868
R361 source.n208 source.n178 5.81868
R362 source.n170 source.n140 5.81868
R363 source.n30 source.n0 5.81868
R364 source.n68 source.n38 5.81868
R365 source.n100 source.n70 5.81868
R366 source.n138 source.n108 5.81868
R367 source.n280 source.n279 5.62119
R368 source.n276 source.n275 5.04292
R369 source.n238 source.n237 5.04292
R370 source.n206 source.n205 5.04292
R371 source.n168 source.n167 5.04292
R372 source.n28 source.n27 5.04292
R373 source.n66 source.n65 5.04292
R374 source.n98 source.n97 5.04292
R375 source.n136 source.n135 5.04292
R376 source.n261 source.n257 4.38594
R377 source.n223 source.n219 4.38594
R378 source.n191 source.n187 4.38594
R379 source.n153 source.n149 4.38594
R380 source.n13 source.n9 4.38594
R381 source.n51 source.n47 4.38594
R382 source.n83 source.n79 4.38594
R383 source.n121 source.n117 4.38594
R384 source.n272 source.n250 4.26717
R385 source.n234 source.n212 4.26717
R386 source.n202 source.n180 4.26717
R387 source.n164 source.n142 4.26717
R388 source.n24 source.n2 4.26717
R389 source.n62 source.n40 4.26717
R390 source.n94 source.n72 4.26717
R391 source.n132 source.n110 4.26717
R392 source.n271 source.n252 3.49141
R393 source.n233 source.n214 3.49141
R394 source.n201 source.n182 3.49141
R395 source.n163 source.n144 3.49141
R396 source.n23 source.n4 3.49141
R397 source.n61 source.n42 3.49141
R398 source.n93 source.n74 3.49141
R399 source.n131 source.n112 3.49141
R400 source.n246 source.t25 3.3005
R401 source.n246 source.t27 3.3005
R402 source.n244 source.t23 3.3005
R403 source.n244 source.t28 3.3005
R404 source.n242 source.t20 3.3005
R405 source.n242 source.t29 3.3005
R406 source.n176 source.t13 3.3005
R407 source.n176 source.t5 3.3005
R408 source.n174 source.t3 3.3005
R409 source.n174 source.t31 3.3005
R410 source.n172 source.t8 3.3005
R411 source.n172 source.t2 3.3005
R412 source.n32 source.t1 3.3005
R413 source.n32 source.t7 3.3005
R414 source.n34 source.t6 3.3005
R415 source.n34 source.t4 3.3005
R416 source.n36 source.t11 3.3005
R417 source.n36 source.t0 3.3005
R418 source.n102 source.t24 3.3005
R419 source.n102 source.t19 3.3005
R420 source.n104 source.t22 3.3005
R421 source.n104 source.t16 3.3005
R422 source.n106 source.t18 3.3005
R423 source.n106 source.t26 3.3005
R424 source.n268 source.n267 2.71565
R425 source.n230 source.n229 2.71565
R426 source.n198 source.n197 2.71565
R427 source.n160 source.n159 2.71565
R428 source.n20 source.n19 2.71565
R429 source.n58 source.n57 2.71565
R430 source.n90 source.n89 2.71565
R431 source.n128 source.n127 2.71565
R432 source.n264 source.n254 1.93989
R433 source.n226 source.n216 1.93989
R434 source.n194 source.n184 1.93989
R435 source.n156 source.n146 1.93989
R436 source.n16 source.n6 1.93989
R437 source.n54 source.n44 1.93989
R438 source.n86 source.n76 1.93989
R439 source.n124 source.n114 1.93989
R440 source.n263 source.n256 1.16414
R441 source.n225 source.n218 1.16414
R442 source.n193 source.n186 1.16414
R443 source.n155 source.n148 1.16414
R444 source.n15 source.n8 1.16414
R445 source.n53 source.n46 1.16414
R446 source.n85 source.n78 1.16414
R447 source.n123 source.n116 1.16414
R448 source.n139 source.n107 0.716017
R449 source.n107 source.n105 0.716017
R450 source.n105 source.n103 0.716017
R451 source.n103 source.n101 0.716017
R452 source.n69 source.n37 0.716017
R453 source.n37 source.n35 0.716017
R454 source.n35 source.n33 0.716017
R455 source.n33 source.n31 0.716017
R456 source.n173 source.n171 0.716017
R457 source.n175 source.n173 0.716017
R458 source.n177 source.n175 0.716017
R459 source.n209 source.n177 0.716017
R460 source.n243 source.n241 0.716017
R461 source.n245 source.n243 0.716017
R462 source.n247 source.n245 0.716017
R463 source.n279 source.n247 0.716017
R464 source.n101 source.n69 0.470328
R465 source.n241 source.n209 0.470328
R466 source.n260 source.n259 0.388379
R467 source.n222 source.n221 0.388379
R468 source.n190 source.n189 0.388379
R469 source.n152 source.n151 0.388379
R470 source.n12 source.n11 0.388379
R471 source.n50 source.n49 0.388379
R472 source.n82 source.n81 0.388379
R473 source.n120 source.n119 0.388379
R474 source source.n280 0.188
R475 source.n262 source.n261 0.155672
R476 source.n262 source.n253 0.155672
R477 source.n269 source.n253 0.155672
R478 source.n270 source.n269 0.155672
R479 source.n270 source.n249 0.155672
R480 source.n277 source.n249 0.155672
R481 source.n224 source.n223 0.155672
R482 source.n224 source.n215 0.155672
R483 source.n231 source.n215 0.155672
R484 source.n232 source.n231 0.155672
R485 source.n232 source.n211 0.155672
R486 source.n239 source.n211 0.155672
R487 source.n192 source.n191 0.155672
R488 source.n192 source.n183 0.155672
R489 source.n199 source.n183 0.155672
R490 source.n200 source.n199 0.155672
R491 source.n200 source.n179 0.155672
R492 source.n207 source.n179 0.155672
R493 source.n154 source.n153 0.155672
R494 source.n154 source.n145 0.155672
R495 source.n161 source.n145 0.155672
R496 source.n162 source.n161 0.155672
R497 source.n162 source.n141 0.155672
R498 source.n169 source.n141 0.155672
R499 source.n29 source.n1 0.155672
R500 source.n22 source.n1 0.155672
R501 source.n22 source.n21 0.155672
R502 source.n21 source.n5 0.155672
R503 source.n14 source.n5 0.155672
R504 source.n14 source.n13 0.155672
R505 source.n67 source.n39 0.155672
R506 source.n60 source.n39 0.155672
R507 source.n60 source.n59 0.155672
R508 source.n59 source.n43 0.155672
R509 source.n52 source.n43 0.155672
R510 source.n52 source.n51 0.155672
R511 source.n99 source.n71 0.155672
R512 source.n92 source.n71 0.155672
R513 source.n92 source.n91 0.155672
R514 source.n91 source.n75 0.155672
R515 source.n84 source.n75 0.155672
R516 source.n84 source.n83 0.155672
R517 source.n137 source.n109 0.155672
R518 source.n130 source.n109 0.155672
R519 source.n130 source.n129 0.155672
R520 source.n129 source.n113 0.155672
R521 source.n122 source.n113 0.155672
R522 source.n122 source.n121 0.155672
R523 drain_right.n5 drain_right.n3 67.9062
R524 drain_right.n2 drain_right.n0 67.9062
R525 drain_right.n9 drain_right.n7 67.9062
R526 drain_right.n9 drain_right.n8 67.1908
R527 drain_right.n11 drain_right.n10 67.1908
R528 drain_right.n13 drain_right.n12 67.1908
R529 drain_right.n5 drain_right.n4 67.1907
R530 drain_right.n2 drain_right.n1 67.1907
R531 drain_right drain_right.n6 26.9193
R532 drain_right drain_right.n13 6.36873
R533 drain_right.n3 drain_right.t11 3.3005
R534 drain_right.n3 drain_right.t0 3.3005
R535 drain_right.n4 drain_right.t1 3.3005
R536 drain_right.n4 drain_right.t10 3.3005
R537 drain_right.n1 drain_right.t13 3.3005
R538 drain_right.n1 drain_right.t14 3.3005
R539 drain_right.n0 drain_right.t3 3.3005
R540 drain_right.n0 drain_right.t4 3.3005
R541 drain_right.n7 drain_right.t12 3.3005
R542 drain_right.n7 drain_right.t5 3.3005
R543 drain_right.n8 drain_right.t2 3.3005
R544 drain_right.n8 drain_right.t8 3.3005
R545 drain_right.n10 drain_right.t7 3.3005
R546 drain_right.n10 drain_right.t9 3.3005
R547 drain_right.n12 drain_right.t6 3.3005
R548 drain_right.n12 drain_right.t15 3.3005
R549 drain_right.n13 drain_right.n11 0.716017
R550 drain_right.n11 drain_right.n9 0.716017
R551 drain_right.n6 drain_right.n5 0.302913
R552 drain_right.n6 drain_right.n2 0.302913
R553 plus.n5 plus.t1 388.748
R554 plus.n27 plus.t4 388.748
R555 plus.n20 plus.t12 367.767
R556 plus.n19 plus.t3 367.767
R557 plus.n1 plus.t15 367.767
R558 plus.n13 plus.t10 367.767
R559 plus.n12 plus.t2 367.767
R560 plus.n4 plus.t13 367.767
R561 plus.n6 plus.t9 367.767
R562 plus.n42 plus.t6 367.767
R563 plus.n41 plus.t11 367.767
R564 plus.n23 plus.t0 367.767
R565 plus.n35 plus.t8 367.767
R566 plus.n34 plus.t7 367.767
R567 plus.n26 plus.t14 367.767
R568 plus.n28 plus.t5 367.767
R569 plus.n8 plus.n7 161.3
R570 plus.n9 plus.n4 161.3
R571 plus.n11 plus.n10 161.3
R572 plus.n12 plus.n3 161.3
R573 plus.n13 plus.n2 161.3
R574 plus.n15 plus.n14 161.3
R575 plus.n16 plus.n1 161.3
R576 plus.n18 plus.n17 161.3
R577 plus.n19 plus.n0 161.3
R578 plus.n21 plus.n20 161.3
R579 plus.n30 plus.n29 161.3
R580 plus.n31 plus.n26 161.3
R581 plus.n33 plus.n32 161.3
R582 plus.n34 plus.n25 161.3
R583 plus.n35 plus.n24 161.3
R584 plus.n37 plus.n36 161.3
R585 plus.n38 plus.n23 161.3
R586 plus.n40 plus.n39 161.3
R587 plus.n41 plus.n22 161.3
R588 plus.n43 plus.n42 161.3
R589 plus.n8 plus.n5 70.4033
R590 plus.n30 plus.n27 70.4033
R591 plus.n20 plus.n19 48.2005
R592 plus.n13 plus.n12 48.2005
R593 plus.n42 plus.n41 48.2005
R594 plus.n35 plus.n34 48.2005
R595 plus.n18 plus.n1 37.246
R596 plus.n7 plus.n4 37.246
R597 plus.n40 plus.n23 37.246
R598 plus.n29 plus.n26 37.246
R599 plus.n14 plus.n1 35.7853
R600 plus.n11 plus.n4 35.7853
R601 plus.n36 plus.n23 35.7853
R602 plus.n33 plus.n26 35.7853
R603 plus plus.n43 29.1619
R604 plus.n6 plus.n5 20.9576
R605 plus.n28 plus.n27 20.9576
R606 plus.n14 plus.n13 12.4157
R607 plus.n12 plus.n11 12.4157
R608 plus.n36 plus.n35 12.4157
R609 plus.n34 plus.n33 12.4157
R610 plus.n19 plus.n18 10.955
R611 plus.n7 plus.n6 10.955
R612 plus.n41 plus.n40 10.955
R613 plus.n29 plus.n28 10.955
R614 plus plus.n21 9.93232
R615 plus.n9 plus.n8 0.189894
R616 plus.n10 plus.n9 0.189894
R617 plus.n10 plus.n3 0.189894
R618 plus.n3 plus.n2 0.189894
R619 plus.n15 plus.n2 0.189894
R620 plus.n16 plus.n15 0.189894
R621 plus.n17 plus.n16 0.189894
R622 plus.n17 plus.n0 0.189894
R623 plus.n21 plus.n0 0.189894
R624 plus.n43 plus.n22 0.189894
R625 plus.n39 plus.n22 0.189894
R626 plus.n39 plus.n38 0.189894
R627 plus.n38 plus.n37 0.189894
R628 plus.n37 plus.n24 0.189894
R629 plus.n25 plus.n24 0.189894
R630 plus.n32 plus.n25 0.189894
R631 plus.n32 plus.n31 0.189894
R632 plus.n31 plus.n30 0.189894
R633 drain_left.n9 drain_left.n7 67.9063
R634 drain_left.n5 drain_left.n3 67.9062
R635 drain_left.n2 drain_left.n0 67.9062
R636 drain_left.n11 drain_left.n10 67.1908
R637 drain_left.n9 drain_left.n8 67.1908
R638 drain_left.n13 drain_left.n12 67.1907
R639 drain_left.n5 drain_left.n4 67.1907
R640 drain_left.n2 drain_left.n1 67.1907
R641 drain_left drain_left.n6 27.4725
R642 drain_left drain_left.n13 6.36873
R643 drain_left.n3 drain_left.t10 3.3005
R644 drain_left.n3 drain_left.t11 3.3005
R645 drain_left.n4 drain_left.t8 3.3005
R646 drain_left.n4 drain_left.t1 3.3005
R647 drain_left.n1 drain_left.t15 3.3005
R648 drain_left.n1 drain_left.t7 3.3005
R649 drain_left.n0 drain_left.t9 3.3005
R650 drain_left.n0 drain_left.t4 3.3005
R651 drain_left.n12 drain_left.t12 3.3005
R652 drain_left.n12 drain_left.t3 3.3005
R653 drain_left.n10 drain_left.t5 3.3005
R654 drain_left.n10 drain_left.t0 3.3005
R655 drain_left.n8 drain_left.t2 3.3005
R656 drain_left.n8 drain_left.t13 3.3005
R657 drain_left.n7 drain_left.t14 3.3005
R658 drain_left.n7 drain_left.t6 3.3005
R659 drain_left.n11 drain_left.n9 0.716017
R660 drain_left.n13 drain_left.n11 0.716017
R661 drain_left.n6 drain_left.n5 0.302913
R662 drain_left.n6 drain_left.n2 0.302913
C0 plus drain_left 4.67512f
C1 drain_left source 13.3261f
C2 drain_left minus 0.172419f
C3 plus drain_right 0.372806f
C4 drain_right source 13.327299f
C5 minus drain_right 4.45794f
C6 plus source 4.66087f
C7 plus minus 4.79552f
C8 minus source 4.64685f
C9 drain_left drain_right 1.15071f
C10 drain_right a_n2210_n2088# 5.35438f
C11 drain_left a_n2210_n2088# 5.68013f
C12 source a_n2210_n2088# 5.512761f
C13 minus a_n2210_n2088# 8.243885f
C14 plus a_n2210_n2088# 9.78162f
C15 drain_left.t9 a_n2210_n2088# 0.137841f
C16 drain_left.t4 a_n2210_n2088# 0.137841f
C17 drain_left.n0 a_n2210_n2088# 1.15362f
C18 drain_left.t15 a_n2210_n2088# 0.137841f
C19 drain_left.t7 a_n2210_n2088# 0.137841f
C20 drain_left.n1 a_n2210_n2088# 1.1496f
C21 drain_left.n2 a_n2210_n2088# 0.711242f
C22 drain_left.t10 a_n2210_n2088# 0.137841f
C23 drain_left.t11 a_n2210_n2088# 0.137841f
C24 drain_left.n3 a_n2210_n2088# 1.15362f
C25 drain_left.t8 a_n2210_n2088# 0.137841f
C26 drain_left.t1 a_n2210_n2088# 0.137841f
C27 drain_left.n4 a_n2210_n2088# 1.1496f
C28 drain_left.n5 a_n2210_n2088# 0.711242f
C29 drain_left.n6 a_n2210_n2088# 1.16666f
C30 drain_left.t14 a_n2210_n2088# 0.137841f
C31 drain_left.t6 a_n2210_n2088# 0.137841f
C32 drain_left.n7 a_n2210_n2088# 1.15362f
C33 drain_left.t2 a_n2210_n2088# 0.137841f
C34 drain_left.t13 a_n2210_n2088# 0.137841f
C35 drain_left.n8 a_n2210_n2088# 1.1496f
C36 drain_left.n9 a_n2210_n2088# 0.747701f
C37 drain_left.t5 a_n2210_n2088# 0.137841f
C38 drain_left.t0 a_n2210_n2088# 0.137841f
C39 drain_left.n10 a_n2210_n2088# 1.1496f
C40 drain_left.n11 a_n2210_n2088# 0.370007f
C41 drain_left.t12 a_n2210_n2088# 0.137841f
C42 drain_left.t3 a_n2210_n2088# 0.137841f
C43 drain_left.n12 a_n2210_n2088# 1.1496f
C44 drain_left.n13 a_n2210_n2088# 0.619781f
C45 plus.n0 a_n2210_n2088# 0.04685f
C46 plus.t12 a_n2210_n2088# 0.407676f
C47 plus.t3 a_n2210_n2088# 0.407676f
C48 plus.t15 a_n2210_n2088# 0.407676f
C49 plus.n1 a_n2210_n2088# 0.19695f
C50 plus.n2 a_n2210_n2088# 0.04685f
C51 plus.t10 a_n2210_n2088# 0.407676f
C52 plus.t2 a_n2210_n2088# 0.407676f
C53 plus.n3 a_n2210_n2088# 0.04685f
C54 plus.t13 a_n2210_n2088# 0.407676f
C55 plus.n4 a_n2210_n2088# 0.19695f
C56 plus.t1 a_n2210_n2088# 0.418044f
C57 plus.n5 a_n2210_n2088# 0.182012f
C58 plus.t9 a_n2210_n2088# 0.407676f
C59 plus.n6 a_n2210_n2088# 0.194206f
C60 plus.n7 a_n2210_n2088# 0.010631f
C61 plus.n8 a_n2210_n2088# 0.149164f
C62 plus.n9 a_n2210_n2088# 0.04685f
C63 plus.n10 a_n2210_n2088# 0.04685f
C64 plus.n11 a_n2210_n2088# 0.010631f
C65 plus.n12 a_n2210_n2088# 0.194495f
C66 plus.n13 a_n2210_n2088# 0.194495f
C67 plus.n14 a_n2210_n2088# 0.010631f
C68 plus.n15 a_n2210_n2088# 0.04685f
C69 plus.n16 a_n2210_n2088# 0.04685f
C70 plus.n17 a_n2210_n2088# 0.04685f
C71 plus.n18 a_n2210_n2088# 0.010631f
C72 plus.n19 a_n2210_n2088# 0.194206f
C73 plus.n20 a_n2210_n2088# 0.192039f
C74 plus.n21 a_n2210_n2088# 0.408478f
C75 plus.n22 a_n2210_n2088# 0.04685f
C76 plus.t6 a_n2210_n2088# 0.407676f
C77 plus.t11 a_n2210_n2088# 0.407676f
C78 plus.t0 a_n2210_n2088# 0.407676f
C79 plus.n23 a_n2210_n2088# 0.19695f
C80 plus.n24 a_n2210_n2088# 0.04685f
C81 plus.t8 a_n2210_n2088# 0.407676f
C82 plus.n25 a_n2210_n2088# 0.04685f
C83 plus.t7 a_n2210_n2088# 0.407676f
C84 plus.t14 a_n2210_n2088# 0.407676f
C85 plus.n26 a_n2210_n2088# 0.19695f
C86 plus.t4 a_n2210_n2088# 0.418044f
C87 plus.n27 a_n2210_n2088# 0.182012f
C88 plus.t5 a_n2210_n2088# 0.407676f
C89 plus.n28 a_n2210_n2088# 0.194206f
C90 plus.n29 a_n2210_n2088# 0.010631f
C91 plus.n30 a_n2210_n2088# 0.149164f
C92 plus.n31 a_n2210_n2088# 0.04685f
C93 plus.n32 a_n2210_n2088# 0.04685f
C94 plus.n33 a_n2210_n2088# 0.010631f
C95 plus.n34 a_n2210_n2088# 0.194495f
C96 plus.n35 a_n2210_n2088# 0.194495f
C97 plus.n36 a_n2210_n2088# 0.010631f
C98 plus.n37 a_n2210_n2088# 0.04685f
C99 plus.n38 a_n2210_n2088# 0.04685f
C100 plus.n39 a_n2210_n2088# 0.04685f
C101 plus.n40 a_n2210_n2088# 0.010631f
C102 plus.n41 a_n2210_n2088# 0.194206f
C103 plus.n42 a_n2210_n2088# 0.192039f
C104 plus.n43 a_n2210_n2088# 1.29442f
C105 drain_right.t3 a_n2210_n2088# 0.137176f
C106 drain_right.t4 a_n2210_n2088# 0.137176f
C107 drain_right.n0 a_n2210_n2088# 1.14805f
C108 drain_right.t13 a_n2210_n2088# 0.137176f
C109 drain_right.t14 a_n2210_n2088# 0.137176f
C110 drain_right.n1 a_n2210_n2088# 1.14405f
C111 drain_right.n2 a_n2210_n2088# 0.707812f
C112 drain_right.t11 a_n2210_n2088# 0.137176f
C113 drain_right.t0 a_n2210_n2088# 0.137176f
C114 drain_right.n3 a_n2210_n2088# 1.14805f
C115 drain_right.t1 a_n2210_n2088# 0.137176f
C116 drain_right.t10 a_n2210_n2088# 0.137176f
C117 drain_right.n4 a_n2210_n2088# 1.14405f
C118 drain_right.n5 a_n2210_n2088# 0.707812f
C119 drain_right.n6 a_n2210_n2088# 1.10265f
C120 drain_right.t12 a_n2210_n2088# 0.137176f
C121 drain_right.t5 a_n2210_n2088# 0.137176f
C122 drain_right.n7 a_n2210_n2088# 1.14805f
C123 drain_right.t2 a_n2210_n2088# 0.137176f
C124 drain_right.t8 a_n2210_n2088# 0.137176f
C125 drain_right.n8 a_n2210_n2088# 1.14406f
C126 drain_right.n9 a_n2210_n2088# 0.7441f
C127 drain_right.t7 a_n2210_n2088# 0.137176f
C128 drain_right.t9 a_n2210_n2088# 0.137176f
C129 drain_right.n10 a_n2210_n2088# 1.14406f
C130 drain_right.n11 a_n2210_n2088# 0.368222f
C131 drain_right.t6 a_n2210_n2088# 0.137176f
C132 drain_right.t15 a_n2210_n2088# 0.137176f
C133 drain_right.n12 a_n2210_n2088# 1.14406f
C134 drain_right.n13 a_n2210_n2088# 0.616786f
C135 source.n0 a_n2210_n2088# 0.03695f
C136 source.n1 a_n2210_n2088# 0.026288f
C137 source.n2 a_n2210_n2088# 0.014126f
C138 source.n3 a_n2210_n2088# 0.033388f
C139 source.n4 a_n2210_n2088# 0.014957f
C140 source.n5 a_n2210_n2088# 0.026288f
C141 source.n6 a_n2210_n2088# 0.014126f
C142 source.n7 a_n2210_n2088# 0.033388f
C143 source.n8 a_n2210_n2088# 0.014957f
C144 source.n9 a_n2210_n2088# 0.112492f
C145 source.t12 a_n2210_n2088# 0.054418f
C146 source.n10 a_n2210_n2088# 0.025041f
C147 source.n11 a_n2210_n2088# 0.019722f
C148 source.n12 a_n2210_n2088# 0.014126f
C149 source.n13 a_n2210_n2088# 0.625487f
C150 source.n14 a_n2210_n2088# 0.026288f
C151 source.n15 a_n2210_n2088# 0.014126f
C152 source.n16 a_n2210_n2088# 0.014957f
C153 source.n17 a_n2210_n2088# 0.033388f
C154 source.n18 a_n2210_n2088# 0.033388f
C155 source.n19 a_n2210_n2088# 0.014957f
C156 source.n20 a_n2210_n2088# 0.014126f
C157 source.n21 a_n2210_n2088# 0.026288f
C158 source.n22 a_n2210_n2088# 0.026288f
C159 source.n23 a_n2210_n2088# 0.014126f
C160 source.n24 a_n2210_n2088# 0.014957f
C161 source.n25 a_n2210_n2088# 0.033388f
C162 source.n26 a_n2210_n2088# 0.07228f
C163 source.n27 a_n2210_n2088# 0.014957f
C164 source.n28 a_n2210_n2088# 0.014126f
C165 source.n29 a_n2210_n2088# 0.060762f
C166 source.n30 a_n2210_n2088# 0.040444f
C167 source.n31 a_n2210_n2088# 0.661753f
C168 source.t1 a_n2210_n2088# 0.124639f
C169 source.t7 a_n2210_n2088# 0.124639f
C170 source.n32 a_n2210_n2088# 0.970701f
C171 source.n33 a_n2210_n2088# 0.367635f
C172 source.t6 a_n2210_n2088# 0.124639f
C173 source.t4 a_n2210_n2088# 0.124639f
C174 source.n34 a_n2210_n2088# 0.970701f
C175 source.n35 a_n2210_n2088# 0.367635f
C176 source.t11 a_n2210_n2088# 0.124639f
C177 source.t0 a_n2210_n2088# 0.124639f
C178 source.n36 a_n2210_n2088# 0.970701f
C179 source.n37 a_n2210_n2088# 0.367635f
C180 source.n38 a_n2210_n2088# 0.03695f
C181 source.n39 a_n2210_n2088# 0.026288f
C182 source.n40 a_n2210_n2088# 0.014126f
C183 source.n41 a_n2210_n2088# 0.033388f
C184 source.n42 a_n2210_n2088# 0.014957f
C185 source.n43 a_n2210_n2088# 0.026288f
C186 source.n44 a_n2210_n2088# 0.014126f
C187 source.n45 a_n2210_n2088# 0.033388f
C188 source.n46 a_n2210_n2088# 0.014957f
C189 source.n47 a_n2210_n2088# 0.112492f
C190 source.t9 a_n2210_n2088# 0.054418f
C191 source.n48 a_n2210_n2088# 0.025041f
C192 source.n49 a_n2210_n2088# 0.019722f
C193 source.n50 a_n2210_n2088# 0.014126f
C194 source.n51 a_n2210_n2088# 0.625487f
C195 source.n52 a_n2210_n2088# 0.026288f
C196 source.n53 a_n2210_n2088# 0.014126f
C197 source.n54 a_n2210_n2088# 0.014957f
C198 source.n55 a_n2210_n2088# 0.033388f
C199 source.n56 a_n2210_n2088# 0.033388f
C200 source.n57 a_n2210_n2088# 0.014957f
C201 source.n58 a_n2210_n2088# 0.014126f
C202 source.n59 a_n2210_n2088# 0.026288f
C203 source.n60 a_n2210_n2088# 0.026288f
C204 source.n61 a_n2210_n2088# 0.014126f
C205 source.n62 a_n2210_n2088# 0.014957f
C206 source.n63 a_n2210_n2088# 0.033388f
C207 source.n64 a_n2210_n2088# 0.07228f
C208 source.n65 a_n2210_n2088# 0.014957f
C209 source.n66 a_n2210_n2088# 0.014126f
C210 source.n67 a_n2210_n2088# 0.060762f
C211 source.n68 a_n2210_n2088# 0.040444f
C212 source.n69 a_n2210_n2088# 0.122855f
C213 source.n70 a_n2210_n2088# 0.03695f
C214 source.n71 a_n2210_n2088# 0.026288f
C215 source.n72 a_n2210_n2088# 0.014126f
C216 source.n73 a_n2210_n2088# 0.033388f
C217 source.n74 a_n2210_n2088# 0.014957f
C218 source.n75 a_n2210_n2088# 0.026288f
C219 source.n76 a_n2210_n2088# 0.014126f
C220 source.n77 a_n2210_n2088# 0.033388f
C221 source.n78 a_n2210_n2088# 0.014957f
C222 source.n79 a_n2210_n2088# 0.112492f
C223 source.t17 a_n2210_n2088# 0.054418f
C224 source.n80 a_n2210_n2088# 0.025041f
C225 source.n81 a_n2210_n2088# 0.019722f
C226 source.n82 a_n2210_n2088# 0.014126f
C227 source.n83 a_n2210_n2088# 0.625487f
C228 source.n84 a_n2210_n2088# 0.026288f
C229 source.n85 a_n2210_n2088# 0.014126f
C230 source.n86 a_n2210_n2088# 0.014957f
C231 source.n87 a_n2210_n2088# 0.033388f
C232 source.n88 a_n2210_n2088# 0.033388f
C233 source.n89 a_n2210_n2088# 0.014957f
C234 source.n90 a_n2210_n2088# 0.014126f
C235 source.n91 a_n2210_n2088# 0.026288f
C236 source.n92 a_n2210_n2088# 0.026288f
C237 source.n93 a_n2210_n2088# 0.014126f
C238 source.n94 a_n2210_n2088# 0.014957f
C239 source.n95 a_n2210_n2088# 0.033388f
C240 source.n96 a_n2210_n2088# 0.07228f
C241 source.n97 a_n2210_n2088# 0.014957f
C242 source.n98 a_n2210_n2088# 0.014126f
C243 source.n99 a_n2210_n2088# 0.060762f
C244 source.n100 a_n2210_n2088# 0.040444f
C245 source.n101 a_n2210_n2088# 0.122855f
C246 source.t24 a_n2210_n2088# 0.124639f
C247 source.t19 a_n2210_n2088# 0.124639f
C248 source.n102 a_n2210_n2088# 0.970701f
C249 source.n103 a_n2210_n2088# 0.367635f
C250 source.t22 a_n2210_n2088# 0.124639f
C251 source.t16 a_n2210_n2088# 0.124639f
C252 source.n104 a_n2210_n2088# 0.970701f
C253 source.n105 a_n2210_n2088# 0.367635f
C254 source.t18 a_n2210_n2088# 0.124639f
C255 source.t26 a_n2210_n2088# 0.124639f
C256 source.n106 a_n2210_n2088# 0.970701f
C257 source.n107 a_n2210_n2088# 0.367635f
C258 source.n108 a_n2210_n2088# 0.03695f
C259 source.n109 a_n2210_n2088# 0.026288f
C260 source.n110 a_n2210_n2088# 0.014126f
C261 source.n111 a_n2210_n2088# 0.033388f
C262 source.n112 a_n2210_n2088# 0.014957f
C263 source.n113 a_n2210_n2088# 0.026288f
C264 source.n114 a_n2210_n2088# 0.014126f
C265 source.n115 a_n2210_n2088# 0.033388f
C266 source.n116 a_n2210_n2088# 0.014957f
C267 source.n117 a_n2210_n2088# 0.112492f
C268 source.t15 a_n2210_n2088# 0.054418f
C269 source.n118 a_n2210_n2088# 0.025041f
C270 source.n119 a_n2210_n2088# 0.019722f
C271 source.n120 a_n2210_n2088# 0.014126f
C272 source.n121 a_n2210_n2088# 0.625487f
C273 source.n122 a_n2210_n2088# 0.026288f
C274 source.n123 a_n2210_n2088# 0.014126f
C275 source.n124 a_n2210_n2088# 0.014957f
C276 source.n125 a_n2210_n2088# 0.033388f
C277 source.n126 a_n2210_n2088# 0.033388f
C278 source.n127 a_n2210_n2088# 0.014957f
C279 source.n128 a_n2210_n2088# 0.014126f
C280 source.n129 a_n2210_n2088# 0.026288f
C281 source.n130 a_n2210_n2088# 0.026288f
C282 source.n131 a_n2210_n2088# 0.014126f
C283 source.n132 a_n2210_n2088# 0.014957f
C284 source.n133 a_n2210_n2088# 0.033388f
C285 source.n134 a_n2210_n2088# 0.07228f
C286 source.n135 a_n2210_n2088# 0.014957f
C287 source.n136 a_n2210_n2088# 0.014126f
C288 source.n137 a_n2210_n2088# 0.060762f
C289 source.n138 a_n2210_n2088# 0.040444f
C290 source.n139 a_n2210_n2088# 1.00437f
C291 source.n140 a_n2210_n2088# 0.03695f
C292 source.n141 a_n2210_n2088# 0.026288f
C293 source.n142 a_n2210_n2088# 0.014126f
C294 source.n143 a_n2210_n2088# 0.033388f
C295 source.n144 a_n2210_n2088# 0.014957f
C296 source.n145 a_n2210_n2088# 0.026288f
C297 source.n146 a_n2210_n2088# 0.014126f
C298 source.n147 a_n2210_n2088# 0.033388f
C299 source.n148 a_n2210_n2088# 0.014957f
C300 source.n149 a_n2210_n2088# 0.112492f
C301 source.t14 a_n2210_n2088# 0.054418f
C302 source.n150 a_n2210_n2088# 0.025041f
C303 source.n151 a_n2210_n2088# 0.019722f
C304 source.n152 a_n2210_n2088# 0.014126f
C305 source.n153 a_n2210_n2088# 0.625487f
C306 source.n154 a_n2210_n2088# 0.026288f
C307 source.n155 a_n2210_n2088# 0.014126f
C308 source.n156 a_n2210_n2088# 0.014957f
C309 source.n157 a_n2210_n2088# 0.033388f
C310 source.n158 a_n2210_n2088# 0.033388f
C311 source.n159 a_n2210_n2088# 0.014957f
C312 source.n160 a_n2210_n2088# 0.014126f
C313 source.n161 a_n2210_n2088# 0.026288f
C314 source.n162 a_n2210_n2088# 0.026288f
C315 source.n163 a_n2210_n2088# 0.014126f
C316 source.n164 a_n2210_n2088# 0.014957f
C317 source.n165 a_n2210_n2088# 0.033388f
C318 source.n166 a_n2210_n2088# 0.07228f
C319 source.n167 a_n2210_n2088# 0.014957f
C320 source.n168 a_n2210_n2088# 0.014126f
C321 source.n169 a_n2210_n2088# 0.060762f
C322 source.n170 a_n2210_n2088# 0.040444f
C323 source.n171 a_n2210_n2088# 1.00437f
C324 source.t8 a_n2210_n2088# 0.124639f
C325 source.t2 a_n2210_n2088# 0.124639f
C326 source.n172 a_n2210_n2088# 0.970695f
C327 source.n173 a_n2210_n2088# 0.367642f
C328 source.t3 a_n2210_n2088# 0.124639f
C329 source.t31 a_n2210_n2088# 0.124639f
C330 source.n174 a_n2210_n2088# 0.970695f
C331 source.n175 a_n2210_n2088# 0.367642f
C332 source.t13 a_n2210_n2088# 0.124639f
C333 source.t5 a_n2210_n2088# 0.124639f
C334 source.n176 a_n2210_n2088# 0.970695f
C335 source.n177 a_n2210_n2088# 0.367642f
C336 source.n178 a_n2210_n2088# 0.03695f
C337 source.n179 a_n2210_n2088# 0.026288f
C338 source.n180 a_n2210_n2088# 0.014126f
C339 source.n181 a_n2210_n2088# 0.033388f
C340 source.n182 a_n2210_n2088# 0.014957f
C341 source.n183 a_n2210_n2088# 0.026288f
C342 source.n184 a_n2210_n2088# 0.014126f
C343 source.n185 a_n2210_n2088# 0.033388f
C344 source.n186 a_n2210_n2088# 0.014957f
C345 source.n187 a_n2210_n2088# 0.112492f
C346 source.t10 a_n2210_n2088# 0.054418f
C347 source.n188 a_n2210_n2088# 0.025041f
C348 source.n189 a_n2210_n2088# 0.019722f
C349 source.n190 a_n2210_n2088# 0.014126f
C350 source.n191 a_n2210_n2088# 0.625487f
C351 source.n192 a_n2210_n2088# 0.026288f
C352 source.n193 a_n2210_n2088# 0.014126f
C353 source.n194 a_n2210_n2088# 0.014957f
C354 source.n195 a_n2210_n2088# 0.033388f
C355 source.n196 a_n2210_n2088# 0.033388f
C356 source.n197 a_n2210_n2088# 0.014957f
C357 source.n198 a_n2210_n2088# 0.014126f
C358 source.n199 a_n2210_n2088# 0.026288f
C359 source.n200 a_n2210_n2088# 0.026288f
C360 source.n201 a_n2210_n2088# 0.014126f
C361 source.n202 a_n2210_n2088# 0.014957f
C362 source.n203 a_n2210_n2088# 0.033388f
C363 source.n204 a_n2210_n2088# 0.07228f
C364 source.n205 a_n2210_n2088# 0.014957f
C365 source.n206 a_n2210_n2088# 0.014126f
C366 source.n207 a_n2210_n2088# 0.060762f
C367 source.n208 a_n2210_n2088# 0.040444f
C368 source.n209 a_n2210_n2088# 0.122855f
C369 source.n210 a_n2210_n2088# 0.03695f
C370 source.n211 a_n2210_n2088# 0.026288f
C371 source.n212 a_n2210_n2088# 0.014126f
C372 source.n213 a_n2210_n2088# 0.033388f
C373 source.n214 a_n2210_n2088# 0.014957f
C374 source.n215 a_n2210_n2088# 0.026288f
C375 source.n216 a_n2210_n2088# 0.014126f
C376 source.n217 a_n2210_n2088# 0.033388f
C377 source.n218 a_n2210_n2088# 0.014957f
C378 source.n219 a_n2210_n2088# 0.112492f
C379 source.t21 a_n2210_n2088# 0.054418f
C380 source.n220 a_n2210_n2088# 0.025041f
C381 source.n221 a_n2210_n2088# 0.019722f
C382 source.n222 a_n2210_n2088# 0.014126f
C383 source.n223 a_n2210_n2088# 0.625487f
C384 source.n224 a_n2210_n2088# 0.026288f
C385 source.n225 a_n2210_n2088# 0.014126f
C386 source.n226 a_n2210_n2088# 0.014957f
C387 source.n227 a_n2210_n2088# 0.033388f
C388 source.n228 a_n2210_n2088# 0.033388f
C389 source.n229 a_n2210_n2088# 0.014957f
C390 source.n230 a_n2210_n2088# 0.014126f
C391 source.n231 a_n2210_n2088# 0.026288f
C392 source.n232 a_n2210_n2088# 0.026288f
C393 source.n233 a_n2210_n2088# 0.014126f
C394 source.n234 a_n2210_n2088# 0.014957f
C395 source.n235 a_n2210_n2088# 0.033388f
C396 source.n236 a_n2210_n2088# 0.07228f
C397 source.n237 a_n2210_n2088# 0.014957f
C398 source.n238 a_n2210_n2088# 0.014126f
C399 source.n239 a_n2210_n2088# 0.060762f
C400 source.n240 a_n2210_n2088# 0.040444f
C401 source.n241 a_n2210_n2088# 0.122855f
C402 source.t20 a_n2210_n2088# 0.124639f
C403 source.t29 a_n2210_n2088# 0.124639f
C404 source.n242 a_n2210_n2088# 0.970695f
C405 source.n243 a_n2210_n2088# 0.367642f
C406 source.t23 a_n2210_n2088# 0.124639f
C407 source.t28 a_n2210_n2088# 0.124639f
C408 source.n244 a_n2210_n2088# 0.970695f
C409 source.n245 a_n2210_n2088# 0.367642f
C410 source.t25 a_n2210_n2088# 0.124639f
C411 source.t27 a_n2210_n2088# 0.124639f
C412 source.n246 a_n2210_n2088# 0.970695f
C413 source.n247 a_n2210_n2088# 0.367642f
C414 source.n248 a_n2210_n2088# 0.03695f
C415 source.n249 a_n2210_n2088# 0.026288f
C416 source.n250 a_n2210_n2088# 0.014126f
C417 source.n251 a_n2210_n2088# 0.033388f
C418 source.n252 a_n2210_n2088# 0.014957f
C419 source.n253 a_n2210_n2088# 0.026288f
C420 source.n254 a_n2210_n2088# 0.014126f
C421 source.n255 a_n2210_n2088# 0.033388f
C422 source.n256 a_n2210_n2088# 0.014957f
C423 source.n257 a_n2210_n2088# 0.112492f
C424 source.t30 a_n2210_n2088# 0.054418f
C425 source.n258 a_n2210_n2088# 0.025041f
C426 source.n259 a_n2210_n2088# 0.019722f
C427 source.n260 a_n2210_n2088# 0.014126f
C428 source.n261 a_n2210_n2088# 0.625487f
C429 source.n262 a_n2210_n2088# 0.026288f
C430 source.n263 a_n2210_n2088# 0.014126f
C431 source.n264 a_n2210_n2088# 0.014957f
C432 source.n265 a_n2210_n2088# 0.033388f
C433 source.n266 a_n2210_n2088# 0.033388f
C434 source.n267 a_n2210_n2088# 0.014957f
C435 source.n268 a_n2210_n2088# 0.014126f
C436 source.n269 a_n2210_n2088# 0.026288f
C437 source.n270 a_n2210_n2088# 0.026288f
C438 source.n271 a_n2210_n2088# 0.014126f
C439 source.n272 a_n2210_n2088# 0.014957f
C440 source.n273 a_n2210_n2088# 0.033388f
C441 source.n274 a_n2210_n2088# 0.07228f
C442 source.n275 a_n2210_n2088# 0.014957f
C443 source.n276 a_n2210_n2088# 0.014126f
C444 source.n277 a_n2210_n2088# 0.060762f
C445 source.n278 a_n2210_n2088# 0.040444f
C446 source.n279 a_n2210_n2088# 0.282854f
C447 source.n280 a_n2210_n2088# 1.08283f
C448 minus.n0 a_n2210_n2088# 0.045557f
C449 minus.t8 a_n2210_n2088# 0.396418f
C450 minus.n1 a_n2210_n2088# 0.191511f
C451 minus.n2 a_n2210_n2088# 0.045557f
C452 minus.n3 a_n2210_n2088# 0.010338f
C453 minus.t13 a_n2210_n2088# 0.396418f
C454 minus.n4 a_n2210_n2088# 0.145045f
C455 minus.t3 a_n2210_n2088# 0.396418f
C456 minus.t10 a_n2210_n2088# 0.4065f
C457 minus.n5 a_n2210_n2088# 0.176986f
C458 minus.n6 a_n2210_n2088# 0.188843f
C459 minus.n7 a_n2210_n2088# 0.010338f
C460 minus.t7 a_n2210_n2088# 0.396418f
C461 minus.n8 a_n2210_n2088# 0.191511f
C462 minus.n9 a_n2210_n2088# 0.045557f
C463 minus.n10 a_n2210_n2088# 0.045557f
C464 minus.n11 a_n2210_n2088# 0.045557f
C465 minus.n12 a_n2210_n2088# 0.189124f
C466 minus.t6 a_n2210_n2088# 0.396418f
C467 minus.n13 a_n2210_n2088# 0.189124f
C468 minus.n14 a_n2210_n2088# 0.010338f
C469 minus.n15 a_n2210_n2088# 0.045557f
C470 minus.n16 a_n2210_n2088# 0.045557f
C471 minus.n17 a_n2210_n2088# 0.045557f
C472 minus.n18 a_n2210_n2088# 0.010338f
C473 minus.t0 a_n2210_n2088# 0.396418f
C474 minus.n19 a_n2210_n2088# 0.188843f
C475 minus.t9 a_n2210_n2088# 0.396418f
C476 minus.n20 a_n2210_n2088# 0.186736f
C477 minus.n21 a_n2210_n2088# 1.39222f
C478 minus.n22 a_n2210_n2088# 0.045557f
C479 minus.t5 a_n2210_n2088# 0.396418f
C480 minus.n23 a_n2210_n2088# 0.191511f
C481 minus.n24 a_n2210_n2088# 0.045557f
C482 minus.n25 a_n2210_n2088# 0.010338f
C483 minus.n26 a_n2210_n2088# 0.145045f
C484 minus.t12 a_n2210_n2088# 0.4065f
C485 minus.n27 a_n2210_n2088# 0.176986f
C486 minus.t11 a_n2210_n2088# 0.396418f
C487 minus.n28 a_n2210_n2088# 0.188843f
C488 minus.n29 a_n2210_n2088# 0.010338f
C489 minus.t2 a_n2210_n2088# 0.396418f
C490 minus.n30 a_n2210_n2088# 0.191511f
C491 minus.n31 a_n2210_n2088# 0.045557f
C492 minus.n32 a_n2210_n2088# 0.045557f
C493 minus.n33 a_n2210_n2088# 0.045557f
C494 minus.t1 a_n2210_n2088# 0.396418f
C495 minus.n34 a_n2210_n2088# 0.189124f
C496 minus.t14 a_n2210_n2088# 0.396418f
C497 minus.n35 a_n2210_n2088# 0.189124f
C498 minus.n36 a_n2210_n2088# 0.010338f
C499 minus.n37 a_n2210_n2088# 0.045557f
C500 minus.n38 a_n2210_n2088# 0.045557f
C501 minus.n39 a_n2210_n2088# 0.045557f
C502 minus.n40 a_n2210_n2088# 0.010338f
C503 minus.t4 a_n2210_n2088# 0.396418f
C504 minus.n41 a_n2210_n2088# 0.188843f
C505 minus.t15 a_n2210_n2088# 0.396418f
C506 minus.n42 a_n2210_n2088# 0.186736f
C507 minus.n43 a_n2210_n2088# 0.304376f
C508 minus.n44 a_n2210_n2088# 1.70359f
.ends

