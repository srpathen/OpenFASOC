* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp output vdd plus minus commonsourceibias outputibias diffpairibias gnd CSoutput
Cload output gnd 0.0p
X0 gnd.t124 gnd.t121 gnd.t123 gnd.t122 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X1 commonsourceibias.t47 commonsourceibias.t46 gnd.t141 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X2 gnd.t153 commonsourceibias.t48 CSoutput.t58 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X3 gnd.t120 gnd.t118 gnd.t119 gnd.t106 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X4 vdd.t282 a_n7636_8799.t36 CSoutput.t111 vdd.t153 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X5 a_n1986_8322.t11 a_n2848_n452.t48 vdd.t293 vdd.t292 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X6 a_n1808_13878.t19 a_n2848_n452.t21 a_n2848_n452.t22 vdd.t11 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X7 a_n7636_8799.t33 plus.t5 a_n3106_n452.t28 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X8 output.t3 outputibias.t8 gnd.t176 gnd.t175 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X9 gnd.t126 commonsourceibias.t49 CSoutput.t57 gnd.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 a_n3106_n452.t27 plus.t6 a_n7636_8799.t15 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X11 vdd.t23 CSoutput.t168 output.t19 gnd.t170 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X12 a_n2848_n452.t24 a_n2848_n452.t23 a_n1808_13878.t18 vdd.t116 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X13 a_n1808_13878.t17 a_n2848_n452.t27 a_n2848_n452.t28 vdd.t283 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X14 vdd.t109 vdd.t107 vdd.t108 vdd.t85 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X15 CSoutput.t83 a_n7636_8799.t37 vdd.t281 vdd.t221 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X16 a_n1808_13878.t7 a_n2848_n452.t49 vdd.t295 vdd.t294 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X17 gnd.t291 commonsourceibias.t44 commonsourceibias.t45 gnd.t137 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 vdd.t22 CSoutput.t169 output.t18 gnd.t171 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X19 CSoutput.t65 a_n7636_8799.t38 vdd.t280 vdd.t133 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X20 vdd.t279 a_n7636_8799.t39 CSoutput.t82 vdd.t215 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 gnd.t138 commonsourceibias.t50 CSoutput.t56 gnd.t137 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 outputibias.t7 outputibias.t6 gnd.t277 gnd.t276 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X23 CSoutput.t154 a_n7636_8799.t40 vdd.t278 vdd.t137 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X24 vdd.t106 vdd.t104 vdd.t105 vdd.t57 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X25 a_n1986_8322.t23 a_n2848_n452.t50 a_n7636_8799.t18 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X26 a_n2848_n452.t12 minus.t5 a_n3106_n452.t43 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X27 a_n7636_8799.t31 plus.t7 a_n3106_n452.t26 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X28 gnd.t204 commonsourceibias.t42 commonsourceibias.t43 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X29 CSoutput.t120 a_n7636_8799.t41 vdd.t277 vdd.t179 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X30 plus.t4 gnd.t115 gnd.t117 gnd.t116 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X31 a_n2848_n452.t11 minus.t6 a_n3106_n452.t42 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X32 vdd.t276 a_n7636_8799.t42 CSoutput.t110 vdd.t208 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X33 CSoutput.t55 commonsourceibias.t51 gnd.t270 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X34 CSoutput.t170 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X35 gnd.t226 commonsourceibias.t40 commonsourceibias.t41 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 vdd.t275 a_n7636_8799.t43 CSoutput.t130 vdd.t231 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X37 CSoutput.t145 a_n7636_8799.t44 vdd.t274 vdd.t181 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X38 vdd.t273 a_n7636_8799.t45 CSoutput.t132 vdd.t235 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X39 a_n3106_n452.t25 plus.t8 a_n7636_8799.t7 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X40 a_n7636_8799.t19 a_n2848_n452.t51 a_n1986_8322.t22 vdd.t11 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X41 CSoutput.t151 a_n7636_8799.t46 vdd.t272 vdd.t123 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X42 vdd.t271 a_n7636_8799.t47 CSoutput.t102 vdd.t260 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X43 a_n3106_n452.t41 minus.t7 a_n2848_n452.t10 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X44 CSoutput.t54 commonsourceibias.t52 gnd.t139 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X45 a_n3106_n452.t36 diffpairibias.t16 gnd.t218 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X46 output.t17 CSoutput.t171 vdd.t31 gnd.t127 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X47 vdd.t21 CSoutput.t172 output.t16 gnd.t128 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X48 CSoutput.t53 commonsourceibias.t53 gnd.t266 gnd.t241 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 CSoutput.t68 a_n7636_8799.t48 vdd.t270 vdd.t171 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X50 CSoutput.t141 a_n7636_8799.t49 vdd.t269 vdd.t221 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X51 vdd.t103 vdd.t101 vdd.t102 vdd.t35 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X52 CSoutput.t52 commonsourceibias.t54 gnd.t268 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X53 gnd.t114 gnd.t112 gnd.t113 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X54 CSoutput.t60 a_n7636_8799.t50 vdd.t268 vdd.t137 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X55 a_n3106_n452.t24 plus.t9 a_n7636_8799.t26 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X56 a_n1808_13878.t16 a_n2848_n452.t29 a_n2848_n452.t30 vdd.t113 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X57 vdd.t100 vdd.t98 vdd.t99 vdd.t57 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X58 vdd.t267 a_n7636_8799.t51 CSoutput.t71 vdd.t260 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X59 a_n3106_n452.t23 plus.t10 a_n7636_8799.t9 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X60 a_n3106_n452.t40 minus.t8 a_n2848_n452.t9 gnd.t222 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X61 diffpairibias.t15 diffpairibias.t14 gnd.t282 gnd.t281 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X62 a_n2848_n452.t40 a_n2848_n452.t39 a_n1808_13878.t15 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X63 CSoutput.t152 a_n7636_8799.t52 vdd.t266 vdd.t213 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X64 gnd.t111 gnd.t109 gnd.t110 gnd.t106 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X65 vdd.t97 vdd.t95 vdd.t96 vdd.t70 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X66 CSoutput.t89 a_n7636_8799.t53 vdd.t265 vdd.t179 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X67 vdd.t264 a_n7636_8799.t54 CSoutput.t150 vdd.t208 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X68 gnd.t272 commonsourceibias.t55 CSoutput.t51 gnd.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X69 gnd.t260 commonsourceibias.t56 CSoutput.t50 gnd.t256 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 diffpairibias.t13 diffpairibias.t12 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X71 CSoutput.t107 a_n7636_8799.t55 vdd.t263 vdd.t217 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 gnd.t269 commonsourceibias.t57 CSoutput.t49 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X73 commonsourceibias.t39 commonsourceibias.t38 gnd.t245 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 vdd.t262 a_n7636_8799.t56 CSoutput.t101 vdd.t231 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X75 vdd.t261 a_n7636_8799.t57 CSoutput.t87 vdd.t260 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X76 vdd.t259 a_n7636_8799.t58 CSoutput.t97 vdd.t145 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X77 vdd.t27 CSoutput.t173 output.t15 gnd.t142 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X78 CSoutput.t163 a_n7636_8799.t59 vdd.t258 vdd.t151 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X79 vdd.t257 a_n7636_8799.t60 CSoutput.t162 vdd.t206 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X80 CSoutput.t92 a_n7636_8799.t61 vdd.t256 vdd.t123 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X81 a_n3106_n452.t39 minus.t9 a_n2848_n452.t8 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X82 a_n3106_n452.t22 plus.t11 a_n7636_8799.t32 gnd.t280 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X83 vdd.t255 a_n7636_8799.t62 CSoutput.t0 vdd.t131 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X84 gnd.t279 commonsourceibias.t58 CSoutput.t48 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 a_n7636_8799.t34 plus.t12 a_n3106_n452.t21 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X86 commonsourceibias.t37 commonsourceibias.t36 gnd.t182 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 CSoutput.t131 a_n7636_8799.t63 vdd.t254 vdd.t189 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X88 CSoutput.t115 a_n7636_8799.t64 vdd.t253 vdd.t171 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X89 CSoutput.t135 a_n7636_8799.t65 vdd.t252 vdd.t239 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X90 a_n3106_n452.t33 diffpairibias.t17 gnd.t192 gnd.t191 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X91 gnd.t275 commonsourceibias.t34 commonsourceibias.t35 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X92 CSoutput.t136 a_n7636_8799.t66 vdd.t251 vdd.t239 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X93 a_n3106_n452.t20 plus.t13 a_n7636_8799.t20 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X94 vdd.t250 a_n7636_8799.t67 CSoutput.t137 vdd.t237 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X95 gnd.t278 commonsourceibias.t32 commonsourceibias.t33 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X96 commonsourceibias.t31 commonsourceibias.t30 gnd.t242 gnd.t241 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X97 vdd.t249 a_n7636_8799.t68 CSoutput.t123 vdd.t203 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X98 a_n2848_n452.t26 a_n2848_n452.t25 a_n1808_13878.t14 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X99 outputibias.t5 outputibias.t4 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X100 a_n2848_n452.t36 a_n2848_n452.t35 a_n1808_13878.t13 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X101 vdd.t248 a_n7636_8799.t69 CSoutput.t6 vdd.t235 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 vdd.t247 a_n7636_8799.t70 CSoutput.t7 vdd.t183 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X103 a_n7636_8799.t4 a_n2848_n452.t52 a_n1986_8322.t21 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X104 CSoutput.t47 commonsourceibias.t59 gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X105 vdd.t246 a_n7636_8799.t71 CSoutput.t161 vdd.t237 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X106 a_n2848_n452.t13 minus.t10 a_n3106_n452.t44 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X107 CSoutput.t46 commonsourceibias.t60 gnd.t186 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 vdd.t245 a_n7636_8799.t72 CSoutput.t138 vdd.t149 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X109 gnd.t12 commonsourceibias.t61 CSoutput.t45 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X110 gnd.t108 gnd.t105 gnd.t107 gnd.t106 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X111 commonsourceibias.t29 commonsourceibias.t28 gnd.t285 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X112 CSoutput.t129 a_n7636_8799.t73 vdd.t244 vdd.t185 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X113 CSoutput.t44 commonsourceibias.t62 gnd.t255 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X114 CSoutput.t174 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X115 outputibias.t3 outputibias.t2 gnd.t287 gnd.t286 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X116 vdd.t243 a_n7636_8799.t74 CSoutput.t126 vdd.t206 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X117 vdd.t94 vdd.t92 vdd.t93 vdd.t78 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X118 CSoutput.t73 a_n7636_8799.t75 vdd.t242 vdd.t151 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X119 vdd.t91 vdd.t88 vdd.t90 vdd.t89 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X120 a_n3106_n452.t0 diffpairibias.t18 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X121 vdd.t87 vdd.t84 vdd.t86 vdd.t85 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X122 gnd.t104 gnd.t102 minus.t4 gnd.t103 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X123 gnd.t101 gnd.t99 gnd.t100 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X124 commonsourceibias.t27 commonsourceibias.t26 gnd.t9 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X125 vdd.t6 a_n2848_n452.t53 a_n1986_8322.t10 vdd.t5 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X126 vdd.t83 vdd.t81 vdd.t82 vdd.t74 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X127 CSoutput.t103 a_n7636_8799.t76 vdd.t241 vdd.t189 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X128 CSoutput.t128 a_n7636_8799.t77 vdd.t240 vdd.t239 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X129 a_n1986_8322.t9 a_n2848_n452.t54 vdd.t13 vdd.t12 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X130 vdd.t238 a_n7636_8799.t78 CSoutput.t134 vdd.t237 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X131 gnd.t284 commonsourceibias.t24 commonsourceibias.t25 gnd.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X132 gnd.t257 commonsourceibias.t63 CSoutput.t43 gnd.t256 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 vdd.t15 a_n2848_n452.t55 a_n1808_13878.t6 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X134 gnd.t98 gnd.t96 plus.t3 gnd.t97 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X135 gnd.t258 commonsourceibias.t64 CSoutput.t42 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X136 a_n2848_n452.t19 minus.t11 a_n3106_n452.t50 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X137 a_n7636_8799.t35 plus.t14 a_n3106_n452.t19 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X138 gnd.t261 commonsourceibias.t65 CSoutput.t41 gnd.t233 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X139 vdd.t80 vdd.t77 vdd.t79 vdd.t78 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X140 a_n7636_8799.t0 plus.t15 a_n3106_n452.t18 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X141 a_n2848_n452.t18 minus.t12 a_n3106_n452.t49 gnd.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X142 diffpairibias.t11 diffpairibias.t10 gnd.t136 gnd.t135 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X143 vdd.t17 CSoutput.t175 output.t14 gnd.t143 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X144 vdd.t76 vdd.t73 vdd.t75 vdd.t74 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X145 vdd.t236 a_n7636_8799.t79 CSoutput.t10 vdd.t235 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X146 gnd.t262 commonsourceibias.t66 CSoutput.t40 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X147 outputibias.t1 outputibias.t0 gnd.t185 gnd.t184 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X148 a_n7636_8799.t21 a_n2848_n452.t56 a_n1986_8322.t20 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X149 a_n1986_8322.t8 a_n2848_n452.t57 vdd.t122 vdd.t121 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X150 vdd.t72 vdd.t69 vdd.t71 vdd.t70 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X151 CSoutput.t4 a_n7636_8799.t80 vdd.t234 vdd.t165 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X152 gnd.t265 commonsourceibias.t67 CSoutput.t39 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X153 vdd.t233 a_n7636_8799.t81 CSoutput.t61 vdd.t149 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X154 vdd.t232 a_n7636_8799.t82 CSoutput.t106 vdd.t231 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X155 a_n2848_n452.t34 a_n2848_n452.t33 a_n1808_13878.t12 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X156 a_n3106_n452.t48 minus.t13 a_n2848_n452.t17 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X157 CSoutput.t176 a_n1986_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X158 CSoutput.t59 a_n7636_8799.t83 vdd.t230 vdd.t185 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 a_n7636_8799.t25 a_n2848_n452.t58 a_n1986_8322.t19 vdd.t283 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X160 CSoutput.t38 commonsourceibias.t68 gnd.t129 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 CSoutput.t177 a_n1986_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X162 a_n1808_13878.t11 a_n2848_n452.t31 a_n2848_n452.t32 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X163 a_n3106_n452.t17 plus.t16 a_n7636_8799.t22 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X164 a_n2848_n452.t16 minus.t14 a_n3106_n452.t47 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X165 vdd.t229 a_n7636_8799.t84 CSoutput.t119 vdd.t215 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X166 CSoutput.t81 a_n7636_8799.t85 vdd.t228 vdd.t217 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X167 vdd.t285 a_n2848_n452.t59 a_n1986_8322.t7 vdd.t284 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X168 gnd.t95 gnd.t92 gnd.t94 gnd.t93 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X169 a_n3106_n452.t38 diffpairibias.t19 gnd.t236 gnd.t235 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X170 CSoutput.t109 a_n7636_8799.t86 vdd.t227 vdd.t213 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X171 CSoutput.t37 commonsourceibias.t69 gnd.t214 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X172 a_n7636_8799.t8 plus.t17 a_n3106_n452.t16 gnd.t160 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X173 CSoutput.t36 commonsourceibias.t70 gnd.t248 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X174 a_n3106_n452.t34 diffpairibias.t20 gnd.t201 gnd.t200 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X175 vdd.t226 a_n7636_8799.t87 CSoutput.t5 vdd.t125 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X176 vdd.t225 a_n7636_8799.t88 CSoutput.t118 vdd.t162 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X177 gnd.t150 commonsourceibias.t71 CSoutput.t35 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X178 CSoutput.t34 commonsourceibias.t72 gnd.t215 gnd.t146 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X179 a_n7636_8799.t11 plus.t18 a_n3106_n452.t15 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X180 vdd.t224 a_n7636_8799.t89 CSoutput.t116 vdd.t203 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X181 vdd.t223 a_n7636_8799.t90 CSoutput.t117 vdd.t173 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X182 minus.t3 gnd.t89 gnd.t91 gnd.t90 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X183 gnd.t88 gnd.t86 gnd.t87 gnd.t42 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X184 diffpairibias.t9 diffpairibias.t8 gnd.t224 gnd.t223 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X185 a_n2848_n452.t15 minus.t15 a_n3106_n452.t46 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X186 CSoutput.t133 a_n7636_8799.t91 vdd.t222 vdd.t221 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X187 CSoutput.t121 a_n7636_8799.t92 vdd.t220 vdd.t127 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X188 a_n3106_n452.t14 plus.t19 a_n7636_8799.t29 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X189 CSoutput.t1 a_n7636_8799.t93 vdd.t219 vdd.t196 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X190 CSoutput.t33 commonsourceibias.t73 gnd.t250 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X191 gnd.t246 commonsourceibias.t74 CSoutput.t32 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X192 vdd.t68 vdd.t66 vdd.t67 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X193 a_n1808_13878.t5 a_n2848_n452.t60 vdd.t289 vdd.t288 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X194 vdd.t291 a_n2848_n452.t61 a_n1808_13878.t4 vdd.t290 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X195 gnd.t228 commonsourceibias.t22 commonsourceibias.t23 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 gnd.t273 commonsourceibias.t75 CSoutput.t31 gnd.t233 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X197 output.t13 CSoutput.t178 vdd.t24 gnd.t161 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X198 vdd.t65 vdd.t63 vdd.t64 vdd.t50 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X199 CSoutput.t148 a_n7636_8799.t94 vdd.t218 vdd.t217 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X200 vdd.t216 a_n7636_8799.t95 CSoutput.t146 vdd.t215 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X201 vdd.t62 vdd.t60 vdd.t61 vdd.t50 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X202 gnd.t187 commonsourceibias.t76 CSoutput.t30 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 a_n3106_n452.t45 minus.t16 a_n2848_n452.t14 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X204 diffpairibias.t7 diffpairibias.t6 gnd.t220 gnd.t219 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X205 CSoutput.t62 a_n7636_8799.t96 vdd.t214 vdd.t213 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X206 gnd.t173 commonsourceibias.t20 commonsourceibias.t21 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 output.t12 CSoutput.t179 vdd.t29 gnd.t162 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X208 vdd.t212 a_n7636_8799.t97 CSoutput.t149 vdd.t125 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X209 vdd.t211 a_n7636_8799.t98 CSoutput.t70 vdd.t162 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X210 CSoutput.t29 commonsourceibias.t77 gnd.t253 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X211 a_n3106_n452.t51 minus.t17 a_n2848_n452.t20 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X212 a_n3106_n452.t13 plus.t20 a_n7636_8799.t24 gnd.t222 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X213 gnd.t85 gnd.t83 gnd.t84 gnd.t42 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X214 gnd.t82 gnd.t80 gnd.t81 gnd.t21 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X215 a_n1986_8322.t18 a_n2848_n452.t62 a_n7636_8799.t27 vdd.t116 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X216 CSoutput.t143 a_n7636_8799.t99 vdd.t210 vdd.t168 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 CSoutput.t28 commonsourceibias.t78 gnd.t14 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 a_n3106_n452.t55 minus.t18 a_n2848_n452.t47 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X219 vdd.t209 a_n7636_8799.t100 CSoutput.t100 vdd.t208 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X220 vdd.t207 a_n7636_8799.t101 CSoutput.t69 vdd.t206 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X221 CSoutput.t158 a_n7636_8799.t102 vdd.t205 vdd.t141 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X222 vdd.t204 a_n7636_8799.t103 CSoutput.t155 vdd.t203 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X223 vdd.t202 a_n7636_8799.t104 CSoutput.t64 vdd.t173 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X224 vdd.t287 a_n2848_n452.t63 a_n1986_8322.t6 vdd.t286 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X225 gnd.t165 commonsourceibias.t18 commonsourceibias.t19 gnd.t164 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 a_n1808_13878.t3 a_n2848_n452.t64 vdd.t2 vdd.t1 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X227 gnd.t79 gnd.t76 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X228 minus.t2 gnd.t73 gnd.t75 gnd.t74 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X229 CSoutput.t27 commonsourceibias.t79 gnd.t213 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X230 a_n3106_n452.t4 diffpairibias.t21 gnd.t167 gnd.t166 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X231 vdd.t201 a_n7636_8799.t105 CSoutput.t108 vdd.t183 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X232 CSoutput.t147 a_n7636_8799.t106 vdd.t200 vdd.t196 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X233 a_n7636_8799.t28 plus.t21 a_n3106_n452.t12 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X234 a_n2848_n452.t7 minus.t19 a_n3106_n452.t37 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X235 CSoutput.t26 commonsourceibias.t80 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X236 output.t11 CSoutput.t180 vdd.t20 gnd.t163 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X237 CSoutput.t142 a_n7636_8799.t107 vdd.t199 vdd.t181 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X238 vdd.t59 vdd.t56 vdd.t58 vdd.t57 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X239 a_n3106_n452.t54 minus.t20 a_n2848_n452.t46 gnd.t280 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X240 CSoutput.t181 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X241 vdd.t55 vdd.t53 vdd.t54 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X242 CSoutput.t25 commonsourceibias.t81 gnd.t147 gnd.t146 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 gnd.t62 gnd.t59 gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X244 a_n1986_8322.t17 a_n2848_n452.t65 a_n7636_8799.t3 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X245 vdd.t8 a_n2848_n452.t66 a_n1986_8322.t5 vdd.t7 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X246 vdd.t52 vdd.t49 vdd.t51 vdd.t50 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X247 vdd.t198 a_n7636_8799.t108 CSoutput.t66 vdd.t153 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X248 CSoutput.t80 a_n7636_8799.t109 vdd.t197 vdd.t196 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X249 gnd.t247 commonsourceibias.t82 CSoutput.t24 gnd.t164 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X250 output.t2 outputibias.t9 gnd.t145 gnd.t144 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X251 CSoutput.t153 a_n7636_8799.t110 vdd.t195 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X252 a_n3106_n452.t52 minus.t21 a_n2848_n452.t45 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X253 gnd.t72 gnd.t70 gnd.t71 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X254 vdd.t30 CSoutput.t182 output.t10 gnd.t188 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X255 vdd.t194 a_n7636_8799.t111 CSoutput.t140 vdd.t176 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X256 vdd.t193 a_n7636_8799.t112 CSoutput.t144 vdd.t135 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X257 a_n3106_n452.t29 minus.t22 a_n2848_n452.t2 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X258 gnd.t69 gnd.t67 gnd.t68 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X259 output.t1 outputibias.t10 gnd.t230 gnd.t229 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X260 diffpairibias.t5 diffpairibias.t4 gnd.t169 gnd.t168 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X261 vdd.t48 vdd.t45 vdd.t47 vdd.t46 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X262 vdd.t192 a_n7636_8799.t113 CSoutput.t79 vdd.t129 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X263 CSoutput.t63 a_n7636_8799.t114 vdd.t191 vdd.t168 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X264 CSoutput.t165 a_n7636_8799.t115 vdd.t190 vdd.t189 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X265 a_n1808_13878.t10 a_n2848_n452.t41 a_n2848_n452.t42 vdd.t110 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X266 gnd.t158 commonsourceibias.t83 CSoutput.t23 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X267 CSoutput.t22 commonsourceibias.t84 gnd.t254 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X268 a_n1986_8322.t16 a_n2848_n452.t67 a_n7636_8799.t5 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X269 gnd.t66 gnd.t63 gnd.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X270 gnd.t149 commonsourceibias.t85 CSoutput.t21 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X271 gnd.t234 commonsourceibias.t16 commonsourceibias.t17 gnd.t233 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X272 CSoutput.t122 a_n7636_8799.t116 vdd.t188 vdd.t165 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 vdd.t187 a_n7636_8799.t117 CSoutput.t167 vdd.t176 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X274 CSoutput.t112 a_n7636_8799.t118 vdd.t186 vdd.t185 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X275 a_n3106_n452.t2 minus.t23 a_n2848_n452.t1 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X276 gnd.t58 gnd.t55 gnd.t57 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X277 vdd.t25 CSoutput.t183 output.t9 gnd.t189 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X278 output.t8 CSoutput.t184 vdd.t32 gnd.t190 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X279 vdd.t184 a_n7636_8799.t119 CSoutput.t95 vdd.t183 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X280 CSoutput.t113 a_n7636_8799.t120 vdd.t182 vdd.t181 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X281 a_n1986_8322.t4 a_n2848_n452.t68 vdd.t118 vdd.t117 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X282 gnd.t54 gnd.t52 plus.t2 gnd.t53 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X283 gnd.t51 gnd.t49 gnd.t50 gnd.t21 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X284 CSoutput.t20 commonsourceibias.t86 gnd.t207 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X285 gnd.t48 gnd.t45 gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X286 CSoutput.t19 commonsourceibias.t87 gnd.t210 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 gnd.t44 gnd.t41 gnd.t43 gnd.t42 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X288 output.t7 CSoutput.t185 vdd.t28 gnd.t194 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X289 vdd.t120 a_n2848_n452.t69 a_n1808_13878.t2 vdd.t119 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X290 CSoutput.t86 a_n7636_8799.t121 vdd.t180 vdd.t179 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X291 CSoutput.t77 a_n7636_8799.t122 vdd.t178 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X292 vdd.t177 a_n7636_8799.t123 CSoutput.t94 vdd.t176 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 vdd.t175 a_n7636_8799.t124 CSoutput.t67 vdd.t135 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X294 vdd.t44 vdd.t41 vdd.t43 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X295 a_n1986_8322.t15 a_n2848_n452.t70 a_n7636_8799.t12 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X296 a_n3106_n452.t11 plus.t22 a_n7636_8799.t6 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X297 output.t0 outputibias.t11 gnd.t155 gnd.t154 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X298 vdd.t40 vdd.t38 vdd.t39 vdd.t35 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X299 a_n7636_8799.t13 a_n2848_n452.t71 a_n1986_8322.t14 vdd.t110 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X300 a_n1808_13878.t1 a_n2848_n452.t72 vdd.t112 vdd.t111 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X301 vdd.t174 a_n7636_8799.t125 CSoutput.t96 vdd.t173 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X302 CSoutput.t2 a_n7636_8799.t126 vdd.t172 vdd.t171 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X303 gnd.t40 gnd.t38 minus.t1 gnd.t39 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X304 a_n2848_n452.t0 minus.t24 a_n3106_n452.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X305 a_n7636_8799.t2 plus.t23 a_n3106_n452.t10 gnd.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X306 CSoutput.t18 commonsourceibias.t88 gnd.t232 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 vdd.t170 a_n7636_8799.t127 CSoutput.t99 vdd.t145 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 a_n2848_n452.t3 minus.t25 a_n3106_n452.t30 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X309 CSoutput.t78 a_n7636_8799.t128 vdd.t169 vdd.t168 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X310 commonsourceibias.t15 commonsourceibias.t14 gnd.t156 gnd.t146 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 gnd.t211 commonsourceibias.t89 CSoutput.t17 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X312 vdd.t18 CSoutput.t186 output.t6 gnd.t195 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X313 gnd.t251 commonsourceibias.t90 CSoutput.t16 gnd.t164 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 CSoutput.t3 a_n7636_8799.t129 vdd.t167 vdd.t143 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X315 CSoutput.t105 a_n7636_8799.t130 vdd.t166 vdd.t165 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X316 CSoutput.t160 a_n7636_8799.t131 vdd.t164 vdd.t143 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X317 vdd.t163 a_n7636_8799.t132 CSoutput.t124 vdd.t162 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 CSoutput.t84 a_n7636_8799.t133 vdd.t161 vdd.t141 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 vdd.t160 a_n7636_8799.t134 CSoutput.t76 vdd.t139 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X320 a_n1808_13878.t9 a_n2848_n452.t43 a_n2848_n452.t44 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X321 gnd.t37 gnd.t34 gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X322 a_n3106_n452.t32 minus.t26 a_n2848_n452.t5 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X323 a_n3106_n452.t3 diffpairibias.t22 gnd.t134 gnd.t133 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X324 gnd.t177 commonsourceibias.t91 CSoutput.t15 gnd.t137 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X325 commonsourceibias.t13 commonsourceibias.t12 gnd.t243 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 a_n7636_8799.t23 plus.t24 a_n3106_n452.t9 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X327 CSoutput.t91 a_n7636_8799.t135 vdd.t159 vdd.t133 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X328 vdd.t158 a_n7636_8799.t136 CSoutput.t139 vdd.t131 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X329 CSoutput.t85 a_n7636_8799.t137 vdd.t157 vdd.t127 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X330 vdd.t156 a_n7636_8799.t138 CSoutput.t159 vdd.t129 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X331 diffpairibias.t3 diffpairibias.t2 gnd.t131 gnd.t130 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X332 a_n7636_8799.t14 a_n2848_n452.t73 a_n1986_8322.t13 vdd.t113 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X333 a_n2848_n452.t38 a_n2848_n452.t37 a_n1808_13878.t8 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X334 vdd.t155 a_n7636_8799.t139 CSoutput.t114 vdd.t139 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X335 gnd.t33 gnd.t31 plus.t1 gnd.t32 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X336 a_n2848_n452.t4 minus.t27 a_n3106_n452.t31 gnd.t160 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X337 vdd.t154 a_n7636_8799.t140 CSoutput.t75 vdd.t153 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X338 CSoutput.t90 a_n7636_8799.t141 vdd.t152 vdd.t151 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 commonsourceibias.t11 commonsourceibias.t10 gnd.t193 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X340 gnd.t252 commonsourceibias.t92 CSoutput.t14 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X341 vdd.t37 vdd.t34 vdd.t36 vdd.t35 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X342 vdd.t150 a_n7636_8799.t142 CSoutput.t156 vdd.t149 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X343 CSoutput.t187 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X344 diffpairibias.t1 diffpairibias.t0 gnd.t203 gnd.t202 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X345 CSoutput.t93 a_n7636_8799.t143 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X346 CSoutput.t13 commonsourceibias.t93 gnd.t267 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X347 gnd.t30 gnd.t27 gnd.t29 gnd.t28 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X348 vdd.t146 a_n7636_8799.t144 CSoutput.t74 vdd.t145 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X349 output.t5 CSoutput.t188 vdd.t19 gnd.t205 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X350 plus.t0 gnd.t24 gnd.t26 gnd.t25 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X351 gnd.t23 gnd.t20 gnd.t22 gnd.t21 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X352 CSoutput.t12 commonsourceibias.t94 gnd.t259 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X353 commonsourceibias.t9 commonsourceibias.t8 gnd.t227 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X354 gnd.t19 gnd.t17 minus.t0 gnd.t18 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X355 a_n7636_8799.t10 plus.t25 a_n3106_n452.t8 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X356 CSoutput.t164 a_n7636_8799.t145 vdd.t144 vdd.t143 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X357 vdd.t115 a_n2848_n452.t74 a_n1808_13878.t0 vdd.t114 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X358 CSoutput.t9 a_n7636_8799.t146 vdd.t142 vdd.t141 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X359 CSoutput.t11 commonsourceibias.t95 gnd.t271 gnd.t241 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X360 a_n7636_8799.t1 plus.t26 a_n3106_n452.t7 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X361 a_n2848_n452.t6 minus.t28 a_n3106_n452.t35 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X362 output.t4 CSoutput.t189 vdd.t26 gnd.t206 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X363 vdd.t140 a_n7636_8799.t147 CSoutput.t157 vdd.t139 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X364 CSoutput.t72 a_n7636_8799.t148 vdd.t138 vdd.t137 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X365 vdd.t136 a_n7636_8799.t149 CSoutput.t127 vdd.t135 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X366 gnd.t290 commonsourceibias.t6 commonsourceibias.t7 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X367 commonsourceibias.t5 commonsourceibias.t4 gnd.t263 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X368 CSoutput.t8 a_n7636_8799.t150 vdd.t134 vdd.t133 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X369 vdd.t132 a_n7636_8799.t151 CSoutput.t88 vdd.t131 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X370 vdd.t130 a_n7636_8799.t152 CSoutput.t166 vdd.t129 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X371 a_n1986_8322.t12 a_n2848_n452.t75 a_n7636_8799.t17 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X372 a_n3106_n452.t6 plus.t27 a_n7636_8799.t16 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X373 commonsourceibias.t3 commonsourceibias.t2 gnd.t283 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X374 CSoutput.t125 a_n7636_8799.t153 vdd.t128 vdd.t127 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X375 vdd.t126 a_n7636_8799.t154 CSoutput.t104 vdd.t125 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X376 CSoutput.t98 a_n7636_8799.t155 vdd.t124 vdd.t123 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X377 a_n3106_n452.t5 plus.t28 a_n7636_8799.t30 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X378 gnd.t274 commonsourceibias.t0 commonsourceibias.t1 gnd.t256 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X379 a_n3106_n452.t53 diffpairibias.t23 gnd.t289 gnd.t288 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
R0 gnd.n6679 gnd.n403 2174.34
R1 gnd.n3841 gnd.n3611 939.716
R2 gnd.n6988 gnd.n84 838.452
R3 gnd.n7151 gnd.n80 838.452
R4 gnd.n5287 gnd.n1128 838.452
R5 gnd.n5206 gnd.n1130 838.452
R6 gnd.n5997 gnd.n997 838.452
R7 gnd.n4196 gnd.n995 838.452
R8 gnd.n3698 gnd.n3639 838.452
R9 gnd.n3843 gnd.n2154 838.452
R10 gnd.n7149 gnd.n86 819.232
R11 gnd.n154 gnd.n82 819.232
R12 gnd.n5605 gnd.n1127 819.232
R13 gnd.n5850 gnd.n1131 819.232
R14 gnd.n5999 gnd.n992 819.232
R15 gnd.n4306 gnd.n994 819.232
R16 gnd.n3763 gnd.n3762 819.232
R17 gnd.n3839 gnd.n2150 819.232
R18 gnd.n4242 gnd.n1002 771.183
R19 gnd.n5868 gnd.n1105 771.183
R20 gnd.n4256 gnd.n2019 771.183
R21 gnd.n5320 gnd.n1107 771.183
R22 gnd.n3519 gnd.n2162 766.379
R23 gnd.n3522 gnd.n3521 766.379
R24 gnd.n2760 gnd.n2663 766.379
R25 gnd.n2756 gnd.n2661 766.379
R26 gnd.n3610 gnd.n2184 756.769
R27 gnd.n3513 gnd.n3512 756.769
R28 gnd.n2853 gnd.n2570 756.769
R29 gnd.n2851 gnd.n2573 756.769
R30 gnd.n6260 gnd.n656 756.769
R31 gnd.n6680 gnd.n404 756.769
R32 gnd.n6893 gnd.n277 756.769
R33 gnd.n6092 gnd.n826 756.769
R34 gnd.n6261 gnd.n6260 585
R35 gnd.n6260 gnd.n6259 585
R36 gnd.n660 gnd.n659 585
R37 gnd.n6258 gnd.n660 585
R38 gnd.n6256 gnd.n6255 585
R39 gnd.n6257 gnd.n6256 585
R40 gnd.n6254 gnd.n662 585
R41 gnd.n662 gnd.n661 585
R42 gnd.n6253 gnd.n6252 585
R43 gnd.n6252 gnd.n6251 585
R44 gnd.n667 gnd.n666 585
R45 gnd.n6250 gnd.n667 585
R46 gnd.n6248 gnd.n6247 585
R47 gnd.n6249 gnd.n6248 585
R48 gnd.n6246 gnd.n669 585
R49 gnd.n669 gnd.n668 585
R50 gnd.n6245 gnd.n6244 585
R51 gnd.n6244 gnd.n6243 585
R52 gnd.n675 gnd.n674 585
R53 gnd.n6242 gnd.n675 585
R54 gnd.n6240 gnd.n6239 585
R55 gnd.n6241 gnd.n6240 585
R56 gnd.n6238 gnd.n677 585
R57 gnd.n677 gnd.n676 585
R58 gnd.n6237 gnd.n6236 585
R59 gnd.n6236 gnd.n6235 585
R60 gnd.n683 gnd.n682 585
R61 gnd.n6234 gnd.n683 585
R62 gnd.n6232 gnd.n6231 585
R63 gnd.n6233 gnd.n6232 585
R64 gnd.n6230 gnd.n685 585
R65 gnd.n685 gnd.n684 585
R66 gnd.n6229 gnd.n6228 585
R67 gnd.n6228 gnd.n6227 585
R68 gnd.n691 gnd.n690 585
R69 gnd.n6226 gnd.n691 585
R70 gnd.n6224 gnd.n6223 585
R71 gnd.n6225 gnd.n6224 585
R72 gnd.n6222 gnd.n693 585
R73 gnd.n693 gnd.n692 585
R74 gnd.n6221 gnd.n6220 585
R75 gnd.n6220 gnd.n6219 585
R76 gnd.n699 gnd.n698 585
R77 gnd.n6218 gnd.n699 585
R78 gnd.n6216 gnd.n6215 585
R79 gnd.n6217 gnd.n6216 585
R80 gnd.n6214 gnd.n701 585
R81 gnd.n701 gnd.n700 585
R82 gnd.n6213 gnd.n6212 585
R83 gnd.n6212 gnd.n6211 585
R84 gnd.n707 gnd.n706 585
R85 gnd.n6210 gnd.n707 585
R86 gnd.n6208 gnd.n6207 585
R87 gnd.n6209 gnd.n6208 585
R88 gnd.n6206 gnd.n709 585
R89 gnd.n709 gnd.n708 585
R90 gnd.n6205 gnd.n6204 585
R91 gnd.n6204 gnd.n6203 585
R92 gnd.n715 gnd.n714 585
R93 gnd.n6202 gnd.n715 585
R94 gnd.n6200 gnd.n6199 585
R95 gnd.n6201 gnd.n6200 585
R96 gnd.n6198 gnd.n717 585
R97 gnd.n717 gnd.n716 585
R98 gnd.n6197 gnd.n6196 585
R99 gnd.n6196 gnd.n6195 585
R100 gnd.n723 gnd.n722 585
R101 gnd.n6194 gnd.n723 585
R102 gnd.n6192 gnd.n6191 585
R103 gnd.n6193 gnd.n6192 585
R104 gnd.n6190 gnd.n725 585
R105 gnd.n725 gnd.n724 585
R106 gnd.n6189 gnd.n6188 585
R107 gnd.n6188 gnd.n6187 585
R108 gnd.n731 gnd.n730 585
R109 gnd.n6186 gnd.n731 585
R110 gnd.n6184 gnd.n6183 585
R111 gnd.n6185 gnd.n6184 585
R112 gnd.n6182 gnd.n733 585
R113 gnd.n733 gnd.n732 585
R114 gnd.n6181 gnd.n6180 585
R115 gnd.n6180 gnd.n6179 585
R116 gnd.n739 gnd.n738 585
R117 gnd.n6178 gnd.n739 585
R118 gnd.n6176 gnd.n6175 585
R119 gnd.n6177 gnd.n6176 585
R120 gnd.n6174 gnd.n741 585
R121 gnd.n741 gnd.n740 585
R122 gnd.n6173 gnd.n6172 585
R123 gnd.n6172 gnd.n6171 585
R124 gnd.n747 gnd.n746 585
R125 gnd.n6170 gnd.n747 585
R126 gnd.n6168 gnd.n6167 585
R127 gnd.n6169 gnd.n6168 585
R128 gnd.n6166 gnd.n749 585
R129 gnd.n749 gnd.n748 585
R130 gnd.n6165 gnd.n6164 585
R131 gnd.n6164 gnd.n6163 585
R132 gnd.n755 gnd.n754 585
R133 gnd.n6162 gnd.n755 585
R134 gnd.n6160 gnd.n6159 585
R135 gnd.n6161 gnd.n6160 585
R136 gnd.n6158 gnd.n757 585
R137 gnd.n757 gnd.n756 585
R138 gnd.n6157 gnd.n6156 585
R139 gnd.n6156 gnd.n6155 585
R140 gnd.n763 gnd.n762 585
R141 gnd.n6154 gnd.n763 585
R142 gnd.n6152 gnd.n6151 585
R143 gnd.n6153 gnd.n6152 585
R144 gnd.n6150 gnd.n765 585
R145 gnd.n765 gnd.n764 585
R146 gnd.n6149 gnd.n6148 585
R147 gnd.n6148 gnd.n6147 585
R148 gnd.n771 gnd.n770 585
R149 gnd.n6146 gnd.n771 585
R150 gnd.n6144 gnd.n6143 585
R151 gnd.n6145 gnd.n6144 585
R152 gnd.n6142 gnd.n773 585
R153 gnd.n773 gnd.n772 585
R154 gnd.n6141 gnd.n6140 585
R155 gnd.n6140 gnd.n6139 585
R156 gnd.n779 gnd.n778 585
R157 gnd.n6138 gnd.n779 585
R158 gnd.n6136 gnd.n6135 585
R159 gnd.n6137 gnd.n6136 585
R160 gnd.n6134 gnd.n781 585
R161 gnd.n781 gnd.n780 585
R162 gnd.n6133 gnd.n6132 585
R163 gnd.n6132 gnd.n6131 585
R164 gnd.n787 gnd.n786 585
R165 gnd.n6130 gnd.n787 585
R166 gnd.n6128 gnd.n6127 585
R167 gnd.n6129 gnd.n6128 585
R168 gnd.n6126 gnd.n789 585
R169 gnd.n789 gnd.n788 585
R170 gnd.n6125 gnd.n6124 585
R171 gnd.n6124 gnd.n6123 585
R172 gnd.n795 gnd.n794 585
R173 gnd.n6122 gnd.n795 585
R174 gnd.n6120 gnd.n6119 585
R175 gnd.n6121 gnd.n6120 585
R176 gnd.n6118 gnd.n797 585
R177 gnd.n797 gnd.n796 585
R178 gnd.n6117 gnd.n6116 585
R179 gnd.n6116 gnd.n6115 585
R180 gnd.n803 gnd.n802 585
R181 gnd.n6114 gnd.n803 585
R182 gnd.n6112 gnd.n6111 585
R183 gnd.n6113 gnd.n6112 585
R184 gnd.n6110 gnd.n805 585
R185 gnd.n805 gnd.n804 585
R186 gnd.n6109 gnd.n6108 585
R187 gnd.n6108 gnd.n6107 585
R188 gnd.n811 gnd.n810 585
R189 gnd.n6106 gnd.n811 585
R190 gnd.n6104 gnd.n6103 585
R191 gnd.n6105 gnd.n6104 585
R192 gnd.n6102 gnd.n813 585
R193 gnd.n813 gnd.n812 585
R194 gnd.n6101 gnd.n6100 585
R195 gnd.n6100 gnd.n6099 585
R196 gnd.n819 gnd.n818 585
R197 gnd.n6098 gnd.n819 585
R198 gnd.n6096 gnd.n6095 585
R199 gnd.n6097 gnd.n6096 585
R200 gnd.n6094 gnd.n821 585
R201 gnd.n821 gnd.n820 585
R202 gnd.n657 gnd.n656 585
R203 gnd.n656 gnd.n655 585
R204 gnd.n6266 gnd.n6265 585
R205 gnd.n6267 gnd.n6266 585
R206 gnd.n654 gnd.n653 585
R207 gnd.n6268 gnd.n654 585
R208 gnd.n6271 gnd.n6270 585
R209 gnd.n6270 gnd.n6269 585
R210 gnd.n651 gnd.n650 585
R211 gnd.n650 gnd.n649 585
R212 gnd.n6276 gnd.n6275 585
R213 gnd.n6277 gnd.n6276 585
R214 gnd.n648 gnd.n647 585
R215 gnd.n6278 gnd.n648 585
R216 gnd.n6281 gnd.n6280 585
R217 gnd.n6280 gnd.n6279 585
R218 gnd.n645 gnd.n644 585
R219 gnd.n644 gnd.n643 585
R220 gnd.n6286 gnd.n6285 585
R221 gnd.n6287 gnd.n6286 585
R222 gnd.n642 gnd.n641 585
R223 gnd.n6288 gnd.n642 585
R224 gnd.n6291 gnd.n6290 585
R225 gnd.n6290 gnd.n6289 585
R226 gnd.n639 gnd.n638 585
R227 gnd.n638 gnd.n637 585
R228 gnd.n6296 gnd.n6295 585
R229 gnd.n6297 gnd.n6296 585
R230 gnd.n636 gnd.n635 585
R231 gnd.n6298 gnd.n636 585
R232 gnd.n6301 gnd.n6300 585
R233 gnd.n6300 gnd.n6299 585
R234 gnd.n633 gnd.n632 585
R235 gnd.n632 gnd.n631 585
R236 gnd.n6306 gnd.n6305 585
R237 gnd.n6307 gnd.n6306 585
R238 gnd.n630 gnd.n629 585
R239 gnd.n6308 gnd.n630 585
R240 gnd.n6311 gnd.n6310 585
R241 gnd.n6310 gnd.n6309 585
R242 gnd.n627 gnd.n626 585
R243 gnd.n626 gnd.n625 585
R244 gnd.n6316 gnd.n6315 585
R245 gnd.n6317 gnd.n6316 585
R246 gnd.n624 gnd.n623 585
R247 gnd.n6318 gnd.n624 585
R248 gnd.n6321 gnd.n6320 585
R249 gnd.n6320 gnd.n6319 585
R250 gnd.n621 gnd.n620 585
R251 gnd.n620 gnd.n619 585
R252 gnd.n6326 gnd.n6325 585
R253 gnd.n6327 gnd.n6326 585
R254 gnd.n618 gnd.n617 585
R255 gnd.n6328 gnd.n618 585
R256 gnd.n6331 gnd.n6330 585
R257 gnd.n6330 gnd.n6329 585
R258 gnd.n615 gnd.n614 585
R259 gnd.n614 gnd.n613 585
R260 gnd.n6336 gnd.n6335 585
R261 gnd.n6337 gnd.n6336 585
R262 gnd.n612 gnd.n611 585
R263 gnd.n6338 gnd.n612 585
R264 gnd.n6341 gnd.n6340 585
R265 gnd.n6340 gnd.n6339 585
R266 gnd.n609 gnd.n608 585
R267 gnd.n608 gnd.n607 585
R268 gnd.n6346 gnd.n6345 585
R269 gnd.n6347 gnd.n6346 585
R270 gnd.n606 gnd.n605 585
R271 gnd.n6348 gnd.n606 585
R272 gnd.n6351 gnd.n6350 585
R273 gnd.n6350 gnd.n6349 585
R274 gnd.n603 gnd.n602 585
R275 gnd.n602 gnd.n601 585
R276 gnd.n6356 gnd.n6355 585
R277 gnd.n6357 gnd.n6356 585
R278 gnd.n600 gnd.n599 585
R279 gnd.n6358 gnd.n600 585
R280 gnd.n6361 gnd.n6360 585
R281 gnd.n6360 gnd.n6359 585
R282 gnd.n597 gnd.n596 585
R283 gnd.n596 gnd.n595 585
R284 gnd.n6366 gnd.n6365 585
R285 gnd.n6367 gnd.n6366 585
R286 gnd.n594 gnd.n593 585
R287 gnd.n6368 gnd.n594 585
R288 gnd.n6371 gnd.n6370 585
R289 gnd.n6370 gnd.n6369 585
R290 gnd.n591 gnd.n590 585
R291 gnd.n590 gnd.n589 585
R292 gnd.n6376 gnd.n6375 585
R293 gnd.n6377 gnd.n6376 585
R294 gnd.n588 gnd.n587 585
R295 gnd.n6378 gnd.n588 585
R296 gnd.n6381 gnd.n6380 585
R297 gnd.n6380 gnd.n6379 585
R298 gnd.n585 gnd.n584 585
R299 gnd.n584 gnd.n583 585
R300 gnd.n6386 gnd.n6385 585
R301 gnd.n6387 gnd.n6386 585
R302 gnd.n582 gnd.n581 585
R303 gnd.n6388 gnd.n582 585
R304 gnd.n6391 gnd.n6390 585
R305 gnd.n6390 gnd.n6389 585
R306 gnd.n579 gnd.n578 585
R307 gnd.n578 gnd.n577 585
R308 gnd.n6396 gnd.n6395 585
R309 gnd.n6397 gnd.n6396 585
R310 gnd.n576 gnd.n575 585
R311 gnd.n6398 gnd.n576 585
R312 gnd.n6401 gnd.n6400 585
R313 gnd.n6400 gnd.n6399 585
R314 gnd.n573 gnd.n572 585
R315 gnd.n572 gnd.n571 585
R316 gnd.n6406 gnd.n6405 585
R317 gnd.n6407 gnd.n6406 585
R318 gnd.n570 gnd.n569 585
R319 gnd.n6408 gnd.n570 585
R320 gnd.n6411 gnd.n6410 585
R321 gnd.n6410 gnd.n6409 585
R322 gnd.n567 gnd.n566 585
R323 gnd.n566 gnd.n565 585
R324 gnd.n6416 gnd.n6415 585
R325 gnd.n6417 gnd.n6416 585
R326 gnd.n564 gnd.n563 585
R327 gnd.n6418 gnd.n564 585
R328 gnd.n6421 gnd.n6420 585
R329 gnd.n6420 gnd.n6419 585
R330 gnd.n561 gnd.n560 585
R331 gnd.n560 gnd.n559 585
R332 gnd.n6426 gnd.n6425 585
R333 gnd.n6427 gnd.n6426 585
R334 gnd.n558 gnd.n557 585
R335 gnd.n6428 gnd.n558 585
R336 gnd.n6431 gnd.n6430 585
R337 gnd.n6430 gnd.n6429 585
R338 gnd.n555 gnd.n554 585
R339 gnd.n554 gnd.n553 585
R340 gnd.n6436 gnd.n6435 585
R341 gnd.n6437 gnd.n6436 585
R342 gnd.n552 gnd.n551 585
R343 gnd.n6438 gnd.n552 585
R344 gnd.n6441 gnd.n6440 585
R345 gnd.n6440 gnd.n6439 585
R346 gnd.n549 gnd.n548 585
R347 gnd.n548 gnd.n547 585
R348 gnd.n6446 gnd.n6445 585
R349 gnd.n6447 gnd.n6446 585
R350 gnd.n546 gnd.n545 585
R351 gnd.n6448 gnd.n546 585
R352 gnd.n6451 gnd.n6450 585
R353 gnd.n6450 gnd.n6449 585
R354 gnd.n543 gnd.n542 585
R355 gnd.n542 gnd.n541 585
R356 gnd.n6456 gnd.n6455 585
R357 gnd.n6457 gnd.n6456 585
R358 gnd.n540 gnd.n539 585
R359 gnd.n6458 gnd.n540 585
R360 gnd.n6461 gnd.n6460 585
R361 gnd.n6460 gnd.n6459 585
R362 gnd.n537 gnd.n536 585
R363 gnd.n536 gnd.n535 585
R364 gnd.n6466 gnd.n6465 585
R365 gnd.n6467 gnd.n6466 585
R366 gnd.n534 gnd.n533 585
R367 gnd.n6468 gnd.n534 585
R368 gnd.n6471 gnd.n6470 585
R369 gnd.n6470 gnd.n6469 585
R370 gnd.n531 gnd.n530 585
R371 gnd.n530 gnd.n529 585
R372 gnd.n6476 gnd.n6475 585
R373 gnd.n6477 gnd.n6476 585
R374 gnd.n528 gnd.n527 585
R375 gnd.n6478 gnd.n528 585
R376 gnd.n6481 gnd.n6480 585
R377 gnd.n6480 gnd.n6479 585
R378 gnd.n525 gnd.n524 585
R379 gnd.n524 gnd.n523 585
R380 gnd.n6486 gnd.n6485 585
R381 gnd.n6487 gnd.n6486 585
R382 gnd.n522 gnd.n521 585
R383 gnd.n6488 gnd.n522 585
R384 gnd.n6491 gnd.n6490 585
R385 gnd.n6490 gnd.n6489 585
R386 gnd.n519 gnd.n518 585
R387 gnd.n518 gnd.n517 585
R388 gnd.n6496 gnd.n6495 585
R389 gnd.n6497 gnd.n6496 585
R390 gnd.n516 gnd.n515 585
R391 gnd.n6498 gnd.n516 585
R392 gnd.n6501 gnd.n6500 585
R393 gnd.n6500 gnd.n6499 585
R394 gnd.n513 gnd.n512 585
R395 gnd.n512 gnd.n511 585
R396 gnd.n6506 gnd.n6505 585
R397 gnd.n6507 gnd.n6506 585
R398 gnd.n510 gnd.n509 585
R399 gnd.n6508 gnd.n510 585
R400 gnd.n6511 gnd.n6510 585
R401 gnd.n6510 gnd.n6509 585
R402 gnd.n507 gnd.n506 585
R403 gnd.n506 gnd.n505 585
R404 gnd.n6516 gnd.n6515 585
R405 gnd.n6517 gnd.n6516 585
R406 gnd.n504 gnd.n503 585
R407 gnd.n6518 gnd.n504 585
R408 gnd.n6521 gnd.n6520 585
R409 gnd.n6520 gnd.n6519 585
R410 gnd.n501 gnd.n500 585
R411 gnd.n500 gnd.n499 585
R412 gnd.n6526 gnd.n6525 585
R413 gnd.n6527 gnd.n6526 585
R414 gnd.n498 gnd.n497 585
R415 gnd.n6528 gnd.n498 585
R416 gnd.n6531 gnd.n6530 585
R417 gnd.n6530 gnd.n6529 585
R418 gnd.n495 gnd.n494 585
R419 gnd.n494 gnd.n493 585
R420 gnd.n6536 gnd.n6535 585
R421 gnd.n6537 gnd.n6536 585
R422 gnd.n492 gnd.n491 585
R423 gnd.n6538 gnd.n492 585
R424 gnd.n6541 gnd.n6540 585
R425 gnd.n6540 gnd.n6539 585
R426 gnd.n489 gnd.n488 585
R427 gnd.n488 gnd.n487 585
R428 gnd.n6546 gnd.n6545 585
R429 gnd.n6547 gnd.n6546 585
R430 gnd.n486 gnd.n485 585
R431 gnd.n6548 gnd.n486 585
R432 gnd.n6551 gnd.n6550 585
R433 gnd.n6550 gnd.n6549 585
R434 gnd.n483 gnd.n482 585
R435 gnd.n482 gnd.n481 585
R436 gnd.n6556 gnd.n6555 585
R437 gnd.n6557 gnd.n6556 585
R438 gnd.n480 gnd.n479 585
R439 gnd.n6558 gnd.n480 585
R440 gnd.n6561 gnd.n6560 585
R441 gnd.n6560 gnd.n6559 585
R442 gnd.n477 gnd.n476 585
R443 gnd.n476 gnd.n475 585
R444 gnd.n6566 gnd.n6565 585
R445 gnd.n6567 gnd.n6566 585
R446 gnd.n474 gnd.n473 585
R447 gnd.n6568 gnd.n474 585
R448 gnd.n6571 gnd.n6570 585
R449 gnd.n6570 gnd.n6569 585
R450 gnd.n471 gnd.n470 585
R451 gnd.n470 gnd.n469 585
R452 gnd.n6576 gnd.n6575 585
R453 gnd.n6577 gnd.n6576 585
R454 gnd.n468 gnd.n467 585
R455 gnd.n6578 gnd.n468 585
R456 gnd.n6581 gnd.n6580 585
R457 gnd.n6580 gnd.n6579 585
R458 gnd.n465 gnd.n464 585
R459 gnd.n464 gnd.n463 585
R460 gnd.n6586 gnd.n6585 585
R461 gnd.n6587 gnd.n6586 585
R462 gnd.n462 gnd.n461 585
R463 gnd.n6588 gnd.n462 585
R464 gnd.n6591 gnd.n6590 585
R465 gnd.n6590 gnd.n6589 585
R466 gnd.n459 gnd.n458 585
R467 gnd.n458 gnd.n457 585
R468 gnd.n6596 gnd.n6595 585
R469 gnd.n6597 gnd.n6596 585
R470 gnd.n456 gnd.n455 585
R471 gnd.n6598 gnd.n456 585
R472 gnd.n6601 gnd.n6600 585
R473 gnd.n6600 gnd.n6599 585
R474 gnd.n453 gnd.n452 585
R475 gnd.n452 gnd.n451 585
R476 gnd.n6606 gnd.n6605 585
R477 gnd.n6607 gnd.n6606 585
R478 gnd.n450 gnd.n449 585
R479 gnd.n6608 gnd.n450 585
R480 gnd.n6611 gnd.n6610 585
R481 gnd.n6610 gnd.n6609 585
R482 gnd.n447 gnd.n446 585
R483 gnd.n446 gnd.n445 585
R484 gnd.n6616 gnd.n6615 585
R485 gnd.n6617 gnd.n6616 585
R486 gnd.n444 gnd.n443 585
R487 gnd.n6618 gnd.n444 585
R488 gnd.n6621 gnd.n6620 585
R489 gnd.n6620 gnd.n6619 585
R490 gnd.n441 gnd.n440 585
R491 gnd.n440 gnd.n439 585
R492 gnd.n6626 gnd.n6625 585
R493 gnd.n6627 gnd.n6626 585
R494 gnd.n438 gnd.n437 585
R495 gnd.n6628 gnd.n438 585
R496 gnd.n6631 gnd.n6630 585
R497 gnd.n6630 gnd.n6629 585
R498 gnd.n435 gnd.n434 585
R499 gnd.n434 gnd.n433 585
R500 gnd.n6636 gnd.n6635 585
R501 gnd.n6637 gnd.n6636 585
R502 gnd.n432 gnd.n431 585
R503 gnd.n6638 gnd.n432 585
R504 gnd.n6641 gnd.n6640 585
R505 gnd.n6640 gnd.n6639 585
R506 gnd.n429 gnd.n428 585
R507 gnd.n428 gnd.n427 585
R508 gnd.n6646 gnd.n6645 585
R509 gnd.n6647 gnd.n6646 585
R510 gnd.n426 gnd.n425 585
R511 gnd.n6648 gnd.n426 585
R512 gnd.n6651 gnd.n6650 585
R513 gnd.n6650 gnd.n6649 585
R514 gnd.n423 gnd.n422 585
R515 gnd.n422 gnd.n421 585
R516 gnd.n6656 gnd.n6655 585
R517 gnd.n6657 gnd.n6656 585
R518 gnd.n420 gnd.n419 585
R519 gnd.n6658 gnd.n420 585
R520 gnd.n6661 gnd.n6660 585
R521 gnd.n6660 gnd.n6659 585
R522 gnd.n417 gnd.n416 585
R523 gnd.n416 gnd.n415 585
R524 gnd.n6666 gnd.n6665 585
R525 gnd.n6667 gnd.n6666 585
R526 gnd.n414 gnd.n413 585
R527 gnd.n6668 gnd.n414 585
R528 gnd.n6671 gnd.n6670 585
R529 gnd.n6670 gnd.n6669 585
R530 gnd.n411 gnd.n410 585
R531 gnd.n410 gnd.n409 585
R532 gnd.n6676 gnd.n6675 585
R533 gnd.n6677 gnd.n6676 585
R534 gnd.n408 gnd.n407 585
R535 gnd.n6678 gnd.n408 585
R536 gnd.n6681 gnd.n6680 585
R537 gnd.n6680 gnd.n6679 585
R538 gnd.n6892 gnd.n281 585
R539 gnd.n6892 gnd.n6891 585
R540 gnd.n6886 gnd.n282 585
R541 gnd.n6890 gnd.n282 585
R542 gnd.n6888 gnd.n6887 585
R543 gnd.n6889 gnd.n6888 585
R544 gnd.n285 gnd.n284 585
R545 gnd.n284 gnd.n283 585
R546 gnd.n6881 gnd.n6880 585
R547 gnd.n6880 gnd.n6879 585
R548 gnd.n288 gnd.n287 585
R549 gnd.n6878 gnd.n288 585
R550 gnd.n6876 gnd.n6875 585
R551 gnd.n6877 gnd.n6876 585
R552 gnd.n291 gnd.n290 585
R553 gnd.n290 gnd.n289 585
R554 gnd.n6871 gnd.n6870 585
R555 gnd.n6870 gnd.n6869 585
R556 gnd.n294 gnd.n293 585
R557 gnd.n6868 gnd.n294 585
R558 gnd.n6866 gnd.n6865 585
R559 gnd.n6867 gnd.n6866 585
R560 gnd.n297 gnd.n296 585
R561 gnd.n296 gnd.n295 585
R562 gnd.n6861 gnd.n6860 585
R563 gnd.n6860 gnd.n6859 585
R564 gnd.n300 gnd.n299 585
R565 gnd.n6858 gnd.n300 585
R566 gnd.n6856 gnd.n6855 585
R567 gnd.n6857 gnd.n6856 585
R568 gnd.n303 gnd.n302 585
R569 gnd.n302 gnd.n301 585
R570 gnd.n6851 gnd.n6850 585
R571 gnd.n6850 gnd.n6849 585
R572 gnd.n306 gnd.n305 585
R573 gnd.n6848 gnd.n306 585
R574 gnd.n6846 gnd.n6845 585
R575 gnd.n6847 gnd.n6846 585
R576 gnd.n309 gnd.n308 585
R577 gnd.n308 gnd.n307 585
R578 gnd.n6841 gnd.n6840 585
R579 gnd.n6840 gnd.n6839 585
R580 gnd.n312 gnd.n311 585
R581 gnd.n6838 gnd.n312 585
R582 gnd.n6836 gnd.n6835 585
R583 gnd.n6837 gnd.n6836 585
R584 gnd.n315 gnd.n314 585
R585 gnd.n314 gnd.n313 585
R586 gnd.n6831 gnd.n6830 585
R587 gnd.n6830 gnd.n6829 585
R588 gnd.n318 gnd.n317 585
R589 gnd.n6828 gnd.n318 585
R590 gnd.n6826 gnd.n6825 585
R591 gnd.n6827 gnd.n6826 585
R592 gnd.n321 gnd.n320 585
R593 gnd.n320 gnd.n319 585
R594 gnd.n6821 gnd.n6820 585
R595 gnd.n6820 gnd.n6819 585
R596 gnd.n324 gnd.n323 585
R597 gnd.n6818 gnd.n324 585
R598 gnd.n6816 gnd.n6815 585
R599 gnd.n6817 gnd.n6816 585
R600 gnd.n327 gnd.n326 585
R601 gnd.n326 gnd.n325 585
R602 gnd.n6811 gnd.n6810 585
R603 gnd.n6810 gnd.n6809 585
R604 gnd.n330 gnd.n329 585
R605 gnd.n6808 gnd.n330 585
R606 gnd.n6806 gnd.n6805 585
R607 gnd.n6807 gnd.n6806 585
R608 gnd.n333 gnd.n332 585
R609 gnd.n332 gnd.n331 585
R610 gnd.n6801 gnd.n6800 585
R611 gnd.n6800 gnd.n6799 585
R612 gnd.n336 gnd.n335 585
R613 gnd.n6798 gnd.n336 585
R614 gnd.n6796 gnd.n6795 585
R615 gnd.n6797 gnd.n6796 585
R616 gnd.n339 gnd.n338 585
R617 gnd.n338 gnd.n337 585
R618 gnd.n6791 gnd.n6790 585
R619 gnd.n6790 gnd.n6789 585
R620 gnd.n342 gnd.n341 585
R621 gnd.n6788 gnd.n342 585
R622 gnd.n6786 gnd.n6785 585
R623 gnd.n6787 gnd.n6786 585
R624 gnd.n345 gnd.n344 585
R625 gnd.n344 gnd.n343 585
R626 gnd.n6781 gnd.n6780 585
R627 gnd.n6780 gnd.n6779 585
R628 gnd.n348 gnd.n347 585
R629 gnd.n6778 gnd.n348 585
R630 gnd.n6776 gnd.n6775 585
R631 gnd.n6777 gnd.n6776 585
R632 gnd.n351 gnd.n350 585
R633 gnd.n350 gnd.n349 585
R634 gnd.n6771 gnd.n6770 585
R635 gnd.n6770 gnd.n6769 585
R636 gnd.n354 gnd.n353 585
R637 gnd.n6768 gnd.n354 585
R638 gnd.n6766 gnd.n6765 585
R639 gnd.n6767 gnd.n6766 585
R640 gnd.n357 gnd.n356 585
R641 gnd.n356 gnd.n355 585
R642 gnd.n6761 gnd.n6760 585
R643 gnd.n6760 gnd.n6759 585
R644 gnd.n360 gnd.n359 585
R645 gnd.n6758 gnd.n360 585
R646 gnd.n6756 gnd.n6755 585
R647 gnd.n6757 gnd.n6756 585
R648 gnd.n363 gnd.n362 585
R649 gnd.n362 gnd.n361 585
R650 gnd.n6751 gnd.n6750 585
R651 gnd.n6750 gnd.n6749 585
R652 gnd.n366 gnd.n365 585
R653 gnd.n6748 gnd.n366 585
R654 gnd.n6746 gnd.n6745 585
R655 gnd.n6747 gnd.n6746 585
R656 gnd.n369 gnd.n368 585
R657 gnd.n368 gnd.n367 585
R658 gnd.n6741 gnd.n6740 585
R659 gnd.n6740 gnd.n6739 585
R660 gnd.n372 gnd.n371 585
R661 gnd.n6738 gnd.n372 585
R662 gnd.n6736 gnd.n6735 585
R663 gnd.n6737 gnd.n6736 585
R664 gnd.n375 gnd.n374 585
R665 gnd.n374 gnd.n373 585
R666 gnd.n6731 gnd.n6730 585
R667 gnd.n6730 gnd.n6729 585
R668 gnd.n378 gnd.n377 585
R669 gnd.n6728 gnd.n378 585
R670 gnd.n6726 gnd.n6725 585
R671 gnd.n6727 gnd.n6726 585
R672 gnd.n381 gnd.n380 585
R673 gnd.n380 gnd.n379 585
R674 gnd.n6721 gnd.n6720 585
R675 gnd.n6720 gnd.n6719 585
R676 gnd.n384 gnd.n383 585
R677 gnd.n6718 gnd.n384 585
R678 gnd.n6716 gnd.n6715 585
R679 gnd.n6717 gnd.n6716 585
R680 gnd.n387 gnd.n386 585
R681 gnd.n386 gnd.n385 585
R682 gnd.n6711 gnd.n6710 585
R683 gnd.n6710 gnd.n6709 585
R684 gnd.n390 gnd.n389 585
R685 gnd.n6708 gnd.n390 585
R686 gnd.n6706 gnd.n6705 585
R687 gnd.n6707 gnd.n6706 585
R688 gnd.n393 gnd.n392 585
R689 gnd.n392 gnd.n391 585
R690 gnd.n6701 gnd.n6700 585
R691 gnd.n6700 gnd.n6699 585
R692 gnd.n396 gnd.n395 585
R693 gnd.n6698 gnd.n396 585
R694 gnd.n6696 gnd.n6695 585
R695 gnd.n6697 gnd.n6696 585
R696 gnd.n399 gnd.n398 585
R697 gnd.n398 gnd.n397 585
R698 gnd.n6691 gnd.n6690 585
R699 gnd.n6690 gnd.n6689 585
R700 gnd.n402 gnd.n401 585
R701 gnd.n6688 gnd.n402 585
R702 gnd.n6686 gnd.n6685 585
R703 gnd.n6687 gnd.n6686 585
R704 gnd.n405 gnd.n404 585
R705 gnd.n404 gnd.n403 585
R706 gnd.n5997 gnd.n5996 585
R707 gnd.n5998 gnd.n5997 585
R708 gnd.n982 gnd.n981 585
R709 gnd.n4299 gnd.n982 585
R710 gnd.n6006 gnd.n6005 585
R711 gnd.n6005 gnd.n6004 585
R712 gnd.n6007 gnd.n976 585
R713 gnd.n4061 gnd.n976 585
R714 gnd.n6009 gnd.n6008 585
R715 gnd.n6010 gnd.n6009 585
R716 gnd.n961 gnd.n960 585
R717 gnd.n4052 gnd.n961 585
R718 gnd.n6018 gnd.n6017 585
R719 gnd.n6017 gnd.n6016 585
R720 gnd.n6019 gnd.n955 585
R721 gnd.n4048 gnd.n955 585
R722 gnd.n6021 gnd.n6020 585
R723 gnd.n6022 gnd.n6021 585
R724 gnd.n939 gnd.n938 585
R725 gnd.n4041 gnd.n939 585
R726 gnd.n6030 gnd.n6029 585
R727 gnd.n6029 gnd.n6028 585
R728 gnd.n6031 gnd.n933 585
R729 gnd.n4078 gnd.n933 585
R730 gnd.n6033 gnd.n6032 585
R731 gnd.n6034 gnd.n6033 585
R732 gnd.n920 gnd.n919 585
R733 gnd.n4033 gnd.n920 585
R734 gnd.n6042 gnd.n6041 585
R735 gnd.n6041 gnd.n6040 585
R736 gnd.n6043 gnd.n914 585
R737 gnd.n4025 gnd.n914 585
R738 gnd.n6045 gnd.n6044 585
R739 gnd.n6046 gnd.n6045 585
R740 gnd.n915 gnd.n913 585
R741 gnd.n4012 gnd.n913 585
R742 gnd.n3994 gnd.n3993 585
R743 gnd.n3993 gnd.n2070 585
R744 gnd.n3995 gnd.n2080 585
R745 gnd.n4004 gnd.n2080 585
R746 gnd.n3997 gnd.n3996 585
R747 gnd.n3998 gnd.n3997 585
R748 gnd.n2087 gnd.n2086 585
R749 gnd.n3984 gnd.n2086 585
R750 gnd.n3972 gnd.n3971 585
R751 gnd.n3973 gnd.n3972 585
R752 gnd.n3970 gnd.n3966 585
R753 gnd.n3976 gnd.n3966 585
R754 gnd.n893 gnd.n892 585
R755 gnd.n3949 gnd.n893 585
R756 gnd.n6056 gnd.n6055 585
R757 gnd.n6055 gnd.n6054 585
R758 gnd.n6057 gnd.n887 585
R759 gnd.n3939 gnd.n887 585
R760 gnd.n6059 gnd.n6058 585
R761 gnd.n6060 gnd.n6059 585
R762 gnd.n872 gnd.n871 585
R763 gnd.n3929 gnd.n872 585
R764 gnd.n6068 gnd.n6067 585
R765 gnd.n6067 gnd.n6066 585
R766 gnd.n6069 gnd.n866 585
R767 gnd.n3895 gnd.n866 585
R768 gnd.n6071 gnd.n6070 585
R769 gnd.n6072 gnd.n6071 585
R770 gnd.n851 gnd.n850 585
R771 gnd.n3901 gnd.n851 585
R772 gnd.n6080 gnd.n6079 585
R773 gnd.n6079 gnd.n6078 585
R774 gnd.n6081 gnd.n845 585
R775 gnd.n3881 gnd.n845 585
R776 gnd.n6083 gnd.n6082 585
R777 gnd.n6084 gnd.n6083 585
R778 gnd.n846 gnd.n844 585
R779 gnd.n844 gnd.n830 585
R780 gnd.n3850 gnd.n831 585
R781 gnd.n6090 gnd.n831 585
R782 gnd.n3852 gnd.n3851 585
R783 gnd.n3851 gnd.n827 585
R784 gnd.n3853 gnd.n2145 585
R785 gnd.n3868 gnd.n2145 585
R786 gnd.n2157 gnd.n2155 585
R787 gnd.n2155 gnd.n2143 585
R788 gnd.n3858 gnd.n3857 585
R789 gnd.n3859 gnd.n3858 585
R790 gnd.n2156 gnd.n2154 585
R791 gnd.n2154 gnd.n2151 585
R792 gnd.n3844 gnd.n3843 585
R793 gnd.n2160 gnd.n2159 585
R794 gnd.n3652 gnd.n3651 585
R795 gnd.n3654 gnd.n3653 585
R796 gnd.n3656 gnd.n3655 585
R797 gnd.n3660 gnd.n3648 585
R798 gnd.n3662 gnd.n3661 585
R799 gnd.n3664 gnd.n3663 585
R800 gnd.n3666 gnd.n3665 585
R801 gnd.n3670 gnd.n3646 585
R802 gnd.n3672 gnd.n3671 585
R803 gnd.n3674 gnd.n3673 585
R804 gnd.n3676 gnd.n3675 585
R805 gnd.n3680 gnd.n3644 585
R806 gnd.n3682 gnd.n3681 585
R807 gnd.n3684 gnd.n3683 585
R808 gnd.n3686 gnd.n3685 585
R809 gnd.n3642 gnd.n3638 585
R810 gnd.n3698 gnd.n3697 585
R811 gnd.n3841 gnd.n3698 585
R812 gnd.n4197 gnd.n4196 585
R813 gnd.n4194 gnd.n4188 585
R814 gnd.n4204 gnd.n4185 585
R815 gnd.n4205 gnd.n4183 585
R816 gnd.n4182 gnd.n4175 585
R817 gnd.n4212 gnd.n4174 585
R818 gnd.n4213 gnd.n4173 585
R819 gnd.n4171 gnd.n4163 585
R820 gnd.n4220 gnd.n4162 585
R821 gnd.n4221 gnd.n4160 585
R822 gnd.n4159 gnd.n4152 585
R823 gnd.n4228 gnd.n4151 585
R824 gnd.n4229 gnd.n4150 585
R825 gnd.n4148 gnd.n4141 585
R826 gnd.n4236 gnd.n4140 585
R827 gnd.n4237 gnd.n4138 585
R828 gnd.n4137 gnd.n4133 585
R829 gnd.n4135 gnd.n4134 585
R830 gnd.n999 gnd.n997 585
R831 gnd.n1961 gnd.n997 585
R832 gnd.n1997 gnd.n995 585
R833 gnd.n5998 gnd.n995 585
R834 gnd.n4298 gnd.n4297 585
R835 gnd.n4299 gnd.n4298 585
R836 gnd.n1996 gnd.n985 585
R837 gnd.n6004 gnd.n985 585
R838 gnd.n4064 gnd.n4062 585
R839 gnd.n4062 gnd.n4061 585
R840 gnd.n4065 gnd.n974 585
R841 gnd.n6010 gnd.n974 585
R842 gnd.n4066 gnd.n2053 585
R843 gnd.n4052 gnd.n2053 585
R844 gnd.n2051 gnd.n963 585
R845 gnd.n6016 gnd.n963 585
R846 gnd.n4070 gnd.n2050 585
R847 gnd.n4048 gnd.n2050 585
R848 gnd.n4071 gnd.n953 585
R849 gnd.n6022 gnd.n953 585
R850 gnd.n4072 gnd.n2049 585
R851 gnd.n4041 gnd.n2049 585
R852 gnd.n2046 gnd.n942 585
R853 gnd.n6028 gnd.n942 585
R854 gnd.n4077 gnd.n4076 585
R855 gnd.n4078 gnd.n4077 585
R856 gnd.n2045 gnd.n932 585
R857 gnd.n6034 gnd.n932 585
R858 gnd.n4032 gnd.n4031 585
R859 gnd.n4033 gnd.n4032 585
R860 gnd.n2061 gnd.n922 585
R861 gnd.n6040 gnd.n922 585
R862 gnd.n4027 gnd.n4026 585
R863 gnd.n4026 gnd.n4025 585
R864 gnd.n2063 gnd.n911 585
R865 gnd.n6046 gnd.n911 585
R866 gnd.n4011 gnd.n4010 585
R867 gnd.n4012 gnd.n4011 585
R868 gnd.n2073 gnd.n2072 585
R869 gnd.n2072 gnd.n2070 585
R870 gnd.n4006 gnd.n4005 585
R871 gnd.n4005 gnd.n4004 585
R872 gnd.n2076 gnd.n2075 585
R873 gnd.n3998 gnd.n2076 585
R874 gnd.n3983 gnd.n3982 585
R875 gnd.n3984 gnd.n3983 585
R876 gnd.n2107 gnd.n2106 585
R877 gnd.n3973 gnd.n2106 585
R878 gnd.n3978 gnd.n3977 585
R879 gnd.n3977 gnd.n3976 585
R880 gnd.n2110 gnd.n2109 585
R881 gnd.n3949 gnd.n2110 585
R882 gnd.n3936 gnd.n896 585
R883 gnd.n6054 gnd.n896 585
R884 gnd.n3938 gnd.n3937 585
R885 gnd.n3939 gnd.n3938 585
R886 gnd.n2120 gnd.n885 585
R887 gnd.n6060 gnd.n885 585
R888 gnd.n3931 gnd.n3930 585
R889 gnd.n3930 gnd.n3929 585
R890 gnd.n2122 gnd.n875 585
R891 gnd.n6066 gnd.n875 585
R892 gnd.n3897 gnd.n3896 585
R893 gnd.n3896 gnd.n3895 585
R894 gnd.n3898 gnd.n864 585
R895 gnd.n6072 gnd.n864 585
R896 gnd.n3900 gnd.n3899 585
R897 gnd.n3901 gnd.n3900 585
R898 gnd.n2130 gnd.n854 585
R899 gnd.n6078 gnd.n854 585
R900 gnd.n3880 gnd.n3879 585
R901 gnd.n3881 gnd.n3880 585
R902 gnd.n2138 gnd.n842 585
R903 gnd.n6084 gnd.n842 585
R904 gnd.n3874 gnd.n3873 585
R905 gnd.n3873 gnd.n830 585
R906 gnd.n3872 gnd.n829 585
R907 gnd.n6090 gnd.n829 585
R908 gnd.n3871 gnd.n3870 585
R909 gnd.n3870 gnd.n827 585
R910 gnd.n3869 gnd.n2140 585
R911 gnd.n3869 gnd.n3868 585
R912 gnd.n3692 gnd.n2142 585
R913 gnd.n2143 gnd.n2142 585
R914 gnd.n3693 gnd.n2153 585
R915 gnd.n3859 gnd.n2153 585
R916 gnd.n3694 gnd.n3639 585
R917 gnd.n3639 gnd.n2151 585
R918 gnd.n7054 gnd.n84 585
R919 gnd.n7150 gnd.n84 585
R920 gnd.n7055 gnd.n6986 585
R921 gnd.n6986 gnd.n81 585
R922 gnd.n7056 gnd.n162 585
R923 gnd.n7070 gnd.n162 585
R924 gnd.n173 gnd.n171 585
R925 gnd.n171 gnd.n161 585
R926 gnd.n7061 gnd.n7060 585
R927 gnd.n7062 gnd.n7061 585
R928 gnd.n172 gnd.n170 585
R929 gnd.n180 gnd.n170 585
R930 gnd.n6982 gnd.n6981 585
R931 gnd.n6981 gnd.n6980 585
R932 gnd.n176 gnd.n175 585
R933 gnd.n261 gnd.n176 585
R934 gnd.n6971 gnd.n6970 585
R935 gnd.n6972 gnd.n6971 585
R936 gnd.n190 gnd.n189 585
R937 gnd.n266 gnd.n189 585
R938 gnd.n6966 gnd.n6965 585
R939 gnd.n6965 gnd.n6964 585
R940 gnd.n193 gnd.n192 585
R941 gnd.n6907 gnd.n193 585
R942 gnd.n6955 gnd.n6954 585
R943 gnd.n6956 gnd.n6955 585
R944 gnd.n205 gnd.n204 585
R945 gnd.n6912 gnd.n204 585
R946 gnd.n6950 gnd.n6949 585
R947 gnd.n6949 gnd.n6948 585
R948 gnd.n208 gnd.n207 585
R949 gnd.n6916 gnd.n208 585
R950 gnd.n6939 gnd.n6938 585
R951 gnd.n6940 gnd.n6939 585
R952 gnd.n227 gnd.n226 585
R953 gnd.n6921 gnd.n226 585
R954 gnd.n6934 gnd.n6933 585
R955 gnd.n6933 gnd.n6932 585
R956 gnd.n230 gnd.n229 585
R957 gnd.n6927 gnd.n230 585
R958 gnd.n5813 gnd.n5811 585
R959 gnd.n5811 gnd.n5810 585
R960 gnd.n5814 gnd.n1169 585
R961 gnd.n1170 gnd.n1169 585
R962 gnd.n5815 gnd.n1168 585
R963 gnd.n5782 gnd.n1168 585
R964 gnd.n1175 gnd.n1166 585
R965 gnd.n1176 gnd.n1175 585
R966 gnd.n5819 gnd.n1165 585
R967 gnd.n5773 gnd.n1165 585
R968 gnd.n5820 gnd.n1164 585
R969 gnd.n5650 gnd.n1164 585
R970 gnd.n5821 gnd.n1163 585
R971 gnd.n5763 gnd.n1163 585
R972 gnd.n1204 gnd.n1161 585
R973 gnd.n1205 gnd.n1204 585
R974 gnd.n5825 gnd.n1160 585
R975 gnd.n5757 gnd.n1160 585
R976 gnd.n5826 gnd.n1159 585
R977 gnd.n5739 gnd.n1159 585
R978 gnd.n5827 gnd.n1158 585
R979 gnd.n1212 gnd.n1158 585
R980 gnd.n1223 gnd.n1156 585
R981 gnd.n5730 gnd.n1223 585
R982 gnd.n5831 gnd.n1155 585
R983 gnd.n1233 gnd.n1155 585
R984 gnd.n5832 gnd.n1154 585
R985 gnd.n5719 gnd.n1154 585
R986 gnd.n5833 gnd.n1153 585
R987 gnd.n5707 gnd.n1153 585
R988 gnd.n1240 gnd.n1151 585
R989 gnd.n1241 gnd.n1240 585
R990 gnd.n5837 gnd.n1150 585
R991 gnd.n5698 gnd.n1150 585
R992 gnd.n5838 gnd.n1149 585
R993 gnd.n5670 gnd.n1149 585
R994 gnd.n5839 gnd.n1148 585
R995 gnd.n5688 gnd.n1148 585
R996 gnd.n1145 gnd.n1143 585
R997 gnd.n5621 gnd.n1143 585
R998 gnd.n5844 gnd.n5843 585
R999 gnd.n5845 gnd.n5844 585
R1000 gnd.n1144 gnd.n1142 585
R1001 gnd.n5612 gnd.n1142 585
R1002 gnd.n5202 gnd.n1130 585
R1003 gnd.n5851 gnd.n1130 585
R1004 gnd.n5206 gnd.n5205 585
R1005 gnd.n5208 gnd.n5199 585
R1006 gnd.n5211 gnd.n5210 585
R1007 gnd.n5192 gnd.n5191 585
R1008 gnd.n5225 gnd.n5224 585
R1009 gnd.n5227 gnd.n5190 585
R1010 gnd.n5230 gnd.n5229 585
R1011 gnd.n5183 gnd.n5182 585
R1012 gnd.n5244 gnd.n5243 585
R1013 gnd.n5246 gnd.n5181 585
R1014 gnd.n5249 gnd.n5248 585
R1015 gnd.n5174 gnd.n5173 585
R1016 gnd.n5263 gnd.n5262 585
R1017 gnd.n5265 gnd.n5172 585
R1018 gnd.n5268 gnd.n5267 585
R1019 gnd.n5165 gnd.n5164 585
R1020 gnd.n5284 gnd.n5283 585
R1021 gnd.n5286 gnd.n5163 585
R1022 gnd.n5288 gnd.n5287 585
R1023 gnd.n5287 gnd.n1118 585
R1024 gnd.n7025 gnd.n80 585
R1025 gnd.n7026 gnd.n7024 585
R1026 gnd.n7027 gnd.n7020 585
R1027 gnd.n7018 gnd.n7016 585
R1028 gnd.n7031 gnd.n7015 585
R1029 gnd.n7032 gnd.n7013 585
R1030 gnd.n7033 gnd.n7012 585
R1031 gnd.n7010 gnd.n7008 585
R1032 gnd.n7037 gnd.n7007 585
R1033 gnd.n7038 gnd.n7005 585
R1034 gnd.n7039 gnd.n7004 585
R1035 gnd.n7002 gnd.n7000 585
R1036 gnd.n7043 gnd.n6999 585
R1037 gnd.n7044 gnd.n6997 585
R1038 gnd.n7045 gnd.n6996 585
R1039 gnd.n6994 gnd.n6992 585
R1040 gnd.n7049 gnd.n6991 585
R1041 gnd.n7050 gnd.n6989 585
R1042 gnd.n7051 gnd.n6988 585
R1043 gnd.n6988 gnd.n83 585
R1044 gnd.n7152 gnd.n7151 585
R1045 gnd.n7151 gnd.n7150 585
R1046 gnd.n79 gnd.n77 585
R1047 gnd.n81 gnd.n79 585
R1048 gnd.n7156 gnd.n76 585
R1049 gnd.n7070 gnd.n76 585
R1050 gnd.n7157 gnd.n75 585
R1051 gnd.n161 gnd.n75 585
R1052 gnd.n7158 gnd.n74 585
R1053 gnd.n7062 gnd.n74 585
R1054 gnd.n179 gnd.n72 585
R1055 gnd.n180 gnd.n179 585
R1056 gnd.n7162 gnd.n71 585
R1057 gnd.n6980 gnd.n71 585
R1058 gnd.n7163 gnd.n70 585
R1059 gnd.n261 gnd.n70 585
R1060 gnd.n7164 gnd.n69 585
R1061 gnd.n6972 gnd.n69 585
R1062 gnd.n265 gnd.n67 585
R1063 gnd.n266 gnd.n265 585
R1064 gnd.n7168 gnd.n66 585
R1065 gnd.n6964 gnd.n66 585
R1066 gnd.n7169 gnd.n65 585
R1067 gnd.n6907 gnd.n65 585
R1068 gnd.n7170 gnd.n64 585
R1069 gnd.n6956 gnd.n64 585
R1070 gnd.n6911 gnd.n62 585
R1071 gnd.n6912 gnd.n6911 585
R1072 gnd.n7174 gnd.n61 585
R1073 gnd.n6948 gnd.n61 585
R1074 gnd.n7175 gnd.n60 585
R1075 gnd.n6916 gnd.n60 585
R1076 gnd.n7176 gnd.n59 585
R1077 gnd.n6940 gnd.n59 585
R1078 gnd.n6920 gnd.n57 585
R1079 gnd.n6921 gnd.n6920 585
R1080 gnd.n7180 gnd.n56 585
R1081 gnd.n6932 gnd.n56 585
R1082 gnd.n7181 gnd.n55 585
R1083 gnd.n6927 gnd.n55 585
R1084 gnd.n7182 gnd.n54 585
R1085 gnd.n5810 gnd.n54 585
R1086 gnd.n1178 gnd.n52 585
R1087 gnd.n1178 gnd.n1170 585
R1088 gnd.n1189 gnd.n1179 585
R1089 gnd.n5782 gnd.n1179 585
R1090 gnd.n1190 gnd.n1187 585
R1091 gnd.n1187 gnd.n1176 585
R1092 gnd.n5771 gnd.n5770 585
R1093 gnd.n5773 gnd.n5771 585
R1094 gnd.n1188 gnd.n1186 585
R1095 gnd.n5650 gnd.n1186 585
R1096 gnd.n5765 gnd.n5764 585
R1097 gnd.n5764 gnd.n5763 585
R1098 gnd.n1193 gnd.n1192 585
R1099 gnd.n1205 gnd.n1193 585
R1100 gnd.n1216 gnd.n1203 585
R1101 gnd.n5757 gnd.n1203 585
R1102 gnd.n5738 gnd.n5737 585
R1103 gnd.n5739 gnd.n5738 585
R1104 gnd.n1215 gnd.n1214 585
R1105 gnd.n1214 gnd.n1212 585
R1106 gnd.n5732 gnd.n5731 585
R1107 gnd.n5731 gnd.n5730 585
R1108 gnd.n1219 gnd.n1218 585
R1109 gnd.n1233 gnd.n1219 585
R1110 gnd.n1245 gnd.n1232 585
R1111 gnd.n5719 gnd.n1232 585
R1112 gnd.n5706 gnd.n5705 585
R1113 gnd.n5707 gnd.n5706 585
R1114 gnd.n1244 gnd.n1243 585
R1115 gnd.n1243 gnd.n1241 585
R1116 gnd.n5700 gnd.n5699 585
R1117 gnd.n5699 gnd.n5698 585
R1118 gnd.n1248 gnd.n1247 585
R1119 gnd.n5670 gnd.n1248 585
R1120 gnd.n1263 gnd.n1258 585
R1121 gnd.n5688 gnd.n1258 585
R1122 gnd.n5620 gnd.n5619 585
R1123 gnd.n5621 gnd.n5620 585
R1124 gnd.n1262 gnd.n1140 585
R1125 gnd.n5845 gnd.n1140 585
R1126 gnd.n5614 gnd.n5613 585
R1127 gnd.n5613 gnd.n5612 585
R1128 gnd.n1265 gnd.n1128 585
R1129 gnd.n5851 gnd.n1128 585
R1130 gnd.n3519 gnd.n3518 585
R1131 gnd.n3520 gnd.n3519 585
R1132 gnd.n2237 gnd.n2236 585
R1133 gnd.n2243 gnd.n2236 585
R1134 gnd.n3494 gnd.n2255 585
R1135 gnd.n2255 gnd.n2242 585
R1136 gnd.n3496 gnd.n3495 585
R1137 gnd.n3497 gnd.n3496 585
R1138 gnd.n2256 gnd.n2254 585
R1139 gnd.n2254 gnd.n2250 585
R1140 gnd.n3228 gnd.n3227 585
R1141 gnd.n3227 gnd.n3226 585
R1142 gnd.n2261 gnd.n2260 585
R1143 gnd.n3197 gnd.n2261 585
R1144 gnd.n3217 gnd.n3216 585
R1145 gnd.n3216 gnd.n3215 585
R1146 gnd.n2268 gnd.n2267 585
R1147 gnd.n3203 gnd.n2268 585
R1148 gnd.n3173 gnd.n2288 585
R1149 gnd.n2288 gnd.n2287 585
R1150 gnd.n3175 gnd.n3174 585
R1151 gnd.n3176 gnd.n3175 585
R1152 gnd.n2289 gnd.n2286 585
R1153 gnd.n2297 gnd.n2286 585
R1154 gnd.n3151 gnd.n2309 585
R1155 gnd.n2309 gnd.n2296 585
R1156 gnd.n3153 gnd.n3152 585
R1157 gnd.n3154 gnd.n3153 585
R1158 gnd.n2310 gnd.n2308 585
R1159 gnd.n2308 gnd.n2304 585
R1160 gnd.n3139 gnd.n3138 585
R1161 gnd.n3138 gnd.n3137 585
R1162 gnd.n2315 gnd.n2314 585
R1163 gnd.n2325 gnd.n2315 585
R1164 gnd.n3127 gnd.n3126 585
R1165 gnd.n3126 gnd.n3125 585
R1166 gnd.n2322 gnd.n2321 585
R1167 gnd.n3113 gnd.n2322 585
R1168 gnd.n3087 gnd.n2343 585
R1169 gnd.n2343 gnd.n2332 585
R1170 gnd.n3089 gnd.n3088 585
R1171 gnd.n3090 gnd.n3089 585
R1172 gnd.n2344 gnd.n2342 585
R1173 gnd.n2352 gnd.n2342 585
R1174 gnd.n3065 gnd.n2364 585
R1175 gnd.n2364 gnd.n2351 585
R1176 gnd.n3067 gnd.n3066 585
R1177 gnd.n3068 gnd.n3067 585
R1178 gnd.n2365 gnd.n2363 585
R1179 gnd.n2363 gnd.n2359 585
R1180 gnd.n3053 gnd.n3052 585
R1181 gnd.n3052 gnd.n3051 585
R1182 gnd.n2370 gnd.n2369 585
R1183 gnd.n2379 gnd.n2370 585
R1184 gnd.n3042 gnd.n3041 585
R1185 gnd.n3041 gnd.n3040 585
R1186 gnd.n2377 gnd.n2376 585
R1187 gnd.n3028 gnd.n2377 585
R1188 gnd.n2466 gnd.n2465 585
R1189 gnd.n2466 gnd.n2386 585
R1190 gnd.n2985 gnd.n2984 585
R1191 gnd.n2984 gnd.n2983 585
R1192 gnd.n2986 gnd.n2460 585
R1193 gnd.n2471 gnd.n2460 585
R1194 gnd.n2988 gnd.n2987 585
R1195 gnd.n2989 gnd.n2988 585
R1196 gnd.n2461 gnd.n2459 585
R1197 gnd.n2484 gnd.n2459 585
R1198 gnd.n2444 gnd.n2443 585
R1199 gnd.n2447 gnd.n2444 585
R1200 gnd.n2999 gnd.n2998 585
R1201 gnd.n2998 gnd.n2997 585
R1202 gnd.n3000 gnd.n2438 585
R1203 gnd.n2959 gnd.n2438 585
R1204 gnd.n3002 gnd.n3001 585
R1205 gnd.n3003 gnd.n3002 585
R1206 gnd.n2439 gnd.n2437 585
R1207 gnd.n2498 gnd.n2437 585
R1208 gnd.n2951 gnd.n2950 585
R1209 gnd.n2950 gnd.n2949 585
R1210 gnd.n2495 gnd.n2494 585
R1211 gnd.n2933 gnd.n2495 585
R1212 gnd.n2920 gnd.n2514 585
R1213 gnd.n2514 gnd.n2513 585
R1214 gnd.n2922 gnd.n2921 585
R1215 gnd.n2923 gnd.n2922 585
R1216 gnd.n2515 gnd.n2512 585
R1217 gnd.n2521 gnd.n2512 585
R1218 gnd.n2901 gnd.n2900 585
R1219 gnd.n2902 gnd.n2901 585
R1220 gnd.n2532 gnd.n2531 585
R1221 gnd.n2531 gnd.n2527 585
R1222 gnd.n2891 gnd.n2890 585
R1223 gnd.n2892 gnd.n2891 585
R1224 gnd.n2542 gnd.n2541 585
R1225 gnd.n2547 gnd.n2541 585
R1226 gnd.n2869 gnd.n2560 585
R1227 gnd.n2560 gnd.n2546 585
R1228 gnd.n2871 gnd.n2870 585
R1229 gnd.n2872 gnd.n2871 585
R1230 gnd.n2561 gnd.n2559 585
R1231 gnd.n2559 gnd.n2555 585
R1232 gnd.n2860 gnd.n2859 585
R1233 gnd.n2861 gnd.n2860 585
R1234 gnd.n2568 gnd.n2567 585
R1235 gnd.n2572 gnd.n2567 585
R1236 gnd.n2837 gnd.n2589 585
R1237 gnd.n2589 gnd.n2571 585
R1238 gnd.n2839 gnd.n2838 585
R1239 gnd.n2840 gnd.n2839 585
R1240 gnd.n2590 gnd.n2588 585
R1241 gnd.n2588 gnd.n2579 585
R1242 gnd.n2832 gnd.n2831 585
R1243 gnd.n2831 gnd.n2830 585
R1244 gnd.n2637 gnd.n2636 585
R1245 gnd.n2638 gnd.n2637 585
R1246 gnd.n2791 gnd.n2790 585
R1247 gnd.n2792 gnd.n2791 585
R1248 gnd.n2647 gnd.n2646 585
R1249 gnd.n2646 gnd.n2645 585
R1250 gnd.n2786 gnd.n2785 585
R1251 gnd.n2785 gnd.n2784 585
R1252 gnd.n2650 gnd.n2649 585
R1253 gnd.n2651 gnd.n2650 585
R1254 gnd.n2775 gnd.n2774 585
R1255 gnd.n2776 gnd.n2775 585
R1256 gnd.n2658 gnd.n2657 585
R1257 gnd.n2767 gnd.n2657 585
R1258 gnd.n2770 gnd.n2769 585
R1259 gnd.n2769 gnd.n2768 585
R1260 gnd.n2661 gnd.n2660 585
R1261 gnd.n2662 gnd.n2661 585
R1262 gnd.n2756 gnd.n2755 585
R1263 gnd.n2754 gnd.n2680 585
R1264 gnd.n2753 gnd.n2679 585
R1265 gnd.n2758 gnd.n2679 585
R1266 gnd.n2752 gnd.n2751 585
R1267 gnd.n2750 gnd.n2749 585
R1268 gnd.n2748 gnd.n2747 585
R1269 gnd.n2746 gnd.n2745 585
R1270 gnd.n2744 gnd.n2743 585
R1271 gnd.n2742 gnd.n2741 585
R1272 gnd.n2740 gnd.n2739 585
R1273 gnd.n2738 gnd.n2737 585
R1274 gnd.n2736 gnd.n2735 585
R1275 gnd.n2734 gnd.n2733 585
R1276 gnd.n2732 gnd.n2731 585
R1277 gnd.n2730 gnd.n2729 585
R1278 gnd.n2728 gnd.n2727 585
R1279 gnd.n2726 gnd.n2725 585
R1280 gnd.n2724 gnd.n2723 585
R1281 gnd.n2722 gnd.n2721 585
R1282 gnd.n2720 gnd.n2719 585
R1283 gnd.n2718 gnd.n2717 585
R1284 gnd.n2716 gnd.n2715 585
R1285 gnd.n2714 gnd.n2713 585
R1286 gnd.n2712 gnd.n2711 585
R1287 gnd.n2710 gnd.n2709 585
R1288 gnd.n2667 gnd.n2666 585
R1289 gnd.n2761 gnd.n2760 585
R1290 gnd.n3523 gnd.n3522 585
R1291 gnd.n3525 gnd.n3524 585
R1292 gnd.n3527 gnd.n3526 585
R1293 gnd.n3529 gnd.n3528 585
R1294 gnd.n3531 gnd.n3530 585
R1295 gnd.n3533 gnd.n3532 585
R1296 gnd.n3535 gnd.n3534 585
R1297 gnd.n3537 gnd.n3536 585
R1298 gnd.n3539 gnd.n3538 585
R1299 gnd.n3541 gnd.n3540 585
R1300 gnd.n3543 gnd.n3542 585
R1301 gnd.n3545 gnd.n3544 585
R1302 gnd.n3547 gnd.n3546 585
R1303 gnd.n3549 gnd.n3548 585
R1304 gnd.n3551 gnd.n3550 585
R1305 gnd.n3553 gnd.n3552 585
R1306 gnd.n3555 gnd.n3554 585
R1307 gnd.n3557 gnd.n3556 585
R1308 gnd.n3559 gnd.n3558 585
R1309 gnd.n3561 gnd.n3560 585
R1310 gnd.n3563 gnd.n3562 585
R1311 gnd.n3565 gnd.n3564 585
R1312 gnd.n3567 gnd.n3566 585
R1313 gnd.n3569 gnd.n3568 585
R1314 gnd.n3571 gnd.n3570 585
R1315 gnd.n3572 gnd.n2204 585
R1316 gnd.n3573 gnd.n2162 585
R1317 gnd.n3611 gnd.n2162 585
R1318 gnd.n3521 gnd.n2234 585
R1319 gnd.n3521 gnd.n3520 585
R1320 gnd.n3190 gnd.n2233 585
R1321 gnd.n2243 gnd.n2233 585
R1322 gnd.n3192 gnd.n3191 585
R1323 gnd.n3191 gnd.n2242 585
R1324 gnd.n3193 gnd.n2252 585
R1325 gnd.n3497 gnd.n2252 585
R1326 gnd.n3195 gnd.n3194 585
R1327 gnd.n3194 gnd.n2250 585
R1328 gnd.n3196 gnd.n2263 585
R1329 gnd.n3226 gnd.n2263 585
R1330 gnd.n3199 gnd.n3198 585
R1331 gnd.n3198 gnd.n3197 585
R1332 gnd.n3200 gnd.n2270 585
R1333 gnd.n3215 gnd.n2270 585
R1334 gnd.n3202 gnd.n3201 585
R1335 gnd.n3203 gnd.n3202 585
R1336 gnd.n2280 gnd.n2279 585
R1337 gnd.n2287 gnd.n2279 585
R1338 gnd.n3178 gnd.n3177 585
R1339 gnd.n3177 gnd.n3176 585
R1340 gnd.n2283 gnd.n2282 585
R1341 gnd.n2297 gnd.n2283 585
R1342 gnd.n3103 gnd.n3102 585
R1343 gnd.n3102 gnd.n2296 585
R1344 gnd.n3104 gnd.n2306 585
R1345 gnd.n3154 gnd.n2306 585
R1346 gnd.n3106 gnd.n3105 585
R1347 gnd.n3105 gnd.n2304 585
R1348 gnd.n3107 gnd.n2317 585
R1349 gnd.n3137 gnd.n2317 585
R1350 gnd.n3109 gnd.n3108 585
R1351 gnd.n3108 gnd.n2325 585
R1352 gnd.n3110 gnd.n2324 585
R1353 gnd.n3125 gnd.n2324 585
R1354 gnd.n3112 gnd.n3111 585
R1355 gnd.n3113 gnd.n3112 585
R1356 gnd.n2336 gnd.n2335 585
R1357 gnd.n2335 gnd.n2332 585
R1358 gnd.n3092 gnd.n3091 585
R1359 gnd.n3091 gnd.n3090 585
R1360 gnd.n2339 gnd.n2338 585
R1361 gnd.n2352 gnd.n2339 585
R1362 gnd.n3016 gnd.n3015 585
R1363 gnd.n3015 gnd.n2351 585
R1364 gnd.n3017 gnd.n2361 585
R1365 gnd.n3068 gnd.n2361 585
R1366 gnd.n3019 gnd.n3018 585
R1367 gnd.n3018 gnd.n2359 585
R1368 gnd.n3020 gnd.n2372 585
R1369 gnd.n3051 gnd.n2372 585
R1370 gnd.n3022 gnd.n3021 585
R1371 gnd.n3021 gnd.n2379 585
R1372 gnd.n3023 gnd.n2378 585
R1373 gnd.n3040 gnd.n2378 585
R1374 gnd.n3025 gnd.n3024 585
R1375 gnd.n3028 gnd.n3025 585
R1376 gnd.n2389 gnd.n2388 585
R1377 gnd.n2388 gnd.n2386 585
R1378 gnd.n2468 gnd.n2467 585
R1379 gnd.n2983 gnd.n2467 585
R1380 gnd.n2470 gnd.n2469 585
R1381 gnd.n2471 gnd.n2470 585
R1382 gnd.n2481 gnd.n2457 585
R1383 gnd.n2989 gnd.n2457 585
R1384 gnd.n2483 gnd.n2482 585
R1385 gnd.n2484 gnd.n2483 585
R1386 gnd.n2480 gnd.n2479 585
R1387 gnd.n2480 gnd.n2447 585
R1388 gnd.n2478 gnd.n2445 585
R1389 gnd.n2997 gnd.n2445 585
R1390 gnd.n2434 gnd.n2432 585
R1391 gnd.n2959 gnd.n2434 585
R1392 gnd.n3005 gnd.n3004 585
R1393 gnd.n3004 gnd.n3003 585
R1394 gnd.n2433 gnd.n2431 585
R1395 gnd.n2498 gnd.n2433 585
R1396 gnd.n2930 gnd.n2497 585
R1397 gnd.n2949 gnd.n2497 585
R1398 gnd.n2932 gnd.n2931 585
R1399 gnd.n2933 gnd.n2932 585
R1400 gnd.n2507 gnd.n2506 585
R1401 gnd.n2513 gnd.n2506 585
R1402 gnd.n2925 gnd.n2924 585
R1403 gnd.n2924 gnd.n2923 585
R1404 gnd.n2510 gnd.n2509 585
R1405 gnd.n2521 gnd.n2510 585
R1406 gnd.n2810 gnd.n2529 585
R1407 gnd.n2902 gnd.n2529 585
R1408 gnd.n2812 gnd.n2811 585
R1409 gnd.n2811 gnd.n2527 585
R1410 gnd.n2813 gnd.n2540 585
R1411 gnd.n2892 gnd.n2540 585
R1412 gnd.n2815 gnd.n2814 585
R1413 gnd.n2815 gnd.n2547 585
R1414 gnd.n2817 gnd.n2816 585
R1415 gnd.n2816 gnd.n2546 585
R1416 gnd.n2818 gnd.n2557 585
R1417 gnd.n2872 gnd.n2557 585
R1418 gnd.n2820 gnd.n2819 585
R1419 gnd.n2819 gnd.n2555 585
R1420 gnd.n2821 gnd.n2566 585
R1421 gnd.n2861 gnd.n2566 585
R1422 gnd.n2823 gnd.n2822 585
R1423 gnd.n2823 gnd.n2572 585
R1424 gnd.n2825 gnd.n2824 585
R1425 gnd.n2824 gnd.n2571 585
R1426 gnd.n2826 gnd.n2587 585
R1427 gnd.n2840 gnd.n2587 585
R1428 gnd.n2827 gnd.n2640 585
R1429 gnd.n2640 gnd.n2579 585
R1430 gnd.n2829 gnd.n2828 585
R1431 gnd.n2830 gnd.n2829 585
R1432 gnd.n2641 gnd.n2639 585
R1433 gnd.n2639 gnd.n2638 585
R1434 gnd.n2794 gnd.n2793 585
R1435 gnd.n2793 gnd.n2792 585
R1436 gnd.n2644 gnd.n2643 585
R1437 gnd.n2645 gnd.n2644 585
R1438 gnd.n2783 gnd.n2782 585
R1439 gnd.n2784 gnd.n2783 585
R1440 gnd.n2653 gnd.n2652 585
R1441 gnd.n2652 gnd.n2651 585
R1442 gnd.n2778 gnd.n2777 585
R1443 gnd.n2777 gnd.n2776 585
R1444 gnd.n2656 gnd.n2655 585
R1445 gnd.n2767 gnd.n2656 585
R1446 gnd.n2766 gnd.n2765 585
R1447 gnd.n2768 gnd.n2766 585
R1448 gnd.n2664 gnd.n2663 585
R1449 gnd.n2663 gnd.n2662 585
R1450 gnd.n3506 gnd.n2184 585
R1451 gnd.n2184 gnd.n2161 585
R1452 gnd.n3507 gnd.n2245 585
R1453 gnd.n2245 gnd.n2235 585
R1454 gnd.n3509 gnd.n3508 585
R1455 gnd.n3510 gnd.n3509 585
R1456 gnd.n2246 gnd.n2244 585
R1457 gnd.n2253 gnd.n2244 585
R1458 gnd.n3500 gnd.n3499 585
R1459 gnd.n3499 gnd.n3498 585
R1460 gnd.n2249 gnd.n2248 585
R1461 gnd.n3225 gnd.n2249 585
R1462 gnd.n3211 gnd.n2272 585
R1463 gnd.n2272 gnd.n2262 585
R1464 gnd.n3213 gnd.n3212 585
R1465 gnd.n3214 gnd.n3213 585
R1466 gnd.n2273 gnd.n2271 585
R1467 gnd.n2271 gnd.n2269 585
R1468 gnd.n3206 gnd.n3205 585
R1469 gnd.n3205 gnd.n3204 585
R1470 gnd.n2276 gnd.n2275 585
R1471 gnd.n2285 gnd.n2276 585
R1472 gnd.n3162 gnd.n2299 585
R1473 gnd.n2299 gnd.n2284 585
R1474 gnd.n3164 gnd.n3163 585
R1475 gnd.n3165 gnd.n3164 585
R1476 gnd.n2300 gnd.n2298 585
R1477 gnd.n2307 gnd.n2298 585
R1478 gnd.n3157 gnd.n3156 585
R1479 gnd.n3156 gnd.n3155 585
R1480 gnd.n2303 gnd.n2302 585
R1481 gnd.n3136 gnd.n2303 585
R1482 gnd.n3121 gnd.n2327 585
R1483 gnd.n2327 gnd.n2316 585
R1484 gnd.n3123 gnd.n3122 585
R1485 gnd.n3124 gnd.n3123 585
R1486 gnd.n2328 gnd.n2326 585
R1487 gnd.n2326 gnd.n2323 585
R1488 gnd.n3116 gnd.n3115 585
R1489 gnd.n3115 gnd.n3114 585
R1490 gnd.n2331 gnd.n2330 585
R1491 gnd.n2341 gnd.n2331 585
R1492 gnd.n3076 gnd.n2354 585
R1493 gnd.n2354 gnd.n2340 585
R1494 gnd.n3078 gnd.n3077 585
R1495 gnd.n3079 gnd.n3078 585
R1496 gnd.n2355 gnd.n2353 585
R1497 gnd.n2362 gnd.n2353 585
R1498 gnd.n3071 gnd.n3070 585
R1499 gnd.n3070 gnd.n3069 585
R1500 gnd.n2358 gnd.n2357 585
R1501 gnd.n3050 gnd.n2358 585
R1502 gnd.n3036 gnd.n2381 585
R1503 gnd.n2381 gnd.n2371 585
R1504 gnd.n3038 gnd.n3037 585
R1505 gnd.n3039 gnd.n3038 585
R1506 gnd.n2382 gnd.n2380 585
R1507 gnd.n3027 gnd.n2380 585
R1508 gnd.n3031 gnd.n3030 585
R1509 gnd.n3030 gnd.n3029 585
R1510 gnd.n2385 gnd.n2384 585
R1511 gnd.n2982 gnd.n2385 585
R1512 gnd.n2475 gnd.n2474 585
R1513 gnd.n2476 gnd.n2475 585
R1514 gnd.n2455 gnd.n2454 585
R1515 gnd.n2458 gnd.n2455 585
R1516 gnd.n2992 gnd.n2991 585
R1517 gnd.n2991 gnd.n2990 585
R1518 gnd.n2993 gnd.n2449 585
R1519 gnd.n2485 gnd.n2449 585
R1520 gnd.n2995 gnd.n2994 585
R1521 gnd.n2996 gnd.n2995 585
R1522 gnd.n2450 gnd.n2448 585
R1523 gnd.n2960 gnd.n2448 585
R1524 gnd.n2944 gnd.n2943 585
R1525 gnd.n2943 gnd.n2436 585
R1526 gnd.n2945 gnd.n2500 585
R1527 gnd.n2500 gnd.n2435 585
R1528 gnd.n2947 gnd.n2946 585
R1529 gnd.n2948 gnd.n2947 585
R1530 gnd.n2501 gnd.n2499 585
R1531 gnd.n2499 gnd.n2496 585
R1532 gnd.n2936 gnd.n2935 585
R1533 gnd.n2935 gnd.n2934 585
R1534 gnd.n2504 gnd.n2503 585
R1535 gnd.n2511 gnd.n2504 585
R1536 gnd.n2910 gnd.n2909 585
R1537 gnd.n2911 gnd.n2910 585
R1538 gnd.n2523 gnd.n2522 585
R1539 gnd.n2530 gnd.n2522 585
R1540 gnd.n2905 gnd.n2904 585
R1541 gnd.n2904 gnd.n2903 585
R1542 gnd.n2526 gnd.n2525 585
R1543 gnd.n2893 gnd.n2526 585
R1544 gnd.n2880 gnd.n2550 585
R1545 gnd.n2550 gnd.n2549 585
R1546 gnd.n2882 gnd.n2881 585
R1547 gnd.n2883 gnd.n2882 585
R1548 gnd.n2551 gnd.n2548 585
R1549 gnd.n2558 gnd.n2548 585
R1550 gnd.n2875 gnd.n2874 585
R1551 gnd.n2874 gnd.n2873 585
R1552 gnd.n2554 gnd.n2553 585
R1553 gnd.n2862 gnd.n2554 585
R1554 gnd.n2849 gnd.n2575 585
R1555 gnd.n2575 gnd.n2574 585
R1556 gnd.n2851 gnd.n2850 585
R1557 gnd.n2852 gnd.n2851 585
R1558 gnd.n2845 gnd.n2573 585
R1559 gnd.n2844 gnd.n2843 585
R1560 gnd.n2578 gnd.n2577 585
R1561 gnd.n2841 gnd.n2578 585
R1562 gnd.n2600 gnd.n2599 585
R1563 gnd.n2603 gnd.n2602 585
R1564 gnd.n2601 gnd.n2596 585
R1565 gnd.n2608 gnd.n2607 585
R1566 gnd.n2610 gnd.n2609 585
R1567 gnd.n2613 gnd.n2612 585
R1568 gnd.n2611 gnd.n2594 585
R1569 gnd.n2618 gnd.n2617 585
R1570 gnd.n2620 gnd.n2619 585
R1571 gnd.n2623 gnd.n2622 585
R1572 gnd.n2621 gnd.n2592 585
R1573 gnd.n2628 gnd.n2627 585
R1574 gnd.n2632 gnd.n2629 585
R1575 gnd.n2633 gnd.n2570 585
R1576 gnd.n3512 gnd.n2199 585
R1577 gnd.n3579 gnd.n3578 585
R1578 gnd.n3581 gnd.n3580 585
R1579 gnd.n3583 gnd.n3582 585
R1580 gnd.n3585 gnd.n3584 585
R1581 gnd.n3587 gnd.n3586 585
R1582 gnd.n3589 gnd.n3588 585
R1583 gnd.n3591 gnd.n3590 585
R1584 gnd.n3593 gnd.n3592 585
R1585 gnd.n3595 gnd.n3594 585
R1586 gnd.n3597 gnd.n3596 585
R1587 gnd.n3599 gnd.n3598 585
R1588 gnd.n3601 gnd.n3600 585
R1589 gnd.n3604 gnd.n3603 585
R1590 gnd.n3602 gnd.n2187 585
R1591 gnd.n3608 gnd.n2185 585
R1592 gnd.n3610 gnd.n3609 585
R1593 gnd.n3611 gnd.n3610 585
R1594 gnd.n3513 gnd.n2240 585
R1595 gnd.n3513 gnd.n2161 585
R1596 gnd.n3515 gnd.n3514 585
R1597 gnd.n3514 gnd.n2235 585
R1598 gnd.n3511 gnd.n2239 585
R1599 gnd.n3511 gnd.n3510 585
R1600 gnd.n3490 gnd.n2241 585
R1601 gnd.n2253 gnd.n2241 585
R1602 gnd.n3489 gnd.n2251 585
R1603 gnd.n3498 gnd.n2251 585
R1604 gnd.n3224 gnd.n2258 585
R1605 gnd.n3225 gnd.n3224 585
R1606 gnd.n3223 gnd.n3222 585
R1607 gnd.n3223 gnd.n2262 585
R1608 gnd.n3221 gnd.n2264 585
R1609 gnd.n3214 gnd.n2264 585
R1610 gnd.n2277 gnd.n2265 585
R1611 gnd.n2277 gnd.n2269 585
R1612 gnd.n3170 gnd.n2278 585
R1613 gnd.n3204 gnd.n2278 585
R1614 gnd.n3169 gnd.n3168 585
R1615 gnd.n3168 gnd.n2285 585
R1616 gnd.n3167 gnd.n2293 585
R1617 gnd.n3167 gnd.n2284 585
R1618 gnd.n3166 gnd.n2295 585
R1619 gnd.n3166 gnd.n3165 585
R1620 gnd.n3145 gnd.n2294 585
R1621 gnd.n2307 gnd.n2294 585
R1622 gnd.n3144 gnd.n2305 585
R1623 gnd.n3155 gnd.n2305 585
R1624 gnd.n3134 gnd.n2312 585
R1625 gnd.n3136 gnd.n3134 585
R1626 gnd.n3133 gnd.n3132 585
R1627 gnd.n3133 gnd.n2316 585
R1628 gnd.n3131 gnd.n2318 585
R1629 gnd.n3124 gnd.n2318 585
R1630 gnd.n2333 gnd.n2319 585
R1631 gnd.n2333 gnd.n2323 585
R1632 gnd.n3084 gnd.n2334 585
R1633 gnd.n3114 gnd.n2334 585
R1634 gnd.n3083 gnd.n3082 585
R1635 gnd.n3082 gnd.n2341 585
R1636 gnd.n3081 gnd.n2348 585
R1637 gnd.n3081 gnd.n2340 585
R1638 gnd.n3080 gnd.n2350 585
R1639 gnd.n3080 gnd.n3079 585
R1640 gnd.n3059 gnd.n2349 585
R1641 gnd.n2362 gnd.n2349 585
R1642 gnd.n3058 gnd.n2360 585
R1643 gnd.n3069 gnd.n2360 585
R1644 gnd.n3049 gnd.n2367 585
R1645 gnd.n3050 gnd.n3049 585
R1646 gnd.n3048 gnd.n3047 585
R1647 gnd.n3048 gnd.n2371 585
R1648 gnd.n3046 gnd.n2373 585
R1649 gnd.n3039 gnd.n2373 585
R1650 gnd.n3026 gnd.n2374 585
R1651 gnd.n3027 gnd.n3026 585
R1652 gnd.n2979 gnd.n2387 585
R1653 gnd.n3029 gnd.n2387 585
R1654 gnd.n2981 gnd.n2980 585
R1655 gnd.n2982 gnd.n2981 585
R1656 gnd.n2974 gnd.n2477 585
R1657 gnd.n2477 gnd.n2476 585
R1658 gnd.n2972 gnd.n2971 585
R1659 gnd.n2971 gnd.n2458 585
R1660 gnd.n2969 gnd.n2456 585
R1661 gnd.n2990 gnd.n2456 585
R1662 gnd.n2487 gnd.n2486 585
R1663 gnd.n2486 gnd.n2485 585
R1664 gnd.n2963 gnd.n2446 585
R1665 gnd.n2996 gnd.n2446 585
R1666 gnd.n2962 gnd.n2961 585
R1667 gnd.n2961 gnd.n2960 585
R1668 gnd.n2958 gnd.n2489 585
R1669 gnd.n2958 gnd.n2436 585
R1670 gnd.n2957 gnd.n2956 585
R1671 gnd.n2957 gnd.n2435 585
R1672 gnd.n2492 gnd.n2491 585
R1673 gnd.n2948 gnd.n2491 585
R1674 gnd.n2916 gnd.n2915 585
R1675 gnd.n2915 gnd.n2496 585
R1676 gnd.n2917 gnd.n2505 585
R1677 gnd.n2934 gnd.n2505 585
R1678 gnd.n2914 gnd.n2913 585
R1679 gnd.n2913 gnd.n2511 585
R1680 gnd.n2912 gnd.n2519 585
R1681 gnd.n2912 gnd.n2911 585
R1682 gnd.n2897 gnd.n2520 585
R1683 gnd.n2530 gnd.n2520 585
R1684 gnd.n2896 gnd.n2528 585
R1685 gnd.n2903 gnd.n2528 585
R1686 gnd.n2895 gnd.n2894 585
R1687 gnd.n2894 gnd.n2893 585
R1688 gnd.n2539 gnd.n2536 585
R1689 gnd.n2549 gnd.n2539 585
R1690 gnd.n2885 gnd.n2884 585
R1691 gnd.n2884 gnd.n2883 585
R1692 gnd.n2545 gnd.n2544 585
R1693 gnd.n2558 gnd.n2545 585
R1694 gnd.n2865 gnd.n2556 585
R1695 gnd.n2873 gnd.n2556 585
R1696 gnd.n2864 gnd.n2863 585
R1697 gnd.n2863 gnd.n2862 585
R1698 gnd.n2565 gnd.n2563 585
R1699 gnd.n2574 gnd.n2565 585
R1700 gnd.n2854 gnd.n2853 585
R1701 gnd.n2853 gnd.n2852 585
R1702 gnd.n6000 gnd.n5999 585
R1703 gnd.n5999 gnd.n5998 585
R1704 gnd.n6001 gnd.n987 585
R1705 gnd.n4299 gnd.n987 585
R1706 gnd.n6003 gnd.n6002 585
R1707 gnd.n6004 gnd.n6003 585
R1708 gnd.n971 gnd.n970 585
R1709 gnd.n4061 gnd.n971 585
R1710 gnd.n6012 gnd.n6011 585
R1711 gnd.n6011 gnd.n6010 585
R1712 gnd.n6013 gnd.n965 585
R1713 gnd.n4052 gnd.n965 585
R1714 gnd.n6015 gnd.n6014 585
R1715 gnd.n6016 gnd.n6015 585
R1716 gnd.n950 gnd.n949 585
R1717 gnd.n4048 gnd.n950 585
R1718 gnd.n6024 gnd.n6023 585
R1719 gnd.n6023 gnd.n6022 585
R1720 gnd.n6025 gnd.n944 585
R1721 gnd.n4041 gnd.n944 585
R1722 gnd.n6027 gnd.n6026 585
R1723 gnd.n6028 gnd.n6027 585
R1724 gnd.n929 gnd.n928 585
R1725 gnd.n4078 gnd.n929 585
R1726 gnd.n6036 gnd.n6035 585
R1727 gnd.n6035 gnd.n6034 585
R1728 gnd.n6037 gnd.n924 585
R1729 gnd.n4033 gnd.n924 585
R1730 gnd.n6039 gnd.n6038 585
R1731 gnd.n6040 gnd.n6039 585
R1732 gnd.n908 gnd.n906 585
R1733 gnd.n4025 gnd.n908 585
R1734 gnd.n6048 gnd.n6047 585
R1735 gnd.n6047 gnd.n6046 585
R1736 gnd.n907 gnd.n905 585
R1737 gnd.n4012 gnd.n907 585
R1738 gnd.n4001 gnd.n4000 585
R1739 gnd.n4000 gnd.n2070 585
R1740 gnd.n4003 gnd.n4002 585
R1741 gnd.n4004 gnd.n4003 585
R1742 gnd.n3999 gnd.n2083 585
R1743 gnd.n3999 gnd.n3998 585
R1744 gnd.n2082 gnd.n2081 585
R1745 gnd.n3984 gnd.n2081 585
R1746 gnd.n3974 gnd.n3967 585
R1747 gnd.n3974 gnd.n3973 585
R1748 gnd.n3975 gnd.n899 585
R1749 gnd.n3976 gnd.n3975 585
R1750 gnd.n6051 gnd.n897 585
R1751 gnd.n3949 gnd.n897 585
R1752 gnd.n6053 gnd.n6052 585
R1753 gnd.n6054 gnd.n6053 585
R1754 gnd.n883 gnd.n882 585
R1755 gnd.n3939 gnd.n883 585
R1756 gnd.n6062 gnd.n6061 585
R1757 gnd.n6061 gnd.n6060 585
R1758 gnd.n6063 gnd.n877 585
R1759 gnd.n3929 gnd.n877 585
R1760 gnd.n6065 gnd.n6064 585
R1761 gnd.n6066 gnd.n6065 585
R1762 gnd.n861 gnd.n860 585
R1763 gnd.n3895 gnd.n861 585
R1764 gnd.n6074 gnd.n6073 585
R1765 gnd.n6073 gnd.n6072 585
R1766 gnd.n6075 gnd.n855 585
R1767 gnd.n3901 gnd.n855 585
R1768 gnd.n6077 gnd.n6076 585
R1769 gnd.n6078 gnd.n6077 585
R1770 gnd.n839 gnd.n838 585
R1771 gnd.n3881 gnd.n839 585
R1772 gnd.n6086 gnd.n6085 585
R1773 gnd.n6085 gnd.n6084 585
R1774 gnd.n6087 gnd.n833 585
R1775 gnd.n833 gnd.n830 585
R1776 gnd.n6089 gnd.n6088 585
R1777 gnd.n6090 gnd.n6089 585
R1778 gnd.n834 gnd.n832 585
R1779 gnd.n832 gnd.n827 585
R1780 gnd.n3867 gnd.n3866 585
R1781 gnd.n3868 gnd.n3867 585
R1782 gnd.n2147 gnd.n2146 585
R1783 gnd.n2146 gnd.n2143 585
R1784 gnd.n3861 gnd.n3860 585
R1785 gnd.n3860 gnd.n3859 585
R1786 gnd.n2150 gnd.n2149 585
R1787 gnd.n2151 gnd.n2150 585
R1788 gnd.n3839 gnd.n3838 585
R1789 gnd.n3837 gnd.n3700 585
R1790 gnd.n3836 gnd.n3699 585
R1791 gnd.n3841 gnd.n3699 585
R1792 gnd.n3835 gnd.n3834 585
R1793 gnd.n3833 gnd.n3832 585
R1794 gnd.n3831 gnd.n3830 585
R1795 gnd.n3829 gnd.n3828 585
R1796 gnd.n3827 gnd.n3826 585
R1797 gnd.n3825 gnd.n3824 585
R1798 gnd.n3823 gnd.n3822 585
R1799 gnd.n3821 gnd.n3820 585
R1800 gnd.n3819 gnd.n3818 585
R1801 gnd.n3817 gnd.n3816 585
R1802 gnd.n3815 gnd.n3814 585
R1803 gnd.n3813 gnd.n3812 585
R1804 gnd.n3811 gnd.n3810 585
R1805 gnd.n3809 gnd.n3808 585
R1806 gnd.n3807 gnd.n3806 585
R1807 gnd.n3804 gnd.n3803 585
R1808 gnd.n3802 gnd.n3801 585
R1809 gnd.n3800 gnd.n3799 585
R1810 gnd.n3798 gnd.n3797 585
R1811 gnd.n3796 gnd.n3795 585
R1812 gnd.n3794 gnd.n3793 585
R1813 gnd.n3792 gnd.n3791 585
R1814 gnd.n3790 gnd.n3789 585
R1815 gnd.n3788 gnd.n3787 585
R1816 gnd.n3786 gnd.n3785 585
R1817 gnd.n3784 gnd.n3783 585
R1818 gnd.n3782 gnd.n3781 585
R1819 gnd.n3780 gnd.n3779 585
R1820 gnd.n3778 gnd.n3777 585
R1821 gnd.n3776 gnd.n3775 585
R1822 gnd.n3774 gnd.n3773 585
R1823 gnd.n3772 gnd.n3771 585
R1824 gnd.n3770 gnd.n3769 585
R1825 gnd.n3768 gnd.n3739 585
R1826 gnd.n3743 gnd.n3740 585
R1827 gnd.n3764 gnd.n3763 585
R1828 gnd.n4306 gnd.n4305 585
R1829 gnd.n4308 gnd.n1991 585
R1830 gnd.n4310 gnd.n4309 585
R1831 gnd.n4311 gnd.n1984 585
R1832 gnd.n4313 gnd.n4312 585
R1833 gnd.n4315 gnd.n1982 585
R1834 gnd.n4317 gnd.n4316 585
R1835 gnd.n4318 gnd.n1977 585
R1836 gnd.n4320 gnd.n4319 585
R1837 gnd.n4322 gnd.n1975 585
R1838 gnd.n4324 gnd.n4323 585
R1839 gnd.n4325 gnd.n1970 585
R1840 gnd.n4327 gnd.n4326 585
R1841 gnd.n4329 gnd.n1968 585
R1842 gnd.n4331 gnd.n4330 585
R1843 gnd.n4332 gnd.n1963 585
R1844 gnd.n4334 gnd.n4333 585
R1845 gnd.n4336 gnd.n1962 585
R1846 gnd.n4337 gnd.n1905 585
R1847 gnd.n4340 gnd.n4339 585
R1848 gnd.n1906 gnd.n1898 585
R1849 gnd.n1934 gnd.n1899 585
R1850 gnd.n1936 gnd.n1935 585
R1851 gnd.n1938 gnd.n1937 585
R1852 gnd.n1940 gnd.n1939 585
R1853 gnd.n1942 gnd.n1941 585
R1854 gnd.n1944 gnd.n1943 585
R1855 gnd.n1946 gnd.n1945 585
R1856 gnd.n1948 gnd.n1947 585
R1857 gnd.n1950 gnd.n1949 585
R1858 gnd.n1952 gnd.n1951 585
R1859 gnd.n1954 gnd.n1953 585
R1860 gnd.n1956 gnd.n1955 585
R1861 gnd.n1957 gnd.n1916 585
R1862 gnd.n1959 gnd.n1958 585
R1863 gnd.n1917 gnd.n1915 585
R1864 gnd.n1918 gnd.n992 585
R1865 gnd.n1961 gnd.n992 585
R1866 gnd.n4302 gnd.n994 585
R1867 gnd.n5998 gnd.n994 585
R1868 gnd.n4301 gnd.n4300 585
R1869 gnd.n4300 gnd.n4299 585
R1870 gnd.n1995 gnd.n984 585
R1871 gnd.n6004 gnd.n984 585
R1872 gnd.n4060 gnd.n4059 585
R1873 gnd.n4061 gnd.n4060 585
R1874 gnd.n2054 gnd.n973 585
R1875 gnd.n6010 gnd.n973 585
R1876 gnd.n4054 gnd.n4053 585
R1877 gnd.n4053 gnd.n4052 585
R1878 gnd.n4051 gnd.n962 585
R1879 gnd.n6016 gnd.n962 585
R1880 gnd.n4050 gnd.n4049 585
R1881 gnd.n4049 gnd.n4048 585
R1882 gnd.n2056 gnd.n952 585
R1883 gnd.n6022 gnd.n952 585
R1884 gnd.n4043 gnd.n4042 585
R1885 gnd.n4042 gnd.n4041 585
R1886 gnd.n4040 gnd.n941 585
R1887 gnd.n6028 gnd.n941 585
R1888 gnd.n4039 gnd.n2044 585
R1889 gnd.n4078 gnd.n2044 585
R1890 gnd.n2058 gnd.n931 585
R1891 gnd.n6034 gnd.n931 585
R1892 gnd.n4035 gnd.n4034 585
R1893 gnd.n4034 gnd.n4033 585
R1894 gnd.n2060 gnd.n921 585
R1895 gnd.n6040 gnd.n921 585
R1896 gnd.n2097 gnd.n2064 585
R1897 gnd.n4025 gnd.n2064 585
R1898 gnd.n2098 gnd.n910 585
R1899 gnd.n6046 gnd.n910 585
R1900 gnd.n2099 gnd.n2071 585
R1901 gnd.n4012 gnd.n2071 585
R1902 gnd.n2101 gnd.n2100 585
R1903 gnd.n2100 gnd.n2070 585
R1904 gnd.n2102 gnd.n2078 585
R1905 gnd.n4004 gnd.n2078 585
R1906 gnd.n2103 gnd.n2085 585
R1907 gnd.n3998 gnd.n2085 585
R1908 gnd.n3986 gnd.n3985 585
R1909 gnd.n3985 gnd.n3984 585
R1910 gnd.n2104 gnd.n2091 585
R1911 gnd.n3973 gnd.n2104 585
R1912 gnd.n3946 gnd.n2112 585
R1913 gnd.n3976 gnd.n2112 585
R1914 gnd.n3948 gnd.n3947 585
R1915 gnd.n3949 gnd.n3948 585
R1916 gnd.n2117 gnd.n895 585
R1917 gnd.n6054 gnd.n895 585
R1918 gnd.n3941 gnd.n3940 585
R1919 gnd.n3940 gnd.n3939 585
R1920 gnd.n2119 gnd.n884 585
R1921 gnd.n6060 gnd.n884 585
R1922 gnd.n3891 gnd.n2123 585
R1923 gnd.n3929 gnd.n2123 585
R1924 gnd.n3892 gnd.n874 585
R1925 gnd.n6066 gnd.n874 585
R1926 gnd.n3894 gnd.n3893 585
R1927 gnd.n3895 gnd.n3894 585
R1928 gnd.n2134 gnd.n863 585
R1929 gnd.n6072 gnd.n863 585
R1930 gnd.n3885 gnd.n2129 585
R1931 gnd.n3901 gnd.n2129 585
R1932 gnd.n3884 gnd.n853 585
R1933 gnd.n6078 gnd.n853 585
R1934 gnd.n3883 gnd.n3882 585
R1935 gnd.n3882 gnd.n3881 585
R1936 gnd.n2136 gnd.n841 585
R1937 gnd.n6084 gnd.n841 585
R1938 gnd.n3752 gnd.n3751 585
R1939 gnd.n3751 gnd.n830 585
R1940 gnd.n3753 gnd.n828 585
R1941 gnd.n6090 gnd.n828 585
R1942 gnd.n3755 gnd.n3754 585
R1943 gnd.n3754 gnd.n827 585
R1944 gnd.n3756 gnd.n2144 585
R1945 gnd.n3868 gnd.n2144 585
R1946 gnd.n3746 gnd.n3745 585
R1947 gnd.n3745 gnd.n2143 585
R1948 gnd.n3760 gnd.n2152 585
R1949 gnd.n3859 gnd.n2152 585
R1950 gnd.n3762 gnd.n3761 585
R1951 gnd.n3762 gnd.n2151 585
R1952 gnd.n7149 gnd.n7148 585
R1953 gnd.n7150 gnd.n7149 585
R1954 gnd.n87 gnd.n85 585
R1955 gnd.n85 gnd.n81 585
R1956 gnd.n7069 gnd.n7068 585
R1957 gnd.n7070 gnd.n7069 585
R1958 gnd.n164 gnd.n163 585
R1959 gnd.n163 gnd.n161 585
R1960 gnd.n7064 gnd.n7063 585
R1961 gnd.n7063 gnd.n7062 585
R1962 gnd.n167 gnd.n166 585
R1963 gnd.n180 gnd.n167 585
R1964 gnd.n6979 gnd.n6978 585
R1965 gnd.n6980 gnd.n6979 585
R1966 gnd.n182 gnd.n181 585
R1967 gnd.n261 gnd.n181 585
R1968 gnd.n6974 gnd.n6973 585
R1969 gnd.n6973 gnd.n6972 585
R1970 gnd.n185 gnd.n184 585
R1971 gnd.n266 gnd.n185 585
R1972 gnd.n6963 gnd.n6962 585
R1973 gnd.n6964 gnd.n6963 585
R1974 gnd.n198 gnd.n197 585
R1975 gnd.n6907 gnd.n197 585
R1976 gnd.n6958 gnd.n6957 585
R1977 gnd.n6957 gnd.n6956 585
R1978 gnd.n201 gnd.n200 585
R1979 gnd.n6912 gnd.n201 585
R1980 gnd.n6947 gnd.n6946 585
R1981 gnd.n6948 gnd.n6947 585
R1982 gnd.n213 gnd.n212 585
R1983 gnd.n6916 gnd.n212 585
R1984 gnd.n6942 gnd.n6941 585
R1985 gnd.n6941 gnd.n6940 585
R1986 gnd.n222 gnd.n221 585
R1987 gnd.n6921 gnd.n222 585
R1988 gnd.n6931 gnd.n6930 585
R1989 gnd.n6932 gnd.n6931 585
R1990 gnd.n6929 gnd.n6928 585
R1991 gnd.n6928 gnd.n6927 585
R1992 gnd.n5776 gnd.n234 585
R1993 gnd.n5810 gnd.n234 585
R1994 gnd.n5778 gnd.n5777 585
R1995 gnd.n5778 gnd.n1170 585
R1996 gnd.n5781 gnd.n5780 585
R1997 gnd.n5782 gnd.n5781 585
R1998 gnd.n5779 gnd.n5775 585
R1999 gnd.n5775 gnd.n1176 585
R2000 gnd.n5774 gnd.n1183 585
R2001 gnd.n5774 gnd.n5773 585
R2002 gnd.n1182 gnd.n1181 585
R2003 gnd.n5650 gnd.n1181 585
R2004 gnd.n5762 gnd.n5761 585
R2005 gnd.n5763 gnd.n5762 585
R2006 gnd.n5760 gnd.n1197 585
R2007 gnd.n1205 gnd.n1197 585
R2008 gnd.n5759 gnd.n5758 585
R2009 gnd.n5758 gnd.n5757 585
R2010 gnd.n1200 gnd.n1198 585
R2011 gnd.n5739 gnd.n1200 585
R2012 gnd.n5727 gnd.n1225 585
R2013 gnd.n1225 gnd.n1212 585
R2014 gnd.n5729 gnd.n5728 585
R2015 gnd.n5730 gnd.n5729 585
R2016 gnd.n1226 gnd.n1224 585
R2017 gnd.n1233 gnd.n1224 585
R2018 gnd.n5721 gnd.n5720 585
R2019 gnd.n5720 gnd.n5719 585
R2020 gnd.n1229 gnd.n1228 585
R2021 gnd.n5707 gnd.n1229 585
R2022 gnd.n5695 gnd.n1253 585
R2023 gnd.n1253 gnd.n1241 585
R2024 gnd.n5697 gnd.n5696 585
R2025 gnd.n5698 gnd.n5697 585
R2026 gnd.n1254 gnd.n1252 585
R2027 gnd.n5670 gnd.n1252 585
R2028 gnd.n5690 gnd.n5689 585
R2029 gnd.n5689 gnd.n5688 585
R2030 gnd.n1137 gnd.n1136 585
R2031 gnd.n5621 gnd.n1137 585
R2032 gnd.n5847 gnd.n5846 585
R2033 gnd.n5846 gnd.n5845 585
R2034 gnd.n5848 gnd.n1132 585
R2035 gnd.n5612 gnd.n1132 585
R2036 gnd.n5850 gnd.n5849 585
R2037 gnd.n5851 gnd.n5850 585
R2038 gnd.n5511 gnd.n1131 585
R2039 gnd.n5516 gnd.n5514 585
R2040 gnd.n5517 gnd.n5510 585
R2041 gnd.n5517 gnd.n1118 585
R2042 gnd.n5520 gnd.n5519 585
R2043 gnd.n5508 gnd.n5507 585
R2044 gnd.n5525 gnd.n5524 585
R2045 gnd.n5527 gnd.n5506 585
R2046 gnd.n5530 gnd.n5529 585
R2047 gnd.n5504 gnd.n5503 585
R2048 gnd.n5535 gnd.n5534 585
R2049 gnd.n5537 gnd.n5502 585
R2050 gnd.n5540 gnd.n5539 585
R2051 gnd.n5500 gnd.n5499 585
R2052 gnd.n5546 gnd.n5545 585
R2053 gnd.n5548 gnd.n5498 585
R2054 gnd.n5549 gnd.n1291 585
R2055 gnd.n1289 gnd.n1288 585
R2056 gnd.n5559 gnd.n5558 585
R2057 gnd.n5561 gnd.n1287 585
R2058 gnd.n5564 gnd.n5563 585
R2059 gnd.n1285 gnd.n1284 585
R2060 gnd.n5569 gnd.n5568 585
R2061 gnd.n5571 gnd.n1283 585
R2062 gnd.n5574 gnd.n5573 585
R2063 gnd.n1281 gnd.n1280 585
R2064 gnd.n5579 gnd.n5578 585
R2065 gnd.n5581 gnd.n1279 585
R2066 gnd.n5584 gnd.n5583 585
R2067 gnd.n1277 gnd.n1276 585
R2068 gnd.n5589 gnd.n5588 585
R2069 gnd.n5591 gnd.n1275 585
R2070 gnd.n5594 gnd.n5593 585
R2071 gnd.n1273 gnd.n1272 585
R2072 gnd.n5600 gnd.n5599 585
R2073 gnd.n5602 gnd.n1271 585
R2074 gnd.n5603 gnd.n1270 585
R2075 gnd.n5606 gnd.n5605 585
R2076 gnd.n155 gnd.n154 585
R2077 gnd.n7078 gnd.n150 585
R2078 gnd.n7080 gnd.n7079 585
R2079 gnd.n7082 gnd.n148 585
R2080 gnd.n7084 gnd.n7083 585
R2081 gnd.n7085 gnd.n143 585
R2082 gnd.n7087 gnd.n7086 585
R2083 gnd.n7089 gnd.n141 585
R2084 gnd.n7091 gnd.n7090 585
R2085 gnd.n7092 gnd.n136 585
R2086 gnd.n7094 gnd.n7093 585
R2087 gnd.n7096 gnd.n134 585
R2088 gnd.n7098 gnd.n7097 585
R2089 gnd.n7099 gnd.n129 585
R2090 gnd.n7101 gnd.n7100 585
R2091 gnd.n7103 gnd.n127 585
R2092 gnd.n7105 gnd.n7104 585
R2093 gnd.n7106 gnd.n122 585
R2094 gnd.n7108 gnd.n7107 585
R2095 gnd.n7110 gnd.n120 585
R2096 gnd.n7112 gnd.n7111 585
R2097 gnd.n7116 gnd.n115 585
R2098 gnd.n7118 gnd.n7117 585
R2099 gnd.n7120 gnd.n113 585
R2100 gnd.n7122 gnd.n7121 585
R2101 gnd.n7123 gnd.n108 585
R2102 gnd.n7125 gnd.n7124 585
R2103 gnd.n7127 gnd.n106 585
R2104 gnd.n7129 gnd.n7128 585
R2105 gnd.n7130 gnd.n101 585
R2106 gnd.n7132 gnd.n7131 585
R2107 gnd.n7134 gnd.n99 585
R2108 gnd.n7136 gnd.n7135 585
R2109 gnd.n7137 gnd.n94 585
R2110 gnd.n7139 gnd.n7138 585
R2111 gnd.n7141 gnd.n92 585
R2112 gnd.n7143 gnd.n7142 585
R2113 gnd.n7144 gnd.n90 585
R2114 gnd.n7145 gnd.n86 585
R2115 gnd.n86 gnd.n83 585
R2116 gnd.n7074 gnd.n82 585
R2117 gnd.n7150 gnd.n82 585
R2118 gnd.n7073 gnd.n7072 585
R2119 gnd.n7072 gnd.n81 585
R2120 gnd.n7071 gnd.n159 585
R2121 gnd.n7071 gnd.n7070 585
R2122 gnd.n256 gnd.n160 585
R2123 gnd.n161 gnd.n160 585
R2124 gnd.n257 gnd.n169 585
R2125 gnd.n7062 gnd.n169 585
R2126 gnd.n259 gnd.n258 585
R2127 gnd.n258 gnd.n180 585
R2128 gnd.n260 gnd.n178 585
R2129 gnd.n6980 gnd.n178 585
R2130 gnd.n263 gnd.n262 585
R2131 gnd.n262 gnd.n261 585
R2132 gnd.n264 gnd.n187 585
R2133 gnd.n6972 gnd.n187 585
R2134 gnd.n268 gnd.n267 585
R2135 gnd.n267 gnd.n266 585
R2136 gnd.n269 gnd.n195 585
R2137 gnd.n6964 gnd.n195 585
R2138 gnd.n6909 gnd.n6908 585
R2139 gnd.n6908 gnd.n6907 585
R2140 gnd.n6910 gnd.n203 585
R2141 gnd.n6956 gnd.n203 585
R2142 gnd.n6914 gnd.n6913 585
R2143 gnd.n6913 gnd.n6912 585
R2144 gnd.n6915 gnd.n210 585
R2145 gnd.n6948 gnd.n210 585
R2146 gnd.n6918 gnd.n6917 585
R2147 gnd.n6917 gnd.n6916 585
R2148 gnd.n6919 gnd.n224 585
R2149 gnd.n6940 gnd.n224 585
R2150 gnd.n6923 gnd.n6922 585
R2151 gnd.n6922 gnd.n6921 585
R2152 gnd.n6924 gnd.n232 585
R2153 gnd.n6932 gnd.n232 585
R2154 gnd.n6926 gnd.n6925 585
R2155 gnd.n6927 gnd.n6926 585
R2156 gnd.n237 gnd.n236 585
R2157 gnd.n5810 gnd.n236 585
R2158 gnd.n5645 gnd.n5644 585
R2159 gnd.n5644 gnd.n1170 585
R2160 gnd.n5646 gnd.n1177 585
R2161 gnd.n5782 gnd.n1177 585
R2162 gnd.n5648 gnd.n5647 585
R2163 gnd.n5647 gnd.n1176 585
R2164 gnd.n5649 gnd.n1185 585
R2165 gnd.n5773 gnd.n1185 585
R2166 gnd.n5652 gnd.n5651 585
R2167 gnd.n5651 gnd.n5650 585
R2168 gnd.n5653 gnd.n1195 585
R2169 gnd.n5763 gnd.n1195 585
R2170 gnd.n5655 gnd.n5654 585
R2171 gnd.n5654 gnd.n1205 585
R2172 gnd.n5656 gnd.n1202 585
R2173 gnd.n5757 gnd.n1202 585
R2174 gnd.n5657 gnd.n1213 585
R2175 gnd.n5739 gnd.n1213 585
R2176 gnd.n5659 gnd.n5658 585
R2177 gnd.n5658 gnd.n1212 585
R2178 gnd.n5660 gnd.n1221 585
R2179 gnd.n5730 gnd.n1221 585
R2180 gnd.n5662 gnd.n5661 585
R2181 gnd.n5661 gnd.n1233 585
R2182 gnd.n5663 gnd.n1231 585
R2183 gnd.n5719 gnd.n1231 585
R2184 gnd.n5664 gnd.n1242 585
R2185 gnd.n5707 gnd.n1242 585
R2186 gnd.n5666 gnd.n5665 585
R2187 gnd.n5665 gnd.n1241 585
R2188 gnd.n5667 gnd.n1250 585
R2189 gnd.n5698 gnd.n1250 585
R2190 gnd.n5669 gnd.n5668 585
R2191 gnd.n5670 gnd.n5669 585
R2192 gnd.n1259 gnd.n1257 585
R2193 gnd.n5688 gnd.n1257 585
R2194 gnd.n5623 gnd.n5622 585
R2195 gnd.n5622 gnd.n5621 585
R2196 gnd.n1261 gnd.n1139 585
R2197 gnd.n5845 gnd.n1139 585
R2198 gnd.n5611 gnd.n5610 585
R2199 gnd.n5612 gnd.n5611 585
R2200 gnd.n1266 gnd.n1127 585
R2201 gnd.n5851 gnd.n1127 585
R2202 gnd.n5425 gnd.n5424 585
R2203 gnd.n5426 gnd.n5425 585
R2204 gnd.n5339 gnd.n1334 585
R2205 gnd.n1340 gnd.n1334 585
R2206 gnd.n5338 gnd.n5337 585
R2207 gnd.n5337 gnd.n5336 585
R2208 gnd.n1337 gnd.n1336 585
R2209 gnd.n1426 gnd.n1337 585
R2210 gnd.n5129 gnd.n1364 585
R2211 gnd.n1428 gnd.n1364 585
R2212 gnd.n5131 gnd.n5130 585
R2213 gnd.n5132 gnd.n5131 585
R2214 gnd.n5128 gnd.n1363 585
R2215 gnd.n5123 gnd.n1363 585
R2216 gnd.n5127 gnd.n5126 585
R2217 gnd.n5126 gnd.n5125 585
R2218 gnd.n1366 gnd.n1365 585
R2219 gnd.n5110 gnd.n1366 585
R2220 gnd.n5095 gnd.n1387 585
R2221 gnd.n1387 gnd.n1376 585
R2222 gnd.n5097 gnd.n5096 585
R2223 gnd.n5098 gnd.n5097 585
R2224 gnd.n5094 gnd.n1386 585
R2225 gnd.n1386 gnd.n1383 585
R2226 gnd.n5093 gnd.n5092 585
R2227 gnd.n5092 gnd.n5091 585
R2228 gnd.n1389 gnd.n1388 585
R2229 gnd.n1442 gnd.n1389 585
R2230 gnd.n5080 gnd.n5079 585
R2231 gnd.n5081 gnd.n5080 585
R2232 gnd.n5078 gnd.n1400 585
R2233 gnd.n1400 gnd.n1397 585
R2234 gnd.n5077 gnd.n5076 585
R2235 gnd.n5076 gnd.n5075 585
R2236 gnd.n1402 gnd.n1401 585
R2237 gnd.n5050 gnd.n1402 585
R2238 gnd.n5063 gnd.n5062 585
R2239 gnd.n5064 gnd.n5063 585
R2240 gnd.n5061 gnd.n1414 585
R2241 gnd.n5056 gnd.n1414 585
R2242 gnd.n5060 gnd.n5059 585
R2243 gnd.n5059 gnd.n5058 585
R2244 gnd.n1416 gnd.n1415 585
R2245 gnd.n5036 gnd.n1416 585
R2246 gnd.n5027 gnd.n1462 585
R2247 gnd.n1462 gnd.n1454 585
R2248 gnd.n5029 gnd.n5028 585
R2249 gnd.n5030 gnd.n5029 585
R2250 gnd.n5026 gnd.n1461 585
R2251 gnd.n4987 gnd.n1461 585
R2252 gnd.n5025 gnd.n5024 585
R2253 gnd.n5024 gnd.n5023 585
R2254 gnd.n1464 gnd.n1463 585
R2255 gnd.n4931 gnd.n1464 585
R2256 gnd.n5009 gnd.n5008 585
R2257 gnd.n5010 gnd.n5009 585
R2258 gnd.n5007 gnd.n1476 585
R2259 gnd.n1476 gnd.n1472 585
R2260 gnd.n5006 gnd.n5005 585
R2261 gnd.n5005 gnd.n5004 585
R2262 gnd.n1478 gnd.n1477 585
R2263 gnd.n4938 gnd.n1478 585
R2264 gnd.n4978 gnd.n4977 585
R2265 gnd.n4979 gnd.n4978 585
R2266 gnd.n4976 gnd.n1490 585
R2267 gnd.n1490 gnd.n1487 585
R2268 gnd.n4975 gnd.n4974 585
R2269 gnd.n4974 gnd.n4973 585
R2270 gnd.n1492 gnd.n1491 585
R2271 gnd.n4946 gnd.n1492 585
R2272 gnd.n4959 gnd.n4958 585
R2273 gnd.n4960 gnd.n4959 585
R2274 gnd.n4957 gnd.n1504 585
R2275 gnd.n4952 gnd.n1504 585
R2276 gnd.n4956 gnd.n4955 585
R2277 gnd.n4955 gnd.n4954 585
R2278 gnd.n1506 gnd.n1505 585
R2279 gnd.n4926 gnd.n1506 585
R2280 gnd.n4908 gnd.n1520 585
R2281 gnd.n4894 gnd.n1520 585
R2282 gnd.n4910 gnd.n4909 585
R2283 gnd.n4911 gnd.n4910 585
R2284 gnd.n4907 gnd.n1519 585
R2285 gnd.n1525 gnd.n1519 585
R2286 gnd.n4906 gnd.n4905 585
R2287 gnd.n4905 gnd.n4904 585
R2288 gnd.n1522 gnd.n1521 585
R2289 gnd.n4884 gnd.n1522 585
R2290 gnd.n4871 gnd.n1539 585
R2291 gnd.n1539 gnd.n1532 585
R2292 gnd.n4873 gnd.n4872 585
R2293 gnd.n4874 gnd.n4873 585
R2294 gnd.n4870 gnd.n1538 585
R2295 gnd.n1544 gnd.n1538 585
R2296 gnd.n4869 gnd.n4868 585
R2297 gnd.n4868 gnd.n4867 585
R2298 gnd.n1541 gnd.n1540 585
R2299 gnd.n4779 gnd.n1541 585
R2300 gnd.n4855 gnd.n4854 585
R2301 gnd.n4856 gnd.n4855 585
R2302 gnd.n4853 gnd.n1556 585
R2303 gnd.n1556 gnd.n1552 585
R2304 gnd.n4852 gnd.n4851 585
R2305 gnd.n4851 gnd.n4850 585
R2306 gnd.n1558 gnd.n1557 585
R2307 gnd.n4788 gnd.n1558 585
R2308 gnd.n4826 gnd.n4825 585
R2309 gnd.n4827 gnd.n4826 585
R2310 gnd.n4824 gnd.n1570 585
R2311 gnd.n1570 gnd.n1567 585
R2312 gnd.n4823 gnd.n4822 585
R2313 gnd.n4822 gnd.n4821 585
R2314 gnd.n1572 gnd.n1571 585
R2315 gnd.n4795 gnd.n1572 585
R2316 gnd.n4808 gnd.n4807 585
R2317 gnd.n4809 gnd.n4808 585
R2318 gnd.n4806 gnd.n1585 585
R2319 gnd.n4801 gnd.n1585 585
R2320 gnd.n4805 gnd.n4804 585
R2321 gnd.n4804 gnd.n4803 585
R2322 gnd.n1587 gnd.n1586 585
R2323 gnd.n4774 gnd.n1587 585
R2324 gnd.n4760 gnd.n4759 585
R2325 gnd.n4759 gnd.n4758 585
R2326 gnd.n4761 gnd.n1603 585
R2327 gnd.n4756 gnd.n1603 585
R2328 gnd.n4763 gnd.n4762 585
R2329 gnd.n4764 gnd.n4763 585
R2330 gnd.n1604 gnd.n1602 585
R2331 gnd.n4750 gnd.n1602 585
R2332 gnd.n4747 gnd.n4746 585
R2333 gnd.n4748 gnd.n4747 585
R2334 gnd.n4745 gnd.n1607 585
R2335 gnd.n1613 gnd.n1607 585
R2336 gnd.n4744 gnd.n4743 585
R2337 gnd.n4743 gnd.n4742 585
R2338 gnd.n1609 gnd.n1608 585
R2339 gnd.n4730 gnd.n1609 585
R2340 gnd.n4718 gnd.n1628 585
R2341 gnd.n1628 gnd.n1619 585
R2342 gnd.n4720 gnd.n4719 585
R2343 gnd.n4721 gnd.n4720 585
R2344 gnd.n4717 gnd.n1627 585
R2345 gnd.n1633 gnd.n1627 585
R2346 gnd.n4716 gnd.n4715 585
R2347 gnd.n4715 gnd.n4714 585
R2348 gnd.n1630 gnd.n1629 585
R2349 gnd.n4602 gnd.n1630 585
R2350 gnd.n4702 gnd.n4701 585
R2351 gnd.n4703 gnd.n4702 585
R2352 gnd.n4700 gnd.n1644 585
R2353 gnd.n1644 gnd.n1640 585
R2354 gnd.n4699 gnd.n4698 585
R2355 gnd.n4698 gnd.n4697 585
R2356 gnd.n1646 gnd.n1645 585
R2357 gnd.n4610 gnd.n1646 585
R2358 gnd.n4649 gnd.n4648 585
R2359 gnd.n4650 gnd.n4649 585
R2360 gnd.n4647 gnd.n1657 585
R2361 gnd.n1661 gnd.n1657 585
R2362 gnd.n4646 gnd.n4645 585
R2363 gnd.n4645 gnd.n4644 585
R2364 gnd.n1659 gnd.n1658 585
R2365 gnd.n4618 gnd.n1659 585
R2366 gnd.n4631 gnd.n4630 585
R2367 gnd.n4632 gnd.n4631 585
R2368 gnd.n4629 gnd.n1672 585
R2369 gnd.n4624 gnd.n1672 585
R2370 gnd.n4628 gnd.n4627 585
R2371 gnd.n4627 gnd.n4626 585
R2372 gnd.n1674 gnd.n1673 585
R2373 gnd.n4597 gnd.n1674 585
R2374 gnd.n4583 gnd.n4582 585
R2375 gnd.n4582 gnd.n4581 585
R2376 gnd.n4584 gnd.n1688 585
R2377 gnd.n4530 gnd.n1688 585
R2378 gnd.n4586 gnd.n4585 585
R2379 gnd.n4587 gnd.n4586 585
R2380 gnd.n1689 gnd.n1687 585
R2381 gnd.n4534 gnd.n1687 585
R2382 gnd.n4562 gnd.n4561 585
R2383 gnd.n4563 gnd.n4562 585
R2384 gnd.n4560 gnd.n1700 585
R2385 gnd.n1704 gnd.n1700 585
R2386 gnd.n4559 gnd.n4558 585
R2387 gnd.n4558 gnd.n4557 585
R2388 gnd.n1702 gnd.n1701 585
R2389 gnd.n4544 gnd.n1702 585
R2390 gnd.n4523 gnd.n1718 585
R2391 gnd.n1718 gnd.n1710 585
R2392 gnd.n4525 gnd.n4524 585
R2393 gnd.n4526 gnd.n4525 585
R2394 gnd.n4522 gnd.n1717 585
R2395 gnd.n1723 gnd.n1717 585
R2396 gnd.n4521 gnd.n4520 585
R2397 gnd.n4520 gnd.n4519 585
R2398 gnd.n1720 gnd.n1719 585
R2399 gnd.n4428 gnd.n1720 585
R2400 gnd.n4506 gnd.n4505 585
R2401 gnd.n4507 gnd.n4506 585
R2402 gnd.n4504 gnd.n1734 585
R2403 gnd.n1734 gnd.n1730 585
R2404 gnd.n4503 gnd.n4502 585
R2405 gnd.n4502 gnd.n4501 585
R2406 gnd.n1736 gnd.n1735 585
R2407 gnd.n4436 gnd.n1736 585
R2408 gnd.n4476 gnd.n4475 585
R2409 gnd.n4477 gnd.n4476 585
R2410 gnd.n4474 gnd.n1748 585
R2411 gnd.n1748 gnd.n1745 585
R2412 gnd.n4473 gnd.n4472 585
R2413 gnd.n4472 gnd.n4471 585
R2414 gnd.n1750 gnd.n1749 585
R2415 gnd.n4444 gnd.n1750 585
R2416 gnd.n4457 gnd.n4456 585
R2417 gnd.n4458 gnd.n4457 585
R2418 gnd.n4455 gnd.n1761 585
R2419 gnd.n4450 gnd.n1761 585
R2420 gnd.n4454 gnd.n4453 585
R2421 gnd.n4453 gnd.n4452 585
R2422 gnd.n1763 gnd.n1762 585
R2423 gnd.n4423 gnd.n1763 585
R2424 gnd.n4410 gnd.n4409 585
R2425 gnd.n4408 gnd.n1809 585
R2426 gnd.n4407 gnd.n1808 585
R2427 gnd.n4412 gnd.n1808 585
R2428 gnd.n4406 gnd.n4405 585
R2429 gnd.n4404 gnd.n4403 585
R2430 gnd.n4402 gnd.n4401 585
R2431 gnd.n4400 gnd.n4399 585
R2432 gnd.n4398 gnd.n4397 585
R2433 gnd.n4396 gnd.n4395 585
R2434 gnd.n4394 gnd.n4393 585
R2435 gnd.n4392 gnd.n4391 585
R2436 gnd.n4390 gnd.n4389 585
R2437 gnd.n4388 gnd.n4387 585
R2438 gnd.n4386 gnd.n4385 585
R2439 gnd.n4384 gnd.n4383 585
R2440 gnd.n4382 gnd.n4381 585
R2441 gnd.n4380 gnd.n4379 585
R2442 gnd.n4378 gnd.n4377 585
R2443 gnd.n4376 gnd.n4375 585
R2444 gnd.n4374 gnd.n4373 585
R2445 gnd.n4372 gnd.n4371 585
R2446 gnd.n4370 gnd.n4369 585
R2447 gnd.n4368 gnd.n4367 585
R2448 gnd.n4366 gnd.n4365 585
R2449 gnd.n4364 gnd.n4363 585
R2450 gnd.n4362 gnd.n4361 585
R2451 gnd.n4360 gnd.n4359 585
R2452 gnd.n4358 gnd.n4357 585
R2453 gnd.n4356 gnd.n4355 585
R2454 gnd.n4354 gnd.n4353 585
R2455 gnd.n4352 gnd.n4351 585
R2456 gnd.n4350 gnd.n4349 585
R2457 gnd.n4348 gnd.n4347 585
R2458 gnd.n4346 gnd.n1897 585
R2459 gnd.n1896 gnd.n1895 585
R2460 gnd.n1894 gnd.n1893 585
R2461 gnd.n1891 gnd.n1890 585
R2462 gnd.n1889 gnd.n1888 585
R2463 gnd.n1887 gnd.n1886 585
R2464 gnd.n1885 gnd.n1884 585
R2465 gnd.n1883 gnd.n1882 585
R2466 gnd.n1881 gnd.n1880 585
R2467 gnd.n1879 gnd.n1878 585
R2468 gnd.n1877 gnd.n1876 585
R2469 gnd.n1875 gnd.n1874 585
R2470 gnd.n1873 gnd.n1872 585
R2471 gnd.n1871 gnd.n1870 585
R2472 gnd.n1869 gnd.n1868 585
R2473 gnd.n1867 gnd.n1866 585
R2474 gnd.n1865 gnd.n1864 585
R2475 gnd.n1863 gnd.n1862 585
R2476 gnd.n1861 gnd.n1860 585
R2477 gnd.n1859 gnd.n1858 585
R2478 gnd.n1857 gnd.n1856 585
R2479 gnd.n1855 gnd.n1854 585
R2480 gnd.n1853 gnd.n1852 585
R2481 gnd.n1851 gnd.n1850 585
R2482 gnd.n1849 gnd.n1848 585
R2483 gnd.n1847 gnd.n1846 585
R2484 gnd.n1845 gnd.n1844 585
R2485 gnd.n1843 gnd.n1842 585
R2486 gnd.n1841 gnd.n1840 585
R2487 gnd.n1839 gnd.n1838 585
R2488 gnd.n1837 gnd.n1836 585
R2489 gnd.n1767 gnd.n1766 585
R2490 gnd.n5429 gnd.n5428 585
R2491 gnd.n5431 gnd.n5430 585
R2492 gnd.n5433 gnd.n5432 585
R2493 gnd.n5435 gnd.n5434 585
R2494 gnd.n5437 gnd.n5436 585
R2495 gnd.n5439 gnd.n5438 585
R2496 gnd.n5441 gnd.n5440 585
R2497 gnd.n5443 gnd.n5442 585
R2498 gnd.n5445 gnd.n5444 585
R2499 gnd.n5447 gnd.n5446 585
R2500 gnd.n5449 gnd.n5448 585
R2501 gnd.n5451 gnd.n5450 585
R2502 gnd.n5453 gnd.n5452 585
R2503 gnd.n5455 gnd.n5454 585
R2504 gnd.n5457 gnd.n5456 585
R2505 gnd.n5459 gnd.n5458 585
R2506 gnd.n5461 gnd.n5460 585
R2507 gnd.n5463 gnd.n5462 585
R2508 gnd.n5465 gnd.n5464 585
R2509 gnd.n5467 gnd.n5466 585
R2510 gnd.n5469 gnd.n5468 585
R2511 gnd.n5471 gnd.n5470 585
R2512 gnd.n5473 gnd.n5472 585
R2513 gnd.n5475 gnd.n5474 585
R2514 gnd.n5477 gnd.n5476 585
R2515 gnd.n5479 gnd.n5478 585
R2516 gnd.n5481 gnd.n5480 585
R2517 gnd.n5483 gnd.n5482 585
R2518 gnd.n5485 gnd.n5484 585
R2519 gnd.n5487 gnd.n1328 585
R2520 gnd.n5489 gnd.n5488 585
R2521 gnd.n5491 gnd.n1292 585
R2522 gnd.n5493 gnd.n5492 585
R2523 gnd.n5496 gnd.n5495 585
R2524 gnd.n1295 gnd.n1293 585
R2525 gnd.n5362 gnd.n5361 585
R2526 gnd.n5364 gnd.n5363 585
R2527 gnd.n5367 gnd.n5366 585
R2528 gnd.n5369 gnd.n5368 585
R2529 gnd.n5371 gnd.n5370 585
R2530 gnd.n5373 gnd.n5372 585
R2531 gnd.n5375 gnd.n5374 585
R2532 gnd.n5377 gnd.n5376 585
R2533 gnd.n5379 gnd.n5378 585
R2534 gnd.n5381 gnd.n5380 585
R2535 gnd.n5383 gnd.n5382 585
R2536 gnd.n5385 gnd.n5384 585
R2537 gnd.n5387 gnd.n5386 585
R2538 gnd.n5389 gnd.n5388 585
R2539 gnd.n5391 gnd.n5390 585
R2540 gnd.n5393 gnd.n5392 585
R2541 gnd.n5395 gnd.n5394 585
R2542 gnd.n5397 gnd.n5396 585
R2543 gnd.n5399 gnd.n5398 585
R2544 gnd.n5401 gnd.n5400 585
R2545 gnd.n5403 gnd.n5402 585
R2546 gnd.n5405 gnd.n5404 585
R2547 gnd.n5407 gnd.n5406 585
R2548 gnd.n5409 gnd.n5408 585
R2549 gnd.n5411 gnd.n5410 585
R2550 gnd.n5413 gnd.n5412 585
R2551 gnd.n5415 gnd.n5414 585
R2552 gnd.n5417 gnd.n5416 585
R2553 gnd.n5419 gnd.n5418 585
R2554 gnd.n5421 gnd.n5420 585
R2555 gnd.n5422 gnd.n1335 585
R2556 gnd.n5427 gnd.n1331 585
R2557 gnd.n5427 gnd.n5426 585
R2558 gnd.n1420 gnd.n1332 585
R2559 gnd.n1340 gnd.n1332 585
R2560 gnd.n1421 gnd.n1339 585
R2561 gnd.n5336 gnd.n1339 585
R2562 gnd.n1423 gnd.n1422 585
R2563 gnd.n1426 gnd.n1423 585
R2564 gnd.n1430 gnd.n1429 585
R2565 gnd.n1429 gnd.n1428 585
R2566 gnd.n1431 gnd.n1361 585
R2567 gnd.n5132 gnd.n1361 585
R2568 gnd.n1432 gnd.n1369 585
R2569 gnd.n5123 gnd.n1369 585
R2570 gnd.n1433 gnd.n1368 585
R2571 gnd.n5125 gnd.n1368 585
R2572 gnd.n1434 gnd.n1377 585
R2573 gnd.n5110 gnd.n1377 585
R2574 gnd.n1436 gnd.n1435 585
R2575 gnd.n1435 gnd.n1376 585
R2576 gnd.n1437 gnd.n1384 585
R2577 gnd.n5098 gnd.n1384 585
R2578 gnd.n1439 gnd.n1438 585
R2579 gnd.n1438 gnd.n1383 585
R2580 gnd.n1440 gnd.n1391 585
R2581 gnd.n5091 gnd.n1391 585
R2582 gnd.n1444 gnd.n1443 585
R2583 gnd.n1443 gnd.n1442 585
R2584 gnd.n1445 gnd.n1398 585
R2585 gnd.n5081 gnd.n1398 585
R2586 gnd.n1447 gnd.n1446 585
R2587 gnd.n1446 gnd.n1397 585
R2588 gnd.n1448 gnd.n1404 585
R2589 gnd.n5075 gnd.n1404 585
R2590 gnd.n5052 gnd.n5051 585
R2591 gnd.n5051 gnd.n5050 585
R2592 gnd.n5053 gnd.n1413 585
R2593 gnd.n5064 gnd.n1413 585
R2594 gnd.n5055 gnd.n5054 585
R2595 gnd.n5056 gnd.n5055 585
R2596 gnd.n1419 gnd.n1418 585
R2597 gnd.n5058 gnd.n1418 585
R2598 gnd.n5035 gnd.n5034 585
R2599 gnd.n5036 gnd.n5035 585
R2600 gnd.n5033 gnd.n1456 585
R2601 gnd.n1456 gnd.n1454 585
R2602 gnd.n5032 gnd.n5031 585
R2603 gnd.n5031 gnd.n5030 585
R2604 gnd.n1458 gnd.n1457 585
R2605 gnd.n4987 gnd.n1458 585
R2606 gnd.n4930 gnd.n1466 585
R2607 gnd.n5023 gnd.n1466 585
R2608 gnd.n4933 gnd.n4932 585
R2609 gnd.n4932 gnd.n4931 585
R2610 gnd.n4934 gnd.n1474 585
R2611 gnd.n5010 gnd.n1474 585
R2612 gnd.n4936 gnd.n4935 585
R2613 gnd.n4935 gnd.n1472 585
R2614 gnd.n4937 gnd.n1480 585
R2615 gnd.n5004 gnd.n1480 585
R2616 gnd.n4940 gnd.n4939 585
R2617 gnd.n4939 gnd.n4938 585
R2618 gnd.n4941 gnd.n1488 585
R2619 gnd.n4979 gnd.n1488 585
R2620 gnd.n4943 gnd.n4942 585
R2621 gnd.n4942 gnd.n1487 585
R2622 gnd.n4944 gnd.n1493 585
R2623 gnd.n4973 gnd.n1493 585
R2624 gnd.n4948 gnd.n4947 585
R2625 gnd.n4947 gnd.n4946 585
R2626 gnd.n4949 gnd.n1501 585
R2627 gnd.n4960 gnd.n1501 585
R2628 gnd.n4951 gnd.n4950 585
R2629 gnd.n4952 gnd.n4951 585
R2630 gnd.n4929 gnd.n1507 585
R2631 gnd.n4954 gnd.n1507 585
R2632 gnd.n4928 gnd.n4927 585
R2633 gnd.n4927 gnd.n4926 585
R2634 gnd.n1509 gnd.n1508 585
R2635 gnd.n4894 gnd.n1509 585
R2636 gnd.n4878 gnd.n1517 585
R2637 gnd.n4911 gnd.n1517 585
R2638 gnd.n4880 gnd.n4879 585
R2639 gnd.n4879 gnd.n1525 585
R2640 gnd.n4881 gnd.n1524 585
R2641 gnd.n4904 gnd.n1524 585
R2642 gnd.n4883 gnd.n4882 585
R2643 gnd.n4884 gnd.n4883 585
R2644 gnd.n4877 gnd.n1534 585
R2645 gnd.n1534 gnd.n1532 585
R2646 gnd.n4876 gnd.n4875 585
R2647 gnd.n4875 gnd.n4874 585
R2648 gnd.n1536 gnd.n1535 585
R2649 gnd.n1544 gnd.n1536 585
R2650 gnd.n4778 gnd.n1543 585
R2651 gnd.n4867 gnd.n1543 585
R2652 gnd.n4781 gnd.n4780 585
R2653 gnd.n4780 gnd.n4779 585
R2654 gnd.n4782 gnd.n1554 585
R2655 gnd.n4856 gnd.n1554 585
R2656 gnd.n4784 gnd.n4783 585
R2657 gnd.n4783 gnd.n1552 585
R2658 gnd.n4785 gnd.n1560 585
R2659 gnd.n4850 gnd.n1560 585
R2660 gnd.n4790 gnd.n4789 585
R2661 gnd.n4789 gnd.n4788 585
R2662 gnd.n4791 gnd.n1568 585
R2663 gnd.n4827 gnd.n1568 585
R2664 gnd.n4793 gnd.n4792 585
R2665 gnd.n4792 gnd.n1567 585
R2666 gnd.n4794 gnd.n1574 585
R2667 gnd.n4821 gnd.n1574 585
R2668 gnd.n4797 gnd.n4796 585
R2669 gnd.n4796 gnd.n4795 585
R2670 gnd.n4798 gnd.n1583 585
R2671 gnd.n4809 gnd.n1583 585
R2672 gnd.n4800 gnd.n4799 585
R2673 gnd.n4801 gnd.n4800 585
R2674 gnd.n4777 gnd.n1589 585
R2675 gnd.n4803 gnd.n1589 585
R2676 gnd.n4776 gnd.n4775 585
R2677 gnd.n4775 gnd.n4774 585
R2678 gnd.n1591 gnd.n1590 585
R2679 gnd.n4758 gnd.n1591 585
R2680 gnd.n4755 gnd.n4754 585
R2681 gnd.n4756 gnd.n4755 585
R2682 gnd.n4753 gnd.n1600 585
R2683 gnd.n4764 gnd.n1600 585
R2684 gnd.n4752 gnd.n4751 585
R2685 gnd.n4751 gnd.n4750 585
R2686 gnd.n1606 gnd.n1605 585
R2687 gnd.n4748 gnd.n1606 585
R2688 gnd.n4726 gnd.n4725 585
R2689 gnd.n4725 gnd.n1613 585
R2690 gnd.n4727 gnd.n1611 585
R2691 gnd.n4742 gnd.n1611 585
R2692 gnd.n4729 gnd.n4728 585
R2693 gnd.n4730 gnd.n4729 585
R2694 gnd.n4724 gnd.n1621 585
R2695 gnd.n1621 gnd.n1619 585
R2696 gnd.n4723 gnd.n4722 585
R2697 gnd.n4722 gnd.n4721 585
R2698 gnd.n1623 gnd.n1622 585
R2699 gnd.n1633 gnd.n1623 585
R2700 gnd.n4601 gnd.n1632 585
R2701 gnd.n4714 gnd.n1632 585
R2702 gnd.n4604 gnd.n4603 585
R2703 gnd.n4603 gnd.n4602 585
R2704 gnd.n4605 gnd.n1642 585
R2705 gnd.n4703 gnd.n1642 585
R2706 gnd.n4607 gnd.n4606 585
R2707 gnd.n4606 gnd.n1640 585
R2708 gnd.n4608 gnd.n1648 585
R2709 gnd.n4697 gnd.n1648 585
R2710 gnd.n4612 gnd.n4611 585
R2711 gnd.n4611 gnd.n4610 585
R2712 gnd.n4613 gnd.n1655 585
R2713 gnd.n4650 gnd.n1655 585
R2714 gnd.n4615 gnd.n4614 585
R2715 gnd.n4614 gnd.n1661 585
R2716 gnd.n4616 gnd.n1660 585
R2717 gnd.n4644 gnd.n1660 585
R2718 gnd.n4620 gnd.n4619 585
R2719 gnd.n4619 gnd.n4618 585
R2720 gnd.n4621 gnd.n1669 585
R2721 gnd.n4632 gnd.n1669 585
R2722 gnd.n4623 gnd.n4622 585
R2723 gnd.n4624 gnd.n4623 585
R2724 gnd.n4600 gnd.n1676 585
R2725 gnd.n4626 gnd.n1676 585
R2726 gnd.n4599 gnd.n4598 585
R2727 gnd.n4598 gnd.n4597 585
R2728 gnd.n1678 gnd.n1677 585
R2729 gnd.n4581 gnd.n1678 585
R2730 gnd.n4532 gnd.n4531 585
R2731 gnd.n4531 gnd.n4530 585
R2732 gnd.n4533 gnd.n1685 585
R2733 gnd.n4587 gnd.n1685 585
R2734 gnd.n4536 gnd.n4535 585
R2735 gnd.n4535 gnd.n4534 585
R2736 gnd.n4537 gnd.n1698 585
R2737 gnd.n4563 gnd.n1698 585
R2738 gnd.n4539 gnd.n4538 585
R2739 gnd.n4538 gnd.n1704 585
R2740 gnd.n4540 gnd.n1703 585
R2741 gnd.n4557 gnd.n1703 585
R2742 gnd.n4542 gnd.n4541 585
R2743 gnd.n4544 gnd.n4542 585
R2744 gnd.n4529 gnd.n1712 585
R2745 gnd.n1712 gnd.n1710 585
R2746 gnd.n4528 gnd.n4527 585
R2747 gnd.n4527 gnd.n4526 585
R2748 gnd.n1714 gnd.n1713 585
R2749 gnd.n1723 gnd.n1714 585
R2750 gnd.n4427 gnd.n1722 585
R2751 gnd.n4519 gnd.n1722 585
R2752 gnd.n4430 gnd.n4429 585
R2753 gnd.n4429 gnd.n4428 585
R2754 gnd.n4431 gnd.n1732 585
R2755 gnd.n4507 gnd.n1732 585
R2756 gnd.n4433 gnd.n4432 585
R2757 gnd.n4432 gnd.n1730 585
R2758 gnd.n4434 gnd.n1738 585
R2759 gnd.n4501 gnd.n1738 585
R2760 gnd.n4438 gnd.n4437 585
R2761 gnd.n4437 gnd.n4436 585
R2762 gnd.n4439 gnd.n1746 585
R2763 gnd.n4477 gnd.n1746 585
R2764 gnd.n4441 gnd.n4440 585
R2765 gnd.n4440 gnd.n1745 585
R2766 gnd.n4442 gnd.n1751 585
R2767 gnd.n4471 gnd.n1751 585
R2768 gnd.n4446 gnd.n4445 585
R2769 gnd.n4445 gnd.n4444 585
R2770 gnd.n4447 gnd.n1759 585
R2771 gnd.n4458 gnd.n1759 585
R2772 gnd.n4449 gnd.n4448 585
R2773 gnd.n4450 gnd.n4449 585
R2774 gnd.n4426 gnd.n1765 585
R2775 gnd.n4452 gnd.n1765 585
R2776 gnd.n4425 gnd.n4424 585
R2777 gnd.n4424 gnd.n4423 585
R2778 gnd.n6093 gnd.n6092 585
R2779 gnd.n6092 gnd.n6091 585
R2780 gnd.n6894 gnd.n6893 585
R2781 gnd.n6893 gnd.n168 585
R2782 gnd.n6897 gnd.n277 585
R2783 gnd.n277 gnd.n177 585
R2784 gnd.n6899 gnd.n6898 585
R2785 gnd.n6899 gnd.n188 585
R2786 gnd.n6900 gnd.n276 585
R2787 gnd.n6900 gnd.n186 585
R2788 gnd.n6902 gnd.n6901 585
R2789 gnd.n6901 gnd.n196 585
R2790 gnd.n6903 gnd.n271 585
R2791 gnd.n271 gnd.n194 585
R2792 gnd.n6905 gnd.n6904 585
R2793 gnd.n6906 gnd.n6905 585
R2794 gnd.n272 gnd.n270 585
R2795 gnd.n270 gnd.n202 585
R2796 gnd.n5796 gnd.n5795 585
R2797 gnd.n5796 gnd.n211 585
R2798 gnd.n5798 gnd.n5797 585
R2799 gnd.n5797 gnd.n209 585
R2800 gnd.n5799 gnd.n5789 585
R2801 gnd.n5789 gnd.n225 585
R2802 gnd.n5801 gnd.n5800 585
R2803 gnd.n5801 gnd.n223 585
R2804 gnd.n5802 gnd.n5788 585
R2805 gnd.n5802 gnd.n233 585
R2806 gnd.n5804 gnd.n5803 585
R2807 gnd.n5803 gnd.n231 585
R2808 gnd.n5806 gnd.n1172 585
R2809 gnd.n1172 gnd.n235 585
R2810 gnd.n5808 gnd.n5807 585
R2811 gnd.n5809 gnd.n5808 585
R2812 gnd.n5786 gnd.n1171 585
R2813 gnd.n1180 gnd.n1171 585
R2814 gnd.n5785 gnd.n5784 585
R2815 gnd.n5784 gnd.n5783 585
R2816 gnd.n5748 gnd.n1174 585
R2817 gnd.n5772 gnd.n1174 585
R2818 gnd.n5750 gnd.n5749 585
R2819 gnd.n5750 gnd.n1184 585
R2820 gnd.n5752 gnd.n5751 585
R2821 gnd.n5751 gnd.n1196 585
R2822 gnd.n5753 gnd.n1207 585
R2823 gnd.n1207 gnd.n1194 585
R2824 gnd.n5755 gnd.n5754 585
R2825 gnd.n5756 gnd.n5755 585
R2826 gnd.n1208 gnd.n1206 585
R2827 gnd.n1206 gnd.n1201 585
R2828 gnd.n5742 gnd.n5741 585
R2829 gnd.n5741 gnd.n5740 585
R2830 gnd.n1211 gnd.n1210 585
R2831 gnd.n1222 gnd.n1211 585
R2832 gnd.n5715 gnd.n1235 585
R2833 gnd.n1235 gnd.n1220 585
R2834 gnd.n5717 gnd.n5716 585
R2835 gnd.n5718 gnd.n5717 585
R2836 gnd.n1236 gnd.n1234 585
R2837 gnd.n1234 gnd.n1230 585
R2838 gnd.n5710 gnd.n5709 585
R2839 gnd.n5709 gnd.n5708 585
R2840 gnd.n1239 gnd.n1238 585
R2841 gnd.n1251 gnd.n1239 585
R2842 gnd.n5684 gnd.n5672 585
R2843 gnd.n5672 gnd.n1249 585
R2844 gnd.n5686 gnd.n5685 585
R2845 gnd.n5687 gnd.n5686 585
R2846 gnd.n5673 gnd.n5671 585
R2847 gnd.n5671 gnd.n1256 585
R2848 gnd.n5679 gnd.n5678 585
R2849 gnd.n5678 gnd.n1141 585
R2850 gnd.n5677 gnd.n5676 585
R2851 gnd.n5677 gnd.n1138 585
R2852 gnd.n1125 gnd.n1124 585
R2853 gnd.n1129 gnd.n1125 585
R2854 gnd.n5854 gnd.n5853 585
R2855 gnd.n5853 gnd.n5852 585
R2856 gnd.n5855 gnd.n1119 585
R2857 gnd.n1126 gnd.n1119 585
R2858 gnd.n5857 gnd.n5856 585
R2859 gnd.n5858 gnd.n5857 585
R2860 gnd.n1116 gnd.n1115 585
R2861 gnd.n5859 gnd.n1116 585
R2862 gnd.n5862 gnd.n5861 585
R2863 gnd.n5861 gnd.n5860 585
R2864 gnd.n5863 gnd.n1110 585
R2865 gnd.n1110 gnd.n1108 585
R2866 gnd.n5865 gnd.n5864 585
R2867 gnd.n5866 gnd.n5865 585
R2868 gnd.n1111 gnd.n1109 585
R2869 gnd.n1109 gnd.n1106 585
R2870 gnd.n5329 gnd.n1349 585
R2871 gnd.n5329 gnd.n5328 585
R2872 gnd.n5331 gnd.n5330 585
R2873 gnd.n5330 gnd.n1296 585
R2874 gnd.n5332 gnd.n1342 585
R2875 gnd.n1342 gnd.n1333 585
R2876 gnd.n5334 gnd.n5333 585
R2877 gnd.n5335 gnd.n5334 585
R2878 gnd.n1343 gnd.n1341 585
R2879 gnd.n1425 gnd.n1341 585
R2880 gnd.n5119 gnd.n1371 585
R2881 gnd.n1424 gnd.n1371 585
R2882 gnd.n5121 gnd.n5120 585
R2883 gnd.n5122 gnd.n5121 585
R2884 gnd.n1372 gnd.n1370 585
R2885 gnd.n1370 gnd.n1367 585
R2886 gnd.n5113 gnd.n5112 585
R2887 gnd.n5112 gnd.n5111 585
R2888 gnd.n1375 gnd.n1374 585
R2889 gnd.n5099 gnd.n1375 585
R2890 gnd.n5089 gnd.n5088 585
R2891 gnd.n5090 gnd.n5089 585
R2892 gnd.n1393 gnd.n1392 585
R2893 gnd.n1441 gnd.n1392 585
R2894 gnd.n5084 gnd.n5083 585
R2895 gnd.n5083 gnd.n5082 585
R2896 gnd.n1396 gnd.n1395 585
R2897 gnd.n1403 gnd.n1396 585
R2898 gnd.n5046 gnd.n5045 585
R2899 gnd.n5047 gnd.n5046 585
R2900 gnd.n1450 gnd.n1449 585
R2901 gnd.n1449 gnd.n1412 585
R2902 gnd.n5041 gnd.n5040 585
R2903 gnd.n5040 gnd.n1417 585
R2904 gnd.n5039 gnd.n1452 585
R2905 gnd.n5039 gnd.n5038 585
R2906 gnd.n5019 gnd.n1453 585
R2907 gnd.n1459 gnd.n1453 585
R2908 gnd.n5021 gnd.n5020 585
R2909 gnd.n5022 gnd.n5021 585
R2910 gnd.n1468 gnd.n1467 585
R2911 gnd.n1475 gnd.n1467 585
R2912 gnd.n5014 gnd.n5013 585
R2913 gnd.n5013 gnd.n5012 585
R2914 gnd.n1471 gnd.n1470 585
R2915 gnd.n1479 gnd.n1471 585
R2916 gnd.n4968 gnd.n1495 585
R2917 gnd.n1495 gnd.n1489 585
R2918 gnd.n4970 gnd.n4969 585
R2919 gnd.n4971 gnd.n4970 585
R2920 gnd.n1496 gnd.n1494 585
R2921 gnd.n4945 gnd.n1494 585
R2922 gnd.n4963 gnd.n4962 585
R2923 gnd.n4962 gnd.n4961 585
R2924 gnd.n1499 gnd.n1498 585
R2925 gnd.n4953 gnd.n1499 585
R2926 gnd.n4898 gnd.n4897 585
R2927 gnd.n4897 gnd.n4896 585
R2928 gnd.n4899 gnd.n1527 585
R2929 gnd.n1527 gnd.n1518 585
R2930 gnd.n4901 gnd.n4900 585
R2931 gnd.n4902 gnd.n4901 585
R2932 gnd.n1528 gnd.n1526 585
R2933 gnd.n1526 gnd.n1523 585
R2934 gnd.n4888 gnd.n4887 585
R2935 gnd.n4887 gnd.n4886 585
R2936 gnd.n1531 gnd.n1530 585
R2937 gnd.n1537 gnd.n1531 585
R2938 gnd.n4865 gnd.n4864 585
R2939 gnd.n4866 gnd.n4865 585
R2940 gnd.n1548 gnd.n1547 585
R2941 gnd.n1555 gnd.n1547 585
R2942 gnd.n4860 gnd.n4859 585
R2943 gnd.n4859 gnd.n4858 585
R2944 gnd.n1551 gnd.n1550 585
R2945 gnd.n1559 gnd.n1551 585
R2946 gnd.n4817 gnd.n1576 585
R2947 gnd.n1576 gnd.n1569 585
R2948 gnd.n4819 gnd.n4818 585
R2949 gnd.n4820 gnd.n4819 585
R2950 gnd.n1577 gnd.n1575 585
R2951 gnd.n1575 gnd.n1573 585
R2952 gnd.n4812 gnd.n4811 585
R2953 gnd.n4811 gnd.n4810 585
R2954 gnd.n1580 gnd.n1579 585
R2955 gnd.n4802 gnd.n1580 585
R2956 gnd.n4772 gnd.n4771 585
R2957 gnd.n4773 gnd.n4772 585
R2958 gnd.n1594 gnd.n1593 585
R2959 gnd.n4757 gnd.n1593 585
R2960 gnd.n4767 gnd.n4766 585
R2961 gnd.n4766 gnd.n4765 585
R2962 gnd.n1597 gnd.n1596 585
R2963 gnd.n4749 gnd.n1597 585
R2964 gnd.n4739 gnd.n4738 585
R2965 gnd.n4740 gnd.n4739 585
R2966 gnd.n1615 gnd.n1614 585
R2967 gnd.n1614 gnd.n1610 585
R2968 gnd.n4734 gnd.n4733 585
R2969 gnd.n4733 gnd.n4732 585
R2970 gnd.n1618 gnd.n1617 585
R2971 gnd.n1624 gnd.n1618 585
R2972 gnd.n4712 gnd.n4711 585
R2973 gnd.n4713 gnd.n4712 585
R2974 gnd.n1636 gnd.n1635 585
R2975 gnd.n1643 gnd.n1635 585
R2976 gnd.n4707 gnd.n4706 585
R2977 gnd.n4706 gnd.n4705 585
R2978 gnd.n1639 gnd.n1638 585
R2979 gnd.n1647 gnd.n1639 585
R2980 gnd.n4640 gnd.n1663 585
R2981 gnd.n1663 gnd.n1656 585
R2982 gnd.n4642 gnd.n4641 585
R2983 gnd.n4643 gnd.n4642 585
R2984 gnd.n1664 gnd.n1662 585
R2985 gnd.n4617 gnd.n1662 585
R2986 gnd.n4635 gnd.n4634 585
R2987 gnd.n4634 gnd.n4633 585
R2988 gnd.n1667 gnd.n1666 585
R2989 gnd.n4625 gnd.n1667 585
R2990 gnd.n4595 gnd.n4594 585
R2991 gnd.n4596 gnd.n4595 585
R2992 gnd.n1680 gnd.n1679 585
R2993 gnd.n1690 gnd.n1679 585
R2994 gnd.n4590 gnd.n4589 585
R2995 gnd.n4589 gnd.n4588 585
R2996 gnd.n1683 gnd.n1682 585
R2997 gnd.n1699 gnd.n1683 585
R2998 gnd.n4554 gnd.n4553 585
R2999 gnd.n4555 gnd.n4554 585
R3000 gnd.n1706 gnd.n1705 585
R3001 gnd.n4543 gnd.n1705 585
R3002 gnd.n4549 gnd.n4548 585
R3003 gnd.n4548 gnd.n4547 585
R3004 gnd.n1709 gnd.n1708 585
R3005 gnd.n1715 gnd.n1709 585
R3006 gnd.n4517 gnd.n4516 585
R3007 gnd.n4518 gnd.n4517 585
R3008 gnd.n1726 gnd.n1725 585
R3009 gnd.n1733 gnd.n1725 585
R3010 gnd.n4512 gnd.n4511 585
R3011 gnd.n4511 gnd.n4510 585
R3012 gnd.n1729 gnd.n1728 585
R3013 gnd.n1737 gnd.n1729 585
R3014 gnd.n4466 gnd.n1753 585
R3015 gnd.n1753 gnd.n1747 585
R3016 gnd.n4468 gnd.n4467 585
R3017 gnd.n4469 gnd.n4468 585
R3018 gnd.n1754 gnd.n1752 585
R3019 gnd.n4443 gnd.n1752 585
R3020 gnd.n4461 gnd.n4460 585
R3021 gnd.n4460 gnd.n4459 585
R3022 gnd.n1757 gnd.n1756 585
R3023 gnd.n4451 gnd.n1757 585
R3024 gnd.n4421 gnd.n4420 585
R3025 gnd.n4422 gnd.n4421 585
R3026 gnd.n1769 gnd.n1768 585
R3027 gnd.n1807 gnd.n1768 585
R3028 gnd.n4416 gnd.n4415 585
R3029 gnd.n4415 gnd.n4414 585
R3030 gnd.n1772 gnd.n1771 585
R3031 gnd.n4254 gnd.n1772 585
R3032 gnd.n4252 gnd.n4251 585
R3033 gnd.n4253 gnd.n4252 585
R3034 gnd.n2022 gnd.n2021 585
R3035 gnd.n2021 gnd.n2020 585
R3036 gnd.n4247 gnd.n4246 585
R3037 gnd.n4246 gnd.n4245 585
R3038 gnd.n2025 gnd.n2024 585
R3039 gnd.n4112 gnd.n2025 585
R3040 gnd.n4110 gnd.n4109 585
R3041 gnd.n4111 gnd.n4110 585
R3042 gnd.n2028 gnd.n2027 585
R3043 gnd.n2027 gnd.n2026 585
R3044 gnd.n4105 gnd.n4104 585
R3045 gnd.n4104 gnd.n996 585
R3046 gnd.n4103 gnd.n2030 585
R3047 gnd.n4103 gnd.n993 585
R3048 gnd.n4102 gnd.n4101 585
R3049 gnd.n4102 gnd.n986 585
R3050 gnd.n2032 gnd.n2031 585
R3051 gnd.n2031 gnd.n983 585
R3052 gnd.n4097 gnd.n4096 585
R3053 gnd.n4096 gnd.n975 585
R3054 gnd.n4095 gnd.n2034 585
R3055 gnd.n4095 gnd.n972 585
R3056 gnd.n4094 gnd.n4093 585
R3057 gnd.n4094 gnd.n964 585
R3058 gnd.n2036 gnd.n2035 585
R3059 gnd.n4047 gnd.n2035 585
R3060 gnd.n4089 gnd.n4088 585
R3061 gnd.n4088 gnd.n954 585
R3062 gnd.n4087 gnd.n2038 585
R3063 gnd.n4087 gnd.n951 585
R3064 gnd.n4086 gnd.n4085 585
R3065 gnd.n4086 gnd.n943 585
R3066 gnd.n2040 gnd.n2039 585
R3067 gnd.n2039 gnd.n940 585
R3068 gnd.n4081 gnd.n4080 585
R3069 gnd.n4080 gnd.n4079 585
R3070 gnd.n2043 gnd.n2042 585
R3071 gnd.n2043 gnd.n930 585
R3072 gnd.n4021 gnd.n2066 585
R3073 gnd.n2066 gnd.n923 585
R3074 gnd.n4023 gnd.n4022 585
R3075 gnd.n4024 gnd.n4023 585
R3076 gnd.n4017 gnd.n2065 585
R3077 gnd.n2065 gnd.n912 585
R3078 gnd.n4016 gnd.n4015 585
R3079 gnd.n4015 gnd.n909 585
R3080 gnd.n4014 gnd.n2069 585
R3081 gnd.n4014 gnd.n4013 585
R3082 gnd.n3955 gnd.n2068 585
R3083 gnd.n2079 gnd.n2068 585
R3084 gnd.n3958 gnd.n3957 585
R3085 gnd.n3958 gnd.n2077 585
R3086 gnd.n3960 gnd.n3959 585
R3087 gnd.n3959 gnd.n2084 585
R3088 gnd.n3962 gnd.n2114 585
R3089 gnd.n2114 gnd.n2105 585
R3090 gnd.n3964 gnd.n3963 585
R3091 gnd.n3965 gnd.n3964 585
R3092 gnd.n3953 gnd.n2113 585
R3093 gnd.n2113 gnd.n2111 585
R3094 gnd.n3952 gnd.n3951 585
R3095 gnd.n3951 gnd.n3950 585
R3096 gnd.n3924 gnd.n2116 585
R3097 gnd.n2116 gnd.n894 585
R3098 gnd.n3925 gnd.n2125 585
R3099 gnd.n2125 gnd.n886 585
R3100 gnd.n3927 gnd.n3926 585
R3101 gnd.n3928 gnd.n3927 585
R3102 gnd.n2126 gnd.n2124 585
R3103 gnd.n2124 gnd.n876 585
R3104 gnd.n3919 gnd.n3918 585
R3105 gnd.n3918 gnd.n873 585
R3106 gnd.n3917 gnd.n2128 585
R3107 gnd.n3917 gnd.n865 585
R3108 gnd.n3916 gnd.n3915 585
R3109 gnd.n3916 gnd.n862 585
R3110 gnd.n3904 gnd.n3903 585
R3111 gnd.n3903 gnd.n3902 585
R3112 gnd.n3911 gnd.n3910 585
R3113 gnd.n3910 gnd.n852 585
R3114 gnd.n3909 gnd.n3908 585
R3115 gnd.n3909 gnd.n843 585
R3116 gnd.n3907 gnd.n826 585
R3117 gnd.n840 gnd.n826 585
R3118 gnd.n5869 gnd.n5868 585
R3119 gnd.n5868 gnd.n5867 585
R3120 gnd.n5870 gnd.n1103 585
R3121 gnd.n5327 gnd.n1103 585
R3122 gnd.n5871 gnd.n1102 585
R3123 gnd.n1350 gnd.n1102 585
R3124 gnd.n5142 gnd.n1100 585
R3125 gnd.n5143 gnd.n5142 585
R3126 gnd.n5875 gnd.n1099 585
R3127 gnd.n5140 gnd.n1099 585
R3128 gnd.n5876 gnd.n1098 585
R3129 gnd.n1338 gnd.n1098 585
R3130 gnd.n5877 gnd.n1097 585
R3131 gnd.n1427 gnd.n1097 585
R3132 gnd.n1362 gnd.n1095 585
R3133 gnd.n5132 gnd.n1362 585
R3134 gnd.n5881 gnd.n1094 585
R3135 gnd.n5124 gnd.n1094 585
R3136 gnd.n5882 gnd.n1093 585
R3137 gnd.n5109 gnd.n1093 585
R3138 gnd.n5883 gnd.n1092 585
R3139 gnd.n1385 gnd.n1092 585
R3140 gnd.n5100 gnd.n1090 585
R3141 gnd.n5101 gnd.n5100 585
R3142 gnd.n5887 gnd.n1089 585
R3143 gnd.n1390 gnd.n1089 585
R3144 gnd.n5888 gnd.n1088 585
R3145 gnd.n1399 gnd.n1088 585
R3146 gnd.n5889 gnd.n1087 585
R3147 gnd.n5074 gnd.n1087 585
R3148 gnd.n5048 gnd.n1085 585
R3149 gnd.n5049 gnd.n5048 585
R3150 gnd.n5893 gnd.n1084 585
R3151 gnd.n5065 gnd.n1084 585
R3152 gnd.n5894 gnd.n1083 585
R3153 gnd.n5057 gnd.n1083 585
R3154 gnd.n5895 gnd.n1082 585
R3155 gnd.n5037 gnd.n1082 585
R3156 gnd.n1460 gnd.n1080 585
R3157 gnd.t178 gnd.n1460 585
R3158 gnd.n5899 gnd.n1079 585
R3159 gnd.n4988 gnd.n1079 585
R3160 gnd.n5900 gnd.n1078 585
R3161 gnd.n1465 gnd.n1078 585
R3162 gnd.n5901 gnd.n1077 585
R3163 gnd.n5011 gnd.n1077 585
R3164 gnd.n5002 gnd.n1075 585
R3165 gnd.n5003 gnd.n5002 585
R3166 gnd.n5905 gnd.n1074 585
R3167 gnd.n4938 gnd.n1074 585
R3168 gnd.n5906 gnd.n1073 585
R3169 gnd.n4980 gnd.n1073 585
R3170 gnd.n5907 gnd.n1072 585
R3171 gnd.n4972 gnd.n1072 585
R3172 gnd.n1502 gnd.n1070 585
R3173 gnd.n1503 gnd.n1502 585
R3174 gnd.n5911 gnd.n1069 585
R3175 gnd.n1500 gnd.n1069 585
R3176 gnd.n5912 gnd.n1068 585
R3177 gnd.n4925 gnd.n1068 585
R3178 gnd.n5913 gnd.n1067 585
R3179 gnd.n4895 gnd.n1067 585
R3180 gnd.n4912 gnd.n1065 585
R3181 gnd.n4913 gnd.n4912 585
R3182 gnd.n5917 gnd.n1064 585
R3183 gnd.n4903 gnd.n1064 585
R3184 gnd.n5918 gnd.n1063 585
R3185 gnd.n4885 gnd.n1063 585
R3186 gnd.n5919 gnd.n1062 585
R3187 gnd.n4836 gnd.n1062 585
R3188 gnd.n1545 gnd.n1060 585
R3189 gnd.n1546 gnd.n1545 585
R3190 gnd.n5923 gnd.n1059 585
R3191 gnd.n1542 gnd.n1059 585
R3192 gnd.n5924 gnd.n1058 585
R3193 gnd.n4857 gnd.n1058 585
R3194 gnd.n5925 gnd.n1057 585
R3195 gnd.n4849 gnd.n1057 585
R3196 gnd.n4786 gnd.n1055 585
R3197 gnd.n4787 gnd.n4786 585
R3198 gnd.n5929 gnd.n1054 585
R3199 gnd.n4828 gnd.n1054 585
R3200 gnd.n5930 gnd.n1053 585
R3201 gnd.n4821 gnd.n1053 585
R3202 gnd.n5931 gnd.n1052 585
R3203 gnd.n1584 gnd.n1052 585
R3204 gnd.n1581 gnd.n1050 585
R3205 gnd.n1582 gnd.n1581 585
R3206 gnd.n5935 gnd.n1049 585
R3207 gnd.n1588 gnd.n1049 585
R3208 gnd.n5936 gnd.n1048 585
R3209 gnd.n1592 gnd.n1048 585
R3210 gnd.n5937 gnd.n1047 585
R3211 gnd.n1601 gnd.n1047 585
R3212 gnd.n1598 gnd.n1045 585
R3213 gnd.n1599 gnd.n1598 585
R3214 gnd.n5941 gnd.n1044 585
R3215 gnd.n4662 gnd.n1044 585
R3216 gnd.n5942 gnd.n1043 585
R3217 gnd.n4741 gnd.n1043 585
R3218 gnd.n5943 gnd.n1042 585
R3219 gnd.n4731 gnd.n1042 585
R3220 gnd.n1625 gnd.n1040 585
R3221 gnd.n1626 gnd.n1625 585
R3222 gnd.n5947 gnd.n1039 585
R3223 gnd.n1634 gnd.n1039 585
R3224 gnd.n5948 gnd.n1038 585
R3225 gnd.n1631 gnd.n1038 585
R3226 gnd.n5949 gnd.n1037 585
R3227 gnd.n4704 gnd.n1037 585
R3228 gnd.n4695 gnd.n1035 585
R3229 gnd.n4696 gnd.n4695 585
R3230 gnd.n5953 gnd.n1034 585
R3231 gnd.n4609 gnd.n1034 585
R3232 gnd.n5954 gnd.n1033 585
R3233 gnd.n4651 gnd.n1033 585
R3234 gnd.n5955 gnd.n1032 585
R3235 gnd.n4644 gnd.n1032 585
R3236 gnd.n1670 gnd.n1030 585
R3237 gnd.n1671 gnd.n1670 585
R3238 gnd.n5959 gnd.n1029 585
R3239 gnd.n1668 gnd.n1029 585
R3240 gnd.n5960 gnd.n1028 585
R3241 gnd.n1675 gnd.n1028 585
R3242 gnd.n5961 gnd.n1027 585
R3243 gnd.n4580 gnd.n1027 585
R3244 gnd.n1686 gnd.n1025 585
R3245 gnd.t174 gnd.n1686 585
R3246 gnd.n5965 gnd.n1024 585
R3247 gnd.n1684 gnd.n1024 585
R3248 gnd.n5966 gnd.n1023 585
R3249 gnd.n4564 gnd.n1023 585
R3250 gnd.n5967 gnd.n1022 585
R3251 gnd.n4556 gnd.n1022 585
R3252 gnd.n4545 gnd.n1020 585
R3253 gnd.n4546 gnd.n4545 585
R3254 gnd.n5971 gnd.n1019 585
R3255 gnd.n1716 gnd.n1019 585
R3256 gnd.n5972 gnd.n1018 585
R3257 gnd.n1724 gnd.n1018 585
R3258 gnd.n5973 gnd.n1017 585
R3259 gnd.n1721 gnd.n1017 585
R3260 gnd.n4508 gnd.n1015 585
R3261 gnd.n4509 gnd.n4508 585
R3262 gnd.n5977 gnd.n1014 585
R3263 gnd.n4500 gnd.n1014 585
R3264 gnd.n5978 gnd.n1013 585
R3265 gnd.n4435 gnd.n1013 585
R3266 gnd.n5979 gnd.n1012 585
R3267 gnd.n4478 gnd.n1012 585
R3268 gnd.n4470 gnd.n1010 585
R3269 gnd.n4471 gnd.n4470 585
R3270 gnd.n5983 gnd.n1009 585
R3271 gnd.n1760 gnd.n1009 585
R3272 gnd.n5984 gnd.n1008 585
R3273 gnd.n1758 gnd.n1008 585
R3274 gnd.n5985 gnd.n1007 585
R3275 gnd.n1764 gnd.n1007 585
R3276 gnd.n4260 gnd.n1005 585
R3277 gnd.n4261 gnd.n4260 585
R3278 gnd.n5989 gnd.n1004 585
R3279 gnd.n4413 gnd.n1004 585
R3280 gnd.n5990 gnd.n1003 585
R3281 gnd.n1773 gnd.n1003 585
R3282 gnd.n5991 gnd.n1002 585
R3283 gnd.n4255 gnd.n1002 585
R3284 gnd.n4242 gnd.n4241 585
R3285 gnd.n4240 gnd.n4128 585
R3286 gnd.n4130 gnd.n4127 585
R3287 gnd.n4244 gnd.n4127 585
R3288 gnd.n4233 gnd.n4143 585
R3289 gnd.n4232 gnd.n4144 585
R3290 gnd.n4146 gnd.n4145 585
R3291 gnd.n4225 gnd.n4154 585
R3292 gnd.n4224 gnd.n4155 585
R3293 gnd.n4165 gnd.n4156 585
R3294 gnd.n4217 gnd.n4166 585
R3295 gnd.n4216 gnd.n4167 585
R3296 gnd.n4169 gnd.n4168 585
R3297 gnd.n4209 gnd.n4177 585
R3298 gnd.n4208 gnd.n4178 585
R3299 gnd.n4190 gnd.n4179 585
R3300 gnd.n4201 gnd.n4191 585
R3301 gnd.n4200 gnd.n4193 585
R3302 gnd.n4192 gnd.n2001 585
R3303 gnd.n4292 gnd.n2002 585
R3304 gnd.n4291 gnd.n2003 585
R3305 gnd.n4290 gnd.n2004 585
R3306 gnd.n4122 gnd.n2005 585
R3307 gnd.n4286 gnd.n2007 585
R3308 gnd.n4285 gnd.n2008 585
R3309 gnd.n4284 gnd.n2009 585
R3310 gnd.n4281 gnd.n2014 585
R3311 gnd.n4280 gnd.n2015 585
R3312 gnd.n4279 gnd.n2016 585
R3313 gnd.n2019 gnd.n2017 585
R3314 gnd.n1353 gnd.n1107 585
R3315 gnd.n5867 gnd.n1107 585
R3316 gnd.n5326 gnd.n5325 585
R3317 gnd.n5327 gnd.n5326 585
R3318 gnd.n1352 gnd.n1351 585
R3319 gnd.n1351 gnd.n1350 585
R3320 gnd.n5145 gnd.n5144 585
R3321 gnd.n5144 gnd.n5143 585
R3322 gnd.n5141 gnd.n1355 585
R3323 gnd.n5141 gnd.n5140 585
R3324 gnd.n5139 gnd.n5138 585
R3325 gnd.n5139 gnd.n1338 585
R3326 gnd.n1357 gnd.n1356 585
R3327 gnd.n1427 gnd.n1356 585
R3328 gnd.n5134 gnd.n5133 585
R3329 gnd.n5133 gnd.n5132 585
R3330 gnd.n1360 gnd.n1359 585
R3331 gnd.n5124 gnd.n1360 585
R3332 gnd.n5108 gnd.n5107 585
R3333 gnd.n5109 gnd.n5108 585
R3334 gnd.n1379 gnd.n1378 585
R3335 gnd.n1385 gnd.n1378 585
R3336 gnd.n5103 gnd.n5102 585
R3337 gnd.n5102 gnd.n5101 585
R3338 gnd.n1382 gnd.n1381 585
R3339 gnd.n1390 gnd.n1382 585
R3340 gnd.n1408 gnd.n1406 585
R3341 gnd.n1406 gnd.n1399 585
R3342 gnd.n5073 gnd.n5072 585
R3343 gnd.n5074 gnd.n5073 585
R3344 gnd.n1407 gnd.n1405 585
R3345 gnd.n5049 gnd.n1405 585
R3346 gnd.n5067 gnd.n5066 585
R3347 gnd.n5066 gnd.n5065 585
R3348 gnd.n1411 gnd.n1410 585
R3349 gnd.n5057 gnd.n1411 585
R3350 gnd.n4991 gnd.n1455 585
R3351 gnd.n5037 gnd.n1455 585
R3352 gnd.n4994 gnd.n4990 585
R3353 gnd.n4990 gnd.t178 585
R3354 gnd.n4995 gnd.n4989 585
R3355 gnd.n4989 gnd.n4988 585
R3356 gnd.n4996 gnd.n4986 585
R3357 gnd.n4986 gnd.n1465 585
R3358 gnd.n1483 gnd.n1473 585
R3359 gnd.n5011 gnd.n1473 585
R3360 gnd.n5001 gnd.n5000 585
R3361 gnd.n5003 gnd.n5001 585
R3362 gnd.n1482 gnd.n1481 585
R3363 gnd.n4938 gnd.n1481 585
R3364 gnd.n4982 gnd.n4981 585
R3365 gnd.n4981 gnd.n4980 585
R3366 gnd.n1486 gnd.n1485 585
R3367 gnd.n4972 gnd.n1486 585
R3368 gnd.n4919 gnd.n4918 585
R3369 gnd.n4918 gnd.n1503 585
R3370 gnd.n1513 gnd.n1511 585
R3371 gnd.n1511 gnd.n1500 585
R3372 gnd.n4924 gnd.n4923 585
R3373 gnd.n4925 gnd.n4924 585
R3374 gnd.n1512 gnd.n1510 585
R3375 gnd.n4895 gnd.n1510 585
R3376 gnd.n4915 gnd.n4914 585
R3377 gnd.n4914 gnd.n4913 585
R3378 gnd.n1516 gnd.n1515 585
R3379 gnd.n4903 gnd.n1516 585
R3380 gnd.n4838 gnd.n1533 585
R3381 gnd.n4885 gnd.n1533 585
R3382 gnd.n4841 gnd.n4837 585
R3383 gnd.n4837 gnd.n4836 585
R3384 gnd.n4842 gnd.n4835 585
R3385 gnd.n4835 gnd.n1546 585
R3386 gnd.n4843 gnd.n4834 585
R3387 gnd.n4834 gnd.n1542 585
R3388 gnd.n1563 gnd.n1553 585
R3389 gnd.n4857 gnd.n1553 585
R3390 gnd.n4848 gnd.n4847 585
R3391 gnd.n4849 gnd.n4848 585
R3392 gnd.n1562 gnd.n1561 585
R3393 gnd.n4787 gnd.n1561 585
R3394 gnd.n4830 gnd.n4829 585
R3395 gnd.n4829 gnd.n4828 585
R3396 gnd.n1566 gnd.n1565 585
R3397 gnd.n4821 gnd.n1566 585
R3398 gnd.n4672 gnd.n4671 585
R3399 gnd.n4671 gnd.n1584 585
R3400 gnd.n4675 gnd.n4670 585
R3401 gnd.n4670 gnd.n1582 585
R3402 gnd.n4676 gnd.n4669 585
R3403 gnd.n4669 gnd.n1588 585
R3404 gnd.n4677 gnd.n4668 585
R3405 gnd.n4668 gnd.n1592 585
R3406 gnd.n4667 gnd.n4665 585
R3407 gnd.n4667 gnd.n1601 585
R3408 gnd.n4681 gnd.n4664 585
R3409 gnd.n4664 gnd.n1599 585
R3410 gnd.n4682 gnd.n4663 585
R3411 gnd.n4663 gnd.n4662 585
R3412 gnd.n4683 gnd.n1612 585
R3413 gnd.n4741 gnd.n1612 585
R3414 gnd.n4660 gnd.n1620 585
R3415 gnd.n4731 gnd.n1620 585
R3416 gnd.n4687 gnd.n4659 585
R3417 gnd.n4659 gnd.n1626 585
R3418 gnd.n4688 gnd.n4658 585
R3419 gnd.n4658 gnd.n1634 585
R3420 gnd.n4689 gnd.n4657 585
R3421 gnd.n4657 gnd.n1631 585
R3422 gnd.n1651 gnd.n1641 585
R3423 gnd.n4704 gnd.n1641 585
R3424 gnd.n4694 gnd.n4693 585
R3425 gnd.n4696 gnd.n4694 585
R3426 gnd.n1650 gnd.n1649 585
R3427 gnd.n4609 gnd.n1649 585
R3428 gnd.n4653 gnd.n4652 585
R3429 gnd.n4652 gnd.n4651 585
R3430 gnd.n1654 gnd.n1653 585
R3431 gnd.n4644 gnd.n1654 585
R3432 gnd.n4573 gnd.n4572 585
R3433 gnd.n4572 gnd.n1671 585
R3434 gnd.n4574 gnd.n4571 585
R3435 gnd.n4571 gnd.n1668 585
R3436 gnd.n1694 gnd.n1692 585
R3437 gnd.n1692 gnd.n1675 585
R3438 gnd.n4579 gnd.n4578 585
R3439 gnd.n4580 gnd.n4579 585
R3440 gnd.n1693 gnd.n1691 585
R3441 gnd.n1691 gnd.t174 585
R3442 gnd.n4567 gnd.n4566 585
R3443 gnd.n4566 gnd.n1684 585
R3444 gnd.n4565 gnd.n1696 585
R3445 gnd.n4565 gnd.n4564 585
R3446 gnd.n4488 gnd.n1697 585
R3447 gnd.n4556 gnd.n1697 585
R3448 gnd.n4487 gnd.n1711 585
R3449 gnd.n4546 gnd.n1711 585
R3450 gnd.n4492 gnd.n4486 585
R3451 gnd.n4486 gnd.n1716 585
R3452 gnd.n4493 gnd.n4485 585
R3453 gnd.n4485 gnd.n1724 585
R3454 gnd.n4494 gnd.n4484 585
R3455 gnd.n4484 gnd.n1721 585
R3456 gnd.n1741 gnd.n1731 585
R3457 gnd.n4509 gnd.n1731 585
R3458 gnd.n4499 gnd.n4498 585
R3459 gnd.n4500 gnd.n4499 585
R3460 gnd.n1740 gnd.n1739 585
R3461 gnd.n4435 gnd.n1739 585
R3462 gnd.n4480 gnd.n4479 585
R3463 gnd.n4479 gnd.n4478 585
R3464 gnd.n1744 gnd.n1743 585
R3465 gnd.n4471 gnd.n1744 585
R3466 gnd.n4267 gnd.n4265 585
R3467 gnd.n4265 gnd.n1760 585
R3468 gnd.n4268 gnd.n4264 585
R3469 gnd.n4264 gnd.n1758 585
R3470 gnd.n4269 gnd.n4263 585
R3471 gnd.n4263 gnd.n1764 585
R3472 gnd.n4262 gnd.n4258 585
R3473 gnd.n4262 gnd.n4261 585
R3474 gnd.n4273 gnd.n1774 585
R3475 gnd.n4413 gnd.n1774 585
R3476 gnd.n4274 gnd.n4257 585
R3477 gnd.n4257 gnd.n1773 585
R3478 gnd.n4275 gnd.n4256 585
R3479 gnd.n4256 gnd.n4255 585
R3480 gnd.n5321 gnd.n5320 585
R3481 gnd.n5320 gnd.n1117 585
R3482 gnd.n5319 gnd.n5149 585
R3483 gnd.n5317 gnd.n5316 585
R3484 gnd.n5151 gnd.n5150 585
R3485 gnd.n5312 gnd.n5308 585
R3486 gnd.n5306 gnd.n5153 585
R3487 gnd.n5304 gnd.n5303 585
R3488 gnd.n5155 gnd.n5154 585
R3489 gnd.n5299 gnd.n5298 585
R3490 gnd.n5296 gnd.n5157 585
R3491 gnd.n5294 gnd.n5293 585
R3492 gnd.n5159 gnd.n5158 585
R3493 gnd.n5279 gnd.n5278 585
R3494 gnd.n5280 gnd.n5276 585
R3495 gnd.n5274 gnd.n5168 585
R3496 gnd.n5273 gnd.n5272 585
R3497 gnd.n5257 gnd.n5170 585
R3498 gnd.n5259 gnd.n5258 585
R3499 gnd.n5255 gnd.n5177 585
R3500 gnd.n5254 gnd.n5253 585
R3501 gnd.n5238 gnd.n5179 585
R3502 gnd.n5240 gnd.n5239 585
R3503 gnd.n5236 gnd.n5186 585
R3504 gnd.n5235 gnd.n5234 585
R3505 gnd.n5219 gnd.n5188 585
R3506 gnd.n5221 gnd.n5220 585
R3507 gnd.n5217 gnd.n5195 585
R3508 gnd.n5216 gnd.n5215 585
R3509 gnd.n5197 gnd.n1105 585
R3510 gnd.n6259 gnd.n655 530.795
R3511 gnd.n5425 gnd.n1335 506.916
R3512 gnd.n5428 gnd.n5427 506.916
R3513 gnd.n4424 gnd.n1767 506.916
R3514 gnd.n4410 gnd.n1763 506.916
R3515 gnd.n1834 gnd.t112 389.64
R3516 gnd.n1329 gnd.t45 389.64
R3517 gnd.n1831 gnd.t63 389.64
R3518 gnd.n5359 gnd.t99 389.64
R3519 gnd.n2010 gnd.t92 371.625
R3520 gnd.n7021 gnd.t80 371.625
R3521 gnd.n5161 gnd.t70 371.625
R3522 gnd.n4186 gnd.t86 371.625
R3523 gnd.n5552 gnd.t67 371.625
R3524 gnd.n1268 gnd.t34 371.625
R3525 gnd.n156 gnd.t20 371.625
R3526 gnd.n7113 gnd.t49 371.625
R3527 gnd.n3719 gnd.t118 371.625
R3528 gnd.n3741 gnd.t109 371.625
R3529 gnd.n3640 gnd.t105 371.625
R3530 gnd.n1989 gnd.t41 371.625
R3531 gnd.n1900 gnd.t83 371.625
R3532 gnd.n5309 gnd.t76 371.625
R3533 gnd.n2630 gnd.t27 323.425
R3534 gnd.n2200 gnd.t59 323.425
R3535 gnd.n3479 gnd.n3453 289.615
R3536 gnd.n3447 gnd.n3421 289.615
R3537 gnd.n3415 gnd.n3389 289.615
R3538 gnd.n3384 gnd.n3358 289.615
R3539 gnd.n3352 gnd.n3326 289.615
R3540 gnd.n3320 gnd.n3294 289.615
R3541 gnd.n3288 gnd.n3262 289.615
R3542 gnd.n3257 gnd.n3231 289.615
R3543 gnd.n2704 gnd.t121 279.217
R3544 gnd.n2226 gnd.t55 279.217
R3545 gnd.n1816 gnd.t98 260.649
R3546 gnd.n5351 gnd.t104 260.649
R3547 gnd.n4412 gnd.n4411 256.663
R3548 gnd.n4412 gnd.n1775 256.663
R3549 gnd.n4412 gnd.n1776 256.663
R3550 gnd.n4412 gnd.n1777 256.663
R3551 gnd.n4412 gnd.n1778 256.663
R3552 gnd.n4412 gnd.n1779 256.663
R3553 gnd.n4412 gnd.n1780 256.663
R3554 gnd.n4412 gnd.n1781 256.663
R3555 gnd.n4412 gnd.n1782 256.663
R3556 gnd.n4412 gnd.n1783 256.663
R3557 gnd.n4412 gnd.n1784 256.663
R3558 gnd.n4412 gnd.n1785 256.663
R3559 gnd.n4412 gnd.n1786 256.663
R3560 gnd.n4412 gnd.n1787 256.663
R3561 gnd.n4412 gnd.n1788 256.663
R3562 gnd.n4412 gnd.n1789 256.663
R3563 gnd.n4348 gnd.n4345 256.663
R3564 gnd.n4412 gnd.n1790 256.663
R3565 gnd.n4412 gnd.n1791 256.663
R3566 gnd.n4412 gnd.n1792 256.663
R3567 gnd.n4412 gnd.n1793 256.663
R3568 gnd.n4412 gnd.n1794 256.663
R3569 gnd.n4412 gnd.n1795 256.663
R3570 gnd.n4412 gnd.n1796 256.663
R3571 gnd.n4412 gnd.n1797 256.663
R3572 gnd.n4412 gnd.n1798 256.663
R3573 gnd.n4412 gnd.n1799 256.663
R3574 gnd.n4412 gnd.n1800 256.663
R3575 gnd.n4412 gnd.n1801 256.663
R3576 gnd.n4412 gnd.n1802 256.663
R3577 gnd.n4412 gnd.n1803 256.663
R3578 gnd.n4412 gnd.n1804 256.663
R3579 gnd.n4412 gnd.n1805 256.663
R3580 gnd.n4412 gnd.n1806 256.663
R3581 gnd.n5493 gnd.n1313 256.663
R3582 gnd.n5493 gnd.n1314 256.663
R3583 gnd.n5493 gnd.n1315 256.663
R3584 gnd.n5493 gnd.n1316 256.663
R3585 gnd.n5493 gnd.n1317 256.663
R3586 gnd.n5493 gnd.n1318 256.663
R3587 gnd.n5493 gnd.n1319 256.663
R3588 gnd.n5493 gnd.n1320 256.663
R3589 gnd.n5493 gnd.n1321 256.663
R3590 gnd.n5493 gnd.n1322 256.663
R3591 gnd.n5493 gnd.n1323 256.663
R3592 gnd.n5493 gnd.n1324 256.663
R3593 gnd.n5493 gnd.n1325 256.663
R3594 gnd.n5493 gnd.n1326 256.663
R3595 gnd.n5493 gnd.n1327 256.663
R3596 gnd.n5493 gnd.n5490 256.663
R3597 gnd.n5496 gnd.n1294 256.663
R3598 gnd.n5494 gnd.n5493 256.663
R3599 gnd.n5493 gnd.n1312 256.663
R3600 gnd.n5493 gnd.n1311 256.663
R3601 gnd.n5493 gnd.n1310 256.663
R3602 gnd.n5493 gnd.n1309 256.663
R3603 gnd.n5493 gnd.n1308 256.663
R3604 gnd.n5493 gnd.n1307 256.663
R3605 gnd.n5493 gnd.n1306 256.663
R3606 gnd.n5493 gnd.n1305 256.663
R3607 gnd.n5493 gnd.n1304 256.663
R3608 gnd.n5493 gnd.n1303 256.663
R3609 gnd.n5493 gnd.n1302 256.663
R3610 gnd.n5493 gnd.n1301 256.663
R3611 gnd.n5493 gnd.n1300 256.663
R3612 gnd.n5493 gnd.n1299 256.663
R3613 gnd.n5493 gnd.n1298 256.663
R3614 gnd.n5493 gnd.n1297 256.663
R3615 gnd.n3842 gnd.n3841 242.672
R3616 gnd.n3841 gnd.n3630 242.672
R3617 gnd.n3841 gnd.n3631 242.672
R3618 gnd.n3841 gnd.n3632 242.672
R3619 gnd.n3841 gnd.n3633 242.672
R3620 gnd.n3841 gnd.n3634 242.672
R3621 gnd.n3841 gnd.n3635 242.672
R3622 gnd.n3841 gnd.n3636 242.672
R3623 gnd.n3841 gnd.n3637 242.672
R3624 gnd.n4195 gnd.n1961 242.672
R3625 gnd.n4184 gnd.n1961 242.672
R3626 gnd.n4181 gnd.n1961 242.672
R3627 gnd.n4172 gnd.n1961 242.672
R3628 gnd.n4161 gnd.n1961 242.672
R3629 gnd.n4158 gnd.n1961 242.672
R3630 gnd.n4149 gnd.n1961 242.672
R3631 gnd.n4139 gnd.n1961 242.672
R3632 gnd.n4136 gnd.n1961 242.672
R3633 gnd.n5207 gnd.n1118 242.672
R3634 gnd.n5209 gnd.n1118 242.672
R3635 gnd.n5226 gnd.n1118 242.672
R3636 gnd.n5228 gnd.n1118 242.672
R3637 gnd.n5245 gnd.n1118 242.672
R3638 gnd.n5247 gnd.n1118 242.672
R3639 gnd.n5264 gnd.n1118 242.672
R3640 gnd.n5266 gnd.n1118 242.672
R3641 gnd.n5285 gnd.n1118 242.672
R3642 gnd.n7023 gnd.n83 242.672
R3643 gnd.n7019 gnd.n83 242.672
R3644 gnd.n7014 gnd.n83 242.672
R3645 gnd.n7011 gnd.n83 242.672
R3646 gnd.n7006 gnd.n83 242.672
R3647 gnd.n7003 gnd.n83 242.672
R3648 gnd.n6998 gnd.n83 242.672
R3649 gnd.n6995 gnd.n83 242.672
R3650 gnd.n6990 gnd.n83 242.672
R3651 gnd.n2758 gnd.n2757 242.672
R3652 gnd.n2758 gnd.n2668 242.672
R3653 gnd.n2758 gnd.n2669 242.672
R3654 gnd.n2758 gnd.n2670 242.672
R3655 gnd.n2758 gnd.n2671 242.672
R3656 gnd.n2758 gnd.n2672 242.672
R3657 gnd.n2758 gnd.n2673 242.672
R3658 gnd.n2758 gnd.n2674 242.672
R3659 gnd.n2758 gnd.n2675 242.672
R3660 gnd.n2758 gnd.n2676 242.672
R3661 gnd.n2758 gnd.n2677 242.672
R3662 gnd.n2758 gnd.n2678 242.672
R3663 gnd.n2759 gnd.n2758 242.672
R3664 gnd.n3611 gnd.n2175 242.672
R3665 gnd.n3611 gnd.n2174 242.672
R3666 gnd.n3611 gnd.n2173 242.672
R3667 gnd.n3611 gnd.n2172 242.672
R3668 gnd.n3611 gnd.n2171 242.672
R3669 gnd.n3611 gnd.n2170 242.672
R3670 gnd.n3611 gnd.n2169 242.672
R3671 gnd.n3611 gnd.n2168 242.672
R3672 gnd.n3611 gnd.n2167 242.672
R3673 gnd.n3611 gnd.n2166 242.672
R3674 gnd.n3611 gnd.n2165 242.672
R3675 gnd.n3611 gnd.n2164 242.672
R3676 gnd.n3611 gnd.n2163 242.672
R3677 gnd.n2842 gnd.n2841 242.672
R3678 gnd.n2841 gnd.n2580 242.672
R3679 gnd.n2841 gnd.n2581 242.672
R3680 gnd.n2841 gnd.n2582 242.672
R3681 gnd.n2841 gnd.n2583 242.672
R3682 gnd.n2841 gnd.n2584 242.672
R3683 gnd.n2841 gnd.n2585 242.672
R3684 gnd.n2841 gnd.n2586 242.672
R3685 gnd.n3611 gnd.n2176 242.672
R3686 gnd.n3611 gnd.n2177 242.672
R3687 gnd.n3611 gnd.n2178 242.672
R3688 gnd.n3611 gnd.n2179 242.672
R3689 gnd.n3611 gnd.n2180 242.672
R3690 gnd.n3611 gnd.n2181 242.672
R3691 gnd.n3611 gnd.n2182 242.672
R3692 gnd.n3611 gnd.n2183 242.672
R3693 gnd.n3841 gnd.n3840 242.672
R3694 gnd.n3841 gnd.n3612 242.672
R3695 gnd.n3841 gnd.n3613 242.672
R3696 gnd.n3841 gnd.n3614 242.672
R3697 gnd.n3841 gnd.n3615 242.672
R3698 gnd.n3841 gnd.n3616 242.672
R3699 gnd.n3841 gnd.n3617 242.672
R3700 gnd.n3841 gnd.n3618 242.672
R3701 gnd.n3841 gnd.n3619 242.672
R3702 gnd.n3841 gnd.n3620 242.672
R3703 gnd.n3841 gnd.n3621 242.672
R3704 gnd.n3841 gnd.n3622 242.672
R3705 gnd.n3841 gnd.n3623 242.672
R3706 gnd.n3841 gnd.n3624 242.672
R3707 gnd.n3841 gnd.n3625 242.672
R3708 gnd.n3841 gnd.n3626 242.672
R3709 gnd.n3841 gnd.n3627 242.672
R3710 gnd.n3841 gnd.n3628 242.672
R3711 gnd.n3841 gnd.n3629 242.672
R3712 gnd.n4307 gnd.n1961 242.672
R3713 gnd.n1992 gnd.n1961 242.672
R3714 gnd.n4314 gnd.n1961 242.672
R3715 gnd.n1983 gnd.n1961 242.672
R3716 gnd.n4321 gnd.n1961 242.672
R3717 gnd.n1976 gnd.n1961 242.672
R3718 gnd.n4328 gnd.n1961 242.672
R3719 gnd.n1969 gnd.n1961 242.672
R3720 gnd.n4335 gnd.n1961 242.672
R3721 gnd.n4338 gnd.n1961 242.672
R3722 gnd.n1961 gnd.n1907 242.672
R3723 gnd.n4344 gnd.n1902 242.672
R3724 gnd.n1961 gnd.n1908 242.672
R3725 gnd.n1961 gnd.n1909 242.672
R3726 gnd.n1961 gnd.n1910 242.672
R3727 gnd.n1961 gnd.n1911 242.672
R3728 gnd.n1961 gnd.n1912 242.672
R3729 gnd.n1961 gnd.n1913 242.672
R3730 gnd.n1961 gnd.n1914 242.672
R3731 gnd.n1961 gnd.n1960 242.672
R3732 gnd.n5515 gnd.n1118 242.672
R3733 gnd.n5518 gnd.n1118 242.672
R3734 gnd.n5526 gnd.n1118 242.672
R3735 gnd.n5528 gnd.n1118 242.672
R3736 gnd.n5536 gnd.n1118 242.672
R3737 gnd.n5538 gnd.n1118 242.672
R3738 gnd.n5547 gnd.n1118 242.672
R3739 gnd.n5550 gnd.n1118 242.672
R3740 gnd.n5554 gnd.n5551 242.672
R3741 gnd.n5497 gnd.n1118 242.672
R3742 gnd.n5560 gnd.n1118 242.672
R3743 gnd.n5562 gnd.n1118 242.672
R3744 gnd.n5570 gnd.n1118 242.672
R3745 gnd.n5572 gnd.n1118 242.672
R3746 gnd.n5580 gnd.n1118 242.672
R3747 gnd.n5582 gnd.n1118 242.672
R3748 gnd.n5590 gnd.n1118 242.672
R3749 gnd.n5592 gnd.n1118 242.672
R3750 gnd.n5601 gnd.n1118 242.672
R3751 gnd.n5604 gnd.n1118 242.672
R3752 gnd.n153 gnd.n83 242.672
R3753 gnd.n7081 gnd.n83 242.672
R3754 gnd.n149 gnd.n83 242.672
R3755 gnd.n7088 gnd.n83 242.672
R3756 gnd.n142 gnd.n83 242.672
R3757 gnd.n7095 gnd.n83 242.672
R3758 gnd.n135 gnd.n83 242.672
R3759 gnd.n7102 gnd.n83 242.672
R3760 gnd.n128 gnd.n83 242.672
R3761 gnd.n7109 gnd.n83 242.672
R3762 gnd.n121 gnd.n83 242.672
R3763 gnd.n7119 gnd.n83 242.672
R3764 gnd.n114 gnd.n83 242.672
R3765 gnd.n7126 gnd.n83 242.672
R3766 gnd.n107 gnd.n83 242.672
R3767 gnd.n7133 gnd.n83 242.672
R3768 gnd.n100 gnd.n83 242.672
R3769 gnd.n7140 gnd.n83 242.672
R3770 gnd.n93 gnd.n83 242.672
R3771 gnd.n4244 gnd.n4243 242.672
R3772 gnd.n4244 gnd.n4113 242.672
R3773 gnd.n4244 gnd.n4114 242.672
R3774 gnd.n4244 gnd.n4115 242.672
R3775 gnd.n4244 gnd.n4116 242.672
R3776 gnd.n4244 gnd.n4117 242.672
R3777 gnd.n4244 gnd.n4118 242.672
R3778 gnd.n4244 gnd.n4119 242.672
R3779 gnd.n4244 gnd.n4120 242.672
R3780 gnd.n4244 gnd.n4121 242.672
R3781 gnd.n4244 gnd.n4123 242.672
R3782 gnd.n4244 gnd.n4124 242.672
R3783 gnd.n4244 gnd.n4125 242.672
R3784 gnd.n4244 gnd.n4126 242.672
R3785 gnd.n5318 gnd.n1117 242.672
R3786 gnd.n5307 gnd.n1117 242.672
R3787 gnd.n5305 gnd.n1117 242.672
R3788 gnd.n5297 gnd.n1117 242.672
R3789 gnd.n5295 gnd.n1117 242.672
R3790 gnd.n5277 gnd.n1117 242.672
R3791 gnd.n5275 gnd.n1117 242.672
R3792 gnd.n5169 gnd.n1117 242.672
R3793 gnd.n5256 gnd.n1117 242.672
R3794 gnd.n5178 gnd.n1117 242.672
R3795 gnd.n5237 gnd.n1117 242.672
R3796 gnd.n5187 gnd.n1117 242.672
R3797 gnd.n5218 gnd.n1117 242.672
R3798 gnd.n5196 gnd.n1117 242.672
R3799 gnd.n90 gnd.n86 240.244
R3800 gnd.n7142 gnd.n7141 240.244
R3801 gnd.n7139 gnd.n94 240.244
R3802 gnd.n7135 gnd.n7134 240.244
R3803 gnd.n7132 gnd.n101 240.244
R3804 gnd.n7128 gnd.n7127 240.244
R3805 gnd.n7125 gnd.n108 240.244
R3806 gnd.n7121 gnd.n7120 240.244
R3807 gnd.n7118 gnd.n115 240.244
R3808 gnd.n7111 gnd.n7110 240.244
R3809 gnd.n7108 gnd.n122 240.244
R3810 gnd.n7104 gnd.n7103 240.244
R3811 gnd.n7101 gnd.n129 240.244
R3812 gnd.n7097 gnd.n7096 240.244
R3813 gnd.n7094 gnd.n136 240.244
R3814 gnd.n7090 gnd.n7089 240.244
R3815 gnd.n7087 gnd.n143 240.244
R3816 gnd.n7083 gnd.n7082 240.244
R3817 gnd.n7080 gnd.n150 240.244
R3818 gnd.n5611 gnd.n1127 240.244
R3819 gnd.n5611 gnd.n1139 240.244
R3820 gnd.n5622 gnd.n1139 240.244
R3821 gnd.n5622 gnd.n1257 240.244
R3822 gnd.n5669 gnd.n1257 240.244
R3823 gnd.n5669 gnd.n1250 240.244
R3824 gnd.n5665 gnd.n1250 240.244
R3825 gnd.n5665 gnd.n1242 240.244
R3826 gnd.n1242 gnd.n1231 240.244
R3827 gnd.n5661 gnd.n1231 240.244
R3828 gnd.n5661 gnd.n1221 240.244
R3829 gnd.n5658 gnd.n1221 240.244
R3830 gnd.n5658 gnd.n1213 240.244
R3831 gnd.n1213 gnd.n1202 240.244
R3832 gnd.n5654 gnd.n1202 240.244
R3833 gnd.n5654 gnd.n1195 240.244
R3834 gnd.n5651 gnd.n1195 240.244
R3835 gnd.n5651 gnd.n1185 240.244
R3836 gnd.n5647 gnd.n1185 240.244
R3837 gnd.n5647 gnd.n1177 240.244
R3838 gnd.n5644 gnd.n1177 240.244
R3839 gnd.n5644 gnd.n236 240.244
R3840 gnd.n6926 gnd.n236 240.244
R3841 gnd.n6926 gnd.n232 240.244
R3842 gnd.n6922 gnd.n232 240.244
R3843 gnd.n6922 gnd.n224 240.244
R3844 gnd.n6917 gnd.n224 240.244
R3845 gnd.n6917 gnd.n210 240.244
R3846 gnd.n6913 gnd.n210 240.244
R3847 gnd.n6913 gnd.n203 240.244
R3848 gnd.n6908 gnd.n203 240.244
R3849 gnd.n6908 gnd.n195 240.244
R3850 gnd.n267 gnd.n195 240.244
R3851 gnd.n267 gnd.n187 240.244
R3852 gnd.n262 gnd.n187 240.244
R3853 gnd.n262 gnd.n178 240.244
R3854 gnd.n258 gnd.n178 240.244
R3855 gnd.n258 gnd.n169 240.244
R3856 gnd.n169 gnd.n160 240.244
R3857 gnd.n7071 gnd.n160 240.244
R3858 gnd.n7072 gnd.n7071 240.244
R3859 gnd.n7072 gnd.n82 240.244
R3860 gnd.n5517 gnd.n5516 240.244
R3861 gnd.n5519 gnd.n5517 240.244
R3862 gnd.n5525 gnd.n5507 240.244
R3863 gnd.n5529 gnd.n5527 240.244
R3864 gnd.n5535 gnd.n5503 240.244
R3865 gnd.n5539 gnd.n5537 240.244
R3866 gnd.n5546 gnd.n5499 240.244
R3867 gnd.n5549 gnd.n5548 240.244
R3868 gnd.n5559 gnd.n1288 240.244
R3869 gnd.n5563 gnd.n5561 240.244
R3870 gnd.n5569 gnd.n1284 240.244
R3871 gnd.n5573 gnd.n5571 240.244
R3872 gnd.n5579 gnd.n1280 240.244
R3873 gnd.n5583 gnd.n5581 240.244
R3874 gnd.n5589 gnd.n1276 240.244
R3875 gnd.n5593 gnd.n5591 240.244
R3876 gnd.n5600 gnd.n1272 240.244
R3877 gnd.n5603 gnd.n5602 240.244
R3878 gnd.n5850 gnd.n1132 240.244
R3879 gnd.n5846 gnd.n1132 240.244
R3880 gnd.n5846 gnd.n1137 240.244
R3881 gnd.n5689 gnd.n1137 240.244
R3882 gnd.n5689 gnd.n1252 240.244
R3883 gnd.n5697 gnd.n1252 240.244
R3884 gnd.n5697 gnd.n1253 240.244
R3885 gnd.n1253 gnd.n1229 240.244
R3886 gnd.n5720 gnd.n1229 240.244
R3887 gnd.n5720 gnd.n1224 240.244
R3888 gnd.n5729 gnd.n1224 240.244
R3889 gnd.n5729 gnd.n1225 240.244
R3890 gnd.n1225 gnd.n1200 240.244
R3891 gnd.n5758 gnd.n1200 240.244
R3892 gnd.n5758 gnd.n1197 240.244
R3893 gnd.n5762 gnd.n1197 240.244
R3894 gnd.n5762 gnd.n1181 240.244
R3895 gnd.n5774 gnd.n1181 240.244
R3896 gnd.n5775 gnd.n5774 240.244
R3897 gnd.n5781 gnd.n5775 240.244
R3898 gnd.n5781 gnd.n5778 240.244
R3899 gnd.n5778 gnd.n234 240.244
R3900 gnd.n6928 gnd.n234 240.244
R3901 gnd.n6931 gnd.n6928 240.244
R3902 gnd.n6931 gnd.n222 240.244
R3903 gnd.n6941 gnd.n222 240.244
R3904 gnd.n6941 gnd.n212 240.244
R3905 gnd.n6947 gnd.n212 240.244
R3906 gnd.n6947 gnd.n201 240.244
R3907 gnd.n6957 gnd.n201 240.244
R3908 gnd.n6957 gnd.n197 240.244
R3909 gnd.n6963 gnd.n197 240.244
R3910 gnd.n6963 gnd.n185 240.244
R3911 gnd.n6973 gnd.n185 240.244
R3912 gnd.n6973 gnd.n181 240.244
R3913 gnd.n6979 gnd.n181 240.244
R3914 gnd.n6979 gnd.n167 240.244
R3915 gnd.n7063 gnd.n167 240.244
R3916 gnd.n7063 gnd.n163 240.244
R3917 gnd.n7069 gnd.n163 240.244
R3918 gnd.n7069 gnd.n85 240.244
R3919 gnd.n7149 gnd.n85 240.244
R3920 gnd.n1915 gnd.n992 240.244
R3921 gnd.n1959 gnd.n1916 240.244
R3922 gnd.n1955 gnd.n1954 240.244
R3923 gnd.n1951 gnd.n1950 240.244
R3924 gnd.n1947 gnd.n1946 240.244
R3925 gnd.n1943 gnd.n1942 240.244
R3926 gnd.n1939 gnd.n1938 240.244
R3927 gnd.n1935 gnd.n1934 240.244
R3928 gnd.n4339 gnd.n1906 240.244
R3929 gnd.n4337 gnd.n4336 240.244
R3930 gnd.n4334 gnd.n1963 240.244
R3931 gnd.n4330 gnd.n4329 240.244
R3932 gnd.n4327 gnd.n1970 240.244
R3933 gnd.n4323 gnd.n4322 240.244
R3934 gnd.n4320 gnd.n1977 240.244
R3935 gnd.n4316 gnd.n4315 240.244
R3936 gnd.n4313 gnd.n1984 240.244
R3937 gnd.n4309 gnd.n4308 240.244
R3938 gnd.n3762 gnd.n2152 240.244
R3939 gnd.n3745 gnd.n2152 240.244
R3940 gnd.n3745 gnd.n2144 240.244
R3941 gnd.n3754 gnd.n2144 240.244
R3942 gnd.n3754 gnd.n828 240.244
R3943 gnd.n3751 gnd.n828 240.244
R3944 gnd.n3751 gnd.n841 240.244
R3945 gnd.n3882 gnd.n841 240.244
R3946 gnd.n3882 gnd.n853 240.244
R3947 gnd.n2129 gnd.n853 240.244
R3948 gnd.n2129 gnd.n863 240.244
R3949 gnd.n3894 gnd.n863 240.244
R3950 gnd.n3894 gnd.n874 240.244
R3951 gnd.n2123 gnd.n874 240.244
R3952 gnd.n2123 gnd.n884 240.244
R3953 gnd.n3940 gnd.n884 240.244
R3954 gnd.n3940 gnd.n895 240.244
R3955 gnd.n3948 gnd.n895 240.244
R3956 gnd.n3948 gnd.n2112 240.244
R3957 gnd.n2112 gnd.n2104 240.244
R3958 gnd.n3985 gnd.n2104 240.244
R3959 gnd.n3985 gnd.n2085 240.244
R3960 gnd.n2085 gnd.n2078 240.244
R3961 gnd.n2100 gnd.n2078 240.244
R3962 gnd.n2100 gnd.n2071 240.244
R3963 gnd.n2071 gnd.n910 240.244
R3964 gnd.n2064 gnd.n910 240.244
R3965 gnd.n2064 gnd.n921 240.244
R3966 gnd.n4034 gnd.n921 240.244
R3967 gnd.n4034 gnd.n931 240.244
R3968 gnd.n2044 gnd.n931 240.244
R3969 gnd.n2044 gnd.n941 240.244
R3970 gnd.n4042 gnd.n941 240.244
R3971 gnd.n4042 gnd.n952 240.244
R3972 gnd.n4049 gnd.n952 240.244
R3973 gnd.n4049 gnd.n962 240.244
R3974 gnd.n4053 gnd.n962 240.244
R3975 gnd.n4053 gnd.n973 240.244
R3976 gnd.n4060 gnd.n973 240.244
R3977 gnd.n4060 gnd.n984 240.244
R3978 gnd.n4300 gnd.n984 240.244
R3979 gnd.n4300 gnd.n994 240.244
R3980 gnd.n3700 gnd.n3699 240.244
R3981 gnd.n3834 gnd.n3699 240.244
R3982 gnd.n3832 gnd.n3831 240.244
R3983 gnd.n3828 gnd.n3827 240.244
R3984 gnd.n3824 gnd.n3823 240.244
R3985 gnd.n3820 gnd.n3819 240.244
R3986 gnd.n3816 gnd.n3815 240.244
R3987 gnd.n3812 gnd.n3811 240.244
R3988 gnd.n3808 gnd.n3807 240.244
R3989 gnd.n3803 gnd.n3802 240.244
R3990 gnd.n3799 gnd.n3798 240.244
R3991 gnd.n3795 gnd.n3794 240.244
R3992 gnd.n3791 gnd.n3790 240.244
R3993 gnd.n3787 gnd.n3786 240.244
R3994 gnd.n3783 gnd.n3782 240.244
R3995 gnd.n3779 gnd.n3778 240.244
R3996 gnd.n3775 gnd.n3774 240.244
R3997 gnd.n3771 gnd.n3770 240.244
R3998 gnd.n3740 gnd.n3739 240.244
R3999 gnd.n3860 gnd.n2150 240.244
R4000 gnd.n3860 gnd.n2146 240.244
R4001 gnd.n3867 gnd.n2146 240.244
R4002 gnd.n3867 gnd.n832 240.244
R4003 gnd.n6089 gnd.n832 240.244
R4004 gnd.n6089 gnd.n833 240.244
R4005 gnd.n6085 gnd.n833 240.244
R4006 gnd.n6085 gnd.n839 240.244
R4007 gnd.n6077 gnd.n839 240.244
R4008 gnd.n6077 gnd.n855 240.244
R4009 gnd.n6073 gnd.n855 240.244
R4010 gnd.n6073 gnd.n861 240.244
R4011 gnd.n6065 gnd.n861 240.244
R4012 gnd.n6065 gnd.n877 240.244
R4013 gnd.n6061 gnd.n877 240.244
R4014 gnd.n6061 gnd.n883 240.244
R4015 gnd.n6053 gnd.n883 240.244
R4016 gnd.n6053 gnd.n897 240.244
R4017 gnd.n3975 gnd.n897 240.244
R4018 gnd.n3975 gnd.n3974 240.244
R4019 gnd.n3974 gnd.n2081 240.244
R4020 gnd.n3999 gnd.n2081 240.244
R4021 gnd.n4003 gnd.n3999 240.244
R4022 gnd.n4003 gnd.n4000 240.244
R4023 gnd.n4000 gnd.n907 240.244
R4024 gnd.n6047 gnd.n907 240.244
R4025 gnd.n6047 gnd.n908 240.244
R4026 gnd.n6039 gnd.n908 240.244
R4027 gnd.n6039 gnd.n924 240.244
R4028 gnd.n6035 gnd.n924 240.244
R4029 gnd.n6035 gnd.n929 240.244
R4030 gnd.n6027 gnd.n929 240.244
R4031 gnd.n6027 gnd.n944 240.244
R4032 gnd.n6023 gnd.n944 240.244
R4033 gnd.n6023 gnd.n950 240.244
R4034 gnd.n6015 gnd.n950 240.244
R4035 gnd.n6015 gnd.n965 240.244
R4036 gnd.n6011 gnd.n965 240.244
R4037 gnd.n6011 gnd.n971 240.244
R4038 gnd.n6003 gnd.n971 240.244
R4039 gnd.n6003 gnd.n987 240.244
R4040 gnd.n5999 gnd.n987 240.244
R4041 gnd.n3610 gnd.n2185 240.244
R4042 gnd.n3603 gnd.n3602 240.244
R4043 gnd.n3600 gnd.n3599 240.244
R4044 gnd.n3596 gnd.n3595 240.244
R4045 gnd.n3592 gnd.n3591 240.244
R4046 gnd.n3588 gnd.n3587 240.244
R4047 gnd.n3584 gnd.n3583 240.244
R4048 gnd.n3580 gnd.n3579 240.244
R4049 gnd.n2853 gnd.n2565 240.244
R4050 gnd.n2863 gnd.n2565 240.244
R4051 gnd.n2863 gnd.n2556 240.244
R4052 gnd.n2556 gnd.n2545 240.244
R4053 gnd.n2884 gnd.n2545 240.244
R4054 gnd.n2884 gnd.n2539 240.244
R4055 gnd.n2894 gnd.n2539 240.244
R4056 gnd.n2894 gnd.n2528 240.244
R4057 gnd.n2528 gnd.n2520 240.244
R4058 gnd.n2912 gnd.n2520 240.244
R4059 gnd.n2913 gnd.n2912 240.244
R4060 gnd.n2913 gnd.n2505 240.244
R4061 gnd.n2915 gnd.n2505 240.244
R4062 gnd.n2915 gnd.n2491 240.244
R4063 gnd.n2957 gnd.n2491 240.244
R4064 gnd.n2958 gnd.n2957 240.244
R4065 gnd.n2961 gnd.n2958 240.244
R4066 gnd.n2961 gnd.n2446 240.244
R4067 gnd.n2486 gnd.n2446 240.244
R4068 gnd.n2486 gnd.n2456 240.244
R4069 gnd.n2971 gnd.n2456 240.244
R4070 gnd.n2971 gnd.n2477 240.244
R4071 gnd.n2981 gnd.n2477 240.244
R4072 gnd.n2981 gnd.n2387 240.244
R4073 gnd.n3026 gnd.n2387 240.244
R4074 gnd.n3026 gnd.n2373 240.244
R4075 gnd.n3048 gnd.n2373 240.244
R4076 gnd.n3049 gnd.n3048 240.244
R4077 gnd.n3049 gnd.n2360 240.244
R4078 gnd.n2360 gnd.n2349 240.244
R4079 gnd.n3080 gnd.n2349 240.244
R4080 gnd.n3081 gnd.n3080 240.244
R4081 gnd.n3082 gnd.n3081 240.244
R4082 gnd.n3082 gnd.n2334 240.244
R4083 gnd.n2334 gnd.n2333 240.244
R4084 gnd.n2333 gnd.n2318 240.244
R4085 gnd.n3133 gnd.n2318 240.244
R4086 gnd.n3134 gnd.n3133 240.244
R4087 gnd.n3134 gnd.n2305 240.244
R4088 gnd.n2305 gnd.n2294 240.244
R4089 gnd.n3166 gnd.n2294 240.244
R4090 gnd.n3167 gnd.n3166 240.244
R4091 gnd.n3168 gnd.n3167 240.244
R4092 gnd.n3168 gnd.n2278 240.244
R4093 gnd.n2278 gnd.n2277 240.244
R4094 gnd.n2277 gnd.n2264 240.244
R4095 gnd.n3223 gnd.n2264 240.244
R4096 gnd.n3224 gnd.n3223 240.244
R4097 gnd.n3224 gnd.n2251 240.244
R4098 gnd.n2251 gnd.n2241 240.244
R4099 gnd.n3511 gnd.n2241 240.244
R4100 gnd.n3514 gnd.n3511 240.244
R4101 gnd.n3514 gnd.n3513 240.244
R4102 gnd.n2843 gnd.n2578 240.244
R4103 gnd.n2599 gnd.n2578 240.244
R4104 gnd.n2602 gnd.n2601 240.244
R4105 gnd.n2609 gnd.n2608 240.244
R4106 gnd.n2612 gnd.n2611 240.244
R4107 gnd.n2619 gnd.n2618 240.244
R4108 gnd.n2622 gnd.n2621 240.244
R4109 gnd.n2629 gnd.n2628 240.244
R4110 gnd.n2851 gnd.n2575 240.244
R4111 gnd.n2575 gnd.n2554 240.244
R4112 gnd.n2874 gnd.n2554 240.244
R4113 gnd.n2874 gnd.n2548 240.244
R4114 gnd.n2882 gnd.n2548 240.244
R4115 gnd.n2882 gnd.n2550 240.244
R4116 gnd.n2550 gnd.n2526 240.244
R4117 gnd.n2904 gnd.n2526 240.244
R4118 gnd.n2904 gnd.n2522 240.244
R4119 gnd.n2910 gnd.n2522 240.244
R4120 gnd.n2910 gnd.n2504 240.244
R4121 gnd.n2935 gnd.n2504 240.244
R4122 gnd.n2935 gnd.n2499 240.244
R4123 gnd.n2947 gnd.n2499 240.244
R4124 gnd.n2947 gnd.n2500 240.244
R4125 gnd.n2943 gnd.n2500 240.244
R4126 gnd.n2943 gnd.n2448 240.244
R4127 gnd.n2995 gnd.n2448 240.244
R4128 gnd.n2995 gnd.n2449 240.244
R4129 gnd.n2991 gnd.n2449 240.244
R4130 gnd.n2991 gnd.n2455 240.244
R4131 gnd.n2475 gnd.n2455 240.244
R4132 gnd.n2475 gnd.n2385 240.244
R4133 gnd.n3030 gnd.n2385 240.244
R4134 gnd.n3030 gnd.n2380 240.244
R4135 gnd.n3038 gnd.n2380 240.244
R4136 gnd.n3038 gnd.n2381 240.244
R4137 gnd.n2381 gnd.n2358 240.244
R4138 gnd.n3070 gnd.n2358 240.244
R4139 gnd.n3070 gnd.n2353 240.244
R4140 gnd.n3078 gnd.n2353 240.244
R4141 gnd.n3078 gnd.n2354 240.244
R4142 gnd.n2354 gnd.n2331 240.244
R4143 gnd.n3115 gnd.n2331 240.244
R4144 gnd.n3115 gnd.n2326 240.244
R4145 gnd.n3123 gnd.n2326 240.244
R4146 gnd.n3123 gnd.n2327 240.244
R4147 gnd.n2327 gnd.n2303 240.244
R4148 gnd.n3156 gnd.n2303 240.244
R4149 gnd.n3156 gnd.n2298 240.244
R4150 gnd.n3164 gnd.n2298 240.244
R4151 gnd.n3164 gnd.n2299 240.244
R4152 gnd.n2299 gnd.n2276 240.244
R4153 gnd.n3205 gnd.n2276 240.244
R4154 gnd.n3205 gnd.n2271 240.244
R4155 gnd.n3213 gnd.n2271 240.244
R4156 gnd.n3213 gnd.n2272 240.244
R4157 gnd.n2272 gnd.n2249 240.244
R4158 gnd.n3499 gnd.n2249 240.244
R4159 gnd.n3499 gnd.n2244 240.244
R4160 gnd.n3509 gnd.n2244 240.244
R4161 gnd.n3509 gnd.n2245 240.244
R4162 gnd.n2245 gnd.n2184 240.244
R4163 gnd.n2204 gnd.n2162 240.244
R4164 gnd.n3570 gnd.n3569 240.244
R4165 gnd.n3566 gnd.n3565 240.244
R4166 gnd.n3562 gnd.n3561 240.244
R4167 gnd.n3558 gnd.n3557 240.244
R4168 gnd.n3554 gnd.n3553 240.244
R4169 gnd.n3550 gnd.n3549 240.244
R4170 gnd.n3546 gnd.n3545 240.244
R4171 gnd.n3542 gnd.n3541 240.244
R4172 gnd.n3538 gnd.n3537 240.244
R4173 gnd.n3534 gnd.n3533 240.244
R4174 gnd.n3530 gnd.n3529 240.244
R4175 gnd.n3526 gnd.n3525 240.244
R4176 gnd.n2766 gnd.n2663 240.244
R4177 gnd.n2766 gnd.n2656 240.244
R4178 gnd.n2777 gnd.n2656 240.244
R4179 gnd.n2777 gnd.n2652 240.244
R4180 gnd.n2783 gnd.n2652 240.244
R4181 gnd.n2783 gnd.n2644 240.244
R4182 gnd.n2793 gnd.n2644 240.244
R4183 gnd.n2793 gnd.n2639 240.244
R4184 gnd.n2829 gnd.n2639 240.244
R4185 gnd.n2829 gnd.n2640 240.244
R4186 gnd.n2640 gnd.n2587 240.244
R4187 gnd.n2824 gnd.n2587 240.244
R4188 gnd.n2824 gnd.n2823 240.244
R4189 gnd.n2823 gnd.n2566 240.244
R4190 gnd.n2819 gnd.n2566 240.244
R4191 gnd.n2819 gnd.n2557 240.244
R4192 gnd.n2816 gnd.n2557 240.244
R4193 gnd.n2816 gnd.n2815 240.244
R4194 gnd.n2815 gnd.n2540 240.244
R4195 gnd.n2811 gnd.n2540 240.244
R4196 gnd.n2811 gnd.n2529 240.244
R4197 gnd.n2529 gnd.n2510 240.244
R4198 gnd.n2924 gnd.n2510 240.244
R4199 gnd.n2924 gnd.n2506 240.244
R4200 gnd.n2932 gnd.n2506 240.244
R4201 gnd.n2932 gnd.n2497 240.244
R4202 gnd.n2497 gnd.n2433 240.244
R4203 gnd.n3004 gnd.n2433 240.244
R4204 gnd.n3004 gnd.n2434 240.244
R4205 gnd.n2445 gnd.n2434 240.244
R4206 gnd.n2480 gnd.n2445 240.244
R4207 gnd.n2483 gnd.n2480 240.244
R4208 gnd.n2483 gnd.n2457 240.244
R4209 gnd.n2470 gnd.n2457 240.244
R4210 gnd.n2470 gnd.n2467 240.244
R4211 gnd.n2467 gnd.n2388 240.244
R4212 gnd.n3025 gnd.n2388 240.244
R4213 gnd.n3025 gnd.n2378 240.244
R4214 gnd.n3021 gnd.n2378 240.244
R4215 gnd.n3021 gnd.n2372 240.244
R4216 gnd.n3018 gnd.n2372 240.244
R4217 gnd.n3018 gnd.n2361 240.244
R4218 gnd.n3015 gnd.n2361 240.244
R4219 gnd.n3015 gnd.n2339 240.244
R4220 gnd.n3091 gnd.n2339 240.244
R4221 gnd.n3091 gnd.n2335 240.244
R4222 gnd.n3112 gnd.n2335 240.244
R4223 gnd.n3112 gnd.n2324 240.244
R4224 gnd.n3108 gnd.n2324 240.244
R4225 gnd.n3108 gnd.n2317 240.244
R4226 gnd.n3105 gnd.n2317 240.244
R4227 gnd.n3105 gnd.n2306 240.244
R4228 gnd.n3102 gnd.n2306 240.244
R4229 gnd.n3102 gnd.n2283 240.244
R4230 gnd.n3177 gnd.n2283 240.244
R4231 gnd.n3177 gnd.n2279 240.244
R4232 gnd.n3202 gnd.n2279 240.244
R4233 gnd.n3202 gnd.n2270 240.244
R4234 gnd.n3198 gnd.n2270 240.244
R4235 gnd.n3198 gnd.n2263 240.244
R4236 gnd.n3194 gnd.n2263 240.244
R4237 gnd.n3194 gnd.n2252 240.244
R4238 gnd.n3191 gnd.n2252 240.244
R4239 gnd.n3191 gnd.n2233 240.244
R4240 gnd.n3521 gnd.n2233 240.244
R4241 gnd.n2680 gnd.n2679 240.244
R4242 gnd.n2751 gnd.n2679 240.244
R4243 gnd.n2749 gnd.n2748 240.244
R4244 gnd.n2745 gnd.n2744 240.244
R4245 gnd.n2741 gnd.n2740 240.244
R4246 gnd.n2737 gnd.n2736 240.244
R4247 gnd.n2733 gnd.n2732 240.244
R4248 gnd.n2729 gnd.n2728 240.244
R4249 gnd.n2725 gnd.n2724 240.244
R4250 gnd.n2721 gnd.n2720 240.244
R4251 gnd.n2717 gnd.n2716 240.244
R4252 gnd.n2713 gnd.n2712 240.244
R4253 gnd.n2709 gnd.n2667 240.244
R4254 gnd.n2769 gnd.n2661 240.244
R4255 gnd.n2769 gnd.n2657 240.244
R4256 gnd.n2775 gnd.n2657 240.244
R4257 gnd.n2775 gnd.n2650 240.244
R4258 gnd.n2785 gnd.n2650 240.244
R4259 gnd.n2785 gnd.n2646 240.244
R4260 gnd.n2791 gnd.n2646 240.244
R4261 gnd.n2791 gnd.n2637 240.244
R4262 gnd.n2831 gnd.n2637 240.244
R4263 gnd.n2831 gnd.n2588 240.244
R4264 gnd.n2839 gnd.n2588 240.244
R4265 gnd.n2839 gnd.n2589 240.244
R4266 gnd.n2589 gnd.n2567 240.244
R4267 gnd.n2860 gnd.n2567 240.244
R4268 gnd.n2860 gnd.n2559 240.244
R4269 gnd.n2871 gnd.n2559 240.244
R4270 gnd.n2871 gnd.n2560 240.244
R4271 gnd.n2560 gnd.n2541 240.244
R4272 gnd.n2891 gnd.n2541 240.244
R4273 gnd.n2891 gnd.n2531 240.244
R4274 gnd.n2901 gnd.n2531 240.244
R4275 gnd.n2901 gnd.n2512 240.244
R4276 gnd.n2922 gnd.n2512 240.244
R4277 gnd.n2922 gnd.n2514 240.244
R4278 gnd.n2514 gnd.n2495 240.244
R4279 gnd.n2950 gnd.n2495 240.244
R4280 gnd.n2950 gnd.n2437 240.244
R4281 gnd.n3002 gnd.n2437 240.244
R4282 gnd.n3002 gnd.n2438 240.244
R4283 gnd.n2998 gnd.n2438 240.244
R4284 gnd.n2998 gnd.n2444 240.244
R4285 gnd.n2459 gnd.n2444 240.244
R4286 gnd.n2988 gnd.n2459 240.244
R4287 gnd.n2988 gnd.n2460 240.244
R4288 gnd.n2984 gnd.n2460 240.244
R4289 gnd.n2984 gnd.n2466 240.244
R4290 gnd.n2466 gnd.n2377 240.244
R4291 gnd.n3041 gnd.n2377 240.244
R4292 gnd.n3041 gnd.n2370 240.244
R4293 gnd.n3052 gnd.n2370 240.244
R4294 gnd.n3052 gnd.n2363 240.244
R4295 gnd.n3067 gnd.n2363 240.244
R4296 gnd.n3067 gnd.n2364 240.244
R4297 gnd.n2364 gnd.n2342 240.244
R4298 gnd.n3089 gnd.n2342 240.244
R4299 gnd.n3089 gnd.n2343 240.244
R4300 gnd.n2343 gnd.n2322 240.244
R4301 gnd.n3126 gnd.n2322 240.244
R4302 gnd.n3126 gnd.n2315 240.244
R4303 gnd.n3138 gnd.n2315 240.244
R4304 gnd.n3138 gnd.n2308 240.244
R4305 gnd.n3153 gnd.n2308 240.244
R4306 gnd.n3153 gnd.n2309 240.244
R4307 gnd.n2309 gnd.n2286 240.244
R4308 gnd.n3175 gnd.n2286 240.244
R4309 gnd.n3175 gnd.n2288 240.244
R4310 gnd.n2288 gnd.n2268 240.244
R4311 gnd.n3216 gnd.n2268 240.244
R4312 gnd.n3216 gnd.n2261 240.244
R4313 gnd.n3227 gnd.n2261 240.244
R4314 gnd.n3227 gnd.n2254 240.244
R4315 gnd.n3496 gnd.n2254 240.244
R4316 gnd.n3496 gnd.n2255 240.244
R4317 gnd.n2255 gnd.n2236 240.244
R4318 gnd.n3519 gnd.n2236 240.244
R4319 gnd.n6989 gnd.n6988 240.244
R4320 gnd.n6994 gnd.n6991 240.244
R4321 gnd.n6997 gnd.n6996 240.244
R4322 gnd.n7002 gnd.n6999 240.244
R4323 gnd.n7005 gnd.n7004 240.244
R4324 gnd.n7010 gnd.n7007 240.244
R4325 gnd.n7013 gnd.n7012 240.244
R4326 gnd.n7018 gnd.n7015 240.244
R4327 gnd.n7024 gnd.n7020 240.244
R4328 gnd.n5613 gnd.n1128 240.244
R4329 gnd.n5613 gnd.n1140 240.244
R4330 gnd.n5620 gnd.n1140 240.244
R4331 gnd.n5620 gnd.n1258 240.244
R4332 gnd.n1258 gnd.n1248 240.244
R4333 gnd.n5699 gnd.n1248 240.244
R4334 gnd.n5699 gnd.n1243 240.244
R4335 gnd.n5706 gnd.n1243 240.244
R4336 gnd.n5706 gnd.n1232 240.244
R4337 gnd.n1232 gnd.n1219 240.244
R4338 gnd.n5731 gnd.n1219 240.244
R4339 gnd.n5731 gnd.n1214 240.244
R4340 gnd.n5738 gnd.n1214 240.244
R4341 gnd.n5738 gnd.n1203 240.244
R4342 gnd.n1203 gnd.n1193 240.244
R4343 gnd.n5764 gnd.n1193 240.244
R4344 gnd.n5764 gnd.n1186 240.244
R4345 gnd.n5771 gnd.n1186 240.244
R4346 gnd.n5771 gnd.n1187 240.244
R4347 gnd.n1187 gnd.n1179 240.244
R4348 gnd.n1179 gnd.n1178 240.244
R4349 gnd.n1178 gnd.n54 240.244
R4350 gnd.n55 gnd.n54 240.244
R4351 gnd.n56 gnd.n55 240.244
R4352 gnd.n6920 gnd.n56 240.244
R4353 gnd.n6920 gnd.n59 240.244
R4354 gnd.n60 gnd.n59 240.244
R4355 gnd.n61 gnd.n60 240.244
R4356 gnd.n6911 gnd.n61 240.244
R4357 gnd.n6911 gnd.n64 240.244
R4358 gnd.n65 gnd.n64 240.244
R4359 gnd.n66 gnd.n65 240.244
R4360 gnd.n265 gnd.n66 240.244
R4361 gnd.n265 gnd.n69 240.244
R4362 gnd.n70 gnd.n69 240.244
R4363 gnd.n71 gnd.n70 240.244
R4364 gnd.n179 gnd.n71 240.244
R4365 gnd.n179 gnd.n74 240.244
R4366 gnd.n75 gnd.n74 240.244
R4367 gnd.n76 gnd.n75 240.244
R4368 gnd.n79 gnd.n76 240.244
R4369 gnd.n7151 gnd.n79 240.244
R4370 gnd.n5210 gnd.n5208 240.244
R4371 gnd.n5225 gnd.n5191 240.244
R4372 gnd.n5229 gnd.n5227 240.244
R4373 gnd.n5244 gnd.n5182 240.244
R4374 gnd.n5248 gnd.n5246 240.244
R4375 gnd.n5263 gnd.n5173 240.244
R4376 gnd.n5267 gnd.n5265 240.244
R4377 gnd.n5284 gnd.n5164 240.244
R4378 gnd.n5287 gnd.n5286 240.244
R4379 gnd.n1142 gnd.n1130 240.244
R4380 gnd.n5844 gnd.n1142 240.244
R4381 gnd.n5844 gnd.n1143 240.244
R4382 gnd.n1148 gnd.n1143 240.244
R4383 gnd.n1149 gnd.n1148 240.244
R4384 gnd.n1150 gnd.n1149 240.244
R4385 gnd.n1240 gnd.n1150 240.244
R4386 gnd.n1240 gnd.n1153 240.244
R4387 gnd.n1154 gnd.n1153 240.244
R4388 gnd.n1155 gnd.n1154 240.244
R4389 gnd.n1223 gnd.n1155 240.244
R4390 gnd.n1223 gnd.n1158 240.244
R4391 gnd.n1159 gnd.n1158 240.244
R4392 gnd.n1160 gnd.n1159 240.244
R4393 gnd.n1204 gnd.n1160 240.244
R4394 gnd.n1204 gnd.n1163 240.244
R4395 gnd.n1164 gnd.n1163 240.244
R4396 gnd.n1165 gnd.n1164 240.244
R4397 gnd.n1175 gnd.n1165 240.244
R4398 gnd.n1175 gnd.n1168 240.244
R4399 gnd.n1169 gnd.n1168 240.244
R4400 gnd.n5811 gnd.n1169 240.244
R4401 gnd.n5811 gnd.n230 240.244
R4402 gnd.n6933 gnd.n230 240.244
R4403 gnd.n6933 gnd.n226 240.244
R4404 gnd.n6939 gnd.n226 240.244
R4405 gnd.n6939 gnd.n208 240.244
R4406 gnd.n6949 gnd.n208 240.244
R4407 gnd.n6949 gnd.n204 240.244
R4408 gnd.n6955 gnd.n204 240.244
R4409 gnd.n6955 gnd.n193 240.244
R4410 gnd.n6965 gnd.n193 240.244
R4411 gnd.n6965 gnd.n189 240.244
R4412 gnd.n6971 gnd.n189 240.244
R4413 gnd.n6971 gnd.n176 240.244
R4414 gnd.n6981 gnd.n176 240.244
R4415 gnd.n6981 gnd.n170 240.244
R4416 gnd.n7061 gnd.n170 240.244
R4417 gnd.n7061 gnd.n171 240.244
R4418 gnd.n171 gnd.n162 240.244
R4419 gnd.n6986 gnd.n162 240.244
R4420 gnd.n6986 gnd.n84 240.244
R4421 gnd.n4135 gnd.n997 240.244
R4422 gnd.n4138 gnd.n4137 240.244
R4423 gnd.n4148 gnd.n4140 240.244
R4424 gnd.n4151 gnd.n4150 240.244
R4425 gnd.n4160 gnd.n4159 240.244
R4426 gnd.n4171 gnd.n4162 240.244
R4427 gnd.n4174 gnd.n4173 240.244
R4428 gnd.n4183 gnd.n4182 240.244
R4429 gnd.n4194 gnd.n4185 240.244
R4430 gnd.n3639 gnd.n2153 240.244
R4431 gnd.n2153 gnd.n2142 240.244
R4432 gnd.n3869 gnd.n2142 240.244
R4433 gnd.n3870 gnd.n3869 240.244
R4434 gnd.n3870 gnd.n829 240.244
R4435 gnd.n3873 gnd.n829 240.244
R4436 gnd.n3873 gnd.n842 240.244
R4437 gnd.n3880 gnd.n842 240.244
R4438 gnd.n3880 gnd.n854 240.244
R4439 gnd.n3900 gnd.n854 240.244
R4440 gnd.n3900 gnd.n864 240.244
R4441 gnd.n3896 gnd.n864 240.244
R4442 gnd.n3896 gnd.n875 240.244
R4443 gnd.n3930 gnd.n875 240.244
R4444 gnd.n3930 gnd.n885 240.244
R4445 gnd.n3938 gnd.n885 240.244
R4446 gnd.n3938 gnd.n896 240.244
R4447 gnd.n2110 gnd.n896 240.244
R4448 gnd.n3977 gnd.n2110 240.244
R4449 gnd.n3977 gnd.n2106 240.244
R4450 gnd.n3983 gnd.n2106 240.244
R4451 gnd.n3983 gnd.n2076 240.244
R4452 gnd.n4005 gnd.n2076 240.244
R4453 gnd.n4005 gnd.n2072 240.244
R4454 gnd.n4011 gnd.n2072 240.244
R4455 gnd.n4011 gnd.n911 240.244
R4456 gnd.n4026 gnd.n911 240.244
R4457 gnd.n4026 gnd.n922 240.244
R4458 gnd.n4032 gnd.n922 240.244
R4459 gnd.n4032 gnd.n932 240.244
R4460 gnd.n4077 gnd.n932 240.244
R4461 gnd.n4077 gnd.n942 240.244
R4462 gnd.n2049 gnd.n942 240.244
R4463 gnd.n2049 gnd.n953 240.244
R4464 gnd.n2050 gnd.n953 240.244
R4465 gnd.n2050 gnd.n963 240.244
R4466 gnd.n2053 gnd.n963 240.244
R4467 gnd.n2053 gnd.n974 240.244
R4468 gnd.n4062 gnd.n974 240.244
R4469 gnd.n4062 gnd.n985 240.244
R4470 gnd.n4298 gnd.n985 240.244
R4471 gnd.n4298 gnd.n995 240.244
R4472 gnd.n3651 gnd.n2160 240.244
R4473 gnd.n3655 gnd.n3654 240.244
R4474 gnd.n3661 gnd.n3660 240.244
R4475 gnd.n3665 gnd.n3664 240.244
R4476 gnd.n3671 gnd.n3670 240.244
R4477 gnd.n3675 gnd.n3674 240.244
R4478 gnd.n3681 gnd.n3680 240.244
R4479 gnd.n3685 gnd.n3684 240.244
R4480 gnd.n3698 gnd.n3638 240.244
R4481 gnd.n3858 gnd.n2154 240.244
R4482 gnd.n3858 gnd.n2155 240.244
R4483 gnd.n2155 gnd.n2145 240.244
R4484 gnd.n3851 gnd.n2145 240.244
R4485 gnd.n3851 gnd.n831 240.244
R4486 gnd.n844 gnd.n831 240.244
R4487 gnd.n6083 gnd.n844 240.244
R4488 gnd.n6083 gnd.n845 240.244
R4489 gnd.n6079 gnd.n845 240.244
R4490 gnd.n6079 gnd.n851 240.244
R4491 gnd.n6071 gnd.n851 240.244
R4492 gnd.n6071 gnd.n866 240.244
R4493 gnd.n6067 gnd.n866 240.244
R4494 gnd.n6067 gnd.n872 240.244
R4495 gnd.n6059 gnd.n872 240.244
R4496 gnd.n6059 gnd.n887 240.244
R4497 gnd.n6055 gnd.n887 240.244
R4498 gnd.n6055 gnd.n893 240.244
R4499 gnd.n3966 gnd.n893 240.244
R4500 gnd.n3972 gnd.n3966 240.244
R4501 gnd.n3972 gnd.n2086 240.244
R4502 gnd.n3997 gnd.n2086 240.244
R4503 gnd.n3997 gnd.n2080 240.244
R4504 gnd.n3993 gnd.n2080 240.244
R4505 gnd.n3993 gnd.n913 240.244
R4506 gnd.n6045 gnd.n913 240.244
R4507 gnd.n6045 gnd.n914 240.244
R4508 gnd.n6041 gnd.n914 240.244
R4509 gnd.n6041 gnd.n920 240.244
R4510 gnd.n6033 gnd.n920 240.244
R4511 gnd.n6033 gnd.n933 240.244
R4512 gnd.n6029 gnd.n933 240.244
R4513 gnd.n6029 gnd.n939 240.244
R4514 gnd.n6021 gnd.n939 240.244
R4515 gnd.n6021 gnd.n955 240.244
R4516 gnd.n6017 gnd.n955 240.244
R4517 gnd.n6017 gnd.n961 240.244
R4518 gnd.n6009 gnd.n961 240.244
R4519 gnd.n6009 gnd.n976 240.244
R4520 gnd.n6005 gnd.n976 240.244
R4521 gnd.n6005 gnd.n982 240.244
R4522 gnd.n5997 gnd.n982 240.244
R4523 gnd.n6266 gnd.n656 240.244
R4524 gnd.n6266 gnd.n654 240.244
R4525 gnd.n6270 gnd.n654 240.244
R4526 gnd.n6270 gnd.n650 240.244
R4527 gnd.n6276 gnd.n650 240.244
R4528 gnd.n6276 gnd.n648 240.244
R4529 gnd.n6280 gnd.n648 240.244
R4530 gnd.n6280 gnd.n644 240.244
R4531 gnd.n6286 gnd.n644 240.244
R4532 gnd.n6286 gnd.n642 240.244
R4533 gnd.n6290 gnd.n642 240.244
R4534 gnd.n6290 gnd.n638 240.244
R4535 gnd.n6296 gnd.n638 240.244
R4536 gnd.n6296 gnd.n636 240.244
R4537 gnd.n6300 gnd.n636 240.244
R4538 gnd.n6300 gnd.n632 240.244
R4539 gnd.n6306 gnd.n632 240.244
R4540 gnd.n6306 gnd.n630 240.244
R4541 gnd.n6310 gnd.n630 240.244
R4542 gnd.n6310 gnd.n626 240.244
R4543 gnd.n6316 gnd.n626 240.244
R4544 gnd.n6316 gnd.n624 240.244
R4545 gnd.n6320 gnd.n624 240.244
R4546 gnd.n6320 gnd.n620 240.244
R4547 gnd.n6326 gnd.n620 240.244
R4548 gnd.n6326 gnd.n618 240.244
R4549 gnd.n6330 gnd.n618 240.244
R4550 gnd.n6330 gnd.n614 240.244
R4551 gnd.n6336 gnd.n614 240.244
R4552 gnd.n6336 gnd.n612 240.244
R4553 gnd.n6340 gnd.n612 240.244
R4554 gnd.n6340 gnd.n608 240.244
R4555 gnd.n6346 gnd.n608 240.244
R4556 gnd.n6346 gnd.n606 240.244
R4557 gnd.n6350 gnd.n606 240.244
R4558 gnd.n6350 gnd.n602 240.244
R4559 gnd.n6356 gnd.n602 240.244
R4560 gnd.n6356 gnd.n600 240.244
R4561 gnd.n6360 gnd.n600 240.244
R4562 gnd.n6360 gnd.n596 240.244
R4563 gnd.n6366 gnd.n596 240.244
R4564 gnd.n6366 gnd.n594 240.244
R4565 gnd.n6370 gnd.n594 240.244
R4566 gnd.n6370 gnd.n590 240.244
R4567 gnd.n6376 gnd.n590 240.244
R4568 gnd.n6376 gnd.n588 240.244
R4569 gnd.n6380 gnd.n588 240.244
R4570 gnd.n6380 gnd.n584 240.244
R4571 gnd.n6386 gnd.n584 240.244
R4572 gnd.n6386 gnd.n582 240.244
R4573 gnd.n6390 gnd.n582 240.244
R4574 gnd.n6390 gnd.n578 240.244
R4575 gnd.n6396 gnd.n578 240.244
R4576 gnd.n6396 gnd.n576 240.244
R4577 gnd.n6400 gnd.n576 240.244
R4578 gnd.n6400 gnd.n572 240.244
R4579 gnd.n6406 gnd.n572 240.244
R4580 gnd.n6406 gnd.n570 240.244
R4581 gnd.n6410 gnd.n570 240.244
R4582 gnd.n6410 gnd.n566 240.244
R4583 gnd.n6416 gnd.n566 240.244
R4584 gnd.n6416 gnd.n564 240.244
R4585 gnd.n6420 gnd.n564 240.244
R4586 gnd.n6420 gnd.n560 240.244
R4587 gnd.n6426 gnd.n560 240.244
R4588 gnd.n6426 gnd.n558 240.244
R4589 gnd.n6430 gnd.n558 240.244
R4590 gnd.n6430 gnd.n554 240.244
R4591 gnd.n6436 gnd.n554 240.244
R4592 gnd.n6436 gnd.n552 240.244
R4593 gnd.n6440 gnd.n552 240.244
R4594 gnd.n6440 gnd.n548 240.244
R4595 gnd.n6446 gnd.n548 240.244
R4596 gnd.n6446 gnd.n546 240.244
R4597 gnd.n6450 gnd.n546 240.244
R4598 gnd.n6450 gnd.n542 240.244
R4599 gnd.n6456 gnd.n542 240.244
R4600 gnd.n6456 gnd.n540 240.244
R4601 gnd.n6460 gnd.n540 240.244
R4602 gnd.n6460 gnd.n536 240.244
R4603 gnd.n6466 gnd.n536 240.244
R4604 gnd.n6466 gnd.n534 240.244
R4605 gnd.n6470 gnd.n534 240.244
R4606 gnd.n6470 gnd.n530 240.244
R4607 gnd.n6476 gnd.n530 240.244
R4608 gnd.n6476 gnd.n528 240.244
R4609 gnd.n6480 gnd.n528 240.244
R4610 gnd.n6480 gnd.n524 240.244
R4611 gnd.n6486 gnd.n524 240.244
R4612 gnd.n6486 gnd.n522 240.244
R4613 gnd.n6490 gnd.n522 240.244
R4614 gnd.n6490 gnd.n518 240.244
R4615 gnd.n6496 gnd.n518 240.244
R4616 gnd.n6496 gnd.n516 240.244
R4617 gnd.n6500 gnd.n516 240.244
R4618 gnd.n6500 gnd.n512 240.244
R4619 gnd.n6506 gnd.n512 240.244
R4620 gnd.n6506 gnd.n510 240.244
R4621 gnd.n6510 gnd.n510 240.244
R4622 gnd.n6510 gnd.n506 240.244
R4623 gnd.n6516 gnd.n506 240.244
R4624 gnd.n6516 gnd.n504 240.244
R4625 gnd.n6520 gnd.n504 240.244
R4626 gnd.n6520 gnd.n500 240.244
R4627 gnd.n6526 gnd.n500 240.244
R4628 gnd.n6526 gnd.n498 240.244
R4629 gnd.n6530 gnd.n498 240.244
R4630 gnd.n6530 gnd.n494 240.244
R4631 gnd.n6536 gnd.n494 240.244
R4632 gnd.n6536 gnd.n492 240.244
R4633 gnd.n6540 gnd.n492 240.244
R4634 gnd.n6540 gnd.n488 240.244
R4635 gnd.n6546 gnd.n488 240.244
R4636 gnd.n6546 gnd.n486 240.244
R4637 gnd.n6550 gnd.n486 240.244
R4638 gnd.n6550 gnd.n482 240.244
R4639 gnd.n6556 gnd.n482 240.244
R4640 gnd.n6556 gnd.n480 240.244
R4641 gnd.n6560 gnd.n480 240.244
R4642 gnd.n6560 gnd.n476 240.244
R4643 gnd.n6566 gnd.n476 240.244
R4644 gnd.n6566 gnd.n474 240.244
R4645 gnd.n6570 gnd.n474 240.244
R4646 gnd.n6570 gnd.n470 240.244
R4647 gnd.n6576 gnd.n470 240.244
R4648 gnd.n6576 gnd.n468 240.244
R4649 gnd.n6580 gnd.n468 240.244
R4650 gnd.n6580 gnd.n464 240.244
R4651 gnd.n6586 gnd.n464 240.244
R4652 gnd.n6586 gnd.n462 240.244
R4653 gnd.n6590 gnd.n462 240.244
R4654 gnd.n6590 gnd.n458 240.244
R4655 gnd.n6596 gnd.n458 240.244
R4656 gnd.n6596 gnd.n456 240.244
R4657 gnd.n6600 gnd.n456 240.244
R4658 gnd.n6600 gnd.n452 240.244
R4659 gnd.n6606 gnd.n452 240.244
R4660 gnd.n6606 gnd.n450 240.244
R4661 gnd.n6610 gnd.n450 240.244
R4662 gnd.n6610 gnd.n446 240.244
R4663 gnd.n6616 gnd.n446 240.244
R4664 gnd.n6616 gnd.n444 240.244
R4665 gnd.n6620 gnd.n444 240.244
R4666 gnd.n6620 gnd.n440 240.244
R4667 gnd.n6626 gnd.n440 240.244
R4668 gnd.n6626 gnd.n438 240.244
R4669 gnd.n6630 gnd.n438 240.244
R4670 gnd.n6630 gnd.n434 240.244
R4671 gnd.n6636 gnd.n434 240.244
R4672 gnd.n6636 gnd.n432 240.244
R4673 gnd.n6640 gnd.n432 240.244
R4674 gnd.n6640 gnd.n428 240.244
R4675 gnd.n6646 gnd.n428 240.244
R4676 gnd.n6646 gnd.n426 240.244
R4677 gnd.n6650 gnd.n426 240.244
R4678 gnd.n6650 gnd.n422 240.244
R4679 gnd.n6656 gnd.n422 240.244
R4680 gnd.n6656 gnd.n420 240.244
R4681 gnd.n6660 gnd.n420 240.244
R4682 gnd.n6660 gnd.n416 240.244
R4683 gnd.n6666 gnd.n416 240.244
R4684 gnd.n6666 gnd.n414 240.244
R4685 gnd.n6670 gnd.n414 240.244
R4686 gnd.n6670 gnd.n410 240.244
R4687 gnd.n6676 gnd.n410 240.244
R4688 gnd.n6676 gnd.n408 240.244
R4689 gnd.n6680 gnd.n408 240.244
R4690 gnd.n6686 gnd.n404 240.244
R4691 gnd.n6686 gnd.n402 240.244
R4692 gnd.n6690 gnd.n402 240.244
R4693 gnd.n6690 gnd.n398 240.244
R4694 gnd.n6696 gnd.n398 240.244
R4695 gnd.n6696 gnd.n396 240.244
R4696 gnd.n6700 gnd.n396 240.244
R4697 gnd.n6700 gnd.n392 240.244
R4698 gnd.n6706 gnd.n392 240.244
R4699 gnd.n6706 gnd.n390 240.244
R4700 gnd.n6710 gnd.n390 240.244
R4701 gnd.n6710 gnd.n386 240.244
R4702 gnd.n6716 gnd.n386 240.244
R4703 gnd.n6716 gnd.n384 240.244
R4704 gnd.n6720 gnd.n384 240.244
R4705 gnd.n6720 gnd.n380 240.244
R4706 gnd.n6726 gnd.n380 240.244
R4707 gnd.n6726 gnd.n378 240.244
R4708 gnd.n6730 gnd.n378 240.244
R4709 gnd.n6730 gnd.n374 240.244
R4710 gnd.n6736 gnd.n374 240.244
R4711 gnd.n6736 gnd.n372 240.244
R4712 gnd.n6740 gnd.n372 240.244
R4713 gnd.n6740 gnd.n368 240.244
R4714 gnd.n6746 gnd.n368 240.244
R4715 gnd.n6746 gnd.n366 240.244
R4716 gnd.n6750 gnd.n366 240.244
R4717 gnd.n6750 gnd.n362 240.244
R4718 gnd.n6756 gnd.n362 240.244
R4719 gnd.n6756 gnd.n360 240.244
R4720 gnd.n6760 gnd.n360 240.244
R4721 gnd.n6760 gnd.n356 240.244
R4722 gnd.n6766 gnd.n356 240.244
R4723 gnd.n6766 gnd.n354 240.244
R4724 gnd.n6770 gnd.n354 240.244
R4725 gnd.n6770 gnd.n350 240.244
R4726 gnd.n6776 gnd.n350 240.244
R4727 gnd.n6776 gnd.n348 240.244
R4728 gnd.n6780 gnd.n348 240.244
R4729 gnd.n6780 gnd.n344 240.244
R4730 gnd.n6786 gnd.n344 240.244
R4731 gnd.n6786 gnd.n342 240.244
R4732 gnd.n6790 gnd.n342 240.244
R4733 gnd.n6790 gnd.n338 240.244
R4734 gnd.n6796 gnd.n338 240.244
R4735 gnd.n6796 gnd.n336 240.244
R4736 gnd.n6800 gnd.n336 240.244
R4737 gnd.n6800 gnd.n332 240.244
R4738 gnd.n6806 gnd.n332 240.244
R4739 gnd.n6806 gnd.n330 240.244
R4740 gnd.n6810 gnd.n330 240.244
R4741 gnd.n6810 gnd.n326 240.244
R4742 gnd.n6816 gnd.n326 240.244
R4743 gnd.n6816 gnd.n324 240.244
R4744 gnd.n6820 gnd.n324 240.244
R4745 gnd.n6820 gnd.n320 240.244
R4746 gnd.n6826 gnd.n320 240.244
R4747 gnd.n6826 gnd.n318 240.244
R4748 gnd.n6830 gnd.n318 240.244
R4749 gnd.n6830 gnd.n314 240.244
R4750 gnd.n6836 gnd.n314 240.244
R4751 gnd.n6836 gnd.n312 240.244
R4752 gnd.n6840 gnd.n312 240.244
R4753 gnd.n6840 gnd.n308 240.244
R4754 gnd.n6846 gnd.n308 240.244
R4755 gnd.n6846 gnd.n306 240.244
R4756 gnd.n6850 gnd.n306 240.244
R4757 gnd.n6850 gnd.n302 240.244
R4758 gnd.n6856 gnd.n302 240.244
R4759 gnd.n6856 gnd.n300 240.244
R4760 gnd.n6860 gnd.n300 240.244
R4761 gnd.n6860 gnd.n296 240.244
R4762 gnd.n6866 gnd.n296 240.244
R4763 gnd.n6866 gnd.n294 240.244
R4764 gnd.n6870 gnd.n294 240.244
R4765 gnd.n6870 gnd.n290 240.244
R4766 gnd.n6876 gnd.n290 240.244
R4767 gnd.n6876 gnd.n288 240.244
R4768 gnd.n6880 gnd.n288 240.244
R4769 gnd.n6880 gnd.n284 240.244
R4770 gnd.n6888 gnd.n284 240.244
R4771 gnd.n6888 gnd.n282 240.244
R4772 gnd.n6892 gnd.n282 240.244
R4773 gnd.n6893 gnd.n6892 240.244
R4774 gnd.n3909 gnd.n826 240.244
R4775 gnd.n3910 gnd.n3909 240.244
R4776 gnd.n3910 gnd.n3903 240.244
R4777 gnd.n3916 gnd.n3903 240.244
R4778 gnd.n3917 gnd.n3916 240.244
R4779 gnd.n3918 gnd.n3917 240.244
R4780 gnd.n3918 gnd.n2124 240.244
R4781 gnd.n3927 gnd.n2124 240.244
R4782 gnd.n3927 gnd.n2125 240.244
R4783 gnd.n2125 gnd.n2116 240.244
R4784 gnd.n3951 gnd.n2116 240.244
R4785 gnd.n3951 gnd.n2113 240.244
R4786 gnd.n3964 gnd.n2113 240.244
R4787 gnd.n3964 gnd.n2114 240.244
R4788 gnd.n3959 gnd.n2114 240.244
R4789 gnd.n3959 gnd.n3958 240.244
R4790 gnd.n3958 gnd.n2068 240.244
R4791 gnd.n4014 gnd.n2068 240.244
R4792 gnd.n4015 gnd.n4014 240.244
R4793 gnd.n4015 gnd.n2065 240.244
R4794 gnd.n4023 gnd.n2065 240.244
R4795 gnd.n4023 gnd.n2066 240.244
R4796 gnd.n2066 gnd.n2043 240.244
R4797 gnd.n4080 gnd.n2043 240.244
R4798 gnd.n4080 gnd.n2039 240.244
R4799 gnd.n4086 gnd.n2039 240.244
R4800 gnd.n4087 gnd.n4086 240.244
R4801 gnd.n4088 gnd.n4087 240.244
R4802 gnd.n4088 gnd.n2035 240.244
R4803 gnd.n4094 gnd.n2035 240.244
R4804 gnd.n4095 gnd.n4094 240.244
R4805 gnd.n4096 gnd.n4095 240.244
R4806 gnd.n4096 gnd.n2031 240.244
R4807 gnd.n4102 gnd.n2031 240.244
R4808 gnd.n4103 gnd.n4102 240.244
R4809 gnd.n4104 gnd.n4103 240.244
R4810 gnd.n4104 gnd.n2027 240.244
R4811 gnd.n4110 gnd.n2027 240.244
R4812 gnd.n4110 gnd.n2025 240.244
R4813 gnd.n4246 gnd.n2025 240.244
R4814 gnd.n4246 gnd.n2021 240.244
R4815 gnd.n4252 gnd.n2021 240.244
R4816 gnd.n4252 gnd.n1772 240.244
R4817 gnd.n4415 gnd.n1772 240.244
R4818 gnd.n4415 gnd.n1768 240.244
R4819 gnd.n4421 gnd.n1768 240.244
R4820 gnd.n4421 gnd.n1757 240.244
R4821 gnd.n4460 gnd.n1757 240.244
R4822 gnd.n4460 gnd.n1752 240.244
R4823 gnd.n4468 gnd.n1752 240.244
R4824 gnd.n4468 gnd.n1753 240.244
R4825 gnd.n1753 gnd.n1729 240.244
R4826 gnd.n4511 gnd.n1729 240.244
R4827 gnd.n4511 gnd.n1725 240.244
R4828 gnd.n4517 gnd.n1725 240.244
R4829 gnd.n4517 gnd.n1709 240.244
R4830 gnd.n4548 gnd.n1709 240.244
R4831 gnd.n4548 gnd.n1705 240.244
R4832 gnd.n4554 gnd.n1705 240.244
R4833 gnd.n4554 gnd.n1683 240.244
R4834 gnd.n4589 gnd.n1683 240.244
R4835 gnd.n4589 gnd.n1679 240.244
R4836 gnd.n4595 gnd.n1679 240.244
R4837 gnd.n4595 gnd.n1667 240.244
R4838 gnd.n4634 gnd.n1667 240.244
R4839 gnd.n4634 gnd.n1662 240.244
R4840 gnd.n4642 gnd.n1662 240.244
R4841 gnd.n4642 gnd.n1663 240.244
R4842 gnd.n1663 gnd.n1639 240.244
R4843 gnd.n4706 gnd.n1639 240.244
R4844 gnd.n4706 gnd.n1635 240.244
R4845 gnd.n4712 gnd.n1635 240.244
R4846 gnd.n4712 gnd.n1618 240.244
R4847 gnd.n4733 gnd.n1618 240.244
R4848 gnd.n4733 gnd.n1614 240.244
R4849 gnd.n4739 gnd.n1614 240.244
R4850 gnd.n4739 gnd.n1597 240.244
R4851 gnd.n4766 gnd.n1597 240.244
R4852 gnd.n4766 gnd.n1593 240.244
R4853 gnd.n4772 gnd.n1593 240.244
R4854 gnd.n4772 gnd.n1580 240.244
R4855 gnd.n4811 gnd.n1580 240.244
R4856 gnd.n4811 gnd.n1575 240.244
R4857 gnd.n4819 gnd.n1575 240.244
R4858 gnd.n4819 gnd.n1576 240.244
R4859 gnd.n1576 gnd.n1551 240.244
R4860 gnd.n4859 gnd.n1551 240.244
R4861 gnd.n4859 gnd.n1547 240.244
R4862 gnd.n4865 gnd.n1547 240.244
R4863 gnd.n4865 gnd.n1531 240.244
R4864 gnd.n4887 gnd.n1531 240.244
R4865 gnd.n4887 gnd.n1526 240.244
R4866 gnd.n4901 gnd.n1526 240.244
R4867 gnd.n4901 gnd.n1527 240.244
R4868 gnd.n4897 gnd.n1527 240.244
R4869 gnd.n4897 gnd.n1499 240.244
R4870 gnd.n4962 gnd.n1499 240.244
R4871 gnd.n4962 gnd.n1494 240.244
R4872 gnd.n4970 gnd.n1494 240.244
R4873 gnd.n4970 gnd.n1495 240.244
R4874 gnd.n1495 gnd.n1471 240.244
R4875 gnd.n5013 gnd.n1471 240.244
R4876 gnd.n5013 gnd.n1467 240.244
R4877 gnd.n5021 gnd.n1467 240.244
R4878 gnd.n5021 gnd.n1453 240.244
R4879 gnd.n5039 gnd.n1453 240.244
R4880 gnd.n5040 gnd.n5039 240.244
R4881 gnd.n5040 gnd.n1449 240.244
R4882 gnd.n5046 gnd.n1449 240.244
R4883 gnd.n5046 gnd.n1396 240.244
R4884 gnd.n5083 gnd.n1396 240.244
R4885 gnd.n5083 gnd.n1392 240.244
R4886 gnd.n5089 gnd.n1392 240.244
R4887 gnd.n5089 gnd.n1375 240.244
R4888 gnd.n5112 gnd.n1375 240.244
R4889 gnd.n5112 gnd.n1370 240.244
R4890 gnd.n5121 gnd.n1370 240.244
R4891 gnd.n5121 gnd.n1371 240.244
R4892 gnd.n1371 gnd.n1341 240.244
R4893 gnd.n5334 gnd.n1341 240.244
R4894 gnd.n5334 gnd.n1342 240.244
R4895 gnd.n5330 gnd.n1342 240.244
R4896 gnd.n5330 gnd.n5329 240.244
R4897 gnd.n5329 gnd.n1109 240.244
R4898 gnd.n5865 gnd.n1109 240.244
R4899 gnd.n5865 gnd.n1110 240.244
R4900 gnd.n5861 gnd.n1110 240.244
R4901 gnd.n5861 gnd.n1116 240.244
R4902 gnd.n5857 gnd.n1116 240.244
R4903 gnd.n5857 gnd.n1119 240.244
R4904 gnd.n5853 gnd.n1119 240.244
R4905 gnd.n5853 gnd.n1125 240.244
R4906 gnd.n5677 gnd.n1125 240.244
R4907 gnd.n5678 gnd.n5677 240.244
R4908 gnd.n5678 gnd.n5671 240.244
R4909 gnd.n5686 gnd.n5671 240.244
R4910 gnd.n5686 gnd.n5672 240.244
R4911 gnd.n5672 gnd.n1239 240.244
R4912 gnd.n5709 gnd.n1239 240.244
R4913 gnd.n5709 gnd.n1234 240.244
R4914 gnd.n5717 gnd.n1234 240.244
R4915 gnd.n5717 gnd.n1235 240.244
R4916 gnd.n1235 gnd.n1211 240.244
R4917 gnd.n5741 gnd.n1211 240.244
R4918 gnd.n5741 gnd.n1206 240.244
R4919 gnd.n5755 gnd.n1206 240.244
R4920 gnd.n5755 gnd.n1207 240.244
R4921 gnd.n5751 gnd.n1207 240.244
R4922 gnd.n5751 gnd.n5750 240.244
R4923 gnd.n5750 gnd.n1174 240.244
R4924 gnd.n5784 gnd.n1174 240.244
R4925 gnd.n5784 gnd.n1171 240.244
R4926 gnd.n5808 gnd.n1171 240.244
R4927 gnd.n5808 gnd.n1172 240.244
R4928 gnd.n5803 gnd.n1172 240.244
R4929 gnd.n5803 gnd.n5802 240.244
R4930 gnd.n5802 gnd.n5801 240.244
R4931 gnd.n5801 gnd.n5789 240.244
R4932 gnd.n5797 gnd.n5789 240.244
R4933 gnd.n5797 gnd.n5796 240.244
R4934 gnd.n5796 gnd.n270 240.244
R4935 gnd.n6905 gnd.n270 240.244
R4936 gnd.n6905 gnd.n271 240.244
R4937 gnd.n6901 gnd.n271 240.244
R4938 gnd.n6901 gnd.n6900 240.244
R4939 gnd.n6900 gnd.n6899 240.244
R4940 gnd.n6899 gnd.n277 240.244
R4941 gnd.n6260 gnd.n660 240.244
R4942 gnd.n6256 gnd.n660 240.244
R4943 gnd.n6256 gnd.n662 240.244
R4944 gnd.n6252 gnd.n662 240.244
R4945 gnd.n6252 gnd.n667 240.244
R4946 gnd.n6248 gnd.n667 240.244
R4947 gnd.n6248 gnd.n669 240.244
R4948 gnd.n6244 gnd.n669 240.244
R4949 gnd.n6244 gnd.n675 240.244
R4950 gnd.n6240 gnd.n675 240.244
R4951 gnd.n6240 gnd.n677 240.244
R4952 gnd.n6236 gnd.n677 240.244
R4953 gnd.n6236 gnd.n683 240.244
R4954 gnd.n6232 gnd.n683 240.244
R4955 gnd.n6232 gnd.n685 240.244
R4956 gnd.n6228 gnd.n685 240.244
R4957 gnd.n6228 gnd.n691 240.244
R4958 gnd.n6224 gnd.n691 240.244
R4959 gnd.n6224 gnd.n693 240.244
R4960 gnd.n6220 gnd.n693 240.244
R4961 gnd.n6220 gnd.n699 240.244
R4962 gnd.n6216 gnd.n699 240.244
R4963 gnd.n6216 gnd.n701 240.244
R4964 gnd.n6212 gnd.n701 240.244
R4965 gnd.n6212 gnd.n707 240.244
R4966 gnd.n6208 gnd.n707 240.244
R4967 gnd.n6208 gnd.n709 240.244
R4968 gnd.n6204 gnd.n709 240.244
R4969 gnd.n6204 gnd.n715 240.244
R4970 gnd.n6200 gnd.n715 240.244
R4971 gnd.n6200 gnd.n717 240.244
R4972 gnd.n6196 gnd.n717 240.244
R4973 gnd.n6196 gnd.n723 240.244
R4974 gnd.n6192 gnd.n723 240.244
R4975 gnd.n6192 gnd.n725 240.244
R4976 gnd.n6188 gnd.n725 240.244
R4977 gnd.n6188 gnd.n731 240.244
R4978 gnd.n6184 gnd.n731 240.244
R4979 gnd.n6184 gnd.n733 240.244
R4980 gnd.n6180 gnd.n733 240.244
R4981 gnd.n6180 gnd.n739 240.244
R4982 gnd.n6176 gnd.n739 240.244
R4983 gnd.n6176 gnd.n741 240.244
R4984 gnd.n6172 gnd.n741 240.244
R4985 gnd.n6172 gnd.n747 240.244
R4986 gnd.n6168 gnd.n747 240.244
R4987 gnd.n6168 gnd.n749 240.244
R4988 gnd.n6164 gnd.n749 240.244
R4989 gnd.n6164 gnd.n755 240.244
R4990 gnd.n6160 gnd.n755 240.244
R4991 gnd.n6160 gnd.n757 240.244
R4992 gnd.n6156 gnd.n757 240.244
R4993 gnd.n6156 gnd.n763 240.244
R4994 gnd.n6152 gnd.n763 240.244
R4995 gnd.n6152 gnd.n765 240.244
R4996 gnd.n6148 gnd.n765 240.244
R4997 gnd.n6148 gnd.n771 240.244
R4998 gnd.n6144 gnd.n771 240.244
R4999 gnd.n6144 gnd.n773 240.244
R5000 gnd.n6140 gnd.n773 240.244
R5001 gnd.n6140 gnd.n779 240.244
R5002 gnd.n6136 gnd.n779 240.244
R5003 gnd.n6136 gnd.n781 240.244
R5004 gnd.n6132 gnd.n781 240.244
R5005 gnd.n6132 gnd.n787 240.244
R5006 gnd.n6128 gnd.n787 240.244
R5007 gnd.n6128 gnd.n789 240.244
R5008 gnd.n6124 gnd.n789 240.244
R5009 gnd.n6124 gnd.n795 240.244
R5010 gnd.n6120 gnd.n795 240.244
R5011 gnd.n6120 gnd.n797 240.244
R5012 gnd.n6116 gnd.n797 240.244
R5013 gnd.n6116 gnd.n803 240.244
R5014 gnd.n6112 gnd.n803 240.244
R5015 gnd.n6112 gnd.n805 240.244
R5016 gnd.n6108 gnd.n805 240.244
R5017 gnd.n6108 gnd.n811 240.244
R5018 gnd.n6104 gnd.n811 240.244
R5019 gnd.n6104 gnd.n813 240.244
R5020 gnd.n6100 gnd.n813 240.244
R5021 gnd.n6100 gnd.n819 240.244
R5022 gnd.n6096 gnd.n819 240.244
R5023 gnd.n6096 gnd.n821 240.244
R5024 gnd.n6092 gnd.n821 240.244
R5025 gnd.n1003 gnd.n1002 240.244
R5026 gnd.n1004 gnd.n1003 240.244
R5027 gnd.n4260 gnd.n1004 240.244
R5028 gnd.n4260 gnd.n1007 240.244
R5029 gnd.n1008 gnd.n1007 240.244
R5030 gnd.n1009 gnd.n1008 240.244
R5031 gnd.n4470 gnd.n1009 240.244
R5032 gnd.n4470 gnd.n1012 240.244
R5033 gnd.n1013 gnd.n1012 240.244
R5034 gnd.n1014 gnd.n1013 240.244
R5035 gnd.n4508 gnd.n1014 240.244
R5036 gnd.n4508 gnd.n1017 240.244
R5037 gnd.n1018 gnd.n1017 240.244
R5038 gnd.n1019 gnd.n1018 240.244
R5039 gnd.n4545 gnd.n1019 240.244
R5040 gnd.n4545 gnd.n1022 240.244
R5041 gnd.n1023 gnd.n1022 240.244
R5042 gnd.n1024 gnd.n1023 240.244
R5043 gnd.n1686 gnd.n1024 240.244
R5044 gnd.n1686 gnd.n1027 240.244
R5045 gnd.n1028 gnd.n1027 240.244
R5046 gnd.n1029 gnd.n1028 240.244
R5047 gnd.n1670 gnd.n1029 240.244
R5048 gnd.n1670 gnd.n1032 240.244
R5049 gnd.n1033 gnd.n1032 240.244
R5050 gnd.n1034 gnd.n1033 240.244
R5051 gnd.n4695 gnd.n1034 240.244
R5052 gnd.n4695 gnd.n1037 240.244
R5053 gnd.n1038 gnd.n1037 240.244
R5054 gnd.n1039 gnd.n1038 240.244
R5055 gnd.n1625 gnd.n1039 240.244
R5056 gnd.n1625 gnd.n1042 240.244
R5057 gnd.n1043 gnd.n1042 240.244
R5058 gnd.n1044 gnd.n1043 240.244
R5059 gnd.n1598 gnd.n1044 240.244
R5060 gnd.n1598 gnd.n1047 240.244
R5061 gnd.n1048 gnd.n1047 240.244
R5062 gnd.n1049 gnd.n1048 240.244
R5063 gnd.n1581 gnd.n1049 240.244
R5064 gnd.n1581 gnd.n1052 240.244
R5065 gnd.n1053 gnd.n1052 240.244
R5066 gnd.n1054 gnd.n1053 240.244
R5067 gnd.n4786 gnd.n1054 240.244
R5068 gnd.n4786 gnd.n1057 240.244
R5069 gnd.n1058 gnd.n1057 240.244
R5070 gnd.n1059 gnd.n1058 240.244
R5071 gnd.n1545 gnd.n1059 240.244
R5072 gnd.n1545 gnd.n1062 240.244
R5073 gnd.n1063 gnd.n1062 240.244
R5074 gnd.n1064 gnd.n1063 240.244
R5075 gnd.n4912 gnd.n1064 240.244
R5076 gnd.n4912 gnd.n1067 240.244
R5077 gnd.n1068 gnd.n1067 240.244
R5078 gnd.n1069 gnd.n1068 240.244
R5079 gnd.n1502 gnd.n1069 240.244
R5080 gnd.n1502 gnd.n1072 240.244
R5081 gnd.n1073 gnd.n1072 240.244
R5082 gnd.n1074 gnd.n1073 240.244
R5083 gnd.n5002 gnd.n1074 240.244
R5084 gnd.n5002 gnd.n1077 240.244
R5085 gnd.n1078 gnd.n1077 240.244
R5086 gnd.n1079 gnd.n1078 240.244
R5087 gnd.n1460 gnd.n1079 240.244
R5088 gnd.n1460 gnd.n1082 240.244
R5089 gnd.n1083 gnd.n1082 240.244
R5090 gnd.n1084 gnd.n1083 240.244
R5091 gnd.n5048 gnd.n1084 240.244
R5092 gnd.n5048 gnd.n1087 240.244
R5093 gnd.n1088 gnd.n1087 240.244
R5094 gnd.n1089 gnd.n1088 240.244
R5095 gnd.n5100 gnd.n1089 240.244
R5096 gnd.n5100 gnd.n1092 240.244
R5097 gnd.n1093 gnd.n1092 240.244
R5098 gnd.n1094 gnd.n1093 240.244
R5099 gnd.n1362 gnd.n1094 240.244
R5100 gnd.n1362 gnd.n1097 240.244
R5101 gnd.n1098 gnd.n1097 240.244
R5102 gnd.n1099 gnd.n1098 240.244
R5103 gnd.n5142 gnd.n1099 240.244
R5104 gnd.n5142 gnd.n1102 240.244
R5105 gnd.n1103 gnd.n1102 240.244
R5106 gnd.n5868 gnd.n1103 240.244
R5107 gnd.n4128 gnd.n4127 240.244
R5108 gnd.n4143 gnd.n4127 240.244
R5109 gnd.n4145 gnd.n4144 240.244
R5110 gnd.n4155 gnd.n4154 240.244
R5111 gnd.n4166 gnd.n4165 240.244
R5112 gnd.n4168 gnd.n4167 240.244
R5113 gnd.n4178 gnd.n4177 240.244
R5114 gnd.n4191 gnd.n4190 240.244
R5115 gnd.n4193 gnd.n4192 240.244
R5116 gnd.n2003 gnd.n2002 240.244
R5117 gnd.n4122 gnd.n2004 240.244
R5118 gnd.n2008 gnd.n2007 240.244
R5119 gnd.n2014 gnd.n2009 240.244
R5120 gnd.n2016 gnd.n2015 240.244
R5121 gnd.n4257 gnd.n4256 240.244
R5122 gnd.n4257 gnd.n1774 240.244
R5123 gnd.n4262 gnd.n1774 240.244
R5124 gnd.n4263 gnd.n4262 240.244
R5125 gnd.n4264 gnd.n4263 240.244
R5126 gnd.n4265 gnd.n4264 240.244
R5127 gnd.n4265 gnd.n1744 240.244
R5128 gnd.n4479 gnd.n1744 240.244
R5129 gnd.n4479 gnd.n1739 240.244
R5130 gnd.n4499 gnd.n1739 240.244
R5131 gnd.n4499 gnd.n1731 240.244
R5132 gnd.n4484 gnd.n1731 240.244
R5133 gnd.n4485 gnd.n4484 240.244
R5134 gnd.n4486 gnd.n4485 240.244
R5135 gnd.n4486 gnd.n1711 240.244
R5136 gnd.n1711 gnd.n1697 240.244
R5137 gnd.n4565 gnd.n1697 240.244
R5138 gnd.n4566 gnd.n4565 240.244
R5139 gnd.n4566 gnd.n1691 240.244
R5140 gnd.n4579 gnd.n1691 240.244
R5141 gnd.n4579 gnd.n1692 240.244
R5142 gnd.n4571 gnd.n1692 240.244
R5143 gnd.n4572 gnd.n4571 240.244
R5144 gnd.n4572 gnd.n1654 240.244
R5145 gnd.n4652 gnd.n1654 240.244
R5146 gnd.n4652 gnd.n1649 240.244
R5147 gnd.n4694 gnd.n1649 240.244
R5148 gnd.n4694 gnd.n1641 240.244
R5149 gnd.n4657 gnd.n1641 240.244
R5150 gnd.n4658 gnd.n4657 240.244
R5151 gnd.n4659 gnd.n4658 240.244
R5152 gnd.n4659 gnd.n1620 240.244
R5153 gnd.n1620 gnd.n1612 240.244
R5154 gnd.n4663 gnd.n1612 240.244
R5155 gnd.n4664 gnd.n4663 240.244
R5156 gnd.n4667 gnd.n4664 240.244
R5157 gnd.n4668 gnd.n4667 240.244
R5158 gnd.n4669 gnd.n4668 240.244
R5159 gnd.n4670 gnd.n4669 240.244
R5160 gnd.n4671 gnd.n4670 240.244
R5161 gnd.n4671 gnd.n1566 240.244
R5162 gnd.n4829 gnd.n1566 240.244
R5163 gnd.n4829 gnd.n1561 240.244
R5164 gnd.n4848 gnd.n1561 240.244
R5165 gnd.n4848 gnd.n1553 240.244
R5166 gnd.n4834 gnd.n1553 240.244
R5167 gnd.n4835 gnd.n4834 240.244
R5168 gnd.n4837 gnd.n4835 240.244
R5169 gnd.n4837 gnd.n1533 240.244
R5170 gnd.n1533 gnd.n1516 240.244
R5171 gnd.n4914 gnd.n1516 240.244
R5172 gnd.n4914 gnd.n1510 240.244
R5173 gnd.n4924 gnd.n1510 240.244
R5174 gnd.n4924 gnd.n1511 240.244
R5175 gnd.n4918 gnd.n1511 240.244
R5176 gnd.n4918 gnd.n1486 240.244
R5177 gnd.n4981 gnd.n1486 240.244
R5178 gnd.n4981 gnd.n1481 240.244
R5179 gnd.n5001 gnd.n1481 240.244
R5180 gnd.n5001 gnd.n1473 240.244
R5181 gnd.n4986 gnd.n1473 240.244
R5182 gnd.n4989 gnd.n4986 240.244
R5183 gnd.n4990 gnd.n4989 240.244
R5184 gnd.n4990 gnd.n1455 240.244
R5185 gnd.n1455 gnd.n1411 240.244
R5186 gnd.n5066 gnd.n1411 240.244
R5187 gnd.n5066 gnd.n1405 240.244
R5188 gnd.n5073 gnd.n1405 240.244
R5189 gnd.n5073 gnd.n1406 240.244
R5190 gnd.n1406 gnd.n1382 240.244
R5191 gnd.n5102 gnd.n1382 240.244
R5192 gnd.n5102 gnd.n1378 240.244
R5193 gnd.n5108 gnd.n1378 240.244
R5194 gnd.n5108 gnd.n1360 240.244
R5195 gnd.n5133 gnd.n1360 240.244
R5196 gnd.n5133 gnd.n1356 240.244
R5197 gnd.n5139 gnd.n1356 240.244
R5198 gnd.n5141 gnd.n5139 240.244
R5199 gnd.n5144 gnd.n5141 240.244
R5200 gnd.n5144 gnd.n1351 240.244
R5201 gnd.n5326 gnd.n1351 240.244
R5202 gnd.n5326 gnd.n1107 240.244
R5203 gnd.n5217 gnd.n5216 240.244
R5204 gnd.n5220 gnd.n5219 240.244
R5205 gnd.n5236 gnd.n5235 240.244
R5206 gnd.n5239 gnd.n5238 240.244
R5207 gnd.n5255 gnd.n5254 240.244
R5208 gnd.n5258 gnd.n5257 240.244
R5209 gnd.n5274 gnd.n5273 240.244
R5210 gnd.n5278 gnd.n5276 240.244
R5211 gnd.n5294 gnd.n5158 240.244
R5212 gnd.n5298 gnd.n5296 240.244
R5213 gnd.n5304 gnd.n5154 240.244
R5214 gnd.n5308 gnd.n5306 240.244
R5215 gnd.n5317 gnd.n5150 240.244
R5216 gnd.n5320 gnd.n5319 240.244
R5217 gnd.n1816 gnd.n1815 240.132
R5218 gnd.n5351 gnd.n5350 240.132
R5219 gnd.n6267 gnd.n655 225.874
R5220 gnd.n6268 gnd.n6267 225.874
R5221 gnd.n6269 gnd.n6268 225.874
R5222 gnd.n6269 gnd.n649 225.874
R5223 gnd.n6277 gnd.n649 225.874
R5224 gnd.n6278 gnd.n6277 225.874
R5225 gnd.n6279 gnd.n6278 225.874
R5226 gnd.n6279 gnd.n643 225.874
R5227 gnd.n6287 gnd.n643 225.874
R5228 gnd.n6288 gnd.n6287 225.874
R5229 gnd.n6289 gnd.n6288 225.874
R5230 gnd.n6289 gnd.n637 225.874
R5231 gnd.n6297 gnd.n637 225.874
R5232 gnd.n6298 gnd.n6297 225.874
R5233 gnd.n6299 gnd.n6298 225.874
R5234 gnd.n6299 gnd.n631 225.874
R5235 gnd.n6307 gnd.n631 225.874
R5236 gnd.n6308 gnd.n6307 225.874
R5237 gnd.n6309 gnd.n6308 225.874
R5238 gnd.n6309 gnd.n625 225.874
R5239 gnd.n6317 gnd.n625 225.874
R5240 gnd.n6318 gnd.n6317 225.874
R5241 gnd.n6319 gnd.n6318 225.874
R5242 gnd.n6319 gnd.n619 225.874
R5243 gnd.n6327 gnd.n619 225.874
R5244 gnd.n6328 gnd.n6327 225.874
R5245 gnd.n6329 gnd.n6328 225.874
R5246 gnd.n6329 gnd.n613 225.874
R5247 gnd.n6337 gnd.n613 225.874
R5248 gnd.n6338 gnd.n6337 225.874
R5249 gnd.n6339 gnd.n6338 225.874
R5250 gnd.n6339 gnd.n607 225.874
R5251 gnd.n6347 gnd.n607 225.874
R5252 gnd.n6348 gnd.n6347 225.874
R5253 gnd.n6349 gnd.n6348 225.874
R5254 gnd.n6349 gnd.n601 225.874
R5255 gnd.n6357 gnd.n601 225.874
R5256 gnd.n6358 gnd.n6357 225.874
R5257 gnd.n6359 gnd.n6358 225.874
R5258 gnd.n6359 gnd.n595 225.874
R5259 gnd.n6367 gnd.n595 225.874
R5260 gnd.n6368 gnd.n6367 225.874
R5261 gnd.n6369 gnd.n6368 225.874
R5262 gnd.n6369 gnd.n589 225.874
R5263 gnd.n6377 gnd.n589 225.874
R5264 gnd.n6378 gnd.n6377 225.874
R5265 gnd.n6379 gnd.n6378 225.874
R5266 gnd.n6379 gnd.n583 225.874
R5267 gnd.n6387 gnd.n583 225.874
R5268 gnd.n6388 gnd.n6387 225.874
R5269 gnd.n6389 gnd.n6388 225.874
R5270 gnd.n6389 gnd.n577 225.874
R5271 gnd.n6397 gnd.n577 225.874
R5272 gnd.n6398 gnd.n6397 225.874
R5273 gnd.n6399 gnd.n6398 225.874
R5274 gnd.n6399 gnd.n571 225.874
R5275 gnd.n6407 gnd.n571 225.874
R5276 gnd.n6408 gnd.n6407 225.874
R5277 gnd.n6409 gnd.n6408 225.874
R5278 gnd.n6409 gnd.n565 225.874
R5279 gnd.n6417 gnd.n565 225.874
R5280 gnd.n6418 gnd.n6417 225.874
R5281 gnd.n6419 gnd.n6418 225.874
R5282 gnd.n6419 gnd.n559 225.874
R5283 gnd.n6427 gnd.n559 225.874
R5284 gnd.n6428 gnd.n6427 225.874
R5285 gnd.n6429 gnd.n6428 225.874
R5286 gnd.n6429 gnd.n553 225.874
R5287 gnd.n6437 gnd.n553 225.874
R5288 gnd.n6438 gnd.n6437 225.874
R5289 gnd.n6439 gnd.n6438 225.874
R5290 gnd.n6439 gnd.n547 225.874
R5291 gnd.n6447 gnd.n547 225.874
R5292 gnd.n6448 gnd.n6447 225.874
R5293 gnd.n6449 gnd.n6448 225.874
R5294 gnd.n6449 gnd.n541 225.874
R5295 gnd.n6457 gnd.n541 225.874
R5296 gnd.n6458 gnd.n6457 225.874
R5297 gnd.n6459 gnd.n6458 225.874
R5298 gnd.n6459 gnd.n535 225.874
R5299 gnd.n6467 gnd.n535 225.874
R5300 gnd.n6468 gnd.n6467 225.874
R5301 gnd.n6469 gnd.n6468 225.874
R5302 gnd.n6469 gnd.n529 225.874
R5303 gnd.n6477 gnd.n529 225.874
R5304 gnd.n6478 gnd.n6477 225.874
R5305 gnd.n6479 gnd.n6478 225.874
R5306 gnd.n6479 gnd.n523 225.874
R5307 gnd.n6487 gnd.n523 225.874
R5308 gnd.n6488 gnd.n6487 225.874
R5309 gnd.n6489 gnd.n6488 225.874
R5310 gnd.n6489 gnd.n517 225.874
R5311 gnd.n6497 gnd.n517 225.874
R5312 gnd.n6498 gnd.n6497 225.874
R5313 gnd.n6499 gnd.n6498 225.874
R5314 gnd.n6499 gnd.n511 225.874
R5315 gnd.n6507 gnd.n511 225.874
R5316 gnd.n6508 gnd.n6507 225.874
R5317 gnd.n6509 gnd.n6508 225.874
R5318 gnd.n6509 gnd.n505 225.874
R5319 gnd.n6517 gnd.n505 225.874
R5320 gnd.n6518 gnd.n6517 225.874
R5321 gnd.n6519 gnd.n6518 225.874
R5322 gnd.n6519 gnd.n499 225.874
R5323 gnd.n6527 gnd.n499 225.874
R5324 gnd.n6528 gnd.n6527 225.874
R5325 gnd.n6529 gnd.n6528 225.874
R5326 gnd.n6529 gnd.n493 225.874
R5327 gnd.n6537 gnd.n493 225.874
R5328 gnd.n6538 gnd.n6537 225.874
R5329 gnd.n6539 gnd.n6538 225.874
R5330 gnd.n6539 gnd.n487 225.874
R5331 gnd.n6547 gnd.n487 225.874
R5332 gnd.n6548 gnd.n6547 225.874
R5333 gnd.n6549 gnd.n6548 225.874
R5334 gnd.n6549 gnd.n481 225.874
R5335 gnd.n6557 gnd.n481 225.874
R5336 gnd.n6558 gnd.n6557 225.874
R5337 gnd.n6559 gnd.n6558 225.874
R5338 gnd.n6559 gnd.n475 225.874
R5339 gnd.n6567 gnd.n475 225.874
R5340 gnd.n6568 gnd.n6567 225.874
R5341 gnd.n6569 gnd.n6568 225.874
R5342 gnd.n6569 gnd.n469 225.874
R5343 gnd.n6577 gnd.n469 225.874
R5344 gnd.n6578 gnd.n6577 225.874
R5345 gnd.n6579 gnd.n6578 225.874
R5346 gnd.n6579 gnd.n463 225.874
R5347 gnd.n6587 gnd.n463 225.874
R5348 gnd.n6588 gnd.n6587 225.874
R5349 gnd.n6589 gnd.n6588 225.874
R5350 gnd.n6589 gnd.n457 225.874
R5351 gnd.n6597 gnd.n457 225.874
R5352 gnd.n6598 gnd.n6597 225.874
R5353 gnd.n6599 gnd.n6598 225.874
R5354 gnd.n6599 gnd.n451 225.874
R5355 gnd.n6607 gnd.n451 225.874
R5356 gnd.n6608 gnd.n6607 225.874
R5357 gnd.n6609 gnd.n6608 225.874
R5358 gnd.n6609 gnd.n445 225.874
R5359 gnd.n6617 gnd.n445 225.874
R5360 gnd.n6618 gnd.n6617 225.874
R5361 gnd.n6619 gnd.n6618 225.874
R5362 gnd.n6619 gnd.n439 225.874
R5363 gnd.n6627 gnd.n439 225.874
R5364 gnd.n6628 gnd.n6627 225.874
R5365 gnd.n6629 gnd.n6628 225.874
R5366 gnd.n6629 gnd.n433 225.874
R5367 gnd.n6637 gnd.n433 225.874
R5368 gnd.n6638 gnd.n6637 225.874
R5369 gnd.n6639 gnd.n6638 225.874
R5370 gnd.n6639 gnd.n427 225.874
R5371 gnd.n6647 gnd.n427 225.874
R5372 gnd.n6648 gnd.n6647 225.874
R5373 gnd.n6649 gnd.n6648 225.874
R5374 gnd.n6649 gnd.n421 225.874
R5375 gnd.n6657 gnd.n421 225.874
R5376 gnd.n6658 gnd.n6657 225.874
R5377 gnd.n6659 gnd.n6658 225.874
R5378 gnd.n6659 gnd.n415 225.874
R5379 gnd.n6667 gnd.n415 225.874
R5380 gnd.n6668 gnd.n6667 225.874
R5381 gnd.n6669 gnd.n6668 225.874
R5382 gnd.n6669 gnd.n409 225.874
R5383 gnd.n6677 gnd.n409 225.874
R5384 gnd.n6678 gnd.n6677 225.874
R5385 gnd.n6679 gnd.n6678 225.874
R5386 gnd.n2704 gnd.t124 224.174
R5387 gnd.n2226 gnd.t57 224.174
R5388 gnd.n6891 gnd.n83 215.659
R5389 gnd.n6687 gnd.n403 206.476
R5390 gnd.n6688 gnd.n6687 206.476
R5391 gnd.n6689 gnd.n6688 206.476
R5392 gnd.n6689 gnd.n397 206.476
R5393 gnd.n6697 gnd.n397 206.476
R5394 gnd.n6698 gnd.n6697 206.476
R5395 gnd.n6699 gnd.n6698 206.476
R5396 gnd.n6699 gnd.n391 206.476
R5397 gnd.n6707 gnd.n391 206.476
R5398 gnd.n6708 gnd.n6707 206.476
R5399 gnd.n6709 gnd.n6708 206.476
R5400 gnd.n6709 gnd.n385 206.476
R5401 gnd.n6717 gnd.n385 206.476
R5402 gnd.n6718 gnd.n6717 206.476
R5403 gnd.n6719 gnd.n6718 206.476
R5404 gnd.n6719 gnd.n379 206.476
R5405 gnd.n6727 gnd.n379 206.476
R5406 gnd.n6728 gnd.n6727 206.476
R5407 gnd.n6729 gnd.n6728 206.476
R5408 gnd.n6729 gnd.n373 206.476
R5409 gnd.n6737 gnd.n373 206.476
R5410 gnd.n6738 gnd.n6737 206.476
R5411 gnd.n6739 gnd.n6738 206.476
R5412 gnd.n6739 gnd.n367 206.476
R5413 gnd.n6747 gnd.n367 206.476
R5414 gnd.n6748 gnd.n6747 206.476
R5415 gnd.n6749 gnd.n6748 206.476
R5416 gnd.n6749 gnd.n361 206.476
R5417 gnd.n6757 gnd.n361 206.476
R5418 gnd.n6758 gnd.n6757 206.476
R5419 gnd.n6759 gnd.n6758 206.476
R5420 gnd.n6759 gnd.n355 206.476
R5421 gnd.n6767 gnd.n355 206.476
R5422 gnd.n6768 gnd.n6767 206.476
R5423 gnd.n6769 gnd.n6768 206.476
R5424 gnd.n6769 gnd.n349 206.476
R5425 gnd.n6777 gnd.n349 206.476
R5426 gnd.n6778 gnd.n6777 206.476
R5427 gnd.n6779 gnd.n6778 206.476
R5428 gnd.n6779 gnd.n343 206.476
R5429 gnd.n6787 gnd.n343 206.476
R5430 gnd.n6788 gnd.n6787 206.476
R5431 gnd.n6789 gnd.n6788 206.476
R5432 gnd.n6789 gnd.n337 206.476
R5433 gnd.n6797 gnd.n337 206.476
R5434 gnd.n6798 gnd.n6797 206.476
R5435 gnd.n6799 gnd.n6798 206.476
R5436 gnd.n6799 gnd.n331 206.476
R5437 gnd.n6807 gnd.n331 206.476
R5438 gnd.n6808 gnd.n6807 206.476
R5439 gnd.n6809 gnd.n6808 206.476
R5440 gnd.n6809 gnd.n325 206.476
R5441 gnd.n6817 gnd.n325 206.476
R5442 gnd.n6818 gnd.n6817 206.476
R5443 gnd.n6819 gnd.n6818 206.476
R5444 gnd.n6819 gnd.n319 206.476
R5445 gnd.n6827 gnd.n319 206.476
R5446 gnd.n6828 gnd.n6827 206.476
R5447 gnd.n6829 gnd.n6828 206.476
R5448 gnd.n6829 gnd.n313 206.476
R5449 gnd.n6837 gnd.n313 206.476
R5450 gnd.n6838 gnd.n6837 206.476
R5451 gnd.n6839 gnd.n6838 206.476
R5452 gnd.n6839 gnd.n307 206.476
R5453 gnd.n6847 gnd.n307 206.476
R5454 gnd.n6848 gnd.n6847 206.476
R5455 gnd.n6849 gnd.n6848 206.476
R5456 gnd.n6849 gnd.n301 206.476
R5457 gnd.n6857 gnd.n301 206.476
R5458 gnd.n6858 gnd.n6857 206.476
R5459 gnd.n6859 gnd.n6858 206.476
R5460 gnd.n6859 gnd.n295 206.476
R5461 gnd.n6867 gnd.n295 206.476
R5462 gnd.n6868 gnd.n6867 206.476
R5463 gnd.n6869 gnd.n6868 206.476
R5464 gnd.n6869 gnd.n289 206.476
R5465 gnd.n6877 gnd.n289 206.476
R5466 gnd.n6878 gnd.n6877 206.476
R5467 gnd.n6879 gnd.n6878 206.476
R5468 gnd.n6879 gnd.n283 206.476
R5469 gnd.n6889 gnd.n283 206.476
R5470 gnd.n6890 gnd.n6889 206.476
R5471 gnd.n6891 gnd.n6890 206.476
R5472 gnd.n5551 gnd.n5550 199.319
R5473 gnd.n5551 gnd.n5497 199.319
R5474 gnd.n1908 gnd.n1902 199.319
R5475 gnd.n1907 gnd.n1902 199.319
R5476 gnd.n1817 gnd.n1814 186.49
R5477 gnd.n5352 gnd.n5349 186.49
R5478 gnd.n3480 gnd.n3479 185
R5479 gnd.n3478 gnd.n3477 185
R5480 gnd.n3457 gnd.n3456 185
R5481 gnd.n3472 gnd.n3471 185
R5482 gnd.n3470 gnd.n3469 185
R5483 gnd.n3461 gnd.n3460 185
R5484 gnd.n3464 gnd.n3463 185
R5485 gnd.n3448 gnd.n3447 185
R5486 gnd.n3446 gnd.n3445 185
R5487 gnd.n3425 gnd.n3424 185
R5488 gnd.n3440 gnd.n3439 185
R5489 gnd.n3438 gnd.n3437 185
R5490 gnd.n3429 gnd.n3428 185
R5491 gnd.n3432 gnd.n3431 185
R5492 gnd.n3416 gnd.n3415 185
R5493 gnd.n3414 gnd.n3413 185
R5494 gnd.n3393 gnd.n3392 185
R5495 gnd.n3408 gnd.n3407 185
R5496 gnd.n3406 gnd.n3405 185
R5497 gnd.n3397 gnd.n3396 185
R5498 gnd.n3400 gnd.n3399 185
R5499 gnd.n3385 gnd.n3384 185
R5500 gnd.n3383 gnd.n3382 185
R5501 gnd.n3362 gnd.n3361 185
R5502 gnd.n3377 gnd.n3376 185
R5503 gnd.n3375 gnd.n3374 185
R5504 gnd.n3366 gnd.n3365 185
R5505 gnd.n3369 gnd.n3368 185
R5506 gnd.n3353 gnd.n3352 185
R5507 gnd.n3351 gnd.n3350 185
R5508 gnd.n3330 gnd.n3329 185
R5509 gnd.n3345 gnd.n3344 185
R5510 gnd.n3343 gnd.n3342 185
R5511 gnd.n3334 gnd.n3333 185
R5512 gnd.n3337 gnd.n3336 185
R5513 gnd.n3321 gnd.n3320 185
R5514 gnd.n3319 gnd.n3318 185
R5515 gnd.n3298 gnd.n3297 185
R5516 gnd.n3313 gnd.n3312 185
R5517 gnd.n3311 gnd.n3310 185
R5518 gnd.n3302 gnd.n3301 185
R5519 gnd.n3305 gnd.n3304 185
R5520 gnd.n3289 gnd.n3288 185
R5521 gnd.n3287 gnd.n3286 185
R5522 gnd.n3266 gnd.n3265 185
R5523 gnd.n3281 gnd.n3280 185
R5524 gnd.n3279 gnd.n3278 185
R5525 gnd.n3270 gnd.n3269 185
R5526 gnd.n3273 gnd.n3272 185
R5527 gnd.n3258 gnd.n3257 185
R5528 gnd.n3256 gnd.n3255 185
R5529 gnd.n3235 gnd.n3234 185
R5530 gnd.n3250 gnd.n3249 185
R5531 gnd.n3248 gnd.n3247 185
R5532 gnd.n3239 gnd.n3238 185
R5533 gnd.n3242 gnd.n3241 185
R5534 gnd.n2705 gnd.t123 178.987
R5535 gnd.n2227 gnd.t58 178.987
R5536 gnd.n1 gnd.t167 170.774
R5537 gnd.n7 gnd.t3 170.103
R5538 gnd.n6 gnd.t134 170.103
R5539 gnd.n5 gnd.t201 170.103
R5540 gnd.n4 gnd.t289 170.103
R5541 gnd.n3 gnd.t236 170.103
R5542 gnd.n2 gnd.t218 170.103
R5543 gnd.n1 gnd.t192 170.103
R5544 gnd.n5420 gnd.n5419 163.367
R5545 gnd.n5416 gnd.n5415 163.367
R5546 gnd.n5412 gnd.n5411 163.367
R5547 gnd.n5408 gnd.n5407 163.367
R5548 gnd.n5404 gnd.n5403 163.367
R5549 gnd.n5400 gnd.n5399 163.367
R5550 gnd.n5396 gnd.n5395 163.367
R5551 gnd.n5392 gnd.n5391 163.367
R5552 gnd.n5388 gnd.n5387 163.367
R5553 gnd.n5384 gnd.n5383 163.367
R5554 gnd.n5380 gnd.n5379 163.367
R5555 gnd.n5376 gnd.n5375 163.367
R5556 gnd.n5372 gnd.n5371 163.367
R5557 gnd.n5368 gnd.n5367 163.367
R5558 gnd.n5363 gnd.n5362 163.367
R5559 gnd.n5495 gnd.n1295 163.367
R5560 gnd.n5492 gnd.n5491 163.367
R5561 gnd.n5489 gnd.n1328 163.367
R5562 gnd.n5484 gnd.n5483 163.367
R5563 gnd.n5480 gnd.n5479 163.367
R5564 gnd.n5476 gnd.n5475 163.367
R5565 gnd.n5472 gnd.n5471 163.367
R5566 gnd.n5468 gnd.n5467 163.367
R5567 gnd.n5464 gnd.n5463 163.367
R5568 gnd.n5460 gnd.n5459 163.367
R5569 gnd.n5456 gnd.n5455 163.367
R5570 gnd.n5452 gnd.n5451 163.367
R5571 gnd.n5448 gnd.n5447 163.367
R5572 gnd.n5444 gnd.n5443 163.367
R5573 gnd.n5440 gnd.n5439 163.367
R5574 gnd.n5436 gnd.n5435 163.367
R5575 gnd.n5432 gnd.n5431 163.367
R5576 gnd.n4424 gnd.n1765 163.367
R5577 gnd.n4449 gnd.n1765 163.367
R5578 gnd.n4449 gnd.n1759 163.367
R5579 gnd.n4445 gnd.n1759 163.367
R5580 gnd.n4445 gnd.n1751 163.367
R5581 gnd.n4440 gnd.n1751 163.367
R5582 gnd.n4440 gnd.n1746 163.367
R5583 gnd.n4437 gnd.n1746 163.367
R5584 gnd.n4437 gnd.n1738 163.367
R5585 gnd.n4432 gnd.n1738 163.367
R5586 gnd.n4432 gnd.n1732 163.367
R5587 gnd.n4429 gnd.n1732 163.367
R5588 gnd.n4429 gnd.n1722 163.367
R5589 gnd.n1722 gnd.n1714 163.367
R5590 gnd.n4527 gnd.n1714 163.367
R5591 gnd.n4527 gnd.n1712 163.367
R5592 gnd.n4542 gnd.n1712 163.367
R5593 gnd.n4542 gnd.n1703 163.367
R5594 gnd.n4538 gnd.n1703 163.367
R5595 gnd.n4538 gnd.n1698 163.367
R5596 gnd.n4535 gnd.n1698 163.367
R5597 gnd.n4535 gnd.n1685 163.367
R5598 gnd.n4531 gnd.n1685 163.367
R5599 gnd.n4531 gnd.n1678 163.367
R5600 gnd.n4598 gnd.n1678 163.367
R5601 gnd.n4598 gnd.n1676 163.367
R5602 gnd.n4623 gnd.n1676 163.367
R5603 gnd.n4623 gnd.n1669 163.367
R5604 gnd.n4619 gnd.n1669 163.367
R5605 gnd.n4619 gnd.n1660 163.367
R5606 gnd.n4614 gnd.n1660 163.367
R5607 gnd.n4614 gnd.n1655 163.367
R5608 gnd.n4611 gnd.n1655 163.367
R5609 gnd.n4611 gnd.n1648 163.367
R5610 gnd.n4606 gnd.n1648 163.367
R5611 gnd.n4606 gnd.n1642 163.367
R5612 gnd.n4603 gnd.n1642 163.367
R5613 gnd.n4603 gnd.n1632 163.367
R5614 gnd.n1632 gnd.n1623 163.367
R5615 gnd.n4722 gnd.n1623 163.367
R5616 gnd.n4722 gnd.n1621 163.367
R5617 gnd.n4729 gnd.n1621 163.367
R5618 gnd.n4729 gnd.n1611 163.367
R5619 gnd.n4725 gnd.n1611 163.367
R5620 gnd.n4725 gnd.n1606 163.367
R5621 gnd.n4751 gnd.n1606 163.367
R5622 gnd.n4751 gnd.n1600 163.367
R5623 gnd.n4755 gnd.n1600 163.367
R5624 gnd.n4755 gnd.n1591 163.367
R5625 gnd.n4775 gnd.n1591 163.367
R5626 gnd.n4775 gnd.n1589 163.367
R5627 gnd.n4800 gnd.n1589 163.367
R5628 gnd.n4800 gnd.n1583 163.367
R5629 gnd.n4796 gnd.n1583 163.367
R5630 gnd.n4796 gnd.n1574 163.367
R5631 gnd.n4792 gnd.n1574 163.367
R5632 gnd.n4792 gnd.n1568 163.367
R5633 gnd.n4789 gnd.n1568 163.367
R5634 gnd.n4789 gnd.n1560 163.367
R5635 gnd.n4783 gnd.n1560 163.367
R5636 gnd.n4783 gnd.n1554 163.367
R5637 gnd.n4780 gnd.n1554 163.367
R5638 gnd.n4780 gnd.n1543 163.367
R5639 gnd.n1543 gnd.n1536 163.367
R5640 gnd.n4875 gnd.n1536 163.367
R5641 gnd.n4875 gnd.n1534 163.367
R5642 gnd.n4883 gnd.n1534 163.367
R5643 gnd.n4883 gnd.n1524 163.367
R5644 gnd.n4879 gnd.n1524 163.367
R5645 gnd.n4879 gnd.n1517 163.367
R5646 gnd.n1517 gnd.n1509 163.367
R5647 gnd.n4927 gnd.n1509 163.367
R5648 gnd.n4927 gnd.n1507 163.367
R5649 gnd.n4951 gnd.n1507 163.367
R5650 gnd.n4951 gnd.n1501 163.367
R5651 gnd.n4947 gnd.n1501 163.367
R5652 gnd.n4947 gnd.n1493 163.367
R5653 gnd.n4942 gnd.n1493 163.367
R5654 gnd.n4942 gnd.n1488 163.367
R5655 gnd.n4939 gnd.n1488 163.367
R5656 gnd.n4939 gnd.n1480 163.367
R5657 gnd.n4935 gnd.n1480 163.367
R5658 gnd.n4935 gnd.n1474 163.367
R5659 gnd.n4932 gnd.n1474 163.367
R5660 gnd.n4932 gnd.n1466 163.367
R5661 gnd.n1466 gnd.n1458 163.367
R5662 gnd.n5031 gnd.n1458 163.367
R5663 gnd.n5031 gnd.n1456 163.367
R5664 gnd.n5035 gnd.n1456 163.367
R5665 gnd.n5035 gnd.n1418 163.367
R5666 gnd.n5055 gnd.n1418 163.367
R5667 gnd.n5055 gnd.n1413 163.367
R5668 gnd.n5051 gnd.n1413 163.367
R5669 gnd.n5051 gnd.n1404 163.367
R5670 gnd.n1446 gnd.n1404 163.367
R5671 gnd.n1446 gnd.n1398 163.367
R5672 gnd.n1443 gnd.n1398 163.367
R5673 gnd.n1443 gnd.n1391 163.367
R5674 gnd.n1438 gnd.n1391 163.367
R5675 gnd.n1438 gnd.n1384 163.367
R5676 gnd.n1435 gnd.n1384 163.367
R5677 gnd.n1435 gnd.n1377 163.367
R5678 gnd.n1377 gnd.n1368 163.367
R5679 gnd.n1369 gnd.n1368 163.367
R5680 gnd.n1369 gnd.n1361 163.367
R5681 gnd.n1429 gnd.n1361 163.367
R5682 gnd.n1429 gnd.n1423 163.367
R5683 gnd.n1423 gnd.n1339 163.367
R5684 gnd.n1339 gnd.n1332 163.367
R5685 gnd.n5427 gnd.n1332 163.367
R5686 gnd.n1809 gnd.n1808 163.367
R5687 gnd.n4405 gnd.n1808 163.367
R5688 gnd.n4403 gnd.n4402 163.367
R5689 gnd.n4399 gnd.n4398 163.367
R5690 gnd.n4395 gnd.n4394 163.367
R5691 gnd.n4391 gnd.n4390 163.367
R5692 gnd.n4387 gnd.n4386 163.367
R5693 gnd.n4383 gnd.n4382 163.367
R5694 gnd.n4379 gnd.n4378 163.367
R5695 gnd.n4375 gnd.n4374 163.367
R5696 gnd.n4371 gnd.n4370 163.367
R5697 gnd.n4367 gnd.n4366 163.367
R5698 gnd.n4363 gnd.n4362 163.367
R5699 gnd.n4359 gnd.n4358 163.367
R5700 gnd.n4355 gnd.n4354 163.367
R5701 gnd.n4351 gnd.n4350 163.367
R5702 gnd.n4347 gnd.n4346 163.367
R5703 gnd.n1895 gnd.n1894 163.367
R5704 gnd.n1890 gnd.n1889 163.367
R5705 gnd.n1886 gnd.n1885 163.367
R5706 gnd.n1882 gnd.n1881 163.367
R5707 gnd.n1878 gnd.n1877 163.367
R5708 gnd.n1874 gnd.n1873 163.367
R5709 gnd.n1870 gnd.n1869 163.367
R5710 gnd.n1866 gnd.n1865 163.367
R5711 gnd.n1862 gnd.n1861 163.367
R5712 gnd.n1858 gnd.n1857 163.367
R5713 gnd.n1854 gnd.n1853 163.367
R5714 gnd.n1850 gnd.n1849 163.367
R5715 gnd.n1846 gnd.n1845 163.367
R5716 gnd.n1842 gnd.n1841 163.367
R5717 gnd.n1838 gnd.n1837 163.367
R5718 gnd.n4453 gnd.n1763 163.367
R5719 gnd.n4453 gnd.n1761 163.367
R5720 gnd.n4457 gnd.n1761 163.367
R5721 gnd.n4457 gnd.n1750 163.367
R5722 gnd.n4472 gnd.n1750 163.367
R5723 gnd.n4472 gnd.n1748 163.367
R5724 gnd.n4476 gnd.n1748 163.367
R5725 gnd.n4476 gnd.n1736 163.367
R5726 gnd.n4502 gnd.n1736 163.367
R5727 gnd.n4502 gnd.n1734 163.367
R5728 gnd.n4506 gnd.n1734 163.367
R5729 gnd.n4506 gnd.n1720 163.367
R5730 gnd.n4520 gnd.n1720 163.367
R5731 gnd.n4520 gnd.n1717 163.367
R5732 gnd.n4525 gnd.n1717 163.367
R5733 gnd.n4525 gnd.n1718 163.367
R5734 gnd.n1718 gnd.n1702 163.367
R5735 gnd.n4558 gnd.n1702 163.367
R5736 gnd.n4558 gnd.n1700 163.367
R5737 gnd.n4562 gnd.n1700 163.367
R5738 gnd.n4562 gnd.n1687 163.367
R5739 gnd.n4586 gnd.n1687 163.367
R5740 gnd.n4586 gnd.n1688 163.367
R5741 gnd.n4582 gnd.n1688 163.367
R5742 gnd.n4582 gnd.n1674 163.367
R5743 gnd.n4627 gnd.n1674 163.367
R5744 gnd.n4627 gnd.n1672 163.367
R5745 gnd.n4631 gnd.n1672 163.367
R5746 gnd.n4631 gnd.n1659 163.367
R5747 gnd.n4645 gnd.n1659 163.367
R5748 gnd.n4645 gnd.n1657 163.367
R5749 gnd.n4649 gnd.n1657 163.367
R5750 gnd.n4649 gnd.n1646 163.367
R5751 gnd.n4698 gnd.n1646 163.367
R5752 gnd.n4698 gnd.n1644 163.367
R5753 gnd.n4702 gnd.n1644 163.367
R5754 gnd.n4702 gnd.n1630 163.367
R5755 gnd.n4715 gnd.n1630 163.367
R5756 gnd.n4715 gnd.n1627 163.367
R5757 gnd.n4720 gnd.n1627 163.367
R5758 gnd.n4720 gnd.n1628 163.367
R5759 gnd.n1628 gnd.n1609 163.367
R5760 gnd.n4743 gnd.n1609 163.367
R5761 gnd.n4743 gnd.n1607 163.367
R5762 gnd.n4747 gnd.n1607 163.367
R5763 gnd.n4747 gnd.n1602 163.367
R5764 gnd.n4763 gnd.n1602 163.367
R5765 gnd.n4763 gnd.n1603 163.367
R5766 gnd.n4759 gnd.n1603 163.367
R5767 gnd.n4759 gnd.n1587 163.367
R5768 gnd.n4804 gnd.n1587 163.367
R5769 gnd.n4804 gnd.n1585 163.367
R5770 gnd.n4808 gnd.n1585 163.367
R5771 gnd.n4808 gnd.n1572 163.367
R5772 gnd.n4822 gnd.n1572 163.367
R5773 gnd.n4822 gnd.n1570 163.367
R5774 gnd.n4826 gnd.n1570 163.367
R5775 gnd.n4826 gnd.n1558 163.367
R5776 gnd.n4851 gnd.n1558 163.367
R5777 gnd.n4851 gnd.n1556 163.367
R5778 gnd.n4855 gnd.n1556 163.367
R5779 gnd.n4855 gnd.n1541 163.367
R5780 gnd.n4868 gnd.n1541 163.367
R5781 gnd.n4868 gnd.n1538 163.367
R5782 gnd.n4873 gnd.n1538 163.367
R5783 gnd.n4873 gnd.n1539 163.367
R5784 gnd.n1539 gnd.n1522 163.367
R5785 gnd.n4905 gnd.n1522 163.367
R5786 gnd.n4905 gnd.n1519 163.367
R5787 gnd.n4910 gnd.n1519 163.367
R5788 gnd.n4910 gnd.n1520 163.367
R5789 gnd.n1520 gnd.n1506 163.367
R5790 gnd.n4955 gnd.n1506 163.367
R5791 gnd.n4955 gnd.n1504 163.367
R5792 gnd.n4959 gnd.n1504 163.367
R5793 gnd.n4959 gnd.n1492 163.367
R5794 gnd.n4974 gnd.n1492 163.367
R5795 gnd.n4974 gnd.n1490 163.367
R5796 gnd.n4978 gnd.n1490 163.367
R5797 gnd.n4978 gnd.n1478 163.367
R5798 gnd.n5005 gnd.n1478 163.367
R5799 gnd.n5005 gnd.n1476 163.367
R5800 gnd.n5009 gnd.n1476 163.367
R5801 gnd.n5009 gnd.n1464 163.367
R5802 gnd.n5024 gnd.n1464 163.367
R5803 gnd.n5024 gnd.n1461 163.367
R5804 gnd.n5029 gnd.n1461 163.367
R5805 gnd.n5029 gnd.n1462 163.367
R5806 gnd.n1462 gnd.n1416 163.367
R5807 gnd.n5059 gnd.n1416 163.367
R5808 gnd.n5059 gnd.n1414 163.367
R5809 gnd.n5063 gnd.n1414 163.367
R5810 gnd.n5063 gnd.n1402 163.367
R5811 gnd.n5076 gnd.n1402 163.367
R5812 gnd.n5076 gnd.n1400 163.367
R5813 gnd.n5080 gnd.n1400 163.367
R5814 gnd.n5080 gnd.n1389 163.367
R5815 gnd.n5092 gnd.n1389 163.367
R5816 gnd.n5092 gnd.n1386 163.367
R5817 gnd.n5097 gnd.n1386 163.367
R5818 gnd.n5097 gnd.n1387 163.367
R5819 gnd.n1387 gnd.n1366 163.367
R5820 gnd.n5126 gnd.n1366 163.367
R5821 gnd.n5126 gnd.n1363 163.367
R5822 gnd.n5131 gnd.n1363 163.367
R5823 gnd.n5131 gnd.n1364 163.367
R5824 gnd.n1364 gnd.n1337 163.367
R5825 gnd.n5337 gnd.n1337 163.367
R5826 gnd.n5337 gnd.n1334 163.367
R5827 gnd.n5425 gnd.n1334 163.367
R5828 gnd.n5358 gnd.n5357 156.462
R5829 gnd.n3420 gnd.n3388 153.042
R5830 gnd.n3484 gnd.n3483 152.079
R5831 gnd.n3452 gnd.n3451 152.079
R5832 gnd.n3420 gnd.n3419 152.079
R5833 gnd.n1822 gnd.n1821 152
R5834 gnd.n1823 gnd.n1812 152
R5835 gnd.n1825 gnd.n1824 152
R5836 gnd.n1827 gnd.n1810 152
R5837 gnd.n1829 gnd.n1828 152
R5838 gnd.n5356 gnd.n5340 152
R5839 gnd.n5348 gnd.n5341 152
R5840 gnd.n5347 gnd.n5346 152
R5841 gnd.n5345 gnd.n5342 152
R5842 gnd.n5343 gnd.t102 150.546
R5843 gnd.t176 gnd.n3462 147.661
R5844 gnd.t145 gnd.n3430 147.661
R5845 gnd.t230 gnd.n3398 147.661
R5846 gnd.t155 gnd.n3367 147.661
R5847 gnd.t199 gnd.n3335 147.661
R5848 gnd.t277 gnd.n3303 147.661
R5849 gnd.t185 gnd.n3271 147.661
R5850 gnd.t287 gnd.n3240 147.661
R5851 gnd.n5494 gnd.n1294 143.351
R5852 gnd.n4345 gnd.n1789 143.351
R5853 gnd.n4345 gnd.n1790 143.351
R5854 gnd.n1819 gnd.t31 130.484
R5855 gnd.n1828 gnd.t96 126.766
R5856 gnd.n1826 gnd.t24 126.766
R5857 gnd.n1812 gnd.t52 126.766
R5858 gnd.n1820 gnd.t115 126.766
R5859 gnd.n5344 gnd.t89 126.766
R5860 gnd.n5346 gnd.t17 126.766
R5861 gnd.n5355 gnd.t73 126.766
R5862 gnd.n5357 gnd.t38 126.766
R5863 gnd.n3479 gnd.n3478 104.615
R5864 gnd.n3478 gnd.n3456 104.615
R5865 gnd.n3471 gnd.n3456 104.615
R5866 gnd.n3471 gnd.n3470 104.615
R5867 gnd.n3470 gnd.n3460 104.615
R5868 gnd.n3463 gnd.n3460 104.615
R5869 gnd.n3447 gnd.n3446 104.615
R5870 gnd.n3446 gnd.n3424 104.615
R5871 gnd.n3439 gnd.n3424 104.615
R5872 gnd.n3439 gnd.n3438 104.615
R5873 gnd.n3438 gnd.n3428 104.615
R5874 gnd.n3431 gnd.n3428 104.615
R5875 gnd.n3415 gnd.n3414 104.615
R5876 gnd.n3414 gnd.n3392 104.615
R5877 gnd.n3407 gnd.n3392 104.615
R5878 gnd.n3407 gnd.n3406 104.615
R5879 gnd.n3406 gnd.n3396 104.615
R5880 gnd.n3399 gnd.n3396 104.615
R5881 gnd.n3384 gnd.n3383 104.615
R5882 gnd.n3383 gnd.n3361 104.615
R5883 gnd.n3376 gnd.n3361 104.615
R5884 gnd.n3376 gnd.n3375 104.615
R5885 gnd.n3375 gnd.n3365 104.615
R5886 gnd.n3368 gnd.n3365 104.615
R5887 gnd.n3352 gnd.n3351 104.615
R5888 gnd.n3351 gnd.n3329 104.615
R5889 gnd.n3344 gnd.n3329 104.615
R5890 gnd.n3344 gnd.n3343 104.615
R5891 gnd.n3343 gnd.n3333 104.615
R5892 gnd.n3336 gnd.n3333 104.615
R5893 gnd.n3320 gnd.n3319 104.615
R5894 gnd.n3319 gnd.n3297 104.615
R5895 gnd.n3312 gnd.n3297 104.615
R5896 gnd.n3312 gnd.n3311 104.615
R5897 gnd.n3311 gnd.n3301 104.615
R5898 gnd.n3304 gnd.n3301 104.615
R5899 gnd.n3288 gnd.n3287 104.615
R5900 gnd.n3287 gnd.n3265 104.615
R5901 gnd.n3280 gnd.n3265 104.615
R5902 gnd.n3280 gnd.n3279 104.615
R5903 gnd.n3279 gnd.n3269 104.615
R5904 gnd.n3272 gnd.n3269 104.615
R5905 gnd.n3257 gnd.n3256 104.615
R5906 gnd.n3256 gnd.n3234 104.615
R5907 gnd.n3249 gnd.n3234 104.615
R5908 gnd.n3249 gnd.n3248 104.615
R5909 gnd.n3248 gnd.n3238 104.615
R5910 gnd.n3241 gnd.n3238 104.615
R5911 gnd.n2630 gnd.t30 100.632
R5912 gnd.n2200 gnd.t61 100.632
R5913 gnd.n7142 gnd.n93 99.6594
R5914 gnd.n7140 gnd.n7139 99.6594
R5915 gnd.n7135 gnd.n100 99.6594
R5916 gnd.n7133 gnd.n7132 99.6594
R5917 gnd.n7128 gnd.n107 99.6594
R5918 gnd.n7126 gnd.n7125 99.6594
R5919 gnd.n7121 gnd.n114 99.6594
R5920 gnd.n7119 gnd.n7118 99.6594
R5921 gnd.n7111 gnd.n121 99.6594
R5922 gnd.n7109 gnd.n7108 99.6594
R5923 gnd.n7104 gnd.n128 99.6594
R5924 gnd.n7102 gnd.n7101 99.6594
R5925 gnd.n7097 gnd.n135 99.6594
R5926 gnd.n7095 gnd.n7094 99.6594
R5927 gnd.n7090 gnd.n142 99.6594
R5928 gnd.n7088 gnd.n7087 99.6594
R5929 gnd.n7083 gnd.n149 99.6594
R5930 gnd.n7081 gnd.n7080 99.6594
R5931 gnd.n154 gnd.n153 99.6594
R5932 gnd.n5515 gnd.n1131 99.6594
R5933 gnd.n5519 gnd.n5518 99.6594
R5934 gnd.n5526 gnd.n5525 99.6594
R5935 gnd.n5529 gnd.n5528 99.6594
R5936 gnd.n5536 gnd.n5535 99.6594
R5937 gnd.n5539 gnd.n5538 99.6594
R5938 gnd.n5547 gnd.n5546 99.6594
R5939 gnd.n5550 gnd.n5549 99.6594
R5940 gnd.n5560 gnd.n5559 99.6594
R5941 gnd.n5563 gnd.n5562 99.6594
R5942 gnd.n5570 gnd.n5569 99.6594
R5943 gnd.n5573 gnd.n5572 99.6594
R5944 gnd.n5580 gnd.n5579 99.6594
R5945 gnd.n5583 gnd.n5582 99.6594
R5946 gnd.n5590 gnd.n5589 99.6594
R5947 gnd.n5593 gnd.n5592 99.6594
R5948 gnd.n5601 gnd.n5600 99.6594
R5949 gnd.n5604 gnd.n5603 99.6594
R5950 gnd.n1960 gnd.n1959 99.6594
R5951 gnd.n1955 gnd.n1914 99.6594
R5952 gnd.n1951 gnd.n1913 99.6594
R5953 gnd.n1947 gnd.n1912 99.6594
R5954 gnd.n1943 gnd.n1911 99.6594
R5955 gnd.n1939 gnd.n1910 99.6594
R5956 gnd.n1935 gnd.n1909 99.6594
R5957 gnd.n1907 gnd.n1906 99.6594
R5958 gnd.n4338 gnd.n4337 99.6594
R5959 gnd.n4335 gnd.n4334 99.6594
R5960 gnd.n4330 gnd.n1969 99.6594
R5961 gnd.n4328 gnd.n4327 99.6594
R5962 gnd.n4323 gnd.n1976 99.6594
R5963 gnd.n4321 gnd.n4320 99.6594
R5964 gnd.n4316 gnd.n1983 99.6594
R5965 gnd.n4314 gnd.n4313 99.6594
R5966 gnd.n4309 gnd.n1992 99.6594
R5967 gnd.n4307 gnd.n4306 99.6594
R5968 gnd.n3840 gnd.n3839 99.6594
R5969 gnd.n3834 gnd.n3612 99.6594
R5970 gnd.n3831 gnd.n3613 99.6594
R5971 gnd.n3827 gnd.n3614 99.6594
R5972 gnd.n3823 gnd.n3615 99.6594
R5973 gnd.n3819 gnd.n3616 99.6594
R5974 gnd.n3815 gnd.n3617 99.6594
R5975 gnd.n3811 gnd.n3618 99.6594
R5976 gnd.n3807 gnd.n3619 99.6594
R5977 gnd.n3802 gnd.n3620 99.6594
R5978 gnd.n3798 gnd.n3621 99.6594
R5979 gnd.n3794 gnd.n3622 99.6594
R5980 gnd.n3790 gnd.n3623 99.6594
R5981 gnd.n3786 gnd.n3624 99.6594
R5982 gnd.n3782 gnd.n3625 99.6594
R5983 gnd.n3778 gnd.n3626 99.6594
R5984 gnd.n3774 gnd.n3627 99.6594
R5985 gnd.n3770 gnd.n3628 99.6594
R5986 gnd.n3740 gnd.n3629 99.6594
R5987 gnd.n3602 gnd.n2183 99.6594
R5988 gnd.n3600 gnd.n2182 99.6594
R5989 gnd.n3596 gnd.n2181 99.6594
R5990 gnd.n3592 gnd.n2180 99.6594
R5991 gnd.n3588 gnd.n2179 99.6594
R5992 gnd.n3584 gnd.n2178 99.6594
R5993 gnd.n3580 gnd.n2177 99.6594
R5994 gnd.n3512 gnd.n2176 99.6594
R5995 gnd.n2842 gnd.n2573 99.6594
R5996 gnd.n2599 gnd.n2580 99.6594
R5997 gnd.n2601 gnd.n2581 99.6594
R5998 gnd.n2609 gnd.n2582 99.6594
R5999 gnd.n2611 gnd.n2583 99.6594
R6000 gnd.n2619 gnd.n2584 99.6594
R6001 gnd.n2621 gnd.n2585 99.6594
R6002 gnd.n2629 gnd.n2586 99.6594
R6003 gnd.n3570 gnd.n2163 99.6594
R6004 gnd.n3566 gnd.n2164 99.6594
R6005 gnd.n3562 gnd.n2165 99.6594
R6006 gnd.n3558 gnd.n2166 99.6594
R6007 gnd.n3554 gnd.n2167 99.6594
R6008 gnd.n3550 gnd.n2168 99.6594
R6009 gnd.n3546 gnd.n2169 99.6594
R6010 gnd.n3542 gnd.n2170 99.6594
R6011 gnd.n3538 gnd.n2171 99.6594
R6012 gnd.n3534 gnd.n2172 99.6594
R6013 gnd.n3530 gnd.n2173 99.6594
R6014 gnd.n3526 gnd.n2174 99.6594
R6015 gnd.n3522 gnd.n2175 99.6594
R6016 gnd.n2757 gnd.n2756 99.6594
R6017 gnd.n2751 gnd.n2668 99.6594
R6018 gnd.n2748 gnd.n2669 99.6594
R6019 gnd.n2744 gnd.n2670 99.6594
R6020 gnd.n2740 gnd.n2671 99.6594
R6021 gnd.n2736 gnd.n2672 99.6594
R6022 gnd.n2732 gnd.n2673 99.6594
R6023 gnd.n2728 gnd.n2674 99.6594
R6024 gnd.n2724 gnd.n2675 99.6594
R6025 gnd.n2720 gnd.n2676 99.6594
R6026 gnd.n2716 gnd.n2677 99.6594
R6027 gnd.n2712 gnd.n2678 99.6594
R6028 gnd.n2759 gnd.n2667 99.6594
R6029 gnd.n6991 gnd.n6990 99.6594
R6030 gnd.n6996 gnd.n6995 99.6594
R6031 gnd.n6999 gnd.n6998 99.6594
R6032 gnd.n7004 gnd.n7003 99.6594
R6033 gnd.n7007 gnd.n7006 99.6594
R6034 gnd.n7012 gnd.n7011 99.6594
R6035 gnd.n7015 gnd.n7014 99.6594
R6036 gnd.n7020 gnd.n7019 99.6594
R6037 gnd.n7023 gnd.n80 99.6594
R6038 gnd.n5207 gnd.n5206 99.6594
R6039 gnd.n5210 gnd.n5209 99.6594
R6040 gnd.n5226 gnd.n5225 99.6594
R6041 gnd.n5229 gnd.n5228 99.6594
R6042 gnd.n5245 gnd.n5244 99.6594
R6043 gnd.n5248 gnd.n5247 99.6594
R6044 gnd.n5264 gnd.n5263 99.6594
R6045 gnd.n5267 gnd.n5266 99.6594
R6046 gnd.n5285 gnd.n5284 99.6594
R6047 gnd.n4137 gnd.n4136 99.6594
R6048 gnd.n4140 gnd.n4139 99.6594
R6049 gnd.n4150 gnd.n4149 99.6594
R6050 gnd.n4159 gnd.n4158 99.6594
R6051 gnd.n4162 gnd.n4161 99.6594
R6052 gnd.n4173 gnd.n4172 99.6594
R6053 gnd.n4182 gnd.n4181 99.6594
R6054 gnd.n4185 gnd.n4184 99.6594
R6055 gnd.n4196 gnd.n4195 99.6594
R6056 gnd.n3843 gnd.n3842 99.6594
R6057 gnd.n3651 gnd.n3630 99.6594
R6058 gnd.n3655 gnd.n3631 99.6594
R6059 gnd.n3661 gnd.n3632 99.6594
R6060 gnd.n3665 gnd.n3633 99.6594
R6061 gnd.n3671 gnd.n3634 99.6594
R6062 gnd.n3675 gnd.n3635 99.6594
R6063 gnd.n3681 gnd.n3636 99.6594
R6064 gnd.n3685 gnd.n3637 99.6594
R6065 gnd.n3842 gnd.n2160 99.6594
R6066 gnd.n3654 gnd.n3630 99.6594
R6067 gnd.n3660 gnd.n3631 99.6594
R6068 gnd.n3664 gnd.n3632 99.6594
R6069 gnd.n3670 gnd.n3633 99.6594
R6070 gnd.n3674 gnd.n3634 99.6594
R6071 gnd.n3680 gnd.n3635 99.6594
R6072 gnd.n3684 gnd.n3636 99.6594
R6073 gnd.n3638 gnd.n3637 99.6594
R6074 gnd.n4195 gnd.n4194 99.6594
R6075 gnd.n4184 gnd.n4183 99.6594
R6076 gnd.n4181 gnd.n4174 99.6594
R6077 gnd.n4172 gnd.n4171 99.6594
R6078 gnd.n4161 gnd.n4160 99.6594
R6079 gnd.n4158 gnd.n4151 99.6594
R6080 gnd.n4149 gnd.n4148 99.6594
R6081 gnd.n4139 gnd.n4138 99.6594
R6082 gnd.n4136 gnd.n4135 99.6594
R6083 gnd.n5208 gnd.n5207 99.6594
R6084 gnd.n5209 gnd.n5191 99.6594
R6085 gnd.n5227 gnd.n5226 99.6594
R6086 gnd.n5228 gnd.n5182 99.6594
R6087 gnd.n5246 gnd.n5245 99.6594
R6088 gnd.n5247 gnd.n5173 99.6594
R6089 gnd.n5265 gnd.n5264 99.6594
R6090 gnd.n5266 gnd.n5164 99.6594
R6091 gnd.n5286 gnd.n5285 99.6594
R6092 gnd.n7024 gnd.n7023 99.6594
R6093 gnd.n7019 gnd.n7018 99.6594
R6094 gnd.n7014 gnd.n7013 99.6594
R6095 gnd.n7011 gnd.n7010 99.6594
R6096 gnd.n7006 gnd.n7005 99.6594
R6097 gnd.n7003 gnd.n7002 99.6594
R6098 gnd.n6998 gnd.n6997 99.6594
R6099 gnd.n6995 gnd.n6994 99.6594
R6100 gnd.n6990 gnd.n6989 99.6594
R6101 gnd.n2757 gnd.n2680 99.6594
R6102 gnd.n2749 gnd.n2668 99.6594
R6103 gnd.n2745 gnd.n2669 99.6594
R6104 gnd.n2741 gnd.n2670 99.6594
R6105 gnd.n2737 gnd.n2671 99.6594
R6106 gnd.n2733 gnd.n2672 99.6594
R6107 gnd.n2729 gnd.n2673 99.6594
R6108 gnd.n2725 gnd.n2674 99.6594
R6109 gnd.n2721 gnd.n2675 99.6594
R6110 gnd.n2717 gnd.n2676 99.6594
R6111 gnd.n2713 gnd.n2677 99.6594
R6112 gnd.n2709 gnd.n2678 99.6594
R6113 gnd.n2760 gnd.n2759 99.6594
R6114 gnd.n3525 gnd.n2175 99.6594
R6115 gnd.n3529 gnd.n2174 99.6594
R6116 gnd.n3533 gnd.n2173 99.6594
R6117 gnd.n3537 gnd.n2172 99.6594
R6118 gnd.n3541 gnd.n2171 99.6594
R6119 gnd.n3545 gnd.n2170 99.6594
R6120 gnd.n3549 gnd.n2169 99.6594
R6121 gnd.n3553 gnd.n2168 99.6594
R6122 gnd.n3557 gnd.n2167 99.6594
R6123 gnd.n3561 gnd.n2166 99.6594
R6124 gnd.n3565 gnd.n2165 99.6594
R6125 gnd.n3569 gnd.n2164 99.6594
R6126 gnd.n2204 gnd.n2163 99.6594
R6127 gnd.n2843 gnd.n2842 99.6594
R6128 gnd.n2602 gnd.n2580 99.6594
R6129 gnd.n2608 gnd.n2581 99.6594
R6130 gnd.n2612 gnd.n2582 99.6594
R6131 gnd.n2618 gnd.n2583 99.6594
R6132 gnd.n2622 gnd.n2584 99.6594
R6133 gnd.n2628 gnd.n2585 99.6594
R6134 gnd.n2586 gnd.n2570 99.6594
R6135 gnd.n3579 gnd.n2176 99.6594
R6136 gnd.n3583 gnd.n2177 99.6594
R6137 gnd.n3587 gnd.n2178 99.6594
R6138 gnd.n3591 gnd.n2179 99.6594
R6139 gnd.n3595 gnd.n2180 99.6594
R6140 gnd.n3599 gnd.n2181 99.6594
R6141 gnd.n3603 gnd.n2182 99.6594
R6142 gnd.n2185 gnd.n2183 99.6594
R6143 gnd.n3840 gnd.n3700 99.6594
R6144 gnd.n3832 gnd.n3612 99.6594
R6145 gnd.n3828 gnd.n3613 99.6594
R6146 gnd.n3824 gnd.n3614 99.6594
R6147 gnd.n3820 gnd.n3615 99.6594
R6148 gnd.n3816 gnd.n3616 99.6594
R6149 gnd.n3812 gnd.n3617 99.6594
R6150 gnd.n3808 gnd.n3618 99.6594
R6151 gnd.n3803 gnd.n3619 99.6594
R6152 gnd.n3799 gnd.n3620 99.6594
R6153 gnd.n3795 gnd.n3621 99.6594
R6154 gnd.n3791 gnd.n3622 99.6594
R6155 gnd.n3787 gnd.n3623 99.6594
R6156 gnd.n3783 gnd.n3624 99.6594
R6157 gnd.n3779 gnd.n3625 99.6594
R6158 gnd.n3775 gnd.n3626 99.6594
R6159 gnd.n3771 gnd.n3627 99.6594
R6160 gnd.n3739 gnd.n3628 99.6594
R6161 gnd.n3763 gnd.n3629 99.6594
R6162 gnd.n4308 gnd.n4307 99.6594
R6163 gnd.n1992 gnd.n1984 99.6594
R6164 gnd.n4315 gnd.n4314 99.6594
R6165 gnd.n1983 gnd.n1977 99.6594
R6166 gnd.n4322 gnd.n4321 99.6594
R6167 gnd.n1976 gnd.n1970 99.6594
R6168 gnd.n4329 gnd.n4328 99.6594
R6169 gnd.n1969 gnd.n1963 99.6594
R6170 gnd.n4336 gnd.n4335 99.6594
R6171 gnd.n4339 gnd.n4338 99.6594
R6172 gnd.n1934 gnd.n1908 99.6594
R6173 gnd.n1938 gnd.n1909 99.6594
R6174 gnd.n1942 gnd.n1910 99.6594
R6175 gnd.n1946 gnd.n1911 99.6594
R6176 gnd.n1950 gnd.n1912 99.6594
R6177 gnd.n1954 gnd.n1913 99.6594
R6178 gnd.n1916 gnd.n1914 99.6594
R6179 gnd.n1960 gnd.n1915 99.6594
R6180 gnd.n5516 gnd.n5515 99.6594
R6181 gnd.n5518 gnd.n5507 99.6594
R6182 gnd.n5527 gnd.n5526 99.6594
R6183 gnd.n5528 gnd.n5503 99.6594
R6184 gnd.n5537 gnd.n5536 99.6594
R6185 gnd.n5538 gnd.n5499 99.6594
R6186 gnd.n5548 gnd.n5547 99.6594
R6187 gnd.n5497 gnd.n1288 99.6594
R6188 gnd.n5561 gnd.n5560 99.6594
R6189 gnd.n5562 gnd.n1284 99.6594
R6190 gnd.n5571 gnd.n5570 99.6594
R6191 gnd.n5572 gnd.n1280 99.6594
R6192 gnd.n5581 gnd.n5580 99.6594
R6193 gnd.n5582 gnd.n1276 99.6594
R6194 gnd.n5591 gnd.n5590 99.6594
R6195 gnd.n5592 gnd.n1272 99.6594
R6196 gnd.n5602 gnd.n5601 99.6594
R6197 gnd.n5605 gnd.n5604 99.6594
R6198 gnd.n153 gnd.n150 99.6594
R6199 gnd.n7082 gnd.n7081 99.6594
R6200 gnd.n149 gnd.n143 99.6594
R6201 gnd.n7089 gnd.n7088 99.6594
R6202 gnd.n142 gnd.n136 99.6594
R6203 gnd.n7096 gnd.n7095 99.6594
R6204 gnd.n135 gnd.n129 99.6594
R6205 gnd.n7103 gnd.n7102 99.6594
R6206 gnd.n128 gnd.n122 99.6594
R6207 gnd.n7110 gnd.n7109 99.6594
R6208 gnd.n121 gnd.n115 99.6594
R6209 gnd.n7120 gnd.n7119 99.6594
R6210 gnd.n114 gnd.n108 99.6594
R6211 gnd.n7127 gnd.n7126 99.6594
R6212 gnd.n107 gnd.n101 99.6594
R6213 gnd.n7134 gnd.n7133 99.6594
R6214 gnd.n100 gnd.n94 99.6594
R6215 gnd.n7141 gnd.n7140 99.6594
R6216 gnd.n93 gnd.n90 99.6594
R6217 gnd.n4243 gnd.n4242 99.6594
R6218 gnd.n4143 gnd.n4113 99.6594
R6219 gnd.n4145 gnd.n4114 99.6594
R6220 gnd.n4155 gnd.n4115 99.6594
R6221 gnd.n4166 gnd.n4116 99.6594
R6222 gnd.n4168 gnd.n4117 99.6594
R6223 gnd.n4178 gnd.n4118 99.6594
R6224 gnd.n4191 gnd.n4119 99.6594
R6225 gnd.n4192 gnd.n4120 99.6594
R6226 gnd.n4121 gnd.n2003 99.6594
R6227 gnd.n4123 gnd.n4122 99.6594
R6228 gnd.n4124 gnd.n2008 99.6594
R6229 gnd.n4125 gnd.n2014 99.6594
R6230 gnd.n4126 gnd.n2016 99.6594
R6231 gnd.n4243 gnd.n4128 99.6594
R6232 gnd.n4144 gnd.n4113 99.6594
R6233 gnd.n4154 gnd.n4114 99.6594
R6234 gnd.n4165 gnd.n4115 99.6594
R6235 gnd.n4167 gnd.n4116 99.6594
R6236 gnd.n4177 gnd.n4117 99.6594
R6237 gnd.n4190 gnd.n4118 99.6594
R6238 gnd.n4193 gnd.n4119 99.6594
R6239 gnd.n4120 gnd.n2002 99.6594
R6240 gnd.n4121 gnd.n2004 99.6594
R6241 gnd.n4123 gnd.n2007 99.6594
R6242 gnd.n4124 gnd.n2009 99.6594
R6243 gnd.n4125 gnd.n2015 99.6594
R6244 gnd.n4126 gnd.n2019 99.6594
R6245 gnd.n5216 gnd.n5196 99.6594
R6246 gnd.n5220 gnd.n5218 99.6594
R6247 gnd.n5235 gnd.n5187 99.6594
R6248 gnd.n5239 gnd.n5237 99.6594
R6249 gnd.n5254 gnd.n5178 99.6594
R6250 gnd.n5258 gnd.n5256 99.6594
R6251 gnd.n5273 gnd.n5169 99.6594
R6252 gnd.n5276 gnd.n5275 99.6594
R6253 gnd.n5277 gnd.n5158 99.6594
R6254 gnd.n5296 gnd.n5295 99.6594
R6255 gnd.n5297 gnd.n5154 99.6594
R6256 gnd.n5306 gnd.n5305 99.6594
R6257 gnd.n5307 gnd.n5150 99.6594
R6258 gnd.n5319 gnd.n5318 99.6594
R6259 gnd.n5318 gnd.n5317 99.6594
R6260 gnd.n5308 gnd.n5307 99.6594
R6261 gnd.n5305 gnd.n5304 99.6594
R6262 gnd.n5298 gnd.n5297 99.6594
R6263 gnd.n5295 gnd.n5294 99.6594
R6264 gnd.n5278 gnd.n5277 99.6594
R6265 gnd.n5275 gnd.n5274 99.6594
R6266 gnd.n5257 gnd.n5169 99.6594
R6267 gnd.n5256 gnd.n5255 99.6594
R6268 gnd.n5238 gnd.n5178 99.6594
R6269 gnd.n5237 gnd.n5236 99.6594
R6270 gnd.n5219 gnd.n5187 99.6594
R6271 gnd.n5218 gnd.n5217 99.6594
R6272 gnd.n5196 gnd.n1105 99.6594
R6273 gnd.n2010 gnd.t95 98.63
R6274 gnd.n7021 gnd.t81 98.63
R6275 gnd.n5161 gnd.t72 98.63
R6276 gnd.n4186 gnd.t87 98.63
R6277 gnd.n5552 gnd.t69 98.63
R6278 gnd.n1268 gnd.t37 98.63
R6279 gnd.n156 gnd.t22 98.63
R6280 gnd.n7113 gnd.t50 98.63
R6281 gnd.n3719 gnd.t120 98.63
R6282 gnd.n3741 gnd.t111 98.63
R6283 gnd.n3640 gnd.t108 98.63
R6284 gnd.n1989 gnd.t43 98.63
R6285 gnd.n1900 gnd.t84 98.63
R6286 gnd.n5309 gnd.t78 98.63
R6287 gnd.n1834 gnd.t114 96.6984
R6288 gnd.n1329 gnd.t47 96.6984
R6289 gnd.n1831 gnd.t66 96.6906
R6290 gnd.n5359 gnd.t100 96.6906
R6291 gnd.n1819 gnd.n1818 81.8399
R6292 gnd.n2631 gnd.t29 74.8376
R6293 gnd.n2201 gnd.t62 74.8376
R6294 gnd.n1835 gnd.t113 72.8438
R6295 gnd.n1330 gnd.t48 72.8438
R6296 gnd.n1820 gnd.n1813 72.8411
R6297 gnd.n1826 gnd.n1811 72.8411
R6298 gnd.n5355 gnd.n5354 72.8411
R6299 gnd.n2011 gnd.t94 72.836
R6300 gnd.n1832 gnd.t65 72.836
R6301 gnd.n5360 gnd.t101 72.836
R6302 gnd.n7022 gnd.t82 72.836
R6303 gnd.n5162 gnd.t71 72.836
R6304 gnd.n4187 gnd.t88 72.836
R6305 gnd.n5553 gnd.t68 72.836
R6306 gnd.n1269 gnd.t36 72.836
R6307 gnd.n157 gnd.t23 72.836
R6308 gnd.n7114 gnd.t51 72.836
R6309 gnd.n3720 gnd.t119 72.836
R6310 gnd.n3742 gnd.t110 72.836
R6311 gnd.n3641 gnd.t107 72.836
R6312 gnd.n1990 gnd.t44 72.836
R6313 gnd.n1901 gnd.t85 72.836
R6314 gnd.n5310 gnd.t79 72.836
R6315 gnd.n5420 gnd.n1297 71.676
R6316 gnd.n5416 gnd.n1298 71.676
R6317 gnd.n5412 gnd.n1299 71.676
R6318 gnd.n5408 gnd.n1300 71.676
R6319 gnd.n5404 gnd.n1301 71.676
R6320 gnd.n5400 gnd.n1302 71.676
R6321 gnd.n5396 gnd.n1303 71.676
R6322 gnd.n5392 gnd.n1304 71.676
R6323 gnd.n5388 gnd.n1305 71.676
R6324 gnd.n5384 gnd.n1306 71.676
R6325 gnd.n5380 gnd.n1307 71.676
R6326 gnd.n5376 gnd.n1308 71.676
R6327 gnd.n5372 gnd.n1309 71.676
R6328 gnd.n5368 gnd.n1310 71.676
R6329 gnd.n5363 gnd.n1311 71.676
R6330 gnd.n1312 gnd.n1295 71.676
R6331 gnd.n5492 gnd.n1294 71.676
R6332 gnd.n5490 gnd.n5489 71.676
R6333 gnd.n5484 gnd.n1327 71.676
R6334 gnd.n5480 gnd.n1326 71.676
R6335 gnd.n5476 gnd.n1325 71.676
R6336 gnd.n5472 gnd.n1324 71.676
R6337 gnd.n5468 gnd.n1323 71.676
R6338 gnd.n5464 gnd.n1322 71.676
R6339 gnd.n5460 gnd.n1321 71.676
R6340 gnd.n5456 gnd.n1320 71.676
R6341 gnd.n5452 gnd.n1319 71.676
R6342 gnd.n5448 gnd.n1318 71.676
R6343 gnd.n5444 gnd.n1317 71.676
R6344 gnd.n5440 gnd.n1316 71.676
R6345 gnd.n5436 gnd.n1315 71.676
R6346 gnd.n5432 gnd.n1314 71.676
R6347 gnd.n5428 gnd.n1313 71.676
R6348 gnd.n4411 gnd.n4410 71.676
R6349 gnd.n4405 gnd.n1775 71.676
R6350 gnd.n4402 gnd.n1776 71.676
R6351 gnd.n4398 gnd.n1777 71.676
R6352 gnd.n4394 gnd.n1778 71.676
R6353 gnd.n4390 gnd.n1779 71.676
R6354 gnd.n4386 gnd.n1780 71.676
R6355 gnd.n4382 gnd.n1781 71.676
R6356 gnd.n4378 gnd.n1782 71.676
R6357 gnd.n4374 gnd.n1783 71.676
R6358 gnd.n4370 gnd.n1784 71.676
R6359 gnd.n4366 gnd.n1785 71.676
R6360 gnd.n4362 gnd.n1786 71.676
R6361 gnd.n4358 gnd.n1787 71.676
R6362 gnd.n4354 gnd.n1788 71.676
R6363 gnd.n4350 gnd.n1789 71.676
R6364 gnd.n4346 gnd.n1791 71.676
R6365 gnd.n1894 gnd.n1792 71.676
R6366 gnd.n1889 gnd.n1793 71.676
R6367 gnd.n1885 gnd.n1794 71.676
R6368 gnd.n1881 gnd.n1795 71.676
R6369 gnd.n1877 gnd.n1796 71.676
R6370 gnd.n1873 gnd.n1797 71.676
R6371 gnd.n1869 gnd.n1798 71.676
R6372 gnd.n1865 gnd.n1799 71.676
R6373 gnd.n1861 gnd.n1800 71.676
R6374 gnd.n1857 gnd.n1801 71.676
R6375 gnd.n1853 gnd.n1802 71.676
R6376 gnd.n1849 gnd.n1803 71.676
R6377 gnd.n1845 gnd.n1804 71.676
R6378 gnd.n1841 gnd.n1805 71.676
R6379 gnd.n1837 gnd.n1806 71.676
R6380 gnd.n4411 gnd.n1809 71.676
R6381 gnd.n4403 gnd.n1775 71.676
R6382 gnd.n4399 gnd.n1776 71.676
R6383 gnd.n4395 gnd.n1777 71.676
R6384 gnd.n4391 gnd.n1778 71.676
R6385 gnd.n4387 gnd.n1779 71.676
R6386 gnd.n4383 gnd.n1780 71.676
R6387 gnd.n4379 gnd.n1781 71.676
R6388 gnd.n4375 gnd.n1782 71.676
R6389 gnd.n4371 gnd.n1783 71.676
R6390 gnd.n4367 gnd.n1784 71.676
R6391 gnd.n4363 gnd.n1785 71.676
R6392 gnd.n4359 gnd.n1786 71.676
R6393 gnd.n4355 gnd.n1787 71.676
R6394 gnd.n4351 gnd.n1788 71.676
R6395 gnd.n4347 gnd.n1790 71.676
R6396 gnd.n1895 gnd.n1791 71.676
R6397 gnd.n1890 gnd.n1792 71.676
R6398 gnd.n1886 gnd.n1793 71.676
R6399 gnd.n1882 gnd.n1794 71.676
R6400 gnd.n1878 gnd.n1795 71.676
R6401 gnd.n1874 gnd.n1796 71.676
R6402 gnd.n1870 gnd.n1797 71.676
R6403 gnd.n1866 gnd.n1798 71.676
R6404 gnd.n1862 gnd.n1799 71.676
R6405 gnd.n1858 gnd.n1800 71.676
R6406 gnd.n1854 gnd.n1801 71.676
R6407 gnd.n1850 gnd.n1802 71.676
R6408 gnd.n1846 gnd.n1803 71.676
R6409 gnd.n1842 gnd.n1804 71.676
R6410 gnd.n1838 gnd.n1805 71.676
R6411 gnd.n1806 gnd.n1767 71.676
R6412 gnd.n5431 gnd.n1313 71.676
R6413 gnd.n5435 gnd.n1314 71.676
R6414 gnd.n5439 gnd.n1315 71.676
R6415 gnd.n5443 gnd.n1316 71.676
R6416 gnd.n5447 gnd.n1317 71.676
R6417 gnd.n5451 gnd.n1318 71.676
R6418 gnd.n5455 gnd.n1319 71.676
R6419 gnd.n5459 gnd.n1320 71.676
R6420 gnd.n5463 gnd.n1321 71.676
R6421 gnd.n5467 gnd.n1322 71.676
R6422 gnd.n5471 gnd.n1323 71.676
R6423 gnd.n5475 gnd.n1324 71.676
R6424 gnd.n5479 gnd.n1325 71.676
R6425 gnd.n5483 gnd.n1326 71.676
R6426 gnd.n1328 gnd.n1327 71.676
R6427 gnd.n5491 gnd.n5490 71.676
R6428 gnd.n5495 gnd.n5494 71.676
R6429 gnd.n5362 gnd.n1312 71.676
R6430 gnd.n5367 gnd.n1311 71.676
R6431 gnd.n5371 gnd.n1310 71.676
R6432 gnd.n5375 gnd.n1309 71.676
R6433 gnd.n5379 gnd.n1308 71.676
R6434 gnd.n5383 gnd.n1307 71.676
R6435 gnd.n5387 gnd.n1306 71.676
R6436 gnd.n5391 gnd.n1305 71.676
R6437 gnd.n5395 gnd.n1304 71.676
R6438 gnd.n5399 gnd.n1303 71.676
R6439 gnd.n5403 gnd.n1302 71.676
R6440 gnd.n5407 gnd.n1301 71.676
R6441 gnd.n5411 gnd.n1300 71.676
R6442 gnd.n5415 gnd.n1299 71.676
R6443 gnd.n5419 gnd.n1298 71.676
R6444 gnd.n1335 gnd.n1297 71.676
R6445 gnd.n8 gnd.t282 69.1507
R6446 gnd.n14 gnd.t203 68.4792
R6447 gnd.n13 gnd.t224 68.4792
R6448 gnd.n12 gnd.t136 68.4792
R6449 gnd.n11 gnd.t220 68.4792
R6450 gnd.n10 gnd.t131 68.4792
R6451 gnd.n9 gnd.t5 68.4792
R6452 gnd.n8 gnd.t169 68.4792
R6453 gnd.n2758 gnd.n2662 64.369
R6454 gnd.n3841 gnd.n2151 63.0944
R6455 gnd.n7150 gnd.n83 63.0944
R6456 gnd.n1892 gnd.n1835 59.5399
R6457 gnd.n5486 gnd.n1330 59.5399
R6458 gnd.n1833 gnd.n1832 59.5399
R6459 gnd.n5365 gnd.n5360 59.5399
R6460 gnd.n1830 gnd.n1829 59.1804
R6461 gnd.n3611 gnd.n2161 57.3586
R6462 gnd.n2417 gnd.t283 56.607
R6463 gnd.n40 gnd.t278 56.607
R6464 gnd.n2394 gnd.t250 56.407
R6465 gnd.n2405 gnd.t254 56.407
R6466 gnd.n17 gnd.t12 56.407
R6467 gnd.n28 gnd.t150 56.407
R6468 gnd.n2426 gnd.t234 55.8337
R6469 gnd.n2403 gnd.t261 55.8337
R6470 gnd.n2414 gnd.t273 55.8337
R6471 gnd.n49 gnd.t141 55.8337
R6472 gnd.n26 gnd.t268 55.8337
R6473 gnd.n37 gnd.t255 55.8337
R6474 gnd.n1817 gnd.n1816 54.358
R6475 gnd.n5352 gnd.n5351 54.358
R6476 gnd.n2417 gnd.n2416 53.0052
R6477 gnd.n2419 gnd.n2418 53.0052
R6478 gnd.n2421 gnd.n2420 53.0052
R6479 gnd.n2423 gnd.n2422 53.0052
R6480 gnd.n2425 gnd.n2424 53.0052
R6481 gnd.n2394 gnd.n2393 53.0052
R6482 gnd.n2396 gnd.n2395 53.0052
R6483 gnd.n2398 gnd.n2397 53.0052
R6484 gnd.n2400 gnd.n2399 53.0052
R6485 gnd.n2402 gnd.n2401 53.0052
R6486 gnd.n2405 gnd.n2404 53.0052
R6487 gnd.n2407 gnd.n2406 53.0052
R6488 gnd.n2409 gnd.n2408 53.0052
R6489 gnd.n2411 gnd.n2410 53.0052
R6490 gnd.n2413 gnd.n2412 53.0052
R6491 gnd.n48 gnd.n47 53.0052
R6492 gnd.n46 gnd.n45 53.0052
R6493 gnd.n44 gnd.n43 53.0052
R6494 gnd.n42 gnd.n41 53.0052
R6495 gnd.n40 gnd.n39 53.0052
R6496 gnd.n25 gnd.n24 53.0052
R6497 gnd.n23 gnd.n22 53.0052
R6498 gnd.n21 gnd.n20 53.0052
R6499 gnd.n19 gnd.n18 53.0052
R6500 gnd.n17 gnd.n16 53.0052
R6501 gnd.n36 gnd.n35 53.0052
R6502 gnd.n34 gnd.n33 53.0052
R6503 gnd.n32 gnd.n31 53.0052
R6504 gnd.n30 gnd.n29 53.0052
R6505 gnd.n28 gnd.n27 53.0052
R6506 gnd.n5343 gnd.n5342 52.4801
R6507 gnd.n3463 gnd.t176 52.3082
R6508 gnd.n3431 gnd.t145 52.3082
R6509 gnd.n3399 gnd.t230 52.3082
R6510 gnd.n3368 gnd.t155 52.3082
R6511 gnd.n3336 gnd.t199 52.3082
R6512 gnd.n3304 gnd.t277 52.3082
R6513 gnd.n3272 gnd.t185 52.3082
R6514 gnd.n3241 gnd.t287 52.3082
R6515 gnd.n3293 gnd.n3261 51.4173
R6516 gnd.n3357 gnd.n3356 50.455
R6517 gnd.n3325 gnd.n3324 50.455
R6518 gnd.n3293 gnd.n3292 50.455
R6519 gnd.n5554 gnd.n5496 45.6325
R6520 gnd.n4348 gnd.n4344 45.6325
R6521 gnd.n2705 gnd.n2704 45.1884
R6522 gnd.n2227 gnd.n2226 45.1884
R6523 gnd.n5423 gnd.n5358 44.3322
R6524 gnd.n1820 gnd.n1819 44.3189
R6525 gnd.n2012 gnd.n2011 42.2793
R6526 gnd.n2706 gnd.n2705 42.2793
R6527 gnd.n2228 gnd.n2227 42.2793
R6528 gnd.n2632 gnd.n2631 42.2793
R6529 gnd.n3578 gnd.n2201 42.2793
R6530 gnd.n7026 gnd.n7022 42.2793
R6531 gnd.n5163 gnd.n5162 42.2793
R6532 gnd.n4188 gnd.n4187 42.2793
R6533 gnd.n1270 gnd.n1269 42.2793
R6534 gnd.n7078 gnd.n157 42.2793
R6535 gnd.n7115 gnd.n7114 42.2793
R6536 gnd.n3805 gnd.n3720 42.2793
R6537 gnd.n3743 gnd.n3742 42.2793
R6538 gnd.n3642 gnd.n3641 42.2793
R6539 gnd.n1991 gnd.n1990 42.2793
R6540 gnd.n5311 gnd.n5310 42.2793
R6541 gnd.n1818 gnd.n1817 41.6274
R6542 gnd.n5353 gnd.n5352 41.6274
R6543 gnd.n6259 gnd.n6258 41.1297
R6544 gnd.n6258 gnd.n6257 41.1297
R6545 gnd.n6257 gnd.n661 41.1297
R6546 gnd.n6251 gnd.n661 41.1297
R6547 gnd.n6251 gnd.n6250 41.1297
R6548 gnd.n6250 gnd.n6249 41.1297
R6549 gnd.n6249 gnd.n668 41.1297
R6550 gnd.n6243 gnd.n668 41.1297
R6551 gnd.n6243 gnd.n6242 41.1297
R6552 gnd.n6242 gnd.n6241 41.1297
R6553 gnd.n6241 gnd.n676 41.1297
R6554 gnd.n6235 gnd.n676 41.1297
R6555 gnd.n6235 gnd.n6234 41.1297
R6556 gnd.n6234 gnd.n6233 41.1297
R6557 gnd.n6233 gnd.n684 41.1297
R6558 gnd.n6227 gnd.n684 41.1297
R6559 gnd.n6227 gnd.n6226 41.1297
R6560 gnd.n6226 gnd.n6225 41.1297
R6561 gnd.n6225 gnd.n692 41.1297
R6562 gnd.n6219 gnd.n692 41.1297
R6563 gnd.n6219 gnd.n6218 41.1297
R6564 gnd.n6218 gnd.n6217 41.1297
R6565 gnd.n6217 gnd.n700 41.1297
R6566 gnd.n6211 gnd.n700 41.1297
R6567 gnd.n6211 gnd.n6210 41.1297
R6568 gnd.n6210 gnd.n6209 41.1297
R6569 gnd.n6209 gnd.n708 41.1297
R6570 gnd.n6203 gnd.n708 41.1297
R6571 gnd.n6203 gnd.n6202 41.1297
R6572 gnd.n6202 gnd.n6201 41.1297
R6573 gnd.n6201 gnd.n716 41.1297
R6574 gnd.n6195 gnd.n716 41.1297
R6575 gnd.n6195 gnd.n6194 41.1297
R6576 gnd.n6194 gnd.n6193 41.1297
R6577 gnd.n6193 gnd.n724 41.1297
R6578 gnd.n6187 gnd.n724 41.1297
R6579 gnd.n6187 gnd.n6186 41.1297
R6580 gnd.n6186 gnd.n6185 41.1297
R6581 gnd.n6185 gnd.n732 41.1297
R6582 gnd.n6179 gnd.n732 41.1297
R6583 gnd.n6179 gnd.n6178 41.1297
R6584 gnd.n6178 gnd.n6177 41.1297
R6585 gnd.n6177 gnd.n740 41.1297
R6586 gnd.n6171 gnd.n740 41.1297
R6587 gnd.n6171 gnd.n6170 41.1297
R6588 gnd.n6170 gnd.n6169 41.1297
R6589 gnd.n6169 gnd.n748 41.1297
R6590 gnd.n6163 gnd.n748 41.1297
R6591 gnd.n6163 gnd.n6162 41.1297
R6592 gnd.n6162 gnd.n6161 41.1297
R6593 gnd.n6161 gnd.n756 41.1297
R6594 gnd.n6155 gnd.n756 41.1297
R6595 gnd.n6155 gnd.n6154 41.1297
R6596 gnd.n6154 gnd.n6153 41.1297
R6597 gnd.n6153 gnd.n764 41.1297
R6598 gnd.n6147 gnd.n764 41.1297
R6599 gnd.n6147 gnd.n6146 41.1297
R6600 gnd.n6146 gnd.n6145 41.1297
R6601 gnd.n6145 gnd.n772 41.1297
R6602 gnd.n6139 gnd.n772 41.1297
R6603 gnd.n6139 gnd.n6138 41.1297
R6604 gnd.n6138 gnd.n6137 41.1297
R6605 gnd.n6137 gnd.n780 41.1297
R6606 gnd.n6131 gnd.n780 41.1297
R6607 gnd.n6131 gnd.n6130 41.1297
R6608 gnd.n6130 gnd.n6129 41.1297
R6609 gnd.n6129 gnd.n788 41.1297
R6610 gnd.n6123 gnd.n788 41.1297
R6611 gnd.n6123 gnd.n6122 41.1297
R6612 gnd.n6122 gnd.n6121 41.1297
R6613 gnd.n6121 gnd.n796 41.1297
R6614 gnd.n6115 gnd.n796 41.1297
R6615 gnd.n6115 gnd.n6114 41.1297
R6616 gnd.n6114 gnd.n6113 41.1297
R6617 gnd.n6113 gnd.n804 41.1297
R6618 gnd.n6107 gnd.n804 41.1297
R6619 gnd.n6107 gnd.n6106 41.1297
R6620 gnd.n6106 gnd.n6105 41.1297
R6621 gnd.n6105 gnd.n812 41.1297
R6622 gnd.n6099 gnd.n812 41.1297
R6623 gnd.n6099 gnd.n6098 41.1297
R6624 gnd.n6098 gnd.n6097 41.1297
R6625 gnd.n6097 gnd.n820 41.1297
R6626 gnd.n1827 gnd.n1826 40.8975
R6627 gnd.n5356 gnd.n5355 40.8975
R6628 gnd.n5554 gnd.n5553 36.9518
R6629 gnd.n4344 gnd.n1901 36.9518
R6630 gnd.n1826 gnd.n1825 35.055
R6631 gnd.n1821 gnd.n1820 35.055
R6632 gnd.n5345 gnd.n5344 35.055
R6633 gnd.n5355 gnd.n5341 35.055
R6634 gnd.n5429 gnd.n1331 32.9371
R6635 gnd.n4425 gnd.n1766 32.9371
R6636 gnd.n2768 gnd.n2662 31.8661
R6637 gnd.n2768 gnd.n2767 31.8661
R6638 gnd.n2776 gnd.n2651 31.8661
R6639 gnd.n2784 gnd.n2651 31.8661
R6640 gnd.n2784 gnd.n2645 31.8661
R6641 gnd.n2792 gnd.n2645 31.8661
R6642 gnd.n2792 gnd.n2638 31.8661
R6643 gnd.n2830 gnd.n2638 31.8661
R6644 gnd.n2840 gnd.n2571 31.8661
R6645 gnd.n3859 gnd.n2151 31.8661
R6646 gnd.n3868 gnd.n2143 31.8661
R6647 gnd.n3868 gnd.n827 31.8661
R6648 gnd.n6090 gnd.n830 31.8661
R6649 gnd.n2026 gnd.n996 31.8661
R6650 gnd.n4112 gnd.n4111 31.8661
R6651 gnd.n4245 gnd.n4112 31.8661
R6652 gnd.n4253 gnd.n2020 31.8661
R6653 gnd.n5866 gnd.n1108 31.8661
R6654 gnd.n5860 gnd.n5859 31.8661
R6655 gnd.n5859 gnd.n5858 31.8661
R6656 gnd.n5852 gnd.n1126 31.8661
R6657 gnd.n6980 gnd.n180 31.8661
R6658 gnd.n7062 gnd.n161 31.8661
R6659 gnd.n7070 gnd.n161 31.8661
R6660 gnd.n7150 gnd.n81 31.8661
R6661 gnd.n2011 gnd.n2010 25.7944
R6662 gnd.n2631 gnd.n2630 25.7944
R6663 gnd.n2201 gnd.n2200 25.7944
R6664 gnd.n7022 gnd.n7021 25.7944
R6665 gnd.n5162 gnd.n5161 25.7944
R6666 gnd.n4187 gnd.n4186 25.7944
R6667 gnd.n5553 gnd.n5552 25.7944
R6668 gnd.n1269 gnd.n1268 25.7944
R6669 gnd.n157 gnd.n156 25.7944
R6670 gnd.n7114 gnd.n7113 25.7944
R6671 gnd.n3720 gnd.n3719 25.7944
R6672 gnd.n3742 gnd.n3741 25.7944
R6673 gnd.n3641 gnd.n3640 25.7944
R6674 gnd.n1990 gnd.n1989 25.7944
R6675 gnd.n1901 gnd.n1900 25.7944
R6676 gnd.n5310 gnd.n5309 25.7944
R6677 gnd.n2852 gnd.n2572 24.8557
R6678 gnd.n2862 gnd.n2555 24.8557
R6679 gnd.n2558 gnd.n2546 24.8557
R6680 gnd.n2883 gnd.n2547 24.8557
R6681 gnd.n2893 gnd.n2527 24.8557
R6682 gnd.n2903 gnd.n2902 24.8557
R6683 gnd.n2513 gnd.n2511 24.8557
R6684 gnd.n2934 gnd.n2933 24.8557
R6685 gnd.n2949 gnd.n2496 24.8557
R6686 gnd.n3003 gnd.n2435 24.8557
R6687 gnd.n2959 gnd.n2436 24.8557
R6688 gnd.n2996 gnd.n2447 24.8557
R6689 gnd.n2485 gnd.n2484 24.8557
R6690 gnd.n2990 gnd.n2989 24.8557
R6691 gnd.n2471 gnd.n2458 24.8557
R6692 gnd.n3029 gnd.n3028 24.8557
R6693 gnd.n3039 gnd.n2379 24.8557
R6694 gnd.n3051 gnd.n2371 24.8557
R6695 gnd.n3050 gnd.n2359 24.8557
R6696 gnd.n3069 gnd.n3068 24.8557
R6697 gnd.n3079 gnd.n2352 24.8557
R6698 gnd.n3090 gnd.n2340 24.8557
R6699 gnd.n3114 gnd.n3113 24.8557
R6700 gnd.n3125 gnd.n2323 24.8557
R6701 gnd.n3124 gnd.n2325 24.8557
R6702 gnd.n3137 gnd.n2316 24.8557
R6703 gnd.n3155 gnd.n3154 24.8557
R6704 gnd.n2307 gnd.n2296 24.8557
R6705 gnd.n3176 gnd.n2284 24.8557
R6706 gnd.n3204 gnd.n3203 24.8557
R6707 gnd.n3215 gnd.n2269 24.8557
R6708 gnd.n3226 gnd.n2262 24.8557
R6709 gnd.n3225 gnd.n2250 24.8557
R6710 gnd.n3498 gnd.n3497 24.8557
R6711 gnd.n3520 gnd.n2235 24.8557
R6712 gnd.n3135 gnd.n820 24.678
R6713 gnd.n1835 gnd.n1834 23.855
R6714 gnd.n1330 gnd.n1329 23.855
R6715 gnd.n1832 gnd.n1831 23.855
R6716 gnd.n5360 gnd.n5359 23.855
R6717 gnd.n2873 gnd.t286 23.2624
R6718 gnd.n2574 gnd.t28 22.6251
R6719 gnd.t154 gnd.n2579 21.3504
R6720 gnd.n3881 gnd.n843 21.0318
R6721 gnd.n6078 gnd.n852 21.0318
R6722 gnd.n3902 gnd.n3901 21.0318
R6723 gnd.n6072 gnd.n862 21.0318
R6724 gnd.n6066 gnd.n873 21.0318
R6725 gnd.n3929 gnd.n876 21.0318
R6726 gnd.n3939 gnd.n886 21.0318
R6727 gnd.n6054 gnd.n894 21.0318
R6728 gnd.n3950 gnd.n3949 21.0318
R6729 gnd.n3976 gnd.n2111 21.0318
R6730 gnd.n3984 gnd.n2105 21.0318
R6731 gnd.n3998 gnd.n2084 21.0318
R6732 gnd.n4004 gnd.n2077 21.0318
R6733 gnd.n2079 gnd.n2070 21.0318
R6734 gnd.n6046 gnd.n909 21.0318
R6735 gnd.n4025 gnd.n912 21.0318
R6736 gnd.n4033 gnd.n923 21.0318
R6737 gnd.n6034 gnd.n930 21.0318
R6738 gnd.n4079 gnd.n4078 21.0318
R6739 gnd.n6028 gnd.n940 21.0318
R6740 gnd.n6022 gnd.n951 21.0318
R6741 gnd.n4048 gnd.n954 21.0318
R6742 gnd.n4052 gnd.n964 21.0318
R6743 gnd.n6010 gnd.n972 21.0318
R6744 gnd.n4061 gnd.n975 21.0318
R6745 gnd.n6004 gnd.n983 21.0318
R6746 gnd.n5998 gnd.n993 21.0318
R6747 gnd.n5851 gnd.n1129 21.0318
R6748 gnd.n5845 gnd.n1141 21.0318
R6749 gnd.n5621 gnd.n1256 21.0318
R6750 gnd.n5688 gnd.n5687 21.0318
R6751 gnd.n5670 gnd.n1249 21.0318
R6752 gnd.n5708 gnd.n1241 21.0318
R6753 gnd.n5707 gnd.n1230 21.0318
R6754 gnd.n1233 gnd.n1220 21.0318
R6755 gnd.n5730 gnd.n1222 21.0318
R6756 gnd.n5740 gnd.n1212 21.0318
R6757 gnd.n5739 gnd.n1201 21.0318
R6758 gnd.n1205 gnd.n1194 21.0318
R6759 gnd.n5763 gnd.n1196 21.0318
R6760 gnd.n5773 gnd.n5772 21.0318
R6761 gnd.n5783 gnd.n1176 21.0318
R6762 gnd.n5782 gnd.n1180 21.0318
R6763 gnd.n5809 gnd.n1170 21.0318
R6764 gnd.n6927 gnd.n231 21.0318
R6765 gnd.n6932 gnd.n233 21.0318
R6766 gnd.n6921 gnd.n223 21.0318
R6767 gnd.n6940 gnd.n225 21.0318
R6768 gnd.n6948 gnd.n211 21.0318
R6769 gnd.n6912 gnd.n202 21.0318
R6770 gnd.n6907 gnd.n194 21.0318
R6771 gnd.n6964 gnd.n196 21.0318
R6772 gnd.n266 gnd.n186 21.0318
R6773 gnd.n6972 gnd.n188 21.0318
R6774 gnd.n1830 gnd.n1762 20.7615
R6775 gnd.n5424 gnd.n5423 20.7615
R6776 gnd.t189 gnd.n2297 20.7131
R6777 gnd.n6060 gnd.t15 20.7131
R6778 gnd.n4013 gnd.t212 20.7131
R6779 gnd.t172 gnd.n1184 20.7131
R6780 gnd.n6916 gnd.t264 20.7131
R6781 gnd.n2026 gnd.n1961 20.3945
R6782 gnd.n1126 gnd.n1118 20.3945
R6783 gnd.t163 gnd.n2332 20.0758
R6784 gnd.n6084 gnd.t233 20.0758
R6785 gnd.t148 gnd.n943 20.0758
R6786 gnd.t146 gnd.n5718 20.0758
R6787 gnd.n261 gnd.t140 20.0758
R6788 gnd.n1814 gnd.t117 19.8005
R6789 gnd.n1814 gnd.t33 19.8005
R6790 gnd.n1815 gnd.t26 19.8005
R6791 gnd.n1815 gnd.t54 19.8005
R6792 gnd.n5349 gnd.t75 19.8005
R6793 gnd.n5349 gnd.t40 19.8005
R6794 gnd.n5350 gnd.t91 19.8005
R6795 gnd.n5350 gnd.t19 19.8005
R6796 gnd.n1811 gnd.n1810 19.5087
R6797 gnd.n1824 gnd.n1811 19.5087
R6798 gnd.n1822 gnd.n1813 19.5087
R6799 gnd.n5354 gnd.n5348 19.5087
R6800 gnd.n3040 gnd.t142 19.4385
R6801 gnd.n6091 gnd.n6090 19.4385
R6802 gnd.n180 gnd.n168 19.4385
R6803 gnd.n4275 gnd.n4274 19.3944
R6804 gnd.n4274 gnd.n4273 19.3944
R6805 gnd.n4273 gnd.n4258 19.3944
R6806 gnd.n4269 gnd.n4258 19.3944
R6807 gnd.n4269 gnd.n4268 19.3944
R6808 gnd.n4268 gnd.n4267 19.3944
R6809 gnd.n4267 gnd.n1743 19.3944
R6810 gnd.n4480 gnd.n1743 19.3944
R6811 gnd.n4480 gnd.n1740 19.3944
R6812 gnd.n4498 gnd.n1740 19.3944
R6813 gnd.n4498 gnd.n1741 19.3944
R6814 gnd.n4494 gnd.n1741 19.3944
R6815 gnd.n4494 gnd.n4493 19.3944
R6816 gnd.n4493 gnd.n4492 19.3944
R6817 gnd.n4492 gnd.n4487 19.3944
R6818 gnd.n4488 gnd.n4487 19.3944
R6819 gnd.n4488 gnd.n1696 19.3944
R6820 gnd.n4567 gnd.n1696 19.3944
R6821 gnd.n4567 gnd.n1693 19.3944
R6822 gnd.n4578 gnd.n1693 19.3944
R6823 gnd.n4578 gnd.n1694 19.3944
R6824 gnd.n4574 gnd.n1694 19.3944
R6825 gnd.n4574 gnd.n4573 19.3944
R6826 gnd.n4573 gnd.n1653 19.3944
R6827 gnd.n4653 gnd.n1653 19.3944
R6828 gnd.n4653 gnd.n1650 19.3944
R6829 gnd.n4693 gnd.n1650 19.3944
R6830 gnd.n4693 gnd.n1651 19.3944
R6831 gnd.n4689 gnd.n1651 19.3944
R6832 gnd.n4689 gnd.n4688 19.3944
R6833 gnd.n4688 gnd.n4687 19.3944
R6834 gnd.n4687 gnd.n4660 19.3944
R6835 gnd.n4683 gnd.n4660 19.3944
R6836 gnd.n4683 gnd.n4682 19.3944
R6837 gnd.n4682 gnd.n4681 19.3944
R6838 gnd.n4681 gnd.n4665 19.3944
R6839 gnd.n4677 gnd.n4665 19.3944
R6840 gnd.n4677 gnd.n4676 19.3944
R6841 gnd.n4676 gnd.n4675 19.3944
R6842 gnd.n4675 gnd.n4672 19.3944
R6843 gnd.n4672 gnd.n1565 19.3944
R6844 gnd.n4830 gnd.n1565 19.3944
R6845 gnd.n4830 gnd.n1562 19.3944
R6846 gnd.n4847 gnd.n1562 19.3944
R6847 gnd.n4847 gnd.n1563 19.3944
R6848 gnd.n4843 gnd.n1563 19.3944
R6849 gnd.n4843 gnd.n4842 19.3944
R6850 gnd.n4842 gnd.n4841 19.3944
R6851 gnd.n4841 gnd.n4838 19.3944
R6852 gnd.n4838 gnd.n1515 19.3944
R6853 gnd.n4915 gnd.n1515 19.3944
R6854 gnd.n4915 gnd.n1512 19.3944
R6855 gnd.n4923 gnd.n1512 19.3944
R6856 gnd.n4923 gnd.n1513 19.3944
R6857 gnd.n4919 gnd.n1513 19.3944
R6858 gnd.n4919 gnd.n1485 19.3944
R6859 gnd.n4982 gnd.n1485 19.3944
R6860 gnd.n4982 gnd.n1482 19.3944
R6861 gnd.n5000 gnd.n1482 19.3944
R6862 gnd.n5000 gnd.n1483 19.3944
R6863 gnd.n4996 gnd.n1483 19.3944
R6864 gnd.n4996 gnd.n4995 19.3944
R6865 gnd.n4995 gnd.n4994 19.3944
R6866 gnd.n4994 gnd.n4991 19.3944
R6867 gnd.n4991 gnd.n1410 19.3944
R6868 gnd.n5067 gnd.n1410 19.3944
R6869 gnd.n5067 gnd.n1407 19.3944
R6870 gnd.n5072 gnd.n1407 19.3944
R6871 gnd.n5072 gnd.n1408 19.3944
R6872 gnd.n1408 gnd.n1381 19.3944
R6873 gnd.n5103 gnd.n1381 19.3944
R6874 gnd.n5103 gnd.n1379 19.3944
R6875 gnd.n5107 gnd.n1379 19.3944
R6876 gnd.n5107 gnd.n1359 19.3944
R6877 gnd.n5134 gnd.n1359 19.3944
R6878 gnd.n5134 gnd.n1357 19.3944
R6879 gnd.n5138 gnd.n1357 19.3944
R6880 gnd.n5138 gnd.n1355 19.3944
R6881 gnd.n5145 gnd.n1355 19.3944
R6882 gnd.n5145 gnd.n1352 19.3944
R6883 gnd.n5325 gnd.n1352 19.3944
R6884 gnd.n5325 gnd.n1353 19.3944
R6885 gnd.n4281 gnd.n4280 19.3944
R6886 gnd.n4280 gnd.n4279 19.3944
R6887 gnd.n4279 gnd.n2017 19.3944
R6888 gnd.n4241 gnd.n4240 19.3944
R6889 gnd.n4240 gnd.n4130 19.3944
R6890 gnd.n4233 gnd.n4130 19.3944
R6891 gnd.n4233 gnd.n4232 19.3944
R6892 gnd.n4232 gnd.n4146 19.3944
R6893 gnd.n4225 gnd.n4146 19.3944
R6894 gnd.n4225 gnd.n4224 19.3944
R6895 gnd.n4224 gnd.n4156 19.3944
R6896 gnd.n4217 gnd.n4156 19.3944
R6897 gnd.n4217 gnd.n4216 19.3944
R6898 gnd.n4216 gnd.n4169 19.3944
R6899 gnd.n4209 gnd.n4169 19.3944
R6900 gnd.n4209 gnd.n4208 19.3944
R6901 gnd.n4208 gnd.n4179 19.3944
R6902 gnd.n4201 gnd.n4179 19.3944
R6903 gnd.n4201 gnd.n4200 19.3944
R6904 gnd.n4200 gnd.n2001 19.3944
R6905 gnd.n4292 gnd.n2001 19.3944
R6906 gnd.n4292 gnd.n4291 19.3944
R6907 gnd.n4291 gnd.n4290 19.3944
R6908 gnd.n4290 gnd.n2005 19.3944
R6909 gnd.n4286 gnd.n2005 19.3944
R6910 gnd.n4286 gnd.n4285 19.3944
R6911 gnd.n4285 gnd.n4284 19.3944
R6912 gnd.n2755 gnd.n2754 19.3944
R6913 gnd.n2754 gnd.n2753 19.3944
R6914 gnd.n2753 gnd.n2752 19.3944
R6915 gnd.n2752 gnd.n2750 19.3944
R6916 gnd.n2750 gnd.n2747 19.3944
R6917 gnd.n2747 gnd.n2746 19.3944
R6918 gnd.n2746 gnd.n2743 19.3944
R6919 gnd.n2743 gnd.n2742 19.3944
R6920 gnd.n2742 gnd.n2739 19.3944
R6921 gnd.n2739 gnd.n2738 19.3944
R6922 gnd.n2738 gnd.n2735 19.3944
R6923 gnd.n2735 gnd.n2734 19.3944
R6924 gnd.n2734 gnd.n2731 19.3944
R6925 gnd.n2731 gnd.n2730 19.3944
R6926 gnd.n2730 gnd.n2727 19.3944
R6927 gnd.n2727 gnd.n2726 19.3944
R6928 gnd.n2726 gnd.n2723 19.3944
R6929 gnd.n2723 gnd.n2722 19.3944
R6930 gnd.n2722 gnd.n2719 19.3944
R6931 gnd.n2719 gnd.n2718 19.3944
R6932 gnd.n2718 gnd.n2715 19.3944
R6933 gnd.n2715 gnd.n2714 19.3944
R6934 gnd.n2711 gnd.n2710 19.3944
R6935 gnd.n2710 gnd.n2666 19.3944
R6936 gnd.n2761 gnd.n2666 19.3944
R6937 gnd.n3528 gnd.n3527 19.3944
R6938 gnd.n3527 gnd.n3524 19.3944
R6939 gnd.n3524 gnd.n3523 19.3944
R6940 gnd.n3573 gnd.n3572 19.3944
R6941 gnd.n3572 gnd.n3571 19.3944
R6942 gnd.n3571 gnd.n3568 19.3944
R6943 gnd.n3568 gnd.n3567 19.3944
R6944 gnd.n3567 gnd.n3564 19.3944
R6945 gnd.n3564 gnd.n3563 19.3944
R6946 gnd.n3563 gnd.n3560 19.3944
R6947 gnd.n3560 gnd.n3559 19.3944
R6948 gnd.n3559 gnd.n3556 19.3944
R6949 gnd.n3556 gnd.n3555 19.3944
R6950 gnd.n3555 gnd.n3552 19.3944
R6951 gnd.n3552 gnd.n3551 19.3944
R6952 gnd.n3551 gnd.n3548 19.3944
R6953 gnd.n3548 gnd.n3547 19.3944
R6954 gnd.n3547 gnd.n3544 19.3944
R6955 gnd.n3544 gnd.n3543 19.3944
R6956 gnd.n3543 gnd.n3540 19.3944
R6957 gnd.n3540 gnd.n3539 19.3944
R6958 gnd.n3539 gnd.n3536 19.3944
R6959 gnd.n3536 gnd.n3535 19.3944
R6960 gnd.n3535 gnd.n3532 19.3944
R6961 gnd.n3532 gnd.n3531 19.3944
R6962 gnd.n2854 gnd.n2563 19.3944
R6963 gnd.n2864 gnd.n2563 19.3944
R6964 gnd.n2865 gnd.n2864 19.3944
R6965 gnd.n2865 gnd.n2544 19.3944
R6966 gnd.n2885 gnd.n2544 19.3944
R6967 gnd.n2885 gnd.n2536 19.3944
R6968 gnd.n2895 gnd.n2536 19.3944
R6969 gnd.n2896 gnd.n2895 19.3944
R6970 gnd.n2897 gnd.n2896 19.3944
R6971 gnd.n2897 gnd.n2519 19.3944
R6972 gnd.n2914 gnd.n2519 19.3944
R6973 gnd.n2917 gnd.n2914 19.3944
R6974 gnd.n2917 gnd.n2916 19.3944
R6975 gnd.n2916 gnd.n2492 19.3944
R6976 gnd.n2956 gnd.n2492 19.3944
R6977 gnd.n2956 gnd.n2489 19.3944
R6978 gnd.n2962 gnd.n2489 19.3944
R6979 gnd.n2963 gnd.n2962 19.3944
R6980 gnd.n2963 gnd.n2487 19.3944
R6981 gnd.n2969 gnd.n2487 19.3944
R6982 gnd.n2972 gnd.n2969 19.3944
R6983 gnd.n2974 gnd.n2972 19.3944
R6984 gnd.n2980 gnd.n2974 19.3944
R6985 gnd.n2980 gnd.n2979 19.3944
R6986 gnd.n2979 gnd.n2374 19.3944
R6987 gnd.n3046 gnd.n2374 19.3944
R6988 gnd.n3047 gnd.n3046 19.3944
R6989 gnd.n3047 gnd.n2367 19.3944
R6990 gnd.n3058 gnd.n2367 19.3944
R6991 gnd.n3059 gnd.n3058 19.3944
R6992 gnd.n3059 gnd.n2350 19.3944
R6993 gnd.n2350 gnd.n2348 19.3944
R6994 gnd.n3083 gnd.n2348 19.3944
R6995 gnd.n3084 gnd.n3083 19.3944
R6996 gnd.n3084 gnd.n2319 19.3944
R6997 gnd.n3131 gnd.n2319 19.3944
R6998 gnd.n3132 gnd.n3131 19.3944
R6999 gnd.n3132 gnd.n2312 19.3944
R7000 gnd.n3144 gnd.n2312 19.3944
R7001 gnd.n3145 gnd.n3144 19.3944
R7002 gnd.n3145 gnd.n2295 19.3944
R7003 gnd.n2295 gnd.n2293 19.3944
R7004 gnd.n3169 gnd.n2293 19.3944
R7005 gnd.n3170 gnd.n3169 19.3944
R7006 gnd.n3170 gnd.n2265 19.3944
R7007 gnd.n3221 gnd.n2265 19.3944
R7008 gnd.n3222 gnd.n3221 19.3944
R7009 gnd.n3222 gnd.n2258 19.3944
R7010 gnd.n3489 gnd.n2258 19.3944
R7011 gnd.n3490 gnd.n3489 19.3944
R7012 gnd.n3490 gnd.n2239 19.3944
R7013 gnd.n3515 gnd.n2239 19.3944
R7014 gnd.n3515 gnd.n2240 19.3944
R7015 gnd.n2845 gnd.n2844 19.3944
R7016 gnd.n2844 gnd.n2577 19.3944
R7017 gnd.n2600 gnd.n2577 19.3944
R7018 gnd.n2603 gnd.n2600 19.3944
R7019 gnd.n2603 gnd.n2596 19.3944
R7020 gnd.n2607 gnd.n2596 19.3944
R7021 gnd.n2610 gnd.n2607 19.3944
R7022 gnd.n2613 gnd.n2610 19.3944
R7023 gnd.n2613 gnd.n2594 19.3944
R7024 gnd.n2617 gnd.n2594 19.3944
R7025 gnd.n2620 gnd.n2617 19.3944
R7026 gnd.n2623 gnd.n2620 19.3944
R7027 gnd.n2623 gnd.n2592 19.3944
R7028 gnd.n2627 gnd.n2592 19.3944
R7029 gnd.n2850 gnd.n2849 19.3944
R7030 gnd.n2849 gnd.n2553 19.3944
R7031 gnd.n2875 gnd.n2553 19.3944
R7032 gnd.n2875 gnd.n2551 19.3944
R7033 gnd.n2881 gnd.n2551 19.3944
R7034 gnd.n2881 gnd.n2880 19.3944
R7035 gnd.n2880 gnd.n2525 19.3944
R7036 gnd.n2905 gnd.n2525 19.3944
R7037 gnd.n2905 gnd.n2523 19.3944
R7038 gnd.n2909 gnd.n2523 19.3944
R7039 gnd.n2909 gnd.n2503 19.3944
R7040 gnd.n2936 gnd.n2503 19.3944
R7041 gnd.n2936 gnd.n2501 19.3944
R7042 gnd.n2946 gnd.n2501 19.3944
R7043 gnd.n2946 gnd.n2945 19.3944
R7044 gnd.n2945 gnd.n2944 19.3944
R7045 gnd.n2944 gnd.n2450 19.3944
R7046 gnd.n2994 gnd.n2450 19.3944
R7047 gnd.n2994 gnd.n2993 19.3944
R7048 gnd.n2993 gnd.n2992 19.3944
R7049 gnd.n2992 gnd.n2454 19.3944
R7050 gnd.n2474 gnd.n2454 19.3944
R7051 gnd.n2474 gnd.n2384 19.3944
R7052 gnd.n3031 gnd.n2384 19.3944
R7053 gnd.n3031 gnd.n2382 19.3944
R7054 gnd.n3037 gnd.n2382 19.3944
R7055 gnd.n3037 gnd.n3036 19.3944
R7056 gnd.n3036 gnd.n2357 19.3944
R7057 gnd.n3071 gnd.n2357 19.3944
R7058 gnd.n3071 gnd.n2355 19.3944
R7059 gnd.n3077 gnd.n2355 19.3944
R7060 gnd.n3077 gnd.n3076 19.3944
R7061 gnd.n3076 gnd.n2330 19.3944
R7062 gnd.n3116 gnd.n2330 19.3944
R7063 gnd.n3116 gnd.n2328 19.3944
R7064 gnd.n3122 gnd.n2328 19.3944
R7065 gnd.n3122 gnd.n3121 19.3944
R7066 gnd.n3121 gnd.n2302 19.3944
R7067 gnd.n3157 gnd.n2302 19.3944
R7068 gnd.n3157 gnd.n2300 19.3944
R7069 gnd.n3163 gnd.n2300 19.3944
R7070 gnd.n3163 gnd.n3162 19.3944
R7071 gnd.n3162 gnd.n2275 19.3944
R7072 gnd.n3206 gnd.n2275 19.3944
R7073 gnd.n3206 gnd.n2273 19.3944
R7074 gnd.n3212 gnd.n2273 19.3944
R7075 gnd.n3212 gnd.n3211 19.3944
R7076 gnd.n3211 gnd.n2248 19.3944
R7077 gnd.n3500 gnd.n2248 19.3944
R7078 gnd.n3500 gnd.n2246 19.3944
R7079 gnd.n3508 gnd.n2246 19.3944
R7080 gnd.n3508 gnd.n3507 19.3944
R7081 gnd.n3507 gnd.n3506 19.3944
R7082 gnd.n3609 gnd.n3608 19.3944
R7083 gnd.n3608 gnd.n2187 19.3944
R7084 gnd.n3604 gnd.n2187 19.3944
R7085 gnd.n3604 gnd.n3601 19.3944
R7086 gnd.n3601 gnd.n3598 19.3944
R7087 gnd.n3598 gnd.n3597 19.3944
R7088 gnd.n3597 gnd.n3594 19.3944
R7089 gnd.n3594 gnd.n3593 19.3944
R7090 gnd.n3593 gnd.n3590 19.3944
R7091 gnd.n3590 gnd.n3589 19.3944
R7092 gnd.n3589 gnd.n3586 19.3944
R7093 gnd.n3586 gnd.n3585 19.3944
R7094 gnd.n3585 gnd.n3582 19.3944
R7095 gnd.n3582 gnd.n3581 19.3944
R7096 gnd.n2765 gnd.n2664 19.3944
R7097 gnd.n2765 gnd.n2655 19.3944
R7098 gnd.n2778 gnd.n2655 19.3944
R7099 gnd.n2778 gnd.n2653 19.3944
R7100 gnd.n2782 gnd.n2653 19.3944
R7101 gnd.n2782 gnd.n2643 19.3944
R7102 gnd.n2794 gnd.n2643 19.3944
R7103 gnd.n2794 gnd.n2641 19.3944
R7104 gnd.n2828 gnd.n2641 19.3944
R7105 gnd.n2828 gnd.n2827 19.3944
R7106 gnd.n2827 gnd.n2826 19.3944
R7107 gnd.n2826 gnd.n2825 19.3944
R7108 gnd.n2825 gnd.n2822 19.3944
R7109 gnd.n2822 gnd.n2821 19.3944
R7110 gnd.n2821 gnd.n2820 19.3944
R7111 gnd.n2820 gnd.n2818 19.3944
R7112 gnd.n2818 gnd.n2817 19.3944
R7113 gnd.n2817 gnd.n2814 19.3944
R7114 gnd.n2814 gnd.n2813 19.3944
R7115 gnd.n2813 gnd.n2812 19.3944
R7116 gnd.n2812 gnd.n2810 19.3944
R7117 gnd.n2810 gnd.n2509 19.3944
R7118 gnd.n2925 gnd.n2509 19.3944
R7119 gnd.n2925 gnd.n2507 19.3944
R7120 gnd.n2931 gnd.n2507 19.3944
R7121 gnd.n2931 gnd.n2930 19.3944
R7122 gnd.n2930 gnd.n2431 19.3944
R7123 gnd.n3005 gnd.n2431 19.3944
R7124 gnd.n3005 gnd.n2432 19.3944
R7125 gnd.n2479 gnd.n2478 19.3944
R7126 gnd.n2482 gnd.n2481 19.3944
R7127 gnd.n2469 gnd.n2468 19.3944
R7128 gnd.n3024 gnd.n2389 19.3944
R7129 gnd.n3024 gnd.n3023 19.3944
R7130 gnd.n3023 gnd.n3022 19.3944
R7131 gnd.n3022 gnd.n3020 19.3944
R7132 gnd.n3020 gnd.n3019 19.3944
R7133 gnd.n3019 gnd.n3017 19.3944
R7134 gnd.n3017 gnd.n3016 19.3944
R7135 gnd.n3016 gnd.n2338 19.3944
R7136 gnd.n3092 gnd.n2338 19.3944
R7137 gnd.n3092 gnd.n2336 19.3944
R7138 gnd.n3111 gnd.n2336 19.3944
R7139 gnd.n3111 gnd.n3110 19.3944
R7140 gnd.n3110 gnd.n3109 19.3944
R7141 gnd.n3109 gnd.n3107 19.3944
R7142 gnd.n3107 gnd.n3106 19.3944
R7143 gnd.n3106 gnd.n3104 19.3944
R7144 gnd.n3104 gnd.n3103 19.3944
R7145 gnd.n3103 gnd.n2282 19.3944
R7146 gnd.n3178 gnd.n2282 19.3944
R7147 gnd.n3178 gnd.n2280 19.3944
R7148 gnd.n3201 gnd.n2280 19.3944
R7149 gnd.n3201 gnd.n3200 19.3944
R7150 gnd.n3200 gnd.n3199 19.3944
R7151 gnd.n3199 gnd.n3196 19.3944
R7152 gnd.n3196 gnd.n3195 19.3944
R7153 gnd.n3195 gnd.n3193 19.3944
R7154 gnd.n3193 gnd.n3192 19.3944
R7155 gnd.n3192 gnd.n3190 19.3944
R7156 gnd.n3190 gnd.n2234 19.3944
R7157 gnd.n2770 gnd.n2660 19.3944
R7158 gnd.n2770 gnd.n2658 19.3944
R7159 gnd.n2774 gnd.n2658 19.3944
R7160 gnd.n2774 gnd.n2649 19.3944
R7161 gnd.n2786 gnd.n2649 19.3944
R7162 gnd.n2786 gnd.n2647 19.3944
R7163 gnd.n2790 gnd.n2647 19.3944
R7164 gnd.n2790 gnd.n2636 19.3944
R7165 gnd.n2832 gnd.n2636 19.3944
R7166 gnd.n2832 gnd.n2590 19.3944
R7167 gnd.n2838 gnd.n2590 19.3944
R7168 gnd.n2838 gnd.n2837 19.3944
R7169 gnd.n2837 gnd.n2568 19.3944
R7170 gnd.n2859 gnd.n2568 19.3944
R7171 gnd.n2859 gnd.n2561 19.3944
R7172 gnd.n2870 gnd.n2561 19.3944
R7173 gnd.n2870 gnd.n2869 19.3944
R7174 gnd.n2869 gnd.n2542 19.3944
R7175 gnd.n2890 gnd.n2542 19.3944
R7176 gnd.n2890 gnd.n2532 19.3944
R7177 gnd.n2900 gnd.n2532 19.3944
R7178 gnd.n2900 gnd.n2515 19.3944
R7179 gnd.n2921 gnd.n2515 19.3944
R7180 gnd.n2921 gnd.n2920 19.3944
R7181 gnd.n2920 gnd.n2494 19.3944
R7182 gnd.n2951 gnd.n2494 19.3944
R7183 gnd.n2951 gnd.n2439 19.3944
R7184 gnd.n3001 gnd.n2439 19.3944
R7185 gnd.n3001 gnd.n3000 19.3944
R7186 gnd.n3000 gnd.n2999 19.3944
R7187 gnd.n2999 gnd.n2443 19.3944
R7188 gnd.n2461 gnd.n2443 19.3944
R7189 gnd.n2987 gnd.n2461 19.3944
R7190 gnd.n2987 gnd.n2986 19.3944
R7191 gnd.n2986 gnd.n2985 19.3944
R7192 gnd.n2985 gnd.n2465 19.3944
R7193 gnd.n2465 gnd.n2376 19.3944
R7194 gnd.n3042 gnd.n2376 19.3944
R7195 gnd.n3042 gnd.n2369 19.3944
R7196 gnd.n3053 gnd.n2369 19.3944
R7197 gnd.n3053 gnd.n2365 19.3944
R7198 gnd.n3066 gnd.n2365 19.3944
R7199 gnd.n3066 gnd.n3065 19.3944
R7200 gnd.n3065 gnd.n2344 19.3944
R7201 gnd.n3088 gnd.n2344 19.3944
R7202 gnd.n3088 gnd.n3087 19.3944
R7203 gnd.n3087 gnd.n2321 19.3944
R7204 gnd.n3127 gnd.n2321 19.3944
R7205 gnd.n3127 gnd.n2314 19.3944
R7206 gnd.n3139 gnd.n2314 19.3944
R7207 gnd.n3139 gnd.n2310 19.3944
R7208 gnd.n3152 gnd.n2310 19.3944
R7209 gnd.n3152 gnd.n3151 19.3944
R7210 gnd.n3151 gnd.n2289 19.3944
R7211 gnd.n3174 gnd.n2289 19.3944
R7212 gnd.n3174 gnd.n3173 19.3944
R7213 gnd.n3173 gnd.n2267 19.3944
R7214 gnd.n3217 gnd.n2267 19.3944
R7215 gnd.n3217 gnd.n2260 19.3944
R7216 gnd.n3228 gnd.n2260 19.3944
R7217 gnd.n3228 gnd.n2256 19.3944
R7218 gnd.n3495 gnd.n2256 19.3944
R7219 gnd.n3495 gnd.n3494 19.3944
R7220 gnd.n3494 gnd.n2237 19.3944
R7221 gnd.n3518 gnd.n2237 19.3944
R7222 gnd.n5614 gnd.n1265 19.3944
R7223 gnd.n5614 gnd.n1262 19.3944
R7224 gnd.n5619 gnd.n1262 19.3944
R7225 gnd.n5619 gnd.n1263 19.3944
R7226 gnd.n1263 gnd.n1247 19.3944
R7227 gnd.n5700 gnd.n1247 19.3944
R7228 gnd.n5700 gnd.n1244 19.3944
R7229 gnd.n5705 gnd.n1244 19.3944
R7230 gnd.n5705 gnd.n1245 19.3944
R7231 gnd.n1245 gnd.n1218 19.3944
R7232 gnd.n5732 gnd.n1218 19.3944
R7233 gnd.n5732 gnd.n1215 19.3944
R7234 gnd.n5737 gnd.n1215 19.3944
R7235 gnd.n5737 gnd.n1216 19.3944
R7236 gnd.n1216 gnd.n1192 19.3944
R7237 gnd.n5765 gnd.n1192 19.3944
R7238 gnd.n5765 gnd.n1188 19.3944
R7239 gnd.n5770 gnd.n1188 19.3944
R7240 gnd.n5770 gnd.n1190 19.3944
R7241 gnd.n1190 gnd.n1189 19.3944
R7242 gnd.n1189 gnd.n52 19.3944
R7243 gnd.n7182 gnd.n52 19.3944
R7244 gnd.n7182 gnd.n7181 19.3944
R7245 gnd.n7181 gnd.n7180 19.3944
R7246 gnd.n7180 gnd.n57 19.3944
R7247 gnd.n7176 gnd.n57 19.3944
R7248 gnd.n7176 gnd.n7175 19.3944
R7249 gnd.n7175 gnd.n7174 19.3944
R7250 gnd.n7174 gnd.n62 19.3944
R7251 gnd.n7170 gnd.n62 19.3944
R7252 gnd.n7170 gnd.n7169 19.3944
R7253 gnd.n7169 gnd.n7168 19.3944
R7254 gnd.n7168 gnd.n67 19.3944
R7255 gnd.n7164 gnd.n67 19.3944
R7256 gnd.n7164 gnd.n7163 19.3944
R7257 gnd.n7163 gnd.n7162 19.3944
R7258 gnd.n7162 gnd.n72 19.3944
R7259 gnd.n7158 gnd.n72 19.3944
R7260 gnd.n7158 gnd.n7157 19.3944
R7261 gnd.n7157 gnd.n7156 19.3944
R7262 gnd.n7156 gnd.n77 19.3944
R7263 gnd.n7152 gnd.n77 19.3944
R7264 gnd.n7051 gnd.n7050 19.3944
R7265 gnd.n7050 gnd.n7049 19.3944
R7266 gnd.n7049 gnd.n6992 19.3944
R7267 gnd.n7045 gnd.n6992 19.3944
R7268 gnd.n7045 gnd.n7044 19.3944
R7269 gnd.n7044 gnd.n7043 19.3944
R7270 gnd.n7043 gnd.n7000 19.3944
R7271 gnd.n7039 gnd.n7000 19.3944
R7272 gnd.n7039 gnd.n7038 19.3944
R7273 gnd.n7038 gnd.n7037 19.3944
R7274 gnd.n7037 gnd.n7008 19.3944
R7275 gnd.n7033 gnd.n7008 19.3944
R7276 gnd.n7033 gnd.n7032 19.3944
R7277 gnd.n7032 gnd.n7031 19.3944
R7278 gnd.n7031 gnd.n7016 19.3944
R7279 gnd.n7027 gnd.n7016 19.3944
R7280 gnd.n5205 gnd.n5199 19.3944
R7281 gnd.n5211 gnd.n5199 19.3944
R7282 gnd.n5211 gnd.n5192 19.3944
R7283 gnd.n5224 gnd.n5192 19.3944
R7284 gnd.n5224 gnd.n5190 19.3944
R7285 gnd.n5230 gnd.n5190 19.3944
R7286 gnd.n5230 gnd.n5183 19.3944
R7287 gnd.n5243 gnd.n5183 19.3944
R7288 gnd.n5243 gnd.n5181 19.3944
R7289 gnd.n5249 gnd.n5181 19.3944
R7290 gnd.n5249 gnd.n5174 19.3944
R7291 gnd.n5262 gnd.n5174 19.3944
R7292 gnd.n5262 gnd.n5172 19.3944
R7293 gnd.n5268 gnd.n5172 19.3944
R7294 gnd.n5268 gnd.n5165 19.3944
R7295 gnd.n5283 gnd.n5165 19.3944
R7296 gnd.n5202 gnd.n1144 19.3944
R7297 gnd.n5843 gnd.n1144 19.3944
R7298 gnd.n5843 gnd.n1145 19.3944
R7299 gnd.n5839 gnd.n1145 19.3944
R7300 gnd.n5839 gnd.n5838 19.3944
R7301 gnd.n5838 gnd.n5837 19.3944
R7302 gnd.n5837 gnd.n1151 19.3944
R7303 gnd.n5833 gnd.n1151 19.3944
R7304 gnd.n5833 gnd.n5832 19.3944
R7305 gnd.n5832 gnd.n5831 19.3944
R7306 gnd.n5831 gnd.n1156 19.3944
R7307 gnd.n5827 gnd.n1156 19.3944
R7308 gnd.n5827 gnd.n5826 19.3944
R7309 gnd.n5826 gnd.n5825 19.3944
R7310 gnd.n5825 gnd.n1161 19.3944
R7311 gnd.n5821 gnd.n1161 19.3944
R7312 gnd.n5821 gnd.n5820 19.3944
R7313 gnd.n5820 gnd.n5819 19.3944
R7314 gnd.n5819 gnd.n1166 19.3944
R7315 gnd.n5815 gnd.n1166 19.3944
R7316 gnd.n5815 gnd.n5814 19.3944
R7317 gnd.n5814 gnd.n5813 19.3944
R7318 gnd.n5813 gnd.n229 19.3944
R7319 gnd.n6934 gnd.n229 19.3944
R7320 gnd.n6934 gnd.n227 19.3944
R7321 gnd.n6938 gnd.n227 19.3944
R7322 gnd.n6938 gnd.n207 19.3944
R7323 gnd.n6950 gnd.n207 19.3944
R7324 gnd.n6950 gnd.n205 19.3944
R7325 gnd.n6954 gnd.n205 19.3944
R7326 gnd.n6954 gnd.n192 19.3944
R7327 gnd.n6966 gnd.n192 19.3944
R7328 gnd.n6966 gnd.n190 19.3944
R7329 gnd.n6970 gnd.n190 19.3944
R7330 gnd.n6970 gnd.n175 19.3944
R7331 gnd.n6982 gnd.n175 19.3944
R7332 gnd.n6982 gnd.n172 19.3944
R7333 gnd.n7060 gnd.n172 19.3944
R7334 gnd.n7060 gnd.n173 19.3944
R7335 gnd.n7056 gnd.n173 19.3944
R7336 gnd.n7056 gnd.n7055 19.3944
R7337 gnd.n7055 gnd.n7054 19.3944
R7338 gnd.n4134 gnd.n999 19.3944
R7339 gnd.n4134 gnd.n4133 19.3944
R7340 gnd.n4237 gnd.n4133 19.3944
R7341 gnd.n4237 gnd.n4236 19.3944
R7342 gnd.n4236 gnd.n4141 19.3944
R7343 gnd.n4229 gnd.n4141 19.3944
R7344 gnd.n4229 gnd.n4228 19.3944
R7345 gnd.n4228 gnd.n4152 19.3944
R7346 gnd.n4221 gnd.n4152 19.3944
R7347 gnd.n4221 gnd.n4220 19.3944
R7348 gnd.n4220 gnd.n4163 19.3944
R7349 gnd.n4213 gnd.n4163 19.3944
R7350 gnd.n4213 gnd.n4212 19.3944
R7351 gnd.n4212 gnd.n4175 19.3944
R7352 gnd.n4205 gnd.n4175 19.3944
R7353 gnd.n4205 gnd.n4204 19.3944
R7354 gnd.n6685 gnd.n405 19.3944
R7355 gnd.n6685 gnd.n401 19.3944
R7356 gnd.n6691 gnd.n401 19.3944
R7357 gnd.n6691 gnd.n399 19.3944
R7358 gnd.n6695 gnd.n399 19.3944
R7359 gnd.n6695 gnd.n395 19.3944
R7360 gnd.n6701 gnd.n395 19.3944
R7361 gnd.n6701 gnd.n393 19.3944
R7362 gnd.n6705 gnd.n393 19.3944
R7363 gnd.n6705 gnd.n389 19.3944
R7364 gnd.n6711 gnd.n389 19.3944
R7365 gnd.n6711 gnd.n387 19.3944
R7366 gnd.n6715 gnd.n387 19.3944
R7367 gnd.n6715 gnd.n383 19.3944
R7368 gnd.n6721 gnd.n383 19.3944
R7369 gnd.n6721 gnd.n381 19.3944
R7370 gnd.n6725 gnd.n381 19.3944
R7371 gnd.n6725 gnd.n377 19.3944
R7372 gnd.n6731 gnd.n377 19.3944
R7373 gnd.n6731 gnd.n375 19.3944
R7374 gnd.n6735 gnd.n375 19.3944
R7375 gnd.n6735 gnd.n371 19.3944
R7376 gnd.n6741 gnd.n371 19.3944
R7377 gnd.n6741 gnd.n369 19.3944
R7378 gnd.n6745 gnd.n369 19.3944
R7379 gnd.n6745 gnd.n365 19.3944
R7380 gnd.n6751 gnd.n365 19.3944
R7381 gnd.n6751 gnd.n363 19.3944
R7382 gnd.n6755 gnd.n363 19.3944
R7383 gnd.n6755 gnd.n359 19.3944
R7384 gnd.n6761 gnd.n359 19.3944
R7385 gnd.n6761 gnd.n357 19.3944
R7386 gnd.n6765 gnd.n357 19.3944
R7387 gnd.n6765 gnd.n353 19.3944
R7388 gnd.n6771 gnd.n353 19.3944
R7389 gnd.n6771 gnd.n351 19.3944
R7390 gnd.n6775 gnd.n351 19.3944
R7391 gnd.n6775 gnd.n347 19.3944
R7392 gnd.n6781 gnd.n347 19.3944
R7393 gnd.n6781 gnd.n345 19.3944
R7394 gnd.n6785 gnd.n345 19.3944
R7395 gnd.n6785 gnd.n341 19.3944
R7396 gnd.n6791 gnd.n341 19.3944
R7397 gnd.n6791 gnd.n339 19.3944
R7398 gnd.n6795 gnd.n339 19.3944
R7399 gnd.n6795 gnd.n335 19.3944
R7400 gnd.n6801 gnd.n335 19.3944
R7401 gnd.n6801 gnd.n333 19.3944
R7402 gnd.n6805 gnd.n333 19.3944
R7403 gnd.n6805 gnd.n329 19.3944
R7404 gnd.n6811 gnd.n329 19.3944
R7405 gnd.n6811 gnd.n327 19.3944
R7406 gnd.n6815 gnd.n327 19.3944
R7407 gnd.n6815 gnd.n323 19.3944
R7408 gnd.n6821 gnd.n323 19.3944
R7409 gnd.n6821 gnd.n321 19.3944
R7410 gnd.n6825 gnd.n321 19.3944
R7411 gnd.n6825 gnd.n317 19.3944
R7412 gnd.n6831 gnd.n317 19.3944
R7413 gnd.n6831 gnd.n315 19.3944
R7414 gnd.n6835 gnd.n315 19.3944
R7415 gnd.n6835 gnd.n311 19.3944
R7416 gnd.n6841 gnd.n311 19.3944
R7417 gnd.n6841 gnd.n309 19.3944
R7418 gnd.n6845 gnd.n309 19.3944
R7419 gnd.n6845 gnd.n305 19.3944
R7420 gnd.n6851 gnd.n305 19.3944
R7421 gnd.n6851 gnd.n303 19.3944
R7422 gnd.n6855 gnd.n303 19.3944
R7423 gnd.n6855 gnd.n299 19.3944
R7424 gnd.n6861 gnd.n299 19.3944
R7425 gnd.n6861 gnd.n297 19.3944
R7426 gnd.n6865 gnd.n297 19.3944
R7427 gnd.n6865 gnd.n293 19.3944
R7428 gnd.n6871 gnd.n293 19.3944
R7429 gnd.n6871 gnd.n291 19.3944
R7430 gnd.n6875 gnd.n291 19.3944
R7431 gnd.n6875 gnd.n287 19.3944
R7432 gnd.n6881 gnd.n287 19.3944
R7433 gnd.n6881 gnd.n285 19.3944
R7434 gnd.n6887 gnd.n285 19.3944
R7435 gnd.n6887 gnd.n6886 19.3944
R7436 gnd.n6886 gnd.n281 19.3944
R7437 gnd.n6894 gnd.n281 19.3944
R7438 gnd.n6265 gnd.n657 19.3944
R7439 gnd.n6265 gnd.n653 19.3944
R7440 gnd.n6271 gnd.n653 19.3944
R7441 gnd.n6271 gnd.n651 19.3944
R7442 gnd.n6275 gnd.n651 19.3944
R7443 gnd.n6275 gnd.n647 19.3944
R7444 gnd.n6281 gnd.n647 19.3944
R7445 gnd.n6281 gnd.n645 19.3944
R7446 gnd.n6285 gnd.n645 19.3944
R7447 gnd.n6285 gnd.n641 19.3944
R7448 gnd.n6291 gnd.n641 19.3944
R7449 gnd.n6291 gnd.n639 19.3944
R7450 gnd.n6295 gnd.n639 19.3944
R7451 gnd.n6295 gnd.n635 19.3944
R7452 gnd.n6301 gnd.n635 19.3944
R7453 gnd.n6301 gnd.n633 19.3944
R7454 gnd.n6305 gnd.n633 19.3944
R7455 gnd.n6305 gnd.n629 19.3944
R7456 gnd.n6311 gnd.n629 19.3944
R7457 gnd.n6311 gnd.n627 19.3944
R7458 gnd.n6315 gnd.n627 19.3944
R7459 gnd.n6315 gnd.n623 19.3944
R7460 gnd.n6321 gnd.n623 19.3944
R7461 gnd.n6321 gnd.n621 19.3944
R7462 gnd.n6325 gnd.n621 19.3944
R7463 gnd.n6325 gnd.n617 19.3944
R7464 gnd.n6331 gnd.n617 19.3944
R7465 gnd.n6331 gnd.n615 19.3944
R7466 gnd.n6335 gnd.n615 19.3944
R7467 gnd.n6335 gnd.n611 19.3944
R7468 gnd.n6341 gnd.n611 19.3944
R7469 gnd.n6341 gnd.n609 19.3944
R7470 gnd.n6345 gnd.n609 19.3944
R7471 gnd.n6345 gnd.n605 19.3944
R7472 gnd.n6351 gnd.n605 19.3944
R7473 gnd.n6351 gnd.n603 19.3944
R7474 gnd.n6355 gnd.n603 19.3944
R7475 gnd.n6355 gnd.n599 19.3944
R7476 gnd.n6361 gnd.n599 19.3944
R7477 gnd.n6361 gnd.n597 19.3944
R7478 gnd.n6365 gnd.n597 19.3944
R7479 gnd.n6365 gnd.n593 19.3944
R7480 gnd.n6371 gnd.n593 19.3944
R7481 gnd.n6371 gnd.n591 19.3944
R7482 gnd.n6375 gnd.n591 19.3944
R7483 gnd.n6375 gnd.n587 19.3944
R7484 gnd.n6381 gnd.n587 19.3944
R7485 gnd.n6381 gnd.n585 19.3944
R7486 gnd.n6385 gnd.n585 19.3944
R7487 gnd.n6385 gnd.n581 19.3944
R7488 gnd.n6391 gnd.n581 19.3944
R7489 gnd.n6391 gnd.n579 19.3944
R7490 gnd.n6395 gnd.n579 19.3944
R7491 gnd.n6395 gnd.n575 19.3944
R7492 gnd.n6401 gnd.n575 19.3944
R7493 gnd.n6401 gnd.n573 19.3944
R7494 gnd.n6405 gnd.n573 19.3944
R7495 gnd.n6405 gnd.n569 19.3944
R7496 gnd.n6411 gnd.n569 19.3944
R7497 gnd.n6411 gnd.n567 19.3944
R7498 gnd.n6415 gnd.n567 19.3944
R7499 gnd.n6415 gnd.n563 19.3944
R7500 gnd.n6421 gnd.n563 19.3944
R7501 gnd.n6421 gnd.n561 19.3944
R7502 gnd.n6425 gnd.n561 19.3944
R7503 gnd.n6425 gnd.n557 19.3944
R7504 gnd.n6431 gnd.n557 19.3944
R7505 gnd.n6431 gnd.n555 19.3944
R7506 gnd.n6435 gnd.n555 19.3944
R7507 gnd.n6435 gnd.n551 19.3944
R7508 gnd.n6441 gnd.n551 19.3944
R7509 gnd.n6441 gnd.n549 19.3944
R7510 gnd.n6445 gnd.n549 19.3944
R7511 gnd.n6445 gnd.n545 19.3944
R7512 gnd.n6451 gnd.n545 19.3944
R7513 gnd.n6451 gnd.n543 19.3944
R7514 gnd.n6455 gnd.n543 19.3944
R7515 gnd.n6455 gnd.n539 19.3944
R7516 gnd.n6461 gnd.n539 19.3944
R7517 gnd.n6461 gnd.n537 19.3944
R7518 gnd.n6465 gnd.n537 19.3944
R7519 gnd.n6465 gnd.n533 19.3944
R7520 gnd.n6471 gnd.n533 19.3944
R7521 gnd.n6471 gnd.n531 19.3944
R7522 gnd.n6475 gnd.n531 19.3944
R7523 gnd.n6475 gnd.n527 19.3944
R7524 gnd.n6481 gnd.n527 19.3944
R7525 gnd.n6481 gnd.n525 19.3944
R7526 gnd.n6485 gnd.n525 19.3944
R7527 gnd.n6485 gnd.n521 19.3944
R7528 gnd.n6491 gnd.n521 19.3944
R7529 gnd.n6491 gnd.n519 19.3944
R7530 gnd.n6495 gnd.n519 19.3944
R7531 gnd.n6495 gnd.n515 19.3944
R7532 gnd.n6501 gnd.n515 19.3944
R7533 gnd.n6501 gnd.n513 19.3944
R7534 gnd.n6505 gnd.n513 19.3944
R7535 gnd.n6505 gnd.n509 19.3944
R7536 gnd.n6511 gnd.n509 19.3944
R7537 gnd.n6511 gnd.n507 19.3944
R7538 gnd.n6515 gnd.n507 19.3944
R7539 gnd.n6515 gnd.n503 19.3944
R7540 gnd.n6521 gnd.n503 19.3944
R7541 gnd.n6521 gnd.n501 19.3944
R7542 gnd.n6525 gnd.n501 19.3944
R7543 gnd.n6525 gnd.n497 19.3944
R7544 gnd.n6531 gnd.n497 19.3944
R7545 gnd.n6531 gnd.n495 19.3944
R7546 gnd.n6535 gnd.n495 19.3944
R7547 gnd.n6535 gnd.n491 19.3944
R7548 gnd.n6541 gnd.n491 19.3944
R7549 gnd.n6541 gnd.n489 19.3944
R7550 gnd.n6545 gnd.n489 19.3944
R7551 gnd.n6545 gnd.n485 19.3944
R7552 gnd.n6551 gnd.n485 19.3944
R7553 gnd.n6551 gnd.n483 19.3944
R7554 gnd.n6555 gnd.n483 19.3944
R7555 gnd.n6555 gnd.n479 19.3944
R7556 gnd.n6561 gnd.n479 19.3944
R7557 gnd.n6561 gnd.n477 19.3944
R7558 gnd.n6565 gnd.n477 19.3944
R7559 gnd.n6565 gnd.n473 19.3944
R7560 gnd.n6571 gnd.n473 19.3944
R7561 gnd.n6571 gnd.n471 19.3944
R7562 gnd.n6575 gnd.n471 19.3944
R7563 gnd.n6575 gnd.n467 19.3944
R7564 gnd.n6581 gnd.n467 19.3944
R7565 gnd.n6581 gnd.n465 19.3944
R7566 gnd.n6585 gnd.n465 19.3944
R7567 gnd.n6585 gnd.n461 19.3944
R7568 gnd.n6591 gnd.n461 19.3944
R7569 gnd.n6591 gnd.n459 19.3944
R7570 gnd.n6595 gnd.n459 19.3944
R7571 gnd.n6595 gnd.n455 19.3944
R7572 gnd.n6601 gnd.n455 19.3944
R7573 gnd.n6601 gnd.n453 19.3944
R7574 gnd.n6605 gnd.n453 19.3944
R7575 gnd.n6605 gnd.n449 19.3944
R7576 gnd.n6611 gnd.n449 19.3944
R7577 gnd.n6611 gnd.n447 19.3944
R7578 gnd.n6615 gnd.n447 19.3944
R7579 gnd.n6615 gnd.n443 19.3944
R7580 gnd.n6621 gnd.n443 19.3944
R7581 gnd.n6621 gnd.n441 19.3944
R7582 gnd.n6625 gnd.n441 19.3944
R7583 gnd.n6625 gnd.n437 19.3944
R7584 gnd.n6631 gnd.n437 19.3944
R7585 gnd.n6631 gnd.n435 19.3944
R7586 gnd.n6635 gnd.n435 19.3944
R7587 gnd.n6635 gnd.n431 19.3944
R7588 gnd.n6641 gnd.n431 19.3944
R7589 gnd.n6641 gnd.n429 19.3944
R7590 gnd.n6645 gnd.n429 19.3944
R7591 gnd.n6645 gnd.n425 19.3944
R7592 gnd.n6651 gnd.n425 19.3944
R7593 gnd.n6651 gnd.n423 19.3944
R7594 gnd.n6655 gnd.n423 19.3944
R7595 gnd.n6655 gnd.n419 19.3944
R7596 gnd.n6661 gnd.n419 19.3944
R7597 gnd.n6661 gnd.n417 19.3944
R7598 gnd.n6665 gnd.n417 19.3944
R7599 gnd.n6665 gnd.n413 19.3944
R7600 gnd.n6671 gnd.n413 19.3944
R7601 gnd.n6671 gnd.n411 19.3944
R7602 gnd.n6675 gnd.n411 19.3944
R7603 gnd.n6675 gnd.n407 19.3944
R7604 gnd.n6681 gnd.n407 19.3944
R7605 gnd.n5514 gnd.n5511 19.3944
R7606 gnd.n5514 gnd.n5510 19.3944
R7607 gnd.n5520 gnd.n5510 19.3944
R7608 gnd.n5520 gnd.n5508 19.3944
R7609 gnd.n5524 gnd.n5508 19.3944
R7610 gnd.n5524 gnd.n5506 19.3944
R7611 gnd.n5530 gnd.n5506 19.3944
R7612 gnd.n5530 gnd.n5504 19.3944
R7613 gnd.n5534 gnd.n5504 19.3944
R7614 gnd.n5534 gnd.n5502 19.3944
R7615 gnd.n5540 gnd.n5502 19.3944
R7616 gnd.n5540 gnd.n5500 19.3944
R7617 gnd.n5545 gnd.n5500 19.3944
R7618 gnd.n5545 gnd.n5498 19.3944
R7619 gnd.n5498 gnd.n1291 19.3944
R7620 gnd.n5558 gnd.n1289 19.3944
R7621 gnd.n5558 gnd.n1287 19.3944
R7622 gnd.n5564 gnd.n1287 19.3944
R7623 gnd.n5564 gnd.n1285 19.3944
R7624 gnd.n5568 gnd.n1285 19.3944
R7625 gnd.n5568 gnd.n1283 19.3944
R7626 gnd.n5574 gnd.n1283 19.3944
R7627 gnd.n5574 gnd.n1281 19.3944
R7628 gnd.n5578 gnd.n1281 19.3944
R7629 gnd.n5578 gnd.n1279 19.3944
R7630 gnd.n5584 gnd.n1279 19.3944
R7631 gnd.n5584 gnd.n1277 19.3944
R7632 gnd.n5588 gnd.n1277 19.3944
R7633 gnd.n5588 gnd.n1275 19.3944
R7634 gnd.n5594 gnd.n1275 19.3944
R7635 gnd.n5594 gnd.n1273 19.3944
R7636 gnd.n5599 gnd.n1273 19.3944
R7637 gnd.n5599 gnd.n1271 19.3944
R7638 gnd.n5610 gnd.n1266 19.3944
R7639 gnd.n5610 gnd.n1261 19.3944
R7640 gnd.n5623 gnd.n1261 19.3944
R7641 gnd.n5623 gnd.n1259 19.3944
R7642 gnd.n5668 gnd.n1259 19.3944
R7643 gnd.n5668 gnd.n5667 19.3944
R7644 gnd.n5667 gnd.n5666 19.3944
R7645 gnd.n5666 gnd.n5664 19.3944
R7646 gnd.n5664 gnd.n5663 19.3944
R7647 gnd.n5663 gnd.n5662 19.3944
R7648 gnd.n5662 gnd.n5660 19.3944
R7649 gnd.n5660 gnd.n5659 19.3944
R7650 gnd.n5659 gnd.n5657 19.3944
R7651 gnd.n5657 gnd.n5656 19.3944
R7652 gnd.n5656 gnd.n5655 19.3944
R7653 gnd.n5655 gnd.n5653 19.3944
R7654 gnd.n5653 gnd.n5652 19.3944
R7655 gnd.n5652 gnd.n5649 19.3944
R7656 gnd.n5649 gnd.n5648 19.3944
R7657 gnd.n5648 gnd.n5646 19.3944
R7658 gnd.n5646 gnd.n5645 19.3944
R7659 gnd.n5645 gnd.n237 19.3944
R7660 gnd.n6925 gnd.n237 19.3944
R7661 gnd.n6925 gnd.n6924 19.3944
R7662 gnd.n6924 gnd.n6923 19.3944
R7663 gnd.n6923 gnd.n6919 19.3944
R7664 gnd.n6919 gnd.n6918 19.3944
R7665 gnd.n6918 gnd.n6915 19.3944
R7666 gnd.n6915 gnd.n6914 19.3944
R7667 gnd.n6914 gnd.n6910 19.3944
R7668 gnd.n6910 gnd.n6909 19.3944
R7669 gnd.n6909 gnd.n269 19.3944
R7670 gnd.n269 gnd.n268 19.3944
R7671 gnd.n268 gnd.n264 19.3944
R7672 gnd.n264 gnd.n263 19.3944
R7673 gnd.n263 gnd.n260 19.3944
R7674 gnd.n260 gnd.n259 19.3944
R7675 gnd.n259 gnd.n257 19.3944
R7676 gnd.n257 gnd.n256 19.3944
R7677 gnd.n256 gnd.n159 19.3944
R7678 gnd.n7073 gnd.n159 19.3944
R7679 gnd.n7074 gnd.n7073 19.3944
R7680 gnd.n7112 gnd.n120 19.3944
R7681 gnd.n7107 gnd.n120 19.3944
R7682 gnd.n7107 gnd.n7106 19.3944
R7683 gnd.n7106 gnd.n7105 19.3944
R7684 gnd.n7105 gnd.n127 19.3944
R7685 gnd.n7100 gnd.n127 19.3944
R7686 gnd.n7100 gnd.n7099 19.3944
R7687 gnd.n7099 gnd.n7098 19.3944
R7688 gnd.n7098 gnd.n134 19.3944
R7689 gnd.n7093 gnd.n134 19.3944
R7690 gnd.n7093 gnd.n7092 19.3944
R7691 gnd.n7092 gnd.n7091 19.3944
R7692 gnd.n7091 gnd.n141 19.3944
R7693 gnd.n7086 gnd.n141 19.3944
R7694 gnd.n7086 gnd.n7085 19.3944
R7695 gnd.n7085 gnd.n7084 19.3944
R7696 gnd.n7084 gnd.n148 19.3944
R7697 gnd.n7079 gnd.n148 19.3944
R7698 gnd.n7145 gnd.n7144 19.3944
R7699 gnd.n7144 gnd.n7143 19.3944
R7700 gnd.n7143 gnd.n92 19.3944
R7701 gnd.n7138 gnd.n92 19.3944
R7702 gnd.n7138 gnd.n7137 19.3944
R7703 gnd.n7137 gnd.n7136 19.3944
R7704 gnd.n7136 gnd.n99 19.3944
R7705 gnd.n7131 gnd.n99 19.3944
R7706 gnd.n7131 gnd.n7130 19.3944
R7707 gnd.n7130 gnd.n7129 19.3944
R7708 gnd.n7129 gnd.n106 19.3944
R7709 gnd.n7124 gnd.n106 19.3944
R7710 gnd.n7124 gnd.n7123 19.3944
R7711 gnd.n7123 gnd.n7122 19.3944
R7712 gnd.n7122 gnd.n113 19.3944
R7713 gnd.n7117 gnd.n113 19.3944
R7714 gnd.n7117 gnd.n7116 19.3944
R7715 gnd.n5849 gnd.n5848 19.3944
R7716 gnd.n5848 gnd.n5847 19.3944
R7717 gnd.n5847 gnd.n1136 19.3944
R7718 gnd.n5690 gnd.n1136 19.3944
R7719 gnd.n5690 gnd.n1254 19.3944
R7720 gnd.n5696 gnd.n1254 19.3944
R7721 gnd.n5696 gnd.n5695 19.3944
R7722 gnd.n5695 gnd.n1228 19.3944
R7723 gnd.n5721 gnd.n1228 19.3944
R7724 gnd.n5721 gnd.n1226 19.3944
R7725 gnd.n5728 gnd.n1226 19.3944
R7726 gnd.n5728 gnd.n5727 19.3944
R7727 gnd.n5727 gnd.n1198 19.3944
R7728 gnd.n5759 gnd.n1198 19.3944
R7729 gnd.n5760 gnd.n5759 19.3944
R7730 gnd.n5761 gnd.n5760 19.3944
R7731 gnd.n1183 gnd.n1182 19.3944
R7732 gnd.n5780 gnd.n5779 19.3944
R7733 gnd.n5777 gnd.n5776 19.3944
R7734 gnd.n6930 gnd.n6929 19.3944
R7735 gnd.n6942 gnd.n221 19.3944
R7736 gnd.n6942 gnd.n213 19.3944
R7737 gnd.n6946 gnd.n213 19.3944
R7738 gnd.n6946 gnd.n200 19.3944
R7739 gnd.n6958 gnd.n200 19.3944
R7740 gnd.n6958 gnd.n198 19.3944
R7741 gnd.n6962 gnd.n198 19.3944
R7742 gnd.n6962 gnd.n184 19.3944
R7743 gnd.n6974 gnd.n184 19.3944
R7744 gnd.n6974 gnd.n182 19.3944
R7745 gnd.n6978 gnd.n182 19.3944
R7746 gnd.n6978 gnd.n166 19.3944
R7747 gnd.n7064 gnd.n166 19.3944
R7748 gnd.n7064 gnd.n164 19.3944
R7749 gnd.n7068 gnd.n164 19.3944
R7750 gnd.n7068 gnd.n87 19.3944
R7751 gnd.n7148 gnd.n87 19.3944
R7752 gnd.n3908 gnd.n3907 19.3944
R7753 gnd.n3911 gnd.n3908 19.3944
R7754 gnd.n3911 gnd.n3904 19.3944
R7755 gnd.n3915 gnd.n3904 19.3944
R7756 gnd.n3915 gnd.n2128 19.3944
R7757 gnd.n3919 gnd.n2128 19.3944
R7758 gnd.n3919 gnd.n2126 19.3944
R7759 gnd.n3926 gnd.n2126 19.3944
R7760 gnd.n3926 gnd.n3925 19.3944
R7761 gnd.n3925 gnd.n3924 19.3944
R7762 gnd.n3953 gnd.n3952 19.3944
R7763 gnd.n3963 gnd.n3962 19.3944
R7764 gnd.n3960 gnd.n3957 19.3944
R7765 gnd.n3955 gnd.n2069 19.3944
R7766 gnd.n4017 gnd.n4016 19.3944
R7767 gnd.n4022 gnd.n4017 19.3944
R7768 gnd.n4022 gnd.n4021 19.3944
R7769 gnd.n4021 gnd.n2042 19.3944
R7770 gnd.n4081 gnd.n2042 19.3944
R7771 gnd.n4081 gnd.n2040 19.3944
R7772 gnd.n4085 gnd.n2040 19.3944
R7773 gnd.n4085 gnd.n2038 19.3944
R7774 gnd.n4089 gnd.n2038 19.3944
R7775 gnd.n4089 gnd.n2036 19.3944
R7776 gnd.n4093 gnd.n2036 19.3944
R7777 gnd.n4093 gnd.n2034 19.3944
R7778 gnd.n4097 gnd.n2034 19.3944
R7779 gnd.n4097 gnd.n2032 19.3944
R7780 gnd.n4101 gnd.n2032 19.3944
R7781 gnd.n4101 gnd.n2030 19.3944
R7782 gnd.n4105 gnd.n2030 19.3944
R7783 gnd.n4105 gnd.n2028 19.3944
R7784 gnd.n4109 gnd.n2028 19.3944
R7785 gnd.n4109 gnd.n2024 19.3944
R7786 gnd.n4247 gnd.n2024 19.3944
R7787 gnd.n4247 gnd.n2022 19.3944
R7788 gnd.n4251 gnd.n2022 19.3944
R7789 gnd.n4251 gnd.n1771 19.3944
R7790 gnd.n4416 gnd.n1771 19.3944
R7791 gnd.n4416 gnd.n1769 19.3944
R7792 gnd.n4420 gnd.n1769 19.3944
R7793 gnd.n4420 gnd.n1756 19.3944
R7794 gnd.n4461 gnd.n1756 19.3944
R7795 gnd.n4461 gnd.n1754 19.3944
R7796 gnd.n4467 gnd.n1754 19.3944
R7797 gnd.n4467 gnd.n4466 19.3944
R7798 gnd.n4466 gnd.n1728 19.3944
R7799 gnd.n4512 gnd.n1728 19.3944
R7800 gnd.n4512 gnd.n1726 19.3944
R7801 gnd.n4516 gnd.n1726 19.3944
R7802 gnd.n4516 gnd.n1708 19.3944
R7803 gnd.n4549 gnd.n1708 19.3944
R7804 gnd.n4549 gnd.n1706 19.3944
R7805 gnd.n4553 gnd.n1706 19.3944
R7806 gnd.n4553 gnd.n1682 19.3944
R7807 gnd.n4590 gnd.n1682 19.3944
R7808 gnd.n4590 gnd.n1680 19.3944
R7809 gnd.n4594 gnd.n1680 19.3944
R7810 gnd.n4594 gnd.n1666 19.3944
R7811 gnd.n4635 gnd.n1666 19.3944
R7812 gnd.n4635 gnd.n1664 19.3944
R7813 gnd.n4641 gnd.n1664 19.3944
R7814 gnd.n4641 gnd.n4640 19.3944
R7815 gnd.n4640 gnd.n1638 19.3944
R7816 gnd.n4707 gnd.n1638 19.3944
R7817 gnd.n4707 gnd.n1636 19.3944
R7818 gnd.n4711 gnd.n1636 19.3944
R7819 gnd.n4711 gnd.n1617 19.3944
R7820 gnd.n4734 gnd.n1617 19.3944
R7821 gnd.n4734 gnd.n1615 19.3944
R7822 gnd.n4738 gnd.n1615 19.3944
R7823 gnd.n4738 gnd.n1596 19.3944
R7824 gnd.n4767 gnd.n1596 19.3944
R7825 gnd.n4767 gnd.n1594 19.3944
R7826 gnd.n4771 gnd.n1594 19.3944
R7827 gnd.n4771 gnd.n1579 19.3944
R7828 gnd.n4812 gnd.n1579 19.3944
R7829 gnd.n4812 gnd.n1577 19.3944
R7830 gnd.n4818 gnd.n1577 19.3944
R7831 gnd.n4818 gnd.n4817 19.3944
R7832 gnd.n4817 gnd.n1550 19.3944
R7833 gnd.n4860 gnd.n1550 19.3944
R7834 gnd.n4860 gnd.n1548 19.3944
R7835 gnd.n4864 gnd.n1548 19.3944
R7836 gnd.n4864 gnd.n1530 19.3944
R7837 gnd.n4888 gnd.n1530 19.3944
R7838 gnd.n4888 gnd.n1528 19.3944
R7839 gnd.n4900 gnd.n1528 19.3944
R7840 gnd.n4900 gnd.n4899 19.3944
R7841 gnd.n4899 gnd.n4898 19.3944
R7842 gnd.n4898 gnd.n1498 19.3944
R7843 gnd.n4963 gnd.n1498 19.3944
R7844 gnd.n4963 gnd.n1496 19.3944
R7845 gnd.n4969 gnd.n1496 19.3944
R7846 gnd.n4969 gnd.n4968 19.3944
R7847 gnd.n4968 gnd.n1470 19.3944
R7848 gnd.n5014 gnd.n1470 19.3944
R7849 gnd.n5014 gnd.n1468 19.3944
R7850 gnd.n5020 gnd.n1468 19.3944
R7851 gnd.n5020 gnd.n5019 19.3944
R7852 gnd.n5019 gnd.n1452 19.3944
R7853 gnd.n5041 gnd.n1452 19.3944
R7854 gnd.n5041 gnd.n1450 19.3944
R7855 gnd.n5045 gnd.n1450 19.3944
R7856 gnd.n5045 gnd.n1395 19.3944
R7857 gnd.n5084 gnd.n1395 19.3944
R7858 gnd.n5084 gnd.n1393 19.3944
R7859 gnd.n5088 gnd.n1393 19.3944
R7860 gnd.n5088 gnd.n1374 19.3944
R7861 gnd.n5113 gnd.n1374 19.3944
R7862 gnd.n5113 gnd.n1372 19.3944
R7863 gnd.n5120 gnd.n1372 19.3944
R7864 gnd.n5120 gnd.n5119 19.3944
R7865 gnd.n5119 gnd.n1343 19.3944
R7866 gnd.n5333 gnd.n1343 19.3944
R7867 gnd.n5333 gnd.n5332 19.3944
R7868 gnd.n5332 gnd.n5331 19.3944
R7869 gnd.n5331 gnd.n1349 19.3944
R7870 gnd.n1349 gnd.n1111 19.3944
R7871 gnd.n5864 gnd.n1111 19.3944
R7872 gnd.n5864 gnd.n5863 19.3944
R7873 gnd.n5863 gnd.n5862 19.3944
R7874 gnd.n5862 gnd.n1115 19.3944
R7875 gnd.n5856 gnd.n1115 19.3944
R7876 gnd.n5856 gnd.n5855 19.3944
R7877 gnd.n5855 gnd.n5854 19.3944
R7878 gnd.n5854 gnd.n1124 19.3944
R7879 gnd.n5676 gnd.n1124 19.3944
R7880 gnd.n5679 gnd.n5676 19.3944
R7881 gnd.n5679 gnd.n5673 19.3944
R7882 gnd.n5685 gnd.n5673 19.3944
R7883 gnd.n5685 gnd.n5684 19.3944
R7884 gnd.n5684 gnd.n1238 19.3944
R7885 gnd.n5710 gnd.n1238 19.3944
R7886 gnd.n5710 gnd.n1236 19.3944
R7887 gnd.n5716 gnd.n1236 19.3944
R7888 gnd.n5716 gnd.n5715 19.3944
R7889 gnd.n5715 gnd.n1210 19.3944
R7890 gnd.n5742 gnd.n1210 19.3944
R7891 gnd.n5742 gnd.n1208 19.3944
R7892 gnd.n5754 gnd.n1208 19.3944
R7893 gnd.n5754 gnd.n5753 19.3944
R7894 gnd.n5753 gnd.n5752 19.3944
R7895 gnd.n5749 gnd.n5748 19.3944
R7896 gnd.n5786 gnd.n5785 19.3944
R7897 gnd.n5807 gnd.n5806 19.3944
R7898 gnd.n5804 gnd.n5788 19.3944
R7899 gnd.n5800 gnd.n5799 19.3944
R7900 gnd.n5799 gnd.n5798 19.3944
R7901 gnd.n5798 gnd.n5795 19.3944
R7902 gnd.n5795 gnd.n272 19.3944
R7903 gnd.n6904 gnd.n272 19.3944
R7904 gnd.n6904 gnd.n6903 19.3944
R7905 gnd.n6903 gnd.n6902 19.3944
R7906 gnd.n6902 gnd.n276 19.3944
R7907 gnd.n6898 gnd.n276 19.3944
R7908 gnd.n6898 gnd.n6897 19.3944
R7909 gnd.n3838 gnd.n3837 19.3944
R7910 gnd.n3837 gnd.n3836 19.3944
R7911 gnd.n3836 gnd.n3835 19.3944
R7912 gnd.n3835 gnd.n3833 19.3944
R7913 gnd.n3833 gnd.n3830 19.3944
R7914 gnd.n3830 gnd.n3829 19.3944
R7915 gnd.n3829 gnd.n3826 19.3944
R7916 gnd.n3826 gnd.n3825 19.3944
R7917 gnd.n3825 gnd.n3822 19.3944
R7918 gnd.n3822 gnd.n3821 19.3944
R7919 gnd.n3821 gnd.n3818 19.3944
R7920 gnd.n3818 gnd.n3817 19.3944
R7921 gnd.n3817 gnd.n3814 19.3944
R7922 gnd.n3814 gnd.n3813 19.3944
R7923 gnd.n3813 gnd.n3810 19.3944
R7924 gnd.n3810 gnd.n3809 19.3944
R7925 gnd.n3809 gnd.n3806 19.3944
R7926 gnd.n3804 gnd.n3801 19.3944
R7927 gnd.n3801 gnd.n3800 19.3944
R7928 gnd.n3800 gnd.n3797 19.3944
R7929 gnd.n3797 gnd.n3796 19.3944
R7930 gnd.n3796 gnd.n3793 19.3944
R7931 gnd.n3793 gnd.n3792 19.3944
R7932 gnd.n3792 gnd.n3789 19.3944
R7933 gnd.n3789 gnd.n3788 19.3944
R7934 gnd.n3788 gnd.n3785 19.3944
R7935 gnd.n3785 gnd.n3784 19.3944
R7936 gnd.n3784 gnd.n3781 19.3944
R7937 gnd.n3781 gnd.n3780 19.3944
R7938 gnd.n3780 gnd.n3777 19.3944
R7939 gnd.n3777 gnd.n3776 19.3944
R7940 gnd.n3776 gnd.n3773 19.3944
R7941 gnd.n3773 gnd.n3772 19.3944
R7942 gnd.n3772 gnd.n3769 19.3944
R7943 gnd.n3769 gnd.n3768 19.3944
R7944 gnd.n3857 gnd.n2156 19.3944
R7945 gnd.n3857 gnd.n2157 19.3944
R7946 gnd.n3853 gnd.n2157 19.3944
R7947 gnd.n3853 gnd.n3852 19.3944
R7948 gnd.n3852 gnd.n3850 19.3944
R7949 gnd.n3850 gnd.n846 19.3944
R7950 gnd.n6082 gnd.n846 19.3944
R7951 gnd.n6082 gnd.n6081 19.3944
R7952 gnd.n6081 gnd.n6080 19.3944
R7953 gnd.n6080 gnd.n850 19.3944
R7954 gnd.n6070 gnd.n850 19.3944
R7955 gnd.n6070 gnd.n6069 19.3944
R7956 gnd.n6069 gnd.n6068 19.3944
R7957 gnd.n6068 gnd.n871 19.3944
R7958 gnd.n6058 gnd.n871 19.3944
R7959 gnd.n6058 gnd.n6057 19.3944
R7960 gnd.n6057 gnd.n6056 19.3944
R7961 gnd.n6056 gnd.n892 19.3944
R7962 gnd.n3970 gnd.n892 19.3944
R7963 gnd.n3971 gnd.n3970 19.3944
R7964 gnd.n3971 gnd.n2087 19.3944
R7965 gnd.n3996 gnd.n2087 19.3944
R7966 gnd.n3996 gnd.n3995 19.3944
R7967 gnd.n3995 gnd.n3994 19.3944
R7968 gnd.n3994 gnd.n915 19.3944
R7969 gnd.n6044 gnd.n915 19.3944
R7970 gnd.n6044 gnd.n6043 19.3944
R7971 gnd.n6043 gnd.n6042 19.3944
R7972 gnd.n6042 gnd.n919 19.3944
R7973 gnd.n6032 gnd.n919 19.3944
R7974 gnd.n6032 gnd.n6031 19.3944
R7975 gnd.n6031 gnd.n6030 19.3944
R7976 gnd.n6030 gnd.n938 19.3944
R7977 gnd.n6020 gnd.n938 19.3944
R7978 gnd.n6020 gnd.n6019 19.3944
R7979 gnd.n6019 gnd.n6018 19.3944
R7980 gnd.n6018 gnd.n960 19.3944
R7981 gnd.n6008 gnd.n960 19.3944
R7982 gnd.n6008 gnd.n6007 19.3944
R7983 gnd.n6007 gnd.n6006 19.3944
R7984 gnd.n6006 gnd.n981 19.3944
R7985 gnd.n5996 gnd.n981 19.3944
R7986 gnd.n3844 gnd.n2159 19.3944
R7987 gnd.n3652 gnd.n2159 19.3944
R7988 gnd.n3653 gnd.n3652 19.3944
R7989 gnd.n3656 gnd.n3653 19.3944
R7990 gnd.n3656 gnd.n3648 19.3944
R7991 gnd.n3662 gnd.n3648 19.3944
R7992 gnd.n3663 gnd.n3662 19.3944
R7993 gnd.n3666 gnd.n3663 19.3944
R7994 gnd.n3666 gnd.n3646 19.3944
R7995 gnd.n3672 gnd.n3646 19.3944
R7996 gnd.n3673 gnd.n3672 19.3944
R7997 gnd.n3676 gnd.n3673 19.3944
R7998 gnd.n3676 gnd.n3644 19.3944
R7999 gnd.n3682 gnd.n3644 19.3944
R8000 gnd.n3683 gnd.n3682 19.3944
R8001 gnd.n3686 gnd.n3683 19.3944
R8002 gnd.n3694 gnd.n3693 19.3944
R8003 gnd.n3693 gnd.n3692 19.3944
R8004 gnd.n3692 gnd.n2140 19.3944
R8005 gnd.n3871 gnd.n2140 19.3944
R8006 gnd.n3872 gnd.n3871 19.3944
R8007 gnd.n3874 gnd.n3872 19.3944
R8008 gnd.n3874 gnd.n2138 19.3944
R8009 gnd.n3879 gnd.n2138 19.3944
R8010 gnd.n3879 gnd.n2130 19.3944
R8011 gnd.n3899 gnd.n2130 19.3944
R8012 gnd.n3899 gnd.n3898 19.3944
R8013 gnd.n3898 gnd.n3897 19.3944
R8014 gnd.n3897 gnd.n2122 19.3944
R8015 gnd.n3931 gnd.n2122 19.3944
R8016 gnd.n3931 gnd.n2120 19.3944
R8017 gnd.n3937 gnd.n2120 19.3944
R8018 gnd.n3937 gnd.n3936 19.3944
R8019 gnd.n3936 gnd.n2109 19.3944
R8020 gnd.n3978 gnd.n2109 19.3944
R8021 gnd.n3978 gnd.n2107 19.3944
R8022 gnd.n3982 gnd.n2107 19.3944
R8023 gnd.n3982 gnd.n2075 19.3944
R8024 gnd.n4006 gnd.n2075 19.3944
R8025 gnd.n4006 gnd.n2073 19.3944
R8026 gnd.n4010 gnd.n2073 19.3944
R8027 gnd.n4010 gnd.n2063 19.3944
R8028 gnd.n4027 gnd.n2063 19.3944
R8029 gnd.n4027 gnd.n2061 19.3944
R8030 gnd.n4031 gnd.n2061 19.3944
R8031 gnd.n4031 gnd.n2045 19.3944
R8032 gnd.n4076 gnd.n2045 19.3944
R8033 gnd.n4076 gnd.n2046 19.3944
R8034 gnd.n4072 gnd.n2046 19.3944
R8035 gnd.n4072 gnd.n4071 19.3944
R8036 gnd.n4071 gnd.n4070 19.3944
R8037 gnd.n4070 gnd.n2051 19.3944
R8038 gnd.n4066 gnd.n2051 19.3944
R8039 gnd.n4066 gnd.n4065 19.3944
R8040 gnd.n4065 gnd.n4064 19.3944
R8041 gnd.n4064 gnd.n1996 19.3944
R8042 gnd.n4297 gnd.n1996 19.3944
R8043 gnd.n4297 gnd.n1997 19.3944
R8044 gnd.n3761 gnd.n3760 19.3944
R8045 gnd.n3760 gnd.n3746 19.3944
R8046 gnd.n3756 gnd.n3746 19.3944
R8047 gnd.n3756 gnd.n3755 19.3944
R8048 gnd.n3755 gnd.n3753 19.3944
R8049 gnd.n3753 gnd.n3752 19.3944
R8050 gnd.n3752 gnd.n2136 19.3944
R8051 gnd.n3883 gnd.n2136 19.3944
R8052 gnd.n3884 gnd.n3883 19.3944
R8053 gnd.n3885 gnd.n3884 19.3944
R8054 gnd.n3885 gnd.n2134 19.3944
R8055 gnd.n3893 gnd.n2134 19.3944
R8056 gnd.n3893 gnd.n3892 19.3944
R8057 gnd.n3892 gnd.n3891 19.3944
R8058 gnd.n3891 gnd.n2119 19.3944
R8059 gnd.n3941 gnd.n2119 19.3944
R8060 gnd.n3941 gnd.n2117 19.3944
R8061 gnd.n3947 gnd.n2117 19.3944
R8062 gnd.n3947 gnd.n3946 19.3944
R8063 gnd.n3946 gnd.n2091 19.3944
R8064 gnd.n3986 gnd.n2091 19.3944
R8065 gnd.n3986 gnd.n2103 19.3944
R8066 gnd.n2103 gnd.n2102 19.3944
R8067 gnd.n2102 gnd.n2101 19.3944
R8068 gnd.n2101 gnd.n2099 19.3944
R8069 gnd.n2099 gnd.n2098 19.3944
R8070 gnd.n2098 gnd.n2097 19.3944
R8071 gnd.n2097 gnd.n2060 19.3944
R8072 gnd.n4035 gnd.n2060 19.3944
R8073 gnd.n4035 gnd.n2058 19.3944
R8074 gnd.n4039 gnd.n2058 19.3944
R8075 gnd.n4040 gnd.n4039 19.3944
R8076 gnd.n4043 gnd.n4040 19.3944
R8077 gnd.n4043 gnd.n2056 19.3944
R8078 gnd.n4050 gnd.n2056 19.3944
R8079 gnd.n4051 gnd.n4050 19.3944
R8080 gnd.n4054 gnd.n4051 19.3944
R8081 gnd.n4054 gnd.n2054 19.3944
R8082 gnd.n4059 gnd.n2054 19.3944
R8083 gnd.n4059 gnd.n1995 19.3944
R8084 gnd.n4301 gnd.n1995 19.3944
R8085 gnd.n4302 gnd.n4301 19.3944
R8086 gnd.n4340 gnd.n1898 19.3944
R8087 gnd.n4340 gnd.n1905 19.3944
R8088 gnd.n1962 gnd.n1905 19.3944
R8089 gnd.n4333 gnd.n1962 19.3944
R8090 gnd.n4333 gnd.n4332 19.3944
R8091 gnd.n4332 gnd.n4331 19.3944
R8092 gnd.n4331 gnd.n1968 19.3944
R8093 gnd.n4326 gnd.n1968 19.3944
R8094 gnd.n4326 gnd.n4325 19.3944
R8095 gnd.n4325 gnd.n4324 19.3944
R8096 gnd.n4324 gnd.n1975 19.3944
R8097 gnd.n4319 gnd.n1975 19.3944
R8098 gnd.n4319 gnd.n4318 19.3944
R8099 gnd.n4318 gnd.n4317 19.3944
R8100 gnd.n4317 gnd.n1982 19.3944
R8101 gnd.n4312 gnd.n1982 19.3944
R8102 gnd.n4312 gnd.n4311 19.3944
R8103 gnd.n4311 gnd.n4310 19.3944
R8104 gnd.n1918 gnd.n1917 19.3944
R8105 gnd.n1958 gnd.n1917 19.3944
R8106 gnd.n1958 gnd.n1957 19.3944
R8107 gnd.n1957 gnd.n1956 19.3944
R8108 gnd.n1956 gnd.n1953 19.3944
R8109 gnd.n1953 gnd.n1952 19.3944
R8110 gnd.n1952 gnd.n1949 19.3944
R8111 gnd.n1949 gnd.n1948 19.3944
R8112 gnd.n1948 gnd.n1945 19.3944
R8113 gnd.n1945 gnd.n1944 19.3944
R8114 gnd.n1944 gnd.n1941 19.3944
R8115 gnd.n1941 gnd.n1940 19.3944
R8116 gnd.n1940 gnd.n1937 19.3944
R8117 gnd.n1937 gnd.n1936 19.3944
R8118 gnd.n1936 gnd.n1899 19.3944
R8119 gnd.n3861 gnd.n2149 19.3944
R8120 gnd.n3861 gnd.n2147 19.3944
R8121 gnd.n3866 gnd.n2147 19.3944
R8122 gnd.n3866 gnd.n834 19.3944
R8123 gnd.n6088 gnd.n834 19.3944
R8124 gnd.n6088 gnd.n6087 19.3944
R8125 gnd.n6087 gnd.n6086 19.3944
R8126 gnd.n6086 gnd.n838 19.3944
R8127 gnd.n6076 gnd.n838 19.3944
R8128 gnd.n6076 gnd.n6075 19.3944
R8129 gnd.n6075 gnd.n6074 19.3944
R8130 gnd.n6074 gnd.n860 19.3944
R8131 gnd.n6064 gnd.n860 19.3944
R8132 gnd.n6064 gnd.n6063 19.3944
R8133 gnd.n6063 gnd.n6062 19.3944
R8134 gnd.n6062 gnd.n882 19.3944
R8135 gnd.n6052 gnd.n6051 19.3944
R8136 gnd.n3967 gnd.n899 19.3944
R8137 gnd.n2083 gnd.n2082 19.3944
R8138 gnd.n4002 gnd.n4001 19.3944
R8139 gnd.n6048 gnd.n905 19.3944
R8140 gnd.n6048 gnd.n906 19.3944
R8141 gnd.n6038 gnd.n906 19.3944
R8142 gnd.n6038 gnd.n6037 19.3944
R8143 gnd.n6037 gnd.n6036 19.3944
R8144 gnd.n6036 gnd.n928 19.3944
R8145 gnd.n6026 gnd.n928 19.3944
R8146 gnd.n6026 gnd.n6025 19.3944
R8147 gnd.n6025 gnd.n6024 19.3944
R8148 gnd.n6024 gnd.n949 19.3944
R8149 gnd.n6014 gnd.n949 19.3944
R8150 gnd.n6014 gnd.n6013 19.3944
R8151 gnd.n6013 gnd.n6012 19.3944
R8152 gnd.n6012 gnd.n970 19.3944
R8153 gnd.n6002 gnd.n970 19.3944
R8154 gnd.n6002 gnd.n6001 19.3944
R8155 gnd.n6001 gnd.n6000 19.3944
R8156 gnd.n6261 gnd.n659 19.3944
R8157 gnd.n6255 gnd.n659 19.3944
R8158 gnd.n6255 gnd.n6254 19.3944
R8159 gnd.n6254 gnd.n6253 19.3944
R8160 gnd.n6253 gnd.n666 19.3944
R8161 gnd.n6247 gnd.n666 19.3944
R8162 gnd.n6247 gnd.n6246 19.3944
R8163 gnd.n6246 gnd.n6245 19.3944
R8164 gnd.n6245 gnd.n674 19.3944
R8165 gnd.n6239 gnd.n674 19.3944
R8166 gnd.n6239 gnd.n6238 19.3944
R8167 gnd.n6238 gnd.n6237 19.3944
R8168 gnd.n6237 gnd.n682 19.3944
R8169 gnd.n6231 gnd.n682 19.3944
R8170 gnd.n6231 gnd.n6230 19.3944
R8171 gnd.n6230 gnd.n6229 19.3944
R8172 gnd.n6229 gnd.n690 19.3944
R8173 gnd.n6223 gnd.n690 19.3944
R8174 gnd.n6223 gnd.n6222 19.3944
R8175 gnd.n6222 gnd.n6221 19.3944
R8176 gnd.n6221 gnd.n698 19.3944
R8177 gnd.n6215 gnd.n698 19.3944
R8178 gnd.n6215 gnd.n6214 19.3944
R8179 gnd.n6214 gnd.n6213 19.3944
R8180 gnd.n6213 gnd.n706 19.3944
R8181 gnd.n6207 gnd.n706 19.3944
R8182 gnd.n6207 gnd.n6206 19.3944
R8183 gnd.n6206 gnd.n6205 19.3944
R8184 gnd.n6205 gnd.n714 19.3944
R8185 gnd.n6199 gnd.n714 19.3944
R8186 gnd.n6199 gnd.n6198 19.3944
R8187 gnd.n6198 gnd.n6197 19.3944
R8188 gnd.n6197 gnd.n722 19.3944
R8189 gnd.n6191 gnd.n722 19.3944
R8190 gnd.n6191 gnd.n6190 19.3944
R8191 gnd.n6190 gnd.n6189 19.3944
R8192 gnd.n6189 gnd.n730 19.3944
R8193 gnd.n6183 gnd.n730 19.3944
R8194 gnd.n6183 gnd.n6182 19.3944
R8195 gnd.n6182 gnd.n6181 19.3944
R8196 gnd.n6181 gnd.n738 19.3944
R8197 gnd.n6175 gnd.n738 19.3944
R8198 gnd.n6175 gnd.n6174 19.3944
R8199 gnd.n6174 gnd.n6173 19.3944
R8200 gnd.n6173 gnd.n746 19.3944
R8201 gnd.n6167 gnd.n746 19.3944
R8202 gnd.n6167 gnd.n6166 19.3944
R8203 gnd.n6166 gnd.n6165 19.3944
R8204 gnd.n6165 gnd.n754 19.3944
R8205 gnd.n6159 gnd.n754 19.3944
R8206 gnd.n6159 gnd.n6158 19.3944
R8207 gnd.n6158 gnd.n6157 19.3944
R8208 gnd.n6157 gnd.n762 19.3944
R8209 gnd.n6151 gnd.n762 19.3944
R8210 gnd.n6151 gnd.n6150 19.3944
R8211 gnd.n6150 gnd.n6149 19.3944
R8212 gnd.n6149 gnd.n770 19.3944
R8213 gnd.n6143 gnd.n770 19.3944
R8214 gnd.n6143 gnd.n6142 19.3944
R8215 gnd.n6142 gnd.n6141 19.3944
R8216 gnd.n6141 gnd.n778 19.3944
R8217 gnd.n6135 gnd.n778 19.3944
R8218 gnd.n6135 gnd.n6134 19.3944
R8219 gnd.n6134 gnd.n6133 19.3944
R8220 gnd.n6133 gnd.n786 19.3944
R8221 gnd.n6127 gnd.n786 19.3944
R8222 gnd.n6127 gnd.n6126 19.3944
R8223 gnd.n6126 gnd.n6125 19.3944
R8224 gnd.n6125 gnd.n794 19.3944
R8225 gnd.n6119 gnd.n794 19.3944
R8226 gnd.n6119 gnd.n6118 19.3944
R8227 gnd.n6118 gnd.n6117 19.3944
R8228 gnd.n6117 gnd.n802 19.3944
R8229 gnd.n6111 gnd.n802 19.3944
R8230 gnd.n6111 gnd.n6110 19.3944
R8231 gnd.n6110 gnd.n6109 19.3944
R8232 gnd.n6109 gnd.n810 19.3944
R8233 gnd.n6103 gnd.n810 19.3944
R8234 gnd.n6103 gnd.n6102 19.3944
R8235 gnd.n6102 gnd.n6101 19.3944
R8236 gnd.n6101 gnd.n818 19.3944
R8237 gnd.n6095 gnd.n818 19.3944
R8238 gnd.n6095 gnd.n6094 19.3944
R8239 gnd.n6094 gnd.n6093 19.3944
R8240 gnd.n5991 gnd.n5990 19.3944
R8241 gnd.n5990 gnd.n5989 19.3944
R8242 gnd.n5989 gnd.n1005 19.3944
R8243 gnd.n5985 gnd.n1005 19.3944
R8244 gnd.n5985 gnd.n5984 19.3944
R8245 gnd.n5984 gnd.n5983 19.3944
R8246 gnd.n5983 gnd.n1010 19.3944
R8247 gnd.n5979 gnd.n1010 19.3944
R8248 gnd.n5979 gnd.n5978 19.3944
R8249 gnd.n5978 gnd.n5977 19.3944
R8250 gnd.n5977 gnd.n1015 19.3944
R8251 gnd.n5973 gnd.n1015 19.3944
R8252 gnd.n5973 gnd.n5972 19.3944
R8253 gnd.n5972 gnd.n5971 19.3944
R8254 gnd.n5971 gnd.n1020 19.3944
R8255 gnd.n5967 gnd.n1020 19.3944
R8256 gnd.n5967 gnd.n5966 19.3944
R8257 gnd.n5966 gnd.n5965 19.3944
R8258 gnd.n5965 gnd.n1025 19.3944
R8259 gnd.n5961 gnd.n1025 19.3944
R8260 gnd.n5961 gnd.n5960 19.3944
R8261 gnd.n5960 gnd.n5959 19.3944
R8262 gnd.n5959 gnd.n1030 19.3944
R8263 gnd.n5955 gnd.n1030 19.3944
R8264 gnd.n5955 gnd.n5954 19.3944
R8265 gnd.n5954 gnd.n5953 19.3944
R8266 gnd.n5953 gnd.n1035 19.3944
R8267 gnd.n5949 gnd.n1035 19.3944
R8268 gnd.n5949 gnd.n5948 19.3944
R8269 gnd.n5948 gnd.n5947 19.3944
R8270 gnd.n5947 gnd.n1040 19.3944
R8271 gnd.n5943 gnd.n1040 19.3944
R8272 gnd.n5943 gnd.n5942 19.3944
R8273 gnd.n5942 gnd.n5941 19.3944
R8274 gnd.n5941 gnd.n1045 19.3944
R8275 gnd.n5937 gnd.n1045 19.3944
R8276 gnd.n5937 gnd.n5936 19.3944
R8277 gnd.n5936 gnd.n5935 19.3944
R8278 gnd.n5935 gnd.n1050 19.3944
R8279 gnd.n5931 gnd.n1050 19.3944
R8280 gnd.n5931 gnd.n5930 19.3944
R8281 gnd.n5930 gnd.n5929 19.3944
R8282 gnd.n5929 gnd.n1055 19.3944
R8283 gnd.n5925 gnd.n1055 19.3944
R8284 gnd.n5925 gnd.n5924 19.3944
R8285 gnd.n5924 gnd.n5923 19.3944
R8286 gnd.n5923 gnd.n1060 19.3944
R8287 gnd.n5919 gnd.n1060 19.3944
R8288 gnd.n5919 gnd.n5918 19.3944
R8289 gnd.n5918 gnd.n5917 19.3944
R8290 gnd.n5917 gnd.n1065 19.3944
R8291 gnd.n5913 gnd.n1065 19.3944
R8292 gnd.n5913 gnd.n5912 19.3944
R8293 gnd.n5912 gnd.n5911 19.3944
R8294 gnd.n5911 gnd.n1070 19.3944
R8295 gnd.n5907 gnd.n1070 19.3944
R8296 gnd.n5907 gnd.n5906 19.3944
R8297 gnd.n5906 gnd.n5905 19.3944
R8298 gnd.n5905 gnd.n1075 19.3944
R8299 gnd.n5901 gnd.n1075 19.3944
R8300 gnd.n5901 gnd.n5900 19.3944
R8301 gnd.n5900 gnd.n5899 19.3944
R8302 gnd.n5899 gnd.n1080 19.3944
R8303 gnd.n5895 gnd.n1080 19.3944
R8304 gnd.n5895 gnd.n5894 19.3944
R8305 gnd.n5894 gnd.n5893 19.3944
R8306 gnd.n5893 gnd.n1085 19.3944
R8307 gnd.n5889 gnd.n1085 19.3944
R8308 gnd.n5889 gnd.n5888 19.3944
R8309 gnd.n5888 gnd.n5887 19.3944
R8310 gnd.n5887 gnd.n1090 19.3944
R8311 gnd.n5883 gnd.n1090 19.3944
R8312 gnd.n5883 gnd.n5882 19.3944
R8313 gnd.n5882 gnd.n5881 19.3944
R8314 gnd.n5881 gnd.n1095 19.3944
R8315 gnd.n5877 gnd.n1095 19.3944
R8316 gnd.n5877 gnd.n5876 19.3944
R8317 gnd.n5876 gnd.n5875 19.3944
R8318 gnd.n5875 gnd.n1100 19.3944
R8319 gnd.n5871 gnd.n1100 19.3944
R8320 gnd.n5871 gnd.n5870 19.3944
R8321 gnd.n5870 gnd.n5869 19.3944
R8322 gnd.n5316 gnd.n5151 19.3944
R8323 gnd.n5316 gnd.n5149 19.3944
R8324 gnd.n5321 gnd.n5149 19.3944
R8325 gnd.n5215 gnd.n5197 19.3944
R8326 gnd.n5215 gnd.n5195 19.3944
R8327 gnd.n5221 gnd.n5195 19.3944
R8328 gnd.n5221 gnd.n5188 19.3944
R8329 gnd.n5234 gnd.n5188 19.3944
R8330 gnd.n5234 gnd.n5186 19.3944
R8331 gnd.n5240 gnd.n5186 19.3944
R8332 gnd.n5240 gnd.n5179 19.3944
R8333 gnd.n5253 gnd.n5179 19.3944
R8334 gnd.n5253 gnd.n5177 19.3944
R8335 gnd.n5259 gnd.n5177 19.3944
R8336 gnd.n5259 gnd.n5170 19.3944
R8337 gnd.n5272 gnd.n5170 19.3944
R8338 gnd.n5272 gnd.n5168 19.3944
R8339 gnd.n5280 gnd.n5168 19.3944
R8340 gnd.n5280 gnd.n5279 19.3944
R8341 gnd.n5279 gnd.n5159 19.3944
R8342 gnd.n5293 gnd.n5159 19.3944
R8343 gnd.n5293 gnd.n5157 19.3944
R8344 gnd.n5299 gnd.n5157 19.3944
R8345 gnd.n5299 gnd.n5155 19.3944
R8346 gnd.n5303 gnd.n5155 19.3944
R8347 gnd.n5303 gnd.n5153 19.3944
R8348 gnd.n5312 gnd.n5153 19.3944
R8349 gnd.n2997 gnd.t127 18.8012
R8350 gnd.n2982 gnd.t144 18.8012
R8351 gnd.n2841 gnd.n2840 18.4825
R8352 gnd.n5554 gnd.n1291 18.4247
R8353 gnd.n4344 gnd.n1899 18.4247
R8354 gnd.n7027 gnd.n7026 18.2308
R8355 gnd.n5283 gnd.n5163 18.2308
R8356 gnd.n4204 gnd.n4188 18.2308
R8357 gnd.n3686 gnd.n3642 18.2308
R8358 gnd.t171 gnd.n2521 18.1639
R8359 gnd.n2549 gnd.t206 17.5266
R8360 gnd.n2948 gnd.t143 16.8893
R8361 gnd.n3859 gnd.t106 16.8893
R8362 gnd.n4299 gnd.t42 16.8893
R8363 gnd.n5612 gnd.t35 16.8893
R8364 gnd.t21 gnd.n81 16.8893
R8365 gnd.n2776 gnd.t122 16.2519
R8366 gnd.n2476 gnd.t190 16.2519
R8367 gnd.n4245 gnd.n4244 15.9333
R8368 gnd.n4244 gnd.n2020 15.9333
R8369 gnd.n4255 gnd.n4253 15.9333
R8370 gnd.n4255 gnd.n4254 15.9333
R8371 gnd.n4254 gnd.n1773 15.9333
R8372 gnd.n4414 gnd.n1773 15.9333
R8373 gnd.n4261 gnd.n1807 15.9333
R8374 gnd.n4459 gnd.n1758 15.9333
R8375 gnd.n4471 gnd.n4469 15.9333
R8376 gnd.n4435 gnd.n1747 15.9333
R8377 gnd.n4518 gnd.n1724 15.9333
R8378 gnd.n4547 gnd.n4546 15.9333
R8379 gnd.n4556 gnd.n4555 15.9333
R8380 gnd.n4588 gnd.n1684 15.9333
R8381 gnd.n4633 gnd.n1668 15.9333
R8382 gnd.n4644 gnd.n4643 15.9333
R8383 gnd.n4609 gnd.n1656 15.9333
R8384 gnd.n4705 gnd.n4704 15.9333
R8385 gnd.n4713 gnd.n1634 15.9333
R8386 gnd.n4732 gnd.n4731 15.9333
R8387 gnd.n4741 gnd.n4740 15.9333
R8388 gnd.n4765 gnd.n1599 15.9333
R8389 gnd.n4773 gnd.n1592 15.9333
R8390 gnd.n4810 gnd.n1582 15.9333
R8391 gnd.n4821 gnd.n1573 15.9333
R8392 gnd.n4821 gnd.n4820 15.9333
R8393 gnd.n4787 gnd.n1569 15.9333
R8394 gnd.n4858 gnd.n4857 15.9333
R8395 gnd.n4866 gnd.n1546 15.9333
R8396 gnd.n4886 gnd.n4885 15.9333
R8397 gnd.n4903 gnd.n4902 15.9333
R8398 gnd.n4896 gnd.n4895 15.9333
R8399 gnd.n4961 gnd.n1500 15.9333
R8400 gnd.n4972 gnd.n4971 15.9333
R8401 gnd.n4938 gnd.n1489 15.9333
R8402 gnd.n5012 gnd.n5011 15.9333
R8403 gnd.n5038 gnd.n5037 15.9333
R8404 gnd.n5065 gnd.n1412 15.9333
R8405 gnd.n5049 gnd.n1403 15.9333
R8406 gnd.n1441 gnd.n1399 15.9333
R8407 gnd.n5143 gnd.n1333 15.9333
R8408 gnd.n5143 gnd.n1296 15.9333
R8409 gnd.n5328 gnd.n5327 15.9333
R8410 gnd.n5327 gnd.n1106 15.9333
R8411 gnd.n5867 gnd.n1106 15.9333
R8412 gnd.n5867 gnd.n5866 15.9333
R8413 gnd.n1117 gnd.n1108 15.9333
R8414 gnd.n5860 gnd.n1117 15.9333
R8415 gnd.n3464 gnd.n3462 15.6674
R8416 gnd.n3432 gnd.n3430 15.6674
R8417 gnd.n3400 gnd.n3398 15.6674
R8418 gnd.n3369 gnd.n3367 15.6674
R8419 gnd.n3337 gnd.n3335 15.6674
R8420 gnd.n3305 gnd.n3303 15.6674
R8421 gnd.n3273 gnd.n3271 15.6674
R8422 gnd.n3242 gnd.n3240 15.6674
R8423 gnd.n2767 gnd.t122 15.6146
R8424 gnd.t56 gnd.n2242 15.6146
R8425 gnd.t60 gnd.n2243 15.6146
R8426 gnd.t93 gnd.n4413 15.6146
R8427 gnd.n1350 gnd.t77 15.6146
R8428 gnd.n1424 gnd.t46 15.296
R8429 gnd.n5344 gnd.n5343 15.0827
R8430 gnd.n1818 gnd.n1813 15.0481
R8431 gnd.n5354 gnd.n5353 15.0481
R8432 gnd.n3136 gnd.t205 14.9773
R8433 gnd.t106 gnd.n2143 14.9773
R8434 gnd.n4510 gnd.t281 14.9773
R8435 gnd.t2 gnd.n5099 14.9773
R8436 gnd.n7070 gnd.t21 14.9773
R8437 gnd.n4436 gnd.n1737 14.6587
R8438 gnd.n4564 gnd.t196 14.6587
R8439 gnd.n4625 gnd.n4624 14.6587
R8440 gnd.n5010 gnd.n1475 14.6587
R8441 gnd.n5057 gnd.t1 14.6587
R8442 gnd.n5111 gnd.n5110 14.6587
R8443 gnd.n5336 gnd.n5335 14.6587
R8444 gnd.t198 gnd.n2285 14.34
R8445 gnd.n3214 gnd.t170 14.34
R8446 gnd.n4519 gnd.n1721 14.0214
R8447 gnd.n4587 gnd.t174 14.0214
R8448 gnd.n4714 gnd.n1631 14.0214
R8449 gnd.n4764 gnd.n1601 14.0214
R8450 gnd.n4867 gnd.n1542 14.0214
R8451 gnd.n4926 gnd.n4925 14.0214
R8452 gnd.t178 gnd.n1454 14.0214
R8453 gnd.n1442 gnd.n1390 14.0214
R8454 gnd.t18 gnd.n1338 14.0214
R8455 gnd.n2923 gnd.t229 13.7027
R8456 gnd.n2633 gnd.n2632 13.5763
R8457 gnd.n3578 gnd.n2199 13.5763
R8458 gnd.n1271 gnd.n1270 13.5763
R8459 gnd.n7079 gnd.n7078 13.5763
R8460 gnd.n3768 gnd.n3743 13.5763
R8461 gnd.n4310 gnd.n1991 13.5763
R8462 gnd.n2841 gnd.n2579 13.384
R8463 gnd.n4451 gnd.t25 13.384
R8464 gnd.n4507 gnd.n1733 13.384
R8465 gnd.n4581 gnd.n1690 13.384
R8466 gnd.n4617 gnd.t231 13.384
R8467 gnd.n4703 gnd.n1643 13.384
R8468 gnd.n4758 gnd.n4757 13.384
R8469 gnd.n4856 gnd.n1555 13.384
R8470 gnd.n4953 gnd.n4952 13.384
R8471 gnd.t216 gnd.n1479 13.384
R8472 gnd.n4987 gnd.n1459 13.384
R8473 gnd.n5090 gnd.n1383 13.384
R8474 gnd.n1829 gnd.n1810 13.1884
R8475 gnd.n1824 gnd.n1823 13.1884
R8476 gnd.n1823 gnd.n1822 13.1884
R8477 gnd.n5347 gnd.n5342 13.1884
R8478 gnd.n5348 gnd.n5347 13.1884
R8479 gnd.n1825 gnd.n1812 13.146
R8480 gnd.n1821 gnd.n1812 13.146
R8481 gnd.n5346 gnd.n5345 13.146
R8482 gnd.n5346 gnd.n5341 13.146
R8483 gnd.n3465 gnd.n3461 12.8005
R8484 gnd.n3433 gnd.n3429 12.8005
R8485 gnd.n3401 gnd.n3397 12.8005
R8486 gnd.n3370 gnd.n3366 12.8005
R8487 gnd.n3338 gnd.n3334 12.8005
R8488 gnd.n3306 gnd.n3302 12.8005
R8489 gnd.n3274 gnd.n3270 12.8005
R8490 gnd.n3243 gnd.n3239 12.8005
R8491 gnd.n4423 gnd.n1764 12.7467
R8492 gnd.t53 gnd.t64 12.7467
R8493 gnd.n4500 gnd.n1730 12.7467
R8494 gnd.t132 gnd.n1710 12.7467
R8495 gnd.n4597 gnd.n1675 12.7467
R8496 gnd.n4696 gnd.n1640 12.7467
R8497 gnd.n4774 gnd.n1588 12.7467
R8498 gnd.n4849 gnd.n1552 12.7467
R8499 gnd.n4960 gnd.n1503 12.7467
R8500 gnd.n5023 gnd.n1465 12.7467
R8501 gnd.n5075 gnd.t240 12.7467
R8502 gnd.n5098 gnd.n1385 12.7467
R8503 gnd.n5122 gnd.t90 12.7467
R8504 gnd.n6091 gnd.n827 12.4281
R8505 gnd.n7062 gnd.n168 12.4281
R8506 gnd.n2632 gnd.n2627 12.4126
R8507 gnd.n3581 gnd.n3578 12.4126
R8508 gnd.n5606 gnd.n1270 12.4126
R8509 gnd.n7078 gnd.n155 12.4126
R8510 gnd.n3764 gnd.n3743 12.4126
R8511 gnd.n4305 gnd.n1991 12.4126
R8512 gnd.n4409 gnd.n1830 12.1761
R8513 gnd.n5423 gnd.n5422 12.1761
R8514 gnd.n1723 gnd.n1715 12.1094
R8515 gnd.n4534 gnd.n1699 12.1094
R8516 gnd.n1633 gnd.n1624 12.1094
R8517 gnd.n4750 gnd.n4749 12.1094
R8518 gnd.n1544 gnd.n1537 12.1094
R8519 gnd.n4894 gnd.n1518 12.1094
R8520 gnd.n5036 gnd.n1417 12.1094
R8521 gnd.n5082 gnd.n5081 12.1094
R8522 gnd.n3469 gnd.n3468 12.0247
R8523 gnd.n3437 gnd.n3436 12.0247
R8524 gnd.n3405 gnd.n3404 12.0247
R8525 gnd.n3374 gnd.n3373 12.0247
R8526 gnd.n3342 gnd.n3341 12.0247
R8527 gnd.n3310 gnd.n3309 12.0247
R8528 gnd.n3278 gnd.n3277 12.0247
R8529 gnd.n3247 gnd.n3246 12.0247
R8530 gnd.n6016 gnd.t249 11.7908
R8531 gnd.n5698 gnd.t11 11.7908
R8532 gnd.n4111 gnd.n1961 11.4721
R8533 gnd.n4458 gnd.n1760 11.4721
R8534 gnd.n4632 gnd.n1671 11.4721
R8535 gnd.n4651 gnd.n4650 11.4721
R8536 gnd.n4809 gnd.n1584 11.4721
R8537 gnd.n4828 gnd.n4827 11.4721
R8538 gnd.n4980 gnd.n1487 11.4721
R8539 gnd.n5003 gnd.n1472 11.4721
R8540 gnd.n5125 gnd.n5124 11.4721
R8541 gnd.n1427 gnd.n1426 11.4721
R8542 gnd.n5858 gnd.n1118 11.4721
R8543 gnd.n3472 gnd.n3459 11.249
R8544 gnd.n3440 gnd.n3427 11.249
R8545 gnd.n3408 gnd.n3395 11.249
R8546 gnd.n3377 gnd.n3364 11.249
R8547 gnd.n3345 gnd.n3332 11.249
R8548 gnd.n3313 gnd.n3300 11.249
R8549 gnd.n3281 gnd.n3268 11.249
R8550 gnd.n3250 gnd.n3237 11.249
R8551 gnd.n2911 gnd.t229 11.1535
R8552 gnd.t164 gnd.n865 11.1535
R8553 gnd.n6040 gnd.t256 11.1535
R8554 gnd.n5757 gnd.t241 11.1535
R8555 gnd.n6906 gnd.t13 11.1535
R8556 gnd.n840 gnd.n830 10.8348
R8557 gnd.n6084 gnd.n843 10.8348
R8558 gnd.n3881 gnd.n852 10.8348
R8559 gnd.n3901 gnd.n862 10.8348
R8560 gnd.n6072 gnd.n865 10.8348
R8561 gnd.n3895 gnd.n873 10.8348
R8562 gnd.n6066 gnd.n876 10.8348
R8563 gnd.n3929 gnd.n3928 10.8348
R8564 gnd.n6060 gnd.n886 10.8348
R8565 gnd.n3939 gnd.n894 10.8348
R8566 gnd.n3949 gnd.n2111 10.8348
R8567 gnd.n3976 gnd.n3965 10.8348
R8568 gnd.n3973 gnd.n2105 10.8348
R8569 gnd.n3984 gnd.n2084 10.8348
R8570 gnd.n4004 gnd.n2079 10.8348
R8571 gnd.n4013 gnd.n2070 10.8348
R8572 gnd.n4012 gnd.n909 10.8348
R8573 gnd.n6046 gnd.n912 10.8348
R8574 gnd.n4025 gnd.n4024 10.8348
R8575 gnd.n6040 gnd.n923 10.8348
R8576 gnd.n4033 gnd.n930 10.8348
R8577 gnd.n4078 gnd.n940 10.8348
R8578 gnd.n6028 gnd.n943 10.8348
R8579 gnd.n4041 gnd.n951 10.8348
R8580 gnd.n6022 gnd.n954 10.8348
R8581 gnd.n4048 gnd.n4047 10.8348
R8582 gnd.n6016 gnd.n964 10.8348
R8583 gnd.n4052 gnd.n972 10.8348
R8584 gnd.n6010 gnd.n975 10.8348
R8585 gnd.n4061 gnd.n983 10.8348
R8586 gnd.n6004 gnd.n986 10.8348
R8587 gnd.n4299 gnd.n993 10.8348
R8588 gnd.n5998 gnd.n996 10.8348
R8589 gnd.n4544 gnd.n4543 10.8348
R8590 gnd.n4610 gnd.t237 10.8348
R8591 gnd.n4730 gnd.n1610 10.8348
R8592 gnd.n4742 gnd.n1610 10.8348
R8593 gnd.n4884 gnd.n1523 10.8348
R8594 gnd.n4904 gnd.n1523 10.8348
R8595 gnd.n4973 gnd.t160 10.8348
R8596 gnd.n5050 gnd.n5047 10.8348
R8597 gnd.n5852 gnd.n5851 10.8348
R8598 gnd.n5612 gnd.n1129 10.8348
R8599 gnd.n5845 gnd.n1138 10.8348
R8600 gnd.n5621 gnd.n1141 10.8348
R8601 gnd.n5688 gnd.n1256 10.8348
R8602 gnd.n5687 gnd.n5670 10.8348
R8603 gnd.n5698 gnd.n1249 10.8348
R8604 gnd.n1251 gnd.n1241 10.8348
R8605 gnd.n5708 gnd.n5707 10.8348
R8606 gnd.n5719 gnd.n1230 10.8348
R8607 gnd.n5718 gnd.n1233 10.8348
R8608 gnd.n5730 gnd.n1220 10.8348
R8609 gnd.n5740 gnd.n5739 10.8348
R8610 gnd.n5757 gnd.n1201 10.8348
R8611 gnd.n5756 gnd.n1205 10.8348
R8612 gnd.n5763 gnd.n1194 10.8348
R8613 gnd.n5650 gnd.n1196 10.8348
R8614 gnd.n5773 gnd.n1184 10.8348
R8615 gnd.n5772 gnd.n1176 10.8348
R8616 gnd.n1180 gnd.n1170 10.8348
R8617 gnd.n5810 gnd.n5809 10.8348
R8618 gnd.n6927 gnd.n235 10.8348
R8619 gnd.n6932 gnd.n231 10.8348
R8620 gnd.n6940 gnd.n223 10.8348
R8621 gnd.n6916 gnd.n225 10.8348
R8622 gnd.n6948 gnd.n209 10.8348
R8623 gnd.n6912 gnd.n211 10.8348
R8624 gnd.n6956 gnd.n202 10.8348
R8625 gnd.n6907 gnd.n6906 10.8348
R8626 gnd.n6964 gnd.n194 10.8348
R8627 gnd.n6972 gnd.n186 10.8348
R8628 gnd.n261 gnd.n188 10.8348
R8629 gnd.n6980 gnd.n177 10.8348
R8630 gnd.n5488 gnd.n1292 10.6151
R8631 gnd.n5488 gnd.n5487 10.6151
R8632 gnd.n5485 gnd.n5482 10.6151
R8633 gnd.n5482 gnd.n5481 10.6151
R8634 gnd.n5481 gnd.n5478 10.6151
R8635 gnd.n5478 gnd.n5477 10.6151
R8636 gnd.n5477 gnd.n5474 10.6151
R8637 gnd.n5474 gnd.n5473 10.6151
R8638 gnd.n5473 gnd.n5470 10.6151
R8639 gnd.n5470 gnd.n5469 10.6151
R8640 gnd.n5469 gnd.n5466 10.6151
R8641 gnd.n5466 gnd.n5465 10.6151
R8642 gnd.n5465 gnd.n5462 10.6151
R8643 gnd.n5462 gnd.n5461 10.6151
R8644 gnd.n5461 gnd.n5458 10.6151
R8645 gnd.n5458 gnd.n5457 10.6151
R8646 gnd.n5457 gnd.n5454 10.6151
R8647 gnd.n5454 gnd.n5453 10.6151
R8648 gnd.n5453 gnd.n5450 10.6151
R8649 gnd.n5450 gnd.n5449 10.6151
R8650 gnd.n5449 gnd.n5446 10.6151
R8651 gnd.n5446 gnd.n5445 10.6151
R8652 gnd.n5445 gnd.n5442 10.6151
R8653 gnd.n5442 gnd.n5441 10.6151
R8654 gnd.n5441 gnd.n5438 10.6151
R8655 gnd.n5438 gnd.n5437 10.6151
R8656 gnd.n5437 gnd.n5434 10.6151
R8657 gnd.n5434 gnd.n5433 10.6151
R8658 gnd.n5433 gnd.n5430 10.6151
R8659 gnd.n5430 gnd.n5429 10.6151
R8660 gnd.n4426 gnd.n4425 10.6151
R8661 gnd.n4448 gnd.n4426 10.6151
R8662 gnd.n4448 gnd.n4447 10.6151
R8663 gnd.n4447 gnd.n4446 10.6151
R8664 gnd.n4446 gnd.n4442 10.6151
R8665 gnd.n4442 gnd.n4441 10.6151
R8666 gnd.n4441 gnd.n4439 10.6151
R8667 gnd.n4439 gnd.n4438 10.6151
R8668 gnd.n4438 gnd.n4434 10.6151
R8669 gnd.n4434 gnd.n4433 10.6151
R8670 gnd.n4433 gnd.n4431 10.6151
R8671 gnd.n4431 gnd.n4430 10.6151
R8672 gnd.n4430 gnd.n4427 10.6151
R8673 gnd.n4427 gnd.n1713 10.6151
R8674 gnd.n4528 gnd.n1713 10.6151
R8675 gnd.n4529 gnd.n4528 10.6151
R8676 gnd.n4541 gnd.n4529 10.6151
R8677 gnd.n4541 gnd.n4540 10.6151
R8678 gnd.n4540 gnd.n4539 10.6151
R8679 gnd.n4539 gnd.n4537 10.6151
R8680 gnd.n4537 gnd.n4536 10.6151
R8681 gnd.n4536 gnd.n4533 10.6151
R8682 gnd.n4533 gnd.n4532 10.6151
R8683 gnd.n4532 gnd.n1677 10.6151
R8684 gnd.n4599 gnd.n1677 10.6151
R8685 gnd.n4600 gnd.n4599 10.6151
R8686 gnd.n4622 gnd.n4600 10.6151
R8687 gnd.n4622 gnd.n4621 10.6151
R8688 gnd.n4621 gnd.n4620 10.6151
R8689 gnd.n4620 gnd.n4616 10.6151
R8690 gnd.n4616 gnd.n4615 10.6151
R8691 gnd.n4615 gnd.n4613 10.6151
R8692 gnd.n4613 gnd.n4612 10.6151
R8693 gnd.n4612 gnd.n4608 10.6151
R8694 gnd.n4608 gnd.n4607 10.6151
R8695 gnd.n4607 gnd.n4605 10.6151
R8696 gnd.n4605 gnd.n4604 10.6151
R8697 gnd.n4604 gnd.n4601 10.6151
R8698 gnd.n4601 gnd.n1622 10.6151
R8699 gnd.n4723 gnd.n1622 10.6151
R8700 gnd.n4724 gnd.n4723 10.6151
R8701 gnd.n4728 gnd.n4724 10.6151
R8702 gnd.n4728 gnd.n4727 10.6151
R8703 gnd.n4727 gnd.n4726 10.6151
R8704 gnd.n4726 gnd.n1605 10.6151
R8705 gnd.n4752 gnd.n1605 10.6151
R8706 gnd.n4753 gnd.n4752 10.6151
R8707 gnd.n4754 gnd.n4753 10.6151
R8708 gnd.n4754 gnd.n1590 10.6151
R8709 gnd.n4776 gnd.n1590 10.6151
R8710 gnd.n4777 gnd.n4776 10.6151
R8711 gnd.n4799 gnd.n4777 10.6151
R8712 gnd.n4799 gnd.n4798 10.6151
R8713 gnd.n4798 gnd.n4797 10.6151
R8714 gnd.n4797 gnd.n4794 10.6151
R8715 gnd.n4794 gnd.n4793 10.6151
R8716 gnd.n4793 gnd.n4791 10.6151
R8717 gnd.n4791 gnd.n4790 10.6151
R8718 gnd.n4790 gnd.n4785 10.6151
R8719 gnd.n4785 gnd.n4784 10.6151
R8720 gnd.n4784 gnd.n4782 10.6151
R8721 gnd.n4782 gnd.n4781 10.6151
R8722 gnd.n4781 gnd.n4778 10.6151
R8723 gnd.n4778 gnd.n1535 10.6151
R8724 gnd.n4876 gnd.n1535 10.6151
R8725 gnd.n4877 gnd.n4876 10.6151
R8726 gnd.n4882 gnd.n4877 10.6151
R8727 gnd.n4882 gnd.n4881 10.6151
R8728 gnd.n4881 gnd.n4880 10.6151
R8729 gnd.n4880 gnd.n4878 10.6151
R8730 gnd.n4878 gnd.n1508 10.6151
R8731 gnd.n4928 gnd.n1508 10.6151
R8732 gnd.n4929 gnd.n4928 10.6151
R8733 gnd.n4950 gnd.n4929 10.6151
R8734 gnd.n4950 gnd.n4949 10.6151
R8735 gnd.n4949 gnd.n4948 10.6151
R8736 gnd.n4948 gnd.n4944 10.6151
R8737 gnd.n4944 gnd.n4943 10.6151
R8738 gnd.n4943 gnd.n4941 10.6151
R8739 gnd.n4941 gnd.n4940 10.6151
R8740 gnd.n4940 gnd.n4937 10.6151
R8741 gnd.n4937 gnd.n4936 10.6151
R8742 gnd.n4936 gnd.n4934 10.6151
R8743 gnd.n4934 gnd.n4933 10.6151
R8744 gnd.n4933 gnd.n4930 10.6151
R8745 gnd.n4930 gnd.n1457 10.6151
R8746 gnd.n5032 gnd.n1457 10.6151
R8747 gnd.n5033 gnd.n5032 10.6151
R8748 gnd.n5034 gnd.n5033 10.6151
R8749 gnd.n5034 gnd.n1419 10.6151
R8750 gnd.n5054 gnd.n1419 10.6151
R8751 gnd.n5054 gnd.n5053 10.6151
R8752 gnd.n5053 gnd.n5052 10.6151
R8753 gnd.n5052 gnd.n1448 10.6151
R8754 gnd.n1448 gnd.n1447 10.6151
R8755 gnd.n1447 gnd.n1445 10.6151
R8756 gnd.n1445 gnd.n1444 10.6151
R8757 gnd.n1444 gnd.n1440 10.6151
R8758 gnd.n1440 gnd.n1439 10.6151
R8759 gnd.n1439 gnd.n1437 10.6151
R8760 gnd.n1437 gnd.n1436 10.6151
R8761 gnd.n1436 gnd.n1434 10.6151
R8762 gnd.n1434 gnd.n1433 10.6151
R8763 gnd.n1433 gnd.n1432 10.6151
R8764 gnd.n1432 gnd.n1431 10.6151
R8765 gnd.n1431 gnd.n1430 10.6151
R8766 gnd.n1430 gnd.n1422 10.6151
R8767 gnd.n1422 gnd.n1421 10.6151
R8768 gnd.n1421 gnd.n1420 10.6151
R8769 gnd.n1420 gnd.n1331 10.6151
R8770 gnd.n1897 gnd.n1896 10.6151
R8771 gnd.n1896 gnd.n1893 10.6151
R8772 gnd.n1891 gnd.n1888 10.6151
R8773 gnd.n1888 gnd.n1887 10.6151
R8774 gnd.n1887 gnd.n1884 10.6151
R8775 gnd.n1884 gnd.n1883 10.6151
R8776 gnd.n1883 gnd.n1880 10.6151
R8777 gnd.n1880 gnd.n1879 10.6151
R8778 gnd.n1879 gnd.n1876 10.6151
R8779 gnd.n1876 gnd.n1875 10.6151
R8780 gnd.n1875 gnd.n1872 10.6151
R8781 gnd.n1872 gnd.n1871 10.6151
R8782 gnd.n1871 gnd.n1868 10.6151
R8783 gnd.n1868 gnd.n1867 10.6151
R8784 gnd.n1867 gnd.n1864 10.6151
R8785 gnd.n1864 gnd.n1863 10.6151
R8786 gnd.n1863 gnd.n1860 10.6151
R8787 gnd.n1860 gnd.n1859 10.6151
R8788 gnd.n1859 gnd.n1856 10.6151
R8789 gnd.n1856 gnd.n1855 10.6151
R8790 gnd.n1855 gnd.n1852 10.6151
R8791 gnd.n1852 gnd.n1851 10.6151
R8792 gnd.n1851 gnd.n1848 10.6151
R8793 gnd.n1848 gnd.n1847 10.6151
R8794 gnd.n1847 gnd.n1844 10.6151
R8795 gnd.n1844 gnd.n1843 10.6151
R8796 gnd.n1843 gnd.n1840 10.6151
R8797 gnd.n1840 gnd.n1839 10.6151
R8798 gnd.n1839 gnd.n1836 10.6151
R8799 gnd.n1836 gnd.n1766 10.6151
R8800 gnd.n4409 gnd.n4408 10.6151
R8801 gnd.n4408 gnd.n4407 10.6151
R8802 gnd.n4407 gnd.n4406 10.6151
R8803 gnd.n4406 gnd.n4404 10.6151
R8804 gnd.n4404 gnd.n4401 10.6151
R8805 gnd.n4401 gnd.n4400 10.6151
R8806 gnd.n4400 gnd.n4397 10.6151
R8807 gnd.n4397 gnd.n4396 10.6151
R8808 gnd.n4396 gnd.n4393 10.6151
R8809 gnd.n4393 gnd.n4392 10.6151
R8810 gnd.n4392 gnd.n4389 10.6151
R8811 gnd.n4389 gnd.n4388 10.6151
R8812 gnd.n4388 gnd.n4385 10.6151
R8813 gnd.n4385 gnd.n4384 10.6151
R8814 gnd.n4384 gnd.n4381 10.6151
R8815 gnd.n4381 gnd.n4380 10.6151
R8816 gnd.n4380 gnd.n4377 10.6151
R8817 gnd.n4377 gnd.n4376 10.6151
R8818 gnd.n4376 gnd.n4373 10.6151
R8819 gnd.n4373 gnd.n4372 10.6151
R8820 gnd.n4372 gnd.n4369 10.6151
R8821 gnd.n4369 gnd.n4368 10.6151
R8822 gnd.n4368 gnd.n4365 10.6151
R8823 gnd.n4365 gnd.n4364 10.6151
R8824 gnd.n4364 gnd.n4361 10.6151
R8825 gnd.n4361 gnd.n4360 10.6151
R8826 gnd.n4360 gnd.n4357 10.6151
R8827 gnd.n4357 gnd.n4356 10.6151
R8828 gnd.n4353 gnd.n4352 10.6151
R8829 gnd.n4352 gnd.n4349 10.6151
R8830 gnd.n5422 gnd.n5421 10.6151
R8831 gnd.n5421 gnd.n5418 10.6151
R8832 gnd.n5418 gnd.n5417 10.6151
R8833 gnd.n5417 gnd.n5414 10.6151
R8834 gnd.n5414 gnd.n5413 10.6151
R8835 gnd.n5413 gnd.n5410 10.6151
R8836 gnd.n5410 gnd.n5409 10.6151
R8837 gnd.n5409 gnd.n5406 10.6151
R8838 gnd.n5406 gnd.n5405 10.6151
R8839 gnd.n5405 gnd.n5402 10.6151
R8840 gnd.n5402 gnd.n5401 10.6151
R8841 gnd.n5401 gnd.n5398 10.6151
R8842 gnd.n5398 gnd.n5397 10.6151
R8843 gnd.n5397 gnd.n5394 10.6151
R8844 gnd.n5394 gnd.n5393 10.6151
R8845 gnd.n5393 gnd.n5390 10.6151
R8846 gnd.n5390 gnd.n5389 10.6151
R8847 gnd.n5389 gnd.n5386 10.6151
R8848 gnd.n5386 gnd.n5385 10.6151
R8849 gnd.n5385 gnd.n5382 10.6151
R8850 gnd.n5382 gnd.n5381 10.6151
R8851 gnd.n5381 gnd.n5378 10.6151
R8852 gnd.n5378 gnd.n5377 10.6151
R8853 gnd.n5377 gnd.n5374 10.6151
R8854 gnd.n5374 gnd.n5373 10.6151
R8855 gnd.n5373 gnd.n5370 10.6151
R8856 gnd.n5370 gnd.n5369 10.6151
R8857 gnd.n5369 gnd.n5366 10.6151
R8858 gnd.n5364 gnd.n5361 10.6151
R8859 gnd.n5361 gnd.n1293 10.6151
R8860 gnd.n4454 gnd.n1762 10.6151
R8861 gnd.n4455 gnd.n4454 10.6151
R8862 gnd.n4456 gnd.n4455 10.6151
R8863 gnd.n4456 gnd.n1749 10.6151
R8864 gnd.n4473 gnd.n1749 10.6151
R8865 gnd.n4474 gnd.n4473 10.6151
R8866 gnd.n4475 gnd.n4474 10.6151
R8867 gnd.n4475 gnd.n1735 10.6151
R8868 gnd.n4503 gnd.n1735 10.6151
R8869 gnd.n4504 gnd.n4503 10.6151
R8870 gnd.n4505 gnd.n4504 10.6151
R8871 gnd.n4505 gnd.n1719 10.6151
R8872 gnd.n4521 gnd.n1719 10.6151
R8873 gnd.n4522 gnd.n4521 10.6151
R8874 gnd.n4524 gnd.n4522 10.6151
R8875 gnd.n4524 gnd.n4523 10.6151
R8876 gnd.n4523 gnd.n1701 10.6151
R8877 gnd.n4559 gnd.n1701 10.6151
R8878 gnd.n4560 gnd.n4559 10.6151
R8879 gnd.n4561 gnd.n4560 10.6151
R8880 gnd.n4561 gnd.n1689 10.6151
R8881 gnd.n4585 gnd.n1689 10.6151
R8882 gnd.n4585 gnd.n4584 10.6151
R8883 gnd.n4584 gnd.n4583 10.6151
R8884 gnd.n4583 gnd.n1673 10.6151
R8885 gnd.n4628 gnd.n1673 10.6151
R8886 gnd.n4629 gnd.n4628 10.6151
R8887 gnd.n4630 gnd.n4629 10.6151
R8888 gnd.n4630 gnd.n1658 10.6151
R8889 gnd.n4646 gnd.n1658 10.6151
R8890 gnd.n4647 gnd.n4646 10.6151
R8891 gnd.n4648 gnd.n4647 10.6151
R8892 gnd.n4648 gnd.n1645 10.6151
R8893 gnd.n4699 gnd.n1645 10.6151
R8894 gnd.n4700 gnd.n4699 10.6151
R8895 gnd.n4701 gnd.n4700 10.6151
R8896 gnd.n4701 gnd.n1629 10.6151
R8897 gnd.n4716 gnd.n1629 10.6151
R8898 gnd.n4717 gnd.n4716 10.6151
R8899 gnd.n4719 gnd.n4717 10.6151
R8900 gnd.n4719 gnd.n4718 10.6151
R8901 gnd.n4718 gnd.n1608 10.6151
R8902 gnd.n4744 gnd.n1608 10.6151
R8903 gnd.n4745 gnd.n4744 10.6151
R8904 gnd.n4746 gnd.n4745 10.6151
R8905 gnd.n4746 gnd.n1604 10.6151
R8906 gnd.n4762 gnd.n1604 10.6151
R8907 gnd.n4762 gnd.n4761 10.6151
R8908 gnd.n4761 gnd.n4760 10.6151
R8909 gnd.n4760 gnd.n1586 10.6151
R8910 gnd.n4805 gnd.n1586 10.6151
R8911 gnd.n4806 gnd.n4805 10.6151
R8912 gnd.n4807 gnd.n4806 10.6151
R8913 gnd.n4807 gnd.n1571 10.6151
R8914 gnd.n4823 gnd.n1571 10.6151
R8915 gnd.n4824 gnd.n4823 10.6151
R8916 gnd.n4825 gnd.n4824 10.6151
R8917 gnd.n4825 gnd.n1557 10.6151
R8918 gnd.n4852 gnd.n1557 10.6151
R8919 gnd.n4853 gnd.n4852 10.6151
R8920 gnd.n4854 gnd.n4853 10.6151
R8921 gnd.n4854 gnd.n1540 10.6151
R8922 gnd.n4869 gnd.n1540 10.6151
R8923 gnd.n4870 gnd.n4869 10.6151
R8924 gnd.n4872 gnd.n4870 10.6151
R8925 gnd.n4872 gnd.n4871 10.6151
R8926 gnd.n4871 gnd.n1521 10.6151
R8927 gnd.n4906 gnd.n1521 10.6151
R8928 gnd.n4907 gnd.n4906 10.6151
R8929 gnd.n4909 gnd.n4907 10.6151
R8930 gnd.n4909 gnd.n4908 10.6151
R8931 gnd.n4908 gnd.n1505 10.6151
R8932 gnd.n4956 gnd.n1505 10.6151
R8933 gnd.n4957 gnd.n4956 10.6151
R8934 gnd.n4958 gnd.n4957 10.6151
R8935 gnd.n4958 gnd.n1491 10.6151
R8936 gnd.n4975 gnd.n1491 10.6151
R8937 gnd.n4976 gnd.n4975 10.6151
R8938 gnd.n4977 gnd.n4976 10.6151
R8939 gnd.n4977 gnd.n1477 10.6151
R8940 gnd.n5006 gnd.n1477 10.6151
R8941 gnd.n5007 gnd.n5006 10.6151
R8942 gnd.n5008 gnd.n5007 10.6151
R8943 gnd.n5008 gnd.n1463 10.6151
R8944 gnd.n5025 gnd.n1463 10.6151
R8945 gnd.n5026 gnd.n5025 10.6151
R8946 gnd.n5028 gnd.n5026 10.6151
R8947 gnd.n5028 gnd.n5027 10.6151
R8948 gnd.n5027 gnd.n1415 10.6151
R8949 gnd.n5060 gnd.n1415 10.6151
R8950 gnd.n5061 gnd.n5060 10.6151
R8951 gnd.n5062 gnd.n5061 10.6151
R8952 gnd.n5062 gnd.n1401 10.6151
R8953 gnd.n5077 gnd.n1401 10.6151
R8954 gnd.n5078 gnd.n5077 10.6151
R8955 gnd.n5079 gnd.n5078 10.6151
R8956 gnd.n5079 gnd.n1388 10.6151
R8957 gnd.n5093 gnd.n1388 10.6151
R8958 gnd.n5094 gnd.n5093 10.6151
R8959 gnd.n5096 gnd.n5094 10.6151
R8960 gnd.n5096 gnd.n5095 10.6151
R8961 gnd.n5095 gnd.n1365 10.6151
R8962 gnd.n5127 gnd.n1365 10.6151
R8963 gnd.n5128 gnd.n5127 10.6151
R8964 gnd.n5130 gnd.n5128 10.6151
R8965 gnd.n5130 gnd.n5129 10.6151
R8966 gnd.n5129 gnd.n1336 10.6151
R8967 gnd.n5338 gnd.n1336 10.6151
R8968 gnd.n5339 gnd.n5338 10.6151
R8969 gnd.n5424 gnd.n5339 10.6151
R8970 gnd.n2830 gnd.t154 10.5161
R8971 gnd.n2287 gnd.t198 10.5161
R8972 gnd.n3197 gnd.t170 10.5161
R8973 gnd.n3950 gnd.t157 10.5161
R8974 gnd.t209 gnd.n3965 10.5161
R8975 gnd.n3973 gnd.t209 10.5161
R8976 gnd.n3998 gnd.t152 10.5161
R8977 gnd.t181 gnd.n5782 10.5161
R8978 gnd.n5810 gnd.t137 10.5161
R8979 gnd.t137 gnd.n235 10.5161
R8980 gnd.t8 gnd.n233 10.5161
R8981 gnd.n3473 gnd.n3457 10.4732
R8982 gnd.n3441 gnd.n3425 10.4732
R8983 gnd.n3409 gnd.n3393 10.4732
R8984 gnd.n3378 gnd.n3362 10.4732
R8985 gnd.n3346 gnd.n3330 10.4732
R8986 gnd.n3314 gnd.n3298 10.4732
R8987 gnd.n3282 gnd.n3266 10.4732
R8988 gnd.n3251 gnd.n3235 10.4732
R8989 gnd.n4444 gnd.n1760 10.1975
R8990 gnd.n4478 gnd.n1745 10.1975
R8991 gnd.n4618 gnd.n1671 10.1975
R8992 gnd.n4795 gnd.n1584 10.1975
R8993 gnd.n4828 gnd.n1567 10.1975
R8994 gnd.n5004 gnd.n5003 10.1975
R8995 gnd.n5124 gnd.n5123 10.1975
R8996 gnd.n1428 gnd.n1427 10.1975
R8997 gnd.n3902 gnd.t6 9.87883
R8998 gnd.n3895 gnd.t164 9.87883
R8999 gnd.n4024 gnd.t256 9.87883
R9000 gnd.n6034 gnd.t244 9.87883
R9001 gnd.t125 gnd.n1212 9.87883
R9002 gnd.t241 gnd.n5756 9.87883
R9003 gnd.n6956 gnd.t13 9.87883
R9004 gnd.t225 gnd.n196 9.87883
R9005 gnd.n3477 gnd.n3476 9.69747
R9006 gnd.n3445 gnd.n3444 9.69747
R9007 gnd.n3413 gnd.n3412 9.69747
R9008 gnd.n3382 gnd.n3381 9.69747
R9009 gnd.n3350 gnd.n3349 9.69747
R9010 gnd.n3318 gnd.n3317 9.69747
R9011 gnd.n3286 gnd.n3285 9.69747
R9012 gnd.n3255 gnd.n3254 9.69747
R9013 gnd.n7185 gnd.n50 9.6512
R9014 gnd.n4526 gnd.n1715 9.56018
R9015 gnd.n4563 gnd.n1699 9.56018
R9016 gnd.n4721 gnd.n1624 9.56018
R9017 gnd.n1626 gnd.t197 9.56018
R9018 gnd.n4749 gnd.n4748 9.56018
R9019 gnd.n4874 gnd.n1537 9.56018
R9020 gnd.n4913 gnd.t238 9.56018
R9021 gnd.n4911 gnd.n1518 9.56018
R9022 gnd.n5058 gnd.n1417 9.56018
R9023 gnd.n5082 gnd.n1397 9.56018
R9024 gnd.n5994 gnd.n999 9.45599
R9025 gnd.n5205 gnd.n5204 9.45599
R9026 gnd.n3483 gnd.n3482 9.45567
R9027 gnd.n3451 gnd.n3450 9.45567
R9028 gnd.n3419 gnd.n3418 9.45567
R9029 gnd.n3388 gnd.n3387 9.45567
R9030 gnd.n3356 gnd.n3355 9.45567
R9031 gnd.n3324 gnd.n3323 9.45567
R9032 gnd.n3292 gnd.n3291 9.45567
R9033 gnd.n3261 gnd.n3260 9.45567
R9034 gnd.n2428 gnd.n2427 9.39724
R9035 gnd.n3482 gnd.n3481 9.3005
R9036 gnd.n3455 gnd.n3454 9.3005
R9037 gnd.n3476 gnd.n3475 9.3005
R9038 gnd.n3474 gnd.n3473 9.3005
R9039 gnd.n3459 gnd.n3458 9.3005
R9040 gnd.n3468 gnd.n3467 9.3005
R9041 gnd.n3466 gnd.n3465 9.3005
R9042 gnd.n3450 gnd.n3449 9.3005
R9043 gnd.n3423 gnd.n3422 9.3005
R9044 gnd.n3444 gnd.n3443 9.3005
R9045 gnd.n3442 gnd.n3441 9.3005
R9046 gnd.n3427 gnd.n3426 9.3005
R9047 gnd.n3436 gnd.n3435 9.3005
R9048 gnd.n3434 gnd.n3433 9.3005
R9049 gnd.n3418 gnd.n3417 9.3005
R9050 gnd.n3391 gnd.n3390 9.3005
R9051 gnd.n3412 gnd.n3411 9.3005
R9052 gnd.n3410 gnd.n3409 9.3005
R9053 gnd.n3395 gnd.n3394 9.3005
R9054 gnd.n3404 gnd.n3403 9.3005
R9055 gnd.n3402 gnd.n3401 9.3005
R9056 gnd.n3387 gnd.n3386 9.3005
R9057 gnd.n3360 gnd.n3359 9.3005
R9058 gnd.n3381 gnd.n3380 9.3005
R9059 gnd.n3379 gnd.n3378 9.3005
R9060 gnd.n3364 gnd.n3363 9.3005
R9061 gnd.n3373 gnd.n3372 9.3005
R9062 gnd.n3371 gnd.n3370 9.3005
R9063 gnd.n3355 gnd.n3354 9.3005
R9064 gnd.n3328 gnd.n3327 9.3005
R9065 gnd.n3349 gnd.n3348 9.3005
R9066 gnd.n3347 gnd.n3346 9.3005
R9067 gnd.n3332 gnd.n3331 9.3005
R9068 gnd.n3341 gnd.n3340 9.3005
R9069 gnd.n3339 gnd.n3338 9.3005
R9070 gnd.n3323 gnd.n3322 9.3005
R9071 gnd.n3296 gnd.n3295 9.3005
R9072 gnd.n3317 gnd.n3316 9.3005
R9073 gnd.n3315 gnd.n3314 9.3005
R9074 gnd.n3300 gnd.n3299 9.3005
R9075 gnd.n3309 gnd.n3308 9.3005
R9076 gnd.n3307 gnd.n3306 9.3005
R9077 gnd.n3291 gnd.n3290 9.3005
R9078 gnd.n3264 gnd.n3263 9.3005
R9079 gnd.n3285 gnd.n3284 9.3005
R9080 gnd.n3283 gnd.n3282 9.3005
R9081 gnd.n3268 gnd.n3267 9.3005
R9082 gnd.n3277 gnd.n3276 9.3005
R9083 gnd.n3275 gnd.n3274 9.3005
R9084 gnd.n3260 gnd.n3259 9.3005
R9085 gnd.n3233 gnd.n3232 9.3005
R9086 gnd.n3254 gnd.n3253 9.3005
R9087 gnd.n3252 gnd.n3251 9.3005
R9088 gnd.n3237 gnd.n3236 9.3005
R9089 gnd.n3246 gnd.n3245 9.3005
R9090 gnd.n3244 gnd.n3243 9.3005
R9091 gnd.n3608 gnd.n3607 9.3005
R9092 gnd.n3606 gnd.n2187 9.3005
R9093 gnd.n3605 gnd.n3604 9.3005
R9094 gnd.n3601 gnd.n2188 9.3005
R9095 gnd.n3598 gnd.n2189 9.3005
R9096 gnd.n3597 gnd.n2190 9.3005
R9097 gnd.n3594 gnd.n2191 9.3005
R9098 gnd.n3593 gnd.n2192 9.3005
R9099 gnd.n3590 gnd.n2193 9.3005
R9100 gnd.n3589 gnd.n2194 9.3005
R9101 gnd.n3586 gnd.n2195 9.3005
R9102 gnd.n3585 gnd.n2196 9.3005
R9103 gnd.n3582 gnd.n2197 9.3005
R9104 gnd.n3581 gnd.n2198 9.3005
R9105 gnd.n3578 gnd.n3577 9.3005
R9106 gnd.n3576 gnd.n2199 9.3005
R9107 gnd.n3609 gnd.n2186 9.3005
R9108 gnd.n2849 gnd.n2848 9.3005
R9109 gnd.n2553 gnd.n2552 9.3005
R9110 gnd.n2876 gnd.n2875 9.3005
R9111 gnd.n2877 gnd.n2551 9.3005
R9112 gnd.n2881 gnd.n2878 9.3005
R9113 gnd.n2880 gnd.n2879 9.3005
R9114 gnd.n2525 gnd.n2524 9.3005
R9115 gnd.n2906 gnd.n2905 9.3005
R9116 gnd.n2907 gnd.n2523 9.3005
R9117 gnd.n2909 gnd.n2908 9.3005
R9118 gnd.n2503 gnd.n2502 9.3005
R9119 gnd.n2937 gnd.n2936 9.3005
R9120 gnd.n2938 gnd.n2501 9.3005
R9121 gnd.n2946 gnd.n2939 9.3005
R9122 gnd.n2945 gnd.n2940 9.3005
R9123 gnd.n2944 gnd.n2942 9.3005
R9124 gnd.n2941 gnd.n2450 9.3005
R9125 gnd.n2994 gnd.n2451 9.3005
R9126 gnd.n2993 gnd.n2452 9.3005
R9127 gnd.n2992 gnd.n2453 9.3005
R9128 gnd.n2472 gnd.n2454 9.3005
R9129 gnd.n2474 gnd.n2473 9.3005
R9130 gnd.n2384 gnd.n2383 9.3005
R9131 gnd.n3032 gnd.n3031 9.3005
R9132 gnd.n3033 gnd.n2382 9.3005
R9133 gnd.n3037 gnd.n3034 9.3005
R9134 gnd.n3036 gnd.n3035 9.3005
R9135 gnd.n2357 gnd.n2356 9.3005
R9136 gnd.n3072 gnd.n3071 9.3005
R9137 gnd.n3073 gnd.n2355 9.3005
R9138 gnd.n3077 gnd.n3074 9.3005
R9139 gnd.n3076 gnd.n3075 9.3005
R9140 gnd.n2330 gnd.n2329 9.3005
R9141 gnd.n3117 gnd.n3116 9.3005
R9142 gnd.n3118 gnd.n2328 9.3005
R9143 gnd.n3122 gnd.n3119 9.3005
R9144 gnd.n3121 gnd.n3120 9.3005
R9145 gnd.n2302 gnd.n2301 9.3005
R9146 gnd.n3158 gnd.n3157 9.3005
R9147 gnd.n3159 gnd.n2300 9.3005
R9148 gnd.n3163 gnd.n3160 9.3005
R9149 gnd.n3162 gnd.n3161 9.3005
R9150 gnd.n2275 gnd.n2274 9.3005
R9151 gnd.n3207 gnd.n3206 9.3005
R9152 gnd.n3208 gnd.n2273 9.3005
R9153 gnd.n3212 gnd.n3209 9.3005
R9154 gnd.n3211 gnd.n3210 9.3005
R9155 gnd.n2248 gnd.n2247 9.3005
R9156 gnd.n3501 gnd.n3500 9.3005
R9157 gnd.n3502 gnd.n2246 9.3005
R9158 gnd.n3508 gnd.n3503 9.3005
R9159 gnd.n3507 gnd.n3504 9.3005
R9160 gnd.n3506 gnd.n3505 9.3005
R9161 gnd.n2850 gnd.n2847 9.3005
R9162 gnd.n2632 gnd.n2591 9.3005
R9163 gnd.n2627 gnd.n2626 9.3005
R9164 gnd.n2625 gnd.n2592 9.3005
R9165 gnd.n2624 gnd.n2623 9.3005
R9166 gnd.n2620 gnd.n2593 9.3005
R9167 gnd.n2617 gnd.n2616 9.3005
R9168 gnd.n2615 gnd.n2594 9.3005
R9169 gnd.n2614 gnd.n2613 9.3005
R9170 gnd.n2610 gnd.n2595 9.3005
R9171 gnd.n2607 gnd.n2606 9.3005
R9172 gnd.n2605 gnd.n2596 9.3005
R9173 gnd.n2604 gnd.n2603 9.3005
R9174 gnd.n2600 gnd.n2598 9.3005
R9175 gnd.n2597 gnd.n2577 9.3005
R9176 gnd.n2844 gnd.n2576 9.3005
R9177 gnd.n2846 gnd.n2845 9.3005
R9178 gnd.n2634 gnd.n2633 9.3005
R9179 gnd.n2857 gnd.n2563 9.3005
R9180 gnd.n2864 gnd.n2564 9.3005
R9181 gnd.n2866 gnd.n2865 9.3005
R9182 gnd.n2867 gnd.n2544 9.3005
R9183 gnd.n2886 gnd.n2885 9.3005
R9184 gnd.n2888 gnd.n2536 9.3005
R9185 gnd.n2895 gnd.n2538 9.3005
R9186 gnd.n2896 gnd.n2533 9.3005
R9187 gnd.n2898 gnd.n2897 9.3005
R9188 gnd.n2534 gnd.n2519 9.3005
R9189 gnd.n2914 gnd.n2517 9.3005
R9190 gnd.n2918 gnd.n2917 9.3005
R9191 gnd.n2916 gnd.n2493 9.3005
R9192 gnd.n2953 gnd.n2492 9.3005
R9193 gnd.n2956 gnd.n2955 9.3005
R9194 gnd.n2489 gnd.n2488 9.3005
R9195 gnd.n2962 gnd.n2490 9.3005
R9196 gnd.n2964 gnd.n2963 9.3005
R9197 gnd.n2966 gnd.n2487 9.3005
R9198 gnd.n2969 gnd.n2968 9.3005
R9199 gnd.n2972 gnd.n2970 9.3005
R9200 gnd.n2974 gnd.n2973 9.3005
R9201 gnd.n2980 gnd.n2975 9.3005
R9202 gnd.n2979 gnd.n2978 9.3005
R9203 gnd.n2375 gnd.n2374 9.3005
R9204 gnd.n3046 gnd.n3045 9.3005
R9205 gnd.n3047 gnd.n2368 9.3005
R9206 gnd.n3055 gnd.n2367 9.3005
R9207 gnd.n3058 gnd.n3057 9.3005
R9208 gnd.n3060 gnd.n3059 9.3005
R9209 gnd.n3063 gnd.n2350 9.3005
R9210 gnd.n3061 gnd.n2348 9.3005
R9211 gnd.n3083 gnd.n2346 9.3005
R9212 gnd.n3085 gnd.n3084 9.3005
R9213 gnd.n2320 gnd.n2319 9.3005
R9214 gnd.n3131 gnd.n3130 9.3005
R9215 gnd.n3132 gnd.n2313 9.3005
R9216 gnd.n3141 gnd.n2312 9.3005
R9217 gnd.n3144 gnd.n3143 9.3005
R9218 gnd.n3146 gnd.n3145 9.3005
R9219 gnd.n3149 gnd.n2295 9.3005
R9220 gnd.n3147 gnd.n2293 9.3005
R9221 gnd.n3169 gnd.n2291 9.3005
R9222 gnd.n3171 gnd.n3170 9.3005
R9223 gnd.n2266 gnd.n2265 9.3005
R9224 gnd.n3221 gnd.n3220 9.3005
R9225 gnd.n3222 gnd.n2259 9.3005
R9226 gnd.n3230 gnd.n2258 9.3005
R9227 gnd.n3489 gnd.n3488 9.3005
R9228 gnd.n3491 gnd.n3490 9.3005
R9229 gnd.n3492 gnd.n2239 9.3005
R9230 gnd.n3516 gnd.n3515 9.3005
R9231 gnd.n2240 gnd.n2202 9.3005
R9232 gnd.n2855 gnd.n2854 9.3005
R9233 gnd.n3572 gnd.n2203 9.3005
R9234 gnd.n3571 gnd.n2205 9.3005
R9235 gnd.n3568 gnd.n2206 9.3005
R9236 gnd.n3567 gnd.n2207 9.3005
R9237 gnd.n3564 gnd.n2208 9.3005
R9238 gnd.n3563 gnd.n2209 9.3005
R9239 gnd.n3560 gnd.n2210 9.3005
R9240 gnd.n3559 gnd.n2211 9.3005
R9241 gnd.n3556 gnd.n2212 9.3005
R9242 gnd.n3555 gnd.n2213 9.3005
R9243 gnd.n3552 gnd.n2214 9.3005
R9244 gnd.n3551 gnd.n2215 9.3005
R9245 gnd.n3548 gnd.n2216 9.3005
R9246 gnd.n3547 gnd.n2217 9.3005
R9247 gnd.n3544 gnd.n2218 9.3005
R9248 gnd.n3543 gnd.n2219 9.3005
R9249 gnd.n3540 gnd.n2220 9.3005
R9250 gnd.n3539 gnd.n2221 9.3005
R9251 gnd.n3536 gnd.n2222 9.3005
R9252 gnd.n3535 gnd.n2223 9.3005
R9253 gnd.n3532 gnd.n2224 9.3005
R9254 gnd.n3531 gnd.n2225 9.3005
R9255 gnd.n3528 gnd.n2229 9.3005
R9256 gnd.n3527 gnd.n2230 9.3005
R9257 gnd.n3524 gnd.n2231 9.3005
R9258 gnd.n3523 gnd.n2232 9.3005
R9259 gnd.n3574 gnd.n3573 9.3005
R9260 gnd.n3024 gnd.n3008 9.3005
R9261 gnd.n3023 gnd.n3009 9.3005
R9262 gnd.n3022 gnd.n3010 9.3005
R9263 gnd.n3020 gnd.n3011 9.3005
R9264 gnd.n3019 gnd.n3012 9.3005
R9265 gnd.n3017 gnd.n3013 9.3005
R9266 gnd.n3016 gnd.n3014 9.3005
R9267 gnd.n2338 gnd.n2337 9.3005
R9268 gnd.n3093 gnd.n3092 9.3005
R9269 gnd.n3094 gnd.n2336 9.3005
R9270 gnd.n3111 gnd.n3095 9.3005
R9271 gnd.n3110 gnd.n3096 9.3005
R9272 gnd.n3109 gnd.n3097 9.3005
R9273 gnd.n3107 gnd.n3098 9.3005
R9274 gnd.n3106 gnd.n3099 9.3005
R9275 gnd.n3104 gnd.n3100 9.3005
R9276 gnd.n3103 gnd.n3101 9.3005
R9277 gnd.n2282 gnd.n2281 9.3005
R9278 gnd.n3179 gnd.n3178 9.3005
R9279 gnd.n3180 gnd.n2280 9.3005
R9280 gnd.n3201 gnd.n3181 9.3005
R9281 gnd.n3200 gnd.n3182 9.3005
R9282 gnd.n3199 gnd.n3183 9.3005
R9283 gnd.n3196 gnd.n3184 9.3005
R9284 gnd.n3195 gnd.n3185 9.3005
R9285 gnd.n3193 gnd.n3186 9.3005
R9286 gnd.n3192 gnd.n3187 9.3005
R9287 gnd.n3190 gnd.n3189 9.3005
R9288 gnd.n3188 gnd.n2234 9.3005
R9289 gnd.n2765 gnd.n2764 9.3005
R9290 gnd.n2655 gnd.n2654 9.3005
R9291 gnd.n2779 gnd.n2778 9.3005
R9292 gnd.n2780 gnd.n2653 9.3005
R9293 gnd.n2782 gnd.n2781 9.3005
R9294 gnd.n2643 gnd.n2642 9.3005
R9295 gnd.n2795 gnd.n2794 9.3005
R9296 gnd.n2796 gnd.n2641 9.3005
R9297 gnd.n2828 gnd.n2797 9.3005
R9298 gnd.n2827 gnd.n2798 9.3005
R9299 gnd.n2826 gnd.n2799 9.3005
R9300 gnd.n2825 gnd.n2800 9.3005
R9301 gnd.n2822 gnd.n2801 9.3005
R9302 gnd.n2821 gnd.n2802 9.3005
R9303 gnd.n2820 gnd.n2803 9.3005
R9304 gnd.n2818 gnd.n2804 9.3005
R9305 gnd.n2817 gnd.n2805 9.3005
R9306 gnd.n2814 gnd.n2806 9.3005
R9307 gnd.n2813 gnd.n2807 9.3005
R9308 gnd.n2812 gnd.n2808 9.3005
R9309 gnd.n2810 gnd.n2809 9.3005
R9310 gnd.n2509 gnd.n2508 9.3005
R9311 gnd.n2926 gnd.n2925 9.3005
R9312 gnd.n2927 gnd.n2507 9.3005
R9313 gnd.n2931 gnd.n2928 9.3005
R9314 gnd.n2930 gnd.n2929 9.3005
R9315 gnd.n2431 gnd.n2430 9.3005
R9316 gnd.n3006 gnd.n3005 9.3005
R9317 gnd.n2763 gnd.n2664 9.3005
R9318 gnd.n2666 gnd.n2665 9.3005
R9319 gnd.n2710 gnd.n2708 9.3005
R9320 gnd.n2711 gnd.n2707 9.3005
R9321 gnd.n2714 gnd.n2703 9.3005
R9322 gnd.n2715 gnd.n2702 9.3005
R9323 gnd.n2718 gnd.n2701 9.3005
R9324 gnd.n2719 gnd.n2700 9.3005
R9325 gnd.n2722 gnd.n2699 9.3005
R9326 gnd.n2723 gnd.n2698 9.3005
R9327 gnd.n2726 gnd.n2697 9.3005
R9328 gnd.n2727 gnd.n2696 9.3005
R9329 gnd.n2730 gnd.n2695 9.3005
R9330 gnd.n2731 gnd.n2694 9.3005
R9331 gnd.n2734 gnd.n2693 9.3005
R9332 gnd.n2735 gnd.n2692 9.3005
R9333 gnd.n2738 gnd.n2691 9.3005
R9334 gnd.n2739 gnd.n2690 9.3005
R9335 gnd.n2742 gnd.n2689 9.3005
R9336 gnd.n2743 gnd.n2688 9.3005
R9337 gnd.n2746 gnd.n2687 9.3005
R9338 gnd.n2747 gnd.n2686 9.3005
R9339 gnd.n2750 gnd.n2685 9.3005
R9340 gnd.n2752 gnd.n2684 9.3005
R9341 gnd.n2753 gnd.n2683 9.3005
R9342 gnd.n2754 gnd.n2682 9.3005
R9343 gnd.n2755 gnd.n2681 9.3005
R9344 gnd.n2762 gnd.n2761 9.3005
R9345 gnd.n2771 gnd.n2770 9.3005
R9346 gnd.n2772 gnd.n2658 9.3005
R9347 gnd.n2774 gnd.n2773 9.3005
R9348 gnd.n2649 gnd.n2648 9.3005
R9349 gnd.n2787 gnd.n2786 9.3005
R9350 gnd.n2788 gnd.n2647 9.3005
R9351 gnd.n2790 gnd.n2789 9.3005
R9352 gnd.n2636 gnd.n2635 9.3005
R9353 gnd.n2833 gnd.n2832 9.3005
R9354 gnd.n2834 gnd.n2590 9.3005
R9355 gnd.n2838 gnd.n2836 9.3005
R9356 gnd.n2837 gnd.n2569 9.3005
R9357 gnd.n2856 gnd.n2568 9.3005
R9358 gnd.n2859 gnd.n2858 9.3005
R9359 gnd.n2562 gnd.n2561 9.3005
R9360 gnd.n2870 gnd.n2868 9.3005
R9361 gnd.n2869 gnd.n2543 9.3005
R9362 gnd.n2887 gnd.n2542 9.3005
R9363 gnd.n2890 gnd.n2889 9.3005
R9364 gnd.n2537 gnd.n2532 9.3005
R9365 gnd.n2900 gnd.n2899 9.3005
R9366 gnd.n2535 gnd.n2515 9.3005
R9367 gnd.n2921 gnd.n2516 9.3005
R9368 gnd.n2920 gnd.n2919 9.3005
R9369 gnd.n2518 gnd.n2494 9.3005
R9370 gnd.n2952 gnd.n2951 9.3005
R9371 gnd.n2954 gnd.n2439 9.3005
R9372 gnd.n3001 gnd.n2440 9.3005
R9373 gnd.n3000 gnd.n2441 9.3005
R9374 gnd.n2999 gnd.n2442 9.3005
R9375 gnd.n2965 gnd.n2443 9.3005
R9376 gnd.n2967 gnd.n2461 9.3005
R9377 gnd.n2987 gnd.n2462 9.3005
R9378 gnd.n2986 gnd.n2463 9.3005
R9379 gnd.n2985 gnd.n2464 9.3005
R9380 gnd.n2976 gnd.n2465 9.3005
R9381 gnd.n2977 gnd.n2376 9.3005
R9382 gnd.n3043 gnd.n3042 9.3005
R9383 gnd.n3044 gnd.n2369 9.3005
R9384 gnd.n3054 gnd.n3053 9.3005
R9385 gnd.n3056 gnd.n2365 9.3005
R9386 gnd.n3066 gnd.n2366 9.3005
R9387 gnd.n3065 gnd.n3064 9.3005
R9388 gnd.n3062 gnd.n2344 9.3005
R9389 gnd.n3088 gnd.n2345 9.3005
R9390 gnd.n3087 gnd.n3086 9.3005
R9391 gnd.n2347 gnd.n2321 9.3005
R9392 gnd.n3128 gnd.n3127 9.3005
R9393 gnd.n3129 gnd.n2314 9.3005
R9394 gnd.n3140 gnd.n3139 9.3005
R9395 gnd.n3142 gnd.n2310 9.3005
R9396 gnd.n3152 gnd.n2311 9.3005
R9397 gnd.n3151 gnd.n3150 9.3005
R9398 gnd.n3148 gnd.n2289 9.3005
R9399 gnd.n3174 gnd.n2290 9.3005
R9400 gnd.n3173 gnd.n3172 9.3005
R9401 gnd.n2292 gnd.n2267 9.3005
R9402 gnd.n3218 gnd.n3217 9.3005
R9403 gnd.n3219 gnd.n2260 9.3005
R9404 gnd.n3229 gnd.n3228 9.3005
R9405 gnd.n3487 gnd.n2256 9.3005
R9406 gnd.n3495 gnd.n2257 9.3005
R9407 gnd.n3494 gnd.n3493 9.3005
R9408 gnd.n2238 gnd.n2237 9.3005
R9409 gnd.n3518 gnd.n3517 9.3005
R9410 gnd.n2660 gnd.n2659 9.3005
R9411 gnd.n6263 gnd.n657 9.3005
R9412 gnd.n6265 gnd.n6264 9.3005
R9413 gnd.n653 gnd.n652 9.3005
R9414 gnd.n6272 gnd.n6271 9.3005
R9415 gnd.n6273 gnd.n651 9.3005
R9416 gnd.n6275 gnd.n6274 9.3005
R9417 gnd.n647 gnd.n646 9.3005
R9418 gnd.n6282 gnd.n6281 9.3005
R9419 gnd.n6283 gnd.n645 9.3005
R9420 gnd.n6285 gnd.n6284 9.3005
R9421 gnd.n641 gnd.n640 9.3005
R9422 gnd.n6292 gnd.n6291 9.3005
R9423 gnd.n6293 gnd.n639 9.3005
R9424 gnd.n6295 gnd.n6294 9.3005
R9425 gnd.n635 gnd.n634 9.3005
R9426 gnd.n6302 gnd.n6301 9.3005
R9427 gnd.n6303 gnd.n633 9.3005
R9428 gnd.n6305 gnd.n6304 9.3005
R9429 gnd.n629 gnd.n628 9.3005
R9430 gnd.n6312 gnd.n6311 9.3005
R9431 gnd.n6313 gnd.n627 9.3005
R9432 gnd.n6315 gnd.n6314 9.3005
R9433 gnd.n623 gnd.n622 9.3005
R9434 gnd.n6322 gnd.n6321 9.3005
R9435 gnd.n6323 gnd.n621 9.3005
R9436 gnd.n6325 gnd.n6324 9.3005
R9437 gnd.n617 gnd.n616 9.3005
R9438 gnd.n6332 gnd.n6331 9.3005
R9439 gnd.n6333 gnd.n615 9.3005
R9440 gnd.n6335 gnd.n6334 9.3005
R9441 gnd.n611 gnd.n610 9.3005
R9442 gnd.n6342 gnd.n6341 9.3005
R9443 gnd.n6343 gnd.n609 9.3005
R9444 gnd.n6345 gnd.n6344 9.3005
R9445 gnd.n605 gnd.n604 9.3005
R9446 gnd.n6352 gnd.n6351 9.3005
R9447 gnd.n6353 gnd.n603 9.3005
R9448 gnd.n6355 gnd.n6354 9.3005
R9449 gnd.n599 gnd.n598 9.3005
R9450 gnd.n6362 gnd.n6361 9.3005
R9451 gnd.n6363 gnd.n597 9.3005
R9452 gnd.n6365 gnd.n6364 9.3005
R9453 gnd.n593 gnd.n592 9.3005
R9454 gnd.n6372 gnd.n6371 9.3005
R9455 gnd.n6373 gnd.n591 9.3005
R9456 gnd.n6375 gnd.n6374 9.3005
R9457 gnd.n587 gnd.n586 9.3005
R9458 gnd.n6382 gnd.n6381 9.3005
R9459 gnd.n6383 gnd.n585 9.3005
R9460 gnd.n6385 gnd.n6384 9.3005
R9461 gnd.n581 gnd.n580 9.3005
R9462 gnd.n6392 gnd.n6391 9.3005
R9463 gnd.n6393 gnd.n579 9.3005
R9464 gnd.n6395 gnd.n6394 9.3005
R9465 gnd.n575 gnd.n574 9.3005
R9466 gnd.n6402 gnd.n6401 9.3005
R9467 gnd.n6403 gnd.n573 9.3005
R9468 gnd.n6405 gnd.n6404 9.3005
R9469 gnd.n569 gnd.n568 9.3005
R9470 gnd.n6412 gnd.n6411 9.3005
R9471 gnd.n6413 gnd.n567 9.3005
R9472 gnd.n6415 gnd.n6414 9.3005
R9473 gnd.n563 gnd.n562 9.3005
R9474 gnd.n6422 gnd.n6421 9.3005
R9475 gnd.n6423 gnd.n561 9.3005
R9476 gnd.n6425 gnd.n6424 9.3005
R9477 gnd.n557 gnd.n556 9.3005
R9478 gnd.n6432 gnd.n6431 9.3005
R9479 gnd.n6433 gnd.n555 9.3005
R9480 gnd.n6435 gnd.n6434 9.3005
R9481 gnd.n551 gnd.n550 9.3005
R9482 gnd.n6442 gnd.n6441 9.3005
R9483 gnd.n6443 gnd.n549 9.3005
R9484 gnd.n6445 gnd.n6444 9.3005
R9485 gnd.n545 gnd.n544 9.3005
R9486 gnd.n6452 gnd.n6451 9.3005
R9487 gnd.n6453 gnd.n543 9.3005
R9488 gnd.n6455 gnd.n6454 9.3005
R9489 gnd.n539 gnd.n538 9.3005
R9490 gnd.n6462 gnd.n6461 9.3005
R9491 gnd.n6463 gnd.n537 9.3005
R9492 gnd.n6465 gnd.n6464 9.3005
R9493 gnd.n533 gnd.n532 9.3005
R9494 gnd.n6472 gnd.n6471 9.3005
R9495 gnd.n6473 gnd.n531 9.3005
R9496 gnd.n6475 gnd.n6474 9.3005
R9497 gnd.n527 gnd.n526 9.3005
R9498 gnd.n6482 gnd.n6481 9.3005
R9499 gnd.n6483 gnd.n525 9.3005
R9500 gnd.n6485 gnd.n6484 9.3005
R9501 gnd.n521 gnd.n520 9.3005
R9502 gnd.n6492 gnd.n6491 9.3005
R9503 gnd.n6493 gnd.n519 9.3005
R9504 gnd.n6495 gnd.n6494 9.3005
R9505 gnd.n515 gnd.n514 9.3005
R9506 gnd.n6502 gnd.n6501 9.3005
R9507 gnd.n6503 gnd.n513 9.3005
R9508 gnd.n6505 gnd.n6504 9.3005
R9509 gnd.n509 gnd.n508 9.3005
R9510 gnd.n6512 gnd.n6511 9.3005
R9511 gnd.n6513 gnd.n507 9.3005
R9512 gnd.n6515 gnd.n6514 9.3005
R9513 gnd.n503 gnd.n502 9.3005
R9514 gnd.n6522 gnd.n6521 9.3005
R9515 gnd.n6523 gnd.n501 9.3005
R9516 gnd.n6525 gnd.n6524 9.3005
R9517 gnd.n497 gnd.n496 9.3005
R9518 gnd.n6532 gnd.n6531 9.3005
R9519 gnd.n6533 gnd.n495 9.3005
R9520 gnd.n6535 gnd.n6534 9.3005
R9521 gnd.n491 gnd.n490 9.3005
R9522 gnd.n6542 gnd.n6541 9.3005
R9523 gnd.n6543 gnd.n489 9.3005
R9524 gnd.n6545 gnd.n6544 9.3005
R9525 gnd.n485 gnd.n484 9.3005
R9526 gnd.n6552 gnd.n6551 9.3005
R9527 gnd.n6553 gnd.n483 9.3005
R9528 gnd.n6555 gnd.n6554 9.3005
R9529 gnd.n479 gnd.n478 9.3005
R9530 gnd.n6562 gnd.n6561 9.3005
R9531 gnd.n6563 gnd.n477 9.3005
R9532 gnd.n6565 gnd.n6564 9.3005
R9533 gnd.n473 gnd.n472 9.3005
R9534 gnd.n6572 gnd.n6571 9.3005
R9535 gnd.n6573 gnd.n471 9.3005
R9536 gnd.n6575 gnd.n6574 9.3005
R9537 gnd.n467 gnd.n466 9.3005
R9538 gnd.n6582 gnd.n6581 9.3005
R9539 gnd.n6583 gnd.n465 9.3005
R9540 gnd.n6585 gnd.n6584 9.3005
R9541 gnd.n461 gnd.n460 9.3005
R9542 gnd.n6592 gnd.n6591 9.3005
R9543 gnd.n6593 gnd.n459 9.3005
R9544 gnd.n6595 gnd.n6594 9.3005
R9545 gnd.n455 gnd.n454 9.3005
R9546 gnd.n6602 gnd.n6601 9.3005
R9547 gnd.n6603 gnd.n453 9.3005
R9548 gnd.n6605 gnd.n6604 9.3005
R9549 gnd.n449 gnd.n448 9.3005
R9550 gnd.n6612 gnd.n6611 9.3005
R9551 gnd.n6613 gnd.n447 9.3005
R9552 gnd.n6615 gnd.n6614 9.3005
R9553 gnd.n443 gnd.n442 9.3005
R9554 gnd.n6622 gnd.n6621 9.3005
R9555 gnd.n6623 gnd.n441 9.3005
R9556 gnd.n6625 gnd.n6624 9.3005
R9557 gnd.n437 gnd.n436 9.3005
R9558 gnd.n6632 gnd.n6631 9.3005
R9559 gnd.n6633 gnd.n435 9.3005
R9560 gnd.n6635 gnd.n6634 9.3005
R9561 gnd.n431 gnd.n430 9.3005
R9562 gnd.n6642 gnd.n6641 9.3005
R9563 gnd.n6643 gnd.n429 9.3005
R9564 gnd.n6645 gnd.n6644 9.3005
R9565 gnd.n425 gnd.n424 9.3005
R9566 gnd.n6652 gnd.n6651 9.3005
R9567 gnd.n6653 gnd.n423 9.3005
R9568 gnd.n6655 gnd.n6654 9.3005
R9569 gnd.n419 gnd.n418 9.3005
R9570 gnd.n6662 gnd.n6661 9.3005
R9571 gnd.n6663 gnd.n417 9.3005
R9572 gnd.n6665 gnd.n6664 9.3005
R9573 gnd.n413 gnd.n412 9.3005
R9574 gnd.n6672 gnd.n6671 9.3005
R9575 gnd.n6673 gnd.n411 9.3005
R9576 gnd.n6675 gnd.n6674 9.3005
R9577 gnd.n407 gnd.n406 9.3005
R9578 gnd.n6682 gnd.n6681 9.3005
R9579 gnd.n6685 gnd.n6684 9.3005
R9580 gnd.n401 gnd.n400 9.3005
R9581 gnd.n6692 gnd.n6691 9.3005
R9582 gnd.n6693 gnd.n399 9.3005
R9583 gnd.n6695 gnd.n6694 9.3005
R9584 gnd.n395 gnd.n394 9.3005
R9585 gnd.n6702 gnd.n6701 9.3005
R9586 gnd.n6703 gnd.n393 9.3005
R9587 gnd.n6705 gnd.n6704 9.3005
R9588 gnd.n389 gnd.n388 9.3005
R9589 gnd.n6712 gnd.n6711 9.3005
R9590 gnd.n6713 gnd.n387 9.3005
R9591 gnd.n6715 gnd.n6714 9.3005
R9592 gnd.n383 gnd.n382 9.3005
R9593 gnd.n6722 gnd.n6721 9.3005
R9594 gnd.n6723 gnd.n381 9.3005
R9595 gnd.n6725 gnd.n6724 9.3005
R9596 gnd.n377 gnd.n376 9.3005
R9597 gnd.n6732 gnd.n6731 9.3005
R9598 gnd.n6733 gnd.n375 9.3005
R9599 gnd.n6735 gnd.n6734 9.3005
R9600 gnd.n371 gnd.n370 9.3005
R9601 gnd.n6742 gnd.n6741 9.3005
R9602 gnd.n6743 gnd.n369 9.3005
R9603 gnd.n6745 gnd.n6744 9.3005
R9604 gnd.n365 gnd.n364 9.3005
R9605 gnd.n6752 gnd.n6751 9.3005
R9606 gnd.n6753 gnd.n363 9.3005
R9607 gnd.n6755 gnd.n6754 9.3005
R9608 gnd.n359 gnd.n358 9.3005
R9609 gnd.n6762 gnd.n6761 9.3005
R9610 gnd.n6763 gnd.n357 9.3005
R9611 gnd.n6765 gnd.n6764 9.3005
R9612 gnd.n353 gnd.n352 9.3005
R9613 gnd.n6772 gnd.n6771 9.3005
R9614 gnd.n6773 gnd.n351 9.3005
R9615 gnd.n6775 gnd.n6774 9.3005
R9616 gnd.n347 gnd.n346 9.3005
R9617 gnd.n6782 gnd.n6781 9.3005
R9618 gnd.n6783 gnd.n345 9.3005
R9619 gnd.n6785 gnd.n6784 9.3005
R9620 gnd.n341 gnd.n340 9.3005
R9621 gnd.n6792 gnd.n6791 9.3005
R9622 gnd.n6793 gnd.n339 9.3005
R9623 gnd.n6795 gnd.n6794 9.3005
R9624 gnd.n335 gnd.n334 9.3005
R9625 gnd.n6802 gnd.n6801 9.3005
R9626 gnd.n6803 gnd.n333 9.3005
R9627 gnd.n6805 gnd.n6804 9.3005
R9628 gnd.n329 gnd.n328 9.3005
R9629 gnd.n6812 gnd.n6811 9.3005
R9630 gnd.n6813 gnd.n327 9.3005
R9631 gnd.n6815 gnd.n6814 9.3005
R9632 gnd.n323 gnd.n322 9.3005
R9633 gnd.n6822 gnd.n6821 9.3005
R9634 gnd.n6823 gnd.n321 9.3005
R9635 gnd.n6825 gnd.n6824 9.3005
R9636 gnd.n317 gnd.n316 9.3005
R9637 gnd.n6832 gnd.n6831 9.3005
R9638 gnd.n6833 gnd.n315 9.3005
R9639 gnd.n6835 gnd.n6834 9.3005
R9640 gnd.n311 gnd.n310 9.3005
R9641 gnd.n6842 gnd.n6841 9.3005
R9642 gnd.n6843 gnd.n309 9.3005
R9643 gnd.n6845 gnd.n6844 9.3005
R9644 gnd.n305 gnd.n304 9.3005
R9645 gnd.n6852 gnd.n6851 9.3005
R9646 gnd.n6853 gnd.n303 9.3005
R9647 gnd.n6855 gnd.n6854 9.3005
R9648 gnd.n299 gnd.n298 9.3005
R9649 gnd.n6862 gnd.n6861 9.3005
R9650 gnd.n6863 gnd.n297 9.3005
R9651 gnd.n6865 gnd.n6864 9.3005
R9652 gnd.n293 gnd.n292 9.3005
R9653 gnd.n6872 gnd.n6871 9.3005
R9654 gnd.n6873 gnd.n291 9.3005
R9655 gnd.n6875 gnd.n6874 9.3005
R9656 gnd.n287 gnd.n286 9.3005
R9657 gnd.n6882 gnd.n6881 9.3005
R9658 gnd.n6883 gnd.n285 9.3005
R9659 gnd.n6887 gnd.n6884 9.3005
R9660 gnd.n6886 gnd.n6885 9.3005
R9661 gnd.n281 gnd.n280 9.3005
R9662 gnd.n6895 gnd.n6894 9.3005
R9663 gnd.n6683 gnd.n405 9.3005
R9664 gnd.n7144 gnd.n89 9.3005
R9665 gnd.n7143 gnd.n91 9.3005
R9666 gnd.n95 gnd.n92 9.3005
R9667 gnd.n7138 gnd.n96 9.3005
R9668 gnd.n7137 gnd.n97 9.3005
R9669 gnd.n7136 gnd.n98 9.3005
R9670 gnd.n102 gnd.n99 9.3005
R9671 gnd.n7131 gnd.n103 9.3005
R9672 gnd.n7130 gnd.n104 9.3005
R9673 gnd.n7129 gnd.n105 9.3005
R9674 gnd.n109 gnd.n106 9.3005
R9675 gnd.n7124 gnd.n110 9.3005
R9676 gnd.n7123 gnd.n111 9.3005
R9677 gnd.n7122 gnd.n112 9.3005
R9678 gnd.n116 gnd.n113 9.3005
R9679 gnd.n7117 gnd.n117 9.3005
R9680 gnd.n7116 gnd.n118 9.3005
R9681 gnd.n7112 gnd.n119 9.3005
R9682 gnd.n123 gnd.n120 9.3005
R9683 gnd.n7107 gnd.n124 9.3005
R9684 gnd.n7106 gnd.n125 9.3005
R9685 gnd.n7105 gnd.n126 9.3005
R9686 gnd.n130 gnd.n127 9.3005
R9687 gnd.n7100 gnd.n131 9.3005
R9688 gnd.n7099 gnd.n132 9.3005
R9689 gnd.n7098 gnd.n133 9.3005
R9690 gnd.n137 gnd.n134 9.3005
R9691 gnd.n7093 gnd.n138 9.3005
R9692 gnd.n7092 gnd.n139 9.3005
R9693 gnd.n7091 gnd.n140 9.3005
R9694 gnd.n144 gnd.n141 9.3005
R9695 gnd.n7086 gnd.n145 9.3005
R9696 gnd.n7085 gnd.n146 9.3005
R9697 gnd.n7084 gnd.n147 9.3005
R9698 gnd.n151 gnd.n148 9.3005
R9699 gnd.n7079 gnd.n152 9.3005
R9700 gnd.n7078 gnd.n7077 9.3005
R9701 gnd.n7076 gnd.n155 9.3005
R9702 gnd.n7146 gnd.n7145 9.3005
R9703 gnd.n5610 gnd.n5609 9.3005
R9704 gnd.n1261 gnd.n1260 9.3005
R9705 gnd.n5624 gnd.n5623 9.3005
R9706 gnd.n5625 gnd.n1259 9.3005
R9707 gnd.n5668 gnd.n5626 9.3005
R9708 gnd.n5667 gnd.n5627 9.3005
R9709 gnd.n5666 gnd.n5628 9.3005
R9710 gnd.n5664 gnd.n5629 9.3005
R9711 gnd.n5663 gnd.n5630 9.3005
R9712 gnd.n5662 gnd.n5631 9.3005
R9713 gnd.n5660 gnd.n5632 9.3005
R9714 gnd.n5659 gnd.n5633 9.3005
R9715 gnd.n5657 gnd.n5634 9.3005
R9716 gnd.n5656 gnd.n5635 9.3005
R9717 gnd.n5655 gnd.n5636 9.3005
R9718 gnd.n5653 gnd.n5637 9.3005
R9719 gnd.n5652 gnd.n5638 9.3005
R9720 gnd.n5649 gnd.n5639 9.3005
R9721 gnd.n5648 gnd.n5640 9.3005
R9722 gnd.n5646 gnd.n5641 9.3005
R9723 gnd.n5645 gnd.n5643 9.3005
R9724 gnd.n5642 gnd.n237 9.3005
R9725 gnd.n6925 gnd.n238 9.3005
R9726 gnd.n6924 gnd.n239 9.3005
R9727 gnd.n6923 gnd.n240 9.3005
R9728 gnd.n6919 gnd.n241 9.3005
R9729 gnd.n6918 gnd.n242 9.3005
R9730 gnd.n6915 gnd.n243 9.3005
R9731 gnd.n6914 gnd.n244 9.3005
R9732 gnd.n6910 gnd.n245 9.3005
R9733 gnd.n6909 gnd.n246 9.3005
R9734 gnd.n269 gnd.n247 9.3005
R9735 gnd.n268 gnd.n248 9.3005
R9736 gnd.n264 gnd.n249 9.3005
R9737 gnd.n263 gnd.n250 9.3005
R9738 gnd.n260 gnd.n251 9.3005
R9739 gnd.n259 gnd.n252 9.3005
R9740 gnd.n257 gnd.n253 9.3005
R9741 gnd.n256 gnd.n255 9.3005
R9742 gnd.n254 gnd.n159 9.3005
R9743 gnd.n7073 gnd.n158 9.3005
R9744 gnd.n7075 gnd.n7074 9.3005
R9745 gnd.n5608 gnd.n1266 9.3005
R9746 gnd.n5597 gnd.n1271 9.3005
R9747 gnd.n5599 gnd.n5598 9.3005
R9748 gnd.n5596 gnd.n1273 9.3005
R9749 gnd.n5595 gnd.n5594 9.3005
R9750 gnd.n1275 gnd.n1274 9.3005
R9751 gnd.n5588 gnd.n5587 9.3005
R9752 gnd.n5586 gnd.n1277 9.3005
R9753 gnd.n5585 gnd.n5584 9.3005
R9754 gnd.n1279 gnd.n1278 9.3005
R9755 gnd.n5578 gnd.n5577 9.3005
R9756 gnd.n5576 gnd.n1281 9.3005
R9757 gnd.n5575 gnd.n5574 9.3005
R9758 gnd.n1283 gnd.n1282 9.3005
R9759 gnd.n5568 gnd.n5567 9.3005
R9760 gnd.n5566 gnd.n1285 9.3005
R9761 gnd.n5565 gnd.n5564 9.3005
R9762 gnd.n1287 gnd.n1286 9.3005
R9763 gnd.n5558 gnd.n5557 9.3005
R9764 gnd.n5556 gnd.n1289 9.3005
R9765 gnd.n1291 gnd.n1290 9.3005
R9766 gnd.n5543 gnd.n5498 9.3005
R9767 gnd.n5545 gnd.n5544 9.3005
R9768 gnd.n5542 gnd.n5500 9.3005
R9769 gnd.n5541 gnd.n5540 9.3005
R9770 gnd.n5502 gnd.n5501 9.3005
R9771 gnd.n5534 gnd.n5533 9.3005
R9772 gnd.n5532 gnd.n5504 9.3005
R9773 gnd.n5531 gnd.n5530 9.3005
R9774 gnd.n5506 gnd.n5505 9.3005
R9775 gnd.n5524 gnd.n5523 9.3005
R9776 gnd.n5522 gnd.n5508 9.3005
R9777 gnd.n5521 gnd.n5520 9.3005
R9778 gnd.n5510 gnd.n5509 9.3005
R9779 gnd.n5514 gnd.n5513 9.3005
R9780 gnd.n5512 gnd.n5511 9.3005
R9781 gnd.n1270 gnd.n1267 9.3005
R9782 gnd.n5607 gnd.n5606 9.3005
R9783 gnd.n5848 gnd.n1134 9.3005
R9784 gnd.n5847 gnd.n1135 9.3005
R9785 gnd.n1255 gnd.n1136 9.3005
R9786 gnd.n5691 gnd.n5690 9.3005
R9787 gnd.n5692 gnd.n1254 9.3005
R9788 gnd.n5696 gnd.n5693 9.3005
R9789 gnd.n5695 gnd.n5694 9.3005
R9790 gnd.n1228 gnd.n1227 9.3005
R9791 gnd.n5722 gnd.n5721 9.3005
R9792 gnd.n5723 gnd.n1226 9.3005
R9793 gnd.n5728 gnd.n5724 9.3005
R9794 gnd.n5727 gnd.n5726 9.3005
R9795 gnd.n5725 gnd.n1198 9.3005
R9796 gnd.n5759 gnd.n1199 9.3005
R9797 gnd.n5760 gnd.n214 9.3005
R9798 gnd.n6944 gnd.n213 9.3005
R9799 gnd.n6946 gnd.n6945 9.3005
R9800 gnd.n200 gnd.n199 9.3005
R9801 gnd.n6959 gnd.n6958 9.3005
R9802 gnd.n6960 gnd.n198 9.3005
R9803 gnd.n6962 gnd.n6961 9.3005
R9804 gnd.n184 gnd.n183 9.3005
R9805 gnd.n6975 gnd.n6974 9.3005
R9806 gnd.n6976 gnd.n182 9.3005
R9807 gnd.n6978 gnd.n6977 9.3005
R9808 gnd.n166 gnd.n165 9.3005
R9809 gnd.n7065 gnd.n7064 9.3005
R9810 gnd.n7066 gnd.n164 9.3005
R9811 gnd.n7068 gnd.n7067 9.3005
R9812 gnd.n88 gnd.n87 9.3005
R9813 gnd.n7148 gnd.n7147 9.3005
R9814 gnd.n5849 gnd.n1133 9.3005
R9815 gnd.n6943 gnd.n6942 9.3005
R9816 gnd.n4018 gnd.n4017 9.3005
R9817 gnd.n4022 gnd.n4019 9.3005
R9818 gnd.n4021 gnd.n4020 9.3005
R9819 gnd.n2042 gnd.n2041 9.3005
R9820 gnd.n4082 gnd.n4081 9.3005
R9821 gnd.n4083 gnd.n2040 9.3005
R9822 gnd.n4085 gnd.n4084 9.3005
R9823 gnd.n2038 gnd.n2037 9.3005
R9824 gnd.n4090 gnd.n4089 9.3005
R9825 gnd.n4091 gnd.n2036 9.3005
R9826 gnd.n4093 gnd.n4092 9.3005
R9827 gnd.n2034 gnd.n2033 9.3005
R9828 gnd.n4098 gnd.n4097 9.3005
R9829 gnd.n4099 gnd.n2032 9.3005
R9830 gnd.n4101 gnd.n4100 9.3005
R9831 gnd.n2030 gnd.n2029 9.3005
R9832 gnd.n4106 gnd.n4105 9.3005
R9833 gnd.n4107 gnd.n2028 9.3005
R9834 gnd.n4109 gnd.n4108 9.3005
R9835 gnd.n2024 gnd.n2023 9.3005
R9836 gnd.n4248 gnd.n4247 9.3005
R9837 gnd.n4249 gnd.n2022 9.3005
R9838 gnd.n4251 gnd.n4250 9.3005
R9839 gnd.n1771 gnd.n1770 9.3005
R9840 gnd.n4417 gnd.n4416 9.3005
R9841 gnd.n4418 gnd.n1769 9.3005
R9842 gnd.n4420 gnd.n4419 9.3005
R9843 gnd.n1756 gnd.n1755 9.3005
R9844 gnd.n4462 gnd.n4461 9.3005
R9845 gnd.n4463 gnd.n1754 9.3005
R9846 gnd.n4467 gnd.n4464 9.3005
R9847 gnd.n4466 gnd.n4465 9.3005
R9848 gnd.n1728 gnd.n1727 9.3005
R9849 gnd.n4513 gnd.n4512 9.3005
R9850 gnd.n4514 gnd.n1726 9.3005
R9851 gnd.n4516 gnd.n4515 9.3005
R9852 gnd.n1708 gnd.n1707 9.3005
R9853 gnd.n4550 gnd.n4549 9.3005
R9854 gnd.n4551 gnd.n1706 9.3005
R9855 gnd.n4553 gnd.n4552 9.3005
R9856 gnd.n1682 gnd.n1681 9.3005
R9857 gnd.n4591 gnd.n4590 9.3005
R9858 gnd.n4592 gnd.n1680 9.3005
R9859 gnd.n4594 gnd.n4593 9.3005
R9860 gnd.n1666 gnd.n1665 9.3005
R9861 gnd.n4636 gnd.n4635 9.3005
R9862 gnd.n4637 gnd.n1664 9.3005
R9863 gnd.n4641 gnd.n4638 9.3005
R9864 gnd.n4640 gnd.n4639 9.3005
R9865 gnd.n1638 gnd.n1637 9.3005
R9866 gnd.n4708 gnd.n4707 9.3005
R9867 gnd.n4709 gnd.n1636 9.3005
R9868 gnd.n4711 gnd.n4710 9.3005
R9869 gnd.n1617 gnd.n1616 9.3005
R9870 gnd.n4735 gnd.n4734 9.3005
R9871 gnd.n4736 gnd.n1615 9.3005
R9872 gnd.n4738 gnd.n4737 9.3005
R9873 gnd.n1596 gnd.n1595 9.3005
R9874 gnd.n4768 gnd.n4767 9.3005
R9875 gnd.n4769 gnd.n1594 9.3005
R9876 gnd.n4771 gnd.n4770 9.3005
R9877 gnd.n1579 gnd.n1578 9.3005
R9878 gnd.n4813 gnd.n4812 9.3005
R9879 gnd.n4814 gnd.n1577 9.3005
R9880 gnd.n4818 gnd.n4815 9.3005
R9881 gnd.n4817 gnd.n4816 9.3005
R9882 gnd.n1550 gnd.n1549 9.3005
R9883 gnd.n4861 gnd.n4860 9.3005
R9884 gnd.n4862 gnd.n1548 9.3005
R9885 gnd.n4864 gnd.n4863 9.3005
R9886 gnd.n1530 gnd.n1529 9.3005
R9887 gnd.n4889 gnd.n4888 9.3005
R9888 gnd.n4890 gnd.n1528 9.3005
R9889 gnd.n4900 gnd.n4891 9.3005
R9890 gnd.n4899 gnd.n4892 9.3005
R9891 gnd.n4898 gnd.n4893 9.3005
R9892 gnd.n1498 gnd.n1497 9.3005
R9893 gnd.n4964 gnd.n4963 9.3005
R9894 gnd.n4965 gnd.n1496 9.3005
R9895 gnd.n4969 gnd.n4966 9.3005
R9896 gnd.n4968 gnd.n4967 9.3005
R9897 gnd.n1470 gnd.n1469 9.3005
R9898 gnd.n5015 gnd.n5014 9.3005
R9899 gnd.n5016 gnd.n1468 9.3005
R9900 gnd.n5020 gnd.n5017 9.3005
R9901 gnd.n5019 gnd.n5018 9.3005
R9902 gnd.n1452 gnd.n1451 9.3005
R9903 gnd.n5042 gnd.n5041 9.3005
R9904 gnd.n5043 gnd.n1450 9.3005
R9905 gnd.n5045 gnd.n5044 9.3005
R9906 gnd.n1395 gnd.n1394 9.3005
R9907 gnd.n5085 gnd.n5084 9.3005
R9908 gnd.n5086 gnd.n1393 9.3005
R9909 gnd.n5088 gnd.n5087 9.3005
R9910 gnd.n1374 gnd.n1373 9.3005
R9911 gnd.n5114 gnd.n5113 9.3005
R9912 gnd.n5115 gnd.n1372 9.3005
R9913 gnd.n5120 gnd.n5116 9.3005
R9914 gnd.n5119 gnd.n5118 9.3005
R9915 gnd.n5117 gnd.n1343 9.3005
R9916 gnd.n5333 gnd.n1344 9.3005
R9917 gnd.n5332 gnd.n1345 9.3005
R9918 gnd.n5331 gnd.n1346 9.3005
R9919 gnd.n1349 gnd.n1348 9.3005
R9920 gnd.n1347 gnd.n1111 9.3005
R9921 gnd.n5864 gnd.n1112 9.3005
R9922 gnd.n5863 gnd.n1113 9.3005
R9923 gnd.n5862 gnd.n1114 9.3005
R9924 gnd.n1120 gnd.n1115 9.3005
R9925 gnd.n5856 gnd.n1121 9.3005
R9926 gnd.n5855 gnd.n1122 9.3005
R9927 gnd.n5854 gnd.n1123 9.3005
R9928 gnd.n5674 gnd.n1124 9.3005
R9929 gnd.n5676 gnd.n5675 9.3005
R9930 gnd.n5680 gnd.n5679 9.3005
R9931 gnd.n5681 gnd.n5673 9.3005
R9932 gnd.n5685 gnd.n5682 9.3005
R9933 gnd.n5684 gnd.n5683 9.3005
R9934 gnd.n1238 gnd.n1237 9.3005
R9935 gnd.n5711 gnd.n5710 9.3005
R9936 gnd.n5712 gnd.n1236 9.3005
R9937 gnd.n5716 gnd.n5713 9.3005
R9938 gnd.n5715 gnd.n5714 9.3005
R9939 gnd.n1210 gnd.n1209 9.3005
R9940 gnd.n5743 gnd.n5742 9.3005
R9941 gnd.n5744 gnd.n1208 9.3005
R9942 gnd.n5754 gnd.n5745 9.3005
R9943 gnd.n5753 gnd.n5746 9.3005
R9944 gnd.n5799 gnd.n5791 9.3005
R9945 gnd.n5798 gnd.n5792 9.3005
R9946 gnd.n5795 gnd.n5794 9.3005
R9947 gnd.n5793 gnd.n272 9.3005
R9948 gnd.n6904 gnd.n273 9.3005
R9949 gnd.n6903 gnd.n274 9.3005
R9950 gnd.n6902 gnd.n275 9.3005
R9951 gnd.n278 gnd.n276 9.3005
R9952 gnd.n6898 gnd.n279 9.3005
R9953 gnd.n6897 gnd.n6896 9.3005
R9954 gnd.n3982 gnd.n3981 9.3005
R9955 gnd.n3693 gnd.n3689 9.3005
R9956 gnd.n3692 gnd.n3691 9.3005
R9957 gnd.n3690 gnd.n2140 9.3005
R9958 gnd.n3871 gnd.n2141 9.3005
R9959 gnd.n3872 gnd.n2139 9.3005
R9960 gnd.n3875 gnd.n3874 9.3005
R9961 gnd.n3876 gnd.n2138 9.3005
R9962 gnd.n3879 gnd.n3878 9.3005
R9963 gnd.n3877 gnd.n2130 9.3005
R9964 gnd.n3899 gnd.n2131 9.3005
R9965 gnd.n3898 gnd.n2132 9.3005
R9966 gnd.n3897 gnd.n2133 9.3005
R9967 gnd.n2122 gnd.n2121 9.3005
R9968 gnd.n3932 gnd.n3931 9.3005
R9969 gnd.n3933 gnd.n2120 9.3005
R9970 gnd.n3937 gnd.n3934 9.3005
R9971 gnd.n3936 gnd.n3935 9.3005
R9972 gnd.n2109 gnd.n2108 9.3005
R9973 gnd.n3979 gnd.n3978 9.3005
R9974 gnd.n3980 gnd.n2107 9.3005
R9975 gnd.n3695 gnd.n3694 9.3005
R9976 gnd.n3687 gnd.n3686 9.3005
R9977 gnd.n3683 gnd.n3643 9.3005
R9978 gnd.n3682 gnd.n3679 9.3005
R9979 gnd.n3678 gnd.n3644 9.3005
R9980 gnd.n3677 gnd.n3676 9.3005
R9981 gnd.n3673 gnd.n3645 9.3005
R9982 gnd.n3672 gnd.n3669 9.3005
R9983 gnd.n3668 gnd.n3646 9.3005
R9984 gnd.n3667 gnd.n3666 9.3005
R9985 gnd.n3663 gnd.n3647 9.3005
R9986 gnd.n3662 gnd.n3659 9.3005
R9987 gnd.n3658 gnd.n3648 9.3005
R9988 gnd.n3657 gnd.n3656 9.3005
R9989 gnd.n3653 gnd.n3649 9.3005
R9990 gnd.n3652 gnd.n3650 9.3005
R9991 gnd.n2159 gnd.n2158 9.3005
R9992 gnd.n3845 gnd.n3844 9.3005
R9993 gnd.n3688 gnd.n3642 9.3005
R9994 gnd.n3697 gnd.n3696 9.3005
R9995 gnd.n3857 gnd.n3856 9.3005
R9996 gnd.n3855 gnd.n2157 9.3005
R9997 gnd.n3854 gnd.n3853 9.3005
R9998 gnd.n3852 gnd.n3847 9.3005
R9999 gnd.n3850 gnd.n3849 9.3005
R10000 gnd.n3848 gnd.n846 9.3005
R10001 gnd.n6082 gnd.n847 9.3005
R10002 gnd.n6081 gnd.n848 9.3005
R10003 gnd.n6080 gnd.n849 9.3005
R10004 gnd.n867 gnd.n850 9.3005
R10005 gnd.n6070 gnd.n868 9.3005
R10006 gnd.n6069 gnd.n869 9.3005
R10007 gnd.n6068 gnd.n870 9.3005
R10008 gnd.n888 gnd.n871 9.3005
R10009 gnd.n6058 gnd.n889 9.3005
R10010 gnd.n6057 gnd.n890 9.3005
R10011 gnd.n6056 gnd.n891 9.3005
R10012 gnd.n3968 gnd.n892 9.3005
R10013 gnd.n3970 gnd.n3969 9.3005
R10014 gnd.n3971 gnd.n2088 9.3005
R10015 gnd.n3988 gnd.n2087 9.3005
R10016 gnd.n3996 gnd.n3989 9.3005
R10017 gnd.n3995 gnd.n3990 9.3005
R10018 gnd.n3994 gnd.n3992 9.3005
R10019 gnd.n3991 gnd.n915 9.3005
R10020 gnd.n6044 gnd.n916 9.3005
R10021 gnd.n6043 gnd.n917 9.3005
R10022 gnd.n6042 gnd.n918 9.3005
R10023 gnd.n934 gnd.n919 9.3005
R10024 gnd.n6032 gnd.n935 9.3005
R10025 gnd.n6031 gnd.n936 9.3005
R10026 gnd.n6030 gnd.n937 9.3005
R10027 gnd.n956 gnd.n938 9.3005
R10028 gnd.n6020 gnd.n957 9.3005
R10029 gnd.n6019 gnd.n958 9.3005
R10030 gnd.n6018 gnd.n959 9.3005
R10031 gnd.n977 gnd.n960 9.3005
R10032 gnd.n6008 gnd.n978 9.3005
R10033 gnd.n6007 gnd.n979 9.3005
R10034 gnd.n6006 gnd.n980 9.3005
R10035 gnd.n998 gnd.n981 9.3005
R10036 gnd.n5996 gnd.n5995 9.3005
R10037 gnd.n3846 gnd.n2156 9.3005
R10038 gnd.n1903 gnd.n1899 9.3005
R10039 gnd.n1936 gnd.n1933 9.3005
R10040 gnd.n1937 gnd.n1932 9.3005
R10041 gnd.n1940 gnd.n1931 9.3005
R10042 gnd.n1941 gnd.n1930 9.3005
R10043 gnd.n1944 gnd.n1929 9.3005
R10044 gnd.n1945 gnd.n1928 9.3005
R10045 gnd.n1948 gnd.n1927 9.3005
R10046 gnd.n1949 gnd.n1926 9.3005
R10047 gnd.n1952 gnd.n1925 9.3005
R10048 gnd.n1953 gnd.n1924 9.3005
R10049 gnd.n1956 gnd.n1923 9.3005
R10050 gnd.n1957 gnd.n1922 9.3005
R10051 gnd.n1958 gnd.n1921 9.3005
R10052 gnd.n1920 gnd.n1917 9.3005
R10053 gnd.n1919 gnd.n1918 9.3005
R10054 gnd.n4341 gnd.n4340 9.3005
R10055 gnd.n1905 gnd.n1904 9.3005
R10056 gnd.n1964 gnd.n1962 9.3005
R10057 gnd.n4333 gnd.n1965 9.3005
R10058 gnd.n4332 gnd.n1966 9.3005
R10059 gnd.n4331 gnd.n1967 9.3005
R10060 gnd.n1971 gnd.n1968 9.3005
R10061 gnd.n4326 gnd.n1972 9.3005
R10062 gnd.n4325 gnd.n1973 9.3005
R10063 gnd.n4324 gnd.n1974 9.3005
R10064 gnd.n1978 gnd.n1975 9.3005
R10065 gnd.n4319 gnd.n1979 9.3005
R10066 gnd.n4318 gnd.n1980 9.3005
R10067 gnd.n4317 gnd.n1981 9.3005
R10068 gnd.n1985 gnd.n1982 9.3005
R10069 gnd.n4312 gnd.n1986 9.3005
R10070 gnd.n4311 gnd.n1987 9.3005
R10071 gnd.n4310 gnd.n1988 9.3005
R10072 gnd.n1993 gnd.n1991 9.3005
R10073 gnd.n4305 gnd.n4304 9.3005
R10074 gnd.n4342 gnd.n1898 9.3005
R10075 gnd.n3760 gnd.n3759 9.3005
R10076 gnd.n3758 gnd.n3746 9.3005
R10077 gnd.n3757 gnd.n3756 9.3005
R10078 gnd.n3755 gnd.n3747 9.3005
R10079 gnd.n3753 gnd.n3748 9.3005
R10080 gnd.n3752 gnd.n3750 9.3005
R10081 gnd.n3749 gnd.n2136 9.3005
R10082 gnd.n3883 gnd.n2137 9.3005
R10083 gnd.n3884 gnd.n2135 9.3005
R10084 gnd.n3886 gnd.n3885 9.3005
R10085 gnd.n3887 gnd.n2134 9.3005
R10086 gnd.n3893 gnd.n3888 9.3005
R10087 gnd.n3892 gnd.n3889 9.3005
R10088 gnd.n3891 gnd.n3890 9.3005
R10089 gnd.n2119 gnd.n2118 9.3005
R10090 gnd.n3942 gnd.n3941 9.3005
R10091 gnd.n3943 gnd.n2117 9.3005
R10092 gnd.n3947 gnd.n3944 9.3005
R10093 gnd.n3946 gnd.n3945 9.3005
R10094 gnd.n2091 gnd.n2089 9.3005
R10095 gnd.n3987 gnd.n3986 9.3005
R10096 gnd.n2103 gnd.n2090 9.3005
R10097 gnd.n2102 gnd.n2092 9.3005
R10098 gnd.n2101 gnd.n2093 9.3005
R10099 gnd.n2099 gnd.n2094 9.3005
R10100 gnd.n2098 gnd.n2095 9.3005
R10101 gnd.n2097 gnd.n2096 9.3005
R10102 gnd.n2060 gnd.n2059 9.3005
R10103 gnd.n4036 gnd.n4035 9.3005
R10104 gnd.n4037 gnd.n2058 9.3005
R10105 gnd.n4039 gnd.n4038 9.3005
R10106 gnd.n4040 gnd.n2057 9.3005
R10107 gnd.n4044 gnd.n4043 9.3005
R10108 gnd.n4045 gnd.n2056 9.3005
R10109 gnd.n4050 gnd.n4046 9.3005
R10110 gnd.n4051 gnd.n2055 9.3005
R10111 gnd.n4055 gnd.n4054 9.3005
R10112 gnd.n4056 gnd.n2054 9.3005
R10113 gnd.n4059 gnd.n4058 9.3005
R10114 gnd.n4057 gnd.n1995 9.3005
R10115 gnd.n4301 gnd.n1994 9.3005
R10116 gnd.n4303 gnd.n4302 9.3005
R10117 gnd.n3761 gnd.n3744 9.3005
R10118 gnd.n3768 gnd.n3767 9.3005
R10119 gnd.n3769 gnd.n3738 9.3005
R10120 gnd.n3772 gnd.n3737 9.3005
R10121 gnd.n3773 gnd.n3736 9.3005
R10122 gnd.n3776 gnd.n3735 9.3005
R10123 gnd.n3777 gnd.n3734 9.3005
R10124 gnd.n3780 gnd.n3733 9.3005
R10125 gnd.n3781 gnd.n3732 9.3005
R10126 gnd.n3784 gnd.n3731 9.3005
R10127 gnd.n3785 gnd.n3730 9.3005
R10128 gnd.n3788 gnd.n3729 9.3005
R10129 gnd.n3789 gnd.n3728 9.3005
R10130 gnd.n3792 gnd.n3727 9.3005
R10131 gnd.n3793 gnd.n3726 9.3005
R10132 gnd.n3796 gnd.n3725 9.3005
R10133 gnd.n3797 gnd.n3724 9.3005
R10134 gnd.n3800 gnd.n3723 9.3005
R10135 gnd.n3801 gnd.n3722 9.3005
R10136 gnd.n3804 gnd.n3721 9.3005
R10137 gnd.n3806 gnd.n3718 9.3005
R10138 gnd.n3809 gnd.n3717 9.3005
R10139 gnd.n3810 gnd.n3716 9.3005
R10140 gnd.n3813 gnd.n3715 9.3005
R10141 gnd.n3814 gnd.n3714 9.3005
R10142 gnd.n3817 gnd.n3713 9.3005
R10143 gnd.n3818 gnd.n3712 9.3005
R10144 gnd.n3821 gnd.n3711 9.3005
R10145 gnd.n3822 gnd.n3710 9.3005
R10146 gnd.n3825 gnd.n3709 9.3005
R10147 gnd.n3826 gnd.n3708 9.3005
R10148 gnd.n3829 gnd.n3707 9.3005
R10149 gnd.n3830 gnd.n3706 9.3005
R10150 gnd.n3833 gnd.n3705 9.3005
R10151 gnd.n3835 gnd.n3704 9.3005
R10152 gnd.n3836 gnd.n3703 9.3005
R10153 gnd.n3837 gnd.n3702 9.3005
R10154 gnd.n3838 gnd.n3701 9.3005
R10155 gnd.n3766 gnd.n3743 9.3005
R10156 gnd.n3765 gnd.n3764 9.3005
R10157 gnd.n3862 gnd.n3861 9.3005
R10158 gnd.n3863 gnd.n2147 9.3005
R10159 gnd.n3866 gnd.n3865 9.3005
R10160 gnd.n3864 gnd.n834 9.3005
R10161 gnd.n6088 gnd.n835 9.3005
R10162 gnd.n6087 gnd.n836 9.3005
R10163 gnd.n6086 gnd.n837 9.3005
R10164 gnd.n856 gnd.n838 9.3005
R10165 gnd.n6076 gnd.n857 9.3005
R10166 gnd.n6075 gnd.n858 9.3005
R10167 gnd.n6074 gnd.n859 9.3005
R10168 gnd.n878 gnd.n860 9.3005
R10169 gnd.n6064 gnd.n879 9.3005
R10170 gnd.n6063 gnd.n880 9.3005
R10171 gnd.n6062 gnd.n881 9.3005
R10172 gnd.n906 gnd.n900 9.3005
R10173 gnd.n6038 gnd.n925 9.3005
R10174 gnd.n6037 gnd.n926 9.3005
R10175 gnd.n6036 gnd.n927 9.3005
R10176 gnd.n945 gnd.n928 9.3005
R10177 gnd.n6026 gnd.n946 9.3005
R10178 gnd.n6025 gnd.n947 9.3005
R10179 gnd.n6024 gnd.n948 9.3005
R10180 gnd.n966 gnd.n949 9.3005
R10181 gnd.n6014 gnd.n967 9.3005
R10182 gnd.n6013 gnd.n968 9.3005
R10183 gnd.n6012 gnd.n969 9.3005
R10184 gnd.n988 gnd.n970 9.3005
R10185 gnd.n6002 gnd.n989 9.3005
R10186 gnd.n6001 gnd.n990 9.3005
R10187 gnd.n6000 gnd.n991 9.3005
R10188 gnd.n2149 gnd.n2148 9.3005
R10189 gnd.n6049 gnd.n6048 9.3005
R10190 gnd.n3908 gnd.n3905 9.3005
R10191 gnd.n3912 gnd.n3911 9.3005
R10192 gnd.n3913 gnd.n3904 9.3005
R10193 gnd.n3915 gnd.n3914 9.3005
R10194 gnd.n2128 gnd.n2127 9.3005
R10195 gnd.n3920 gnd.n3919 9.3005
R10196 gnd.n3921 gnd.n2126 9.3005
R10197 gnd.n3926 gnd.n3922 9.3005
R10198 gnd.n3925 gnd.n3923 9.3005
R10199 gnd.n3907 gnd.n3906 9.3005
R10200 gnd.n6094 gnd.n824 9.3005
R10201 gnd.n6095 gnd.n823 9.3005
R10202 gnd.n822 gnd.n818 9.3005
R10203 gnd.n6101 gnd.n817 9.3005
R10204 gnd.n6102 gnd.n816 9.3005
R10205 gnd.n6103 gnd.n815 9.3005
R10206 gnd.n814 gnd.n810 9.3005
R10207 gnd.n6109 gnd.n809 9.3005
R10208 gnd.n6110 gnd.n808 9.3005
R10209 gnd.n6111 gnd.n807 9.3005
R10210 gnd.n806 gnd.n802 9.3005
R10211 gnd.n6117 gnd.n801 9.3005
R10212 gnd.n6118 gnd.n800 9.3005
R10213 gnd.n6119 gnd.n799 9.3005
R10214 gnd.n798 gnd.n794 9.3005
R10215 gnd.n6125 gnd.n793 9.3005
R10216 gnd.n6126 gnd.n792 9.3005
R10217 gnd.n6127 gnd.n791 9.3005
R10218 gnd.n790 gnd.n786 9.3005
R10219 gnd.n6133 gnd.n785 9.3005
R10220 gnd.n6134 gnd.n784 9.3005
R10221 gnd.n6135 gnd.n783 9.3005
R10222 gnd.n782 gnd.n778 9.3005
R10223 gnd.n6141 gnd.n777 9.3005
R10224 gnd.n6142 gnd.n776 9.3005
R10225 gnd.n6143 gnd.n775 9.3005
R10226 gnd.n774 gnd.n770 9.3005
R10227 gnd.n6149 gnd.n769 9.3005
R10228 gnd.n6150 gnd.n768 9.3005
R10229 gnd.n6151 gnd.n767 9.3005
R10230 gnd.n766 gnd.n762 9.3005
R10231 gnd.n6157 gnd.n761 9.3005
R10232 gnd.n6158 gnd.n760 9.3005
R10233 gnd.n6159 gnd.n759 9.3005
R10234 gnd.n758 gnd.n754 9.3005
R10235 gnd.n6165 gnd.n753 9.3005
R10236 gnd.n6166 gnd.n752 9.3005
R10237 gnd.n6167 gnd.n751 9.3005
R10238 gnd.n750 gnd.n746 9.3005
R10239 gnd.n6173 gnd.n745 9.3005
R10240 gnd.n6174 gnd.n744 9.3005
R10241 gnd.n6175 gnd.n743 9.3005
R10242 gnd.n742 gnd.n738 9.3005
R10243 gnd.n6181 gnd.n737 9.3005
R10244 gnd.n6182 gnd.n736 9.3005
R10245 gnd.n6183 gnd.n735 9.3005
R10246 gnd.n734 gnd.n730 9.3005
R10247 gnd.n6189 gnd.n729 9.3005
R10248 gnd.n6190 gnd.n728 9.3005
R10249 gnd.n6191 gnd.n727 9.3005
R10250 gnd.n726 gnd.n722 9.3005
R10251 gnd.n6197 gnd.n721 9.3005
R10252 gnd.n6198 gnd.n720 9.3005
R10253 gnd.n6199 gnd.n719 9.3005
R10254 gnd.n718 gnd.n714 9.3005
R10255 gnd.n6205 gnd.n713 9.3005
R10256 gnd.n6206 gnd.n712 9.3005
R10257 gnd.n6207 gnd.n711 9.3005
R10258 gnd.n710 gnd.n706 9.3005
R10259 gnd.n6213 gnd.n705 9.3005
R10260 gnd.n6214 gnd.n704 9.3005
R10261 gnd.n6215 gnd.n703 9.3005
R10262 gnd.n702 gnd.n698 9.3005
R10263 gnd.n6221 gnd.n697 9.3005
R10264 gnd.n6222 gnd.n696 9.3005
R10265 gnd.n6223 gnd.n695 9.3005
R10266 gnd.n694 gnd.n690 9.3005
R10267 gnd.n6229 gnd.n689 9.3005
R10268 gnd.n6230 gnd.n688 9.3005
R10269 gnd.n6231 gnd.n687 9.3005
R10270 gnd.n686 gnd.n682 9.3005
R10271 gnd.n6237 gnd.n681 9.3005
R10272 gnd.n6238 gnd.n680 9.3005
R10273 gnd.n6239 gnd.n679 9.3005
R10274 gnd.n678 gnd.n674 9.3005
R10275 gnd.n6245 gnd.n673 9.3005
R10276 gnd.n6246 gnd.n672 9.3005
R10277 gnd.n6247 gnd.n671 9.3005
R10278 gnd.n670 gnd.n666 9.3005
R10279 gnd.n6253 gnd.n665 9.3005
R10280 gnd.n6254 gnd.n664 9.3005
R10281 gnd.n6255 gnd.n663 9.3005
R10282 gnd.n659 gnd.n658 9.3005
R10283 gnd.n6262 gnd.n6261 9.3005
R10284 gnd.n6093 gnd.n825 9.3005
R10285 gnd.n5215 gnd.n5214 9.3005
R10286 gnd.n5195 gnd.n5193 9.3005
R10287 gnd.n5222 gnd.n5221 9.3005
R10288 gnd.n5189 gnd.n5188 9.3005
R10289 gnd.n5234 gnd.n5233 9.3005
R10290 gnd.n5186 gnd.n5184 9.3005
R10291 gnd.n5241 gnd.n5240 9.3005
R10292 gnd.n5180 gnd.n5179 9.3005
R10293 gnd.n5253 gnd.n5252 9.3005
R10294 gnd.n5177 gnd.n5175 9.3005
R10295 gnd.n5260 gnd.n5259 9.3005
R10296 gnd.n5171 gnd.n5170 9.3005
R10297 gnd.n5272 gnd.n5271 9.3005
R10298 gnd.n5168 gnd.n5166 9.3005
R10299 gnd.n5281 gnd.n5280 9.3005
R10300 gnd.n5279 gnd.n5160 9.3005
R10301 gnd.n5290 gnd.n5159 9.3005
R10302 gnd.n5293 gnd.n5292 9.3005
R10303 gnd.n5198 gnd.n5197 9.3005
R10304 gnd.n5283 gnd.n5282 9.3005
R10305 gnd.n5270 gnd.n5165 9.3005
R10306 gnd.n5269 gnd.n5268 9.3005
R10307 gnd.n5176 gnd.n5172 9.3005
R10308 gnd.n5262 gnd.n5261 9.3005
R10309 gnd.n5251 gnd.n5174 9.3005
R10310 gnd.n5250 gnd.n5249 9.3005
R10311 gnd.n5185 gnd.n5181 9.3005
R10312 gnd.n5243 gnd.n5242 9.3005
R10313 gnd.n5232 gnd.n5183 9.3005
R10314 gnd.n5231 gnd.n5230 9.3005
R10315 gnd.n5194 gnd.n5190 9.3005
R10316 gnd.n5224 gnd.n5223 9.3005
R10317 gnd.n5213 gnd.n5192 9.3005
R10318 gnd.n5212 gnd.n5211 9.3005
R10319 gnd.n5200 gnd.n5199 9.3005
R10320 gnd.n5167 gnd.n5163 9.3005
R10321 gnd.n5289 gnd.n5288 9.3005
R10322 gnd.n5157 gnd.n5156 9.3005
R10323 gnd.n5300 gnd.n5299 9.3005
R10324 gnd.n5301 gnd.n5155 9.3005
R10325 gnd.n5303 gnd.n5302 9.3005
R10326 gnd.n5153 gnd.n5152 9.3005
R10327 gnd.n5313 gnd.n5312 9.3005
R10328 gnd.n5314 gnd.n5151 9.3005
R10329 gnd.n5316 gnd.n5315 9.3005
R10330 gnd.n5149 gnd.n5148 9.3005
R10331 gnd.n5322 gnd.n5321 9.3005
R10332 gnd.n4274 gnd.n2018 9.3005
R10333 gnd.n4273 gnd.n4272 9.3005
R10334 gnd.n4271 gnd.n4258 9.3005
R10335 gnd.n4270 gnd.n4269 9.3005
R10336 gnd.n4268 gnd.n4259 9.3005
R10337 gnd.n4267 gnd.n4266 9.3005
R10338 gnd.n1743 gnd.n1742 9.3005
R10339 gnd.n4481 gnd.n4480 9.3005
R10340 gnd.n4482 gnd.n1740 9.3005
R10341 gnd.n4498 gnd.n4497 9.3005
R10342 gnd.n4496 gnd.n1741 9.3005
R10343 gnd.n4495 gnd.n4494 9.3005
R10344 gnd.n4493 gnd.n4483 9.3005
R10345 gnd.n4492 gnd.n4491 9.3005
R10346 gnd.n4490 gnd.n4487 9.3005
R10347 gnd.n4489 gnd.n4488 9.3005
R10348 gnd.n1696 gnd.n1695 9.3005
R10349 gnd.n4568 gnd.n4567 9.3005
R10350 gnd.n4569 gnd.n1693 9.3005
R10351 gnd.n4578 gnd.n4577 9.3005
R10352 gnd.n4576 gnd.n1694 9.3005
R10353 gnd.n4575 gnd.n4574 9.3005
R10354 gnd.n4573 gnd.n4570 9.3005
R10355 gnd.n1653 gnd.n1652 9.3005
R10356 gnd.n4654 gnd.n4653 9.3005
R10357 gnd.n4655 gnd.n1650 9.3005
R10358 gnd.n4693 gnd.n4692 9.3005
R10359 gnd.n4691 gnd.n1651 9.3005
R10360 gnd.n4690 gnd.n4689 9.3005
R10361 gnd.n4688 gnd.n4656 9.3005
R10362 gnd.n4687 gnd.n4686 9.3005
R10363 gnd.n4685 gnd.n4660 9.3005
R10364 gnd.n4684 gnd.n4683 9.3005
R10365 gnd.n4682 gnd.n4661 9.3005
R10366 gnd.n4681 gnd.n4680 9.3005
R10367 gnd.n4679 gnd.n4665 9.3005
R10368 gnd.n4678 gnd.n4677 9.3005
R10369 gnd.n4676 gnd.n4666 9.3005
R10370 gnd.n4675 gnd.n4674 9.3005
R10371 gnd.n4673 gnd.n4672 9.3005
R10372 gnd.n1565 gnd.n1564 9.3005
R10373 gnd.n4831 gnd.n4830 9.3005
R10374 gnd.n4832 gnd.n1562 9.3005
R10375 gnd.n4847 gnd.n4846 9.3005
R10376 gnd.n4845 gnd.n1563 9.3005
R10377 gnd.n4844 gnd.n4843 9.3005
R10378 gnd.n4842 gnd.n4833 9.3005
R10379 gnd.n4841 gnd.n4840 9.3005
R10380 gnd.n4839 gnd.n4838 9.3005
R10381 gnd.n1515 gnd.n1514 9.3005
R10382 gnd.n4916 gnd.n4915 9.3005
R10383 gnd.n4917 gnd.n1512 9.3005
R10384 gnd.n4923 gnd.n4922 9.3005
R10385 gnd.n4921 gnd.n1513 9.3005
R10386 gnd.n4920 gnd.n4919 9.3005
R10387 gnd.n1485 gnd.n1484 9.3005
R10388 gnd.n4983 gnd.n4982 9.3005
R10389 gnd.n4984 gnd.n1482 9.3005
R10390 gnd.n5000 gnd.n4999 9.3005
R10391 gnd.n4998 gnd.n1483 9.3005
R10392 gnd.n4997 gnd.n4996 9.3005
R10393 gnd.n4995 gnd.n4985 9.3005
R10394 gnd.n4994 gnd.n4993 9.3005
R10395 gnd.n4992 gnd.n4991 9.3005
R10396 gnd.n1410 gnd.n1409 9.3005
R10397 gnd.n5068 gnd.n5067 9.3005
R10398 gnd.n5069 gnd.n1407 9.3005
R10399 gnd.n5072 gnd.n5071 9.3005
R10400 gnd.n5070 gnd.n1408 9.3005
R10401 gnd.n1381 gnd.n1380 9.3005
R10402 gnd.n5104 gnd.n5103 9.3005
R10403 gnd.n5105 gnd.n1379 9.3005
R10404 gnd.n5107 gnd.n5106 9.3005
R10405 gnd.n1359 gnd.n1358 9.3005
R10406 gnd.n5135 gnd.n5134 9.3005
R10407 gnd.n5136 gnd.n1357 9.3005
R10408 gnd.n5138 gnd.n5137 9.3005
R10409 gnd.n1355 gnd.n1354 9.3005
R10410 gnd.n5146 gnd.n5145 9.3005
R10411 gnd.n5147 gnd.n1352 9.3005
R10412 gnd.n5325 gnd.n5324 9.3005
R10413 gnd.n5323 gnd.n1353 9.3005
R10414 gnd.n4276 gnd.n4275 9.3005
R10415 gnd.n4279 gnd.n4278 9.3005
R10416 gnd.n4280 gnd.n2013 9.3005
R10417 gnd.n4282 gnd.n4281 9.3005
R10418 gnd.n4284 gnd.n4283 9.3005
R10419 gnd.n4285 gnd.n2006 9.3005
R10420 gnd.n4287 gnd.n4286 9.3005
R10421 gnd.n4288 gnd.n2005 9.3005
R10422 gnd.n4290 gnd.n4289 9.3005
R10423 gnd.n4291 gnd.n1999 9.3005
R10424 gnd.n4277 gnd.n2017 9.3005
R10425 gnd.n2075 gnd.n2074 9.3005
R10426 gnd.n4007 gnd.n4006 9.3005
R10427 gnd.n4008 gnd.n2073 9.3005
R10428 gnd.n4010 gnd.n4009 9.3005
R10429 gnd.n2063 gnd.n2062 9.3005
R10430 gnd.n4028 gnd.n4027 9.3005
R10431 gnd.n4029 gnd.n2061 9.3005
R10432 gnd.n4031 gnd.n4030 9.3005
R10433 gnd.n2047 gnd.n2045 9.3005
R10434 gnd.n4076 gnd.n4075 9.3005
R10435 gnd.n4074 gnd.n2046 9.3005
R10436 gnd.n4073 gnd.n4072 9.3005
R10437 gnd.n4071 gnd.n2048 9.3005
R10438 gnd.n4070 gnd.n4069 9.3005
R10439 gnd.n4068 gnd.n2051 9.3005
R10440 gnd.n4067 gnd.n4066 9.3005
R10441 gnd.n4065 gnd.n2052 9.3005
R10442 gnd.n4064 gnd.n4063 9.3005
R10443 gnd.n1998 gnd.n1996 9.3005
R10444 gnd.n4297 gnd.n4296 9.3005
R10445 gnd.n4295 gnd.n1997 9.3005
R10446 gnd.n4293 gnd.n4292 9.3005
R10447 gnd.n2001 gnd.n2000 9.3005
R10448 gnd.n4200 gnd.n4199 9.3005
R10449 gnd.n4202 gnd.n4201 9.3005
R10450 gnd.n4180 gnd.n4179 9.3005
R10451 gnd.n4208 gnd.n4207 9.3005
R10452 gnd.n4210 gnd.n4209 9.3005
R10453 gnd.n4170 gnd.n4169 9.3005
R10454 gnd.n4216 gnd.n4215 9.3005
R10455 gnd.n4218 gnd.n4217 9.3005
R10456 gnd.n4157 gnd.n4156 9.3005
R10457 gnd.n4224 gnd.n4223 9.3005
R10458 gnd.n4226 gnd.n4225 9.3005
R10459 gnd.n4147 gnd.n4146 9.3005
R10460 gnd.n4232 gnd.n4231 9.3005
R10461 gnd.n4234 gnd.n4233 9.3005
R10462 gnd.n4132 gnd.n4130 9.3005
R10463 gnd.n4240 gnd.n4239 9.3005
R10464 gnd.n4241 gnd.n4129 9.3005
R10465 gnd.n4134 gnd.n1000 9.3005
R10466 gnd.n4133 gnd.n4131 9.3005
R10467 gnd.n4238 gnd.n4237 9.3005
R10468 gnd.n4236 gnd.n4235 9.3005
R10469 gnd.n4142 gnd.n4141 9.3005
R10470 gnd.n4230 gnd.n4229 9.3005
R10471 gnd.n4228 gnd.n4227 9.3005
R10472 gnd.n4153 gnd.n4152 9.3005
R10473 gnd.n4222 gnd.n4221 9.3005
R10474 gnd.n4220 gnd.n4219 9.3005
R10475 gnd.n4164 gnd.n4163 9.3005
R10476 gnd.n4214 gnd.n4213 9.3005
R10477 gnd.n4212 gnd.n4211 9.3005
R10478 gnd.n4176 gnd.n4175 9.3005
R10479 gnd.n4206 gnd.n4205 9.3005
R10480 gnd.n4204 gnd.n4203 9.3005
R10481 gnd.n4189 gnd.n4188 9.3005
R10482 gnd.n4198 gnd.n4197 9.3005
R10483 gnd.n5990 gnd.n1001 9.3005
R10484 gnd.n5989 gnd.n5988 9.3005
R10485 gnd.n5987 gnd.n1005 9.3005
R10486 gnd.n5986 gnd.n5985 9.3005
R10487 gnd.n5984 gnd.n1006 9.3005
R10488 gnd.n5983 gnd.n5982 9.3005
R10489 gnd.n5981 gnd.n1010 9.3005
R10490 gnd.n5980 gnd.n5979 9.3005
R10491 gnd.n5978 gnd.n1011 9.3005
R10492 gnd.n5977 gnd.n5976 9.3005
R10493 gnd.n5975 gnd.n1015 9.3005
R10494 gnd.n5974 gnd.n5973 9.3005
R10495 gnd.n5972 gnd.n1016 9.3005
R10496 gnd.n5971 gnd.n5970 9.3005
R10497 gnd.n5969 gnd.n1020 9.3005
R10498 gnd.n5968 gnd.n5967 9.3005
R10499 gnd.n5966 gnd.n1021 9.3005
R10500 gnd.n5965 gnd.n5964 9.3005
R10501 gnd.n5963 gnd.n1025 9.3005
R10502 gnd.n5962 gnd.n5961 9.3005
R10503 gnd.n5960 gnd.n1026 9.3005
R10504 gnd.n5959 gnd.n5958 9.3005
R10505 gnd.n5957 gnd.n1030 9.3005
R10506 gnd.n5956 gnd.n5955 9.3005
R10507 gnd.n5954 gnd.n1031 9.3005
R10508 gnd.n5953 gnd.n5952 9.3005
R10509 gnd.n5951 gnd.n1035 9.3005
R10510 gnd.n5950 gnd.n5949 9.3005
R10511 gnd.n5948 gnd.n1036 9.3005
R10512 gnd.n5947 gnd.n5946 9.3005
R10513 gnd.n5945 gnd.n1040 9.3005
R10514 gnd.n5944 gnd.n5943 9.3005
R10515 gnd.n5942 gnd.n1041 9.3005
R10516 gnd.n5941 gnd.n5940 9.3005
R10517 gnd.n5939 gnd.n1045 9.3005
R10518 gnd.n5938 gnd.n5937 9.3005
R10519 gnd.n5936 gnd.n1046 9.3005
R10520 gnd.n5935 gnd.n5934 9.3005
R10521 gnd.n5933 gnd.n1050 9.3005
R10522 gnd.n5932 gnd.n5931 9.3005
R10523 gnd.n5930 gnd.n1051 9.3005
R10524 gnd.n5929 gnd.n5928 9.3005
R10525 gnd.n5927 gnd.n1055 9.3005
R10526 gnd.n5926 gnd.n5925 9.3005
R10527 gnd.n5924 gnd.n1056 9.3005
R10528 gnd.n5923 gnd.n5922 9.3005
R10529 gnd.n5921 gnd.n1060 9.3005
R10530 gnd.n5920 gnd.n5919 9.3005
R10531 gnd.n5918 gnd.n1061 9.3005
R10532 gnd.n5917 gnd.n5916 9.3005
R10533 gnd.n5915 gnd.n1065 9.3005
R10534 gnd.n5914 gnd.n5913 9.3005
R10535 gnd.n5912 gnd.n1066 9.3005
R10536 gnd.n5911 gnd.n5910 9.3005
R10537 gnd.n5909 gnd.n1070 9.3005
R10538 gnd.n5908 gnd.n5907 9.3005
R10539 gnd.n5906 gnd.n1071 9.3005
R10540 gnd.n5905 gnd.n5904 9.3005
R10541 gnd.n5903 gnd.n1075 9.3005
R10542 gnd.n5902 gnd.n5901 9.3005
R10543 gnd.n5900 gnd.n1076 9.3005
R10544 gnd.n5899 gnd.n5898 9.3005
R10545 gnd.n5897 gnd.n1080 9.3005
R10546 gnd.n5896 gnd.n5895 9.3005
R10547 gnd.n5894 gnd.n1081 9.3005
R10548 gnd.n5893 gnd.n5892 9.3005
R10549 gnd.n5891 gnd.n1085 9.3005
R10550 gnd.n5890 gnd.n5889 9.3005
R10551 gnd.n5888 gnd.n1086 9.3005
R10552 gnd.n5887 gnd.n5886 9.3005
R10553 gnd.n5885 gnd.n1090 9.3005
R10554 gnd.n5884 gnd.n5883 9.3005
R10555 gnd.n5882 gnd.n1091 9.3005
R10556 gnd.n5881 gnd.n5880 9.3005
R10557 gnd.n5879 gnd.n1095 9.3005
R10558 gnd.n5878 gnd.n5877 9.3005
R10559 gnd.n5876 gnd.n1096 9.3005
R10560 gnd.n5875 gnd.n5874 9.3005
R10561 gnd.n5873 gnd.n1100 9.3005
R10562 gnd.n5872 gnd.n5871 9.3005
R10563 gnd.n5870 gnd.n1101 9.3005
R10564 gnd.n5869 gnd.n1104 9.3005
R10565 gnd.n5992 gnd.n5991 9.3005
R10566 gnd.n1146 gnd.n1144 9.3005
R10567 gnd.n5843 gnd.n5842 9.3005
R10568 gnd.n5841 gnd.n1145 9.3005
R10569 gnd.n5840 gnd.n5839 9.3005
R10570 gnd.n5838 gnd.n1147 9.3005
R10571 gnd.n5837 gnd.n5836 9.3005
R10572 gnd.n5835 gnd.n1151 9.3005
R10573 gnd.n5834 gnd.n5833 9.3005
R10574 gnd.n5832 gnd.n1152 9.3005
R10575 gnd.n5831 gnd.n5830 9.3005
R10576 gnd.n5829 gnd.n1156 9.3005
R10577 gnd.n5828 gnd.n5827 9.3005
R10578 gnd.n5826 gnd.n1157 9.3005
R10579 gnd.n5825 gnd.n5824 9.3005
R10580 gnd.n5823 gnd.n1161 9.3005
R10581 gnd.n5822 gnd.n5821 9.3005
R10582 gnd.n5820 gnd.n1162 9.3005
R10583 gnd.n5819 gnd.n5818 9.3005
R10584 gnd.n5817 gnd.n1166 9.3005
R10585 gnd.n5816 gnd.n5815 9.3005
R10586 gnd.n5814 gnd.n1167 9.3005
R10587 gnd.n5813 gnd.n5812 9.3005
R10588 gnd.n229 gnd.n228 9.3005
R10589 gnd.n6935 gnd.n6934 9.3005
R10590 gnd.n6936 gnd.n227 9.3005
R10591 gnd.n6938 gnd.n6937 9.3005
R10592 gnd.n207 gnd.n206 9.3005
R10593 gnd.n6951 gnd.n6950 9.3005
R10594 gnd.n6952 gnd.n205 9.3005
R10595 gnd.n6954 gnd.n6953 9.3005
R10596 gnd.n192 gnd.n191 9.3005
R10597 gnd.n6967 gnd.n6966 9.3005
R10598 gnd.n6968 gnd.n190 9.3005
R10599 gnd.n6970 gnd.n6969 9.3005
R10600 gnd.n175 gnd.n174 9.3005
R10601 gnd.n6983 gnd.n6982 9.3005
R10602 gnd.n6984 gnd.n172 9.3005
R10603 gnd.n7060 gnd.n7059 9.3005
R10604 gnd.n7058 gnd.n173 9.3005
R10605 gnd.n7057 gnd.n7056 9.3005
R10606 gnd.n7055 gnd.n6985 9.3005
R10607 gnd.n7054 gnd.n7053 9.3005
R10608 gnd.n5203 gnd.n5202 9.3005
R10609 gnd.n7050 gnd.n6987 9.3005
R10610 gnd.n7049 gnd.n7048 9.3005
R10611 gnd.n7047 gnd.n6992 9.3005
R10612 gnd.n7046 gnd.n7045 9.3005
R10613 gnd.n7044 gnd.n6993 9.3005
R10614 gnd.n7043 gnd.n7042 9.3005
R10615 gnd.n7041 gnd.n7000 9.3005
R10616 gnd.n7040 gnd.n7039 9.3005
R10617 gnd.n7038 gnd.n7001 9.3005
R10618 gnd.n7037 gnd.n7036 9.3005
R10619 gnd.n7035 gnd.n7008 9.3005
R10620 gnd.n7034 gnd.n7033 9.3005
R10621 gnd.n7032 gnd.n7009 9.3005
R10622 gnd.n7031 gnd.n7030 9.3005
R10623 gnd.n7029 gnd.n7016 9.3005
R10624 gnd.n7028 gnd.n7027 9.3005
R10625 gnd.n7026 gnd.n7017 9.3005
R10626 gnd.n7025 gnd.n78 9.3005
R10627 gnd.n7052 gnd.n7051 9.3005
R10628 gnd.n5615 gnd.n5614 9.3005
R10629 gnd.n5616 gnd.n1262 9.3005
R10630 gnd.n5619 gnd.n5618 9.3005
R10631 gnd.n5617 gnd.n1263 9.3005
R10632 gnd.n1247 gnd.n1246 9.3005
R10633 gnd.n5701 gnd.n5700 9.3005
R10634 gnd.n5702 gnd.n1244 9.3005
R10635 gnd.n5705 gnd.n5704 9.3005
R10636 gnd.n5703 gnd.n1245 9.3005
R10637 gnd.n1218 gnd.n1217 9.3005
R10638 gnd.n5733 gnd.n5732 9.3005
R10639 gnd.n5734 gnd.n1215 9.3005
R10640 gnd.n5737 gnd.n5736 9.3005
R10641 gnd.n5735 gnd.n1216 9.3005
R10642 gnd.n1192 gnd.n1191 9.3005
R10643 gnd.n5766 gnd.n5765 9.3005
R10644 gnd.n5767 gnd.n1188 9.3005
R10645 gnd.n5770 gnd.n5769 9.3005
R10646 gnd.n5768 gnd.n1190 9.3005
R10647 gnd.n1189 gnd.n51 9.3005
R10648 gnd.n7184 gnd.n52 9.3005
R10649 gnd.n7183 gnd.n7182 9.3005
R10650 gnd.n7181 gnd.n53 9.3005
R10651 gnd.n7180 gnd.n7179 9.3005
R10652 gnd.n7178 gnd.n57 9.3005
R10653 gnd.n7177 gnd.n7176 9.3005
R10654 gnd.n7175 gnd.n58 9.3005
R10655 gnd.n7174 gnd.n7173 9.3005
R10656 gnd.n7172 gnd.n62 9.3005
R10657 gnd.n7171 gnd.n7170 9.3005
R10658 gnd.n7169 gnd.n63 9.3005
R10659 gnd.n7168 gnd.n7167 9.3005
R10660 gnd.n7166 gnd.n67 9.3005
R10661 gnd.n7165 gnd.n7164 9.3005
R10662 gnd.n7163 gnd.n68 9.3005
R10663 gnd.n7162 gnd.n7161 9.3005
R10664 gnd.n7160 gnd.n72 9.3005
R10665 gnd.n7159 gnd.n7158 9.3005
R10666 gnd.n7157 gnd.n73 9.3005
R10667 gnd.n7156 gnd.n7155 9.3005
R10668 gnd.n7154 gnd.n77 9.3005
R10669 gnd.n7153 gnd.n7152 9.3005
R10670 gnd.n1265 gnd.n1264 9.3005
R10671 gnd.t195 gnd.n2351 9.24152
R10672 gnd.n2253 gnd.t56 9.24152
R10673 gnd.n3510 gnd.t60 9.24152
R10674 gnd.n4047 gnd.t249 9.24152
R10675 gnd.n4596 gnd.t168 9.24152
R10676 gnd.n5022 gnd.t133 9.24152
R10677 gnd.t11 gnd.n1251 9.24152
R10678 gnd.t276 gnd.t195 8.92286
R10679 gnd.n4452 gnd.n1764 8.92286
R10680 gnd.n4626 gnd.n1675 8.92286
R10681 gnd.n4697 gnd.n4696 8.92286
R10682 gnd.n4803 gnd.n1588 8.92286
R10683 gnd.n4850 gnd.n4849 8.92286
R10684 gnd.n4946 gnd.n1503 8.92286
R10685 gnd.n4931 gnd.n1465 8.92286
R10686 gnd.n1385 gnd.n1376 8.92286
R10687 gnd.n5140 gnd.n1340 8.92286
R10688 gnd.n3480 gnd.n3455 8.92171
R10689 gnd.n3448 gnd.n3423 8.92171
R10690 gnd.n3416 gnd.n3391 8.92171
R10691 gnd.n3385 gnd.n3360 8.92171
R10692 gnd.n3353 gnd.n3328 8.92171
R10693 gnd.n3321 gnd.n3296 8.92171
R10694 gnd.n3289 gnd.n3264 8.92171
R10695 gnd.n3258 gnd.n3233 8.92171
R10696 gnd.n5358 gnd.n5340 8.72777
R10697 gnd.n2983 gnd.t190 8.60421
R10698 gnd.n4413 gnd.n4412 8.60421
R10699 gnd.t130 gnd.n4801 8.60421
R10700 gnd.n4788 gnd.t288 8.60421
R10701 gnd.n2415 gnd.n2403 8.43467
R10702 gnd.n38 gnd.n26 8.43467
R10703 gnd.n3981 gnd.n0 8.41456
R10704 gnd.n7185 gnd.n7184 8.41456
R10705 gnd.n4261 gnd.t97 8.28555
R10706 gnd.n4530 gnd.n1690 8.28555
R10707 gnd.n4602 gnd.n1643 8.28555
R10708 gnd.n4757 gnd.n4756 8.28555
R10709 gnd.n4779 gnd.n1555 8.28555
R10710 gnd.n4954 gnd.n4953 8.28555
R10711 gnd.n5030 gnd.n1459 8.28555
R10712 gnd.t103 gnd.n1367 8.28555
R10713 gnd.n3481 gnd.n3453 8.14595
R10714 gnd.n3449 gnd.n3421 8.14595
R10715 gnd.n3417 gnd.n3389 8.14595
R10716 gnd.n3386 gnd.n3358 8.14595
R10717 gnd.n3354 gnd.n3326 8.14595
R10718 gnd.n3322 gnd.n3294 8.14595
R10719 gnd.n3290 gnd.n3262 8.14595
R10720 gnd.n3259 gnd.n3231 8.14595
R10721 gnd.n3486 gnd.n3485 7.97301
R10722 gnd.t143 gnd.n2498 7.9669
R10723 gnd.n4557 gnd.t191 7.9669
R10724 gnd.n5064 gnd.t223 7.9669
R10725 gnd.n7026 gnd.n7025 7.75808
R10726 gnd.n5288 gnd.n5163 7.75808
R10727 gnd.n4197 gnd.n4188 7.75808
R10728 gnd.n3697 gnd.n3642 7.75808
R10729 gnd.n4422 gnd.t97 7.64824
R10730 gnd.n4478 gnd.t116 7.64824
R10731 gnd.n4428 gnd.n1721 7.64824
R10732 gnd.n4530 gnd.t174 7.64824
R10733 gnd.t179 gnd.n1613 7.64824
R10734 gnd.n4662 gnd.t179 7.64824
R10735 gnd.n4836 gnd.t151 7.64824
R10736 gnd.t151 gnd.n1532 7.64824
R10737 gnd.n5030 gnd.t178 7.64824
R10738 gnd.n5091 gnd.n1390 7.64824
R10739 gnd.n5109 gnd.t103 7.64824
R10740 gnd.n2892 gnd.t206 7.32958
R10741 gnd.n4412 gnd.n1807 7.32958
R10742 gnd.n5493 gnd.n1296 7.32958
R10743 gnd.n1828 gnd.n1827 7.30353
R10744 gnd.n5357 gnd.n5356 7.30353
R10745 gnd.n2852 gnd.n2571 7.01093
R10746 gnd.n2574 gnd.n2572 7.01093
R10747 gnd.n2862 gnd.n2861 7.01093
R10748 gnd.n2873 gnd.n2555 7.01093
R10749 gnd.n2872 gnd.n2558 7.01093
R10750 gnd.n2883 gnd.n2546 7.01093
R10751 gnd.n2549 gnd.n2547 7.01093
R10752 gnd.n2893 gnd.n2892 7.01093
R10753 gnd.n2903 gnd.n2527 7.01093
R10754 gnd.n2902 gnd.n2530 7.01093
R10755 gnd.n2911 gnd.n2521 7.01093
R10756 gnd.n2923 gnd.n2511 7.01093
R10757 gnd.n2933 gnd.n2496 7.01093
R10758 gnd.n2949 gnd.n2948 7.01093
R10759 gnd.n2498 gnd.n2435 7.01093
R10760 gnd.n3003 gnd.n2436 7.01093
R10761 gnd.n2997 gnd.n2996 7.01093
R10762 gnd.n2485 gnd.n2447 7.01093
R10763 gnd.n2989 gnd.n2458 7.01093
R10764 gnd.n2476 gnd.n2471 7.01093
R10765 gnd.n2983 gnd.n2982 7.01093
R10766 gnd.n3029 gnd.n2386 7.01093
R10767 gnd.n3028 gnd.n3027 7.01093
R10768 gnd.n3040 gnd.n3039 7.01093
R10769 gnd.n2379 gnd.n2371 7.01093
R10770 gnd.n3069 gnd.n2359 7.01093
R10771 gnd.n3068 gnd.n2362 7.01093
R10772 gnd.n3079 gnd.n2351 7.01093
R10773 gnd.n2352 gnd.n2340 7.01093
R10774 gnd.n3090 gnd.n2341 7.01093
R10775 gnd.n3114 gnd.n2332 7.01093
R10776 gnd.n3113 gnd.n2323 7.01093
R10777 gnd.n3137 gnd.n3136 7.01093
R10778 gnd.n3155 gnd.n2304 7.01093
R10779 gnd.n3154 gnd.n2307 7.01093
R10780 gnd.n3165 gnd.n2296 7.01093
R10781 gnd.n2297 gnd.n2284 7.01093
R10782 gnd.n3176 gnd.n2285 7.01093
R10783 gnd.n3203 gnd.n2269 7.01093
R10784 gnd.n3215 gnd.n3214 7.01093
R10785 gnd.n3197 gnd.n2262 7.01093
R10786 gnd.n3226 gnd.n3225 7.01093
R10787 gnd.n3498 gnd.n2250 7.01093
R10788 gnd.n3497 gnd.n2253 7.01093
R10789 gnd.n3510 gnd.n2242 7.01093
R10790 gnd.n2243 gnd.n2235 7.01093
R10791 gnd.n3520 gnd.n2161 7.01093
R10792 gnd.n4452 gnd.n4451 7.01093
R10793 gnd.n4501 gnd.n1737 7.01093
R10794 gnd.n4697 gnd.n1647 7.01093
R10795 gnd.t10 gnd.n1601 7.01093
R10796 gnd.n4803 gnd.n4802 7.01093
R10797 gnd.n4850 gnd.n1559 7.01093
R10798 gnd.t239 gnd.n1542 7.01093
R10799 gnd.n4946 gnd.n4945 7.01093
R10800 gnd.n5111 gnd.n1376 7.01093
R10801 gnd.n5335 gnd.n1340 7.01093
R10802 gnd.n5140 gnd.t74 7.01093
R10803 gnd.n2530 gnd.t171 6.69227
R10804 gnd.n2362 gnd.t276 6.69227
R10805 gnd.n3204 gnd.t161 6.69227
R10806 gnd.n4580 gnd.t168 6.69227
R10807 gnd.n4988 gnd.t133 6.69227
R10808 gnd.n5487 gnd.n5486 6.5566
R10809 gnd.n1893 gnd.n1892 6.5566
R10810 gnd.n4353 gnd.n1833 6.5566
R10811 gnd.n5365 gnd.n5364 6.5566
R10812 gnd.n3135 gnd.n2304 6.37362
R10813 gnd.n4526 gnd.n1716 6.37362
R10814 gnd.n4564 gnd.n4563 6.37362
R10815 gnd.n4721 gnd.n1626 6.37362
R10816 gnd.n4913 gnd.n4911 6.37362
R10817 gnd.n5058 gnd.n5057 6.37362
R10818 gnd.n5074 gnd.n1397 6.37362
R10819 gnd.n4281 gnd.n2012 6.20656
R10820 gnd.n7115 gnd.n7112 6.20656
R10821 gnd.n3805 gnd.n3804 6.20656
R10822 gnd.n5311 gnd.n5151 6.20656
R10823 gnd.t184 gnd.n2959 6.05496
R10824 gnd.n2960 gnd.t127 6.05496
R10825 gnd.t144 gnd.n2386 6.05496
R10826 gnd.t128 gnd.n3124 6.05496
R10827 gnd.n3483 gnd.n3453 5.81868
R10828 gnd.n3451 gnd.n3421 5.81868
R10829 gnd.n3419 gnd.n3389 5.81868
R10830 gnd.n3388 gnd.n3358 5.81868
R10831 gnd.n3356 gnd.n3326 5.81868
R10832 gnd.n3324 gnd.n3294 5.81868
R10833 gnd.n3292 gnd.n3262 5.81868
R10834 gnd.n3261 gnd.n3231 5.81868
R10835 gnd.n4469 gnd.n1745 5.73631
R10836 gnd.n4501 gnd.t32 5.73631
R10837 gnd.n4626 gnd.t159 5.73631
R10838 gnd.n4618 gnd.n4617 5.73631
R10839 gnd.n4643 gnd.n1661 5.73631
R10840 gnd.t197 gnd.n1619 5.73631
R10841 gnd.n4802 gnd.t208 5.73631
R10842 gnd.n4795 gnd.n1573 5.73631
R10843 gnd.n4820 gnd.n1567 5.73631
R10844 gnd.t280 gnd.n1559 5.73631
R10845 gnd.n1525 gnd.t238 5.73631
R10846 gnd.n4979 gnd.n1489 5.73631
R10847 gnd.n5004 gnd.n1479 5.73631
R10848 gnd.n4931 gnd.t0 5.73631
R10849 gnd.n5123 gnd.n5122 5.73631
R10850 gnd.n5426 gnd.t74 5.73631
R10851 gnd.n5496 gnd.n1292 5.62001
R10852 gnd.n4348 gnd.n1897 5.62001
R10853 gnd.n4349 gnd.n4348 5.62001
R10854 gnd.n5496 gnd.n1293 5.62001
R10855 gnd.n2711 gnd.n2706 5.4308
R10856 gnd.n3528 gnd.n2228 5.4308
R10857 gnd.n3027 gnd.t142 5.41765
R10858 gnd.t194 gnd.n3050 5.41765
R10859 gnd.t175 gnd.n2316 5.41765
R10860 gnd.n4651 gnd.t217 5.41765
R10861 gnd.n4980 gnd.t135 5.41765
R10862 gnd.n4546 gnd.n4544 5.09899
R10863 gnd.n4557 gnd.n4556 5.09899
R10864 gnd.t180 gnd.n1631 5.09899
R10865 gnd.n4731 gnd.n4730 5.09899
R10866 gnd.n4742 gnd.n4741 5.09899
R10867 gnd.n4885 gnd.n4884 5.09899
R10868 gnd.n4904 gnd.n4903 5.09899
R10869 gnd.n4925 gnd.t183 5.09899
R10870 gnd.n5065 gnd.n5064 5.09899
R10871 gnd.n5050 gnd.n5049 5.09899
R10872 gnd.n3481 gnd.n3480 5.04292
R10873 gnd.n3449 gnd.n3448 5.04292
R10874 gnd.n3417 gnd.n3416 5.04292
R10875 gnd.n3386 gnd.n3385 5.04292
R10876 gnd.n3354 gnd.n3353 5.04292
R10877 gnd.n3322 gnd.n3321 5.04292
R10878 gnd.n3290 gnd.n3289 5.04292
R10879 gnd.n3259 gnd.n3258 5.04292
R10880 gnd.n2427 gnd.n2426 4.82753
R10881 gnd.n50 gnd.n49 4.82753
R10882 gnd.n2990 gnd.t188 4.78034
R10883 gnd.n2341 gnd.t163 4.78034
R10884 gnd.t166 gnd.n4443 4.78034
R10885 gnd.n1661 gnd.t217 4.78034
R10886 gnd.t135 gnd.n4979 4.78034
R10887 gnd.t202 gnd.n1424 4.78034
R10888 gnd.n5493 gnd.t39 4.78034
R10889 gnd.n2432 gnd.n2429 4.74817
R10890 gnd.n2482 gnd.n2392 4.74817
R10891 gnd.n2469 gnd.n2391 4.74817
R10892 gnd.n2390 gnd.n2389 4.74817
R10893 gnd.n2478 gnd.n2429 4.74817
R10894 gnd.n2479 gnd.n2392 4.74817
R10895 gnd.n2481 gnd.n2391 4.74817
R10896 gnd.n2468 gnd.n2390 4.74817
R10897 gnd.n1182 gnd.n220 4.74817
R10898 gnd.n5779 gnd.n219 4.74817
R10899 gnd.n5777 gnd.n218 4.74817
R10900 gnd.n6929 gnd.n217 4.74817
R10901 gnd.n221 gnd.n216 4.74817
R10902 gnd.n5761 gnd.n220 4.74817
R10903 gnd.n1183 gnd.n219 4.74817
R10904 gnd.n5780 gnd.n218 4.74817
R10905 gnd.n5776 gnd.n217 4.74817
R10906 gnd.n6930 gnd.n216 4.74817
R10907 gnd.n3924 gnd.n2115 4.74817
R10908 gnd.n3963 gnd.n3954 4.74817
R10909 gnd.n3961 gnd.n3960 4.74817
R10910 gnd.n3956 gnd.n3955 4.74817
R10911 gnd.n4016 gnd.n2067 4.74817
R10912 gnd.n5749 gnd.n5747 4.74817
R10913 gnd.n5785 gnd.n1173 4.74817
R10914 gnd.n5807 gnd.n5787 4.74817
R10915 gnd.n5805 gnd.n5804 4.74817
R10916 gnd.n5800 gnd.n5790 4.74817
R10917 gnd.n5752 gnd.n5747 4.74817
R10918 gnd.n5748 gnd.n1173 4.74817
R10919 gnd.n5787 gnd.n5786 4.74817
R10920 gnd.n5806 gnd.n5805 4.74817
R10921 gnd.n5790 gnd.n5788 4.74817
R10922 gnd.n6052 gnd.n898 4.74817
R10923 gnd.n6050 gnd.n899 4.74817
R10924 gnd.n2082 gnd.n904 4.74817
R10925 gnd.n4002 gnd.n903 4.74817
R10926 gnd.n905 gnd.n902 4.74817
R10927 gnd.n898 gnd.n882 4.74817
R10928 gnd.n6051 gnd.n6050 4.74817
R10929 gnd.n3967 gnd.n904 4.74817
R10930 gnd.n2083 gnd.n903 4.74817
R10931 gnd.n4001 gnd.n902 4.74817
R10932 gnd.n3952 gnd.n2115 4.74817
R10933 gnd.n3954 gnd.n3953 4.74817
R10934 gnd.n3962 gnd.n3961 4.74817
R10935 gnd.n3957 gnd.n3956 4.74817
R10936 gnd.n2069 gnd.n2067 4.74817
R10937 gnd.n2415 gnd.n2414 4.7074
R10938 gnd.n38 gnd.n37 4.7074
R10939 gnd.n2427 gnd.n2415 4.65959
R10940 gnd.n50 gnd.n38 4.65959
R10941 gnd.n5555 gnd.n5554 4.6132
R10942 gnd.n4344 gnd.n4343 4.6132
R10943 gnd.n4459 gnd.n4458 4.46168
R10944 gnd.n4477 gnd.n1747 4.46168
R10945 gnd.n4428 gnd.t222 4.46168
R10946 gnd.n4633 gnd.n4632 4.46168
R10947 gnd.n4650 gnd.n1656 4.46168
R10948 gnd.n4810 gnd.n4809 4.46168
R10949 gnd.n4827 gnd.n1569 4.46168
R10950 gnd.n4971 gnd.n1487 4.46168
R10951 gnd.n5012 gnd.n1472 4.46168
R10952 gnd.n5091 gnd.t221 4.46168
R10953 gnd.n5125 gnd.n1367 4.46168
R10954 gnd.n1426 gnd.n1425 4.46168
R10955 gnd.n5353 gnd.n5340 4.46111
R10956 gnd.n3466 gnd.n3462 4.38594
R10957 gnd.n3434 gnd.n3430 4.38594
R10958 gnd.n3402 gnd.n3398 4.38594
R10959 gnd.n3371 gnd.n3367 4.38594
R10960 gnd.n3339 gnd.n3335 4.38594
R10961 gnd.n3307 gnd.n3303 4.38594
R10962 gnd.n3275 gnd.n3271 4.38594
R10963 gnd.n3244 gnd.n3240 4.38594
R10964 gnd.n3477 gnd.n3455 4.26717
R10965 gnd.n3445 gnd.n3423 4.26717
R10966 gnd.n3413 gnd.n3391 4.26717
R10967 gnd.n3382 gnd.n3360 4.26717
R10968 gnd.n3350 gnd.n3328 4.26717
R10969 gnd.n3318 gnd.n3296 4.26717
R10970 gnd.n3286 gnd.n3264 4.26717
R10971 gnd.n3255 gnd.n3233 4.26717
R10972 gnd.n2934 gnd.t162 4.14303
R10973 gnd.n3165 gnd.t189 4.14303
R10974 gnd.t42 gnd.n986 4.14303
R10975 gnd.n4748 gnd.t235 4.14303
R10976 gnd.n4874 gnd.t219 4.14303
R10977 gnd.t35 gnd.n1138 4.14303
R10978 gnd.n3485 gnd.n3484 4.08274
R10979 gnd.n5486 gnd.n5485 4.05904
R10980 gnd.n1892 gnd.n1891 4.05904
R10981 gnd.n4356 gnd.n1833 4.05904
R10982 gnd.n5366 gnd.n5365 4.05904
R10983 gnd.n15 gnd.n7 3.99943
R10984 gnd.t116 gnd.n4477 3.82437
R10985 gnd.t222 gnd.n1733 3.82437
R10986 gnd.n1724 gnd.n1723 3.82437
R10987 gnd.n4534 gnd.n1684 3.82437
R10988 gnd.t237 gnd.n1647 3.82437
R10989 gnd.n1634 gnd.n1633 3.82437
R10990 gnd.n4750 gnd.n1599 3.82437
R10991 gnd.n1546 gnd.n1544 3.82437
R10992 gnd.n4895 gnd.n4894 3.82437
R10993 gnd.n4945 gnd.t160 3.82437
R10994 gnd.n5037 gnd.n5036 3.82437
R10995 gnd.n5081 gnd.n1399 3.82437
R10996 gnd.t221 gnd.n5090 3.82437
R10997 gnd.n1350 gnd.t39 3.82437
R10998 gnd.n3485 gnd.n3357 3.70378
R10999 gnd.n3007 gnd.n2428 3.65935
R11000 gnd.n15 gnd.n14 3.60163
R11001 gnd.t205 gnd.n3135 3.50571
R11002 gnd.n3476 gnd.n3457 3.49141
R11003 gnd.n3444 gnd.n3425 3.49141
R11004 gnd.n3412 gnd.n3393 3.49141
R11005 gnd.n3381 gnd.n3362 3.49141
R11006 gnd.n3349 gnd.n3330 3.49141
R11007 gnd.n3317 gnd.n3298 3.49141
R11008 gnd.n3285 gnd.n3266 3.49141
R11009 gnd.n3254 gnd.n3235 3.49141
R11010 gnd.n4423 gnd.n4422 3.18706
R11011 gnd.t32 gnd.n4500 3.18706
R11012 gnd.n4510 gnd.n1730 3.18706
R11013 gnd.n4597 gnd.n4596 3.18706
R11014 gnd.n4705 gnd.n1640 3.18706
R11015 gnd.n4774 gnd.n4773 3.18706
R11016 gnd.n4858 gnd.n1552 3.18706
R11017 gnd.n4961 gnd.n4960 3.18706
R11018 gnd.n5023 gnd.n5022 3.18706
R11019 gnd.n5099 gnd.n5098 3.18706
R11020 gnd.n5132 gnd.t90 3.18706
R11021 gnd.n5426 gnd.n1333 3.18706
R11022 gnd.n2513 gnd.t162 2.8684
R11023 gnd.n4543 gnd.t191 2.8684
R11024 gnd.n5047 gnd.t223 2.8684
R11025 gnd.n2416 gnd.t245 2.82907
R11026 gnd.n2416 gnd.t228 2.82907
R11027 gnd.n2418 gnd.t285 2.82907
R11028 gnd.n2418 gnd.t274 2.82907
R11029 gnd.n2420 gnd.t243 2.82907
R11030 gnd.n2420 gnd.t290 2.82907
R11031 gnd.n2422 gnd.t263 2.82907
R11032 gnd.n2422 gnd.t204 2.82907
R11033 gnd.n2424 gnd.t227 2.82907
R11034 gnd.n2424 gnd.t165 2.82907
R11035 gnd.n2393 gnd.t267 2.82907
R11036 gnd.n2393 gnd.t149 2.82907
R11037 gnd.n2395 gnd.t213 2.82907
R11038 gnd.n2395 gnd.t260 2.82907
R11039 gnd.n2397 gnd.t210 2.82907
R11040 gnd.n2397 gnd.t211 2.82907
R11041 gnd.n2399 gnd.t248 2.82907
R11042 gnd.n2399 gnd.t246 2.82907
R11043 gnd.n2401 gnd.t139 2.82907
R11044 gnd.n2401 gnd.t247 2.82907
R11045 gnd.n2404 gnd.t270 2.82907
R11046 gnd.n2404 gnd.t252 2.82907
R11047 gnd.n2406 gnd.t232 2.82907
R11048 gnd.n2406 gnd.t257 2.82907
R11049 gnd.n2408 gnd.t259 2.82907
R11050 gnd.n2408 gnd.t153 2.82907
R11051 gnd.n2410 gnd.t16 2.82907
R11052 gnd.n2410 gnd.t158 2.82907
R11053 gnd.n2412 gnd.t7 2.82907
R11054 gnd.n2412 gnd.t251 2.82907
R11055 gnd.n47 gnd.t193 2.82907
R11056 gnd.n47 gnd.t226 2.82907
R11057 gnd.n45 gnd.t9 2.82907
R11058 gnd.n45 gnd.t275 2.82907
R11059 gnd.n43 gnd.t182 2.82907
R11060 gnd.n43 gnd.t291 2.82907
R11061 gnd.n41 gnd.t242 2.82907
R11062 gnd.n41 gnd.t173 2.82907
R11063 gnd.n39 gnd.t156 2.82907
R11064 gnd.n39 gnd.t284 2.82907
R11065 gnd.n24 gnd.t129 2.82907
R11066 gnd.n24 gnd.t269 2.82907
R11067 gnd.n22 gnd.t186 2.82907
R11068 gnd.n22 gnd.t279 2.82907
R11069 gnd.n20 gnd.t253 2.82907
R11070 gnd.n20 gnd.t177 2.82907
R11071 gnd.n18 gnd.t271 2.82907
R11072 gnd.n18 gnd.t262 2.82907
R11073 gnd.n16 gnd.t215 2.82907
R11074 gnd.n16 gnd.t126 2.82907
R11075 gnd.n35 gnd.t14 2.82907
R11076 gnd.n35 gnd.t258 2.82907
R11077 gnd.n33 gnd.t214 2.82907
R11078 gnd.n33 gnd.t265 2.82907
R11079 gnd.n31 gnd.t207 2.82907
R11080 gnd.n31 gnd.t138 2.82907
R11081 gnd.n29 gnd.t266 2.82907
R11082 gnd.n29 gnd.t187 2.82907
R11083 gnd.n27 gnd.t147 2.82907
R11084 gnd.n27 gnd.t272 2.82907
R11085 gnd.n3473 gnd.n3472 2.71565
R11086 gnd.n3441 gnd.n3440 2.71565
R11087 gnd.n3409 gnd.n3408 2.71565
R11088 gnd.n3378 gnd.n3377 2.71565
R11089 gnd.n3346 gnd.n3345 2.71565
R11090 gnd.n3314 gnd.n3313 2.71565
R11091 gnd.n3282 gnd.n3281 2.71565
R11092 gnd.n3251 gnd.n3250 2.71565
R11093 gnd.n4443 gnd.t53 2.54975
R11094 gnd.n4509 gnd.n4507 2.54975
R11095 gnd.n1716 gnd.t132 2.54975
R11096 gnd.n4581 gnd.n4580 2.54975
R11097 gnd.n4644 gnd.t231 2.54975
R11098 gnd.n4704 gnd.n4703 2.54975
R11099 gnd.n4602 gnd.t180 2.54975
R11100 gnd.n4758 gnd.n1592 2.54975
R11101 gnd.n4857 gnd.n4856 2.54975
R11102 gnd.n4954 gnd.t183 2.54975
R11103 gnd.n4952 gnd.n1500 2.54975
R11104 gnd.n4938 gnd.t216 2.54975
R11105 gnd.n4988 gnd.n4987 2.54975
R11106 gnd.t240 gnd.n5074 2.54975
R11107 gnd.n5101 gnd.n1383 2.54975
R11108 gnd.n3007 gnd.n2429 2.27742
R11109 gnd.n3007 gnd.n2392 2.27742
R11110 gnd.n3007 gnd.n2391 2.27742
R11111 gnd.n3007 gnd.n2390 2.27742
R11112 gnd.n6943 gnd.n220 2.27742
R11113 gnd.n6943 gnd.n219 2.27742
R11114 gnd.n6943 gnd.n218 2.27742
R11115 gnd.n6943 gnd.n217 2.27742
R11116 gnd.n6943 gnd.n216 2.27742
R11117 gnd.n5747 gnd.n215 2.27742
R11118 gnd.n1173 gnd.n215 2.27742
R11119 gnd.n5787 gnd.n215 2.27742
R11120 gnd.n5805 gnd.n215 2.27742
R11121 gnd.n5790 gnd.n215 2.27742
R11122 gnd.n6049 gnd.n898 2.27742
R11123 gnd.n6050 gnd.n6049 2.27742
R11124 gnd.n6049 gnd.n904 2.27742
R11125 gnd.n6049 gnd.n903 2.27742
R11126 gnd.n6049 gnd.n902 2.27742
R11127 gnd.n2115 gnd.n901 2.27742
R11128 gnd.n3954 gnd.n901 2.27742
R11129 gnd.n3961 gnd.n901 2.27742
R11130 gnd.n3956 gnd.n901 2.27742
R11131 gnd.n2067 gnd.n901 2.27742
R11132 gnd.n2861 gnd.t28 2.23109
R11133 gnd.n2484 gnd.t188 2.23109
R11134 gnd.n4662 gnd.t235 2.23109
R11135 gnd.n4836 gnd.t219 2.23109
R11136 gnd.n3469 gnd.n3459 1.93989
R11137 gnd.n3437 gnd.n3427 1.93989
R11138 gnd.n3405 gnd.n3395 1.93989
R11139 gnd.n3374 gnd.n3364 1.93989
R11140 gnd.n3342 gnd.n3332 1.93989
R11141 gnd.n3310 gnd.n3300 1.93989
R11142 gnd.n3278 gnd.n3268 1.93989
R11143 gnd.n3247 gnd.n3237 1.93989
R11144 gnd.n4519 gnd.n4518 1.91244
R11145 gnd.n4588 gnd.n4587 1.91244
R11146 gnd.n4765 gnd.n4764 1.91244
R11147 gnd.n4867 gnd.n4866 1.91244
R11148 gnd.n5038 gnd.n1454 1.91244
R11149 gnd.n1442 gnd.n1441 1.91244
R11150 gnd.n1425 gnd.t18 1.91244
R11151 gnd.t286 gnd.n2872 1.59378
R11152 gnd.n3051 gnd.t194 1.59378
R11153 gnd.n2325 gnd.t175 1.59378
R11154 gnd.t4 gnd.n4713 1.59378
R11155 gnd.n4896 gnd.t200 1.59378
R11156 gnd.t25 gnd.n4450 1.27512
R11157 gnd.n4450 gnd.n1758 1.27512
R11158 gnd.n4436 gnd.n4435 1.27512
R11159 gnd.t159 gnd.n4625 1.27512
R11160 gnd.n4624 gnd.n1668 1.27512
R11161 gnd.n4610 gnd.n4609 1.27512
R11162 gnd.n4801 gnd.n1582 1.27512
R11163 gnd.n4788 gnd.n4787 1.27512
R11164 gnd.n4973 gnd.n4972 1.27512
R11165 gnd.n5011 gnd.n5010 1.27512
R11166 gnd.t0 gnd.n1475 1.27512
R11167 gnd.n5110 gnd.n5109 1.27512
R11168 gnd.n5336 gnd.n1338 1.27512
R11169 gnd.n2714 gnd.n2706 1.16414
R11170 gnd.n3531 gnd.n2228 1.16414
R11171 gnd.n3468 gnd.n3461 1.16414
R11172 gnd.n3436 gnd.n3429 1.16414
R11173 gnd.n3404 gnd.n3397 1.16414
R11174 gnd.n3373 gnd.n3366 1.16414
R11175 gnd.n3341 gnd.n3334 1.16414
R11176 gnd.n3309 gnd.n3302 1.16414
R11177 gnd.n3277 gnd.n3270 1.16414
R11178 gnd.n3246 gnd.n3239 1.16414
R11179 gnd.n5554 gnd.n1289 0.970197
R11180 gnd.n4344 gnd.n1898 0.970197
R11181 gnd.n3452 gnd.n3420 0.962709
R11182 gnd.n3484 gnd.n3452 0.962709
R11183 gnd.n3325 gnd.n3293 0.962709
R11184 gnd.n3357 gnd.n3325 0.962709
R11185 gnd.n2960 gnd.t184 0.956468
R11186 gnd.n3125 gnd.t128 0.956468
R11187 gnd.t233 gnd.n840 0.956468
R11188 gnd.n6078 gnd.t6 0.956468
R11189 gnd.n4079 gnd.t244 0.956468
R11190 gnd.n4041 gnd.t148 0.956468
R11191 gnd.n4444 gnd.t166 0.956468
R11192 gnd.t281 gnd.n4509 0.956468
R11193 gnd.n5101 gnd.t2 0.956468
R11194 gnd.n1428 gnd.t202 0.956468
R11195 gnd.n5719 gnd.t146 0.956468
R11196 gnd.n1222 gnd.t125 0.956468
R11197 gnd.n266 gnd.t225 0.956468
R11198 gnd.t140 gnd.n177 0.956468
R11199 gnd.n2423 gnd.n2421 0.773756
R11200 gnd.n46 gnd.n44 0.773756
R11201 gnd.n2426 gnd.n2425 0.773756
R11202 gnd.n2425 gnd.n2423 0.773756
R11203 gnd.n2421 gnd.n2419 0.773756
R11204 gnd.n2419 gnd.n2417 0.773756
R11205 gnd.n42 gnd.n40 0.773756
R11206 gnd.n44 gnd.n42 0.773756
R11207 gnd.n48 gnd.n46 0.773756
R11208 gnd.n49 gnd.n48 0.773756
R11209 gnd.n2 gnd.n1 0.672012
R11210 gnd.n3 gnd.n2 0.672012
R11211 gnd.n4 gnd.n3 0.672012
R11212 gnd.n5 gnd.n4 0.672012
R11213 gnd.n6 gnd.n5 0.672012
R11214 gnd.n7 gnd.n6 0.672012
R11215 gnd.n9 gnd.n8 0.672012
R11216 gnd.n10 gnd.n9 0.672012
R11217 gnd.n11 gnd.n10 0.672012
R11218 gnd.n12 gnd.n11 0.672012
R11219 gnd.n13 gnd.n12 0.672012
R11220 gnd.n14 gnd.n13 0.672012
R11221 gnd.n4471 gnd.t64 0.637812
R11222 gnd.n4547 gnd.n1710 0.637812
R11223 gnd.n4555 gnd.n1704 0.637812
R11224 gnd.n1704 gnd.t196 0.637812
R11225 gnd.n4732 gnd.n1619 0.637812
R11226 gnd.n4740 gnd.n1613 0.637812
R11227 gnd.n4756 gnd.t10 0.637812
R11228 gnd.n4779 gnd.t239 0.637812
R11229 gnd.n4886 gnd.n1532 0.637812
R11230 gnd.n4902 gnd.n1525 0.637812
R11231 gnd.t1 gnd.n5056 0.637812
R11232 gnd.n5056 gnd.n1412 0.637812
R11233 gnd.n5075 gnd.n1403 0.637812
R11234 gnd.n5132 gnd.t46 0.637812
R11235 gnd.n2403 gnd.n2402 0.573776
R11236 gnd.n2402 gnd.n2400 0.573776
R11237 gnd.n2400 gnd.n2398 0.573776
R11238 gnd.n2398 gnd.n2396 0.573776
R11239 gnd.n2396 gnd.n2394 0.573776
R11240 gnd.n2414 gnd.n2413 0.573776
R11241 gnd.n2413 gnd.n2411 0.573776
R11242 gnd.n2411 gnd.n2409 0.573776
R11243 gnd.n2409 gnd.n2407 0.573776
R11244 gnd.n2407 gnd.n2405 0.573776
R11245 gnd.n19 gnd.n17 0.573776
R11246 gnd.n21 gnd.n19 0.573776
R11247 gnd.n23 gnd.n21 0.573776
R11248 gnd.n25 gnd.n23 0.573776
R11249 gnd.n26 gnd.n25 0.573776
R11250 gnd.n30 gnd.n28 0.573776
R11251 gnd.n32 gnd.n30 0.573776
R11252 gnd.n34 gnd.n32 0.573776
R11253 gnd.n36 gnd.n34 0.573776
R11254 gnd.n37 gnd.n36 0.573776
R11255 gnd gnd.n0 0.551497
R11256 gnd.n6943 gnd.n215 0.548625
R11257 gnd.n6049 gnd.n901 0.548625
R11258 gnd.n3696 gnd.n3695 0.532512
R11259 gnd.n3846 gnd.n3845 0.532512
R11260 gnd.n7053 gnd.n7052 0.532512
R11261 gnd.n7153 gnd.n78 0.532512
R11262 gnd.n5993 gnd.n5992 0.523366
R11263 gnd.n5201 gnd.n1104 0.523366
R11264 gnd.n7147 gnd.n7146 0.520317
R11265 gnd.n7076 gnd.n7075 0.520317
R11266 gnd.n5608 gnd.n5607 0.520317
R11267 gnd.n5512 gnd.n1133 0.520317
R11268 gnd.n1919 gnd.n991 0.520317
R11269 gnd.n4304 gnd.n4303 0.520317
R11270 gnd.n3765 gnd.n3744 0.520317
R11271 gnd.n3701 gnd.n2148 0.520317
R11272 gnd.n5323 gnd.n5322 0.489829
R11273 gnd.n4277 gnd.n4276 0.489829
R11274 gnd.n3188 gnd.n2232 0.486781
R11275 gnd.n2763 gnd.n2762 0.48678
R11276 gnd.n3505 gnd.n2186 0.480683
R11277 gnd.n2847 gnd.n2846 0.480683
R11278 gnd.n6263 gnd.n6262 0.480683
R11279 gnd.n6683 gnd.n6682 0.480683
R11280 gnd.n6896 gnd.n6895 0.480683
R11281 gnd.n3906 gnd.n825 0.480683
R11282 gnd.n7186 gnd.n7185 0.470187
R11283 gnd.n5995 gnd.n5994 0.432431
R11284 gnd.n5204 gnd.n5203 0.432431
R11285 gnd.n4284 gnd.n2012 0.388379
R11286 gnd.n3465 gnd.n3464 0.388379
R11287 gnd.n3433 gnd.n3432 0.388379
R11288 gnd.n3401 gnd.n3400 0.388379
R11289 gnd.n3370 gnd.n3369 0.388379
R11290 gnd.n3338 gnd.n3337 0.388379
R11291 gnd.n3306 gnd.n3305 0.388379
R11292 gnd.n3274 gnd.n3273 0.388379
R11293 gnd.n3243 gnd.n3242 0.388379
R11294 gnd.n7116 gnd.n7115 0.388379
R11295 gnd.n3806 gnd.n3805 0.388379
R11296 gnd.n5312 gnd.n5311 0.388379
R11297 gnd.n7186 gnd.n15 0.374463
R11298 gnd.n2287 gnd.t161 0.319156
R11299 gnd.n3928 gnd.t15 0.319156
R11300 gnd.n6054 gnd.t157 0.319156
R11301 gnd.t152 gnd.n2077 0.319156
R11302 gnd.t212 gnd.n4012 0.319156
R11303 gnd.n4414 gnd.t93 0.319156
R11304 gnd.n4714 gnd.t4 0.319156
R11305 gnd.t208 gnd.t130 0.319156
R11306 gnd.t288 gnd.t280 0.319156
R11307 gnd.n4926 gnd.t200 0.319156
R11308 gnd.n5328 gnd.t77 0.319156
R11309 gnd.n5650 gnd.t172 0.319156
R11310 gnd.n5783 gnd.t181 0.319156
R11311 gnd.n6921 gnd.t8 0.319156
R11312 gnd.t264 gnd.n209 0.319156
R11313 gnd.n2681 gnd.n2659 0.311721
R11314 gnd.n4295 gnd.n4294 0.302329
R11315 gnd.n5291 gnd.n1264 0.302329
R11316 gnd gnd.n7186 0.295112
R11317 gnd.n3576 gnd.n3575 0.268793
R11318 gnd.n3575 gnd.n3574 0.241354
R11319 gnd.n5555 gnd.n1290 0.229039
R11320 gnd.n5556 gnd.n5555 0.229039
R11321 gnd.n4343 gnd.n1903 0.229039
R11322 gnd.n4343 gnd.n4342 0.229039
R11323 gnd.n2835 gnd.n2634 0.206293
R11324 gnd.n3482 gnd.n3454 0.155672
R11325 gnd.n3475 gnd.n3454 0.155672
R11326 gnd.n3475 gnd.n3474 0.155672
R11327 gnd.n3474 gnd.n3458 0.155672
R11328 gnd.n3467 gnd.n3458 0.155672
R11329 gnd.n3467 gnd.n3466 0.155672
R11330 gnd.n3450 gnd.n3422 0.155672
R11331 gnd.n3443 gnd.n3422 0.155672
R11332 gnd.n3443 gnd.n3442 0.155672
R11333 gnd.n3442 gnd.n3426 0.155672
R11334 gnd.n3435 gnd.n3426 0.155672
R11335 gnd.n3435 gnd.n3434 0.155672
R11336 gnd.n3418 gnd.n3390 0.155672
R11337 gnd.n3411 gnd.n3390 0.155672
R11338 gnd.n3411 gnd.n3410 0.155672
R11339 gnd.n3410 gnd.n3394 0.155672
R11340 gnd.n3403 gnd.n3394 0.155672
R11341 gnd.n3403 gnd.n3402 0.155672
R11342 gnd.n3387 gnd.n3359 0.155672
R11343 gnd.n3380 gnd.n3359 0.155672
R11344 gnd.n3380 gnd.n3379 0.155672
R11345 gnd.n3379 gnd.n3363 0.155672
R11346 gnd.n3372 gnd.n3363 0.155672
R11347 gnd.n3372 gnd.n3371 0.155672
R11348 gnd.n3355 gnd.n3327 0.155672
R11349 gnd.n3348 gnd.n3327 0.155672
R11350 gnd.n3348 gnd.n3347 0.155672
R11351 gnd.n3347 gnd.n3331 0.155672
R11352 gnd.n3340 gnd.n3331 0.155672
R11353 gnd.n3340 gnd.n3339 0.155672
R11354 gnd.n3323 gnd.n3295 0.155672
R11355 gnd.n3316 gnd.n3295 0.155672
R11356 gnd.n3316 gnd.n3315 0.155672
R11357 gnd.n3315 gnd.n3299 0.155672
R11358 gnd.n3308 gnd.n3299 0.155672
R11359 gnd.n3308 gnd.n3307 0.155672
R11360 gnd.n3291 gnd.n3263 0.155672
R11361 gnd.n3284 gnd.n3263 0.155672
R11362 gnd.n3284 gnd.n3283 0.155672
R11363 gnd.n3283 gnd.n3267 0.155672
R11364 gnd.n3276 gnd.n3267 0.155672
R11365 gnd.n3276 gnd.n3275 0.155672
R11366 gnd.n3260 gnd.n3232 0.155672
R11367 gnd.n3253 gnd.n3232 0.155672
R11368 gnd.n3253 gnd.n3252 0.155672
R11369 gnd.n3252 gnd.n3236 0.155672
R11370 gnd.n3245 gnd.n3236 0.155672
R11371 gnd.n3245 gnd.n3244 0.155672
R11372 gnd.n3607 gnd.n2186 0.152939
R11373 gnd.n3607 gnd.n3606 0.152939
R11374 gnd.n3606 gnd.n3605 0.152939
R11375 gnd.n3605 gnd.n2188 0.152939
R11376 gnd.n2189 gnd.n2188 0.152939
R11377 gnd.n2190 gnd.n2189 0.152939
R11378 gnd.n2191 gnd.n2190 0.152939
R11379 gnd.n2192 gnd.n2191 0.152939
R11380 gnd.n2193 gnd.n2192 0.152939
R11381 gnd.n2194 gnd.n2193 0.152939
R11382 gnd.n2195 gnd.n2194 0.152939
R11383 gnd.n2196 gnd.n2195 0.152939
R11384 gnd.n2197 gnd.n2196 0.152939
R11385 gnd.n2198 gnd.n2197 0.152939
R11386 gnd.n3577 gnd.n2198 0.152939
R11387 gnd.n3577 gnd.n3576 0.152939
R11388 gnd.n2848 gnd.n2847 0.152939
R11389 gnd.n2848 gnd.n2552 0.152939
R11390 gnd.n2876 gnd.n2552 0.152939
R11391 gnd.n2877 gnd.n2876 0.152939
R11392 gnd.n2878 gnd.n2877 0.152939
R11393 gnd.n2879 gnd.n2878 0.152939
R11394 gnd.n2879 gnd.n2524 0.152939
R11395 gnd.n2906 gnd.n2524 0.152939
R11396 gnd.n2907 gnd.n2906 0.152939
R11397 gnd.n2908 gnd.n2907 0.152939
R11398 gnd.n2908 gnd.n2502 0.152939
R11399 gnd.n2937 gnd.n2502 0.152939
R11400 gnd.n2938 gnd.n2937 0.152939
R11401 gnd.n2939 gnd.n2938 0.152939
R11402 gnd.n2940 gnd.n2939 0.152939
R11403 gnd.n2942 gnd.n2940 0.152939
R11404 gnd.n2942 gnd.n2941 0.152939
R11405 gnd.n2941 gnd.n2451 0.152939
R11406 gnd.n2452 gnd.n2451 0.152939
R11407 gnd.n2453 gnd.n2452 0.152939
R11408 gnd.n2472 gnd.n2453 0.152939
R11409 gnd.n2473 gnd.n2472 0.152939
R11410 gnd.n2473 gnd.n2383 0.152939
R11411 gnd.n3032 gnd.n2383 0.152939
R11412 gnd.n3033 gnd.n3032 0.152939
R11413 gnd.n3034 gnd.n3033 0.152939
R11414 gnd.n3035 gnd.n3034 0.152939
R11415 gnd.n3035 gnd.n2356 0.152939
R11416 gnd.n3072 gnd.n2356 0.152939
R11417 gnd.n3073 gnd.n3072 0.152939
R11418 gnd.n3074 gnd.n3073 0.152939
R11419 gnd.n3075 gnd.n3074 0.152939
R11420 gnd.n3075 gnd.n2329 0.152939
R11421 gnd.n3117 gnd.n2329 0.152939
R11422 gnd.n3118 gnd.n3117 0.152939
R11423 gnd.n3119 gnd.n3118 0.152939
R11424 gnd.n3120 gnd.n3119 0.152939
R11425 gnd.n3120 gnd.n2301 0.152939
R11426 gnd.n3158 gnd.n2301 0.152939
R11427 gnd.n3159 gnd.n3158 0.152939
R11428 gnd.n3160 gnd.n3159 0.152939
R11429 gnd.n3161 gnd.n3160 0.152939
R11430 gnd.n3161 gnd.n2274 0.152939
R11431 gnd.n3207 gnd.n2274 0.152939
R11432 gnd.n3208 gnd.n3207 0.152939
R11433 gnd.n3209 gnd.n3208 0.152939
R11434 gnd.n3210 gnd.n3209 0.152939
R11435 gnd.n3210 gnd.n2247 0.152939
R11436 gnd.n3501 gnd.n2247 0.152939
R11437 gnd.n3502 gnd.n3501 0.152939
R11438 gnd.n3503 gnd.n3502 0.152939
R11439 gnd.n3504 gnd.n3503 0.152939
R11440 gnd.n3505 gnd.n3504 0.152939
R11441 gnd.n2846 gnd.n2576 0.152939
R11442 gnd.n2597 gnd.n2576 0.152939
R11443 gnd.n2598 gnd.n2597 0.152939
R11444 gnd.n2604 gnd.n2598 0.152939
R11445 gnd.n2605 gnd.n2604 0.152939
R11446 gnd.n2606 gnd.n2605 0.152939
R11447 gnd.n2606 gnd.n2595 0.152939
R11448 gnd.n2614 gnd.n2595 0.152939
R11449 gnd.n2615 gnd.n2614 0.152939
R11450 gnd.n2616 gnd.n2615 0.152939
R11451 gnd.n2616 gnd.n2593 0.152939
R11452 gnd.n2624 gnd.n2593 0.152939
R11453 gnd.n2625 gnd.n2624 0.152939
R11454 gnd.n2626 gnd.n2625 0.152939
R11455 gnd.n2626 gnd.n2591 0.152939
R11456 gnd.n2634 gnd.n2591 0.152939
R11457 gnd.n3574 gnd.n2203 0.152939
R11458 gnd.n2205 gnd.n2203 0.152939
R11459 gnd.n2206 gnd.n2205 0.152939
R11460 gnd.n2207 gnd.n2206 0.152939
R11461 gnd.n2208 gnd.n2207 0.152939
R11462 gnd.n2209 gnd.n2208 0.152939
R11463 gnd.n2210 gnd.n2209 0.152939
R11464 gnd.n2211 gnd.n2210 0.152939
R11465 gnd.n2212 gnd.n2211 0.152939
R11466 gnd.n2213 gnd.n2212 0.152939
R11467 gnd.n2214 gnd.n2213 0.152939
R11468 gnd.n2215 gnd.n2214 0.152939
R11469 gnd.n2216 gnd.n2215 0.152939
R11470 gnd.n2217 gnd.n2216 0.152939
R11471 gnd.n2218 gnd.n2217 0.152939
R11472 gnd.n2219 gnd.n2218 0.152939
R11473 gnd.n2220 gnd.n2219 0.152939
R11474 gnd.n2221 gnd.n2220 0.152939
R11475 gnd.n2222 gnd.n2221 0.152939
R11476 gnd.n2223 gnd.n2222 0.152939
R11477 gnd.n2224 gnd.n2223 0.152939
R11478 gnd.n2225 gnd.n2224 0.152939
R11479 gnd.n2229 gnd.n2225 0.152939
R11480 gnd.n2230 gnd.n2229 0.152939
R11481 gnd.n2231 gnd.n2230 0.152939
R11482 gnd.n2232 gnd.n2231 0.152939
R11483 gnd.n3009 gnd.n3008 0.152939
R11484 gnd.n3010 gnd.n3009 0.152939
R11485 gnd.n3011 gnd.n3010 0.152939
R11486 gnd.n3012 gnd.n3011 0.152939
R11487 gnd.n3013 gnd.n3012 0.152939
R11488 gnd.n3014 gnd.n3013 0.152939
R11489 gnd.n3014 gnd.n2337 0.152939
R11490 gnd.n3093 gnd.n2337 0.152939
R11491 gnd.n3094 gnd.n3093 0.152939
R11492 gnd.n3095 gnd.n3094 0.152939
R11493 gnd.n3096 gnd.n3095 0.152939
R11494 gnd.n3097 gnd.n3096 0.152939
R11495 gnd.n3098 gnd.n3097 0.152939
R11496 gnd.n3099 gnd.n3098 0.152939
R11497 gnd.n3100 gnd.n3099 0.152939
R11498 gnd.n3101 gnd.n3100 0.152939
R11499 gnd.n3101 gnd.n2281 0.152939
R11500 gnd.n3179 gnd.n2281 0.152939
R11501 gnd.n3180 gnd.n3179 0.152939
R11502 gnd.n3181 gnd.n3180 0.152939
R11503 gnd.n3182 gnd.n3181 0.152939
R11504 gnd.n3183 gnd.n3182 0.152939
R11505 gnd.n3184 gnd.n3183 0.152939
R11506 gnd.n3185 gnd.n3184 0.152939
R11507 gnd.n3186 gnd.n3185 0.152939
R11508 gnd.n3187 gnd.n3186 0.152939
R11509 gnd.n3189 gnd.n3187 0.152939
R11510 gnd.n3189 gnd.n3188 0.152939
R11511 gnd.n2764 gnd.n2763 0.152939
R11512 gnd.n2764 gnd.n2654 0.152939
R11513 gnd.n2779 gnd.n2654 0.152939
R11514 gnd.n2780 gnd.n2779 0.152939
R11515 gnd.n2781 gnd.n2780 0.152939
R11516 gnd.n2781 gnd.n2642 0.152939
R11517 gnd.n2795 gnd.n2642 0.152939
R11518 gnd.n2796 gnd.n2795 0.152939
R11519 gnd.n2797 gnd.n2796 0.152939
R11520 gnd.n2798 gnd.n2797 0.152939
R11521 gnd.n2799 gnd.n2798 0.152939
R11522 gnd.n2800 gnd.n2799 0.152939
R11523 gnd.n2801 gnd.n2800 0.152939
R11524 gnd.n2802 gnd.n2801 0.152939
R11525 gnd.n2803 gnd.n2802 0.152939
R11526 gnd.n2804 gnd.n2803 0.152939
R11527 gnd.n2805 gnd.n2804 0.152939
R11528 gnd.n2806 gnd.n2805 0.152939
R11529 gnd.n2807 gnd.n2806 0.152939
R11530 gnd.n2808 gnd.n2807 0.152939
R11531 gnd.n2809 gnd.n2808 0.152939
R11532 gnd.n2809 gnd.n2508 0.152939
R11533 gnd.n2926 gnd.n2508 0.152939
R11534 gnd.n2927 gnd.n2926 0.152939
R11535 gnd.n2928 gnd.n2927 0.152939
R11536 gnd.n2929 gnd.n2928 0.152939
R11537 gnd.n2929 gnd.n2430 0.152939
R11538 gnd.n3006 gnd.n2430 0.152939
R11539 gnd.n2682 gnd.n2681 0.152939
R11540 gnd.n2683 gnd.n2682 0.152939
R11541 gnd.n2684 gnd.n2683 0.152939
R11542 gnd.n2685 gnd.n2684 0.152939
R11543 gnd.n2686 gnd.n2685 0.152939
R11544 gnd.n2687 gnd.n2686 0.152939
R11545 gnd.n2688 gnd.n2687 0.152939
R11546 gnd.n2689 gnd.n2688 0.152939
R11547 gnd.n2690 gnd.n2689 0.152939
R11548 gnd.n2691 gnd.n2690 0.152939
R11549 gnd.n2692 gnd.n2691 0.152939
R11550 gnd.n2693 gnd.n2692 0.152939
R11551 gnd.n2694 gnd.n2693 0.152939
R11552 gnd.n2695 gnd.n2694 0.152939
R11553 gnd.n2696 gnd.n2695 0.152939
R11554 gnd.n2697 gnd.n2696 0.152939
R11555 gnd.n2698 gnd.n2697 0.152939
R11556 gnd.n2699 gnd.n2698 0.152939
R11557 gnd.n2700 gnd.n2699 0.152939
R11558 gnd.n2701 gnd.n2700 0.152939
R11559 gnd.n2702 gnd.n2701 0.152939
R11560 gnd.n2703 gnd.n2702 0.152939
R11561 gnd.n2707 gnd.n2703 0.152939
R11562 gnd.n2708 gnd.n2707 0.152939
R11563 gnd.n2708 gnd.n2665 0.152939
R11564 gnd.n2762 gnd.n2665 0.152939
R11565 gnd.n6264 gnd.n6263 0.152939
R11566 gnd.n6264 gnd.n652 0.152939
R11567 gnd.n6272 gnd.n652 0.152939
R11568 gnd.n6273 gnd.n6272 0.152939
R11569 gnd.n6274 gnd.n6273 0.152939
R11570 gnd.n6274 gnd.n646 0.152939
R11571 gnd.n6282 gnd.n646 0.152939
R11572 gnd.n6283 gnd.n6282 0.152939
R11573 gnd.n6284 gnd.n6283 0.152939
R11574 gnd.n6284 gnd.n640 0.152939
R11575 gnd.n6292 gnd.n640 0.152939
R11576 gnd.n6293 gnd.n6292 0.152939
R11577 gnd.n6294 gnd.n6293 0.152939
R11578 gnd.n6294 gnd.n634 0.152939
R11579 gnd.n6302 gnd.n634 0.152939
R11580 gnd.n6303 gnd.n6302 0.152939
R11581 gnd.n6304 gnd.n6303 0.152939
R11582 gnd.n6304 gnd.n628 0.152939
R11583 gnd.n6312 gnd.n628 0.152939
R11584 gnd.n6313 gnd.n6312 0.152939
R11585 gnd.n6314 gnd.n6313 0.152939
R11586 gnd.n6314 gnd.n622 0.152939
R11587 gnd.n6322 gnd.n622 0.152939
R11588 gnd.n6323 gnd.n6322 0.152939
R11589 gnd.n6324 gnd.n6323 0.152939
R11590 gnd.n6324 gnd.n616 0.152939
R11591 gnd.n6332 gnd.n616 0.152939
R11592 gnd.n6333 gnd.n6332 0.152939
R11593 gnd.n6334 gnd.n6333 0.152939
R11594 gnd.n6334 gnd.n610 0.152939
R11595 gnd.n6342 gnd.n610 0.152939
R11596 gnd.n6343 gnd.n6342 0.152939
R11597 gnd.n6344 gnd.n6343 0.152939
R11598 gnd.n6344 gnd.n604 0.152939
R11599 gnd.n6352 gnd.n604 0.152939
R11600 gnd.n6353 gnd.n6352 0.152939
R11601 gnd.n6354 gnd.n6353 0.152939
R11602 gnd.n6354 gnd.n598 0.152939
R11603 gnd.n6362 gnd.n598 0.152939
R11604 gnd.n6363 gnd.n6362 0.152939
R11605 gnd.n6364 gnd.n6363 0.152939
R11606 gnd.n6364 gnd.n592 0.152939
R11607 gnd.n6372 gnd.n592 0.152939
R11608 gnd.n6373 gnd.n6372 0.152939
R11609 gnd.n6374 gnd.n6373 0.152939
R11610 gnd.n6374 gnd.n586 0.152939
R11611 gnd.n6382 gnd.n586 0.152939
R11612 gnd.n6383 gnd.n6382 0.152939
R11613 gnd.n6384 gnd.n6383 0.152939
R11614 gnd.n6384 gnd.n580 0.152939
R11615 gnd.n6392 gnd.n580 0.152939
R11616 gnd.n6393 gnd.n6392 0.152939
R11617 gnd.n6394 gnd.n6393 0.152939
R11618 gnd.n6394 gnd.n574 0.152939
R11619 gnd.n6402 gnd.n574 0.152939
R11620 gnd.n6403 gnd.n6402 0.152939
R11621 gnd.n6404 gnd.n6403 0.152939
R11622 gnd.n6404 gnd.n568 0.152939
R11623 gnd.n6412 gnd.n568 0.152939
R11624 gnd.n6413 gnd.n6412 0.152939
R11625 gnd.n6414 gnd.n6413 0.152939
R11626 gnd.n6414 gnd.n562 0.152939
R11627 gnd.n6422 gnd.n562 0.152939
R11628 gnd.n6423 gnd.n6422 0.152939
R11629 gnd.n6424 gnd.n6423 0.152939
R11630 gnd.n6424 gnd.n556 0.152939
R11631 gnd.n6432 gnd.n556 0.152939
R11632 gnd.n6433 gnd.n6432 0.152939
R11633 gnd.n6434 gnd.n6433 0.152939
R11634 gnd.n6434 gnd.n550 0.152939
R11635 gnd.n6442 gnd.n550 0.152939
R11636 gnd.n6443 gnd.n6442 0.152939
R11637 gnd.n6444 gnd.n6443 0.152939
R11638 gnd.n6444 gnd.n544 0.152939
R11639 gnd.n6452 gnd.n544 0.152939
R11640 gnd.n6453 gnd.n6452 0.152939
R11641 gnd.n6454 gnd.n6453 0.152939
R11642 gnd.n6454 gnd.n538 0.152939
R11643 gnd.n6462 gnd.n538 0.152939
R11644 gnd.n6463 gnd.n6462 0.152939
R11645 gnd.n6464 gnd.n6463 0.152939
R11646 gnd.n6464 gnd.n532 0.152939
R11647 gnd.n6472 gnd.n532 0.152939
R11648 gnd.n6473 gnd.n6472 0.152939
R11649 gnd.n6474 gnd.n6473 0.152939
R11650 gnd.n6474 gnd.n526 0.152939
R11651 gnd.n6482 gnd.n526 0.152939
R11652 gnd.n6483 gnd.n6482 0.152939
R11653 gnd.n6484 gnd.n6483 0.152939
R11654 gnd.n6484 gnd.n520 0.152939
R11655 gnd.n6492 gnd.n520 0.152939
R11656 gnd.n6493 gnd.n6492 0.152939
R11657 gnd.n6494 gnd.n6493 0.152939
R11658 gnd.n6494 gnd.n514 0.152939
R11659 gnd.n6502 gnd.n514 0.152939
R11660 gnd.n6503 gnd.n6502 0.152939
R11661 gnd.n6504 gnd.n6503 0.152939
R11662 gnd.n6504 gnd.n508 0.152939
R11663 gnd.n6512 gnd.n508 0.152939
R11664 gnd.n6513 gnd.n6512 0.152939
R11665 gnd.n6514 gnd.n6513 0.152939
R11666 gnd.n6514 gnd.n502 0.152939
R11667 gnd.n6522 gnd.n502 0.152939
R11668 gnd.n6523 gnd.n6522 0.152939
R11669 gnd.n6524 gnd.n6523 0.152939
R11670 gnd.n6524 gnd.n496 0.152939
R11671 gnd.n6532 gnd.n496 0.152939
R11672 gnd.n6533 gnd.n6532 0.152939
R11673 gnd.n6534 gnd.n6533 0.152939
R11674 gnd.n6534 gnd.n490 0.152939
R11675 gnd.n6542 gnd.n490 0.152939
R11676 gnd.n6543 gnd.n6542 0.152939
R11677 gnd.n6544 gnd.n6543 0.152939
R11678 gnd.n6544 gnd.n484 0.152939
R11679 gnd.n6552 gnd.n484 0.152939
R11680 gnd.n6553 gnd.n6552 0.152939
R11681 gnd.n6554 gnd.n6553 0.152939
R11682 gnd.n6554 gnd.n478 0.152939
R11683 gnd.n6562 gnd.n478 0.152939
R11684 gnd.n6563 gnd.n6562 0.152939
R11685 gnd.n6564 gnd.n6563 0.152939
R11686 gnd.n6564 gnd.n472 0.152939
R11687 gnd.n6572 gnd.n472 0.152939
R11688 gnd.n6573 gnd.n6572 0.152939
R11689 gnd.n6574 gnd.n6573 0.152939
R11690 gnd.n6574 gnd.n466 0.152939
R11691 gnd.n6582 gnd.n466 0.152939
R11692 gnd.n6583 gnd.n6582 0.152939
R11693 gnd.n6584 gnd.n6583 0.152939
R11694 gnd.n6584 gnd.n460 0.152939
R11695 gnd.n6592 gnd.n460 0.152939
R11696 gnd.n6593 gnd.n6592 0.152939
R11697 gnd.n6594 gnd.n6593 0.152939
R11698 gnd.n6594 gnd.n454 0.152939
R11699 gnd.n6602 gnd.n454 0.152939
R11700 gnd.n6603 gnd.n6602 0.152939
R11701 gnd.n6604 gnd.n6603 0.152939
R11702 gnd.n6604 gnd.n448 0.152939
R11703 gnd.n6612 gnd.n448 0.152939
R11704 gnd.n6613 gnd.n6612 0.152939
R11705 gnd.n6614 gnd.n6613 0.152939
R11706 gnd.n6614 gnd.n442 0.152939
R11707 gnd.n6622 gnd.n442 0.152939
R11708 gnd.n6623 gnd.n6622 0.152939
R11709 gnd.n6624 gnd.n6623 0.152939
R11710 gnd.n6624 gnd.n436 0.152939
R11711 gnd.n6632 gnd.n436 0.152939
R11712 gnd.n6633 gnd.n6632 0.152939
R11713 gnd.n6634 gnd.n6633 0.152939
R11714 gnd.n6634 gnd.n430 0.152939
R11715 gnd.n6642 gnd.n430 0.152939
R11716 gnd.n6643 gnd.n6642 0.152939
R11717 gnd.n6644 gnd.n6643 0.152939
R11718 gnd.n6644 gnd.n424 0.152939
R11719 gnd.n6652 gnd.n424 0.152939
R11720 gnd.n6653 gnd.n6652 0.152939
R11721 gnd.n6654 gnd.n6653 0.152939
R11722 gnd.n6654 gnd.n418 0.152939
R11723 gnd.n6662 gnd.n418 0.152939
R11724 gnd.n6663 gnd.n6662 0.152939
R11725 gnd.n6664 gnd.n6663 0.152939
R11726 gnd.n6664 gnd.n412 0.152939
R11727 gnd.n6672 gnd.n412 0.152939
R11728 gnd.n6673 gnd.n6672 0.152939
R11729 gnd.n6674 gnd.n6673 0.152939
R11730 gnd.n6674 gnd.n406 0.152939
R11731 gnd.n6682 gnd.n406 0.152939
R11732 gnd.n6684 gnd.n6683 0.152939
R11733 gnd.n6684 gnd.n400 0.152939
R11734 gnd.n6692 gnd.n400 0.152939
R11735 gnd.n6693 gnd.n6692 0.152939
R11736 gnd.n6694 gnd.n6693 0.152939
R11737 gnd.n6694 gnd.n394 0.152939
R11738 gnd.n6702 gnd.n394 0.152939
R11739 gnd.n6703 gnd.n6702 0.152939
R11740 gnd.n6704 gnd.n6703 0.152939
R11741 gnd.n6704 gnd.n388 0.152939
R11742 gnd.n6712 gnd.n388 0.152939
R11743 gnd.n6713 gnd.n6712 0.152939
R11744 gnd.n6714 gnd.n6713 0.152939
R11745 gnd.n6714 gnd.n382 0.152939
R11746 gnd.n6722 gnd.n382 0.152939
R11747 gnd.n6723 gnd.n6722 0.152939
R11748 gnd.n6724 gnd.n6723 0.152939
R11749 gnd.n6724 gnd.n376 0.152939
R11750 gnd.n6732 gnd.n376 0.152939
R11751 gnd.n6733 gnd.n6732 0.152939
R11752 gnd.n6734 gnd.n6733 0.152939
R11753 gnd.n6734 gnd.n370 0.152939
R11754 gnd.n6742 gnd.n370 0.152939
R11755 gnd.n6743 gnd.n6742 0.152939
R11756 gnd.n6744 gnd.n6743 0.152939
R11757 gnd.n6744 gnd.n364 0.152939
R11758 gnd.n6752 gnd.n364 0.152939
R11759 gnd.n6753 gnd.n6752 0.152939
R11760 gnd.n6754 gnd.n6753 0.152939
R11761 gnd.n6754 gnd.n358 0.152939
R11762 gnd.n6762 gnd.n358 0.152939
R11763 gnd.n6763 gnd.n6762 0.152939
R11764 gnd.n6764 gnd.n6763 0.152939
R11765 gnd.n6764 gnd.n352 0.152939
R11766 gnd.n6772 gnd.n352 0.152939
R11767 gnd.n6773 gnd.n6772 0.152939
R11768 gnd.n6774 gnd.n6773 0.152939
R11769 gnd.n6774 gnd.n346 0.152939
R11770 gnd.n6782 gnd.n346 0.152939
R11771 gnd.n6783 gnd.n6782 0.152939
R11772 gnd.n6784 gnd.n6783 0.152939
R11773 gnd.n6784 gnd.n340 0.152939
R11774 gnd.n6792 gnd.n340 0.152939
R11775 gnd.n6793 gnd.n6792 0.152939
R11776 gnd.n6794 gnd.n6793 0.152939
R11777 gnd.n6794 gnd.n334 0.152939
R11778 gnd.n6802 gnd.n334 0.152939
R11779 gnd.n6803 gnd.n6802 0.152939
R11780 gnd.n6804 gnd.n6803 0.152939
R11781 gnd.n6804 gnd.n328 0.152939
R11782 gnd.n6812 gnd.n328 0.152939
R11783 gnd.n6813 gnd.n6812 0.152939
R11784 gnd.n6814 gnd.n6813 0.152939
R11785 gnd.n6814 gnd.n322 0.152939
R11786 gnd.n6822 gnd.n322 0.152939
R11787 gnd.n6823 gnd.n6822 0.152939
R11788 gnd.n6824 gnd.n6823 0.152939
R11789 gnd.n6824 gnd.n316 0.152939
R11790 gnd.n6832 gnd.n316 0.152939
R11791 gnd.n6833 gnd.n6832 0.152939
R11792 gnd.n6834 gnd.n6833 0.152939
R11793 gnd.n6834 gnd.n310 0.152939
R11794 gnd.n6842 gnd.n310 0.152939
R11795 gnd.n6843 gnd.n6842 0.152939
R11796 gnd.n6844 gnd.n6843 0.152939
R11797 gnd.n6844 gnd.n304 0.152939
R11798 gnd.n6852 gnd.n304 0.152939
R11799 gnd.n6853 gnd.n6852 0.152939
R11800 gnd.n6854 gnd.n6853 0.152939
R11801 gnd.n6854 gnd.n298 0.152939
R11802 gnd.n6862 gnd.n298 0.152939
R11803 gnd.n6863 gnd.n6862 0.152939
R11804 gnd.n6864 gnd.n6863 0.152939
R11805 gnd.n6864 gnd.n292 0.152939
R11806 gnd.n6872 gnd.n292 0.152939
R11807 gnd.n6873 gnd.n6872 0.152939
R11808 gnd.n6874 gnd.n6873 0.152939
R11809 gnd.n6874 gnd.n286 0.152939
R11810 gnd.n6882 gnd.n286 0.152939
R11811 gnd.n6883 gnd.n6882 0.152939
R11812 gnd.n6884 gnd.n6883 0.152939
R11813 gnd.n6885 gnd.n6884 0.152939
R11814 gnd.n6885 gnd.n280 0.152939
R11815 gnd.n6895 gnd.n280 0.152939
R11816 gnd.n5792 gnd.n5791 0.152939
R11817 gnd.n5794 gnd.n5792 0.152939
R11818 gnd.n5794 gnd.n5793 0.152939
R11819 gnd.n5793 gnd.n273 0.152939
R11820 gnd.n274 gnd.n273 0.152939
R11821 gnd.n275 gnd.n274 0.152939
R11822 gnd.n278 gnd.n275 0.152939
R11823 gnd.n279 gnd.n278 0.152939
R11824 gnd.n6896 gnd.n279 0.152939
R11825 gnd.n6944 gnd.n6943 0.152939
R11826 gnd.n6945 gnd.n6944 0.152939
R11827 gnd.n6945 gnd.n199 0.152939
R11828 gnd.n6959 gnd.n199 0.152939
R11829 gnd.n6960 gnd.n6959 0.152939
R11830 gnd.n6961 gnd.n6960 0.152939
R11831 gnd.n6961 gnd.n183 0.152939
R11832 gnd.n6975 gnd.n183 0.152939
R11833 gnd.n6976 gnd.n6975 0.152939
R11834 gnd.n6977 gnd.n6976 0.152939
R11835 gnd.n6977 gnd.n165 0.152939
R11836 gnd.n7065 gnd.n165 0.152939
R11837 gnd.n7066 gnd.n7065 0.152939
R11838 gnd.n7067 gnd.n7066 0.152939
R11839 gnd.n7067 gnd.n88 0.152939
R11840 gnd.n7147 gnd.n88 0.152939
R11841 gnd.n7146 gnd.n89 0.152939
R11842 gnd.n91 gnd.n89 0.152939
R11843 gnd.n95 gnd.n91 0.152939
R11844 gnd.n96 gnd.n95 0.152939
R11845 gnd.n97 gnd.n96 0.152939
R11846 gnd.n98 gnd.n97 0.152939
R11847 gnd.n102 gnd.n98 0.152939
R11848 gnd.n103 gnd.n102 0.152939
R11849 gnd.n104 gnd.n103 0.152939
R11850 gnd.n105 gnd.n104 0.152939
R11851 gnd.n109 gnd.n105 0.152939
R11852 gnd.n110 gnd.n109 0.152939
R11853 gnd.n111 gnd.n110 0.152939
R11854 gnd.n112 gnd.n111 0.152939
R11855 gnd.n116 gnd.n112 0.152939
R11856 gnd.n117 gnd.n116 0.152939
R11857 gnd.n118 gnd.n117 0.152939
R11858 gnd.n119 gnd.n118 0.152939
R11859 gnd.n123 gnd.n119 0.152939
R11860 gnd.n124 gnd.n123 0.152939
R11861 gnd.n125 gnd.n124 0.152939
R11862 gnd.n126 gnd.n125 0.152939
R11863 gnd.n130 gnd.n126 0.152939
R11864 gnd.n131 gnd.n130 0.152939
R11865 gnd.n132 gnd.n131 0.152939
R11866 gnd.n133 gnd.n132 0.152939
R11867 gnd.n137 gnd.n133 0.152939
R11868 gnd.n138 gnd.n137 0.152939
R11869 gnd.n139 gnd.n138 0.152939
R11870 gnd.n140 gnd.n139 0.152939
R11871 gnd.n144 gnd.n140 0.152939
R11872 gnd.n145 gnd.n144 0.152939
R11873 gnd.n146 gnd.n145 0.152939
R11874 gnd.n147 gnd.n146 0.152939
R11875 gnd.n151 gnd.n147 0.152939
R11876 gnd.n152 gnd.n151 0.152939
R11877 gnd.n7077 gnd.n152 0.152939
R11878 gnd.n7077 gnd.n7076 0.152939
R11879 gnd.n5609 gnd.n5608 0.152939
R11880 gnd.n5609 gnd.n1260 0.152939
R11881 gnd.n5624 gnd.n1260 0.152939
R11882 gnd.n5625 gnd.n5624 0.152939
R11883 gnd.n5626 gnd.n5625 0.152939
R11884 gnd.n5627 gnd.n5626 0.152939
R11885 gnd.n5628 gnd.n5627 0.152939
R11886 gnd.n5629 gnd.n5628 0.152939
R11887 gnd.n5630 gnd.n5629 0.152939
R11888 gnd.n5631 gnd.n5630 0.152939
R11889 gnd.n5632 gnd.n5631 0.152939
R11890 gnd.n5633 gnd.n5632 0.152939
R11891 gnd.n5634 gnd.n5633 0.152939
R11892 gnd.n5635 gnd.n5634 0.152939
R11893 gnd.n5636 gnd.n5635 0.152939
R11894 gnd.n5637 gnd.n5636 0.152939
R11895 gnd.n5638 gnd.n5637 0.152939
R11896 gnd.n5639 gnd.n5638 0.152939
R11897 gnd.n5640 gnd.n5639 0.152939
R11898 gnd.n5641 gnd.n5640 0.152939
R11899 gnd.n5643 gnd.n5641 0.152939
R11900 gnd.n5643 gnd.n5642 0.152939
R11901 gnd.n5642 gnd.n238 0.152939
R11902 gnd.n239 gnd.n238 0.152939
R11903 gnd.n240 gnd.n239 0.152939
R11904 gnd.n241 gnd.n240 0.152939
R11905 gnd.n242 gnd.n241 0.152939
R11906 gnd.n243 gnd.n242 0.152939
R11907 gnd.n244 gnd.n243 0.152939
R11908 gnd.n245 gnd.n244 0.152939
R11909 gnd.n246 gnd.n245 0.152939
R11910 gnd.n247 gnd.n246 0.152939
R11911 gnd.n248 gnd.n247 0.152939
R11912 gnd.n249 gnd.n248 0.152939
R11913 gnd.n250 gnd.n249 0.152939
R11914 gnd.n251 gnd.n250 0.152939
R11915 gnd.n252 gnd.n251 0.152939
R11916 gnd.n253 gnd.n252 0.152939
R11917 gnd.n255 gnd.n253 0.152939
R11918 gnd.n255 gnd.n254 0.152939
R11919 gnd.n254 gnd.n158 0.152939
R11920 gnd.n7075 gnd.n158 0.152939
R11921 gnd.n5513 gnd.n5512 0.152939
R11922 gnd.n5513 gnd.n5509 0.152939
R11923 gnd.n5521 gnd.n5509 0.152939
R11924 gnd.n5522 gnd.n5521 0.152939
R11925 gnd.n5523 gnd.n5522 0.152939
R11926 gnd.n5523 gnd.n5505 0.152939
R11927 gnd.n5531 gnd.n5505 0.152939
R11928 gnd.n5532 gnd.n5531 0.152939
R11929 gnd.n5533 gnd.n5532 0.152939
R11930 gnd.n5533 gnd.n5501 0.152939
R11931 gnd.n5541 gnd.n5501 0.152939
R11932 gnd.n5542 gnd.n5541 0.152939
R11933 gnd.n5544 gnd.n5542 0.152939
R11934 gnd.n5544 gnd.n5543 0.152939
R11935 gnd.n5543 gnd.n1290 0.152939
R11936 gnd.n5557 gnd.n5556 0.152939
R11937 gnd.n5557 gnd.n1286 0.152939
R11938 gnd.n5565 gnd.n1286 0.152939
R11939 gnd.n5566 gnd.n5565 0.152939
R11940 gnd.n5567 gnd.n5566 0.152939
R11941 gnd.n5567 gnd.n1282 0.152939
R11942 gnd.n5575 gnd.n1282 0.152939
R11943 gnd.n5576 gnd.n5575 0.152939
R11944 gnd.n5577 gnd.n5576 0.152939
R11945 gnd.n5577 gnd.n1278 0.152939
R11946 gnd.n5585 gnd.n1278 0.152939
R11947 gnd.n5586 gnd.n5585 0.152939
R11948 gnd.n5587 gnd.n5586 0.152939
R11949 gnd.n5587 gnd.n1274 0.152939
R11950 gnd.n5595 gnd.n1274 0.152939
R11951 gnd.n5596 gnd.n5595 0.152939
R11952 gnd.n5598 gnd.n5596 0.152939
R11953 gnd.n5598 gnd.n5597 0.152939
R11954 gnd.n5597 gnd.n1267 0.152939
R11955 gnd.n5607 gnd.n1267 0.152939
R11956 gnd.n1134 gnd.n1133 0.152939
R11957 gnd.n1135 gnd.n1134 0.152939
R11958 gnd.n1255 gnd.n1135 0.152939
R11959 gnd.n5691 gnd.n1255 0.152939
R11960 gnd.n5692 gnd.n5691 0.152939
R11961 gnd.n5693 gnd.n5692 0.152939
R11962 gnd.n5694 gnd.n5693 0.152939
R11963 gnd.n5694 gnd.n1227 0.152939
R11964 gnd.n5722 gnd.n1227 0.152939
R11965 gnd.n5723 gnd.n5722 0.152939
R11966 gnd.n5724 gnd.n5723 0.152939
R11967 gnd.n5726 gnd.n5724 0.152939
R11968 gnd.n5726 gnd.n5725 0.152939
R11969 gnd.n5725 gnd.n1199 0.152939
R11970 gnd.n1199 gnd.n214 0.152939
R11971 gnd.n6943 gnd.n214 0.152939
R11972 gnd.n4019 gnd.n4018 0.152939
R11973 gnd.n4020 gnd.n4019 0.152939
R11974 gnd.n4020 gnd.n2041 0.152939
R11975 gnd.n4082 gnd.n2041 0.152939
R11976 gnd.n4083 gnd.n4082 0.152939
R11977 gnd.n4084 gnd.n4083 0.152939
R11978 gnd.n4084 gnd.n2037 0.152939
R11979 gnd.n4090 gnd.n2037 0.152939
R11980 gnd.n4091 gnd.n4090 0.152939
R11981 gnd.n4092 gnd.n4091 0.152939
R11982 gnd.n4092 gnd.n2033 0.152939
R11983 gnd.n4098 gnd.n2033 0.152939
R11984 gnd.n4099 gnd.n4098 0.152939
R11985 gnd.n4100 gnd.n4099 0.152939
R11986 gnd.n4100 gnd.n2029 0.152939
R11987 gnd.n4106 gnd.n2029 0.152939
R11988 gnd.n4107 gnd.n4106 0.152939
R11989 gnd.n4108 gnd.n4107 0.152939
R11990 gnd.n4108 gnd.n2023 0.152939
R11991 gnd.n4248 gnd.n2023 0.152939
R11992 gnd.n4249 gnd.n4248 0.152939
R11993 gnd.n4250 gnd.n4249 0.152939
R11994 gnd.n4250 gnd.n1770 0.152939
R11995 gnd.n4417 gnd.n1770 0.152939
R11996 gnd.n4418 gnd.n4417 0.152939
R11997 gnd.n4419 gnd.n4418 0.152939
R11998 gnd.n4419 gnd.n1755 0.152939
R11999 gnd.n4462 gnd.n1755 0.152939
R12000 gnd.n4463 gnd.n4462 0.152939
R12001 gnd.n4464 gnd.n4463 0.152939
R12002 gnd.n4465 gnd.n4464 0.152939
R12003 gnd.n4465 gnd.n1727 0.152939
R12004 gnd.n4513 gnd.n1727 0.152939
R12005 gnd.n4514 gnd.n4513 0.152939
R12006 gnd.n4515 gnd.n4514 0.152939
R12007 gnd.n4515 gnd.n1707 0.152939
R12008 gnd.n4550 gnd.n1707 0.152939
R12009 gnd.n4551 gnd.n4550 0.152939
R12010 gnd.n4552 gnd.n4551 0.152939
R12011 gnd.n4552 gnd.n1681 0.152939
R12012 gnd.n4591 gnd.n1681 0.152939
R12013 gnd.n4592 gnd.n4591 0.152939
R12014 gnd.n4593 gnd.n4592 0.152939
R12015 gnd.n4593 gnd.n1665 0.152939
R12016 gnd.n4636 gnd.n1665 0.152939
R12017 gnd.n4637 gnd.n4636 0.152939
R12018 gnd.n4638 gnd.n4637 0.152939
R12019 gnd.n4639 gnd.n4638 0.152939
R12020 gnd.n4639 gnd.n1637 0.152939
R12021 gnd.n4708 gnd.n1637 0.152939
R12022 gnd.n4709 gnd.n4708 0.152939
R12023 gnd.n4710 gnd.n4709 0.152939
R12024 gnd.n4710 gnd.n1616 0.152939
R12025 gnd.n4735 gnd.n1616 0.152939
R12026 gnd.n4736 gnd.n4735 0.152939
R12027 gnd.n4737 gnd.n4736 0.152939
R12028 gnd.n4737 gnd.n1595 0.152939
R12029 gnd.n4768 gnd.n1595 0.152939
R12030 gnd.n4769 gnd.n4768 0.152939
R12031 gnd.n4770 gnd.n4769 0.152939
R12032 gnd.n4770 gnd.n1578 0.152939
R12033 gnd.n4813 gnd.n1578 0.152939
R12034 gnd.n4814 gnd.n4813 0.152939
R12035 gnd.n4815 gnd.n4814 0.152939
R12036 gnd.n4816 gnd.n4815 0.152939
R12037 gnd.n4816 gnd.n1549 0.152939
R12038 gnd.n4861 gnd.n1549 0.152939
R12039 gnd.n4862 gnd.n4861 0.152939
R12040 gnd.n4863 gnd.n4862 0.152939
R12041 gnd.n4863 gnd.n1529 0.152939
R12042 gnd.n4889 gnd.n1529 0.152939
R12043 gnd.n4890 gnd.n4889 0.152939
R12044 gnd.n4891 gnd.n4890 0.152939
R12045 gnd.n4892 gnd.n4891 0.152939
R12046 gnd.n4893 gnd.n4892 0.152939
R12047 gnd.n4893 gnd.n1497 0.152939
R12048 gnd.n4964 gnd.n1497 0.152939
R12049 gnd.n4965 gnd.n4964 0.152939
R12050 gnd.n4966 gnd.n4965 0.152939
R12051 gnd.n4967 gnd.n4966 0.152939
R12052 gnd.n4967 gnd.n1469 0.152939
R12053 gnd.n5015 gnd.n1469 0.152939
R12054 gnd.n5016 gnd.n5015 0.152939
R12055 gnd.n5017 gnd.n5016 0.152939
R12056 gnd.n5018 gnd.n5017 0.152939
R12057 gnd.n5018 gnd.n1451 0.152939
R12058 gnd.n5042 gnd.n1451 0.152939
R12059 gnd.n5043 gnd.n5042 0.152939
R12060 gnd.n5044 gnd.n5043 0.152939
R12061 gnd.n5044 gnd.n1394 0.152939
R12062 gnd.n5085 gnd.n1394 0.152939
R12063 gnd.n5086 gnd.n5085 0.152939
R12064 gnd.n5087 gnd.n5086 0.152939
R12065 gnd.n5087 gnd.n1373 0.152939
R12066 gnd.n5114 gnd.n1373 0.152939
R12067 gnd.n5115 gnd.n5114 0.152939
R12068 gnd.n5116 gnd.n5115 0.152939
R12069 gnd.n5118 gnd.n5116 0.152939
R12070 gnd.n5118 gnd.n5117 0.152939
R12071 gnd.n5117 gnd.n1344 0.152939
R12072 gnd.n1345 gnd.n1344 0.152939
R12073 gnd.n1346 gnd.n1345 0.152939
R12074 gnd.n1348 gnd.n1346 0.152939
R12075 gnd.n1348 gnd.n1347 0.152939
R12076 gnd.n1347 gnd.n1112 0.152939
R12077 gnd.n1113 gnd.n1112 0.152939
R12078 gnd.n1114 gnd.n1113 0.152939
R12079 gnd.n1120 gnd.n1114 0.152939
R12080 gnd.n1121 gnd.n1120 0.152939
R12081 gnd.n1122 gnd.n1121 0.152939
R12082 gnd.n1123 gnd.n1122 0.152939
R12083 gnd.n5674 gnd.n1123 0.152939
R12084 gnd.n5675 gnd.n5674 0.152939
R12085 gnd.n5680 gnd.n5675 0.152939
R12086 gnd.n5681 gnd.n5680 0.152939
R12087 gnd.n5682 gnd.n5681 0.152939
R12088 gnd.n5683 gnd.n5682 0.152939
R12089 gnd.n5683 gnd.n1237 0.152939
R12090 gnd.n5711 gnd.n1237 0.152939
R12091 gnd.n5712 gnd.n5711 0.152939
R12092 gnd.n5713 gnd.n5712 0.152939
R12093 gnd.n5714 gnd.n5713 0.152939
R12094 gnd.n5714 gnd.n1209 0.152939
R12095 gnd.n5743 gnd.n1209 0.152939
R12096 gnd.n5744 gnd.n5743 0.152939
R12097 gnd.n5745 gnd.n5744 0.152939
R12098 gnd.n5746 gnd.n5745 0.152939
R12099 gnd.n3695 gnd.n3689 0.152939
R12100 gnd.n3691 gnd.n3689 0.152939
R12101 gnd.n3691 gnd.n3690 0.152939
R12102 gnd.n3690 gnd.n2141 0.152939
R12103 gnd.n2141 gnd.n2139 0.152939
R12104 gnd.n3875 gnd.n2139 0.152939
R12105 gnd.n3876 gnd.n3875 0.152939
R12106 gnd.n3878 gnd.n3876 0.152939
R12107 gnd.n3878 gnd.n3877 0.152939
R12108 gnd.n3877 gnd.n2131 0.152939
R12109 gnd.n2132 gnd.n2131 0.152939
R12110 gnd.n2133 gnd.n2132 0.152939
R12111 gnd.n2133 gnd.n2121 0.152939
R12112 gnd.n3932 gnd.n2121 0.152939
R12113 gnd.n3933 gnd.n3932 0.152939
R12114 gnd.n3934 gnd.n3933 0.152939
R12115 gnd.n3935 gnd.n3934 0.152939
R12116 gnd.n3935 gnd.n2108 0.152939
R12117 gnd.n3979 gnd.n2108 0.152939
R12118 gnd.n3980 gnd.n3979 0.152939
R12119 gnd.n3845 gnd.n2158 0.152939
R12120 gnd.n3650 gnd.n2158 0.152939
R12121 gnd.n3650 gnd.n3649 0.152939
R12122 gnd.n3657 gnd.n3649 0.152939
R12123 gnd.n3658 gnd.n3657 0.152939
R12124 gnd.n3659 gnd.n3658 0.152939
R12125 gnd.n3659 gnd.n3647 0.152939
R12126 gnd.n3667 gnd.n3647 0.152939
R12127 gnd.n3668 gnd.n3667 0.152939
R12128 gnd.n3669 gnd.n3668 0.152939
R12129 gnd.n3669 gnd.n3645 0.152939
R12130 gnd.n3677 gnd.n3645 0.152939
R12131 gnd.n3678 gnd.n3677 0.152939
R12132 gnd.n3679 gnd.n3678 0.152939
R12133 gnd.n3679 gnd.n3643 0.152939
R12134 gnd.n3687 gnd.n3643 0.152939
R12135 gnd.n3688 gnd.n3687 0.152939
R12136 gnd.n3696 gnd.n3688 0.152939
R12137 gnd.n3856 gnd.n3846 0.152939
R12138 gnd.n3856 gnd.n3855 0.152939
R12139 gnd.n3855 gnd.n3854 0.152939
R12140 gnd.n3854 gnd.n3847 0.152939
R12141 gnd.n3849 gnd.n3847 0.152939
R12142 gnd.n3849 gnd.n3848 0.152939
R12143 gnd.n3848 gnd.n847 0.152939
R12144 gnd.n848 gnd.n847 0.152939
R12145 gnd.n849 gnd.n848 0.152939
R12146 gnd.n867 gnd.n849 0.152939
R12147 gnd.n868 gnd.n867 0.152939
R12148 gnd.n869 gnd.n868 0.152939
R12149 gnd.n870 gnd.n869 0.152939
R12150 gnd.n888 gnd.n870 0.152939
R12151 gnd.n889 gnd.n888 0.152939
R12152 gnd.n890 gnd.n889 0.152939
R12153 gnd.n891 gnd.n890 0.152939
R12154 gnd.n3968 gnd.n891 0.152939
R12155 gnd.n3969 gnd.n3968 0.152939
R12156 gnd.n3969 gnd.n2088 0.152939
R12157 gnd.n3988 gnd.n2088 0.152939
R12158 gnd.n3989 gnd.n3988 0.152939
R12159 gnd.n3990 gnd.n3989 0.152939
R12160 gnd.n3992 gnd.n3990 0.152939
R12161 gnd.n3992 gnd.n3991 0.152939
R12162 gnd.n3991 gnd.n916 0.152939
R12163 gnd.n917 gnd.n916 0.152939
R12164 gnd.n918 gnd.n917 0.152939
R12165 gnd.n934 gnd.n918 0.152939
R12166 gnd.n935 gnd.n934 0.152939
R12167 gnd.n936 gnd.n935 0.152939
R12168 gnd.n937 gnd.n936 0.152939
R12169 gnd.n956 gnd.n937 0.152939
R12170 gnd.n957 gnd.n956 0.152939
R12171 gnd.n958 gnd.n957 0.152939
R12172 gnd.n959 gnd.n958 0.152939
R12173 gnd.n977 gnd.n959 0.152939
R12174 gnd.n978 gnd.n977 0.152939
R12175 gnd.n979 gnd.n978 0.152939
R12176 gnd.n980 gnd.n979 0.152939
R12177 gnd.n998 gnd.n980 0.152939
R12178 gnd.n5995 gnd.n998 0.152939
R12179 gnd.n6049 gnd.n900 0.152939
R12180 gnd.n925 gnd.n900 0.152939
R12181 gnd.n926 gnd.n925 0.152939
R12182 gnd.n927 gnd.n926 0.152939
R12183 gnd.n945 gnd.n927 0.152939
R12184 gnd.n946 gnd.n945 0.152939
R12185 gnd.n947 gnd.n946 0.152939
R12186 gnd.n948 gnd.n947 0.152939
R12187 gnd.n966 gnd.n948 0.152939
R12188 gnd.n967 gnd.n966 0.152939
R12189 gnd.n968 gnd.n967 0.152939
R12190 gnd.n969 gnd.n968 0.152939
R12191 gnd.n988 gnd.n969 0.152939
R12192 gnd.n989 gnd.n988 0.152939
R12193 gnd.n990 gnd.n989 0.152939
R12194 gnd.n991 gnd.n990 0.152939
R12195 gnd.n1920 gnd.n1919 0.152939
R12196 gnd.n1921 gnd.n1920 0.152939
R12197 gnd.n1922 gnd.n1921 0.152939
R12198 gnd.n1923 gnd.n1922 0.152939
R12199 gnd.n1924 gnd.n1923 0.152939
R12200 gnd.n1925 gnd.n1924 0.152939
R12201 gnd.n1926 gnd.n1925 0.152939
R12202 gnd.n1927 gnd.n1926 0.152939
R12203 gnd.n1928 gnd.n1927 0.152939
R12204 gnd.n1929 gnd.n1928 0.152939
R12205 gnd.n1930 gnd.n1929 0.152939
R12206 gnd.n1931 gnd.n1930 0.152939
R12207 gnd.n1932 gnd.n1931 0.152939
R12208 gnd.n1933 gnd.n1932 0.152939
R12209 gnd.n1933 gnd.n1903 0.152939
R12210 gnd.n4342 gnd.n4341 0.152939
R12211 gnd.n4341 gnd.n1904 0.152939
R12212 gnd.n1964 gnd.n1904 0.152939
R12213 gnd.n1965 gnd.n1964 0.152939
R12214 gnd.n1966 gnd.n1965 0.152939
R12215 gnd.n1967 gnd.n1966 0.152939
R12216 gnd.n1971 gnd.n1967 0.152939
R12217 gnd.n1972 gnd.n1971 0.152939
R12218 gnd.n1973 gnd.n1972 0.152939
R12219 gnd.n1974 gnd.n1973 0.152939
R12220 gnd.n1978 gnd.n1974 0.152939
R12221 gnd.n1979 gnd.n1978 0.152939
R12222 gnd.n1980 gnd.n1979 0.152939
R12223 gnd.n1981 gnd.n1980 0.152939
R12224 gnd.n1985 gnd.n1981 0.152939
R12225 gnd.n1986 gnd.n1985 0.152939
R12226 gnd.n1987 gnd.n1986 0.152939
R12227 gnd.n1988 gnd.n1987 0.152939
R12228 gnd.n1993 gnd.n1988 0.152939
R12229 gnd.n4304 gnd.n1993 0.152939
R12230 gnd.n3759 gnd.n3744 0.152939
R12231 gnd.n3759 gnd.n3758 0.152939
R12232 gnd.n3758 gnd.n3757 0.152939
R12233 gnd.n3757 gnd.n3747 0.152939
R12234 gnd.n3748 gnd.n3747 0.152939
R12235 gnd.n3750 gnd.n3748 0.152939
R12236 gnd.n3750 gnd.n3749 0.152939
R12237 gnd.n3749 gnd.n2137 0.152939
R12238 gnd.n2137 gnd.n2135 0.152939
R12239 gnd.n3886 gnd.n2135 0.152939
R12240 gnd.n3887 gnd.n3886 0.152939
R12241 gnd.n3888 gnd.n3887 0.152939
R12242 gnd.n3889 gnd.n3888 0.152939
R12243 gnd.n3890 gnd.n3889 0.152939
R12244 gnd.n3890 gnd.n2118 0.152939
R12245 gnd.n3942 gnd.n2118 0.152939
R12246 gnd.n3943 gnd.n3942 0.152939
R12247 gnd.n3944 gnd.n3943 0.152939
R12248 gnd.n3945 gnd.n3944 0.152939
R12249 gnd.n3945 gnd.n2089 0.152939
R12250 gnd.n3987 gnd.n2089 0.152939
R12251 gnd.n3987 gnd.n2090 0.152939
R12252 gnd.n2092 gnd.n2090 0.152939
R12253 gnd.n2093 gnd.n2092 0.152939
R12254 gnd.n2094 gnd.n2093 0.152939
R12255 gnd.n2095 gnd.n2094 0.152939
R12256 gnd.n2096 gnd.n2095 0.152939
R12257 gnd.n2096 gnd.n2059 0.152939
R12258 gnd.n4036 gnd.n2059 0.152939
R12259 gnd.n4037 gnd.n4036 0.152939
R12260 gnd.n4038 gnd.n4037 0.152939
R12261 gnd.n4038 gnd.n2057 0.152939
R12262 gnd.n4044 gnd.n2057 0.152939
R12263 gnd.n4045 gnd.n4044 0.152939
R12264 gnd.n4046 gnd.n4045 0.152939
R12265 gnd.n4046 gnd.n2055 0.152939
R12266 gnd.n4055 gnd.n2055 0.152939
R12267 gnd.n4056 gnd.n4055 0.152939
R12268 gnd.n4058 gnd.n4056 0.152939
R12269 gnd.n4058 gnd.n4057 0.152939
R12270 gnd.n4057 gnd.n1994 0.152939
R12271 gnd.n4303 gnd.n1994 0.152939
R12272 gnd.n3702 gnd.n3701 0.152939
R12273 gnd.n3703 gnd.n3702 0.152939
R12274 gnd.n3704 gnd.n3703 0.152939
R12275 gnd.n3705 gnd.n3704 0.152939
R12276 gnd.n3706 gnd.n3705 0.152939
R12277 gnd.n3707 gnd.n3706 0.152939
R12278 gnd.n3708 gnd.n3707 0.152939
R12279 gnd.n3709 gnd.n3708 0.152939
R12280 gnd.n3710 gnd.n3709 0.152939
R12281 gnd.n3711 gnd.n3710 0.152939
R12282 gnd.n3712 gnd.n3711 0.152939
R12283 gnd.n3713 gnd.n3712 0.152939
R12284 gnd.n3714 gnd.n3713 0.152939
R12285 gnd.n3715 gnd.n3714 0.152939
R12286 gnd.n3716 gnd.n3715 0.152939
R12287 gnd.n3717 gnd.n3716 0.152939
R12288 gnd.n3718 gnd.n3717 0.152939
R12289 gnd.n3721 gnd.n3718 0.152939
R12290 gnd.n3722 gnd.n3721 0.152939
R12291 gnd.n3723 gnd.n3722 0.152939
R12292 gnd.n3724 gnd.n3723 0.152939
R12293 gnd.n3725 gnd.n3724 0.152939
R12294 gnd.n3726 gnd.n3725 0.152939
R12295 gnd.n3727 gnd.n3726 0.152939
R12296 gnd.n3728 gnd.n3727 0.152939
R12297 gnd.n3729 gnd.n3728 0.152939
R12298 gnd.n3730 gnd.n3729 0.152939
R12299 gnd.n3731 gnd.n3730 0.152939
R12300 gnd.n3732 gnd.n3731 0.152939
R12301 gnd.n3733 gnd.n3732 0.152939
R12302 gnd.n3734 gnd.n3733 0.152939
R12303 gnd.n3735 gnd.n3734 0.152939
R12304 gnd.n3736 gnd.n3735 0.152939
R12305 gnd.n3737 gnd.n3736 0.152939
R12306 gnd.n3738 gnd.n3737 0.152939
R12307 gnd.n3767 gnd.n3738 0.152939
R12308 gnd.n3767 gnd.n3766 0.152939
R12309 gnd.n3766 gnd.n3765 0.152939
R12310 gnd.n3862 gnd.n2148 0.152939
R12311 gnd.n3863 gnd.n3862 0.152939
R12312 gnd.n3865 gnd.n3863 0.152939
R12313 gnd.n3865 gnd.n3864 0.152939
R12314 gnd.n3864 gnd.n835 0.152939
R12315 gnd.n836 gnd.n835 0.152939
R12316 gnd.n837 gnd.n836 0.152939
R12317 gnd.n856 gnd.n837 0.152939
R12318 gnd.n857 gnd.n856 0.152939
R12319 gnd.n858 gnd.n857 0.152939
R12320 gnd.n859 gnd.n858 0.152939
R12321 gnd.n878 gnd.n859 0.152939
R12322 gnd.n879 gnd.n878 0.152939
R12323 gnd.n880 gnd.n879 0.152939
R12324 gnd.n881 gnd.n880 0.152939
R12325 gnd.n6049 gnd.n881 0.152939
R12326 gnd.n3906 gnd.n3905 0.152939
R12327 gnd.n3912 gnd.n3905 0.152939
R12328 gnd.n3913 gnd.n3912 0.152939
R12329 gnd.n3914 gnd.n3913 0.152939
R12330 gnd.n3914 gnd.n2127 0.152939
R12331 gnd.n3920 gnd.n2127 0.152939
R12332 gnd.n3921 gnd.n3920 0.152939
R12333 gnd.n3922 gnd.n3921 0.152939
R12334 gnd.n3923 gnd.n3922 0.152939
R12335 gnd.n6262 gnd.n658 0.152939
R12336 gnd.n663 gnd.n658 0.152939
R12337 gnd.n664 gnd.n663 0.152939
R12338 gnd.n665 gnd.n664 0.152939
R12339 gnd.n670 gnd.n665 0.152939
R12340 gnd.n671 gnd.n670 0.152939
R12341 gnd.n672 gnd.n671 0.152939
R12342 gnd.n673 gnd.n672 0.152939
R12343 gnd.n678 gnd.n673 0.152939
R12344 gnd.n679 gnd.n678 0.152939
R12345 gnd.n680 gnd.n679 0.152939
R12346 gnd.n681 gnd.n680 0.152939
R12347 gnd.n686 gnd.n681 0.152939
R12348 gnd.n687 gnd.n686 0.152939
R12349 gnd.n688 gnd.n687 0.152939
R12350 gnd.n689 gnd.n688 0.152939
R12351 gnd.n694 gnd.n689 0.152939
R12352 gnd.n695 gnd.n694 0.152939
R12353 gnd.n696 gnd.n695 0.152939
R12354 gnd.n697 gnd.n696 0.152939
R12355 gnd.n702 gnd.n697 0.152939
R12356 gnd.n703 gnd.n702 0.152939
R12357 gnd.n704 gnd.n703 0.152939
R12358 gnd.n705 gnd.n704 0.152939
R12359 gnd.n710 gnd.n705 0.152939
R12360 gnd.n711 gnd.n710 0.152939
R12361 gnd.n712 gnd.n711 0.152939
R12362 gnd.n713 gnd.n712 0.152939
R12363 gnd.n718 gnd.n713 0.152939
R12364 gnd.n719 gnd.n718 0.152939
R12365 gnd.n720 gnd.n719 0.152939
R12366 gnd.n721 gnd.n720 0.152939
R12367 gnd.n726 gnd.n721 0.152939
R12368 gnd.n727 gnd.n726 0.152939
R12369 gnd.n728 gnd.n727 0.152939
R12370 gnd.n729 gnd.n728 0.152939
R12371 gnd.n734 gnd.n729 0.152939
R12372 gnd.n735 gnd.n734 0.152939
R12373 gnd.n736 gnd.n735 0.152939
R12374 gnd.n737 gnd.n736 0.152939
R12375 gnd.n742 gnd.n737 0.152939
R12376 gnd.n743 gnd.n742 0.152939
R12377 gnd.n744 gnd.n743 0.152939
R12378 gnd.n745 gnd.n744 0.152939
R12379 gnd.n750 gnd.n745 0.152939
R12380 gnd.n751 gnd.n750 0.152939
R12381 gnd.n752 gnd.n751 0.152939
R12382 gnd.n753 gnd.n752 0.152939
R12383 gnd.n758 gnd.n753 0.152939
R12384 gnd.n759 gnd.n758 0.152939
R12385 gnd.n760 gnd.n759 0.152939
R12386 gnd.n761 gnd.n760 0.152939
R12387 gnd.n766 gnd.n761 0.152939
R12388 gnd.n767 gnd.n766 0.152939
R12389 gnd.n768 gnd.n767 0.152939
R12390 gnd.n769 gnd.n768 0.152939
R12391 gnd.n774 gnd.n769 0.152939
R12392 gnd.n775 gnd.n774 0.152939
R12393 gnd.n776 gnd.n775 0.152939
R12394 gnd.n777 gnd.n776 0.152939
R12395 gnd.n782 gnd.n777 0.152939
R12396 gnd.n783 gnd.n782 0.152939
R12397 gnd.n784 gnd.n783 0.152939
R12398 gnd.n785 gnd.n784 0.152939
R12399 gnd.n790 gnd.n785 0.152939
R12400 gnd.n791 gnd.n790 0.152939
R12401 gnd.n792 gnd.n791 0.152939
R12402 gnd.n793 gnd.n792 0.152939
R12403 gnd.n798 gnd.n793 0.152939
R12404 gnd.n799 gnd.n798 0.152939
R12405 gnd.n800 gnd.n799 0.152939
R12406 gnd.n801 gnd.n800 0.152939
R12407 gnd.n806 gnd.n801 0.152939
R12408 gnd.n807 gnd.n806 0.152939
R12409 gnd.n808 gnd.n807 0.152939
R12410 gnd.n809 gnd.n808 0.152939
R12411 gnd.n814 gnd.n809 0.152939
R12412 gnd.n815 gnd.n814 0.152939
R12413 gnd.n816 gnd.n815 0.152939
R12414 gnd.n817 gnd.n816 0.152939
R12415 gnd.n822 gnd.n817 0.152939
R12416 gnd.n823 gnd.n822 0.152939
R12417 gnd.n824 gnd.n823 0.152939
R12418 gnd.n825 gnd.n824 0.152939
R12419 gnd.n5300 gnd.n5156 0.152939
R12420 gnd.n5301 gnd.n5300 0.152939
R12421 gnd.n5302 gnd.n5301 0.152939
R12422 gnd.n5302 gnd.n5152 0.152939
R12423 gnd.n5313 gnd.n5152 0.152939
R12424 gnd.n5314 gnd.n5313 0.152939
R12425 gnd.n5315 gnd.n5314 0.152939
R12426 gnd.n5315 gnd.n5148 0.152939
R12427 gnd.n5322 gnd.n5148 0.152939
R12428 gnd.n4276 gnd.n2018 0.152939
R12429 gnd.n4272 gnd.n2018 0.152939
R12430 gnd.n4272 gnd.n4271 0.152939
R12431 gnd.n4271 gnd.n4270 0.152939
R12432 gnd.n4270 gnd.n4259 0.152939
R12433 gnd.n4266 gnd.n4259 0.152939
R12434 gnd.n4266 gnd.n1742 0.152939
R12435 gnd.n4481 gnd.n1742 0.152939
R12436 gnd.n4482 gnd.n4481 0.152939
R12437 gnd.n4497 gnd.n4482 0.152939
R12438 gnd.n4497 gnd.n4496 0.152939
R12439 gnd.n4496 gnd.n4495 0.152939
R12440 gnd.n4495 gnd.n4483 0.152939
R12441 gnd.n4491 gnd.n4483 0.152939
R12442 gnd.n4491 gnd.n4490 0.152939
R12443 gnd.n4490 gnd.n4489 0.152939
R12444 gnd.n4489 gnd.n1695 0.152939
R12445 gnd.n4568 gnd.n1695 0.152939
R12446 gnd.n4569 gnd.n4568 0.152939
R12447 gnd.n4577 gnd.n4569 0.152939
R12448 gnd.n4577 gnd.n4576 0.152939
R12449 gnd.n4576 gnd.n4575 0.152939
R12450 gnd.n4575 gnd.n4570 0.152939
R12451 gnd.n4570 gnd.n1652 0.152939
R12452 gnd.n4654 gnd.n1652 0.152939
R12453 gnd.n4655 gnd.n4654 0.152939
R12454 gnd.n4692 gnd.n4655 0.152939
R12455 gnd.n4692 gnd.n4691 0.152939
R12456 gnd.n4691 gnd.n4690 0.152939
R12457 gnd.n4690 gnd.n4656 0.152939
R12458 gnd.n4686 gnd.n4656 0.152939
R12459 gnd.n4686 gnd.n4685 0.152939
R12460 gnd.n4685 gnd.n4684 0.152939
R12461 gnd.n4684 gnd.n4661 0.152939
R12462 gnd.n4680 gnd.n4661 0.152939
R12463 gnd.n4680 gnd.n4679 0.152939
R12464 gnd.n4679 gnd.n4678 0.152939
R12465 gnd.n4678 gnd.n4666 0.152939
R12466 gnd.n4674 gnd.n4666 0.152939
R12467 gnd.n4674 gnd.n4673 0.152939
R12468 gnd.n4673 gnd.n1564 0.152939
R12469 gnd.n4831 gnd.n1564 0.152939
R12470 gnd.n4832 gnd.n4831 0.152939
R12471 gnd.n4846 gnd.n4832 0.152939
R12472 gnd.n4846 gnd.n4845 0.152939
R12473 gnd.n4845 gnd.n4844 0.152939
R12474 gnd.n4844 gnd.n4833 0.152939
R12475 gnd.n4840 gnd.n4833 0.152939
R12476 gnd.n4840 gnd.n4839 0.152939
R12477 gnd.n4839 gnd.n1514 0.152939
R12478 gnd.n4916 gnd.n1514 0.152939
R12479 gnd.n4917 gnd.n4916 0.152939
R12480 gnd.n4922 gnd.n4917 0.152939
R12481 gnd.n4922 gnd.n4921 0.152939
R12482 gnd.n4921 gnd.n4920 0.152939
R12483 gnd.n4920 gnd.n1484 0.152939
R12484 gnd.n4983 gnd.n1484 0.152939
R12485 gnd.n4984 gnd.n4983 0.152939
R12486 gnd.n4999 gnd.n4984 0.152939
R12487 gnd.n4999 gnd.n4998 0.152939
R12488 gnd.n4998 gnd.n4997 0.152939
R12489 gnd.n4997 gnd.n4985 0.152939
R12490 gnd.n4993 gnd.n4985 0.152939
R12491 gnd.n4993 gnd.n4992 0.152939
R12492 gnd.n4992 gnd.n1409 0.152939
R12493 gnd.n5068 gnd.n1409 0.152939
R12494 gnd.n5069 gnd.n5068 0.152939
R12495 gnd.n5071 gnd.n5069 0.152939
R12496 gnd.n5071 gnd.n5070 0.152939
R12497 gnd.n5070 gnd.n1380 0.152939
R12498 gnd.n5104 gnd.n1380 0.152939
R12499 gnd.n5105 gnd.n5104 0.152939
R12500 gnd.n5106 gnd.n5105 0.152939
R12501 gnd.n5106 gnd.n1358 0.152939
R12502 gnd.n5135 gnd.n1358 0.152939
R12503 gnd.n5136 gnd.n5135 0.152939
R12504 gnd.n5137 gnd.n5136 0.152939
R12505 gnd.n5137 gnd.n1354 0.152939
R12506 gnd.n5146 gnd.n1354 0.152939
R12507 gnd.n5147 gnd.n5146 0.152939
R12508 gnd.n5324 gnd.n5147 0.152939
R12509 gnd.n5324 gnd.n5323 0.152939
R12510 gnd.n4289 gnd.n1999 0.152939
R12511 gnd.n4289 gnd.n4288 0.152939
R12512 gnd.n4288 gnd.n4287 0.152939
R12513 gnd.n4287 gnd.n2006 0.152939
R12514 gnd.n4283 gnd.n2006 0.152939
R12515 gnd.n4283 gnd.n4282 0.152939
R12516 gnd.n4282 gnd.n2013 0.152939
R12517 gnd.n4278 gnd.n2013 0.152939
R12518 gnd.n4278 gnd.n4277 0.152939
R12519 gnd.n4007 gnd.n2074 0.152939
R12520 gnd.n4008 gnd.n4007 0.152939
R12521 gnd.n4009 gnd.n4008 0.152939
R12522 gnd.n4009 gnd.n2062 0.152939
R12523 gnd.n4028 gnd.n2062 0.152939
R12524 gnd.n4029 gnd.n4028 0.152939
R12525 gnd.n4030 gnd.n4029 0.152939
R12526 gnd.n4030 gnd.n2047 0.152939
R12527 gnd.n4075 gnd.n2047 0.152939
R12528 gnd.n4075 gnd.n4074 0.152939
R12529 gnd.n4074 gnd.n4073 0.152939
R12530 gnd.n4073 gnd.n2048 0.152939
R12531 gnd.n4069 gnd.n2048 0.152939
R12532 gnd.n4069 gnd.n4068 0.152939
R12533 gnd.n4068 gnd.n4067 0.152939
R12534 gnd.n4067 gnd.n2052 0.152939
R12535 gnd.n4063 gnd.n2052 0.152939
R12536 gnd.n4063 gnd.n1998 0.152939
R12537 gnd.n4296 gnd.n1998 0.152939
R12538 gnd.n4296 gnd.n4295 0.152939
R12539 gnd.n5992 gnd.n1001 0.152939
R12540 gnd.n5988 gnd.n1001 0.152939
R12541 gnd.n5988 gnd.n5987 0.152939
R12542 gnd.n5987 gnd.n5986 0.152939
R12543 gnd.n5986 gnd.n1006 0.152939
R12544 gnd.n5982 gnd.n1006 0.152939
R12545 gnd.n5982 gnd.n5981 0.152939
R12546 gnd.n5981 gnd.n5980 0.152939
R12547 gnd.n5980 gnd.n1011 0.152939
R12548 gnd.n5976 gnd.n1011 0.152939
R12549 gnd.n5976 gnd.n5975 0.152939
R12550 gnd.n5975 gnd.n5974 0.152939
R12551 gnd.n5974 gnd.n1016 0.152939
R12552 gnd.n5970 gnd.n1016 0.152939
R12553 gnd.n5970 gnd.n5969 0.152939
R12554 gnd.n5969 gnd.n5968 0.152939
R12555 gnd.n5968 gnd.n1021 0.152939
R12556 gnd.n5964 gnd.n1021 0.152939
R12557 gnd.n5964 gnd.n5963 0.152939
R12558 gnd.n5963 gnd.n5962 0.152939
R12559 gnd.n5962 gnd.n1026 0.152939
R12560 gnd.n5958 gnd.n1026 0.152939
R12561 gnd.n5958 gnd.n5957 0.152939
R12562 gnd.n5957 gnd.n5956 0.152939
R12563 gnd.n5956 gnd.n1031 0.152939
R12564 gnd.n5952 gnd.n1031 0.152939
R12565 gnd.n5952 gnd.n5951 0.152939
R12566 gnd.n5951 gnd.n5950 0.152939
R12567 gnd.n5950 gnd.n1036 0.152939
R12568 gnd.n5946 gnd.n1036 0.152939
R12569 gnd.n5946 gnd.n5945 0.152939
R12570 gnd.n5945 gnd.n5944 0.152939
R12571 gnd.n5944 gnd.n1041 0.152939
R12572 gnd.n5940 gnd.n1041 0.152939
R12573 gnd.n5940 gnd.n5939 0.152939
R12574 gnd.n5939 gnd.n5938 0.152939
R12575 gnd.n5938 gnd.n1046 0.152939
R12576 gnd.n5934 gnd.n1046 0.152939
R12577 gnd.n5934 gnd.n5933 0.152939
R12578 gnd.n5933 gnd.n5932 0.152939
R12579 gnd.n5932 gnd.n1051 0.152939
R12580 gnd.n5928 gnd.n1051 0.152939
R12581 gnd.n5928 gnd.n5927 0.152939
R12582 gnd.n5927 gnd.n5926 0.152939
R12583 gnd.n5926 gnd.n1056 0.152939
R12584 gnd.n5922 gnd.n1056 0.152939
R12585 gnd.n5922 gnd.n5921 0.152939
R12586 gnd.n5921 gnd.n5920 0.152939
R12587 gnd.n5920 gnd.n1061 0.152939
R12588 gnd.n5916 gnd.n1061 0.152939
R12589 gnd.n5916 gnd.n5915 0.152939
R12590 gnd.n5915 gnd.n5914 0.152939
R12591 gnd.n5914 gnd.n1066 0.152939
R12592 gnd.n5910 gnd.n1066 0.152939
R12593 gnd.n5910 gnd.n5909 0.152939
R12594 gnd.n5909 gnd.n5908 0.152939
R12595 gnd.n5908 gnd.n1071 0.152939
R12596 gnd.n5904 gnd.n1071 0.152939
R12597 gnd.n5904 gnd.n5903 0.152939
R12598 gnd.n5903 gnd.n5902 0.152939
R12599 gnd.n5902 gnd.n1076 0.152939
R12600 gnd.n5898 gnd.n1076 0.152939
R12601 gnd.n5898 gnd.n5897 0.152939
R12602 gnd.n5897 gnd.n5896 0.152939
R12603 gnd.n5896 gnd.n1081 0.152939
R12604 gnd.n5892 gnd.n1081 0.152939
R12605 gnd.n5892 gnd.n5891 0.152939
R12606 gnd.n5891 gnd.n5890 0.152939
R12607 gnd.n5890 gnd.n1086 0.152939
R12608 gnd.n5886 gnd.n1086 0.152939
R12609 gnd.n5886 gnd.n5885 0.152939
R12610 gnd.n5885 gnd.n5884 0.152939
R12611 gnd.n5884 gnd.n1091 0.152939
R12612 gnd.n5880 gnd.n1091 0.152939
R12613 gnd.n5880 gnd.n5879 0.152939
R12614 gnd.n5879 gnd.n5878 0.152939
R12615 gnd.n5878 gnd.n1096 0.152939
R12616 gnd.n5874 gnd.n1096 0.152939
R12617 gnd.n5874 gnd.n5873 0.152939
R12618 gnd.n5873 gnd.n5872 0.152939
R12619 gnd.n5872 gnd.n1101 0.152939
R12620 gnd.n1104 gnd.n1101 0.152939
R12621 gnd.n5203 gnd.n1146 0.152939
R12622 gnd.n5842 gnd.n1146 0.152939
R12623 gnd.n5842 gnd.n5841 0.152939
R12624 gnd.n5841 gnd.n5840 0.152939
R12625 gnd.n5840 gnd.n1147 0.152939
R12626 gnd.n5836 gnd.n1147 0.152939
R12627 gnd.n5836 gnd.n5835 0.152939
R12628 gnd.n5835 gnd.n5834 0.152939
R12629 gnd.n5834 gnd.n1152 0.152939
R12630 gnd.n5830 gnd.n1152 0.152939
R12631 gnd.n5830 gnd.n5829 0.152939
R12632 gnd.n5829 gnd.n5828 0.152939
R12633 gnd.n5828 gnd.n1157 0.152939
R12634 gnd.n5824 gnd.n1157 0.152939
R12635 gnd.n5824 gnd.n5823 0.152939
R12636 gnd.n5823 gnd.n5822 0.152939
R12637 gnd.n5822 gnd.n1162 0.152939
R12638 gnd.n5818 gnd.n1162 0.152939
R12639 gnd.n5818 gnd.n5817 0.152939
R12640 gnd.n5817 gnd.n5816 0.152939
R12641 gnd.n5816 gnd.n1167 0.152939
R12642 gnd.n5812 gnd.n1167 0.152939
R12643 gnd.n5812 gnd.n228 0.152939
R12644 gnd.n6935 gnd.n228 0.152939
R12645 gnd.n6936 gnd.n6935 0.152939
R12646 gnd.n6937 gnd.n6936 0.152939
R12647 gnd.n6937 gnd.n206 0.152939
R12648 gnd.n6951 gnd.n206 0.152939
R12649 gnd.n6952 gnd.n6951 0.152939
R12650 gnd.n6953 gnd.n6952 0.152939
R12651 gnd.n6953 gnd.n191 0.152939
R12652 gnd.n6967 gnd.n191 0.152939
R12653 gnd.n6968 gnd.n6967 0.152939
R12654 gnd.n6969 gnd.n6968 0.152939
R12655 gnd.n6969 gnd.n174 0.152939
R12656 gnd.n6983 gnd.n174 0.152939
R12657 gnd.n6984 gnd.n6983 0.152939
R12658 gnd.n7059 gnd.n6984 0.152939
R12659 gnd.n7059 gnd.n7058 0.152939
R12660 gnd.n7058 gnd.n7057 0.152939
R12661 gnd.n7057 gnd.n6985 0.152939
R12662 gnd.n7053 gnd.n6985 0.152939
R12663 gnd.n7052 gnd.n6987 0.152939
R12664 gnd.n7048 gnd.n6987 0.152939
R12665 gnd.n7048 gnd.n7047 0.152939
R12666 gnd.n7047 gnd.n7046 0.152939
R12667 gnd.n7046 gnd.n6993 0.152939
R12668 gnd.n7042 gnd.n6993 0.152939
R12669 gnd.n7042 gnd.n7041 0.152939
R12670 gnd.n7041 gnd.n7040 0.152939
R12671 gnd.n7040 gnd.n7001 0.152939
R12672 gnd.n7036 gnd.n7001 0.152939
R12673 gnd.n7036 gnd.n7035 0.152939
R12674 gnd.n7035 gnd.n7034 0.152939
R12675 gnd.n7034 gnd.n7009 0.152939
R12676 gnd.n7030 gnd.n7009 0.152939
R12677 gnd.n7030 gnd.n7029 0.152939
R12678 gnd.n7029 gnd.n7028 0.152939
R12679 gnd.n7028 gnd.n7017 0.152939
R12680 gnd.n7017 gnd.n78 0.152939
R12681 gnd.n5615 gnd.n1264 0.152939
R12682 gnd.n5616 gnd.n5615 0.152939
R12683 gnd.n5618 gnd.n5616 0.152939
R12684 gnd.n5618 gnd.n5617 0.152939
R12685 gnd.n5617 gnd.n1246 0.152939
R12686 gnd.n5701 gnd.n1246 0.152939
R12687 gnd.n5702 gnd.n5701 0.152939
R12688 gnd.n5704 gnd.n5702 0.152939
R12689 gnd.n5704 gnd.n5703 0.152939
R12690 gnd.n5703 gnd.n1217 0.152939
R12691 gnd.n5733 gnd.n1217 0.152939
R12692 gnd.n5734 gnd.n5733 0.152939
R12693 gnd.n5736 gnd.n5734 0.152939
R12694 gnd.n5736 gnd.n5735 0.152939
R12695 gnd.n5735 gnd.n1191 0.152939
R12696 gnd.n5766 gnd.n1191 0.152939
R12697 gnd.n5767 gnd.n5766 0.152939
R12698 gnd.n5769 gnd.n5767 0.152939
R12699 gnd.n5769 gnd.n5768 0.152939
R12700 gnd.n5768 gnd.n51 0.152939
R12701 gnd.n7184 gnd.n51 0.152939
R12702 gnd.n7184 gnd.n7183 0.152939
R12703 gnd.n7183 gnd.n53 0.152939
R12704 gnd.n7179 gnd.n53 0.152939
R12705 gnd.n7179 gnd.n7178 0.152939
R12706 gnd.n7178 gnd.n7177 0.152939
R12707 gnd.n7177 gnd.n58 0.152939
R12708 gnd.n7173 gnd.n58 0.152939
R12709 gnd.n7173 gnd.n7172 0.152939
R12710 gnd.n7172 gnd.n7171 0.152939
R12711 gnd.n7171 gnd.n63 0.152939
R12712 gnd.n7167 gnd.n63 0.152939
R12713 gnd.n7167 gnd.n7166 0.152939
R12714 gnd.n7166 gnd.n7165 0.152939
R12715 gnd.n7165 gnd.n68 0.152939
R12716 gnd.n7161 gnd.n68 0.152939
R12717 gnd.n7161 gnd.n7160 0.152939
R12718 gnd.n7160 gnd.n7159 0.152939
R12719 gnd.n7159 gnd.n73 0.152939
R12720 gnd.n7155 gnd.n73 0.152939
R12721 gnd.n7155 gnd.n7154 0.152939
R12722 gnd.n7154 gnd.n7153 0.152939
R12723 gnd.n5291 gnd.n5156 0.151415
R12724 gnd.n4294 gnd.n1999 0.151415
R12725 gnd.n3981 gnd.n3980 0.145814
R12726 gnd.n3981 gnd.n2074 0.145814
R12727 gnd.n2428 gnd.n0 0.127478
R12728 gnd.n5791 gnd.n215 0.10111
R12729 gnd.n3923 gnd.n901 0.10111
R12730 gnd.n3008 gnd.n3007 0.0767195
R12731 gnd.n3007 gnd.n3006 0.0767195
R12732 gnd.n5994 gnd.n5993 0.063
R12733 gnd.n5204 gnd.n5201 0.063
R12734 gnd.n4018 gnd.n901 0.0523293
R12735 gnd.n5746 gnd.n215 0.0523293
R12736 gnd.n3575 gnd.n2202 0.0477147
R12737 gnd.n2771 gnd.n2659 0.0442063
R12738 gnd.n2772 gnd.n2771 0.0442063
R12739 gnd.n2773 gnd.n2772 0.0442063
R12740 gnd.n2773 gnd.n2648 0.0442063
R12741 gnd.n2787 gnd.n2648 0.0442063
R12742 gnd.n2788 gnd.n2787 0.0442063
R12743 gnd.n2789 gnd.n2788 0.0442063
R12744 gnd.n2789 gnd.n2635 0.0442063
R12745 gnd.n2833 gnd.n2635 0.0442063
R12746 gnd.n2834 gnd.n2833 0.0442063
R12747 gnd.n2836 gnd.n2569 0.0344674
R12748 gnd.n5292 gnd.n5290 0.0344674
R12749 gnd.n4293 gnd.n2000 0.0344674
R12750 gnd.n2856 gnd.n2855 0.0269946
R12751 gnd.n2858 gnd.n2857 0.0269946
R12752 gnd.n2564 gnd.n2562 0.0269946
R12753 gnd.n2868 gnd.n2866 0.0269946
R12754 gnd.n2867 gnd.n2543 0.0269946
R12755 gnd.n2887 gnd.n2886 0.0269946
R12756 gnd.n2889 gnd.n2888 0.0269946
R12757 gnd.n2538 gnd.n2537 0.0269946
R12758 gnd.n2899 gnd.n2533 0.0269946
R12759 gnd.n2898 gnd.n2535 0.0269946
R12760 gnd.n2534 gnd.n2516 0.0269946
R12761 gnd.n2919 gnd.n2517 0.0269946
R12762 gnd.n2918 gnd.n2518 0.0269946
R12763 gnd.n2952 gnd.n2493 0.0269946
R12764 gnd.n2954 gnd.n2953 0.0269946
R12765 gnd.n2955 gnd.n2440 0.0269946
R12766 gnd.n2488 gnd.n2441 0.0269946
R12767 gnd.n2490 gnd.n2442 0.0269946
R12768 gnd.n2965 gnd.n2964 0.0269946
R12769 gnd.n2967 gnd.n2966 0.0269946
R12770 gnd.n2968 gnd.n2462 0.0269946
R12771 gnd.n2970 gnd.n2463 0.0269946
R12772 gnd.n2973 gnd.n2464 0.0269946
R12773 gnd.n2976 gnd.n2975 0.0269946
R12774 gnd.n2978 gnd.n2977 0.0269946
R12775 gnd.n3043 gnd.n2375 0.0269946
R12776 gnd.n3045 gnd.n3044 0.0269946
R12777 gnd.n3054 gnd.n2368 0.0269946
R12778 gnd.n3056 gnd.n3055 0.0269946
R12779 gnd.n3057 gnd.n2366 0.0269946
R12780 gnd.n3064 gnd.n3060 0.0269946
R12781 gnd.n3063 gnd.n3062 0.0269946
R12782 gnd.n3061 gnd.n2345 0.0269946
R12783 gnd.n3086 gnd.n2346 0.0269946
R12784 gnd.n3085 gnd.n2347 0.0269946
R12785 gnd.n3128 gnd.n2320 0.0269946
R12786 gnd.n3130 gnd.n3129 0.0269946
R12787 gnd.n3140 gnd.n2313 0.0269946
R12788 gnd.n3142 gnd.n3141 0.0269946
R12789 gnd.n3143 gnd.n2311 0.0269946
R12790 gnd.n3150 gnd.n3146 0.0269946
R12791 gnd.n3149 gnd.n3148 0.0269946
R12792 gnd.n3147 gnd.n2290 0.0269946
R12793 gnd.n3172 gnd.n2291 0.0269946
R12794 gnd.n3171 gnd.n2292 0.0269946
R12795 gnd.n3218 gnd.n2266 0.0269946
R12796 gnd.n3220 gnd.n3219 0.0269946
R12797 gnd.n3229 gnd.n2259 0.0269946
R12798 gnd.n3488 gnd.n2257 0.0269946
R12799 gnd.n3493 gnd.n3491 0.0269946
R12800 gnd.n3492 gnd.n2238 0.0269946
R12801 gnd.n3517 gnd.n3516 0.0269946
R12802 gnd.n5201 gnd.n5200 0.0246168
R12803 gnd.n5993 gnd.n1000 0.0246168
R12804 gnd.n2836 gnd.n2835 0.0202011
R12805 gnd.n5200 gnd.n5198 0.0174837
R12806 gnd.n5212 gnd.n5198 0.0174837
R12807 gnd.n5214 gnd.n5212 0.0174837
R12808 gnd.n5214 gnd.n5213 0.0174837
R12809 gnd.n5213 gnd.n5193 0.0174837
R12810 gnd.n5223 gnd.n5193 0.0174837
R12811 gnd.n5223 gnd.n5222 0.0174837
R12812 gnd.n5222 gnd.n5194 0.0174837
R12813 gnd.n5194 gnd.n5189 0.0174837
R12814 gnd.n5231 gnd.n5189 0.0174837
R12815 gnd.n5233 gnd.n5231 0.0174837
R12816 gnd.n5233 gnd.n5232 0.0174837
R12817 gnd.n5232 gnd.n5184 0.0174837
R12818 gnd.n5242 gnd.n5184 0.0174837
R12819 gnd.n5242 gnd.n5241 0.0174837
R12820 gnd.n5241 gnd.n5185 0.0174837
R12821 gnd.n5185 gnd.n5180 0.0174837
R12822 gnd.n5250 gnd.n5180 0.0174837
R12823 gnd.n5252 gnd.n5250 0.0174837
R12824 gnd.n5252 gnd.n5251 0.0174837
R12825 gnd.n5251 gnd.n5175 0.0174837
R12826 gnd.n5261 gnd.n5175 0.0174837
R12827 gnd.n5261 gnd.n5260 0.0174837
R12828 gnd.n5260 gnd.n5176 0.0174837
R12829 gnd.n5176 gnd.n5171 0.0174837
R12830 gnd.n5269 gnd.n5171 0.0174837
R12831 gnd.n5271 gnd.n5269 0.0174837
R12832 gnd.n5271 gnd.n5270 0.0174837
R12833 gnd.n5270 gnd.n5166 0.0174837
R12834 gnd.n5282 gnd.n5166 0.0174837
R12835 gnd.n5282 gnd.n5281 0.0174837
R12836 gnd.n5281 gnd.n5167 0.0174837
R12837 gnd.n5167 gnd.n5160 0.0174837
R12838 gnd.n5289 gnd.n5160 0.0174837
R12839 gnd.n5290 gnd.n5289 0.0174837
R12840 gnd.n4129 gnd.n1000 0.0174837
R12841 gnd.n4131 gnd.n4129 0.0174837
R12842 gnd.n4239 gnd.n4131 0.0174837
R12843 gnd.n4239 gnd.n4238 0.0174837
R12844 gnd.n4238 gnd.n4132 0.0174837
R12845 gnd.n4235 gnd.n4132 0.0174837
R12846 gnd.n4235 gnd.n4234 0.0174837
R12847 gnd.n4234 gnd.n4142 0.0174837
R12848 gnd.n4231 gnd.n4142 0.0174837
R12849 gnd.n4231 gnd.n4230 0.0174837
R12850 gnd.n4230 gnd.n4147 0.0174837
R12851 gnd.n4227 gnd.n4147 0.0174837
R12852 gnd.n4227 gnd.n4226 0.0174837
R12853 gnd.n4226 gnd.n4153 0.0174837
R12854 gnd.n4223 gnd.n4153 0.0174837
R12855 gnd.n4223 gnd.n4222 0.0174837
R12856 gnd.n4222 gnd.n4157 0.0174837
R12857 gnd.n4219 gnd.n4157 0.0174837
R12858 gnd.n4219 gnd.n4218 0.0174837
R12859 gnd.n4218 gnd.n4164 0.0174837
R12860 gnd.n4215 gnd.n4164 0.0174837
R12861 gnd.n4215 gnd.n4214 0.0174837
R12862 gnd.n4214 gnd.n4170 0.0174837
R12863 gnd.n4211 gnd.n4170 0.0174837
R12864 gnd.n4211 gnd.n4210 0.0174837
R12865 gnd.n4210 gnd.n4176 0.0174837
R12866 gnd.n4207 gnd.n4176 0.0174837
R12867 gnd.n4207 gnd.n4206 0.0174837
R12868 gnd.n4206 gnd.n4180 0.0174837
R12869 gnd.n4203 gnd.n4180 0.0174837
R12870 gnd.n4203 gnd.n4202 0.0174837
R12871 gnd.n4202 gnd.n4189 0.0174837
R12872 gnd.n4199 gnd.n4189 0.0174837
R12873 gnd.n4199 gnd.n4198 0.0174837
R12874 gnd.n4198 gnd.n2000 0.0174837
R12875 gnd.n2835 gnd.n2834 0.0148637
R12876 gnd.n3486 gnd.n3230 0.0144266
R12877 gnd.n3487 gnd.n3486 0.0130679
R12878 gnd.n2855 gnd.n2569 0.00797283
R12879 gnd.n2857 gnd.n2856 0.00797283
R12880 gnd.n2858 gnd.n2564 0.00797283
R12881 gnd.n2866 gnd.n2562 0.00797283
R12882 gnd.n2868 gnd.n2867 0.00797283
R12883 gnd.n2886 gnd.n2543 0.00797283
R12884 gnd.n2888 gnd.n2887 0.00797283
R12885 gnd.n2889 gnd.n2538 0.00797283
R12886 gnd.n2537 gnd.n2533 0.00797283
R12887 gnd.n2899 gnd.n2898 0.00797283
R12888 gnd.n2535 gnd.n2534 0.00797283
R12889 gnd.n2517 gnd.n2516 0.00797283
R12890 gnd.n2919 gnd.n2918 0.00797283
R12891 gnd.n2518 gnd.n2493 0.00797283
R12892 gnd.n2953 gnd.n2952 0.00797283
R12893 gnd.n2955 gnd.n2954 0.00797283
R12894 gnd.n2488 gnd.n2440 0.00797283
R12895 gnd.n2490 gnd.n2441 0.00797283
R12896 gnd.n2964 gnd.n2442 0.00797283
R12897 gnd.n2966 gnd.n2965 0.00797283
R12898 gnd.n2968 gnd.n2967 0.00797283
R12899 gnd.n2970 gnd.n2462 0.00797283
R12900 gnd.n2973 gnd.n2463 0.00797283
R12901 gnd.n2975 gnd.n2464 0.00797283
R12902 gnd.n2978 gnd.n2976 0.00797283
R12903 gnd.n2977 gnd.n2375 0.00797283
R12904 gnd.n3045 gnd.n3043 0.00797283
R12905 gnd.n3044 gnd.n2368 0.00797283
R12906 gnd.n3055 gnd.n3054 0.00797283
R12907 gnd.n3057 gnd.n3056 0.00797283
R12908 gnd.n3060 gnd.n2366 0.00797283
R12909 gnd.n3064 gnd.n3063 0.00797283
R12910 gnd.n3062 gnd.n3061 0.00797283
R12911 gnd.n2346 gnd.n2345 0.00797283
R12912 gnd.n3086 gnd.n3085 0.00797283
R12913 gnd.n2347 gnd.n2320 0.00797283
R12914 gnd.n3130 gnd.n3128 0.00797283
R12915 gnd.n3129 gnd.n2313 0.00797283
R12916 gnd.n3141 gnd.n3140 0.00797283
R12917 gnd.n3143 gnd.n3142 0.00797283
R12918 gnd.n3146 gnd.n2311 0.00797283
R12919 gnd.n3150 gnd.n3149 0.00797283
R12920 gnd.n3148 gnd.n3147 0.00797283
R12921 gnd.n2291 gnd.n2290 0.00797283
R12922 gnd.n3172 gnd.n3171 0.00797283
R12923 gnd.n2292 gnd.n2266 0.00797283
R12924 gnd.n3220 gnd.n3218 0.00797283
R12925 gnd.n3219 gnd.n2259 0.00797283
R12926 gnd.n3230 gnd.n3229 0.00797283
R12927 gnd.n3488 gnd.n3487 0.00797283
R12928 gnd.n3491 gnd.n2257 0.00797283
R12929 gnd.n3493 gnd.n3492 0.00797283
R12930 gnd.n3516 gnd.n2238 0.00797283
R12931 gnd.n3517 gnd.n2202 0.00797283
R12932 gnd.n5643 gnd.n1167 0.00614909
R12933 gnd.n3988 gnd.n3987 0.00614909
R12934 gnd.n5292 gnd.n5291 0.000839674
R12935 gnd.n4294 gnd.n4293 0.000839674
R12936 commonsourceibias.n25 commonsourceibias.t46 230.006
R12937 commonsourceibias.n91 commonsourceibias.t62 230.006
R12938 commonsourceibias.n154 commonsourceibias.t54 230.006
R12939 commonsourceibias.n258 commonsourceibias.t16 230.006
R12940 commonsourceibias.n217 commonsourceibias.t75 230.006
R12941 commonsourceibias.n355 commonsourceibias.t65 230.006
R12942 commonsourceibias.n70 commonsourceibias.t32 207.983
R12943 commonsourceibias.n136 commonsourceibias.t71 207.983
R12944 commonsourceibias.n199 commonsourceibias.t61 207.983
R12945 commonsourceibias.n304 commonsourceibias.t2 207.983
R12946 commonsourceibias.n338 commonsourceibias.t84 207.983
R12947 commonsourceibias.n401 commonsourceibias.t73 207.983
R12948 commonsourceibias.n10 commonsourceibias.t14 168.701
R12949 commonsourceibias.n63 commonsourceibias.t24 168.701
R12950 commonsourceibias.n57 commonsourceibias.t30 168.701
R12951 commonsourceibias.n16 commonsourceibias.t20 168.701
R12952 commonsourceibias.n49 commonsourceibias.t36 168.701
R12953 commonsourceibias.n43 commonsourceibias.t44 168.701
R12954 commonsourceibias.n19 commonsourceibias.t26 168.701
R12955 commonsourceibias.n21 commonsourceibias.t34 168.701
R12956 commonsourceibias.n23 commonsourceibias.t10 168.701
R12957 commonsourceibias.n26 commonsourceibias.t40 168.701
R12958 commonsourceibias.n1 commonsourceibias.t81 168.701
R12959 commonsourceibias.n129 commonsourceibias.t55 168.701
R12960 commonsourceibias.n123 commonsourceibias.t53 168.701
R12961 commonsourceibias.n7 commonsourceibias.t76 168.701
R12962 commonsourceibias.n115 commonsourceibias.t86 168.701
R12963 commonsourceibias.n109 commonsourceibias.t50 168.701
R12964 commonsourceibias.n85 commonsourceibias.t69 168.701
R12965 commonsourceibias.n87 commonsourceibias.t67 168.701
R12966 commonsourceibias.n89 commonsourceibias.t78 168.701
R12967 commonsourceibias.n92 commonsourceibias.t64 168.701
R12968 commonsourceibias.n155 commonsourceibias.t57 168.701
R12969 commonsourceibias.n152 commonsourceibias.t68 168.701
R12970 commonsourceibias.n150 commonsourceibias.t58 168.701
R12971 commonsourceibias.n148 commonsourceibias.t60 168.701
R12972 commonsourceibias.n172 commonsourceibias.t91 168.701
R12973 commonsourceibias.n178 commonsourceibias.t77 168.701
R12974 commonsourceibias.n145 commonsourceibias.t66 168.701
R12975 commonsourceibias.n186 commonsourceibias.t95 168.701
R12976 commonsourceibias.n192 commonsourceibias.t49 168.701
R12977 commonsourceibias.n139 commonsourceibias.t72 168.701
R12978 commonsourceibias.n259 commonsourceibias.t8 168.701
R12979 commonsourceibias.n256 commonsourceibias.t18 168.701
R12980 commonsourceibias.n254 commonsourceibias.t4 168.701
R12981 commonsourceibias.n252 commonsourceibias.t42 168.701
R12982 commonsourceibias.n276 commonsourceibias.t12 168.701
R12983 commonsourceibias.n282 commonsourceibias.t6 168.701
R12984 commonsourceibias.n284 commonsourceibias.t28 168.701
R12985 commonsourceibias.n291 commonsourceibias.t0 168.701
R12986 commonsourceibias.n297 commonsourceibias.t38 168.701
R12987 commonsourceibias.n244 commonsourceibias.t22 168.701
R12988 commonsourceibias.n203 commonsourceibias.t92 168.701
R12989 commonsourceibias.n331 commonsourceibias.t51 168.701
R12990 commonsourceibias.n325 commonsourceibias.t63 168.701
R12991 commonsourceibias.n318 commonsourceibias.t88 168.701
R12992 commonsourceibias.n316 commonsourceibias.t48 168.701
R12993 commonsourceibias.n218 commonsourceibias.t59 168.701
R12994 commonsourceibias.n215 commonsourceibias.t90 168.701
R12995 commonsourceibias.n213 commonsourceibias.t80 168.701
R12996 commonsourceibias.n211 commonsourceibias.t83 168.701
R12997 commonsourceibias.n235 commonsourceibias.t94 168.701
R12998 commonsourceibias.n356 commonsourceibias.t52 168.701
R12999 commonsourceibias.n353 commonsourceibias.t82 168.701
R13000 commonsourceibias.n351 commonsourceibias.t70 168.701
R13001 commonsourceibias.n349 commonsourceibias.t74 168.701
R13002 commonsourceibias.n373 commonsourceibias.t87 168.701
R13003 commonsourceibias.n379 commonsourceibias.t89 168.701
R13004 commonsourceibias.n381 commonsourceibias.t79 168.701
R13005 commonsourceibias.n388 commonsourceibias.t56 168.701
R13006 commonsourceibias.n394 commonsourceibias.t93 168.701
R13007 commonsourceibias.n341 commonsourceibias.t85 168.701
R13008 commonsourceibias.n27 commonsourceibias.n24 161.3
R13009 commonsourceibias.n29 commonsourceibias.n28 161.3
R13010 commonsourceibias.n31 commonsourceibias.n30 161.3
R13011 commonsourceibias.n32 commonsourceibias.n22 161.3
R13012 commonsourceibias.n34 commonsourceibias.n33 161.3
R13013 commonsourceibias.n36 commonsourceibias.n35 161.3
R13014 commonsourceibias.n37 commonsourceibias.n20 161.3
R13015 commonsourceibias.n39 commonsourceibias.n38 161.3
R13016 commonsourceibias.n41 commonsourceibias.n40 161.3
R13017 commonsourceibias.n42 commonsourceibias.n18 161.3
R13018 commonsourceibias.n45 commonsourceibias.n44 161.3
R13019 commonsourceibias.n46 commonsourceibias.n17 161.3
R13020 commonsourceibias.n48 commonsourceibias.n47 161.3
R13021 commonsourceibias.n50 commonsourceibias.n15 161.3
R13022 commonsourceibias.n52 commonsourceibias.n51 161.3
R13023 commonsourceibias.n53 commonsourceibias.n14 161.3
R13024 commonsourceibias.n55 commonsourceibias.n54 161.3
R13025 commonsourceibias.n56 commonsourceibias.n13 161.3
R13026 commonsourceibias.n59 commonsourceibias.n58 161.3
R13027 commonsourceibias.n60 commonsourceibias.n12 161.3
R13028 commonsourceibias.n62 commonsourceibias.n61 161.3
R13029 commonsourceibias.n64 commonsourceibias.n11 161.3
R13030 commonsourceibias.n66 commonsourceibias.n65 161.3
R13031 commonsourceibias.n68 commonsourceibias.n67 161.3
R13032 commonsourceibias.n69 commonsourceibias.n9 161.3
R13033 commonsourceibias.n93 commonsourceibias.n90 161.3
R13034 commonsourceibias.n95 commonsourceibias.n94 161.3
R13035 commonsourceibias.n97 commonsourceibias.n96 161.3
R13036 commonsourceibias.n98 commonsourceibias.n88 161.3
R13037 commonsourceibias.n100 commonsourceibias.n99 161.3
R13038 commonsourceibias.n102 commonsourceibias.n101 161.3
R13039 commonsourceibias.n103 commonsourceibias.n86 161.3
R13040 commonsourceibias.n105 commonsourceibias.n104 161.3
R13041 commonsourceibias.n107 commonsourceibias.n106 161.3
R13042 commonsourceibias.n108 commonsourceibias.n84 161.3
R13043 commonsourceibias.n111 commonsourceibias.n110 161.3
R13044 commonsourceibias.n112 commonsourceibias.n8 161.3
R13045 commonsourceibias.n114 commonsourceibias.n113 161.3
R13046 commonsourceibias.n116 commonsourceibias.n6 161.3
R13047 commonsourceibias.n118 commonsourceibias.n117 161.3
R13048 commonsourceibias.n119 commonsourceibias.n5 161.3
R13049 commonsourceibias.n121 commonsourceibias.n120 161.3
R13050 commonsourceibias.n122 commonsourceibias.n4 161.3
R13051 commonsourceibias.n125 commonsourceibias.n124 161.3
R13052 commonsourceibias.n126 commonsourceibias.n3 161.3
R13053 commonsourceibias.n128 commonsourceibias.n127 161.3
R13054 commonsourceibias.n130 commonsourceibias.n2 161.3
R13055 commonsourceibias.n132 commonsourceibias.n131 161.3
R13056 commonsourceibias.n134 commonsourceibias.n133 161.3
R13057 commonsourceibias.n135 commonsourceibias.n0 161.3
R13058 commonsourceibias.n198 commonsourceibias.n138 161.3
R13059 commonsourceibias.n197 commonsourceibias.n196 161.3
R13060 commonsourceibias.n195 commonsourceibias.n194 161.3
R13061 commonsourceibias.n193 commonsourceibias.n140 161.3
R13062 commonsourceibias.n191 commonsourceibias.n190 161.3
R13063 commonsourceibias.n189 commonsourceibias.n141 161.3
R13064 commonsourceibias.n188 commonsourceibias.n187 161.3
R13065 commonsourceibias.n185 commonsourceibias.n142 161.3
R13066 commonsourceibias.n184 commonsourceibias.n183 161.3
R13067 commonsourceibias.n182 commonsourceibias.n143 161.3
R13068 commonsourceibias.n181 commonsourceibias.n180 161.3
R13069 commonsourceibias.n179 commonsourceibias.n144 161.3
R13070 commonsourceibias.n177 commonsourceibias.n176 161.3
R13071 commonsourceibias.n175 commonsourceibias.n146 161.3
R13072 commonsourceibias.n174 commonsourceibias.n173 161.3
R13073 commonsourceibias.n171 commonsourceibias.n147 161.3
R13074 commonsourceibias.n170 commonsourceibias.n169 161.3
R13075 commonsourceibias.n168 commonsourceibias.n167 161.3
R13076 commonsourceibias.n166 commonsourceibias.n149 161.3
R13077 commonsourceibias.n165 commonsourceibias.n164 161.3
R13078 commonsourceibias.n163 commonsourceibias.n162 161.3
R13079 commonsourceibias.n161 commonsourceibias.n151 161.3
R13080 commonsourceibias.n160 commonsourceibias.n159 161.3
R13081 commonsourceibias.n158 commonsourceibias.n157 161.3
R13082 commonsourceibias.n156 commonsourceibias.n153 161.3
R13083 commonsourceibias.n303 commonsourceibias.n243 161.3
R13084 commonsourceibias.n302 commonsourceibias.n301 161.3
R13085 commonsourceibias.n300 commonsourceibias.n299 161.3
R13086 commonsourceibias.n298 commonsourceibias.n245 161.3
R13087 commonsourceibias.n296 commonsourceibias.n295 161.3
R13088 commonsourceibias.n294 commonsourceibias.n246 161.3
R13089 commonsourceibias.n293 commonsourceibias.n292 161.3
R13090 commonsourceibias.n290 commonsourceibias.n247 161.3
R13091 commonsourceibias.n289 commonsourceibias.n288 161.3
R13092 commonsourceibias.n287 commonsourceibias.n248 161.3
R13093 commonsourceibias.n286 commonsourceibias.n285 161.3
R13094 commonsourceibias.n283 commonsourceibias.n249 161.3
R13095 commonsourceibias.n281 commonsourceibias.n280 161.3
R13096 commonsourceibias.n279 commonsourceibias.n250 161.3
R13097 commonsourceibias.n278 commonsourceibias.n277 161.3
R13098 commonsourceibias.n275 commonsourceibias.n251 161.3
R13099 commonsourceibias.n274 commonsourceibias.n273 161.3
R13100 commonsourceibias.n272 commonsourceibias.n271 161.3
R13101 commonsourceibias.n270 commonsourceibias.n253 161.3
R13102 commonsourceibias.n269 commonsourceibias.n268 161.3
R13103 commonsourceibias.n267 commonsourceibias.n266 161.3
R13104 commonsourceibias.n265 commonsourceibias.n255 161.3
R13105 commonsourceibias.n264 commonsourceibias.n263 161.3
R13106 commonsourceibias.n262 commonsourceibias.n261 161.3
R13107 commonsourceibias.n260 commonsourceibias.n257 161.3
R13108 commonsourceibias.n237 commonsourceibias.n236 161.3
R13109 commonsourceibias.n234 commonsourceibias.n210 161.3
R13110 commonsourceibias.n233 commonsourceibias.n232 161.3
R13111 commonsourceibias.n231 commonsourceibias.n230 161.3
R13112 commonsourceibias.n229 commonsourceibias.n212 161.3
R13113 commonsourceibias.n228 commonsourceibias.n227 161.3
R13114 commonsourceibias.n226 commonsourceibias.n225 161.3
R13115 commonsourceibias.n224 commonsourceibias.n214 161.3
R13116 commonsourceibias.n223 commonsourceibias.n222 161.3
R13117 commonsourceibias.n221 commonsourceibias.n220 161.3
R13118 commonsourceibias.n219 commonsourceibias.n216 161.3
R13119 commonsourceibias.n313 commonsourceibias.n209 161.3
R13120 commonsourceibias.n337 commonsourceibias.n202 161.3
R13121 commonsourceibias.n336 commonsourceibias.n335 161.3
R13122 commonsourceibias.n334 commonsourceibias.n333 161.3
R13123 commonsourceibias.n332 commonsourceibias.n204 161.3
R13124 commonsourceibias.n330 commonsourceibias.n329 161.3
R13125 commonsourceibias.n328 commonsourceibias.n205 161.3
R13126 commonsourceibias.n327 commonsourceibias.n326 161.3
R13127 commonsourceibias.n324 commonsourceibias.n206 161.3
R13128 commonsourceibias.n323 commonsourceibias.n322 161.3
R13129 commonsourceibias.n321 commonsourceibias.n207 161.3
R13130 commonsourceibias.n320 commonsourceibias.n319 161.3
R13131 commonsourceibias.n317 commonsourceibias.n208 161.3
R13132 commonsourceibias.n315 commonsourceibias.n314 161.3
R13133 commonsourceibias.n400 commonsourceibias.n340 161.3
R13134 commonsourceibias.n399 commonsourceibias.n398 161.3
R13135 commonsourceibias.n397 commonsourceibias.n396 161.3
R13136 commonsourceibias.n395 commonsourceibias.n342 161.3
R13137 commonsourceibias.n393 commonsourceibias.n392 161.3
R13138 commonsourceibias.n391 commonsourceibias.n343 161.3
R13139 commonsourceibias.n390 commonsourceibias.n389 161.3
R13140 commonsourceibias.n387 commonsourceibias.n344 161.3
R13141 commonsourceibias.n386 commonsourceibias.n385 161.3
R13142 commonsourceibias.n384 commonsourceibias.n345 161.3
R13143 commonsourceibias.n383 commonsourceibias.n382 161.3
R13144 commonsourceibias.n380 commonsourceibias.n346 161.3
R13145 commonsourceibias.n378 commonsourceibias.n377 161.3
R13146 commonsourceibias.n376 commonsourceibias.n347 161.3
R13147 commonsourceibias.n375 commonsourceibias.n374 161.3
R13148 commonsourceibias.n372 commonsourceibias.n348 161.3
R13149 commonsourceibias.n371 commonsourceibias.n370 161.3
R13150 commonsourceibias.n369 commonsourceibias.n368 161.3
R13151 commonsourceibias.n367 commonsourceibias.n350 161.3
R13152 commonsourceibias.n366 commonsourceibias.n365 161.3
R13153 commonsourceibias.n364 commonsourceibias.n363 161.3
R13154 commonsourceibias.n362 commonsourceibias.n352 161.3
R13155 commonsourceibias.n361 commonsourceibias.n360 161.3
R13156 commonsourceibias.n359 commonsourceibias.n358 161.3
R13157 commonsourceibias.n357 commonsourceibias.n354 161.3
R13158 commonsourceibias.n80 commonsourceibias.n78 81.5057
R13159 commonsourceibias.n240 commonsourceibias.n238 81.5057
R13160 commonsourceibias.n80 commonsourceibias.n79 80.9324
R13161 commonsourceibias.n82 commonsourceibias.n81 80.9324
R13162 commonsourceibias.n77 commonsourceibias.n76 80.9324
R13163 commonsourceibias.n75 commonsourceibias.n74 80.9324
R13164 commonsourceibias.n73 commonsourceibias.n72 80.9324
R13165 commonsourceibias.n307 commonsourceibias.n306 80.9324
R13166 commonsourceibias.n309 commonsourceibias.n308 80.9324
R13167 commonsourceibias.n311 commonsourceibias.n310 80.9324
R13168 commonsourceibias.n242 commonsourceibias.n241 80.9324
R13169 commonsourceibias.n240 commonsourceibias.n239 80.9324
R13170 commonsourceibias.n71 commonsourceibias.n70 80.6037
R13171 commonsourceibias.n137 commonsourceibias.n136 80.6037
R13172 commonsourceibias.n200 commonsourceibias.n199 80.6037
R13173 commonsourceibias.n305 commonsourceibias.n304 80.6037
R13174 commonsourceibias.n339 commonsourceibias.n338 80.6037
R13175 commonsourceibias.n402 commonsourceibias.n401 80.6037
R13176 commonsourceibias.n65 commonsourceibias.n64 56.5617
R13177 commonsourceibias.n51 commonsourceibias.n50 56.5617
R13178 commonsourceibias.n42 commonsourceibias.n41 56.5617
R13179 commonsourceibias.n28 commonsourceibias.n27 56.5617
R13180 commonsourceibias.n131 commonsourceibias.n130 56.5617
R13181 commonsourceibias.n117 commonsourceibias.n116 56.5617
R13182 commonsourceibias.n108 commonsourceibias.n107 56.5617
R13183 commonsourceibias.n94 commonsourceibias.n93 56.5617
R13184 commonsourceibias.n157 commonsourceibias.n156 56.5617
R13185 commonsourceibias.n171 commonsourceibias.n170 56.5617
R13186 commonsourceibias.n180 commonsourceibias.n179 56.5617
R13187 commonsourceibias.n194 commonsourceibias.n193 56.5617
R13188 commonsourceibias.n261 commonsourceibias.n260 56.5617
R13189 commonsourceibias.n275 commonsourceibias.n274 56.5617
R13190 commonsourceibias.n285 commonsourceibias.n283 56.5617
R13191 commonsourceibias.n299 commonsourceibias.n298 56.5617
R13192 commonsourceibias.n333 commonsourceibias.n332 56.5617
R13193 commonsourceibias.n319 commonsourceibias.n317 56.5617
R13194 commonsourceibias.n220 commonsourceibias.n219 56.5617
R13195 commonsourceibias.n234 commonsourceibias.n233 56.5617
R13196 commonsourceibias.n358 commonsourceibias.n357 56.5617
R13197 commonsourceibias.n372 commonsourceibias.n371 56.5617
R13198 commonsourceibias.n382 commonsourceibias.n380 56.5617
R13199 commonsourceibias.n396 commonsourceibias.n395 56.5617
R13200 commonsourceibias.n56 commonsourceibias.n55 56.0773
R13201 commonsourceibias.n37 commonsourceibias.n36 56.0773
R13202 commonsourceibias.n122 commonsourceibias.n121 56.0773
R13203 commonsourceibias.n103 commonsourceibias.n102 56.0773
R13204 commonsourceibias.n166 commonsourceibias.n165 56.0773
R13205 commonsourceibias.n185 commonsourceibias.n184 56.0773
R13206 commonsourceibias.n270 commonsourceibias.n269 56.0773
R13207 commonsourceibias.n290 commonsourceibias.n289 56.0773
R13208 commonsourceibias.n324 commonsourceibias.n323 56.0773
R13209 commonsourceibias.n229 commonsourceibias.n228 56.0773
R13210 commonsourceibias.n367 commonsourceibias.n366 56.0773
R13211 commonsourceibias.n387 commonsourceibias.n386 56.0773
R13212 commonsourceibias.n70 commonsourceibias.n69 46.0096
R13213 commonsourceibias.n136 commonsourceibias.n135 46.0096
R13214 commonsourceibias.n199 commonsourceibias.n198 46.0096
R13215 commonsourceibias.n304 commonsourceibias.n303 46.0096
R13216 commonsourceibias.n338 commonsourceibias.n337 46.0096
R13217 commonsourceibias.n401 commonsourceibias.n400 46.0096
R13218 commonsourceibias.n58 commonsourceibias.n12 41.5458
R13219 commonsourceibias.n33 commonsourceibias.n32 41.5458
R13220 commonsourceibias.n124 commonsourceibias.n3 41.5458
R13221 commonsourceibias.n99 commonsourceibias.n98 41.5458
R13222 commonsourceibias.n162 commonsourceibias.n161 41.5458
R13223 commonsourceibias.n187 commonsourceibias.n141 41.5458
R13224 commonsourceibias.n266 commonsourceibias.n265 41.5458
R13225 commonsourceibias.n292 commonsourceibias.n246 41.5458
R13226 commonsourceibias.n326 commonsourceibias.n205 41.5458
R13227 commonsourceibias.n225 commonsourceibias.n224 41.5458
R13228 commonsourceibias.n363 commonsourceibias.n362 41.5458
R13229 commonsourceibias.n389 commonsourceibias.n343 41.5458
R13230 commonsourceibias.n48 commonsourceibias.n17 40.577
R13231 commonsourceibias.n44 commonsourceibias.n17 40.577
R13232 commonsourceibias.n114 commonsourceibias.n8 40.577
R13233 commonsourceibias.n110 commonsourceibias.n8 40.577
R13234 commonsourceibias.n173 commonsourceibias.n146 40.577
R13235 commonsourceibias.n177 commonsourceibias.n146 40.577
R13236 commonsourceibias.n277 commonsourceibias.n250 40.577
R13237 commonsourceibias.n281 commonsourceibias.n250 40.577
R13238 commonsourceibias.n315 commonsourceibias.n209 40.577
R13239 commonsourceibias.n236 commonsourceibias.n209 40.577
R13240 commonsourceibias.n374 commonsourceibias.n347 40.577
R13241 commonsourceibias.n378 commonsourceibias.n347 40.577
R13242 commonsourceibias.n62 commonsourceibias.n12 39.6083
R13243 commonsourceibias.n32 commonsourceibias.n31 39.6083
R13244 commonsourceibias.n128 commonsourceibias.n3 39.6083
R13245 commonsourceibias.n98 commonsourceibias.n97 39.6083
R13246 commonsourceibias.n161 commonsourceibias.n160 39.6083
R13247 commonsourceibias.n191 commonsourceibias.n141 39.6083
R13248 commonsourceibias.n265 commonsourceibias.n264 39.6083
R13249 commonsourceibias.n296 commonsourceibias.n246 39.6083
R13250 commonsourceibias.n330 commonsourceibias.n205 39.6083
R13251 commonsourceibias.n224 commonsourceibias.n223 39.6083
R13252 commonsourceibias.n362 commonsourceibias.n361 39.6083
R13253 commonsourceibias.n393 commonsourceibias.n343 39.6083
R13254 commonsourceibias.n26 commonsourceibias.n25 33.0515
R13255 commonsourceibias.n92 commonsourceibias.n91 33.0515
R13256 commonsourceibias.n155 commonsourceibias.n154 33.0515
R13257 commonsourceibias.n259 commonsourceibias.n258 33.0515
R13258 commonsourceibias.n218 commonsourceibias.n217 33.0515
R13259 commonsourceibias.n356 commonsourceibias.n355 33.0515
R13260 commonsourceibias.n25 commonsourceibias.n24 28.5514
R13261 commonsourceibias.n91 commonsourceibias.n90 28.5514
R13262 commonsourceibias.n154 commonsourceibias.n153 28.5514
R13263 commonsourceibias.n258 commonsourceibias.n257 28.5514
R13264 commonsourceibias.n217 commonsourceibias.n216 28.5514
R13265 commonsourceibias.n355 commonsourceibias.n354 28.5514
R13266 commonsourceibias.n69 commonsourceibias.n68 26.0455
R13267 commonsourceibias.n135 commonsourceibias.n134 26.0455
R13268 commonsourceibias.n198 commonsourceibias.n197 26.0455
R13269 commonsourceibias.n303 commonsourceibias.n302 26.0455
R13270 commonsourceibias.n337 commonsourceibias.n336 26.0455
R13271 commonsourceibias.n400 commonsourceibias.n399 26.0455
R13272 commonsourceibias.n55 commonsourceibias.n14 25.0767
R13273 commonsourceibias.n38 commonsourceibias.n37 25.0767
R13274 commonsourceibias.n121 commonsourceibias.n5 25.0767
R13275 commonsourceibias.n104 commonsourceibias.n103 25.0767
R13276 commonsourceibias.n167 commonsourceibias.n166 25.0767
R13277 commonsourceibias.n184 commonsourceibias.n143 25.0767
R13278 commonsourceibias.n271 commonsourceibias.n270 25.0767
R13279 commonsourceibias.n289 commonsourceibias.n248 25.0767
R13280 commonsourceibias.n323 commonsourceibias.n207 25.0767
R13281 commonsourceibias.n230 commonsourceibias.n229 25.0767
R13282 commonsourceibias.n368 commonsourceibias.n367 25.0767
R13283 commonsourceibias.n386 commonsourceibias.n345 25.0767
R13284 commonsourceibias.n51 commonsourceibias.n16 24.3464
R13285 commonsourceibias.n41 commonsourceibias.n19 24.3464
R13286 commonsourceibias.n117 commonsourceibias.n7 24.3464
R13287 commonsourceibias.n107 commonsourceibias.n85 24.3464
R13288 commonsourceibias.n170 commonsourceibias.n148 24.3464
R13289 commonsourceibias.n180 commonsourceibias.n145 24.3464
R13290 commonsourceibias.n274 commonsourceibias.n252 24.3464
R13291 commonsourceibias.n285 commonsourceibias.n284 24.3464
R13292 commonsourceibias.n319 commonsourceibias.n318 24.3464
R13293 commonsourceibias.n233 commonsourceibias.n211 24.3464
R13294 commonsourceibias.n371 commonsourceibias.n349 24.3464
R13295 commonsourceibias.n382 commonsourceibias.n381 24.3464
R13296 commonsourceibias.n65 commonsourceibias.n10 23.8546
R13297 commonsourceibias.n27 commonsourceibias.n26 23.8546
R13298 commonsourceibias.n131 commonsourceibias.n1 23.8546
R13299 commonsourceibias.n93 commonsourceibias.n92 23.8546
R13300 commonsourceibias.n156 commonsourceibias.n155 23.8546
R13301 commonsourceibias.n194 commonsourceibias.n139 23.8546
R13302 commonsourceibias.n260 commonsourceibias.n259 23.8546
R13303 commonsourceibias.n299 commonsourceibias.n244 23.8546
R13304 commonsourceibias.n333 commonsourceibias.n203 23.8546
R13305 commonsourceibias.n219 commonsourceibias.n218 23.8546
R13306 commonsourceibias.n357 commonsourceibias.n356 23.8546
R13307 commonsourceibias.n396 commonsourceibias.n341 23.8546
R13308 commonsourceibias.n64 commonsourceibias.n63 16.9689
R13309 commonsourceibias.n28 commonsourceibias.n23 16.9689
R13310 commonsourceibias.n130 commonsourceibias.n129 16.9689
R13311 commonsourceibias.n94 commonsourceibias.n89 16.9689
R13312 commonsourceibias.n157 commonsourceibias.n152 16.9689
R13313 commonsourceibias.n193 commonsourceibias.n192 16.9689
R13314 commonsourceibias.n261 commonsourceibias.n256 16.9689
R13315 commonsourceibias.n298 commonsourceibias.n297 16.9689
R13316 commonsourceibias.n332 commonsourceibias.n331 16.9689
R13317 commonsourceibias.n220 commonsourceibias.n215 16.9689
R13318 commonsourceibias.n358 commonsourceibias.n353 16.9689
R13319 commonsourceibias.n395 commonsourceibias.n394 16.9689
R13320 commonsourceibias.n50 commonsourceibias.n49 16.477
R13321 commonsourceibias.n43 commonsourceibias.n42 16.477
R13322 commonsourceibias.n116 commonsourceibias.n115 16.477
R13323 commonsourceibias.n109 commonsourceibias.n108 16.477
R13324 commonsourceibias.n172 commonsourceibias.n171 16.477
R13325 commonsourceibias.n179 commonsourceibias.n178 16.477
R13326 commonsourceibias.n276 commonsourceibias.n275 16.477
R13327 commonsourceibias.n283 commonsourceibias.n282 16.477
R13328 commonsourceibias.n317 commonsourceibias.n316 16.477
R13329 commonsourceibias.n235 commonsourceibias.n234 16.477
R13330 commonsourceibias.n373 commonsourceibias.n372 16.477
R13331 commonsourceibias.n380 commonsourceibias.n379 16.477
R13332 commonsourceibias.n57 commonsourceibias.n56 15.9852
R13333 commonsourceibias.n36 commonsourceibias.n21 15.9852
R13334 commonsourceibias.n123 commonsourceibias.n122 15.9852
R13335 commonsourceibias.n102 commonsourceibias.n87 15.9852
R13336 commonsourceibias.n165 commonsourceibias.n150 15.9852
R13337 commonsourceibias.n186 commonsourceibias.n185 15.9852
R13338 commonsourceibias.n269 commonsourceibias.n254 15.9852
R13339 commonsourceibias.n291 commonsourceibias.n290 15.9852
R13340 commonsourceibias.n325 commonsourceibias.n324 15.9852
R13341 commonsourceibias.n228 commonsourceibias.n213 15.9852
R13342 commonsourceibias.n366 commonsourceibias.n351 15.9852
R13343 commonsourceibias.n388 commonsourceibias.n387 15.9852
R13344 commonsourceibias.n73 commonsourceibias.n71 13.2057
R13345 commonsourceibias.n307 commonsourceibias.n305 13.2057
R13346 commonsourceibias.n404 commonsourceibias.n201 11.9876
R13347 commonsourceibias.n404 commonsourceibias.n403 10.3347
R13348 commonsourceibias.n112 commonsourceibias.n83 9.50363
R13349 commonsourceibias.n313 commonsourceibias.n312 9.50363
R13350 commonsourceibias.n201 commonsourceibias.n137 8.732
R13351 commonsourceibias.n403 commonsourceibias.n339 8.732
R13352 commonsourceibias.n58 commonsourceibias.n57 8.60764
R13353 commonsourceibias.n33 commonsourceibias.n21 8.60764
R13354 commonsourceibias.n124 commonsourceibias.n123 8.60764
R13355 commonsourceibias.n99 commonsourceibias.n87 8.60764
R13356 commonsourceibias.n162 commonsourceibias.n150 8.60764
R13357 commonsourceibias.n187 commonsourceibias.n186 8.60764
R13358 commonsourceibias.n266 commonsourceibias.n254 8.60764
R13359 commonsourceibias.n292 commonsourceibias.n291 8.60764
R13360 commonsourceibias.n326 commonsourceibias.n325 8.60764
R13361 commonsourceibias.n225 commonsourceibias.n213 8.60764
R13362 commonsourceibias.n363 commonsourceibias.n351 8.60764
R13363 commonsourceibias.n389 commonsourceibias.n388 8.60764
R13364 commonsourceibias.n49 commonsourceibias.n48 8.11581
R13365 commonsourceibias.n44 commonsourceibias.n43 8.11581
R13366 commonsourceibias.n115 commonsourceibias.n114 8.11581
R13367 commonsourceibias.n110 commonsourceibias.n109 8.11581
R13368 commonsourceibias.n173 commonsourceibias.n172 8.11581
R13369 commonsourceibias.n178 commonsourceibias.n177 8.11581
R13370 commonsourceibias.n277 commonsourceibias.n276 8.11581
R13371 commonsourceibias.n282 commonsourceibias.n281 8.11581
R13372 commonsourceibias.n316 commonsourceibias.n315 8.11581
R13373 commonsourceibias.n236 commonsourceibias.n235 8.11581
R13374 commonsourceibias.n374 commonsourceibias.n373 8.11581
R13375 commonsourceibias.n379 commonsourceibias.n378 8.11581
R13376 commonsourceibias.n63 commonsourceibias.n62 7.62397
R13377 commonsourceibias.n31 commonsourceibias.n23 7.62397
R13378 commonsourceibias.n129 commonsourceibias.n128 7.62397
R13379 commonsourceibias.n97 commonsourceibias.n89 7.62397
R13380 commonsourceibias.n160 commonsourceibias.n152 7.62397
R13381 commonsourceibias.n192 commonsourceibias.n191 7.62397
R13382 commonsourceibias.n264 commonsourceibias.n256 7.62397
R13383 commonsourceibias.n297 commonsourceibias.n296 7.62397
R13384 commonsourceibias.n331 commonsourceibias.n330 7.62397
R13385 commonsourceibias.n223 commonsourceibias.n215 7.62397
R13386 commonsourceibias.n361 commonsourceibias.n353 7.62397
R13387 commonsourceibias.n394 commonsourceibias.n393 7.62397
R13388 commonsourceibias.n201 commonsourceibias.n200 5.00473
R13389 commonsourceibias.n403 commonsourceibias.n402 5.00473
R13390 commonsourceibias commonsourceibias.n404 3.87639
R13391 commonsourceibias.n78 commonsourceibias.t41 2.82907
R13392 commonsourceibias.n78 commonsourceibias.t47 2.82907
R13393 commonsourceibias.n79 commonsourceibias.t35 2.82907
R13394 commonsourceibias.n79 commonsourceibias.t11 2.82907
R13395 commonsourceibias.n81 commonsourceibias.t45 2.82907
R13396 commonsourceibias.n81 commonsourceibias.t27 2.82907
R13397 commonsourceibias.n76 commonsourceibias.t21 2.82907
R13398 commonsourceibias.n76 commonsourceibias.t37 2.82907
R13399 commonsourceibias.n74 commonsourceibias.t25 2.82907
R13400 commonsourceibias.n74 commonsourceibias.t31 2.82907
R13401 commonsourceibias.n72 commonsourceibias.t33 2.82907
R13402 commonsourceibias.n72 commonsourceibias.t15 2.82907
R13403 commonsourceibias.n306 commonsourceibias.t23 2.82907
R13404 commonsourceibias.n306 commonsourceibias.t3 2.82907
R13405 commonsourceibias.n308 commonsourceibias.t1 2.82907
R13406 commonsourceibias.n308 commonsourceibias.t39 2.82907
R13407 commonsourceibias.n310 commonsourceibias.t7 2.82907
R13408 commonsourceibias.n310 commonsourceibias.t29 2.82907
R13409 commonsourceibias.n241 commonsourceibias.t43 2.82907
R13410 commonsourceibias.n241 commonsourceibias.t13 2.82907
R13411 commonsourceibias.n239 commonsourceibias.t19 2.82907
R13412 commonsourceibias.n239 commonsourceibias.t5 2.82907
R13413 commonsourceibias.n238 commonsourceibias.t17 2.82907
R13414 commonsourceibias.n238 commonsourceibias.t9 2.82907
R13415 commonsourceibias.n68 commonsourceibias.n10 0.738255
R13416 commonsourceibias.n134 commonsourceibias.n1 0.738255
R13417 commonsourceibias.n197 commonsourceibias.n139 0.738255
R13418 commonsourceibias.n302 commonsourceibias.n244 0.738255
R13419 commonsourceibias.n336 commonsourceibias.n203 0.738255
R13420 commonsourceibias.n399 commonsourceibias.n341 0.738255
R13421 commonsourceibias.n75 commonsourceibias.n73 0.573776
R13422 commonsourceibias.n77 commonsourceibias.n75 0.573776
R13423 commonsourceibias.n82 commonsourceibias.n80 0.573776
R13424 commonsourceibias.n242 commonsourceibias.n240 0.573776
R13425 commonsourceibias.n311 commonsourceibias.n309 0.573776
R13426 commonsourceibias.n309 commonsourceibias.n307 0.573776
R13427 commonsourceibias.n83 commonsourceibias.n77 0.287138
R13428 commonsourceibias.n83 commonsourceibias.n82 0.287138
R13429 commonsourceibias.n312 commonsourceibias.n242 0.287138
R13430 commonsourceibias.n312 commonsourceibias.n311 0.287138
R13431 commonsourceibias.n71 commonsourceibias.n9 0.285035
R13432 commonsourceibias.n137 commonsourceibias.n0 0.285035
R13433 commonsourceibias.n200 commonsourceibias.n138 0.285035
R13434 commonsourceibias.n305 commonsourceibias.n243 0.285035
R13435 commonsourceibias.n339 commonsourceibias.n202 0.285035
R13436 commonsourceibias.n402 commonsourceibias.n340 0.285035
R13437 commonsourceibias.n16 commonsourceibias.n14 0.246418
R13438 commonsourceibias.n38 commonsourceibias.n19 0.246418
R13439 commonsourceibias.n7 commonsourceibias.n5 0.246418
R13440 commonsourceibias.n104 commonsourceibias.n85 0.246418
R13441 commonsourceibias.n167 commonsourceibias.n148 0.246418
R13442 commonsourceibias.n145 commonsourceibias.n143 0.246418
R13443 commonsourceibias.n271 commonsourceibias.n252 0.246418
R13444 commonsourceibias.n284 commonsourceibias.n248 0.246418
R13445 commonsourceibias.n318 commonsourceibias.n207 0.246418
R13446 commonsourceibias.n230 commonsourceibias.n211 0.246418
R13447 commonsourceibias.n368 commonsourceibias.n349 0.246418
R13448 commonsourceibias.n381 commonsourceibias.n345 0.246418
R13449 commonsourceibias.n67 commonsourceibias.n9 0.189894
R13450 commonsourceibias.n67 commonsourceibias.n66 0.189894
R13451 commonsourceibias.n66 commonsourceibias.n11 0.189894
R13452 commonsourceibias.n61 commonsourceibias.n11 0.189894
R13453 commonsourceibias.n61 commonsourceibias.n60 0.189894
R13454 commonsourceibias.n60 commonsourceibias.n59 0.189894
R13455 commonsourceibias.n59 commonsourceibias.n13 0.189894
R13456 commonsourceibias.n54 commonsourceibias.n13 0.189894
R13457 commonsourceibias.n54 commonsourceibias.n53 0.189894
R13458 commonsourceibias.n53 commonsourceibias.n52 0.189894
R13459 commonsourceibias.n52 commonsourceibias.n15 0.189894
R13460 commonsourceibias.n47 commonsourceibias.n15 0.189894
R13461 commonsourceibias.n47 commonsourceibias.n46 0.189894
R13462 commonsourceibias.n46 commonsourceibias.n45 0.189894
R13463 commonsourceibias.n45 commonsourceibias.n18 0.189894
R13464 commonsourceibias.n40 commonsourceibias.n18 0.189894
R13465 commonsourceibias.n40 commonsourceibias.n39 0.189894
R13466 commonsourceibias.n39 commonsourceibias.n20 0.189894
R13467 commonsourceibias.n35 commonsourceibias.n20 0.189894
R13468 commonsourceibias.n35 commonsourceibias.n34 0.189894
R13469 commonsourceibias.n34 commonsourceibias.n22 0.189894
R13470 commonsourceibias.n30 commonsourceibias.n22 0.189894
R13471 commonsourceibias.n30 commonsourceibias.n29 0.189894
R13472 commonsourceibias.n29 commonsourceibias.n24 0.189894
R13473 commonsourceibias.n111 commonsourceibias.n84 0.189894
R13474 commonsourceibias.n106 commonsourceibias.n84 0.189894
R13475 commonsourceibias.n106 commonsourceibias.n105 0.189894
R13476 commonsourceibias.n105 commonsourceibias.n86 0.189894
R13477 commonsourceibias.n101 commonsourceibias.n86 0.189894
R13478 commonsourceibias.n101 commonsourceibias.n100 0.189894
R13479 commonsourceibias.n100 commonsourceibias.n88 0.189894
R13480 commonsourceibias.n96 commonsourceibias.n88 0.189894
R13481 commonsourceibias.n96 commonsourceibias.n95 0.189894
R13482 commonsourceibias.n95 commonsourceibias.n90 0.189894
R13483 commonsourceibias.n133 commonsourceibias.n0 0.189894
R13484 commonsourceibias.n133 commonsourceibias.n132 0.189894
R13485 commonsourceibias.n132 commonsourceibias.n2 0.189894
R13486 commonsourceibias.n127 commonsourceibias.n2 0.189894
R13487 commonsourceibias.n127 commonsourceibias.n126 0.189894
R13488 commonsourceibias.n126 commonsourceibias.n125 0.189894
R13489 commonsourceibias.n125 commonsourceibias.n4 0.189894
R13490 commonsourceibias.n120 commonsourceibias.n4 0.189894
R13491 commonsourceibias.n120 commonsourceibias.n119 0.189894
R13492 commonsourceibias.n119 commonsourceibias.n118 0.189894
R13493 commonsourceibias.n118 commonsourceibias.n6 0.189894
R13494 commonsourceibias.n113 commonsourceibias.n6 0.189894
R13495 commonsourceibias.n196 commonsourceibias.n138 0.189894
R13496 commonsourceibias.n196 commonsourceibias.n195 0.189894
R13497 commonsourceibias.n195 commonsourceibias.n140 0.189894
R13498 commonsourceibias.n190 commonsourceibias.n140 0.189894
R13499 commonsourceibias.n190 commonsourceibias.n189 0.189894
R13500 commonsourceibias.n189 commonsourceibias.n188 0.189894
R13501 commonsourceibias.n188 commonsourceibias.n142 0.189894
R13502 commonsourceibias.n183 commonsourceibias.n142 0.189894
R13503 commonsourceibias.n183 commonsourceibias.n182 0.189894
R13504 commonsourceibias.n182 commonsourceibias.n181 0.189894
R13505 commonsourceibias.n181 commonsourceibias.n144 0.189894
R13506 commonsourceibias.n176 commonsourceibias.n144 0.189894
R13507 commonsourceibias.n176 commonsourceibias.n175 0.189894
R13508 commonsourceibias.n175 commonsourceibias.n174 0.189894
R13509 commonsourceibias.n174 commonsourceibias.n147 0.189894
R13510 commonsourceibias.n169 commonsourceibias.n147 0.189894
R13511 commonsourceibias.n169 commonsourceibias.n168 0.189894
R13512 commonsourceibias.n168 commonsourceibias.n149 0.189894
R13513 commonsourceibias.n164 commonsourceibias.n149 0.189894
R13514 commonsourceibias.n164 commonsourceibias.n163 0.189894
R13515 commonsourceibias.n163 commonsourceibias.n151 0.189894
R13516 commonsourceibias.n159 commonsourceibias.n151 0.189894
R13517 commonsourceibias.n159 commonsourceibias.n158 0.189894
R13518 commonsourceibias.n158 commonsourceibias.n153 0.189894
R13519 commonsourceibias.n262 commonsourceibias.n257 0.189894
R13520 commonsourceibias.n263 commonsourceibias.n262 0.189894
R13521 commonsourceibias.n263 commonsourceibias.n255 0.189894
R13522 commonsourceibias.n267 commonsourceibias.n255 0.189894
R13523 commonsourceibias.n268 commonsourceibias.n267 0.189894
R13524 commonsourceibias.n268 commonsourceibias.n253 0.189894
R13525 commonsourceibias.n272 commonsourceibias.n253 0.189894
R13526 commonsourceibias.n273 commonsourceibias.n272 0.189894
R13527 commonsourceibias.n273 commonsourceibias.n251 0.189894
R13528 commonsourceibias.n278 commonsourceibias.n251 0.189894
R13529 commonsourceibias.n279 commonsourceibias.n278 0.189894
R13530 commonsourceibias.n280 commonsourceibias.n279 0.189894
R13531 commonsourceibias.n280 commonsourceibias.n249 0.189894
R13532 commonsourceibias.n286 commonsourceibias.n249 0.189894
R13533 commonsourceibias.n287 commonsourceibias.n286 0.189894
R13534 commonsourceibias.n288 commonsourceibias.n287 0.189894
R13535 commonsourceibias.n288 commonsourceibias.n247 0.189894
R13536 commonsourceibias.n293 commonsourceibias.n247 0.189894
R13537 commonsourceibias.n294 commonsourceibias.n293 0.189894
R13538 commonsourceibias.n295 commonsourceibias.n294 0.189894
R13539 commonsourceibias.n295 commonsourceibias.n245 0.189894
R13540 commonsourceibias.n300 commonsourceibias.n245 0.189894
R13541 commonsourceibias.n301 commonsourceibias.n300 0.189894
R13542 commonsourceibias.n301 commonsourceibias.n243 0.189894
R13543 commonsourceibias.n221 commonsourceibias.n216 0.189894
R13544 commonsourceibias.n222 commonsourceibias.n221 0.189894
R13545 commonsourceibias.n222 commonsourceibias.n214 0.189894
R13546 commonsourceibias.n226 commonsourceibias.n214 0.189894
R13547 commonsourceibias.n227 commonsourceibias.n226 0.189894
R13548 commonsourceibias.n227 commonsourceibias.n212 0.189894
R13549 commonsourceibias.n231 commonsourceibias.n212 0.189894
R13550 commonsourceibias.n232 commonsourceibias.n231 0.189894
R13551 commonsourceibias.n232 commonsourceibias.n210 0.189894
R13552 commonsourceibias.n237 commonsourceibias.n210 0.189894
R13553 commonsourceibias.n314 commonsourceibias.n208 0.189894
R13554 commonsourceibias.n320 commonsourceibias.n208 0.189894
R13555 commonsourceibias.n321 commonsourceibias.n320 0.189894
R13556 commonsourceibias.n322 commonsourceibias.n321 0.189894
R13557 commonsourceibias.n322 commonsourceibias.n206 0.189894
R13558 commonsourceibias.n327 commonsourceibias.n206 0.189894
R13559 commonsourceibias.n328 commonsourceibias.n327 0.189894
R13560 commonsourceibias.n329 commonsourceibias.n328 0.189894
R13561 commonsourceibias.n329 commonsourceibias.n204 0.189894
R13562 commonsourceibias.n334 commonsourceibias.n204 0.189894
R13563 commonsourceibias.n335 commonsourceibias.n334 0.189894
R13564 commonsourceibias.n335 commonsourceibias.n202 0.189894
R13565 commonsourceibias.n359 commonsourceibias.n354 0.189894
R13566 commonsourceibias.n360 commonsourceibias.n359 0.189894
R13567 commonsourceibias.n360 commonsourceibias.n352 0.189894
R13568 commonsourceibias.n364 commonsourceibias.n352 0.189894
R13569 commonsourceibias.n365 commonsourceibias.n364 0.189894
R13570 commonsourceibias.n365 commonsourceibias.n350 0.189894
R13571 commonsourceibias.n369 commonsourceibias.n350 0.189894
R13572 commonsourceibias.n370 commonsourceibias.n369 0.189894
R13573 commonsourceibias.n370 commonsourceibias.n348 0.189894
R13574 commonsourceibias.n375 commonsourceibias.n348 0.189894
R13575 commonsourceibias.n376 commonsourceibias.n375 0.189894
R13576 commonsourceibias.n377 commonsourceibias.n376 0.189894
R13577 commonsourceibias.n377 commonsourceibias.n346 0.189894
R13578 commonsourceibias.n383 commonsourceibias.n346 0.189894
R13579 commonsourceibias.n384 commonsourceibias.n383 0.189894
R13580 commonsourceibias.n385 commonsourceibias.n384 0.189894
R13581 commonsourceibias.n385 commonsourceibias.n344 0.189894
R13582 commonsourceibias.n390 commonsourceibias.n344 0.189894
R13583 commonsourceibias.n391 commonsourceibias.n390 0.189894
R13584 commonsourceibias.n392 commonsourceibias.n391 0.189894
R13585 commonsourceibias.n392 commonsourceibias.n342 0.189894
R13586 commonsourceibias.n397 commonsourceibias.n342 0.189894
R13587 commonsourceibias.n398 commonsourceibias.n397 0.189894
R13588 commonsourceibias.n398 commonsourceibias.n340 0.189894
R13589 commonsourceibias.n112 commonsourceibias.n111 0.170955
R13590 commonsourceibias.n113 commonsourceibias.n112 0.170955
R13591 commonsourceibias.n313 commonsourceibias.n237 0.170955
R13592 commonsourceibias.n314 commonsourceibias.n313 0.170955
R13593 CSoutput.n19 CSoutput.t189 184.661
R13594 CSoutput.n78 CSoutput.n77 165.8
R13595 CSoutput.n76 CSoutput.n0 165.8
R13596 CSoutput.n75 CSoutput.n74 165.8
R13597 CSoutput.n73 CSoutput.n72 165.8
R13598 CSoutput.n71 CSoutput.n2 165.8
R13599 CSoutput.n69 CSoutput.n68 165.8
R13600 CSoutput.n67 CSoutput.n3 165.8
R13601 CSoutput.n66 CSoutput.n65 165.8
R13602 CSoutput.n63 CSoutput.n4 165.8
R13603 CSoutput.n61 CSoutput.n60 165.8
R13604 CSoutput.n59 CSoutput.n5 165.8
R13605 CSoutput.n58 CSoutput.n57 165.8
R13606 CSoutput.n55 CSoutput.n6 165.8
R13607 CSoutput.n54 CSoutput.n53 165.8
R13608 CSoutput.n52 CSoutput.n51 165.8
R13609 CSoutput.n50 CSoutput.n8 165.8
R13610 CSoutput.n48 CSoutput.n47 165.8
R13611 CSoutput.n46 CSoutput.n9 165.8
R13612 CSoutput.n45 CSoutput.n44 165.8
R13613 CSoutput.n42 CSoutput.n10 165.8
R13614 CSoutput.n41 CSoutput.n40 165.8
R13615 CSoutput.n39 CSoutput.n38 165.8
R13616 CSoutput.n37 CSoutput.n12 165.8
R13617 CSoutput.n35 CSoutput.n34 165.8
R13618 CSoutput.n33 CSoutput.n13 165.8
R13619 CSoutput.n32 CSoutput.n31 165.8
R13620 CSoutput.n29 CSoutput.n14 165.8
R13621 CSoutput.n28 CSoutput.n27 165.8
R13622 CSoutput.n26 CSoutput.n25 165.8
R13623 CSoutput.n24 CSoutput.n16 165.8
R13624 CSoutput.n22 CSoutput.n21 165.8
R13625 CSoutput.n20 CSoutput.n17 165.8
R13626 CSoutput.n77 CSoutput.t168 162.194
R13627 CSoutput.n18 CSoutput.t169 120.501
R13628 CSoutput.n23 CSoutput.t179 120.501
R13629 CSoutput.n15 CSoutput.t175 120.501
R13630 CSoutput.n30 CSoutput.t171 120.501
R13631 CSoutput.n36 CSoutput.t182 120.501
R13632 CSoutput.n11 CSoutput.t184 120.501
R13633 CSoutput.n43 CSoutput.t173 120.501
R13634 CSoutput.n49 CSoutput.t185 120.501
R13635 CSoutput.n7 CSoutput.t186 120.501
R13636 CSoutput.n56 CSoutput.t180 120.501
R13637 CSoutput.n62 CSoutput.t172 120.501
R13638 CSoutput.n64 CSoutput.t188 120.501
R13639 CSoutput.n70 CSoutput.t183 120.501
R13640 CSoutput.n1 CSoutput.t178 120.501
R13641 CSoutput.n330 CSoutput.n328 103.469
R13642 CSoutput.n310 CSoutput.n308 103.469
R13643 CSoutput.n291 CSoutput.n289 103.469
R13644 CSoutput.n120 CSoutput.n118 103.469
R13645 CSoutput.n100 CSoutput.n98 103.469
R13646 CSoutput.n81 CSoutput.n79 103.469
R13647 CSoutput.n344 CSoutput.n343 103.111
R13648 CSoutput.n342 CSoutput.n341 103.111
R13649 CSoutput.n340 CSoutput.n339 103.111
R13650 CSoutput.n338 CSoutput.n337 103.111
R13651 CSoutput.n336 CSoutput.n335 103.111
R13652 CSoutput.n334 CSoutput.n333 103.111
R13653 CSoutput.n332 CSoutput.n331 103.111
R13654 CSoutput.n330 CSoutput.n329 103.111
R13655 CSoutput.n326 CSoutput.n325 103.111
R13656 CSoutput.n324 CSoutput.n323 103.111
R13657 CSoutput.n322 CSoutput.n321 103.111
R13658 CSoutput.n320 CSoutput.n319 103.111
R13659 CSoutput.n318 CSoutput.n317 103.111
R13660 CSoutput.n316 CSoutput.n315 103.111
R13661 CSoutput.n314 CSoutput.n313 103.111
R13662 CSoutput.n312 CSoutput.n311 103.111
R13663 CSoutput.n310 CSoutput.n309 103.111
R13664 CSoutput.n307 CSoutput.n306 103.111
R13665 CSoutput.n305 CSoutput.n304 103.111
R13666 CSoutput.n303 CSoutput.n302 103.111
R13667 CSoutput.n301 CSoutput.n300 103.111
R13668 CSoutput.n299 CSoutput.n298 103.111
R13669 CSoutput.n297 CSoutput.n296 103.111
R13670 CSoutput.n295 CSoutput.n294 103.111
R13671 CSoutput.n293 CSoutput.n292 103.111
R13672 CSoutput.n291 CSoutput.n290 103.111
R13673 CSoutput.n120 CSoutput.n119 103.111
R13674 CSoutput.n122 CSoutput.n121 103.111
R13675 CSoutput.n124 CSoutput.n123 103.111
R13676 CSoutput.n126 CSoutput.n125 103.111
R13677 CSoutput.n128 CSoutput.n127 103.111
R13678 CSoutput.n130 CSoutput.n129 103.111
R13679 CSoutput.n132 CSoutput.n131 103.111
R13680 CSoutput.n134 CSoutput.n133 103.111
R13681 CSoutput.n136 CSoutput.n135 103.111
R13682 CSoutput.n100 CSoutput.n99 103.111
R13683 CSoutput.n102 CSoutput.n101 103.111
R13684 CSoutput.n104 CSoutput.n103 103.111
R13685 CSoutput.n106 CSoutput.n105 103.111
R13686 CSoutput.n108 CSoutput.n107 103.111
R13687 CSoutput.n110 CSoutput.n109 103.111
R13688 CSoutput.n112 CSoutput.n111 103.111
R13689 CSoutput.n114 CSoutput.n113 103.111
R13690 CSoutput.n116 CSoutput.n115 103.111
R13691 CSoutput.n81 CSoutput.n80 103.111
R13692 CSoutput.n83 CSoutput.n82 103.111
R13693 CSoutput.n85 CSoutput.n84 103.111
R13694 CSoutput.n87 CSoutput.n86 103.111
R13695 CSoutput.n89 CSoutput.n88 103.111
R13696 CSoutput.n91 CSoutput.n90 103.111
R13697 CSoutput.n93 CSoutput.n92 103.111
R13698 CSoutput.n95 CSoutput.n94 103.111
R13699 CSoutput.n97 CSoutput.n96 103.111
R13700 CSoutput.n346 CSoutput.n345 103.111
R13701 CSoutput.n362 CSoutput.n360 81.5057
R13702 CSoutput.n351 CSoutput.n349 81.5057
R13703 CSoutput.n386 CSoutput.n384 81.5057
R13704 CSoutput.n375 CSoutput.n373 81.5057
R13705 CSoutput.n370 CSoutput.n369 80.9324
R13706 CSoutput.n368 CSoutput.n367 80.9324
R13707 CSoutput.n366 CSoutput.n365 80.9324
R13708 CSoutput.n364 CSoutput.n363 80.9324
R13709 CSoutput.n362 CSoutput.n361 80.9324
R13710 CSoutput.n359 CSoutput.n358 80.9324
R13711 CSoutput.n357 CSoutput.n356 80.9324
R13712 CSoutput.n355 CSoutput.n354 80.9324
R13713 CSoutput.n353 CSoutput.n352 80.9324
R13714 CSoutput.n351 CSoutput.n350 80.9324
R13715 CSoutput.n386 CSoutput.n385 80.9324
R13716 CSoutput.n388 CSoutput.n387 80.9324
R13717 CSoutput.n390 CSoutput.n389 80.9324
R13718 CSoutput.n392 CSoutput.n391 80.9324
R13719 CSoutput.n394 CSoutput.n393 80.9324
R13720 CSoutput.n375 CSoutput.n374 80.9324
R13721 CSoutput.n377 CSoutput.n376 80.9324
R13722 CSoutput.n379 CSoutput.n378 80.9324
R13723 CSoutput.n381 CSoutput.n380 80.9324
R13724 CSoutput.n383 CSoutput.n382 80.9324
R13725 CSoutput.n25 CSoutput.n24 48.1486
R13726 CSoutput.n69 CSoutput.n3 48.1486
R13727 CSoutput.n38 CSoutput.n37 48.1486
R13728 CSoutput.n42 CSoutput.n41 48.1486
R13729 CSoutput.n51 CSoutput.n50 48.1486
R13730 CSoutput.n55 CSoutput.n54 48.1486
R13731 CSoutput.n22 CSoutput.n17 46.462
R13732 CSoutput.n72 CSoutput.n71 46.462
R13733 CSoutput.n20 CSoutput.n19 44.9055
R13734 CSoutput.n29 CSoutput.n28 43.7635
R13735 CSoutput.n65 CSoutput.n63 43.7635
R13736 CSoutput.n35 CSoutput.n13 41.7396
R13737 CSoutput.n57 CSoutput.n5 41.7396
R13738 CSoutput.n44 CSoutput.n9 37.0171
R13739 CSoutput.n48 CSoutput.n9 37.0171
R13740 CSoutput.n76 CSoutput.n75 34.9932
R13741 CSoutput.n31 CSoutput.n13 32.2947
R13742 CSoutput.n61 CSoutput.n5 32.2947
R13743 CSoutput.n30 CSoutput.n29 29.6014
R13744 CSoutput.n63 CSoutput.n62 29.6014
R13745 CSoutput.n19 CSoutput.n18 28.4085
R13746 CSoutput.n18 CSoutput.n17 25.1176
R13747 CSoutput.n72 CSoutput.n1 25.1176
R13748 CSoutput.n43 CSoutput.n42 22.0922
R13749 CSoutput.n50 CSoutput.n49 22.0922
R13750 CSoutput.n77 CSoutput.n76 21.8586
R13751 CSoutput.n37 CSoutput.n36 18.9681
R13752 CSoutput.n56 CSoutput.n55 18.9681
R13753 CSoutput.n25 CSoutput.n15 17.6292
R13754 CSoutput.n64 CSoutput.n3 17.6292
R13755 CSoutput.n24 CSoutput.n23 15.844
R13756 CSoutput.n70 CSoutput.n69 15.844
R13757 CSoutput.n38 CSoutput.n11 14.5051
R13758 CSoutput.n54 CSoutput.n7 14.5051
R13759 CSoutput.n397 CSoutput.n78 11.6139
R13760 CSoutput.n41 CSoutput.n11 11.3811
R13761 CSoutput.n51 CSoutput.n7 11.3811
R13762 CSoutput.n23 CSoutput.n22 10.0422
R13763 CSoutput.n71 CSoutput.n70 10.0422
R13764 CSoutput.n327 CSoutput.n307 9.25285
R13765 CSoutput.n117 CSoutput.n97 9.25285
R13766 CSoutput.n371 CSoutput.n359 8.97993
R13767 CSoutput.n395 CSoutput.n383 8.97993
R13768 CSoutput.n372 CSoutput.n348 8.61621
R13769 CSoutput.n28 CSoutput.n15 8.25698
R13770 CSoutput.n65 CSoutput.n64 8.25698
R13771 CSoutput.n372 CSoutput.n371 7.89345
R13772 CSoutput.n396 CSoutput.n395 7.89345
R13773 CSoutput.n348 CSoutput.n347 7.12641
R13774 CSoutput.n138 CSoutput.n137 7.12641
R13775 CSoutput.n36 CSoutput.n35 6.91809
R13776 CSoutput.n57 CSoutput.n56 6.91809
R13777 CSoutput.n371 CSoutput.n370 5.25266
R13778 CSoutput.n395 CSoutput.n394 5.25266
R13779 CSoutput.n347 CSoutput.n346 5.1449
R13780 CSoutput.n327 CSoutput.n326 5.1449
R13781 CSoutput.n137 CSoutput.n136 5.1449
R13782 CSoutput.n117 CSoutput.n116 5.1449
R13783 CSoutput.n397 CSoutput.n138 5.02377
R13784 CSoutput.n229 CSoutput.n182 4.5005
R13785 CSoutput.n198 CSoutput.n182 4.5005
R13786 CSoutput.n193 CSoutput.n177 4.5005
R13787 CSoutput.n193 CSoutput.n179 4.5005
R13788 CSoutput.n193 CSoutput.n176 4.5005
R13789 CSoutput.n193 CSoutput.n180 4.5005
R13790 CSoutput.n193 CSoutput.n175 4.5005
R13791 CSoutput.n193 CSoutput.t174 4.5005
R13792 CSoutput.n193 CSoutput.n174 4.5005
R13793 CSoutput.n193 CSoutput.n181 4.5005
R13794 CSoutput.n193 CSoutput.n182 4.5005
R13795 CSoutput.n191 CSoutput.n177 4.5005
R13796 CSoutput.n191 CSoutput.n179 4.5005
R13797 CSoutput.n191 CSoutput.n176 4.5005
R13798 CSoutput.n191 CSoutput.n180 4.5005
R13799 CSoutput.n191 CSoutput.n175 4.5005
R13800 CSoutput.n191 CSoutput.t174 4.5005
R13801 CSoutput.n191 CSoutput.n174 4.5005
R13802 CSoutput.n191 CSoutput.n181 4.5005
R13803 CSoutput.n191 CSoutput.n182 4.5005
R13804 CSoutput.n190 CSoutput.n177 4.5005
R13805 CSoutput.n190 CSoutput.n179 4.5005
R13806 CSoutput.n190 CSoutput.n176 4.5005
R13807 CSoutput.n190 CSoutput.n180 4.5005
R13808 CSoutput.n190 CSoutput.n175 4.5005
R13809 CSoutput.n190 CSoutput.t174 4.5005
R13810 CSoutput.n190 CSoutput.n174 4.5005
R13811 CSoutput.n190 CSoutput.n181 4.5005
R13812 CSoutput.n190 CSoutput.n182 4.5005
R13813 CSoutput.n275 CSoutput.n177 4.5005
R13814 CSoutput.n275 CSoutput.n179 4.5005
R13815 CSoutput.n275 CSoutput.n176 4.5005
R13816 CSoutput.n275 CSoutput.n180 4.5005
R13817 CSoutput.n275 CSoutput.n175 4.5005
R13818 CSoutput.n275 CSoutput.t174 4.5005
R13819 CSoutput.n275 CSoutput.n174 4.5005
R13820 CSoutput.n275 CSoutput.n181 4.5005
R13821 CSoutput.n275 CSoutput.n182 4.5005
R13822 CSoutput.n273 CSoutput.n177 4.5005
R13823 CSoutput.n273 CSoutput.n179 4.5005
R13824 CSoutput.n273 CSoutput.n176 4.5005
R13825 CSoutput.n273 CSoutput.n180 4.5005
R13826 CSoutput.n273 CSoutput.n175 4.5005
R13827 CSoutput.n273 CSoutput.t174 4.5005
R13828 CSoutput.n273 CSoutput.n174 4.5005
R13829 CSoutput.n273 CSoutput.n181 4.5005
R13830 CSoutput.n271 CSoutput.n177 4.5005
R13831 CSoutput.n271 CSoutput.n179 4.5005
R13832 CSoutput.n271 CSoutput.n176 4.5005
R13833 CSoutput.n271 CSoutput.n180 4.5005
R13834 CSoutput.n271 CSoutput.n175 4.5005
R13835 CSoutput.n271 CSoutput.t174 4.5005
R13836 CSoutput.n271 CSoutput.n174 4.5005
R13837 CSoutput.n271 CSoutput.n181 4.5005
R13838 CSoutput.n201 CSoutput.n177 4.5005
R13839 CSoutput.n201 CSoutput.n179 4.5005
R13840 CSoutput.n201 CSoutput.n176 4.5005
R13841 CSoutput.n201 CSoutput.n180 4.5005
R13842 CSoutput.n201 CSoutput.n175 4.5005
R13843 CSoutput.n201 CSoutput.t174 4.5005
R13844 CSoutput.n201 CSoutput.n174 4.5005
R13845 CSoutput.n201 CSoutput.n181 4.5005
R13846 CSoutput.n201 CSoutput.n182 4.5005
R13847 CSoutput.n200 CSoutput.n177 4.5005
R13848 CSoutput.n200 CSoutput.n179 4.5005
R13849 CSoutput.n200 CSoutput.n176 4.5005
R13850 CSoutput.n200 CSoutput.n180 4.5005
R13851 CSoutput.n200 CSoutput.n175 4.5005
R13852 CSoutput.n200 CSoutput.t174 4.5005
R13853 CSoutput.n200 CSoutput.n174 4.5005
R13854 CSoutput.n200 CSoutput.n181 4.5005
R13855 CSoutput.n200 CSoutput.n182 4.5005
R13856 CSoutput.n204 CSoutput.n177 4.5005
R13857 CSoutput.n204 CSoutput.n179 4.5005
R13858 CSoutput.n204 CSoutput.n176 4.5005
R13859 CSoutput.n204 CSoutput.n180 4.5005
R13860 CSoutput.n204 CSoutput.n175 4.5005
R13861 CSoutput.n204 CSoutput.t174 4.5005
R13862 CSoutput.n204 CSoutput.n174 4.5005
R13863 CSoutput.n204 CSoutput.n181 4.5005
R13864 CSoutput.n204 CSoutput.n182 4.5005
R13865 CSoutput.n203 CSoutput.n177 4.5005
R13866 CSoutput.n203 CSoutput.n179 4.5005
R13867 CSoutput.n203 CSoutput.n176 4.5005
R13868 CSoutput.n203 CSoutput.n180 4.5005
R13869 CSoutput.n203 CSoutput.n175 4.5005
R13870 CSoutput.n203 CSoutput.t174 4.5005
R13871 CSoutput.n203 CSoutput.n174 4.5005
R13872 CSoutput.n203 CSoutput.n181 4.5005
R13873 CSoutput.n203 CSoutput.n182 4.5005
R13874 CSoutput.n186 CSoutput.n177 4.5005
R13875 CSoutput.n186 CSoutput.n179 4.5005
R13876 CSoutput.n186 CSoutput.n176 4.5005
R13877 CSoutput.n186 CSoutput.n180 4.5005
R13878 CSoutput.n186 CSoutput.n175 4.5005
R13879 CSoutput.n186 CSoutput.t174 4.5005
R13880 CSoutput.n186 CSoutput.n174 4.5005
R13881 CSoutput.n186 CSoutput.n181 4.5005
R13882 CSoutput.n186 CSoutput.n182 4.5005
R13883 CSoutput.n278 CSoutput.n177 4.5005
R13884 CSoutput.n278 CSoutput.n179 4.5005
R13885 CSoutput.n278 CSoutput.n176 4.5005
R13886 CSoutput.n278 CSoutput.n180 4.5005
R13887 CSoutput.n278 CSoutput.n175 4.5005
R13888 CSoutput.n278 CSoutput.t174 4.5005
R13889 CSoutput.n278 CSoutput.n174 4.5005
R13890 CSoutput.n278 CSoutput.n181 4.5005
R13891 CSoutput.n278 CSoutput.n182 4.5005
R13892 CSoutput.n265 CSoutput.n236 4.5005
R13893 CSoutput.n265 CSoutput.n242 4.5005
R13894 CSoutput.n223 CSoutput.n212 4.5005
R13895 CSoutput.n223 CSoutput.n214 4.5005
R13896 CSoutput.n223 CSoutput.n211 4.5005
R13897 CSoutput.n223 CSoutput.n215 4.5005
R13898 CSoutput.n223 CSoutput.n210 4.5005
R13899 CSoutput.n223 CSoutput.t170 4.5005
R13900 CSoutput.n223 CSoutput.n209 4.5005
R13901 CSoutput.n223 CSoutput.n216 4.5005
R13902 CSoutput.n265 CSoutput.n223 4.5005
R13903 CSoutput.n244 CSoutput.n212 4.5005
R13904 CSoutput.n244 CSoutput.n214 4.5005
R13905 CSoutput.n244 CSoutput.n211 4.5005
R13906 CSoutput.n244 CSoutput.n215 4.5005
R13907 CSoutput.n244 CSoutput.n210 4.5005
R13908 CSoutput.n244 CSoutput.t170 4.5005
R13909 CSoutput.n244 CSoutput.n209 4.5005
R13910 CSoutput.n244 CSoutput.n216 4.5005
R13911 CSoutput.n265 CSoutput.n244 4.5005
R13912 CSoutput.n222 CSoutput.n212 4.5005
R13913 CSoutput.n222 CSoutput.n214 4.5005
R13914 CSoutput.n222 CSoutput.n211 4.5005
R13915 CSoutput.n222 CSoutput.n215 4.5005
R13916 CSoutput.n222 CSoutput.n210 4.5005
R13917 CSoutput.n222 CSoutput.t170 4.5005
R13918 CSoutput.n222 CSoutput.n209 4.5005
R13919 CSoutput.n222 CSoutput.n216 4.5005
R13920 CSoutput.n265 CSoutput.n222 4.5005
R13921 CSoutput.n246 CSoutput.n212 4.5005
R13922 CSoutput.n246 CSoutput.n214 4.5005
R13923 CSoutput.n246 CSoutput.n211 4.5005
R13924 CSoutput.n246 CSoutput.n215 4.5005
R13925 CSoutput.n246 CSoutput.n210 4.5005
R13926 CSoutput.n246 CSoutput.t170 4.5005
R13927 CSoutput.n246 CSoutput.n209 4.5005
R13928 CSoutput.n246 CSoutput.n216 4.5005
R13929 CSoutput.n265 CSoutput.n246 4.5005
R13930 CSoutput.n212 CSoutput.n207 4.5005
R13931 CSoutput.n214 CSoutput.n207 4.5005
R13932 CSoutput.n211 CSoutput.n207 4.5005
R13933 CSoutput.n215 CSoutput.n207 4.5005
R13934 CSoutput.n210 CSoutput.n207 4.5005
R13935 CSoutput.t170 CSoutput.n207 4.5005
R13936 CSoutput.n209 CSoutput.n207 4.5005
R13937 CSoutput.n216 CSoutput.n207 4.5005
R13938 CSoutput.n268 CSoutput.n212 4.5005
R13939 CSoutput.n268 CSoutput.n214 4.5005
R13940 CSoutput.n268 CSoutput.n211 4.5005
R13941 CSoutput.n268 CSoutput.n215 4.5005
R13942 CSoutput.n268 CSoutput.n210 4.5005
R13943 CSoutput.n268 CSoutput.t170 4.5005
R13944 CSoutput.n268 CSoutput.n209 4.5005
R13945 CSoutput.n268 CSoutput.n216 4.5005
R13946 CSoutput.n266 CSoutput.n212 4.5005
R13947 CSoutput.n266 CSoutput.n214 4.5005
R13948 CSoutput.n266 CSoutput.n211 4.5005
R13949 CSoutput.n266 CSoutput.n215 4.5005
R13950 CSoutput.n266 CSoutput.n210 4.5005
R13951 CSoutput.n266 CSoutput.t170 4.5005
R13952 CSoutput.n266 CSoutput.n209 4.5005
R13953 CSoutput.n266 CSoutput.n216 4.5005
R13954 CSoutput.n266 CSoutput.n265 4.5005
R13955 CSoutput.n248 CSoutput.n212 4.5005
R13956 CSoutput.n248 CSoutput.n214 4.5005
R13957 CSoutput.n248 CSoutput.n211 4.5005
R13958 CSoutput.n248 CSoutput.n215 4.5005
R13959 CSoutput.n248 CSoutput.n210 4.5005
R13960 CSoutput.n248 CSoutput.t170 4.5005
R13961 CSoutput.n248 CSoutput.n209 4.5005
R13962 CSoutput.n248 CSoutput.n216 4.5005
R13963 CSoutput.n265 CSoutput.n248 4.5005
R13964 CSoutput.n220 CSoutput.n212 4.5005
R13965 CSoutput.n220 CSoutput.n214 4.5005
R13966 CSoutput.n220 CSoutput.n211 4.5005
R13967 CSoutput.n220 CSoutput.n215 4.5005
R13968 CSoutput.n220 CSoutput.n210 4.5005
R13969 CSoutput.n220 CSoutput.t170 4.5005
R13970 CSoutput.n220 CSoutput.n209 4.5005
R13971 CSoutput.n220 CSoutput.n216 4.5005
R13972 CSoutput.n265 CSoutput.n220 4.5005
R13973 CSoutput.n250 CSoutput.n212 4.5005
R13974 CSoutput.n250 CSoutput.n214 4.5005
R13975 CSoutput.n250 CSoutput.n211 4.5005
R13976 CSoutput.n250 CSoutput.n215 4.5005
R13977 CSoutput.n250 CSoutput.n210 4.5005
R13978 CSoutput.n250 CSoutput.t170 4.5005
R13979 CSoutput.n250 CSoutput.n209 4.5005
R13980 CSoutput.n250 CSoutput.n216 4.5005
R13981 CSoutput.n265 CSoutput.n250 4.5005
R13982 CSoutput.n219 CSoutput.n212 4.5005
R13983 CSoutput.n219 CSoutput.n214 4.5005
R13984 CSoutput.n219 CSoutput.n211 4.5005
R13985 CSoutput.n219 CSoutput.n215 4.5005
R13986 CSoutput.n219 CSoutput.n210 4.5005
R13987 CSoutput.n219 CSoutput.t170 4.5005
R13988 CSoutput.n219 CSoutput.n209 4.5005
R13989 CSoutput.n219 CSoutput.n216 4.5005
R13990 CSoutput.n265 CSoutput.n219 4.5005
R13991 CSoutput.n264 CSoutput.n212 4.5005
R13992 CSoutput.n264 CSoutput.n214 4.5005
R13993 CSoutput.n264 CSoutput.n211 4.5005
R13994 CSoutput.n264 CSoutput.n215 4.5005
R13995 CSoutput.n264 CSoutput.n210 4.5005
R13996 CSoutput.n264 CSoutput.t170 4.5005
R13997 CSoutput.n264 CSoutput.n209 4.5005
R13998 CSoutput.n264 CSoutput.n216 4.5005
R13999 CSoutput.n265 CSoutput.n264 4.5005
R14000 CSoutput.n263 CSoutput.n148 4.5005
R14001 CSoutput.n164 CSoutput.n148 4.5005
R14002 CSoutput.n159 CSoutput.n143 4.5005
R14003 CSoutput.n159 CSoutput.n145 4.5005
R14004 CSoutput.n159 CSoutput.n142 4.5005
R14005 CSoutput.n159 CSoutput.n146 4.5005
R14006 CSoutput.n159 CSoutput.n141 4.5005
R14007 CSoutput.n159 CSoutput.t187 4.5005
R14008 CSoutput.n159 CSoutput.n140 4.5005
R14009 CSoutput.n159 CSoutput.n147 4.5005
R14010 CSoutput.n159 CSoutput.n148 4.5005
R14011 CSoutput.n157 CSoutput.n143 4.5005
R14012 CSoutput.n157 CSoutput.n145 4.5005
R14013 CSoutput.n157 CSoutput.n142 4.5005
R14014 CSoutput.n157 CSoutput.n146 4.5005
R14015 CSoutput.n157 CSoutput.n141 4.5005
R14016 CSoutput.n157 CSoutput.t187 4.5005
R14017 CSoutput.n157 CSoutput.n140 4.5005
R14018 CSoutput.n157 CSoutput.n147 4.5005
R14019 CSoutput.n157 CSoutput.n148 4.5005
R14020 CSoutput.n156 CSoutput.n143 4.5005
R14021 CSoutput.n156 CSoutput.n145 4.5005
R14022 CSoutput.n156 CSoutput.n142 4.5005
R14023 CSoutput.n156 CSoutput.n146 4.5005
R14024 CSoutput.n156 CSoutput.n141 4.5005
R14025 CSoutput.n156 CSoutput.t187 4.5005
R14026 CSoutput.n156 CSoutput.n140 4.5005
R14027 CSoutput.n156 CSoutput.n147 4.5005
R14028 CSoutput.n156 CSoutput.n148 4.5005
R14029 CSoutput.n285 CSoutput.n143 4.5005
R14030 CSoutput.n285 CSoutput.n145 4.5005
R14031 CSoutput.n285 CSoutput.n142 4.5005
R14032 CSoutput.n285 CSoutput.n146 4.5005
R14033 CSoutput.n285 CSoutput.n141 4.5005
R14034 CSoutput.n285 CSoutput.t187 4.5005
R14035 CSoutput.n285 CSoutput.n140 4.5005
R14036 CSoutput.n285 CSoutput.n147 4.5005
R14037 CSoutput.n285 CSoutput.n148 4.5005
R14038 CSoutput.n283 CSoutput.n143 4.5005
R14039 CSoutput.n283 CSoutput.n145 4.5005
R14040 CSoutput.n283 CSoutput.n142 4.5005
R14041 CSoutput.n283 CSoutput.n146 4.5005
R14042 CSoutput.n283 CSoutput.n141 4.5005
R14043 CSoutput.n283 CSoutput.t187 4.5005
R14044 CSoutput.n283 CSoutput.n140 4.5005
R14045 CSoutput.n283 CSoutput.n147 4.5005
R14046 CSoutput.n281 CSoutput.n143 4.5005
R14047 CSoutput.n281 CSoutput.n145 4.5005
R14048 CSoutput.n281 CSoutput.n142 4.5005
R14049 CSoutput.n281 CSoutput.n146 4.5005
R14050 CSoutput.n281 CSoutput.n141 4.5005
R14051 CSoutput.n281 CSoutput.t187 4.5005
R14052 CSoutput.n281 CSoutput.n140 4.5005
R14053 CSoutput.n281 CSoutput.n147 4.5005
R14054 CSoutput.n167 CSoutput.n143 4.5005
R14055 CSoutput.n167 CSoutput.n145 4.5005
R14056 CSoutput.n167 CSoutput.n142 4.5005
R14057 CSoutput.n167 CSoutput.n146 4.5005
R14058 CSoutput.n167 CSoutput.n141 4.5005
R14059 CSoutput.n167 CSoutput.t187 4.5005
R14060 CSoutput.n167 CSoutput.n140 4.5005
R14061 CSoutput.n167 CSoutput.n147 4.5005
R14062 CSoutput.n167 CSoutput.n148 4.5005
R14063 CSoutput.n166 CSoutput.n143 4.5005
R14064 CSoutput.n166 CSoutput.n145 4.5005
R14065 CSoutput.n166 CSoutput.n142 4.5005
R14066 CSoutput.n166 CSoutput.n146 4.5005
R14067 CSoutput.n166 CSoutput.n141 4.5005
R14068 CSoutput.n166 CSoutput.t187 4.5005
R14069 CSoutput.n166 CSoutput.n140 4.5005
R14070 CSoutput.n166 CSoutput.n147 4.5005
R14071 CSoutput.n166 CSoutput.n148 4.5005
R14072 CSoutput.n170 CSoutput.n143 4.5005
R14073 CSoutput.n170 CSoutput.n145 4.5005
R14074 CSoutput.n170 CSoutput.n142 4.5005
R14075 CSoutput.n170 CSoutput.n146 4.5005
R14076 CSoutput.n170 CSoutput.n141 4.5005
R14077 CSoutput.n170 CSoutput.t187 4.5005
R14078 CSoutput.n170 CSoutput.n140 4.5005
R14079 CSoutput.n170 CSoutput.n147 4.5005
R14080 CSoutput.n170 CSoutput.n148 4.5005
R14081 CSoutput.n169 CSoutput.n143 4.5005
R14082 CSoutput.n169 CSoutput.n145 4.5005
R14083 CSoutput.n169 CSoutput.n142 4.5005
R14084 CSoutput.n169 CSoutput.n146 4.5005
R14085 CSoutput.n169 CSoutput.n141 4.5005
R14086 CSoutput.n169 CSoutput.t187 4.5005
R14087 CSoutput.n169 CSoutput.n140 4.5005
R14088 CSoutput.n169 CSoutput.n147 4.5005
R14089 CSoutput.n169 CSoutput.n148 4.5005
R14090 CSoutput.n152 CSoutput.n143 4.5005
R14091 CSoutput.n152 CSoutput.n145 4.5005
R14092 CSoutput.n152 CSoutput.n142 4.5005
R14093 CSoutput.n152 CSoutput.n146 4.5005
R14094 CSoutput.n152 CSoutput.n141 4.5005
R14095 CSoutput.n152 CSoutput.t187 4.5005
R14096 CSoutput.n152 CSoutput.n140 4.5005
R14097 CSoutput.n152 CSoutput.n147 4.5005
R14098 CSoutput.n152 CSoutput.n148 4.5005
R14099 CSoutput.n288 CSoutput.n143 4.5005
R14100 CSoutput.n288 CSoutput.n145 4.5005
R14101 CSoutput.n288 CSoutput.n142 4.5005
R14102 CSoutput.n288 CSoutput.n146 4.5005
R14103 CSoutput.n288 CSoutput.n141 4.5005
R14104 CSoutput.n288 CSoutput.t187 4.5005
R14105 CSoutput.n288 CSoutput.n140 4.5005
R14106 CSoutput.n288 CSoutput.n147 4.5005
R14107 CSoutput.n288 CSoutput.n148 4.5005
R14108 CSoutput.n347 CSoutput.n327 4.10845
R14109 CSoutput.n137 CSoutput.n117 4.10845
R14110 CSoutput.n345 CSoutput.t116 4.06363
R14111 CSoutput.n345 CSoutput.t131 4.06363
R14112 CSoutput.n343 CSoutput.t130 4.06363
R14113 CSoutput.n343 CSoutput.t3 4.06363
R14114 CSoutput.n341 CSoutput.t99 4.06363
R14115 CSoutput.n341 CSoutput.t163 4.06363
R14116 CSoutput.n339 CSoutput.t110 4.06363
R14117 CSoutput.n339 CSoutput.t120 4.06363
R14118 CSoutput.n337 CSoutput.t140 4.06363
R14119 CSoutput.n337 CSoutput.t153 4.06363
R14120 CSoutput.n335 CSoutput.t108 4.06363
R14121 CSoutput.n335 CSoutput.t154 4.06363
R14122 CSoutput.n333 CSoutput.t75 4.06363
R14123 CSoutput.n333 CSoutput.t142 4.06363
R14124 CSoutput.n331 CSoutput.t117 4.06363
R14125 CSoutput.n331 CSoutput.t136 4.06363
R14126 CSoutput.n329 CSoutput.t162 4.06363
R14127 CSoutput.n329 CSoutput.t91 4.06363
R14128 CSoutput.n328 CSoutput.t5 4.06363
R14129 CSoutput.n328 CSoutput.t109 4.06363
R14130 CSoutput.n325 CSoutput.t155 4.06363
R14131 CSoutput.n325 CSoutput.t103 4.06363
R14132 CSoutput.n323 CSoutput.t101 4.06363
R14133 CSoutput.n323 CSoutput.t164 4.06363
R14134 CSoutput.n321 CSoutput.t74 4.06363
R14135 CSoutput.n321 CSoutput.t73 4.06363
R14136 CSoutput.n319 CSoutput.t150 4.06363
R14137 CSoutput.n319 CSoutput.t89 4.06363
R14138 CSoutput.n317 CSoutput.t94 4.06363
R14139 CSoutput.n317 CSoutput.t77 4.06363
R14140 CSoutput.n315 CSoutput.t95 4.06363
R14141 CSoutput.n315 CSoutput.t60 4.06363
R14142 CSoutput.n313 CSoutput.t111 4.06363
R14143 CSoutput.n313 CSoutput.t113 4.06363
R14144 CSoutput.n311 CSoutput.t64 4.06363
R14145 CSoutput.n311 CSoutput.t128 4.06363
R14146 CSoutput.n309 CSoutput.t126 4.06363
R14147 CSoutput.n309 CSoutput.t8 4.06363
R14148 CSoutput.n308 CSoutput.t149 4.06363
R14149 CSoutput.n308 CSoutput.t62 4.06363
R14150 CSoutput.n306 CSoutput.t123 4.06363
R14151 CSoutput.n306 CSoutput.t165 4.06363
R14152 CSoutput.n304 CSoutput.t106 4.06363
R14153 CSoutput.n304 CSoutput.t160 4.06363
R14154 CSoutput.n302 CSoutput.t97 4.06363
R14155 CSoutput.n302 CSoutput.t90 4.06363
R14156 CSoutput.n300 CSoutput.t100 4.06363
R14157 CSoutput.n300 CSoutput.t86 4.06363
R14158 CSoutput.n298 CSoutput.t167 4.06363
R14159 CSoutput.n298 CSoutput.t93 4.06363
R14160 CSoutput.n296 CSoutput.t7 4.06363
R14161 CSoutput.n296 CSoutput.t72 4.06363
R14162 CSoutput.n294 CSoutput.t66 4.06363
R14163 CSoutput.n294 CSoutput.t145 4.06363
R14164 CSoutput.n292 CSoutput.t96 4.06363
R14165 CSoutput.n292 CSoutput.t135 4.06363
R14166 CSoutput.n290 CSoutput.t69 4.06363
R14167 CSoutput.n290 CSoutput.t65 4.06363
R14168 CSoutput.n289 CSoutput.t104 4.06363
R14169 CSoutput.n289 CSoutput.t152 4.06363
R14170 CSoutput.n118 CSoutput.t102 4.06363
R14171 CSoutput.n118 CSoutput.t151 4.06363
R14172 CSoutput.n119 CSoutput.t137 4.06363
R14173 CSoutput.n119 CSoutput.t84 4.06363
R14174 CSoutput.n121 CSoutput.t139 4.06363
R14175 CSoutput.n121 CSoutput.t68 4.06363
R14176 CSoutput.n123 CSoutput.t6 4.06363
R14177 CSoutput.n123 CSoutput.t1 4.06363
R14178 CSoutput.n125 CSoutput.t144 4.06363
R14179 CSoutput.n125 CSoutput.t83 4.06363
R14180 CSoutput.n127 CSoutput.t138 4.06363
R14181 CSoutput.n127 CSoutput.t129 4.06363
R14182 CSoutput.n129 CSoutput.t119 4.06363
R14183 CSoutput.n129 CSoutput.t63 4.06363
R14184 CSoutput.n131 CSoutput.t76 4.06363
R14185 CSoutput.n131 CSoutput.t81 4.06363
R14186 CSoutput.n133 CSoutput.t118 4.06363
R14187 CSoutput.n133 CSoutput.t122 4.06363
R14188 CSoutput.n135 CSoutput.t159 4.06363
R14189 CSoutput.n135 CSoutput.t85 4.06363
R14190 CSoutput.n98 CSoutput.t87 4.06363
R14191 CSoutput.n98 CSoutput.t92 4.06363
R14192 CSoutput.n99 CSoutput.t134 4.06363
R14193 CSoutput.n99 CSoutput.t9 4.06363
R14194 CSoutput.n101 CSoutput.t88 4.06363
R14195 CSoutput.n101 CSoutput.t115 4.06363
R14196 CSoutput.n103 CSoutput.t10 4.06363
R14197 CSoutput.n103 CSoutput.t147 4.06363
R14198 CSoutput.n105 CSoutput.t67 4.06363
R14199 CSoutput.n105 CSoutput.t141 4.06363
R14200 CSoutput.n107 CSoutput.t61 4.06363
R14201 CSoutput.n107 CSoutput.t59 4.06363
R14202 CSoutput.n109 CSoutput.t146 4.06363
R14203 CSoutput.n109 CSoutput.t78 4.06363
R14204 CSoutput.n111 CSoutput.t157 4.06363
R14205 CSoutput.n111 CSoutput.t148 4.06363
R14206 CSoutput.n113 CSoutput.t70 4.06363
R14207 CSoutput.n113 CSoutput.t105 4.06363
R14208 CSoutput.n115 CSoutput.t166 4.06363
R14209 CSoutput.n115 CSoutput.t125 4.06363
R14210 CSoutput.n79 CSoutput.t71 4.06363
R14211 CSoutput.n79 CSoutput.t98 4.06363
R14212 CSoutput.n80 CSoutput.t161 4.06363
R14213 CSoutput.n80 CSoutput.t158 4.06363
R14214 CSoutput.n82 CSoutput.t0 4.06363
R14215 CSoutput.n82 CSoutput.t2 4.06363
R14216 CSoutput.n84 CSoutput.t132 4.06363
R14217 CSoutput.n84 CSoutput.t80 4.06363
R14218 CSoutput.n86 CSoutput.t127 4.06363
R14219 CSoutput.n86 CSoutput.t133 4.06363
R14220 CSoutput.n88 CSoutput.t156 4.06363
R14221 CSoutput.n88 CSoutput.t112 4.06363
R14222 CSoutput.n90 CSoutput.t82 4.06363
R14223 CSoutput.n90 CSoutput.t143 4.06363
R14224 CSoutput.n92 CSoutput.t114 4.06363
R14225 CSoutput.n92 CSoutput.t107 4.06363
R14226 CSoutput.n94 CSoutput.t124 4.06363
R14227 CSoutput.n94 CSoutput.t4 4.06363
R14228 CSoutput.n96 CSoutput.t79 4.06363
R14229 CSoutput.n96 CSoutput.t121 4.06363
R14230 CSoutput.n44 CSoutput.n43 3.79402
R14231 CSoutput.n49 CSoutput.n48 3.79402
R14232 CSoutput.n397 CSoutput.n396 3.57343
R14233 CSoutput.n369 CSoutput.t49 2.82907
R14234 CSoutput.n369 CSoutput.t52 2.82907
R14235 CSoutput.n367 CSoutput.t48 2.82907
R14236 CSoutput.n367 CSoutput.t38 2.82907
R14237 CSoutput.n365 CSoutput.t15 2.82907
R14238 CSoutput.n365 CSoutput.t46 2.82907
R14239 CSoutput.n363 CSoutput.t40 2.82907
R14240 CSoutput.n363 CSoutput.t29 2.82907
R14241 CSoutput.n361 CSoutput.t57 2.82907
R14242 CSoutput.n361 CSoutput.t11 2.82907
R14243 CSoutput.n360 CSoutput.t45 2.82907
R14244 CSoutput.n360 CSoutput.t34 2.82907
R14245 CSoutput.n358 CSoutput.t42 2.82907
R14246 CSoutput.n358 CSoutput.t44 2.82907
R14247 CSoutput.n356 CSoutput.t39 2.82907
R14248 CSoutput.n356 CSoutput.t28 2.82907
R14249 CSoutput.n354 CSoutput.t56 2.82907
R14250 CSoutput.n354 CSoutput.t37 2.82907
R14251 CSoutput.n352 CSoutput.t30 2.82907
R14252 CSoutput.n352 CSoutput.t20 2.82907
R14253 CSoutput.n350 CSoutput.t51 2.82907
R14254 CSoutput.n350 CSoutput.t53 2.82907
R14255 CSoutput.n349 CSoutput.t35 2.82907
R14256 CSoutput.n349 CSoutput.t25 2.82907
R14257 CSoutput.n384 CSoutput.t21 2.82907
R14258 CSoutput.n384 CSoutput.t33 2.82907
R14259 CSoutput.n385 CSoutput.t50 2.82907
R14260 CSoutput.n385 CSoutput.t13 2.82907
R14261 CSoutput.n387 CSoutput.t17 2.82907
R14262 CSoutput.n387 CSoutput.t27 2.82907
R14263 CSoutput.n389 CSoutput.t32 2.82907
R14264 CSoutput.n389 CSoutput.t19 2.82907
R14265 CSoutput.n391 CSoutput.t24 2.82907
R14266 CSoutput.n391 CSoutput.t36 2.82907
R14267 CSoutput.n393 CSoutput.t41 2.82907
R14268 CSoutput.n393 CSoutput.t54 2.82907
R14269 CSoutput.n373 CSoutput.t14 2.82907
R14270 CSoutput.n373 CSoutput.t22 2.82907
R14271 CSoutput.n374 CSoutput.t43 2.82907
R14272 CSoutput.n374 CSoutput.t55 2.82907
R14273 CSoutput.n376 CSoutput.t58 2.82907
R14274 CSoutput.n376 CSoutput.t18 2.82907
R14275 CSoutput.n378 CSoutput.t23 2.82907
R14276 CSoutput.n378 CSoutput.t12 2.82907
R14277 CSoutput.n380 CSoutput.t16 2.82907
R14278 CSoutput.n380 CSoutput.t26 2.82907
R14279 CSoutput.n382 CSoutput.t31 2.82907
R14280 CSoutput.n382 CSoutput.t47 2.82907
R14281 CSoutput.n396 CSoutput.n372 2.75627
R14282 CSoutput.n348 CSoutput.n138 2.57547
R14283 CSoutput.n75 CSoutput.n1 2.45513
R14284 CSoutput.n229 CSoutput.n227 2.251
R14285 CSoutput.n229 CSoutput.n226 2.251
R14286 CSoutput.n229 CSoutput.n225 2.251
R14287 CSoutput.n229 CSoutput.n224 2.251
R14288 CSoutput.n198 CSoutput.n197 2.251
R14289 CSoutput.n198 CSoutput.n196 2.251
R14290 CSoutput.n198 CSoutput.n195 2.251
R14291 CSoutput.n198 CSoutput.n194 2.251
R14292 CSoutput.n271 CSoutput.n270 2.251
R14293 CSoutput.n236 CSoutput.n234 2.251
R14294 CSoutput.n236 CSoutput.n233 2.251
R14295 CSoutput.n236 CSoutput.n232 2.251
R14296 CSoutput.n254 CSoutput.n236 2.251
R14297 CSoutput.n242 CSoutput.n241 2.251
R14298 CSoutput.n242 CSoutput.n240 2.251
R14299 CSoutput.n242 CSoutput.n239 2.251
R14300 CSoutput.n242 CSoutput.n238 2.251
R14301 CSoutput.n268 CSoutput.n208 2.251
R14302 CSoutput.n263 CSoutput.n261 2.251
R14303 CSoutput.n263 CSoutput.n260 2.251
R14304 CSoutput.n263 CSoutput.n259 2.251
R14305 CSoutput.n263 CSoutput.n258 2.251
R14306 CSoutput.n164 CSoutput.n163 2.251
R14307 CSoutput.n164 CSoutput.n162 2.251
R14308 CSoutput.n164 CSoutput.n161 2.251
R14309 CSoutput.n164 CSoutput.n160 2.251
R14310 CSoutput.n281 CSoutput.n280 2.251
R14311 CSoutput.n198 CSoutput.n178 2.2505
R14312 CSoutput.n193 CSoutput.n178 2.2505
R14313 CSoutput.n191 CSoutput.n178 2.2505
R14314 CSoutput.n190 CSoutput.n178 2.2505
R14315 CSoutput.n275 CSoutput.n178 2.2505
R14316 CSoutput.n273 CSoutput.n178 2.2505
R14317 CSoutput.n271 CSoutput.n178 2.2505
R14318 CSoutput.n201 CSoutput.n178 2.2505
R14319 CSoutput.n200 CSoutput.n178 2.2505
R14320 CSoutput.n204 CSoutput.n178 2.2505
R14321 CSoutput.n203 CSoutput.n178 2.2505
R14322 CSoutput.n186 CSoutput.n178 2.2505
R14323 CSoutput.n278 CSoutput.n178 2.2505
R14324 CSoutput.n278 CSoutput.n277 2.2505
R14325 CSoutput.n242 CSoutput.n213 2.2505
R14326 CSoutput.n223 CSoutput.n213 2.2505
R14327 CSoutput.n244 CSoutput.n213 2.2505
R14328 CSoutput.n222 CSoutput.n213 2.2505
R14329 CSoutput.n246 CSoutput.n213 2.2505
R14330 CSoutput.n213 CSoutput.n207 2.2505
R14331 CSoutput.n268 CSoutput.n213 2.2505
R14332 CSoutput.n266 CSoutput.n213 2.2505
R14333 CSoutput.n248 CSoutput.n213 2.2505
R14334 CSoutput.n220 CSoutput.n213 2.2505
R14335 CSoutput.n250 CSoutput.n213 2.2505
R14336 CSoutput.n219 CSoutput.n213 2.2505
R14337 CSoutput.n264 CSoutput.n213 2.2505
R14338 CSoutput.n264 CSoutput.n217 2.2505
R14339 CSoutput.n164 CSoutput.n144 2.2505
R14340 CSoutput.n159 CSoutput.n144 2.2505
R14341 CSoutput.n157 CSoutput.n144 2.2505
R14342 CSoutput.n156 CSoutput.n144 2.2505
R14343 CSoutput.n285 CSoutput.n144 2.2505
R14344 CSoutput.n283 CSoutput.n144 2.2505
R14345 CSoutput.n281 CSoutput.n144 2.2505
R14346 CSoutput.n167 CSoutput.n144 2.2505
R14347 CSoutput.n166 CSoutput.n144 2.2505
R14348 CSoutput.n170 CSoutput.n144 2.2505
R14349 CSoutput.n169 CSoutput.n144 2.2505
R14350 CSoutput.n152 CSoutput.n144 2.2505
R14351 CSoutput.n288 CSoutput.n144 2.2505
R14352 CSoutput.n288 CSoutput.n287 2.2505
R14353 CSoutput.n206 CSoutput.n199 2.25024
R14354 CSoutput.n206 CSoutput.n192 2.25024
R14355 CSoutput.n274 CSoutput.n206 2.25024
R14356 CSoutput.n206 CSoutput.n202 2.25024
R14357 CSoutput.n206 CSoutput.n205 2.25024
R14358 CSoutput.n206 CSoutput.n173 2.25024
R14359 CSoutput.n256 CSoutput.n253 2.25024
R14360 CSoutput.n256 CSoutput.n252 2.25024
R14361 CSoutput.n256 CSoutput.n251 2.25024
R14362 CSoutput.n256 CSoutput.n218 2.25024
R14363 CSoutput.n256 CSoutput.n255 2.25024
R14364 CSoutput.n257 CSoutput.n256 2.25024
R14365 CSoutput.n172 CSoutput.n165 2.25024
R14366 CSoutput.n172 CSoutput.n158 2.25024
R14367 CSoutput.n284 CSoutput.n172 2.25024
R14368 CSoutput.n172 CSoutput.n168 2.25024
R14369 CSoutput.n172 CSoutput.n171 2.25024
R14370 CSoutput.n172 CSoutput.n139 2.25024
R14371 CSoutput.n273 CSoutput.n183 1.50111
R14372 CSoutput.n221 CSoutput.n207 1.50111
R14373 CSoutput.n283 CSoutput.n149 1.50111
R14374 CSoutput.n229 CSoutput.n228 1.501
R14375 CSoutput.n236 CSoutput.n235 1.501
R14376 CSoutput.n263 CSoutput.n262 1.501
R14377 CSoutput.n277 CSoutput.n188 1.12536
R14378 CSoutput.n277 CSoutput.n189 1.12536
R14379 CSoutput.n277 CSoutput.n276 1.12536
R14380 CSoutput.n237 CSoutput.n217 1.12536
R14381 CSoutput.n243 CSoutput.n217 1.12536
R14382 CSoutput.n245 CSoutput.n217 1.12536
R14383 CSoutput.n287 CSoutput.n154 1.12536
R14384 CSoutput.n287 CSoutput.n155 1.12536
R14385 CSoutput.n287 CSoutput.n286 1.12536
R14386 CSoutput.n277 CSoutput.n184 1.12536
R14387 CSoutput.n277 CSoutput.n185 1.12536
R14388 CSoutput.n277 CSoutput.n187 1.12536
R14389 CSoutput.n267 CSoutput.n217 1.12536
R14390 CSoutput.n247 CSoutput.n217 1.12536
R14391 CSoutput.n249 CSoutput.n217 1.12536
R14392 CSoutput.n287 CSoutput.n150 1.12536
R14393 CSoutput.n287 CSoutput.n151 1.12536
R14394 CSoutput.n287 CSoutput.n153 1.12536
R14395 CSoutput.n31 CSoutput.n30 0.669944
R14396 CSoutput.n62 CSoutput.n61 0.669944
R14397 CSoutput.n364 CSoutput.n362 0.573776
R14398 CSoutput.n366 CSoutput.n364 0.573776
R14399 CSoutput.n368 CSoutput.n366 0.573776
R14400 CSoutput.n370 CSoutput.n368 0.573776
R14401 CSoutput.n353 CSoutput.n351 0.573776
R14402 CSoutput.n355 CSoutput.n353 0.573776
R14403 CSoutput.n357 CSoutput.n355 0.573776
R14404 CSoutput.n359 CSoutput.n357 0.573776
R14405 CSoutput.n394 CSoutput.n392 0.573776
R14406 CSoutput.n392 CSoutput.n390 0.573776
R14407 CSoutput.n390 CSoutput.n388 0.573776
R14408 CSoutput.n388 CSoutput.n386 0.573776
R14409 CSoutput.n383 CSoutput.n381 0.573776
R14410 CSoutput.n381 CSoutput.n379 0.573776
R14411 CSoutput.n379 CSoutput.n377 0.573776
R14412 CSoutput.n377 CSoutput.n375 0.573776
R14413 CSoutput.n397 CSoutput.n288 0.53442
R14414 CSoutput.n332 CSoutput.n330 0.358259
R14415 CSoutput.n334 CSoutput.n332 0.358259
R14416 CSoutput.n336 CSoutput.n334 0.358259
R14417 CSoutput.n338 CSoutput.n336 0.358259
R14418 CSoutput.n340 CSoutput.n338 0.358259
R14419 CSoutput.n342 CSoutput.n340 0.358259
R14420 CSoutput.n344 CSoutput.n342 0.358259
R14421 CSoutput.n346 CSoutput.n344 0.358259
R14422 CSoutput.n312 CSoutput.n310 0.358259
R14423 CSoutput.n314 CSoutput.n312 0.358259
R14424 CSoutput.n316 CSoutput.n314 0.358259
R14425 CSoutput.n318 CSoutput.n316 0.358259
R14426 CSoutput.n320 CSoutput.n318 0.358259
R14427 CSoutput.n322 CSoutput.n320 0.358259
R14428 CSoutput.n324 CSoutput.n322 0.358259
R14429 CSoutput.n326 CSoutput.n324 0.358259
R14430 CSoutput.n293 CSoutput.n291 0.358259
R14431 CSoutput.n295 CSoutput.n293 0.358259
R14432 CSoutput.n297 CSoutput.n295 0.358259
R14433 CSoutput.n299 CSoutput.n297 0.358259
R14434 CSoutput.n301 CSoutput.n299 0.358259
R14435 CSoutput.n303 CSoutput.n301 0.358259
R14436 CSoutput.n305 CSoutput.n303 0.358259
R14437 CSoutput.n307 CSoutput.n305 0.358259
R14438 CSoutput.n136 CSoutput.n134 0.358259
R14439 CSoutput.n134 CSoutput.n132 0.358259
R14440 CSoutput.n132 CSoutput.n130 0.358259
R14441 CSoutput.n130 CSoutput.n128 0.358259
R14442 CSoutput.n128 CSoutput.n126 0.358259
R14443 CSoutput.n126 CSoutput.n124 0.358259
R14444 CSoutput.n124 CSoutput.n122 0.358259
R14445 CSoutput.n122 CSoutput.n120 0.358259
R14446 CSoutput.n116 CSoutput.n114 0.358259
R14447 CSoutput.n114 CSoutput.n112 0.358259
R14448 CSoutput.n112 CSoutput.n110 0.358259
R14449 CSoutput.n110 CSoutput.n108 0.358259
R14450 CSoutput.n108 CSoutput.n106 0.358259
R14451 CSoutput.n106 CSoutput.n104 0.358259
R14452 CSoutput.n104 CSoutput.n102 0.358259
R14453 CSoutput.n102 CSoutput.n100 0.358259
R14454 CSoutput.n97 CSoutput.n95 0.358259
R14455 CSoutput.n95 CSoutput.n93 0.358259
R14456 CSoutput.n93 CSoutput.n91 0.358259
R14457 CSoutput.n91 CSoutput.n89 0.358259
R14458 CSoutput.n89 CSoutput.n87 0.358259
R14459 CSoutput.n87 CSoutput.n85 0.358259
R14460 CSoutput.n85 CSoutput.n83 0.358259
R14461 CSoutput.n83 CSoutput.n81 0.358259
R14462 CSoutput.n21 CSoutput.n20 0.169105
R14463 CSoutput.n21 CSoutput.n16 0.169105
R14464 CSoutput.n26 CSoutput.n16 0.169105
R14465 CSoutput.n27 CSoutput.n26 0.169105
R14466 CSoutput.n27 CSoutput.n14 0.169105
R14467 CSoutput.n32 CSoutput.n14 0.169105
R14468 CSoutput.n33 CSoutput.n32 0.169105
R14469 CSoutput.n34 CSoutput.n33 0.169105
R14470 CSoutput.n34 CSoutput.n12 0.169105
R14471 CSoutput.n39 CSoutput.n12 0.169105
R14472 CSoutput.n40 CSoutput.n39 0.169105
R14473 CSoutput.n40 CSoutput.n10 0.169105
R14474 CSoutput.n45 CSoutput.n10 0.169105
R14475 CSoutput.n46 CSoutput.n45 0.169105
R14476 CSoutput.n47 CSoutput.n46 0.169105
R14477 CSoutput.n47 CSoutput.n8 0.169105
R14478 CSoutput.n52 CSoutput.n8 0.169105
R14479 CSoutput.n53 CSoutput.n52 0.169105
R14480 CSoutput.n53 CSoutput.n6 0.169105
R14481 CSoutput.n58 CSoutput.n6 0.169105
R14482 CSoutput.n59 CSoutput.n58 0.169105
R14483 CSoutput.n60 CSoutput.n59 0.169105
R14484 CSoutput.n60 CSoutput.n4 0.169105
R14485 CSoutput.n66 CSoutput.n4 0.169105
R14486 CSoutput.n67 CSoutput.n66 0.169105
R14487 CSoutput.n68 CSoutput.n67 0.169105
R14488 CSoutput.n68 CSoutput.n2 0.169105
R14489 CSoutput.n73 CSoutput.n2 0.169105
R14490 CSoutput.n74 CSoutput.n73 0.169105
R14491 CSoutput.n74 CSoutput.n0 0.169105
R14492 CSoutput.n78 CSoutput.n0 0.169105
R14493 CSoutput.n231 CSoutput.n230 0.0910737
R14494 CSoutput.n282 CSoutput.n279 0.0723685
R14495 CSoutput.n236 CSoutput.n231 0.0522944
R14496 CSoutput.n279 CSoutput.n278 0.0499135
R14497 CSoutput.n230 CSoutput.n229 0.0499135
R14498 CSoutput.n264 CSoutput.n263 0.0464294
R14499 CSoutput.n272 CSoutput.n269 0.0391444
R14500 CSoutput.n231 CSoutput.t177 0.023435
R14501 CSoutput.n279 CSoutput.t176 0.02262
R14502 CSoutput.n230 CSoutput.t181 0.02262
R14503 CSoutput CSoutput.n397 0.0052
R14504 CSoutput.n201 CSoutput.n184 0.00365111
R14505 CSoutput.n204 CSoutput.n185 0.00365111
R14506 CSoutput.n187 CSoutput.n186 0.00365111
R14507 CSoutput.n229 CSoutput.n188 0.00365111
R14508 CSoutput.n193 CSoutput.n189 0.00365111
R14509 CSoutput.n276 CSoutput.n190 0.00365111
R14510 CSoutput.n267 CSoutput.n266 0.00365111
R14511 CSoutput.n247 CSoutput.n220 0.00365111
R14512 CSoutput.n249 CSoutput.n219 0.00365111
R14513 CSoutput.n237 CSoutput.n236 0.00365111
R14514 CSoutput.n243 CSoutput.n223 0.00365111
R14515 CSoutput.n245 CSoutput.n222 0.00365111
R14516 CSoutput.n167 CSoutput.n150 0.00365111
R14517 CSoutput.n170 CSoutput.n151 0.00365111
R14518 CSoutput.n153 CSoutput.n152 0.00365111
R14519 CSoutput.n263 CSoutput.n154 0.00365111
R14520 CSoutput.n159 CSoutput.n155 0.00365111
R14521 CSoutput.n286 CSoutput.n156 0.00365111
R14522 CSoutput.n198 CSoutput.n188 0.00340054
R14523 CSoutput.n191 CSoutput.n189 0.00340054
R14524 CSoutput.n276 CSoutput.n275 0.00340054
R14525 CSoutput.n271 CSoutput.n184 0.00340054
R14526 CSoutput.n200 CSoutput.n185 0.00340054
R14527 CSoutput.n203 CSoutput.n187 0.00340054
R14528 CSoutput.n242 CSoutput.n237 0.00340054
R14529 CSoutput.n244 CSoutput.n243 0.00340054
R14530 CSoutput.n246 CSoutput.n245 0.00340054
R14531 CSoutput.n268 CSoutput.n267 0.00340054
R14532 CSoutput.n248 CSoutput.n247 0.00340054
R14533 CSoutput.n250 CSoutput.n249 0.00340054
R14534 CSoutput.n164 CSoutput.n154 0.00340054
R14535 CSoutput.n157 CSoutput.n155 0.00340054
R14536 CSoutput.n286 CSoutput.n285 0.00340054
R14537 CSoutput.n281 CSoutput.n150 0.00340054
R14538 CSoutput.n166 CSoutput.n151 0.00340054
R14539 CSoutput.n169 CSoutput.n153 0.00340054
R14540 CSoutput.n199 CSoutput.n193 0.00252698
R14541 CSoutput.n192 CSoutput.n190 0.00252698
R14542 CSoutput.n274 CSoutput.n273 0.00252698
R14543 CSoutput.n202 CSoutput.n200 0.00252698
R14544 CSoutput.n205 CSoutput.n203 0.00252698
R14545 CSoutput.n278 CSoutput.n173 0.00252698
R14546 CSoutput.n199 CSoutput.n198 0.00252698
R14547 CSoutput.n192 CSoutput.n191 0.00252698
R14548 CSoutput.n275 CSoutput.n274 0.00252698
R14549 CSoutput.n202 CSoutput.n201 0.00252698
R14550 CSoutput.n205 CSoutput.n204 0.00252698
R14551 CSoutput.n186 CSoutput.n173 0.00252698
R14552 CSoutput.n253 CSoutput.n223 0.00252698
R14553 CSoutput.n252 CSoutput.n222 0.00252698
R14554 CSoutput.n251 CSoutput.n207 0.00252698
R14555 CSoutput.n248 CSoutput.n218 0.00252698
R14556 CSoutput.n255 CSoutput.n250 0.00252698
R14557 CSoutput.n264 CSoutput.n257 0.00252698
R14558 CSoutput.n253 CSoutput.n242 0.00252698
R14559 CSoutput.n252 CSoutput.n244 0.00252698
R14560 CSoutput.n251 CSoutput.n246 0.00252698
R14561 CSoutput.n266 CSoutput.n218 0.00252698
R14562 CSoutput.n255 CSoutput.n220 0.00252698
R14563 CSoutput.n257 CSoutput.n219 0.00252698
R14564 CSoutput.n165 CSoutput.n159 0.00252698
R14565 CSoutput.n158 CSoutput.n156 0.00252698
R14566 CSoutput.n284 CSoutput.n283 0.00252698
R14567 CSoutput.n168 CSoutput.n166 0.00252698
R14568 CSoutput.n171 CSoutput.n169 0.00252698
R14569 CSoutput.n288 CSoutput.n139 0.00252698
R14570 CSoutput.n165 CSoutput.n164 0.00252698
R14571 CSoutput.n158 CSoutput.n157 0.00252698
R14572 CSoutput.n285 CSoutput.n284 0.00252698
R14573 CSoutput.n168 CSoutput.n167 0.00252698
R14574 CSoutput.n171 CSoutput.n170 0.00252698
R14575 CSoutput.n152 CSoutput.n139 0.00252698
R14576 CSoutput.n273 CSoutput.n272 0.0020275
R14577 CSoutput.n272 CSoutput.n271 0.0020275
R14578 CSoutput.n269 CSoutput.n207 0.0020275
R14579 CSoutput.n269 CSoutput.n268 0.0020275
R14580 CSoutput.n283 CSoutput.n282 0.0020275
R14581 CSoutput.n282 CSoutput.n281 0.0020275
R14582 CSoutput.n183 CSoutput.n182 0.00166668
R14583 CSoutput.n265 CSoutput.n221 0.00166668
R14584 CSoutput.n149 CSoutput.n148 0.00166668
R14585 CSoutput.n287 CSoutput.n149 0.00133328
R14586 CSoutput.n221 CSoutput.n217 0.00133328
R14587 CSoutput.n277 CSoutput.n183 0.00133328
R14588 CSoutput.n280 CSoutput.n172 0.001
R14589 CSoutput.n258 CSoutput.n172 0.001
R14590 CSoutput.n160 CSoutput.n140 0.001
R14591 CSoutput.n259 CSoutput.n140 0.001
R14592 CSoutput.n161 CSoutput.n141 0.001
R14593 CSoutput.n260 CSoutput.n141 0.001
R14594 CSoutput.n162 CSoutput.n142 0.001
R14595 CSoutput.n261 CSoutput.n142 0.001
R14596 CSoutput.n163 CSoutput.n143 0.001
R14597 CSoutput.n262 CSoutput.n143 0.001
R14598 CSoutput.n256 CSoutput.n208 0.001
R14599 CSoutput.n256 CSoutput.n254 0.001
R14600 CSoutput.n238 CSoutput.n209 0.001
R14601 CSoutput.n232 CSoutput.n209 0.001
R14602 CSoutput.n239 CSoutput.n210 0.001
R14603 CSoutput.n233 CSoutput.n210 0.001
R14604 CSoutput.n240 CSoutput.n211 0.001
R14605 CSoutput.n234 CSoutput.n211 0.001
R14606 CSoutput.n241 CSoutput.n212 0.001
R14607 CSoutput.n235 CSoutput.n212 0.001
R14608 CSoutput.n270 CSoutput.n206 0.001
R14609 CSoutput.n224 CSoutput.n206 0.001
R14610 CSoutput.n194 CSoutput.n174 0.001
R14611 CSoutput.n225 CSoutput.n174 0.001
R14612 CSoutput.n195 CSoutput.n175 0.001
R14613 CSoutput.n226 CSoutput.n175 0.001
R14614 CSoutput.n196 CSoutput.n176 0.001
R14615 CSoutput.n227 CSoutput.n176 0.001
R14616 CSoutput.n197 CSoutput.n177 0.001
R14617 CSoutput.n228 CSoutput.n177 0.001
R14618 CSoutput.n228 CSoutput.n178 0.001
R14619 CSoutput.n227 CSoutput.n179 0.001
R14620 CSoutput.n226 CSoutput.n180 0.001
R14621 CSoutput.n225 CSoutput.t174 0.001
R14622 CSoutput.n224 CSoutput.n181 0.001
R14623 CSoutput.n197 CSoutput.n179 0.001
R14624 CSoutput.n196 CSoutput.n180 0.001
R14625 CSoutput.n195 CSoutput.t174 0.001
R14626 CSoutput.n194 CSoutput.n181 0.001
R14627 CSoutput.n270 CSoutput.n182 0.001
R14628 CSoutput.n235 CSoutput.n213 0.001
R14629 CSoutput.n234 CSoutput.n214 0.001
R14630 CSoutput.n233 CSoutput.n215 0.001
R14631 CSoutput.n232 CSoutput.t170 0.001
R14632 CSoutput.n254 CSoutput.n216 0.001
R14633 CSoutput.n241 CSoutput.n214 0.001
R14634 CSoutput.n240 CSoutput.n215 0.001
R14635 CSoutput.n239 CSoutput.t170 0.001
R14636 CSoutput.n238 CSoutput.n216 0.001
R14637 CSoutput.n265 CSoutput.n208 0.001
R14638 CSoutput.n262 CSoutput.n144 0.001
R14639 CSoutput.n261 CSoutput.n145 0.001
R14640 CSoutput.n260 CSoutput.n146 0.001
R14641 CSoutput.n259 CSoutput.t187 0.001
R14642 CSoutput.n258 CSoutput.n147 0.001
R14643 CSoutput.n163 CSoutput.n145 0.001
R14644 CSoutput.n162 CSoutput.n146 0.001
R14645 CSoutput.n161 CSoutput.t187 0.001
R14646 CSoutput.n160 CSoutput.n147 0.001
R14647 CSoutput.n280 CSoutput.n148 0.001
R14648 a_n7636_8799.n229 a_n7636_8799.t63 485.149
R14649 a_n7636_8799.n248 a_n7636_8799.t76 485.149
R14650 a_n7636_8799.n268 a_n7636_8799.t115 485.149
R14651 a_n7636_8799.n168 a_n7636_8799.t138 485.149
R14652 a_n7636_8799.n187 a_n7636_8799.t152 485.149
R14653 a_n7636_8799.n207 a_n7636_8799.t113 485.149
R14654 a_n7636_8799.n54 a_n7636_8799.t87 485.135
R14655 a_n7636_8799.n241 a_n7636_8799.t86 464.166
R14656 a_n7636_8799.n223 a_n7636_8799.t60 464.166
R14657 a_n7636_8799.n240 a_n7636_8799.t135 464.166
R14658 a_n7636_8799.n239 a_n7636_8799.t90 464.166
R14659 a_n7636_8799.n224 a_n7636_8799.t66 464.166
R14660 a_n7636_8799.n238 a_n7636_8799.t140 464.166
R14661 a_n7636_8799.n237 a_n7636_8799.t107 464.166
R14662 a_n7636_8799.n225 a_n7636_8799.t105 464.166
R14663 a_n7636_8799.n236 a_n7636_8799.t40 464.166
R14664 a_n7636_8799.n235 a_n7636_8799.t111 464.166
R14665 a_n7636_8799.n226 a_n7636_8799.t110 464.166
R14666 a_n7636_8799.n234 a_n7636_8799.t42 464.166
R14667 a_n7636_8799.n233 a_n7636_8799.t41 464.166
R14668 a_n7636_8799.n227 a_n7636_8799.t127 464.166
R14669 a_n7636_8799.n232 a_n7636_8799.t59 464.166
R14670 a_n7636_8799.n231 a_n7636_8799.t43 464.166
R14671 a_n7636_8799.n228 a_n7636_8799.t129 464.166
R14672 a_n7636_8799.n230 a_n7636_8799.t89 464.166
R14673 a_n7636_8799.n69 a_n7636_8799.t97 485.135
R14674 a_n7636_8799.n260 a_n7636_8799.t96 464.166
R14675 a_n7636_8799.n242 a_n7636_8799.t74 464.166
R14676 a_n7636_8799.n259 a_n7636_8799.t150 464.166
R14677 a_n7636_8799.n258 a_n7636_8799.t104 464.166
R14678 a_n7636_8799.n243 a_n7636_8799.t77 464.166
R14679 a_n7636_8799.n257 a_n7636_8799.t36 464.166
R14680 a_n7636_8799.n256 a_n7636_8799.t120 464.166
R14681 a_n7636_8799.n244 a_n7636_8799.t119 464.166
R14682 a_n7636_8799.n255 a_n7636_8799.t50 464.166
R14683 a_n7636_8799.n254 a_n7636_8799.t123 464.166
R14684 a_n7636_8799.n245 a_n7636_8799.t122 464.166
R14685 a_n7636_8799.n253 a_n7636_8799.t54 464.166
R14686 a_n7636_8799.n252 a_n7636_8799.t53 464.166
R14687 a_n7636_8799.n246 a_n7636_8799.t144 464.166
R14688 a_n7636_8799.n251 a_n7636_8799.t75 464.166
R14689 a_n7636_8799.n250 a_n7636_8799.t56 464.166
R14690 a_n7636_8799.n247 a_n7636_8799.t145 464.166
R14691 a_n7636_8799.n249 a_n7636_8799.t103 464.166
R14692 a_n7636_8799.n84 a_n7636_8799.t154 485.135
R14693 a_n7636_8799.n280 a_n7636_8799.t52 464.166
R14694 a_n7636_8799.n262 a_n7636_8799.t101 464.166
R14695 a_n7636_8799.n279 a_n7636_8799.t38 464.166
R14696 a_n7636_8799.n278 a_n7636_8799.t125 464.166
R14697 a_n7636_8799.n263 a_n7636_8799.t65 464.166
R14698 a_n7636_8799.n277 a_n7636_8799.t108 464.166
R14699 a_n7636_8799.n276 a_n7636_8799.t44 464.166
R14700 a_n7636_8799.n264 a_n7636_8799.t70 464.166
R14701 a_n7636_8799.n275 a_n7636_8799.t148 464.166
R14702 a_n7636_8799.n274 a_n7636_8799.t117 464.166
R14703 a_n7636_8799.n265 a_n7636_8799.t143 464.166
R14704 a_n7636_8799.n273 a_n7636_8799.t100 464.166
R14705 a_n7636_8799.n272 a_n7636_8799.t121 464.166
R14706 a_n7636_8799.n266 a_n7636_8799.t58 464.166
R14707 a_n7636_8799.n271 a_n7636_8799.t141 464.166
R14708 a_n7636_8799.n270 a_n7636_8799.t82 464.166
R14709 a_n7636_8799.n267 a_n7636_8799.t131 464.166
R14710 a_n7636_8799.n269 a_n7636_8799.t68 464.166
R14711 a_n7636_8799.n169 a_n7636_8799.t137 464.166
R14712 a_n7636_8799.n170 a_n7636_8799.t88 464.166
R14713 a_n7636_8799.n171 a_n7636_8799.t116 464.166
R14714 a_n7636_8799.n172 a_n7636_8799.t134 464.166
R14715 a_n7636_8799.n167 a_n7636_8799.t85 464.166
R14716 a_n7636_8799.n173 a_n7636_8799.t84 464.166
R14717 a_n7636_8799.n174 a_n7636_8799.t114 464.166
R14718 a_n7636_8799.n175 a_n7636_8799.t72 464.166
R14719 a_n7636_8799.n176 a_n7636_8799.t73 464.166
R14720 a_n7636_8799.n166 a_n7636_8799.t112 464.166
R14721 a_n7636_8799.n177 a_n7636_8799.t37 464.166
R14722 a_n7636_8799.n165 a_n7636_8799.t69 464.166
R14723 a_n7636_8799.n178 a_n7636_8799.t93 464.166
R14724 a_n7636_8799.n179 a_n7636_8799.t136 464.166
R14725 a_n7636_8799.n180 a_n7636_8799.t48 464.166
R14726 a_n7636_8799.n181 a_n7636_8799.t67 464.166
R14727 a_n7636_8799.n164 a_n7636_8799.t133 464.166
R14728 a_n7636_8799.n182 a_n7636_8799.t47 464.166
R14729 a_n7636_8799.n188 a_n7636_8799.t153 464.166
R14730 a_n7636_8799.n189 a_n7636_8799.t98 464.166
R14731 a_n7636_8799.n190 a_n7636_8799.t130 464.166
R14732 a_n7636_8799.n191 a_n7636_8799.t147 464.166
R14733 a_n7636_8799.n186 a_n7636_8799.t94 464.166
R14734 a_n7636_8799.n192 a_n7636_8799.t95 464.166
R14735 a_n7636_8799.n193 a_n7636_8799.t128 464.166
R14736 a_n7636_8799.n194 a_n7636_8799.t81 464.166
R14737 a_n7636_8799.n195 a_n7636_8799.t83 464.166
R14738 a_n7636_8799.n185 a_n7636_8799.t124 464.166
R14739 a_n7636_8799.n196 a_n7636_8799.t49 464.166
R14740 a_n7636_8799.n184 a_n7636_8799.t79 464.166
R14741 a_n7636_8799.n197 a_n7636_8799.t106 464.166
R14742 a_n7636_8799.n198 a_n7636_8799.t151 464.166
R14743 a_n7636_8799.n199 a_n7636_8799.t64 464.166
R14744 a_n7636_8799.n200 a_n7636_8799.t78 464.166
R14745 a_n7636_8799.n183 a_n7636_8799.t146 464.166
R14746 a_n7636_8799.n201 a_n7636_8799.t57 464.166
R14747 a_n7636_8799.n208 a_n7636_8799.t92 464.166
R14748 a_n7636_8799.n209 a_n7636_8799.t132 464.166
R14749 a_n7636_8799.n210 a_n7636_8799.t80 464.166
R14750 a_n7636_8799.n211 a_n7636_8799.t139 464.166
R14751 a_n7636_8799.n206 a_n7636_8799.t55 464.166
R14752 a_n7636_8799.n212 a_n7636_8799.t39 464.166
R14753 a_n7636_8799.n213 a_n7636_8799.t99 464.166
R14754 a_n7636_8799.n214 a_n7636_8799.t142 464.166
R14755 a_n7636_8799.n215 a_n7636_8799.t118 464.166
R14756 a_n7636_8799.n205 a_n7636_8799.t149 464.166
R14757 a_n7636_8799.n216 a_n7636_8799.t91 464.166
R14758 a_n7636_8799.n204 a_n7636_8799.t45 464.166
R14759 a_n7636_8799.n217 a_n7636_8799.t109 464.166
R14760 a_n7636_8799.n218 a_n7636_8799.t62 464.166
R14761 a_n7636_8799.n219 a_n7636_8799.t126 464.166
R14762 a_n7636_8799.n220 a_n7636_8799.t71 464.166
R14763 a_n7636_8799.n203 a_n7636_8799.t102 464.166
R14764 a_n7636_8799.n221 a_n7636_8799.t51 464.166
R14765 a_n7636_8799.n41 a_n7636_8799.n68 71.7212
R14766 a_n7636_8799.n68 a_n7636_8799.n228 17.8606
R14767 a_n7636_8799.n67 a_n7636_8799.n41 76.9909
R14768 a_n7636_8799.n231 a_n7636_8799.n67 7.32118
R14769 a_n7636_8799.n66 a_n7636_8799.n40 78.3454
R14770 a_n7636_8799.n40 a_n7636_8799.n65 72.8951
R14771 a_n7636_8799.n64 a_n7636_8799.n42 70.1674
R14772 a_n7636_8799.n234 a_n7636_8799.n64 20.9683
R14773 a_n7636_8799.n42 a_n7636_8799.n63 72.3034
R14774 a_n7636_8799.n63 a_n7636_8799.n226 16.6962
R14775 a_n7636_8799.n62 a_n7636_8799.n43 77.6622
R14776 a_n7636_8799.n235 a_n7636_8799.n62 5.97853
R14777 a_n7636_8799.n61 a_n7636_8799.n43 77.6622
R14778 a_n7636_8799.n44 a_n7636_8799.n60 72.3034
R14779 a_n7636_8799.n59 a_n7636_8799.n44 70.1674
R14780 a_n7636_8799.n238 a_n7636_8799.n59 20.9683
R14781 a_n7636_8799.n46 a_n7636_8799.n58 72.8951
R14782 a_n7636_8799.n58 a_n7636_8799.n224 15.5127
R14783 a_n7636_8799.n57 a_n7636_8799.n46 78.3454
R14784 a_n7636_8799.n239 a_n7636_8799.n57 4.61226
R14785 a_n7636_8799.n56 a_n7636_8799.n45 76.9909
R14786 a_n7636_8799.n45 a_n7636_8799.n55 71.7212
R14787 a_n7636_8799.n241 a_n7636_8799.n54 20.9683
R14788 a_n7636_8799.n47 a_n7636_8799.n54 70.1674
R14789 a_n7636_8799.n33 a_n7636_8799.n83 71.7212
R14790 a_n7636_8799.n83 a_n7636_8799.n247 17.8606
R14791 a_n7636_8799.n82 a_n7636_8799.n33 76.9909
R14792 a_n7636_8799.n250 a_n7636_8799.n82 7.32118
R14793 a_n7636_8799.n81 a_n7636_8799.n32 78.3454
R14794 a_n7636_8799.n32 a_n7636_8799.n80 72.8951
R14795 a_n7636_8799.n79 a_n7636_8799.n34 70.1674
R14796 a_n7636_8799.n253 a_n7636_8799.n79 20.9683
R14797 a_n7636_8799.n34 a_n7636_8799.n78 72.3034
R14798 a_n7636_8799.n78 a_n7636_8799.n245 16.6962
R14799 a_n7636_8799.n77 a_n7636_8799.n35 77.6622
R14800 a_n7636_8799.n254 a_n7636_8799.n77 5.97853
R14801 a_n7636_8799.n76 a_n7636_8799.n35 77.6622
R14802 a_n7636_8799.n36 a_n7636_8799.n75 72.3034
R14803 a_n7636_8799.n74 a_n7636_8799.n36 70.1674
R14804 a_n7636_8799.n257 a_n7636_8799.n74 20.9683
R14805 a_n7636_8799.n38 a_n7636_8799.n73 72.8951
R14806 a_n7636_8799.n73 a_n7636_8799.n243 15.5127
R14807 a_n7636_8799.n72 a_n7636_8799.n38 78.3454
R14808 a_n7636_8799.n258 a_n7636_8799.n72 4.61226
R14809 a_n7636_8799.n71 a_n7636_8799.n37 76.9909
R14810 a_n7636_8799.n37 a_n7636_8799.n70 71.7212
R14811 a_n7636_8799.n260 a_n7636_8799.n69 20.9683
R14812 a_n7636_8799.n39 a_n7636_8799.n69 70.1674
R14813 a_n7636_8799.n25 a_n7636_8799.n98 71.7212
R14814 a_n7636_8799.n98 a_n7636_8799.n267 17.8606
R14815 a_n7636_8799.n97 a_n7636_8799.n25 76.9909
R14816 a_n7636_8799.n270 a_n7636_8799.n97 7.32118
R14817 a_n7636_8799.n96 a_n7636_8799.n24 78.3454
R14818 a_n7636_8799.n24 a_n7636_8799.n95 72.8951
R14819 a_n7636_8799.n94 a_n7636_8799.n26 70.1674
R14820 a_n7636_8799.n273 a_n7636_8799.n94 20.9683
R14821 a_n7636_8799.n26 a_n7636_8799.n93 72.3034
R14822 a_n7636_8799.n93 a_n7636_8799.n265 16.6962
R14823 a_n7636_8799.n92 a_n7636_8799.n27 77.6622
R14824 a_n7636_8799.n274 a_n7636_8799.n92 5.97853
R14825 a_n7636_8799.n91 a_n7636_8799.n27 77.6622
R14826 a_n7636_8799.n28 a_n7636_8799.n90 72.3034
R14827 a_n7636_8799.n89 a_n7636_8799.n28 70.1674
R14828 a_n7636_8799.n277 a_n7636_8799.n89 20.9683
R14829 a_n7636_8799.n30 a_n7636_8799.n88 72.8951
R14830 a_n7636_8799.n88 a_n7636_8799.n263 15.5127
R14831 a_n7636_8799.n87 a_n7636_8799.n30 78.3454
R14832 a_n7636_8799.n278 a_n7636_8799.n87 4.61226
R14833 a_n7636_8799.n86 a_n7636_8799.n29 76.9909
R14834 a_n7636_8799.n29 a_n7636_8799.n85 71.7212
R14835 a_n7636_8799.n280 a_n7636_8799.n84 20.9683
R14836 a_n7636_8799.n31 a_n7636_8799.n84 70.1674
R14837 a_n7636_8799.n17 a_n7636_8799.n113 70.1674
R14838 a_n7636_8799.n182 a_n7636_8799.n113 20.9683
R14839 a_n7636_8799.n112 a_n7636_8799.n17 71.7212
R14840 a_n7636_8799.n112 a_n7636_8799.n164 17.8606
R14841 a_n7636_8799.n16 a_n7636_8799.n111 76.9909
R14842 a_n7636_8799.n181 a_n7636_8799.n111 7.32118
R14843 a_n7636_8799.n110 a_n7636_8799.n16 78.3454
R14844 a_n7636_8799.n18 a_n7636_8799.n109 72.8951
R14845 a_n7636_8799.n108 a_n7636_8799.n18 70.1674
R14846 a_n7636_8799.n108 a_n7636_8799.n165 20.9683
R14847 a_n7636_8799.n19 a_n7636_8799.n107 72.3034
R14848 a_n7636_8799.n177 a_n7636_8799.n107 16.6962
R14849 a_n7636_8799.n106 a_n7636_8799.n19 77.6622
R14850 a_n7636_8799.n106 a_n7636_8799.n166 5.97853
R14851 a_n7636_8799.n20 a_n7636_8799.n105 77.6622
R14852 a_n7636_8799.n104 a_n7636_8799.n20 72.3034
R14853 a_n7636_8799.n21 a_n7636_8799.n103 70.1674
R14854 a_n7636_8799.n173 a_n7636_8799.n103 20.9683
R14855 a_n7636_8799.n102 a_n7636_8799.n21 72.8951
R14856 a_n7636_8799.n102 a_n7636_8799.n167 15.5127
R14857 a_n7636_8799.n22 a_n7636_8799.n101 78.3454
R14858 a_n7636_8799.n172 a_n7636_8799.n101 4.61226
R14859 a_n7636_8799.n100 a_n7636_8799.n22 76.9909
R14860 a_n7636_8799.n99 a_n7636_8799.n170 17.8606
R14861 a_n7636_8799.n99 a_n7636_8799.n23 71.7212
R14862 a_n7636_8799.n9 a_n7636_8799.n128 70.1674
R14863 a_n7636_8799.n201 a_n7636_8799.n128 20.9683
R14864 a_n7636_8799.n127 a_n7636_8799.n9 71.7212
R14865 a_n7636_8799.n127 a_n7636_8799.n183 17.8606
R14866 a_n7636_8799.n8 a_n7636_8799.n126 76.9909
R14867 a_n7636_8799.n200 a_n7636_8799.n126 7.32118
R14868 a_n7636_8799.n125 a_n7636_8799.n8 78.3454
R14869 a_n7636_8799.n10 a_n7636_8799.n124 72.8951
R14870 a_n7636_8799.n123 a_n7636_8799.n10 70.1674
R14871 a_n7636_8799.n123 a_n7636_8799.n184 20.9683
R14872 a_n7636_8799.n11 a_n7636_8799.n122 72.3034
R14873 a_n7636_8799.n196 a_n7636_8799.n122 16.6962
R14874 a_n7636_8799.n121 a_n7636_8799.n11 77.6622
R14875 a_n7636_8799.n121 a_n7636_8799.n185 5.97853
R14876 a_n7636_8799.n12 a_n7636_8799.n120 77.6622
R14877 a_n7636_8799.n119 a_n7636_8799.n12 72.3034
R14878 a_n7636_8799.n13 a_n7636_8799.n118 70.1674
R14879 a_n7636_8799.n192 a_n7636_8799.n118 20.9683
R14880 a_n7636_8799.n117 a_n7636_8799.n13 72.8951
R14881 a_n7636_8799.n117 a_n7636_8799.n186 15.5127
R14882 a_n7636_8799.n14 a_n7636_8799.n116 78.3454
R14883 a_n7636_8799.n191 a_n7636_8799.n116 4.61226
R14884 a_n7636_8799.n115 a_n7636_8799.n14 76.9909
R14885 a_n7636_8799.n114 a_n7636_8799.n189 17.8606
R14886 a_n7636_8799.n114 a_n7636_8799.n15 71.7212
R14887 a_n7636_8799.n1 a_n7636_8799.n143 70.1674
R14888 a_n7636_8799.n221 a_n7636_8799.n143 20.9683
R14889 a_n7636_8799.n142 a_n7636_8799.n1 71.7212
R14890 a_n7636_8799.n142 a_n7636_8799.n203 17.8606
R14891 a_n7636_8799.n0 a_n7636_8799.n141 76.9909
R14892 a_n7636_8799.n220 a_n7636_8799.n141 7.32118
R14893 a_n7636_8799.n140 a_n7636_8799.n0 78.3454
R14894 a_n7636_8799.n2 a_n7636_8799.n139 72.8951
R14895 a_n7636_8799.n138 a_n7636_8799.n2 70.1674
R14896 a_n7636_8799.n138 a_n7636_8799.n204 20.9683
R14897 a_n7636_8799.n3 a_n7636_8799.n137 72.3034
R14898 a_n7636_8799.n216 a_n7636_8799.n137 16.6962
R14899 a_n7636_8799.n136 a_n7636_8799.n3 77.6622
R14900 a_n7636_8799.n136 a_n7636_8799.n205 5.97853
R14901 a_n7636_8799.n4 a_n7636_8799.n135 77.6622
R14902 a_n7636_8799.n134 a_n7636_8799.n4 72.3034
R14903 a_n7636_8799.n5 a_n7636_8799.n133 70.1674
R14904 a_n7636_8799.n212 a_n7636_8799.n133 20.9683
R14905 a_n7636_8799.n132 a_n7636_8799.n5 72.8951
R14906 a_n7636_8799.n132 a_n7636_8799.n206 15.5127
R14907 a_n7636_8799.n6 a_n7636_8799.n131 78.3454
R14908 a_n7636_8799.n211 a_n7636_8799.n131 4.61226
R14909 a_n7636_8799.n130 a_n7636_8799.n6 76.9909
R14910 a_n7636_8799.n129 a_n7636_8799.n209 17.8606
R14911 a_n7636_8799.n129 a_n7636_8799.n7 71.7212
R14912 a_n7636_8799.n48 a_n7636_8799.n144 98.9633
R14913 a_n7636_8799.n287 a_n7636_8799.n49 98.9632
R14914 a_n7636_8799.n49 a_n7636_8799.n286 98.6055
R14915 a_n7636_8799.n49 a_n7636_8799.n285 98.6055
R14916 a_n7636_8799.n48 a_n7636_8799.n146 98.6055
R14917 a_n7636_8799.n48 a_n7636_8799.n145 98.6055
R14918 a_n7636_8799.n149 a_n7636_8799.n147 81.4626
R14919 a_n7636_8799.n157 a_n7636_8799.n155 81.4626
R14920 a_n7636_8799.n153 a_n7636_8799.n151 81.4626
R14921 a_n7636_8799.n160 a_n7636_8799.n159 80.9324
R14922 a_n7636_8799.n162 a_n7636_8799.n161 80.9324
R14923 a_n7636_8799.n53 a_n7636_8799.n163 80.9324
R14924 a_n7636_8799.n52 a_n7636_8799.n150 80.9324
R14925 a_n7636_8799.n149 a_n7636_8799.n148 80.9324
R14926 a_n7636_8799.n157 a_n7636_8799.n156 80.9324
R14927 a_n7636_8799.n51 a_n7636_8799.n158 80.9324
R14928 a_n7636_8799.n50 a_n7636_8799.n154 80.9324
R14929 a_n7636_8799.n153 a_n7636_8799.n152 80.9324
R14930 a_n7636_8799.n41 a_n7636_8799.n229 70.4033
R14931 a_n7636_8799.n33 a_n7636_8799.n248 70.4033
R14932 a_n7636_8799.n25 a_n7636_8799.n268 70.4033
R14933 a_n7636_8799.n168 a_n7636_8799.n23 70.4033
R14934 a_n7636_8799.n187 a_n7636_8799.n15 70.4033
R14935 a_n7636_8799.n207 a_n7636_8799.n7 70.4033
R14936 a_n7636_8799.n240 a_n7636_8799.n239 48.2005
R14937 a_n7636_8799.n59 a_n7636_8799.n237 20.9683
R14938 a_n7636_8799.n236 a_n7636_8799.n235 48.2005
R14939 a_n7636_8799.n64 a_n7636_8799.n233 20.9683
R14940 a_n7636_8799.n232 a_n7636_8799.n231 48.2005
R14941 a_n7636_8799.n259 a_n7636_8799.n258 48.2005
R14942 a_n7636_8799.n74 a_n7636_8799.n256 20.9683
R14943 a_n7636_8799.n255 a_n7636_8799.n254 48.2005
R14944 a_n7636_8799.n79 a_n7636_8799.n252 20.9683
R14945 a_n7636_8799.n251 a_n7636_8799.n250 48.2005
R14946 a_n7636_8799.n279 a_n7636_8799.n278 48.2005
R14947 a_n7636_8799.n89 a_n7636_8799.n276 20.9683
R14948 a_n7636_8799.n275 a_n7636_8799.n274 48.2005
R14949 a_n7636_8799.n94 a_n7636_8799.n272 20.9683
R14950 a_n7636_8799.n271 a_n7636_8799.n270 48.2005
R14951 a_n7636_8799.n172 a_n7636_8799.n171 48.2005
R14952 a_n7636_8799.n174 a_n7636_8799.n103 20.9683
R14953 a_n7636_8799.n176 a_n7636_8799.n166 48.2005
R14954 a_n7636_8799.n178 a_n7636_8799.n108 20.9683
R14955 a_n7636_8799.n181 a_n7636_8799.n180 48.2005
R14956 a_n7636_8799.t46 a_n7636_8799.n113 485.135
R14957 a_n7636_8799.n191 a_n7636_8799.n190 48.2005
R14958 a_n7636_8799.n193 a_n7636_8799.n118 20.9683
R14959 a_n7636_8799.n195 a_n7636_8799.n185 48.2005
R14960 a_n7636_8799.n197 a_n7636_8799.n123 20.9683
R14961 a_n7636_8799.n200 a_n7636_8799.n199 48.2005
R14962 a_n7636_8799.t61 a_n7636_8799.n128 485.135
R14963 a_n7636_8799.n211 a_n7636_8799.n210 48.2005
R14964 a_n7636_8799.n213 a_n7636_8799.n133 20.9683
R14965 a_n7636_8799.n215 a_n7636_8799.n205 48.2005
R14966 a_n7636_8799.n217 a_n7636_8799.n138 20.9683
R14967 a_n7636_8799.n220 a_n7636_8799.n219 48.2005
R14968 a_n7636_8799.t155 a_n7636_8799.n143 485.135
R14969 a_n7636_8799.n55 a_n7636_8799.n223 17.8606
R14970 a_n7636_8799.n230 a_n7636_8799.n68 25.894
R14971 a_n7636_8799.n70 a_n7636_8799.n242 17.8606
R14972 a_n7636_8799.n249 a_n7636_8799.n83 25.894
R14973 a_n7636_8799.n85 a_n7636_8799.n262 17.8606
R14974 a_n7636_8799.n269 a_n7636_8799.n98 25.894
R14975 a_n7636_8799.n182 a_n7636_8799.n112 25.894
R14976 a_n7636_8799.n201 a_n7636_8799.n127 25.894
R14977 a_n7636_8799.n221 a_n7636_8799.n142 25.894
R14978 a_n7636_8799.n66 a_n7636_8799.n227 43.3183
R14979 a_n7636_8799.n81 a_n7636_8799.n246 43.3183
R14980 a_n7636_8799.n96 a_n7636_8799.n266 43.3183
R14981 a_n7636_8799.n179 a_n7636_8799.n110 43.3183
R14982 a_n7636_8799.n198 a_n7636_8799.n125 43.3183
R14983 a_n7636_8799.n218 a_n7636_8799.n140 43.3183
R14984 a_n7636_8799.n60 a_n7636_8799.n225 16.6962
R14985 a_n7636_8799.n234 a_n7636_8799.n63 27.6507
R14986 a_n7636_8799.n75 a_n7636_8799.n244 16.6962
R14987 a_n7636_8799.n253 a_n7636_8799.n78 27.6507
R14988 a_n7636_8799.n90 a_n7636_8799.n264 16.6962
R14989 a_n7636_8799.n273 a_n7636_8799.n93 27.6507
R14990 a_n7636_8799.n175 a_n7636_8799.n104 16.6962
R14991 a_n7636_8799.n165 a_n7636_8799.n107 27.6507
R14992 a_n7636_8799.n194 a_n7636_8799.n119 16.6962
R14993 a_n7636_8799.n184 a_n7636_8799.n122 27.6507
R14994 a_n7636_8799.n214 a_n7636_8799.n134 16.6962
R14995 a_n7636_8799.n204 a_n7636_8799.n137 27.6507
R14996 a_n7636_8799.n61 a_n7636_8799.n225 41.7634
R14997 a_n7636_8799.n76 a_n7636_8799.n244 41.7634
R14998 a_n7636_8799.n91 a_n7636_8799.n264 41.7634
R14999 a_n7636_8799.n105 a_n7636_8799.n175 41.7634
R15000 a_n7636_8799.n120 a_n7636_8799.n194 41.7634
R15001 a_n7636_8799.n135 a_n7636_8799.n214 41.7634
R15002 a_n7636_8799.n238 a_n7636_8799.n58 29.3885
R15003 a_n7636_8799.n65 a_n7636_8799.n227 15.5127
R15004 a_n7636_8799.n257 a_n7636_8799.n73 29.3885
R15005 a_n7636_8799.n80 a_n7636_8799.n246 15.5127
R15006 a_n7636_8799.n277 a_n7636_8799.n88 29.3885
R15007 a_n7636_8799.n95 a_n7636_8799.n266 15.5127
R15008 a_n7636_8799.n173 a_n7636_8799.n102 29.3885
R15009 a_n7636_8799.n179 a_n7636_8799.n109 15.5127
R15010 a_n7636_8799.n192 a_n7636_8799.n117 29.3885
R15011 a_n7636_8799.n198 a_n7636_8799.n124 15.5127
R15012 a_n7636_8799.n212 a_n7636_8799.n132 29.3885
R15013 a_n7636_8799.n218 a_n7636_8799.n139 15.5127
R15014 a_n7636_8799.n160 a_n7636_8799.n51 34.3237
R15015 a_n7636_8799.n56 a_n7636_8799.n223 40.1848
R15016 a_n7636_8799.n71 a_n7636_8799.n242 40.1848
R15017 a_n7636_8799.n86 a_n7636_8799.n262 40.1848
R15018 a_n7636_8799.n170 a_n7636_8799.n100 40.1848
R15019 a_n7636_8799.n189 a_n7636_8799.n115 40.1848
R15020 a_n7636_8799.n209 a_n7636_8799.n130 40.1848
R15021 a_n7636_8799.n230 a_n7636_8799.n229 20.9576
R15022 a_n7636_8799.n249 a_n7636_8799.n248 20.9576
R15023 a_n7636_8799.n269 a_n7636_8799.n268 20.9576
R15024 a_n7636_8799.n169 a_n7636_8799.n168 20.9576
R15025 a_n7636_8799.n188 a_n7636_8799.n187 20.9576
R15026 a_n7636_8799.n208 a_n7636_8799.n207 20.9576
R15027 a_n7636_8799.n56 a_n7636_8799.n240 7.32118
R15028 a_n7636_8799.n67 a_n7636_8799.n228 40.1848
R15029 a_n7636_8799.n71 a_n7636_8799.n259 7.32118
R15030 a_n7636_8799.n82 a_n7636_8799.n247 40.1848
R15031 a_n7636_8799.n86 a_n7636_8799.n279 7.32118
R15032 a_n7636_8799.n97 a_n7636_8799.n267 40.1848
R15033 a_n7636_8799.n171 a_n7636_8799.n100 7.32118
R15034 a_n7636_8799.n164 a_n7636_8799.n111 40.1848
R15035 a_n7636_8799.n190 a_n7636_8799.n115 7.32118
R15036 a_n7636_8799.n183 a_n7636_8799.n126 40.1848
R15037 a_n7636_8799.n210 a_n7636_8799.n130 7.32118
R15038 a_n7636_8799.n203 a_n7636_8799.n141 40.1848
R15039 a_n7636_8799.n233 a_n7636_8799.n65 29.3885
R15040 a_n7636_8799.n252 a_n7636_8799.n80 29.3885
R15041 a_n7636_8799.n272 a_n7636_8799.n95 29.3885
R15042 a_n7636_8799.n109 a_n7636_8799.n178 29.3885
R15043 a_n7636_8799.n124 a_n7636_8799.n197 29.3885
R15044 a_n7636_8799.n139 a_n7636_8799.n217 29.3885
R15045 a_n7636_8799.n61 a_n7636_8799.n236 5.97853
R15046 a_n7636_8799.n62 a_n7636_8799.n226 41.7634
R15047 a_n7636_8799.n76 a_n7636_8799.n255 5.97853
R15048 a_n7636_8799.n77 a_n7636_8799.n245 41.7634
R15049 a_n7636_8799.n91 a_n7636_8799.n275 5.97853
R15050 a_n7636_8799.n92 a_n7636_8799.n265 41.7634
R15051 a_n7636_8799.n176 a_n7636_8799.n105 5.97853
R15052 a_n7636_8799.n177 a_n7636_8799.n106 41.7634
R15053 a_n7636_8799.n195 a_n7636_8799.n120 5.97853
R15054 a_n7636_8799.n196 a_n7636_8799.n121 41.7634
R15055 a_n7636_8799.n215 a_n7636_8799.n135 5.97853
R15056 a_n7636_8799.n216 a_n7636_8799.n136 41.7634
R15057 a_n7636_8799.n283 a_n7636_8799.n53 12.3339
R15058 a_n7636_8799.n284 a_n7636_8799.n283 11.4887
R15059 a_n7636_8799.n237 a_n7636_8799.n60 27.6507
R15060 a_n7636_8799.n256 a_n7636_8799.n75 27.6507
R15061 a_n7636_8799.n276 a_n7636_8799.n90 27.6507
R15062 a_n7636_8799.n174 a_n7636_8799.n104 27.6507
R15063 a_n7636_8799.n193 a_n7636_8799.n119 27.6507
R15064 a_n7636_8799.n213 a_n7636_8799.n134 27.6507
R15065 a_n7636_8799.n57 a_n7636_8799.n224 43.3183
R15066 a_n7636_8799.n66 a_n7636_8799.n232 4.61226
R15067 a_n7636_8799.n72 a_n7636_8799.n243 43.3183
R15068 a_n7636_8799.n81 a_n7636_8799.n251 4.61226
R15069 a_n7636_8799.n87 a_n7636_8799.n263 43.3183
R15070 a_n7636_8799.n96 a_n7636_8799.n271 4.61226
R15071 a_n7636_8799.n167 a_n7636_8799.n101 43.3183
R15072 a_n7636_8799.n180 a_n7636_8799.n110 4.61226
R15073 a_n7636_8799.n186 a_n7636_8799.n116 43.3183
R15074 a_n7636_8799.n199 a_n7636_8799.n125 4.61226
R15075 a_n7636_8799.n206 a_n7636_8799.n131 43.3183
R15076 a_n7636_8799.n49 a_n7636_8799.n284 31.5519
R15077 a_n7636_8799.n219 a_n7636_8799.n140 4.61226
R15078 a_n7636_8799.n261 a_n7636_8799.n47 9.04406
R15079 a_n7636_8799.n202 a_n7636_8799.n17 9.04406
R15080 a_n7636_8799.n241 a_n7636_8799.n55 25.894
R15081 a_n7636_8799.n260 a_n7636_8799.n70 25.894
R15082 a_n7636_8799.n280 a_n7636_8799.n85 25.894
R15083 a_n7636_8799.n99 a_n7636_8799.n169 25.894
R15084 a_n7636_8799.n114 a_n7636_8799.n188 25.894
R15085 a_n7636_8799.n129 a_n7636_8799.n208 25.894
R15086 a_n7636_8799.n284 a_n7636_8799.n48 17.6132
R15087 a_n7636_8799.n282 a_n7636_8799.n222 6.93972
R15088 a_n7636_8799.n282 a_n7636_8799.n281 6.44309
R15089 a_n7636_8799.n261 a_n7636_8799.n39 4.93611
R15090 a_n7636_8799.n281 a_n7636_8799.n31 4.93611
R15091 a_n7636_8799.n202 a_n7636_8799.n9 4.93611
R15092 a_n7636_8799.n222 a_n7636_8799.n1 4.93611
R15093 a_n7636_8799.n281 a_n7636_8799.n261 4.10845
R15094 a_n7636_8799.n222 a_n7636_8799.n202 4.10845
R15095 a_n7636_8799.n286 a_n7636_8799.t18 3.61217
R15096 a_n7636_8799.n286 a_n7636_8799.t21 3.61217
R15097 a_n7636_8799.n285 a_n7636_8799.t12 3.61217
R15098 a_n7636_8799.n285 a_n7636_8799.t13 3.61217
R15099 a_n7636_8799.n146 a_n7636_8799.t5 3.61217
R15100 a_n7636_8799.n146 a_n7636_8799.t14 3.61217
R15101 a_n7636_8799.n145 a_n7636_8799.t27 3.61217
R15102 a_n7636_8799.n145 a_n7636_8799.t4 3.61217
R15103 a_n7636_8799.n144 a_n7636_8799.t17 3.61217
R15104 a_n7636_8799.n144 a_n7636_8799.t25 3.61217
R15105 a_n7636_8799.t3 a_n7636_8799.n287 3.61217
R15106 a_n7636_8799.n287 a_n7636_8799.t19 3.61217
R15107 a_n7636_8799.n283 a_n7636_8799.n282 3.4105
R15108 a_n7636_8799.n159 a_n7636_8799.t30 2.82907
R15109 a_n7636_8799.n159 a_n7636_8799.t23 2.82907
R15110 a_n7636_8799.n161 a_n7636_8799.t9 2.82907
R15111 a_n7636_8799.n161 a_n7636_8799.t1 2.82907
R15112 a_n7636_8799.n163 a_n7636_8799.t20 2.82907
R15113 a_n7636_8799.n163 a_n7636_8799.t0 2.82907
R15114 a_n7636_8799.n150 a_n7636_8799.t22 2.82907
R15115 a_n7636_8799.n150 a_n7636_8799.t8 2.82907
R15116 a_n7636_8799.n148 a_n7636_8799.t6 2.82907
R15117 a_n7636_8799.n148 a_n7636_8799.t28 2.82907
R15118 a_n7636_8799.n147 a_n7636_8799.t32 2.82907
R15119 a_n7636_8799.n147 a_n7636_8799.t33 2.82907
R15120 a_n7636_8799.n155 a_n7636_8799.t26 2.82907
R15121 a_n7636_8799.n155 a_n7636_8799.t35 2.82907
R15122 a_n7636_8799.n156 a_n7636_8799.t16 2.82907
R15123 a_n7636_8799.n156 a_n7636_8799.t10 2.82907
R15124 a_n7636_8799.n158 a_n7636_8799.t29 2.82907
R15125 a_n7636_8799.n158 a_n7636_8799.t11 2.82907
R15126 a_n7636_8799.n154 a_n7636_8799.t7 2.82907
R15127 a_n7636_8799.n154 a_n7636_8799.t31 2.82907
R15128 a_n7636_8799.n152 a_n7636_8799.t15 2.82907
R15129 a_n7636_8799.n152 a_n7636_8799.t34 2.82907
R15130 a_n7636_8799.n151 a_n7636_8799.t24 2.82907
R15131 a_n7636_8799.n151 a_n7636_8799.t2 2.82907
R15132 a_n7636_8799.n41 a_n7636_8799.n40 1.13686
R15133 a_n7636_8799.n33 a_n7636_8799.n32 1.13686
R15134 a_n7636_8799.n25 a_n7636_8799.n24 1.13686
R15135 a_n7636_8799.n17 a_n7636_8799.n16 1.13686
R15136 a_n7636_8799.n9 a_n7636_8799.n8 1.13686
R15137 a_n7636_8799.n1 a_n7636_8799.n0 1.13686
R15138 a_n7636_8799.n46 a_n7636_8799.n45 0.758076
R15139 a_n7636_8799.n46 a_n7636_8799.n44 0.758076
R15140 a_n7636_8799.n44 a_n7636_8799.n43 0.758076
R15141 a_n7636_8799.n43 a_n7636_8799.n42 0.758076
R15142 a_n7636_8799.n40 a_n7636_8799.n42 0.758076
R15143 a_n7636_8799.n38 a_n7636_8799.n37 0.758076
R15144 a_n7636_8799.n38 a_n7636_8799.n36 0.758076
R15145 a_n7636_8799.n36 a_n7636_8799.n35 0.758076
R15146 a_n7636_8799.n35 a_n7636_8799.n34 0.758076
R15147 a_n7636_8799.n32 a_n7636_8799.n34 0.758076
R15148 a_n7636_8799.n30 a_n7636_8799.n29 0.758076
R15149 a_n7636_8799.n30 a_n7636_8799.n28 0.758076
R15150 a_n7636_8799.n28 a_n7636_8799.n27 0.758076
R15151 a_n7636_8799.n27 a_n7636_8799.n26 0.758076
R15152 a_n7636_8799.n24 a_n7636_8799.n26 0.758076
R15153 a_n7636_8799.n21 a_n7636_8799.n22 0.758076
R15154 a_n7636_8799.n20 a_n7636_8799.n21 0.758076
R15155 a_n7636_8799.n19 a_n7636_8799.n20 0.758076
R15156 a_n7636_8799.n18 a_n7636_8799.n19 0.758076
R15157 a_n7636_8799.n16 a_n7636_8799.n18 0.758076
R15158 a_n7636_8799.n13 a_n7636_8799.n14 0.758076
R15159 a_n7636_8799.n12 a_n7636_8799.n13 0.758076
R15160 a_n7636_8799.n11 a_n7636_8799.n12 0.758076
R15161 a_n7636_8799.n10 a_n7636_8799.n11 0.758076
R15162 a_n7636_8799.n8 a_n7636_8799.n10 0.758076
R15163 a_n7636_8799.n5 a_n7636_8799.n6 0.758076
R15164 a_n7636_8799.n4 a_n7636_8799.n5 0.758076
R15165 a_n7636_8799.n3 a_n7636_8799.n4 0.758076
R15166 a_n7636_8799.n2 a_n7636_8799.n3 0.758076
R15167 a_n7636_8799.n0 a_n7636_8799.n2 0.758076
R15168 a_n7636_8799.n6 a_n7636_8799.n7 0.568682
R15169 a_n7636_8799.n14 a_n7636_8799.n15 0.568682
R15170 a_n7636_8799.n22 a_n7636_8799.n23 0.568682
R15171 a_n7636_8799.n29 a_n7636_8799.n31 0.568682
R15172 a_n7636_8799.n37 a_n7636_8799.n39 0.568682
R15173 a_n7636_8799.n45 a_n7636_8799.n47 0.568682
R15174 a_n7636_8799.n50 a_n7636_8799.n153 0.530672
R15175 a_n7636_8799.n51 a_n7636_8799.n157 0.530672
R15176 a_n7636_8799.n52 a_n7636_8799.n149 0.530672
R15177 a_n7636_8799.n53 a_n7636_8799.n162 0.530672
R15178 a_n7636_8799.n162 a_n7636_8799.n160 0.530672
R15179 a_n7636_8799.n53 a_n7636_8799.n52 0.530672
R15180 a_n7636_8799.n51 a_n7636_8799.n50 0.530672
R15181 vdd.n327 vdd.n291 756.745
R15182 vdd.n268 vdd.n232 756.745
R15183 vdd.n225 vdd.n189 756.745
R15184 vdd.n166 vdd.n130 756.745
R15185 vdd.n124 vdd.n88 756.745
R15186 vdd.n65 vdd.n29 756.745
R15187 vdd.n1746 vdd.n1710 756.745
R15188 vdd.n1805 vdd.n1769 756.745
R15189 vdd.n1644 vdd.n1608 756.745
R15190 vdd.n1703 vdd.n1667 756.745
R15191 vdd.n1543 vdd.n1507 756.745
R15192 vdd.n1602 vdd.n1566 756.745
R15193 vdd.n2177 vdd.t84 640.208
R15194 vdd.n965 vdd.t69 640.208
R15195 vdd.n2151 vdd.t107 640.208
R15196 vdd.n957 vdd.t95 640.208
R15197 vdd.n2922 vdd.t45 640.208
R15198 vdd.n2642 vdd.t92 640.208
R15199 vdd.n832 vdd.t73 640.208
R15200 vdd.n2639 vdd.t77 640.208
R15201 vdd.n799 vdd.t81 640.208
R15202 vdd.n1027 vdd.t88 640.208
R15203 vdd.n1317 vdd.t60 592.009
R15204 vdd.n1355 vdd.t49 592.009
R15205 vdd.n1251 vdd.t63 592.009
R15206 vdd.n2333 vdd.t41 592.009
R15207 vdd.n1970 vdd.t53 592.009
R15208 vdd.n1930 vdd.t66 592.009
R15209 vdd.n426 vdd.t56 592.009
R15210 vdd.n440 vdd.t98 592.009
R15211 vdd.n452 vdd.t104 592.009
R15212 vdd.n768 vdd.t34 592.009
R15213 vdd.n3184 vdd.t38 592.009
R15214 vdd.n688 vdd.t101 592.009
R15215 vdd.n328 vdd.n327 585
R15216 vdd.n326 vdd.n293 585
R15217 vdd.n325 vdd.n324 585
R15218 vdd.n296 vdd.n294 585
R15219 vdd.n319 vdd.n318 585
R15220 vdd.n317 vdd.n316 585
R15221 vdd.n300 vdd.n299 585
R15222 vdd.n311 vdd.n310 585
R15223 vdd.n309 vdd.n308 585
R15224 vdd.n304 vdd.n303 585
R15225 vdd.n269 vdd.n268 585
R15226 vdd.n267 vdd.n234 585
R15227 vdd.n266 vdd.n265 585
R15228 vdd.n237 vdd.n235 585
R15229 vdd.n260 vdd.n259 585
R15230 vdd.n258 vdd.n257 585
R15231 vdd.n241 vdd.n240 585
R15232 vdd.n252 vdd.n251 585
R15233 vdd.n250 vdd.n249 585
R15234 vdd.n245 vdd.n244 585
R15235 vdd.n226 vdd.n225 585
R15236 vdd.n224 vdd.n191 585
R15237 vdd.n223 vdd.n222 585
R15238 vdd.n194 vdd.n192 585
R15239 vdd.n217 vdd.n216 585
R15240 vdd.n215 vdd.n214 585
R15241 vdd.n198 vdd.n197 585
R15242 vdd.n209 vdd.n208 585
R15243 vdd.n207 vdd.n206 585
R15244 vdd.n202 vdd.n201 585
R15245 vdd.n167 vdd.n166 585
R15246 vdd.n165 vdd.n132 585
R15247 vdd.n164 vdd.n163 585
R15248 vdd.n135 vdd.n133 585
R15249 vdd.n158 vdd.n157 585
R15250 vdd.n156 vdd.n155 585
R15251 vdd.n139 vdd.n138 585
R15252 vdd.n150 vdd.n149 585
R15253 vdd.n148 vdd.n147 585
R15254 vdd.n143 vdd.n142 585
R15255 vdd.n125 vdd.n124 585
R15256 vdd.n123 vdd.n90 585
R15257 vdd.n122 vdd.n121 585
R15258 vdd.n93 vdd.n91 585
R15259 vdd.n116 vdd.n115 585
R15260 vdd.n114 vdd.n113 585
R15261 vdd.n97 vdd.n96 585
R15262 vdd.n108 vdd.n107 585
R15263 vdd.n106 vdd.n105 585
R15264 vdd.n101 vdd.n100 585
R15265 vdd.n66 vdd.n65 585
R15266 vdd.n64 vdd.n31 585
R15267 vdd.n63 vdd.n62 585
R15268 vdd.n34 vdd.n32 585
R15269 vdd.n57 vdd.n56 585
R15270 vdd.n55 vdd.n54 585
R15271 vdd.n38 vdd.n37 585
R15272 vdd.n49 vdd.n48 585
R15273 vdd.n47 vdd.n46 585
R15274 vdd.n42 vdd.n41 585
R15275 vdd.n1747 vdd.n1746 585
R15276 vdd.n1745 vdd.n1712 585
R15277 vdd.n1744 vdd.n1743 585
R15278 vdd.n1715 vdd.n1713 585
R15279 vdd.n1738 vdd.n1737 585
R15280 vdd.n1736 vdd.n1735 585
R15281 vdd.n1719 vdd.n1718 585
R15282 vdd.n1730 vdd.n1729 585
R15283 vdd.n1728 vdd.n1727 585
R15284 vdd.n1723 vdd.n1722 585
R15285 vdd.n1806 vdd.n1805 585
R15286 vdd.n1804 vdd.n1771 585
R15287 vdd.n1803 vdd.n1802 585
R15288 vdd.n1774 vdd.n1772 585
R15289 vdd.n1797 vdd.n1796 585
R15290 vdd.n1795 vdd.n1794 585
R15291 vdd.n1778 vdd.n1777 585
R15292 vdd.n1789 vdd.n1788 585
R15293 vdd.n1787 vdd.n1786 585
R15294 vdd.n1782 vdd.n1781 585
R15295 vdd.n1645 vdd.n1644 585
R15296 vdd.n1643 vdd.n1610 585
R15297 vdd.n1642 vdd.n1641 585
R15298 vdd.n1613 vdd.n1611 585
R15299 vdd.n1636 vdd.n1635 585
R15300 vdd.n1634 vdd.n1633 585
R15301 vdd.n1617 vdd.n1616 585
R15302 vdd.n1628 vdd.n1627 585
R15303 vdd.n1626 vdd.n1625 585
R15304 vdd.n1621 vdd.n1620 585
R15305 vdd.n1704 vdd.n1703 585
R15306 vdd.n1702 vdd.n1669 585
R15307 vdd.n1701 vdd.n1700 585
R15308 vdd.n1672 vdd.n1670 585
R15309 vdd.n1695 vdd.n1694 585
R15310 vdd.n1693 vdd.n1692 585
R15311 vdd.n1676 vdd.n1675 585
R15312 vdd.n1687 vdd.n1686 585
R15313 vdd.n1685 vdd.n1684 585
R15314 vdd.n1680 vdd.n1679 585
R15315 vdd.n1544 vdd.n1543 585
R15316 vdd.n1542 vdd.n1509 585
R15317 vdd.n1541 vdd.n1540 585
R15318 vdd.n1512 vdd.n1510 585
R15319 vdd.n1535 vdd.n1534 585
R15320 vdd.n1533 vdd.n1532 585
R15321 vdd.n1516 vdd.n1515 585
R15322 vdd.n1527 vdd.n1526 585
R15323 vdd.n1525 vdd.n1524 585
R15324 vdd.n1520 vdd.n1519 585
R15325 vdd.n1603 vdd.n1602 585
R15326 vdd.n1601 vdd.n1568 585
R15327 vdd.n1600 vdd.n1599 585
R15328 vdd.n1571 vdd.n1569 585
R15329 vdd.n1594 vdd.n1593 585
R15330 vdd.n1592 vdd.n1591 585
R15331 vdd.n1575 vdd.n1574 585
R15332 vdd.n1586 vdd.n1585 585
R15333 vdd.n1584 vdd.n1583 585
R15334 vdd.n1579 vdd.n1578 585
R15335 vdd.n3356 vdd.n392 509.269
R15336 vdd.n3352 vdd.n393 509.269
R15337 vdd.n3224 vdd.n685 509.269
R15338 vdd.n3221 vdd.n684 509.269
R15339 vdd.n2328 vdd.n1075 509.269
R15340 vdd.n2331 vdd.n2330 509.269
R15341 vdd.n1224 vdd.n1188 509.269
R15342 vdd.n1420 vdd.n1189 509.269
R15343 vdd.n305 vdd.t254 329.043
R15344 vdd.n246 vdd.t226 329.043
R15345 vdd.n203 vdd.t241 329.043
R15346 vdd.n144 vdd.t212 329.043
R15347 vdd.n102 vdd.t190 329.043
R15348 vdd.n43 vdd.t126 329.043
R15349 vdd.n1724 vdd.t272 329.043
R15350 vdd.n1783 vdd.t156 329.043
R15351 vdd.n1622 vdd.t256 329.043
R15352 vdd.n1681 vdd.t130 329.043
R15353 vdd.n1521 vdd.t124 329.043
R15354 vdd.n1580 vdd.t192 329.043
R15355 vdd.n1317 vdd.t62 319.788
R15356 vdd.n1355 vdd.t52 319.788
R15357 vdd.n1251 vdd.t65 319.788
R15358 vdd.n2333 vdd.t43 319.788
R15359 vdd.n1970 vdd.t54 319.788
R15360 vdd.n1930 vdd.t67 319.788
R15361 vdd.n426 vdd.t58 319.788
R15362 vdd.n440 vdd.t99 319.788
R15363 vdd.n452 vdd.t105 319.788
R15364 vdd.n768 vdd.t37 319.788
R15365 vdd.n3184 vdd.t40 319.788
R15366 vdd.n688 vdd.t103 319.788
R15367 vdd.n1318 vdd.t61 303.69
R15368 vdd.n1356 vdd.t51 303.69
R15369 vdd.n1252 vdd.t64 303.69
R15370 vdd.n2334 vdd.t44 303.69
R15371 vdd.n1971 vdd.t55 303.69
R15372 vdd.n1931 vdd.t68 303.69
R15373 vdd.n427 vdd.t59 303.69
R15374 vdd.n441 vdd.t100 303.69
R15375 vdd.n453 vdd.t106 303.69
R15376 vdd.n769 vdd.t36 303.69
R15377 vdd.n3185 vdd.t39 303.69
R15378 vdd.n689 vdd.t102 303.69
R15379 vdd.n2865 vdd.n913 297.074
R15380 vdd.n3058 vdd.n809 297.074
R15381 vdd.n2995 vdd.n806 297.074
R15382 vdd.n2788 vdd.n914 297.074
R15383 vdd.n2603 vdd.n954 297.074
R15384 vdd.n2534 vdd.n2533 297.074
R15385 vdd.n2280 vdd.n1050 297.074
R15386 vdd.n2376 vdd.n1048 297.074
R15387 vdd.n2974 vdd.n807 297.074
R15388 vdd.n3061 vdd.n3060 297.074
R15389 vdd.n2637 vdd.n915 297.074
R15390 vdd.n2863 vdd.n916 297.074
R15391 vdd.n2531 vdd.n963 297.074
R15392 vdd.n961 vdd.n936 297.074
R15393 vdd.n2217 vdd.n1051 297.074
R15394 vdd.n2374 vdd.n1052 297.074
R15395 vdd.n2976 vdd.n807 185
R15396 vdd.n3059 vdd.n807 185
R15397 vdd.n2978 vdd.n2977 185
R15398 vdd.n2977 vdd.n805 185
R15399 vdd.n2979 vdd.n839 185
R15400 vdd.n2989 vdd.n839 185
R15401 vdd.n2980 vdd.n848 185
R15402 vdd.n848 vdd.n846 185
R15403 vdd.n2982 vdd.n2981 185
R15404 vdd.n2983 vdd.n2982 185
R15405 vdd.n2935 vdd.n847 185
R15406 vdd.n847 vdd.n843 185
R15407 vdd.n2934 vdd.n2933 185
R15408 vdd.n2933 vdd.n2932 185
R15409 vdd.n850 vdd.n849 185
R15410 vdd.n851 vdd.n850 185
R15411 vdd.n2925 vdd.n2924 185
R15412 vdd.n2926 vdd.n2925 185
R15413 vdd.n2921 vdd.n860 185
R15414 vdd.n860 vdd.n857 185
R15415 vdd.n2920 vdd.n2919 185
R15416 vdd.n2919 vdd.n2918 185
R15417 vdd.n862 vdd.n861 185
R15418 vdd.n870 vdd.n862 185
R15419 vdd.n2911 vdd.n2910 185
R15420 vdd.n2912 vdd.n2911 185
R15421 vdd.n2909 vdd.n871 185
R15422 vdd.n2760 vdd.n871 185
R15423 vdd.n2908 vdd.n2907 185
R15424 vdd.n2907 vdd.n2906 185
R15425 vdd.n873 vdd.n872 185
R15426 vdd.n874 vdd.n873 185
R15427 vdd.n2899 vdd.n2898 185
R15428 vdd.n2900 vdd.n2899 185
R15429 vdd.n2897 vdd.n883 185
R15430 vdd.n883 vdd.n880 185
R15431 vdd.n2896 vdd.n2895 185
R15432 vdd.n2895 vdd.n2894 185
R15433 vdd.n885 vdd.n884 185
R15434 vdd.n893 vdd.n885 185
R15435 vdd.n2887 vdd.n2886 185
R15436 vdd.n2888 vdd.n2887 185
R15437 vdd.n2885 vdd.n894 185
R15438 vdd.n900 vdd.n894 185
R15439 vdd.n2884 vdd.n2883 185
R15440 vdd.n2883 vdd.n2882 185
R15441 vdd.n896 vdd.n895 185
R15442 vdd.n897 vdd.n896 185
R15443 vdd.n2875 vdd.n2874 185
R15444 vdd.n2876 vdd.n2875 185
R15445 vdd.n2873 vdd.n906 185
R15446 vdd.n2781 vdd.n906 185
R15447 vdd.n2872 vdd.n2871 185
R15448 vdd.n2871 vdd.n2870 185
R15449 vdd.n908 vdd.n907 185
R15450 vdd.t288 vdd.n908 185
R15451 vdd.n2863 vdd.n2862 185
R15452 vdd.n2864 vdd.n2863 185
R15453 vdd.n2861 vdd.n916 185
R15454 vdd.n2860 vdd.n2859 185
R15455 vdd.n918 vdd.n917 185
R15456 vdd.n2646 vdd.n2645 185
R15457 vdd.n2648 vdd.n2647 185
R15458 vdd.n2650 vdd.n2649 185
R15459 vdd.n2652 vdd.n2651 185
R15460 vdd.n2654 vdd.n2653 185
R15461 vdd.n2656 vdd.n2655 185
R15462 vdd.n2658 vdd.n2657 185
R15463 vdd.n2660 vdd.n2659 185
R15464 vdd.n2662 vdd.n2661 185
R15465 vdd.n2664 vdd.n2663 185
R15466 vdd.n2666 vdd.n2665 185
R15467 vdd.n2668 vdd.n2667 185
R15468 vdd.n2670 vdd.n2669 185
R15469 vdd.n2672 vdd.n2671 185
R15470 vdd.n2674 vdd.n2673 185
R15471 vdd.n2676 vdd.n2675 185
R15472 vdd.n2678 vdd.n2677 185
R15473 vdd.n2680 vdd.n2679 185
R15474 vdd.n2682 vdd.n2681 185
R15475 vdd.n2684 vdd.n2683 185
R15476 vdd.n2686 vdd.n2685 185
R15477 vdd.n2688 vdd.n2687 185
R15478 vdd.n2690 vdd.n2689 185
R15479 vdd.n2692 vdd.n2691 185
R15480 vdd.n2694 vdd.n2693 185
R15481 vdd.n2696 vdd.n2695 185
R15482 vdd.n2698 vdd.n2697 185
R15483 vdd.n2700 vdd.n2699 185
R15484 vdd.n2702 vdd.n2701 185
R15485 vdd.n2704 vdd.n2703 185
R15486 vdd.n2706 vdd.n2705 185
R15487 vdd.n2707 vdd.n2637 185
R15488 vdd.n2857 vdd.n2637 185
R15489 vdd.n3062 vdd.n3061 185
R15490 vdd.n3063 vdd.n798 185
R15491 vdd.n3065 vdd.n3064 185
R15492 vdd.n3067 vdd.n796 185
R15493 vdd.n3069 vdd.n3068 185
R15494 vdd.n3070 vdd.n795 185
R15495 vdd.n3072 vdd.n3071 185
R15496 vdd.n3074 vdd.n793 185
R15497 vdd.n3076 vdd.n3075 185
R15498 vdd.n3077 vdd.n792 185
R15499 vdd.n3079 vdd.n3078 185
R15500 vdd.n3081 vdd.n790 185
R15501 vdd.n3083 vdd.n3082 185
R15502 vdd.n3084 vdd.n789 185
R15503 vdd.n3086 vdd.n3085 185
R15504 vdd.n3088 vdd.n788 185
R15505 vdd.n3089 vdd.n786 185
R15506 vdd.n3092 vdd.n3091 185
R15507 vdd.n787 vdd.n785 185
R15508 vdd.n2948 vdd.n2947 185
R15509 vdd.n2950 vdd.n2949 185
R15510 vdd.n2952 vdd.n2944 185
R15511 vdd.n2954 vdd.n2953 185
R15512 vdd.n2955 vdd.n2943 185
R15513 vdd.n2957 vdd.n2956 185
R15514 vdd.n2959 vdd.n2941 185
R15515 vdd.n2961 vdd.n2960 185
R15516 vdd.n2962 vdd.n2940 185
R15517 vdd.n2964 vdd.n2963 185
R15518 vdd.n2966 vdd.n2938 185
R15519 vdd.n2968 vdd.n2967 185
R15520 vdd.n2969 vdd.n2937 185
R15521 vdd.n2971 vdd.n2970 185
R15522 vdd.n2973 vdd.n2936 185
R15523 vdd.n2975 vdd.n2974 185
R15524 vdd.n2974 vdd.n692 185
R15525 vdd.n3060 vdd.n802 185
R15526 vdd.n3060 vdd.n3059 185
R15527 vdd.n2712 vdd.n804 185
R15528 vdd.n805 vdd.n804 185
R15529 vdd.n2713 vdd.n838 185
R15530 vdd.n2989 vdd.n838 185
R15531 vdd.n2715 vdd.n2714 185
R15532 vdd.n2714 vdd.n846 185
R15533 vdd.n2716 vdd.n845 185
R15534 vdd.n2983 vdd.n845 185
R15535 vdd.n2718 vdd.n2717 185
R15536 vdd.n2717 vdd.n843 185
R15537 vdd.n2719 vdd.n853 185
R15538 vdd.n2932 vdd.n853 185
R15539 vdd.n2721 vdd.n2720 185
R15540 vdd.n2720 vdd.n851 185
R15541 vdd.n2722 vdd.n859 185
R15542 vdd.n2926 vdd.n859 185
R15543 vdd.n2724 vdd.n2723 185
R15544 vdd.n2723 vdd.n857 185
R15545 vdd.n2725 vdd.n864 185
R15546 vdd.n2918 vdd.n864 185
R15547 vdd.n2727 vdd.n2726 185
R15548 vdd.n2726 vdd.n870 185
R15549 vdd.n2728 vdd.n869 185
R15550 vdd.n2912 vdd.n869 185
R15551 vdd.n2762 vdd.n2761 185
R15552 vdd.n2761 vdd.n2760 185
R15553 vdd.n2763 vdd.n876 185
R15554 vdd.n2906 vdd.n876 185
R15555 vdd.n2765 vdd.n2764 185
R15556 vdd.n2764 vdd.n874 185
R15557 vdd.n2766 vdd.n882 185
R15558 vdd.n2900 vdd.n882 185
R15559 vdd.n2768 vdd.n2767 185
R15560 vdd.n2767 vdd.n880 185
R15561 vdd.n2769 vdd.n887 185
R15562 vdd.n2894 vdd.n887 185
R15563 vdd.n2771 vdd.n2770 185
R15564 vdd.n2770 vdd.n893 185
R15565 vdd.n2772 vdd.n892 185
R15566 vdd.n2888 vdd.n892 185
R15567 vdd.n2774 vdd.n2773 185
R15568 vdd.n2773 vdd.n900 185
R15569 vdd.n2775 vdd.n899 185
R15570 vdd.n2882 vdd.n899 185
R15571 vdd.n2777 vdd.n2776 185
R15572 vdd.n2776 vdd.n897 185
R15573 vdd.n2778 vdd.n905 185
R15574 vdd.n2876 vdd.n905 185
R15575 vdd.n2780 vdd.n2779 185
R15576 vdd.n2781 vdd.n2780 185
R15577 vdd.n2711 vdd.n910 185
R15578 vdd.n2870 vdd.n910 185
R15579 vdd.n2710 vdd.n2709 185
R15580 vdd.n2709 vdd.t288 185
R15581 vdd.n2708 vdd.n915 185
R15582 vdd.n2864 vdd.n915 185
R15583 vdd.n2328 vdd.n2327 185
R15584 vdd.n2329 vdd.n2328 185
R15585 vdd.n1076 vdd.n1074 185
R15586 vdd.n1894 vdd.n1074 185
R15587 vdd.n1897 vdd.n1896 185
R15588 vdd.n1896 vdd.n1895 185
R15589 vdd.n1079 vdd.n1078 185
R15590 vdd.n1080 vdd.n1079 185
R15591 vdd.n1883 vdd.n1882 185
R15592 vdd.n1884 vdd.n1883 185
R15593 vdd.n1088 vdd.n1087 185
R15594 vdd.n1875 vdd.n1087 185
R15595 vdd.n1878 vdd.n1877 185
R15596 vdd.n1877 vdd.n1876 185
R15597 vdd.n1091 vdd.n1090 185
R15598 vdd.n1098 vdd.n1091 185
R15599 vdd.n1866 vdd.n1865 185
R15600 vdd.n1867 vdd.n1866 185
R15601 vdd.n1100 vdd.n1099 185
R15602 vdd.n1099 vdd.n1097 185
R15603 vdd.n1861 vdd.n1860 185
R15604 vdd.n1860 vdd.n1859 185
R15605 vdd.n1103 vdd.n1102 185
R15606 vdd.n1104 vdd.n1103 185
R15607 vdd.n1850 vdd.n1849 185
R15608 vdd.n1851 vdd.n1850 185
R15609 vdd.n1111 vdd.n1110 185
R15610 vdd.n1842 vdd.n1110 185
R15611 vdd.n1845 vdd.n1844 185
R15612 vdd.n1844 vdd.n1843 185
R15613 vdd.n1114 vdd.n1113 185
R15614 vdd.n1120 vdd.n1114 185
R15615 vdd.n1833 vdd.n1832 185
R15616 vdd.n1834 vdd.n1833 185
R15617 vdd.n1122 vdd.n1121 185
R15618 vdd.n1825 vdd.n1121 185
R15619 vdd.n1828 vdd.n1827 185
R15620 vdd.n1827 vdd.n1826 185
R15621 vdd.n1125 vdd.n1124 185
R15622 vdd.n1126 vdd.n1125 185
R15623 vdd.n1816 vdd.n1815 185
R15624 vdd.n1817 vdd.n1816 185
R15625 vdd.n1134 vdd.n1133 185
R15626 vdd.n1133 vdd.n1132 185
R15627 vdd.n1504 vdd.n1503 185
R15628 vdd.n1503 vdd.n1502 185
R15629 vdd.n1137 vdd.n1136 185
R15630 vdd.n1143 vdd.n1137 185
R15631 vdd.n1493 vdd.n1492 185
R15632 vdd.n1494 vdd.n1493 185
R15633 vdd.n1145 vdd.n1144 185
R15634 vdd.n1485 vdd.n1144 185
R15635 vdd.n1488 vdd.n1487 185
R15636 vdd.n1487 vdd.n1486 185
R15637 vdd.n1148 vdd.n1147 185
R15638 vdd.n1155 vdd.n1148 185
R15639 vdd.n1476 vdd.n1475 185
R15640 vdd.n1477 vdd.n1476 185
R15641 vdd.n1157 vdd.n1156 185
R15642 vdd.n1156 vdd.n1154 185
R15643 vdd.n1471 vdd.n1470 185
R15644 vdd.n1470 vdd.n1469 185
R15645 vdd.n1160 vdd.n1159 185
R15646 vdd.n1161 vdd.n1160 185
R15647 vdd.n1460 vdd.n1459 185
R15648 vdd.n1461 vdd.n1460 185
R15649 vdd.n1168 vdd.n1167 185
R15650 vdd.n1452 vdd.n1167 185
R15651 vdd.n1455 vdd.n1454 185
R15652 vdd.n1454 vdd.n1453 185
R15653 vdd.n1171 vdd.n1170 185
R15654 vdd.n1177 vdd.n1171 185
R15655 vdd.n1443 vdd.n1442 185
R15656 vdd.n1444 vdd.n1443 185
R15657 vdd.n1179 vdd.n1178 185
R15658 vdd.n1435 vdd.n1178 185
R15659 vdd.n1438 vdd.n1437 185
R15660 vdd.n1437 vdd.n1436 185
R15661 vdd.n1182 vdd.n1181 185
R15662 vdd.n1183 vdd.n1182 185
R15663 vdd.n1426 vdd.n1425 185
R15664 vdd.n1427 vdd.n1426 185
R15665 vdd.n1190 vdd.n1189 185
R15666 vdd.n1225 vdd.n1189 185
R15667 vdd.n1421 vdd.n1420 185
R15668 vdd.n1193 vdd.n1192 185
R15669 vdd.n1417 vdd.n1416 185
R15670 vdd.n1418 vdd.n1417 185
R15671 vdd.n1227 vdd.n1226 185
R15672 vdd.n1412 vdd.n1229 185
R15673 vdd.n1411 vdd.n1230 185
R15674 vdd.n1410 vdd.n1231 185
R15675 vdd.n1233 vdd.n1232 185
R15676 vdd.n1406 vdd.n1235 185
R15677 vdd.n1405 vdd.n1236 185
R15678 vdd.n1404 vdd.n1237 185
R15679 vdd.n1239 vdd.n1238 185
R15680 vdd.n1400 vdd.n1241 185
R15681 vdd.n1399 vdd.n1242 185
R15682 vdd.n1398 vdd.n1243 185
R15683 vdd.n1245 vdd.n1244 185
R15684 vdd.n1394 vdd.n1247 185
R15685 vdd.n1393 vdd.n1248 185
R15686 vdd.n1392 vdd.n1249 185
R15687 vdd.n1253 vdd.n1250 185
R15688 vdd.n1388 vdd.n1255 185
R15689 vdd.n1387 vdd.n1256 185
R15690 vdd.n1386 vdd.n1257 185
R15691 vdd.n1259 vdd.n1258 185
R15692 vdd.n1382 vdd.n1261 185
R15693 vdd.n1381 vdd.n1262 185
R15694 vdd.n1380 vdd.n1263 185
R15695 vdd.n1265 vdd.n1264 185
R15696 vdd.n1376 vdd.n1267 185
R15697 vdd.n1375 vdd.n1268 185
R15698 vdd.n1374 vdd.n1269 185
R15699 vdd.n1271 vdd.n1270 185
R15700 vdd.n1370 vdd.n1273 185
R15701 vdd.n1369 vdd.n1274 185
R15702 vdd.n1368 vdd.n1275 185
R15703 vdd.n1277 vdd.n1276 185
R15704 vdd.n1364 vdd.n1279 185
R15705 vdd.n1363 vdd.n1280 185
R15706 vdd.n1362 vdd.n1281 185
R15707 vdd.n1283 vdd.n1282 185
R15708 vdd.n1358 vdd.n1285 185
R15709 vdd.n1357 vdd.n1354 185
R15710 vdd.n1353 vdd.n1286 185
R15711 vdd.n1288 vdd.n1287 185
R15712 vdd.n1349 vdd.n1290 185
R15713 vdd.n1348 vdd.n1291 185
R15714 vdd.n1347 vdd.n1292 185
R15715 vdd.n1294 vdd.n1293 185
R15716 vdd.n1343 vdd.n1296 185
R15717 vdd.n1342 vdd.n1297 185
R15718 vdd.n1341 vdd.n1298 185
R15719 vdd.n1300 vdd.n1299 185
R15720 vdd.n1337 vdd.n1302 185
R15721 vdd.n1336 vdd.n1303 185
R15722 vdd.n1335 vdd.n1304 185
R15723 vdd.n1306 vdd.n1305 185
R15724 vdd.n1331 vdd.n1308 185
R15725 vdd.n1330 vdd.n1309 185
R15726 vdd.n1329 vdd.n1310 185
R15727 vdd.n1312 vdd.n1311 185
R15728 vdd.n1325 vdd.n1314 185
R15729 vdd.n1324 vdd.n1315 185
R15730 vdd.n1323 vdd.n1316 185
R15731 vdd.n1320 vdd.n1224 185
R15732 vdd.n1418 vdd.n1224 185
R15733 vdd.n2332 vdd.n2331 185
R15734 vdd.n2336 vdd.n1069 185
R15735 vdd.n1999 vdd.n1068 185
R15736 vdd.n2002 vdd.n2001 185
R15737 vdd.n2004 vdd.n2003 185
R15738 vdd.n2007 vdd.n2006 185
R15739 vdd.n2009 vdd.n2008 185
R15740 vdd.n2011 vdd.n1997 185
R15741 vdd.n2013 vdd.n2012 185
R15742 vdd.n2014 vdd.n1991 185
R15743 vdd.n2016 vdd.n2015 185
R15744 vdd.n2018 vdd.n1989 185
R15745 vdd.n2020 vdd.n2019 185
R15746 vdd.n2021 vdd.n1984 185
R15747 vdd.n2023 vdd.n2022 185
R15748 vdd.n2025 vdd.n1982 185
R15749 vdd.n2027 vdd.n2026 185
R15750 vdd.n2028 vdd.n1978 185
R15751 vdd.n2030 vdd.n2029 185
R15752 vdd.n2032 vdd.n1975 185
R15753 vdd.n2034 vdd.n2033 185
R15754 vdd.n1976 vdd.n1969 185
R15755 vdd.n2038 vdd.n1973 185
R15756 vdd.n2039 vdd.n1965 185
R15757 vdd.n2041 vdd.n2040 185
R15758 vdd.n2043 vdd.n1963 185
R15759 vdd.n2045 vdd.n2044 185
R15760 vdd.n2046 vdd.n1958 185
R15761 vdd.n2048 vdd.n2047 185
R15762 vdd.n2050 vdd.n1956 185
R15763 vdd.n2052 vdd.n2051 185
R15764 vdd.n2053 vdd.n1951 185
R15765 vdd.n2055 vdd.n2054 185
R15766 vdd.n2057 vdd.n1949 185
R15767 vdd.n2059 vdd.n2058 185
R15768 vdd.n2060 vdd.n1944 185
R15769 vdd.n2062 vdd.n2061 185
R15770 vdd.n2064 vdd.n1942 185
R15771 vdd.n2066 vdd.n2065 185
R15772 vdd.n2067 vdd.n1938 185
R15773 vdd.n2069 vdd.n2068 185
R15774 vdd.n2071 vdd.n1935 185
R15775 vdd.n2073 vdd.n2072 185
R15776 vdd.n1936 vdd.n1929 185
R15777 vdd.n2077 vdd.n1933 185
R15778 vdd.n2078 vdd.n1925 185
R15779 vdd.n2080 vdd.n2079 185
R15780 vdd.n2082 vdd.n1923 185
R15781 vdd.n2084 vdd.n2083 185
R15782 vdd.n2085 vdd.n1918 185
R15783 vdd.n2087 vdd.n2086 185
R15784 vdd.n2089 vdd.n1916 185
R15785 vdd.n2091 vdd.n2090 185
R15786 vdd.n2092 vdd.n1911 185
R15787 vdd.n2094 vdd.n2093 185
R15788 vdd.n2096 vdd.n1910 185
R15789 vdd.n2097 vdd.n1907 185
R15790 vdd.n2100 vdd.n2099 185
R15791 vdd.n1909 vdd.n1905 185
R15792 vdd.n2317 vdd.n1903 185
R15793 vdd.n2319 vdd.n2318 185
R15794 vdd.n2321 vdd.n1901 185
R15795 vdd.n2323 vdd.n2322 185
R15796 vdd.n2324 vdd.n1075 185
R15797 vdd.n2330 vdd.n1072 185
R15798 vdd.n2330 vdd.n2329 185
R15799 vdd.n1083 vdd.n1071 185
R15800 vdd.n1894 vdd.n1071 185
R15801 vdd.n1893 vdd.n1892 185
R15802 vdd.n1895 vdd.n1893 185
R15803 vdd.n1082 vdd.n1081 185
R15804 vdd.n1081 vdd.n1080 185
R15805 vdd.n1886 vdd.n1885 185
R15806 vdd.n1885 vdd.n1884 185
R15807 vdd.n1086 vdd.n1085 185
R15808 vdd.n1875 vdd.n1086 185
R15809 vdd.n1874 vdd.n1873 185
R15810 vdd.n1876 vdd.n1874 185
R15811 vdd.n1093 vdd.n1092 185
R15812 vdd.n1098 vdd.n1092 185
R15813 vdd.n1869 vdd.n1868 185
R15814 vdd.n1868 vdd.n1867 185
R15815 vdd.n1096 vdd.n1095 185
R15816 vdd.n1097 vdd.n1096 185
R15817 vdd.n1858 vdd.n1857 185
R15818 vdd.n1859 vdd.n1858 185
R15819 vdd.n1106 vdd.n1105 185
R15820 vdd.n1105 vdd.n1104 185
R15821 vdd.n1853 vdd.n1852 185
R15822 vdd.n1852 vdd.n1851 185
R15823 vdd.n1109 vdd.n1108 185
R15824 vdd.n1842 vdd.n1109 185
R15825 vdd.n1841 vdd.n1840 185
R15826 vdd.n1843 vdd.n1841 185
R15827 vdd.n1116 vdd.n1115 185
R15828 vdd.n1120 vdd.n1115 185
R15829 vdd.n1836 vdd.n1835 185
R15830 vdd.n1835 vdd.n1834 185
R15831 vdd.n1119 vdd.n1118 185
R15832 vdd.n1825 vdd.n1119 185
R15833 vdd.n1824 vdd.n1823 185
R15834 vdd.n1826 vdd.n1824 185
R15835 vdd.n1128 vdd.n1127 185
R15836 vdd.n1127 vdd.n1126 185
R15837 vdd.n1819 vdd.n1818 185
R15838 vdd.n1818 vdd.n1817 185
R15839 vdd.n1131 vdd.n1130 185
R15840 vdd.n1132 vdd.n1131 185
R15841 vdd.n1501 vdd.n1500 185
R15842 vdd.n1502 vdd.n1501 185
R15843 vdd.n1139 vdd.n1138 185
R15844 vdd.n1143 vdd.n1138 185
R15845 vdd.n1496 vdd.n1495 185
R15846 vdd.n1495 vdd.n1494 185
R15847 vdd.n1142 vdd.n1141 185
R15848 vdd.n1485 vdd.n1142 185
R15849 vdd.n1484 vdd.n1483 185
R15850 vdd.n1486 vdd.n1484 185
R15851 vdd.n1150 vdd.n1149 185
R15852 vdd.n1155 vdd.n1149 185
R15853 vdd.n1479 vdd.n1478 185
R15854 vdd.n1478 vdd.n1477 185
R15855 vdd.n1153 vdd.n1152 185
R15856 vdd.n1154 vdd.n1153 185
R15857 vdd.n1468 vdd.n1467 185
R15858 vdd.n1469 vdd.n1468 185
R15859 vdd.n1163 vdd.n1162 185
R15860 vdd.n1162 vdd.n1161 185
R15861 vdd.n1463 vdd.n1462 185
R15862 vdd.n1462 vdd.n1461 185
R15863 vdd.n1166 vdd.n1165 185
R15864 vdd.n1452 vdd.n1166 185
R15865 vdd.n1451 vdd.n1450 185
R15866 vdd.n1453 vdd.n1451 185
R15867 vdd.n1173 vdd.n1172 185
R15868 vdd.n1177 vdd.n1172 185
R15869 vdd.n1446 vdd.n1445 185
R15870 vdd.n1445 vdd.n1444 185
R15871 vdd.n1176 vdd.n1175 185
R15872 vdd.n1435 vdd.n1176 185
R15873 vdd.n1434 vdd.n1433 185
R15874 vdd.n1436 vdd.n1434 185
R15875 vdd.n1185 vdd.n1184 185
R15876 vdd.n1184 vdd.n1183 185
R15877 vdd.n1429 vdd.n1428 185
R15878 vdd.n1428 vdd.n1427 185
R15879 vdd.n1188 vdd.n1187 185
R15880 vdd.n1225 vdd.n1188 185
R15881 vdd.n956 vdd.n954 185
R15882 vdd.n2532 vdd.n954 185
R15883 vdd.n2454 vdd.n973 185
R15884 vdd.n973 vdd.t5 185
R15885 vdd.n2456 vdd.n2455 185
R15886 vdd.n2457 vdd.n2456 185
R15887 vdd.n2453 vdd.n972 185
R15888 vdd.n2156 vdd.n972 185
R15889 vdd.n2452 vdd.n2451 185
R15890 vdd.n2451 vdd.n2450 185
R15891 vdd.n975 vdd.n974 185
R15892 vdd.n976 vdd.n975 185
R15893 vdd.n2441 vdd.n2440 185
R15894 vdd.n2442 vdd.n2441 185
R15895 vdd.n2439 vdd.n986 185
R15896 vdd.n986 vdd.n983 185
R15897 vdd.n2438 vdd.n2437 185
R15898 vdd.n2437 vdd.n2436 185
R15899 vdd.n988 vdd.n987 185
R15900 vdd.n989 vdd.n988 185
R15901 vdd.n2429 vdd.n2428 185
R15902 vdd.n2430 vdd.n2429 185
R15903 vdd.n2427 vdd.n997 185
R15904 vdd.n1002 vdd.n997 185
R15905 vdd.n2426 vdd.n2425 185
R15906 vdd.n2425 vdd.n2424 185
R15907 vdd.n999 vdd.n998 185
R15908 vdd.n1008 vdd.n999 185
R15909 vdd.n2417 vdd.n2416 185
R15910 vdd.n2418 vdd.n2417 185
R15911 vdd.n2415 vdd.n1009 185
R15912 vdd.n2257 vdd.n1009 185
R15913 vdd.n2414 vdd.n2413 185
R15914 vdd.n2413 vdd.n2412 185
R15915 vdd.n1011 vdd.n1010 185
R15916 vdd.n1012 vdd.n1011 185
R15917 vdd.n2405 vdd.n2404 185
R15918 vdd.n2406 vdd.n2405 185
R15919 vdd.n2403 vdd.n1021 185
R15920 vdd.n1021 vdd.n1018 185
R15921 vdd.n2402 vdd.n2401 185
R15922 vdd.n2401 vdd.n2400 185
R15923 vdd.n1023 vdd.n1022 185
R15924 vdd.n1033 vdd.n1023 185
R15925 vdd.n2392 vdd.n2391 185
R15926 vdd.n2393 vdd.n2392 185
R15927 vdd.n2390 vdd.n1034 185
R15928 vdd.n1034 vdd.n1030 185
R15929 vdd.n2389 vdd.n2388 185
R15930 vdd.n2388 vdd.n2387 185
R15931 vdd.n1036 vdd.n1035 185
R15932 vdd.n1037 vdd.n1036 185
R15933 vdd.n2380 vdd.n2379 185
R15934 vdd.n2381 vdd.n2380 185
R15935 vdd.n2378 vdd.n1046 185
R15936 vdd.n1046 vdd.n1043 185
R15937 vdd.n2377 vdd.n2376 185
R15938 vdd.n2376 vdd.n2375 185
R15939 vdd.n1048 vdd.n1047 185
R15940 vdd.n2112 vdd.n2111 185
R15941 vdd.n2113 vdd.n2109 185
R15942 vdd.n2109 vdd.n1049 185
R15943 vdd.n2115 vdd.n2114 185
R15944 vdd.n2117 vdd.n2108 185
R15945 vdd.n2120 vdd.n2119 185
R15946 vdd.n2121 vdd.n2107 185
R15947 vdd.n2123 vdd.n2122 185
R15948 vdd.n2125 vdd.n2106 185
R15949 vdd.n2128 vdd.n2127 185
R15950 vdd.n2129 vdd.n2105 185
R15951 vdd.n2131 vdd.n2130 185
R15952 vdd.n2133 vdd.n2104 185
R15953 vdd.n2136 vdd.n2135 185
R15954 vdd.n2137 vdd.n2103 185
R15955 vdd.n2139 vdd.n2138 185
R15956 vdd.n2141 vdd.n2102 185
R15957 vdd.n2314 vdd.n2142 185
R15958 vdd.n2313 vdd.n2312 185
R15959 vdd.n2310 vdd.n2143 185
R15960 vdd.n2308 vdd.n2307 185
R15961 vdd.n2306 vdd.n2144 185
R15962 vdd.n2305 vdd.n2304 185
R15963 vdd.n2302 vdd.n2145 185
R15964 vdd.n2300 vdd.n2299 185
R15965 vdd.n2298 vdd.n2146 185
R15966 vdd.n2297 vdd.n2296 185
R15967 vdd.n2294 vdd.n2147 185
R15968 vdd.n2292 vdd.n2291 185
R15969 vdd.n2290 vdd.n2148 185
R15970 vdd.n2289 vdd.n2288 185
R15971 vdd.n2286 vdd.n2149 185
R15972 vdd.n2284 vdd.n2283 185
R15973 vdd.n2282 vdd.n2150 185
R15974 vdd.n2281 vdd.n2280 185
R15975 vdd.n2535 vdd.n2534 185
R15976 vdd.n2537 vdd.n2536 185
R15977 vdd.n2539 vdd.n2538 185
R15978 vdd.n2542 vdd.n2541 185
R15979 vdd.n2544 vdd.n2543 185
R15980 vdd.n2546 vdd.n2545 185
R15981 vdd.n2548 vdd.n2547 185
R15982 vdd.n2550 vdd.n2549 185
R15983 vdd.n2552 vdd.n2551 185
R15984 vdd.n2554 vdd.n2553 185
R15985 vdd.n2556 vdd.n2555 185
R15986 vdd.n2558 vdd.n2557 185
R15987 vdd.n2560 vdd.n2559 185
R15988 vdd.n2562 vdd.n2561 185
R15989 vdd.n2564 vdd.n2563 185
R15990 vdd.n2566 vdd.n2565 185
R15991 vdd.n2568 vdd.n2567 185
R15992 vdd.n2570 vdd.n2569 185
R15993 vdd.n2572 vdd.n2571 185
R15994 vdd.n2574 vdd.n2573 185
R15995 vdd.n2576 vdd.n2575 185
R15996 vdd.n2578 vdd.n2577 185
R15997 vdd.n2580 vdd.n2579 185
R15998 vdd.n2582 vdd.n2581 185
R15999 vdd.n2584 vdd.n2583 185
R16000 vdd.n2586 vdd.n2585 185
R16001 vdd.n2588 vdd.n2587 185
R16002 vdd.n2590 vdd.n2589 185
R16003 vdd.n2592 vdd.n2591 185
R16004 vdd.n2594 vdd.n2593 185
R16005 vdd.n2596 vdd.n2595 185
R16006 vdd.n2598 vdd.n2597 185
R16007 vdd.n2600 vdd.n2599 185
R16008 vdd.n2601 vdd.n955 185
R16009 vdd.n2603 vdd.n2602 185
R16010 vdd.n2604 vdd.n2603 185
R16011 vdd.n2533 vdd.n959 185
R16012 vdd.n2533 vdd.n2532 185
R16013 vdd.n2154 vdd.n960 185
R16014 vdd.t5 vdd.n960 185
R16015 vdd.n2155 vdd.n970 185
R16016 vdd.n2457 vdd.n970 185
R16017 vdd.n2158 vdd.n2157 185
R16018 vdd.n2157 vdd.n2156 185
R16019 vdd.n2159 vdd.n977 185
R16020 vdd.n2450 vdd.n977 185
R16021 vdd.n2161 vdd.n2160 185
R16022 vdd.n2160 vdd.n976 185
R16023 vdd.n2162 vdd.n984 185
R16024 vdd.n2442 vdd.n984 185
R16025 vdd.n2164 vdd.n2163 185
R16026 vdd.n2163 vdd.n983 185
R16027 vdd.n2165 vdd.n990 185
R16028 vdd.n2436 vdd.n990 185
R16029 vdd.n2167 vdd.n2166 185
R16030 vdd.n2166 vdd.n989 185
R16031 vdd.n2168 vdd.n995 185
R16032 vdd.n2430 vdd.n995 185
R16033 vdd.n2170 vdd.n2169 185
R16034 vdd.n2169 vdd.n1002 185
R16035 vdd.n2171 vdd.n1000 185
R16036 vdd.n2424 vdd.n1000 185
R16037 vdd.n2173 vdd.n2172 185
R16038 vdd.n2172 vdd.n1008 185
R16039 vdd.n2174 vdd.n1006 185
R16040 vdd.n2418 vdd.n1006 185
R16041 vdd.n2259 vdd.n2258 185
R16042 vdd.n2258 vdd.n2257 185
R16043 vdd.n2260 vdd.n1013 185
R16044 vdd.n2412 vdd.n1013 185
R16045 vdd.n2262 vdd.n2261 185
R16046 vdd.n2261 vdd.n1012 185
R16047 vdd.n2263 vdd.n1019 185
R16048 vdd.n2406 vdd.n1019 185
R16049 vdd.n2265 vdd.n2264 185
R16050 vdd.n2264 vdd.n1018 185
R16051 vdd.n2266 vdd.n1024 185
R16052 vdd.n2400 vdd.n1024 185
R16053 vdd.n2268 vdd.n2267 185
R16054 vdd.n2267 vdd.n1033 185
R16055 vdd.n2269 vdd.n1031 185
R16056 vdd.n2393 vdd.n1031 185
R16057 vdd.n2271 vdd.n2270 185
R16058 vdd.n2270 vdd.n1030 185
R16059 vdd.n2272 vdd.n1038 185
R16060 vdd.n2387 vdd.n1038 185
R16061 vdd.n2274 vdd.n2273 185
R16062 vdd.n2273 vdd.n1037 185
R16063 vdd.n2275 vdd.n1044 185
R16064 vdd.n2381 vdd.n1044 185
R16065 vdd.n2277 vdd.n2276 185
R16066 vdd.n2276 vdd.n1043 185
R16067 vdd.n2278 vdd.n1050 185
R16068 vdd.n2375 vdd.n1050 185
R16069 vdd.n3357 vdd.n3356 185
R16070 vdd.n3356 vdd.n3355 185
R16071 vdd.n3358 vdd.n387 185
R16072 vdd.n387 vdd.n386 185
R16073 vdd.n3360 vdd.n3359 185
R16074 vdd.n3361 vdd.n3360 185
R16075 vdd.n382 vdd.n381 185
R16076 vdd.n3362 vdd.n382 185
R16077 vdd.n3365 vdd.n3364 185
R16078 vdd.n3364 vdd.n3363 185
R16079 vdd.n3366 vdd.n376 185
R16080 vdd.n376 vdd.n375 185
R16081 vdd.n3368 vdd.n3367 185
R16082 vdd.n3369 vdd.n3368 185
R16083 vdd.n371 vdd.n370 185
R16084 vdd.n3370 vdd.n371 185
R16085 vdd.n3373 vdd.n3372 185
R16086 vdd.n3372 vdd.n3371 185
R16087 vdd.n3374 vdd.n365 185
R16088 vdd.n3331 vdd.n365 185
R16089 vdd.n3376 vdd.n3375 185
R16090 vdd.n3377 vdd.n3376 185
R16091 vdd.n360 vdd.n359 185
R16092 vdd.n3378 vdd.n360 185
R16093 vdd.n3381 vdd.n3380 185
R16094 vdd.n3380 vdd.n3379 185
R16095 vdd.n3382 vdd.n354 185
R16096 vdd.n361 vdd.n354 185
R16097 vdd.n3384 vdd.n3383 185
R16098 vdd.n3385 vdd.n3384 185
R16099 vdd.n350 vdd.n349 185
R16100 vdd.n3386 vdd.n350 185
R16101 vdd.n3389 vdd.n3388 185
R16102 vdd.n3388 vdd.n3387 185
R16103 vdd.n3390 vdd.n345 185
R16104 vdd.n345 vdd.n344 185
R16105 vdd.n3392 vdd.n3391 185
R16106 vdd.n3393 vdd.n3392 185
R16107 vdd.n339 vdd.n337 185
R16108 vdd.n3394 vdd.n339 185
R16109 vdd.n3397 vdd.n3396 185
R16110 vdd.n3396 vdd.n3395 185
R16111 vdd.n338 vdd.n336 185
R16112 vdd.n340 vdd.n338 185
R16113 vdd.n3307 vdd.n3306 185
R16114 vdd.n3308 vdd.n3307 185
R16115 vdd.n635 vdd.n634 185
R16116 vdd.n634 vdd.n633 185
R16117 vdd.n3302 vdd.n3301 185
R16118 vdd.n3301 vdd.n3300 185
R16119 vdd.n638 vdd.n637 185
R16120 vdd.n644 vdd.n638 185
R16121 vdd.n3288 vdd.n3287 185
R16122 vdd.n3289 vdd.n3288 185
R16123 vdd.n646 vdd.n645 185
R16124 vdd.n3280 vdd.n645 185
R16125 vdd.n3283 vdd.n3282 185
R16126 vdd.n3282 vdd.n3281 185
R16127 vdd.n649 vdd.n648 185
R16128 vdd.n656 vdd.n649 185
R16129 vdd.n3271 vdd.n3270 185
R16130 vdd.n3272 vdd.n3271 185
R16131 vdd.n658 vdd.n657 185
R16132 vdd.n657 vdd.n655 185
R16133 vdd.n3266 vdd.n3265 185
R16134 vdd.n3265 vdd.n3264 185
R16135 vdd.n661 vdd.n660 185
R16136 vdd.n662 vdd.n661 185
R16137 vdd.n3255 vdd.n3254 185
R16138 vdd.n3256 vdd.n3255 185
R16139 vdd.n669 vdd.n668 185
R16140 vdd.n3247 vdd.n668 185
R16141 vdd.n3250 vdd.n3249 185
R16142 vdd.n3249 vdd.n3248 185
R16143 vdd.n672 vdd.n671 185
R16144 vdd.n679 vdd.n672 185
R16145 vdd.n3238 vdd.n3237 185
R16146 vdd.n3239 vdd.n3238 185
R16147 vdd.n681 vdd.n680 185
R16148 vdd.n680 vdd.n678 185
R16149 vdd.n3233 vdd.n3232 185
R16150 vdd.n3232 vdd.n3231 185
R16151 vdd.n684 vdd.n683 185
R16152 vdd.n723 vdd.n684 185
R16153 vdd.n3221 vdd.n3220 185
R16154 vdd.n3219 vdd.n725 185
R16155 vdd.n3218 vdd.n724 185
R16156 vdd.n3223 vdd.n724 185
R16157 vdd.n729 vdd.n728 185
R16158 vdd.n733 vdd.n732 185
R16159 vdd.n3214 vdd.n734 185
R16160 vdd.n3213 vdd.n3212 185
R16161 vdd.n3211 vdd.n3210 185
R16162 vdd.n3209 vdd.n3208 185
R16163 vdd.n3207 vdd.n3206 185
R16164 vdd.n3205 vdd.n3204 185
R16165 vdd.n3203 vdd.n3202 185
R16166 vdd.n3201 vdd.n3200 185
R16167 vdd.n3199 vdd.n3198 185
R16168 vdd.n3197 vdd.n3196 185
R16169 vdd.n3195 vdd.n3194 185
R16170 vdd.n3193 vdd.n3192 185
R16171 vdd.n3191 vdd.n3190 185
R16172 vdd.n3189 vdd.n3188 185
R16173 vdd.n3187 vdd.n3186 185
R16174 vdd.n3178 vdd.n747 185
R16175 vdd.n3180 vdd.n3179 185
R16176 vdd.n3177 vdd.n3176 185
R16177 vdd.n3175 vdd.n3174 185
R16178 vdd.n3173 vdd.n3172 185
R16179 vdd.n3171 vdd.n3170 185
R16180 vdd.n3169 vdd.n3168 185
R16181 vdd.n3167 vdd.n3166 185
R16182 vdd.n3165 vdd.n3164 185
R16183 vdd.n3163 vdd.n3162 185
R16184 vdd.n3161 vdd.n3160 185
R16185 vdd.n3159 vdd.n3158 185
R16186 vdd.n3157 vdd.n3156 185
R16187 vdd.n3155 vdd.n3154 185
R16188 vdd.n3153 vdd.n3152 185
R16189 vdd.n3151 vdd.n3150 185
R16190 vdd.n3149 vdd.n3148 185
R16191 vdd.n3147 vdd.n3146 185
R16192 vdd.n3145 vdd.n3144 185
R16193 vdd.n3143 vdd.n3142 185
R16194 vdd.n3141 vdd.n3140 185
R16195 vdd.n3139 vdd.n3138 185
R16196 vdd.n3132 vdd.n767 185
R16197 vdd.n3134 vdd.n3133 185
R16198 vdd.n3131 vdd.n3130 185
R16199 vdd.n3129 vdd.n3128 185
R16200 vdd.n3127 vdd.n3126 185
R16201 vdd.n3125 vdd.n3124 185
R16202 vdd.n3123 vdd.n3122 185
R16203 vdd.n3121 vdd.n3120 185
R16204 vdd.n3119 vdd.n3118 185
R16205 vdd.n3117 vdd.n3116 185
R16206 vdd.n3115 vdd.n3114 185
R16207 vdd.n3113 vdd.n3112 185
R16208 vdd.n3111 vdd.n3110 185
R16209 vdd.n3109 vdd.n3108 185
R16210 vdd.n3107 vdd.n3106 185
R16211 vdd.n3105 vdd.n3104 185
R16212 vdd.n3103 vdd.n3102 185
R16213 vdd.n3101 vdd.n3100 185
R16214 vdd.n3099 vdd.n3098 185
R16215 vdd.n3097 vdd.n3096 185
R16216 vdd.n3095 vdd.n691 185
R16217 vdd.n3225 vdd.n3224 185
R16218 vdd.n3224 vdd.n3223 185
R16219 vdd.n3352 vdd.n3351 185
R16220 vdd.n618 vdd.n425 185
R16221 vdd.n617 vdd.n616 185
R16222 vdd.n615 vdd.n614 185
R16223 vdd.n613 vdd.n430 185
R16224 vdd.n609 vdd.n608 185
R16225 vdd.n607 vdd.n606 185
R16226 vdd.n605 vdd.n604 185
R16227 vdd.n603 vdd.n432 185
R16228 vdd.n599 vdd.n598 185
R16229 vdd.n597 vdd.n596 185
R16230 vdd.n595 vdd.n594 185
R16231 vdd.n593 vdd.n434 185
R16232 vdd.n589 vdd.n588 185
R16233 vdd.n587 vdd.n586 185
R16234 vdd.n585 vdd.n584 185
R16235 vdd.n583 vdd.n436 185
R16236 vdd.n579 vdd.n578 185
R16237 vdd.n577 vdd.n576 185
R16238 vdd.n575 vdd.n574 185
R16239 vdd.n573 vdd.n438 185
R16240 vdd.n569 vdd.n568 185
R16241 vdd.n567 vdd.n566 185
R16242 vdd.n565 vdd.n564 185
R16243 vdd.n563 vdd.n442 185
R16244 vdd.n559 vdd.n558 185
R16245 vdd.n557 vdd.n556 185
R16246 vdd.n555 vdd.n554 185
R16247 vdd.n553 vdd.n444 185
R16248 vdd.n549 vdd.n548 185
R16249 vdd.n547 vdd.n546 185
R16250 vdd.n545 vdd.n544 185
R16251 vdd.n543 vdd.n446 185
R16252 vdd.n539 vdd.n538 185
R16253 vdd.n537 vdd.n536 185
R16254 vdd.n535 vdd.n534 185
R16255 vdd.n533 vdd.n448 185
R16256 vdd.n529 vdd.n528 185
R16257 vdd.n527 vdd.n526 185
R16258 vdd.n525 vdd.n524 185
R16259 vdd.n523 vdd.n450 185
R16260 vdd.n519 vdd.n518 185
R16261 vdd.n517 vdd.n516 185
R16262 vdd.n515 vdd.n514 185
R16263 vdd.n513 vdd.n454 185
R16264 vdd.n509 vdd.n508 185
R16265 vdd.n507 vdd.n506 185
R16266 vdd.n505 vdd.n504 185
R16267 vdd.n503 vdd.n456 185
R16268 vdd.n499 vdd.n498 185
R16269 vdd.n497 vdd.n496 185
R16270 vdd.n495 vdd.n494 185
R16271 vdd.n493 vdd.n458 185
R16272 vdd.n489 vdd.n488 185
R16273 vdd.n487 vdd.n486 185
R16274 vdd.n485 vdd.n484 185
R16275 vdd.n483 vdd.n460 185
R16276 vdd.n479 vdd.n478 185
R16277 vdd.n477 vdd.n476 185
R16278 vdd.n475 vdd.n474 185
R16279 vdd.n473 vdd.n462 185
R16280 vdd.n469 vdd.n468 185
R16281 vdd.n467 vdd.n466 185
R16282 vdd.n465 vdd.n392 185
R16283 vdd.n3348 vdd.n393 185
R16284 vdd.n3355 vdd.n393 185
R16285 vdd.n3347 vdd.n3346 185
R16286 vdd.n3346 vdd.n386 185
R16287 vdd.n3345 vdd.n385 185
R16288 vdd.n3361 vdd.n385 185
R16289 vdd.n621 vdd.n384 185
R16290 vdd.n3362 vdd.n384 185
R16291 vdd.n3341 vdd.n383 185
R16292 vdd.n3363 vdd.n383 185
R16293 vdd.n3340 vdd.n3339 185
R16294 vdd.n3339 vdd.n375 185
R16295 vdd.n3338 vdd.n374 185
R16296 vdd.n3369 vdd.n374 185
R16297 vdd.n623 vdd.n373 185
R16298 vdd.n3370 vdd.n373 185
R16299 vdd.n3334 vdd.n372 185
R16300 vdd.n3371 vdd.n372 185
R16301 vdd.n3333 vdd.n3332 185
R16302 vdd.n3332 vdd.n3331 185
R16303 vdd.n3330 vdd.n364 185
R16304 vdd.n3377 vdd.n364 185
R16305 vdd.n625 vdd.n363 185
R16306 vdd.n3378 vdd.n363 185
R16307 vdd.n3326 vdd.n362 185
R16308 vdd.n3379 vdd.n362 185
R16309 vdd.n3325 vdd.n3324 185
R16310 vdd.n3324 vdd.n361 185
R16311 vdd.n3323 vdd.n353 185
R16312 vdd.n3385 vdd.n353 185
R16313 vdd.n627 vdd.n352 185
R16314 vdd.n3386 vdd.n352 185
R16315 vdd.n3319 vdd.n351 185
R16316 vdd.n3387 vdd.n351 185
R16317 vdd.n3318 vdd.n3317 185
R16318 vdd.n3317 vdd.n344 185
R16319 vdd.n3316 vdd.n343 185
R16320 vdd.n3393 vdd.n343 185
R16321 vdd.n629 vdd.n342 185
R16322 vdd.n3394 vdd.n342 185
R16323 vdd.n3312 vdd.n341 185
R16324 vdd.n3395 vdd.n341 185
R16325 vdd.n3311 vdd.n3310 185
R16326 vdd.n3310 vdd.n340 185
R16327 vdd.n3309 vdd.n631 185
R16328 vdd.n3309 vdd.n3308 185
R16329 vdd.n3297 vdd.n632 185
R16330 vdd.n633 vdd.n632 185
R16331 vdd.n3299 vdd.n3298 185
R16332 vdd.n3300 vdd.n3299 185
R16333 vdd.n640 vdd.n639 185
R16334 vdd.n644 vdd.n639 185
R16335 vdd.n3291 vdd.n3290 185
R16336 vdd.n3290 vdd.n3289 185
R16337 vdd.n643 vdd.n642 185
R16338 vdd.n3280 vdd.n643 185
R16339 vdd.n3279 vdd.n3278 185
R16340 vdd.n3281 vdd.n3279 185
R16341 vdd.n651 vdd.n650 185
R16342 vdd.n656 vdd.n650 185
R16343 vdd.n3274 vdd.n3273 185
R16344 vdd.n3273 vdd.n3272 185
R16345 vdd.n654 vdd.n653 185
R16346 vdd.n655 vdd.n654 185
R16347 vdd.n3263 vdd.n3262 185
R16348 vdd.n3264 vdd.n3263 185
R16349 vdd.n664 vdd.n663 185
R16350 vdd.n663 vdd.n662 185
R16351 vdd.n3258 vdd.n3257 185
R16352 vdd.n3257 vdd.n3256 185
R16353 vdd.n667 vdd.n666 185
R16354 vdd.n3247 vdd.n667 185
R16355 vdd.n3246 vdd.n3245 185
R16356 vdd.n3248 vdd.n3246 185
R16357 vdd.n674 vdd.n673 185
R16358 vdd.n679 vdd.n673 185
R16359 vdd.n3241 vdd.n3240 185
R16360 vdd.n3240 vdd.n3239 185
R16361 vdd.n677 vdd.n676 185
R16362 vdd.n678 vdd.n677 185
R16363 vdd.n3230 vdd.n3229 185
R16364 vdd.n3231 vdd.n3230 185
R16365 vdd.n686 vdd.n685 185
R16366 vdd.n723 vdd.n685 185
R16367 vdd.n913 vdd.n912 185
R16368 vdd.n2855 vdd.n2854 185
R16369 vdd.n2853 vdd.n2638 185
R16370 vdd.n2857 vdd.n2638 185
R16371 vdd.n2852 vdd.n2851 185
R16372 vdd.n2850 vdd.n2849 185
R16373 vdd.n2848 vdd.n2847 185
R16374 vdd.n2846 vdd.n2845 185
R16375 vdd.n2844 vdd.n2843 185
R16376 vdd.n2842 vdd.n2841 185
R16377 vdd.n2840 vdd.n2839 185
R16378 vdd.n2838 vdd.n2837 185
R16379 vdd.n2836 vdd.n2835 185
R16380 vdd.n2834 vdd.n2833 185
R16381 vdd.n2832 vdd.n2831 185
R16382 vdd.n2830 vdd.n2829 185
R16383 vdd.n2828 vdd.n2827 185
R16384 vdd.n2826 vdd.n2825 185
R16385 vdd.n2824 vdd.n2823 185
R16386 vdd.n2822 vdd.n2821 185
R16387 vdd.n2820 vdd.n2819 185
R16388 vdd.n2818 vdd.n2817 185
R16389 vdd.n2816 vdd.n2815 185
R16390 vdd.n2814 vdd.n2813 185
R16391 vdd.n2812 vdd.n2811 185
R16392 vdd.n2810 vdd.n2809 185
R16393 vdd.n2808 vdd.n2807 185
R16394 vdd.n2806 vdd.n2805 185
R16395 vdd.n2804 vdd.n2803 185
R16396 vdd.n2802 vdd.n2801 185
R16397 vdd.n2800 vdd.n2799 185
R16398 vdd.n2798 vdd.n2797 185
R16399 vdd.n2796 vdd.n2795 185
R16400 vdd.n2793 vdd.n2792 185
R16401 vdd.n2791 vdd.n2790 185
R16402 vdd.n2789 vdd.n2788 185
R16403 vdd.n2995 vdd.n2994 185
R16404 vdd.n2997 vdd.n834 185
R16405 vdd.n2999 vdd.n2998 185
R16406 vdd.n3001 vdd.n831 185
R16407 vdd.n3003 vdd.n3002 185
R16408 vdd.n3005 vdd.n829 185
R16409 vdd.n3007 vdd.n3006 185
R16410 vdd.n3008 vdd.n828 185
R16411 vdd.n3010 vdd.n3009 185
R16412 vdd.n3012 vdd.n826 185
R16413 vdd.n3014 vdd.n3013 185
R16414 vdd.n3015 vdd.n825 185
R16415 vdd.n3017 vdd.n3016 185
R16416 vdd.n3019 vdd.n823 185
R16417 vdd.n3021 vdd.n3020 185
R16418 vdd.n3022 vdd.n822 185
R16419 vdd.n3024 vdd.n3023 185
R16420 vdd.n3026 vdd.n731 185
R16421 vdd.n3028 vdd.n3027 185
R16422 vdd.n3030 vdd.n820 185
R16423 vdd.n3032 vdd.n3031 185
R16424 vdd.n3033 vdd.n819 185
R16425 vdd.n3035 vdd.n3034 185
R16426 vdd.n3037 vdd.n817 185
R16427 vdd.n3039 vdd.n3038 185
R16428 vdd.n3040 vdd.n816 185
R16429 vdd.n3042 vdd.n3041 185
R16430 vdd.n3044 vdd.n814 185
R16431 vdd.n3046 vdd.n3045 185
R16432 vdd.n3047 vdd.n813 185
R16433 vdd.n3049 vdd.n3048 185
R16434 vdd.n3051 vdd.n812 185
R16435 vdd.n3052 vdd.n811 185
R16436 vdd.n3055 vdd.n3054 185
R16437 vdd.n3056 vdd.n809 185
R16438 vdd.n809 vdd.n692 185
R16439 vdd.n2993 vdd.n806 185
R16440 vdd.n3059 vdd.n806 185
R16441 vdd.n2992 vdd.n2991 185
R16442 vdd.n2991 vdd.n805 185
R16443 vdd.n2990 vdd.n836 185
R16444 vdd.n2990 vdd.n2989 185
R16445 vdd.n2744 vdd.n837 185
R16446 vdd.n846 vdd.n837 185
R16447 vdd.n2745 vdd.n844 185
R16448 vdd.n2983 vdd.n844 185
R16449 vdd.n2747 vdd.n2746 185
R16450 vdd.n2746 vdd.n843 185
R16451 vdd.n2748 vdd.n852 185
R16452 vdd.n2932 vdd.n852 185
R16453 vdd.n2750 vdd.n2749 185
R16454 vdd.n2749 vdd.n851 185
R16455 vdd.n2751 vdd.n858 185
R16456 vdd.n2926 vdd.n858 185
R16457 vdd.n2753 vdd.n2752 185
R16458 vdd.n2752 vdd.n857 185
R16459 vdd.n2754 vdd.n863 185
R16460 vdd.n2918 vdd.n863 185
R16461 vdd.n2756 vdd.n2755 185
R16462 vdd.n2755 vdd.n870 185
R16463 vdd.n2757 vdd.n868 185
R16464 vdd.n2912 vdd.n868 185
R16465 vdd.n2759 vdd.n2758 185
R16466 vdd.n2760 vdd.n2759 185
R16467 vdd.n2743 vdd.n875 185
R16468 vdd.n2906 vdd.n875 185
R16469 vdd.n2742 vdd.n2741 185
R16470 vdd.n2741 vdd.n874 185
R16471 vdd.n2740 vdd.n881 185
R16472 vdd.n2900 vdd.n881 185
R16473 vdd.n2739 vdd.n2738 185
R16474 vdd.n2738 vdd.n880 185
R16475 vdd.n2737 vdd.n886 185
R16476 vdd.n2894 vdd.n886 185
R16477 vdd.n2736 vdd.n2735 185
R16478 vdd.n2735 vdd.n893 185
R16479 vdd.n2734 vdd.n891 185
R16480 vdd.n2888 vdd.n891 185
R16481 vdd.n2733 vdd.n2732 185
R16482 vdd.n2732 vdd.n900 185
R16483 vdd.n2731 vdd.n898 185
R16484 vdd.n2882 vdd.n898 185
R16485 vdd.n2730 vdd.n2729 185
R16486 vdd.n2729 vdd.n897 185
R16487 vdd.n2641 vdd.n904 185
R16488 vdd.n2876 vdd.n904 185
R16489 vdd.n2783 vdd.n2782 185
R16490 vdd.n2782 vdd.n2781 185
R16491 vdd.n2784 vdd.n909 185
R16492 vdd.n2870 vdd.n909 185
R16493 vdd.n2786 vdd.n2785 185
R16494 vdd.n2785 vdd.t288 185
R16495 vdd.n2787 vdd.n914 185
R16496 vdd.n2864 vdd.n914 185
R16497 vdd.n2866 vdd.n2865 185
R16498 vdd.n2865 vdd.n2864 185
R16499 vdd.n2867 vdd.n911 185
R16500 vdd.n911 vdd.t288 185
R16501 vdd.n2869 vdd.n2868 185
R16502 vdd.n2870 vdd.n2869 185
R16503 vdd.n903 vdd.n902 185
R16504 vdd.n2781 vdd.n903 185
R16505 vdd.n2878 vdd.n2877 185
R16506 vdd.n2877 vdd.n2876 185
R16507 vdd.n2879 vdd.n901 185
R16508 vdd.n901 vdd.n897 185
R16509 vdd.n2881 vdd.n2880 185
R16510 vdd.n2882 vdd.n2881 185
R16511 vdd.n890 vdd.n889 185
R16512 vdd.n900 vdd.n890 185
R16513 vdd.n2890 vdd.n2889 185
R16514 vdd.n2889 vdd.n2888 185
R16515 vdd.n2891 vdd.n888 185
R16516 vdd.n893 vdd.n888 185
R16517 vdd.n2893 vdd.n2892 185
R16518 vdd.n2894 vdd.n2893 185
R16519 vdd.n879 vdd.n878 185
R16520 vdd.n880 vdd.n879 185
R16521 vdd.n2902 vdd.n2901 185
R16522 vdd.n2901 vdd.n2900 185
R16523 vdd.n2903 vdd.n877 185
R16524 vdd.n877 vdd.n874 185
R16525 vdd.n2905 vdd.n2904 185
R16526 vdd.n2906 vdd.n2905 185
R16527 vdd.n867 vdd.n866 185
R16528 vdd.n2760 vdd.n867 185
R16529 vdd.n2914 vdd.n2913 185
R16530 vdd.n2913 vdd.n2912 185
R16531 vdd.n2915 vdd.n865 185
R16532 vdd.n870 vdd.n865 185
R16533 vdd.n2917 vdd.n2916 185
R16534 vdd.n2918 vdd.n2917 185
R16535 vdd.n856 vdd.n855 185
R16536 vdd.n857 vdd.n856 185
R16537 vdd.n2928 vdd.n2927 185
R16538 vdd.n2927 vdd.n2926 185
R16539 vdd.n2929 vdd.n854 185
R16540 vdd.n854 vdd.n851 185
R16541 vdd.n2931 vdd.n2930 185
R16542 vdd.n2932 vdd.n2931 185
R16543 vdd.n842 vdd.n841 185
R16544 vdd.n843 vdd.n842 185
R16545 vdd.n2985 vdd.n2984 185
R16546 vdd.n2984 vdd.n2983 185
R16547 vdd.n2986 vdd.n840 185
R16548 vdd.n846 vdd.n840 185
R16549 vdd.n2988 vdd.n2987 185
R16550 vdd.n2989 vdd.n2988 185
R16551 vdd.n810 vdd.n808 185
R16552 vdd.n808 vdd.n805 185
R16553 vdd.n3058 vdd.n3057 185
R16554 vdd.n3059 vdd.n3058 185
R16555 vdd.n2531 vdd.n2530 185
R16556 vdd.n2532 vdd.n2531 185
R16557 vdd.n964 vdd.n962 185
R16558 vdd.n962 vdd.t5 185
R16559 vdd.n2446 vdd.n971 185
R16560 vdd.n2457 vdd.n971 185
R16561 vdd.n2447 vdd.n980 185
R16562 vdd.n2156 vdd.n980 185
R16563 vdd.n2449 vdd.n2448 185
R16564 vdd.n2450 vdd.n2449 185
R16565 vdd.n2445 vdd.n979 185
R16566 vdd.n979 vdd.n976 185
R16567 vdd.n2444 vdd.n2443 185
R16568 vdd.n2443 vdd.n2442 185
R16569 vdd.n982 vdd.n981 185
R16570 vdd.n983 vdd.n982 185
R16571 vdd.n2435 vdd.n2434 185
R16572 vdd.n2436 vdd.n2435 185
R16573 vdd.n2433 vdd.n992 185
R16574 vdd.n992 vdd.n989 185
R16575 vdd.n2432 vdd.n2431 185
R16576 vdd.n2431 vdd.n2430 185
R16577 vdd.n994 vdd.n993 185
R16578 vdd.n1002 vdd.n994 185
R16579 vdd.n2423 vdd.n2422 185
R16580 vdd.n2424 vdd.n2423 185
R16581 vdd.n2421 vdd.n1003 185
R16582 vdd.n1008 vdd.n1003 185
R16583 vdd.n2420 vdd.n2419 185
R16584 vdd.n2419 vdd.n2418 185
R16585 vdd.n1005 vdd.n1004 185
R16586 vdd.n2257 vdd.n1005 185
R16587 vdd.n2411 vdd.n2410 185
R16588 vdd.n2412 vdd.n2411 185
R16589 vdd.n2409 vdd.n1015 185
R16590 vdd.n1015 vdd.n1012 185
R16591 vdd.n2408 vdd.n2407 185
R16592 vdd.n2407 vdd.n2406 185
R16593 vdd.n1017 vdd.n1016 185
R16594 vdd.n1018 vdd.n1017 185
R16595 vdd.n2399 vdd.n2398 185
R16596 vdd.n2400 vdd.n2399 185
R16597 vdd.n2396 vdd.n1026 185
R16598 vdd.n1033 vdd.n1026 185
R16599 vdd.n2395 vdd.n2394 185
R16600 vdd.n2394 vdd.n2393 185
R16601 vdd.n1029 vdd.n1028 185
R16602 vdd.n1030 vdd.n1029 185
R16603 vdd.n2386 vdd.n2385 185
R16604 vdd.n2387 vdd.n2386 185
R16605 vdd.n2384 vdd.n1040 185
R16606 vdd.n1040 vdd.n1037 185
R16607 vdd.n2383 vdd.n2382 185
R16608 vdd.n2382 vdd.n2381 185
R16609 vdd.n1042 vdd.n1041 185
R16610 vdd.n1043 vdd.n1042 185
R16611 vdd.n2374 vdd.n2373 185
R16612 vdd.n2375 vdd.n2374 185
R16613 vdd.n2462 vdd.n936 185
R16614 vdd.n2604 vdd.n936 185
R16615 vdd.n2464 vdd.n2463 185
R16616 vdd.n2466 vdd.n2465 185
R16617 vdd.n2468 vdd.n2467 185
R16618 vdd.n2470 vdd.n2469 185
R16619 vdd.n2472 vdd.n2471 185
R16620 vdd.n2474 vdd.n2473 185
R16621 vdd.n2476 vdd.n2475 185
R16622 vdd.n2478 vdd.n2477 185
R16623 vdd.n2480 vdd.n2479 185
R16624 vdd.n2482 vdd.n2481 185
R16625 vdd.n2484 vdd.n2483 185
R16626 vdd.n2486 vdd.n2485 185
R16627 vdd.n2488 vdd.n2487 185
R16628 vdd.n2490 vdd.n2489 185
R16629 vdd.n2492 vdd.n2491 185
R16630 vdd.n2494 vdd.n2493 185
R16631 vdd.n2496 vdd.n2495 185
R16632 vdd.n2498 vdd.n2497 185
R16633 vdd.n2500 vdd.n2499 185
R16634 vdd.n2502 vdd.n2501 185
R16635 vdd.n2504 vdd.n2503 185
R16636 vdd.n2506 vdd.n2505 185
R16637 vdd.n2508 vdd.n2507 185
R16638 vdd.n2510 vdd.n2509 185
R16639 vdd.n2512 vdd.n2511 185
R16640 vdd.n2514 vdd.n2513 185
R16641 vdd.n2516 vdd.n2515 185
R16642 vdd.n2518 vdd.n2517 185
R16643 vdd.n2520 vdd.n2519 185
R16644 vdd.n2522 vdd.n2521 185
R16645 vdd.n2524 vdd.n2523 185
R16646 vdd.n2526 vdd.n2525 185
R16647 vdd.n2528 vdd.n2527 185
R16648 vdd.n2529 vdd.n963 185
R16649 vdd.n2461 vdd.n961 185
R16650 vdd.n2532 vdd.n961 185
R16651 vdd.n2460 vdd.n2459 185
R16652 vdd.n2459 vdd.t5 185
R16653 vdd.n2458 vdd.n968 185
R16654 vdd.n2458 vdd.n2457 185
R16655 vdd.n2238 vdd.n969 185
R16656 vdd.n2156 vdd.n969 185
R16657 vdd.n2239 vdd.n978 185
R16658 vdd.n2450 vdd.n978 185
R16659 vdd.n2241 vdd.n2240 185
R16660 vdd.n2240 vdd.n976 185
R16661 vdd.n2242 vdd.n985 185
R16662 vdd.n2442 vdd.n985 185
R16663 vdd.n2244 vdd.n2243 185
R16664 vdd.n2243 vdd.n983 185
R16665 vdd.n2245 vdd.n991 185
R16666 vdd.n2436 vdd.n991 185
R16667 vdd.n2247 vdd.n2246 185
R16668 vdd.n2246 vdd.n989 185
R16669 vdd.n2248 vdd.n996 185
R16670 vdd.n2430 vdd.n996 185
R16671 vdd.n2250 vdd.n2249 185
R16672 vdd.n2249 vdd.n1002 185
R16673 vdd.n2251 vdd.n1001 185
R16674 vdd.n2424 vdd.n1001 185
R16675 vdd.n2253 vdd.n2252 185
R16676 vdd.n2252 vdd.n1008 185
R16677 vdd.n2254 vdd.n1007 185
R16678 vdd.n2418 vdd.n1007 185
R16679 vdd.n2256 vdd.n2255 185
R16680 vdd.n2257 vdd.n2256 185
R16681 vdd.n2237 vdd.n1014 185
R16682 vdd.n2412 vdd.n1014 185
R16683 vdd.n2236 vdd.n2235 185
R16684 vdd.n2235 vdd.n1012 185
R16685 vdd.n2234 vdd.n1020 185
R16686 vdd.n2406 vdd.n1020 185
R16687 vdd.n2233 vdd.n2232 185
R16688 vdd.n2232 vdd.n1018 185
R16689 vdd.n2231 vdd.n1025 185
R16690 vdd.n2400 vdd.n1025 185
R16691 vdd.n2230 vdd.n2229 185
R16692 vdd.n2229 vdd.n1033 185
R16693 vdd.n2228 vdd.n1032 185
R16694 vdd.n2393 vdd.n1032 185
R16695 vdd.n2227 vdd.n2226 185
R16696 vdd.n2226 vdd.n1030 185
R16697 vdd.n2225 vdd.n1039 185
R16698 vdd.n2387 vdd.n1039 185
R16699 vdd.n2224 vdd.n2223 185
R16700 vdd.n2223 vdd.n1037 185
R16701 vdd.n2222 vdd.n1045 185
R16702 vdd.n2381 vdd.n1045 185
R16703 vdd.n2221 vdd.n2220 185
R16704 vdd.n2220 vdd.n1043 185
R16705 vdd.n2219 vdd.n1051 185
R16706 vdd.n2375 vdd.n1051 185
R16707 vdd.n2372 vdd.n1052 185
R16708 vdd.n2371 vdd.n2370 185
R16709 vdd.n2368 vdd.n1053 185
R16710 vdd.n2366 vdd.n2365 185
R16711 vdd.n2364 vdd.n1054 185
R16712 vdd.n2363 vdd.n2362 185
R16713 vdd.n2360 vdd.n1055 185
R16714 vdd.n2358 vdd.n2357 185
R16715 vdd.n2356 vdd.n1056 185
R16716 vdd.n2355 vdd.n2354 185
R16717 vdd.n2352 vdd.n1057 185
R16718 vdd.n2350 vdd.n2349 185
R16719 vdd.n2348 vdd.n1058 185
R16720 vdd.n2347 vdd.n2346 185
R16721 vdd.n2344 vdd.n1059 185
R16722 vdd.n2342 vdd.n2341 185
R16723 vdd.n2340 vdd.n1060 185
R16724 vdd.n2339 vdd.n1062 185
R16725 vdd.n2184 vdd.n1063 185
R16726 vdd.n2187 vdd.n2186 185
R16727 vdd.n2189 vdd.n2188 185
R16728 vdd.n2191 vdd.n2183 185
R16729 vdd.n2194 vdd.n2193 185
R16730 vdd.n2195 vdd.n2182 185
R16731 vdd.n2197 vdd.n2196 185
R16732 vdd.n2199 vdd.n2181 185
R16733 vdd.n2202 vdd.n2201 185
R16734 vdd.n2203 vdd.n2180 185
R16735 vdd.n2205 vdd.n2204 185
R16736 vdd.n2207 vdd.n2179 185
R16737 vdd.n2210 vdd.n2209 185
R16738 vdd.n2211 vdd.n2176 185
R16739 vdd.n2214 vdd.n2213 185
R16740 vdd.n2216 vdd.n2175 185
R16741 vdd.n2218 vdd.n2217 185
R16742 vdd.n2217 vdd.n1049 185
R16743 vdd.n327 vdd.n326 171.744
R16744 vdd.n326 vdd.n325 171.744
R16745 vdd.n325 vdd.n294 171.744
R16746 vdd.n318 vdd.n294 171.744
R16747 vdd.n318 vdd.n317 171.744
R16748 vdd.n317 vdd.n299 171.744
R16749 vdd.n310 vdd.n299 171.744
R16750 vdd.n310 vdd.n309 171.744
R16751 vdd.n309 vdd.n303 171.744
R16752 vdd.n268 vdd.n267 171.744
R16753 vdd.n267 vdd.n266 171.744
R16754 vdd.n266 vdd.n235 171.744
R16755 vdd.n259 vdd.n235 171.744
R16756 vdd.n259 vdd.n258 171.744
R16757 vdd.n258 vdd.n240 171.744
R16758 vdd.n251 vdd.n240 171.744
R16759 vdd.n251 vdd.n250 171.744
R16760 vdd.n250 vdd.n244 171.744
R16761 vdd.n225 vdd.n224 171.744
R16762 vdd.n224 vdd.n223 171.744
R16763 vdd.n223 vdd.n192 171.744
R16764 vdd.n216 vdd.n192 171.744
R16765 vdd.n216 vdd.n215 171.744
R16766 vdd.n215 vdd.n197 171.744
R16767 vdd.n208 vdd.n197 171.744
R16768 vdd.n208 vdd.n207 171.744
R16769 vdd.n207 vdd.n201 171.744
R16770 vdd.n166 vdd.n165 171.744
R16771 vdd.n165 vdd.n164 171.744
R16772 vdd.n164 vdd.n133 171.744
R16773 vdd.n157 vdd.n133 171.744
R16774 vdd.n157 vdd.n156 171.744
R16775 vdd.n156 vdd.n138 171.744
R16776 vdd.n149 vdd.n138 171.744
R16777 vdd.n149 vdd.n148 171.744
R16778 vdd.n148 vdd.n142 171.744
R16779 vdd.n124 vdd.n123 171.744
R16780 vdd.n123 vdd.n122 171.744
R16781 vdd.n122 vdd.n91 171.744
R16782 vdd.n115 vdd.n91 171.744
R16783 vdd.n115 vdd.n114 171.744
R16784 vdd.n114 vdd.n96 171.744
R16785 vdd.n107 vdd.n96 171.744
R16786 vdd.n107 vdd.n106 171.744
R16787 vdd.n106 vdd.n100 171.744
R16788 vdd.n65 vdd.n64 171.744
R16789 vdd.n64 vdd.n63 171.744
R16790 vdd.n63 vdd.n32 171.744
R16791 vdd.n56 vdd.n32 171.744
R16792 vdd.n56 vdd.n55 171.744
R16793 vdd.n55 vdd.n37 171.744
R16794 vdd.n48 vdd.n37 171.744
R16795 vdd.n48 vdd.n47 171.744
R16796 vdd.n47 vdd.n41 171.744
R16797 vdd.n1746 vdd.n1745 171.744
R16798 vdd.n1745 vdd.n1744 171.744
R16799 vdd.n1744 vdd.n1713 171.744
R16800 vdd.n1737 vdd.n1713 171.744
R16801 vdd.n1737 vdd.n1736 171.744
R16802 vdd.n1736 vdd.n1718 171.744
R16803 vdd.n1729 vdd.n1718 171.744
R16804 vdd.n1729 vdd.n1728 171.744
R16805 vdd.n1728 vdd.n1722 171.744
R16806 vdd.n1805 vdd.n1804 171.744
R16807 vdd.n1804 vdd.n1803 171.744
R16808 vdd.n1803 vdd.n1772 171.744
R16809 vdd.n1796 vdd.n1772 171.744
R16810 vdd.n1796 vdd.n1795 171.744
R16811 vdd.n1795 vdd.n1777 171.744
R16812 vdd.n1788 vdd.n1777 171.744
R16813 vdd.n1788 vdd.n1787 171.744
R16814 vdd.n1787 vdd.n1781 171.744
R16815 vdd.n1644 vdd.n1643 171.744
R16816 vdd.n1643 vdd.n1642 171.744
R16817 vdd.n1642 vdd.n1611 171.744
R16818 vdd.n1635 vdd.n1611 171.744
R16819 vdd.n1635 vdd.n1634 171.744
R16820 vdd.n1634 vdd.n1616 171.744
R16821 vdd.n1627 vdd.n1616 171.744
R16822 vdd.n1627 vdd.n1626 171.744
R16823 vdd.n1626 vdd.n1620 171.744
R16824 vdd.n1703 vdd.n1702 171.744
R16825 vdd.n1702 vdd.n1701 171.744
R16826 vdd.n1701 vdd.n1670 171.744
R16827 vdd.n1694 vdd.n1670 171.744
R16828 vdd.n1694 vdd.n1693 171.744
R16829 vdd.n1693 vdd.n1675 171.744
R16830 vdd.n1686 vdd.n1675 171.744
R16831 vdd.n1686 vdd.n1685 171.744
R16832 vdd.n1685 vdd.n1679 171.744
R16833 vdd.n1543 vdd.n1542 171.744
R16834 vdd.n1542 vdd.n1541 171.744
R16835 vdd.n1541 vdd.n1510 171.744
R16836 vdd.n1534 vdd.n1510 171.744
R16837 vdd.n1534 vdd.n1533 171.744
R16838 vdd.n1533 vdd.n1515 171.744
R16839 vdd.n1526 vdd.n1515 171.744
R16840 vdd.n1526 vdd.n1525 171.744
R16841 vdd.n1525 vdd.n1519 171.744
R16842 vdd.n1602 vdd.n1601 171.744
R16843 vdd.n1601 vdd.n1600 171.744
R16844 vdd.n1600 vdd.n1569 171.744
R16845 vdd.n1593 vdd.n1569 171.744
R16846 vdd.n1593 vdd.n1592 171.744
R16847 vdd.n1592 vdd.n1574 171.744
R16848 vdd.n1585 vdd.n1574 171.744
R16849 vdd.n1585 vdd.n1584 171.744
R16850 vdd.n1584 vdd.n1578 171.744
R16851 vdd.n468 vdd.n467 146.341
R16852 vdd.n474 vdd.n473 146.341
R16853 vdd.n478 vdd.n477 146.341
R16854 vdd.n484 vdd.n483 146.341
R16855 vdd.n488 vdd.n487 146.341
R16856 vdd.n494 vdd.n493 146.341
R16857 vdd.n498 vdd.n497 146.341
R16858 vdd.n504 vdd.n503 146.341
R16859 vdd.n508 vdd.n507 146.341
R16860 vdd.n514 vdd.n513 146.341
R16861 vdd.n518 vdd.n517 146.341
R16862 vdd.n524 vdd.n523 146.341
R16863 vdd.n528 vdd.n527 146.341
R16864 vdd.n534 vdd.n533 146.341
R16865 vdd.n538 vdd.n537 146.341
R16866 vdd.n544 vdd.n543 146.341
R16867 vdd.n548 vdd.n547 146.341
R16868 vdd.n554 vdd.n553 146.341
R16869 vdd.n558 vdd.n557 146.341
R16870 vdd.n564 vdd.n563 146.341
R16871 vdd.n568 vdd.n567 146.341
R16872 vdd.n574 vdd.n573 146.341
R16873 vdd.n578 vdd.n577 146.341
R16874 vdd.n584 vdd.n583 146.341
R16875 vdd.n588 vdd.n587 146.341
R16876 vdd.n594 vdd.n593 146.341
R16877 vdd.n598 vdd.n597 146.341
R16878 vdd.n604 vdd.n603 146.341
R16879 vdd.n608 vdd.n607 146.341
R16880 vdd.n614 vdd.n613 146.341
R16881 vdd.n616 vdd.n425 146.341
R16882 vdd.n3230 vdd.n685 146.341
R16883 vdd.n3230 vdd.n677 146.341
R16884 vdd.n3240 vdd.n677 146.341
R16885 vdd.n3240 vdd.n673 146.341
R16886 vdd.n3246 vdd.n673 146.341
R16887 vdd.n3246 vdd.n667 146.341
R16888 vdd.n3257 vdd.n667 146.341
R16889 vdd.n3257 vdd.n663 146.341
R16890 vdd.n3263 vdd.n663 146.341
R16891 vdd.n3263 vdd.n654 146.341
R16892 vdd.n3273 vdd.n654 146.341
R16893 vdd.n3273 vdd.n650 146.341
R16894 vdd.n3279 vdd.n650 146.341
R16895 vdd.n3279 vdd.n643 146.341
R16896 vdd.n3290 vdd.n643 146.341
R16897 vdd.n3290 vdd.n639 146.341
R16898 vdd.n3299 vdd.n639 146.341
R16899 vdd.n3299 vdd.n632 146.341
R16900 vdd.n3309 vdd.n632 146.341
R16901 vdd.n3310 vdd.n3309 146.341
R16902 vdd.n3310 vdd.n341 146.341
R16903 vdd.n342 vdd.n341 146.341
R16904 vdd.n343 vdd.n342 146.341
R16905 vdd.n3317 vdd.n343 146.341
R16906 vdd.n3317 vdd.n351 146.341
R16907 vdd.n352 vdd.n351 146.341
R16908 vdd.n353 vdd.n352 146.341
R16909 vdd.n3324 vdd.n353 146.341
R16910 vdd.n3324 vdd.n362 146.341
R16911 vdd.n363 vdd.n362 146.341
R16912 vdd.n364 vdd.n363 146.341
R16913 vdd.n3332 vdd.n364 146.341
R16914 vdd.n3332 vdd.n372 146.341
R16915 vdd.n373 vdd.n372 146.341
R16916 vdd.n374 vdd.n373 146.341
R16917 vdd.n3339 vdd.n374 146.341
R16918 vdd.n3339 vdd.n383 146.341
R16919 vdd.n384 vdd.n383 146.341
R16920 vdd.n385 vdd.n384 146.341
R16921 vdd.n3346 vdd.n385 146.341
R16922 vdd.n3346 vdd.n393 146.341
R16923 vdd.n725 vdd.n724 146.341
R16924 vdd.n728 vdd.n724 146.341
R16925 vdd.n734 vdd.n733 146.341
R16926 vdd.n3212 vdd.n3211 146.341
R16927 vdd.n3208 vdd.n3207 146.341
R16928 vdd.n3204 vdd.n3203 146.341
R16929 vdd.n3200 vdd.n3199 146.341
R16930 vdd.n3196 vdd.n3195 146.341
R16931 vdd.n3192 vdd.n3191 146.341
R16932 vdd.n3188 vdd.n3187 146.341
R16933 vdd.n3179 vdd.n3178 146.341
R16934 vdd.n3176 vdd.n3175 146.341
R16935 vdd.n3172 vdd.n3171 146.341
R16936 vdd.n3168 vdd.n3167 146.341
R16937 vdd.n3164 vdd.n3163 146.341
R16938 vdd.n3160 vdd.n3159 146.341
R16939 vdd.n3156 vdd.n3155 146.341
R16940 vdd.n3152 vdd.n3151 146.341
R16941 vdd.n3148 vdd.n3147 146.341
R16942 vdd.n3144 vdd.n3143 146.341
R16943 vdd.n3140 vdd.n3139 146.341
R16944 vdd.n3133 vdd.n3132 146.341
R16945 vdd.n3130 vdd.n3129 146.341
R16946 vdd.n3126 vdd.n3125 146.341
R16947 vdd.n3122 vdd.n3121 146.341
R16948 vdd.n3118 vdd.n3117 146.341
R16949 vdd.n3114 vdd.n3113 146.341
R16950 vdd.n3110 vdd.n3109 146.341
R16951 vdd.n3106 vdd.n3105 146.341
R16952 vdd.n3102 vdd.n3101 146.341
R16953 vdd.n3098 vdd.n3097 146.341
R16954 vdd.n3224 vdd.n691 146.341
R16955 vdd.n3232 vdd.n684 146.341
R16956 vdd.n3232 vdd.n680 146.341
R16957 vdd.n3238 vdd.n680 146.341
R16958 vdd.n3238 vdd.n672 146.341
R16959 vdd.n3249 vdd.n672 146.341
R16960 vdd.n3249 vdd.n668 146.341
R16961 vdd.n3255 vdd.n668 146.341
R16962 vdd.n3255 vdd.n661 146.341
R16963 vdd.n3265 vdd.n661 146.341
R16964 vdd.n3265 vdd.n657 146.341
R16965 vdd.n3271 vdd.n657 146.341
R16966 vdd.n3271 vdd.n649 146.341
R16967 vdd.n3282 vdd.n649 146.341
R16968 vdd.n3282 vdd.n645 146.341
R16969 vdd.n3288 vdd.n645 146.341
R16970 vdd.n3288 vdd.n638 146.341
R16971 vdd.n3301 vdd.n638 146.341
R16972 vdd.n3301 vdd.n634 146.341
R16973 vdd.n3307 vdd.n634 146.341
R16974 vdd.n3307 vdd.n338 146.341
R16975 vdd.n3396 vdd.n338 146.341
R16976 vdd.n3396 vdd.n339 146.341
R16977 vdd.n3392 vdd.n339 146.341
R16978 vdd.n3392 vdd.n345 146.341
R16979 vdd.n3388 vdd.n345 146.341
R16980 vdd.n3388 vdd.n350 146.341
R16981 vdd.n3384 vdd.n350 146.341
R16982 vdd.n3384 vdd.n354 146.341
R16983 vdd.n3380 vdd.n354 146.341
R16984 vdd.n3380 vdd.n360 146.341
R16985 vdd.n3376 vdd.n360 146.341
R16986 vdd.n3376 vdd.n365 146.341
R16987 vdd.n3372 vdd.n365 146.341
R16988 vdd.n3372 vdd.n371 146.341
R16989 vdd.n3368 vdd.n371 146.341
R16990 vdd.n3368 vdd.n376 146.341
R16991 vdd.n3364 vdd.n376 146.341
R16992 vdd.n3364 vdd.n382 146.341
R16993 vdd.n3360 vdd.n382 146.341
R16994 vdd.n3360 vdd.n387 146.341
R16995 vdd.n3356 vdd.n387 146.341
R16996 vdd.n2322 vdd.n2321 146.341
R16997 vdd.n2319 vdd.n1903 146.341
R16998 vdd.n2099 vdd.n1909 146.341
R16999 vdd.n2097 vdd.n2096 146.341
R17000 vdd.n2094 vdd.n1911 146.341
R17001 vdd.n2090 vdd.n2089 146.341
R17002 vdd.n2087 vdd.n1918 146.341
R17003 vdd.n2083 vdd.n2082 146.341
R17004 vdd.n2080 vdd.n1925 146.341
R17005 vdd.n1936 vdd.n1933 146.341
R17006 vdd.n2072 vdd.n2071 146.341
R17007 vdd.n2069 vdd.n1938 146.341
R17008 vdd.n2065 vdd.n2064 146.341
R17009 vdd.n2062 vdd.n1944 146.341
R17010 vdd.n2058 vdd.n2057 146.341
R17011 vdd.n2055 vdd.n1951 146.341
R17012 vdd.n2051 vdd.n2050 146.341
R17013 vdd.n2048 vdd.n1958 146.341
R17014 vdd.n2044 vdd.n2043 146.341
R17015 vdd.n2041 vdd.n1965 146.341
R17016 vdd.n1976 vdd.n1973 146.341
R17017 vdd.n2033 vdd.n2032 146.341
R17018 vdd.n2030 vdd.n1978 146.341
R17019 vdd.n2026 vdd.n2025 146.341
R17020 vdd.n2023 vdd.n1984 146.341
R17021 vdd.n2019 vdd.n2018 146.341
R17022 vdd.n2016 vdd.n1991 146.341
R17023 vdd.n2012 vdd.n2011 146.341
R17024 vdd.n2009 vdd.n2006 146.341
R17025 vdd.n2004 vdd.n2001 146.341
R17026 vdd.n1999 vdd.n1069 146.341
R17027 vdd.n1428 vdd.n1188 146.341
R17028 vdd.n1428 vdd.n1184 146.341
R17029 vdd.n1434 vdd.n1184 146.341
R17030 vdd.n1434 vdd.n1176 146.341
R17031 vdd.n1445 vdd.n1176 146.341
R17032 vdd.n1445 vdd.n1172 146.341
R17033 vdd.n1451 vdd.n1172 146.341
R17034 vdd.n1451 vdd.n1166 146.341
R17035 vdd.n1462 vdd.n1166 146.341
R17036 vdd.n1462 vdd.n1162 146.341
R17037 vdd.n1468 vdd.n1162 146.341
R17038 vdd.n1468 vdd.n1153 146.341
R17039 vdd.n1478 vdd.n1153 146.341
R17040 vdd.n1478 vdd.n1149 146.341
R17041 vdd.n1484 vdd.n1149 146.341
R17042 vdd.n1484 vdd.n1142 146.341
R17043 vdd.n1495 vdd.n1142 146.341
R17044 vdd.n1495 vdd.n1138 146.341
R17045 vdd.n1501 vdd.n1138 146.341
R17046 vdd.n1501 vdd.n1131 146.341
R17047 vdd.n1818 vdd.n1131 146.341
R17048 vdd.n1818 vdd.n1127 146.341
R17049 vdd.n1824 vdd.n1127 146.341
R17050 vdd.n1824 vdd.n1119 146.341
R17051 vdd.n1835 vdd.n1119 146.341
R17052 vdd.n1835 vdd.n1115 146.341
R17053 vdd.n1841 vdd.n1115 146.341
R17054 vdd.n1841 vdd.n1109 146.341
R17055 vdd.n1852 vdd.n1109 146.341
R17056 vdd.n1852 vdd.n1105 146.341
R17057 vdd.n1858 vdd.n1105 146.341
R17058 vdd.n1858 vdd.n1096 146.341
R17059 vdd.n1868 vdd.n1096 146.341
R17060 vdd.n1868 vdd.n1092 146.341
R17061 vdd.n1874 vdd.n1092 146.341
R17062 vdd.n1874 vdd.n1086 146.341
R17063 vdd.n1885 vdd.n1086 146.341
R17064 vdd.n1885 vdd.n1081 146.341
R17065 vdd.n1893 vdd.n1081 146.341
R17066 vdd.n1893 vdd.n1071 146.341
R17067 vdd.n2330 vdd.n1071 146.341
R17068 vdd.n1417 vdd.n1193 146.341
R17069 vdd.n1417 vdd.n1226 146.341
R17070 vdd.n1230 vdd.n1229 146.341
R17071 vdd.n1232 vdd.n1231 146.341
R17072 vdd.n1236 vdd.n1235 146.341
R17073 vdd.n1238 vdd.n1237 146.341
R17074 vdd.n1242 vdd.n1241 146.341
R17075 vdd.n1244 vdd.n1243 146.341
R17076 vdd.n1248 vdd.n1247 146.341
R17077 vdd.n1250 vdd.n1249 146.341
R17078 vdd.n1256 vdd.n1255 146.341
R17079 vdd.n1258 vdd.n1257 146.341
R17080 vdd.n1262 vdd.n1261 146.341
R17081 vdd.n1264 vdd.n1263 146.341
R17082 vdd.n1268 vdd.n1267 146.341
R17083 vdd.n1270 vdd.n1269 146.341
R17084 vdd.n1274 vdd.n1273 146.341
R17085 vdd.n1276 vdd.n1275 146.341
R17086 vdd.n1280 vdd.n1279 146.341
R17087 vdd.n1282 vdd.n1281 146.341
R17088 vdd.n1354 vdd.n1285 146.341
R17089 vdd.n1287 vdd.n1286 146.341
R17090 vdd.n1291 vdd.n1290 146.341
R17091 vdd.n1293 vdd.n1292 146.341
R17092 vdd.n1297 vdd.n1296 146.341
R17093 vdd.n1299 vdd.n1298 146.341
R17094 vdd.n1303 vdd.n1302 146.341
R17095 vdd.n1305 vdd.n1304 146.341
R17096 vdd.n1309 vdd.n1308 146.341
R17097 vdd.n1311 vdd.n1310 146.341
R17098 vdd.n1315 vdd.n1314 146.341
R17099 vdd.n1316 vdd.n1224 146.341
R17100 vdd.n1426 vdd.n1189 146.341
R17101 vdd.n1426 vdd.n1182 146.341
R17102 vdd.n1437 vdd.n1182 146.341
R17103 vdd.n1437 vdd.n1178 146.341
R17104 vdd.n1443 vdd.n1178 146.341
R17105 vdd.n1443 vdd.n1171 146.341
R17106 vdd.n1454 vdd.n1171 146.341
R17107 vdd.n1454 vdd.n1167 146.341
R17108 vdd.n1460 vdd.n1167 146.341
R17109 vdd.n1460 vdd.n1160 146.341
R17110 vdd.n1470 vdd.n1160 146.341
R17111 vdd.n1470 vdd.n1156 146.341
R17112 vdd.n1476 vdd.n1156 146.341
R17113 vdd.n1476 vdd.n1148 146.341
R17114 vdd.n1487 vdd.n1148 146.341
R17115 vdd.n1487 vdd.n1144 146.341
R17116 vdd.n1493 vdd.n1144 146.341
R17117 vdd.n1493 vdd.n1137 146.341
R17118 vdd.n1503 vdd.n1137 146.341
R17119 vdd.n1503 vdd.n1133 146.341
R17120 vdd.n1816 vdd.n1133 146.341
R17121 vdd.n1816 vdd.n1125 146.341
R17122 vdd.n1827 vdd.n1125 146.341
R17123 vdd.n1827 vdd.n1121 146.341
R17124 vdd.n1833 vdd.n1121 146.341
R17125 vdd.n1833 vdd.n1114 146.341
R17126 vdd.n1844 vdd.n1114 146.341
R17127 vdd.n1844 vdd.n1110 146.341
R17128 vdd.n1850 vdd.n1110 146.341
R17129 vdd.n1850 vdd.n1103 146.341
R17130 vdd.n1860 vdd.n1103 146.341
R17131 vdd.n1860 vdd.n1099 146.341
R17132 vdd.n1866 vdd.n1099 146.341
R17133 vdd.n1866 vdd.n1091 146.341
R17134 vdd.n1877 vdd.n1091 146.341
R17135 vdd.n1877 vdd.n1087 146.341
R17136 vdd.n1883 vdd.n1087 146.341
R17137 vdd.n1883 vdd.n1079 146.341
R17138 vdd.n1896 vdd.n1079 146.341
R17139 vdd.n1896 vdd.n1074 146.341
R17140 vdd.n2328 vdd.n1074 146.341
R17141 vdd.n1073 vdd.n1049 141.707
R17142 vdd.n3223 vdd.n692 141.707
R17143 vdd.n2177 vdd.t87 127.284
R17144 vdd.n965 vdd.t71 127.284
R17145 vdd.n2151 vdd.t109 127.284
R17146 vdd.n957 vdd.t96 127.284
R17147 vdd.n2922 vdd.t47 127.284
R17148 vdd.n2922 vdd.t48 127.284
R17149 vdd.n2642 vdd.t94 127.284
R17150 vdd.n832 vdd.t75 127.284
R17151 vdd.n2639 vdd.t80 127.284
R17152 vdd.n799 vdd.t82 127.284
R17153 vdd.n1027 vdd.t90 127.284
R17154 vdd.n1027 vdd.t91 127.284
R17155 vdd.n22 vdd.n20 117.314
R17156 vdd.n17 vdd.n15 117.314
R17157 vdd.n27 vdd.n26 116.927
R17158 vdd.n24 vdd.n23 116.927
R17159 vdd.n22 vdd.n21 116.927
R17160 vdd.n17 vdd.n16 116.927
R17161 vdd.n19 vdd.n18 116.927
R17162 vdd.n27 vdd.n25 116.927
R17163 vdd.n2178 vdd.t86 111.188
R17164 vdd.n966 vdd.t72 111.188
R17165 vdd.n2152 vdd.t108 111.188
R17166 vdd.n958 vdd.t97 111.188
R17167 vdd.n2643 vdd.t93 111.188
R17168 vdd.n833 vdd.t76 111.188
R17169 vdd.n2640 vdd.t79 111.188
R17170 vdd.n800 vdd.t83 111.188
R17171 vdd.n2865 vdd.n911 99.5127
R17172 vdd.n2869 vdd.n911 99.5127
R17173 vdd.n2869 vdd.n903 99.5127
R17174 vdd.n2877 vdd.n903 99.5127
R17175 vdd.n2877 vdd.n901 99.5127
R17176 vdd.n2881 vdd.n901 99.5127
R17177 vdd.n2881 vdd.n890 99.5127
R17178 vdd.n2889 vdd.n890 99.5127
R17179 vdd.n2889 vdd.n888 99.5127
R17180 vdd.n2893 vdd.n888 99.5127
R17181 vdd.n2893 vdd.n879 99.5127
R17182 vdd.n2901 vdd.n879 99.5127
R17183 vdd.n2901 vdd.n877 99.5127
R17184 vdd.n2905 vdd.n877 99.5127
R17185 vdd.n2905 vdd.n867 99.5127
R17186 vdd.n2913 vdd.n867 99.5127
R17187 vdd.n2913 vdd.n865 99.5127
R17188 vdd.n2917 vdd.n865 99.5127
R17189 vdd.n2917 vdd.n856 99.5127
R17190 vdd.n2927 vdd.n856 99.5127
R17191 vdd.n2927 vdd.n854 99.5127
R17192 vdd.n2931 vdd.n854 99.5127
R17193 vdd.n2931 vdd.n842 99.5127
R17194 vdd.n2984 vdd.n842 99.5127
R17195 vdd.n2984 vdd.n840 99.5127
R17196 vdd.n2988 vdd.n840 99.5127
R17197 vdd.n2988 vdd.n808 99.5127
R17198 vdd.n3058 vdd.n808 99.5127
R17199 vdd.n3054 vdd.n809 99.5127
R17200 vdd.n3052 vdd.n3051 99.5127
R17201 vdd.n3049 vdd.n813 99.5127
R17202 vdd.n3045 vdd.n3044 99.5127
R17203 vdd.n3042 vdd.n816 99.5127
R17204 vdd.n3038 vdd.n3037 99.5127
R17205 vdd.n3035 vdd.n819 99.5127
R17206 vdd.n3031 vdd.n3030 99.5127
R17207 vdd.n3028 vdd.n3026 99.5127
R17208 vdd.n3024 vdd.n822 99.5127
R17209 vdd.n3020 vdd.n3019 99.5127
R17210 vdd.n3017 vdd.n825 99.5127
R17211 vdd.n3013 vdd.n3012 99.5127
R17212 vdd.n3010 vdd.n828 99.5127
R17213 vdd.n3006 vdd.n3005 99.5127
R17214 vdd.n3003 vdd.n831 99.5127
R17215 vdd.n2998 vdd.n2997 99.5127
R17216 vdd.n2785 vdd.n914 99.5127
R17217 vdd.n2785 vdd.n909 99.5127
R17218 vdd.n2782 vdd.n909 99.5127
R17219 vdd.n2782 vdd.n904 99.5127
R17220 vdd.n2729 vdd.n904 99.5127
R17221 vdd.n2729 vdd.n898 99.5127
R17222 vdd.n2732 vdd.n898 99.5127
R17223 vdd.n2732 vdd.n891 99.5127
R17224 vdd.n2735 vdd.n891 99.5127
R17225 vdd.n2735 vdd.n886 99.5127
R17226 vdd.n2738 vdd.n886 99.5127
R17227 vdd.n2738 vdd.n881 99.5127
R17228 vdd.n2741 vdd.n881 99.5127
R17229 vdd.n2741 vdd.n875 99.5127
R17230 vdd.n2759 vdd.n875 99.5127
R17231 vdd.n2759 vdd.n868 99.5127
R17232 vdd.n2755 vdd.n868 99.5127
R17233 vdd.n2755 vdd.n863 99.5127
R17234 vdd.n2752 vdd.n863 99.5127
R17235 vdd.n2752 vdd.n858 99.5127
R17236 vdd.n2749 vdd.n858 99.5127
R17237 vdd.n2749 vdd.n852 99.5127
R17238 vdd.n2746 vdd.n852 99.5127
R17239 vdd.n2746 vdd.n844 99.5127
R17240 vdd.n844 vdd.n837 99.5127
R17241 vdd.n2990 vdd.n837 99.5127
R17242 vdd.n2991 vdd.n2990 99.5127
R17243 vdd.n2991 vdd.n806 99.5127
R17244 vdd.n2855 vdd.n2638 99.5127
R17245 vdd.n2851 vdd.n2638 99.5127
R17246 vdd.n2849 vdd.n2848 99.5127
R17247 vdd.n2845 vdd.n2844 99.5127
R17248 vdd.n2841 vdd.n2840 99.5127
R17249 vdd.n2837 vdd.n2836 99.5127
R17250 vdd.n2833 vdd.n2832 99.5127
R17251 vdd.n2829 vdd.n2828 99.5127
R17252 vdd.n2825 vdd.n2824 99.5127
R17253 vdd.n2821 vdd.n2820 99.5127
R17254 vdd.n2817 vdd.n2816 99.5127
R17255 vdd.n2813 vdd.n2812 99.5127
R17256 vdd.n2809 vdd.n2808 99.5127
R17257 vdd.n2805 vdd.n2804 99.5127
R17258 vdd.n2801 vdd.n2800 99.5127
R17259 vdd.n2797 vdd.n2796 99.5127
R17260 vdd.n2792 vdd.n2791 99.5127
R17261 vdd.n2603 vdd.n955 99.5127
R17262 vdd.n2599 vdd.n2598 99.5127
R17263 vdd.n2595 vdd.n2594 99.5127
R17264 vdd.n2591 vdd.n2590 99.5127
R17265 vdd.n2587 vdd.n2586 99.5127
R17266 vdd.n2583 vdd.n2582 99.5127
R17267 vdd.n2579 vdd.n2578 99.5127
R17268 vdd.n2575 vdd.n2574 99.5127
R17269 vdd.n2571 vdd.n2570 99.5127
R17270 vdd.n2567 vdd.n2566 99.5127
R17271 vdd.n2563 vdd.n2562 99.5127
R17272 vdd.n2559 vdd.n2558 99.5127
R17273 vdd.n2555 vdd.n2554 99.5127
R17274 vdd.n2551 vdd.n2550 99.5127
R17275 vdd.n2547 vdd.n2546 99.5127
R17276 vdd.n2543 vdd.n2542 99.5127
R17277 vdd.n2538 vdd.n2537 99.5127
R17278 vdd.n2276 vdd.n1050 99.5127
R17279 vdd.n2276 vdd.n1044 99.5127
R17280 vdd.n2273 vdd.n1044 99.5127
R17281 vdd.n2273 vdd.n1038 99.5127
R17282 vdd.n2270 vdd.n1038 99.5127
R17283 vdd.n2270 vdd.n1031 99.5127
R17284 vdd.n2267 vdd.n1031 99.5127
R17285 vdd.n2267 vdd.n1024 99.5127
R17286 vdd.n2264 vdd.n1024 99.5127
R17287 vdd.n2264 vdd.n1019 99.5127
R17288 vdd.n2261 vdd.n1019 99.5127
R17289 vdd.n2261 vdd.n1013 99.5127
R17290 vdd.n2258 vdd.n1013 99.5127
R17291 vdd.n2258 vdd.n1006 99.5127
R17292 vdd.n2172 vdd.n1006 99.5127
R17293 vdd.n2172 vdd.n1000 99.5127
R17294 vdd.n2169 vdd.n1000 99.5127
R17295 vdd.n2169 vdd.n995 99.5127
R17296 vdd.n2166 vdd.n995 99.5127
R17297 vdd.n2166 vdd.n990 99.5127
R17298 vdd.n2163 vdd.n990 99.5127
R17299 vdd.n2163 vdd.n984 99.5127
R17300 vdd.n2160 vdd.n984 99.5127
R17301 vdd.n2160 vdd.n977 99.5127
R17302 vdd.n2157 vdd.n977 99.5127
R17303 vdd.n2157 vdd.n970 99.5127
R17304 vdd.n970 vdd.n960 99.5127
R17305 vdd.n2533 vdd.n960 99.5127
R17306 vdd.n2111 vdd.n2109 99.5127
R17307 vdd.n2115 vdd.n2109 99.5127
R17308 vdd.n2119 vdd.n2117 99.5127
R17309 vdd.n2123 vdd.n2107 99.5127
R17310 vdd.n2127 vdd.n2125 99.5127
R17311 vdd.n2131 vdd.n2105 99.5127
R17312 vdd.n2135 vdd.n2133 99.5127
R17313 vdd.n2139 vdd.n2103 99.5127
R17314 vdd.n2142 vdd.n2141 99.5127
R17315 vdd.n2312 vdd.n2310 99.5127
R17316 vdd.n2308 vdd.n2144 99.5127
R17317 vdd.n2304 vdd.n2302 99.5127
R17318 vdd.n2300 vdd.n2146 99.5127
R17319 vdd.n2296 vdd.n2294 99.5127
R17320 vdd.n2292 vdd.n2148 99.5127
R17321 vdd.n2288 vdd.n2286 99.5127
R17322 vdd.n2284 vdd.n2150 99.5127
R17323 vdd.n2376 vdd.n1046 99.5127
R17324 vdd.n2380 vdd.n1046 99.5127
R17325 vdd.n2380 vdd.n1036 99.5127
R17326 vdd.n2388 vdd.n1036 99.5127
R17327 vdd.n2388 vdd.n1034 99.5127
R17328 vdd.n2392 vdd.n1034 99.5127
R17329 vdd.n2392 vdd.n1023 99.5127
R17330 vdd.n2401 vdd.n1023 99.5127
R17331 vdd.n2401 vdd.n1021 99.5127
R17332 vdd.n2405 vdd.n1021 99.5127
R17333 vdd.n2405 vdd.n1011 99.5127
R17334 vdd.n2413 vdd.n1011 99.5127
R17335 vdd.n2413 vdd.n1009 99.5127
R17336 vdd.n2417 vdd.n1009 99.5127
R17337 vdd.n2417 vdd.n999 99.5127
R17338 vdd.n2425 vdd.n999 99.5127
R17339 vdd.n2425 vdd.n997 99.5127
R17340 vdd.n2429 vdd.n997 99.5127
R17341 vdd.n2429 vdd.n988 99.5127
R17342 vdd.n2437 vdd.n988 99.5127
R17343 vdd.n2437 vdd.n986 99.5127
R17344 vdd.n2441 vdd.n986 99.5127
R17345 vdd.n2441 vdd.n975 99.5127
R17346 vdd.n2451 vdd.n975 99.5127
R17347 vdd.n2451 vdd.n972 99.5127
R17348 vdd.n2456 vdd.n972 99.5127
R17349 vdd.n2456 vdd.n973 99.5127
R17350 vdd.n973 vdd.n954 99.5127
R17351 vdd.n2974 vdd.n2973 99.5127
R17352 vdd.n2971 vdd.n2937 99.5127
R17353 vdd.n2967 vdd.n2966 99.5127
R17354 vdd.n2964 vdd.n2940 99.5127
R17355 vdd.n2960 vdd.n2959 99.5127
R17356 vdd.n2957 vdd.n2943 99.5127
R17357 vdd.n2953 vdd.n2952 99.5127
R17358 vdd.n2950 vdd.n2947 99.5127
R17359 vdd.n3091 vdd.n787 99.5127
R17360 vdd.n3089 vdd.n3088 99.5127
R17361 vdd.n3086 vdd.n789 99.5127
R17362 vdd.n3082 vdd.n3081 99.5127
R17363 vdd.n3079 vdd.n792 99.5127
R17364 vdd.n3075 vdd.n3074 99.5127
R17365 vdd.n3072 vdd.n795 99.5127
R17366 vdd.n3068 vdd.n3067 99.5127
R17367 vdd.n3065 vdd.n798 99.5127
R17368 vdd.n2709 vdd.n915 99.5127
R17369 vdd.n2709 vdd.n910 99.5127
R17370 vdd.n2780 vdd.n910 99.5127
R17371 vdd.n2780 vdd.n905 99.5127
R17372 vdd.n2776 vdd.n905 99.5127
R17373 vdd.n2776 vdd.n899 99.5127
R17374 vdd.n2773 vdd.n899 99.5127
R17375 vdd.n2773 vdd.n892 99.5127
R17376 vdd.n2770 vdd.n892 99.5127
R17377 vdd.n2770 vdd.n887 99.5127
R17378 vdd.n2767 vdd.n887 99.5127
R17379 vdd.n2767 vdd.n882 99.5127
R17380 vdd.n2764 vdd.n882 99.5127
R17381 vdd.n2764 vdd.n876 99.5127
R17382 vdd.n2761 vdd.n876 99.5127
R17383 vdd.n2761 vdd.n869 99.5127
R17384 vdd.n2726 vdd.n869 99.5127
R17385 vdd.n2726 vdd.n864 99.5127
R17386 vdd.n2723 vdd.n864 99.5127
R17387 vdd.n2723 vdd.n859 99.5127
R17388 vdd.n2720 vdd.n859 99.5127
R17389 vdd.n2720 vdd.n853 99.5127
R17390 vdd.n2717 vdd.n853 99.5127
R17391 vdd.n2717 vdd.n845 99.5127
R17392 vdd.n2714 vdd.n845 99.5127
R17393 vdd.n2714 vdd.n838 99.5127
R17394 vdd.n838 vdd.n804 99.5127
R17395 vdd.n3060 vdd.n804 99.5127
R17396 vdd.n2859 vdd.n918 99.5127
R17397 vdd.n2647 vdd.n2646 99.5127
R17398 vdd.n2651 vdd.n2650 99.5127
R17399 vdd.n2655 vdd.n2654 99.5127
R17400 vdd.n2659 vdd.n2658 99.5127
R17401 vdd.n2663 vdd.n2662 99.5127
R17402 vdd.n2667 vdd.n2666 99.5127
R17403 vdd.n2671 vdd.n2670 99.5127
R17404 vdd.n2675 vdd.n2674 99.5127
R17405 vdd.n2679 vdd.n2678 99.5127
R17406 vdd.n2683 vdd.n2682 99.5127
R17407 vdd.n2687 vdd.n2686 99.5127
R17408 vdd.n2691 vdd.n2690 99.5127
R17409 vdd.n2695 vdd.n2694 99.5127
R17410 vdd.n2699 vdd.n2698 99.5127
R17411 vdd.n2703 vdd.n2702 99.5127
R17412 vdd.n2705 vdd.n2637 99.5127
R17413 vdd.n2863 vdd.n908 99.5127
R17414 vdd.n2871 vdd.n908 99.5127
R17415 vdd.n2871 vdd.n906 99.5127
R17416 vdd.n2875 vdd.n906 99.5127
R17417 vdd.n2875 vdd.n896 99.5127
R17418 vdd.n2883 vdd.n896 99.5127
R17419 vdd.n2883 vdd.n894 99.5127
R17420 vdd.n2887 vdd.n894 99.5127
R17421 vdd.n2887 vdd.n885 99.5127
R17422 vdd.n2895 vdd.n885 99.5127
R17423 vdd.n2895 vdd.n883 99.5127
R17424 vdd.n2899 vdd.n883 99.5127
R17425 vdd.n2899 vdd.n873 99.5127
R17426 vdd.n2907 vdd.n873 99.5127
R17427 vdd.n2907 vdd.n871 99.5127
R17428 vdd.n2911 vdd.n871 99.5127
R17429 vdd.n2911 vdd.n862 99.5127
R17430 vdd.n2919 vdd.n862 99.5127
R17431 vdd.n2919 vdd.n860 99.5127
R17432 vdd.n2925 vdd.n860 99.5127
R17433 vdd.n2925 vdd.n850 99.5127
R17434 vdd.n2933 vdd.n850 99.5127
R17435 vdd.n2933 vdd.n847 99.5127
R17436 vdd.n2982 vdd.n847 99.5127
R17437 vdd.n2982 vdd.n848 99.5127
R17438 vdd.n848 vdd.n839 99.5127
R17439 vdd.n2977 vdd.n839 99.5127
R17440 vdd.n2977 vdd.n807 99.5127
R17441 vdd.n2527 vdd.n2526 99.5127
R17442 vdd.n2523 vdd.n2522 99.5127
R17443 vdd.n2519 vdd.n2518 99.5127
R17444 vdd.n2515 vdd.n2514 99.5127
R17445 vdd.n2511 vdd.n2510 99.5127
R17446 vdd.n2507 vdd.n2506 99.5127
R17447 vdd.n2503 vdd.n2502 99.5127
R17448 vdd.n2499 vdd.n2498 99.5127
R17449 vdd.n2495 vdd.n2494 99.5127
R17450 vdd.n2491 vdd.n2490 99.5127
R17451 vdd.n2487 vdd.n2486 99.5127
R17452 vdd.n2483 vdd.n2482 99.5127
R17453 vdd.n2479 vdd.n2478 99.5127
R17454 vdd.n2475 vdd.n2474 99.5127
R17455 vdd.n2471 vdd.n2470 99.5127
R17456 vdd.n2467 vdd.n2466 99.5127
R17457 vdd.n2463 vdd.n936 99.5127
R17458 vdd.n2220 vdd.n1051 99.5127
R17459 vdd.n2220 vdd.n1045 99.5127
R17460 vdd.n2223 vdd.n1045 99.5127
R17461 vdd.n2223 vdd.n1039 99.5127
R17462 vdd.n2226 vdd.n1039 99.5127
R17463 vdd.n2226 vdd.n1032 99.5127
R17464 vdd.n2229 vdd.n1032 99.5127
R17465 vdd.n2229 vdd.n1025 99.5127
R17466 vdd.n2232 vdd.n1025 99.5127
R17467 vdd.n2232 vdd.n1020 99.5127
R17468 vdd.n2235 vdd.n1020 99.5127
R17469 vdd.n2235 vdd.n1014 99.5127
R17470 vdd.n2256 vdd.n1014 99.5127
R17471 vdd.n2256 vdd.n1007 99.5127
R17472 vdd.n2252 vdd.n1007 99.5127
R17473 vdd.n2252 vdd.n1001 99.5127
R17474 vdd.n2249 vdd.n1001 99.5127
R17475 vdd.n2249 vdd.n996 99.5127
R17476 vdd.n2246 vdd.n996 99.5127
R17477 vdd.n2246 vdd.n991 99.5127
R17478 vdd.n2243 vdd.n991 99.5127
R17479 vdd.n2243 vdd.n985 99.5127
R17480 vdd.n2240 vdd.n985 99.5127
R17481 vdd.n2240 vdd.n978 99.5127
R17482 vdd.n978 vdd.n969 99.5127
R17483 vdd.n2458 vdd.n969 99.5127
R17484 vdd.n2459 vdd.n2458 99.5127
R17485 vdd.n2459 vdd.n961 99.5127
R17486 vdd.n2370 vdd.n2368 99.5127
R17487 vdd.n2366 vdd.n1054 99.5127
R17488 vdd.n2362 vdd.n2360 99.5127
R17489 vdd.n2358 vdd.n1056 99.5127
R17490 vdd.n2354 vdd.n2352 99.5127
R17491 vdd.n2350 vdd.n1058 99.5127
R17492 vdd.n2346 vdd.n2344 99.5127
R17493 vdd.n2342 vdd.n1060 99.5127
R17494 vdd.n2184 vdd.n1062 99.5127
R17495 vdd.n2189 vdd.n2186 99.5127
R17496 vdd.n2193 vdd.n2191 99.5127
R17497 vdd.n2197 vdd.n2182 99.5127
R17498 vdd.n2201 vdd.n2199 99.5127
R17499 vdd.n2205 vdd.n2180 99.5127
R17500 vdd.n2209 vdd.n2207 99.5127
R17501 vdd.n2214 vdd.n2176 99.5127
R17502 vdd.n2217 vdd.n2216 99.5127
R17503 vdd.n2374 vdd.n1042 99.5127
R17504 vdd.n2382 vdd.n1042 99.5127
R17505 vdd.n2382 vdd.n1040 99.5127
R17506 vdd.n2386 vdd.n1040 99.5127
R17507 vdd.n2386 vdd.n1029 99.5127
R17508 vdd.n2394 vdd.n1029 99.5127
R17509 vdd.n2394 vdd.n1026 99.5127
R17510 vdd.n2399 vdd.n1026 99.5127
R17511 vdd.n2399 vdd.n1017 99.5127
R17512 vdd.n2407 vdd.n1017 99.5127
R17513 vdd.n2407 vdd.n1015 99.5127
R17514 vdd.n2411 vdd.n1015 99.5127
R17515 vdd.n2411 vdd.n1005 99.5127
R17516 vdd.n2419 vdd.n1005 99.5127
R17517 vdd.n2419 vdd.n1003 99.5127
R17518 vdd.n2423 vdd.n1003 99.5127
R17519 vdd.n2423 vdd.n994 99.5127
R17520 vdd.n2431 vdd.n994 99.5127
R17521 vdd.n2431 vdd.n992 99.5127
R17522 vdd.n2435 vdd.n992 99.5127
R17523 vdd.n2435 vdd.n982 99.5127
R17524 vdd.n2443 vdd.n982 99.5127
R17525 vdd.n2443 vdd.n979 99.5127
R17526 vdd.n2449 vdd.n979 99.5127
R17527 vdd.n2449 vdd.n980 99.5127
R17528 vdd.n980 vdd.n971 99.5127
R17529 vdd.n971 vdd.n962 99.5127
R17530 vdd.n2531 vdd.n962 99.5127
R17531 vdd.n9 vdd.n7 98.9633
R17532 vdd.n2 vdd.n0 98.9633
R17533 vdd.n9 vdd.n8 98.6055
R17534 vdd.n11 vdd.n10 98.6055
R17535 vdd.n13 vdd.n12 98.6055
R17536 vdd.n6 vdd.n5 98.6055
R17537 vdd.n4 vdd.n3 98.6055
R17538 vdd.n2 vdd.n1 98.6055
R17539 vdd.t254 vdd.n303 85.8723
R17540 vdd.t226 vdd.n244 85.8723
R17541 vdd.t241 vdd.n201 85.8723
R17542 vdd.t212 vdd.n142 85.8723
R17543 vdd.t190 vdd.n100 85.8723
R17544 vdd.t126 vdd.n41 85.8723
R17545 vdd.t272 vdd.n1722 85.8723
R17546 vdd.t156 vdd.n1781 85.8723
R17547 vdd.t256 vdd.n1620 85.8723
R17548 vdd.t130 vdd.n1679 85.8723
R17549 vdd.t124 vdd.n1519 85.8723
R17550 vdd.t192 vdd.n1578 85.8723
R17551 vdd.n2923 vdd.n2922 78.546
R17552 vdd.n2397 vdd.n1027 78.546
R17553 vdd.n290 vdd.n289 75.1835
R17554 vdd.n288 vdd.n287 75.1835
R17555 vdd.n286 vdd.n285 75.1835
R17556 vdd.n284 vdd.n283 75.1835
R17557 vdd.n282 vdd.n281 75.1835
R17558 vdd.n280 vdd.n279 75.1835
R17559 vdd.n278 vdd.n277 75.1835
R17560 vdd.n276 vdd.n275 75.1835
R17561 vdd.n274 vdd.n273 75.1835
R17562 vdd.n188 vdd.n187 75.1835
R17563 vdd.n186 vdd.n185 75.1835
R17564 vdd.n184 vdd.n183 75.1835
R17565 vdd.n182 vdd.n181 75.1835
R17566 vdd.n180 vdd.n179 75.1835
R17567 vdd.n178 vdd.n177 75.1835
R17568 vdd.n176 vdd.n175 75.1835
R17569 vdd.n174 vdd.n173 75.1835
R17570 vdd.n172 vdd.n171 75.1835
R17571 vdd.n87 vdd.n86 75.1835
R17572 vdd.n85 vdd.n84 75.1835
R17573 vdd.n83 vdd.n82 75.1835
R17574 vdd.n81 vdd.n80 75.1835
R17575 vdd.n79 vdd.n78 75.1835
R17576 vdd.n77 vdd.n76 75.1835
R17577 vdd.n75 vdd.n74 75.1835
R17578 vdd.n73 vdd.n72 75.1835
R17579 vdd.n71 vdd.n70 75.1835
R17580 vdd.n1752 vdd.n1751 75.1835
R17581 vdd.n1754 vdd.n1753 75.1835
R17582 vdd.n1756 vdd.n1755 75.1835
R17583 vdd.n1758 vdd.n1757 75.1835
R17584 vdd.n1760 vdd.n1759 75.1835
R17585 vdd.n1762 vdd.n1761 75.1835
R17586 vdd.n1764 vdd.n1763 75.1835
R17587 vdd.n1766 vdd.n1765 75.1835
R17588 vdd.n1768 vdd.n1767 75.1835
R17589 vdd.n1650 vdd.n1649 75.1835
R17590 vdd.n1652 vdd.n1651 75.1835
R17591 vdd.n1654 vdd.n1653 75.1835
R17592 vdd.n1656 vdd.n1655 75.1835
R17593 vdd.n1658 vdd.n1657 75.1835
R17594 vdd.n1660 vdd.n1659 75.1835
R17595 vdd.n1662 vdd.n1661 75.1835
R17596 vdd.n1664 vdd.n1663 75.1835
R17597 vdd.n1666 vdd.n1665 75.1835
R17598 vdd.n1549 vdd.n1548 75.1835
R17599 vdd.n1551 vdd.n1550 75.1835
R17600 vdd.n1553 vdd.n1552 75.1835
R17601 vdd.n1555 vdd.n1554 75.1835
R17602 vdd.n1557 vdd.n1556 75.1835
R17603 vdd.n1559 vdd.n1558 75.1835
R17604 vdd.n1561 vdd.n1560 75.1835
R17605 vdd.n1563 vdd.n1562 75.1835
R17606 vdd.n1565 vdd.n1564 75.1835
R17607 vdd.n2858 vdd.n2857 72.8958
R17608 vdd.n2857 vdd.n2621 72.8958
R17609 vdd.n2857 vdd.n2622 72.8958
R17610 vdd.n2857 vdd.n2623 72.8958
R17611 vdd.n2857 vdd.n2624 72.8958
R17612 vdd.n2857 vdd.n2625 72.8958
R17613 vdd.n2857 vdd.n2626 72.8958
R17614 vdd.n2857 vdd.n2627 72.8958
R17615 vdd.n2857 vdd.n2628 72.8958
R17616 vdd.n2857 vdd.n2629 72.8958
R17617 vdd.n2857 vdd.n2630 72.8958
R17618 vdd.n2857 vdd.n2631 72.8958
R17619 vdd.n2857 vdd.n2632 72.8958
R17620 vdd.n2857 vdd.n2633 72.8958
R17621 vdd.n2857 vdd.n2634 72.8958
R17622 vdd.n2857 vdd.n2635 72.8958
R17623 vdd.n2857 vdd.n2636 72.8958
R17624 vdd.n803 vdd.n692 72.8958
R17625 vdd.n3066 vdd.n692 72.8958
R17626 vdd.n797 vdd.n692 72.8958
R17627 vdd.n3073 vdd.n692 72.8958
R17628 vdd.n794 vdd.n692 72.8958
R17629 vdd.n3080 vdd.n692 72.8958
R17630 vdd.n791 vdd.n692 72.8958
R17631 vdd.n3087 vdd.n692 72.8958
R17632 vdd.n3090 vdd.n692 72.8958
R17633 vdd.n2946 vdd.n692 72.8958
R17634 vdd.n2951 vdd.n692 72.8958
R17635 vdd.n2945 vdd.n692 72.8958
R17636 vdd.n2958 vdd.n692 72.8958
R17637 vdd.n2942 vdd.n692 72.8958
R17638 vdd.n2965 vdd.n692 72.8958
R17639 vdd.n2939 vdd.n692 72.8958
R17640 vdd.n2972 vdd.n692 72.8958
R17641 vdd.n2110 vdd.n1049 72.8958
R17642 vdd.n2116 vdd.n1049 72.8958
R17643 vdd.n2118 vdd.n1049 72.8958
R17644 vdd.n2124 vdd.n1049 72.8958
R17645 vdd.n2126 vdd.n1049 72.8958
R17646 vdd.n2132 vdd.n1049 72.8958
R17647 vdd.n2134 vdd.n1049 72.8958
R17648 vdd.n2140 vdd.n1049 72.8958
R17649 vdd.n2311 vdd.n1049 72.8958
R17650 vdd.n2309 vdd.n1049 72.8958
R17651 vdd.n2303 vdd.n1049 72.8958
R17652 vdd.n2301 vdd.n1049 72.8958
R17653 vdd.n2295 vdd.n1049 72.8958
R17654 vdd.n2293 vdd.n1049 72.8958
R17655 vdd.n2287 vdd.n1049 72.8958
R17656 vdd.n2285 vdd.n1049 72.8958
R17657 vdd.n2279 vdd.n1049 72.8958
R17658 vdd.n2604 vdd.n937 72.8958
R17659 vdd.n2604 vdd.n938 72.8958
R17660 vdd.n2604 vdd.n939 72.8958
R17661 vdd.n2604 vdd.n940 72.8958
R17662 vdd.n2604 vdd.n941 72.8958
R17663 vdd.n2604 vdd.n942 72.8958
R17664 vdd.n2604 vdd.n943 72.8958
R17665 vdd.n2604 vdd.n944 72.8958
R17666 vdd.n2604 vdd.n945 72.8958
R17667 vdd.n2604 vdd.n946 72.8958
R17668 vdd.n2604 vdd.n947 72.8958
R17669 vdd.n2604 vdd.n948 72.8958
R17670 vdd.n2604 vdd.n949 72.8958
R17671 vdd.n2604 vdd.n950 72.8958
R17672 vdd.n2604 vdd.n951 72.8958
R17673 vdd.n2604 vdd.n952 72.8958
R17674 vdd.n2604 vdd.n953 72.8958
R17675 vdd.n2857 vdd.n2856 72.8958
R17676 vdd.n2857 vdd.n2605 72.8958
R17677 vdd.n2857 vdd.n2606 72.8958
R17678 vdd.n2857 vdd.n2607 72.8958
R17679 vdd.n2857 vdd.n2608 72.8958
R17680 vdd.n2857 vdd.n2609 72.8958
R17681 vdd.n2857 vdd.n2610 72.8958
R17682 vdd.n2857 vdd.n2611 72.8958
R17683 vdd.n2857 vdd.n2612 72.8958
R17684 vdd.n2857 vdd.n2613 72.8958
R17685 vdd.n2857 vdd.n2614 72.8958
R17686 vdd.n2857 vdd.n2615 72.8958
R17687 vdd.n2857 vdd.n2616 72.8958
R17688 vdd.n2857 vdd.n2617 72.8958
R17689 vdd.n2857 vdd.n2618 72.8958
R17690 vdd.n2857 vdd.n2619 72.8958
R17691 vdd.n2857 vdd.n2620 72.8958
R17692 vdd.n2996 vdd.n692 72.8958
R17693 vdd.n835 vdd.n692 72.8958
R17694 vdd.n3004 vdd.n692 72.8958
R17695 vdd.n830 vdd.n692 72.8958
R17696 vdd.n3011 vdd.n692 72.8958
R17697 vdd.n827 vdd.n692 72.8958
R17698 vdd.n3018 vdd.n692 72.8958
R17699 vdd.n824 vdd.n692 72.8958
R17700 vdd.n3025 vdd.n692 72.8958
R17701 vdd.n3029 vdd.n692 72.8958
R17702 vdd.n821 vdd.n692 72.8958
R17703 vdd.n3036 vdd.n692 72.8958
R17704 vdd.n818 vdd.n692 72.8958
R17705 vdd.n3043 vdd.n692 72.8958
R17706 vdd.n815 vdd.n692 72.8958
R17707 vdd.n3050 vdd.n692 72.8958
R17708 vdd.n3053 vdd.n692 72.8958
R17709 vdd.n2604 vdd.n935 72.8958
R17710 vdd.n2604 vdd.n934 72.8958
R17711 vdd.n2604 vdd.n933 72.8958
R17712 vdd.n2604 vdd.n932 72.8958
R17713 vdd.n2604 vdd.n931 72.8958
R17714 vdd.n2604 vdd.n930 72.8958
R17715 vdd.n2604 vdd.n929 72.8958
R17716 vdd.n2604 vdd.n928 72.8958
R17717 vdd.n2604 vdd.n927 72.8958
R17718 vdd.n2604 vdd.n926 72.8958
R17719 vdd.n2604 vdd.n925 72.8958
R17720 vdd.n2604 vdd.n924 72.8958
R17721 vdd.n2604 vdd.n923 72.8958
R17722 vdd.n2604 vdd.n922 72.8958
R17723 vdd.n2604 vdd.n921 72.8958
R17724 vdd.n2604 vdd.n920 72.8958
R17725 vdd.n2604 vdd.n919 72.8958
R17726 vdd.n2369 vdd.n1049 72.8958
R17727 vdd.n2367 vdd.n1049 72.8958
R17728 vdd.n2361 vdd.n1049 72.8958
R17729 vdd.n2359 vdd.n1049 72.8958
R17730 vdd.n2353 vdd.n1049 72.8958
R17731 vdd.n2351 vdd.n1049 72.8958
R17732 vdd.n2345 vdd.n1049 72.8958
R17733 vdd.n2343 vdd.n1049 72.8958
R17734 vdd.n1061 vdd.n1049 72.8958
R17735 vdd.n2185 vdd.n1049 72.8958
R17736 vdd.n2190 vdd.n1049 72.8958
R17737 vdd.n2192 vdd.n1049 72.8958
R17738 vdd.n2198 vdd.n1049 72.8958
R17739 vdd.n2200 vdd.n1049 72.8958
R17740 vdd.n2206 vdd.n1049 72.8958
R17741 vdd.n2208 vdd.n1049 72.8958
R17742 vdd.n2215 vdd.n1049 72.8958
R17743 vdd.n1419 vdd.n1418 66.2847
R17744 vdd.n1418 vdd.n1194 66.2847
R17745 vdd.n1418 vdd.n1195 66.2847
R17746 vdd.n1418 vdd.n1196 66.2847
R17747 vdd.n1418 vdd.n1197 66.2847
R17748 vdd.n1418 vdd.n1198 66.2847
R17749 vdd.n1418 vdd.n1199 66.2847
R17750 vdd.n1418 vdd.n1200 66.2847
R17751 vdd.n1418 vdd.n1201 66.2847
R17752 vdd.n1418 vdd.n1202 66.2847
R17753 vdd.n1418 vdd.n1203 66.2847
R17754 vdd.n1418 vdd.n1204 66.2847
R17755 vdd.n1418 vdd.n1205 66.2847
R17756 vdd.n1418 vdd.n1206 66.2847
R17757 vdd.n1418 vdd.n1207 66.2847
R17758 vdd.n1418 vdd.n1208 66.2847
R17759 vdd.n1418 vdd.n1209 66.2847
R17760 vdd.n1418 vdd.n1210 66.2847
R17761 vdd.n1418 vdd.n1211 66.2847
R17762 vdd.n1418 vdd.n1212 66.2847
R17763 vdd.n1418 vdd.n1213 66.2847
R17764 vdd.n1418 vdd.n1214 66.2847
R17765 vdd.n1418 vdd.n1215 66.2847
R17766 vdd.n1418 vdd.n1216 66.2847
R17767 vdd.n1418 vdd.n1217 66.2847
R17768 vdd.n1418 vdd.n1218 66.2847
R17769 vdd.n1418 vdd.n1219 66.2847
R17770 vdd.n1418 vdd.n1220 66.2847
R17771 vdd.n1418 vdd.n1221 66.2847
R17772 vdd.n1418 vdd.n1222 66.2847
R17773 vdd.n1418 vdd.n1223 66.2847
R17774 vdd.n1073 vdd.n1070 66.2847
R17775 vdd.n2000 vdd.n1073 66.2847
R17776 vdd.n2005 vdd.n1073 66.2847
R17777 vdd.n2010 vdd.n1073 66.2847
R17778 vdd.n1998 vdd.n1073 66.2847
R17779 vdd.n2017 vdd.n1073 66.2847
R17780 vdd.n1990 vdd.n1073 66.2847
R17781 vdd.n2024 vdd.n1073 66.2847
R17782 vdd.n1983 vdd.n1073 66.2847
R17783 vdd.n2031 vdd.n1073 66.2847
R17784 vdd.n1977 vdd.n1073 66.2847
R17785 vdd.n1972 vdd.n1073 66.2847
R17786 vdd.n2042 vdd.n1073 66.2847
R17787 vdd.n1964 vdd.n1073 66.2847
R17788 vdd.n2049 vdd.n1073 66.2847
R17789 vdd.n1957 vdd.n1073 66.2847
R17790 vdd.n2056 vdd.n1073 66.2847
R17791 vdd.n1950 vdd.n1073 66.2847
R17792 vdd.n2063 vdd.n1073 66.2847
R17793 vdd.n1943 vdd.n1073 66.2847
R17794 vdd.n2070 vdd.n1073 66.2847
R17795 vdd.n1937 vdd.n1073 66.2847
R17796 vdd.n1932 vdd.n1073 66.2847
R17797 vdd.n2081 vdd.n1073 66.2847
R17798 vdd.n1924 vdd.n1073 66.2847
R17799 vdd.n2088 vdd.n1073 66.2847
R17800 vdd.n1917 vdd.n1073 66.2847
R17801 vdd.n2095 vdd.n1073 66.2847
R17802 vdd.n2098 vdd.n1073 66.2847
R17803 vdd.n1908 vdd.n1073 66.2847
R17804 vdd.n2320 vdd.n1073 66.2847
R17805 vdd.n1902 vdd.n1073 66.2847
R17806 vdd.n3223 vdd.n3222 66.2847
R17807 vdd.n3223 vdd.n693 66.2847
R17808 vdd.n3223 vdd.n694 66.2847
R17809 vdd.n3223 vdd.n695 66.2847
R17810 vdd.n3223 vdd.n696 66.2847
R17811 vdd.n3223 vdd.n697 66.2847
R17812 vdd.n3223 vdd.n698 66.2847
R17813 vdd.n3223 vdd.n699 66.2847
R17814 vdd.n3223 vdd.n700 66.2847
R17815 vdd.n3223 vdd.n701 66.2847
R17816 vdd.n3223 vdd.n702 66.2847
R17817 vdd.n3223 vdd.n703 66.2847
R17818 vdd.n3223 vdd.n704 66.2847
R17819 vdd.n3223 vdd.n705 66.2847
R17820 vdd.n3223 vdd.n706 66.2847
R17821 vdd.n3223 vdd.n707 66.2847
R17822 vdd.n3223 vdd.n708 66.2847
R17823 vdd.n3223 vdd.n709 66.2847
R17824 vdd.n3223 vdd.n710 66.2847
R17825 vdd.n3223 vdd.n711 66.2847
R17826 vdd.n3223 vdd.n712 66.2847
R17827 vdd.n3223 vdd.n713 66.2847
R17828 vdd.n3223 vdd.n714 66.2847
R17829 vdd.n3223 vdd.n715 66.2847
R17830 vdd.n3223 vdd.n716 66.2847
R17831 vdd.n3223 vdd.n717 66.2847
R17832 vdd.n3223 vdd.n718 66.2847
R17833 vdd.n3223 vdd.n719 66.2847
R17834 vdd.n3223 vdd.n720 66.2847
R17835 vdd.n3223 vdd.n721 66.2847
R17836 vdd.n3223 vdd.n722 66.2847
R17837 vdd.n3354 vdd.n3353 66.2847
R17838 vdd.n3354 vdd.n424 66.2847
R17839 vdd.n3354 vdd.n423 66.2847
R17840 vdd.n3354 vdd.n422 66.2847
R17841 vdd.n3354 vdd.n421 66.2847
R17842 vdd.n3354 vdd.n420 66.2847
R17843 vdd.n3354 vdd.n419 66.2847
R17844 vdd.n3354 vdd.n418 66.2847
R17845 vdd.n3354 vdd.n417 66.2847
R17846 vdd.n3354 vdd.n416 66.2847
R17847 vdd.n3354 vdd.n415 66.2847
R17848 vdd.n3354 vdd.n414 66.2847
R17849 vdd.n3354 vdd.n413 66.2847
R17850 vdd.n3354 vdd.n412 66.2847
R17851 vdd.n3354 vdd.n411 66.2847
R17852 vdd.n3354 vdd.n410 66.2847
R17853 vdd.n3354 vdd.n409 66.2847
R17854 vdd.n3354 vdd.n408 66.2847
R17855 vdd.n3354 vdd.n407 66.2847
R17856 vdd.n3354 vdd.n406 66.2847
R17857 vdd.n3354 vdd.n405 66.2847
R17858 vdd.n3354 vdd.n404 66.2847
R17859 vdd.n3354 vdd.n403 66.2847
R17860 vdd.n3354 vdd.n402 66.2847
R17861 vdd.n3354 vdd.n401 66.2847
R17862 vdd.n3354 vdd.n400 66.2847
R17863 vdd.n3354 vdd.n399 66.2847
R17864 vdd.n3354 vdd.n398 66.2847
R17865 vdd.n3354 vdd.n397 66.2847
R17866 vdd.n3354 vdd.n396 66.2847
R17867 vdd.n3354 vdd.n395 66.2847
R17868 vdd.n3354 vdd.n394 66.2847
R17869 vdd.n467 vdd.n394 52.4337
R17870 vdd.n473 vdd.n395 52.4337
R17871 vdd.n477 vdd.n396 52.4337
R17872 vdd.n483 vdd.n397 52.4337
R17873 vdd.n487 vdd.n398 52.4337
R17874 vdd.n493 vdd.n399 52.4337
R17875 vdd.n497 vdd.n400 52.4337
R17876 vdd.n503 vdd.n401 52.4337
R17877 vdd.n507 vdd.n402 52.4337
R17878 vdd.n513 vdd.n403 52.4337
R17879 vdd.n517 vdd.n404 52.4337
R17880 vdd.n523 vdd.n405 52.4337
R17881 vdd.n527 vdd.n406 52.4337
R17882 vdd.n533 vdd.n407 52.4337
R17883 vdd.n537 vdd.n408 52.4337
R17884 vdd.n543 vdd.n409 52.4337
R17885 vdd.n547 vdd.n410 52.4337
R17886 vdd.n553 vdd.n411 52.4337
R17887 vdd.n557 vdd.n412 52.4337
R17888 vdd.n563 vdd.n413 52.4337
R17889 vdd.n567 vdd.n414 52.4337
R17890 vdd.n573 vdd.n415 52.4337
R17891 vdd.n577 vdd.n416 52.4337
R17892 vdd.n583 vdd.n417 52.4337
R17893 vdd.n587 vdd.n418 52.4337
R17894 vdd.n593 vdd.n419 52.4337
R17895 vdd.n597 vdd.n420 52.4337
R17896 vdd.n603 vdd.n421 52.4337
R17897 vdd.n607 vdd.n422 52.4337
R17898 vdd.n613 vdd.n423 52.4337
R17899 vdd.n616 vdd.n424 52.4337
R17900 vdd.n3353 vdd.n3352 52.4337
R17901 vdd.n3222 vdd.n3221 52.4337
R17902 vdd.n728 vdd.n693 52.4337
R17903 vdd.n734 vdd.n694 52.4337
R17904 vdd.n3211 vdd.n695 52.4337
R17905 vdd.n3207 vdd.n696 52.4337
R17906 vdd.n3203 vdd.n697 52.4337
R17907 vdd.n3199 vdd.n698 52.4337
R17908 vdd.n3195 vdd.n699 52.4337
R17909 vdd.n3191 vdd.n700 52.4337
R17910 vdd.n3187 vdd.n701 52.4337
R17911 vdd.n3179 vdd.n702 52.4337
R17912 vdd.n3175 vdd.n703 52.4337
R17913 vdd.n3171 vdd.n704 52.4337
R17914 vdd.n3167 vdd.n705 52.4337
R17915 vdd.n3163 vdd.n706 52.4337
R17916 vdd.n3159 vdd.n707 52.4337
R17917 vdd.n3155 vdd.n708 52.4337
R17918 vdd.n3151 vdd.n709 52.4337
R17919 vdd.n3147 vdd.n710 52.4337
R17920 vdd.n3143 vdd.n711 52.4337
R17921 vdd.n3139 vdd.n712 52.4337
R17922 vdd.n3133 vdd.n713 52.4337
R17923 vdd.n3129 vdd.n714 52.4337
R17924 vdd.n3125 vdd.n715 52.4337
R17925 vdd.n3121 vdd.n716 52.4337
R17926 vdd.n3117 vdd.n717 52.4337
R17927 vdd.n3113 vdd.n718 52.4337
R17928 vdd.n3109 vdd.n719 52.4337
R17929 vdd.n3105 vdd.n720 52.4337
R17930 vdd.n3101 vdd.n721 52.4337
R17931 vdd.n3097 vdd.n722 52.4337
R17932 vdd.n2322 vdd.n1902 52.4337
R17933 vdd.n2320 vdd.n2319 52.4337
R17934 vdd.n1909 vdd.n1908 52.4337
R17935 vdd.n2098 vdd.n2097 52.4337
R17936 vdd.n2095 vdd.n2094 52.4337
R17937 vdd.n2090 vdd.n1917 52.4337
R17938 vdd.n2088 vdd.n2087 52.4337
R17939 vdd.n2083 vdd.n1924 52.4337
R17940 vdd.n2081 vdd.n2080 52.4337
R17941 vdd.n1933 vdd.n1932 52.4337
R17942 vdd.n2072 vdd.n1937 52.4337
R17943 vdd.n2070 vdd.n2069 52.4337
R17944 vdd.n2065 vdd.n1943 52.4337
R17945 vdd.n2063 vdd.n2062 52.4337
R17946 vdd.n2058 vdd.n1950 52.4337
R17947 vdd.n2056 vdd.n2055 52.4337
R17948 vdd.n2051 vdd.n1957 52.4337
R17949 vdd.n2049 vdd.n2048 52.4337
R17950 vdd.n2044 vdd.n1964 52.4337
R17951 vdd.n2042 vdd.n2041 52.4337
R17952 vdd.n1973 vdd.n1972 52.4337
R17953 vdd.n2033 vdd.n1977 52.4337
R17954 vdd.n2031 vdd.n2030 52.4337
R17955 vdd.n2026 vdd.n1983 52.4337
R17956 vdd.n2024 vdd.n2023 52.4337
R17957 vdd.n2019 vdd.n1990 52.4337
R17958 vdd.n2017 vdd.n2016 52.4337
R17959 vdd.n2012 vdd.n1998 52.4337
R17960 vdd.n2010 vdd.n2009 52.4337
R17961 vdd.n2005 vdd.n2004 52.4337
R17962 vdd.n2000 vdd.n1999 52.4337
R17963 vdd.n2331 vdd.n1070 52.4337
R17964 vdd.n1420 vdd.n1419 52.4337
R17965 vdd.n1226 vdd.n1194 52.4337
R17966 vdd.n1230 vdd.n1195 52.4337
R17967 vdd.n1232 vdd.n1196 52.4337
R17968 vdd.n1236 vdd.n1197 52.4337
R17969 vdd.n1238 vdd.n1198 52.4337
R17970 vdd.n1242 vdd.n1199 52.4337
R17971 vdd.n1244 vdd.n1200 52.4337
R17972 vdd.n1248 vdd.n1201 52.4337
R17973 vdd.n1250 vdd.n1202 52.4337
R17974 vdd.n1256 vdd.n1203 52.4337
R17975 vdd.n1258 vdd.n1204 52.4337
R17976 vdd.n1262 vdd.n1205 52.4337
R17977 vdd.n1264 vdd.n1206 52.4337
R17978 vdd.n1268 vdd.n1207 52.4337
R17979 vdd.n1270 vdd.n1208 52.4337
R17980 vdd.n1274 vdd.n1209 52.4337
R17981 vdd.n1276 vdd.n1210 52.4337
R17982 vdd.n1280 vdd.n1211 52.4337
R17983 vdd.n1282 vdd.n1212 52.4337
R17984 vdd.n1354 vdd.n1213 52.4337
R17985 vdd.n1287 vdd.n1214 52.4337
R17986 vdd.n1291 vdd.n1215 52.4337
R17987 vdd.n1293 vdd.n1216 52.4337
R17988 vdd.n1297 vdd.n1217 52.4337
R17989 vdd.n1299 vdd.n1218 52.4337
R17990 vdd.n1303 vdd.n1219 52.4337
R17991 vdd.n1305 vdd.n1220 52.4337
R17992 vdd.n1309 vdd.n1221 52.4337
R17993 vdd.n1311 vdd.n1222 52.4337
R17994 vdd.n1315 vdd.n1223 52.4337
R17995 vdd.n1419 vdd.n1193 52.4337
R17996 vdd.n1229 vdd.n1194 52.4337
R17997 vdd.n1231 vdd.n1195 52.4337
R17998 vdd.n1235 vdd.n1196 52.4337
R17999 vdd.n1237 vdd.n1197 52.4337
R18000 vdd.n1241 vdd.n1198 52.4337
R18001 vdd.n1243 vdd.n1199 52.4337
R18002 vdd.n1247 vdd.n1200 52.4337
R18003 vdd.n1249 vdd.n1201 52.4337
R18004 vdd.n1255 vdd.n1202 52.4337
R18005 vdd.n1257 vdd.n1203 52.4337
R18006 vdd.n1261 vdd.n1204 52.4337
R18007 vdd.n1263 vdd.n1205 52.4337
R18008 vdd.n1267 vdd.n1206 52.4337
R18009 vdd.n1269 vdd.n1207 52.4337
R18010 vdd.n1273 vdd.n1208 52.4337
R18011 vdd.n1275 vdd.n1209 52.4337
R18012 vdd.n1279 vdd.n1210 52.4337
R18013 vdd.n1281 vdd.n1211 52.4337
R18014 vdd.n1285 vdd.n1212 52.4337
R18015 vdd.n1286 vdd.n1213 52.4337
R18016 vdd.n1290 vdd.n1214 52.4337
R18017 vdd.n1292 vdd.n1215 52.4337
R18018 vdd.n1296 vdd.n1216 52.4337
R18019 vdd.n1298 vdd.n1217 52.4337
R18020 vdd.n1302 vdd.n1218 52.4337
R18021 vdd.n1304 vdd.n1219 52.4337
R18022 vdd.n1308 vdd.n1220 52.4337
R18023 vdd.n1310 vdd.n1221 52.4337
R18024 vdd.n1314 vdd.n1222 52.4337
R18025 vdd.n1316 vdd.n1223 52.4337
R18026 vdd.n1070 vdd.n1069 52.4337
R18027 vdd.n2001 vdd.n2000 52.4337
R18028 vdd.n2006 vdd.n2005 52.4337
R18029 vdd.n2011 vdd.n2010 52.4337
R18030 vdd.n1998 vdd.n1991 52.4337
R18031 vdd.n2018 vdd.n2017 52.4337
R18032 vdd.n1990 vdd.n1984 52.4337
R18033 vdd.n2025 vdd.n2024 52.4337
R18034 vdd.n1983 vdd.n1978 52.4337
R18035 vdd.n2032 vdd.n2031 52.4337
R18036 vdd.n1977 vdd.n1976 52.4337
R18037 vdd.n1972 vdd.n1965 52.4337
R18038 vdd.n2043 vdd.n2042 52.4337
R18039 vdd.n1964 vdd.n1958 52.4337
R18040 vdd.n2050 vdd.n2049 52.4337
R18041 vdd.n1957 vdd.n1951 52.4337
R18042 vdd.n2057 vdd.n2056 52.4337
R18043 vdd.n1950 vdd.n1944 52.4337
R18044 vdd.n2064 vdd.n2063 52.4337
R18045 vdd.n1943 vdd.n1938 52.4337
R18046 vdd.n2071 vdd.n2070 52.4337
R18047 vdd.n1937 vdd.n1936 52.4337
R18048 vdd.n1932 vdd.n1925 52.4337
R18049 vdd.n2082 vdd.n2081 52.4337
R18050 vdd.n1924 vdd.n1918 52.4337
R18051 vdd.n2089 vdd.n2088 52.4337
R18052 vdd.n1917 vdd.n1911 52.4337
R18053 vdd.n2096 vdd.n2095 52.4337
R18054 vdd.n2099 vdd.n2098 52.4337
R18055 vdd.n1908 vdd.n1903 52.4337
R18056 vdd.n2321 vdd.n2320 52.4337
R18057 vdd.n1902 vdd.n1075 52.4337
R18058 vdd.n3222 vdd.n725 52.4337
R18059 vdd.n733 vdd.n693 52.4337
R18060 vdd.n3212 vdd.n694 52.4337
R18061 vdd.n3208 vdd.n695 52.4337
R18062 vdd.n3204 vdd.n696 52.4337
R18063 vdd.n3200 vdd.n697 52.4337
R18064 vdd.n3196 vdd.n698 52.4337
R18065 vdd.n3192 vdd.n699 52.4337
R18066 vdd.n3188 vdd.n700 52.4337
R18067 vdd.n3178 vdd.n701 52.4337
R18068 vdd.n3176 vdd.n702 52.4337
R18069 vdd.n3172 vdd.n703 52.4337
R18070 vdd.n3168 vdd.n704 52.4337
R18071 vdd.n3164 vdd.n705 52.4337
R18072 vdd.n3160 vdd.n706 52.4337
R18073 vdd.n3156 vdd.n707 52.4337
R18074 vdd.n3152 vdd.n708 52.4337
R18075 vdd.n3148 vdd.n709 52.4337
R18076 vdd.n3144 vdd.n710 52.4337
R18077 vdd.n3140 vdd.n711 52.4337
R18078 vdd.n3132 vdd.n712 52.4337
R18079 vdd.n3130 vdd.n713 52.4337
R18080 vdd.n3126 vdd.n714 52.4337
R18081 vdd.n3122 vdd.n715 52.4337
R18082 vdd.n3118 vdd.n716 52.4337
R18083 vdd.n3114 vdd.n717 52.4337
R18084 vdd.n3110 vdd.n718 52.4337
R18085 vdd.n3106 vdd.n719 52.4337
R18086 vdd.n3102 vdd.n720 52.4337
R18087 vdd.n3098 vdd.n721 52.4337
R18088 vdd.n722 vdd.n691 52.4337
R18089 vdd.n3353 vdd.n425 52.4337
R18090 vdd.n614 vdd.n424 52.4337
R18091 vdd.n608 vdd.n423 52.4337
R18092 vdd.n604 vdd.n422 52.4337
R18093 vdd.n598 vdd.n421 52.4337
R18094 vdd.n594 vdd.n420 52.4337
R18095 vdd.n588 vdd.n419 52.4337
R18096 vdd.n584 vdd.n418 52.4337
R18097 vdd.n578 vdd.n417 52.4337
R18098 vdd.n574 vdd.n416 52.4337
R18099 vdd.n568 vdd.n415 52.4337
R18100 vdd.n564 vdd.n414 52.4337
R18101 vdd.n558 vdd.n413 52.4337
R18102 vdd.n554 vdd.n412 52.4337
R18103 vdd.n548 vdd.n411 52.4337
R18104 vdd.n544 vdd.n410 52.4337
R18105 vdd.n538 vdd.n409 52.4337
R18106 vdd.n534 vdd.n408 52.4337
R18107 vdd.n528 vdd.n407 52.4337
R18108 vdd.n524 vdd.n406 52.4337
R18109 vdd.n518 vdd.n405 52.4337
R18110 vdd.n514 vdd.n404 52.4337
R18111 vdd.n508 vdd.n403 52.4337
R18112 vdd.n504 vdd.n402 52.4337
R18113 vdd.n498 vdd.n401 52.4337
R18114 vdd.n494 vdd.n400 52.4337
R18115 vdd.n488 vdd.n399 52.4337
R18116 vdd.n484 vdd.n398 52.4337
R18117 vdd.n478 vdd.n397 52.4337
R18118 vdd.n474 vdd.n396 52.4337
R18119 vdd.n468 vdd.n395 52.4337
R18120 vdd.n394 vdd.n392 52.4337
R18121 vdd.t111 vdd.t286 51.4683
R18122 vdd.n274 vdd.n272 42.0461
R18123 vdd.n172 vdd.n170 42.0461
R18124 vdd.n71 vdd.n69 42.0461
R18125 vdd.n1752 vdd.n1750 42.0461
R18126 vdd.n1650 vdd.n1648 42.0461
R18127 vdd.n1549 vdd.n1547 42.0461
R18128 vdd.n332 vdd.n331 41.6884
R18129 vdd.n230 vdd.n229 41.6884
R18130 vdd.n129 vdd.n128 41.6884
R18131 vdd.n1810 vdd.n1809 41.6884
R18132 vdd.n1708 vdd.n1707 41.6884
R18133 vdd.n1607 vdd.n1606 41.6884
R18134 vdd.n1319 vdd.n1318 41.1157
R18135 vdd.n1357 vdd.n1356 41.1157
R18136 vdd.n1253 vdd.n1252 41.1157
R18137 vdd.n428 vdd.n427 41.1157
R18138 vdd.n566 vdd.n441 41.1157
R18139 vdd.n454 vdd.n453 41.1157
R18140 vdd.n3053 vdd.n3052 39.2114
R18141 vdd.n3050 vdd.n3049 39.2114
R18142 vdd.n3045 vdd.n815 39.2114
R18143 vdd.n3043 vdd.n3042 39.2114
R18144 vdd.n3038 vdd.n818 39.2114
R18145 vdd.n3036 vdd.n3035 39.2114
R18146 vdd.n3031 vdd.n821 39.2114
R18147 vdd.n3029 vdd.n3028 39.2114
R18148 vdd.n3025 vdd.n3024 39.2114
R18149 vdd.n3020 vdd.n824 39.2114
R18150 vdd.n3018 vdd.n3017 39.2114
R18151 vdd.n3013 vdd.n827 39.2114
R18152 vdd.n3011 vdd.n3010 39.2114
R18153 vdd.n3006 vdd.n830 39.2114
R18154 vdd.n3004 vdd.n3003 39.2114
R18155 vdd.n2998 vdd.n835 39.2114
R18156 vdd.n2996 vdd.n2995 39.2114
R18157 vdd.n2856 vdd.n913 39.2114
R18158 vdd.n2851 vdd.n2605 39.2114
R18159 vdd.n2848 vdd.n2606 39.2114
R18160 vdd.n2844 vdd.n2607 39.2114
R18161 vdd.n2840 vdd.n2608 39.2114
R18162 vdd.n2836 vdd.n2609 39.2114
R18163 vdd.n2832 vdd.n2610 39.2114
R18164 vdd.n2828 vdd.n2611 39.2114
R18165 vdd.n2824 vdd.n2612 39.2114
R18166 vdd.n2820 vdd.n2613 39.2114
R18167 vdd.n2816 vdd.n2614 39.2114
R18168 vdd.n2812 vdd.n2615 39.2114
R18169 vdd.n2808 vdd.n2616 39.2114
R18170 vdd.n2804 vdd.n2617 39.2114
R18171 vdd.n2800 vdd.n2618 39.2114
R18172 vdd.n2796 vdd.n2619 39.2114
R18173 vdd.n2791 vdd.n2620 39.2114
R18174 vdd.n2599 vdd.n953 39.2114
R18175 vdd.n2595 vdd.n952 39.2114
R18176 vdd.n2591 vdd.n951 39.2114
R18177 vdd.n2587 vdd.n950 39.2114
R18178 vdd.n2583 vdd.n949 39.2114
R18179 vdd.n2579 vdd.n948 39.2114
R18180 vdd.n2575 vdd.n947 39.2114
R18181 vdd.n2571 vdd.n946 39.2114
R18182 vdd.n2567 vdd.n945 39.2114
R18183 vdd.n2563 vdd.n944 39.2114
R18184 vdd.n2559 vdd.n943 39.2114
R18185 vdd.n2555 vdd.n942 39.2114
R18186 vdd.n2551 vdd.n941 39.2114
R18187 vdd.n2547 vdd.n940 39.2114
R18188 vdd.n2543 vdd.n939 39.2114
R18189 vdd.n2538 vdd.n938 39.2114
R18190 vdd.n2534 vdd.n937 39.2114
R18191 vdd.n2110 vdd.n1048 39.2114
R18192 vdd.n2116 vdd.n2115 39.2114
R18193 vdd.n2119 vdd.n2118 39.2114
R18194 vdd.n2124 vdd.n2123 39.2114
R18195 vdd.n2127 vdd.n2126 39.2114
R18196 vdd.n2132 vdd.n2131 39.2114
R18197 vdd.n2135 vdd.n2134 39.2114
R18198 vdd.n2140 vdd.n2139 39.2114
R18199 vdd.n2311 vdd.n2142 39.2114
R18200 vdd.n2310 vdd.n2309 39.2114
R18201 vdd.n2303 vdd.n2144 39.2114
R18202 vdd.n2302 vdd.n2301 39.2114
R18203 vdd.n2295 vdd.n2146 39.2114
R18204 vdd.n2294 vdd.n2293 39.2114
R18205 vdd.n2287 vdd.n2148 39.2114
R18206 vdd.n2286 vdd.n2285 39.2114
R18207 vdd.n2279 vdd.n2150 39.2114
R18208 vdd.n2972 vdd.n2971 39.2114
R18209 vdd.n2967 vdd.n2939 39.2114
R18210 vdd.n2965 vdd.n2964 39.2114
R18211 vdd.n2960 vdd.n2942 39.2114
R18212 vdd.n2958 vdd.n2957 39.2114
R18213 vdd.n2953 vdd.n2945 39.2114
R18214 vdd.n2951 vdd.n2950 39.2114
R18215 vdd.n2946 vdd.n787 39.2114
R18216 vdd.n3090 vdd.n3089 39.2114
R18217 vdd.n3087 vdd.n3086 39.2114
R18218 vdd.n3082 vdd.n791 39.2114
R18219 vdd.n3080 vdd.n3079 39.2114
R18220 vdd.n3075 vdd.n794 39.2114
R18221 vdd.n3073 vdd.n3072 39.2114
R18222 vdd.n3068 vdd.n797 39.2114
R18223 vdd.n3066 vdd.n3065 39.2114
R18224 vdd.n3061 vdd.n803 39.2114
R18225 vdd.n2858 vdd.n916 39.2114
R18226 vdd.n2621 vdd.n918 39.2114
R18227 vdd.n2647 vdd.n2622 39.2114
R18228 vdd.n2651 vdd.n2623 39.2114
R18229 vdd.n2655 vdd.n2624 39.2114
R18230 vdd.n2659 vdd.n2625 39.2114
R18231 vdd.n2663 vdd.n2626 39.2114
R18232 vdd.n2667 vdd.n2627 39.2114
R18233 vdd.n2671 vdd.n2628 39.2114
R18234 vdd.n2675 vdd.n2629 39.2114
R18235 vdd.n2679 vdd.n2630 39.2114
R18236 vdd.n2683 vdd.n2631 39.2114
R18237 vdd.n2687 vdd.n2632 39.2114
R18238 vdd.n2691 vdd.n2633 39.2114
R18239 vdd.n2695 vdd.n2634 39.2114
R18240 vdd.n2699 vdd.n2635 39.2114
R18241 vdd.n2703 vdd.n2636 39.2114
R18242 vdd.n2859 vdd.n2858 39.2114
R18243 vdd.n2646 vdd.n2621 39.2114
R18244 vdd.n2650 vdd.n2622 39.2114
R18245 vdd.n2654 vdd.n2623 39.2114
R18246 vdd.n2658 vdd.n2624 39.2114
R18247 vdd.n2662 vdd.n2625 39.2114
R18248 vdd.n2666 vdd.n2626 39.2114
R18249 vdd.n2670 vdd.n2627 39.2114
R18250 vdd.n2674 vdd.n2628 39.2114
R18251 vdd.n2678 vdd.n2629 39.2114
R18252 vdd.n2682 vdd.n2630 39.2114
R18253 vdd.n2686 vdd.n2631 39.2114
R18254 vdd.n2690 vdd.n2632 39.2114
R18255 vdd.n2694 vdd.n2633 39.2114
R18256 vdd.n2698 vdd.n2634 39.2114
R18257 vdd.n2702 vdd.n2635 39.2114
R18258 vdd.n2705 vdd.n2636 39.2114
R18259 vdd.n803 vdd.n798 39.2114
R18260 vdd.n3067 vdd.n3066 39.2114
R18261 vdd.n797 vdd.n795 39.2114
R18262 vdd.n3074 vdd.n3073 39.2114
R18263 vdd.n794 vdd.n792 39.2114
R18264 vdd.n3081 vdd.n3080 39.2114
R18265 vdd.n791 vdd.n789 39.2114
R18266 vdd.n3088 vdd.n3087 39.2114
R18267 vdd.n3091 vdd.n3090 39.2114
R18268 vdd.n2947 vdd.n2946 39.2114
R18269 vdd.n2952 vdd.n2951 39.2114
R18270 vdd.n2945 vdd.n2943 39.2114
R18271 vdd.n2959 vdd.n2958 39.2114
R18272 vdd.n2942 vdd.n2940 39.2114
R18273 vdd.n2966 vdd.n2965 39.2114
R18274 vdd.n2939 vdd.n2937 39.2114
R18275 vdd.n2973 vdd.n2972 39.2114
R18276 vdd.n2111 vdd.n2110 39.2114
R18277 vdd.n2117 vdd.n2116 39.2114
R18278 vdd.n2118 vdd.n2107 39.2114
R18279 vdd.n2125 vdd.n2124 39.2114
R18280 vdd.n2126 vdd.n2105 39.2114
R18281 vdd.n2133 vdd.n2132 39.2114
R18282 vdd.n2134 vdd.n2103 39.2114
R18283 vdd.n2141 vdd.n2140 39.2114
R18284 vdd.n2312 vdd.n2311 39.2114
R18285 vdd.n2309 vdd.n2308 39.2114
R18286 vdd.n2304 vdd.n2303 39.2114
R18287 vdd.n2301 vdd.n2300 39.2114
R18288 vdd.n2296 vdd.n2295 39.2114
R18289 vdd.n2293 vdd.n2292 39.2114
R18290 vdd.n2288 vdd.n2287 39.2114
R18291 vdd.n2285 vdd.n2284 39.2114
R18292 vdd.n2280 vdd.n2279 39.2114
R18293 vdd.n2537 vdd.n937 39.2114
R18294 vdd.n2542 vdd.n938 39.2114
R18295 vdd.n2546 vdd.n939 39.2114
R18296 vdd.n2550 vdd.n940 39.2114
R18297 vdd.n2554 vdd.n941 39.2114
R18298 vdd.n2558 vdd.n942 39.2114
R18299 vdd.n2562 vdd.n943 39.2114
R18300 vdd.n2566 vdd.n944 39.2114
R18301 vdd.n2570 vdd.n945 39.2114
R18302 vdd.n2574 vdd.n946 39.2114
R18303 vdd.n2578 vdd.n947 39.2114
R18304 vdd.n2582 vdd.n948 39.2114
R18305 vdd.n2586 vdd.n949 39.2114
R18306 vdd.n2590 vdd.n950 39.2114
R18307 vdd.n2594 vdd.n951 39.2114
R18308 vdd.n2598 vdd.n952 39.2114
R18309 vdd.n955 vdd.n953 39.2114
R18310 vdd.n2856 vdd.n2855 39.2114
R18311 vdd.n2849 vdd.n2605 39.2114
R18312 vdd.n2845 vdd.n2606 39.2114
R18313 vdd.n2841 vdd.n2607 39.2114
R18314 vdd.n2837 vdd.n2608 39.2114
R18315 vdd.n2833 vdd.n2609 39.2114
R18316 vdd.n2829 vdd.n2610 39.2114
R18317 vdd.n2825 vdd.n2611 39.2114
R18318 vdd.n2821 vdd.n2612 39.2114
R18319 vdd.n2817 vdd.n2613 39.2114
R18320 vdd.n2813 vdd.n2614 39.2114
R18321 vdd.n2809 vdd.n2615 39.2114
R18322 vdd.n2805 vdd.n2616 39.2114
R18323 vdd.n2801 vdd.n2617 39.2114
R18324 vdd.n2797 vdd.n2618 39.2114
R18325 vdd.n2792 vdd.n2619 39.2114
R18326 vdd.n2788 vdd.n2620 39.2114
R18327 vdd.n2997 vdd.n2996 39.2114
R18328 vdd.n835 vdd.n831 39.2114
R18329 vdd.n3005 vdd.n3004 39.2114
R18330 vdd.n830 vdd.n828 39.2114
R18331 vdd.n3012 vdd.n3011 39.2114
R18332 vdd.n827 vdd.n825 39.2114
R18333 vdd.n3019 vdd.n3018 39.2114
R18334 vdd.n824 vdd.n822 39.2114
R18335 vdd.n3026 vdd.n3025 39.2114
R18336 vdd.n3030 vdd.n3029 39.2114
R18337 vdd.n821 vdd.n819 39.2114
R18338 vdd.n3037 vdd.n3036 39.2114
R18339 vdd.n818 vdd.n816 39.2114
R18340 vdd.n3044 vdd.n3043 39.2114
R18341 vdd.n815 vdd.n813 39.2114
R18342 vdd.n3051 vdd.n3050 39.2114
R18343 vdd.n3054 vdd.n3053 39.2114
R18344 vdd.n963 vdd.n919 39.2114
R18345 vdd.n2526 vdd.n920 39.2114
R18346 vdd.n2522 vdd.n921 39.2114
R18347 vdd.n2518 vdd.n922 39.2114
R18348 vdd.n2514 vdd.n923 39.2114
R18349 vdd.n2510 vdd.n924 39.2114
R18350 vdd.n2506 vdd.n925 39.2114
R18351 vdd.n2502 vdd.n926 39.2114
R18352 vdd.n2498 vdd.n927 39.2114
R18353 vdd.n2494 vdd.n928 39.2114
R18354 vdd.n2490 vdd.n929 39.2114
R18355 vdd.n2486 vdd.n930 39.2114
R18356 vdd.n2482 vdd.n931 39.2114
R18357 vdd.n2478 vdd.n932 39.2114
R18358 vdd.n2474 vdd.n933 39.2114
R18359 vdd.n2470 vdd.n934 39.2114
R18360 vdd.n2466 vdd.n935 39.2114
R18361 vdd.n2369 vdd.n1052 39.2114
R18362 vdd.n2368 vdd.n2367 39.2114
R18363 vdd.n2361 vdd.n1054 39.2114
R18364 vdd.n2360 vdd.n2359 39.2114
R18365 vdd.n2353 vdd.n1056 39.2114
R18366 vdd.n2352 vdd.n2351 39.2114
R18367 vdd.n2345 vdd.n1058 39.2114
R18368 vdd.n2344 vdd.n2343 39.2114
R18369 vdd.n1061 vdd.n1060 39.2114
R18370 vdd.n2185 vdd.n2184 39.2114
R18371 vdd.n2190 vdd.n2189 39.2114
R18372 vdd.n2193 vdd.n2192 39.2114
R18373 vdd.n2198 vdd.n2197 39.2114
R18374 vdd.n2201 vdd.n2200 39.2114
R18375 vdd.n2206 vdd.n2205 39.2114
R18376 vdd.n2209 vdd.n2208 39.2114
R18377 vdd.n2215 vdd.n2214 39.2114
R18378 vdd.n2463 vdd.n935 39.2114
R18379 vdd.n2467 vdd.n934 39.2114
R18380 vdd.n2471 vdd.n933 39.2114
R18381 vdd.n2475 vdd.n932 39.2114
R18382 vdd.n2479 vdd.n931 39.2114
R18383 vdd.n2483 vdd.n930 39.2114
R18384 vdd.n2487 vdd.n929 39.2114
R18385 vdd.n2491 vdd.n928 39.2114
R18386 vdd.n2495 vdd.n927 39.2114
R18387 vdd.n2499 vdd.n926 39.2114
R18388 vdd.n2503 vdd.n925 39.2114
R18389 vdd.n2507 vdd.n924 39.2114
R18390 vdd.n2511 vdd.n923 39.2114
R18391 vdd.n2515 vdd.n922 39.2114
R18392 vdd.n2519 vdd.n921 39.2114
R18393 vdd.n2523 vdd.n920 39.2114
R18394 vdd.n2527 vdd.n919 39.2114
R18395 vdd.n2370 vdd.n2369 39.2114
R18396 vdd.n2367 vdd.n2366 39.2114
R18397 vdd.n2362 vdd.n2361 39.2114
R18398 vdd.n2359 vdd.n2358 39.2114
R18399 vdd.n2354 vdd.n2353 39.2114
R18400 vdd.n2351 vdd.n2350 39.2114
R18401 vdd.n2346 vdd.n2345 39.2114
R18402 vdd.n2343 vdd.n2342 39.2114
R18403 vdd.n1062 vdd.n1061 39.2114
R18404 vdd.n2186 vdd.n2185 39.2114
R18405 vdd.n2191 vdd.n2190 39.2114
R18406 vdd.n2192 vdd.n2182 39.2114
R18407 vdd.n2199 vdd.n2198 39.2114
R18408 vdd.n2200 vdd.n2180 39.2114
R18409 vdd.n2207 vdd.n2206 39.2114
R18410 vdd.n2208 vdd.n2176 39.2114
R18411 vdd.n2216 vdd.n2215 39.2114
R18412 vdd.n2335 vdd.n2334 37.2369
R18413 vdd.n2038 vdd.n1971 37.2369
R18414 vdd.n2077 vdd.n1931 37.2369
R18415 vdd.n3138 vdd.n769 37.2369
R18416 vdd.n3186 vdd.n3185 37.2369
R18417 vdd.n690 vdd.n689 37.2369
R18418 vdd.n2377 vdd.n1047 31.6883
R18419 vdd.n2602 vdd.n956 31.6883
R18420 vdd.n2535 vdd.n959 31.6883
R18421 vdd.n2281 vdd.n2278 31.6883
R18422 vdd.n2789 vdd.n2787 31.6883
R18423 vdd.n2994 vdd.n2993 31.6883
R18424 vdd.n2866 vdd.n912 31.6883
R18425 vdd.n3057 vdd.n3056 31.6883
R18426 vdd.n2976 vdd.n2975 31.6883
R18427 vdd.n3062 vdd.n802 31.6883
R18428 vdd.n2708 vdd.n2707 31.6883
R18429 vdd.n2862 vdd.n2861 31.6883
R18430 vdd.n2373 vdd.n2372 31.6883
R18431 vdd.n2530 vdd.n2529 31.6883
R18432 vdd.n2462 vdd.n2461 31.6883
R18433 vdd.n2219 vdd.n2218 31.6883
R18434 vdd.n2212 vdd.n2178 30.449
R18435 vdd.n967 vdd.n966 30.449
R18436 vdd.n2153 vdd.n2152 30.449
R18437 vdd.n2540 vdd.n958 30.449
R18438 vdd.n2644 vdd.n2643 30.449
R18439 vdd.n3000 vdd.n833 30.449
R18440 vdd.n2794 vdd.n2640 30.449
R18441 vdd.n801 vdd.n800 30.449
R18442 vdd.n1418 vdd.n1225 22.2201
R18443 vdd.n2329 vdd.n1073 22.2201
R18444 vdd.n3223 vdd.n723 22.2201
R18445 vdd.n3355 vdd.n3354 22.2201
R18446 vdd.n1429 vdd.n1187 19.3944
R18447 vdd.n1429 vdd.n1185 19.3944
R18448 vdd.n1433 vdd.n1185 19.3944
R18449 vdd.n1433 vdd.n1175 19.3944
R18450 vdd.n1446 vdd.n1175 19.3944
R18451 vdd.n1446 vdd.n1173 19.3944
R18452 vdd.n1450 vdd.n1173 19.3944
R18453 vdd.n1450 vdd.n1165 19.3944
R18454 vdd.n1463 vdd.n1165 19.3944
R18455 vdd.n1463 vdd.n1163 19.3944
R18456 vdd.n1467 vdd.n1163 19.3944
R18457 vdd.n1467 vdd.n1152 19.3944
R18458 vdd.n1479 vdd.n1152 19.3944
R18459 vdd.n1479 vdd.n1150 19.3944
R18460 vdd.n1483 vdd.n1150 19.3944
R18461 vdd.n1483 vdd.n1141 19.3944
R18462 vdd.n1496 vdd.n1141 19.3944
R18463 vdd.n1496 vdd.n1139 19.3944
R18464 vdd.n1500 vdd.n1139 19.3944
R18465 vdd.n1500 vdd.n1130 19.3944
R18466 vdd.n1819 vdd.n1130 19.3944
R18467 vdd.n1819 vdd.n1128 19.3944
R18468 vdd.n1823 vdd.n1128 19.3944
R18469 vdd.n1823 vdd.n1118 19.3944
R18470 vdd.n1836 vdd.n1118 19.3944
R18471 vdd.n1836 vdd.n1116 19.3944
R18472 vdd.n1840 vdd.n1116 19.3944
R18473 vdd.n1840 vdd.n1108 19.3944
R18474 vdd.n1853 vdd.n1108 19.3944
R18475 vdd.n1853 vdd.n1106 19.3944
R18476 vdd.n1857 vdd.n1106 19.3944
R18477 vdd.n1857 vdd.n1095 19.3944
R18478 vdd.n1869 vdd.n1095 19.3944
R18479 vdd.n1869 vdd.n1093 19.3944
R18480 vdd.n1873 vdd.n1093 19.3944
R18481 vdd.n1873 vdd.n1085 19.3944
R18482 vdd.n1886 vdd.n1085 19.3944
R18483 vdd.n1886 vdd.n1082 19.3944
R18484 vdd.n1892 vdd.n1082 19.3944
R18485 vdd.n1892 vdd.n1083 19.3944
R18486 vdd.n1083 vdd.n1072 19.3944
R18487 vdd.n1353 vdd.n1288 19.3944
R18488 vdd.n1349 vdd.n1288 19.3944
R18489 vdd.n1349 vdd.n1348 19.3944
R18490 vdd.n1348 vdd.n1347 19.3944
R18491 vdd.n1347 vdd.n1294 19.3944
R18492 vdd.n1343 vdd.n1294 19.3944
R18493 vdd.n1343 vdd.n1342 19.3944
R18494 vdd.n1342 vdd.n1341 19.3944
R18495 vdd.n1341 vdd.n1300 19.3944
R18496 vdd.n1337 vdd.n1300 19.3944
R18497 vdd.n1337 vdd.n1336 19.3944
R18498 vdd.n1336 vdd.n1335 19.3944
R18499 vdd.n1335 vdd.n1306 19.3944
R18500 vdd.n1331 vdd.n1306 19.3944
R18501 vdd.n1331 vdd.n1330 19.3944
R18502 vdd.n1330 vdd.n1329 19.3944
R18503 vdd.n1329 vdd.n1312 19.3944
R18504 vdd.n1325 vdd.n1312 19.3944
R18505 vdd.n1325 vdd.n1324 19.3944
R18506 vdd.n1324 vdd.n1323 19.3944
R18507 vdd.n1388 vdd.n1387 19.3944
R18508 vdd.n1387 vdd.n1386 19.3944
R18509 vdd.n1386 vdd.n1259 19.3944
R18510 vdd.n1382 vdd.n1259 19.3944
R18511 vdd.n1382 vdd.n1381 19.3944
R18512 vdd.n1381 vdd.n1380 19.3944
R18513 vdd.n1380 vdd.n1265 19.3944
R18514 vdd.n1376 vdd.n1265 19.3944
R18515 vdd.n1376 vdd.n1375 19.3944
R18516 vdd.n1375 vdd.n1374 19.3944
R18517 vdd.n1374 vdd.n1271 19.3944
R18518 vdd.n1370 vdd.n1271 19.3944
R18519 vdd.n1370 vdd.n1369 19.3944
R18520 vdd.n1369 vdd.n1368 19.3944
R18521 vdd.n1368 vdd.n1277 19.3944
R18522 vdd.n1364 vdd.n1277 19.3944
R18523 vdd.n1364 vdd.n1363 19.3944
R18524 vdd.n1363 vdd.n1362 19.3944
R18525 vdd.n1362 vdd.n1283 19.3944
R18526 vdd.n1358 vdd.n1283 19.3944
R18527 vdd.n1421 vdd.n1192 19.3944
R18528 vdd.n1416 vdd.n1192 19.3944
R18529 vdd.n1416 vdd.n1227 19.3944
R18530 vdd.n1412 vdd.n1227 19.3944
R18531 vdd.n1412 vdd.n1411 19.3944
R18532 vdd.n1411 vdd.n1410 19.3944
R18533 vdd.n1410 vdd.n1233 19.3944
R18534 vdd.n1406 vdd.n1233 19.3944
R18535 vdd.n1406 vdd.n1405 19.3944
R18536 vdd.n1405 vdd.n1404 19.3944
R18537 vdd.n1404 vdd.n1239 19.3944
R18538 vdd.n1400 vdd.n1239 19.3944
R18539 vdd.n1400 vdd.n1399 19.3944
R18540 vdd.n1399 vdd.n1398 19.3944
R18541 vdd.n1398 vdd.n1245 19.3944
R18542 vdd.n1394 vdd.n1245 19.3944
R18543 vdd.n1394 vdd.n1393 19.3944
R18544 vdd.n1393 vdd.n1392 19.3944
R18545 vdd.n2034 vdd.n1969 19.3944
R18546 vdd.n2034 vdd.n1975 19.3944
R18547 vdd.n2029 vdd.n1975 19.3944
R18548 vdd.n2029 vdd.n2028 19.3944
R18549 vdd.n2028 vdd.n2027 19.3944
R18550 vdd.n2027 vdd.n1982 19.3944
R18551 vdd.n2022 vdd.n1982 19.3944
R18552 vdd.n2022 vdd.n2021 19.3944
R18553 vdd.n2021 vdd.n2020 19.3944
R18554 vdd.n2020 vdd.n1989 19.3944
R18555 vdd.n2015 vdd.n1989 19.3944
R18556 vdd.n2015 vdd.n2014 19.3944
R18557 vdd.n2014 vdd.n2013 19.3944
R18558 vdd.n2013 vdd.n1997 19.3944
R18559 vdd.n2008 vdd.n1997 19.3944
R18560 vdd.n2008 vdd.n2007 19.3944
R18561 vdd.n2003 vdd.n2002 19.3944
R18562 vdd.n2336 vdd.n1068 19.3944
R18563 vdd.n2073 vdd.n1929 19.3944
R18564 vdd.n2073 vdd.n1935 19.3944
R18565 vdd.n2068 vdd.n1935 19.3944
R18566 vdd.n2068 vdd.n2067 19.3944
R18567 vdd.n2067 vdd.n2066 19.3944
R18568 vdd.n2066 vdd.n1942 19.3944
R18569 vdd.n2061 vdd.n1942 19.3944
R18570 vdd.n2061 vdd.n2060 19.3944
R18571 vdd.n2060 vdd.n2059 19.3944
R18572 vdd.n2059 vdd.n1949 19.3944
R18573 vdd.n2054 vdd.n1949 19.3944
R18574 vdd.n2054 vdd.n2053 19.3944
R18575 vdd.n2053 vdd.n2052 19.3944
R18576 vdd.n2052 vdd.n1956 19.3944
R18577 vdd.n2047 vdd.n1956 19.3944
R18578 vdd.n2047 vdd.n2046 19.3944
R18579 vdd.n2046 vdd.n2045 19.3944
R18580 vdd.n2045 vdd.n1963 19.3944
R18581 vdd.n2040 vdd.n1963 19.3944
R18582 vdd.n2040 vdd.n2039 19.3944
R18583 vdd.n2324 vdd.n2323 19.3944
R18584 vdd.n2323 vdd.n1901 19.3944
R18585 vdd.n2318 vdd.n2317 19.3944
R18586 vdd.n2100 vdd.n1905 19.3944
R18587 vdd.n2100 vdd.n1907 19.3944
R18588 vdd.n1910 vdd.n1907 19.3944
R18589 vdd.n2093 vdd.n1910 19.3944
R18590 vdd.n2093 vdd.n2092 19.3944
R18591 vdd.n2092 vdd.n2091 19.3944
R18592 vdd.n2091 vdd.n1916 19.3944
R18593 vdd.n2086 vdd.n1916 19.3944
R18594 vdd.n2086 vdd.n2085 19.3944
R18595 vdd.n2085 vdd.n2084 19.3944
R18596 vdd.n2084 vdd.n1923 19.3944
R18597 vdd.n2079 vdd.n1923 19.3944
R18598 vdd.n2079 vdd.n2078 19.3944
R18599 vdd.n1425 vdd.n1190 19.3944
R18600 vdd.n1425 vdd.n1181 19.3944
R18601 vdd.n1438 vdd.n1181 19.3944
R18602 vdd.n1438 vdd.n1179 19.3944
R18603 vdd.n1442 vdd.n1179 19.3944
R18604 vdd.n1442 vdd.n1170 19.3944
R18605 vdd.n1455 vdd.n1170 19.3944
R18606 vdd.n1455 vdd.n1168 19.3944
R18607 vdd.n1459 vdd.n1168 19.3944
R18608 vdd.n1459 vdd.n1159 19.3944
R18609 vdd.n1471 vdd.n1159 19.3944
R18610 vdd.n1471 vdd.n1157 19.3944
R18611 vdd.n1475 vdd.n1157 19.3944
R18612 vdd.n1475 vdd.n1147 19.3944
R18613 vdd.n1488 vdd.n1147 19.3944
R18614 vdd.n1488 vdd.n1145 19.3944
R18615 vdd.n1492 vdd.n1145 19.3944
R18616 vdd.n1492 vdd.n1136 19.3944
R18617 vdd.n1504 vdd.n1136 19.3944
R18618 vdd.n1504 vdd.n1134 19.3944
R18619 vdd.n1815 vdd.n1134 19.3944
R18620 vdd.n1815 vdd.n1124 19.3944
R18621 vdd.n1828 vdd.n1124 19.3944
R18622 vdd.n1828 vdd.n1122 19.3944
R18623 vdd.n1832 vdd.n1122 19.3944
R18624 vdd.n1832 vdd.n1113 19.3944
R18625 vdd.n1845 vdd.n1113 19.3944
R18626 vdd.n1845 vdd.n1111 19.3944
R18627 vdd.n1849 vdd.n1111 19.3944
R18628 vdd.n1849 vdd.n1102 19.3944
R18629 vdd.n1861 vdd.n1102 19.3944
R18630 vdd.n1861 vdd.n1100 19.3944
R18631 vdd.n1865 vdd.n1100 19.3944
R18632 vdd.n1865 vdd.n1090 19.3944
R18633 vdd.n1878 vdd.n1090 19.3944
R18634 vdd.n1878 vdd.n1088 19.3944
R18635 vdd.n1882 vdd.n1088 19.3944
R18636 vdd.n1882 vdd.n1078 19.3944
R18637 vdd.n1897 vdd.n1078 19.3944
R18638 vdd.n1897 vdd.n1076 19.3944
R18639 vdd.n2327 vdd.n1076 19.3944
R18640 vdd.n3229 vdd.n686 19.3944
R18641 vdd.n3229 vdd.n676 19.3944
R18642 vdd.n3241 vdd.n676 19.3944
R18643 vdd.n3241 vdd.n674 19.3944
R18644 vdd.n3245 vdd.n674 19.3944
R18645 vdd.n3245 vdd.n666 19.3944
R18646 vdd.n3258 vdd.n666 19.3944
R18647 vdd.n3258 vdd.n664 19.3944
R18648 vdd.n3262 vdd.n664 19.3944
R18649 vdd.n3262 vdd.n653 19.3944
R18650 vdd.n3274 vdd.n653 19.3944
R18651 vdd.n3274 vdd.n651 19.3944
R18652 vdd.n3278 vdd.n651 19.3944
R18653 vdd.n3278 vdd.n642 19.3944
R18654 vdd.n3291 vdd.n642 19.3944
R18655 vdd.n3291 vdd.n640 19.3944
R18656 vdd.n3298 vdd.n640 19.3944
R18657 vdd.n3298 vdd.n3297 19.3944
R18658 vdd.n3297 vdd.n631 19.3944
R18659 vdd.n3311 vdd.n631 19.3944
R18660 vdd.n3312 vdd.n3311 19.3944
R18661 vdd.n3312 vdd.n629 19.3944
R18662 vdd.n3316 vdd.n629 19.3944
R18663 vdd.n3318 vdd.n3316 19.3944
R18664 vdd.n3319 vdd.n3318 19.3944
R18665 vdd.n3319 vdd.n627 19.3944
R18666 vdd.n3323 vdd.n627 19.3944
R18667 vdd.n3325 vdd.n3323 19.3944
R18668 vdd.n3326 vdd.n3325 19.3944
R18669 vdd.n3326 vdd.n625 19.3944
R18670 vdd.n3330 vdd.n625 19.3944
R18671 vdd.n3333 vdd.n3330 19.3944
R18672 vdd.n3334 vdd.n3333 19.3944
R18673 vdd.n3334 vdd.n623 19.3944
R18674 vdd.n3338 vdd.n623 19.3944
R18675 vdd.n3340 vdd.n3338 19.3944
R18676 vdd.n3341 vdd.n3340 19.3944
R18677 vdd.n3341 vdd.n621 19.3944
R18678 vdd.n3345 vdd.n621 19.3944
R18679 vdd.n3347 vdd.n3345 19.3944
R18680 vdd.n3348 vdd.n3347 19.3944
R18681 vdd.n569 vdd.n438 19.3944
R18682 vdd.n575 vdd.n438 19.3944
R18683 vdd.n576 vdd.n575 19.3944
R18684 vdd.n579 vdd.n576 19.3944
R18685 vdd.n579 vdd.n436 19.3944
R18686 vdd.n585 vdd.n436 19.3944
R18687 vdd.n586 vdd.n585 19.3944
R18688 vdd.n589 vdd.n586 19.3944
R18689 vdd.n589 vdd.n434 19.3944
R18690 vdd.n595 vdd.n434 19.3944
R18691 vdd.n596 vdd.n595 19.3944
R18692 vdd.n599 vdd.n596 19.3944
R18693 vdd.n599 vdd.n432 19.3944
R18694 vdd.n605 vdd.n432 19.3944
R18695 vdd.n606 vdd.n605 19.3944
R18696 vdd.n609 vdd.n606 19.3944
R18697 vdd.n609 vdd.n430 19.3944
R18698 vdd.n615 vdd.n430 19.3944
R18699 vdd.n617 vdd.n615 19.3944
R18700 vdd.n618 vdd.n617 19.3944
R18701 vdd.n516 vdd.n515 19.3944
R18702 vdd.n519 vdd.n516 19.3944
R18703 vdd.n519 vdd.n450 19.3944
R18704 vdd.n525 vdd.n450 19.3944
R18705 vdd.n526 vdd.n525 19.3944
R18706 vdd.n529 vdd.n526 19.3944
R18707 vdd.n529 vdd.n448 19.3944
R18708 vdd.n535 vdd.n448 19.3944
R18709 vdd.n536 vdd.n535 19.3944
R18710 vdd.n539 vdd.n536 19.3944
R18711 vdd.n539 vdd.n446 19.3944
R18712 vdd.n545 vdd.n446 19.3944
R18713 vdd.n546 vdd.n545 19.3944
R18714 vdd.n549 vdd.n546 19.3944
R18715 vdd.n549 vdd.n444 19.3944
R18716 vdd.n555 vdd.n444 19.3944
R18717 vdd.n556 vdd.n555 19.3944
R18718 vdd.n559 vdd.n556 19.3944
R18719 vdd.n559 vdd.n442 19.3944
R18720 vdd.n565 vdd.n442 19.3944
R18721 vdd.n466 vdd.n465 19.3944
R18722 vdd.n469 vdd.n466 19.3944
R18723 vdd.n469 vdd.n462 19.3944
R18724 vdd.n475 vdd.n462 19.3944
R18725 vdd.n476 vdd.n475 19.3944
R18726 vdd.n479 vdd.n476 19.3944
R18727 vdd.n479 vdd.n460 19.3944
R18728 vdd.n485 vdd.n460 19.3944
R18729 vdd.n486 vdd.n485 19.3944
R18730 vdd.n489 vdd.n486 19.3944
R18731 vdd.n489 vdd.n458 19.3944
R18732 vdd.n495 vdd.n458 19.3944
R18733 vdd.n496 vdd.n495 19.3944
R18734 vdd.n499 vdd.n496 19.3944
R18735 vdd.n499 vdd.n456 19.3944
R18736 vdd.n505 vdd.n456 19.3944
R18737 vdd.n506 vdd.n505 19.3944
R18738 vdd.n509 vdd.n506 19.3944
R18739 vdd.n3233 vdd.n683 19.3944
R18740 vdd.n3233 vdd.n681 19.3944
R18741 vdd.n3237 vdd.n681 19.3944
R18742 vdd.n3237 vdd.n671 19.3944
R18743 vdd.n3250 vdd.n671 19.3944
R18744 vdd.n3250 vdd.n669 19.3944
R18745 vdd.n3254 vdd.n669 19.3944
R18746 vdd.n3254 vdd.n660 19.3944
R18747 vdd.n3266 vdd.n660 19.3944
R18748 vdd.n3266 vdd.n658 19.3944
R18749 vdd.n3270 vdd.n658 19.3944
R18750 vdd.n3270 vdd.n648 19.3944
R18751 vdd.n3283 vdd.n648 19.3944
R18752 vdd.n3283 vdd.n646 19.3944
R18753 vdd.n3287 vdd.n646 19.3944
R18754 vdd.n3287 vdd.n637 19.3944
R18755 vdd.n3302 vdd.n637 19.3944
R18756 vdd.n3302 vdd.n635 19.3944
R18757 vdd.n3306 vdd.n635 19.3944
R18758 vdd.n3306 vdd.n336 19.3944
R18759 vdd.n3397 vdd.n336 19.3944
R18760 vdd.n3397 vdd.n337 19.3944
R18761 vdd.n3391 vdd.n337 19.3944
R18762 vdd.n3391 vdd.n3390 19.3944
R18763 vdd.n3390 vdd.n3389 19.3944
R18764 vdd.n3389 vdd.n349 19.3944
R18765 vdd.n3383 vdd.n349 19.3944
R18766 vdd.n3383 vdd.n3382 19.3944
R18767 vdd.n3382 vdd.n3381 19.3944
R18768 vdd.n3381 vdd.n359 19.3944
R18769 vdd.n3375 vdd.n359 19.3944
R18770 vdd.n3375 vdd.n3374 19.3944
R18771 vdd.n3374 vdd.n3373 19.3944
R18772 vdd.n3373 vdd.n370 19.3944
R18773 vdd.n3367 vdd.n370 19.3944
R18774 vdd.n3367 vdd.n3366 19.3944
R18775 vdd.n3366 vdd.n3365 19.3944
R18776 vdd.n3365 vdd.n381 19.3944
R18777 vdd.n3359 vdd.n381 19.3944
R18778 vdd.n3359 vdd.n3358 19.3944
R18779 vdd.n3358 vdd.n3357 19.3944
R18780 vdd.n3180 vdd.n747 19.3944
R18781 vdd.n3180 vdd.n3177 19.3944
R18782 vdd.n3177 vdd.n3174 19.3944
R18783 vdd.n3174 vdd.n3173 19.3944
R18784 vdd.n3173 vdd.n3170 19.3944
R18785 vdd.n3170 vdd.n3169 19.3944
R18786 vdd.n3169 vdd.n3166 19.3944
R18787 vdd.n3166 vdd.n3165 19.3944
R18788 vdd.n3165 vdd.n3162 19.3944
R18789 vdd.n3162 vdd.n3161 19.3944
R18790 vdd.n3161 vdd.n3158 19.3944
R18791 vdd.n3158 vdd.n3157 19.3944
R18792 vdd.n3157 vdd.n3154 19.3944
R18793 vdd.n3154 vdd.n3153 19.3944
R18794 vdd.n3153 vdd.n3150 19.3944
R18795 vdd.n3150 vdd.n3149 19.3944
R18796 vdd.n3149 vdd.n3146 19.3944
R18797 vdd.n3146 vdd.n3145 19.3944
R18798 vdd.n3145 vdd.n3142 19.3944
R18799 vdd.n3142 vdd.n3141 19.3944
R18800 vdd.n3220 vdd.n3219 19.3944
R18801 vdd.n3219 vdd.n3218 19.3944
R18802 vdd.n732 vdd.n729 19.3944
R18803 vdd.n3214 vdd.n3213 19.3944
R18804 vdd.n3213 vdd.n3210 19.3944
R18805 vdd.n3210 vdd.n3209 19.3944
R18806 vdd.n3209 vdd.n3206 19.3944
R18807 vdd.n3206 vdd.n3205 19.3944
R18808 vdd.n3205 vdd.n3202 19.3944
R18809 vdd.n3202 vdd.n3201 19.3944
R18810 vdd.n3201 vdd.n3198 19.3944
R18811 vdd.n3198 vdd.n3197 19.3944
R18812 vdd.n3197 vdd.n3194 19.3944
R18813 vdd.n3194 vdd.n3193 19.3944
R18814 vdd.n3193 vdd.n3190 19.3944
R18815 vdd.n3190 vdd.n3189 19.3944
R18816 vdd.n3134 vdd.n767 19.3944
R18817 vdd.n3134 vdd.n3131 19.3944
R18818 vdd.n3131 vdd.n3128 19.3944
R18819 vdd.n3128 vdd.n3127 19.3944
R18820 vdd.n3127 vdd.n3124 19.3944
R18821 vdd.n3124 vdd.n3123 19.3944
R18822 vdd.n3123 vdd.n3120 19.3944
R18823 vdd.n3120 vdd.n3119 19.3944
R18824 vdd.n3119 vdd.n3116 19.3944
R18825 vdd.n3116 vdd.n3115 19.3944
R18826 vdd.n3115 vdd.n3112 19.3944
R18827 vdd.n3112 vdd.n3111 19.3944
R18828 vdd.n3111 vdd.n3108 19.3944
R18829 vdd.n3108 vdd.n3107 19.3944
R18830 vdd.n3107 vdd.n3104 19.3944
R18831 vdd.n3104 vdd.n3103 19.3944
R18832 vdd.n3100 vdd.n3099 19.3944
R18833 vdd.n3096 vdd.n3095 19.3944
R18834 vdd.n1357 vdd.n1353 19.0066
R18835 vdd.n2038 vdd.n1969 19.0066
R18836 vdd.n569 vdd.n566 19.0066
R18837 vdd.n3138 vdd.n767 19.0066
R18838 vdd.n2178 vdd.n2177 16.0975
R18839 vdd.n966 vdd.n965 16.0975
R18840 vdd.n1318 vdd.n1317 16.0975
R18841 vdd.n1356 vdd.n1355 16.0975
R18842 vdd.n1252 vdd.n1251 16.0975
R18843 vdd.n2334 vdd.n2333 16.0975
R18844 vdd.n1971 vdd.n1970 16.0975
R18845 vdd.n1931 vdd.n1930 16.0975
R18846 vdd.n2152 vdd.n2151 16.0975
R18847 vdd.n958 vdd.n957 16.0975
R18848 vdd.n2643 vdd.n2642 16.0975
R18849 vdd.n427 vdd.n426 16.0975
R18850 vdd.n441 vdd.n440 16.0975
R18851 vdd.n453 vdd.n452 16.0975
R18852 vdd.n769 vdd.n768 16.0975
R18853 vdd.n3185 vdd.n3184 16.0975
R18854 vdd.n833 vdd.n832 16.0975
R18855 vdd.n2640 vdd.n2639 16.0975
R18856 vdd.n689 vdd.n688 16.0975
R18857 vdd.n800 vdd.n799 16.0975
R18858 vdd.t286 vdd.n2604 15.4182
R18859 vdd.n2857 vdd.t111 15.4182
R18860 vdd.n28 vdd.n27 14.5238
R18861 vdd.n2375 vdd.n1049 14.5112
R18862 vdd.n3059 vdd.n692 14.5112
R18863 vdd.n328 vdd.n293 13.1884
R18864 vdd.n269 vdd.n234 13.1884
R18865 vdd.n226 vdd.n191 13.1884
R18866 vdd.n167 vdd.n132 13.1884
R18867 vdd.n125 vdd.n90 13.1884
R18868 vdd.n66 vdd.n31 13.1884
R18869 vdd.n1747 vdd.n1712 13.1884
R18870 vdd.n1806 vdd.n1771 13.1884
R18871 vdd.n1645 vdd.n1610 13.1884
R18872 vdd.n1704 vdd.n1669 13.1884
R18873 vdd.n1544 vdd.n1509 13.1884
R18874 vdd.n1603 vdd.n1568 13.1884
R18875 vdd.n1388 vdd.n1253 12.9944
R18876 vdd.n1392 vdd.n1253 12.9944
R18877 vdd.n2077 vdd.n1929 12.9944
R18878 vdd.n2078 vdd.n2077 12.9944
R18879 vdd.n515 vdd.n454 12.9944
R18880 vdd.n509 vdd.n454 12.9944
R18881 vdd.n3186 vdd.n747 12.9944
R18882 vdd.n3189 vdd.n3186 12.9944
R18883 vdd.n329 vdd.n291 12.8005
R18884 vdd.n324 vdd.n295 12.8005
R18885 vdd.n270 vdd.n232 12.8005
R18886 vdd.n265 vdd.n236 12.8005
R18887 vdd.n227 vdd.n189 12.8005
R18888 vdd.n222 vdd.n193 12.8005
R18889 vdd.n168 vdd.n130 12.8005
R18890 vdd.n163 vdd.n134 12.8005
R18891 vdd.n126 vdd.n88 12.8005
R18892 vdd.n121 vdd.n92 12.8005
R18893 vdd.n67 vdd.n29 12.8005
R18894 vdd.n62 vdd.n33 12.8005
R18895 vdd.n1748 vdd.n1710 12.8005
R18896 vdd.n1743 vdd.n1714 12.8005
R18897 vdd.n1807 vdd.n1769 12.8005
R18898 vdd.n1802 vdd.n1773 12.8005
R18899 vdd.n1646 vdd.n1608 12.8005
R18900 vdd.n1641 vdd.n1612 12.8005
R18901 vdd.n1705 vdd.n1667 12.8005
R18902 vdd.n1700 vdd.n1671 12.8005
R18903 vdd.n1545 vdd.n1507 12.8005
R18904 vdd.n1540 vdd.n1511 12.8005
R18905 vdd.n1604 vdd.n1566 12.8005
R18906 vdd.n1599 vdd.n1570 12.8005
R18907 vdd.n323 vdd.n296 12.0247
R18908 vdd.n264 vdd.n237 12.0247
R18909 vdd.n221 vdd.n194 12.0247
R18910 vdd.n162 vdd.n135 12.0247
R18911 vdd.n120 vdd.n93 12.0247
R18912 vdd.n61 vdd.n34 12.0247
R18913 vdd.n1742 vdd.n1715 12.0247
R18914 vdd.n1801 vdd.n1774 12.0247
R18915 vdd.n1640 vdd.n1613 12.0247
R18916 vdd.n1699 vdd.n1672 12.0247
R18917 vdd.n1539 vdd.n1512 12.0247
R18918 vdd.n1598 vdd.n1571 12.0247
R18919 vdd.n1427 vdd.n1183 11.337
R18920 vdd.n1436 vdd.n1183 11.337
R18921 vdd.n1436 vdd.n1435 11.337
R18922 vdd.n1444 vdd.n1177 11.337
R18923 vdd.n1453 vdd.n1452 11.337
R18924 vdd.n1469 vdd.n1161 11.337
R18925 vdd.n1477 vdd.n1154 11.337
R18926 vdd.n1486 vdd.n1485 11.337
R18927 vdd.n1494 vdd.n1143 11.337
R18928 vdd.n1817 vdd.n1132 11.337
R18929 vdd.n1826 vdd.n1126 11.337
R18930 vdd.n1834 vdd.n1120 11.337
R18931 vdd.n1843 vdd.n1842 11.337
R18932 vdd.n1859 vdd.n1104 11.337
R18933 vdd.n1867 vdd.n1097 11.337
R18934 vdd.n1876 vdd.n1875 11.337
R18935 vdd.n1884 vdd.n1080 11.337
R18936 vdd.n1895 vdd.n1080 11.337
R18937 vdd.n1895 vdd.n1894 11.337
R18938 vdd.n3231 vdd.n678 11.337
R18939 vdd.n3239 vdd.n678 11.337
R18940 vdd.n3239 vdd.n679 11.337
R18941 vdd.n3248 vdd.n3247 11.337
R18942 vdd.n3264 vdd.n662 11.337
R18943 vdd.n3272 vdd.n655 11.337
R18944 vdd.n3281 vdd.n3280 11.337
R18945 vdd.n3289 vdd.n644 11.337
R18946 vdd.n3308 vdd.n633 11.337
R18947 vdd.n3395 vdd.n340 11.337
R18948 vdd.n3393 vdd.n344 11.337
R18949 vdd.n3387 vdd.n3386 11.337
R18950 vdd.n3379 vdd.n361 11.337
R18951 vdd.n3378 vdd.n3377 11.337
R18952 vdd.n3371 vdd.n3370 11.337
R18953 vdd.n3369 vdd.n375 11.337
R18954 vdd.n3363 vdd.n3362 11.337
R18955 vdd.n3362 vdd.n3361 11.337
R18956 vdd.n3361 vdd.n386 11.337
R18957 vdd.n320 vdd.n319 11.249
R18958 vdd.n261 vdd.n260 11.249
R18959 vdd.n218 vdd.n217 11.249
R18960 vdd.n159 vdd.n158 11.249
R18961 vdd.n117 vdd.n116 11.249
R18962 vdd.n58 vdd.n57 11.249
R18963 vdd.n1739 vdd.n1738 11.249
R18964 vdd.n1798 vdd.n1797 11.249
R18965 vdd.n1637 vdd.n1636 11.249
R18966 vdd.n1696 vdd.n1695 11.249
R18967 vdd.n1536 vdd.n1535 11.249
R18968 vdd.n1595 vdd.n1594 11.249
R18969 vdd.n1225 vdd.t50 11.2237
R18970 vdd.n3355 vdd.t57 11.2237
R18971 vdd.n2532 vdd.t12 11.1103
R18972 vdd.n2864 vdd.t290 11.1103
R18973 vdd.t141 vdd.n1098 10.7702
R18974 vdd.n3256 vdd.t206 10.7702
R18975 vdd.n305 vdd.n304 10.7238
R18976 vdd.n246 vdd.n245 10.7238
R18977 vdd.n203 vdd.n202 10.7238
R18978 vdd.n144 vdd.n143 10.7238
R18979 vdd.n102 vdd.n101 10.7238
R18980 vdd.n43 vdd.n42 10.7238
R18981 vdd.n1724 vdd.n1723 10.7238
R18982 vdd.n1783 vdd.n1782 10.7238
R18983 vdd.n1622 vdd.n1621 10.7238
R18984 vdd.n1681 vdd.n1680 10.7238
R18985 vdd.n1521 vdd.n1520 10.7238
R18986 vdd.n1580 vdd.n1579 10.7238
R18987 vdd.n2378 vdd.n2377 10.6151
R18988 vdd.n2379 vdd.n2378 10.6151
R18989 vdd.n2379 vdd.n1035 10.6151
R18990 vdd.n2389 vdd.n1035 10.6151
R18991 vdd.n2390 vdd.n2389 10.6151
R18992 vdd.n2391 vdd.n2390 10.6151
R18993 vdd.n2391 vdd.n1022 10.6151
R18994 vdd.n2402 vdd.n1022 10.6151
R18995 vdd.n2403 vdd.n2402 10.6151
R18996 vdd.n2404 vdd.n2403 10.6151
R18997 vdd.n2404 vdd.n1010 10.6151
R18998 vdd.n2414 vdd.n1010 10.6151
R18999 vdd.n2415 vdd.n2414 10.6151
R19000 vdd.n2416 vdd.n2415 10.6151
R19001 vdd.n2416 vdd.n998 10.6151
R19002 vdd.n2426 vdd.n998 10.6151
R19003 vdd.n2427 vdd.n2426 10.6151
R19004 vdd.n2428 vdd.n2427 10.6151
R19005 vdd.n2428 vdd.n987 10.6151
R19006 vdd.n2438 vdd.n987 10.6151
R19007 vdd.n2439 vdd.n2438 10.6151
R19008 vdd.n2440 vdd.n2439 10.6151
R19009 vdd.n2440 vdd.n974 10.6151
R19010 vdd.n2452 vdd.n974 10.6151
R19011 vdd.n2453 vdd.n2452 10.6151
R19012 vdd.n2455 vdd.n2453 10.6151
R19013 vdd.n2455 vdd.n2454 10.6151
R19014 vdd.n2454 vdd.n956 10.6151
R19015 vdd.n2602 vdd.n2601 10.6151
R19016 vdd.n2601 vdd.n2600 10.6151
R19017 vdd.n2600 vdd.n2597 10.6151
R19018 vdd.n2597 vdd.n2596 10.6151
R19019 vdd.n2596 vdd.n2593 10.6151
R19020 vdd.n2593 vdd.n2592 10.6151
R19021 vdd.n2592 vdd.n2589 10.6151
R19022 vdd.n2589 vdd.n2588 10.6151
R19023 vdd.n2588 vdd.n2585 10.6151
R19024 vdd.n2585 vdd.n2584 10.6151
R19025 vdd.n2584 vdd.n2581 10.6151
R19026 vdd.n2581 vdd.n2580 10.6151
R19027 vdd.n2580 vdd.n2577 10.6151
R19028 vdd.n2577 vdd.n2576 10.6151
R19029 vdd.n2576 vdd.n2573 10.6151
R19030 vdd.n2573 vdd.n2572 10.6151
R19031 vdd.n2572 vdd.n2569 10.6151
R19032 vdd.n2569 vdd.n2568 10.6151
R19033 vdd.n2568 vdd.n2565 10.6151
R19034 vdd.n2565 vdd.n2564 10.6151
R19035 vdd.n2564 vdd.n2561 10.6151
R19036 vdd.n2561 vdd.n2560 10.6151
R19037 vdd.n2560 vdd.n2557 10.6151
R19038 vdd.n2557 vdd.n2556 10.6151
R19039 vdd.n2556 vdd.n2553 10.6151
R19040 vdd.n2553 vdd.n2552 10.6151
R19041 vdd.n2552 vdd.n2549 10.6151
R19042 vdd.n2549 vdd.n2548 10.6151
R19043 vdd.n2548 vdd.n2545 10.6151
R19044 vdd.n2545 vdd.n2544 10.6151
R19045 vdd.n2544 vdd.n2541 10.6151
R19046 vdd.n2539 vdd.n2536 10.6151
R19047 vdd.n2536 vdd.n2535 10.6151
R19048 vdd.n2278 vdd.n2277 10.6151
R19049 vdd.n2277 vdd.n2275 10.6151
R19050 vdd.n2275 vdd.n2274 10.6151
R19051 vdd.n2274 vdd.n2272 10.6151
R19052 vdd.n2272 vdd.n2271 10.6151
R19053 vdd.n2271 vdd.n2269 10.6151
R19054 vdd.n2269 vdd.n2268 10.6151
R19055 vdd.n2268 vdd.n2266 10.6151
R19056 vdd.n2266 vdd.n2265 10.6151
R19057 vdd.n2265 vdd.n2263 10.6151
R19058 vdd.n2263 vdd.n2262 10.6151
R19059 vdd.n2262 vdd.n2260 10.6151
R19060 vdd.n2260 vdd.n2259 10.6151
R19061 vdd.n2259 vdd.n2174 10.6151
R19062 vdd.n2174 vdd.n2173 10.6151
R19063 vdd.n2173 vdd.n2171 10.6151
R19064 vdd.n2171 vdd.n2170 10.6151
R19065 vdd.n2170 vdd.n2168 10.6151
R19066 vdd.n2168 vdd.n2167 10.6151
R19067 vdd.n2167 vdd.n2165 10.6151
R19068 vdd.n2165 vdd.n2164 10.6151
R19069 vdd.n2164 vdd.n2162 10.6151
R19070 vdd.n2162 vdd.n2161 10.6151
R19071 vdd.n2161 vdd.n2159 10.6151
R19072 vdd.n2159 vdd.n2158 10.6151
R19073 vdd.n2158 vdd.n2155 10.6151
R19074 vdd.n2155 vdd.n2154 10.6151
R19075 vdd.n2154 vdd.n959 10.6151
R19076 vdd.n2112 vdd.n1047 10.6151
R19077 vdd.n2113 vdd.n2112 10.6151
R19078 vdd.n2114 vdd.n2113 10.6151
R19079 vdd.n2114 vdd.n2108 10.6151
R19080 vdd.n2120 vdd.n2108 10.6151
R19081 vdd.n2121 vdd.n2120 10.6151
R19082 vdd.n2122 vdd.n2121 10.6151
R19083 vdd.n2122 vdd.n2106 10.6151
R19084 vdd.n2128 vdd.n2106 10.6151
R19085 vdd.n2129 vdd.n2128 10.6151
R19086 vdd.n2130 vdd.n2129 10.6151
R19087 vdd.n2130 vdd.n2104 10.6151
R19088 vdd.n2136 vdd.n2104 10.6151
R19089 vdd.n2137 vdd.n2136 10.6151
R19090 vdd.n2138 vdd.n2137 10.6151
R19091 vdd.n2138 vdd.n2102 10.6151
R19092 vdd.n2314 vdd.n2102 10.6151
R19093 vdd.n2314 vdd.n2313 10.6151
R19094 vdd.n2313 vdd.n2143 10.6151
R19095 vdd.n2307 vdd.n2143 10.6151
R19096 vdd.n2307 vdd.n2306 10.6151
R19097 vdd.n2306 vdd.n2305 10.6151
R19098 vdd.n2305 vdd.n2145 10.6151
R19099 vdd.n2299 vdd.n2145 10.6151
R19100 vdd.n2299 vdd.n2298 10.6151
R19101 vdd.n2298 vdd.n2297 10.6151
R19102 vdd.n2297 vdd.n2147 10.6151
R19103 vdd.n2291 vdd.n2147 10.6151
R19104 vdd.n2291 vdd.n2290 10.6151
R19105 vdd.n2290 vdd.n2289 10.6151
R19106 vdd.n2289 vdd.n2149 10.6151
R19107 vdd.n2283 vdd.n2282 10.6151
R19108 vdd.n2282 vdd.n2281 10.6151
R19109 vdd.n2787 vdd.n2786 10.6151
R19110 vdd.n2786 vdd.n2784 10.6151
R19111 vdd.n2784 vdd.n2783 10.6151
R19112 vdd.n2783 vdd.n2641 10.6151
R19113 vdd.n2730 vdd.n2641 10.6151
R19114 vdd.n2731 vdd.n2730 10.6151
R19115 vdd.n2733 vdd.n2731 10.6151
R19116 vdd.n2734 vdd.n2733 10.6151
R19117 vdd.n2736 vdd.n2734 10.6151
R19118 vdd.n2737 vdd.n2736 10.6151
R19119 vdd.n2739 vdd.n2737 10.6151
R19120 vdd.n2740 vdd.n2739 10.6151
R19121 vdd.n2742 vdd.n2740 10.6151
R19122 vdd.n2743 vdd.n2742 10.6151
R19123 vdd.n2758 vdd.n2743 10.6151
R19124 vdd.n2758 vdd.n2757 10.6151
R19125 vdd.n2757 vdd.n2756 10.6151
R19126 vdd.n2756 vdd.n2754 10.6151
R19127 vdd.n2754 vdd.n2753 10.6151
R19128 vdd.n2753 vdd.n2751 10.6151
R19129 vdd.n2751 vdd.n2750 10.6151
R19130 vdd.n2750 vdd.n2748 10.6151
R19131 vdd.n2748 vdd.n2747 10.6151
R19132 vdd.n2747 vdd.n2745 10.6151
R19133 vdd.n2745 vdd.n2744 10.6151
R19134 vdd.n2744 vdd.n836 10.6151
R19135 vdd.n2992 vdd.n836 10.6151
R19136 vdd.n2993 vdd.n2992 10.6151
R19137 vdd.n2854 vdd.n912 10.6151
R19138 vdd.n2854 vdd.n2853 10.6151
R19139 vdd.n2853 vdd.n2852 10.6151
R19140 vdd.n2852 vdd.n2850 10.6151
R19141 vdd.n2850 vdd.n2847 10.6151
R19142 vdd.n2847 vdd.n2846 10.6151
R19143 vdd.n2846 vdd.n2843 10.6151
R19144 vdd.n2843 vdd.n2842 10.6151
R19145 vdd.n2842 vdd.n2839 10.6151
R19146 vdd.n2839 vdd.n2838 10.6151
R19147 vdd.n2838 vdd.n2835 10.6151
R19148 vdd.n2835 vdd.n2834 10.6151
R19149 vdd.n2834 vdd.n2831 10.6151
R19150 vdd.n2831 vdd.n2830 10.6151
R19151 vdd.n2830 vdd.n2827 10.6151
R19152 vdd.n2827 vdd.n2826 10.6151
R19153 vdd.n2826 vdd.n2823 10.6151
R19154 vdd.n2823 vdd.n2822 10.6151
R19155 vdd.n2822 vdd.n2819 10.6151
R19156 vdd.n2819 vdd.n2818 10.6151
R19157 vdd.n2818 vdd.n2815 10.6151
R19158 vdd.n2815 vdd.n2814 10.6151
R19159 vdd.n2814 vdd.n2811 10.6151
R19160 vdd.n2811 vdd.n2810 10.6151
R19161 vdd.n2810 vdd.n2807 10.6151
R19162 vdd.n2807 vdd.n2806 10.6151
R19163 vdd.n2806 vdd.n2803 10.6151
R19164 vdd.n2803 vdd.n2802 10.6151
R19165 vdd.n2802 vdd.n2799 10.6151
R19166 vdd.n2799 vdd.n2798 10.6151
R19167 vdd.n2798 vdd.n2795 10.6151
R19168 vdd.n2793 vdd.n2790 10.6151
R19169 vdd.n2790 vdd.n2789 10.6151
R19170 vdd.n2867 vdd.n2866 10.6151
R19171 vdd.n2868 vdd.n2867 10.6151
R19172 vdd.n2868 vdd.n902 10.6151
R19173 vdd.n2878 vdd.n902 10.6151
R19174 vdd.n2879 vdd.n2878 10.6151
R19175 vdd.n2880 vdd.n2879 10.6151
R19176 vdd.n2880 vdd.n889 10.6151
R19177 vdd.n2890 vdd.n889 10.6151
R19178 vdd.n2891 vdd.n2890 10.6151
R19179 vdd.n2892 vdd.n2891 10.6151
R19180 vdd.n2892 vdd.n878 10.6151
R19181 vdd.n2902 vdd.n878 10.6151
R19182 vdd.n2903 vdd.n2902 10.6151
R19183 vdd.n2904 vdd.n2903 10.6151
R19184 vdd.n2904 vdd.n866 10.6151
R19185 vdd.n2914 vdd.n866 10.6151
R19186 vdd.n2915 vdd.n2914 10.6151
R19187 vdd.n2916 vdd.n2915 10.6151
R19188 vdd.n2916 vdd.n855 10.6151
R19189 vdd.n2928 vdd.n855 10.6151
R19190 vdd.n2929 vdd.n2928 10.6151
R19191 vdd.n2930 vdd.n2929 10.6151
R19192 vdd.n2930 vdd.n841 10.6151
R19193 vdd.n2985 vdd.n841 10.6151
R19194 vdd.n2986 vdd.n2985 10.6151
R19195 vdd.n2987 vdd.n2986 10.6151
R19196 vdd.n2987 vdd.n810 10.6151
R19197 vdd.n3057 vdd.n810 10.6151
R19198 vdd.n3056 vdd.n3055 10.6151
R19199 vdd.n3055 vdd.n811 10.6151
R19200 vdd.n812 vdd.n811 10.6151
R19201 vdd.n3048 vdd.n812 10.6151
R19202 vdd.n3048 vdd.n3047 10.6151
R19203 vdd.n3047 vdd.n3046 10.6151
R19204 vdd.n3046 vdd.n814 10.6151
R19205 vdd.n3041 vdd.n814 10.6151
R19206 vdd.n3041 vdd.n3040 10.6151
R19207 vdd.n3040 vdd.n3039 10.6151
R19208 vdd.n3039 vdd.n817 10.6151
R19209 vdd.n3034 vdd.n817 10.6151
R19210 vdd.n3034 vdd.n3033 10.6151
R19211 vdd.n3033 vdd.n3032 10.6151
R19212 vdd.n3032 vdd.n820 10.6151
R19213 vdd.n3027 vdd.n820 10.6151
R19214 vdd.n3027 vdd.n731 10.6151
R19215 vdd.n3023 vdd.n731 10.6151
R19216 vdd.n3023 vdd.n3022 10.6151
R19217 vdd.n3022 vdd.n3021 10.6151
R19218 vdd.n3021 vdd.n823 10.6151
R19219 vdd.n3016 vdd.n823 10.6151
R19220 vdd.n3016 vdd.n3015 10.6151
R19221 vdd.n3015 vdd.n3014 10.6151
R19222 vdd.n3014 vdd.n826 10.6151
R19223 vdd.n3009 vdd.n826 10.6151
R19224 vdd.n3009 vdd.n3008 10.6151
R19225 vdd.n3008 vdd.n3007 10.6151
R19226 vdd.n3007 vdd.n829 10.6151
R19227 vdd.n3002 vdd.n829 10.6151
R19228 vdd.n3002 vdd.n3001 10.6151
R19229 vdd.n2999 vdd.n834 10.6151
R19230 vdd.n2994 vdd.n834 10.6151
R19231 vdd.n2975 vdd.n2936 10.6151
R19232 vdd.n2970 vdd.n2936 10.6151
R19233 vdd.n2970 vdd.n2969 10.6151
R19234 vdd.n2969 vdd.n2968 10.6151
R19235 vdd.n2968 vdd.n2938 10.6151
R19236 vdd.n2963 vdd.n2938 10.6151
R19237 vdd.n2963 vdd.n2962 10.6151
R19238 vdd.n2962 vdd.n2961 10.6151
R19239 vdd.n2961 vdd.n2941 10.6151
R19240 vdd.n2956 vdd.n2941 10.6151
R19241 vdd.n2956 vdd.n2955 10.6151
R19242 vdd.n2955 vdd.n2954 10.6151
R19243 vdd.n2954 vdd.n2944 10.6151
R19244 vdd.n2949 vdd.n2944 10.6151
R19245 vdd.n2949 vdd.n2948 10.6151
R19246 vdd.n2948 vdd.n785 10.6151
R19247 vdd.n3092 vdd.n785 10.6151
R19248 vdd.n3092 vdd.n786 10.6151
R19249 vdd.n788 vdd.n786 10.6151
R19250 vdd.n3085 vdd.n788 10.6151
R19251 vdd.n3085 vdd.n3084 10.6151
R19252 vdd.n3084 vdd.n3083 10.6151
R19253 vdd.n3083 vdd.n790 10.6151
R19254 vdd.n3078 vdd.n790 10.6151
R19255 vdd.n3078 vdd.n3077 10.6151
R19256 vdd.n3077 vdd.n3076 10.6151
R19257 vdd.n3076 vdd.n793 10.6151
R19258 vdd.n3071 vdd.n793 10.6151
R19259 vdd.n3071 vdd.n3070 10.6151
R19260 vdd.n3070 vdd.n3069 10.6151
R19261 vdd.n3069 vdd.n796 10.6151
R19262 vdd.n3064 vdd.n3063 10.6151
R19263 vdd.n3063 vdd.n3062 10.6151
R19264 vdd.n2710 vdd.n2708 10.6151
R19265 vdd.n2711 vdd.n2710 10.6151
R19266 vdd.n2779 vdd.n2711 10.6151
R19267 vdd.n2779 vdd.n2778 10.6151
R19268 vdd.n2778 vdd.n2777 10.6151
R19269 vdd.n2777 vdd.n2775 10.6151
R19270 vdd.n2775 vdd.n2774 10.6151
R19271 vdd.n2774 vdd.n2772 10.6151
R19272 vdd.n2772 vdd.n2771 10.6151
R19273 vdd.n2771 vdd.n2769 10.6151
R19274 vdd.n2769 vdd.n2768 10.6151
R19275 vdd.n2768 vdd.n2766 10.6151
R19276 vdd.n2766 vdd.n2765 10.6151
R19277 vdd.n2765 vdd.n2763 10.6151
R19278 vdd.n2763 vdd.n2762 10.6151
R19279 vdd.n2762 vdd.n2728 10.6151
R19280 vdd.n2728 vdd.n2727 10.6151
R19281 vdd.n2727 vdd.n2725 10.6151
R19282 vdd.n2725 vdd.n2724 10.6151
R19283 vdd.n2724 vdd.n2722 10.6151
R19284 vdd.n2722 vdd.n2721 10.6151
R19285 vdd.n2721 vdd.n2719 10.6151
R19286 vdd.n2719 vdd.n2718 10.6151
R19287 vdd.n2718 vdd.n2716 10.6151
R19288 vdd.n2716 vdd.n2715 10.6151
R19289 vdd.n2715 vdd.n2713 10.6151
R19290 vdd.n2713 vdd.n2712 10.6151
R19291 vdd.n2712 vdd.n802 10.6151
R19292 vdd.n2861 vdd.n2860 10.6151
R19293 vdd.n2860 vdd.n917 10.6151
R19294 vdd.n2645 vdd.n917 10.6151
R19295 vdd.n2648 vdd.n2645 10.6151
R19296 vdd.n2649 vdd.n2648 10.6151
R19297 vdd.n2652 vdd.n2649 10.6151
R19298 vdd.n2653 vdd.n2652 10.6151
R19299 vdd.n2656 vdd.n2653 10.6151
R19300 vdd.n2657 vdd.n2656 10.6151
R19301 vdd.n2660 vdd.n2657 10.6151
R19302 vdd.n2661 vdd.n2660 10.6151
R19303 vdd.n2664 vdd.n2661 10.6151
R19304 vdd.n2665 vdd.n2664 10.6151
R19305 vdd.n2668 vdd.n2665 10.6151
R19306 vdd.n2669 vdd.n2668 10.6151
R19307 vdd.n2672 vdd.n2669 10.6151
R19308 vdd.n2673 vdd.n2672 10.6151
R19309 vdd.n2676 vdd.n2673 10.6151
R19310 vdd.n2677 vdd.n2676 10.6151
R19311 vdd.n2680 vdd.n2677 10.6151
R19312 vdd.n2681 vdd.n2680 10.6151
R19313 vdd.n2684 vdd.n2681 10.6151
R19314 vdd.n2685 vdd.n2684 10.6151
R19315 vdd.n2688 vdd.n2685 10.6151
R19316 vdd.n2689 vdd.n2688 10.6151
R19317 vdd.n2692 vdd.n2689 10.6151
R19318 vdd.n2693 vdd.n2692 10.6151
R19319 vdd.n2696 vdd.n2693 10.6151
R19320 vdd.n2697 vdd.n2696 10.6151
R19321 vdd.n2700 vdd.n2697 10.6151
R19322 vdd.n2701 vdd.n2700 10.6151
R19323 vdd.n2706 vdd.n2704 10.6151
R19324 vdd.n2707 vdd.n2706 10.6151
R19325 vdd.n2862 vdd.n907 10.6151
R19326 vdd.n2872 vdd.n907 10.6151
R19327 vdd.n2873 vdd.n2872 10.6151
R19328 vdd.n2874 vdd.n2873 10.6151
R19329 vdd.n2874 vdd.n895 10.6151
R19330 vdd.n2884 vdd.n895 10.6151
R19331 vdd.n2885 vdd.n2884 10.6151
R19332 vdd.n2886 vdd.n2885 10.6151
R19333 vdd.n2886 vdd.n884 10.6151
R19334 vdd.n2896 vdd.n884 10.6151
R19335 vdd.n2897 vdd.n2896 10.6151
R19336 vdd.n2898 vdd.n2897 10.6151
R19337 vdd.n2898 vdd.n872 10.6151
R19338 vdd.n2908 vdd.n872 10.6151
R19339 vdd.n2909 vdd.n2908 10.6151
R19340 vdd.n2910 vdd.n2909 10.6151
R19341 vdd.n2910 vdd.n861 10.6151
R19342 vdd.n2920 vdd.n861 10.6151
R19343 vdd.n2921 vdd.n2920 10.6151
R19344 vdd.n2924 vdd.n2921 10.6151
R19345 vdd.n2934 vdd.n849 10.6151
R19346 vdd.n2935 vdd.n2934 10.6151
R19347 vdd.n2981 vdd.n2935 10.6151
R19348 vdd.n2981 vdd.n2980 10.6151
R19349 vdd.n2980 vdd.n2979 10.6151
R19350 vdd.n2979 vdd.n2978 10.6151
R19351 vdd.n2978 vdd.n2976 10.6151
R19352 vdd.n2373 vdd.n1041 10.6151
R19353 vdd.n2383 vdd.n1041 10.6151
R19354 vdd.n2384 vdd.n2383 10.6151
R19355 vdd.n2385 vdd.n2384 10.6151
R19356 vdd.n2385 vdd.n1028 10.6151
R19357 vdd.n2395 vdd.n1028 10.6151
R19358 vdd.n2396 vdd.n2395 10.6151
R19359 vdd.n2398 vdd.n1016 10.6151
R19360 vdd.n2408 vdd.n1016 10.6151
R19361 vdd.n2409 vdd.n2408 10.6151
R19362 vdd.n2410 vdd.n2409 10.6151
R19363 vdd.n2410 vdd.n1004 10.6151
R19364 vdd.n2420 vdd.n1004 10.6151
R19365 vdd.n2421 vdd.n2420 10.6151
R19366 vdd.n2422 vdd.n2421 10.6151
R19367 vdd.n2422 vdd.n993 10.6151
R19368 vdd.n2432 vdd.n993 10.6151
R19369 vdd.n2433 vdd.n2432 10.6151
R19370 vdd.n2434 vdd.n2433 10.6151
R19371 vdd.n2434 vdd.n981 10.6151
R19372 vdd.n2444 vdd.n981 10.6151
R19373 vdd.n2445 vdd.n2444 10.6151
R19374 vdd.n2448 vdd.n2445 10.6151
R19375 vdd.n2448 vdd.n2447 10.6151
R19376 vdd.n2447 vdd.n2446 10.6151
R19377 vdd.n2446 vdd.n964 10.6151
R19378 vdd.n2530 vdd.n964 10.6151
R19379 vdd.n2529 vdd.n2528 10.6151
R19380 vdd.n2528 vdd.n2525 10.6151
R19381 vdd.n2525 vdd.n2524 10.6151
R19382 vdd.n2524 vdd.n2521 10.6151
R19383 vdd.n2521 vdd.n2520 10.6151
R19384 vdd.n2520 vdd.n2517 10.6151
R19385 vdd.n2517 vdd.n2516 10.6151
R19386 vdd.n2516 vdd.n2513 10.6151
R19387 vdd.n2513 vdd.n2512 10.6151
R19388 vdd.n2512 vdd.n2509 10.6151
R19389 vdd.n2509 vdd.n2508 10.6151
R19390 vdd.n2508 vdd.n2505 10.6151
R19391 vdd.n2505 vdd.n2504 10.6151
R19392 vdd.n2504 vdd.n2501 10.6151
R19393 vdd.n2501 vdd.n2500 10.6151
R19394 vdd.n2500 vdd.n2497 10.6151
R19395 vdd.n2497 vdd.n2496 10.6151
R19396 vdd.n2496 vdd.n2493 10.6151
R19397 vdd.n2493 vdd.n2492 10.6151
R19398 vdd.n2492 vdd.n2489 10.6151
R19399 vdd.n2489 vdd.n2488 10.6151
R19400 vdd.n2488 vdd.n2485 10.6151
R19401 vdd.n2485 vdd.n2484 10.6151
R19402 vdd.n2484 vdd.n2481 10.6151
R19403 vdd.n2481 vdd.n2480 10.6151
R19404 vdd.n2480 vdd.n2477 10.6151
R19405 vdd.n2477 vdd.n2476 10.6151
R19406 vdd.n2476 vdd.n2473 10.6151
R19407 vdd.n2473 vdd.n2472 10.6151
R19408 vdd.n2472 vdd.n2469 10.6151
R19409 vdd.n2469 vdd.n2468 10.6151
R19410 vdd.n2465 vdd.n2464 10.6151
R19411 vdd.n2464 vdd.n2462 10.6151
R19412 vdd.n2221 vdd.n2219 10.6151
R19413 vdd.n2222 vdd.n2221 10.6151
R19414 vdd.n2224 vdd.n2222 10.6151
R19415 vdd.n2225 vdd.n2224 10.6151
R19416 vdd.n2227 vdd.n2225 10.6151
R19417 vdd.n2228 vdd.n2227 10.6151
R19418 vdd.n2230 vdd.n2228 10.6151
R19419 vdd.n2231 vdd.n2230 10.6151
R19420 vdd.n2233 vdd.n2231 10.6151
R19421 vdd.n2234 vdd.n2233 10.6151
R19422 vdd.n2236 vdd.n2234 10.6151
R19423 vdd.n2237 vdd.n2236 10.6151
R19424 vdd.n2255 vdd.n2237 10.6151
R19425 vdd.n2255 vdd.n2254 10.6151
R19426 vdd.n2254 vdd.n2253 10.6151
R19427 vdd.n2253 vdd.n2251 10.6151
R19428 vdd.n2251 vdd.n2250 10.6151
R19429 vdd.n2250 vdd.n2248 10.6151
R19430 vdd.n2248 vdd.n2247 10.6151
R19431 vdd.n2247 vdd.n2245 10.6151
R19432 vdd.n2245 vdd.n2244 10.6151
R19433 vdd.n2244 vdd.n2242 10.6151
R19434 vdd.n2242 vdd.n2241 10.6151
R19435 vdd.n2241 vdd.n2239 10.6151
R19436 vdd.n2239 vdd.n2238 10.6151
R19437 vdd.n2238 vdd.n968 10.6151
R19438 vdd.n2460 vdd.n968 10.6151
R19439 vdd.n2461 vdd.n2460 10.6151
R19440 vdd.n2372 vdd.n2371 10.6151
R19441 vdd.n2371 vdd.n1053 10.6151
R19442 vdd.n2365 vdd.n1053 10.6151
R19443 vdd.n2365 vdd.n2364 10.6151
R19444 vdd.n2364 vdd.n2363 10.6151
R19445 vdd.n2363 vdd.n1055 10.6151
R19446 vdd.n2357 vdd.n1055 10.6151
R19447 vdd.n2357 vdd.n2356 10.6151
R19448 vdd.n2356 vdd.n2355 10.6151
R19449 vdd.n2355 vdd.n1057 10.6151
R19450 vdd.n2349 vdd.n1057 10.6151
R19451 vdd.n2349 vdd.n2348 10.6151
R19452 vdd.n2348 vdd.n2347 10.6151
R19453 vdd.n2347 vdd.n1059 10.6151
R19454 vdd.n2341 vdd.n1059 10.6151
R19455 vdd.n2341 vdd.n2340 10.6151
R19456 vdd.n2340 vdd.n2339 10.6151
R19457 vdd.n2339 vdd.n1063 10.6151
R19458 vdd.n2187 vdd.n1063 10.6151
R19459 vdd.n2188 vdd.n2187 10.6151
R19460 vdd.n2188 vdd.n2183 10.6151
R19461 vdd.n2194 vdd.n2183 10.6151
R19462 vdd.n2195 vdd.n2194 10.6151
R19463 vdd.n2196 vdd.n2195 10.6151
R19464 vdd.n2196 vdd.n2181 10.6151
R19465 vdd.n2202 vdd.n2181 10.6151
R19466 vdd.n2203 vdd.n2202 10.6151
R19467 vdd.n2204 vdd.n2203 10.6151
R19468 vdd.n2204 vdd.n2179 10.6151
R19469 vdd.n2210 vdd.n2179 10.6151
R19470 vdd.n2211 vdd.n2210 10.6151
R19471 vdd.n2213 vdd.n2175 10.6151
R19472 vdd.n2218 vdd.n2175 10.6151
R19473 vdd.n1851 vdd.t131 10.5435
R19474 vdd.n656 vdd.t239 10.5435
R19475 vdd.n316 vdd.n298 10.4732
R19476 vdd.n257 vdd.n239 10.4732
R19477 vdd.n214 vdd.n196 10.4732
R19478 vdd.n155 vdd.n137 10.4732
R19479 vdd.n113 vdd.n95 10.4732
R19480 vdd.n54 vdd.n36 10.4732
R19481 vdd.n1735 vdd.n1717 10.4732
R19482 vdd.n1794 vdd.n1776 10.4732
R19483 vdd.n1633 vdd.n1615 10.4732
R19484 vdd.n1692 vdd.n1674 10.4732
R19485 vdd.n1532 vdd.n1514 10.4732
R19486 vdd.n1591 vdd.n1573 10.4732
R19487 vdd.t221 vdd.n1825 10.3167
R19488 vdd.n3300 vdd.t183 10.3167
R19489 vdd.n1502 vdd.t149 10.09
R19490 vdd.n3394 vdd.t147 10.09
R19491 vdd.t217 vdd.n1155 9.86327
R19492 vdd.n3385 vdd.t145 9.86327
R19493 vdd.n315 vdd.n300 9.69747
R19494 vdd.n256 vdd.n241 9.69747
R19495 vdd.n213 vdd.n198 9.69747
R19496 vdd.n154 vdd.n139 9.69747
R19497 vdd.n112 vdd.n97 9.69747
R19498 vdd.n53 vdd.n38 9.69747
R19499 vdd.n1734 vdd.n1719 9.69747
R19500 vdd.n1793 vdd.n1778 9.69747
R19501 vdd.n1632 vdd.n1617 9.69747
R19502 vdd.n1691 vdd.n1676 9.69747
R19503 vdd.n1531 vdd.n1516 9.69747
R19504 vdd.n1590 vdd.n1575 9.69747
R19505 vdd.n2315 vdd.n2314 9.67831
R19506 vdd.n3216 vdd.n731 9.67831
R19507 vdd.n3093 vdd.n3092 9.67831
R19508 vdd.n2339 vdd.n2338 9.67831
R19509 vdd.n1461 vdd.t162 9.63654
R19510 vdd.n3331 vdd.t143 9.63654
R19511 vdd.n331 vdd.n330 9.45567
R19512 vdd.n272 vdd.n271 9.45567
R19513 vdd.n229 vdd.n228 9.45567
R19514 vdd.n170 vdd.n169 9.45567
R19515 vdd.n128 vdd.n127 9.45567
R19516 vdd.n69 vdd.n68 9.45567
R19517 vdd.n1750 vdd.n1749 9.45567
R19518 vdd.n1809 vdd.n1808 9.45567
R19519 vdd.n1648 vdd.n1647 9.45567
R19520 vdd.n1707 vdd.n1706 9.45567
R19521 vdd.n1547 vdd.n1546 9.45567
R19522 vdd.n1606 vdd.n1605 9.45567
R19523 vdd.n1435 vdd.t129 9.40981
R19524 vdd.n3363 vdd.t189 9.40981
R19525 vdd.n2075 vdd.n1929 9.3005
R19526 vdd.n2074 vdd.n2073 9.3005
R19527 vdd.n1935 vdd.n1934 9.3005
R19528 vdd.n2068 vdd.n1939 9.3005
R19529 vdd.n2067 vdd.n1940 9.3005
R19530 vdd.n2066 vdd.n1941 9.3005
R19531 vdd.n1945 vdd.n1942 9.3005
R19532 vdd.n2061 vdd.n1946 9.3005
R19533 vdd.n2060 vdd.n1947 9.3005
R19534 vdd.n2059 vdd.n1948 9.3005
R19535 vdd.n1952 vdd.n1949 9.3005
R19536 vdd.n2054 vdd.n1953 9.3005
R19537 vdd.n2053 vdd.n1954 9.3005
R19538 vdd.n2052 vdd.n1955 9.3005
R19539 vdd.n1959 vdd.n1956 9.3005
R19540 vdd.n2047 vdd.n1960 9.3005
R19541 vdd.n2046 vdd.n1961 9.3005
R19542 vdd.n2045 vdd.n1962 9.3005
R19543 vdd.n1966 vdd.n1963 9.3005
R19544 vdd.n2040 vdd.n1967 9.3005
R19545 vdd.n2039 vdd.n1968 9.3005
R19546 vdd.n2038 vdd.n2037 9.3005
R19547 vdd.n2036 vdd.n1969 9.3005
R19548 vdd.n2035 vdd.n2034 9.3005
R19549 vdd.n1975 vdd.n1974 9.3005
R19550 vdd.n2029 vdd.n1979 9.3005
R19551 vdd.n2028 vdd.n1980 9.3005
R19552 vdd.n2027 vdd.n1981 9.3005
R19553 vdd.n1985 vdd.n1982 9.3005
R19554 vdd.n2022 vdd.n1986 9.3005
R19555 vdd.n2021 vdd.n1987 9.3005
R19556 vdd.n2020 vdd.n1988 9.3005
R19557 vdd.n1992 vdd.n1989 9.3005
R19558 vdd.n2015 vdd.n1993 9.3005
R19559 vdd.n2014 vdd.n1994 9.3005
R19560 vdd.n2013 vdd.n1995 9.3005
R19561 vdd.n1997 vdd.n1996 9.3005
R19562 vdd.n2008 vdd.n1064 9.3005
R19563 vdd.n2077 vdd.n2076 9.3005
R19564 vdd.n2101 vdd.n2100 9.3005
R19565 vdd.n1907 vdd.n1906 9.3005
R19566 vdd.n1912 vdd.n1910 9.3005
R19567 vdd.n2093 vdd.n1913 9.3005
R19568 vdd.n2092 vdd.n1914 9.3005
R19569 vdd.n2091 vdd.n1915 9.3005
R19570 vdd.n1919 vdd.n1916 9.3005
R19571 vdd.n2086 vdd.n1920 9.3005
R19572 vdd.n2085 vdd.n1921 9.3005
R19573 vdd.n2084 vdd.n1922 9.3005
R19574 vdd.n1926 vdd.n1923 9.3005
R19575 vdd.n2079 vdd.n1927 9.3005
R19576 vdd.n2078 vdd.n1928 9.3005
R19577 vdd.n2323 vdd.n1900 9.3005
R19578 vdd.n2325 vdd.n2324 9.3005
R19579 vdd.n1815 vdd.n1814 9.3005
R19580 vdd.n1124 vdd.n1123 9.3005
R19581 vdd.n1829 vdd.n1828 9.3005
R19582 vdd.n1830 vdd.n1122 9.3005
R19583 vdd.n1832 vdd.n1831 9.3005
R19584 vdd.n1113 vdd.n1112 9.3005
R19585 vdd.n1846 vdd.n1845 9.3005
R19586 vdd.n1847 vdd.n1111 9.3005
R19587 vdd.n1849 vdd.n1848 9.3005
R19588 vdd.n1102 vdd.n1101 9.3005
R19589 vdd.n1862 vdd.n1861 9.3005
R19590 vdd.n1863 vdd.n1100 9.3005
R19591 vdd.n1865 vdd.n1864 9.3005
R19592 vdd.n1090 vdd.n1089 9.3005
R19593 vdd.n1879 vdd.n1878 9.3005
R19594 vdd.n1880 vdd.n1088 9.3005
R19595 vdd.n1882 vdd.n1881 9.3005
R19596 vdd.n1078 vdd.n1077 9.3005
R19597 vdd.n1898 vdd.n1897 9.3005
R19598 vdd.n1899 vdd.n1076 9.3005
R19599 vdd.n2327 vdd.n2326 9.3005
R19600 vdd.n307 vdd.n306 9.3005
R19601 vdd.n302 vdd.n301 9.3005
R19602 vdd.n313 vdd.n312 9.3005
R19603 vdd.n315 vdd.n314 9.3005
R19604 vdd.n298 vdd.n297 9.3005
R19605 vdd.n321 vdd.n320 9.3005
R19606 vdd.n323 vdd.n322 9.3005
R19607 vdd.n295 vdd.n292 9.3005
R19608 vdd.n330 vdd.n329 9.3005
R19609 vdd.n248 vdd.n247 9.3005
R19610 vdd.n243 vdd.n242 9.3005
R19611 vdd.n254 vdd.n253 9.3005
R19612 vdd.n256 vdd.n255 9.3005
R19613 vdd.n239 vdd.n238 9.3005
R19614 vdd.n262 vdd.n261 9.3005
R19615 vdd.n264 vdd.n263 9.3005
R19616 vdd.n236 vdd.n233 9.3005
R19617 vdd.n271 vdd.n270 9.3005
R19618 vdd.n205 vdd.n204 9.3005
R19619 vdd.n200 vdd.n199 9.3005
R19620 vdd.n211 vdd.n210 9.3005
R19621 vdd.n213 vdd.n212 9.3005
R19622 vdd.n196 vdd.n195 9.3005
R19623 vdd.n219 vdd.n218 9.3005
R19624 vdd.n221 vdd.n220 9.3005
R19625 vdd.n193 vdd.n190 9.3005
R19626 vdd.n228 vdd.n227 9.3005
R19627 vdd.n146 vdd.n145 9.3005
R19628 vdd.n141 vdd.n140 9.3005
R19629 vdd.n152 vdd.n151 9.3005
R19630 vdd.n154 vdd.n153 9.3005
R19631 vdd.n137 vdd.n136 9.3005
R19632 vdd.n160 vdd.n159 9.3005
R19633 vdd.n162 vdd.n161 9.3005
R19634 vdd.n134 vdd.n131 9.3005
R19635 vdd.n169 vdd.n168 9.3005
R19636 vdd.n104 vdd.n103 9.3005
R19637 vdd.n99 vdd.n98 9.3005
R19638 vdd.n110 vdd.n109 9.3005
R19639 vdd.n112 vdd.n111 9.3005
R19640 vdd.n95 vdd.n94 9.3005
R19641 vdd.n118 vdd.n117 9.3005
R19642 vdd.n120 vdd.n119 9.3005
R19643 vdd.n92 vdd.n89 9.3005
R19644 vdd.n127 vdd.n126 9.3005
R19645 vdd.n45 vdd.n44 9.3005
R19646 vdd.n40 vdd.n39 9.3005
R19647 vdd.n51 vdd.n50 9.3005
R19648 vdd.n53 vdd.n52 9.3005
R19649 vdd.n36 vdd.n35 9.3005
R19650 vdd.n59 vdd.n58 9.3005
R19651 vdd.n61 vdd.n60 9.3005
R19652 vdd.n33 vdd.n30 9.3005
R19653 vdd.n68 vdd.n67 9.3005
R19654 vdd.n3138 vdd.n3137 9.3005
R19655 vdd.n3141 vdd.n766 9.3005
R19656 vdd.n3142 vdd.n765 9.3005
R19657 vdd.n3145 vdd.n764 9.3005
R19658 vdd.n3146 vdd.n763 9.3005
R19659 vdd.n3149 vdd.n762 9.3005
R19660 vdd.n3150 vdd.n761 9.3005
R19661 vdd.n3153 vdd.n760 9.3005
R19662 vdd.n3154 vdd.n759 9.3005
R19663 vdd.n3157 vdd.n758 9.3005
R19664 vdd.n3158 vdd.n757 9.3005
R19665 vdd.n3161 vdd.n756 9.3005
R19666 vdd.n3162 vdd.n755 9.3005
R19667 vdd.n3165 vdd.n754 9.3005
R19668 vdd.n3166 vdd.n753 9.3005
R19669 vdd.n3169 vdd.n752 9.3005
R19670 vdd.n3170 vdd.n751 9.3005
R19671 vdd.n3173 vdd.n750 9.3005
R19672 vdd.n3174 vdd.n749 9.3005
R19673 vdd.n3177 vdd.n748 9.3005
R19674 vdd.n3181 vdd.n3180 9.3005
R19675 vdd.n3182 vdd.n747 9.3005
R19676 vdd.n3186 vdd.n3183 9.3005
R19677 vdd.n3189 vdd.n746 9.3005
R19678 vdd.n3190 vdd.n745 9.3005
R19679 vdd.n3193 vdd.n744 9.3005
R19680 vdd.n3194 vdd.n743 9.3005
R19681 vdd.n3197 vdd.n742 9.3005
R19682 vdd.n3198 vdd.n741 9.3005
R19683 vdd.n3201 vdd.n740 9.3005
R19684 vdd.n3202 vdd.n739 9.3005
R19685 vdd.n3205 vdd.n738 9.3005
R19686 vdd.n3206 vdd.n737 9.3005
R19687 vdd.n3209 vdd.n736 9.3005
R19688 vdd.n3210 vdd.n735 9.3005
R19689 vdd.n3213 vdd.n730 9.3005
R19690 vdd.n3219 vdd.n727 9.3005
R19691 vdd.n3220 vdd.n726 9.3005
R19692 vdd.n3234 vdd.n3233 9.3005
R19693 vdd.n3235 vdd.n681 9.3005
R19694 vdd.n3237 vdd.n3236 9.3005
R19695 vdd.n671 vdd.n670 9.3005
R19696 vdd.n3251 vdd.n3250 9.3005
R19697 vdd.n3252 vdd.n669 9.3005
R19698 vdd.n3254 vdd.n3253 9.3005
R19699 vdd.n660 vdd.n659 9.3005
R19700 vdd.n3267 vdd.n3266 9.3005
R19701 vdd.n3268 vdd.n658 9.3005
R19702 vdd.n3270 vdd.n3269 9.3005
R19703 vdd.n648 vdd.n647 9.3005
R19704 vdd.n3284 vdd.n3283 9.3005
R19705 vdd.n3285 vdd.n646 9.3005
R19706 vdd.n3287 vdd.n3286 9.3005
R19707 vdd.n637 vdd.n636 9.3005
R19708 vdd.n3303 vdd.n3302 9.3005
R19709 vdd.n3304 vdd.n635 9.3005
R19710 vdd.n3306 vdd.n3305 9.3005
R19711 vdd.n336 vdd.n334 9.3005
R19712 vdd.n683 vdd.n682 9.3005
R19713 vdd.n3398 vdd.n3397 9.3005
R19714 vdd.n337 vdd.n335 9.3005
R19715 vdd.n3391 vdd.n346 9.3005
R19716 vdd.n3390 vdd.n347 9.3005
R19717 vdd.n3389 vdd.n348 9.3005
R19718 vdd.n355 vdd.n349 9.3005
R19719 vdd.n3383 vdd.n356 9.3005
R19720 vdd.n3382 vdd.n357 9.3005
R19721 vdd.n3381 vdd.n358 9.3005
R19722 vdd.n366 vdd.n359 9.3005
R19723 vdd.n3375 vdd.n367 9.3005
R19724 vdd.n3374 vdd.n368 9.3005
R19725 vdd.n3373 vdd.n369 9.3005
R19726 vdd.n377 vdd.n370 9.3005
R19727 vdd.n3367 vdd.n378 9.3005
R19728 vdd.n3366 vdd.n379 9.3005
R19729 vdd.n3365 vdd.n380 9.3005
R19730 vdd.n388 vdd.n381 9.3005
R19731 vdd.n3359 vdd.n389 9.3005
R19732 vdd.n3358 vdd.n390 9.3005
R19733 vdd.n3357 vdd.n391 9.3005
R19734 vdd.n466 vdd.n463 9.3005
R19735 vdd.n470 vdd.n469 9.3005
R19736 vdd.n471 vdd.n462 9.3005
R19737 vdd.n475 vdd.n472 9.3005
R19738 vdd.n476 vdd.n461 9.3005
R19739 vdd.n480 vdd.n479 9.3005
R19740 vdd.n481 vdd.n460 9.3005
R19741 vdd.n485 vdd.n482 9.3005
R19742 vdd.n486 vdd.n459 9.3005
R19743 vdd.n490 vdd.n489 9.3005
R19744 vdd.n491 vdd.n458 9.3005
R19745 vdd.n495 vdd.n492 9.3005
R19746 vdd.n496 vdd.n457 9.3005
R19747 vdd.n500 vdd.n499 9.3005
R19748 vdd.n501 vdd.n456 9.3005
R19749 vdd.n505 vdd.n502 9.3005
R19750 vdd.n506 vdd.n455 9.3005
R19751 vdd.n510 vdd.n509 9.3005
R19752 vdd.n511 vdd.n454 9.3005
R19753 vdd.n515 vdd.n512 9.3005
R19754 vdd.n516 vdd.n451 9.3005
R19755 vdd.n520 vdd.n519 9.3005
R19756 vdd.n521 vdd.n450 9.3005
R19757 vdd.n525 vdd.n522 9.3005
R19758 vdd.n526 vdd.n449 9.3005
R19759 vdd.n530 vdd.n529 9.3005
R19760 vdd.n531 vdd.n448 9.3005
R19761 vdd.n535 vdd.n532 9.3005
R19762 vdd.n536 vdd.n447 9.3005
R19763 vdd.n540 vdd.n539 9.3005
R19764 vdd.n541 vdd.n446 9.3005
R19765 vdd.n545 vdd.n542 9.3005
R19766 vdd.n546 vdd.n445 9.3005
R19767 vdd.n550 vdd.n549 9.3005
R19768 vdd.n551 vdd.n444 9.3005
R19769 vdd.n555 vdd.n552 9.3005
R19770 vdd.n556 vdd.n443 9.3005
R19771 vdd.n560 vdd.n559 9.3005
R19772 vdd.n561 vdd.n442 9.3005
R19773 vdd.n565 vdd.n562 9.3005
R19774 vdd.n566 vdd.n439 9.3005
R19775 vdd.n570 vdd.n569 9.3005
R19776 vdd.n571 vdd.n438 9.3005
R19777 vdd.n575 vdd.n572 9.3005
R19778 vdd.n576 vdd.n437 9.3005
R19779 vdd.n580 vdd.n579 9.3005
R19780 vdd.n581 vdd.n436 9.3005
R19781 vdd.n585 vdd.n582 9.3005
R19782 vdd.n586 vdd.n435 9.3005
R19783 vdd.n590 vdd.n589 9.3005
R19784 vdd.n591 vdd.n434 9.3005
R19785 vdd.n595 vdd.n592 9.3005
R19786 vdd.n596 vdd.n433 9.3005
R19787 vdd.n600 vdd.n599 9.3005
R19788 vdd.n601 vdd.n432 9.3005
R19789 vdd.n605 vdd.n602 9.3005
R19790 vdd.n606 vdd.n431 9.3005
R19791 vdd.n610 vdd.n609 9.3005
R19792 vdd.n611 vdd.n430 9.3005
R19793 vdd.n615 vdd.n612 9.3005
R19794 vdd.n617 vdd.n429 9.3005
R19795 vdd.n619 vdd.n618 9.3005
R19796 vdd.n3351 vdd.n3350 9.3005
R19797 vdd.n465 vdd.n464 9.3005
R19798 vdd.n3229 vdd.n3228 9.3005
R19799 vdd.n676 vdd.n675 9.3005
R19800 vdd.n3242 vdd.n3241 9.3005
R19801 vdd.n3243 vdd.n674 9.3005
R19802 vdd.n3245 vdd.n3244 9.3005
R19803 vdd.n666 vdd.n665 9.3005
R19804 vdd.n3259 vdd.n3258 9.3005
R19805 vdd.n3260 vdd.n664 9.3005
R19806 vdd.n3262 vdd.n3261 9.3005
R19807 vdd.n653 vdd.n652 9.3005
R19808 vdd.n3275 vdd.n3274 9.3005
R19809 vdd.n3276 vdd.n651 9.3005
R19810 vdd.n3278 vdd.n3277 9.3005
R19811 vdd.n642 vdd.n641 9.3005
R19812 vdd.n3292 vdd.n3291 9.3005
R19813 vdd.n3293 vdd.n640 9.3005
R19814 vdd.n3298 vdd.n3294 9.3005
R19815 vdd.n3297 vdd.n3296 9.3005
R19816 vdd.n3295 vdd.n631 9.3005
R19817 vdd.n3311 vdd.n630 9.3005
R19818 vdd.n3313 vdd.n3312 9.3005
R19819 vdd.n3314 vdd.n629 9.3005
R19820 vdd.n3316 vdd.n3315 9.3005
R19821 vdd.n3318 vdd.n628 9.3005
R19822 vdd.n3320 vdd.n3319 9.3005
R19823 vdd.n3321 vdd.n627 9.3005
R19824 vdd.n3323 vdd.n3322 9.3005
R19825 vdd.n3325 vdd.n626 9.3005
R19826 vdd.n3327 vdd.n3326 9.3005
R19827 vdd.n3328 vdd.n625 9.3005
R19828 vdd.n3330 vdd.n3329 9.3005
R19829 vdd.n3333 vdd.n624 9.3005
R19830 vdd.n3335 vdd.n3334 9.3005
R19831 vdd.n3336 vdd.n623 9.3005
R19832 vdd.n3338 vdd.n3337 9.3005
R19833 vdd.n3340 vdd.n622 9.3005
R19834 vdd.n3342 vdd.n3341 9.3005
R19835 vdd.n3343 vdd.n621 9.3005
R19836 vdd.n3345 vdd.n3344 9.3005
R19837 vdd.n3347 vdd.n620 9.3005
R19838 vdd.n3349 vdd.n3348 9.3005
R19839 vdd.n3227 vdd.n686 9.3005
R19840 vdd.n3226 vdd.n3225 9.3005
R19841 vdd.n3095 vdd.n687 9.3005
R19842 vdd.n3104 vdd.n783 9.3005
R19843 vdd.n3107 vdd.n782 9.3005
R19844 vdd.n3108 vdd.n781 9.3005
R19845 vdd.n3111 vdd.n780 9.3005
R19846 vdd.n3112 vdd.n779 9.3005
R19847 vdd.n3115 vdd.n778 9.3005
R19848 vdd.n3116 vdd.n777 9.3005
R19849 vdd.n3119 vdd.n776 9.3005
R19850 vdd.n3120 vdd.n775 9.3005
R19851 vdd.n3123 vdd.n774 9.3005
R19852 vdd.n3124 vdd.n773 9.3005
R19853 vdd.n3127 vdd.n772 9.3005
R19854 vdd.n3128 vdd.n771 9.3005
R19855 vdd.n3131 vdd.n770 9.3005
R19856 vdd.n3135 vdd.n3134 9.3005
R19857 vdd.n3136 vdd.n767 9.3005
R19858 vdd.n2337 vdd.n2336 9.3005
R19859 vdd.n2332 vdd.n1067 9.3005
R19860 vdd.n1430 vdd.n1429 9.3005
R19861 vdd.n1431 vdd.n1185 9.3005
R19862 vdd.n1433 vdd.n1432 9.3005
R19863 vdd.n1175 vdd.n1174 9.3005
R19864 vdd.n1447 vdd.n1446 9.3005
R19865 vdd.n1448 vdd.n1173 9.3005
R19866 vdd.n1450 vdd.n1449 9.3005
R19867 vdd.n1165 vdd.n1164 9.3005
R19868 vdd.n1464 vdd.n1463 9.3005
R19869 vdd.n1465 vdd.n1163 9.3005
R19870 vdd.n1467 vdd.n1466 9.3005
R19871 vdd.n1152 vdd.n1151 9.3005
R19872 vdd.n1480 vdd.n1479 9.3005
R19873 vdd.n1481 vdd.n1150 9.3005
R19874 vdd.n1483 vdd.n1482 9.3005
R19875 vdd.n1141 vdd.n1140 9.3005
R19876 vdd.n1497 vdd.n1496 9.3005
R19877 vdd.n1498 vdd.n1139 9.3005
R19878 vdd.n1500 vdd.n1499 9.3005
R19879 vdd.n1130 vdd.n1129 9.3005
R19880 vdd.n1820 vdd.n1819 9.3005
R19881 vdd.n1821 vdd.n1128 9.3005
R19882 vdd.n1823 vdd.n1822 9.3005
R19883 vdd.n1118 vdd.n1117 9.3005
R19884 vdd.n1837 vdd.n1836 9.3005
R19885 vdd.n1838 vdd.n1116 9.3005
R19886 vdd.n1840 vdd.n1839 9.3005
R19887 vdd.n1108 vdd.n1107 9.3005
R19888 vdd.n1854 vdd.n1853 9.3005
R19889 vdd.n1855 vdd.n1106 9.3005
R19890 vdd.n1857 vdd.n1856 9.3005
R19891 vdd.n1095 vdd.n1094 9.3005
R19892 vdd.n1870 vdd.n1869 9.3005
R19893 vdd.n1871 vdd.n1093 9.3005
R19894 vdd.n1873 vdd.n1872 9.3005
R19895 vdd.n1085 vdd.n1084 9.3005
R19896 vdd.n1887 vdd.n1886 9.3005
R19897 vdd.n1888 vdd.n1082 9.3005
R19898 vdd.n1892 vdd.n1891 9.3005
R19899 vdd.n1890 vdd.n1083 9.3005
R19900 vdd.n1889 vdd.n1072 9.3005
R19901 vdd.n1187 vdd.n1186 9.3005
R19902 vdd.n1323 vdd.n1322 9.3005
R19903 vdd.n1324 vdd.n1313 9.3005
R19904 vdd.n1326 vdd.n1325 9.3005
R19905 vdd.n1327 vdd.n1312 9.3005
R19906 vdd.n1329 vdd.n1328 9.3005
R19907 vdd.n1330 vdd.n1307 9.3005
R19908 vdd.n1332 vdd.n1331 9.3005
R19909 vdd.n1333 vdd.n1306 9.3005
R19910 vdd.n1335 vdd.n1334 9.3005
R19911 vdd.n1336 vdd.n1301 9.3005
R19912 vdd.n1338 vdd.n1337 9.3005
R19913 vdd.n1339 vdd.n1300 9.3005
R19914 vdd.n1341 vdd.n1340 9.3005
R19915 vdd.n1342 vdd.n1295 9.3005
R19916 vdd.n1344 vdd.n1343 9.3005
R19917 vdd.n1345 vdd.n1294 9.3005
R19918 vdd.n1347 vdd.n1346 9.3005
R19919 vdd.n1348 vdd.n1289 9.3005
R19920 vdd.n1350 vdd.n1349 9.3005
R19921 vdd.n1351 vdd.n1288 9.3005
R19922 vdd.n1353 vdd.n1352 9.3005
R19923 vdd.n1357 vdd.n1284 9.3005
R19924 vdd.n1359 vdd.n1358 9.3005
R19925 vdd.n1360 vdd.n1283 9.3005
R19926 vdd.n1362 vdd.n1361 9.3005
R19927 vdd.n1363 vdd.n1278 9.3005
R19928 vdd.n1365 vdd.n1364 9.3005
R19929 vdd.n1366 vdd.n1277 9.3005
R19930 vdd.n1368 vdd.n1367 9.3005
R19931 vdd.n1369 vdd.n1272 9.3005
R19932 vdd.n1371 vdd.n1370 9.3005
R19933 vdd.n1372 vdd.n1271 9.3005
R19934 vdd.n1374 vdd.n1373 9.3005
R19935 vdd.n1375 vdd.n1266 9.3005
R19936 vdd.n1377 vdd.n1376 9.3005
R19937 vdd.n1378 vdd.n1265 9.3005
R19938 vdd.n1380 vdd.n1379 9.3005
R19939 vdd.n1381 vdd.n1260 9.3005
R19940 vdd.n1383 vdd.n1382 9.3005
R19941 vdd.n1384 vdd.n1259 9.3005
R19942 vdd.n1386 vdd.n1385 9.3005
R19943 vdd.n1387 vdd.n1254 9.3005
R19944 vdd.n1389 vdd.n1388 9.3005
R19945 vdd.n1390 vdd.n1253 9.3005
R19946 vdd.n1392 vdd.n1391 9.3005
R19947 vdd.n1393 vdd.n1246 9.3005
R19948 vdd.n1395 vdd.n1394 9.3005
R19949 vdd.n1396 vdd.n1245 9.3005
R19950 vdd.n1398 vdd.n1397 9.3005
R19951 vdd.n1399 vdd.n1240 9.3005
R19952 vdd.n1401 vdd.n1400 9.3005
R19953 vdd.n1402 vdd.n1239 9.3005
R19954 vdd.n1404 vdd.n1403 9.3005
R19955 vdd.n1405 vdd.n1234 9.3005
R19956 vdd.n1407 vdd.n1406 9.3005
R19957 vdd.n1408 vdd.n1233 9.3005
R19958 vdd.n1410 vdd.n1409 9.3005
R19959 vdd.n1411 vdd.n1228 9.3005
R19960 vdd.n1413 vdd.n1412 9.3005
R19961 vdd.n1414 vdd.n1227 9.3005
R19962 vdd.n1416 vdd.n1415 9.3005
R19963 vdd.n1192 vdd.n1191 9.3005
R19964 vdd.n1422 vdd.n1421 9.3005
R19965 vdd.n1321 vdd.n1320 9.3005
R19966 vdd.n1425 vdd.n1424 9.3005
R19967 vdd.n1181 vdd.n1180 9.3005
R19968 vdd.n1439 vdd.n1438 9.3005
R19969 vdd.n1440 vdd.n1179 9.3005
R19970 vdd.n1442 vdd.n1441 9.3005
R19971 vdd.n1170 vdd.n1169 9.3005
R19972 vdd.n1456 vdd.n1455 9.3005
R19973 vdd.n1457 vdd.n1168 9.3005
R19974 vdd.n1459 vdd.n1458 9.3005
R19975 vdd.n1159 vdd.n1158 9.3005
R19976 vdd.n1472 vdd.n1471 9.3005
R19977 vdd.n1473 vdd.n1157 9.3005
R19978 vdd.n1475 vdd.n1474 9.3005
R19979 vdd.n1147 vdd.n1146 9.3005
R19980 vdd.n1489 vdd.n1488 9.3005
R19981 vdd.n1490 vdd.n1145 9.3005
R19982 vdd.n1492 vdd.n1491 9.3005
R19983 vdd.n1136 vdd.n1135 9.3005
R19984 vdd.n1505 vdd.n1504 9.3005
R19985 vdd.n1506 vdd.n1134 9.3005
R19986 vdd.n1423 vdd.n1190 9.3005
R19987 vdd.n1726 vdd.n1725 9.3005
R19988 vdd.n1721 vdd.n1720 9.3005
R19989 vdd.n1732 vdd.n1731 9.3005
R19990 vdd.n1734 vdd.n1733 9.3005
R19991 vdd.n1717 vdd.n1716 9.3005
R19992 vdd.n1740 vdd.n1739 9.3005
R19993 vdd.n1742 vdd.n1741 9.3005
R19994 vdd.n1714 vdd.n1711 9.3005
R19995 vdd.n1749 vdd.n1748 9.3005
R19996 vdd.n1785 vdd.n1784 9.3005
R19997 vdd.n1780 vdd.n1779 9.3005
R19998 vdd.n1791 vdd.n1790 9.3005
R19999 vdd.n1793 vdd.n1792 9.3005
R20000 vdd.n1776 vdd.n1775 9.3005
R20001 vdd.n1799 vdd.n1798 9.3005
R20002 vdd.n1801 vdd.n1800 9.3005
R20003 vdd.n1773 vdd.n1770 9.3005
R20004 vdd.n1808 vdd.n1807 9.3005
R20005 vdd.n1624 vdd.n1623 9.3005
R20006 vdd.n1619 vdd.n1618 9.3005
R20007 vdd.n1630 vdd.n1629 9.3005
R20008 vdd.n1632 vdd.n1631 9.3005
R20009 vdd.n1615 vdd.n1614 9.3005
R20010 vdd.n1638 vdd.n1637 9.3005
R20011 vdd.n1640 vdd.n1639 9.3005
R20012 vdd.n1612 vdd.n1609 9.3005
R20013 vdd.n1647 vdd.n1646 9.3005
R20014 vdd.n1683 vdd.n1682 9.3005
R20015 vdd.n1678 vdd.n1677 9.3005
R20016 vdd.n1689 vdd.n1688 9.3005
R20017 vdd.n1691 vdd.n1690 9.3005
R20018 vdd.n1674 vdd.n1673 9.3005
R20019 vdd.n1697 vdd.n1696 9.3005
R20020 vdd.n1699 vdd.n1698 9.3005
R20021 vdd.n1671 vdd.n1668 9.3005
R20022 vdd.n1706 vdd.n1705 9.3005
R20023 vdd.n1523 vdd.n1522 9.3005
R20024 vdd.n1518 vdd.n1517 9.3005
R20025 vdd.n1529 vdd.n1528 9.3005
R20026 vdd.n1531 vdd.n1530 9.3005
R20027 vdd.n1514 vdd.n1513 9.3005
R20028 vdd.n1537 vdd.n1536 9.3005
R20029 vdd.n1539 vdd.n1538 9.3005
R20030 vdd.n1511 vdd.n1508 9.3005
R20031 vdd.n1546 vdd.n1545 9.3005
R20032 vdd.n1582 vdd.n1581 9.3005
R20033 vdd.n1577 vdd.n1576 9.3005
R20034 vdd.n1588 vdd.n1587 9.3005
R20035 vdd.n1590 vdd.n1589 9.3005
R20036 vdd.n1573 vdd.n1572 9.3005
R20037 vdd.n1596 vdd.n1595 9.3005
R20038 vdd.n1598 vdd.n1597 9.3005
R20039 vdd.n1570 vdd.n1567 9.3005
R20040 vdd.n1605 vdd.n1604 9.3005
R20041 vdd.n1461 vdd.t165 9.18308
R20042 vdd.n3331 vdd.t231 9.18308
R20043 vdd.n1155 vdd.t215 8.95635
R20044 vdd.n2329 vdd.t42 8.95635
R20045 vdd.n723 vdd.t35 8.95635
R20046 vdd.t179 vdd.n3385 8.95635
R20047 vdd.n312 vdd.n311 8.92171
R20048 vdd.n253 vdd.n252 8.92171
R20049 vdd.n210 vdd.n209 8.92171
R20050 vdd.n151 vdd.n150 8.92171
R20051 vdd.n109 vdd.n108 8.92171
R20052 vdd.n50 vdd.n49 8.92171
R20053 vdd.n1731 vdd.n1730 8.92171
R20054 vdd.n1790 vdd.n1789 8.92171
R20055 vdd.n1629 vdd.n1628 8.92171
R20056 vdd.n1688 vdd.n1687 8.92171
R20057 vdd.n1528 vdd.n1527 8.92171
R20058 vdd.n1587 vdd.n1586 8.92171
R20059 vdd.n231 vdd.n129 8.81535
R20060 vdd.n1709 vdd.n1607 8.81535
R20061 vdd.n1502 vdd.t185 8.72962
R20062 vdd.t176 vdd.n3394 8.72962
R20063 vdd.n1825 vdd.t235 8.50289
R20064 vdd.n3300 vdd.t181 8.50289
R20065 vdd.n28 vdd.n14 8.42249
R20066 vdd.n1851 vdd.t171 8.27616
R20067 vdd.t173 vdd.n656 8.27616
R20068 vdd.n3400 vdd.n3399 8.16225
R20069 vdd.n1813 vdd.n1812 8.16225
R20070 vdd.n308 vdd.n302 8.14595
R20071 vdd.n249 vdd.n243 8.14595
R20072 vdd.n206 vdd.n200 8.14595
R20073 vdd.n147 vdd.n141 8.14595
R20074 vdd.n105 vdd.n99 8.14595
R20075 vdd.n46 vdd.n40 8.14595
R20076 vdd.n1727 vdd.n1721 8.14595
R20077 vdd.n1786 vdd.n1780 8.14595
R20078 vdd.n1625 vdd.n1619 8.14595
R20079 vdd.n1684 vdd.n1678 8.14595
R20080 vdd.n1524 vdd.n1518 8.14595
R20081 vdd.n1583 vdd.n1577 8.14595
R20082 vdd.n2923 vdd.n849 8.11757
R20083 vdd.n2397 vdd.n2396 8.11757
R20084 vdd.n1098 vdd.t260 8.04943
R20085 vdd.n3256 vdd.t213 8.04943
R20086 vdd.n2375 vdd.n1043 7.70933
R20087 vdd.n2381 vdd.n1043 7.70933
R20088 vdd.n2387 vdd.n1037 7.70933
R20089 vdd.n2387 vdd.n1030 7.70933
R20090 vdd.n2393 vdd.n1030 7.70933
R20091 vdd.n2393 vdd.n1033 7.70933
R20092 vdd.n2400 vdd.n1018 7.70933
R20093 vdd.n2406 vdd.n1018 7.70933
R20094 vdd.n2412 vdd.n1012 7.70933
R20095 vdd.n2418 vdd.n1008 7.70933
R20096 vdd.n2424 vdd.n1002 7.70933
R20097 vdd.n2436 vdd.n989 7.70933
R20098 vdd.n2442 vdd.n983 7.70933
R20099 vdd.n2442 vdd.n976 7.70933
R20100 vdd.n2450 vdd.n976 7.70933
R20101 vdd.n2457 vdd.t5 7.70933
R20102 vdd.n2532 vdd.t5 7.70933
R20103 vdd.n2864 vdd.t288 7.70933
R20104 vdd.n2870 vdd.t288 7.70933
R20105 vdd.n2876 vdd.n897 7.70933
R20106 vdd.n2882 vdd.n897 7.70933
R20107 vdd.n2882 vdd.n900 7.70933
R20108 vdd.n2888 vdd.n893 7.70933
R20109 vdd.n2900 vdd.n880 7.70933
R20110 vdd.n2906 vdd.n874 7.70933
R20111 vdd.n2912 vdd.n870 7.70933
R20112 vdd.n2918 vdd.n857 7.70933
R20113 vdd.n2926 vdd.n857 7.70933
R20114 vdd.n2932 vdd.n851 7.70933
R20115 vdd.n2932 vdd.n843 7.70933
R20116 vdd.n2983 vdd.n843 7.70933
R20117 vdd.n2983 vdd.n846 7.70933
R20118 vdd.n2989 vdd.n805 7.70933
R20119 vdd.n3059 vdd.n805 7.70933
R20120 vdd.n307 vdd.n304 7.3702
R20121 vdd.n248 vdd.n245 7.3702
R20122 vdd.n205 vdd.n202 7.3702
R20123 vdd.n146 vdd.n143 7.3702
R20124 vdd.n104 vdd.n101 7.3702
R20125 vdd.n45 vdd.n42 7.3702
R20126 vdd.n1726 vdd.n1723 7.3702
R20127 vdd.n1785 vdd.n1782 7.3702
R20128 vdd.n1624 vdd.n1621 7.3702
R20129 vdd.n1683 vdd.n1680 7.3702
R20130 vdd.n1523 vdd.n1520 7.3702
R20131 vdd.n1582 vdd.n1579 7.3702
R20132 vdd.n1884 vdd.t123 7.1425
R20133 vdd.n679 vdd.t125 7.1425
R20134 vdd.n1358 vdd.n1357 6.98232
R20135 vdd.n2039 vdd.n2038 6.98232
R20136 vdd.n566 vdd.n565 6.98232
R20137 vdd.n3141 vdd.n3138 6.98232
R20138 vdd.t237 vdd.n1097 6.91577
R20139 vdd.n3264 vdd.t133 6.91577
R20140 vdd.n1843 vdd.t196 6.68904
R20141 vdd.n3280 vdd.t153 6.68904
R20142 vdd.t135 vdd.n1126 6.46231
R20143 vdd.n3308 vdd.t137 6.46231
R20144 vdd.n3400 vdd.n333 6.38151
R20145 vdd.n1812 vdd.n1811 6.38151
R20146 vdd.n1494 vdd.t168 6.23558
R20147 vdd.t208 vdd.n344 6.23558
R20148 vdd.t139 vdd.n1154 6.00885
R20149 vdd.n2412 vdd.t0 6.00885
R20150 vdd.n2912 vdd.t4 6.00885
R20151 vdd.n3379 vdd.t151 6.00885
R20152 vdd.n1033 vdd.t89 5.89549
R20153 vdd.t46 vdd.n851 5.89549
R20154 vdd.n308 vdd.n307 5.81868
R20155 vdd.n249 vdd.n248 5.81868
R20156 vdd.n206 vdd.n205 5.81868
R20157 vdd.n147 vdd.n146 5.81868
R20158 vdd.n105 vdd.n104 5.81868
R20159 vdd.n46 vdd.n45 5.81868
R20160 vdd.n1727 vdd.n1726 5.81868
R20161 vdd.n1786 vdd.n1785 5.81868
R20162 vdd.n1625 vdd.n1624 5.81868
R20163 vdd.n1684 vdd.n1683 5.81868
R20164 vdd.n1524 vdd.n1523 5.81868
R20165 vdd.n1583 vdd.n1582 5.81868
R20166 vdd.n1453 vdd.t127 5.78212
R20167 vdd.t85 vdd.n1037 5.78212
R20168 vdd.n2156 vdd.t70 5.78212
R20169 vdd.n2781 vdd.t78 5.78212
R20170 vdd.n846 vdd.t74 5.78212
R20171 vdd.n3370 vdd.t203 5.78212
R20172 vdd.n2540 vdd.n2539 5.77611
R20173 vdd.n2283 vdd.n2153 5.77611
R20174 vdd.n2794 vdd.n2793 5.77611
R20175 vdd.n3000 vdd.n2999 5.77611
R20176 vdd.n3064 vdd.n801 5.77611
R20177 vdd.n2704 vdd.n2644 5.77611
R20178 vdd.n2465 vdd.n967 5.77611
R20179 vdd.n2213 vdd.n2212 5.77611
R20180 vdd.n1320 vdd.n1319 5.62474
R20181 vdd.n2335 vdd.n2332 5.62474
R20182 vdd.n3351 vdd.n428 5.62474
R20183 vdd.n3225 vdd.n690 5.62474
R20184 vdd.n1177 vdd.t127 5.55539
R20185 vdd.t203 vdd.n3369 5.55539
R20186 vdd.t292 vdd.n989 5.44203
R20187 vdd.n893 vdd.t14 5.44203
R20188 vdd.n1469 vdd.t139 5.32866
R20189 vdd.t151 vdd.n3378 5.32866
R20190 vdd.n1485 vdd.t168 5.10193
R20191 vdd.t110 vdd.n1012 5.10193
R20192 vdd.n1002 vdd.t3 5.10193
R20193 vdd.t283 vdd.n880 5.10193
R20194 vdd.n870 vdd.t9 5.10193
R20195 vdd.n3387 vdd.t208 5.10193
R20196 vdd.n311 vdd.n302 5.04292
R20197 vdd.n252 vdd.n243 5.04292
R20198 vdd.n209 vdd.n200 5.04292
R20199 vdd.n150 vdd.n141 5.04292
R20200 vdd.n108 vdd.n99 5.04292
R20201 vdd.n49 vdd.n40 5.04292
R20202 vdd.n1730 vdd.n1721 5.04292
R20203 vdd.n1789 vdd.n1780 5.04292
R20204 vdd.n1628 vdd.n1619 5.04292
R20205 vdd.n1687 vdd.n1678 5.04292
R20206 vdd.n1527 vdd.n1518 5.04292
R20207 vdd.n1586 vdd.n1577 5.04292
R20208 vdd.n1817 vdd.t135 4.8752
R20209 vdd.t33 vdd.t7 4.8752
R20210 vdd.t11 vdd.t284 4.8752
R20211 vdd.t1 vdd.t16 4.8752
R20212 vdd.t294 vdd.t116 4.8752
R20213 vdd.t137 vdd.n340 4.8752
R20214 vdd.n2541 vdd.n2540 4.83952
R20215 vdd.n2153 vdd.n2149 4.83952
R20216 vdd.n2795 vdd.n2794 4.83952
R20217 vdd.n3001 vdd.n3000 4.83952
R20218 vdd.n801 vdd.n796 4.83952
R20219 vdd.n2701 vdd.n2644 4.83952
R20220 vdd.n2468 vdd.n967 4.83952
R20221 vdd.n2212 vdd.n2211 4.83952
R20222 vdd.n2007 vdd.n1065 4.74817
R20223 vdd.n2002 vdd.n1066 4.74817
R20224 vdd.n1904 vdd.n1901 4.74817
R20225 vdd.n2316 vdd.n1905 4.74817
R20226 vdd.n2318 vdd.n1904 4.74817
R20227 vdd.n2317 vdd.n2316 4.74817
R20228 vdd.n3218 vdd.n3217 4.74817
R20229 vdd.n3215 vdd.n3214 4.74817
R20230 vdd.n3215 vdd.n732 4.74817
R20231 vdd.n3217 vdd.n729 4.74817
R20232 vdd.n3100 vdd.n784 4.74817
R20233 vdd.n3096 vdd.n3094 4.74817
R20234 vdd.n3099 vdd.n3094 4.74817
R20235 vdd.n3103 vdd.n784 4.74817
R20236 vdd.n2003 vdd.n1065 4.74817
R20237 vdd.n1068 vdd.n1066 4.74817
R20238 vdd.n333 vdd.n332 4.7074
R20239 vdd.n231 vdd.n230 4.7074
R20240 vdd.n1811 vdd.n1810 4.7074
R20241 vdd.n1709 vdd.n1708 4.7074
R20242 vdd.n1120 vdd.t196 4.64847
R20243 vdd.n3289 vdd.t153 4.64847
R20244 vdd.n2418 vdd.t121 4.53511
R20245 vdd.n2906 vdd.t119 4.53511
R20246 vdd.n1859 vdd.t237 4.42174
R20247 vdd.t133 vdd.n655 4.42174
R20248 vdd.n2450 vdd.t117 4.30838
R20249 vdd.n2876 vdd.t114 4.30838
R20250 vdd.n312 vdd.n300 4.26717
R20251 vdd.n253 vdd.n241 4.26717
R20252 vdd.n210 vdd.n198 4.26717
R20253 vdd.n151 vdd.n139 4.26717
R20254 vdd.n109 vdd.n97 4.26717
R20255 vdd.n50 vdd.n38 4.26717
R20256 vdd.n1731 vdd.n1719 4.26717
R20257 vdd.n1790 vdd.n1778 4.26717
R20258 vdd.n1629 vdd.n1617 4.26717
R20259 vdd.n1688 vdd.n1676 4.26717
R20260 vdd.n1528 vdd.n1516 4.26717
R20261 vdd.n1587 vdd.n1575 4.26717
R20262 vdd.n1875 vdd.t123 4.19501
R20263 vdd.n3248 vdd.t125 4.19501
R20264 vdd.n333 vdd.n231 4.10845
R20265 vdd.n1811 vdd.n1709 4.10845
R20266 vdd.n289 vdd.t167 4.06363
R20267 vdd.n289 vdd.t224 4.06363
R20268 vdd.n287 vdd.t258 4.06363
R20269 vdd.n287 vdd.t275 4.06363
R20270 vdd.n285 vdd.t277 4.06363
R20271 vdd.n285 vdd.t170 4.06363
R20272 vdd.n283 vdd.t195 4.06363
R20273 vdd.n283 vdd.t276 4.06363
R20274 vdd.n281 vdd.t278 4.06363
R20275 vdd.n281 vdd.t194 4.06363
R20276 vdd.n279 vdd.t199 4.06363
R20277 vdd.n279 vdd.t201 4.06363
R20278 vdd.n277 vdd.t251 4.06363
R20279 vdd.n277 vdd.t154 4.06363
R20280 vdd.n275 vdd.t159 4.06363
R20281 vdd.n275 vdd.t223 4.06363
R20282 vdd.n273 vdd.t227 4.06363
R20283 vdd.n273 vdd.t257 4.06363
R20284 vdd.n187 vdd.t144 4.06363
R20285 vdd.n187 vdd.t204 4.06363
R20286 vdd.n185 vdd.t242 4.06363
R20287 vdd.n185 vdd.t262 4.06363
R20288 vdd.n183 vdd.t265 4.06363
R20289 vdd.n183 vdd.t146 4.06363
R20290 vdd.n181 vdd.t178 4.06363
R20291 vdd.n181 vdd.t264 4.06363
R20292 vdd.n179 vdd.t268 4.06363
R20293 vdd.n179 vdd.t177 4.06363
R20294 vdd.n177 vdd.t182 4.06363
R20295 vdd.n177 vdd.t184 4.06363
R20296 vdd.n175 vdd.t240 4.06363
R20297 vdd.n175 vdd.t282 4.06363
R20298 vdd.n173 vdd.t134 4.06363
R20299 vdd.n173 vdd.t202 4.06363
R20300 vdd.n171 vdd.t214 4.06363
R20301 vdd.n171 vdd.t243 4.06363
R20302 vdd.n86 vdd.t164 4.06363
R20303 vdd.n86 vdd.t249 4.06363
R20304 vdd.n84 vdd.t152 4.06363
R20305 vdd.n84 vdd.t232 4.06363
R20306 vdd.n82 vdd.t180 4.06363
R20307 vdd.n82 vdd.t259 4.06363
R20308 vdd.n80 vdd.t148 4.06363
R20309 vdd.n80 vdd.t209 4.06363
R20310 vdd.n78 vdd.t138 4.06363
R20311 vdd.n78 vdd.t187 4.06363
R20312 vdd.n76 vdd.t274 4.06363
R20313 vdd.n76 vdd.t247 4.06363
R20314 vdd.n74 vdd.t252 4.06363
R20315 vdd.n74 vdd.t198 4.06363
R20316 vdd.n72 vdd.t280 4.06363
R20317 vdd.n72 vdd.t174 4.06363
R20318 vdd.n70 vdd.t266 4.06363
R20319 vdd.n70 vdd.t207 4.06363
R20320 vdd.n1751 vdd.t161 4.06363
R20321 vdd.n1751 vdd.t271 4.06363
R20322 vdd.n1753 vdd.t270 4.06363
R20323 vdd.n1753 vdd.t250 4.06363
R20324 vdd.n1755 vdd.t219 4.06363
R20325 vdd.n1755 vdd.t158 4.06363
R20326 vdd.n1757 vdd.t281 4.06363
R20327 vdd.n1757 vdd.t248 4.06363
R20328 vdd.n1759 vdd.t244 4.06363
R20329 vdd.n1759 vdd.t193 4.06363
R20330 vdd.n1761 vdd.t191 4.06363
R20331 vdd.n1761 vdd.t245 4.06363
R20332 vdd.n1763 vdd.t228 4.06363
R20333 vdd.n1763 vdd.t229 4.06363
R20334 vdd.n1765 vdd.t188 4.06363
R20335 vdd.n1765 vdd.t160 4.06363
R20336 vdd.n1767 vdd.t157 4.06363
R20337 vdd.n1767 vdd.t225 4.06363
R20338 vdd.n1649 vdd.t142 4.06363
R20339 vdd.n1649 vdd.t261 4.06363
R20340 vdd.n1651 vdd.t253 4.06363
R20341 vdd.n1651 vdd.t238 4.06363
R20342 vdd.n1653 vdd.t200 4.06363
R20343 vdd.n1653 vdd.t132 4.06363
R20344 vdd.n1655 vdd.t269 4.06363
R20345 vdd.n1655 vdd.t236 4.06363
R20346 vdd.n1657 vdd.t230 4.06363
R20347 vdd.n1657 vdd.t175 4.06363
R20348 vdd.n1659 vdd.t169 4.06363
R20349 vdd.n1659 vdd.t233 4.06363
R20350 vdd.n1661 vdd.t218 4.06363
R20351 vdd.n1661 vdd.t216 4.06363
R20352 vdd.n1663 vdd.t166 4.06363
R20353 vdd.n1663 vdd.t140 4.06363
R20354 vdd.n1665 vdd.t128 4.06363
R20355 vdd.n1665 vdd.t211 4.06363
R20356 vdd.n1548 vdd.t205 4.06363
R20357 vdd.n1548 vdd.t267 4.06363
R20358 vdd.n1550 vdd.t172 4.06363
R20359 vdd.n1550 vdd.t246 4.06363
R20360 vdd.n1552 vdd.t197 4.06363
R20361 vdd.n1552 vdd.t255 4.06363
R20362 vdd.n1554 vdd.t222 4.06363
R20363 vdd.n1554 vdd.t273 4.06363
R20364 vdd.n1556 vdd.t186 4.06363
R20365 vdd.n1556 vdd.t136 4.06363
R20366 vdd.n1558 vdd.t210 4.06363
R20367 vdd.n1558 vdd.t150 4.06363
R20368 vdd.n1560 vdd.t263 4.06363
R20369 vdd.n1560 vdd.t279 4.06363
R20370 vdd.n1562 vdd.t234 4.06363
R20371 vdd.n1562 vdd.t155 4.06363
R20372 vdd.n1564 vdd.t220 4.06363
R20373 vdd.n1564 vdd.t163 4.06363
R20374 vdd.n26 vdd.t28 3.9605
R20375 vdd.n26 vdd.t18 3.9605
R20376 vdd.n23 vdd.t31 3.9605
R20377 vdd.n23 vdd.t30 3.9605
R20378 vdd.n21 vdd.t29 3.9605
R20379 vdd.n21 vdd.t17 3.9605
R20380 vdd.n20 vdd.t26 3.9605
R20381 vdd.n20 vdd.t22 3.9605
R20382 vdd.n15 vdd.t24 3.9605
R20383 vdd.n15 vdd.t23 3.9605
R20384 vdd.n16 vdd.t19 3.9605
R20385 vdd.n16 vdd.t25 3.9605
R20386 vdd.n18 vdd.t20 3.9605
R20387 vdd.n18 vdd.t21 3.9605
R20388 vdd.n25 vdd.t32 3.9605
R20389 vdd.n25 vdd.t27 3.9605
R20390 vdd.n7 vdd.t295 3.61217
R20391 vdd.n7 vdd.t120 3.61217
R20392 vdd.n8 vdd.t2 3.61217
R20393 vdd.n8 vdd.t15 3.61217
R20394 vdd.n10 vdd.t289 3.61217
R20395 vdd.n10 vdd.t115 3.61217
R20396 vdd.n12 vdd.t112 3.61217
R20397 vdd.n12 vdd.t291 3.61217
R20398 vdd.n5 vdd.t13 3.61217
R20399 vdd.n5 vdd.t287 3.61217
R20400 vdd.n3 vdd.t118 3.61217
R20401 vdd.n3 vdd.t6 3.61217
R20402 vdd.n1 vdd.t293 3.61217
R20403 vdd.n1 vdd.t285 3.61217
R20404 vdd.n0 vdd.t122 3.61217
R20405 vdd.n0 vdd.t8 3.61217
R20406 vdd.n316 vdd.n315 3.49141
R20407 vdd.n257 vdd.n256 3.49141
R20408 vdd.n214 vdd.n213 3.49141
R20409 vdd.n155 vdd.n154 3.49141
R20410 vdd.n113 vdd.n112 3.49141
R20411 vdd.n54 vdd.n53 3.49141
R20412 vdd.n1735 vdd.n1734 3.49141
R20413 vdd.n1794 vdd.n1793 3.49141
R20414 vdd.n1633 vdd.n1632 3.49141
R20415 vdd.n1692 vdd.n1691 3.49141
R20416 vdd.n1532 vdd.n1531 3.49141
R20417 vdd.n1591 vdd.n1590 3.49141
R20418 vdd.n2156 vdd.t117 3.40145
R20419 vdd.n2604 vdd.t12 3.40145
R20420 vdd.n2857 vdd.t290 3.40145
R20421 vdd.n2781 vdd.t114 3.40145
R20422 vdd.n1876 vdd.t260 3.28809
R20423 vdd.n3247 vdd.t213 3.28809
R20424 vdd.n2257 vdd.t121 3.17472
R20425 vdd.n2760 vdd.t119 3.17472
R20426 vdd.t171 vdd.n1104 3.06136
R20427 vdd.n3272 vdd.t173 3.06136
R20428 vdd.n1834 vdd.t235 2.83463
R20429 vdd.n644 vdd.t181 2.83463
R20430 vdd.n319 vdd.n298 2.71565
R20431 vdd.n260 vdd.n239 2.71565
R20432 vdd.n217 vdd.n196 2.71565
R20433 vdd.n158 vdd.n137 2.71565
R20434 vdd.n116 vdd.n95 2.71565
R20435 vdd.n57 vdd.n36 2.71565
R20436 vdd.n1738 vdd.n1717 2.71565
R20437 vdd.n1797 vdd.n1776 2.71565
R20438 vdd.n1636 vdd.n1615 2.71565
R20439 vdd.n1695 vdd.n1674 2.71565
R20440 vdd.n1535 vdd.n1514 2.71565
R20441 vdd.n1594 vdd.n1573 2.71565
R20442 vdd.t185 vdd.n1132 2.6079
R20443 vdd.n2406 vdd.t110 2.6079
R20444 vdd.n2430 vdd.t3 2.6079
R20445 vdd.n2894 vdd.t283 2.6079
R20446 vdd.n2918 vdd.t9 2.6079
R20447 vdd.n3395 vdd.t176 2.6079
R20448 vdd.n2924 vdd.n2923 2.49806
R20449 vdd.n2398 vdd.n2397 2.49806
R20450 vdd.n306 vdd.n305 2.4129
R20451 vdd.n247 vdd.n246 2.4129
R20452 vdd.n204 vdd.n203 2.4129
R20453 vdd.n145 vdd.n144 2.4129
R20454 vdd.n103 vdd.n102 2.4129
R20455 vdd.n44 vdd.n43 2.4129
R20456 vdd.n1725 vdd.n1724 2.4129
R20457 vdd.n1784 vdd.n1783 2.4129
R20458 vdd.n1623 vdd.n1622 2.4129
R20459 vdd.n1682 vdd.n1681 2.4129
R20460 vdd.n1522 vdd.n1521 2.4129
R20461 vdd.n1581 vdd.n1580 2.4129
R20462 vdd.n1486 vdd.t215 2.38117
R20463 vdd.n1894 vdd.t42 2.38117
R20464 vdd.n3231 vdd.t35 2.38117
R20465 vdd.n3386 vdd.t179 2.38117
R20466 vdd.n2315 vdd.n1904 2.27742
R20467 vdd.n2316 vdd.n2315 2.27742
R20468 vdd.n3216 vdd.n3215 2.27742
R20469 vdd.n3217 vdd.n3216 2.27742
R20470 vdd.n3094 vdd.n3093 2.27742
R20471 vdd.n3093 vdd.n784 2.27742
R20472 vdd.n2338 vdd.n1065 2.27742
R20473 vdd.n2338 vdd.n1066 2.27742
R20474 vdd.n2430 vdd.t292 2.2678
R20475 vdd.n2894 vdd.t14 2.2678
R20476 vdd.t165 vdd.n1161 2.15444
R20477 vdd.n3377 vdd.t231 2.15444
R20478 vdd.t284 vdd.n983 2.04107
R20479 vdd.n900 vdd.t1 2.04107
R20480 vdd.n320 vdd.n296 1.93989
R20481 vdd.n261 vdd.n237 1.93989
R20482 vdd.n218 vdd.n194 1.93989
R20483 vdd.n159 vdd.n135 1.93989
R20484 vdd.n117 vdd.n93 1.93989
R20485 vdd.n58 vdd.n34 1.93989
R20486 vdd.n1739 vdd.n1715 1.93989
R20487 vdd.n1798 vdd.n1774 1.93989
R20488 vdd.n1637 vdd.n1613 1.93989
R20489 vdd.n1696 vdd.n1672 1.93989
R20490 vdd.n1536 vdd.n1512 1.93989
R20491 vdd.n1595 vdd.n1571 1.93989
R20492 vdd.n1444 vdd.t129 1.92771
R20493 vdd.n2381 vdd.t85 1.92771
R20494 vdd.n2457 vdd.t70 1.92771
R20495 vdd.n2870 vdd.t78 1.92771
R20496 vdd.n2989 vdd.t74 1.92771
R20497 vdd.t189 vdd.n375 1.92771
R20498 vdd.n1452 vdd.t162 1.70098
R20499 vdd.n2257 vdd.t0 1.70098
R20500 vdd.n1008 vdd.t33 1.70098
R20501 vdd.t116 vdd.n874 1.70098
R20502 vdd.n2760 vdd.t4 1.70098
R20503 vdd.n3371 vdd.t143 1.70098
R20504 vdd.n1477 vdd.t217 1.47425
R20505 vdd.n361 vdd.t145 1.47425
R20506 vdd.n1143 vdd.t149 1.24752
R20507 vdd.t147 vdd.n3393 1.24752
R20508 vdd.n331 vdd.n291 1.16414
R20509 vdd.n324 vdd.n323 1.16414
R20510 vdd.n272 vdd.n232 1.16414
R20511 vdd.n265 vdd.n264 1.16414
R20512 vdd.n229 vdd.n189 1.16414
R20513 vdd.n222 vdd.n221 1.16414
R20514 vdd.n170 vdd.n130 1.16414
R20515 vdd.n163 vdd.n162 1.16414
R20516 vdd.n128 vdd.n88 1.16414
R20517 vdd.n121 vdd.n120 1.16414
R20518 vdd.n69 vdd.n29 1.16414
R20519 vdd.n62 vdd.n61 1.16414
R20520 vdd.n1750 vdd.n1710 1.16414
R20521 vdd.n1743 vdd.n1742 1.16414
R20522 vdd.n1809 vdd.n1769 1.16414
R20523 vdd.n1802 vdd.n1801 1.16414
R20524 vdd.n1648 vdd.n1608 1.16414
R20525 vdd.n1641 vdd.n1640 1.16414
R20526 vdd.n1707 vdd.n1667 1.16414
R20527 vdd.n1700 vdd.n1699 1.16414
R20528 vdd.n1547 vdd.n1507 1.16414
R20529 vdd.n1540 vdd.n1539 1.16414
R20530 vdd.n1606 vdd.n1566 1.16414
R20531 vdd.n1599 vdd.n1598 1.16414
R20532 vdd.n2424 vdd.t7 1.13415
R20533 vdd.n2900 vdd.t294 1.13415
R20534 vdd.n1826 vdd.t221 1.02079
R20535 vdd.t89 vdd.t10 1.02079
R20536 vdd.t113 vdd.t46 1.02079
R20537 vdd.t183 vdd.n633 1.02079
R20538 vdd.n1323 vdd.n1319 0.970197
R20539 vdd.n2336 vdd.n2335 0.970197
R20540 vdd.n618 vdd.n428 0.970197
R20541 vdd.n3095 vdd.n690 0.970197
R20542 vdd.n1812 vdd.n28 0.90431
R20543 vdd vdd.n3400 0.896477
R20544 vdd.n1842 vdd.t131 0.794056
R20545 vdd.n2400 vdd.t10 0.794056
R20546 vdd.n2436 vdd.t11 0.794056
R20547 vdd.n2888 vdd.t16 0.794056
R20548 vdd.n2926 vdd.t113 0.794056
R20549 vdd.n3281 vdd.t239 0.794056
R20550 vdd.n1867 vdd.t141 0.567326
R20551 vdd.t206 vdd.n662 0.567326
R20552 vdd.n2326 vdd.n2325 0.530988
R20553 vdd.n726 vdd.n682 0.530988
R20554 vdd.n464 vdd.n391 0.530988
R20555 vdd.n3350 vdd.n3349 0.530988
R20556 vdd.n3227 vdd.n3226 0.530988
R20557 vdd.n1889 vdd.n1067 0.530988
R20558 vdd.n1321 vdd.n1186 0.530988
R20559 vdd.n1423 vdd.n1422 0.530988
R20560 vdd.n4 vdd.n2 0.459552
R20561 vdd.n11 vdd.n9 0.459552
R20562 vdd.n329 vdd.n328 0.388379
R20563 vdd.n295 vdd.n293 0.388379
R20564 vdd.n270 vdd.n269 0.388379
R20565 vdd.n236 vdd.n234 0.388379
R20566 vdd.n227 vdd.n226 0.388379
R20567 vdd.n193 vdd.n191 0.388379
R20568 vdd.n168 vdd.n167 0.388379
R20569 vdd.n134 vdd.n132 0.388379
R20570 vdd.n126 vdd.n125 0.388379
R20571 vdd.n92 vdd.n90 0.388379
R20572 vdd.n67 vdd.n66 0.388379
R20573 vdd.n33 vdd.n31 0.388379
R20574 vdd.n1748 vdd.n1747 0.388379
R20575 vdd.n1714 vdd.n1712 0.388379
R20576 vdd.n1807 vdd.n1806 0.388379
R20577 vdd.n1773 vdd.n1771 0.388379
R20578 vdd.n1646 vdd.n1645 0.388379
R20579 vdd.n1612 vdd.n1610 0.388379
R20580 vdd.n1705 vdd.n1704 0.388379
R20581 vdd.n1671 vdd.n1669 0.388379
R20582 vdd.n1545 vdd.n1544 0.388379
R20583 vdd.n1511 vdd.n1509 0.388379
R20584 vdd.n1604 vdd.n1603 0.388379
R20585 vdd.n1570 vdd.n1568 0.388379
R20586 vdd.n19 vdd.n17 0.387128
R20587 vdd.n24 vdd.n22 0.387128
R20588 vdd.n6 vdd.n4 0.358259
R20589 vdd.n13 vdd.n11 0.358259
R20590 vdd.n276 vdd.n274 0.358259
R20591 vdd.n278 vdd.n276 0.358259
R20592 vdd.n280 vdd.n278 0.358259
R20593 vdd.n282 vdd.n280 0.358259
R20594 vdd.n284 vdd.n282 0.358259
R20595 vdd.n286 vdd.n284 0.358259
R20596 vdd.n288 vdd.n286 0.358259
R20597 vdd.n290 vdd.n288 0.358259
R20598 vdd.n332 vdd.n290 0.358259
R20599 vdd.n174 vdd.n172 0.358259
R20600 vdd.n176 vdd.n174 0.358259
R20601 vdd.n178 vdd.n176 0.358259
R20602 vdd.n180 vdd.n178 0.358259
R20603 vdd.n182 vdd.n180 0.358259
R20604 vdd.n184 vdd.n182 0.358259
R20605 vdd.n186 vdd.n184 0.358259
R20606 vdd.n188 vdd.n186 0.358259
R20607 vdd.n230 vdd.n188 0.358259
R20608 vdd.n73 vdd.n71 0.358259
R20609 vdd.n75 vdd.n73 0.358259
R20610 vdd.n77 vdd.n75 0.358259
R20611 vdd.n79 vdd.n77 0.358259
R20612 vdd.n81 vdd.n79 0.358259
R20613 vdd.n83 vdd.n81 0.358259
R20614 vdd.n85 vdd.n83 0.358259
R20615 vdd.n87 vdd.n85 0.358259
R20616 vdd.n129 vdd.n87 0.358259
R20617 vdd.n1810 vdd.n1768 0.358259
R20618 vdd.n1768 vdd.n1766 0.358259
R20619 vdd.n1766 vdd.n1764 0.358259
R20620 vdd.n1764 vdd.n1762 0.358259
R20621 vdd.n1762 vdd.n1760 0.358259
R20622 vdd.n1760 vdd.n1758 0.358259
R20623 vdd.n1758 vdd.n1756 0.358259
R20624 vdd.n1756 vdd.n1754 0.358259
R20625 vdd.n1754 vdd.n1752 0.358259
R20626 vdd.n1708 vdd.n1666 0.358259
R20627 vdd.n1666 vdd.n1664 0.358259
R20628 vdd.n1664 vdd.n1662 0.358259
R20629 vdd.n1662 vdd.n1660 0.358259
R20630 vdd.n1660 vdd.n1658 0.358259
R20631 vdd.n1658 vdd.n1656 0.358259
R20632 vdd.n1656 vdd.n1654 0.358259
R20633 vdd.n1654 vdd.n1652 0.358259
R20634 vdd.n1652 vdd.n1650 0.358259
R20635 vdd.n1607 vdd.n1565 0.358259
R20636 vdd.n1565 vdd.n1563 0.358259
R20637 vdd.n1563 vdd.n1561 0.358259
R20638 vdd.n1561 vdd.n1559 0.358259
R20639 vdd.n1559 vdd.n1557 0.358259
R20640 vdd.n1557 vdd.n1555 0.358259
R20641 vdd.n1555 vdd.n1553 0.358259
R20642 vdd.n1553 vdd.n1551 0.358259
R20643 vdd.n1551 vdd.n1549 0.358259
R20644 vdd.n14 vdd.n6 0.334552
R20645 vdd.n14 vdd.n13 0.334552
R20646 vdd.n27 vdd.n19 0.21707
R20647 vdd.n27 vdd.n24 0.21707
R20648 vdd.n330 vdd.n292 0.155672
R20649 vdd.n322 vdd.n292 0.155672
R20650 vdd.n322 vdd.n321 0.155672
R20651 vdd.n321 vdd.n297 0.155672
R20652 vdd.n314 vdd.n297 0.155672
R20653 vdd.n314 vdd.n313 0.155672
R20654 vdd.n313 vdd.n301 0.155672
R20655 vdd.n306 vdd.n301 0.155672
R20656 vdd.n271 vdd.n233 0.155672
R20657 vdd.n263 vdd.n233 0.155672
R20658 vdd.n263 vdd.n262 0.155672
R20659 vdd.n262 vdd.n238 0.155672
R20660 vdd.n255 vdd.n238 0.155672
R20661 vdd.n255 vdd.n254 0.155672
R20662 vdd.n254 vdd.n242 0.155672
R20663 vdd.n247 vdd.n242 0.155672
R20664 vdd.n228 vdd.n190 0.155672
R20665 vdd.n220 vdd.n190 0.155672
R20666 vdd.n220 vdd.n219 0.155672
R20667 vdd.n219 vdd.n195 0.155672
R20668 vdd.n212 vdd.n195 0.155672
R20669 vdd.n212 vdd.n211 0.155672
R20670 vdd.n211 vdd.n199 0.155672
R20671 vdd.n204 vdd.n199 0.155672
R20672 vdd.n169 vdd.n131 0.155672
R20673 vdd.n161 vdd.n131 0.155672
R20674 vdd.n161 vdd.n160 0.155672
R20675 vdd.n160 vdd.n136 0.155672
R20676 vdd.n153 vdd.n136 0.155672
R20677 vdd.n153 vdd.n152 0.155672
R20678 vdd.n152 vdd.n140 0.155672
R20679 vdd.n145 vdd.n140 0.155672
R20680 vdd.n127 vdd.n89 0.155672
R20681 vdd.n119 vdd.n89 0.155672
R20682 vdd.n119 vdd.n118 0.155672
R20683 vdd.n118 vdd.n94 0.155672
R20684 vdd.n111 vdd.n94 0.155672
R20685 vdd.n111 vdd.n110 0.155672
R20686 vdd.n110 vdd.n98 0.155672
R20687 vdd.n103 vdd.n98 0.155672
R20688 vdd.n68 vdd.n30 0.155672
R20689 vdd.n60 vdd.n30 0.155672
R20690 vdd.n60 vdd.n59 0.155672
R20691 vdd.n59 vdd.n35 0.155672
R20692 vdd.n52 vdd.n35 0.155672
R20693 vdd.n52 vdd.n51 0.155672
R20694 vdd.n51 vdd.n39 0.155672
R20695 vdd.n44 vdd.n39 0.155672
R20696 vdd.n1749 vdd.n1711 0.155672
R20697 vdd.n1741 vdd.n1711 0.155672
R20698 vdd.n1741 vdd.n1740 0.155672
R20699 vdd.n1740 vdd.n1716 0.155672
R20700 vdd.n1733 vdd.n1716 0.155672
R20701 vdd.n1733 vdd.n1732 0.155672
R20702 vdd.n1732 vdd.n1720 0.155672
R20703 vdd.n1725 vdd.n1720 0.155672
R20704 vdd.n1808 vdd.n1770 0.155672
R20705 vdd.n1800 vdd.n1770 0.155672
R20706 vdd.n1800 vdd.n1799 0.155672
R20707 vdd.n1799 vdd.n1775 0.155672
R20708 vdd.n1792 vdd.n1775 0.155672
R20709 vdd.n1792 vdd.n1791 0.155672
R20710 vdd.n1791 vdd.n1779 0.155672
R20711 vdd.n1784 vdd.n1779 0.155672
R20712 vdd.n1647 vdd.n1609 0.155672
R20713 vdd.n1639 vdd.n1609 0.155672
R20714 vdd.n1639 vdd.n1638 0.155672
R20715 vdd.n1638 vdd.n1614 0.155672
R20716 vdd.n1631 vdd.n1614 0.155672
R20717 vdd.n1631 vdd.n1630 0.155672
R20718 vdd.n1630 vdd.n1618 0.155672
R20719 vdd.n1623 vdd.n1618 0.155672
R20720 vdd.n1706 vdd.n1668 0.155672
R20721 vdd.n1698 vdd.n1668 0.155672
R20722 vdd.n1698 vdd.n1697 0.155672
R20723 vdd.n1697 vdd.n1673 0.155672
R20724 vdd.n1690 vdd.n1673 0.155672
R20725 vdd.n1690 vdd.n1689 0.155672
R20726 vdd.n1689 vdd.n1677 0.155672
R20727 vdd.n1682 vdd.n1677 0.155672
R20728 vdd.n1546 vdd.n1508 0.155672
R20729 vdd.n1538 vdd.n1508 0.155672
R20730 vdd.n1538 vdd.n1537 0.155672
R20731 vdd.n1537 vdd.n1513 0.155672
R20732 vdd.n1530 vdd.n1513 0.155672
R20733 vdd.n1530 vdd.n1529 0.155672
R20734 vdd.n1529 vdd.n1517 0.155672
R20735 vdd.n1522 vdd.n1517 0.155672
R20736 vdd.n1605 vdd.n1567 0.155672
R20737 vdd.n1597 vdd.n1567 0.155672
R20738 vdd.n1597 vdd.n1596 0.155672
R20739 vdd.n1596 vdd.n1572 0.155672
R20740 vdd.n1589 vdd.n1572 0.155672
R20741 vdd.n1589 vdd.n1588 0.155672
R20742 vdd.n1588 vdd.n1576 0.155672
R20743 vdd.n1581 vdd.n1576 0.155672
R20744 vdd.n2101 vdd.n1906 0.152939
R20745 vdd.n1912 vdd.n1906 0.152939
R20746 vdd.n1913 vdd.n1912 0.152939
R20747 vdd.n1914 vdd.n1913 0.152939
R20748 vdd.n1915 vdd.n1914 0.152939
R20749 vdd.n1919 vdd.n1915 0.152939
R20750 vdd.n1920 vdd.n1919 0.152939
R20751 vdd.n1921 vdd.n1920 0.152939
R20752 vdd.n1922 vdd.n1921 0.152939
R20753 vdd.n1926 vdd.n1922 0.152939
R20754 vdd.n1927 vdd.n1926 0.152939
R20755 vdd.n1928 vdd.n1927 0.152939
R20756 vdd.n2076 vdd.n1928 0.152939
R20757 vdd.n2076 vdd.n2075 0.152939
R20758 vdd.n2075 vdd.n2074 0.152939
R20759 vdd.n2074 vdd.n1934 0.152939
R20760 vdd.n1939 vdd.n1934 0.152939
R20761 vdd.n1940 vdd.n1939 0.152939
R20762 vdd.n1941 vdd.n1940 0.152939
R20763 vdd.n1945 vdd.n1941 0.152939
R20764 vdd.n1946 vdd.n1945 0.152939
R20765 vdd.n1947 vdd.n1946 0.152939
R20766 vdd.n1948 vdd.n1947 0.152939
R20767 vdd.n1952 vdd.n1948 0.152939
R20768 vdd.n1953 vdd.n1952 0.152939
R20769 vdd.n1954 vdd.n1953 0.152939
R20770 vdd.n1955 vdd.n1954 0.152939
R20771 vdd.n1959 vdd.n1955 0.152939
R20772 vdd.n1960 vdd.n1959 0.152939
R20773 vdd.n1961 vdd.n1960 0.152939
R20774 vdd.n1962 vdd.n1961 0.152939
R20775 vdd.n1966 vdd.n1962 0.152939
R20776 vdd.n1967 vdd.n1966 0.152939
R20777 vdd.n1968 vdd.n1967 0.152939
R20778 vdd.n2037 vdd.n1968 0.152939
R20779 vdd.n2037 vdd.n2036 0.152939
R20780 vdd.n2036 vdd.n2035 0.152939
R20781 vdd.n2035 vdd.n1974 0.152939
R20782 vdd.n1979 vdd.n1974 0.152939
R20783 vdd.n1980 vdd.n1979 0.152939
R20784 vdd.n1981 vdd.n1980 0.152939
R20785 vdd.n1985 vdd.n1981 0.152939
R20786 vdd.n1986 vdd.n1985 0.152939
R20787 vdd.n1987 vdd.n1986 0.152939
R20788 vdd.n1988 vdd.n1987 0.152939
R20789 vdd.n1992 vdd.n1988 0.152939
R20790 vdd.n1993 vdd.n1992 0.152939
R20791 vdd.n1994 vdd.n1993 0.152939
R20792 vdd.n1995 vdd.n1994 0.152939
R20793 vdd.n1996 vdd.n1995 0.152939
R20794 vdd.n1996 vdd.n1064 0.152939
R20795 vdd.n2325 vdd.n1900 0.152939
R20796 vdd.n1814 vdd.n1123 0.152939
R20797 vdd.n1829 vdd.n1123 0.152939
R20798 vdd.n1830 vdd.n1829 0.152939
R20799 vdd.n1831 vdd.n1830 0.152939
R20800 vdd.n1831 vdd.n1112 0.152939
R20801 vdd.n1846 vdd.n1112 0.152939
R20802 vdd.n1847 vdd.n1846 0.152939
R20803 vdd.n1848 vdd.n1847 0.152939
R20804 vdd.n1848 vdd.n1101 0.152939
R20805 vdd.n1862 vdd.n1101 0.152939
R20806 vdd.n1863 vdd.n1862 0.152939
R20807 vdd.n1864 vdd.n1863 0.152939
R20808 vdd.n1864 vdd.n1089 0.152939
R20809 vdd.n1879 vdd.n1089 0.152939
R20810 vdd.n1880 vdd.n1879 0.152939
R20811 vdd.n1881 vdd.n1880 0.152939
R20812 vdd.n1881 vdd.n1077 0.152939
R20813 vdd.n1898 vdd.n1077 0.152939
R20814 vdd.n1899 vdd.n1898 0.152939
R20815 vdd.n2326 vdd.n1899 0.152939
R20816 vdd.n735 vdd.n730 0.152939
R20817 vdd.n736 vdd.n735 0.152939
R20818 vdd.n737 vdd.n736 0.152939
R20819 vdd.n738 vdd.n737 0.152939
R20820 vdd.n739 vdd.n738 0.152939
R20821 vdd.n740 vdd.n739 0.152939
R20822 vdd.n741 vdd.n740 0.152939
R20823 vdd.n742 vdd.n741 0.152939
R20824 vdd.n743 vdd.n742 0.152939
R20825 vdd.n744 vdd.n743 0.152939
R20826 vdd.n745 vdd.n744 0.152939
R20827 vdd.n746 vdd.n745 0.152939
R20828 vdd.n3183 vdd.n746 0.152939
R20829 vdd.n3183 vdd.n3182 0.152939
R20830 vdd.n3182 vdd.n3181 0.152939
R20831 vdd.n3181 vdd.n748 0.152939
R20832 vdd.n749 vdd.n748 0.152939
R20833 vdd.n750 vdd.n749 0.152939
R20834 vdd.n751 vdd.n750 0.152939
R20835 vdd.n752 vdd.n751 0.152939
R20836 vdd.n753 vdd.n752 0.152939
R20837 vdd.n754 vdd.n753 0.152939
R20838 vdd.n755 vdd.n754 0.152939
R20839 vdd.n756 vdd.n755 0.152939
R20840 vdd.n757 vdd.n756 0.152939
R20841 vdd.n758 vdd.n757 0.152939
R20842 vdd.n759 vdd.n758 0.152939
R20843 vdd.n760 vdd.n759 0.152939
R20844 vdd.n761 vdd.n760 0.152939
R20845 vdd.n762 vdd.n761 0.152939
R20846 vdd.n763 vdd.n762 0.152939
R20847 vdd.n764 vdd.n763 0.152939
R20848 vdd.n765 vdd.n764 0.152939
R20849 vdd.n766 vdd.n765 0.152939
R20850 vdd.n3137 vdd.n766 0.152939
R20851 vdd.n3137 vdd.n3136 0.152939
R20852 vdd.n3136 vdd.n3135 0.152939
R20853 vdd.n3135 vdd.n770 0.152939
R20854 vdd.n771 vdd.n770 0.152939
R20855 vdd.n772 vdd.n771 0.152939
R20856 vdd.n773 vdd.n772 0.152939
R20857 vdd.n774 vdd.n773 0.152939
R20858 vdd.n775 vdd.n774 0.152939
R20859 vdd.n776 vdd.n775 0.152939
R20860 vdd.n777 vdd.n776 0.152939
R20861 vdd.n778 vdd.n777 0.152939
R20862 vdd.n779 vdd.n778 0.152939
R20863 vdd.n780 vdd.n779 0.152939
R20864 vdd.n781 vdd.n780 0.152939
R20865 vdd.n782 vdd.n781 0.152939
R20866 vdd.n783 vdd.n782 0.152939
R20867 vdd.n727 vdd.n726 0.152939
R20868 vdd.n3234 vdd.n682 0.152939
R20869 vdd.n3235 vdd.n3234 0.152939
R20870 vdd.n3236 vdd.n3235 0.152939
R20871 vdd.n3236 vdd.n670 0.152939
R20872 vdd.n3251 vdd.n670 0.152939
R20873 vdd.n3252 vdd.n3251 0.152939
R20874 vdd.n3253 vdd.n3252 0.152939
R20875 vdd.n3253 vdd.n659 0.152939
R20876 vdd.n3267 vdd.n659 0.152939
R20877 vdd.n3268 vdd.n3267 0.152939
R20878 vdd.n3269 vdd.n3268 0.152939
R20879 vdd.n3269 vdd.n647 0.152939
R20880 vdd.n3284 vdd.n647 0.152939
R20881 vdd.n3285 vdd.n3284 0.152939
R20882 vdd.n3286 vdd.n3285 0.152939
R20883 vdd.n3286 vdd.n636 0.152939
R20884 vdd.n3303 vdd.n636 0.152939
R20885 vdd.n3304 vdd.n3303 0.152939
R20886 vdd.n3305 vdd.n3304 0.152939
R20887 vdd.n3305 vdd.n334 0.152939
R20888 vdd.n3398 vdd.n335 0.152939
R20889 vdd.n346 vdd.n335 0.152939
R20890 vdd.n347 vdd.n346 0.152939
R20891 vdd.n348 vdd.n347 0.152939
R20892 vdd.n355 vdd.n348 0.152939
R20893 vdd.n356 vdd.n355 0.152939
R20894 vdd.n357 vdd.n356 0.152939
R20895 vdd.n358 vdd.n357 0.152939
R20896 vdd.n366 vdd.n358 0.152939
R20897 vdd.n367 vdd.n366 0.152939
R20898 vdd.n368 vdd.n367 0.152939
R20899 vdd.n369 vdd.n368 0.152939
R20900 vdd.n377 vdd.n369 0.152939
R20901 vdd.n378 vdd.n377 0.152939
R20902 vdd.n379 vdd.n378 0.152939
R20903 vdd.n380 vdd.n379 0.152939
R20904 vdd.n388 vdd.n380 0.152939
R20905 vdd.n389 vdd.n388 0.152939
R20906 vdd.n390 vdd.n389 0.152939
R20907 vdd.n391 vdd.n390 0.152939
R20908 vdd.n464 vdd.n463 0.152939
R20909 vdd.n470 vdd.n463 0.152939
R20910 vdd.n471 vdd.n470 0.152939
R20911 vdd.n472 vdd.n471 0.152939
R20912 vdd.n472 vdd.n461 0.152939
R20913 vdd.n480 vdd.n461 0.152939
R20914 vdd.n481 vdd.n480 0.152939
R20915 vdd.n482 vdd.n481 0.152939
R20916 vdd.n482 vdd.n459 0.152939
R20917 vdd.n490 vdd.n459 0.152939
R20918 vdd.n491 vdd.n490 0.152939
R20919 vdd.n492 vdd.n491 0.152939
R20920 vdd.n492 vdd.n457 0.152939
R20921 vdd.n500 vdd.n457 0.152939
R20922 vdd.n501 vdd.n500 0.152939
R20923 vdd.n502 vdd.n501 0.152939
R20924 vdd.n502 vdd.n455 0.152939
R20925 vdd.n510 vdd.n455 0.152939
R20926 vdd.n511 vdd.n510 0.152939
R20927 vdd.n512 vdd.n511 0.152939
R20928 vdd.n512 vdd.n451 0.152939
R20929 vdd.n520 vdd.n451 0.152939
R20930 vdd.n521 vdd.n520 0.152939
R20931 vdd.n522 vdd.n521 0.152939
R20932 vdd.n522 vdd.n449 0.152939
R20933 vdd.n530 vdd.n449 0.152939
R20934 vdd.n531 vdd.n530 0.152939
R20935 vdd.n532 vdd.n531 0.152939
R20936 vdd.n532 vdd.n447 0.152939
R20937 vdd.n540 vdd.n447 0.152939
R20938 vdd.n541 vdd.n540 0.152939
R20939 vdd.n542 vdd.n541 0.152939
R20940 vdd.n542 vdd.n445 0.152939
R20941 vdd.n550 vdd.n445 0.152939
R20942 vdd.n551 vdd.n550 0.152939
R20943 vdd.n552 vdd.n551 0.152939
R20944 vdd.n552 vdd.n443 0.152939
R20945 vdd.n560 vdd.n443 0.152939
R20946 vdd.n561 vdd.n560 0.152939
R20947 vdd.n562 vdd.n561 0.152939
R20948 vdd.n562 vdd.n439 0.152939
R20949 vdd.n570 vdd.n439 0.152939
R20950 vdd.n571 vdd.n570 0.152939
R20951 vdd.n572 vdd.n571 0.152939
R20952 vdd.n572 vdd.n437 0.152939
R20953 vdd.n580 vdd.n437 0.152939
R20954 vdd.n581 vdd.n580 0.152939
R20955 vdd.n582 vdd.n581 0.152939
R20956 vdd.n582 vdd.n435 0.152939
R20957 vdd.n590 vdd.n435 0.152939
R20958 vdd.n591 vdd.n590 0.152939
R20959 vdd.n592 vdd.n591 0.152939
R20960 vdd.n592 vdd.n433 0.152939
R20961 vdd.n600 vdd.n433 0.152939
R20962 vdd.n601 vdd.n600 0.152939
R20963 vdd.n602 vdd.n601 0.152939
R20964 vdd.n602 vdd.n431 0.152939
R20965 vdd.n610 vdd.n431 0.152939
R20966 vdd.n611 vdd.n610 0.152939
R20967 vdd.n612 vdd.n611 0.152939
R20968 vdd.n612 vdd.n429 0.152939
R20969 vdd.n619 vdd.n429 0.152939
R20970 vdd.n3350 vdd.n619 0.152939
R20971 vdd.n3228 vdd.n3227 0.152939
R20972 vdd.n3228 vdd.n675 0.152939
R20973 vdd.n3242 vdd.n675 0.152939
R20974 vdd.n3243 vdd.n3242 0.152939
R20975 vdd.n3244 vdd.n3243 0.152939
R20976 vdd.n3244 vdd.n665 0.152939
R20977 vdd.n3259 vdd.n665 0.152939
R20978 vdd.n3260 vdd.n3259 0.152939
R20979 vdd.n3261 vdd.n3260 0.152939
R20980 vdd.n3261 vdd.n652 0.152939
R20981 vdd.n3275 vdd.n652 0.152939
R20982 vdd.n3276 vdd.n3275 0.152939
R20983 vdd.n3277 vdd.n3276 0.152939
R20984 vdd.n3277 vdd.n641 0.152939
R20985 vdd.n3292 vdd.n641 0.152939
R20986 vdd.n3293 vdd.n3292 0.152939
R20987 vdd.n3294 vdd.n3293 0.152939
R20988 vdd.n3296 vdd.n3294 0.152939
R20989 vdd.n3296 vdd.n3295 0.152939
R20990 vdd.n3295 vdd.n630 0.152939
R20991 vdd.n3313 vdd.n630 0.152939
R20992 vdd.n3314 vdd.n3313 0.152939
R20993 vdd.n3315 vdd.n3314 0.152939
R20994 vdd.n3315 vdd.n628 0.152939
R20995 vdd.n3320 vdd.n628 0.152939
R20996 vdd.n3321 vdd.n3320 0.152939
R20997 vdd.n3322 vdd.n3321 0.152939
R20998 vdd.n3322 vdd.n626 0.152939
R20999 vdd.n3327 vdd.n626 0.152939
R21000 vdd.n3328 vdd.n3327 0.152939
R21001 vdd.n3329 vdd.n3328 0.152939
R21002 vdd.n3329 vdd.n624 0.152939
R21003 vdd.n3335 vdd.n624 0.152939
R21004 vdd.n3336 vdd.n3335 0.152939
R21005 vdd.n3337 vdd.n3336 0.152939
R21006 vdd.n3337 vdd.n622 0.152939
R21007 vdd.n3342 vdd.n622 0.152939
R21008 vdd.n3343 vdd.n3342 0.152939
R21009 vdd.n3344 vdd.n3343 0.152939
R21010 vdd.n3344 vdd.n620 0.152939
R21011 vdd.n3349 vdd.n620 0.152939
R21012 vdd.n3226 vdd.n687 0.152939
R21013 vdd.n2337 vdd.n1067 0.152939
R21014 vdd.n1430 vdd.n1186 0.152939
R21015 vdd.n1431 vdd.n1430 0.152939
R21016 vdd.n1432 vdd.n1431 0.152939
R21017 vdd.n1432 vdd.n1174 0.152939
R21018 vdd.n1447 vdd.n1174 0.152939
R21019 vdd.n1448 vdd.n1447 0.152939
R21020 vdd.n1449 vdd.n1448 0.152939
R21021 vdd.n1449 vdd.n1164 0.152939
R21022 vdd.n1464 vdd.n1164 0.152939
R21023 vdd.n1465 vdd.n1464 0.152939
R21024 vdd.n1466 vdd.n1465 0.152939
R21025 vdd.n1466 vdd.n1151 0.152939
R21026 vdd.n1480 vdd.n1151 0.152939
R21027 vdd.n1481 vdd.n1480 0.152939
R21028 vdd.n1482 vdd.n1481 0.152939
R21029 vdd.n1482 vdd.n1140 0.152939
R21030 vdd.n1497 vdd.n1140 0.152939
R21031 vdd.n1498 vdd.n1497 0.152939
R21032 vdd.n1499 vdd.n1498 0.152939
R21033 vdd.n1499 vdd.n1129 0.152939
R21034 vdd.n1820 vdd.n1129 0.152939
R21035 vdd.n1821 vdd.n1820 0.152939
R21036 vdd.n1822 vdd.n1821 0.152939
R21037 vdd.n1822 vdd.n1117 0.152939
R21038 vdd.n1837 vdd.n1117 0.152939
R21039 vdd.n1838 vdd.n1837 0.152939
R21040 vdd.n1839 vdd.n1838 0.152939
R21041 vdd.n1839 vdd.n1107 0.152939
R21042 vdd.n1854 vdd.n1107 0.152939
R21043 vdd.n1855 vdd.n1854 0.152939
R21044 vdd.n1856 vdd.n1855 0.152939
R21045 vdd.n1856 vdd.n1094 0.152939
R21046 vdd.n1870 vdd.n1094 0.152939
R21047 vdd.n1871 vdd.n1870 0.152939
R21048 vdd.n1872 vdd.n1871 0.152939
R21049 vdd.n1872 vdd.n1084 0.152939
R21050 vdd.n1887 vdd.n1084 0.152939
R21051 vdd.n1888 vdd.n1887 0.152939
R21052 vdd.n1891 vdd.n1888 0.152939
R21053 vdd.n1891 vdd.n1890 0.152939
R21054 vdd.n1890 vdd.n1889 0.152939
R21055 vdd.n1422 vdd.n1191 0.152939
R21056 vdd.n1415 vdd.n1191 0.152939
R21057 vdd.n1415 vdd.n1414 0.152939
R21058 vdd.n1414 vdd.n1413 0.152939
R21059 vdd.n1413 vdd.n1228 0.152939
R21060 vdd.n1409 vdd.n1228 0.152939
R21061 vdd.n1409 vdd.n1408 0.152939
R21062 vdd.n1408 vdd.n1407 0.152939
R21063 vdd.n1407 vdd.n1234 0.152939
R21064 vdd.n1403 vdd.n1234 0.152939
R21065 vdd.n1403 vdd.n1402 0.152939
R21066 vdd.n1402 vdd.n1401 0.152939
R21067 vdd.n1401 vdd.n1240 0.152939
R21068 vdd.n1397 vdd.n1240 0.152939
R21069 vdd.n1397 vdd.n1396 0.152939
R21070 vdd.n1396 vdd.n1395 0.152939
R21071 vdd.n1395 vdd.n1246 0.152939
R21072 vdd.n1391 vdd.n1246 0.152939
R21073 vdd.n1391 vdd.n1390 0.152939
R21074 vdd.n1390 vdd.n1389 0.152939
R21075 vdd.n1389 vdd.n1254 0.152939
R21076 vdd.n1385 vdd.n1254 0.152939
R21077 vdd.n1385 vdd.n1384 0.152939
R21078 vdd.n1384 vdd.n1383 0.152939
R21079 vdd.n1383 vdd.n1260 0.152939
R21080 vdd.n1379 vdd.n1260 0.152939
R21081 vdd.n1379 vdd.n1378 0.152939
R21082 vdd.n1378 vdd.n1377 0.152939
R21083 vdd.n1377 vdd.n1266 0.152939
R21084 vdd.n1373 vdd.n1266 0.152939
R21085 vdd.n1373 vdd.n1372 0.152939
R21086 vdd.n1372 vdd.n1371 0.152939
R21087 vdd.n1371 vdd.n1272 0.152939
R21088 vdd.n1367 vdd.n1272 0.152939
R21089 vdd.n1367 vdd.n1366 0.152939
R21090 vdd.n1366 vdd.n1365 0.152939
R21091 vdd.n1365 vdd.n1278 0.152939
R21092 vdd.n1361 vdd.n1278 0.152939
R21093 vdd.n1361 vdd.n1360 0.152939
R21094 vdd.n1360 vdd.n1359 0.152939
R21095 vdd.n1359 vdd.n1284 0.152939
R21096 vdd.n1352 vdd.n1284 0.152939
R21097 vdd.n1352 vdd.n1351 0.152939
R21098 vdd.n1351 vdd.n1350 0.152939
R21099 vdd.n1350 vdd.n1289 0.152939
R21100 vdd.n1346 vdd.n1289 0.152939
R21101 vdd.n1346 vdd.n1345 0.152939
R21102 vdd.n1345 vdd.n1344 0.152939
R21103 vdd.n1344 vdd.n1295 0.152939
R21104 vdd.n1340 vdd.n1295 0.152939
R21105 vdd.n1340 vdd.n1339 0.152939
R21106 vdd.n1339 vdd.n1338 0.152939
R21107 vdd.n1338 vdd.n1301 0.152939
R21108 vdd.n1334 vdd.n1301 0.152939
R21109 vdd.n1334 vdd.n1333 0.152939
R21110 vdd.n1333 vdd.n1332 0.152939
R21111 vdd.n1332 vdd.n1307 0.152939
R21112 vdd.n1328 vdd.n1307 0.152939
R21113 vdd.n1328 vdd.n1327 0.152939
R21114 vdd.n1327 vdd.n1326 0.152939
R21115 vdd.n1326 vdd.n1313 0.152939
R21116 vdd.n1322 vdd.n1313 0.152939
R21117 vdd.n1322 vdd.n1321 0.152939
R21118 vdd.n1424 vdd.n1423 0.152939
R21119 vdd.n1424 vdd.n1180 0.152939
R21120 vdd.n1439 vdd.n1180 0.152939
R21121 vdd.n1440 vdd.n1439 0.152939
R21122 vdd.n1441 vdd.n1440 0.152939
R21123 vdd.n1441 vdd.n1169 0.152939
R21124 vdd.n1456 vdd.n1169 0.152939
R21125 vdd.n1457 vdd.n1456 0.152939
R21126 vdd.n1458 vdd.n1457 0.152939
R21127 vdd.n1458 vdd.n1158 0.152939
R21128 vdd.n1472 vdd.n1158 0.152939
R21129 vdd.n1473 vdd.n1472 0.152939
R21130 vdd.n1474 vdd.n1473 0.152939
R21131 vdd.n1474 vdd.n1146 0.152939
R21132 vdd.n1489 vdd.n1146 0.152939
R21133 vdd.n1490 vdd.n1489 0.152939
R21134 vdd.n1491 vdd.n1490 0.152939
R21135 vdd.n1491 vdd.n1135 0.152939
R21136 vdd.n1505 vdd.n1135 0.152939
R21137 vdd.n1506 vdd.n1505 0.152939
R21138 vdd.n1427 vdd.t50 0.113865
R21139 vdd.t57 vdd.n386 0.113865
R21140 vdd.n2315 vdd.n1900 0.110256
R21141 vdd.n3216 vdd.n727 0.110256
R21142 vdd.n3093 vdd.n687 0.110256
R21143 vdd.n2338 vdd.n2337 0.110256
R21144 vdd.n1814 vdd.n1813 0.0695946
R21145 vdd.n3399 vdd.n334 0.0695946
R21146 vdd.n3399 vdd.n3398 0.0695946
R21147 vdd.n1813 vdd.n1506 0.0695946
R21148 vdd.n2315 vdd.n2101 0.0431829
R21149 vdd.n2338 vdd.n1064 0.0431829
R21150 vdd.n3216 vdd.n730 0.0431829
R21151 vdd.n3093 vdd.n783 0.0431829
R21152 vdd vdd.n28 0.00833333
R21153 a_n2848_n452.n5 a_n2848_n452.t75 539.01
R21154 a_n2848_n452.n97 a_n2848_n452.t58 512.366
R21155 a_n2848_n452.n96 a_n2848_n452.t62 512.366
R21156 a_n2848_n452.n70 a_n2848_n452.t52 512.366
R21157 a_n2848_n452.n95 a_n2848_n452.t67 512.366
R21158 a_n2848_n452.n1 a_n2848_n452.t37 533.058
R21159 a_n2848_n452.n101 a_n2848_n452.t41 512.366
R21160 a_n2848_n452.n100 a_n2848_n452.t25 512.366
R21161 a_n2848_n452.n69 a_n2848_n452.t43 512.366
R21162 a_n2848_n452.n98 a_n2848_n452.t33 512.366
R21163 a_n2848_n452.n19 a_n2848_n452.t35 539.01
R21164 a_n2848_n452.n78 a_n2848_n452.t27 512.366
R21165 a_n2848_n452.n79 a_n2848_n452.t23 512.366
R21166 a_n2848_n452.n73 a_n2848_n452.t31 512.366
R21167 a_n2848_n452.n80 a_n2848_n452.t39 512.366
R21168 a_n2848_n452.n23 a_n2848_n452.t70 539.01
R21169 a_n2848_n452.n75 a_n2848_n452.t71 512.366
R21170 a_n2848_n452.n76 a_n2848_n452.t50 512.366
R21171 a_n2848_n452.n74 a_n2848_n452.t56 512.366
R21172 a_n2848_n452.n77 a_n2848_n452.t65 512.366
R21173 a_n2848_n452.n92 a_n2848_n452.t64 512.366
R21174 a_n2848_n452.n82 a_n2848_n452.t55 512.366
R21175 a_n2848_n452.n93 a_n2848_n452.t49 512.366
R21176 a_n2848_n452.n90 a_n2848_n452.t72 512.366
R21177 a_n2848_n452.n83 a_n2848_n452.t61 512.366
R21178 a_n2848_n452.n91 a_n2848_n452.t60 512.366
R21179 a_n2848_n452.n88 a_n2848_n452.t68 512.366
R21180 a_n2848_n452.n84 a_n2848_n452.t53 512.366
R21181 a_n2848_n452.n89 a_n2848_n452.t54 512.366
R21182 a_n2848_n452.n86 a_n2848_n452.t57 512.366
R21183 a_n2848_n452.n85 a_n2848_n452.t66 512.366
R21184 a_n2848_n452.n87 a_n2848_n452.t48 512.366
R21185 a_n2848_n452.n50 a_n2848_n452.n3 70.3058
R21186 a_n2848_n452.n47 a_n2848_n452.n6 70.3058
R21187 a_n2848_n452.n16 a_n2848_n452.n37 70.3058
R21188 a_n2848_n452.n20 a_n2848_n452.n34 70.3058
R21189 a_n2848_n452.n33 a_n2848_n452.n21 70.1674
R21190 a_n2848_n452.n33 a_n2848_n452.n74 20.9683
R21191 a_n2848_n452.n21 a_n2848_n452.n32 75.0448
R21192 a_n2848_n452.n76 a_n2848_n452.n32 11.2134
R21193 a_n2848_n452.n22 a_n2848_n452.n23 44.8194
R21194 a_n2848_n452.n36 a_n2848_n452.n17 70.1674
R21195 a_n2848_n452.n36 a_n2848_n452.n73 20.9683
R21196 a_n2848_n452.n17 a_n2848_n452.n35 75.0448
R21197 a_n2848_n452.n79 a_n2848_n452.n35 11.2134
R21198 a_n2848_n452.n18 a_n2848_n452.n19 44.8194
R21199 a_n2848_n452.n7 a_n2848_n452.n45 70.1674
R21200 a_n2848_n452.n9 a_n2848_n452.n43 70.1674
R21201 a_n2848_n452.n11 a_n2848_n452.n41 70.1674
R21202 a_n2848_n452.n14 a_n2848_n452.n39 70.1674
R21203 a_n2848_n452.n87 a_n2848_n452.n39 20.9683
R21204 a_n2848_n452.n38 a_n2848_n452.n15 75.0448
R21205 a_n2848_n452.n38 a_n2848_n452.n85 11.2134
R21206 a_n2848_n452.n15 a_n2848_n452.n86 161.3
R21207 a_n2848_n452.n89 a_n2848_n452.n41 20.9683
R21208 a_n2848_n452.n40 a_n2848_n452.n12 75.0448
R21209 a_n2848_n452.n40 a_n2848_n452.n84 11.2134
R21210 a_n2848_n452.n12 a_n2848_n452.n88 161.3
R21211 a_n2848_n452.n91 a_n2848_n452.n43 20.9683
R21212 a_n2848_n452.n42 a_n2848_n452.n10 75.0448
R21213 a_n2848_n452.n42 a_n2848_n452.n83 11.2134
R21214 a_n2848_n452.n10 a_n2848_n452.n90 161.3
R21215 a_n2848_n452.n93 a_n2848_n452.n45 20.9683
R21216 a_n2848_n452.n44 a_n2848_n452.n8 75.0448
R21217 a_n2848_n452.n44 a_n2848_n452.n82 11.2134
R21218 a_n2848_n452.n8 a_n2848_n452.n92 161.3
R21219 a_n2848_n452.n6 a_n2848_n452.n46 70.1674
R21220 a_n2848_n452.n46 a_n2848_n452.n69 20.9683
R21221 a_n2848_n452.n99 a_n2848_n452.n0 161.3
R21222 a_n2848_n452.n4 a_n2848_n452.n49 70.1674
R21223 a_n2848_n452.n49 a_n2848_n452.n70 20.9683
R21224 a_n2848_n452.n48 a_n2848_n452.n4 75.0448
R21225 a_n2848_n452.n96 a_n2848_n452.n48 11.2134
R21226 a_n2848_n452.n2 a_n2848_n452.n5 44.8194
R21227 a_n2848_n452.n100 a_n2848_n452.n51 20.9683
R21228 a_n2848_n452.n51 a_n2848_n452.n0 70.1674
R21229 a_n2848_n452.n0 a_n2848_n452.n1 70.3058
R21230 a_n2848_n452.n67 a_n2848_n452.n65 81.4626
R21231 a_n2848_n452.n58 a_n2848_n452.n56 81.4626
R21232 a_n2848_n452.n54 a_n2848_n452.n52 81.4626
R21233 a_n2848_n452.n67 a_n2848_n452.n66 80.9324
R21234 a_n2848_n452.n31 a_n2848_n452.n68 80.9324
R21235 a_n2848_n452.n30 a_n2848_n452.n64 80.9324
R21236 a_n2848_n452.n63 a_n2848_n452.n62 80.9324
R21237 a_n2848_n452.n61 a_n2848_n452.n60 80.9324
R21238 a_n2848_n452.n58 a_n2848_n452.n57 80.9324
R21239 a_n2848_n452.n29 a_n2848_n452.n59 80.9324
R21240 a_n2848_n452.n28 a_n2848_n452.n55 80.9324
R21241 a_n2848_n452.n54 a_n2848_n452.n53 80.9324
R21242 a_n2848_n452.n24 a_n2848_n452.t36 74.6477
R21243 a_n2848_n452.t22 a_n2848_n452.n27 74.6477
R21244 a_n2848_n452.n26 a_n2848_n452.t38 74.2899
R21245 a_n2848_n452.n25 a_n2848_n452.t30 74.2897
R21246 a_n2848_n452.n27 a_n2848_n452.n104 70.6783
R21247 a_n2848_n452.n27 a_n2848_n452.n103 70.6783
R21248 a_n2848_n452.n25 a_n2848_n452.n72 70.6783
R21249 a_n2848_n452.n24 a_n2848_n452.n71 70.6783
R21250 a_n2848_n452.n97 a_n2848_n452.n96 48.2005
R21251 a_n2848_n452.n95 a_n2848_n452.n49 20.9683
R21252 a_n2848_n452.n101 a_n2848_n452.n51 20.9683
R21253 a_n2848_n452.n98 a_n2848_n452.n46 20.9683
R21254 a_n2848_n452.n79 a_n2848_n452.n78 48.2005
R21255 a_n2848_n452.n80 a_n2848_n452.n36 20.9683
R21256 a_n2848_n452.n76 a_n2848_n452.n75 48.2005
R21257 a_n2848_n452.n77 a_n2848_n452.n33 20.9683
R21258 a_n2848_n452.n92 a_n2848_n452.n82 48.2005
R21259 a_n2848_n452.t69 a_n2848_n452.n45 533.335
R21260 a_n2848_n452.n90 a_n2848_n452.n83 48.2005
R21261 a_n2848_n452.t74 a_n2848_n452.n43 533.335
R21262 a_n2848_n452.n88 a_n2848_n452.n84 48.2005
R21263 a_n2848_n452.t63 a_n2848_n452.n41 533.335
R21264 a_n2848_n452.n86 a_n2848_n452.n85 48.2005
R21265 a_n2848_n452.t59 a_n2848_n452.n39 533.335
R21266 a_n2848_n452.n50 a_n2848_n452.t73 533.058
R21267 a_n2848_n452.n47 a_n2848_n452.t21 533.058
R21268 a_n2848_n452.t29 a_n2848_n452.n37 533.058
R21269 a_n2848_n452.t51 a_n2848_n452.n34 533.058
R21270 a_n2848_n452.n61 a_n2848_n452.n29 33.585
R21271 a_n2848_n452.n48 a_n2848_n452.n70 35.3134
R21272 a_n2848_n452.n100 a_n2848_n452.n99 24.1005
R21273 a_n2848_n452.n99 a_n2848_n452.n69 24.1005
R21274 a_n2848_n452.n73 a_n2848_n452.n35 35.3134
R21275 a_n2848_n452.n74 a_n2848_n452.n32 35.3134
R21276 a_n2848_n452.n93 a_n2848_n452.n44 35.3134
R21277 a_n2848_n452.n91 a_n2848_n452.n42 35.3134
R21278 a_n2848_n452.n89 a_n2848_n452.n40 35.3134
R21279 a_n2848_n452.n87 a_n2848_n452.n38 35.3134
R21280 a_n2848_n452.n0 a_n2848_n452.n31 23.891
R21281 a_n2848_n452.n22 a_n2848_n452.n13 12.046
R21282 a_n2848_n452.n3 a_n2848_n452.n94 11.8414
R21283 a_n2848_n452.n102 a_n2848_n452.n0 10.5365
R21284 a_n2848_n452.n81 a_n2848_n452.n25 9.50122
R21285 a_n2848_n452.n15 a_n2848_n452.n13 7.47588
R21286 a_n2848_n452.n94 a_n2848_n452.n7 7.47588
R21287 a_n2848_n452.n81 a_n2848_n452.n16 6.70126
R21288 a_n2848_n452.n26 a_n2848_n452.n102 5.65783
R21289 a_n2848_n452.n94 a_n2848_n452.n81 5.3452
R21290 a_n2848_n452.n18 a_n2848_n452.n20 3.95126
R21291 a_n2848_n452.n6 a_n2848_n452.n2 3.95126
R21292 a_n2848_n452.n104 a_n2848_n452.t44 3.61217
R21293 a_n2848_n452.n104 a_n2848_n452.t34 3.61217
R21294 a_n2848_n452.n103 a_n2848_n452.t42 3.61217
R21295 a_n2848_n452.n103 a_n2848_n452.t26 3.61217
R21296 a_n2848_n452.n72 a_n2848_n452.t32 3.61217
R21297 a_n2848_n452.n72 a_n2848_n452.t40 3.61217
R21298 a_n2848_n452.n71 a_n2848_n452.t28 3.61217
R21299 a_n2848_n452.n71 a_n2848_n452.t24 3.61217
R21300 a_n2848_n452.n65 a_n2848_n452.t1 2.82907
R21301 a_n2848_n452.n65 a_n2848_n452.t6 2.82907
R21302 a_n2848_n452.n66 a_n2848_n452.t14 2.82907
R21303 a_n2848_n452.n66 a_n2848_n452.t15 2.82907
R21304 a_n2848_n452.n68 a_n2848_n452.t10 2.82907
R21305 a_n2848_n452.n68 a_n2848_n452.t11 2.82907
R21306 a_n2848_n452.n64 a_n2848_n452.t2 2.82907
R21307 a_n2848_n452.n64 a_n2848_n452.t7 2.82907
R21308 a_n2848_n452.n62 a_n2848_n452.t47 2.82907
R21309 a_n2848_n452.n62 a_n2848_n452.t3 2.82907
R21310 a_n2848_n452.n60 a_n2848_n452.t9 2.82907
R21311 a_n2848_n452.n60 a_n2848_n452.t18 2.82907
R21312 a_n2848_n452.n56 a_n2848_n452.t17 2.82907
R21313 a_n2848_n452.n56 a_n2848_n452.t13 2.82907
R21314 a_n2848_n452.n57 a_n2848_n452.t20 2.82907
R21315 a_n2848_n452.n57 a_n2848_n452.t19 2.82907
R21316 a_n2848_n452.n59 a_n2848_n452.t45 2.82907
R21317 a_n2848_n452.n59 a_n2848_n452.t0 2.82907
R21318 a_n2848_n452.n55 a_n2848_n452.t5 2.82907
R21319 a_n2848_n452.n55 a_n2848_n452.t4 2.82907
R21320 a_n2848_n452.n53 a_n2848_n452.t8 2.82907
R21321 a_n2848_n452.n53 a_n2848_n452.t12 2.82907
R21322 a_n2848_n452.n52 a_n2848_n452.t46 2.82907
R21323 a_n2848_n452.n52 a_n2848_n452.t16 2.82907
R21324 a_n2848_n452.n102 a_n2848_n452.n13 1.30542
R21325 a_n2848_n452.n10 a_n2848_n452.n11 1.04595
R21326 a_n2848_n452.n5 a_n2848_n452.n97 13.657
R21327 a_n2848_n452.n95 a_n2848_n452.n50 21.4216
R21328 a_n2848_n452.n1 a_n2848_n452.n101 21.4216
R21329 a_n2848_n452.n98 a_n2848_n452.n47 21.4216
R21330 a_n2848_n452.n78 a_n2848_n452.n19 13.657
R21331 a_n2848_n452.n37 a_n2848_n452.n80 21.4216
R21332 a_n2848_n452.n75 a_n2848_n452.n23 13.657
R21333 a_n2848_n452.n34 a_n2848_n452.n77 21.4216
R21334 a_n2848_n452.n0 a_n2848_n452.n6 1.47777
R21335 a_n2848_n452.n22 a_n2848_n452.n21 0.758076
R21336 a_n2848_n452.n21 a_n2848_n452.n20 0.758076
R21337 a_n2848_n452.n18 a_n2848_n452.n17 0.758076
R21338 a_n2848_n452.n17 a_n2848_n452.n16 0.758076
R21339 a_n2848_n452.n15 a_n2848_n452.n14 0.758076
R21340 a_n2848_n452.n12 a_n2848_n452.n11 0.758076
R21341 a_n2848_n452.n10 a_n2848_n452.n9 0.758076
R21342 a_n2848_n452.n8 a_n2848_n452.n7 0.758076
R21343 a_n2848_n452.n4 a_n2848_n452.n2 0.758076
R21344 a_n2848_n452.n4 a_n2848_n452.n3 0.758076
R21345 a_n2848_n452.n27 a_n2848_n452.n26 0.716017
R21346 a_n2848_n452.n25 a_n2848_n452.n24 0.716017
R21347 a_n2848_n452.n12 a_n2848_n452.n14 0.67853
R21348 a_n2848_n452.n8 a_n2848_n452.n9 0.67853
R21349 a_n2848_n452.n28 a_n2848_n452.n54 0.530672
R21350 a_n2848_n452.n29 a_n2848_n452.n58 0.530672
R21351 a_n2848_n452.n63 a_n2848_n452.n61 0.530672
R21352 a_n2848_n452.n30 a_n2848_n452.n63 0.530672
R21353 a_n2848_n452.n31 a_n2848_n452.n67 0.530672
R21354 a_n2848_n452.n31 a_n2848_n452.n30 0.530672
R21355 a_n2848_n452.n29 a_n2848_n452.n28 0.530672
R21356 a_n1986_8322.n6 a_n1986_8322.t6 74.6477
R21357 a_n1986_8322.n1 a_n1986_8322.t13 74.6477
R21358 a_n1986_8322.t22 a_n1986_8322.n18 74.6476
R21359 a_n1986_8322.n14 a_n1986_8322.t15 74.2899
R21360 a_n1986_8322.n7 a_n1986_8322.t4 74.2899
R21361 a_n1986_8322.n8 a_n1986_8322.t7 74.2899
R21362 a_n1986_8322.n11 a_n1986_8322.t8 74.2899
R21363 a_n1986_8322.n4 a_n1986_8322.t12 74.2899
R21364 a_n1986_8322.n18 a_n1986_8322.n17 70.6783
R21365 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R21366 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R21367 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R21368 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R21369 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R21370 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R21371 a_n1986_8322.n13 a_n1986_8322.t2 9.7972
R21372 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R21373 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R21374 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R21375 a_n1986_8322.n17 a_n1986_8322.t20 3.61217
R21376 a_n1986_8322.n17 a_n1986_8322.t17 3.61217
R21377 a_n1986_8322.n15 a_n1986_8322.t14 3.61217
R21378 a_n1986_8322.n15 a_n1986_8322.t23 3.61217
R21379 a_n1986_8322.n5 a_n1986_8322.t10 3.61217
R21380 a_n1986_8322.n5 a_n1986_8322.t9 3.61217
R21381 a_n1986_8322.n9 a_n1986_8322.t5 3.61217
R21382 a_n1986_8322.n9 a_n1986_8322.t11 3.61217
R21383 a_n1986_8322.n0 a_n1986_8322.t21 3.61217
R21384 a_n1986_8322.n0 a_n1986_8322.t16 3.61217
R21385 a_n1986_8322.n2 a_n1986_8322.t19 3.61217
R21386 a_n1986_8322.n2 a_n1986_8322.t18 3.61217
R21387 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R21388 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R21389 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R21390 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R21391 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R21392 a_n1986_8322.n16 a_n1986_8322.n14 0.358259
R21393 a_n1986_8322.n18 a_n1986_8322.n16 0.358259
R21394 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R21395 a_n1986_8322.t3 a_n1986_8322.t0 0.0788333
R21396 a_n1986_8322.t1 a_n1986_8322.t3 0.0631667
R21397 a_n1986_8322.t2 a_n1986_8322.t1 0.0471944
R21398 a_n1986_8322.t2 a_n1986_8322.t0 0.0453889
R21399 a_n1808_13878.n16 a_n1808_13878.n0 98.9633
R21400 a_n1808_13878.n3 a_n1808_13878.n1 98.7517
R21401 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R21402 a_n1808_13878.n3 a_n1808_13878.n2 98.6055
R21403 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R21404 a_n1808_13878.n15 a_n1808_13878.n14 98.6054
R21405 a_n1808_13878.n7 a_n1808_13878.t1 74.6477
R21406 a_n1808_13878.n12 a_n1808_13878.t2 74.2899
R21407 a_n1808_13878.n9 a_n1808_13878.t3 74.2899
R21408 a_n1808_13878.n8 a_n1808_13878.t0 74.2899
R21409 a_n1808_13878.n11 a_n1808_13878.n10 70.6783
R21410 a_n1808_13878.n7 a_n1808_13878.n6 70.6783
R21411 a_n1808_13878.n13 a_n1808_13878.n5 13.5694
R21412 a_n1808_13878.n15 a_n1808_13878.n13 11.5762
R21413 a_n1808_13878.n13 a_n1808_13878.n12 6.2408
R21414 a_n1808_13878.n14 a_n1808_13878.t15 3.61217
R21415 a_n1808_13878.n14 a_n1808_13878.t16 3.61217
R21416 a_n1808_13878.n0 a_n1808_13878.t13 3.61217
R21417 a_n1808_13878.n0 a_n1808_13878.t17 3.61217
R21418 a_n1808_13878.n10 a_n1808_13878.t6 3.61217
R21419 a_n1808_13878.n10 a_n1808_13878.t7 3.61217
R21420 a_n1808_13878.n6 a_n1808_13878.t4 3.61217
R21421 a_n1808_13878.n6 a_n1808_13878.t5 3.61217
R21422 a_n1808_13878.n4 a_n1808_13878.t12 3.61217
R21423 a_n1808_13878.n4 a_n1808_13878.t19 3.61217
R21424 a_n1808_13878.n2 a_n1808_13878.t14 3.61217
R21425 a_n1808_13878.n2 a_n1808_13878.t9 3.61217
R21426 a_n1808_13878.n1 a_n1808_13878.t8 3.61217
R21427 a_n1808_13878.n1 a_n1808_13878.t10 3.61217
R21428 a_n1808_13878.t18 a_n1808_13878.n17 3.61217
R21429 a_n1808_13878.n17 a_n1808_13878.t11 3.61217
R21430 a_n1808_13878.n8 a_n1808_13878.n7 0.358259
R21431 a_n1808_13878.n11 a_n1808_13878.n9 0.358259
R21432 a_n1808_13878.n12 a_n1808_13878.n11 0.358259
R21433 a_n1808_13878.n16 a_n1808_13878.n15 0.358259
R21434 a_n1808_13878.n5 a_n1808_13878.n3 0.146627
R21435 a_n1808_13878.n9 a_n1808_13878.n8 0.101793
R21436 plus.n76 plus.t11 250.337
R21437 plus.n15 plus.t14 250.337
R21438 plus.n124 plus.t1 243.97
R21439 plus.n120 plus.t24 231.093
R21440 plus.n59 plus.t20 231.093
R21441 plus.n124 plus.n123 223.454
R21442 plus.n126 plus.n125 223.454
R21443 plus.n77 plus.t5 187.445
R21444 plus.n74 plus.t22 187.445
R21445 plus.n72 plus.t21 187.445
R21446 plus.n89 plus.t16 187.445
R21447 plus.n95 plus.t17 187.445
R21448 plus.n68 plus.t13 187.445
R21449 plus.n66 plus.t15 187.445
R21450 plus.n107 plus.t10 187.445
R21451 plus.n113 plus.t26 187.445
R21452 plus.n62 plus.t28 187.445
R21453 plus.n1 plus.t23 187.445
R21454 plus.n52 plus.t6 187.445
R21455 plus.n46 plus.t12 187.445
R21456 plus.n5 plus.t8 187.445
R21457 plus.n7 plus.t7 187.445
R21458 plus.n34 plus.t19 187.445
R21459 plus.n28 plus.t18 187.445
R21460 plus.n11 plus.t27 187.445
R21461 plus.n13 plus.t25 187.445
R21462 plus.n16 plus.t9 187.445
R21463 plus.n121 plus.n120 161.3
R21464 plus.n119 plus.n61 161.3
R21465 plus.n118 plus.n117 161.3
R21466 plus.n116 plus.n115 161.3
R21467 plus.n114 plus.n63 161.3
R21468 plus.n112 plus.n111 161.3
R21469 plus.n110 plus.n64 161.3
R21470 plus.n109 plus.n108 161.3
R21471 plus.n106 plus.n65 161.3
R21472 plus.n105 plus.n104 161.3
R21473 plus.n103 plus.n102 161.3
R21474 plus.n101 plus.n67 161.3
R21475 plus.n100 plus.n99 161.3
R21476 plus.n98 plus.n97 161.3
R21477 plus.n96 plus.n69 161.3
R21478 plus.n94 plus.n93 161.3
R21479 plus.n92 plus.n70 161.3
R21480 plus.n91 plus.n90 161.3
R21481 plus.n88 plus.n71 161.3
R21482 plus.n87 plus.n86 161.3
R21483 plus.n85 plus.n84 161.3
R21484 plus.n83 plus.n73 161.3
R21485 plus.n82 plus.n81 161.3
R21486 plus.n80 plus.n79 161.3
R21487 plus.n78 plus.n75 161.3
R21488 plus.n17 plus.n14 161.3
R21489 plus.n19 plus.n18 161.3
R21490 plus.n21 plus.n20 161.3
R21491 plus.n22 plus.n12 161.3
R21492 plus.n24 plus.n23 161.3
R21493 plus.n26 plus.n25 161.3
R21494 plus.n27 plus.n10 161.3
R21495 plus.n30 plus.n29 161.3
R21496 plus.n31 plus.n9 161.3
R21497 plus.n33 plus.n32 161.3
R21498 plus.n35 plus.n8 161.3
R21499 plus.n37 plus.n36 161.3
R21500 plus.n39 plus.n38 161.3
R21501 plus.n40 plus.n6 161.3
R21502 plus.n42 plus.n41 161.3
R21503 plus.n44 plus.n43 161.3
R21504 plus.n45 plus.n4 161.3
R21505 plus.n48 plus.n47 161.3
R21506 plus.n49 plus.n3 161.3
R21507 plus.n51 plus.n50 161.3
R21508 plus.n53 plus.n2 161.3
R21509 plus.n55 plus.n54 161.3
R21510 plus.n57 plus.n56 161.3
R21511 plus.n58 plus.n0 161.3
R21512 plus.n60 plus.n59 161.3
R21513 plus.n88 plus.n87 56.5617
R21514 plus.n97 plus.n96 56.5617
R21515 plus.n106 plus.n105 56.5617
R21516 plus.n45 plus.n44 56.5617
R21517 plus.n36 plus.n35 56.5617
R21518 plus.n27 plus.n26 56.5617
R21519 plus.n79 plus.n78 56.5617
R21520 plus.n115 plus.n114 56.5617
R21521 plus.n54 plus.n53 56.5617
R21522 plus.n18 plus.n17 56.5617
R21523 plus.n119 plus.n118 50.2647
R21524 plus.n58 plus.n57 50.2647
R21525 plus.n84 plus.n83 46.3896
R21526 plus.n108 plus.n64 46.3896
R21527 plus.n47 plus.n3 46.3896
R21528 plus.n23 plus.n22 46.3896
R21529 plus.n76 plus.n75 43.1929
R21530 plus.n15 plus.n14 43.1929
R21531 plus.n94 plus.n70 42.5146
R21532 plus.n101 plus.n100 42.5146
R21533 plus.n40 plus.n39 42.5146
R21534 plus.n33 plus.n9 42.5146
R21535 plus.n77 plus.n76 40.6041
R21536 plus.n16 plus.n15 40.6041
R21537 plus.n90 plus.n70 38.6395
R21538 plus.n102 plus.n101 38.6395
R21539 plus.n41 plus.n40 38.6395
R21540 plus.n29 plus.n9 38.6395
R21541 plus.n122 plus.n121 35.2031
R21542 plus.n83 plus.n82 34.7644
R21543 plus.n112 plus.n64 34.7644
R21544 plus.n51 plus.n3 34.7644
R21545 plus.n22 plus.n21 34.7644
R21546 plus.n79 plus.n74 21.8872
R21547 plus.n114 plus.n113 21.8872
R21548 plus.n53 plus.n52 21.8872
R21549 plus.n18 plus.n13 21.8872
R21550 plus.n89 plus.n88 19.9199
R21551 plus.n105 plus.n66 19.9199
R21552 plus.n44 plus.n5 19.9199
R21553 plus.n28 plus.n27 19.9199
R21554 plus.n123 plus.t2 19.8005
R21555 plus.n123 plus.t4 19.8005
R21556 plus.n125 plus.t3 19.8005
R21557 plus.n125 plus.t0 19.8005
R21558 plus.n96 plus.n95 17.9525
R21559 plus.n97 plus.n68 17.9525
R21560 plus.n36 plus.n7 17.9525
R21561 plus.n35 plus.n34 17.9525
R21562 plus.n87 plus.n72 15.9852
R21563 plus.n107 plus.n106 15.9852
R21564 plus.n46 plus.n45 15.9852
R21565 plus.n26 plus.n11 15.9852
R21566 plus plus.n127 14.4034
R21567 plus.n78 plus.n77 14.0178
R21568 plus.n115 plus.n62 14.0178
R21569 plus.n54 plus.n1 14.0178
R21570 plus.n17 plus.n16 14.0178
R21571 plus.n122 plus.n60 11.9342
R21572 plus.n118 plus.n62 10.575
R21573 plus.n57 plus.n1 10.575
R21574 plus.n120 plus.n119 9.49444
R21575 plus.n59 plus.n58 9.49444
R21576 plus.n84 plus.n72 8.60764
R21577 plus.n108 plus.n107 8.60764
R21578 plus.n47 plus.n46 8.60764
R21579 plus.n23 plus.n11 8.60764
R21580 plus.n95 plus.n94 6.6403
R21581 plus.n100 plus.n68 6.6403
R21582 plus.n39 plus.n7 6.6403
R21583 plus.n34 plus.n33 6.6403
R21584 plus.n127 plus.n126 5.40567
R21585 plus.n90 plus.n89 4.67295
R21586 plus.n102 plus.n66 4.67295
R21587 plus.n41 plus.n5 4.67295
R21588 plus.n29 plus.n28 4.67295
R21589 plus.n82 plus.n74 2.7056
R21590 plus.n113 plus.n112 2.7056
R21591 plus.n52 plus.n51 2.7056
R21592 plus.n21 plus.n13 2.7056
R21593 plus.n127 plus.n122 1.188
R21594 plus.n126 plus.n124 0.716017
R21595 plus.n80 plus.n75 0.189894
R21596 plus.n81 plus.n80 0.189894
R21597 plus.n81 plus.n73 0.189894
R21598 plus.n85 plus.n73 0.189894
R21599 plus.n86 plus.n85 0.189894
R21600 plus.n86 plus.n71 0.189894
R21601 plus.n91 plus.n71 0.189894
R21602 plus.n92 plus.n91 0.189894
R21603 plus.n93 plus.n92 0.189894
R21604 plus.n93 plus.n69 0.189894
R21605 plus.n98 plus.n69 0.189894
R21606 plus.n99 plus.n98 0.189894
R21607 plus.n99 plus.n67 0.189894
R21608 plus.n103 plus.n67 0.189894
R21609 plus.n104 plus.n103 0.189894
R21610 plus.n104 plus.n65 0.189894
R21611 plus.n109 plus.n65 0.189894
R21612 plus.n110 plus.n109 0.189894
R21613 plus.n111 plus.n110 0.189894
R21614 plus.n111 plus.n63 0.189894
R21615 plus.n116 plus.n63 0.189894
R21616 plus.n117 plus.n116 0.189894
R21617 plus.n117 plus.n61 0.189894
R21618 plus.n121 plus.n61 0.189894
R21619 plus.n60 plus.n0 0.189894
R21620 plus.n56 plus.n0 0.189894
R21621 plus.n56 plus.n55 0.189894
R21622 plus.n55 plus.n2 0.189894
R21623 plus.n50 plus.n2 0.189894
R21624 plus.n50 plus.n49 0.189894
R21625 plus.n49 plus.n48 0.189894
R21626 plus.n48 plus.n4 0.189894
R21627 plus.n43 plus.n4 0.189894
R21628 plus.n43 plus.n42 0.189894
R21629 plus.n42 plus.n6 0.189894
R21630 plus.n38 plus.n6 0.189894
R21631 plus.n38 plus.n37 0.189894
R21632 plus.n37 plus.n8 0.189894
R21633 plus.n32 plus.n8 0.189894
R21634 plus.n32 plus.n31 0.189894
R21635 plus.n31 plus.n30 0.189894
R21636 plus.n30 plus.n10 0.189894
R21637 plus.n25 plus.n10 0.189894
R21638 plus.n25 plus.n24 0.189894
R21639 plus.n24 plus.n12 0.189894
R21640 plus.n20 plus.n12 0.189894
R21641 plus.n20 plus.n19 0.189894
R21642 plus.n19 plus.n14 0.189894
R21643 a_n3106_n452.n1 a_n3106_n452.t0 214.321
R21644 a_n3106_n452.n14 a_n3106_n452.t3 214.321
R21645 a_n3106_n452.n15 a_n3106_n452.t34 214.321
R21646 a_n3106_n452.n16 a_n3106_n452.t53 214.321
R21647 a_n3106_n452.n17 a_n3106_n452.t38 214.321
R21648 a_n3106_n452.n18 a_n3106_n452.t36 214.321
R21649 a_n3106_n452.n19 a_n3106_n452.t33 214.321
R21650 a_n3106_n452.n20 a_n3106_n452.t4 214.321
R21651 a_n3106_n452.n0 a_n3106_n452.t22 55.8337
R21652 a_n3106_n452.n2 a_n3106_n452.t35 55.8337
R21653 a_n3106_n452.n13 a_n3106_n452.t40 55.8337
R21654 a_n3106_n452.n47 a_n3106_n452.t9 55.8335
R21655 a_n3106_n452.n45 a_n3106_n452.t44 55.8335
R21656 a_n3106_n452.n34 a_n3106_n452.t54 55.8335
R21657 a_n3106_n452.n33 a_n3106_n452.t19 55.8335
R21658 a_n3106_n452.n22 a_n3106_n452.t13 55.8335
R21659 a_n3106_n452.n49 a_n3106_n452.n48 53.0052
R21660 a_n3106_n452.n51 a_n3106_n452.n50 53.0052
R21661 a_n3106_n452.n53 a_n3106_n452.n52 53.0052
R21662 a_n3106_n452.n55 a_n3106_n452.n54 53.0052
R21663 a_n3106_n452.n4 a_n3106_n452.n3 53.0052
R21664 a_n3106_n452.n6 a_n3106_n452.n5 53.0052
R21665 a_n3106_n452.n8 a_n3106_n452.n7 53.0052
R21666 a_n3106_n452.n10 a_n3106_n452.n9 53.0052
R21667 a_n3106_n452.n12 a_n3106_n452.n11 53.0052
R21668 a_n3106_n452.n44 a_n3106_n452.n43 53.0051
R21669 a_n3106_n452.n42 a_n3106_n452.n41 53.0051
R21670 a_n3106_n452.n40 a_n3106_n452.n39 53.0051
R21671 a_n3106_n452.n38 a_n3106_n452.n37 53.0051
R21672 a_n3106_n452.n36 a_n3106_n452.n35 53.0051
R21673 a_n3106_n452.n32 a_n3106_n452.n31 53.0051
R21674 a_n3106_n452.n30 a_n3106_n452.n29 53.0051
R21675 a_n3106_n452.n28 a_n3106_n452.n27 53.0051
R21676 a_n3106_n452.n26 a_n3106_n452.n25 53.0051
R21677 a_n3106_n452.n24 a_n3106_n452.n23 53.0051
R21678 a_n3106_n452.n57 a_n3106_n452.n56 53.0051
R21679 a_n3106_n452.n21 a_n3106_n452.n13 12.2417
R21680 a_n3106_n452.n47 a_n3106_n452.n46 12.2417
R21681 a_n3106_n452.n22 a_n3106_n452.n21 5.16214
R21682 a_n3106_n452.n46 a_n3106_n452.n45 5.16214
R21683 a_n3106_n452.n48 a_n3106_n452.t7 2.82907
R21684 a_n3106_n452.n48 a_n3106_n452.t5 2.82907
R21685 a_n3106_n452.n50 a_n3106_n452.t18 2.82907
R21686 a_n3106_n452.n50 a_n3106_n452.t23 2.82907
R21687 a_n3106_n452.n52 a_n3106_n452.t16 2.82907
R21688 a_n3106_n452.n52 a_n3106_n452.t20 2.82907
R21689 a_n3106_n452.n54 a_n3106_n452.t12 2.82907
R21690 a_n3106_n452.n54 a_n3106_n452.t17 2.82907
R21691 a_n3106_n452.n3 a_n3106_n452.t46 2.82907
R21692 a_n3106_n452.n3 a_n3106_n452.t2 2.82907
R21693 a_n3106_n452.n5 a_n3106_n452.t42 2.82907
R21694 a_n3106_n452.n5 a_n3106_n452.t45 2.82907
R21695 a_n3106_n452.n7 a_n3106_n452.t37 2.82907
R21696 a_n3106_n452.n7 a_n3106_n452.t41 2.82907
R21697 a_n3106_n452.n9 a_n3106_n452.t30 2.82907
R21698 a_n3106_n452.n9 a_n3106_n452.t29 2.82907
R21699 a_n3106_n452.n11 a_n3106_n452.t49 2.82907
R21700 a_n3106_n452.n11 a_n3106_n452.t55 2.82907
R21701 a_n3106_n452.n43 a_n3106_n452.t50 2.82907
R21702 a_n3106_n452.n43 a_n3106_n452.t48 2.82907
R21703 a_n3106_n452.n41 a_n3106_n452.t1 2.82907
R21704 a_n3106_n452.n41 a_n3106_n452.t51 2.82907
R21705 a_n3106_n452.n39 a_n3106_n452.t31 2.82907
R21706 a_n3106_n452.n39 a_n3106_n452.t52 2.82907
R21707 a_n3106_n452.n37 a_n3106_n452.t43 2.82907
R21708 a_n3106_n452.n37 a_n3106_n452.t32 2.82907
R21709 a_n3106_n452.n35 a_n3106_n452.t47 2.82907
R21710 a_n3106_n452.n35 a_n3106_n452.t39 2.82907
R21711 a_n3106_n452.n31 a_n3106_n452.t8 2.82907
R21712 a_n3106_n452.n31 a_n3106_n452.t24 2.82907
R21713 a_n3106_n452.n29 a_n3106_n452.t15 2.82907
R21714 a_n3106_n452.n29 a_n3106_n452.t6 2.82907
R21715 a_n3106_n452.n27 a_n3106_n452.t26 2.82907
R21716 a_n3106_n452.n27 a_n3106_n452.t14 2.82907
R21717 a_n3106_n452.n25 a_n3106_n452.t21 2.82907
R21718 a_n3106_n452.n25 a_n3106_n452.t25 2.82907
R21719 a_n3106_n452.n23 a_n3106_n452.t10 2.82907
R21720 a_n3106_n452.n23 a_n3106_n452.t27 2.82907
R21721 a_n3106_n452.t28 a_n3106_n452.n57 2.82907
R21722 a_n3106_n452.n57 a_n3106_n452.t11 2.82907
R21723 a_n3106_n452.n46 a_n3106_n452.n1 2.54197
R21724 a_n3106_n452.n21 a_n3106_n452.n20 2.0129
R21725 a_n3106_n452.n20 a_n3106_n452.n19 0.672012
R21726 a_n3106_n452.n19 a_n3106_n452.n18 0.672012
R21727 a_n3106_n452.n18 a_n3106_n452.n17 0.672012
R21728 a_n3106_n452.n17 a_n3106_n452.n16 0.672012
R21729 a_n3106_n452.n16 a_n3106_n452.n15 0.672012
R21730 a_n3106_n452.n15 a_n3106_n452.n14 0.672012
R21731 a_n3106_n452.n14 a_n3106_n452.n1 0.672012
R21732 a_n3106_n452.n24 a_n3106_n452.n22 0.530672
R21733 a_n3106_n452.n26 a_n3106_n452.n24 0.530672
R21734 a_n3106_n452.n28 a_n3106_n452.n26 0.530672
R21735 a_n3106_n452.n30 a_n3106_n452.n28 0.530672
R21736 a_n3106_n452.n32 a_n3106_n452.n30 0.530672
R21737 a_n3106_n452.n33 a_n3106_n452.n32 0.530672
R21738 a_n3106_n452.n36 a_n3106_n452.n34 0.530672
R21739 a_n3106_n452.n38 a_n3106_n452.n36 0.530672
R21740 a_n3106_n452.n40 a_n3106_n452.n38 0.530672
R21741 a_n3106_n452.n42 a_n3106_n452.n40 0.530672
R21742 a_n3106_n452.n44 a_n3106_n452.n42 0.530672
R21743 a_n3106_n452.n45 a_n3106_n452.n44 0.530672
R21744 a_n3106_n452.n13 a_n3106_n452.n12 0.530672
R21745 a_n3106_n452.n12 a_n3106_n452.n10 0.530672
R21746 a_n3106_n452.n10 a_n3106_n452.n8 0.530672
R21747 a_n3106_n452.n8 a_n3106_n452.n6 0.530672
R21748 a_n3106_n452.n6 a_n3106_n452.n4 0.530672
R21749 a_n3106_n452.n4 a_n3106_n452.n2 0.530672
R21750 a_n3106_n452.n56 a_n3106_n452.n0 0.530672
R21751 a_n3106_n452.n56 a_n3106_n452.n55 0.530672
R21752 a_n3106_n452.n55 a_n3106_n452.n53 0.530672
R21753 a_n3106_n452.n53 a_n3106_n452.n51 0.530672
R21754 a_n3106_n452.n51 a_n3106_n452.n49 0.530672
R21755 a_n3106_n452.n49 a_n3106_n452.n47 0.530672
R21756 a_n3106_n452.n34 a_n3106_n452.n33 0.235414
R21757 a_n3106_n452.n2 a_n3106_n452.n0 0.235414
R21758 outputibias.n27 outputibias.n1 289.615
R21759 outputibias.n58 outputibias.n32 289.615
R21760 outputibias.n90 outputibias.n64 289.615
R21761 outputibias.n122 outputibias.n96 289.615
R21762 outputibias.n28 outputibias.n27 185
R21763 outputibias.n26 outputibias.n25 185
R21764 outputibias.n5 outputibias.n4 185
R21765 outputibias.n20 outputibias.n19 185
R21766 outputibias.n18 outputibias.n17 185
R21767 outputibias.n9 outputibias.n8 185
R21768 outputibias.n12 outputibias.n11 185
R21769 outputibias.n59 outputibias.n58 185
R21770 outputibias.n57 outputibias.n56 185
R21771 outputibias.n36 outputibias.n35 185
R21772 outputibias.n51 outputibias.n50 185
R21773 outputibias.n49 outputibias.n48 185
R21774 outputibias.n40 outputibias.n39 185
R21775 outputibias.n43 outputibias.n42 185
R21776 outputibias.n91 outputibias.n90 185
R21777 outputibias.n89 outputibias.n88 185
R21778 outputibias.n68 outputibias.n67 185
R21779 outputibias.n83 outputibias.n82 185
R21780 outputibias.n81 outputibias.n80 185
R21781 outputibias.n72 outputibias.n71 185
R21782 outputibias.n75 outputibias.n74 185
R21783 outputibias.n123 outputibias.n122 185
R21784 outputibias.n121 outputibias.n120 185
R21785 outputibias.n100 outputibias.n99 185
R21786 outputibias.n115 outputibias.n114 185
R21787 outputibias.n113 outputibias.n112 185
R21788 outputibias.n104 outputibias.n103 185
R21789 outputibias.n107 outputibias.n106 185
R21790 outputibias.n0 outputibias.t8 178.945
R21791 outputibias.n133 outputibias.t10 177.018
R21792 outputibias.n132 outputibias.t11 177.018
R21793 outputibias.n0 outputibias.t9 177.018
R21794 outputibias.t5 outputibias.n10 147.661
R21795 outputibias.t7 outputibias.n41 147.661
R21796 outputibias.t1 outputibias.n73 147.661
R21797 outputibias.t3 outputibias.n105 147.661
R21798 outputibias.n128 outputibias.t4 132.363
R21799 outputibias.n128 outputibias.t6 130.436
R21800 outputibias.n129 outputibias.t0 130.436
R21801 outputibias.n130 outputibias.t2 130.436
R21802 outputibias.n27 outputibias.n26 104.615
R21803 outputibias.n26 outputibias.n4 104.615
R21804 outputibias.n19 outputibias.n4 104.615
R21805 outputibias.n19 outputibias.n18 104.615
R21806 outputibias.n18 outputibias.n8 104.615
R21807 outputibias.n11 outputibias.n8 104.615
R21808 outputibias.n58 outputibias.n57 104.615
R21809 outputibias.n57 outputibias.n35 104.615
R21810 outputibias.n50 outputibias.n35 104.615
R21811 outputibias.n50 outputibias.n49 104.615
R21812 outputibias.n49 outputibias.n39 104.615
R21813 outputibias.n42 outputibias.n39 104.615
R21814 outputibias.n90 outputibias.n89 104.615
R21815 outputibias.n89 outputibias.n67 104.615
R21816 outputibias.n82 outputibias.n67 104.615
R21817 outputibias.n82 outputibias.n81 104.615
R21818 outputibias.n81 outputibias.n71 104.615
R21819 outputibias.n74 outputibias.n71 104.615
R21820 outputibias.n122 outputibias.n121 104.615
R21821 outputibias.n121 outputibias.n99 104.615
R21822 outputibias.n114 outputibias.n99 104.615
R21823 outputibias.n114 outputibias.n113 104.615
R21824 outputibias.n113 outputibias.n103 104.615
R21825 outputibias.n106 outputibias.n103 104.615
R21826 outputibias.n63 outputibias.n31 95.6354
R21827 outputibias.n63 outputibias.n62 94.6732
R21828 outputibias.n95 outputibias.n94 94.6732
R21829 outputibias.n127 outputibias.n126 94.6732
R21830 outputibias.n11 outputibias.t5 52.3082
R21831 outputibias.n42 outputibias.t7 52.3082
R21832 outputibias.n74 outputibias.t1 52.3082
R21833 outputibias.n106 outputibias.t3 52.3082
R21834 outputibias.n12 outputibias.n10 15.6674
R21835 outputibias.n43 outputibias.n41 15.6674
R21836 outputibias.n75 outputibias.n73 15.6674
R21837 outputibias.n107 outputibias.n105 15.6674
R21838 outputibias.n13 outputibias.n9 12.8005
R21839 outputibias.n44 outputibias.n40 12.8005
R21840 outputibias.n76 outputibias.n72 12.8005
R21841 outputibias.n108 outputibias.n104 12.8005
R21842 outputibias.n17 outputibias.n16 12.0247
R21843 outputibias.n48 outputibias.n47 12.0247
R21844 outputibias.n80 outputibias.n79 12.0247
R21845 outputibias.n112 outputibias.n111 12.0247
R21846 outputibias.n20 outputibias.n7 11.249
R21847 outputibias.n51 outputibias.n38 11.249
R21848 outputibias.n83 outputibias.n70 11.249
R21849 outputibias.n115 outputibias.n102 11.249
R21850 outputibias.n21 outputibias.n5 10.4732
R21851 outputibias.n52 outputibias.n36 10.4732
R21852 outputibias.n84 outputibias.n68 10.4732
R21853 outputibias.n116 outputibias.n100 10.4732
R21854 outputibias.n25 outputibias.n24 9.69747
R21855 outputibias.n56 outputibias.n55 9.69747
R21856 outputibias.n88 outputibias.n87 9.69747
R21857 outputibias.n120 outputibias.n119 9.69747
R21858 outputibias.n31 outputibias.n30 9.45567
R21859 outputibias.n62 outputibias.n61 9.45567
R21860 outputibias.n94 outputibias.n93 9.45567
R21861 outputibias.n126 outputibias.n125 9.45567
R21862 outputibias.n30 outputibias.n29 9.3005
R21863 outputibias.n3 outputibias.n2 9.3005
R21864 outputibias.n24 outputibias.n23 9.3005
R21865 outputibias.n22 outputibias.n21 9.3005
R21866 outputibias.n7 outputibias.n6 9.3005
R21867 outputibias.n16 outputibias.n15 9.3005
R21868 outputibias.n14 outputibias.n13 9.3005
R21869 outputibias.n61 outputibias.n60 9.3005
R21870 outputibias.n34 outputibias.n33 9.3005
R21871 outputibias.n55 outputibias.n54 9.3005
R21872 outputibias.n53 outputibias.n52 9.3005
R21873 outputibias.n38 outputibias.n37 9.3005
R21874 outputibias.n47 outputibias.n46 9.3005
R21875 outputibias.n45 outputibias.n44 9.3005
R21876 outputibias.n93 outputibias.n92 9.3005
R21877 outputibias.n66 outputibias.n65 9.3005
R21878 outputibias.n87 outputibias.n86 9.3005
R21879 outputibias.n85 outputibias.n84 9.3005
R21880 outputibias.n70 outputibias.n69 9.3005
R21881 outputibias.n79 outputibias.n78 9.3005
R21882 outputibias.n77 outputibias.n76 9.3005
R21883 outputibias.n125 outputibias.n124 9.3005
R21884 outputibias.n98 outputibias.n97 9.3005
R21885 outputibias.n119 outputibias.n118 9.3005
R21886 outputibias.n117 outputibias.n116 9.3005
R21887 outputibias.n102 outputibias.n101 9.3005
R21888 outputibias.n111 outputibias.n110 9.3005
R21889 outputibias.n109 outputibias.n108 9.3005
R21890 outputibias.n28 outputibias.n3 8.92171
R21891 outputibias.n59 outputibias.n34 8.92171
R21892 outputibias.n91 outputibias.n66 8.92171
R21893 outputibias.n123 outputibias.n98 8.92171
R21894 outputibias.n29 outputibias.n1 8.14595
R21895 outputibias.n60 outputibias.n32 8.14595
R21896 outputibias.n92 outputibias.n64 8.14595
R21897 outputibias.n124 outputibias.n96 8.14595
R21898 outputibias.n31 outputibias.n1 5.81868
R21899 outputibias.n62 outputibias.n32 5.81868
R21900 outputibias.n94 outputibias.n64 5.81868
R21901 outputibias.n126 outputibias.n96 5.81868
R21902 outputibias.n131 outputibias.n130 5.20947
R21903 outputibias.n29 outputibias.n28 5.04292
R21904 outputibias.n60 outputibias.n59 5.04292
R21905 outputibias.n92 outputibias.n91 5.04292
R21906 outputibias.n124 outputibias.n123 5.04292
R21907 outputibias.n131 outputibias.n127 4.42209
R21908 outputibias.n14 outputibias.n10 4.38594
R21909 outputibias.n45 outputibias.n41 4.38594
R21910 outputibias.n77 outputibias.n73 4.38594
R21911 outputibias.n109 outputibias.n105 4.38594
R21912 outputibias.n132 outputibias.n131 4.28454
R21913 outputibias.n25 outputibias.n3 4.26717
R21914 outputibias.n56 outputibias.n34 4.26717
R21915 outputibias.n88 outputibias.n66 4.26717
R21916 outputibias.n120 outputibias.n98 4.26717
R21917 outputibias.n24 outputibias.n5 3.49141
R21918 outputibias.n55 outputibias.n36 3.49141
R21919 outputibias.n87 outputibias.n68 3.49141
R21920 outputibias.n119 outputibias.n100 3.49141
R21921 outputibias.n21 outputibias.n20 2.71565
R21922 outputibias.n52 outputibias.n51 2.71565
R21923 outputibias.n84 outputibias.n83 2.71565
R21924 outputibias.n116 outputibias.n115 2.71565
R21925 outputibias.n17 outputibias.n7 1.93989
R21926 outputibias.n48 outputibias.n38 1.93989
R21927 outputibias.n80 outputibias.n70 1.93989
R21928 outputibias.n112 outputibias.n102 1.93989
R21929 outputibias.n130 outputibias.n129 1.9266
R21930 outputibias.n129 outputibias.n128 1.9266
R21931 outputibias.n133 outputibias.n132 1.92658
R21932 outputibias.n134 outputibias.n133 1.29913
R21933 outputibias.n16 outputibias.n9 1.16414
R21934 outputibias.n47 outputibias.n40 1.16414
R21935 outputibias.n79 outputibias.n72 1.16414
R21936 outputibias.n111 outputibias.n104 1.16414
R21937 outputibias.n127 outputibias.n95 0.962709
R21938 outputibias.n95 outputibias.n63 0.962709
R21939 outputibias.n13 outputibias.n12 0.388379
R21940 outputibias.n44 outputibias.n43 0.388379
R21941 outputibias.n76 outputibias.n75 0.388379
R21942 outputibias.n108 outputibias.n107 0.388379
R21943 outputibias.n134 outputibias.n0 0.337251
R21944 outputibias outputibias.n134 0.302375
R21945 outputibias.n30 outputibias.n2 0.155672
R21946 outputibias.n23 outputibias.n2 0.155672
R21947 outputibias.n23 outputibias.n22 0.155672
R21948 outputibias.n22 outputibias.n6 0.155672
R21949 outputibias.n15 outputibias.n6 0.155672
R21950 outputibias.n15 outputibias.n14 0.155672
R21951 outputibias.n61 outputibias.n33 0.155672
R21952 outputibias.n54 outputibias.n33 0.155672
R21953 outputibias.n54 outputibias.n53 0.155672
R21954 outputibias.n53 outputibias.n37 0.155672
R21955 outputibias.n46 outputibias.n37 0.155672
R21956 outputibias.n46 outputibias.n45 0.155672
R21957 outputibias.n93 outputibias.n65 0.155672
R21958 outputibias.n86 outputibias.n65 0.155672
R21959 outputibias.n86 outputibias.n85 0.155672
R21960 outputibias.n85 outputibias.n69 0.155672
R21961 outputibias.n78 outputibias.n69 0.155672
R21962 outputibias.n78 outputibias.n77 0.155672
R21963 outputibias.n125 outputibias.n97 0.155672
R21964 outputibias.n118 outputibias.n97 0.155672
R21965 outputibias.n118 outputibias.n117 0.155672
R21966 outputibias.n117 outputibias.n101 0.155672
R21967 outputibias.n110 outputibias.n101 0.155672
R21968 outputibias.n110 outputibias.n109 0.155672
R21969 output.n41 output.n15 289.615
R21970 output.n72 output.n46 289.615
R21971 output.n104 output.n78 289.615
R21972 output.n136 output.n110 289.615
R21973 output.n77 output.n45 197.26
R21974 output.n77 output.n76 196.298
R21975 output.n109 output.n108 196.298
R21976 output.n141 output.n140 196.298
R21977 output.n42 output.n41 185
R21978 output.n40 output.n39 185
R21979 output.n19 output.n18 185
R21980 output.n34 output.n33 185
R21981 output.n32 output.n31 185
R21982 output.n23 output.n22 185
R21983 output.n26 output.n25 185
R21984 output.n73 output.n72 185
R21985 output.n71 output.n70 185
R21986 output.n50 output.n49 185
R21987 output.n65 output.n64 185
R21988 output.n63 output.n62 185
R21989 output.n54 output.n53 185
R21990 output.n57 output.n56 185
R21991 output.n105 output.n104 185
R21992 output.n103 output.n102 185
R21993 output.n82 output.n81 185
R21994 output.n97 output.n96 185
R21995 output.n95 output.n94 185
R21996 output.n86 output.n85 185
R21997 output.n89 output.n88 185
R21998 output.n137 output.n136 185
R21999 output.n135 output.n134 185
R22000 output.n114 output.n113 185
R22001 output.n129 output.n128 185
R22002 output.n127 output.n126 185
R22003 output.n118 output.n117 185
R22004 output.n121 output.n120 185
R22005 output.t3 output.n24 147.661
R22006 output.t2 output.n55 147.661
R22007 output.t1 output.n87 147.661
R22008 output.t0 output.n119 147.661
R22009 output.n41 output.n40 104.615
R22010 output.n40 output.n18 104.615
R22011 output.n33 output.n18 104.615
R22012 output.n33 output.n32 104.615
R22013 output.n32 output.n22 104.615
R22014 output.n25 output.n22 104.615
R22015 output.n72 output.n71 104.615
R22016 output.n71 output.n49 104.615
R22017 output.n64 output.n49 104.615
R22018 output.n64 output.n63 104.615
R22019 output.n63 output.n53 104.615
R22020 output.n56 output.n53 104.615
R22021 output.n104 output.n103 104.615
R22022 output.n103 output.n81 104.615
R22023 output.n96 output.n81 104.615
R22024 output.n96 output.n95 104.615
R22025 output.n95 output.n85 104.615
R22026 output.n88 output.n85 104.615
R22027 output.n136 output.n135 104.615
R22028 output.n135 output.n113 104.615
R22029 output.n128 output.n113 104.615
R22030 output.n128 output.n127 104.615
R22031 output.n127 output.n117 104.615
R22032 output.n120 output.n117 104.615
R22033 output.n1 output.t19 77.056
R22034 output.n14 output.t4 76.6694
R22035 output.n1 output.n0 72.7095
R22036 output.n3 output.n2 72.7095
R22037 output.n5 output.n4 72.7095
R22038 output.n7 output.n6 72.7095
R22039 output.n9 output.n8 72.7095
R22040 output.n11 output.n10 72.7095
R22041 output.n13 output.n12 72.7095
R22042 output.n25 output.t3 52.3082
R22043 output.n56 output.t2 52.3082
R22044 output.n88 output.t1 52.3082
R22045 output.n120 output.t0 52.3082
R22046 output.n26 output.n24 15.6674
R22047 output.n57 output.n55 15.6674
R22048 output.n89 output.n87 15.6674
R22049 output.n121 output.n119 15.6674
R22050 output.n27 output.n23 12.8005
R22051 output.n58 output.n54 12.8005
R22052 output.n90 output.n86 12.8005
R22053 output.n122 output.n118 12.8005
R22054 output.n31 output.n30 12.0247
R22055 output.n62 output.n61 12.0247
R22056 output.n94 output.n93 12.0247
R22057 output.n126 output.n125 12.0247
R22058 output.n34 output.n21 11.249
R22059 output.n65 output.n52 11.249
R22060 output.n97 output.n84 11.249
R22061 output.n129 output.n116 11.249
R22062 output.n35 output.n19 10.4732
R22063 output.n66 output.n50 10.4732
R22064 output.n98 output.n82 10.4732
R22065 output.n130 output.n114 10.4732
R22066 output.n39 output.n38 9.69747
R22067 output.n70 output.n69 9.69747
R22068 output.n102 output.n101 9.69747
R22069 output.n134 output.n133 9.69747
R22070 output.n45 output.n44 9.45567
R22071 output.n76 output.n75 9.45567
R22072 output.n108 output.n107 9.45567
R22073 output.n140 output.n139 9.45567
R22074 output.n44 output.n43 9.3005
R22075 output.n17 output.n16 9.3005
R22076 output.n38 output.n37 9.3005
R22077 output.n36 output.n35 9.3005
R22078 output.n21 output.n20 9.3005
R22079 output.n30 output.n29 9.3005
R22080 output.n28 output.n27 9.3005
R22081 output.n75 output.n74 9.3005
R22082 output.n48 output.n47 9.3005
R22083 output.n69 output.n68 9.3005
R22084 output.n67 output.n66 9.3005
R22085 output.n52 output.n51 9.3005
R22086 output.n61 output.n60 9.3005
R22087 output.n59 output.n58 9.3005
R22088 output.n107 output.n106 9.3005
R22089 output.n80 output.n79 9.3005
R22090 output.n101 output.n100 9.3005
R22091 output.n99 output.n98 9.3005
R22092 output.n84 output.n83 9.3005
R22093 output.n93 output.n92 9.3005
R22094 output.n91 output.n90 9.3005
R22095 output.n139 output.n138 9.3005
R22096 output.n112 output.n111 9.3005
R22097 output.n133 output.n132 9.3005
R22098 output.n131 output.n130 9.3005
R22099 output.n116 output.n115 9.3005
R22100 output.n125 output.n124 9.3005
R22101 output.n123 output.n122 9.3005
R22102 output.n42 output.n17 8.92171
R22103 output.n73 output.n48 8.92171
R22104 output.n105 output.n80 8.92171
R22105 output.n137 output.n112 8.92171
R22106 output output.n141 8.15037
R22107 output.n43 output.n15 8.14595
R22108 output.n74 output.n46 8.14595
R22109 output.n106 output.n78 8.14595
R22110 output.n138 output.n110 8.14595
R22111 output.n45 output.n15 5.81868
R22112 output.n76 output.n46 5.81868
R22113 output.n108 output.n78 5.81868
R22114 output.n140 output.n110 5.81868
R22115 output.n43 output.n42 5.04292
R22116 output.n74 output.n73 5.04292
R22117 output.n106 output.n105 5.04292
R22118 output.n138 output.n137 5.04292
R22119 output.n28 output.n24 4.38594
R22120 output.n59 output.n55 4.38594
R22121 output.n91 output.n87 4.38594
R22122 output.n123 output.n119 4.38594
R22123 output.n39 output.n17 4.26717
R22124 output.n70 output.n48 4.26717
R22125 output.n102 output.n80 4.26717
R22126 output.n134 output.n112 4.26717
R22127 output.n0 output.t9 3.9605
R22128 output.n0 output.t13 3.9605
R22129 output.n2 output.t16 3.9605
R22130 output.n2 output.t5 3.9605
R22131 output.n4 output.t6 3.9605
R22132 output.n4 output.t11 3.9605
R22133 output.n6 output.t15 3.9605
R22134 output.n6 output.t7 3.9605
R22135 output.n8 output.t10 3.9605
R22136 output.n8 output.t8 3.9605
R22137 output.n10 output.t14 3.9605
R22138 output.n10 output.t17 3.9605
R22139 output.n12 output.t18 3.9605
R22140 output.n12 output.t12 3.9605
R22141 output.n38 output.n19 3.49141
R22142 output.n69 output.n50 3.49141
R22143 output.n101 output.n82 3.49141
R22144 output.n133 output.n114 3.49141
R22145 output.n35 output.n34 2.71565
R22146 output.n66 output.n65 2.71565
R22147 output.n98 output.n97 2.71565
R22148 output.n130 output.n129 2.71565
R22149 output.n31 output.n21 1.93989
R22150 output.n62 output.n52 1.93989
R22151 output.n94 output.n84 1.93989
R22152 output.n126 output.n116 1.93989
R22153 output.n30 output.n23 1.16414
R22154 output.n61 output.n54 1.16414
R22155 output.n93 output.n86 1.16414
R22156 output.n125 output.n118 1.16414
R22157 output.n141 output.n109 0.962709
R22158 output.n109 output.n77 0.962709
R22159 output.n27 output.n26 0.388379
R22160 output.n58 output.n57 0.388379
R22161 output.n90 output.n89 0.388379
R22162 output.n122 output.n121 0.388379
R22163 output.n14 output.n13 0.387128
R22164 output.n13 output.n11 0.387128
R22165 output.n11 output.n9 0.387128
R22166 output.n9 output.n7 0.387128
R22167 output.n7 output.n5 0.387128
R22168 output.n5 output.n3 0.387128
R22169 output.n3 output.n1 0.387128
R22170 output.n44 output.n16 0.155672
R22171 output.n37 output.n16 0.155672
R22172 output.n37 output.n36 0.155672
R22173 output.n36 output.n20 0.155672
R22174 output.n29 output.n20 0.155672
R22175 output.n29 output.n28 0.155672
R22176 output.n75 output.n47 0.155672
R22177 output.n68 output.n47 0.155672
R22178 output.n68 output.n67 0.155672
R22179 output.n67 output.n51 0.155672
R22180 output.n60 output.n51 0.155672
R22181 output.n60 output.n59 0.155672
R22182 output.n107 output.n79 0.155672
R22183 output.n100 output.n79 0.155672
R22184 output.n100 output.n99 0.155672
R22185 output.n99 output.n83 0.155672
R22186 output.n92 output.n83 0.155672
R22187 output.n92 output.n91 0.155672
R22188 output.n139 output.n111 0.155672
R22189 output.n132 output.n111 0.155672
R22190 output.n132 output.n131 0.155672
R22191 output.n131 output.n115 0.155672
R22192 output.n124 output.n115 0.155672
R22193 output.n124 output.n123 0.155672
R22194 output output.n14 0.126227
R22195 minus.n76 minus.t28 250.337
R22196 minus.n15 minus.t20 250.337
R22197 minus.n126 minus.t1 243.255
R22198 minus.n120 minus.t8 231.093
R22199 minus.n59 minus.t10 231.093
R22200 minus.n125 minus.n123 224.169
R22201 minus.n125 minus.n124 223.454
R22202 minus.n62 minus.t12 187.445
R22203 minus.n113 minus.t18 187.445
R22204 minus.n107 minus.t25 187.445
R22205 minus.n66 minus.t22 187.445
R22206 minus.n68 minus.t19 187.445
R22207 minus.n95 minus.t7 187.445
R22208 minus.n89 minus.t6 187.445
R22209 minus.n72 minus.t16 187.445
R22210 minus.n74 minus.t15 187.445
R22211 minus.n77 minus.t23 187.445
R22212 minus.n16 minus.t14 187.445
R22213 minus.n13 minus.t9 187.445
R22214 minus.n11 minus.t5 187.445
R22215 minus.n28 minus.t26 187.445
R22216 minus.n34 minus.t27 187.445
R22217 minus.n7 minus.t21 187.445
R22218 minus.n5 minus.t24 187.445
R22219 minus.n46 minus.t17 187.445
R22220 minus.n52 minus.t11 187.445
R22221 minus.n1 minus.t13 187.445
R22222 minus.n78 minus.n75 161.3
R22223 minus.n80 minus.n79 161.3
R22224 minus.n82 minus.n81 161.3
R22225 minus.n83 minus.n73 161.3
R22226 minus.n85 minus.n84 161.3
R22227 minus.n87 minus.n86 161.3
R22228 minus.n88 minus.n71 161.3
R22229 minus.n91 minus.n90 161.3
R22230 minus.n92 minus.n70 161.3
R22231 minus.n94 minus.n93 161.3
R22232 minus.n96 minus.n69 161.3
R22233 minus.n98 minus.n97 161.3
R22234 minus.n100 minus.n99 161.3
R22235 minus.n101 minus.n67 161.3
R22236 minus.n103 minus.n102 161.3
R22237 minus.n105 minus.n104 161.3
R22238 minus.n106 minus.n65 161.3
R22239 minus.n109 minus.n108 161.3
R22240 minus.n110 minus.n64 161.3
R22241 minus.n112 minus.n111 161.3
R22242 minus.n114 minus.n63 161.3
R22243 minus.n116 minus.n115 161.3
R22244 minus.n118 minus.n117 161.3
R22245 minus.n119 minus.n61 161.3
R22246 minus.n121 minus.n120 161.3
R22247 minus.n60 minus.n59 161.3
R22248 minus.n58 minus.n0 161.3
R22249 minus.n57 minus.n56 161.3
R22250 minus.n55 minus.n54 161.3
R22251 minus.n53 minus.n2 161.3
R22252 minus.n51 minus.n50 161.3
R22253 minus.n49 minus.n3 161.3
R22254 minus.n48 minus.n47 161.3
R22255 minus.n45 minus.n4 161.3
R22256 minus.n44 minus.n43 161.3
R22257 minus.n42 minus.n41 161.3
R22258 minus.n40 minus.n6 161.3
R22259 minus.n39 minus.n38 161.3
R22260 minus.n37 minus.n36 161.3
R22261 minus.n35 minus.n8 161.3
R22262 minus.n33 minus.n32 161.3
R22263 minus.n31 minus.n9 161.3
R22264 minus.n30 minus.n29 161.3
R22265 minus.n27 minus.n10 161.3
R22266 minus.n26 minus.n25 161.3
R22267 minus.n24 minus.n23 161.3
R22268 minus.n22 minus.n12 161.3
R22269 minus.n21 minus.n20 161.3
R22270 minus.n19 minus.n18 161.3
R22271 minus.n17 minus.n14 161.3
R22272 minus.n106 minus.n105 56.5617
R22273 minus.n97 minus.n96 56.5617
R22274 minus.n88 minus.n87 56.5617
R22275 minus.n27 minus.n26 56.5617
R22276 minus.n36 minus.n35 56.5617
R22277 minus.n45 minus.n44 56.5617
R22278 minus.n115 minus.n114 56.5617
R22279 minus.n79 minus.n78 56.5617
R22280 minus.n18 minus.n17 56.5617
R22281 minus.n54 minus.n53 56.5617
R22282 minus.n119 minus.n118 50.2647
R22283 minus.n58 minus.n57 50.2647
R22284 minus.n108 minus.n64 46.3896
R22285 minus.n84 minus.n83 46.3896
R22286 minus.n23 minus.n22 46.3896
R22287 minus.n47 minus.n3 46.3896
R22288 minus.n76 minus.n75 43.1929
R22289 minus.n15 minus.n14 43.1929
R22290 minus.n101 minus.n100 42.5146
R22291 minus.n94 minus.n70 42.5146
R22292 minus.n33 minus.n9 42.5146
R22293 minus.n40 minus.n39 42.5146
R22294 minus.n77 minus.n76 40.6041
R22295 minus.n16 minus.n15 40.6041
R22296 minus.n102 minus.n101 38.6395
R22297 minus.n90 minus.n70 38.6395
R22298 minus.n29 minus.n9 38.6395
R22299 minus.n41 minus.n40 38.6395
R22300 minus.n122 minus.n121 35.4191
R22301 minus.n112 minus.n64 34.7644
R22302 minus.n83 minus.n82 34.7644
R22303 minus.n22 minus.n21 34.7644
R22304 minus.n51 minus.n3 34.7644
R22305 minus.n114 minus.n113 21.8872
R22306 minus.n79 minus.n74 21.8872
R22307 minus.n18 minus.n13 21.8872
R22308 minus.n53 minus.n52 21.8872
R22309 minus.n105 minus.n66 19.9199
R22310 minus.n89 minus.n88 19.9199
R22311 minus.n28 minus.n27 19.9199
R22312 minus.n44 minus.n5 19.9199
R22313 minus.n124 minus.t0 19.8005
R22314 minus.n124 minus.t2 19.8005
R22315 minus.n123 minus.t4 19.8005
R22316 minus.n123 minus.t3 19.8005
R22317 minus.n97 minus.n68 17.9525
R22318 minus.n96 minus.n95 17.9525
R22319 minus.n35 minus.n34 17.9525
R22320 minus.n36 minus.n7 17.9525
R22321 minus.n107 minus.n106 15.9852
R22322 minus.n87 minus.n72 15.9852
R22323 minus.n26 minus.n11 15.9852
R22324 minus.n46 minus.n45 15.9852
R22325 minus.n115 minus.n62 14.0178
R22326 minus.n78 minus.n77 14.0178
R22327 minus.n17 minus.n16 14.0178
R22328 minus.n54 minus.n1 14.0178
R22329 minus.n122 minus.n60 12.1501
R22330 minus minus.n127 10.9162
R22331 minus.n118 minus.n62 10.575
R22332 minus.n57 minus.n1 10.575
R22333 minus.n120 minus.n119 9.49444
R22334 minus.n59 minus.n58 9.49444
R22335 minus.n108 minus.n107 8.60764
R22336 minus.n84 minus.n72 8.60764
R22337 minus.n23 minus.n11 8.60764
R22338 minus.n47 minus.n46 8.60764
R22339 minus.n100 minus.n68 6.6403
R22340 minus.n95 minus.n94 6.6403
R22341 minus.n34 minus.n33 6.6403
R22342 minus.n39 minus.n7 6.6403
R22343 minus.n127 minus.n126 4.80222
R22344 minus.n102 minus.n66 4.67295
R22345 minus.n90 minus.n89 4.67295
R22346 minus.n29 minus.n28 4.67295
R22347 minus.n41 minus.n5 4.67295
R22348 minus.n113 minus.n112 2.7056
R22349 minus.n82 minus.n74 2.7056
R22350 minus.n21 minus.n13 2.7056
R22351 minus.n52 minus.n51 2.7056
R22352 minus.n127 minus.n122 0.972091
R22353 minus.n126 minus.n125 0.716017
R22354 minus.n121 minus.n61 0.189894
R22355 minus.n117 minus.n61 0.189894
R22356 minus.n117 minus.n116 0.189894
R22357 minus.n116 minus.n63 0.189894
R22358 minus.n111 minus.n63 0.189894
R22359 minus.n111 minus.n110 0.189894
R22360 minus.n110 minus.n109 0.189894
R22361 minus.n109 minus.n65 0.189894
R22362 minus.n104 minus.n65 0.189894
R22363 minus.n104 minus.n103 0.189894
R22364 minus.n103 minus.n67 0.189894
R22365 minus.n99 minus.n67 0.189894
R22366 minus.n99 minus.n98 0.189894
R22367 minus.n98 minus.n69 0.189894
R22368 minus.n93 minus.n69 0.189894
R22369 minus.n93 minus.n92 0.189894
R22370 minus.n92 minus.n91 0.189894
R22371 minus.n91 minus.n71 0.189894
R22372 minus.n86 minus.n71 0.189894
R22373 minus.n86 minus.n85 0.189894
R22374 minus.n85 minus.n73 0.189894
R22375 minus.n81 minus.n73 0.189894
R22376 minus.n81 minus.n80 0.189894
R22377 minus.n80 minus.n75 0.189894
R22378 minus.n19 minus.n14 0.189894
R22379 minus.n20 minus.n19 0.189894
R22380 minus.n20 minus.n12 0.189894
R22381 minus.n24 minus.n12 0.189894
R22382 minus.n25 minus.n24 0.189894
R22383 minus.n25 minus.n10 0.189894
R22384 minus.n30 minus.n10 0.189894
R22385 minus.n31 minus.n30 0.189894
R22386 minus.n32 minus.n31 0.189894
R22387 minus.n32 minus.n8 0.189894
R22388 minus.n37 minus.n8 0.189894
R22389 minus.n38 minus.n37 0.189894
R22390 minus.n38 minus.n6 0.189894
R22391 minus.n42 minus.n6 0.189894
R22392 minus.n43 minus.n42 0.189894
R22393 minus.n43 minus.n4 0.189894
R22394 minus.n48 minus.n4 0.189894
R22395 minus.n49 minus.n48 0.189894
R22396 minus.n50 minus.n49 0.189894
R22397 minus.n50 minus.n2 0.189894
R22398 minus.n55 minus.n2 0.189894
R22399 minus.n56 minus.n55 0.189894
R22400 minus.n56 minus.n0 0.189894
R22401 minus.n60 minus.n0 0.189894
R22402 diffpairibias.n0 diffpairibias.t18 436.822
R22403 diffpairibias.n21 diffpairibias.t19 435.479
R22404 diffpairibias.n20 diffpairibias.t16 435.479
R22405 diffpairibias.n19 diffpairibias.t17 435.479
R22406 diffpairibias.n18 diffpairibias.t21 435.479
R22407 diffpairibias.n0 diffpairibias.t22 435.479
R22408 diffpairibias.n1 diffpairibias.t20 435.479
R22409 diffpairibias.n2 diffpairibias.t23 435.479
R22410 diffpairibias.n10 diffpairibias.t0 377.536
R22411 diffpairibias.n10 diffpairibias.t8 376.193
R22412 diffpairibias.n11 diffpairibias.t10 376.193
R22413 diffpairibias.n12 diffpairibias.t6 376.193
R22414 diffpairibias.n13 diffpairibias.t2 376.193
R22415 diffpairibias.n14 diffpairibias.t12 376.193
R22416 diffpairibias.n15 diffpairibias.t4 376.193
R22417 diffpairibias.n16 diffpairibias.t14 376.193
R22418 diffpairibias.n3 diffpairibias.t1 113.368
R22419 diffpairibias.n3 diffpairibias.t9 112.698
R22420 diffpairibias.n4 diffpairibias.t11 112.698
R22421 diffpairibias.n5 diffpairibias.t7 112.698
R22422 diffpairibias.n6 diffpairibias.t3 112.698
R22423 diffpairibias.n7 diffpairibias.t13 112.698
R22424 diffpairibias.n8 diffpairibias.t5 112.698
R22425 diffpairibias.n9 diffpairibias.t15 112.698
R22426 diffpairibias.n17 diffpairibias.n16 4.77242
R22427 diffpairibias.n17 diffpairibias.n9 4.30807
R22428 diffpairibias.n18 diffpairibias.n17 4.13945
R22429 diffpairibias.n16 diffpairibias.n15 1.34352
R22430 diffpairibias.n15 diffpairibias.n14 1.34352
R22431 diffpairibias.n14 diffpairibias.n13 1.34352
R22432 diffpairibias.n13 diffpairibias.n12 1.34352
R22433 diffpairibias.n12 diffpairibias.n11 1.34352
R22434 diffpairibias.n11 diffpairibias.n10 1.34352
R22435 diffpairibias.n2 diffpairibias.n1 1.34352
R22436 diffpairibias.n1 diffpairibias.n0 1.34352
R22437 diffpairibias.n19 diffpairibias.n18 1.34352
R22438 diffpairibias.n20 diffpairibias.n19 1.34352
R22439 diffpairibias.n21 diffpairibias.n20 1.34352
R22440 diffpairibias.n22 diffpairibias.n21 0.862419
R22441 diffpairibias diffpairibias.n22 0.684875
R22442 diffpairibias.n9 diffpairibias.n8 0.672012
R22443 diffpairibias.n8 diffpairibias.n7 0.672012
R22444 diffpairibias.n7 diffpairibias.n6 0.672012
R22445 diffpairibias.n6 diffpairibias.n5 0.672012
R22446 diffpairibias.n5 diffpairibias.n4 0.672012
R22447 diffpairibias.n4 diffpairibias.n3 0.672012
R22448 diffpairibias.n22 diffpairibias.n2 0.190907
C0 minus commonsourceibias 0.515369f
C1 plus commonsourceibias 0.498793f
C2 output outputibias 2.34152f
C3 vdd output 7.23429f
C4 CSoutput output 6.13571f
C5 CSoutput outputibias 0.032386f
C6 vdd CSoutput 0.140826p
C7 minus diffpairibias 5.39e-19
C8 commonsourceibias output 0.006808f
C9 vdd plus 0.096191f
C10 CSoutput minus 2.25384f
C11 plus diffpairibias 4.4e-19
C12 commonsourceibias outputibias 0.003832f
C13 vdd commonsourceibias 0.004218f
C14 CSoutput plus 0.874948f
C15 commonsourceibias diffpairibias 0.052851f
C16 CSoutput commonsourceibias 29.0223f
C17 minus plus 9.674179f
C18 diffpairibias gnd 48.95304f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.118072p
C22 plus gnd 37.535206f
C23 minus gnd 28.66781f
C24 CSoutput gnd 88.04513f
C25 vdd gnd 0.439193p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 minus.n0 gnd 0.031832f
C74 minus.t13 gnd 0.535246f
C75 minus.n1 gnd 0.216477f
C76 minus.n2 gnd 0.031832f
C77 minus.t11 gnd 0.535246f
C78 minus.n3 gnd 0.027201f
C79 minus.n4 gnd 0.031832f
C80 minus.t17 gnd 0.535246f
C81 minus.t24 gnd 0.535246f
C82 minus.n5 gnd 0.216477f
C83 minus.n6 gnd 0.031832f
C84 minus.t21 gnd 0.535246f
C85 minus.n7 gnd 0.216477f
C86 minus.n8 gnd 0.031832f
C87 minus.t27 gnd 0.535246f
C88 minus.n9 gnd 0.025872f
C89 minus.n10 gnd 0.031832f
C90 minus.t26 gnd 0.535246f
C91 minus.t5 gnd 0.535246f
C92 minus.n11 gnd 0.216477f
C93 minus.n12 gnd 0.031832f
C94 minus.t9 gnd 0.535246f
C95 minus.n13 gnd 0.216477f
C96 minus.n14 gnd 0.135091f
C97 minus.t14 gnd 0.535246f
C98 minus.t20 gnd 0.59877f
C99 minus.n15 gnd 0.253084f
C100 minus.n16 gnd 0.247907f
C101 minus.n17 gnd 0.040787f
C102 minus.n18 gnd 0.036021f
C103 minus.n19 gnd 0.031832f
C104 minus.n20 gnd 0.031832f
C105 minus.n21 gnd 0.038039f
C106 minus.n22 gnd 0.027201f
C107 minus.n23 gnd 0.041457f
C108 minus.n24 gnd 0.031832f
C109 minus.n25 gnd 0.031832f
C110 minus.n26 gnd 0.039596f
C111 minus.n27 gnd 0.037213f
C112 minus.n28 gnd 0.216477f
C113 minus.n29 gnd 0.039874f
C114 minus.n30 gnd 0.031832f
C115 minus.n31 gnd 0.031832f
C116 minus.n32 gnd 0.031832f
C117 minus.n33 gnd 0.04095f
C118 minus.n34 gnd 0.216477f
C119 minus.n35 gnd 0.038404f
C120 minus.n36 gnd 0.038404f
C121 minus.n37 gnd 0.031832f
C122 minus.n38 gnd 0.031832f
C123 minus.n39 gnd 0.04095f
C124 minus.n40 gnd 0.025872f
C125 minus.n41 gnd 0.039874f
C126 minus.n42 gnd 0.031832f
C127 minus.n43 gnd 0.031832f
C128 minus.n44 gnd 0.037213f
C129 minus.n45 gnd 0.039596f
C130 minus.n46 gnd 0.216477f
C131 minus.n47 gnd 0.041457f
C132 minus.n48 gnd 0.031832f
C133 minus.n49 gnd 0.031832f
C134 minus.n50 gnd 0.031832f
C135 minus.n51 gnd 0.038039f
C136 minus.n52 gnd 0.216477f
C137 minus.n53 gnd 0.036021f
C138 minus.n54 gnd 0.040787f
C139 minus.n55 gnd 0.031832f
C140 minus.n56 gnd 0.031832f
C141 minus.n57 gnd 0.041526f
C142 minus.n58 gnd 0.011569f
C143 minus.t10 gnd 0.578869f
C144 minus.n59 gnd 0.250644f
C145 minus.n60 gnd 0.372897f
C146 minus.n61 gnd 0.031832f
C147 minus.t8 gnd 0.578869f
C148 minus.t12 gnd 0.535246f
C149 minus.n62 gnd 0.216477f
C150 minus.n63 gnd 0.031832f
C151 minus.t18 gnd 0.535246f
C152 minus.n64 gnd 0.027201f
C153 minus.n65 gnd 0.031832f
C154 minus.t25 gnd 0.535246f
C155 minus.t22 gnd 0.535246f
C156 minus.n66 gnd 0.216477f
C157 minus.n67 gnd 0.031832f
C158 minus.t19 gnd 0.535246f
C159 minus.n68 gnd 0.216477f
C160 minus.n69 gnd 0.031832f
C161 minus.t7 gnd 0.535246f
C162 minus.n70 gnd 0.025872f
C163 minus.n71 gnd 0.031832f
C164 minus.t6 gnd 0.535246f
C165 minus.t16 gnd 0.535246f
C166 minus.n72 gnd 0.216477f
C167 minus.n73 gnd 0.031832f
C168 minus.t15 gnd 0.535246f
C169 minus.n74 gnd 0.216477f
C170 minus.n75 gnd 0.135091f
C171 minus.t23 gnd 0.535246f
C172 minus.t28 gnd 0.59877f
C173 minus.n76 gnd 0.253084f
C174 minus.n77 gnd 0.247907f
C175 minus.n78 gnd 0.040787f
C176 minus.n79 gnd 0.036021f
C177 minus.n80 gnd 0.031832f
C178 minus.n81 gnd 0.031832f
C179 minus.n82 gnd 0.038039f
C180 minus.n83 gnd 0.027201f
C181 minus.n84 gnd 0.041457f
C182 minus.n85 gnd 0.031832f
C183 minus.n86 gnd 0.031832f
C184 minus.n87 gnd 0.039596f
C185 minus.n88 gnd 0.037213f
C186 minus.n89 gnd 0.216477f
C187 minus.n90 gnd 0.039874f
C188 minus.n91 gnd 0.031832f
C189 minus.n92 gnd 0.031832f
C190 minus.n93 gnd 0.031832f
C191 minus.n94 gnd 0.04095f
C192 minus.n95 gnd 0.216477f
C193 minus.n96 gnd 0.038404f
C194 minus.n97 gnd 0.038404f
C195 minus.n98 gnd 0.031832f
C196 minus.n99 gnd 0.031832f
C197 minus.n100 gnd 0.04095f
C198 minus.n101 gnd 0.025872f
C199 minus.n102 gnd 0.039874f
C200 minus.n103 gnd 0.031832f
C201 minus.n104 gnd 0.031832f
C202 minus.n105 gnd 0.037213f
C203 minus.n106 gnd 0.039596f
C204 minus.n107 gnd 0.216477f
C205 minus.n108 gnd 0.041457f
C206 minus.n109 gnd 0.031832f
C207 minus.n110 gnd 0.031832f
C208 minus.n111 gnd 0.031832f
C209 minus.n112 gnd 0.038039f
C210 minus.n113 gnd 0.216477f
C211 minus.n114 gnd 0.036021f
C212 minus.n115 gnd 0.040787f
C213 minus.n116 gnd 0.031832f
C214 minus.n117 gnd 0.031832f
C215 minus.n118 gnd 0.041526f
C216 minus.n119 gnd 0.011569f
C217 minus.n120 gnd 0.250644f
C218 minus.n121 gnd 1.16121f
C219 minus.n122 gnd 1.70573f
C220 minus.t4 gnd 0.009813f
C221 minus.t3 gnd 0.009813f
C222 minus.n123 gnd 0.032267f
C223 minus.t0 gnd 0.009813f
C224 minus.t2 gnd 0.009813f
C225 minus.n124 gnd 0.031825f
C226 minus.n125 gnd 0.271609f
C227 minus.t1 gnd 0.054617f
C228 minus.n126 gnd 0.148215f
C229 minus.n127 gnd 1.6183f
C230 output.t19 gnd 0.464308f
C231 output.t9 gnd 0.044422f
C232 output.t13 gnd 0.044422f
C233 output.n0 gnd 0.364624f
C234 output.n1 gnd 0.614102f
C235 output.t16 gnd 0.044422f
C236 output.t5 gnd 0.044422f
C237 output.n2 gnd 0.364624f
C238 output.n3 gnd 0.350265f
C239 output.t6 gnd 0.044422f
C240 output.t11 gnd 0.044422f
C241 output.n4 gnd 0.364624f
C242 output.n5 gnd 0.350265f
C243 output.t15 gnd 0.044422f
C244 output.t7 gnd 0.044422f
C245 output.n6 gnd 0.364624f
C246 output.n7 gnd 0.350265f
C247 output.t10 gnd 0.044422f
C248 output.t8 gnd 0.044422f
C249 output.n8 gnd 0.364624f
C250 output.n9 gnd 0.350265f
C251 output.t14 gnd 0.044422f
C252 output.t17 gnd 0.044422f
C253 output.n10 gnd 0.364624f
C254 output.n11 gnd 0.350265f
C255 output.t18 gnd 0.044422f
C256 output.t12 gnd 0.044422f
C257 output.n12 gnd 0.364624f
C258 output.n13 gnd 0.350265f
C259 output.t4 gnd 0.462979f
C260 output.n14 gnd 0.28994f
C261 output.n15 gnd 0.015803f
C262 output.n16 gnd 0.011243f
C263 output.n17 gnd 0.006041f
C264 output.n18 gnd 0.01428f
C265 output.n19 gnd 0.006397f
C266 output.n20 gnd 0.011243f
C267 output.n21 gnd 0.006041f
C268 output.n22 gnd 0.01428f
C269 output.n23 gnd 0.006397f
C270 output.n24 gnd 0.048111f
C271 output.t3 gnd 0.023274f
C272 output.n25 gnd 0.01071f
C273 output.n26 gnd 0.008435f
C274 output.n27 gnd 0.006041f
C275 output.n28 gnd 0.267512f
C276 output.n29 gnd 0.011243f
C277 output.n30 gnd 0.006041f
C278 output.n31 gnd 0.006397f
C279 output.n32 gnd 0.01428f
C280 output.n33 gnd 0.01428f
C281 output.n34 gnd 0.006397f
C282 output.n35 gnd 0.006041f
C283 output.n36 gnd 0.011243f
C284 output.n37 gnd 0.011243f
C285 output.n38 gnd 0.006041f
C286 output.n39 gnd 0.006397f
C287 output.n40 gnd 0.01428f
C288 output.n41 gnd 0.030913f
C289 output.n42 gnd 0.006397f
C290 output.n43 gnd 0.006041f
C291 output.n44 gnd 0.025987f
C292 output.n45 gnd 0.097665f
C293 output.n46 gnd 0.015803f
C294 output.n47 gnd 0.011243f
C295 output.n48 gnd 0.006041f
C296 output.n49 gnd 0.01428f
C297 output.n50 gnd 0.006397f
C298 output.n51 gnd 0.011243f
C299 output.n52 gnd 0.006041f
C300 output.n53 gnd 0.01428f
C301 output.n54 gnd 0.006397f
C302 output.n55 gnd 0.048111f
C303 output.t2 gnd 0.023274f
C304 output.n56 gnd 0.01071f
C305 output.n57 gnd 0.008435f
C306 output.n58 gnd 0.006041f
C307 output.n59 gnd 0.267512f
C308 output.n60 gnd 0.011243f
C309 output.n61 gnd 0.006041f
C310 output.n62 gnd 0.006397f
C311 output.n63 gnd 0.01428f
C312 output.n64 gnd 0.01428f
C313 output.n65 gnd 0.006397f
C314 output.n66 gnd 0.006041f
C315 output.n67 gnd 0.011243f
C316 output.n68 gnd 0.011243f
C317 output.n69 gnd 0.006041f
C318 output.n70 gnd 0.006397f
C319 output.n71 gnd 0.01428f
C320 output.n72 gnd 0.030913f
C321 output.n73 gnd 0.006397f
C322 output.n74 gnd 0.006041f
C323 output.n75 gnd 0.025987f
C324 output.n76 gnd 0.09306f
C325 output.n77 gnd 1.65264f
C326 output.n78 gnd 0.015803f
C327 output.n79 gnd 0.011243f
C328 output.n80 gnd 0.006041f
C329 output.n81 gnd 0.01428f
C330 output.n82 gnd 0.006397f
C331 output.n83 gnd 0.011243f
C332 output.n84 gnd 0.006041f
C333 output.n85 gnd 0.01428f
C334 output.n86 gnd 0.006397f
C335 output.n87 gnd 0.048111f
C336 output.t1 gnd 0.023274f
C337 output.n88 gnd 0.01071f
C338 output.n89 gnd 0.008435f
C339 output.n90 gnd 0.006041f
C340 output.n91 gnd 0.267512f
C341 output.n92 gnd 0.011243f
C342 output.n93 gnd 0.006041f
C343 output.n94 gnd 0.006397f
C344 output.n95 gnd 0.01428f
C345 output.n96 gnd 0.01428f
C346 output.n97 gnd 0.006397f
C347 output.n98 gnd 0.006041f
C348 output.n99 gnd 0.011243f
C349 output.n100 gnd 0.011243f
C350 output.n101 gnd 0.006041f
C351 output.n102 gnd 0.006397f
C352 output.n103 gnd 0.01428f
C353 output.n104 gnd 0.030913f
C354 output.n105 gnd 0.006397f
C355 output.n106 gnd 0.006041f
C356 output.n107 gnd 0.025987f
C357 output.n108 gnd 0.09306f
C358 output.n109 gnd 0.713089f
C359 output.n110 gnd 0.015803f
C360 output.n111 gnd 0.011243f
C361 output.n112 gnd 0.006041f
C362 output.n113 gnd 0.01428f
C363 output.n114 gnd 0.006397f
C364 output.n115 gnd 0.011243f
C365 output.n116 gnd 0.006041f
C366 output.n117 gnd 0.01428f
C367 output.n118 gnd 0.006397f
C368 output.n119 gnd 0.048111f
C369 output.t0 gnd 0.023274f
C370 output.n120 gnd 0.01071f
C371 output.n121 gnd 0.008435f
C372 output.n122 gnd 0.006041f
C373 output.n123 gnd 0.267512f
C374 output.n124 gnd 0.011243f
C375 output.n125 gnd 0.006041f
C376 output.n126 gnd 0.006397f
C377 output.n127 gnd 0.01428f
C378 output.n128 gnd 0.01428f
C379 output.n129 gnd 0.006397f
C380 output.n130 gnd 0.006041f
C381 output.n131 gnd 0.011243f
C382 output.n132 gnd 0.011243f
C383 output.n133 gnd 0.006041f
C384 output.n134 gnd 0.006397f
C385 output.n135 gnd 0.01428f
C386 output.n136 gnd 0.030913f
C387 output.n137 gnd 0.006397f
C388 output.n138 gnd 0.006041f
C389 output.n139 gnd 0.025987f
C390 output.n140 gnd 0.09306f
C391 output.n141 gnd 1.67353f
C392 outputibias.t9 gnd 0.11477f
C393 outputibias.t8 gnd 0.115567f
C394 outputibias.n0 gnd 0.130108f
C395 outputibias.n1 gnd 0.001372f
C396 outputibias.n2 gnd 9.76e-19
C397 outputibias.n3 gnd 5.24e-19
C398 outputibias.n4 gnd 0.001239f
C399 outputibias.n5 gnd 5.55e-19
C400 outputibias.n6 gnd 9.76e-19
C401 outputibias.n7 gnd 5.24e-19
C402 outputibias.n8 gnd 0.001239f
C403 outputibias.n9 gnd 5.55e-19
C404 outputibias.n10 gnd 0.004176f
C405 outputibias.t5 gnd 0.00202f
C406 outputibias.n11 gnd 9.3e-19
C407 outputibias.n12 gnd 7.32e-19
C408 outputibias.n13 gnd 5.24e-19
C409 outputibias.n14 gnd 0.02322f
C410 outputibias.n15 gnd 9.76e-19
C411 outputibias.n16 gnd 5.24e-19
C412 outputibias.n17 gnd 5.55e-19
C413 outputibias.n18 gnd 0.001239f
C414 outputibias.n19 gnd 0.001239f
C415 outputibias.n20 gnd 5.55e-19
C416 outputibias.n21 gnd 5.24e-19
C417 outputibias.n22 gnd 9.76e-19
C418 outputibias.n23 gnd 9.76e-19
C419 outputibias.n24 gnd 5.24e-19
C420 outputibias.n25 gnd 5.55e-19
C421 outputibias.n26 gnd 0.001239f
C422 outputibias.n27 gnd 0.002683f
C423 outputibias.n28 gnd 5.55e-19
C424 outputibias.n29 gnd 5.24e-19
C425 outputibias.n30 gnd 0.002256f
C426 outputibias.n31 gnd 0.005781f
C427 outputibias.n32 gnd 0.001372f
C428 outputibias.n33 gnd 9.76e-19
C429 outputibias.n34 gnd 5.24e-19
C430 outputibias.n35 gnd 0.001239f
C431 outputibias.n36 gnd 5.55e-19
C432 outputibias.n37 gnd 9.76e-19
C433 outputibias.n38 gnd 5.24e-19
C434 outputibias.n39 gnd 0.001239f
C435 outputibias.n40 gnd 5.55e-19
C436 outputibias.n41 gnd 0.004176f
C437 outputibias.t7 gnd 0.00202f
C438 outputibias.n42 gnd 9.3e-19
C439 outputibias.n43 gnd 7.32e-19
C440 outputibias.n44 gnd 5.24e-19
C441 outputibias.n45 gnd 0.02322f
C442 outputibias.n46 gnd 9.76e-19
C443 outputibias.n47 gnd 5.24e-19
C444 outputibias.n48 gnd 5.55e-19
C445 outputibias.n49 gnd 0.001239f
C446 outputibias.n50 gnd 0.001239f
C447 outputibias.n51 gnd 5.55e-19
C448 outputibias.n52 gnd 5.24e-19
C449 outputibias.n53 gnd 9.76e-19
C450 outputibias.n54 gnd 9.76e-19
C451 outputibias.n55 gnd 5.24e-19
C452 outputibias.n56 gnd 5.55e-19
C453 outputibias.n57 gnd 0.001239f
C454 outputibias.n58 gnd 0.002683f
C455 outputibias.n59 gnd 5.55e-19
C456 outputibias.n60 gnd 5.24e-19
C457 outputibias.n61 gnd 0.002256f
C458 outputibias.n62 gnd 0.005197f
C459 outputibias.n63 gnd 0.121892f
C460 outputibias.n64 gnd 0.001372f
C461 outputibias.n65 gnd 9.76e-19
C462 outputibias.n66 gnd 5.24e-19
C463 outputibias.n67 gnd 0.001239f
C464 outputibias.n68 gnd 5.55e-19
C465 outputibias.n69 gnd 9.76e-19
C466 outputibias.n70 gnd 5.24e-19
C467 outputibias.n71 gnd 0.001239f
C468 outputibias.n72 gnd 5.55e-19
C469 outputibias.n73 gnd 0.004176f
C470 outputibias.t1 gnd 0.00202f
C471 outputibias.n74 gnd 9.3e-19
C472 outputibias.n75 gnd 7.32e-19
C473 outputibias.n76 gnd 5.24e-19
C474 outputibias.n77 gnd 0.02322f
C475 outputibias.n78 gnd 9.76e-19
C476 outputibias.n79 gnd 5.24e-19
C477 outputibias.n80 gnd 5.55e-19
C478 outputibias.n81 gnd 0.001239f
C479 outputibias.n82 gnd 0.001239f
C480 outputibias.n83 gnd 5.55e-19
C481 outputibias.n84 gnd 5.24e-19
C482 outputibias.n85 gnd 9.76e-19
C483 outputibias.n86 gnd 9.76e-19
C484 outputibias.n87 gnd 5.24e-19
C485 outputibias.n88 gnd 5.55e-19
C486 outputibias.n89 gnd 0.001239f
C487 outputibias.n90 gnd 0.002683f
C488 outputibias.n91 gnd 5.55e-19
C489 outputibias.n92 gnd 5.24e-19
C490 outputibias.n93 gnd 0.002256f
C491 outputibias.n94 gnd 0.005197f
C492 outputibias.n95 gnd 0.064513f
C493 outputibias.n96 gnd 0.001372f
C494 outputibias.n97 gnd 9.76e-19
C495 outputibias.n98 gnd 5.24e-19
C496 outputibias.n99 gnd 0.001239f
C497 outputibias.n100 gnd 5.55e-19
C498 outputibias.n101 gnd 9.76e-19
C499 outputibias.n102 gnd 5.24e-19
C500 outputibias.n103 gnd 0.001239f
C501 outputibias.n104 gnd 5.55e-19
C502 outputibias.n105 gnd 0.004176f
C503 outputibias.t3 gnd 0.00202f
C504 outputibias.n106 gnd 9.3e-19
C505 outputibias.n107 gnd 7.32e-19
C506 outputibias.n108 gnd 5.24e-19
C507 outputibias.n109 gnd 0.02322f
C508 outputibias.n110 gnd 9.76e-19
C509 outputibias.n111 gnd 5.24e-19
C510 outputibias.n112 gnd 5.55e-19
C511 outputibias.n113 gnd 0.001239f
C512 outputibias.n114 gnd 0.001239f
C513 outputibias.n115 gnd 5.55e-19
C514 outputibias.n116 gnd 5.24e-19
C515 outputibias.n117 gnd 9.76e-19
C516 outputibias.n118 gnd 9.76e-19
C517 outputibias.n119 gnd 5.24e-19
C518 outputibias.n120 gnd 5.55e-19
C519 outputibias.n121 gnd 0.001239f
C520 outputibias.n122 gnd 0.002683f
C521 outputibias.n123 gnd 5.55e-19
C522 outputibias.n124 gnd 5.24e-19
C523 outputibias.n125 gnd 0.002256f
C524 outputibias.n126 gnd 0.005197f
C525 outputibias.n127 gnd 0.084814f
C526 outputibias.t2 gnd 0.108319f
C527 outputibias.t0 gnd 0.108319f
C528 outputibias.t6 gnd 0.108319f
C529 outputibias.t4 gnd 0.109238f
C530 outputibias.n128 gnd 0.134674f
C531 outputibias.n129 gnd 0.07244f
C532 outputibias.n130 gnd 0.079818f
C533 outputibias.n131 gnd 0.164901f
C534 outputibias.t11 gnd 0.11477f
C535 outputibias.n132 gnd 0.067481f
C536 outputibias.t10 gnd 0.11477f
C537 outputibias.n133 gnd 0.065115f
C538 outputibias.n134 gnd 0.029159f
C539 a_n3106_n452.t11 gnd 0.10001f
C540 a_n3106_n452.t22 gnd 1.03942f
C541 a_n3106_n452.n0 gnd 0.392946f
C542 a_n3106_n452.t0 gnd 1.29145f
C543 a_n3106_n452.n1 gnd 1.22854f
C544 a_n3106_n452.t35 gnd 1.03942f
C545 a_n3106_n452.n2 gnd 0.392946f
C546 a_n3106_n452.t46 gnd 0.10001f
C547 a_n3106_n452.t2 gnd 0.10001f
C548 a_n3106_n452.n3 gnd 0.816794f
C549 a_n3106_n452.n4 gnd 0.411618f
C550 a_n3106_n452.t42 gnd 0.10001f
C551 a_n3106_n452.t45 gnd 0.10001f
C552 a_n3106_n452.n5 gnd 0.816794f
C553 a_n3106_n452.n6 gnd 0.411618f
C554 a_n3106_n452.t37 gnd 0.10001f
C555 a_n3106_n452.t41 gnd 0.10001f
C556 a_n3106_n452.n7 gnd 0.816794f
C557 a_n3106_n452.n8 gnd 0.411618f
C558 a_n3106_n452.t30 gnd 0.10001f
C559 a_n3106_n452.t29 gnd 0.10001f
C560 a_n3106_n452.n9 gnd 0.816794f
C561 a_n3106_n452.n10 gnd 0.411618f
C562 a_n3106_n452.t49 gnd 0.10001f
C563 a_n3106_n452.t55 gnd 0.10001f
C564 a_n3106_n452.n11 gnd 0.816794f
C565 a_n3106_n452.n12 gnd 0.411618f
C566 a_n3106_n452.t40 gnd 1.03942f
C567 a_n3106_n452.n13 gnd 0.972974f
C568 a_n3106_n452.t3 gnd 1.29145f
C569 a_n3106_n452.n14 gnd 0.909591f
C570 a_n3106_n452.t34 gnd 1.29145f
C571 a_n3106_n452.n15 gnd 0.909591f
C572 a_n3106_n452.t53 gnd 1.29145f
C573 a_n3106_n452.n16 gnd 0.909591f
C574 a_n3106_n452.t38 gnd 1.29145f
C575 a_n3106_n452.n17 gnd 0.909591f
C576 a_n3106_n452.t36 gnd 1.29145f
C577 a_n3106_n452.n18 gnd 0.909591f
C578 a_n3106_n452.t33 gnd 1.29145f
C579 a_n3106_n452.n19 gnd 0.909591f
C580 a_n3106_n452.t4 gnd 1.29145f
C581 a_n3106_n452.n20 gnd 0.789472f
C582 a_n3106_n452.n21 gnd 0.948419f
C583 a_n3106_n452.t13 gnd 1.03941f
C584 a_n3106_n452.n22 gnd 0.645631f
C585 a_n3106_n452.t10 gnd 0.10001f
C586 a_n3106_n452.t27 gnd 0.10001f
C587 a_n3106_n452.n23 gnd 0.816793f
C588 a_n3106_n452.n24 gnd 0.41162f
C589 a_n3106_n452.t21 gnd 0.10001f
C590 a_n3106_n452.t25 gnd 0.10001f
C591 a_n3106_n452.n25 gnd 0.816793f
C592 a_n3106_n452.n26 gnd 0.41162f
C593 a_n3106_n452.t26 gnd 0.10001f
C594 a_n3106_n452.t14 gnd 0.10001f
C595 a_n3106_n452.n27 gnd 0.816793f
C596 a_n3106_n452.n28 gnd 0.41162f
C597 a_n3106_n452.t15 gnd 0.10001f
C598 a_n3106_n452.t6 gnd 0.10001f
C599 a_n3106_n452.n29 gnd 0.816793f
C600 a_n3106_n452.n30 gnd 0.41162f
C601 a_n3106_n452.t8 gnd 0.10001f
C602 a_n3106_n452.t24 gnd 0.10001f
C603 a_n3106_n452.n31 gnd 0.816793f
C604 a_n3106_n452.n32 gnd 0.41162f
C605 a_n3106_n452.t19 gnd 1.03941f
C606 a_n3106_n452.n33 gnd 0.39295f
C607 a_n3106_n452.t54 gnd 1.03941f
C608 a_n3106_n452.n34 gnd 0.39295f
C609 a_n3106_n452.t47 gnd 0.10001f
C610 a_n3106_n452.t39 gnd 0.10001f
C611 a_n3106_n452.n35 gnd 0.816793f
C612 a_n3106_n452.n36 gnd 0.41162f
C613 a_n3106_n452.t43 gnd 0.10001f
C614 a_n3106_n452.t32 gnd 0.10001f
C615 a_n3106_n452.n37 gnd 0.816793f
C616 a_n3106_n452.n38 gnd 0.41162f
C617 a_n3106_n452.t31 gnd 0.10001f
C618 a_n3106_n452.t52 gnd 0.10001f
C619 a_n3106_n452.n39 gnd 0.816793f
C620 a_n3106_n452.n40 gnd 0.41162f
C621 a_n3106_n452.t1 gnd 0.10001f
C622 a_n3106_n452.t51 gnd 0.10001f
C623 a_n3106_n452.n41 gnd 0.816793f
C624 a_n3106_n452.n42 gnd 0.41162f
C625 a_n3106_n452.t50 gnd 0.10001f
C626 a_n3106_n452.t48 gnd 0.10001f
C627 a_n3106_n452.n43 gnd 0.816793f
C628 a_n3106_n452.n44 gnd 0.41162f
C629 a_n3106_n452.t44 gnd 1.03941f
C630 a_n3106_n452.n45 gnd 0.645631f
C631 a_n3106_n452.n46 gnd 1.05146f
C632 a_n3106_n452.t9 gnd 1.03941f
C633 a_n3106_n452.n47 gnd 0.972978f
C634 a_n3106_n452.t7 gnd 0.10001f
C635 a_n3106_n452.t5 gnd 0.10001f
C636 a_n3106_n452.n48 gnd 0.816794f
C637 a_n3106_n452.n49 gnd 0.411618f
C638 a_n3106_n452.t18 gnd 0.10001f
C639 a_n3106_n452.t23 gnd 0.10001f
C640 a_n3106_n452.n50 gnd 0.816794f
C641 a_n3106_n452.n51 gnd 0.411618f
C642 a_n3106_n452.t16 gnd 0.10001f
C643 a_n3106_n452.t20 gnd 0.10001f
C644 a_n3106_n452.n52 gnd 0.816794f
C645 a_n3106_n452.n53 gnd 0.411618f
C646 a_n3106_n452.t12 gnd 0.10001f
C647 a_n3106_n452.t17 gnd 0.10001f
C648 a_n3106_n452.n54 gnd 0.816794f
C649 a_n3106_n452.n55 gnd 0.411618f
C650 a_n3106_n452.n56 gnd 0.411617f
C651 a_n3106_n452.n57 gnd 0.816796f
C652 a_n3106_n452.t28 gnd 0.10001f
C653 plus.n0 gnd 0.023652f
C654 plus.t20 gnd 0.430126f
C655 plus.t23 gnd 0.397712f
C656 plus.n1 gnd 0.160852f
C657 plus.n2 gnd 0.023652f
C658 plus.t6 gnd 0.397712f
C659 plus.n3 gnd 0.020211f
C660 plus.n4 gnd 0.023652f
C661 plus.t12 gnd 0.397712f
C662 plus.t8 gnd 0.397712f
C663 plus.n5 gnd 0.160852f
C664 plus.n6 gnd 0.023652f
C665 plus.t7 gnd 0.397712f
C666 plus.n7 gnd 0.160852f
C667 plus.n8 gnd 0.023652f
C668 plus.t19 gnd 0.397712f
C669 plus.n9 gnd 0.019224f
C670 plus.n10 gnd 0.023652f
C671 plus.t18 gnd 0.397712f
C672 plus.t27 gnd 0.397712f
C673 plus.n11 gnd 0.160852f
C674 plus.n12 gnd 0.023652f
C675 plus.t25 gnd 0.397712f
C676 plus.n13 gnd 0.160852f
C677 plus.n14 gnd 0.100378f
C678 plus.t9 gnd 0.397712f
C679 plus.t14 gnd 0.444913f
C680 plus.n15 gnd 0.188053f
C681 plus.n16 gnd 0.184206f
C682 plus.n17 gnd 0.030307f
C683 plus.n18 gnd 0.026765f
C684 plus.n19 gnd 0.023652f
C685 plus.n20 gnd 0.023652f
C686 plus.n21 gnd 0.028265f
C687 plus.n22 gnd 0.020211f
C688 plus.n23 gnd 0.030804f
C689 plus.n24 gnd 0.023652f
C690 plus.n25 gnd 0.023652f
C691 plus.n26 gnd 0.029422f
C692 plus.n27 gnd 0.027651f
C693 plus.n28 gnd 0.160852f
C694 plus.n29 gnd 0.029629f
C695 plus.n30 gnd 0.023652f
C696 plus.n31 gnd 0.023652f
C697 plus.n32 gnd 0.023652f
C698 plus.n33 gnd 0.030428f
C699 plus.n34 gnd 0.160852f
C700 plus.n35 gnd 0.028536f
C701 plus.n36 gnd 0.028536f
C702 plus.n37 gnd 0.023652f
C703 plus.n38 gnd 0.023652f
C704 plus.n39 gnd 0.030428f
C705 plus.n40 gnd 0.019224f
C706 plus.n41 gnd 0.029629f
C707 plus.n42 gnd 0.023652f
C708 plus.n43 gnd 0.023652f
C709 plus.n44 gnd 0.027651f
C710 plus.n45 gnd 0.029422f
C711 plus.n46 gnd 0.160852f
C712 plus.n47 gnd 0.030804f
C713 plus.n48 gnd 0.023652f
C714 plus.n49 gnd 0.023652f
C715 plus.n50 gnd 0.023652f
C716 plus.n51 gnd 0.028265f
C717 plus.n52 gnd 0.160852f
C718 plus.n53 gnd 0.026765f
C719 plus.n54 gnd 0.030307f
C720 plus.n55 gnd 0.023652f
C721 plus.n56 gnd 0.023652f
C722 plus.n57 gnd 0.030855f
C723 plus.n58 gnd 0.008596f
C724 plus.n59 gnd 0.18624f
C725 plus.n60 gnd 0.270994f
C726 plus.n61 gnd 0.023652f
C727 plus.t28 gnd 0.397712f
C728 plus.n62 gnd 0.160852f
C729 plus.n63 gnd 0.023652f
C730 plus.t26 gnd 0.397712f
C731 plus.n64 gnd 0.020211f
C732 plus.n65 gnd 0.023652f
C733 plus.t10 gnd 0.397712f
C734 plus.t15 gnd 0.397712f
C735 plus.n66 gnd 0.160852f
C736 plus.n67 gnd 0.023652f
C737 plus.t13 gnd 0.397712f
C738 plus.n68 gnd 0.160852f
C739 plus.n69 gnd 0.023652f
C740 plus.t17 gnd 0.397712f
C741 plus.n70 gnd 0.019224f
C742 plus.n71 gnd 0.023652f
C743 plus.t16 gnd 0.397712f
C744 plus.t21 gnd 0.397712f
C745 plus.n72 gnd 0.160852f
C746 plus.n73 gnd 0.023652f
C747 plus.t22 gnd 0.397712f
C748 plus.n74 gnd 0.160852f
C749 plus.n75 gnd 0.100378f
C750 plus.t5 gnd 0.397712f
C751 plus.t11 gnd 0.444913f
C752 plus.n76 gnd 0.188053f
C753 plus.n77 gnd 0.184206f
C754 plus.n78 gnd 0.030307f
C755 plus.n79 gnd 0.026765f
C756 plus.n80 gnd 0.023652f
C757 plus.n81 gnd 0.023652f
C758 plus.n82 gnd 0.028265f
C759 plus.n83 gnd 0.020211f
C760 plus.n84 gnd 0.030804f
C761 plus.n85 gnd 0.023652f
C762 plus.n86 gnd 0.023652f
C763 plus.n87 gnd 0.029422f
C764 plus.n88 gnd 0.027651f
C765 plus.n89 gnd 0.160852f
C766 plus.n90 gnd 0.029629f
C767 plus.n91 gnd 0.023652f
C768 plus.n92 gnd 0.023652f
C769 plus.n93 gnd 0.023652f
C770 plus.n94 gnd 0.030428f
C771 plus.n95 gnd 0.160852f
C772 plus.n96 gnd 0.028536f
C773 plus.n97 gnd 0.028536f
C774 plus.n98 gnd 0.023652f
C775 plus.n99 gnd 0.023652f
C776 plus.n100 gnd 0.030428f
C777 plus.n101 gnd 0.019224f
C778 plus.n102 gnd 0.029629f
C779 plus.n103 gnd 0.023652f
C780 plus.n104 gnd 0.023652f
C781 plus.n105 gnd 0.027651f
C782 plus.n106 gnd 0.029422f
C783 plus.n107 gnd 0.160852f
C784 plus.n108 gnd 0.030804f
C785 plus.n109 gnd 0.023652f
C786 plus.n110 gnd 0.023652f
C787 plus.n111 gnd 0.023652f
C788 plus.n112 gnd 0.028265f
C789 plus.n113 gnd 0.160852f
C790 plus.n114 gnd 0.026765f
C791 plus.n115 gnd 0.030307f
C792 plus.n116 gnd 0.023652f
C793 plus.n117 gnd 0.023652f
C794 plus.n118 gnd 0.030855f
C795 plus.n119 gnd 0.008596f
C796 plus.t24 gnd 0.430126f
C797 plus.n120 gnd 0.18624f
C798 plus.n121 gnd 0.853371f
C799 plus.n122 gnd 1.25804f
C800 plus.t1 gnd 0.040831f
C801 plus.t2 gnd 0.007291f
C802 plus.t4 gnd 0.007291f
C803 plus.n123 gnd 0.023647f
C804 plus.n124 gnd 0.183575f
C805 plus.t3 gnd 0.007291f
C806 plus.t0 gnd 0.007291f
C807 plus.n125 gnd 0.023647f
C808 plus.n126 gnd 0.137795f
C809 plus.n127 gnd 2.64316f
C810 a_n1808_13878.t11 gnd 0.185195f
C811 a_n1808_13878.t13 gnd 0.185195f
C812 a_n1808_13878.t17 gnd 0.185195f
C813 a_n1808_13878.n0 gnd 1.46067f
C814 a_n1808_13878.t8 gnd 0.185195f
C815 a_n1808_13878.t10 gnd 0.185195f
C816 a_n1808_13878.n1 gnd 1.4598f
C817 a_n1808_13878.t14 gnd 0.185195f
C818 a_n1808_13878.t9 gnd 0.185195f
C819 a_n1808_13878.n2 gnd 1.45825f
C820 a_n1808_13878.n3 gnd 2.03762f
C821 a_n1808_13878.t12 gnd 0.185195f
C822 a_n1808_13878.t19 gnd 0.185195f
C823 a_n1808_13878.n4 gnd 1.45825f
C824 a_n1808_13878.n5 gnd 3.69301f
C825 a_n1808_13878.t1 gnd 1.73408f
C826 a_n1808_13878.t4 gnd 0.185195f
C827 a_n1808_13878.t5 gnd 0.185195f
C828 a_n1808_13878.n6 gnd 1.30452f
C829 a_n1808_13878.n7 gnd 1.4576f
C830 a_n1808_13878.t0 gnd 1.73062f
C831 a_n1808_13878.n8 gnd 0.733487f
C832 a_n1808_13878.t3 gnd 1.73062f
C833 a_n1808_13878.n9 gnd 0.733487f
C834 a_n1808_13878.t6 gnd 0.185195f
C835 a_n1808_13878.t7 gnd 0.185195f
C836 a_n1808_13878.n10 gnd 1.30452f
C837 a_n1808_13878.n11 gnd 0.74059f
C838 a_n1808_13878.t2 gnd 1.73062f
C839 a_n1808_13878.n12 gnd 1.7272f
C840 a_n1808_13878.n13 gnd 2.51438f
C841 a_n1808_13878.t15 gnd 0.185195f
C842 a_n1808_13878.t16 gnd 0.185195f
C843 a_n1808_13878.n14 gnd 1.45825f
C844 a_n1808_13878.n15 gnd 1.80025f
C845 a_n1808_13878.n16 gnd 1.31079f
C846 a_n1808_13878.n17 gnd 1.45826f
C847 a_n1808_13878.t18 gnd 0.185195f
C848 a_n1986_8322.t0 gnd 38.672398f
C849 a_n1986_8322.t2 gnd 27.512402f
C850 a_n1986_8322.t3 gnd 19.268198f
C851 a_n1986_8322.t1 gnd 38.672398f
C852 a_n1986_8322.t13 gnd 0.875792f
C853 a_n1986_8322.t21 gnd 0.093533f
C854 a_n1986_8322.t16 gnd 0.093533f
C855 a_n1986_8322.n0 gnd 0.658844f
C856 a_n1986_8322.n1 gnd 0.736161f
C857 a_n1986_8322.t19 gnd 0.093533f
C858 a_n1986_8322.t18 gnd 0.093533f
C859 a_n1986_8322.n2 gnd 0.658844f
C860 a_n1986_8322.n3 gnd 0.374034f
C861 a_n1986_8322.t12 gnd 0.874048f
C862 a_n1986_8322.n4 gnd 1.39896f
C863 a_n1986_8322.t6 gnd 0.875792f
C864 a_n1986_8322.t10 gnd 0.093533f
C865 a_n1986_8322.t9 gnd 0.093533f
C866 a_n1986_8322.n5 gnd 0.658844f
C867 a_n1986_8322.n6 gnd 0.736161f
C868 a_n1986_8322.t4 gnd 0.874048f
C869 a_n1986_8322.n7 gnd 0.370446f
C870 a_n1986_8322.t7 gnd 0.874048f
C871 a_n1986_8322.n8 gnd 0.370446f
C872 a_n1986_8322.t5 gnd 0.093533f
C873 a_n1986_8322.t11 gnd 0.093533f
C874 a_n1986_8322.n9 gnd 0.658844f
C875 a_n1986_8322.n10 gnd 0.374034f
C876 a_n1986_8322.t8 gnd 0.874048f
C877 a_n1986_8322.n11 gnd 0.872317f
C878 a_n1986_8322.n12 gnd 1.59071f
C879 a_n1986_8322.n13 gnd 3.20172f
C880 a_n1986_8322.t15 gnd 0.874048f
C881 a_n1986_8322.n14 gnd 0.76652f
C882 a_n1986_8322.t14 gnd 0.093533f
C883 a_n1986_8322.t23 gnd 0.093533f
C884 a_n1986_8322.n15 gnd 0.658844f
C885 a_n1986_8322.n16 gnd 0.374034f
C886 a_n1986_8322.t20 gnd 0.093533f
C887 a_n1986_8322.t17 gnd 0.093533f
C888 a_n1986_8322.n17 gnd 0.658844f
C889 a_n1986_8322.n18 gnd 0.736159f
C890 a_n1986_8322.t22 gnd 0.875794f
C891 a_n2848_n452.n0 gnd 3.415f
C892 a_n2848_n452.n1 gnd 0.285666f
C893 a_n2848_n452.n2 gnd 0.492471f
C894 a_n2848_n452.n3 gnd 0.664435f
C895 a_n2848_n452.n4 gnd 0.215942f
C896 a_n2848_n452.n5 gnd 0.282512f
C897 a_n2848_n452.n6 gnd 0.546457f
C898 a_n2848_n452.n7 gnd 0.526038f
C899 a_n2848_n452.n8 gnd 0.204894f
C900 a_n2848_n452.n9 gnd 0.150908f
C901 a_n2848_n452.n10 gnd 0.23718f
C902 a_n2848_n452.n11 gnd 0.183194f
C903 a_n2848_n452.n12 gnd 0.204894f
C904 a_n2848_n452.n13 gnd 1.0063f
C905 a_n2848_n452.n14 gnd 0.150908f
C906 a_n2848_n452.n15 gnd 0.580023f
C907 a_n2848_n452.n16 gnd 0.432289f
C908 a_n2848_n452.n17 gnd 0.215942f
C909 a_n2848_n452.n18 gnd 0.492471f
C910 a_n2848_n452.n19 gnd 0.282512f
C911 a_n2848_n452.n20 gnd 0.438486f
C912 a_n2848_n452.n21 gnd 0.215942f
C913 a_n2848_n452.n22 gnd 0.731535f
C914 a_n2848_n452.n23 gnd 0.282512f
C915 a_n2848_n452.n24 gnd 1.17886f
C916 a_n2848_n452.n25 gnd 1.91568f
C917 a_n2848_n452.n26 gnd 1.14458f
C918 a_n2848_n452.n27 gnd 1.77783f
C919 a_n2848_n452.n28 gnd 0.377489f
C920 a_n2848_n452.n29 gnd 3.11576f
C921 a_n2848_n452.n30 gnd 0.377488f
C922 a_n2848_n452.n31 gnd 3.20158f
C923 a_n2848_n452.n32 gnd 0.008361f
C924 a_n2848_n452.n34 gnd 0.285666f
C925 a_n2848_n452.n35 gnd 0.008361f
C926 a_n2848_n452.n37 gnd 0.285666f
C927 a_n2848_n452.n38 gnd 0.008361f
C928 a_n2848_n452.n39 gnd 0.28526f
C929 a_n2848_n452.n40 gnd 0.008361f
C930 a_n2848_n452.n41 gnd 0.28526f
C931 a_n2848_n452.n42 gnd 0.008361f
C932 a_n2848_n452.n43 gnd 0.28526f
C933 a_n2848_n452.n44 gnd 0.008361f
C934 a_n2848_n452.n45 gnd 0.28526f
C935 a_n2848_n452.n47 gnd 0.285666f
C936 a_n2848_n452.n48 gnd 0.008361f
C937 a_n2848_n452.n50 gnd 0.285666f
C938 a_n2848_n452.t37 gnd 0.708223f
C939 a_n2848_n452.t41 gnd 0.696704f
C940 a_n2848_n452.t25 gnd 0.696704f
C941 a_n2848_n452.t46 gnd 0.116496f
C942 a_n2848_n452.t16 gnd 0.116496f
C943 a_n2848_n452.n52 gnd 1.03243f
C944 a_n2848_n452.t8 gnd 0.116496f
C945 a_n2848_n452.t12 gnd 0.116496f
C946 a_n2848_n452.n53 gnd 1.0294f
C947 a_n2848_n452.n54 gnd 0.912817f
C948 a_n2848_n452.t5 gnd 0.116496f
C949 a_n2848_n452.t4 gnd 0.116496f
C950 a_n2848_n452.n55 gnd 1.0294f
C951 a_n2848_n452.t17 gnd 0.116496f
C952 a_n2848_n452.t13 gnd 0.116496f
C953 a_n2848_n452.n56 gnd 1.03243f
C954 a_n2848_n452.t20 gnd 0.116496f
C955 a_n2848_n452.t19 gnd 0.116496f
C956 a_n2848_n452.n57 gnd 1.0294f
C957 a_n2848_n452.n58 gnd 0.912817f
C958 a_n2848_n452.t45 gnd 0.116496f
C959 a_n2848_n452.t0 gnd 0.116496f
C960 a_n2848_n452.n59 gnd 1.0294f
C961 a_n2848_n452.t9 gnd 0.116496f
C962 a_n2848_n452.t18 gnd 0.116496f
C963 a_n2848_n452.n60 gnd 1.0294f
C964 a_n2848_n452.n61 gnd 3.15028f
C965 a_n2848_n452.t47 gnd 0.116496f
C966 a_n2848_n452.t3 gnd 0.116496f
C967 a_n2848_n452.n62 gnd 1.0294f
C968 a_n2848_n452.n63 gnd 0.449443f
C969 a_n2848_n452.t2 gnd 0.116496f
C970 a_n2848_n452.t7 gnd 0.116496f
C971 a_n2848_n452.n64 gnd 1.0294f
C972 a_n2848_n452.t1 gnd 0.116496f
C973 a_n2848_n452.t6 gnd 0.116496f
C974 a_n2848_n452.n65 gnd 1.03243f
C975 a_n2848_n452.t14 gnd 0.116496f
C976 a_n2848_n452.t15 gnd 0.116496f
C977 a_n2848_n452.n66 gnd 1.0294f
C978 a_n2848_n452.n67 gnd 0.912814f
C979 a_n2848_n452.t10 gnd 0.116496f
C980 a_n2848_n452.t11 gnd 0.116496f
C981 a_n2848_n452.n68 gnd 1.0294f
C982 a_n2848_n452.t43 gnd 0.696704f
C983 a_n2848_n452.n69 gnd 0.302425f
C984 a_n2848_n452.t33 gnd 0.696704f
C985 a_n2848_n452.t21 gnd 0.708223f
C986 a_n2848_n452.t75 gnd 0.711378f
C987 a_n2848_n452.t58 gnd 0.696704f
C988 a_n2848_n452.t62 gnd 0.696704f
C989 a_n2848_n452.t52 gnd 0.696704f
C990 a_n2848_n452.n70 gnd 0.306315f
C991 a_n2848_n452.t67 gnd 0.696704f
C992 a_n2848_n452.t73 gnd 0.708223f
C993 a_n2848_n452.t36 gnd 1.40246f
C994 a_n2848_n452.t28 gnd 0.14978f
C995 a_n2848_n452.t24 gnd 0.14978f
C996 a_n2848_n452.n71 gnd 1.05505f
C997 a_n2848_n452.t32 gnd 0.14978f
C998 a_n2848_n452.t40 gnd 0.14978f
C999 a_n2848_n452.n72 gnd 1.05505f
C1000 a_n2848_n452.t30 gnd 1.39967f
C1001 a_n2848_n452.t31 gnd 0.696704f
C1002 a_n2848_n452.n73 gnd 0.306315f
C1003 a_n2848_n452.t39 gnd 0.696704f
C1004 a_n2848_n452.t27 gnd 0.696704f
C1005 a_n2848_n452.t56 gnd 0.696704f
C1006 a_n2848_n452.n74 gnd 0.306315f
C1007 a_n2848_n452.t65 gnd 0.696704f
C1008 a_n2848_n452.t71 gnd 0.696704f
C1009 a_n2848_n452.t70 gnd 0.711378f
C1010 a_n2848_n452.n75 gnd 0.308932f
C1011 a_n2848_n452.t50 gnd 0.696704f
C1012 a_n2848_n452.n76 gnd 0.302425f
C1013 a_n2848_n452.n77 gnd 0.308933f
C1014 a_n2848_n452.t51 gnd 0.708223f
C1015 a_n2848_n452.t35 gnd 0.711378f
C1016 a_n2848_n452.n78 gnd 0.308932f
C1017 a_n2848_n452.t23 gnd 0.696704f
C1018 a_n2848_n452.n79 gnd 0.302425f
C1019 a_n2848_n452.n80 gnd 0.308933f
C1020 a_n2848_n452.t29 gnd 0.708223f
C1021 a_n2848_n452.n81 gnd 1.13204f
C1022 a_n2848_n452.t55 gnd 0.696704f
C1023 a_n2848_n452.n82 gnd 0.302425f
C1024 a_n2848_n452.t61 gnd 0.696704f
C1025 a_n2848_n452.n83 gnd 0.302425f
C1026 a_n2848_n452.t53 gnd 0.696704f
C1027 a_n2848_n452.n84 gnd 0.302425f
C1028 a_n2848_n452.t66 gnd 0.696704f
C1029 a_n2848_n452.n85 gnd 0.302425f
C1030 a_n2848_n452.t57 gnd 0.696704f
C1031 a_n2848_n452.n86 gnd 0.296933f
C1032 a_n2848_n452.t48 gnd 0.696704f
C1033 a_n2848_n452.n87 gnd 0.306315f
C1034 a_n2848_n452.t59 gnd 0.708378f
C1035 a_n2848_n452.t68 gnd 0.696704f
C1036 a_n2848_n452.n88 gnd 0.296933f
C1037 a_n2848_n452.t54 gnd 0.696704f
C1038 a_n2848_n452.n89 gnd 0.306315f
C1039 a_n2848_n452.t63 gnd 0.708378f
C1040 a_n2848_n452.t72 gnd 0.696704f
C1041 a_n2848_n452.n90 gnd 0.296933f
C1042 a_n2848_n452.t60 gnd 0.696704f
C1043 a_n2848_n452.n91 gnd 0.306315f
C1044 a_n2848_n452.t74 gnd 0.708378f
C1045 a_n2848_n452.t64 gnd 0.696704f
C1046 a_n2848_n452.n92 gnd 0.296933f
C1047 a_n2848_n452.t49 gnd 0.696704f
C1048 a_n2848_n452.n93 gnd 0.306315f
C1049 a_n2848_n452.t69 gnd 0.708378f
C1050 a_n2848_n452.n94 gnd 1.33845f
C1051 a_n2848_n452.n95 gnd 0.308933f
C1052 a_n2848_n452.n96 gnd 0.302425f
C1053 a_n2848_n452.n97 gnd 0.308932f
C1054 a_n2848_n452.n98 gnd 0.308933f
C1055 a_n2848_n452.n99 gnd 0.01225f
C1056 a_n2848_n452.n100 gnd 0.302425f
C1057 a_n2848_n452.n101 gnd 0.308933f
C1058 a_n2848_n452.n102 gnd 0.786935f
C1059 a_n2848_n452.t38 gnd 1.39967f
C1060 a_n2848_n452.t42 gnd 0.14978f
C1061 a_n2848_n452.t26 gnd 0.14978f
C1062 a_n2848_n452.n103 gnd 1.05505f
C1063 a_n2848_n452.t44 gnd 0.14978f
C1064 a_n2848_n452.t34 gnd 0.14978f
C1065 a_n2848_n452.n104 gnd 1.05505f
C1066 a_n2848_n452.t22 gnd 1.40246f
C1067 vdd.t122 gnd 0.040594f
C1068 vdd.t8 gnd 0.040594f
C1069 vdd.n0 gnd 0.320175f
C1070 vdd.t293 gnd 0.040594f
C1071 vdd.t285 gnd 0.040594f
C1072 vdd.n1 gnd 0.319647f
C1073 vdd.n2 gnd 0.294775f
C1074 vdd.t118 gnd 0.040594f
C1075 vdd.t6 gnd 0.040594f
C1076 vdd.n3 gnd 0.319647f
C1077 vdd.n4 gnd 0.149079f
C1078 vdd.t13 gnd 0.040594f
C1079 vdd.t287 gnd 0.040594f
C1080 vdd.n5 gnd 0.319647f
C1081 vdd.n6 gnd 0.139883f
C1082 vdd.t295 gnd 0.040594f
C1083 vdd.t120 gnd 0.040594f
C1084 vdd.n7 gnd 0.320175f
C1085 vdd.t2 gnd 0.040594f
C1086 vdd.t15 gnd 0.040594f
C1087 vdd.n8 gnd 0.319647f
C1088 vdd.n9 gnd 0.294775f
C1089 vdd.t289 gnd 0.040594f
C1090 vdd.t115 gnd 0.040594f
C1091 vdd.n10 gnd 0.319647f
C1092 vdd.n11 gnd 0.149079f
C1093 vdd.t112 gnd 0.040594f
C1094 vdd.t291 gnd 0.040594f
C1095 vdd.n12 gnd 0.319647f
C1096 vdd.n13 gnd 0.139883f
C1097 vdd.n14 gnd 0.098895f
C1098 vdd.t24 gnd 0.022552f
C1099 vdd.t23 gnd 0.022552f
C1100 vdd.n15 gnd 0.207586f
C1101 vdd.t19 gnd 0.022552f
C1102 vdd.t25 gnd 0.022552f
C1103 vdd.n16 gnd 0.206979f
C1104 vdd.n17 gnd 0.360208f
C1105 vdd.t20 gnd 0.022552f
C1106 vdd.t21 gnd 0.022552f
C1107 vdd.n18 gnd 0.206979f
C1108 vdd.n19 gnd 0.149023f
C1109 vdd.t26 gnd 0.022552f
C1110 vdd.t22 gnd 0.022552f
C1111 vdd.n20 gnd 0.207586f
C1112 vdd.t29 gnd 0.022552f
C1113 vdd.t17 gnd 0.022552f
C1114 vdd.n21 gnd 0.206979f
C1115 vdd.n22 gnd 0.360208f
C1116 vdd.t31 gnd 0.022552f
C1117 vdd.t30 gnd 0.022552f
C1118 vdd.n23 gnd 0.206979f
C1119 vdd.n24 gnd 0.149023f
C1120 vdd.t32 gnd 0.022552f
C1121 vdd.t27 gnd 0.022552f
C1122 vdd.n25 gnd 0.206979f
C1123 vdd.t28 gnd 0.022552f
C1124 vdd.t18 gnd 0.022552f
C1125 vdd.n26 gnd 0.206979f
C1126 vdd.n27 gnd 23.597301f
C1127 vdd.n28 gnd 8.68612f
C1128 vdd.n29 gnd 0.006151f
C1129 vdd.n30 gnd 0.005708f
C1130 vdd.n31 gnd 0.003157f
C1131 vdd.n32 gnd 0.00725f
C1132 vdd.n33 gnd 0.003067f
C1133 vdd.n34 gnd 0.003248f
C1134 vdd.n35 gnd 0.005708f
C1135 vdd.n36 gnd 0.003067f
C1136 vdd.n37 gnd 0.00725f
C1137 vdd.n38 gnd 0.003248f
C1138 vdd.n39 gnd 0.005708f
C1139 vdd.n40 gnd 0.003067f
C1140 vdd.n41 gnd 0.005437f
C1141 vdd.n42 gnd 0.005453f
C1142 vdd.t126 gnd 0.015575f
C1143 vdd.n43 gnd 0.034655f
C1144 vdd.n44 gnd 0.18035f
C1145 vdd.n45 gnd 0.003067f
C1146 vdd.n46 gnd 0.003248f
C1147 vdd.n47 gnd 0.00725f
C1148 vdd.n48 gnd 0.00725f
C1149 vdd.n49 gnd 0.003248f
C1150 vdd.n50 gnd 0.003067f
C1151 vdd.n51 gnd 0.005708f
C1152 vdd.n52 gnd 0.005708f
C1153 vdd.n53 gnd 0.003067f
C1154 vdd.n54 gnd 0.003248f
C1155 vdd.n55 gnd 0.00725f
C1156 vdd.n56 gnd 0.00725f
C1157 vdd.n57 gnd 0.003248f
C1158 vdd.n58 gnd 0.003067f
C1159 vdd.n59 gnd 0.005708f
C1160 vdd.n60 gnd 0.005708f
C1161 vdd.n61 gnd 0.003067f
C1162 vdd.n62 gnd 0.003248f
C1163 vdd.n63 gnd 0.00725f
C1164 vdd.n64 gnd 0.00725f
C1165 vdd.n65 gnd 0.01714f
C1166 vdd.n66 gnd 0.003157f
C1167 vdd.n67 gnd 0.003067f
C1168 vdd.n68 gnd 0.014753f
C1169 vdd.n69 gnd 0.0103f
C1170 vdd.t266 gnd 0.036084f
C1171 vdd.t207 gnd 0.036084f
C1172 vdd.n70 gnd 0.247994f
C1173 vdd.n71 gnd 0.195009f
C1174 vdd.t280 gnd 0.036084f
C1175 vdd.t174 gnd 0.036084f
C1176 vdd.n72 gnd 0.247994f
C1177 vdd.n73 gnd 0.157371f
C1178 vdd.t252 gnd 0.036084f
C1179 vdd.t198 gnd 0.036084f
C1180 vdd.n74 gnd 0.247994f
C1181 vdd.n75 gnd 0.157371f
C1182 vdd.t274 gnd 0.036084f
C1183 vdd.t247 gnd 0.036084f
C1184 vdd.n76 gnd 0.247994f
C1185 vdd.n77 gnd 0.157371f
C1186 vdd.t138 gnd 0.036084f
C1187 vdd.t187 gnd 0.036084f
C1188 vdd.n78 gnd 0.247994f
C1189 vdd.n79 gnd 0.157371f
C1190 vdd.t148 gnd 0.036084f
C1191 vdd.t209 gnd 0.036084f
C1192 vdd.n80 gnd 0.247994f
C1193 vdd.n81 gnd 0.157371f
C1194 vdd.t180 gnd 0.036084f
C1195 vdd.t259 gnd 0.036084f
C1196 vdd.n82 gnd 0.247994f
C1197 vdd.n83 gnd 0.157371f
C1198 vdd.t152 gnd 0.036084f
C1199 vdd.t232 gnd 0.036084f
C1200 vdd.n84 gnd 0.247994f
C1201 vdd.n85 gnd 0.157371f
C1202 vdd.t164 gnd 0.036084f
C1203 vdd.t249 gnd 0.036084f
C1204 vdd.n86 gnd 0.247994f
C1205 vdd.n87 gnd 0.157371f
C1206 vdd.n88 gnd 0.006151f
C1207 vdd.n89 gnd 0.005708f
C1208 vdd.n90 gnd 0.003157f
C1209 vdd.n91 gnd 0.00725f
C1210 vdd.n92 gnd 0.003067f
C1211 vdd.n93 gnd 0.003248f
C1212 vdd.n94 gnd 0.005708f
C1213 vdd.n95 gnd 0.003067f
C1214 vdd.n96 gnd 0.00725f
C1215 vdd.n97 gnd 0.003248f
C1216 vdd.n98 gnd 0.005708f
C1217 vdd.n99 gnd 0.003067f
C1218 vdd.n100 gnd 0.005437f
C1219 vdd.n101 gnd 0.005453f
C1220 vdd.t190 gnd 0.015575f
C1221 vdd.n102 gnd 0.034655f
C1222 vdd.n103 gnd 0.18035f
C1223 vdd.n104 gnd 0.003067f
C1224 vdd.n105 gnd 0.003248f
C1225 vdd.n106 gnd 0.00725f
C1226 vdd.n107 gnd 0.00725f
C1227 vdd.n108 gnd 0.003248f
C1228 vdd.n109 gnd 0.003067f
C1229 vdd.n110 gnd 0.005708f
C1230 vdd.n111 gnd 0.005708f
C1231 vdd.n112 gnd 0.003067f
C1232 vdd.n113 gnd 0.003248f
C1233 vdd.n114 gnd 0.00725f
C1234 vdd.n115 gnd 0.00725f
C1235 vdd.n116 gnd 0.003248f
C1236 vdd.n117 gnd 0.003067f
C1237 vdd.n118 gnd 0.005708f
C1238 vdd.n119 gnd 0.005708f
C1239 vdd.n120 gnd 0.003067f
C1240 vdd.n121 gnd 0.003248f
C1241 vdd.n122 gnd 0.00725f
C1242 vdd.n123 gnd 0.00725f
C1243 vdd.n124 gnd 0.01714f
C1244 vdd.n125 gnd 0.003157f
C1245 vdd.n126 gnd 0.003067f
C1246 vdd.n127 gnd 0.014753f
C1247 vdd.n128 gnd 0.009977f
C1248 vdd.n129 gnd 0.117085f
C1249 vdd.n130 gnd 0.006151f
C1250 vdd.n131 gnd 0.005708f
C1251 vdd.n132 gnd 0.003157f
C1252 vdd.n133 gnd 0.00725f
C1253 vdd.n134 gnd 0.003067f
C1254 vdd.n135 gnd 0.003248f
C1255 vdd.n136 gnd 0.005708f
C1256 vdd.n137 gnd 0.003067f
C1257 vdd.n138 gnd 0.00725f
C1258 vdd.n139 gnd 0.003248f
C1259 vdd.n140 gnd 0.005708f
C1260 vdd.n141 gnd 0.003067f
C1261 vdd.n142 gnd 0.005437f
C1262 vdd.n143 gnd 0.005453f
C1263 vdd.t212 gnd 0.015575f
C1264 vdd.n144 gnd 0.034655f
C1265 vdd.n145 gnd 0.18035f
C1266 vdd.n146 gnd 0.003067f
C1267 vdd.n147 gnd 0.003248f
C1268 vdd.n148 gnd 0.00725f
C1269 vdd.n149 gnd 0.00725f
C1270 vdd.n150 gnd 0.003248f
C1271 vdd.n151 gnd 0.003067f
C1272 vdd.n152 gnd 0.005708f
C1273 vdd.n153 gnd 0.005708f
C1274 vdd.n154 gnd 0.003067f
C1275 vdd.n155 gnd 0.003248f
C1276 vdd.n156 gnd 0.00725f
C1277 vdd.n157 gnd 0.00725f
C1278 vdd.n158 gnd 0.003248f
C1279 vdd.n159 gnd 0.003067f
C1280 vdd.n160 gnd 0.005708f
C1281 vdd.n161 gnd 0.005708f
C1282 vdd.n162 gnd 0.003067f
C1283 vdd.n163 gnd 0.003248f
C1284 vdd.n164 gnd 0.00725f
C1285 vdd.n165 gnd 0.00725f
C1286 vdd.n166 gnd 0.01714f
C1287 vdd.n167 gnd 0.003157f
C1288 vdd.n168 gnd 0.003067f
C1289 vdd.n169 gnd 0.014753f
C1290 vdd.n170 gnd 0.0103f
C1291 vdd.t214 gnd 0.036084f
C1292 vdd.t243 gnd 0.036084f
C1293 vdd.n171 gnd 0.247994f
C1294 vdd.n172 gnd 0.195009f
C1295 vdd.t134 gnd 0.036084f
C1296 vdd.t202 gnd 0.036084f
C1297 vdd.n173 gnd 0.247994f
C1298 vdd.n174 gnd 0.157371f
C1299 vdd.t240 gnd 0.036084f
C1300 vdd.t282 gnd 0.036084f
C1301 vdd.n175 gnd 0.247994f
C1302 vdd.n176 gnd 0.157371f
C1303 vdd.t182 gnd 0.036084f
C1304 vdd.t184 gnd 0.036084f
C1305 vdd.n177 gnd 0.247994f
C1306 vdd.n178 gnd 0.157371f
C1307 vdd.t268 gnd 0.036084f
C1308 vdd.t177 gnd 0.036084f
C1309 vdd.n179 gnd 0.247994f
C1310 vdd.n180 gnd 0.157371f
C1311 vdd.t178 gnd 0.036084f
C1312 vdd.t264 gnd 0.036084f
C1313 vdd.n181 gnd 0.247994f
C1314 vdd.n182 gnd 0.157371f
C1315 vdd.t265 gnd 0.036084f
C1316 vdd.t146 gnd 0.036084f
C1317 vdd.n183 gnd 0.247994f
C1318 vdd.n184 gnd 0.157371f
C1319 vdd.t242 gnd 0.036084f
C1320 vdd.t262 gnd 0.036084f
C1321 vdd.n185 gnd 0.247994f
C1322 vdd.n186 gnd 0.157371f
C1323 vdd.t144 gnd 0.036084f
C1324 vdd.t204 gnd 0.036084f
C1325 vdd.n187 gnd 0.247994f
C1326 vdd.n188 gnd 0.157371f
C1327 vdd.n189 gnd 0.006151f
C1328 vdd.n190 gnd 0.005708f
C1329 vdd.n191 gnd 0.003157f
C1330 vdd.n192 gnd 0.00725f
C1331 vdd.n193 gnd 0.003067f
C1332 vdd.n194 gnd 0.003248f
C1333 vdd.n195 gnd 0.005708f
C1334 vdd.n196 gnd 0.003067f
C1335 vdd.n197 gnd 0.00725f
C1336 vdd.n198 gnd 0.003248f
C1337 vdd.n199 gnd 0.005708f
C1338 vdd.n200 gnd 0.003067f
C1339 vdd.n201 gnd 0.005437f
C1340 vdd.n202 gnd 0.005453f
C1341 vdd.t241 gnd 0.015575f
C1342 vdd.n203 gnd 0.034655f
C1343 vdd.n204 gnd 0.18035f
C1344 vdd.n205 gnd 0.003067f
C1345 vdd.n206 gnd 0.003248f
C1346 vdd.n207 gnd 0.00725f
C1347 vdd.n208 gnd 0.00725f
C1348 vdd.n209 gnd 0.003248f
C1349 vdd.n210 gnd 0.003067f
C1350 vdd.n211 gnd 0.005708f
C1351 vdd.n212 gnd 0.005708f
C1352 vdd.n213 gnd 0.003067f
C1353 vdd.n214 gnd 0.003248f
C1354 vdd.n215 gnd 0.00725f
C1355 vdd.n216 gnd 0.00725f
C1356 vdd.n217 gnd 0.003248f
C1357 vdd.n218 gnd 0.003067f
C1358 vdd.n219 gnd 0.005708f
C1359 vdd.n220 gnd 0.005708f
C1360 vdd.n221 gnd 0.003067f
C1361 vdd.n222 gnd 0.003248f
C1362 vdd.n223 gnd 0.00725f
C1363 vdd.n224 gnd 0.00725f
C1364 vdd.n225 gnd 0.01714f
C1365 vdd.n226 gnd 0.003157f
C1366 vdd.n227 gnd 0.003067f
C1367 vdd.n228 gnd 0.014753f
C1368 vdd.n229 gnd 0.009977f
C1369 vdd.n230 gnd 0.069654f
C1370 vdd.n231 gnd 0.250981f
C1371 vdd.n232 gnd 0.006151f
C1372 vdd.n233 gnd 0.005708f
C1373 vdd.n234 gnd 0.003157f
C1374 vdd.n235 gnd 0.00725f
C1375 vdd.n236 gnd 0.003067f
C1376 vdd.n237 gnd 0.003248f
C1377 vdd.n238 gnd 0.005708f
C1378 vdd.n239 gnd 0.003067f
C1379 vdd.n240 gnd 0.00725f
C1380 vdd.n241 gnd 0.003248f
C1381 vdd.n242 gnd 0.005708f
C1382 vdd.n243 gnd 0.003067f
C1383 vdd.n244 gnd 0.005437f
C1384 vdd.n245 gnd 0.005453f
C1385 vdd.t226 gnd 0.015575f
C1386 vdd.n246 gnd 0.034655f
C1387 vdd.n247 gnd 0.18035f
C1388 vdd.n248 gnd 0.003067f
C1389 vdd.n249 gnd 0.003248f
C1390 vdd.n250 gnd 0.00725f
C1391 vdd.n251 gnd 0.00725f
C1392 vdd.n252 gnd 0.003248f
C1393 vdd.n253 gnd 0.003067f
C1394 vdd.n254 gnd 0.005708f
C1395 vdd.n255 gnd 0.005708f
C1396 vdd.n256 gnd 0.003067f
C1397 vdd.n257 gnd 0.003248f
C1398 vdd.n258 gnd 0.00725f
C1399 vdd.n259 gnd 0.00725f
C1400 vdd.n260 gnd 0.003248f
C1401 vdd.n261 gnd 0.003067f
C1402 vdd.n262 gnd 0.005708f
C1403 vdd.n263 gnd 0.005708f
C1404 vdd.n264 gnd 0.003067f
C1405 vdd.n265 gnd 0.003248f
C1406 vdd.n266 gnd 0.00725f
C1407 vdd.n267 gnd 0.00725f
C1408 vdd.n268 gnd 0.01714f
C1409 vdd.n269 gnd 0.003157f
C1410 vdd.n270 gnd 0.003067f
C1411 vdd.n271 gnd 0.014753f
C1412 vdd.n272 gnd 0.0103f
C1413 vdd.t227 gnd 0.036084f
C1414 vdd.t257 gnd 0.036084f
C1415 vdd.n273 gnd 0.247994f
C1416 vdd.n274 gnd 0.195009f
C1417 vdd.t159 gnd 0.036084f
C1418 vdd.t223 gnd 0.036084f
C1419 vdd.n275 gnd 0.247994f
C1420 vdd.n276 gnd 0.157371f
C1421 vdd.t251 gnd 0.036084f
C1422 vdd.t154 gnd 0.036084f
C1423 vdd.n277 gnd 0.247994f
C1424 vdd.n278 gnd 0.157371f
C1425 vdd.t199 gnd 0.036084f
C1426 vdd.t201 gnd 0.036084f
C1427 vdd.n279 gnd 0.247994f
C1428 vdd.n280 gnd 0.157371f
C1429 vdd.t278 gnd 0.036084f
C1430 vdd.t194 gnd 0.036084f
C1431 vdd.n281 gnd 0.247994f
C1432 vdd.n282 gnd 0.157371f
C1433 vdd.t195 gnd 0.036084f
C1434 vdd.t276 gnd 0.036084f
C1435 vdd.n283 gnd 0.247994f
C1436 vdd.n284 gnd 0.157371f
C1437 vdd.t277 gnd 0.036084f
C1438 vdd.t170 gnd 0.036084f
C1439 vdd.n285 gnd 0.247994f
C1440 vdd.n286 gnd 0.157371f
C1441 vdd.t258 gnd 0.036084f
C1442 vdd.t275 gnd 0.036084f
C1443 vdd.n287 gnd 0.247994f
C1444 vdd.n288 gnd 0.157371f
C1445 vdd.t167 gnd 0.036084f
C1446 vdd.t224 gnd 0.036084f
C1447 vdd.n289 gnd 0.247994f
C1448 vdd.n290 gnd 0.157371f
C1449 vdd.n291 gnd 0.006151f
C1450 vdd.n292 gnd 0.005708f
C1451 vdd.n293 gnd 0.003157f
C1452 vdd.n294 gnd 0.00725f
C1453 vdd.n295 gnd 0.003067f
C1454 vdd.n296 gnd 0.003248f
C1455 vdd.n297 gnd 0.005708f
C1456 vdd.n298 gnd 0.003067f
C1457 vdd.n299 gnd 0.00725f
C1458 vdd.n300 gnd 0.003248f
C1459 vdd.n301 gnd 0.005708f
C1460 vdd.n302 gnd 0.003067f
C1461 vdd.n303 gnd 0.005437f
C1462 vdd.n304 gnd 0.005453f
C1463 vdd.t254 gnd 0.015575f
C1464 vdd.n305 gnd 0.034655f
C1465 vdd.n306 gnd 0.18035f
C1466 vdd.n307 gnd 0.003067f
C1467 vdd.n308 gnd 0.003248f
C1468 vdd.n309 gnd 0.00725f
C1469 vdd.n310 gnd 0.00725f
C1470 vdd.n311 gnd 0.003248f
C1471 vdd.n312 gnd 0.003067f
C1472 vdd.n313 gnd 0.005708f
C1473 vdd.n314 gnd 0.005708f
C1474 vdd.n315 gnd 0.003067f
C1475 vdd.n316 gnd 0.003248f
C1476 vdd.n317 gnd 0.00725f
C1477 vdd.n318 gnd 0.00725f
C1478 vdd.n319 gnd 0.003248f
C1479 vdd.n320 gnd 0.003067f
C1480 vdd.n321 gnd 0.005708f
C1481 vdd.n322 gnd 0.005708f
C1482 vdd.n323 gnd 0.003067f
C1483 vdd.n324 gnd 0.003248f
C1484 vdd.n325 gnd 0.00725f
C1485 vdd.n326 gnd 0.00725f
C1486 vdd.n327 gnd 0.01714f
C1487 vdd.n328 gnd 0.003157f
C1488 vdd.n329 gnd 0.003067f
C1489 vdd.n330 gnd 0.014753f
C1490 vdd.n331 gnd 0.009977f
C1491 vdd.n332 gnd 0.069654f
C1492 vdd.n333 gnd 0.287319f
C1493 vdd.n334 gnd 0.008614f
C1494 vdd.n335 gnd 0.011208f
C1495 vdd.n336 gnd 0.009021f
C1496 vdd.n337 gnd 0.009021f
C1497 vdd.n338 gnd 0.011208f
C1498 vdd.n339 gnd 0.011208f
C1499 vdd.n340 gnd 0.818956f
C1500 vdd.n341 gnd 0.011208f
C1501 vdd.n342 gnd 0.011208f
C1502 vdd.n343 gnd 0.011208f
C1503 vdd.n344 gnd 0.88768f
C1504 vdd.n345 gnd 0.011208f
C1505 vdd.n346 gnd 0.011208f
C1506 vdd.n347 gnd 0.011208f
C1507 vdd.n348 gnd 0.011208f
C1508 vdd.n349 gnd 0.009021f
C1509 vdd.n350 gnd 0.011208f
C1510 vdd.t208 gnd 0.572697f
C1511 vdd.n351 gnd 0.011208f
C1512 vdd.n352 gnd 0.011208f
C1513 vdd.n353 gnd 0.011208f
C1514 vdd.t145 gnd 0.572697f
C1515 vdd.n354 gnd 0.011208f
C1516 vdd.n355 gnd 0.011208f
C1517 vdd.n356 gnd 0.011208f
C1518 vdd.n357 gnd 0.011208f
C1519 vdd.n358 gnd 0.011208f
C1520 vdd.n359 gnd 0.009021f
C1521 vdd.n360 gnd 0.011208f
C1522 vdd.n361 gnd 0.647147f
C1523 vdd.n362 gnd 0.011208f
C1524 vdd.n363 gnd 0.011208f
C1525 vdd.n364 gnd 0.011208f
C1526 vdd.t231 gnd 0.572697f
C1527 vdd.n365 gnd 0.011208f
C1528 vdd.n366 gnd 0.011208f
C1529 vdd.n367 gnd 0.011208f
C1530 vdd.n368 gnd 0.011208f
C1531 vdd.n369 gnd 0.011208f
C1532 vdd.n370 gnd 0.009021f
C1533 vdd.n371 gnd 0.011208f
C1534 vdd.t143 gnd 0.572697f
C1535 vdd.n372 gnd 0.011208f
C1536 vdd.n373 gnd 0.011208f
C1537 vdd.n374 gnd 0.011208f
C1538 vdd.n375 gnd 0.670055f
C1539 vdd.n376 gnd 0.011208f
C1540 vdd.n377 gnd 0.011208f
C1541 vdd.n378 gnd 0.011208f
C1542 vdd.n379 gnd 0.011208f
C1543 vdd.n380 gnd 0.011208f
C1544 vdd.n381 gnd 0.009021f
C1545 vdd.n382 gnd 0.011208f
C1546 vdd.t189 gnd 0.572697f
C1547 vdd.n383 gnd 0.011208f
C1548 vdd.n384 gnd 0.011208f
C1549 vdd.n385 gnd 0.011208f
C1550 vdd.n386 gnd 0.578424f
C1551 vdd.n387 gnd 0.011208f
C1552 vdd.n388 gnd 0.011208f
C1553 vdd.n389 gnd 0.011208f
C1554 vdd.n390 gnd 0.011208f
C1555 vdd.n391 gnd 0.027113f
C1556 vdd.n392 gnd 0.027694f
C1557 vdd.t57 gnd 0.572697f
C1558 vdd.n393 gnd 0.027113f
C1559 vdd.n425 gnd 0.011208f
C1560 vdd.t59 gnd 0.137886f
C1561 vdd.t58 gnd 0.147363f
C1562 vdd.t56 gnd 0.180078f
C1563 vdd.n426 gnd 0.230835f
C1564 vdd.n427 gnd 0.194845f
C1565 vdd.n428 gnd 0.014794f
C1566 vdd.n429 gnd 0.011208f
C1567 vdd.n430 gnd 0.009021f
C1568 vdd.n431 gnd 0.011208f
C1569 vdd.n432 gnd 0.009021f
C1570 vdd.n433 gnd 0.011208f
C1571 vdd.n434 gnd 0.009021f
C1572 vdd.n435 gnd 0.011208f
C1573 vdd.n436 gnd 0.009021f
C1574 vdd.n437 gnd 0.011208f
C1575 vdd.n438 gnd 0.009021f
C1576 vdd.n439 gnd 0.011208f
C1577 vdd.t100 gnd 0.137886f
C1578 vdd.t99 gnd 0.147363f
C1579 vdd.t98 gnd 0.180078f
C1580 vdd.n440 gnd 0.230835f
C1581 vdd.n441 gnd 0.194845f
C1582 vdd.n442 gnd 0.009021f
C1583 vdd.n443 gnd 0.011208f
C1584 vdd.n444 gnd 0.009021f
C1585 vdd.n445 gnd 0.011208f
C1586 vdd.n446 gnd 0.009021f
C1587 vdd.n447 gnd 0.011208f
C1588 vdd.n448 gnd 0.009021f
C1589 vdd.n449 gnd 0.011208f
C1590 vdd.n450 gnd 0.009021f
C1591 vdd.n451 gnd 0.011208f
C1592 vdd.t106 gnd 0.137886f
C1593 vdd.t105 gnd 0.147363f
C1594 vdd.t104 gnd 0.180078f
C1595 vdd.n452 gnd 0.230835f
C1596 vdd.n453 gnd 0.194845f
C1597 vdd.n454 gnd 0.019305f
C1598 vdd.n455 gnd 0.011208f
C1599 vdd.n456 gnd 0.009021f
C1600 vdd.n457 gnd 0.011208f
C1601 vdd.n458 gnd 0.009021f
C1602 vdd.n459 gnd 0.011208f
C1603 vdd.n460 gnd 0.009021f
C1604 vdd.n461 gnd 0.011208f
C1605 vdd.n462 gnd 0.009021f
C1606 vdd.n463 gnd 0.011208f
C1607 vdd.n464 gnd 0.027694f
C1608 vdd.n465 gnd 0.007487f
C1609 vdd.n466 gnd 0.009021f
C1610 vdd.n467 gnd 0.011208f
C1611 vdd.n468 gnd 0.011208f
C1612 vdd.n469 gnd 0.009021f
C1613 vdd.n470 gnd 0.011208f
C1614 vdd.n471 gnd 0.011208f
C1615 vdd.n472 gnd 0.011208f
C1616 vdd.n473 gnd 0.011208f
C1617 vdd.n474 gnd 0.011208f
C1618 vdd.n475 gnd 0.009021f
C1619 vdd.n476 gnd 0.009021f
C1620 vdd.n477 gnd 0.011208f
C1621 vdd.n478 gnd 0.011208f
C1622 vdd.n479 gnd 0.009021f
C1623 vdd.n480 gnd 0.011208f
C1624 vdd.n481 gnd 0.011208f
C1625 vdd.n482 gnd 0.011208f
C1626 vdd.n483 gnd 0.011208f
C1627 vdd.n484 gnd 0.011208f
C1628 vdd.n485 gnd 0.009021f
C1629 vdd.n486 gnd 0.009021f
C1630 vdd.n487 gnd 0.011208f
C1631 vdd.n488 gnd 0.011208f
C1632 vdd.n489 gnd 0.009021f
C1633 vdd.n490 gnd 0.011208f
C1634 vdd.n491 gnd 0.011208f
C1635 vdd.n492 gnd 0.011208f
C1636 vdd.n493 gnd 0.011208f
C1637 vdd.n494 gnd 0.011208f
C1638 vdd.n495 gnd 0.009021f
C1639 vdd.n496 gnd 0.009021f
C1640 vdd.n497 gnd 0.011208f
C1641 vdd.n498 gnd 0.011208f
C1642 vdd.n499 gnd 0.009021f
C1643 vdd.n500 gnd 0.011208f
C1644 vdd.n501 gnd 0.011208f
C1645 vdd.n502 gnd 0.011208f
C1646 vdd.n503 gnd 0.011208f
C1647 vdd.n504 gnd 0.011208f
C1648 vdd.n505 gnd 0.009021f
C1649 vdd.n506 gnd 0.009021f
C1650 vdd.n507 gnd 0.011208f
C1651 vdd.n508 gnd 0.011208f
C1652 vdd.n509 gnd 0.007533f
C1653 vdd.n510 gnd 0.011208f
C1654 vdd.n511 gnd 0.011208f
C1655 vdd.n512 gnd 0.011208f
C1656 vdd.n513 gnd 0.011208f
C1657 vdd.n514 gnd 0.011208f
C1658 vdd.n515 gnd 0.007533f
C1659 vdd.n516 gnd 0.009021f
C1660 vdd.n517 gnd 0.011208f
C1661 vdd.n518 gnd 0.011208f
C1662 vdd.n519 gnd 0.009021f
C1663 vdd.n520 gnd 0.011208f
C1664 vdd.n521 gnd 0.011208f
C1665 vdd.n522 gnd 0.011208f
C1666 vdd.n523 gnd 0.011208f
C1667 vdd.n524 gnd 0.011208f
C1668 vdd.n525 gnd 0.009021f
C1669 vdd.n526 gnd 0.009021f
C1670 vdd.n527 gnd 0.011208f
C1671 vdd.n528 gnd 0.011208f
C1672 vdd.n529 gnd 0.009021f
C1673 vdd.n530 gnd 0.011208f
C1674 vdd.n531 gnd 0.011208f
C1675 vdd.n532 gnd 0.011208f
C1676 vdd.n533 gnd 0.011208f
C1677 vdd.n534 gnd 0.011208f
C1678 vdd.n535 gnd 0.009021f
C1679 vdd.n536 gnd 0.009021f
C1680 vdd.n537 gnd 0.011208f
C1681 vdd.n538 gnd 0.011208f
C1682 vdd.n539 gnd 0.009021f
C1683 vdd.n540 gnd 0.011208f
C1684 vdd.n541 gnd 0.011208f
C1685 vdd.n542 gnd 0.011208f
C1686 vdd.n543 gnd 0.011208f
C1687 vdd.n544 gnd 0.011208f
C1688 vdd.n545 gnd 0.009021f
C1689 vdd.n546 gnd 0.009021f
C1690 vdd.n547 gnd 0.011208f
C1691 vdd.n548 gnd 0.011208f
C1692 vdd.n549 gnd 0.009021f
C1693 vdd.n550 gnd 0.011208f
C1694 vdd.n551 gnd 0.011208f
C1695 vdd.n552 gnd 0.011208f
C1696 vdd.n553 gnd 0.011208f
C1697 vdd.n554 gnd 0.011208f
C1698 vdd.n555 gnd 0.009021f
C1699 vdd.n556 gnd 0.009021f
C1700 vdd.n557 gnd 0.011208f
C1701 vdd.n558 gnd 0.011208f
C1702 vdd.n559 gnd 0.009021f
C1703 vdd.n560 gnd 0.011208f
C1704 vdd.n561 gnd 0.011208f
C1705 vdd.n562 gnd 0.011208f
C1706 vdd.n563 gnd 0.011208f
C1707 vdd.n564 gnd 0.011208f
C1708 vdd.n565 gnd 0.006134f
C1709 vdd.n566 gnd 0.019305f
C1710 vdd.n567 gnd 0.011208f
C1711 vdd.n568 gnd 0.011208f
C1712 vdd.n569 gnd 0.008931f
C1713 vdd.n570 gnd 0.011208f
C1714 vdd.n571 gnd 0.011208f
C1715 vdd.n572 gnd 0.011208f
C1716 vdd.n573 gnd 0.011208f
C1717 vdd.n574 gnd 0.011208f
C1718 vdd.n575 gnd 0.009021f
C1719 vdd.n576 gnd 0.009021f
C1720 vdd.n577 gnd 0.011208f
C1721 vdd.n578 gnd 0.011208f
C1722 vdd.n579 gnd 0.009021f
C1723 vdd.n580 gnd 0.011208f
C1724 vdd.n581 gnd 0.011208f
C1725 vdd.n582 gnd 0.011208f
C1726 vdd.n583 gnd 0.011208f
C1727 vdd.n584 gnd 0.011208f
C1728 vdd.n585 gnd 0.009021f
C1729 vdd.n586 gnd 0.009021f
C1730 vdd.n587 gnd 0.011208f
C1731 vdd.n588 gnd 0.011208f
C1732 vdd.n589 gnd 0.009021f
C1733 vdd.n590 gnd 0.011208f
C1734 vdd.n591 gnd 0.011208f
C1735 vdd.n592 gnd 0.011208f
C1736 vdd.n593 gnd 0.011208f
C1737 vdd.n594 gnd 0.011208f
C1738 vdd.n595 gnd 0.009021f
C1739 vdd.n596 gnd 0.009021f
C1740 vdd.n597 gnd 0.011208f
C1741 vdd.n598 gnd 0.011208f
C1742 vdd.n599 gnd 0.009021f
C1743 vdd.n600 gnd 0.011208f
C1744 vdd.n601 gnd 0.011208f
C1745 vdd.n602 gnd 0.011208f
C1746 vdd.n603 gnd 0.011208f
C1747 vdd.n604 gnd 0.011208f
C1748 vdd.n605 gnd 0.009021f
C1749 vdd.n606 gnd 0.009021f
C1750 vdd.n607 gnd 0.011208f
C1751 vdd.n608 gnd 0.011208f
C1752 vdd.n609 gnd 0.009021f
C1753 vdd.n610 gnd 0.011208f
C1754 vdd.n611 gnd 0.011208f
C1755 vdd.n612 gnd 0.011208f
C1756 vdd.n613 gnd 0.011208f
C1757 vdd.n614 gnd 0.011208f
C1758 vdd.n615 gnd 0.009021f
C1759 vdd.n616 gnd 0.011208f
C1760 vdd.n617 gnd 0.009021f
C1761 vdd.n618 gnd 0.004736f
C1762 vdd.n619 gnd 0.011208f
C1763 vdd.n620 gnd 0.011208f
C1764 vdd.n621 gnd 0.009021f
C1765 vdd.n622 gnd 0.011208f
C1766 vdd.n623 gnd 0.009021f
C1767 vdd.n624 gnd 0.011208f
C1768 vdd.n625 gnd 0.009021f
C1769 vdd.n626 gnd 0.011208f
C1770 vdd.n627 gnd 0.009021f
C1771 vdd.n628 gnd 0.011208f
C1772 vdd.n629 gnd 0.009021f
C1773 vdd.n630 gnd 0.011208f
C1774 vdd.n631 gnd 0.009021f
C1775 vdd.n632 gnd 0.011208f
C1776 vdd.n633 gnd 0.624239f
C1777 vdd.t137 gnd 0.572697f
C1778 vdd.n634 gnd 0.011208f
C1779 vdd.n635 gnd 0.009021f
C1780 vdd.n636 gnd 0.011208f
C1781 vdd.n637 gnd 0.009021f
C1782 vdd.n638 gnd 0.011208f
C1783 vdd.t181 gnd 0.572697f
C1784 vdd.n639 gnd 0.011208f
C1785 vdd.n640 gnd 0.009021f
C1786 vdd.n641 gnd 0.011208f
C1787 vdd.n642 gnd 0.009021f
C1788 vdd.n643 gnd 0.011208f
C1789 vdd.t153 gnd 0.572697f
C1790 vdd.n644 gnd 0.715871f
C1791 vdd.n645 gnd 0.011208f
C1792 vdd.n646 gnd 0.009021f
C1793 vdd.n647 gnd 0.011208f
C1794 vdd.n648 gnd 0.009021f
C1795 vdd.n649 gnd 0.011208f
C1796 vdd.t239 gnd 0.572697f
C1797 vdd.n650 gnd 0.011208f
C1798 vdd.n651 gnd 0.009021f
C1799 vdd.n652 gnd 0.011208f
C1800 vdd.n653 gnd 0.009021f
C1801 vdd.n654 gnd 0.011208f
C1802 vdd.n655 gnd 0.796048f
C1803 vdd.n656 gnd 0.950677f
C1804 vdd.t173 gnd 0.572697f
C1805 vdd.n657 gnd 0.011208f
C1806 vdd.n658 gnd 0.009021f
C1807 vdd.n659 gnd 0.011208f
C1808 vdd.n660 gnd 0.009021f
C1809 vdd.n661 gnd 0.011208f
C1810 vdd.n662 gnd 0.601332f
C1811 vdd.n663 gnd 0.011208f
C1812 vdd.n664 gnd 0.009021f
C1813 vdd.n665 gnd 0.011208f
C1814 vdd.n666 gnd 0.009021f
C1815 vdd.n667 gnd 0.011208f
C1816 vdd.t213 gnd 0.572697f
C1817 vdd.t206 gnd 0.572697f
C1818 vdd.n668 gnd 0.011208f
C1819 vdd.n669 gnd 0.009021f
C1820 vdd.n670 gnd 0.011208f
C1821 vdd.n671 gnd 0.009021f
C1822 vdd.n672 gnd 0.011208f
C1823 vdd.t125 gnd 0.572697f
C1824 vdd.n673 gnd 0.011208f
C1825 vdd.n674 gnd 0.009021f
C1826 vdd.n675 gnd 0.011208f
C1827 vdd.n676 gnd 0.009021f
C1828 vdd.n677 gnd 0.011208f
C1829 vdd.n678 gnd 1.14539f
C1830 vdd.n679 gnd 0.933496f
C1831 vdd.n680 gnd 0.011208f
C1832 vdd.n681 gnd 0.009021f
C1833 vdd.n682 gnd 0.027113f
C1834 vdd.n683 gnd 0.007487f
C1835 vdd.n684 gnd 0.027113f
C1836 vdd.t35 gnd 0.572697f
C1837 vdd.n685 gnd 0.027113f
C1838 vdd.n686 gnd 0.007487f
C1839 vdd.n687 gnd 0.009639f
C1840 vdd.t102 gnd 0.137886f
C1841 vdd.t103 gnd 0.147363f
C1842 vdd.t101 gnd 0.180078f
C1843 vdd.n688 gnd 0.230835f
C1844 vdd.n689 gnd 0.193943f
C1845 vdd.n690 gnd 0.013892f
C1846 vdd.n691 gnd 0.011208f
C1847 vdd.n692 gnd 7.891759f
C1848 vdd.n723 gnd 1.57492f
C1849 vdd.n724 gnd 0.011208f
C1850 vdd.n725 gnd 0.011208f
C1851 vdd.n726 gnd 0.027694f
C1852 vdd.n727 gnd 0.009639f
C1853 vdd.n728 gnd 0.011208f
C1854 vdd.n729 gnd 0.009021f
C1855 vdd.n730 gnd 0.007173f
C1856 vdd.n731 gnd 0.018314f
C1857 vdd.n732 gnd 0.009021f
C1858 vdd.n733 gnd 0.011208f
C1859 vdd.n734 gnd 0.011208f
C1860 vdd.n735 gnd 0.011208f
C1861 vdd.n736 gnd 0.011208f
C1862 vdd.n737 gnd 0.011208f
C1863 vdd.n738 gnd 0.011208f
C1864 vdd.n739 gnd 0.011208f
C1865 vdd.n740 gnd 0.011208f
C1866 vdd.n741 gnd 0.011208f
C1867 vdd.n742 gnd 0.011208f
C1868 vdd.n743 gnd 0.011208f
C1869 vdd.n744 gnd 0.011208f
C1870 vdd.n745 gnd 0.011208f
C1871 vdd.n746 gnd 0.011208f
C1872 vdd.n747 gnd 0.007533f
C1873 vdd.n748 gnd 0.011208f
C1874 vdd.n749 gnd 0.011208f
C1875 vdd.n750 gnd 0.011208f
C1876 vdd.n751 gnd 0.011208f
C1877 vdd.n752 gnd 0.011208f
C1878 vdd.n753 gnd 0.011208f
C1879 vdd.n754 gnd 0.011208f
C1880 vdd.n755 gnd 0.011208f
C1881 vdd.n756 gnd 0.011208f
C1882 vdd.n757 gnd 0.011208f
C1883 vdd.n758 gnd 0.011208f
C1884 vdd.n759 gnd 0.011208f
C1885 vdd.n760 gnd 0.011208f
C1886 vdd.n761 gnd 0.011208f
C1887 vdd.n762 gnd 0.011208f
C1888 vdd.n763 gnd 0.011208f
C1889 vdd.n764 gnd 0.011208f
C1890 vdd.n765 gnd 0.011208f
C1891 vdd.n766 gnd 0.011208f
C1892 vdd.n767 gnd 0.008931f
C1893 vdd.t36 gnd 0.137886f
C1894 vdd.t37 gnd 0.147363f
C1895 vdd.t34 gnd 0.180078f
C1896 vdd.n768 gnd 0.230835f
C1897 vdd.n769 gnd 0.193943f
C1898 vdd.n770 gnd 0.011208f
C1899 vdd.n771 gnd 0.011208f
C1900 vdd.n772 gnd 0.011208f
C1901 vdd.n773 gnd 0.011208f
C1902 vdd.n774 gnd 0.011208f
C1903 vdd.n775 gnd 0.011208f
C1904 vdd.n776 gnd 0.011208f
C1905 vdd.n777 gnd 0.011208f
C1906 vdd.n778 gnd 0.011208f
C1907 vdd.n779 gnd 0.011208f
C1908 vdd.n780 gnd 0.011208f
C1909 vdd.n781 gnd 0.011208f
C1910 vdd.n782 gnd 0.011208f
C1911 vdd.n783 gnd 0.007173f
C1912 vdd.n785 gnd 0.007621f
C1913 vdd.n786 gnd 0.007621f
C1914 vdd.n787 gnd 0.007621f
C1915 vdd.n788 gnd 0.007621f
C1916 vdd.n789 gnd 0.007621f
C1917 vdd.n790 gnd 0.007621f
C1918 vdd.n792 gnd 0.007621f
C1919 vdd.n793 gnd 0.007621f
C1920 vdd.n795 gnd 0.007621f
C1921 vdd.n796 gnd 0.005548f
C1922 vdd.n798 gnd 0.007621f
C1923 vdd.t83 gnd 0.307978f
C1924 vdd.t82 gnd 0.315254f
C1925 vdd.t81 gnd 0.20106f
C1926 vdd.n799 gnd 0.108662f
C1927 vdd.n800 gnd 0.061637f
C1928 vdd.n801 gnd 0.010892f
C1929 vdd.n802 gnd 0.017813f
C1930 vdd.n804 gnd 0.007621f
C1931 vdd.n805 gnd 0.778867f
C1932 vdd.n806 gnd 0.016885f
C1933 vdd.n807 gnd 0.016885f
C1934 vdd.n808 gnd 0.007621f
C1935 vdd.n809 gnd 0.018084f
C1936 vdd.n810 gnd 0.007621f
C1937 vdd.n811 gnd 0.007621f
C1938 vdd.n812 gnd 0.007621f
C1939 vdd.n813 gnd 0.007621f
C1940 vdd.n814 gnd 0.007621f
C1941 vdd.n816 gnd 0.007621f
C1942 vdd.n817 gnd 0.007621f
C1943 vdd.n819 gnd 0.007621f
C1944 vdd.n820 gnd 0.007621f
C1945 vdd.n822 gnd 0.007621f
C1946 vdd.n823 gnd 0.007621f
C1947 vdd.n825 gnd 0.007621f
C1948 vdd.n826 gnd 0.007621f
C1949 vdd.n828 gnd 0.007621f
C1950 vdd.n829 gnd 0.007621f
C1951 vdd.n831 gnd 0.007621f
C1952 vdd.t76 gnd 0.307978f
C1953 vdd.t75 gnd 0.315254f
C1954 vdd.t73 gnd 0.20106f
C1955 vdd.n832 gnd 0.108662f
C1956 vdd.n833 gnd 0.061637f
C1957 vdd.n834 gnd 0.007621f
C1958 vdd.n836 gnd 0.007621f
C1959 vdd.n837 gnd 0.007621f
C1960 vdd.t74 gnd 0.389434f
C1961 vdd.n838 gnd 0.007621f
C1962 vdd.n839 gnd 0.007621f
C1963 vdd.n840 gnd 0.007621f
C1964 vdd.n841 gnd 0.007621f
C1965 vdd.n842 gnd 0.007621f
C1966 vdd.n843 gnd 0.778867f
C1967 vdd.n844 gnd 0.007621f
C1968 vdd.n845 gnd 0.007621f
C1969 vdd.n846 gnd 0.681509f
C1970 vdd.n847 gnd 0.007621f
C1971 vdd.n848 gnd 0.007621f
C1972 vdd.n849 gnd 0.006725f
C1973 vdd.n850 gnd 0.007621f
C1974 vdd.n851 gnd 0.687236f
C1975 vdd.n852 gnd 0.007621f
C1976 vdd.n853 gnd 0.007621f
C1977 vdd.n854 gnd 0.007621f
C1978 vdd.n855 gnd 0.007621f
C1979 vdd.n856 gnd 0.007621f
C1980 vdd.n857 gnd 0.778867f
C1981 vdd.n858 gnd 0.007621f
C1982 vdd.n859 gnd 0.007621f
C1983 vdd.t46 gnd 0.349345f
C1984 vdd.t113 gnd 0.091632f
C1985 vdd.n860 gnd 0.007621f
C1986 vdd.n861 gnd 0.007621f
C1987 vdd.n862 gnd 0.007621f
C1988 vdd.t9 gnd 0.389434f
C1989 vdd.n863 gnd 0.007621f
C1990 vdd.n864 gnd 0.007621f
C1991 vdd.n865 gnd 0.007621f
C1992 vdd.n866 gnd 0.007621f
C1993 vdd.n867 gnd 0.007621f
C1994 vdd.t4 gnd 0.389434f
C1995 vdd.n868 gnd 0.007621f
C1996 vdd.n869 gnd 0.007621f
C1997 vdd.n870 gnd 0.647147f
C1998 vdd.n871 gnd 0.007621f
C1999 vdd.n872 gnd 0.007621f
C2000 vdd.n873 gnd 0.007621f
C2001 vdd.n874 gnd 0.475338f
C2002 vdd.n875 gnd 0.007621f
C2003 vdd.n876 gnd 0.007621f
C2004 vdd.t119 gnd 0.389434f
C2005 vdd.n877 gnd 0.007621f
C2006 vdd.n878 gnd 0.007621f
C2007 vdd.n879 gnd 0.007621f
C2008 vdd.n880 gnd 0.647147f
C2009 vdd.n881 gnd 0.007621f
C2010 vdd.n882 gnd 0.007621f
C2011 vdd.t116 gnd 0.332164f
C2012 vdd.t294 gnd 0.303529f
C2013 vdd.n883 gnd 0.007621f
C2014 vdd.n884 gnd 0.007621f
C2015 vdd.n885 gnd 0.007621f
C2016 vdd.t14 gnd 0.389434f
C2017 vdd.n886 gnd 0.007621f
C2018 vdd.n887 gnd 0.007621f
C2019 vdd.t283 gnd 0.389434f
C2020 vdd.n888 gnd 0.007621f
C2021 vdd.n889 gnd 0.007621f
C2022 vdd.n890 gnd 0.007621f
C2023 vdd.t16 gnd 0.286348f
C2024 vdd.n891 gnd 0.007621f
C2025 vdd.n892 gnd 0.007621f
C2026 vdd.n893 gnd 0.664328f
C2027 vdd.n894 gnd 0.007621f
C2028 vdd.n895 gnd 0.007621f
C2029 vdd.n896 gnd 0.007621f
C2030 vdd.n897 gnd 0.778867f
C2031 vdd.n898 gnd 0.007621f
C2032 vdd.n899 gnd 0.007621f
C2033 vdd.t1 gnd 0.349345f
C2034 vdd.n900 gnd 0.492519f
C2035 vdd.n901 gnd 0.007621f
C2036 vdd.n902 gnd 0.007621f
C2037 vdd.n903 gnd 0.007621f
C2038 vdd.t114 gnd 0.389434f
C2039 vdd.n904 gnd 0.007621f
C2040 vdd.n905 gnd 0.007621f
C2041 vdd.n906 gnd 0.007621f
C2042 vdd.n907 gnd 0.007621f
C2043 vdd.n908 gnd 0.007621f
C2044 vdd.t288 gnd 0.778867f
C2045 vdd.n909 gnd 0.007621f
C2046 vdd.n910 gnd 0.007621f
C2047 vdd.t78 gnd 0.389434f
C2048 vdd.n911 gnd 0.007621f
C2049 vdd.n912 gnd 0.018084f
C2050 vdd.n913 gnd 0.018084f
C2051 vdd.t290 gnd 0.733052f
C2052 vdd.n914 gnd 0.016885f
C2053 vdd.n915 gnd 0.016885f
C2054 vdd.n916 gnd 0.018084f
C2055 vdd.n917 gnd 0.007621f
C2056 vdd.n918 gnd 0.007621f
C2057 vdd.t12 gnd 0.733052f
C2058 vdd.n936 gnd 0.018084f
C2059 vdd.n954 gnd 0.016885f
C2060 vdd.n955 gnd 0.007621f
C2061 vdd.n956 gnd 0.016885f
C2062 vdd.t97 gnd 0.307978f
C2063 vdd.t96 gnd 0.315254f
C2064 vdd.t95 gnd 0.20106f
C2065 vdd.n957 gnd 0.108662f
C2066 vdd.n958 gnd 0.061637f
C2067 vdd.n959 gnd 0.017813f
C2068 vdd.n960 gnd 0.007621f
C2069 vdd.t5 gnd 0.778867f
C2070 vdd.n961 gnd 0.016885f
C2071 vdd.n962 gnd 0.007621f
C2072 vdd.n963 gnd 0.018084f
C2073 vdd.n964 gnd 0.007621f
C2074 vdd.t72 gnd 0.307978f
C2075 vdd.t71 gnd 0.315254f
C2076 vdd.t69 gnd 0.20106f
C2077 vdd.n965 gnd 0.108662f
C2078 vdd.n966 gnd 0.061637f
C2079 vdd.n967 gnd 0.010892f
C2080 vdd.n968 gnd 0.007621f
C2081 vdd.n969 gnd 0.007621f
C2082 vdd.t70 gnd 0.389434f
C2083 vdd.n970 gnd 0.007621f
C2084 vdd.n971 gnd 0.007621f
C2085 vdd.n972 gnd 0.007621f
C2086 vdd.n973 gnd 0.007621f
C2087 vdd.n974 gnd 0.007621f
C2088 vdd.n975 gnd 0.007621f
C2089 vdd.n976 gnd 0.778867f
C2090 vdd.n977 gnd 0.007621f
C2091 vdd.n978 gnd 0.007621f
C2092 vdd.t117 gnd 0.389434f
C2093 vdd.n979 gnd 0.007621f
C2094 vdd.n980 gnd 0.007621f
C2095 vdd.n981 gnd 0.007621f
C2096 vdd.n982 gnd 0.007621f
C2097 vdd.n983 gnd 0.492519f
C2098 vdd.n984 gnd 0.007621f
C2099 vdd.n985 gnd 0.007621f
C2100 vdd.n986 gnd 0.007621f
C2101 vdd.n987 gnd 0.007621f
C2102 vdd.n988 gnd 0.007621f
C2103 vdd.n989 gnd 0.664328f
C2104 vdd.n990 gnd 0.007621f
C2105 vdd.n991 gnd 0.007621f
C2106 vdd.t284 gnd 0.349345f
C2107 vdd.t11 gnd 0.286348f
C2108 vdd.n992 gnd 0.007621f
C2109 vdd.n993 gnd 0.007621f
C2110 vdd.n994 gnd 0.007621f
C2111 vdd.t3 gnd 0.389434f
C2112 vdd.n995 gnd 0.007621f
C2113 vdd.n996 gnd 0.007621f
C2114 vdd.t292 gnd 0.389434f
C2115 vdd.n997 gnd 0.007621f
C2116 vdd.n998 gnd 0.007621f
C2117 vdd.n999 gnd 0.007621f
C2118 vdd.t7 gnd 0.303529f
C2119 vdd.n1000 gnd 0.007621f
C2120 vdd.n1001 gnd 0.007621f
C2121 vdd.n1002 gnd 0.647147f
C2122 vdd.n1003 gnd 0.007621f
C2123 vdd.n1004 gnd 0.007621f
C2124 vdd.n1005 gnd 0.007621f
C2125 vdd.t121 gnd 0.389434f
C2126 vdd.n1006 gnd 0.007621f
C2127 vdd.n1007 gnd 0.007621f
C2128 vdd.t33 gnd 0.332164f
C2129 vdd.n1008 gnd 0.475338f
C2130 vdd.n1009 gnd 0.007621f
C2131 vdd.n1010 gnd 0.007621f
C2132 vdd.n1011 gnd 0.007621f
C2133 vdd.n1012 gnd 0.647147f
C2134 vdd.n1013 gnd 0.007621f
C2135 vdd.n1014 gnd 0.007621f
C2136 vdd.t0 gnd 0.389434f
C2137 vdd.n1015 gnd 0.007621f
C2138 vdd.n1016 gnd 0.007621f
C2139 vdd.n1017 gnd 0.007621f
C2140 vdd.n1018 gnd 0.778867f
C2141 vdd.n1019 gnd 0.007621f
C2142 vdd.n1020 gnd 0.007621f
C2143 vdd.t110 gnd 0.389434f
C2144 vdd.n1021 gnd 0.007621f
C2145 vdd.n1022 gnd 0.007621f
C2146 vdd.n1023 gnd 0.007621f
C2147 vdd.t10 gnd 0.091632f
C2148 vdd.n1024 gnd 0.007621f
C2149 vdd.n1025 gnd 0.007621f
C2150 vdd.n1026 gnd 0.007621f
C2151 vdd.t90 gnd 0.315254f
C2152 vdd.t88 gnd 0.20106f
C2153 vdd.t91 gnd 0.315254f
C2154 vdd.n1027 gnd 0.177186f
C2155 vdd.n1028 gnd 0.007621f
C2156 vdd.n1029 gnd 0.007621f
C2157 vdd.n1030 gnd 0.778867f
C2158 vdd.n1031 gnd 0.007621f
C2159 vdd.n1032 gnd 0.007621f
C2160 vdd.t89 gnd 0.349345f
C2161 vdd.n1033 gnd 0.687236f
C2162 vdd.n1034 gnd 0.007621f
C2163 vdd.n1035 gnd 0.007621f
C2164 vdd.n1036 gnd 0.007621f
C2165 vdd.n1037 gnd 0.681509f
C2166 vdd.n1038 gnd 0.007621f
C2167 vdd.n1039 gnd 0.007621f
C2168 vdd.n1040 gnd 0.007621f
C2169 vdd.n1041 gnd 0.007621f
C2170 vdd.n1042 gnd 0.007621f
C2171 vdd.n1043 gnd 0.778867f
C2172 vdd.n1044 gnd 0.007621f
C2173 vdd.n1045 gnd 0.007621f
C2174 vdd.t85 gnd 0.389434f
C2175 vdd.n1046 gnd 0.007621f
C2176 vdd.n1047 gnd 0.018084f
C2177 vdd.n1048 gnd 0.018084f
C2178 vdd.n1049 gnd 7.891759f
C2179 vdd.n1050 gnd 0.016885f
C2180 vdd.n1051 gnd 0.016885f
C2181 vdd.n1052 gnd 0.018084f
C2182 vdd.n1053 gnd 0.007621f
C2183 vdd.n1054 gnd 0.007621f
C2184 vdd.n1055 gnd 0.007621f
C2185 vdd.n1056 gnd 0.007621f
C2186 vdd.n1057 gnd 0.007621f
C2187 vdd.n1058 gnd 0.007621f
C2188 vdd.n1059 gnd 0.007621f
C2189 vdd.n1060 gnd 0.007621f
C2190 vdd.n1062 gnd 0.007621f
C2191 vdd.n1063 gnd 0.007621f
C2192 vdd.n1064 gnd 0.007173f
C2193 vdd.n1067 gnd 0.027694f
C2194 vdd.n1068 gnd 0.009021f
C2195 vdd.n1069 gnd 0.011208f
C2196 vdd.n1071 gnd 0.011208f
C2197 vdd.n1072 gnd 0.007487f
C2198 vdd.t42 gnd 0.572697f
C2199 vdd.n1073 gnd 8.281191f
C2200 vdd.n1074 gnd 0.011208f
C2201 vdd.n1075 gnd 0.027694f
C2202 vdd.n1076 gnd 0.009021f
C2203 vdd.n1077 gnd 0.011208f
C2204 vdd.n1078 gnd 0.009021f
C2205 vdd.n1079 gnd 0.011208f
C2206 vdd.n1080 gnd 1.14539f
C2207 vdd.n1081 gnd 0.011208f
C2208 vdd.n1082 gnd 0.009021f
C2209 vdd.n1083 gnd 0.009021f
C2210 vdd.n1084 gnd 0.011208f
C2211 vdd.n1085 gnd 0.009021f
C2212 vdd.n1086 gnd 0.011208f
C2213 vdd.t123 gnd 0.572697f
C2214 vdd.n1087 gnd 0.011208f
C2215 vdd.n1088 gnd 0.009021f
C2216 vdd.n1089 gnd 0.011208f
C2217 vdd.n1090 gnd 0.009021f
C2218 vdd.n1091 gnd 0.011208f
C2219 vdd.t260 gnd 0.572697f
C2220 vdd.n1092 gnd 0.011208f
C2221 vdd.n1093 gnd 0.009021f
C2222 vdd.n1094 gnd 0.011208f
C2223 vdd.n1095 gnd 0.009021f
C2224 vdd.n1096 gnd 0.011208f
C2225 vdd.n1097 gnd 0.922042f
C2226 vdd.n1098 gnd 0.950677f
C2227 vdd.t141 gnd 0.572697f
C2228 vdd.n1099 gnd 0.011208f
C2229 vdd.n1100 gnd 0.009021f
C2230 vdd.n1101 gnd 0.011208f
C2231 vdd.n1102 gnd 0.009021f
C2232 vdd.n1103 gnd 0.011208f
C2233 vdd.n1104 gnd 0.727325f
C2234 vdd.n1105 gnd 0.011208f
C2235 vdd.n1106 gnd 0.009021f
C2236 vdd.n1107 gnd 0.011208f
C2237 vdd.n1108 gnd 0.009021f
C2238 vdd.n1109 gnd 0.011208f
C2239 vdd.t131 gnd 0.572697f
C2240 vdd.t171 gnd 0.572697f
C2241 vdd.n1110 gnd 0.011208f
C2242 vdd.n1111 gnd 0.009021f
C2243 vdd.n1112 gnd 0.011208f
C2244 vdd.n1113 gnd 0.009021f
C2245 vdd.n1114 gnd 0.011208f
C2246 vdd.t196 gnd 0.572697f
C2247 vdd.n1115 gnd 0.011208f
C2248 vdd.n1116 gnd 0.009021f
C2249 vdd.n1117 gnd 0.011208f
C2250 vdd.n1118 gnd 0.009021f
C2251 vdd.n1119 gnd 0.011208f
C2252 vdd.t235 gnd 0.572697f
C2253 vdd.n1120 gnd 0.807502f
C2254 vdd.n1121 gnd 0.011208f
C2255 vdd.n1122 gnd 0.009021f
C2256 vdd.n1123 gnd 0.011208f
C2257 vdd.n1124 gnd 0.009021f
C2258 vdd.n1125 gnd 0.011208f
C2259 vdd.n1126 gnd 0.899134f
C2260 vdd.n1127 gnd 0.011208f
C2261 vdd.n1128 gnd 0.009021f
C2262 vdd.n1129 gnd 0.011208f
C2263 vdd.n1130 gnd 0.009021f
C2264 vdd.n1131 gnd 0.011208f
C2265 vdd.n1132 gnd 0.704417f
C2266 vdd.t135 gnd 0.572697f
C2267 vdd.n1133 gnd 0.011208f
C2268 vdd.n1134 gnd 0.009021f
C2269 vdd.n1135 gnd 0.011208f
C2270 vdd.n1136 gnd 0.009021f
C2271 vdd.n1137 gnd 0.011208f
C2272 vdd.t149 gnd 0.572697f
C2273 vdd.n1138 gnd 0.011208f
C2274 vdd.n1139 gnd 0.009021f
C2275 vdd.n1140 gnd 0.011208f
C2276 vdd.n1141 gnd 0.009021f
C2277 vdd.n1142 gnd 0.011208f
C2278 vdd.t168 gnd 0.572697f
C2279 vdd.n1143 gnd 0.635693f
C2280 vdd.n1144 gnd 0.011208f
C2281 vdd.n1145 gnd 0.009021f
C2282 vdd.n1146 gnd 0.011208f
C2283 vdd.n1147 gnd 0.009021f
C2284 vdd.n1148 gnd 0.011208f
C2285 vdd.t215 gnd 0.572697f
C2286 vdd.n1149 gnd 0.011208f
C2287 vdd.n1150 gnd 0.009021f
C2288 vdd.n1151 gnd 0.011208f
C2289 vdd.n1152 gnd 0.009021f
C2290 vdd.n1153 gnd 0.011208f
C2291 vdd.n1154 gnd 0.876226f
C2292 vdd.n1155 gnd 0.950677f
C2293 vdd.t217 gnd 0.572697f
C2294 vdd.n1156 gnd 0.011208f
C2295 vdd.n1157 gnd 0.009021f
C2296 vdd.n1158 gnd 0.011208f
C2297 vdd.n1159 gnd 0.009021f
C2298 vdd.n1160 gnd 0.011208f
C2299 vdd.n1161 gnd 0.681509f
C2300 vdd.n1162 gnd 0.011208f
C2301 vdd.n1163 gnd 0.009021f
C2302 vdd.n1164 gnd 0.011208f
C2303 vdd.n1165 gnd 0.009021f
C2304 vdd.n1166 gnd 0.011208f
C2305 vdd.t162 gnd 0.572697f
C2306 vdd.t165 gnd 0.572697f
C2307 vdd.n1167 gnd 0.011208f
C2308 vdd.n1168 gnd 0.009021f
C2309 vdd.n1169 gnd 0.011208f
C2310 vdd.n1170 gnd 0.009021f
C2311 vdd.n1171 gnd 0.011208f
C2312 vdd.t127 gnd 0.572697f
C2313 vdd.n1172 gnd 0.011208f
C2314 vdd.n1173 gnd 0.009021f
C2315 vdd.n1174 gnd 0.011208f
C2316 vdd.n1175 gnd 0.009021f
C2317 vdd.n1176 gnd 0.011208f
C2318 vdd.t129 gnd 0.572697f
C2319 vdd.n1177 gnd 0.853318f
C2320 vdd.n1178 gnd 0.011208f
C2321 vdd.n1179 gnd 0.009021f
C2322 vdd.n1180 gnd 0.011208f
C2323 vdd.n1181 gnd 0.009021f
C2324 vdd.n1182 gnd 0.011208f
C2325 vdd.n1183 gnd 1.14539f
C2326 vdd.n1184 gnd 0.011208f
C2327 vdd.n1185 gnd 0.009021f
C2328 vdd.n1186 gnd 0.027113f
C2329 vdd.n1187 gnd 0.007487f
C2330 vdd.n1188 gnd 0.027113f
C2331 vdd.t50 gnd 0.572697f
C2332 vdd.n1189 gnd 0.027113f
C2333 vdd.n1190 gnd 0.007487f
C2334 vdd.n1191 gnd 0.011208f
C2335 vdd.n1192 gnd 0.009021f
C2336 vdd.n1193 gnd 0.011208f
C2337 vdd.n1224 gnd 0.027694f
C2338 vdd.n1225 gnd 1.68946f
C2339 vdd.n1226 gnd 0.011208f
C2340 vdd.n1227 gnd 0.009021f
C2341 vdd.n1228 gnd 0.011208f
C2342 vdd.n1229 gnd 0.011208f
C2343 vdd.n1230 gnd 0.011208f
C2344 vdd.n1231 gnd 0.011208f
C2345 vdd.n1232 gnd 0.011208f
C2346 vdd.n1233 gnd 0.009021f
C2347 vdd.n1234 gnd 0.011208f
C2348 vdd.n1235 gnd 0.011208f
C2349 vdd.n1236 gnd 0.011208f
C2350 vdd.n1237 gnd 0.011208f
C2351 vdd.n1238 gnd 0.011208f
C2352 vdd.n1239 gnd 0.009021f
C2353 vdd.n1240 gnd 0.011208f
C2354 vdd.n1241 gnd 0.011208f
C2355 vdd.n1242 gnd 0.011208f
C2356 vdd.n1243 gnd 0.011208f
C2357 vdd.n1244 gnd 0.011208f
C2358 vdd.n1245 gnd 0.009021f
C2359 vdd.n1246 gnd 0.011208f
C2360 vdd.n1247 gnd 0.011208f
C2361 vdd.n1248 gnd 0.011208f
C2362 vdd.n1249 gnd 0.011208f
C2363 vdd.n1250 gnd 0.011208f
C2364 vdd.t64 gnd 0.137886f
C2365 vdd.t65 gnd 0.147363f
C2366 vdd.t63 gnd 0.180078f
C2367 vdd.n1251 gnd 0.230835f
C2368 vdd.n1252 gnd 0.194845f
C2369 vdd.n1253 gnd 0.019305f
C2370 vdd.n1254 gnd 0.011208f
C2371 vdd.n1255 gnd 0.011208f
C2372 vdd.n1256 gnd 0.011208f
C2373 vdd.n1257 gnd 0.011208f
C2374 vdd.n1258 gnd 0.011208f
C2375 vdd.n1259 gnd 0.009021f
C2376 vdd.n1260 gnd 0.011208f
C2377 vdd.n1261 gnd 0.011208f
C2378 vdd.n1262 gnd 0.011208f
C2379 vdd.n1263 gnd 0.011208f
C2380 vdd.n1264 gnd 0.011208f
C2381 vdd.n1265 gnd 0.009021f
C2382 vdd.n1266 gnd 0.011208f
C2383 vdd.n1267 gnd 0.011208f
C2384 vdd.n1268 gnd 0.011208f
C2385 vdd.n1269 gnd 0.011208f
C2386 vdd.n1270 gnd 0.011208f
C2387 vdd.n1271 gnd 0.009021f
C2388 vdd.n1272 gnd 0.011208f
C2389 vdd.n1273 gnd 0.011208f
C2390 vdd.n1274 gnd 0.011208f
C2391 vdd.n1275 gnd 0.011208f
C2392 vdd.n1276 gnd 0.011208f
C2393 vdd.n1277 gnd 0.009021f
C2394 vdd.n1278 gnd 0.011208f
C2395 vdd.n1279 gnd 0.011208f
C2396 vdd.n1280 gnd 0.011208f
C2397 vdd.n1281 gnd 0.011208f
C2398 vdd.n1282 gnd 0.011208f
C2399 vdd.n1283 gnd 0.009021f
C2400 vdd.n1284 gnd 0.011208f
C2401 vdd.n1285 gnd 0.011208f
C2402 vdd.n1286 gnd 0.011208f
C2403 vdd.n1287 gnd 0.011208f
C2404 vdd.n1288 gnd 0.009021f
C2405 vdd.n1289 gnd 0.011208f
C2406 vdd.n1290 gnd 0.011208f
C2407 vdd.n1291 gnd 0.011208f
C2408 vdd.n1292 gnd 0.011208f
C2409 vdd.n1293 gnd 0.011208f
C2410 vdd.n1294 gnd 0.009021f
C2411 vdd.n1295 gnd 0.011208f
C2412 vdd.n1296 gnd 0.011208f
C2413 vdd.n1297 gnd 0.011208f
C2414 vdd.n1298 gnd 0.011208f
C2415 vdd.n1299 gnd 0.011208f
C2416 vdd.n1300 gnd 0.009021f
C2417 vdd.n1301 gnd 0.011208f
C2418 vdd.n1302 gnd 0.011208f
C2419 vdd.n1303 gnd 0.011208f
C2420 vdd.n1304 gnd 0.011208f
C2421 vdd.n1305 gnd 0.011208f
C2422 vdd.n1306 gnd 0.009021f
C2423 vdd.n1307 gnd 0.011208f
C2424 vdd.n1308 gnd 0.011208f
C2425 vdd.n1309 gnd 0.011208f
C2426 vdd.n1310 gnd 0.011208f
C2427 vdd.n1311 gnd 0.011208f
C2428 vdd.n1312 gnd 0.009021f
C2429 vdd.n1313 gnd 0.011208f
C2430 vdd.n1314 gnd 0.011208f
C2431 vdd.n1315 gnd 0.011208f
C2432 vdd.n1316 gnd 0.011208f
C2433 vdd.t61 gnd 0.137886f
C2434 vdd.t62 gnd 0.147363f
C2435 vdd.t60 gnd 0.180078f
C2436 vdd.n1317 gnd 0.230835f
C2437 vdd.n1318 gnd 0.194845f
C2438 vdd.n1319 gnd 0.014794f
C2439 vdd.n1320 gnd 0.004285f
C2440 vdd.n1321 gnd 0.027694f
C2441 vdd.n1322 gnd 0.011208f
C2442 vdd.n1323 gnd 0.004736f
C2443 vdd.n1324 gnd 0.009021f
C2444 vdd.n1325 gnd 0.009021f
C2445 vdd.n1326 gnd 0.011208f
C2446 vdd.n1327 gnd 0.011208f
C2447 vdd.n1328 gnd 0.011208f
C2448 vdd.n1329 gnd 0.009021f
C2449 vdd.n1330 gnd 0.009021f
C2450 vdd.n1331 gnd 0.009021f
C2451 vdd.n1332 gnd 0.011208f
C2452 vdd.n1333 gnd 0.011208f
C2453 vdd.n1334 gnd 0.011208f
C2454 vdd.n1335 gnd 0.009021f
C2455 vdd.n1336 gnd 0.009021f
C2456 vdd.n1337 gnd 0.009021f
C2457 vdd.n1338 gnd 0.011208f
C2458 vdd.n1339 gnd 0.011208f
C2459 vdd.n1340 gnd 0.011208f
C2460 vdd.n1341 gnd 0.009021f
C2461 vdd.n1342 gnd 0.009021f
C2462 vdd.n1343 gnd 0.009021f
C2463 vdd.n1344 gnd 0.011208f
C2464 vdd.n1345 gnd 0.011208f
C2465 vdd.n1346 gnd 0.011208f
C2466 vdd.n1347 gnd 0.009021f
C2467 vdd.n1348 gnd 0.009021f
C2468 vdd.n1349 gnd 0.009021f
C2469 vdd.n1350 gnd 0.011208f
C2470 vdd.n1351 gnd 0.011208f
C2471 vdd.n1352 gnd 0.011208f
C2472 vdd.n1353 gnd 0.008931f
C2473 vdd.n1354 gnd 0.011208f
C2474 vdd.t51 gnd 0.137886f
C2475 vdd.t52 gnd 0.147363f
C2476 vdd.t49 gnd 0.180078f
C2477 vdd.n1355 gnd 0.230835f
C2478 vdd.n1356 gnd 0.194845f
C2479 vdd.n1357 gnd 0.019305f
C2480 vdd.n1358 gnd 0.006134f
C2481 vdd.n1359 gnd 0.011208f
C2482 vdd.n1360 gnd 0.011208f
C2483 vdd.n1361 gnd 0.011208f
C2484 vdd.n1362 gnd 0.009021f
C2485 vdd.n1363 gnd 0.009021f
C2486 vdd.n1364 gnd 0.009021f
C2487 vdd.n1365 gnd 0.011208f
C2488 vdd.n1366 gnd 0.011208f
C2489 vdd.n1367 gnd 0.011208f
C2490 vdd.n1368 gnd 0.009021f
C2491 vdd.n1369 gnd 0.009021f
C2492 vdd.n1370 gnd 0.009021f
C2493 vdd.n1371 gnd 0.011208f
C2494 vdd.n1372 gnd 0.011208f
C2495 vdd.n1373 gnd 0.011208f
C2496 vdd.n1374 gnd 0.009021f
C2497 vdd.n1375 gnd 0.009021f
C2498 vdd.n1376 gnd 0.009021f
C2499 vdd.n1377 gnd 0.011208f
C2500 vdd.n1378 gnd 0.011208f
C2501 vdd.n1379 gnd 0.011208f
C2502 vdd.n1380 gnd 0.009021f
C2503 vdd.n1381 gnd 0.009021f
C2504 vdd.n1382 gnd 0.009021f
C2505 vdd.n1383 gnd 0.011208f
C2506 vdd.n1384 gnd 0.011208f
C2507 vdd.n1385 gnd 0.011208f
C2508 vdd.n1386 gnd 0.009021f
C2509 vdd.n1387 gnd 0.009021f
C2510 vdd.n1388 gnd 0.007533f
C2511 vdd.n1389 gnd 0.011208f
C2512 vdd.n1390 gnd 0.011208f
C2513 vdd.n1391 gnd 0.011208f
C2514 vdd.n1392 gnd 0.007533f
C2515 vdd.n1393 gnd 0.009021f
C2516 vdd.n1394 gnd 0.009021f
C2517 vdd.n1395 gnd 0.011208f
C2518 vdd.n1396 gnd 0.011208f
C2519 vdd.n1397 gnd 0.011208f
C2520 vdd.n1398 gnd 0.009021f
C2521 vdd.n1399 gnd 0.009021f
C2522 vdd.n1400 gnd 0.009021f
C2523 vdd.n1401 gnd 0.011208f
C2524 vdd.n1402 gnd 0.011208f
C2525 vdd.n1403 gnd 0.011208f
C2526 vdd.n1404 gnd 0.009021f
C2527 vdd.n1405 gnd 0.009021f
C2528 vdd.n1406 gnd 0.009021f
C2529 vdd.n1407 gnd 0.011208f
C2530 vdd.n1408 gnd 0.011208f
C2531 vdd.n1409 gnd 0.011208f
C2532 vdd.n1410 gnd 0.009021f
C2533 vdd.n1411 gnd 0.009021f
C2534 vdd.n1412 gnd 0.009021f
C2535 vdd.n1413 gnd 0.011208f
C2536 vdd.n1414 gnd 0.011208f
C2537 vdd.n1415 gnd 0.011208f
C2538 vdd.n1416 gnd 0.009021f
C2539 vdd.n1417 gnd 0.011208f
C2540 vdd.n1418 gnd 2.71458f
C2541 vdd.n1420 gnd 0.027694f
C2542 vdd.n1421 gnd 0.007487f
C2543 vdd.n1422 gnd 0.027694f
C2544 vdd.n1423 gnd 0.027113f
C2545 vdd.n1424 gnd 0.011208f
C2546 vdd.n1425 gnd 0.009021f
C2547 vdd.n1426 gnd 0.011208f
C2548 vdd.n1427 gnd 0.578424f
C2549 vdd.n1428 gnd 0.011208f
C2550 vdd.n1429 gnd 0.009021f
C2551 vdd.n1430 gnd 0.011208f
C2552 vdd.n1431 gnd 0.011208f
C2553 vdd.n1432 gnd 0.011208f
C2554 vdd.n1433 gnd 0.009021f
C2555 vdd.n1434 gnd 0.011208f
C2556 vdd.n1435 gnd 1.04803f
C2557 vdd.n1436 gnd 1.14539f
C2558 vdd.n1437 gnd 0.011208f
C2559 vdd.n1438 gnd 0.009021f
C2560 vdd.n1439 gnd 0.011208f
C2561 vdd.n1440 gnd 0.011208f
C2562 vdd.n1441 gnd 0.011208f
C2563 vdd.n1442 gnd 0.009021f
C2564 vdd.n1443 gnd 0.011208f
C2565 vdd.n1444 gnd 0.670055f
C2566 vdd.n1445 gnd 0.011208f
C2567 vdd.n1446 gnd 0.009021f
C2568 vdd.n1447 gnd 0.011208f
C2569 vdd.n1448 gnd 0.011208f
C2570 vdd.n1449 gnd 0.011208f
C2571 vdd.n1450 gnd 0.009021f
C2572 vdd.n1451 gnd 0.011208f
C2573 vdd.n1452 gnd 0.658601f
C2574 vdd.n1453 gnd 0.864772f
C2575 vdd.n1454 gnd 0.011208f
C2576 vdd.n1455 gnd 0.009021f
C2577 vdd.n1456 gnd 0.011208f
C2578 vdd.n1457 gnd 0.011208f
C2579 vdd.n1458 gnd 0.011208f
C2580 vdd.n1459 gnd 0.009021f
C2581 vdd.n1460 gnd 0.011208f
C2582 vdd.n1461 gnd 0.950677f
C2583 vdd.n1462 gnd 0.011208f
C2584 vdd.n1463 gnd 0.009021f
C2585 vdd.n1464 gnd 0.011208f
C2586 vdd.n1465 gnd 0.011208f
C2587 vdd.n1466 gnd 0.011208f
C2588 vdd.n1467 gnd 0.009021f
C2589 vdd.n1468 gnd 0.011208f
C2590 vdd.t139 gnd 0.572697f
C2591 vdd.n1469 gnd 0.841864f
C2592 vdd.n1470 gnd 0.011208f
C2593 vdd.n1471 gnd 0.009021f
C2594 vdd.n1472 gnd 0.011208f
C2595 vdd.n1473 gnd 0.011208f
C2596 vdd.n1474 gnd 0.011208f
C2597 vdd.n1475 gnd 0.009021f
C2598 vdd.n1476 gnd 0.011208f
C2599 vdd.n1477 gnd 0.647147f
C2600 vdd.n1478 gnd 0.011208f
C2601 vdd.n1479 gnd 0.009021f
C2602 vdd.n1480 gnd 0.011208f
C2603 vdd.n1481 gnd 0.011208f
C2604 vdd.n1482 gnd 0.011208f
C2605 vdd.n1483 gnd 0.009021f
C2606 vdd.n1484 gnd 0.011208f
C2607 vdd.n1485 gnd 0.83041f
C2608 vdd.n1486 gnd 0.692963f
C2609 vdd.n1487 gnd 0.011208f
C2610 vdd.n1488 gnd 0.009021f
C2611 vdd.n1489 gnd 0.011208f
C2612 vdd.n1490 gnd 0.011208f
C2613 vdd.n1491 gnd 0.011208f
C2614 vdd.n1492 gnd 0.009021f
C2615 vdd.n1493 gnd 0.011208f
C2616 vdd.n1494 gnd 0.88768f
C2617 vdd.n1495 gnd 0.011208f
C2618 vdd.n1496 gnd 0.009021f
C2619 vdd.n1497 gnd 0.011208f
C2620 vdd.n1498 gnd 0.011208f
C2621 vdd.n1499 gnd 0.011208f
C2622 vdd.n1500 gnd 0.009021f
C2623 vdd.n1501 gnd 0.011208f
C2624 vdd.t185 gnd 0.572697f
C2625 vdd.n1502 gnd 0.950677f
C2626 vdd.n1503 gnd 0.011208f
C2627 vdd.n1504 gnd 0.009021f
C2628 vdd.n1505 gnd 0.011208f
C2629 vdd.n1506 gnd 0.008614f
C2630 vdd.n1507 gnd 0.006151f
C2631 vdd.n1508 gnd 0.005708f
C2632 vdd.n1509 gnd 0.003157f
C2633 vdd.n1510 gnd 0.00725f
C2634 vdd.n1511 gnd 0.003067f
C2635 vdd.n1512 gnd 0.003248f
C2636 vdd.n1513 gnd 0.005708f
C2637 vdd.n1514 gnd 0.003067f
C2638 vdd.n1515 gnd 0.00725f
C2639 vdd.n1516 gnd 0.003248f
C2640 vdd.n1517 gnd 0.005708f
C2641 vdd.n1518 gnd 0.003067f
C2642 vdd.n1519 gnd 0.005437f
C2643 vdd.n1520 gnd 0.005453f
C2644 vdd.t124 gnd 0.015575f
C2645 vdd.n1521 gnd 0.034655f
C2646 vdd.n1522 gnd 0.18035f
C2647 vdd.n1523 gnd 0.003067f
C2648 vdd.n1524 gnd 0.003248f
C2649 vdd.n1525 gnd 0.00725f
C2650 vdd.n1526 gnd 0.00725f
C2651 vdd.n1527 gnd 0.003248f
C2652 vdd.n1528 gnd 0.003067f
C2653 vdd.n1529 gnd 0.005708f
C2654 vdd.n1530 gnd 0.005708f
C2655 vdd.n1531 gnd 0.003067f
C2656 vdd.n1532 gnd 0.003248f
C2657 vdd.n1533 gnd 0.00725f
C2658 vdd.n1534 gnd 0.00725f
C2659 vdd.n1535 gnd 0.003248f
C2660 vdd.n1536 gnd 0.003067f
C2661 vdd.n1537 gnd 0.005708f
C2662 vdd.n1538 gnd 0.005708f
C2663 vdd.n1539 gnd 0.003067f
C2664 vdd.n1540 gnd 0.003248f
C2665 vdd.n1541 gnd 0.00725f
C2666 vdd.n1542 gnd 0.00725f
C2667 vdd.n1543 gnd 0.01714f
C2668 vdd.n1544 gnd 0.003157f
C2669 vdd.n1545 gnd 0.003067f
C2670 vdd.n1546 gnd 0.014753f
C2671 vdd.n1547 gnd 0.0103f
C2672 vdd.t205 gnd 0.036084f
C2673 vdd.t267 gnd 0.036084f
C2674 vdd.n1548 gnd 0.247994f
C2675 vdd.n1549 gnd 0.195009f
C2676 vdd.t172 gnd 0.036084f
C2677 vdd.t246 gnd 0.036084f
C2678 vdd.n1550 gnd 0.247994f
C2679 vdd.n1551 gnd 0.157371f
C2680 vdd.t197 gnd 0.036084f
C2681 vdd.t255 gnd 0.036084f
C2682 vdd.n1552 gnd 0.247994f
C2683 vdd.n1553 gnd 0.157371f
C2684 vdd.t222 gnd 0.036084f
C2685 vdd.t273 gnd 0.036084f
C2686 vdd.n1554 gnd 0.247994f
C2687 vdd.n1555 gnd 0.157371f
C2688 vdd.t186 gnd 0.036084f
C2689 vdd.t136 gnd 0.036084f
C2690 vdd.n1556 gnd 0.247994f
C2691 vdd.n1557 gnd 0.157371f
C2692 vdd.t210 gnd 0.036084f
C2693 vdd.t150 gnd 0.036084f
C2694 vdd.n1558 gnd 0.247994f
C2695 vdd.n1559 gnd 0.157371f
C2696 vdd.t263 gnd 0.036084f
C2697 vdd.t279 gnd 0.036084f
C2698 vdd.n1560 gnd 0.247994f
C2699 vdd.n1561 gnd 0.157371f
C2700 vdd.t234 gnd 0.036084f
C2701 vdd.t155 gnd 0.036084f
C2702 vdd.n1562 gnd 0.247994f
C2703 vdd.n1563 gnd 0.157371f
C2704 vdd.t220 gnd 0.036084f
C2705 vdd.t163 gnd 0.036084f
C2706 vdd.n1564 gnd 0.247994f
C2707 vdd.n1565 gnd 0.157371f
C2708 vdd.n1566 gnd 0.006151f
C2709 vdd.n1567 gnd 0.005708f
C2710 vdd.n1568 gnd 0.003157f
C2711 vdd.n1569 gnd 0.00725f
C2712 vdd.n1570 gnd 0.003067f
C2713 vdd.n1571 gnd 0.003248f
C2714 vdd.n1572 gnd 0.005708f
C2715 vdd.n1573 gnd 0.003067f
C2716 vdd.n1574 gnd 0.00725f
C2717 vdd.n1575 gnd 0.003248f
C2718 vdd.n1576 gnd 0.005708f
C2719 vdd.n1577 gnd 0.003067f
C2720 vdd.n1578 gnd 0.005437f
C2721 vdd.n1579 gnd 0.005453f
C2722 vdd.t192 gnd 0.015575f
C2723 vdd.n1580 gnd 0.034655f
C2724 vdd.n1581 gnd 0.18035f
C2725 vdd.n1582 gnd 0.003067f
C2726 vdd.n1583 gnd 0.003248f
C2727 vdd.n1584 gnd 0.00725f
C2728 vdd.n1585 gnd 0.00725f
C2729 vdd.n1586 gnd 0.003248f
C2730 vdd.n1587 gnd 0.003067f
C2731 vdd.n1588 gnd 0.005708f
C2732 vdd.n1589 gnd 0.005708f
C2733 vdd.n1590 gnd 0.003067f
C2734 vdd.n1591 gnd 0.003248f
C2735 vdd.n1592 gnd 0.00725f
C2736 vdd.n1593 gnd 0.00725f
C2737 vdd.n1594 gnd 0.003248f
C2738 vdd.n1595 gnd 0.003067f
C2739 vdd.n1596 gnd 0.005708f
C2740 vdd.n1597 gnd 0.005708f
C2741 vdd.n1598 gnd 0.003067f
C2742 vdd.n1599 gnd 0.003248f
C2743 vdd.n1600 gnd 0.00725f
C2744 vdd.n1601 gnd 0.00725f
C2745 vdd.n1602 gnd 0.01714f
C2746 vdd.n1603 gnd 0.003157f
C2747 vdd.n1604 gnd 0.003067f
C2748 vdd.n1605 gnd 0.014753f
C2749 vdd.n1606 gnd 0.009977f
C2750 vdd.n1607 gnd 0.117085f
C2751 vdd.n1608 gnd 0.006151f
C2752 vdd.n1609 gnd 0.005708f
C2753 vdd.n1610 gnd 0.003157f
C2754 vdd.n1611 gnd 0.00725f
C2755 vdd.n1612 gnd 0.003067f
C2756 vdd.n1613 gnd 0.003248f
C2757 vdd.n1614 gnd 0.005708f
C2758 vdd.n1615 gnd 0.003067f
C2759 vdd.n1616 gnd 0.00725f
C2760 vdd.n1617 gnd 0.003248f
C2761 vdd.n1618 gnd 0.005708f
C2762 vdd.n1619 gnd 0.003067f
C2763 vdd.n1620 gnd 0.005437f
C2764 vdd.n1621 gnd 0.005453f
C2765 vdd.t256 gnd 0.015575f
C2766 vdd.n1622 gnd 0.034655f
C2767 vdd.n1623 gnd 0.18035f
C2768 vdd.n1624 gnd 0.003067f
C2769 vdd.n1625 gnd 0.003248f
C2770 vdd.n1626 gnd 0.00725f
C2771 vdd.n1627 gnd 0.00725f
C2772 vdd.n1628 gnd 0.003248f
C2773 vdd.n1629 gnd 0.003067f
C2774 vdd.n1630 gnd 0.005708f
C2775 vdd.n1631 gnd 0.005708f
C2776 vdd.n1632 gnd 0.003067f
C2777 vdd.n1633 gnd 0.003248f
C2778 vdd.n1634 gnd 0.00725f
C2779 vdd.n1635 gnd 0.00725f
C2780 vdd.n1636 gnd 0.003248f
C2781 vdd.n1637 gnd 0.003067f
C2782 vdd.n1638 gnd 0.005708f
C2783 vdd.n1639 gnd 0.005708f
C2784 vdd.n1640 gnd 0.003067f
C2785 vdd.n1641 gnd 0.003248f
C2786 vdd.n1642 gnd 0.00725f
C2787 vdd.n1643 gnd 0.00725f
C2788 vdd.n1644 gnd 0.01714f
C2789 vdd.n1645 gnd 0.003157f
C2790 vdd.n1646 gnd 0.003067f
C2791 vdd.n1647 gnd 0.014753f
C2792 vdd.n1648 gnd 0.0103f
C2793 vdd.t142 gnd 0.036084f
C2794 vdd.t261 gnd 0.036084f
C2795 vdd.n1649 gnd 0.247994f
C2796 vdd.n1650 gnd 0.195009f
C2797 vdd.t253 gnd 0.036084f
C2798 vdd.t238 gnd 0.036084f
C2799 vdd.n1651 gnd 0.247994f
C2800 vdd.n1652 gnd 0.157371f
C2801 vdd.t200 gnd 0.036084f
C2802 vdd.t132 gnd 0.036084f
C2803 vdd.n1653 gnd 0.247994f
C2804 vdd.n1654 gnd 0.157371f
C2805 vdd.t269 gnd 0.036084f
C2806 vdd.t236 gnd 0.036084f
C2807 vdd.n1655 gnd 0.247994f
C2808 vdd.n1656 gnd 0.157371f
C2809 vdd.t230 gnd 0.036084f
C2810 vdd.t175 gnd 0.036084f
C2811 vdd.n1657 gnd 0.247994f
C2812 vdd.n1658 gnd 0.157371f
C2813 vdd.t169 gnd 0.036084f
C2814 vdd.t233 gnd 0.036084f
C2815 vdd.n1659 gnd 0.247994f
C2816 vdd.n1660 gnd 0.157371f
C2817 vdd.t218 gnd 0.036084f
C2818 vdd.t216 gnd 0.036084f
C2819 vdd.n1661 gnd 0.247994f
C2820 vdd.n1662 gnd 0.157371f
C2821 vdd.t166 gnd 0.036084f
C2822 vdd.t140 gnd 0.036084f
C2823 vdd.n1663 gnd 0.247994f
C2824 vdd.n1664 gnd 0.157371f
C2825 vdd.t128 gnd 0.036084f
C2826 vdd.t211 gnd 0.036084f
C2827 vdd.n1665 gnd 0.247994f
C2828 vdd.n1666 gnd 0.157371f
C2829 vdd.n1667 gnd 0.006151f
C2830 vdd.n1668 gnd 0.005708f
C2831 vdd.n1669 gnd 0.003157f
C2832 vdd.n1670 gnd 0.00725f
C2833 vdd.n1671 gnd 0.003067f
C2834 vdd.n1672 gnd 0.003248f
C2835 vdd.n1673 gnd 0.005708f
C2836 vdd.n1674 gnd 0.003067f
C2837 vdd.n1675 gnd 0.00725f
C2838 vdd.n1676 gnd 0.003248f
C2839 vdd.n1677 gnd 0.005708f
C2840 vdd.n1678 gnd 0.003067f
C2841 vdd.n1679 gnd 0.005437f
C2842 vdd.n1680 gnd 0.005453f
C2843 vdd.t130 gnd 0.015575f
C2844 vdd.n1681 gnd 0.034655f
C2845 vdd.n1682 gnd 0.18035f
C2846 vdd.n1683 gnd 0.003067f
C2847 vdd.n1684 gnd 0.003248f
C2848 vdd.n1685 gnd 0.00725f
C2849 vdd.n1686 gnd 0.00725f
C2850 vdd.n1687 gnd 0.003248f
C2851 vdd.n1688 gnd 0.003067f
C2852 vdd.n1689 gnd 0.005708f
C2853 vdd.n1690 gnd 0.005708f
C2854 vdd.n1691 gnd 0.003067f
C2855 vdd.n1692 gnd 0.003248f
C2856 vdd.n1693 gnd 0.00725f
C2857 vdd.n1694 gnd 0.00725f
C2858 vdd.n1695 gnd 0.003248f
C2859 vdd.n1696 gnd 0.003067f
C2860 vdd.n1697 gnd 0.005708f
C2861 vdd.n1698 gnd 0.005708f
C2862 vdd.n1699 gnd 0.003067f
C2863 vdd.n1700 gnd 0.003248f
C2864 vdd.n1701 gnd 0.00725f
C2865 vdd.n1702 gnd 0.00725f
C2866 vdd.n1703 gnd 0.01714f
C2867 vdd.n1704 gnd 0.003157f
C2868 vdd.n1705 gnd 0.003067f
C2869 vdd.n1706 gnd 0.014753f
C2870 vdd.n1707 gnd 0.009977f
C2871 vdd.n1708 gnd 0.069654f
C2872 vdd.n1709 gnd 0.250981f
C2873 vdd.n1710 gnd 0.006151f
C2874 vdd.n1711 gnd 0.005708f
C2875 vdd.n1712 gnd 0.003157f
C2876 vdd.n1713 gnd 0.00725f
C2877 vdd.n1714 gnd 0.003067f
C2878 vdd.n1715 gnd 0.003248f
C2879 vdd.n1716 gnd 0.005708f
C2880 vdd.n1717 gnd 0.003067f
C2881 vdd.n1718 gnd 0.00725f
C2882 vdd.n1719 gnd 0.003248f
C2883 vdd.n1720 gnd 0.005708f
C2884 vdd.n1721 gnd 0.003067f
C2885 vdd.n1722 gnd 0.005437f
C2886 vdd.n1723 gnd 0.005453f
C2887 vdd.t272 gnd 0.015575f
C2888 vdd.n1724 gnd 0.034655f
C2889 vdd.n1725 gnd 0.18035f
C2890 vdd.n1726 gnd 0.003067f
C2891 vdd.n1727 gnd 0.003248f
C2892 vdd.n1728 gnd 0.00725f
C2893 vdd.n1729 gnd 0.00725f
C2894 vdd.n1730 gnd 0.003248f
C2895 vdd.n1731 gnd 0.003067f
C2896 vdd.n1732 gnd 0.005708f
C2897 vdd.n1733 gnd 0.005708f
C2898 vdd.n1734 gnd 0.003067f
C2899 vdd.n1735 gnd 0.003248f
C2900 vdd.n1736 gnd 0.00725f
C2901 vdd.n1737 gnd 0.00725f
C2902 vdd.n1738 gnd 0.003248f
C2903 vdd.n1739 gnd 0.003067f
C2904 vdd.n1740 gnd 0.005708f
C2905 vdd.n1741 gnd 0.005708f
C2906 vdd.n1742 gnd 0.003067f
C2907 vdd.n1743 gnd 0.003248f
C2908 vdd.n1744 gnd 0.00725f
C2909 vdd.n1745 gnd 0.00725f
C2910 vdd.n1746 gnd 0.01714f
C2911 vdd.n1747 gnd 0.003157f
C2912 vdd.n1748 gnd 0.003067f
C2913 vdd.n1749 gnd 0.014753f
C2914 vdd.n1750 gnd 0.0103f
C2915 vdd.t161 gnd 0.036084f
C2916 vdd.t271 gnd 0.036084f
C2917 vdd.n1751 gnd 0.247994f
C2918 vdd.n1752 gnd 0.195009f
C2919 vdd.t270 gnd 0.036084f
C2920 vdd.t250 gnd 0.036084f
C2921 vdd.n1753 gnd 0.247994f
C2922 vdd.n1754 gnd 0.157371f
C2923 vdd.t219 gnd 0.036084f
C2924 vdd.t158 gnd 0.036084f
C2925 vdd.n1755 gnd 0.247994f
C2926 vdd.n1756 gnd 0.157371f
C2927 vdd.t281 gnd 0.036084f
C2928 vdd.t248 gnd 0.036084f
C2929 vdd.n1757 gnd 0.247994f
C2930 vdd.n1758 gnd 0.157371f
C2931 vdd.t244 gnd 0.036084f
C2932 vdd.t193 gnd 0.036084f
C2933 vdd.n1759 gnd 0.247994f
C2934 vdd.n1760 gnd 0.157371f
C2935 vdd.t191 gnd 0.036084f
C2936 vdd.t245 gnd 0.036084f
C2937 vdd.n1761 gnd 0.247994f
C2938 vdd.n1762 gnd 0.157371f
C2939 vdd.t228 gnd 0.036084f
C2940 vdd.t229 gnd 0.036084f
C2941 vdd.n1763 gnd 0.247994f
C2942 vdd.n1764 gnd 0.157371f
C2943 vdd.t188 gnd 0.036084f
C2944 vdd.t160 gnd 0.036084f
C2945 vdd.n1765 gnd 0.247994f
C2946 vdd.n1766 gnd 0.157371f
C2947 vdd.t157 gnd 0.036084f
C2948 vdd.t225 gnd 0.036084f
C2949 vdd.n1767 gnd 0.247994f
C2950 vdd.n1768 gnd 0.157371f
C2951 vdd.n1769 gnd 0.006151f
C2952 vdd.n1770 gnd 0.005708f
C2953 vdd.n1771 gnd 0.003157f
C2954 vdd.n1772 gnd 0.00725f
C2955 vdd.n1773 gnd 0.003067f
C2956 vdd.n1774 gnd 0.003248f
C2957 vdd.n1775 gnd 0.005708f
C2958 vdd.n1776 gnd 0.003067f
C2959 vdd.n1777 gnd 0.00725f
C2960 vdd.n1778 gnd 0.003248f
C2961 vdd.n1779 gnd 0.005708f
C2962 vdd.n1780 gnd 0.003067f
C2963 vdd.n1781 gnd 0.005437f
C2964 vdd.n1782 gnd 0.005453f
C2965 vdd.t156 gnd 0.015575f
C2966 vdd.n1783 gnd 0.034655f
C2967 vdd.n1784 gnd 0.18035f
C2968 vdd.n1785 gnd 0.003067f
C2969 vdd.n1786 gnd 0.003248f
C2970 vdd.n1787 gnd 0.00725f
C2971 vdd.n1788 gnd 0.00725f
C2972 vdd.n1789 gnd 0.003248f
C2973 vdd.n1790 gnd 0.003067f
C2974 vdd.n1791 gnd 0.005708f
C2975 vdd.n1792 gnd 0.005708f
C2976 vdd.n1793 gnd 0.003067f
C2977 vdd.n1794 gnd 0.003248f
C2978 vdd.n1795 gnd 0.00725f
C2979 vdd.n1796 gnd 0.00725f
C2980 vdd.n1797 gnd 0.003248f
C2981 vdd.n1798 gnd 0.003067f
C2982 vdd.n1799 gnd 0.005708f
C2983 vdd.n1800 gnd 0.005708f
C2984 vdd.n1801 gnd 0.003067f
C2985 vdd.n1802 gnd 0.003248f
C2986 vdd.n1803 gnd 0.00725f
C2987 vdd.n1804 gnd 0.00725f
C2988 vdd.n1805 gnd 0.01714f
C2989 vdd.n1806 gnd 0.003157f
C2990 vdd.n1807 gnd 0.003067f
C2991 vdd.n1808 gnd 0.014753f
C2992 vdd.n1809 gnd 0.009977f
C2993 vdd.n1810 gnd 0.069654f
C2994 vdd.n1811 gnd 0.287319f
C2995 vdd.n1812 gnd 2.87863f
C2996 vdd.n1813 gnd 0.661084f
C2997 vdd.n1814 gnd 0.008614f
C2998 vdd.n1815 gnd 0.009021f
C2999 vdd.n1816 gnd 0.011208f
C3000 vdd.n1817 gnd 0.818956f
C3001 vdd.n1818 gnd 0.011208f
C3002 vdd.n1819 gnd 0.009021f
C3003 vdd.n1820 gnd 0.011208f
C3004 vdd.n1821 gnd 0.011208f
C3005 vdd.n1822 gnd 0.011208f
C3006 vdd.n1823 gnd 0.009021f
C3007 vdd.n1824 gnd 0.011208f
C3008 vdd.n1825 gnd 0.950677f
C3009 vdd.t221 gnd 0.572697f
C3010 vdd.n1826 gnd 0.624239f
C3011 vdd.n1827 gnd 0.011208f
C3012 vdd.n1828 gnd 0.009021f
C3013 vdd.n1829 gnd 0.011208f
C3014 vdd.n1830 gnd 0.011208f
C3015 vdd.n1831 gnd 0.011208f
C3016 vdd.n1832 gnd 0.009021f
C3017 vdd.n1833 gnd 0.011208f
C3018 vdd.n1834 gnd 0.715871f
C3019 vdd.n1835 gnd 0.011208f
C3020 vdd.n1836 gnd 0.009021f
C3021 vdd.n1837 gnd 0.011208f
C3022 vdd.n1838 gnd 0.011208f
C3023 vdd.n1839 gnd 0.011208f
C3024 vdd.n1840 gnd 0.009021f
C3025 vdd.n1841 gnd 0.011208f
C3026 vdd.n1842 gnd 0.612785f
C3027 vdd.n1843 gnd 0.910588f
C3028 vdd.n1844 gnd 0.011208f
C3029 vdd.n1845 gnd 0.009021f
C3030 vdd.n1846 gnd 0.011208f
C3031 vdd.n1847 gnd 0.011208f
C3032 vdd.n1848 gnd 0.011208f
C3033 vdd.n1849 gnd 0.009021f
C3034 vdd.n1850 gnd 0.011208f
C3035 vdd.n1851 gnd 0.950677f
C3036 vdd.n1852 gnd 0.011208f
C3037 vdd.n1853 gnd 0.009021f
C3038 vdd.n1854 gnd 0.011208f
C3039 vdd.n1855 gnd 0.011208f
C3040 vdd.n1856 gnd 0.011208f
C3041 vdd.n1857 gnd 0.009021f
C3042 vdd.n1858 gnd 0.011208f
C3043 vdd.t237 gnd 0.572697f
C3044 vdd.n1859 gnd 0.796048f
C3045 vdd.n1860 gnd 0.011208f
C3046 vdd.n1861 gnd 0.009021f
C3047 vdd.n1862 gnd 0.011208f
C3048 vdd.n1863 gnd 0.011208f
C3049 vdd.n1864 gnd 0.011208f
C3050 vdd.n1865 gnd 0.009021f
C3051 vdd.n1866 gnd 0.011208f
C3052 vdd.n1867 gnd 0.601332f
C3053 vdd.n1868 gnd 0.011208f
C3054 vdd.n1869 gnd 0.009021f
C3055 vdd.n1870 gnd 0.011208f
C3056 vdd.n1871 gnd 0.011208f
C3057 vdd.n1872 gnd 0.011208f
C3058 vdd.n1873 gnd 0.009021f
C3059 vdd.n1874 gnd 0.011208f
C3060 vdd.n1875 gnd 0.784594f
C3061 vdd.n1876 gnd 0.738779f
C3062 vdd.n1877 gnd 0.011208f
C3063 vdd.n1878 gnd 0.009021f
C3064 vdd.n1879 gnd 0.011208f
C3065 vdd.n1880 gnd 0.011208f
C3066 vdd.n1881 gnd 0.011208f
C3067 vdd.n1882 gnd 0.009021f
C3068 vdd.n1883 gnd 0.011208f
C3069 vdd.n1884 gnd 0.933496f
C3070 vdd.n1885 gnd 0.011208f
C3071 vdd.n1886 gnd 0.009021f
C3072 vdd.n1887 gnd 0.011208f
C3073 vdd.n1888 gnd 0.011208f
C3074 vdd.n1889 gnd 0.027113f
C3075 vdd.n1890 gnd 0.011208f
C3076 vdd.n1891 gnd 0.011208f
C3077 vdd.n1892 gnd 0.009021f
C3078 vdd.n1893 gnd 0.011208f
C3079 vdd.n1894 gnd 0.692963f
C3080 vdd.n1895 gnd 1.14539f
C3081 vdd.n1896 gnd 0.011208f
C3082 vdd.n1897 gnd 0.009021f
C3083 vdd.n1898 gnd 0.011208f
C3084 vdd.n1899 gnd 0.011208f
C3085 vdd.n1900 gnd 0.009639f
C3086 vdd.n1901 gnd 0.009021f
C3087 vdd.n1903 gnd 0.011208f
C3088 vdd.n1905 gnd 0.009021f
C3089 vdd.n1906 gnd 0.011208f
C3090 vdd.n1907 gnd 0.009021f
C3091 vdd.n1909 gnd 0.011208f
C3092 vdd.n1910 gnd 0.009021f
C3093 vdd.n1911 gnd 0.011208f
C3094 vdd.n1912 gnd 0.011208f
C3095 vdd.n1913 gnd 0.011208f
C3096 vdd.n1914 gnd 0.011208f
C3097 vdd.n1915 gnd 0.011208f
C3098 vdd.n1916 gnd 0.009021f
C3099 vdd.n1918 gnd 0.011208f
C3100 vdd.n1919 gnd 0.011208f
C3101 vdd.n1920 gnd 0.011208f
C3102 vdd.n1921 gnd 0.011208f
C3103 vdd.n1922 gnd 0.011208f
C3104 vdd.n1923 gnd 0.009021f
C3105 vdd.n1925 gnd 0.011208f
C3106 vdd.n1926 gnd 0.011208f
C3107 vdd.n1927 gnd 0.011208f
C3108 vdd.n1928 gnd 0.011208f
C3109 vdd.n1929 gnd 0.007533f
C3110 vdd.t68 gnd 0.137886f
C3111 vdd.t67 gnd 0.147363f
C3112 vdd.t66 gnd 0.180078f
C3113 vdd.n1930 gnd 0.230835f
C3114 vdd.n1931 gnd 0.193943f
C3115 vdd.n1933 gnd 0.011208f
C3116 vdd.n1934 gnd 0.011208f
C3117 vdd.n1935 gnd 0.009021f
C3118 vdd.n1936 gnd 0.011208f
C3119 vdd.n1938 gnd 0.011208f
C3120 vdd.n1939 gnd 0.011208f
C3121 vdd.n1940 gnd 0.011208f
C3122 vdd.n1941 gnd 0.011208f
C3123 vdd.n1942 gnd 0.009021f
C3124 vdd.n1944 gnd 0.011208f
C3125 vdd.n1945 gnd 0.011208f
C3126 vdd.n1946 gnd 0.011208f
C3127 vdd.n1947 gnd 0.011208f
C3128 vdd.n1948 gnd 0.011208f
C3129 vdd.n1949 gnd 0.009021f
C3130 vdd.n1951 gnd 0.011208f
C3131 vdd.n1952 gnd 0.011208f
C3132 vdd.n1953 gnd 0.011208f
C3133 vdd.n1954 gnd 0.011208f
C3134 vdd.n1955 gnd 0.011208f
C3135 vdd.n1956 gnd 0.009021f
C3136 vdd.n1958 gnd 0.011208f
C3137 vdd.n1959 gnd 0.011208f
C3138 vdd.n1960 gnd 0.011208f
C3139 vdd.n1961 gnd 0.011208f
C3140 vdd.n1962 gnd 0.011208f
C3141 vdd.n1963 gnd 0.009021f
C3142 vdd.n1965 gnd 0.011208f
C3143 vdd.n1966 gnd 0.011208f
C3144 vdd.n1967 gnd 0.011208f
C3145 vdd.n1968 gnd 0.011208f
C3146 vdd.n1969 gnd 0.008931f
C3147 vdd.t55 gnd 0.137886f
C3148 vdd.t54 gnd 0.147363f
C3149 vdd.t53 gnd 0.180078f
C3150 vdd.n1970 gnd 0.230835f
C3151 vdd.n1971 gnd 0.193943f
C3152 vdd.n1973 gnd 0.011208f
C3153 vdd.n1974 gnd 0.011208f
C3154 vdd.n1975 gnd 0.009021f
C3155 vdd.n1976 gnd 0.011208f
C3156 vdd.n1978 gnd 0.011208f
C3157 vdd.n1979 gnd 0.011208f
C3158 vdd.n1980 gnd 0.011208f
C3159 vdd.n1981 gnd 0.011208f
C3160 vdd.n1982 gnd 0.009021f
C3161 vdd.n1984 gnd 0.011208f
C3162 vdd.n1985 gnd 0.011208f
C3163 vdd.n1986 gnd 0.011208f
C3164 vdd.n1987 gnd 0.011208f
C3165 vdd.n1988 gnd 0.011208f
C3166 vdd.n1989 gnd 0.009021f
C3167 vdd.n1991 gnd 0.011208f
C3168 vdd.n1992 gnd 0.011208f
C3169 vdd.n1993 gnd 0.011208f
C3170 vdd.n1994 gnd 0.011208f
C3171 vdd.n1995 gnd 0.011208f
C3172 vdd.n1996 gnd 0.011208f
C3173 vdd.n1997 gnd 0.009021f
C3174 vdd.n1999 gnd 0.011208f
C3175 vdd.n2001 gnd 0.011208f
C3176 vdd.n2002 gnd 0.009021f
C3177 vdd.n2003 gnd 0.009021f
C3178 vdd.n2004 gnd 0.011208f
C3179 vdd.n2006 gnd 0.011208f
C3180 vdd.n2007 gnd 0.009021f
C3181 vdd.n2008 gnd 0.009021f
C3182 vdd.n2009 gnd 0.011208f
C3183 vdd.n2011 gnd 0.011208f
C3184 vdd.n2012 gnd 0.011208f
C3185 vdd.n2013 gnd 0.009021f
C3186 vdd.n2014 gnd 0.009021f
C3187 vdd.n2015 gnd 0.009021f
C3188 vdd.n2016 gnd 0.011208f
C3189 vdd.n2018 gnd 0.011208f
C3190 vdd.n2019 gnd 0.011208f
C3191 vdd.n2020 gnd 0.009021f
C3192 vdd.n2021 gnd 0.009021f
C3193 vdd.n2022 gnd 0.009021f
C3194 vdd.n2023 gnd 0.011208f
C3195 vdd.n2025 gnd 0.011208f
C3196 vdd.n2026 gnd 0.011208f
C3197 vdd.n2027 gnd 0.009021f
C3198 vdd.n2028 gnd 0.009021f
C3199 vdd.n2029 gnd 0.009021f
C3200 vdd.n2030 gnd 0.011208f
C3201 vdd.n2032 gnd 0.011208f
C3202 vdd.n2033 gnd 0.011208f
C3203 vdd.n2034 gnd 0.009021f
C3204 vdd.n2035 gnd 0.011208f
C3205 vdd.n2036 gnd 0.011208f
C3206 vdd.n2037 gnd 0.011208f
C3207 vdd.n2038 gnd 0.018403f
C3208 vdd.n2039 gnd 0.006134f
C3209 vdd.n2040 gnd 0.009021f
C3210 vdd.n2041 gnd 0.011208f
C3211 vdd.n2043 gnd 0.011208f
C3212 vdd.n2044 gnd 0.011208f
C3213 vdd.n2045 gnd 0.009021f
C3214 vdd.n2046 gnd 0.009021f
C3215 vdd.n2047 gnd 0.009021f
C3216 vdd.n2048 gnd 0.011208f
C3217 vdd.n2050 gnd 0.011208f
C3218 vdd.n2051 gnd 0.011208f
C3219 vdd.n2052 gnd 0.009021f
C3220 vdd.n2053 gnd 0.009021f
C3221 vdd.n2054 gnd 0.009021f
C3222 vdd.n2055 gnd 0.011208f
C3223 vdd.n2057 gnd 0.011208f
C3224 vdd.n2058 gnd 0.011208f
C3225 vdd.n2059 gnd 0.009021f
C3226 vdd.n2060 gnd 0.009021f
C3227 vdd.n2061 gnd 0.009021f
C3228 vdd.n2062 gnd 0.011208f
C3229 vdd.n2064 gnd 0.011208f
C3230 vdd.n2065 gnd 0.011208f
C3231 vdd.n2066 gnd 0.009021f
C3232 vdd.n2067 gnd 0.009021f
C3233 vdd.n2068 gnd 0.009021f
C3234 vdd.n2069 gnd 0.011208f
C3235 vdd.n2071 gnd 0.011208f
C3236 vdd.n2072 gnd 0.011208f
C3237 vdd.n2073 gnd 0.009021f
C3238 vdd.n2074 gnd 0.011208f
C3239 vdd.n2075 gnd 0.011208f
C3240 vdd.n2076 gnd 0.011208f
C3241 vdd.n2077 gnd 0.018403f
C3242 vdd.n2078 gnd 0.007533f
C3243 vdd.n2079 gnd 0.009021f
C3244 vdd.n2080 gnd 0.011208f
C3245 vdd.n2082 gnd 0.011208f
C3246 vdd.n2083 gnd 0.011208f
C3247 vdd.n2084 gnd 0.009021f
C3248 vdd.n2085 gnd 0.009021f
C3249 vdd.n2086 gnd 0.009021f
C3250 vdd.n2087 gnd 0.011208f
C3251 vdd.n2089 gnd 0.011208f
C3252 vdd.n2090 gnd 0.011208f
C3253 vdd.n2091 gnd 0.009021f
C3254 vdd.n2092 gnd 0.009021f
C3255 vdd.n2093 gnd 0.009021f
C3256 vdd.n2094 gnd 0.011208f
C3257 vdd.n2096 gnd 0.011208f
C3258 vdd.n2097 gnd 0.011208f
C3259 vdd.n2099 gnd 0.011208f
C3260 vdd.n2100 gnd 0.009021f
C3261 vdd.n2101 gnd 0.007173f
C3262 vdd.n2102 gnd 0.007621f
C3263 vdd.n2103 gnd 0.007621f
C3264 vdd.n2104 gnd 0.007621f
C3265 vdd.n2105 gnd 0.007621f
C3266 vdd.n2106 gnd 0.007621f
C3267 vdd.n2107 gnd 0.007621f
C3268 vdd.n2108 gnd 0.007621f
C3269 vdd.n2109 gnd 0.007621f
C3270 vdd.n2111 gnd 0.007621f
C3271 vdd.n2112 gnd 0.007621f
C3272 vdd.n2113 gnd 0.007621f
C3273 vdd.n2114 gnd 0.007621f
C3274 vdd.n2115 gnd 0.007621f
C3275 vdd.n2117 gnd 0.007621f
C3276 vdd.n2119 gnd 0.007621f
C3277 vdd.n2120 gnd 0.007621f
C3278 vdd.n2121 gnd 0.007621f
C3279 vdd.n2122 gnd 0.007621f
C3280 vdd.n2123 gnd 0.007621f
C3281 vdd.n2125 gnd 0.007621f
C3282 vdd.n2127 gnd 0.007621f
C3283 vdd.n2128 gnd 0.007621f
C3284 vdd.n2129 gnd 0.007621f
C3285 vdd.n2130 gnd 0.007621f
C3286 vdd.n2131 gnd 0.007621f
C3287 vdd.n2133 gnd 0.007621f
C3288 vdd.n2135 gnd 0.007621f
C3289 vdd.n2136 gnd 0.007621f
C3290 vdd.n2137 gnd 0.007621f
C3291 vdd.n2138 gnd 0.007621f
C3292 vdd.n2139 gnd 0.007621f
C3293 vdd.n2141 gnd 0.007621f
C3294 vdd.n2142 gnd 0.007621f
C3295 vdd.n2143 gnd 0.007621f
C3296 vdd.n2144 gnd 0.007621f
C3297 vdd.n2145 gnd 0.007621f
C3298 vdd.n2146 gnd 0.007621f
C3299 vdd.n2147 gnd 0.007621f
C3300 vdd.n2148 gnd 0.007621f
C3301 vdd.n2149 gnd 0.005548f
C3302 vdd.n2150 gnd 0.007621f
C3303 vdd.t108 gnd 0.307978f
C3304 vdd.t109 gnd 0.315254f
C3305 vdd.t107 gnd 0.20106f
C3306 vdd.n2151 gnd 0.108662f
C3307 vdd.n2152 gnd 0.061637f
C3308 vdd.n2153 gnd 0.010892f
C3309 vdd.n2154 gnd 0.007621f
C3310 vdd.n2155 gnd 0.007621f
C3311 vdd.n2156 gnd 0.463884f
C3312 vdd.n2157 gnd 0.007621f
C3313 vdd.n2158 gnd 0.007621f
C3314 vdd.n2159 gnd 0.007621f
C3315 vdd.n2160 gnd 0.007621f
C3316 vdd.n2161 gnd 0.007621f
C3317 vdd.n2162 gnd 0.007621f
C3318 vdd.n2163 gnd 0.007621f
C3319 vdd.n2164 gnd 0.007621f
C3320 vdd.n2165 gnd 0.007621f
C3321 vdd.n2166 gnd 0.007621f
C3322 vdd.n2167 gnd 0.007621f
C3323 vdd.n2168 gnd 0.007621f
C3324 vdd.n2169 gnd 0.007621f
C3325 vdd.n2170 gnd 0.007621f
C3326 vdd.n2171 gnd 0.007621f
C3327 vdd.n2172 gnd 0.007621f
C3328 vdd.n2173 gnd 0.007621f
C3329 vdd.n2174 gnd 0.007621f
C3330 vdd.n2175 gnd 0.007621f
C3331 vdd.n2176 gnd 0.007621f
C3332 vdd.t86 gnd 0.307978f
C3333 vdd.t87 gnd 0.315254f
C3334 vdd.t84 gnd 0.20106f
C3335 vdd.n2177 gnd 0.108662f
C3336 vdd.n2178 gnd 0.061637f
C3337 vdd.n2179 gnd 0.007621f
C3338 vdd.n2180 gnd 0.007621f
C3339 vdd.n2181 gnd 0.007621f
C3340 vdd.n2182 gnd 0.007621f
C3341 vdd.n2183 gnd 0.007621f
C3342 vdd.n2184 gnd 0.007621f
C3343 vdd.n2186 gnd 0.007621f
C3344 vdd.n2187 gnd 0.007621f
C3345 vdd.n2188 gnd 0.007621f
C3346 vdd.n2189 gnd 0.007621f
C3347 vdd.n2191 gnd 0.007621f
C3348 vdd.n2193 gnd 0.007621f
C3349 vdd.n2194 gnd 0.007621f
C3350 vdd.n2195 gnd 0.007621f
C3351 vdd.n2196 gnd 0.007621f
C3352 vdd.n2197 gnd 0.007621f
C3353 vdd.n2199 gnd 0.007621f
C3354 vdd.n2201 gnd 0.007621f
C3355 vdd.n2202 gnd 0.007621f
C3356 vdd.n2203 gnd 0.007621f
C3357 vdd.n2204 gnd 0.007621f
C3358 vdd.n2205 gnd 0.007621f
C3359 vdd.n2207 gnd 0.007621f
C3360 vdd.n2209 gnd 0.007621f
C3361 vdd.n2210 gnd 0.007621f
C3362 vdd.n2211 gnd 0.005548f
C3363 vdd.n2212 gnd 0.010892f
C3364 vdd.n2213 gnd 0.005884f
C3365 vdd.n2214 gnd 0.007621f
C3366 vdd.n2216 gnd 0.007621f
C3367 vdd.n2217 gnd 0.018084f
C3368 vdd.n2218 gnd 0.018084f
C3369 vdd.n2219 gnd 0.016885f
C3370 vdd.n2220 gnd 0.007621f
C3371 vdd.n2221 gnd 0.007621f
C3372 vdd.n2222 gnd 0.007621f
C3373 vdd.n2223 gnd 0.007621f
C3374 vdd.n2224 gnd 0.007621f
C3375 vdd.n2225 gnd 0.007621f
C3376 vdd.n2226 gnd 0.007621f
C3377 vdd.n2227 gnd 0.007621f
C3378 vdd.n2228 gnd 0.007621f
C3379 vdd.n2229 gnd 0.007621f
C3380 vdd.n2230 gnd 0.007621f
C3381 vdd.n2231 gnd 0.007621f
C3382 vdd.n2232 gnd 0.007621f
C3383 vdd.n2233 gnd 0.007621f
C3384 vdd.n2234 gnd 0.007621f
C3385 vdd.n2235 gnd 0.007621f
C3386 vdd.n2236 gnd 0.007621f
C3387 vdd.n2237 gnd 0.007621f
C3388 vdd.n2238 gnd 0.007621f
C3389 vdd.n2239 gnd 0.007621f
C3390 vdd.n2240 gnd 0.007621f
C3391 vdd.n2241 gnd 0.007621f
C3392 vdd.n2242 gnd 0.007621f
C3393 vdd.n2243 gnd 0.007621f
C3394 vdd.n2244 gnd 0.007621f
C3395 vdd.n2245 gnd 0.007621f
C3396 vdd.n2246 gnd 0.007621f
C3397 vdd.n2247 gnd 0.007621f
C3398 vdd.n2248 gnd 0.007621f
C3399 vdd.n2249 gnd 0.007621f
C3400 vdd.n2250 gnd 0.007621f
C3401 vdd.n2251 gnd 0.007621f
C3402 vdd.n2252 gnd 0.007621f
C3403 vdd.n2253 gnd 0.007621f
C3404 vdd.n2254 gnd 0.007621f
C3405 vdd.n2255 gnd 0.007621f
C3406 vdd.n2256 gnd 0.007621f
C3407 vdd.n2257 gnd 0.24626f
C3408 vdd.n2258 gnd 0.007621f
C3409 vdd.n2259 gnd 0.007621f
C3410 vdd.n2260 gnd 0.007621f
C3411 vdd.n2261 gnd 0.007621f
C3412 vdd.n2262 gnd 0.007621f
C3413 vdd.n2263 gnd 0.007621f
C3414 vdd.n2264 gnd 0.007621f
C3415 vdd.n2265 gnd 0.007621f
C3416 vdd.n2266 gnd 0.007621f
C3417 vdd.n2267 gnd 0.007621f
C3418 vdd.n2268 gnd 0.007621f
C3419 vdd.n2269 gnd 0.007621f
C3420 vdd.n2270 gnd 0.007621f
C3421 vdd.n2271 gnd 0.007621f
C3422 vdd.n2272 gnd 0.007621f
C3423 vdd.n2273 gnd 0.007621f
C3424 vdd.n2274 gnd 0.007621f
C3425 vdd.n2275 gnd 0.007621f
C3426 vdd.n2276 gnd 0.007621f
C3427 vdd.n2277 gnd 0.007621f
C3428 vdd.n2278 gnd 0.016885f
C3429 vdd.n2280 gnd 0.018084f
C3430 vdd.n2281 gnd 0.018084f
C3431 vdd.n2282 gnd 0.007621f
C3432 vdd.n2283 gnd 0.005884f
C3433 vdd.n2284 gnd 0.007621f
C3434 vdd.n2286 gnd 0.007621f
C3435 vdd.n2288 gnd 0.007621f
C3436 vdd.n2289 gnd 0.007621f
C3437 vdd.n2290 gnd 0.007621f
C3438 vdd.n2291 gnd 0.007621f
C3439 vdd.n2292 gnd 0.007621f
C3440 vdd.n2294 gnd 0.007621f
C3441 vdd.n2296 gnd 0.007621f
C3442 vdd.n2297 gnd 0.007621f
C3443 vdd.n2298 gnd 0.007621f
C3444 vdd.n2299 gnd 0.007621f
C3445 vdd.n2300 gnd 0.007621f
C3446 vdd.n2302 gnd 0.007621f
C3447 vdd.n2304 gnd 0.007621f
C3448 vdd.n2305 gnd 0.007621f
C3449 vdd.n2306 gnd 0.007621f
C3450 vdd.n2307 gnd 0.007621f
C3451 vdd.n2308 gnd 0.007621f
C3452 vdd.n2310 gnd 0.007621f
C3453 vdd.n2312 gnd 0.007621f
C3454 vdd.n2313 gnd 0.007621f
C3455 vdd.n2314 gnd 0.022733f
C3456 vdd.n2315 gnd 0.673901f
C3457 vdd.n2317 gnd 0.009021f
C3458 vdd.n2318 gnd 0.009021f
C3459 vdd.n2319 gnd 0.011208f
C3460 vdd.n2321 gnd 0.011208f
C3461 vdd.n2322 gnd 0.011208f
C3462 vdd.n2323 gnd 0.009021f
C3463 vdd.n2324 gnd 0.007487f
C3464 vdd.n2325 gnd 0.027694f
C3465 vdd.n2326 gnd 0.027113f
C3466 vdd.n2327 gnd 0.007487f
C3467 vdd.n2328 gnd 0.027113f
C3468 vdd.n2329 gnd 1.57492f
C3469 vdd.n2330 gnd 0.027113f
C3470 vdd.n2331 gnd 0.027694f
C3471 vdd.n2332 gnd 0.004285f
C3472 vdd.t44 gnd 0.137886f
C3473 vdd.t43 gnd 0.147363f
C3474 vdd.t41 gnd 0.180078f
C3475 vdd.n2333 gnd 0.230835f
C3476 vdd.n2334 gnd 0.193943f
C3477 vdd.n2335 gnd 0.013892f
C3478 vdd.n2336 gnd 0.004736f
C3479 vdd.n2337 gnd 0.009639f
C3480 vdd.n2338 gnd 0.673901f
C3481 vdd.n2339 gnd 0.022733f
C3482 vdd.n2340 gnd 0.007621f
C3483 vdd.n2341 gnd 0.007621f
C3484 vdd.n2342 gnd 0.007621f
C3485 vdd.n2344 gnd 0.007621f
C3486 vdd.n2346 gnd 0.007621f
C3487 vdd.n2347 gnd 0.007621f
C3488 vdd.n2348 gnd 0.007621f
C3489 vdd.n2349 gnd 0.007621f
C3490 vdd.n2350 gnd 0.007621f
C3491 vdd.n2352 gnd 0.007621f
C3492 vdd.n2354 gnd 0.007621f
C3493 vdd.n2355 gnd 0.007621f
C3494 vdd.n2356 gnd 0.007621f
C3495 vdd.n2357 gnd 0.007621f
C3496 vdd.n2358 gnd 0.007621f
C3497 vdd.n2360 gnd 0.007621f
C3498 vdd.n2362 gnd 0.007621f
C3499 vdd.n2363 gnd 0.007621f
C3500 vdd.n2364 gnd 0.007621f
C3501 vdd.n2365 gnd 0.007621f
C3502 vdd.n2366 gnd 0.007621f
C3503 vdd.n2368 gnd 0.007621f
C3504 vdd.n2370 gnd 0.007621f
C3505 vdd.n2371 gnd 0.007621f
C3506 vdd.n2372 gnd 0.018084f
C3507 vdd.n2373 gnd 0.016885f
C3508 vdd.n2374 gnd 0.016885f
C3509 vdd.n2375 gnd 1.12249f
C3510 vdd.n2376 gnd 0.016885f
C3511 vdd.n2377 gnd 0.016885f
C3512 vdd.n2378 gnd 0.007621f
C3513 vdd.n2379 gnd 0.007621f
C3514 vdd.n2380 gnd 0.007621f
C3515 vdd.n2381 gnd 0.486792f
C3516 vdd.n2382 gnd 0.007621f
C3517 vdd.n2383 gnd 0.007621f
C3518 vdd.n2384 gnd 0.007621f
C3519 vdd.n2385 gnd 0.007621f
C3520 vdd.n2386 gnd 0.007621f
C3521 vdd.n2387 gnd 0.778867f
C3522 vdd.n2388 gnd 0.007621f
C3523 vdd.n2389 gnd 0.007621f
C3524 vdd.n2390 gnd 0.007621f
C3525 vdd.n2391 gnd 0.007621f
C3526 vdd.n2392 gnd 0.007621f
C3527 vdd.n2393 gnd 0.778867f
C3528 vdd.n2394 gnd 0.007621f
C3529 vdd.n2395 gnd 0.007621f
C3530 vdd.n2396 gnd 0.006725f
C3531 vdd.n2397 gnd 0.022078f
C3532 vdd.n2398 gnd 0.004707f
C3533 vdd.n2399 gnd 0.007621f
C3534 vdd.n2400 gnd 0.429523f
C3535 vdd.n2401 gnd 0.007621f
C3536 vdd.n2402 gnd 0.007621f
C3537 vdd.n2403 gnd 0.007621f
C3538 vdd.n2404 gnd 0.007621f
C3539 vdd.n2405 gnd 0.007621f
C3540 vdd.n2406 gnd 0.521154f
C3541 vdd.n2407 gnd 0.007621f
C3542 vdd.n2408 gnd 0.007621f
C3543 vdd.n2409 gnd 0.007621f
C3544 vdd.n2410 gnd 0.007621f
C3545 vdd.n2411 gnd 0.007621f
C3546 vdd.n2412 gnd 0.692963f
C3547 vdd.n2413 gnd 0.007621f
C3548 vdd.n2414 gnd 0.007621f
C3549 vdd.n2415 gnd 0.007621f
C3550 vdd.n2416 gnd 0.007621f
C3551 vdd.n2417 gnd 0.007621f
C3552 vdd.n2418 gnd 0.618512f
C3553 vdd.n2419 gnd 0.007621f
C3554 vdd.n2420 gnd 0.007621f
C3555 vdd.n2421 gnd 0.007621f
C3556 vdd.n2422 gnd 0.007621f
C3557 vdd.n2423 gnd 0.007621f
C3558 vdd.n2424 gnd 0.446703f
C3559 vdd.n2425 gnd 0.007621f
C3560 vdd.n2426 gnd 0.007621f
C3561 vdd.n2427 gnd 0.007621f
C3562 vdd.n2428 gnd 0.007621f
C3563 vdd.n2429 gnd 0.007621f
C3564 vdd.n2430 gnd 0.24626f
C3565 vdd.n2431 gnd 0.007621f
C3566 vdd.n2432 gnd 0.007621f
C3567 vdd.n2433 gnd 0.007621f
C3568 vdd.n2434 gnd 0.007621f
C3569 vdd.n2435 gnd 0.007621f
C3570 vdd.n2436 gnd 0.429523f
C3571 vdd.n2437 gnd 0.007621f
C3572 vdd.n2438 gnd 0.007621f
C3573 vdd.n2439 gnd 0.007621f
C3574 vdd.n2440 gnd 0.007621f
C3575 vdd.n2441 gnd 0.007621f
C3576 vdd.n2442 gnd 0.778867f
C3577 vdd.n2443 gnd 0.007621f
C3578 vdd.n2444 gnd 0.007621f
C3579 vdd.n2445 gnd 0.007621f
C3580 vdd.n2446 gnd 0.007621f
C3581 vdd.n2447 gnd 0.007621f
C3582 vdd.n2448 gnd 0.007621f
C3583 vdd.n2449 gnd 0.007621f
C3584 vdd.n2450 gnd 0.607058f
C3585 vdd.n2451 gnd 0.007621f
C3586 vdd.n2452 gnd 0.007621f
C3587 vdd.n2453 gnd 0.007621f
C3588 vdd.n2454 gnd 0.007621f
C3589 vdd.n2455 gnd 0.007621f
C3590 vdd.n2456 gnd 0.007621f
C3591 vdd.n2457 gnd 0.486792f
C3592 vdd.n2458 gnd 0.007621f
C3593 vdd.n2459 gnd 0.007621f
C3594 vdd.n2460 gnd 0.007621f
C3595 vdd.n2461 gnd 0.017813f
C3596 vdd.n2462 gnd 0.017156f
C3597 vdd.n2463 gnd 0.007621f
C3598 vdd.n2464 gnd 0.007621f
C3599 vdd.n2465 gnd 0.005884f
C3600 vdd.n2466 gnd 0.007621f
C3601 vdd.n2467 gnd 0.007621f
C3602 vdd.n2468 gnd 0.005548f
C3603 vdd.n2469 gnd 0.007621f
C3604 vdd.n2470 gnd 0.007621f
C3605 vdd.n2471 gnd 0.007621f
C3606 vdd.n2472 gnd 0.007621f
C3607 vdd.n2473 gnd 0.007621f
C3608 vdd.n2474 gnd 0.007621f
C3609 vdd.n2475 gnd 0.007621f
C3610 vdd.n2476 gnd 0.007621f
C3611 vdd.n2477 gnd 0.007621f
C3612 vdd.n2478 gnd 0.007621f
C3613 vdd.n2479 gnd 0.007621f
C3614 vdd.n2480 gnd 0.007621f
C3615 vdd.n2481 gnd 0.007621f
C3616 vdd.n2482 gnd 0.007621f
C3617 vdd.n2483 gnd 0.007621f
C3618 vdd.n2484 gnd 0.007621f
C3619 vdd.n2485 gnd 0.007621f
C3620 vdd.n2486 gnd 0.007621f
C3621 vdd.n2487 gnd 0.007621f
C3622 vdd.n2488 gnd 0.007621f
C3623 vdd.n2489 gnd 0.007621f
C3624 vdd.n2490 gnd 0.007621f
C3625 vdd.n2491 gnd 0.007621f
C3626 vdd.n2492 gnd 0.007621f
C3627 vdd.n2493 gnd 0.007621f
C3628 vdd.n2494 gnd 0.007621f
C3629 vdd.n2495 gnd 0.007621f
C3630 vdd.n2496 gnd 0.007621f
C3631 vdd.n2497 gnd 0.007621f
C3632 vdd.n2498 gnd 0.007621f
C3633 vdd.n2499 gnd 0.007621f
C3634 vdd.n2500 gnd 0.007621f
C3635 vdd.n2501 gnd 0.007621f
C3636 vdd.n2502 gnd 0.007621f
C3637 vdd.n2503 gnd 0.007621f
C3638 vdd.n2504 gnd 0.007621f
C3639 vdd.n2505 gnd 0.007621f
C3640 vdd.n2506 gnd 0.007621f
C3641 vdd.n2507 gnd 0.007621f
C3642 vdd.n2508 gnd 0.007621f
C3643 vdd.n2509 gnd 0.007621f
C3644 vdd.n2510 gnd 0.007621f
C3645 vdd.n2511 gnd 0.007621f
C3646 vdd.n2512 gnd 0.007621f
C3647 vdd.n2513 gnd 0.007621f
C3648 vdd.n2514 gnd 0.007621f
C3649 vdd.n2515 gnd 0.007621f
C3650 vdd.n2516 gnd 0.007621f
C3651 vdd.n2517 gnd 0.007621f
C3652 vdd.n2518 gnd 0.007621f
C3653 vdd.n2519 gnd 0.007621f
C3654 vdd.n2520 gnd 0.007621f
C3655 vdd.n2521 gnd 0.007621f
C3656 vdd.n2522 gnd 0.007621f
C3657 vdd.n2523 gnd 0.007621f
C3658 vdd.n2524 gnd 0.007621f
C3659 vdd.n2525 gnd 0.007621f
C3660 vdd.n2526 gnd 0.007621f
C3661 vdd.n2527 gnd 0.007621f
C3662 vdd.n2528 gnd 0.007621f
C3663 vdd.n2529 gnd 0.018084f
C3664 vdd.n2530 gnd 0.016885f
C3665 vdd.n2531 gnd 0.016885f
C3666 vdd.n2532 gnd 0.950677f
C3667 vdd.n2533 gnd 0.016885f
C3668 vdd.n2534 gnd 0.018084f
C3669 vdd.n2535 gnd 0.017156f
C3670 vdd.n2536 gnd 0.007621f
C3671 vdd.n2537 gnd 0.007621f
C3672 vdd.n2538 gnd 0.007621f
C3673 vdd.n2539 gnd 0.005884f
C3674 vdd.n2540 gnd 0.010892f
C3675 vdd.n2541 gnd 0.005548f
C3676 vdd.n2542 gnd 0.007621f
C3677 vdd.n2543 gnd 0.007621f
C3678 vdd.n2544 gnd 0.007621f
C3679 vdd.n2545 gnd 0.007621f
C3680 vdd.n2546 gnd 0.007621f
C3681 vdd.n2547 gnd 0.007621f
C3682 vdd.n2548 gnd 0.007621f
C3683 vdd.n2549 gnd 0.007621f
C3684 vdd.n2550 gnd 0.007621f
C3685 vdd.n2551 gnd 0.007621f
C3686 vdd.n2552 gnd 0.007621f
C3687 vdd.n2553 gnd 0.007621f
C3688 vdd.n2554 gnd 0.007621f
C3689 vdd.n2555 gnd 0.007621f
C3690 vdd.n2556 gnd 0.007621f
C3691 vdd.n2557 gnd 0.007621f
C3692 vdd.n2558 gnd 0.007621f
C3693 vdd.n2559 gnd 0.007621f
C3694 vdd.n2560 gnd 0.007621f
C3695 vdd.n2561 gnd 0.007621f
C3696 vdd.n2562 gnd 0.007621f
C3697 vdd.n2563 gnd 0.007621f
C3698 vdd.n2564 gnd 0.007621f
C3699 vdd.n2565 gnd 0.007621f
C3700 vdd.n2566 gnd 0.007621f
C3701 vdd.n2567 gnd 0.007621f
C3702 vdd.n2568 gnd 0.007621f
C3703 vdd.n2569 gnd 0.007621f
C3704 vdd.n2570 gnd 0.007621f
C3705 vdd.n2571 gnd 0.007621f
C3706 vdd.n2572 gnd 0.007621f
C3707 vdd.n2573 gnd 0.007621f
C3708 vdd.n2574 gnd 0.007621f
C3709 vdd.n2575 gnd 0.007621f
C3710 vdd.n2576 gnd 0.007621f
C3711 vdd.n2577 gnd 0.007621f
C3712 vdd.n2578 gnd 0.007621f
C3713 vdd.n2579 gnd 0.007621f
C3714 vdd.n2580 gnd 0.007621f
C3715 vdd.n2581 gnd 0.007621f
C3716 vdd.n2582 gnd 0.007621f
C3717 vdd.n2583 gnd 0.007621f
C3718 vdd.n2584 gnd 0.007621f
C3719 vdd.n2585 gnd 0.007621f
C3720 vdd.n2586 gnd 0.007621f
C3721 vdd.n2587 gnd 0.007621f
C3722 vdd.n2588 gnd 0.007621f
C3723 vdd.n2589 gnd 0.007621f
C3724 vdd.n2590 gnd 0.007621f
C3725 vdd.n2591 gnd 0.007621f
C3726 vdd.n2592 gnd 0.007621f
C3727 vdd.n2593 gnd 0.007621f
C3728 vdd.n2594 gnd 0.007621f
C3729 vdd.n2595 gnd 0.007621f
C3730 vdd.n2596 gnd 0.007621f
C3731 vdd.n2597 gnd 0.007621f
C3732 vdd.n2598 gnd 0.007621f
C3733 vdd.n2599 gnd 0.007621f
C3734 vdd.n2600 gnd 0.007621f
C3735 vdd.n2601 gnd 0.007621f
C3736 vdd.n2602 gnd 0.018084f
C3737 vdd.n2603 gnd 0.018084f
C3738 vdd.n2604 gnd 0.950677f
C3739 vdd.t286 gnd 3.37891f
C3740 vdd.t111 gnd 3.37891f
C3741 vdd.n2637 gnd 0.018084f
C3742 vdd.n2638 gnd 0.007621f
C3743 vdd.t79 gnd 0.307978f
C3744 vdd.t80 gnd 0.315254f
C3745 vdd.t77 gnd 0.20106f
C3746 vdd.n2639 gnd 0.108662f
C3747 vdd.n2640 gnd 0.061637f
C3748 vdd.n2641 gnd 0.007621f
C3749 vdd.t93 gnd 0.307978f
C3750 vdd.t94 gnd 0.315254f
C3751 vdd.t92 gnd 0.20106f
C3752 vdd.n2642 gnd 0.108662f
C3753 vdd.n2643 gnd 0.061637f
C3754 vdd.n2644 gnd 0.010892f
C3755 vdd.n2645 gnd 0.007621f
C3756 vdd.n2646 gnd 0.007621f
C3757 vdd.n2647 gnd 0.007621f
C3758 vdd.n2648 gnd 0.007621f
C3759 vdd.n2649 gnd 0.007621f
C3760 vdd.n2650 gnd 0.007621f
C3761 vdd.n2651 gnd 0.007621f
C3762 vdd.n2652 gnd 0.007621f
C3763 vdd.n2653 gnd 0.007621f
C3764 vdd.n2654 gnd 0.007621f
C3765 vdd.n2655 gnd 0.007621f
C3766 vdd.n2656 gnd 0.007621f
C3767 vdd.n2657 gnd 0.007621f
C3768 vdd.n2658 gnd 0.007621f
C3769 vdd.n2659 gnd 0.007621f
C3770 vdd.n2660 gnd 0.007621f
C3771 vdd.n2661 gnd 0.007621f
C3772 vdd.n2662 gnd 0.007621f
C3773 vdd.n2663 gnd 0.007621f
C3774 vdd.n2664 gnd 0.007621f
C3775 vdd.n2665 gnd 0.007621f
C3776 vdd.n2666 gnd 0.007621f
C3777 vdd.n2667 gnd 0.007621f
C3778 vdd.n2668 gnd 0.007621f
C3779 vdd.n2669 gnd 0.007621f
C3780 vdd.n2670 gnd 0.007621f
C3781 vdd.n2671 gnd 0.007621f
C3782 vdd.n2672 gnd 0.007621f
C3783 vdd.n2673 gnd 0.007621f
C3784 vdd.n2674 gnd 0.007621f
C3785 vdd.n2675 gnd 0.007621f
C3786 vdd.n2676 gnd 0.007621f
C3787 vdd.n2677 gnd 0.007621f
C3788 vdd.n2678 gnd 0.007621f
C3789 vdd.n2679 gnd 0.007621f
C3790 vdd.n2680 gnd 0.007621f
C3791 vdd.n2681 gnd 0.007621f
C3792 vdd.n2682 gnd 0.007621f
C3793 vdd.n2683 gnd 0.007621f
C3794 vdd.n2684 gnd 0.007621f
C3795 vdd.n2685 gnd 0.007621f
C3796 vdd.n2686 gnd 0.007621f
C3797 vdd.n2687 gnd 0.007621f
C3798 vdd.n2688 gnd 0.007621f
C3799 vdd.n2689 gnd 0.007621f
C3800 vdd.n2690 gnd 0.007621f
C3801 vdd.n2691 gnd 0.007621f
C3802 vdd.n2692 gnd 0.007621f
C3803 vdd.n2693 gnd 0.007621f
C3804 vdd.n2694 gnd 0.007621f
C3805 vdd.n2695 gnd 0.007621f
C3806 vdd.n2696 gnd 0.007621f
C3807 vdd.n2697 gnd 0.007621f
C3808 vdd.n2698 gnd 0.007621f
C3809 vdd.n2699 gnd 0.007621f
C3810 vdd.n2700 gnd 0.007621f
C3811 vdd.n2701 gnd 0.005548f
C3812 vdd.n2702 gnd 0.007621f
C3813 vdd.n2703 gnd 0.007621f
C3814 vdd.n2704 gnd 0.005884f
C3815 vdd.n2705 gnd 0.007621f
C3816 vdd.n2706 gnd 0.007621f
C3817 vdd.n2707 gnd 0.018084f
C3818 vdd.n2708 gnd 0.016885f
C3819 vdd.n2709 gnd 0.007621f
C3820 vdd.n2710 gnd 0.007621f
C3821 vdd.n2711 gnd 0.007621f
C3822 vdd.n2712 gnd 0.007621f
C3823 vdd.n2713 gnd 0.007621f
C3824 vdd.n2714 gnd 0.007621f
C3825 vdd.n2715 gnd 0.007621f
C3826 vdd.n2716 gnd 0.007621f
C3827 vdd.n2717 gnd 0.007621f
C3828 vdd.n2718 gnd 0.007621f
C3829 vdd.n2719 gnd 0.007621f
C3830 vdd.n2720 gnd 0.007621f
C3831 vdd.n2721 gnd 0.007621f
C3832 vdd.n2722 gnd 0.007621f
C3833 vdd.n2723 gnd 0.007621f
C3834 vdd.n2724 gnd 0.007621f
C3835 vdd.n2725 gnd 0.007621f
C3836 vdd.n2726 gnd 0.007621f
C3837 vdd.n2727 gnd 0.007621f
C3838 vdd.n2728 gnd 0.007621f
C3839 vdd.n2729 gnd 0.007621f
C3840 vdd.n2730 gnd 0.007621f
C3841 vdd.n2731 gnd 0.007621f
C3842 vdd.n2732 gnd 0.007621f
C3843 vdd.n2733 gnd 0.007621f
C3844 vdd.n2734 gnd 0.007621f
C3845 vdd.n2735 gnd 0.007621f
C3846 vdd.n2736 gnd 0.007621f
C3847 vdd.n2737 gnd 0.007621f
C3848 vdd.n2738 gnd 0.007621f
C3849 vdd.n2739 gnd 0.007621f
C3850 vdd.n2740 gnd 0.007621f
C3851 vdd.n2741 gnd 0.007621f
C3852 vdd.n2742 gnd 0.007621f
C3853 vdd.n2743 gnd 0.007621f
C3854 vdd.n2744 gnd 0.007621f
C3855 vdd.n2745 gnd 0.007621f
C3856 vdd.n2746 gnd 0.007621f
C3857 vdd.n2747 gnd 0.007621f
C3858 vdd.n2748 gnd 0.007621f
C3859 vdd.n2749 gnd 0.007621f
C3860 vdd.n2750 gnd 0.007621f
C3861 vdd.n2751 gnd 0.007621f
C3862 vdd.n2752 gnd 0.007621f
C3863 vdd.n2753 gnd 0.007621f
C3864 vdd.n2754 gnd 0.007621f
C3865 vdd.n2755 gnd 0.007621f
C3866 vdd.n2756 gnd 0.007621f
C3867 vdd.n2757 gnd 0.007621f
C3868 vdd.n2758 gnd 0.007621f
C3869 vdd.n2759 gnd 0.007621f
C3870 vdd.n2760 gnd 0.24626f
C3871 vdd.n2761 gnd 0.007621f
C3872 vdd.n2762 gnd 0.007621f
C3873 vdd.n2763 gnd 0.007621f
C3874 vdd.n2764 gnd 0.007621f
C3875 vdd.n2765 gnd 0.007621f
C3876 vdd.n2766 gnd 0.007621f
C3877 vdd.n2767 gnd 0.007621f
C3878 vdd.n2768 gnd 0.007621f
C3879 vdd.n2769 gnd 0.007621f
C3880 vdd.n2770 gnd 0.007621f
C3881 vdd.n2771 gnd 0.007621f
C3882 vdd.n2772 gnd 0.007621f
C3883 vdd.n2773 gnd 0.007621f
C3884 vdd.n2774 gnd 0.007621f
C3885 vdd.n2775 gnd 0.007621f
C3886 vdd.n2776 gnd 0.007621f
C3887 vdd.n2777 gnd 0.007621f
C3888 vdd.n2778 gnd 0.007621f
C3889 vdd.n2779 gnd 0.007621f
C3890 vdd.n2780 gnd 0.007621f
C3891 vdd.n2781 gnd 0.463884f
C3892 vdd.n2782 gnd 0.007621f
C3893 vdd.n2783 gnd 0.007621f
C3894 vdd.n2784 gnd 0.007621f
C3895 vdd.n2785 gnd 0.007621f
C3896 vdd.n2786 gnd 0.007621f
C3897 vdd.n2787 gnd 0.016885f
C3898 vdd.n2788 gnd 0.018084f
C3899 vdd.n2789 gnd 0.018084f
C3900 vdd.n2790 gnd 0.007621f
C3901 vdd.n2791 gnd 0.007621f
C3902 vdd.n2792 gnd 0.007621f
C3903 vdd.n2793 gnd 0.005884f
C3904 vdd.n2794 gnd 0.010892f
C3905 vdd.n2795 gnd 0.005548f
C3906 vdd.n2796 gnd 0.007621f
C3907 vdd.n2797 gnd 0.007621f
C3908 vdd.n2798 gnd 0.007621f
C3909 vdd.n2799 gnd 0.007621f
C3910 vdd.n2800 gnd 0.007621f
C3911 vdd.n2801 gnd 0.007621f
C3912 vdd.n2802 gnd 0.007621f
C3913 vdd.n2803 gnd 0.007621f
C3914 vdd.n2804 gnd 0.007621f
C3915 vdd.n2805 gnd 0.007621f
C3916 vdd.n2806 gnd 0.007621f
C3917 vdd.n2807 gnd 0.007621f
C3918 vdd.n2808 gnd 0.007621f
C3919 vdd.n2809 gnd 0.007621f
C3920 vdd.n2810 gnd 0.007621f
C3921 vdd.n2811 gnd 0.007621f
C3922 vdd.n2812 gnd 0.007621f
C3923 vdd.n2813 gnd 0.007621f
C3924 vdd.n2814 gnd 0.007621f
C3925 vdd.n2815 gnd 0.007621f
C3926 vdd.n2816 gnd 0.007621f
C3927 vdd.n2817 gnd 0.007621f
C3928 vdd.n2818 gnd 0.007621f
C3929 vdd.n2819 gnd 0.007621f
C3930 vdd.n2820 gnd 0.007621f
C3931 vdd.n2821 gnd 0.007621f
C3932 vdd.n2822 gnd 0.007621f
C3933 vdd.n2823 gnd 0.007621f
C3934 vdd.n2824 gnd 0.007621f
C3935 vdd.n2825 gnd 0.007621f
C3936 vdd.n2826 gnd 0.007621f
C3937 vdd.n2827 gnd 0.007621f
C3938 vdd.n2828 gnd 0.007621f
C3939 vdd.n2829 gnd 0.007621f
C3940 vdd.n2830 gnd 0.007621f
C3941 vdd.n2831 gnd 0.007621f
C3942 vdd.n2832 gnd 0.007621f
C3943 vdd.n2833 gnd 0.007621f
C3944 vdd.n2834 gnd 0.007621f
C3945 vdd.n2835 gnd 0.007621f
C3946 vdd.n2836 gnd 0.007621f
C3947 vdd.n2837 gnd 0.007621f
C3948 vdd.n2838 gnd 0.007621f
C3949 vdd.n2839 gnd 0.007621f
C3950 vdd.n2840 gnd 0.007621f
C3951 vdd.n2841 gnd 0.007621f
C3952 vdd.n2842 gnd 0.007621f
C3953 vdd.n2843 gnd 0.007621f
C3954 vdd.n2844 gnd 0.007621f
C3955 vdd.n2845 gnd 0.007621f
C3956 vdd.n2846 gnd 0.007621f
C3957 vdd.n2847 gnd 0.007621f
C3958 vdd.n2848 gnd 0.007621f
C3959 vdd.n2849 gnd 0.007621f
C3960 vdd.n2850 gnd 0.007621f
C3961 vdd.n2851 gnd 0.007621f
C3962 vdd.n2852 gnd 0.007621f
C3963 vdd.n2853 gnd 0.007621f
C3964 vdd.n2854 gnd 0.007621f
C3965 vdd.n2855 gnd 0.007621f
C3966 vdd.n2857 gnd 0.950677f
C3967 vdd.n2859 gnd 0.007621f
C3968 vdd.n2860 gnd 0.007621f
C3969 vdd.n2861 gnd 0.018084f
C3970 vdd.n2862 gnd 0.016885f
C3971 vdd.n2863 gnd 0.016885f
C3972 vdd.n2864 gnd 0.950677f
C3973 vdd.n2865 gnd 0.016885f
C3974 vdd.n2866 gnd 0.016885f
C3975 vdd.n2867 gnd 0.007621f
C3976 vdd.n2868 gnd 0.007621f
C3977 vdd.n2869 gnd 0.007621f
C3978 vdd.n2870 gnd 0.486792f
C3979 vdd.n2871 gnd 0.007621f
C3980 vdd.n2872 gnd 0.007621f
C3981 vdd.n2873 gnd 0.007621f
C3982 vdd.n2874 gnd 0.007621f
C3983 vdd.n2875 gnd 0.007621f
C3984 vdd.n2876 gnd 0.607058f
C3985 vdd.n2877 gnd 0.007621f
C3986 vdd.n2878 gnd 0.007621f
C3987 vdd.n2879 gnd 0.007621f
C3988 vdd.n2880 gnd 0.007621f
C3989 vdd.n2881 gnd 0.007621f
C3990 vdd.n2882 gnd 0.778867f
C3991 vdd.n2883 gnd 0.007621f
C3992 vdd.n2884 gnd 0.007621f
C3993 vdd.n2885 gnd 0.007621f
C3994 vdd.n2886 gnd 0.007621f
C3995 vdd.n2887 gnd 0.007621f
C3996 vdd.n2888 gnd 0.429523f
C3997 vdd.n2889 gnd 0.007621f
C3998 vdd.n2890 gnd 0.007621f
C3999 vdd.n2891 gnd 0.007621f
C4000 vdd.n2892 gnd 0.007621f
C4001 vdd.n2893 gnd 0.007621f
C4002 vdd.n2894 gnd 0.24626f
C4003 vdd.n2895 gnd 0.007621f
C4004 vdd.n2896 gnd 0.007621f
C4005 vdd.n2897 gnd 0.007621f
C4006 vdd.n2898 gnd 0.007621f
C4007 vdd.n2899 gnd 0.007621f
C4008 vdd.n2900 gnd 0.446703f
C4009 vdd.n2901 gnd 0.007621f
C4010 vdd.n2902 gnd 0.007621f
C4011 vdd.n2903 gnd 0.007621f
C4012 vdd.n2904 gnd 0.007621f
C4013 vdd.n2905 gnd 0.007621f
C4014 vdd.n2906 gnd 0.618512f
C4015 vdd.n2907 gnd 0.007621f
C4016 vdd.n2908 gnd 0.007621f
C4017 vdd.n2909 gnd 0.007621f
C4018 vdd.n2910 gnd 0.007621f
C4019 vdd.n2911 gnd 0.007621f
C4020 vdd.n2912 gnd 0.692963f
C4021 vdd.n2913 gnd 0.007621f
C4022 vdd.n2914 gnd 0.007621f
C4023 vdd.n2915 gnd 0.007621f
C4024 vdd.n2916 gnd 0.007621f
C4025 vdd.n2917 gnd 0.007621f
C4026 vdd.n2918 gnd 0.521154f
C4027 vdd.n2919 gnd 0.007621f
C4028 vdd.n2920 gnd 0.007621f
C4029 vdd.n2921 gnd 0.007621f
C4030 vdd.t47 gnd 0.315254f
C4031 vdd.t45 gnd 0.20106f
C4032 vdd.t48 gnd 0.315254f
C4033 vdd.n2922 gnd 0.177186f
C4034 vdd.n2923 gnd 0.022078f
C4035 vdd.n2924 gnd 0.004707f
C4036 vdd.n2925 gnd 0.007621f
C4037 vdd.n2926 gnd 0.429523f
C4038 vdd.n2927 gnd 0.007621f
C4039 vdd.n2928 gnd 0.007621f
C4040 vdd.n2929 gnd 0.007621f
C4041 vdd.n2930 gnd 0.007621f
C4042 vdd.n2931 gnd 0.007621f
C4043 vdd.n2932 gnd 0.778867f
C4044 vdd.n2933 gnd 0.007621f
C4045 vdd.n2934 gnd 0.007621f
C4046 vdd.n2935 gnd 0.007621f
C4047 vdd.n2936 gnd 0.007621f
C4048 vdd.n2937 gnd 0.007621f
C4049 vdd.n2938 gnd 0.007621f
C4050 vdd.n2940 gnd 0.007621f
C4051 vdd.n2941 gnd 0.007621f
C4052 vdd.n2943 gnd 0.007621f
C4053 vdd.n2944 gnd 0.007621f
C4054 vdd.n2947 gnd 0.007621f
C4055 vdd.n2948 gnd 0.007621f
C4056 vdd.n2949 gnd 0.007621f
C4057 vdd.n2950 gnd 0.007621f
C4058 vdd.n2952 gnd 0.007621f
C4059 vdd.n2953 gnd 0.007621f
C4060 vdd.n2954 gnd 0.007621f
C4061 vdd.n2955 gnd 0.007621f
C4062 vdd.n2956 gnd 0.007621f
C4063 vdd.n2957 gnd 0.007621f
C4064 vdd.n2959 gnd 0.007621f
C4065 vdd.n2960 gnd 0.007621f
C4066 vdd.n2961 gnd 0.007621f
C4067 vdd.n2962 gnd 0.007621f
C4068 vdd.n2963 gnd 0.007621f
C4069 vdd.n2964 gnd 0.007621f
C4070 vdd.n2966 gnd 0.007621f
C4071 vdd.n2967 gnd 0.007621f
C4072 vdd.n2968 gnd 0.007621f
C4073 vdd.n2969 gnd 0.007621f
C4074 vdd.n2970 gnd 0.007621f
C4075 vdd.n2971 gnd 0.007621f
C4076 vdd.n2973 gnd 0.007621f
C4077 vdd.n2974 gnd 0.018084f
C4078 vdd.n2975 gnd 0.018084f
C4079 vdd.n2976 gnd 0.016885f
C4080 vdd.n2977 gnd 0.007621f
C4081 vdd.n2978 gnd 0.007621f
C4082 vdd.n2979 gnd 0.007621f
C4083 vdd.n2980 gnd 0.007621f
C4084 vdd.n2981 gnd 0.007621f
C4085 vdd.n2982 gnd 0.007621f
C4086 vdd.n2983 gnd 0.778867f
C4087 vdd.n2984 gnd 0.007621f
C4088 vdd.n2985 gnd 0.007621f
C4089 vdd.n2986 gnd 0.007621f
C4090 vdd.n2987 gnd 0.007621f
C4091 vdd.n2988 gnd 0.007621f
C4092 vdd.n2989 gnd 0.486792f
C4093 vdd.n2990 gnd 0.007621f
C4094 vdd.n2991 gnd 0.007621f
C4095 vdd.n2992 gnd 0.007621f
C4096 vdd.n2993 gnd 0.017813f
C4097 vdd.n2994 gnd 0.017156f
C4098 vdd.n2995 gnd 0.018084f
C4099 vdd.n2997 gnd 0.007621f
C4100 vdd.n2998 gnd 0.007621f
C4101 vdd.n2999 gnd 0.005884f
C4102 vdd.n3000 gnd 0.010892f
C4103 vdd.n3001 gnd 0.005548f
C4104 vdd.n3002 gnd 0.007621f
C4105 vdd.n3003 gnd 0.007621f
C4106 vdd.n3005 gnd 0.007621f
C4107 vdd.n3006 gnd 0.007621f
C4108 vdd.n3007 gnd 0.007621f
C4109 vdd.n3008 gnd 0.007621f
C4110 vdd.n3009 gnd 0.007621f
C4111 vdd.n3010 gnd 0.007621f
C4112 vdd.n3012 gnd 0.007621f
C4113 vdd.n3013 gnd 0.007621f
C4114 vdd.n3014 gnd 0.007621f
C4115 vdd.n3015 gnd 0.007621f
C4116 vdd.n3016 gnd 0.007621f
C4117 vdd.n3017 gnd 0.007621f
C4118 vdd.n3019 gnd 0.007621f
C4119 vdd.n3020 gnd 0.007621f
C4120 vdd.n3021 gnd 0.007621f
C4121 vdd.n3022 gnd 0.007621f
C4122 vdd.n3023 gnd 0.007621f
C4123 vdd.n3024 gnd 0.007621f
C4124 vdd.n3026 gnd 0.007621f
C4125 vdd.n3027 gnd 0.007621f
C4126 vdd.n3028 gnd 0.007621f
C4127 vdd.n3030 gnd 0.007621f
C4128 vdd.n3031 gnd 0.007621f
C4129 vdd.n3032 gnd 0.007621f
C4130 vdd.n3033 gnd 0.007621f
C4131 vdd.n3034 gnd 0.007621f
C4132 vdd.n3035 gnd 0.007621f
C4133 vdd.n3037 gnd 0.007621f
C4134 vdd.n3038 gnd 0.007621f
C4135 vdd.n3039 gnd 0.007621f
C4136 vdd.n3040 gnd 0.007621f
C4137 vdd.n3041 gnd 0.007621f
C4138 vdd.n3042 gnd 0.007621f
C4139 vdd.n3044 gnd 0.007621f
C4140 vdd.n3045 gnd 0.007621f
C4141 vdd.n3046 gnd 0.007621f
C4142 vdd.n3047 gnd 0.007621f
C4143 vdd.n3048 gnd 0.007621f
C4144 vdd.n3049 gnd 0.007621f
C4145 vdd.n3051 gnd 0.007621f
C4146 vdd.n3052 gnd 0.007621f
C4147 vdd.n3054 gnd 0.007621f
C4148 vdd.n3055 gnd 0.007621f
C4149 vdd.n3056 gnd 0.018084f
C4150 vdd.n3057 gnd 0.016885f
C4151 vdd.n3058 gnd 0.016885f
C4152 vdd.n3059 gnd 1.12249f
C4153 vdd.n3060 gnd 0.016885f
C4154 vdd.n3061 gnd 0.018084f
C4155 vdd.n3062 gnd 0.017156f
C4156 vdd.n3063 gnd 0.007621f
C4157 vdd.n3064 gnd 0.005884f
C4158 vdd.n3065 gnd 0.007621f
C4159 vdd.n3067 gnd 0.007621f
C4160 vdd.n3068 gnd 0.007621f
C4161 vdd.n3069 gnd 0.007621f
C4162 vdd.n3070 gnd 0.007621f
C4163 vdd.n3071 gnd 0.007621f
C4164 vdd.n3072 gnd 0.007621f
C4165 vdd.n3074 gnd 0.007621f
C4166 vdd.n3075 gnd 0.007621f
C4167 vdd.n3076 gnd 0.007621f
C4168 vdd.n3077 gnd 0.007621f
C4169 vdd.n3078 gnd 0.007621f
C4170 vdd.n3079 gnd 0.007621f
C4171 vdd.n3081 gnd 0.007621f
C4172 vdd.n3082 gnd 0.007621f
C4173 vdd.n3083 gnd 0.007621f
C4174 vdd.n3084 gnd 0.007621f
C4175 vdd.n3085 gnd 0.007621f
C4176 vdd.n3086 gnd 0.007621f
C4177 vdd.n3088 gnd 0.007621f
C4178 vdd.n3089 gnd 0.007621f
C4179 vdd.n3091 gnd 0.007621f
C4180 vdd.n3092 gnd 0.018314f
C4181 vdd.n3093 gnd 0.67832f
C4182 vdd.n3095 gnd 0.004736f
C4183 vdd.n3096 gnd 0.009021f
C4184 vdd.n3097 gnd 0.011208f
C4185 vdd.n3098 gnd 0.011208f
C4186 vdd.n3099 gnd 0.009021f
C4187 vdd.n3100 gnd 0.009021f
C4188 vdd.n3101 gnd 0.011208f
C4189 vdd.n3102 gnd 0.011208f
C4190 vdd.n3103 gnd 0.009021f
C4191 vdd.n3104 gnd 0.009021f
C4192 vdd.n3105 gnd 0.011208f
C4193 vdd.n3106 gnd 0.011208f
C4194 vdd.n3107 gnd 0.009021f
C4195 vdd.n3108 gnd 0.009021f
C4196 vdd.n3109 gnd 0.011208f
C4197 vdd.n3110 gnd 0.011208f
C4198 vdd.n3111 gnd 0.009021f
C4199 vdd.n3112 gnd 0.009021f
C4200 vdd.n3113 gnd 0.011208f
C4201 vdd.n3114 gnd 0.011208f
C4202 vdd.n3115 gnd 0.009021f
C4203 vdd.n3116 gnd 0.009021f
C4204 vdd.n3117 gnd 0.011208f
C4205 vdd.n3118 gnd 0.011208f
C4206 vdd.n3119 gnd 0.009021f
C4207 vdd.n3120 gnd 0.009021f
C4208 vdd.n3121 gnd 0.011208f
C4209 vdd.n3122 gnd 0.011208f
C4210 vdd.n3123 gnd 0.009021f
C4211 vdd.n3124 gnd 0.009021f
C4212 vdd.n3125 gnd 0.011208f
C4213 vdd.n3126 gnd 0.011208f
C4214 vdd.n3127 gnd 0.009021f
C4215 vdd.n3128 gnd 0.009021f
C4216 vdd.n3129 gnd 0.011208f
C4217 vdd.n3130 gnd 0.011208f
C4218 vdd.n3131 gnd 0.009021f
C4219 vdd.n3132 gnd 0.011208f
C4220 vdd.n3133 gnd 0.011208f
C4221 vdd.n3134 gnd 0.009021f
C4222 vdd.n3135 gnd 0.011208f
C4223 vdd.n3136 gnd 0.011208f
C4224 vdd.n3137 gnd 0.011208f
C4225 vdd.n3138 gnd 0.018403f
C4226 vdd.n3139 gnd 0.011208f
C4227 vdd.n3140 gnd 0.011208f
C4228 vdd.n3141 gnd 0.006134f
C4229 vdd.n3142 gnd 0.009021f
C4230 vdd.n3143 gnd 0.011208f
C4231 vdd.n3144 gnd 0.011208f
C4232 vdd.n3145 gnd 0.009021f
C4233 vdd.n3146 gnd 0.009021f
C4234 vdd.n3147 gnd 0.011208f
C4235 vdd.n3148 gnd 0.011208f
C4236 vdd.n3149 gnd 0.009021f
C4237 vdd.n3150 gnd 0.009021f
C4238 vdd.n3151 gnd 0.011208f
C4239 vdd.n3152 gnd 0.011208f
C4240 vdd.n3153 gnd 0.009021f
C4241 vdd.n3154 gnd 0.009021f
C4242 vdd.n3155 gnd 0.011208f
C4243 vdd.n3156 gnd 0.011208f
C4244 vdd.n3157 gnd 0.009021f
C4245 vdd.n3158 gnd 0.009021f
C4246 vdd.n3159 gnd 0.011208f
C4247 vdd.n3160 gnd 0.011208f
C4248 vdd.n3161 gnd 0.009021f
C4249 vdd.n3162 gnd 0.009021f
C4250 vdd.n3163 gnd 0.011208f
C4251 vdd.n3164 gnd 0.011208f
C4252 vdd.n3165 gnd 0.009021f
C4253 vdd.n3166 gnd 0.009021f
C4254 vdd.n3167 gnd 0.011208f
C4255 vdd.n3168 gnd 0.011208f
C4256 vdd.n3169 gnd 0.009021f
C4257 vdd.n3170 gnd 0.009021f
C4258 vdd.n3171 gnd 0.011208f
C4259 vdd.n3172 gnd 0.011208f
C4260 vdd.n3173 gnd 0.009021f
C4261 vdd.n3174 gnd 0.009021f
C4262 vdd.n3175 gnd 0.011208f
C4263 vdd.n3176 gnd 0.011208f
C4264 vdd.n3177 gnd 0.009021f
C4265 vdd.n3178 gnd 0.011208f
C4266 vdd.n3179 gnd 0.011208f
C4267 vdd.n3180 gnd 0.009021f
C4268 vdd.n3181 gnd 0.011208f
C4269 vdd.n3182 gnd 0.011208f
C4270 vdd.n3183 gnd 0.011208f
C4271 vdd.t39 gnd 0.137886f
C4272 vdd.t40 gnd 0.147363f
C4273 vdd.t38 gnd 0.180078f
C4274 vdd.n3184 gnd 0.230835f
C4275 vdd.n3185 gnd 0.193943f
C4276 vdd.n3186 gnd 0.018403f
C4277 vdd.n3187 gnd 0.011208f
C4278 vdd.n3188 gnd 0.011208f
C4279 vdd.n3189 gnd 0.007533f
C4280 vdd.n3190 gnd 0.009021f
C4281 vdd.n3191 gnd 0.011208f
C4282 vdd.n3192 gnd 0.011208f
C4283 vdd.n3193 gnd 0.009021f
C4284 vdd.n3194 gnd 0.009021f
C4285 vdd.n3195 gnd 0.011208f
C4286 vdd.n3196 gnd 0.011208f
C4287 vdd.n3197 gnd 0.009021f
C4288 vdd.n3198 gnd 0.009021f
C4289 vdd.n3199 gnd 0.011208f
C4290 vdd.n3200 gnd 0.011208f
C4291 vdd.n3201 gnd 0.009021f
C4292 vdd.n3202 gnd 0.009021f
C4293 vdd.n3203 gnd 0.011208f
C4294 vdd.n3204 gnd 0.011208f
C4295 vdd.n3205 gnd 0.009021f
C4296 vdd.n3206 gnd 0.009021f
C4297 vdd.n3207 gnd 0.011208f
C4298 vdd.n3208 gnd 0.011208f
C4299 vdd.n3209 gnd 0.009021f
C4300 vdd.n3210 gnd 0.009021f
C4301 vdd.n3211 gnd 0.011208f
C4302 vdd.n3212 gnd 0.011208f
C4303 vdd.n3213 gnd 0.009021f
C4304 vdd.n3214 gnd 0.009021f
C4305 vdd.n3216 gnd 0.67832f
C4306 vdd.n3218 gnd 0.009021f
C4307 vdd.n3219 gnd 0.009021f
C4308 vdd.n3220 gnd 0.007487f
C4309 vdd.n3221 gnd 0.027694f
C4310 vdd.n3223 gnd 8.281191f
C4311 vdd.n3224 gnd 0.027694f
C4312 vdd.n3225 gnd 0.004285f
C4313 vdd.n3226 gnd 0.027694f
C4314 vdd.n3227 gnd 0.027113f
C4315 vdd.n3228 gnd 0.011208f
C4316 vdd.n3229 gnd 0.009021f
C4317 vdd.n3230 gnd 0.011208f
C4318 vdd.n3231 gnd 0.692963f
C4319 vdd.n3232 gnd 0.011208f
C4320 vdd.n3233 gnd 0.009021f
C4321 vdd.n3234 gnd 0.011208f
C4322 vdd.n3235 gnd 0.011208f
C4323 vdd.n3236 gnd 0.011208f
C4324 vdd.n3237 gnd 0.009021f
C4325 vdd.n3238 gnd 0.011208f
C4326 vdd.n3239 gnd 1.14539f
C4327 vdd.n3240 gnd 0.011208f
C4328 vdd.n3241 gnd 0.009021f
C4329 vdd.n3242 gnd 0.011208f
C4330 vdd.n3243 gnd 0.011208f
C4331 vdd.n3244 gnd 0.011208f
C4332 vdd.n3245 gnd 0.009021f
C4333 vdd.n3246 gnd 0.011208f
C4334 vdd.n3247 gnd 0.738779f
C4335 vdd.n3248 gnd 0.784594f
C4336 vdd.n3249 gnd 0.011208f
C4337 vdd.n3250 gnd 0.009021f
C4338 vdd.n3251 gnd 0.011208f
C4339 vdd.n3252 gnd 0.011208f
C4340 vdd.n3253 gnd 0.011208f
C4341 vdd.n3254 gnd 0.009021f
C4342 vdd.n3255 gnd 0.011208f
C4343 vdd.n3256 gnd 0.950677f
C4344 vdd.n3257 gnd 0.011208f
C4345 vdd.n3258 gnd 0.009021f
C4346 vdd.n3259 gnd 0.011208f
C4347 vdd.n3260 gnd 0.011208f
C4348 vdd.n3261 gnd 0.011208f
C4349 vdd.n3262 gnd 0.009021f
C4350 vdd.n3263 gnd 0.011208f
C4351 vdd.t133 gnd 0.572697f
C4352 vdd.n3264 gnd 0.922042f
C4353 vdd.n3265 gnd 0.011208f
C4354 vdd.n3266 gnd 0.009021f
C4355 vdd.n3267 gnd 0.011208f
C4356 vdd.n3268 gnd 0.011208f
C4357 vdd.n3269 gnd 0.011208f
C4358 vdd.n3270 gnd 0.009021f
C4359 vdd.n3271 gnd 0.011208f
C4360 vdd.n3272 gnd 0.727325f
C4361 vdd.n3273 gnd 0.011208f
C4362 vdd.n3274 gnd 0.009021f
C4363 vdd.n3275 gnd 0.011208f
C4364 vdd.n3276 gnd 0.011208f
C4365 vdd.n3277 gnd 0.011208f
C4366 vdd.n3278 gnd 0.009021f
C4367 vdd.n3279 gnd 0.011208f
C4368 vdd.n3280 gnd 0.910588f
C4369 vdd.n3281 gnd 0.612785f
C4370 vdd.n3282 gnd 0.011208f
C4371 vdd.n3283 gnd 0.009021f
C4372 vdd.n3284 gnd 0.011208f
C4373 vdd.n3285 gnd 0.011208f
C4374 vdd.n3286 gnd 0.011208f
C4375 vdd.n3287 gnd 0.009021f
C4376 vdd.n3288 gnd 0.011208f
C4377 vdd.n3289 gnd 0.807502f
C4378 vdd.n3290 gnd 0.011208f
C4379 vdd.n3291 gnd 0.009021f
C4380 vdd.n3292 gnd 0.011208f
C4381 vdd.n3293 gnd 0.011208f
C4382 vdd.n3294 gnd 0.011208f
C4383 vdd.n3295 gnd 0.011208f
C4384 vdd.n3296 gnd 0.011208f
C4385 vdd.n3297 gnd 0.009021f
C4386 vdd.n3298 gnd 0.009021f
C4387 vdd.n3299 gnd 0.011208f
C4388 vdd.t183 gnd 0.572697f
C4389 vdd.n3300 gnd 0.950677f
C4390 vdd.n3301 gnd 0.011208f
C4391 vdd.n3302 gnd 0.009021f
C4392 vdd.n3303 gnd 0.011208f
C4393 vdd.n3304 gnd 0.011208f
C4394 vdd.n3305 gnd 0.011208f
C4395 vdd.n3306 gnd 0.009021f
C4396 vdd.n3307 gnd 0.011208f
C4397 vdd.n3308 gnd 0.899134f
C4398 vdd.n3309 gnd 0.011208f
C4399 vdd.n3310 gnd 0.011208f
C4400 vdd.n3311 gnd 0.009021f
C4401 vdd.n3312 gnd 0.009021f
C4402 vdd.n3313 gnd 0.011208f
C4403 vdd.n3314 gnd 0.011208f
C4404 vdd.n3315 gnd 0.011208f
C4405 vdd.n3316 gnd 0.009021f
C4406 vdd.n3317 gnd 0.011208f
C4407 vdd.n3318 gnd 0.009021f
C4408 vdd.n3319 gnd 0.009021f
C4409 vdd.n3320 gnd 0.011208f
C4410 vdd.n3321 gnd 0.011208f
C4411 vdd.n3322 gnd 0.011208f
C4412 vdd.n3323 gnd 0.009021f
C4413 vdd.n3324 gnd 0.011208f
C4414 vdd.n3325 gnd 0.009021f
C4415 vdd.n3326 gnd 0.009021f
C4416 vdd.n3327 gnd 0.011208f
C4417 vdd.n3328 gnd 0.011208f
C4418 vdd.n3329 gnd 0.011208f
C4419 vdd.n3330 gnd 0.009021f
C4420 vdd.n3331 gnd 0.950677f
C4421 vdd.n3332 gnd 0.011208f
C4422 vdd.n3333 gnd 0.009021f
C4423 vdd.n3334 gnd 0.009021f
C4424 vdd.n3335 gnd 0.011208f
C4425 vdd.n3336 gnd 0.011208f
C4426 vdd.n3337 gnd 0.011208f
C4427 vdd.n3338 gnd 0.009021f
C4428 vdd.n3339 gnd 0.011208f
C4429 vdd.n3340 gnd 0.009021f
C4430 vdd.n3341 gnd 0.009021f
C4431 vdd.n3342 gnd 0.011208f
C4432 vdd.n3343 gnd 0.011208f
C4433 vdd.n3344 gnd 0.011208f
C4434 vdd.n3345 gnd 0.009021f
C4435 vdd.n3346 gnd 0.011208f
C4436 vdd.n3347 gnd 0.009021f
C4437 vdd.n3348 gnd 0.007487f
C4438 vdd.n3349 gnd 0.027113f
C4439 vdd.n3350 gnd 0.027694f
C4440 vdd.n3351 gnd 0.004285f
C4441 vdd.n3352 gnd 0.027694f
C4442 vdd.n3354 gnd 2.71458f
C4443 vdd.n3355 gnd 1.68946f
C4444 vdd.n3356 gnd 0.027113f
C4445 vdd.n3357 gnd 0.007487f
C4446 vdd.n3358 gnd 0.009021f
C4447 vdd.n3359 gnd 0.009021f
C4448 vdd.n3360 gnd 0.011208f
C4449 vdd.n3361 gnd 1.14539f
C4450 vdd.n3362 gnd 1.14539f
C4451 vdd.n3363 gnd 1.04803f
C4452 vdd.n3364 gnd 0.011208f
C4453 vdd.n3365 gnd 0.009021f
C4454 vdd.n3366 gnd 0.009021f
C4455 vdd.n3367 gnd 0.009021f
C4456 vdd.n3368 gnd 0.011208f
C4457 vdd.n3369 gnd 0.853318f
C4458 vdd.t203 gnd 0.572697f
C4459 vdd.n3370 gnd 0.864772f
C4460 vdd.n3371 gnd 0.658601f
C4461 vdd.n3372 gnd 0.011208f
C4462 vdd.n3373 gnd 0.009021f
C4463 vdd.n3374 gnd 0.009021f
C4464 vdd.n3375 gnd 0.009021f
C4465 vdd.n3376 gnd 0.011208f
C4466 vdd.n3377 gnd 0.681509f
C4467 vdd.n3378 gnd 0.841864f
C4468 vdd.t151 gnd 0.572697f
C4469 vdd.n3379 gnd 0.876226f
C4470 vdd.n3380 gnd 0.011208f
C4471 vdd.n3381 gnd 0.009021f
C4472 vdd.n3382 gnd 0.009021f
C4473 vdd.n3383 gnd 0.009021f
C4474 vdd.n3384 gnd 0.011208f
C4475 vdd.n3385 gnd 0.950677f
C4476 vdd.t179 gnd 0.572697f
C4477 vdd.n3386 gnd 0.692963f
C4478 vdd.n3387 gnd 0.83041f
C4479 vdd.n3388 gnd 0.011208f
C4480 vdd.n3389 gnd 0.009021f
C4481 vdd.n3390 gnd 0.009021f
C4482 vdd.n3391 gnd 0.009021f
C4483 vdd.n3392 gnd 0.011208f
C4484 vdd.n3393 gnd 0.635693f
C4485 vdd.t147 gnd 0.572697f
C4486 vdd.n3394 gnd 0.950677f
C4487 vdd.t176 gnd 0.572697f
C4488 vdd.n3395 gnd 0.704417f
C4489 vdd.n3396 gnd 0.011208f
C4490 vdd.n3397 gnd 0.009021f
C4491 vdd.n3398 gnd 0.008614f
C4492 vdd.n3399 gnd 0.661084f
C4493 vdd.n3400 gnd 2.86602f
C4494 a_n7636_8799.n0 gnd 0.207851f
C4495 a_n7636_8799.n1 gnd 0.285406f
C4496 a_n7636_8799.n2 gnd 0.207851f
C4497 a_n7636_8799.n3 gnd 0.207851f
C4498 a_n7636_8799.n4 gnd 0.207851f
C4499 a_n7636_8799.n5 gnd 0.207851f
C4500 a_n7636_8799.n6 gnd 0.207851f
C4501 a_n7636_8799.n7 gnd 0.216127f
C4502 a_n7636_8799.n8 gnd 0.207851f
C4503 a_n7636_8799.n9 gnd 0.285406f
C4504 a_n7636_8799.n10 gnd 0.207851f
C4505 a_n7636_8799.n11 gnd 0.207851f
C4506 a_n7636_8799.n12 gnd 0.207851f
C4507 a_n7636_8799.n13 gnd 0.207851f
C4508 a_n7636_8799.n14 gnd 0.207851f
C4509 a_n7636_8799.n15 gnd 0.216127f
C4510 a_n7636_8799.n16 gnd 0.207851f
C4511 a_n7636_8799.n17 gnd 0.450503f
C4512 a_n7636_8799.n18 gnd 0.207851f
C4513 a_n7636_8799.n19 gnd 0.207851f
C4514 a_n7636_8799.n20 gnd 0.207851f
C4515 a_n7636_8799.n21 gnd 0.207851f
C4516 a_n7636_8799.n22 gnd 0.207851f
C4517 a_n7636_8799.n23 gnd 0.216127f
C4518 a_n7636_8799.n24 gnd 0.207851f
C4519 a_n7636_8799.n25 gnd 0.320053f
C4520 a_n7636_8799.n26 gnd 0.207851f
C4521 a_n7636_8799.n27 gnd 0.207851f
C4522 a_n7636_8799.n28 gnd 0.207851f
C4523 a_n7636_8799.n29 gnd 0.207851f
C4524 a_n7636_8799.n30 gnd 0.207851f
C4525 a_n7636_8799.n31 gnd 0.181481f
C4526 a_n7636_8799.n32 gnd 0.207851f
C4527 a_n7636_8799.n33 gnd 0.320053f
C4528 a_n7636_8799.n34 gnd 0.207851f
C4529 a_n7636_8799.n35 gnd 0.207851f
C4530 a_n7636_8799.n36 gnd 0.207851f
C4531 a_n7636_8799.n37 gnd 0.207851f
C4532 a_n7636_8799.n38 gnd 0.207851f
C4533 a_n7636_8799.n39 gnd 0.181481f
C4534 a_n7636_8799.n40 gnd 0.207851f
C4535 a_n7636_8799.n41 gnd 0.320053f
C4536 a_n7636_8799.n42 gnd 0.207851f
C4537 a_n7636_8799.n43 gnd 0.207851f
C4538 a_n7636_8799.n44 gnd 0.207851f
C4539 a_n7636_8799.n45 gnd 0.207851f
C4540 a_n7636_8799.n46 gnd 0.207851f
C4541 a_n7636_8799.n47 gnd 0.346578f
C4542 a_n7636_8799.n48 gnd 2.79182f
C4543 a_n7636_8799.n49 gnd 4.03031f
C4544 a_n7636_8799.n50 gnd 0.363344f
C4545 a_n7636_8799.n51 gnd 3.04515f
C4546 a_n7636_8799.n52 gnd 0.363343f
C4547 a_n7636_8799.n53 gnd 0.856369f
C4548 a_n7636_8799.n54 gnd 0.250233f
C4549 a_n7636_8799.n55 gnd 0.003658f
C4550 a_n7636_8799.n56 gnd 0.009643f
C4551 a_n7636_8799.n57 gnd 0.010536f
C4552 a_n7636_8799.n58 gnd 0.005567f
C4553 a_n7636_8799.n60 gnd 0.004672f
C4554 a_n7636_8799.n61 gnd 0.010104f
C4555 a_n7636_8799.n62 gnd 0.010104f
C4556 a_n7636_8799.n63 gnd 0.004672f
C4557 a_n7636_8799.n65 gnd 0.005567f
C4558 a_n7636_8799.n66 gnd 0.010536f
C4559 a_n7636_8799.n67 gnd 0.009643f
C4560 a_n7636_8799.n68 gnd 0.003658f
C4561 a_n7636_8799.n69 gnd 0.250233f
C4562 a_n7636_8799.n70 gnd 0.003658f
C4563 a_n7636_8799.n71 gnd 0.009643f
C4564 a_n7636_8799.n72 gnd 0.010536f
C4565 a_n7636_8799.n73 gnd 0.005567f
C4566 a_n7636_8799.n75 gnd 0.004672f
C4567 a_n7636_8799.n76 gnd 0.010104f
C4568 a_n7636_8799.n77 gnd 0.010104f
C4569 a_n7636_8799.n78 gnd 0.004672f
C4570 a_n7636_8799.n80 gnd 0.005567f
C4571 a_n7636_8799.n81 gnd 0.010536f
C4572 a_n7636_8799.n82 gnd 0.009643f
C4573 a_n7636_8799.n83 gnd 0.003658f
C4574 a_n7636_8799.n84 gnd 0.250233f
C4575 a_n7636_8799.n85 gnd 0.003658f
C4576 a_n7636_8799.n86 gnd 0.009643f
C4577 a_n7636_8799.n87 gnd 0.010536f
C4578 a_n7636_8799.n88 gnd 0.005567f
C4579 a_n7636_8799.n90 gnd 0.004672f
C4580 a_n7636_8799.n91 gnd 0.010104f
C4581 a_n7636_8799.n92 gnd 0.010104f
C4582 a_n7636_8799.n93 gnd 0.004672f
C4583 a_n7636_8799.n95 gnd 0.005567f
C4584 a_n7636_8799.n96 gnd 0.010536f
C4585 a_n7636_8799.n97 gnd 0.009643f
C4586 a_n7636_8799.n98 gnd 0.003658f
C4587 a_n7636_8799.n99 gnd 0.003658f
C4588 a_n7636_8799.n100 gnd 0.009643f
C4589 a_n7636_8799.n101 gnd 0.010536f
C4590 a_n7636_8799.n102 gnd 0.005567f
C4591 a_n7636_8799.n104 gnd 0.004672f
C4592 a_n7636_8799.n105 gnd 0.010104f
C4593 a_n7636_8799.n106 gnd 0.010104f
C4594 a_n7636_8799.n107 gnd 0.004672f
C4595 a_n7636_8799.n109 gnd 0.005567f
C4596 a_n7636_8799.n110 gnd 0.010536f
C4597 a_n7636_8799.n111 gnd 0.009643f
C4598 a_n7636_8799.n112 gnd 0.003658f
C4599 a_n7636_8799.n113 gnd 0.250233f
C4600 a_n7636_8799.n114 gnd 0.003658f
C4601 a_n7636_8799.n115 gnd 0.009643f
C4602 a_n7636_8799.n116 gnd 0.010536f
C4603 a_n7636_8799.n117 gnd 0.005567f
C4604 a_n7636_8799.n119 gnd 0.004672f
C4605 a_n7636_8799.n120 gnd 0.010104f
C4606 a_n7636_8799.n121 gnd 0.010104f
C4607 a_n7636_8799.n122 gnd 0.004672f
C4608 a_n7636_8799.n124 gnd 0.005567f
C4609 a_n7636_8799.n125 gnd 0.010536f
C4610 a_n7636_8799.n126 gnd 0.009643f
C4611 a_n7636_8799.n127 gnd 0.003658f
C4612 a_n7636_8799.n128 gnd 0.250233f
C4613 a_n7636_8799.n129 gnd 0.003658f
C4614 a_n7636_8799.n130 gnd 0.009643f
C4615 a_n7636_8799.n131 gnd 0.010536f
C4616 a_n7636_8799.n132 gnd 0.005567f
C4617 a_n7636_8799.n134 gnd 0.004672f
C4618 a_n7636_8799.n135 gnd 0.010104f
C4619 a_n7636_8799.n136 gnd 0.010104f
C4620 a_n7636_8799.n137 gnd 0.004672f
C4621 a_n7636_8799.n139 gnd 0.005567f
C4622 a_n7636_8799.n140 gnd 0.010536f
C4623 a_n7636_8799.n141 gnd 0.009643f
C4624 a_n7636_8799.n142 gnd 0.003658f
C4625 a_n7636_8799.n143 gnd 0.250233f
C4626 a_n7636_8799.t19 gnd 0.144168f
C4627 a_n7636_8799.t17 gnd 0.144168f
C4628 a_n7636_8799.t25 gnd 0.144168f
C4629 a_n7636_8799.n144 gnd 1.13707f
C4630 a_n7636_8799.t27 gnd 0.144168f
C4631 a_n7636_8799.t4 gnd 0.144168f
C4632 a_n7636_8799.n145 gnd 1.1352f
C4633 a_n7636_8799.t5 gnd 0.144168f
C4634 a_n7636_8799.t14 gnd 0.144168f
C4635 a_n7636_8799.n146 gnd 1.1352f
C4636 a_n7636_8799.t32 gnd 0.11213f
C4637 a_n7636_8799.t33 gnd 0.11213f
C4638 a_n7636_8799.n147 gnd 0.993745f
C4639 a_n7636_8799.t6 gnd 0.11213f
C4640 a_n7636_8799.t28 gnd 0.11213f
C4641 a_n7636_8799.n148 gnd 0.990823f
C4642 a_n7636_8799.n149 gnd 0.87861f
C4643 a_n7636_8799.t22 gnd 0.11213f
C4644 a_n7636_8799.t8 gnd 0.11213f
C4645 a_n7636_8799.n150 gnd 0.990823f
C4646 a_n7636_8799.t24 gnd 0.11213f
C4647 a_n7636_8799.t2 gnd 0.11213f
C4648 a_n7636_8799.n151 gnd 0.993744f
C4649 a_n7636_8799.t15 gnd 0.11213f
C4650 a_n7636_8799.t34 gnd 0.11213f
C4651 a_n7636_8799.n152 gnd 0.990822f
C4652 a_n7636_8799.n153 gnd 0.878612f
C4653 a_n7636_8799.t7 gnd 0.11213f
C4654 a_n7636_8799.t31 gnd 0.11213f
C4655 a_n7636_8799.n154 gnd 0.990822f
C4656 a_n7636_8799.t26 gnd 0.11213f
C4657 a_n7636_8799.t35 gnd 0.11213f
C4658 a_n7636_8799.n155 gnd 0.993744f
C4659 a_n7636_8799.t16 gnd 0.11213f
C4660 a_n7636_8799.t10 gnd 0.11213f
C4661 a_n7636_8799.n156 gnd 0.990822f
C4662 a_n7636_8799.n157 gnd 0.878612f
C4663 a_n7636_8799.t29 gnd 0.11213f
C4664 a_n7636_8799.t11 gnd 0.11213f
C4665 a_n7636_8799.n158 gnd 0.990822f
C4666 a_n7636_8799.t30 gnd 0.11213f
C4667 a_n7636_8799.t23 gnd 0.11213f
C4668 a_n7636_8799.n159 gnd 0.990823f
C4669 a_n7636_8799.n160 gnd 3.09086f
C4670 a_n7636_8799.t9 gnd 0.11213f
C4671 a_n7636_8799.t1 gnd 0.11213f
C4672 a_n7636_8799.n161 gnd 0.990823f
C4673 a_n7636_8799.n162 gnd 0.432601f
C4674 a_n7636_8799.t20 gnd 0.11213f
C4675 a_n7636_8799.t0 gnd 0.11213f
C4676 a_n7636_8799.n163 gnd 0.990823f
C4677 a_n7636_8799.t133 gnd 0.597786f
C4678 a_n7636_8799.n164 gnd 0.269131f
C4679 a_n7636_8799.t48 gnd 0.597786f
C4680 a_n7636_8799.t69 gnd 0.597786f
C4681 a_n7636_8799.n165 gnd 0.271059f
C4682 a_n7636_8799.t93 gnd 0.597786f
C4683 a_n7636_8799.t112 gnd 0.597786f
C4684 a_n7636_8799.n166 gnd 0.264259f
C4685 a_n7636_8799.t72 gnd 0.597786f
C4686 a_n7636_8799.t85 gnd 0.597786f
C4687 a_n7636_8799.n167 gnd 0.268238f
C4688 a_n7636_8799.t116 gnd 0.597786f
C4689 a_n7636_8799.t137 gnd 0.597786f
C4690 a_n7636_8799.t138 gnd 0.6091f
C4691 a_n7636_8799.n168 gnd 0.250596f
C4692 a_n7636_8799.n169 gnd 0.271432f
C4693 a_n7636_8799.t88 gnd 0.597786f
C4694 a_n7636_8799.n170 gnd 0.269131f
C4695 a_n7636_8799.n171 gnd 0.2649f
C4696 a_n7636_8799.t134 gnd 0.597786f
C4697 a_n7636_8799.n172 gnd 0.263619f
C4698 a_n7636_8799.t84 gnd 0.597786f
C4699 a_n7636_8799.n173 gnd 0.270804f
C4700 a_n7636_8799.t114 gnd 0.597786f
C4701 a_n7636_8799.n174 gnd 0.271059f
C4702 a_n7636_8799.n175 gnd 0.268671f
C4703 a_n7636_8799.t73 gnd 0.597786f
C4704 a_n7636_8799.n176 gnd 0.264259f
C4705 a_n7636_8799.t37 gnd 0.597786f
C4706 a_n7636_8799.n177 gnd 0.268671f
C4707 a_n7636_8799.n178 gnd 0.270804f
C4708 a_n7636_8799.t136 gnd 0.597786f
C4709 a_n7636_8799.n179 gnd 0.268238f
C4710 a_n7636_8799.n180 gnd 0.263619f
C4711 a_n7636_8799.t67 gnd 0.597786f
C4712 a_n7636_8799.n181 gnd 0.2649f
C4713 a_n7636_8799.t47 gnd 0.597786f
C4714 a_n7636_8799.n182 gnd 0.271432f
C4715 a_n7636_8799.t46 gnd 0.60909f
C4716 a_n7636_8799.t146 gnd 0.597786f
C4717 a_n7636_8799.n183 gnd 0.269131f
C4718 a_n7636_8799.t64 gnd 0.597786f
C4719 a_n7636_8799.t79 gnd 0.597786f
C4720 a_n7636_8799.n184 gnd 0.271059f
C4721 a_n7636_8799.t106 gnd 0.597786f
C4722 a_n7636_8799.t124 gnd 0.597786f
C4723 a_n7636_8799.n185 gnd 0.264259f
C4724 a_n7636_8799.t81 gnd 0.597786f
C4725 a_n7636_8799.t94 gnd 0.597786f
C4726 a_n7636_8799.n186 gnd 0.268238f
C4727 a_n7636_8799.t130 gnd 0.597786f
C4728 a_n7636_8799.t153 gnd 0.597786f
C4729 a_n7636_8799.t152 gnd 0.6091f
C4730 a_n7636_8799.n187 gnd 0.250596f
C4731 a_n7636_8799.n188 gnd 0.271432f
C4732 a_n7636_8799.t98 gnd 0.597786f
C4733 a_n7636_8799.n189 gnd 0.269131f
C4734 a_n7636_8799.n190 gnd 0.2649f
C4735 a_n7636_8799.t147 gnd 0.597786f
C4736 a_n7636_8799.n191 gnd 0.263619f
C4737 a_n7636_8799.t95 gnd 0.597786f
C4738 a_n7636_8799.n192 gnd 0.270804f
C4739 a_n7636_8799.t128 gnd 0.597786f
C4740 a_n7636_8799.n193 gnd 0.271059f
C4741 a_n7636_8799.n194 gnd 0.268671f
C4742 a_n7636_8799.t83 gnd 0.597786f
C4743 a_n7636_8799.n195 gnd 0.264259f
C4744 a_n7636_8799.t49 gnd 0.597786f
C4745 a_n7636_8799.n196 gnd 0.268671f
C4746 a_n7636_8799.n197 gnd 0.270804f
C4747 a_n7636_8799.t151 gnd 0.597786f
C4748 a_n7636_8799.n198 gnd 0.268238f
C4749 a_n7636_8799.n199 gnd 0.263619f
C4750 a_n7636_8799.t78 gnd 0.597786f
C4751 a_n7636_8799.n200 gnd 0.2649f
C4752 a_n7636_8799.t57 gnd 0.597786f
C4753 a_n7636_8799.n201 gnd 0.271432f
C4754 a_n7636_8799.t61 gnd 0.60909f
C4755 a_n7636_8799.n202 gnd 0.898688f
C4756 a_n7636_8799.t102 gnd 0.597786f
C4757 a_n7636_8799.n203 gnd 0.269131f
C4758 a_n7636_8799.t126 gnd 0.597786f
C4759 a_n7636_8799.t45 gnd 0.597786f
C4760 a_n7636_8799.n204 gnd 0.271059f
C4761 a_n7636_8799.t109 gnd 0.597786f
C4762 a_n7636_8799.t149 gnd 0.597786f
C4763 a_n7636_8799.n205 gnd 0.264259f
C4764 a_n7636_8799.t142 gnd 0.597786f
C4765 a_n7636_8799.t55 gnd 0.597786f
C4766 a_n7636_8799.n206 gnd 0.268238f
C4767 a_n7636_8799.t80 gnd 0.597786f
C4768 a_n7636_8799.t92 gnd 0.597786f
C4769 a_n7636_8799.t113 gnd 0.6091f
C4770 a_n7636_8799.n207 gnd 0.250596f
C4771 a_n7636_8799.n208 gnd 0.271432f
C4772 a_n7636_8799.t132 gnd 0.597786f
C4773 a_n7636_8799.n209 gnd 0.269131f
C4774 a_n7636_8799.n210 gnd 0.2649f
C4775 a_n7636_8799.t139 gnd 0.597786f
C4776 a_n7636_8799.n211 gnd 0.263619f
C4777 a_n7636_8799.t39 gnd 0.597786f
C4778 a_n7636_8799.n212 gnd 0.270804f
C4779 a_n7636_8799.t99 gnd 0.597786f
C4780 a_n7636_8799.n213 gnd 0.271059f
C4781 a_n7636_8799.n214 gnd 0.268671f
C4782 a_n7636_8799.t118 gnd 0.597786f
C4783 a_n7636_8799.n215 gnd 0.264259f
C4784 a_n7636_8799.t91 gnd 0.597786f
C4785 a_n7636_8799.n216 gnd 0.268671f
C4786 a_n7636_8799.n217 gnd 0.270804f
C4787 a_n7636_8799.t62 gnd 0.597786f
C4788 a_n7636_8799.n218 gnd 0.268238f
C4789 a_n7636_8799.n219 gnd 0.263619f
C4790 a_n7636_8799.t71 gnd 0.597786f
C4791 a_n7636_8799.n220 gnd 0.2649f
C4792 a_n7636_8799.t51 gnd 0.597786f
C4793 a_n7636_8799.n221 gnd 0.271432f
C4794 a_n7636_8799.t155 gnd 0.60909f
C4795 a_n7636_8799.n222 gnd 1.53919f
C4796 a_n7636_8799.t87 gnd 0.60909f
C4797 a_n7636_8799.t86 gnd 0.597786f
C4798 a_n7636_8799.t60 gnd 0.597786f
C4799 a_n7636_8799.n223 gnd 0.269131f
C4800 a_n7636_8799.t135 gnd 0.597786f
C4801 a_n7636_8799.t90 gnd 0.597786f
C4802 a_n7636_8799.t66 gnd 0.597786f
C4803 a_n7636_8799.n224 gnd 0.268238f
C4804 a_n7636_8799.t140 gnd 0.597786f
C4805 a_n7636_8799.t107 gnd 0.597786f
C4806 a_n7636_8799.t105 gnd 0.597786f
C4807 a_n7636_8799.n225 gnd 0.268671f
C4808 a_n7636_8799.t40 gnd 0.597786f
C4809 a_n7636_8799.t111 gnd 0.597786f
C4810 a_n7636_8799.t110 gnd 0.597786f
C4811 a_n7636_8799.n226 gnd 0.268671f
C4812 a_n7636_8799.t42 gnd 0.597786f
C4813 a_n7636_8799.t41 gnd 0.597786f
C4814 a_n7636_8799.t127 gnd 0.597786f
C4815 a_n7636_8799.n227 gnd 0.268238f
C4816 a_n7636_8799.t59 gnd 0.597786f
C4817 a_n7636_8799.t43 gnd 0.597786f
C4818 a_n7636_8799.t129 gnd 0.597786f
C4819 a_n7636_8799.n228 gnd 0.269131f
C4820 a_n7636_8799.t63 gnd 0.6091f
C4821 a_n7636_8799.n229 gnd 0.250596f
C4822 a_n7636_8799.t89 gnd 0.597786f
C4823 a_n7636_8799.n230 gnd 0.271432f
C4824 a_n7636_8799.n231 gnd 0.2649f
C4825 a_n7636_8799.n232 gnd 0.263619f
C4826 a_n7636_8799.n233 gnd 0.270804f
C4827 a_n7636_8799.n234 gnd 0.271059f
C4828 a_n7636_8799.n235 gnd 0.264259f
C4829 a_n7636_8799.n236 gnd 0.264259f
C4830 a_n7636_8799.n237 gnd 0.271059f
C4831 a_n7636_8799.n238 gnd 0.270804f
C4832 a_n7636_8799.n239 gnd 0.263619f
C4833 a_n7636_8799.n240 gnd 0.2649f
C4834 a_n7636_8799.n241 gnd 0.271432f
C4835 a_n7636_8799.t97 gnd 0.60909f
C4836 a_n7636_8799.t96 gnd 0.597786f
C4837 a_n7636_8799.t74 gnd 0.597786f
C4838 a_n7636_8799.n242 gnd 0.269131f
C4839 a_n7636_8799.t150 gnd 0.597786f
C4840 a_n7636_8799.t104 gnd 0.597786f
C4841 a_n7636_8799.t77 gnd 0.597786f
C4842 a_n7636_8799.n243 gnd 0.268238f
C4843 a_n7636_8799.t36 gnd 0.597786f
C4844 a_n7636_8799.t120 gnd 0.597786f
C4845 a_n7636_8799.t119 gnd 0.597786f
C4846 a_n7636_8799.n244 gnd 0.268671f
C4847 a_n7636_8799.t50 gnd 0.597786f
C4848 a_n7636_8799.t123 gnd 0.597786f
C4849 a_n7636_8799.t122 gnd 0.597786f
C4850 a_n7636_8799.n245 gnd 0.268671f
C4851 a_n7636_8799.t54 gnd 0.597786f
C4852 a_n7636_8799.t53 gnd 0.597786f
C4853 a_n7636_8799.t144 gnd 0.597786f
C4854 a_n7636_8799.n246 gnd 0.268238f
C4855 a_n7636_8799.t75 gnd 0.597786f
C4856 a_n7636_8799.t56 gnd 0.597786f
C4857 a_n7636_8799.t145 gnd 0.597786f
C4858 a_n7636_8799.n247 gnd 0.269131f
C4859 a_n7636_8799.t76 gnd 0.6091f
C4860 a_n7636_8799.n248 gnd 0.250596f
C4861 a_n7636_8799.t103 gnd 0.597786f
C4862 a_n7636_8799.n249 gnd 0.271432f
C4863 a_n7636_8799.n250 gnd 0.2649f
C4864 a_n7636_8799.n251 gnd 0.263619f
C4865 a_n7636_8799.n252 gnd 0.270804f
C4866 a_n7636_8799.n253 gnd 0.271059f
C4867 a_n7636_8799.n254 gnd 0.264259f
C4868 a_n7636_8799.n255 gnd 0.264259f
C4869 a_n7636_8799.n256 gnd 0.271059f
C4870 a_n7636_8799.n257 gnd 0.270804f
C4871 a_n7636_8799.n258 gnd 0.263619f
C4872 a_n7636_8799.n259 gnd 0.2649f
C4873 a_n7636_8799.n260 gnd 0.271432f
C4874 a_n7636_8799.n261 gnd 0.898688f
C4875 a_n7636_8799.t154 gnd 0.60909f
C4876 a_n7636_8799.t52 gnd 0.597786f
C4877 a_n7636_8799.t101 gnd 0.597786f
C4878 a_n7636_8799.n262 gnd 0.269131f
C4879 a_n7636_8799.t38 gnd 0.597786f
C4880 a_n7636_8799.t125 gnd 0.597786f
C4881 a_n7636_8799.t65 gnd 0.597786f
C4882 a_n7636_8799.n263 gnd 0.268238f
C4883 a_n7636_8799.t108 gnd 0.597786f
C4884 a_n7636_8799.t44 gnd 0.597786f
C4885 a_n7636_8799.t70 gnd 0.597786f
C4886 a_n7636_8799.n264 gnd 0.268671f
C4887 a_n7636_8799.t148 gnd 0.597786f
C4888 a_n7636_8799.t117 gnd 0.597786f
C4889 a_n7636_8799.t143 gnd 0.597786f
C4890 a_n7636_8799.n265 gnd 0.268671f
C4891 a_n7636_8799.t100 gnd 0.597786f
C4892 a_n7636_8799.t121 gnd 0.597786f
C4893 a_n7636_8799.t58 gnd 0.597786f
C4894 a_n7636_8799.n266 gnd 0.268238f
C4895 a_n7636_8799.t141 gnd 0.597786f
C4896 a_n7636_8799.t82 gnd 0.597786f
C4897 a_n7636_8799.t131 gnd 0.597786f
C4898 a_n7636_8799.n267 gnd 0.269131f
C4899 a_n7636_8799.t115 gnd 0.6091f
C4900 a_n7636_8799.n268 gnd 0.250596f
C4901 a_n7636_8799.t68 gnd 0.597786f
C4902 a_n7636_8799.n269 gnd 0.271432f
C4903 a_n7636_8799.n270 gnd 0.2649f
C4904 a_n7636_8799.n271 gnd 0.263619f
C4905 a_n7636_8799.n272 gnd 0.270804f
C4906 a_n7636_8799.n273 gnd 0.271059f
C4907 a_n7636_8799.n274 gnd 0.264259f
C4908 a_n7636_8799.n275 gnd 0.264259f
C4909 a_n7636_8799.n276 gnd 0.271059f
C4910 a_n7636_8799.n277 gnd 0.270804f
C4911 a_n7636_8799.n278 gnd 0.263619f
C4912 a_n7636_8799.n279 gnd 0.2649f
C4913 a_n7636_8799.n280 gnd 0.271432f
C4914 a_n7636_8799.n281 gnd 1.08607f
C4915 a_n7636_8799.n282 gnd 12.209499f
C4916 a_n7636_8799.n283 gnd 4.37493f
C4917 a_n7636_8799.n284 gnd 5.67621f
C4918 a_n7636_8799.t12 gnd 0.144168f
C4919 a_n7636_8799.t13 gnd 0.144168f
C4920 a_n7636_8799.n285 gnd 1.1352f
C4921 a_n7636_8799.t18 gnd 0.144168f
C4922 a_n7636_8799.t21 gnd 0.144168f
C4923 a_n7636_8799.n286 gnd 1.1352f
C4924 a_n7636_8799.n287 gnd 1.13708f
C4925 a_n7636_8799.t3 gnd 0.144168f
C4926 CSoutput.n0 gnd 0.048568f
C4927 CSoutput.t178 gnd 0.321267f
C4928 CSoutput.n1 gnd 0.145068f
C4929 CSoutput.n2 gnd 0.048568f
C4930 CSoutput.t183 gnd 0.321267f
C4931 CSoutput.n3 gnd 0.038494f
C4932 CSoutput.n4 gnd 0.048568f
C4933 CSoutput.t172 gnd 0.321267f
C4934 CSoutput.n5 gnd 0.033194f
C4935 CSoutput.n6 gnd 0.048568f
C4936 CSoutput.t180 gnd 0.321267f
C4937 CSoutput.t186 gnd 0.321267f
C4938 CSoutput.n7 gnd 0.143487f
C4939 CSoutput.n8 gnd 0.048568f
C4940 CSoutput.t185 gnd 0.321267f
C4941 CSoutput.n9 gnd 0.031648f
C4942 CSoutput.n10 gnd 0.048568f
C4943 CSoutput.t173 gnd 0.321267f
C4944 CSoutput.t184 gnd 0.321267f
C4945 CSoutput.n11 gnd 0.143487f
C4946 CSoutput.n12 gnd 0.048568f
C4947 CSoutput.t182 gnd 0.321267f
C4948 CSoutput.n13 gnd 0.033194f
C4949 CSoutput.n14 gnd 0.048568f
C4950 CSoutput.t171 gnd 0.321267f
C4951 CSoutput.t175 gnd 0.321267f
C4952 CSoutput.n15 gnd 0.143487f
C4953 CSoutput.n16 gnd 0.048568f
C4954 CSoutput.t179 gnd 0.321267f
C4955 CSoutput.n17 gnd 0.035452f
C4956 CSoutput.t189 gnd 0.383922f
C4957 CSoutput.t169 gnd 0.321267f
C4958 CSoutput.n18 gnd 0.183177f
C4959 CSoutput.n19 gnd 0.177745f
C4960 CSoutput.n20 gnd 0.206206f
C4961 CSoutput.n21 gnd 0.048568f
C4962 CSoutput.n22 gnd 0.040535f
C4963 CSoutput.n23 gnd 0.143487f
C4964 CSoutput.n24 gnd 0.039075f
C4965 CSoutput.n25 gnd 0.038494f
C4966 CSoutput.n26 gnd 0.048568f
C4967 CSoutput.n27 gnd 0.048568f
C4968 CSoutput.n28 gnd 0.040224f
C4969 CSoutput.n29 gnd 0.034151f
C4970 CSoutput.n30 gnd 0.146681f
C4971 CSoutput.n31 gnd 0.034621f
C4972 CSoutput.n32 gnd 0.048568f
C4973 CSoutput.n33 gnd 0.048568f
C4974 CSoutput.n34 gnd 0.048568f
C4975 CSoutput.n35 gnd 0.039795f
C4976 CSoutput.n36 gnd 0.143487f
C4977 CSoutput.n37 gnd 0.038058f
C4978 CSoutput.n38 gnd 0.03951f
C4979 CSoutput.n39 gnd 0.048568f
C4980 CSoutput.n40 gnd 0.048568f
C4981 CSoutput.n41 gnd 0.040527f
C4982 CSoutput.n42 gnd 0.037042f
C4983 CSoutput.n43 gnd 0.143487f
C4984 CSoutput.n44 gnd 0.037981f
C4985 CSoutput.n45 gnd 0.048568f
C4986 CSoutput.n46 gnd 0.048568f
C4987 CSoutput.n47 gnd 0.048568f
C4988 CSoutput.n48 gnd 0.037981f
C4989 CSoutput.n49 gnd 0.143487f
C4990 CSoutput.n50 gnd 0.037042f
C4991 CSoutput.n51 gnd 0.040527f
C4992 CSoutput.n52 gnd 0.048568f
C4993 CSoutput.n53 gnd 0.048568f
C4994 CSoutput.n54 gnd 0.03951f
C4995 CSoutput.n55 gnd 0.038058f
C4996 CSoutput.n56 gnd 0.143487f
C4997 CSoutput.n57 gnd 0.039795f
C4998 CSoutput.n58 gnd 0.048568f
C4999 CSoutput.n59 gnd 0.048568f
C5000 CSoutput.n60 gnd 0.048568f
C5001 CSoutput.n61 gnd 0.034621f
C5002 CSoutput.n62 gnd 0.146681f
C5003 CSoutput.n63 gnd 0.034151f
C5004 CSoutput.t188 gnd 0.321267f
C5005 CSoutput.n64 gnd 0.143487f
C5006 CSoutput.n65 gnd 0.040224f
C5007 CSoutput.n66 gnd 0.048568f
C5008 CSoutput.n67 gnd 0.048568f
C5009 CSoutput.n68 gnd 0.048568f
C5010 CSoutput.n69 gnd 0.039075f
C5011 CSoutput.n70 gnd 0.143487f
C5012 CSoutput.n71 gnd 0.040535f
C5013 CSoutput.n72 gnd 0.035452f
C5014 CSoutput.n73 gnd 0.048568f
C5015 CSoutput.n74 gnd 0.048568f
C5016 CSoutput.n75 gnd 0.036767f
C5017 CSoutput.n76 gnd 0.021836f
C5018 CSoutput.t168 gnd 0.360966f
C5019 CSoutput.n77 gnd 0.179313f
C5020 CSoutput.n78 gnd 0.767266f
C5021 CSoutput.t71 gnd 0.060582f
C5022 CSoutput.t98 gnd 0.060582f
C5023 CSoutput.n79 gnd 0.469044f
C5024 CSoutput.t161 gnd 0.060582f
C5025 CSoutput.t158 gnd 0.060582f
C5026 CSoutput.n80 gnd 0.468208f
C5027 CSoutput.n81 gnd 0.47523f
C5028 CSoutput.t0 gnd 0.060582f
C5029 CSoutput.t2 gnd 0.060582f
C5030 CSoutput.n82 gnd 0.468208f
C5031 CSoutput.n83 gnd 0.234173f
C5032 CSoutput.t132 gnd 0.060582f
C5033 CSoutput.t80 gnd 0.060582f
C5034 CSoutput.n84 gnd 0.468208f
C5035 CSoutput.n85 gnd 0.234173f
C5036 CSoutput.t127 gnd 0.060582f
C5037 CSoutput.t133 gnd 0.060582f
C5038 CSoutput.n86 gnd 0.468208f
C5039 CSoutput.n87 gnd 0.234173f
C5040 CSoutput.t156 gnd 0.060582f
C5041 CSoutput.t112 gnd 0.060582f
C5042 CSoutput.n88 gnd 0.468208f
C5043 CSoutput.n89 gnd 0.234173f
C5044 CSoutput.t82 gnd 0.060582f
C5045 CSoutput.t143 gnd 0.060582f
C5046 CSoutput.n90 gnd 0.468208f
C5047 CSoutput.n91 gnd 0.234173f
C5048 CSoutput.t114 gnd 0.060582f
C5049 CSoutput.t107 gnd 0.060582f
C5050 CSoutput.n92 gnd 0.468208f
C5051 CSoutput.n93 gnd 0.234173f
C5052 CSoutput.t124 gnd 0.060582f
C5053 CSoutput.t4 gnd 0.060582f
C5054 CSoutput.n94 gnd 0.468208f
C5055 CSoutput.n95 gnd 0.234173f
C5056 CSoutput.t79 gnd 0.060582f
C5057 CSoutput.t121 gnd 0.060582f
C5058 CSoutput.n96 gnd 0.468208f
C5059 CSoutput.n97 gnd 0.42942f
C5060 CSoutput.t87 gnd 0.060582f
C5061 CSoutput.t92 gnd 0.060582f
C5062 CSoutput.n98 gnd 0.469044f
C5063 CSoutput.t134 gnd 0.060582f
C5064 CSoutput.t9 gnd 0.060582f
C5065 CSoutput.n99 gnd 0.468208f
C5066 CSoutput.n100 gnd 0.47523f
C5067 CSoutput.t88 gnd 0.060582f
C5068 CSoutput.t115 gnd 0.060582f
C5069 CSoutput.n101 gnd 0.468208f
C5070 CSoutput.n102 gnd 0.234173f
C5071 CSoutput.t10 gnd 0.060582f
C5072 CSoutput.t147 gnd 0.060582f
C5073 CSoutput.n103 gnd 0.468208f
C5074 CSoutput.n104 gnd 0.234173f
C5075 CSoutput.t67 gnd 0.060582f
C5076 CSoutput.t141 gnd 0.060582f
C5077 CSoutput.n105 gnd 0.468208f
C5078 CSoutput.n106 gnd 0.234173f
C5079 CSoutput.t61 gnd 0.060582f
C5080 CSoutput.t59 gnd 0.060582f
C5081 CSoutput.n107 gnd 0.468208f
C5082 CSoutput.n108 gnd 0.234173f
C5083 CSoutput.t146 gnd 0.060582f
C5084 CSoutput.t78 gnd 0.060582f
C5085 CSoutput.n109 gnd 0.468208f
C5086 CSoutput.n110 gnd 0.234173f
C5087 CSoutput.t157 gnd 0.060582f
C5088 CSoutput.t148 gnd 0.060582f
C5089 CSoutput.n111 gnd 0.468208f
C5090 CSoutput.n112 gnd 0.234173f
C5091 CSoutput.t70 gnd 0.060582f
C5092 CSoutput.t105 gnd 0.060582f
C5093 CSoutput.n113 gnd 0.468208f
C5094 CSoutput.n114 gnd 0.234173f
C5095 CSoutput.t166 gnd 0.060582f
C5096 CSoutput.t125 gnd 0.060582f
C5097 CSoutput.n115 gnd 0.468208f
C5098 CSoutput.n116 gnd 0.349211f
C5099 CSoutput.n117 gnd 0.440353f
C5100 CSoutput.t102 gnd 0.060582f
C5101 CSoutput.t151 gnd 0.060582f
C5102 CSoutput.n118 gnd 0.469044f
C5103 CSoutput.t137 gnd 0.060582f
C5104 CSoutput.t84 gnd 0.060582f
C5105 CSoutput.n119 gnd 0.468208f
C5106 CSoutput.n120 gnd 0.47523f
C5107 CSoutput.t139 gnd 0.060582f
C5108 CSoutput.t68 gnd 0.060582f
C5109 CSoutput.n121 gnd 0.468208f
C5110 CSoutput.n122 gnd 0.234173f
C5111 CSoutput.t6 gnd 0.060582f
C5112 CSoutput.t1 gnd 0.060582f
C5113 CSoutput.n123 gnd 0.468208f
C5114 CSoutput.n124 gnd 0.234173f
C5115 CSoutput.t144 gnd 0.060582f
C5116 CSoutput.t83 gnd 0.060582f
C5117 CSoutput.n125 gnd 0.468208f
C5118 CSoutput.n126 gnd 0.234173f
C5119 CSoutput.t138 gnd 0.060582f
C5120 CSoutput.t129 gnd 0.060582f
C5121 CSoutput.n127 gnd 0.468208f
C5122 CSoutput.n128 gnd 0.234173f
C5123 CSoutput.t119 gnd 0.060582f
C5124 CSoutput.t63 gnd 0.060582f
C5125 CSoutput.n129 gnd 0.468208f
C5126 CSoutput.n130 gnd 0.234173f
C5127 CSoutput.t76 gnd 0.060582f
C5128 CSoutput.t81 gnd 0.060582f
C5129 CSoutput.n131 gnd 0.468208f
C5130 CSoutput.n132 gnd 0.234173f
C5131 CSoutput.t118 gnd 0.060582f
C5132 CSoutput.t122 gnd 0.060582f
C5133 CSoutput.n133 gnd 0.468208f
C5134 CSoutput.n134 gnd 0.234173f
C5135 CSoutput.t159 gnd 0.060582f
C5136 CSoutput.t85 gnd 0.060582f
C5137 CSoutput.n135 gnd 0.468208f
C5138 CSoutput.n136 gnd 0.349211f
C5139 CSoutput.n137 gnd 0.492202f
C5140 CSoutput.n138 gnd 8.46936f
C5141 CSoutput.n140 gnd 0.859159f
C5142 CSoutput.n141 gnd 0.644369f
C5143 CSoutput.n142 gnd 0.859159f
C5144 CSoutput.n143 gnd 0.859159f
C5145 CSoutput.n144 gnd 2.31312f
C5146 CSoutput.n145 gnd 0.859159f
C5147 CSoutput.n146 gnd 0.859159f
C5148 CSoutput.t187 gnd 1.07395f
C5149 CSoutput.n147 gnd 0.859159f
C5150 CSoutput.n148 gnd 0.859159f
C5151 CSoutput.n152 gnd 0.859159f
C5152 CSoutput.n156 gnd 0.859159f
C5153 CSoutput.n157 gnd 0.859159f
C5154 CSoutput.n159 gnd 0.859159f
C5155 CSoutput.n164 gnd 0.859159f
C5156 CSoutput.n166 gnd 0.859159f
C5157 CSoutput.n167 gnd 0.859159f
C5158 CSoutput.n169 gnd 0.859159f
C5159 CSoutput.n170 gnd 0.859159f
C5160 CSoutput.n172 gnd 0.859159f
C5161 CSoutput.t176 gnd 14.356501f
C5162 CSoutput.n174 gnd 0.859159f
C5163 CSoutput.n175 gnd 0.644369f
C5164 CSoutput.n176 gnd 0.859159f
C5165 CSoutput.n177 gnd 0.859159f
C5166 CSoutput.n178 gnd 2.31312f
C5167 CSoutput.n179 gnd 0.859159f
C5168 CSoutput.n180 gnd 0.859159f
C5169 CSoutput.t174 gnd 1.07395f
C5170 CSoutput.n181 gnd 0.859159f
C5171 CSoutput.n182 gnd 0.859159f
C5172 CSoutput.n186 gnd 0.859159f
C5173 CSoutput.n190 gnd 0.859159f
C5174 CSoutput.n191 gnd 0.859159f
C5175 CSoutput.n193 gnd 0.859159f
C5176 CSoutput.n198 gnd 0.859159f
C5177 CSoutput.n200 gnd 0.859159f
C5178 CSoutput.n201 gnd 0.859159f
C5179 CSoutput.n203 gnd 0.859159f
C5180 CSoutput.n204 gnd 0.859159f
C5181 CSoutput.n206 gnd 0.859159f
C5182 CSoutput.n207 gnd 0.644369f
C5183 CSoutput.n209 gnd 0.859159f
C5184 CSoutput.n210 gnd 0.644369f
C5185 CSoutput.n211 gnd 0.859159f
C5186 CSoutput.n212 gnd 0.859159f
C5187 CSoutput.n213 gnd 2.31312f
C5188 CSoutput.n214 gnd 0.859159f
C5189 CSoutput.n215 gnd 0.859159f
C5190 CSoutput.t170 gnd 1.07395f
C5191 CSoutput.n216 gnd 0.859159f
C5192 CSoutput.n217 gnd 2.31312f
C5193 CSoutput.n219 gnd 0.859159f
C5194 CSoutput.n220 gnd 0.859159f
C5195 CSoutput.n222 gnd 0.859159f
C5196 CSoutput.n223 gnd 0.859159f
C5197 CSoutput.t177 gnd 14.122499f
C5198 CSoutput.t181 gnd 14.356501f
C5199 CSoutput.n229 gnd 2.69531f
C5200 CSoutput.n230 gnd 10.9797f
C5201 CSoutput.n231 gnd 11.439099f
C5202 CSoutput.n236 gnd 2.91974f
C5203 CSoutput.n242 gnd 0.859159f
C5204 CSoutput.n244 gnd 0.859159f
C5205 CSoutput.n246 gnd 0.859159f
C5206 CSoutput.n248 gnd 0.859159f
C5207 CSoutput.n250 gnd 0.859159f
C5208 CSoutput.n256 gnd 0.859159f
C5209 CSoutput.n263 gnd 1.57623f
C5210 CSoutput.n264 gnd 1.57623f
C5211 CSoutput.n265 gnd 0.859159f
C5212 CSoutput.n266 gnd 0.859159f
C5213 CSoutput.n268 gnd 0.644369f
C5214 CSoutput.n269 gnd 0.551844f
C5215 CSoutput.n271 gnd 0.644369f
C5216 CSoutput.n272 gnd 0.551844f
C5217 CSoutput.n273 gnd 0.644369f
C5218 CSoutput.n275 gnd 0.859159f
C5219 CSoutput.n277 gnd 2.31312f
C5220 CSoutput.n278 gnd 2.69531f
C5221 CSoutput.n279 gnd 10.098499f
C5222 CSoutput.n281 gnd 0.644369f
C5223 CSoutput.n282 gnd 1.658f
C5224 CSoutput.n283 gnd 0.644369f
C5225 CSoutput.n285 gnd 0.859159f
C5226 CSoutput.n287 gnd 2.31312f
C5227 CSoutput.n288 gnd 5.03835f
C5228 CSoutput.t104 gnd 0.060582f
C5229 CSoutput.t152 gnd 0.060582f
C5230 CSoutput.n289 gnd 0.469044f
C5231 CSoutput.t69 gnd 0.060582f
C5232 CSoutput.t65 gnd 0.060582f
C5233 CSoutput.n290 gnd 0.468208f
C5234 CSoutput.n291 gnd 0.47523f
C5235 CSoutput.t96 gnd 0.060582f
C5236 CSoutput.t135 gnd 0.060582f
C5237 CSoutput.n292 gnd 0.468208f
C5238 CSoutput.n293 gnd 0.234173f
C5239 CSoutput.t66 gnd 0.060582f
C5240 CSoutput.t145 gnd 0.060582f
C5241 CSoutput.n294 gnd 0.468208f
C5242 CSoutput.n295 gnd 0.234173f
C5243 CSoutput.t7 gnd 0.060582f
C5244 CSoutput.t72 gnd 0.060582f
C5245 CSoutput.n296 gnd 0.468208f
C5246 CSoutput.n297 gnd 0.234173f
C5247 CSoutput.t167 gnd 0.060582f
C5248 CSoutput.t93 gnd 0.060582f
C5249 CSoutput.n298 gnd 0.468208f
C5250 CSoutput.n299 gnd 0.234173f
C5251 CSoutput.t100 gnd 0.060582f
C5252 CSoutput.t86 gnd 0.060582f
C5253 CSoutput.n300 gnd 0.468208f
C5254 CSoutput.n301 gnd 0.234173f
C5255 CSoutput.t97 gnd 0.060582f
C5256 CSoutput.t90 gnd 0.060582f
C5257 CSoutput.n302 gnd 0.468208f
C5258 CSoutput.n303 gnd 0.234173f
C5259 CSoutput.t106 gnd 0.060582f
C5260 CSoutput.t160 gnd 0.060582f
C5261 CSoutput.n304 gnd 0.468208f
C5262 CSoutput.n305 gnd 0.234173f
C5263 CSoutput.t123 gnd 0.060582f
C5264 CSoutput.t165 gnd 0.060582f
C5265 CSoutput.n306 gnd 0.468208f
C5266 CSoutput.n307 gnd 0.42942f
C5267 CSoutput.t149 gnd 0.060582f
C5268 CSoutput.t62 gnd 0.060582f
C5269 CSoutput.n308 gnd 0.469044f
C5270 CSoutput.t126 gnd 0.060582f
C5271 CSoutput.t8 gnd 0.060582f
C5272 CSoutput.n309 gnd 0.468208f
C5273 CSoutput.n310 gnd 0.47523f
C5274 CSoutput.t64 gnd 0.060582f
C5275 CSoutput.t128 gnd 0.060582f
C5276 CSoutput.n311 gnd 0.468208f
C5277 CSoutput.n312 gnd 0.234173f
C5278 CSoutput.t111 gnd 0.060582f
C5279 CSoutput.t113 gnd 0.060582f
C5280 CSoutput.n313 gnd 0.468208f
C5281 CSoutput.n314 gnd 0.234173f
C5282 CSoutput.t95 gnd 0.060582f
C5283 CSoutput.t60 gnd 0.060582f
C5284 CSoutput.n315 gnd 0.468208f
C5285 CSoutput.n316 gnd 0.234173f
C5286 CSoutput.t94 gnd 0.060582f
C5287 CSoutput.t77 gnd 0.060582f
C5288 CSoutput.n317 gnd 0.468208f
C5289 CSoutput.n318 gnd 0.234173f
C5290 CSoutput.t150 gnd 0.060582f
C5291 CSoutput.t89 gnd 0.060582f
C5292 CSoutput.n319 gnd 0.468208f
C5293 CSoutput.n320 gnd 0.234173f
C5294 CSoutput.t74 gnd 0.060582f
C5295 CSoutput.t73 gnd 0.060582f
C5296 CSoutput.n321 gnd 0.468208f
C5297 CSoutput.n322 gnd 0.234173f
C5298 CSoutput.t101 gnd 0.060582f
C5299 CSoutput.t164 gnd 0.060582f
C5300 CSoutput.n323 gnd 0.468208f
C5301 CSoutput.n324 gnd 0.234173f
C5302 CSoutput.t155 gnd 0.060582f
C5303 CSoutput.t103 gnd 0.060582f
C5304 CSoutput.n325 gnd 0.468208f
C5305 CSoutput.n326 gnd 0.349211f
C5306 CSoutput.n327 gnd 0.440353f
C5307 CSoutput.t5 gnd 0.060582f
C5308 CSoutput.t109 gnd 0.060582f
C5309 CSoutput.n328 gnd 0.469044f
C5310 CSoutput.t162 gnd 0.060582f
C5311 CSoutput.t91 gnd 0.060582f
C5312 CSoutput.n329 gnd 0.468208f
C5313 CSoutput.n330 gnd 0.47523f
C5314 CSoutput.t117 gnd 0.060582f
C5315 CSoutput.t136 gnd 0.060582f
C5316 CSoutput.n331 gnd 0.468208f
C5317 CSoutput.n332 gnd 0.234173f
C5318 CSoutput.t75 gnd 0.060582f
C5319 CSoutput.t142 gnd 0.060582f
C5320 CSoutput.n333 gnd 0.468208f
C5321 CSoutput.n334 gnd 0.234173f
C5322 CSoutput.t108 gnd 0.060582f
C5323 CSoutput.t154 gnd 0.060582f
C5324 CSoutput.n335 gnd 0.468208f
C5325 CSoutput.n336 gnd 0.234173f
C5326 CSoutput.t140 gnd 0.060582f
C5327 CSoutput.t153 gnd 0.060582f
C5328 CSoutput.n337 gnd 0.468208f
C5329 CSoutput.n338 gnd 0.234173f
C5330 CSoutput.t110 gnd 0.060582f
C5331 CSoutput.t120 gnd 0.060582f
C5332 CSoutput.n339 gnd 0.468208f
C5333 CSoutput.n340 gnd 0.234173f
C5334 CSoutput.t99 gnd 0.060582f
C5335 CSoutput.t163 gnd 0.060582f
C5336 CSoutput.n341 gnd 0.468208f
C5337 CSoutput.n342 gnd 0.234173f
C5338 CSoutput.t130 gnd 0.060582f
C5339 CSoutput.t3 gnd 0.060582f
C5340 CSoutput.n343 gnd 0.468208f
C5341 CSoutput.n344 gnd 0.234173f
C5342 CSoutput.t116 gnd 0.060582f
C5343 CSoutput.t131 gnd 0.060582f
C5344 CSoutput.n345 gnd 0.468206f
C5345 CSoutput.n346 gnd 0.349213f
C5346 CSoutput.n347 gnd 0.492202f
C5347 CSoutput.n348 gnd 12.4079f
C5348 CSoutput.t35 gnd 0.053009f
C5349 CSoutput.t25 gnd 0.053009f
C5350 CSoutput.n349 gnd 0.469974f
C5351 CSoutput.t51 gnd 0.053009f
C5352 CSoutput.t53 gnd 0.053009f
C5353 CSoutput.n350 gnd 0.468406f
C5354 CSoutput.n351 gnd 0.436467f
C5355 CSoutput.t30 gnd 0.053009f
C5356 CSoutput.t20 gnd 0.053009f
C5357 CSoutput.n352 gnd 0.468406f
C5358 CSoutput.n353 gnd 0.215158f
C5359 CSoutput.t56 gnd 0.053009f
C5360 CSoutput.t37 gnd 0.053009f
C5361 CSoutput.n354 gnd 0.468406f
C5362 CSoutput.n355 gnd 0.215158f
C5363 CSoutput.t39 gnd 0.053009f
C5364 CSoutput.t28 gnd 0.053009f
C5365 CSoutput.n356 gnd 0.468406f
C5366 CSoutput.n357 gnd 0.215158f
C5367 CSoutput.t42 gnd 0.053009f
C5368 CSoutput.t44 gnd 0.053009f
C5369 CSoutput.n358 gnd 0.468406f
C5370 CSoutput.n359 gnd 0.396794f
C5371 CSoutput.t45 gnd 0.053009f
C5372 CSoutput.t34 gnd 0.053009f
C5373 CSoutput.n360 gnd 0.469974f
C5374 CSoutput.t57 gnd 0.053009f
C5375 CSoutput.t11 gnd 0.053009f
C5376 CSoutput.n361 gnd 0.468406f
C5377 CSoutput.n362 gnd 0.436467f
C5378 CSoutput.t40 gnd 0.053009f
C5379 CSoutput.t29 gnd 0.053009f
C5380 CSoutput.n363 gnd 0.468406f
C5381 CSoutput.n364 gnd 0.215158f
C5382 CSoutput.t15 gnd 0.053009f
C5383 CSoutput.t46 gnd 0.053009f
C5384 CSoutput.n365 gnd 0.468406f
C5385 CSoutput.n366 gnd 0.215158f
C5386 CSoutput.t48 gnd 0.053009f
C5387 CSoutput.t38 gnd 0.053009f
C5388 CSoutput.n367 gnd 0.468406f
C5389 CSoutput.n368 gnd 0.215158f
C5390 CSoutput.t49 gnd 0.053009f
C5391 CSoutput.t52 gnd 0.053009f
C5392 CSoutput.n369 gnd 0.468406f
C5393 CSoutput.n370 gnd 0.326656f
C5394 CSoutput.n371 gnd 0.606951f
C5395 CSoutput.n372 gnd 12.5767f
C5396 CSoutput.t14 gnd 0.053009f
C5397 CSoutput.t22 gnd 0.053009f
C5398 CSoutput.n373 gnd 0.469974f
C5399 CSoutput.t43 gnd 0.053009f
C5400 CSoutput.t55 gnd 0.053009f
C5401 CSoutput.n374 gnd 0.468406f
C5402 CSoutput.n375 gnd 0.436467f
C5403 CSoutput.t58 gnd 0.053009f
C5404 CSoutput.t18 gnd 0.053009f
C5405 CSoutput.n376 gnd 0.468406f
C5406 CSoutput.n377 gnd 0.215158f
C5407 CSoutput.t23 gnd 0.053009f
C5408 CSoutput.t12 gnd 0.053009f
C5409 CSoutput.n378 gnd 0.468406f
C5410 CSoutput.n379 gnd 0.215158f
C5411 CSoutput.t16 gnd 0.053009f
C5412 CSoutput.t26 gnd 0.053009f
C5413 CSoutput.n380 gnd 0.468406f
C5414 CSoutput.n381 gnd 0.215158f
C5415 CSoutput.t31 gnd 0.053009f
C5416 CSoutput.t47 gnd 0.053009f
C5417 CSoutput.n382 gnd 0.468406f
C5418 CSoutput.n383 gnd 0.396794f
C5419 CSoutput.t21 gnd 0.053009f
C5420 CSoutput.t33 gnd 0.053009f
C5421 CSoutput.n384 gnd 0.469974f
C5422 CSoutput.t50 gnd 0.053009f
C5423 CSoutput.t13 gnd 0.053009f
C5424 CSoutput.n385 gnd 0.468406f
C5425 CSoutput.n386 gnd 0.436467f
C5426 CSoutput.t17 gnd 0.053009f
C5427 CSoutput.t27 gnd 0.053009f
C5428 CSoutput.n387 gnd 0.468406f
C5429 CSoutput.n388 gnd 0.215158f
C5430 CSoutput.t32 gnd 0.053009f
C5431 CSoutput.t19 gnd 0.053009f
C5432 CSoutput.n389 gnd 0.468406f
C5433 CSoutput.n390 gnd 0.215158f
C5434 CSoutput.t24 gnd 0.053009f
C5435 CSoutput.t36 gnd 0.053009f
C5436 CSoutput.n391 gnd 0.468406f
C5437 CSoutput.n392 gnd 0.215158f
C5438 CSoutput.t41 gnd 0.053009f
C5439 CSoutput.t54 gnd 0.053009f
C5440 CSoutput.n393 gnd 0.468406f
C5441 CSoutput.n394 gnd 0.326656f
C5442 CSoutput.n395 gnd 0.606951f
C5443 CSoutput.n396 gnd 7.06881f
C5444 CSoutput.n397 gnd 15.512099f
C5445 commonsourceibias.n0 gnd 0.010301f
C5446 commonsourceibias.t71 gnd 0.155981f
C5447 commonsourceibias.t81 gnd 0.144227f
C5448 commonsourceibias.n1 gnd 0.057546f
C5449 commonsourceibias.n2 gnd 0.00772f
C5450 commonsourceibias.t55 gnd 0.144227f
C5451 commonsourceibias.n3 gnd 0.006245f
C5452 commonsourceibias.n4 gnd 0.00772f
C5453 commonsourceibias.t53 gnd 0.144227f
C5454 commonsourceibias.n5 gnd 0.007453f
C5455 commonsourceibias.n6 gnd 0.00772f
C5456 commonsourceibias.t76 gnd 0.144227f
C5457 commonsourceibias.n7 gnd 0.057546f
C5458 commonsourceibias.t86 gnd 0.144227f
C5459 commonsourceibias.n8 gnd 0.006235f
C5460 commonsourceibias.n9 gnd 0.010301f
C5461 commonsourceibias.t32 gnd 0.155981f
C5462 commonsourceibias.t14 gnd 0.144227f
C5463 commonsourceibias.n10 gnd 0.057546f
C5464 commonsourceibias.n11 gnd 0.00772f
C5465 commonsourceibias.t24 gnd 0.144227f
C5466 commonsourceibias.n12 gnd 0.006245f
C5467 commonsourceibias.n13 gnd 0.00772f
C5468 commonsourceibias.t30 gnd 0.144227f
C5469 commonsourceibias.n14 gnd 0.007453f
C5470 commonsourceibias.n15 gnd 0.00772f
C5471 commonsourceibias.t20 gnd 0.144227f
C5472 commonsourceibias.n16 gnd 0.057546f
C5473 commonsourceibias.t36 gnd 0.144227f
C5474 commonsourceibias.n17 gnd 0.006235f
C5475 commonsourceibias.n18 gnd 0.00772f
C5476 commonsourceibias.t44 gnd 0.144227f
C5477 commonsourceibias.t26 gnd 0.144227f
C5478 commonsourceibias.n19 gnd 0.057546f
C5479 commonsourceibias.n20 gnd 0.00772f
C5480 commonsourceibias.t34 gnd 0.144227f
C5481 commonsourceibias.n21 gnd 0.057546f
C5482 commonsourceibias.n22 gnd 0.00772f
C5483 commonsourceibias.t10 gnd 0.144227f
C5484 commonsourceibias.n23 gnd 0.057546f
C5485 commonsourceibias.n24 gnd 0.038863f
C5486 commonsourceibias.t40 gnd 0.144227f
C5487 commonsourceibias.t46 gnd 0.162743f
C5488 commonsourceibias.n25 gnd 0.066782f
C5489 commonsourceibias.n26 gnd 0.069137f
C5490 commonsourceibias.n27 gnd 0.009515f
C5491 commonsourceibias.n28 gnd 0.010526f
C5492 commonsourceibias.n29 gnd 0.00772f
C5493 commonsourceibias.n30 gnd 0.00772f
C5494 commonsourceibias.n31 gnd 0.010457f
C5495 commonsourceibias.n32 gnd 0.006245f
C5496 commonsourceibias.n33 gnd 0.010587f
C5497 commonsourceibias.n34 gnd 0.00772f
C5498 commonsourceibias.n35 gnd 0.00772f
C5499 commonsourceibias.n36 gnd 0.010651f
C5500 commonsourceibias.n37 gnd 0.009185f
C5501 commonsourceibias.n38 gnd 0.007453f
C5502 commonsourceibias.n39 gnd 0.00772f
C5503 commonsourceibias.n40 gnd 0.00772f
C5504 commonsourceibias.n41 gnd 0.009442f
C5505 commonsourceibias.n42 gnd 0.010598f
C5506 commonsourceibias.n43 gnd 0.057546f
C5507 commonsourceibias.n44 gnd 0.010527f
C5508 commonsourceibias.n45 gnd 0.00772f
C5509 commonsourceibias.n46 gnd 0.00772f
C5510 commonsourceibias.n47 gnd 0.00772f
C5511 commonsourceibias.n48 gnd 0.010527f
C5512 commonsourceibias.n49 gnd 0.057546f
C5513 commonsourceibias.n50 gnd 0.010598f
C5514 commonsourceibias.n51 gnd 0.009442f
C5515 commonsourceibias.n52 gnd 0.00772f
C5516 commonsourceibias.n53 gnd 0.00772f
C5517 commonsourceibias.n54 gnd 0.00772f
C5518 commonsourceibias.n55 gnd 0.009185f
C5519 commonsourceibias.n56 gnd 0.010651f
C5520 commonsourceibias.n57 gnd 0.057546f
C5521 commonsourceibias.n58 gnd 0.010587f
C5522 commonsourceibias.n59 gnd 0.00772f
C5523 commonsourceibias.n60 gnd 0.00772f
C5524 commonsourceibias.n61 gnd 0.00772f
C5525 commonsourceibias.n62 gnd 0.010457f
C5526 commonsourceibias.n63 gnd 0.057546f
C5527 commonsourceibias.n64 gnd 0.010526f
C5528 commonsourceibias.n65 gnd 0.009515f
C5529 commonsourceibias.n66 gnd 0.00772f
C5530 commonsourceibias.n67 gnd 0.00772f
C5531 commonsourceibias.n68 gnd 0.007831f
C5532 commonsourceibias.n69 gnd 0.008096f
C5533 commonsourceibias.n70 gnd 0.068855f
C5534 commonsourceibias.n71 gnd 0.076384f
C5535 commonsourceibias.t33 gnd 0.016658f
C5536 commonsourceibias.t15 gnd 0.016658f
C5537 commonsourceibias.n72 gnd 0.147197f
C5538 commonsourceibias.n73 gnd 0.12719f
C5539 commonsourceibias.t25 gnd 0.016658f
C5540 commonsourceibias.t31 gnd 0.016658f
C5541 commonsourceibias.n74 gnd 0.147197f
C5542 commonsourceibias.n75 gnd 0.067614f
C5543 commonsourceibias.t21 gnd 0.016658f
C5544 commonsourceibias.t37 gnd 0.016658f
C5545 commonsourceibias.n76 gnd 0.147197f
C5546 commonsourceibias.n77 gnd 0.056488f
C5547 commonsourceibias.t41 gnd 0.016658f
C5548 commonsourceibias.t47 gnd 0.016658f
C5549 commonsourceibias.n78 gnd 0.14769f
C5550 commonsourceibias.t35 gnd 0.016658f
C5551 commonsourceibias.t11 gnd 0.016658f
C5552 commonsourceibias.n79 gnd 0.147197f
C5553 commonsourceibias.n80 gnd 0.13716f
C5554 commonsourceibias.t45 gnd 0.016658f
C5555 commonsourceibias.t27 gnd 0.016658f
C5556 commonsourceibias.n81 gnd 0.147197f
C5557 commonsourceibias.n82 gnd 0.056488f
C5558 commonsourceibias.n83 gnd 0.068401f
C5559 commonsourceibias.n84 gnd 0.00772f
C5560 commonsourceibias.t50 gnd 0.144227f
C5561 commonsourceibias.t69 gnd 0.144227f
C5562 commonsourceibias.n85 gnd 0.057546f
C5563 commonsourceibias.n86 gnd 0.00772f
C5564 commonsourceibias.t67 gnd 0.144227f
C5565 commonsourceibias.n87 gnd 0.057546f
C5566 commonsourceibias.n88 gnd 0.00772f
C5567 commonsourceibias.t78 gnd 0.144227f
C5568 commonsourceibias.n89 gnd 0.057546f
C5569 commonsourceibias.n90 gnd 0.038863f
C5570 commonsourceibias.t64 gnd 0.144227f
C5571 commonsourceibias.t62 gnd 0.162743f
C5572 commonsourceibias.n91 gnd 0.066782f
C5573 commonsourceibias.n92 gnd 0.069137f
C5574 commonsourceibias.n93 gnd 0.009515f
C5575 commonsourceibias.n94 gnd 0.010526f
C5576 commonsourceibias.n95 gnd 0.00772f
C5577 commonsourceibias.n96 gnd 0.00772f
C5578 commonsourceibias.n97 gnd 0.010457f
C5579 commonsourceibias.n98 gnd 0.006245f
C5580 commonsourceibias.n99 gnd 0.010587f
C5581 commonsourceibias.n100 gnd 0.00772f
C5582 commonsourceibias.n101 gnd 0.00772f
C5583 commonsourceibias.n102 gnd 0.010651f
C5584 commonsourceibias.n103 gnd 0.009185f
C5585 commonsourceibias.n104 gnd 0.007453f
C5586 commonsourceibias.n105 gnd 0.00772f
C5587 commonsourceibias.n106 gnd 0.00772f
C5588 commonsourceibias.n107 gnd 0.009442f
C5589 commonsourceibias.n108 gnd 0.010598f
C5590 commonsourceibias.n109 gnd 0.057546f
C5591 commonsourceibias.n110 gnd 0.010527f
C5592 commonsourceibias.n111 gnd 0.007683f
C5593 commonsourceibias.n112 gnd 0.055804f
C5594 commonsourceibias.n113 gnd 0.007683f
C5595 commonsourceibias.n114 gnd 0.010527f
C5596 commonsourceibias.n115 gnd 0.057546f
C5597 commonsourceibias.n116 gnd 0.010598f
C5598 commonsourceibias.n117 gnd 0.009442f
C5599 commonsourceibias.n118 gnd 0.00772f
C5600 commonsourceibias.n119 gnd 0.00772f
C5601 commonsourceibias.n120 gnd 0.00772f
C5602 commonsourceibias.n121 gnd 0.009185f
C5603 commonsourceibias.n122 gnd 0.010651f
C5604 commonsourceibias.n123 gnd 0.057546f
C5605 commonsourceibias.n124 gnd 0.010587f
C5606 commonsourceibias.n125 gnd 0.00772f
C5607 commonsourceibias.n126 gnd 0.00772f
C5608 commonsourceibias.n127 gnd 0.00772f
C5609 commonsourceibias.n128 gnd 0.010457f
C5610 commonsourceibias.n129 gnd 0.057546f
C5611 commonsourceibias.n130 gnd 0.010526f
C5612 commonsourceibias.n131 gnd 0.009515f
C5613 commonsourceibias.n132 gnd 0.00772f
C5614 commonsourceibias.n133 gnd 0.00772f
C5615 commonsourceibias.n134 gnd 0.007831f
C5616 commonsourceibias.n135 gnd 0.008096f
C5617 commonsourceibias.n136 gnd 0.068855f
C5618 commonsourceibias.n137 gnd 0.04456f
C5619 commonsourceibias.n138 gnd 0.010301f
C5620 commonsourceibias.t72 gnd 0.144227f
C5621 commonsourceibias.n139 gnd 0.057546f
C5622 commonsourceibias.n140 gnd 0.00772f
C5623 commonsourceibias.t49 gnd 0.144227f
C5624 commonsourceibias.n141 gnd 0.006245f
C5625 commonsourceibias.n142 gnd 0.00772f
C5626 commonsourceibias.t95 gnd 0.144227f
C5627 commonsourceibias.n143 gnd 0.007453f
C5628 commonsourceibias.n144 gnd 0.00772f
C5629 commonsourceibias.t66 gnd 0.144227f
C5630 commonsourceibias.n145 gnd 0.057546f
C5631 commonsourceibias.t77 gnd 0.144227f
C5632 commonsourceibias.n146 gnd 0.006235f
C5633 commonsourceibias.n147 gnd 0.00772f
C5634 commonsourceibias.t91 gnd 0.144227f
C5635 commonsourceibias.t60 gnd 0.144227f
C5636 commonsourceibias.n148 gnd 0.057546f
C5637 commonsourceibias.n149 gnd 0.00772f
C5638 commonsourceibias.t58 gnd 0.144227f
C5639 commonsourceibias.n150 gnd 0.057546f
C5640 commonsourceibias.n151 gnd 0.00772f
C5641 commonsourceibias.t68 gnd 0.144227f
C5642 commonsourceibias.n152 gnd 0.057546f
C5643 commonsourceibias.n153 gnd 0.038863f
C5644 commonsourceibias.t57 gnd 0.144227f
C5645 commonsourceibias.t54 gnd 0.162743f
C5646 commonsourceibias.n154 gnd 0.066782f
C5647 commonsourceibias.n155 gnd 0.069137f
C5648 commonsourceibias.n156 gnd 0.009515f
C5649 commonsourceibias.n157 gnd 0.010526f
C5650 commonsourceibias.n158 gnd 0.00772f
C5651 commonsourceibias.n159 gnd 0.00772f
C5652 commonsourceibias.n160 gnd 0.010457f
C5653 commonsourceibias.n161 gnd 0.006245f
C5654 commonsourceibias.n162 gnd 0.010587f
C5655 commonsourceibias.n163 gnd 0.00772f
C5656 commonsourceibias.n164 gnd 0.00772f
C5657 commonsourceibias.n165 gnd 0.010651f
C5658 commonsourceibias.n166 gnd 0.009185f
C5659 commonsourceibias.n167 gnd 0.007453f
C5660 commonsourceibias.n168 gnd 0.00772f
C5661 commonsourceibias.n169 gnd 0.00772f
C5662 commonsourceibias.n170 gnd 0.009442f
C5663 commonsourceibias.n171 gnd 0.010598f
C5664 commonsourceibias.n172 gnd 0.057546f
C5665 commonsourceibias.n173 gnd 0.010527f
C5666 commonsourceibias.n174 gnd 0.00772f
C5667 commonsourceibias.n175 gnd 0.00772f
C5668 commonsourceibias.n176 gnd 0.00772f
C5669 commonsourceibias.n177 gnd 0.010527f
C5670 commonsourceibias.n178 gnd 0.057546f
C5671 commonsourceibias.n179 gnd 0.010598f
C5672 commonsourceibias.n180 gnd 0.009442f
C5673 commonsourceibias.n181 gnd 0.00772f
C5674 commonsourceibias.n182 gnd 0.00772f
C5675 commonsourceibias.n183 gnd 0.00772f
C5676 commonsourceibias.n184 gnd 0.009185f
C5677 commonsourceibias.n185 gnd 0.010651f
C5678 commonsourceibias.n186 gnd 0.057546f
C5679 commonsourceibias.n187 gnd 0.010587f
C5680 commonsourceibias.n188 gnd 0.00772f
C5681 commonsourceibias.n189 gnd 0.00772f
C5682 commonsourceibias.n190 gnd 0.00772f
C5683 commonsourceibias.n191 gnd 0.010457f
C5684 commonsourceibias.n192 gnd 0.057546f
C5685 commonsourceibias.n193 gnd 0.010526f
C5686 commonsourceibias.n194 gnd 0.009515f
C5687 commonsourceibias.n195 gnd 0.00772f
C5688 commonsourceibias.n196 gnd 0.00772f
C5689 commonsourceibias.n197 gnd 0.007831f
C5690 commonsourceibias.n198 gnd 0.008096f
C5691 commonsourceibias.t61 gnd 0.155981f
C5692 commonsourceibias.n199 gnd 0.068855f
C5693 commonsourceibias.n200 gnd 0.023432f
C5694 commonsourceibias.n201 gnd 0.388694f
C5695 commonsourceibias.n202 gnd 0.010301f
C5696 commonsourceibias.t84 gnd 0.155981f
C5697 commonsourceibias.t92 gnd 0.144227f
C5698 commonsourceibias.n203 gnd 0.057546f
C5699 commonsourceibias.n204 gnd 0.00772f
C5700 commonsourceibias.t51 gnd 0.144227f
C5701 commonsourceibias.n205 gnd 0.006245f
C5702 commonsourceibias.n206 gnd 0.00772f
C5703 commonsourceibias.t63 gnd 0.144227f
C5704 commonsourceibias.n207 gnd 0.007453f
C5705 commonsourceibias.n208 gnd 0.00772f
C5706 commonsourceibias.t48 gnd 0.144227f
C5707 commonsourceibias.n209 gnd 0.006235f
C5708 commonsourceibias.n210 gnd 0.00772f
C5709 commonsourceibias.t94 gnd 0.144227f
C5710 commonsourceibias.t83 gnd 0.144227f
C5711 commonsourceibias.n211 gnd 0.057546f
C5712 commonsourceibias.n212 gnd 0.00772f
C5713 commonsourceibias.t80 gnd 0.144227f
C5714 commonsourceibias.n213 gnd 0.057546f
C5715 commonsourceibias.n214 gnd 0.00772f
C5716 commonsourceibias.t90 gnd 0.144227f
C5717 commonsourceibias.n215 gnd 0.057546f
C5718 commonsourceibias.n216 gnd 0.038863f
C5719 commonsourceibias.t59 gnd 0.144227f
C5720 commonsourceibias.t75 gnd 0.162743f
C5721 commonsourceibias.n217 gnd 0.066782f
C5722 commonsourceibias.n218 gnd 0.069137f
C5723 commonsourceibias.n219 gnd 0.009515f
C5724 commonsourceibias.n220 gnd 0.010526f
C5725 commonsourceibias.n221 gnd 0.00772f
C5726 commonsourceibias.n222 gnd 0.00772f
C5727 commonsourceibias.n223 gnd 0.010457f
C5728 commonsourceibias.n224 gnd 0.006245f
C5729 commonsourceibias.n225 gnd 0.010587f
C5730 commonsourceibias.n226 gnd 0.00772f
C5731 commonsourceibias.n227 gnd 0.00772f
C5732 commonsourceibias.n228 gnd 0.010651f
C5733 commonsourceibias.n229 gnd 0.009185f
C5734 commonsourceibias.n230 gnd 0.007453f
C5735 commonsourceibias.n231 gnd 0.00772f
C5736 commonsourceibias.n232 gnd 0.00772f
C5737 commonsourceibias.n233 gnd 0.009442f
C5738 commonsourceibias.n234 gnd 0.010598f
C5739 commonsourceibias.n235 gnd 0.057546f
C5740 commonsourceibias.n236 gnd 0.010527f
C5741 commonsourceibias.n237 gnd 0.007683f
C5742 commonsourceibias.t17 gnd 0.016658f
C5743 commonsourceibias.t9 gnd 0.016658f
C5744 commonsourceibias.n238 gnd 0.14769f
C5745 commonsourceibias.t19 gnd 0.016658f
C5746 commonsourceibias.t5 gnd 0.016658f
C5747 commonsourceibias.n239 gnd 0.147197f
C5748 commonsourceibias.n240 gnd 0.13716f
C5749 commonsourceibias.t43 gnd 0.016658f
C5750 commonsourceibias.t13 gnd 0.016658f
C5751 commonsourceibias.n241 gnd 0.147197f
C5752 commonsourceibias.n242 gnd 0.056488f
C5753 commonsourceibias.n243 gnd 0.010301f
C5754 commonsourceibias.t22 gnd 0.144227f
C5755 commonsourceibias.n244 gnd 0.057546f
C5756 commonsourceibias.n245 gnd 0.00772f
C5757 commonsourceibias.t38 gnd 0.144227f
C5758 commonsourceibias.n246 gnd 0.006245f
C5759 commonsourceibias.n247 gnd 0.00772f
C5760 commonsourceibias.t0 gnd 0.144227f
C5761 commonsourceibias.n248 gnd 0.007453f
C5762 commonsourceibias.n249 gnd 0.00772f
C5763 commonsourceibias.t6 gnd 0.144227f
C5764 commonsourceibias.n250 gnd 0.006235f
C5765 commonsourceibias.n251 gnd 0.00772f
C5766 commonsourceibias.t12 gnd 0.144227f
C5767 commonsourceibias.t42 gnd 0.144227f
C5768 commonsourceibias.n252 gnd 0.057546f
C5769 commonsourceibias.n253 gnd 0.00772f
C5770 commonsourceibias.t4 gnd 0.144227f
C5771 commonsourceibias.n254 gnd 0.057546f
C5772 commonsourceibias.n255 gnd 0.00772f
C5773 commonsourceibias.t18 gnd 0.144227f
C5774 commonsourceibias.n256 gnd 0.057546f
C5775 commonsourceibias.n257 gnd 0.038863f
C5776 commonsourceibias.t8 gnd 0.144227f
C5777 commonsourceibias.t16 gnd 0.162743f
C5778 commonsourceibias.n258 gnd 0.066782f
C5779 commonsourceibias.n259 gnd 0.069137f
C5780 commonsourceibias.n260 gnd 0.009515f
C5781 commonsourceibias.n261 gnd 0.010526f
C5782 commonsourceibias.n262 gnd 0.00772f
C5783 commonsourceibias.n263 gnd 0.00772f
C5784 commonsourceibias.n264 gnd 0.010457f
C5785 commonsourceibias.n265 gnd 0.006245f
C5786 commonsourceibias.n266 gnd 0.010587f
C5787 commonsourceibias.n267 gnd 0.00772f
C5788 commonsourceibias.n268 gnd 0.00772f
C5789 commonsourceibias.n269 gnd 0.010651f
C5790 commonsourceibias.n270 gnd 0.009185f
C5791 commonsourceibias.n271 gnd 0.007453f
C5792 commonsourceibias.n272 gnd 0.00772f
C5793 commonsourceibias.n273 gnd 0.00772f
C5794 commonsourceibias.n274 gnd 0.009442f
C5795 commonsourceibias.n275 gnd 0.010598f
C5796 commonsourceibias.n276 gnd 0.057546f
C5797 commonsourceibias.n277 gnd 0.010527f
C5798 commonsourceibias.n278 gnd 0.00772f
C5799 commonsourceibias.n279 gnd 0.00772f
C5800 commonsourceibias.n280 gnd 0.00772f
C5801 commonsourceibias.n281 gnd 0.010527f
C5802 commonsourceibias.n282 gnd 0.057546f
C5803 commonsourceibias.n283 gnd 0.010598f
C5804 commonsourceibias.t28 gnd 0.144227f
C5805 commonsourceibias.n284 gnd 0.057546f
C5806 commonsourceibias.n285 gnd 0.009442f
C5807 commonsourceibias.n286 gnd 0.00772f
C5808 commonsourceibias.n287 gnd 0.00772f
C5809 commonsourceibias.n288 gnd 0.00772f
C5810 commonsourceibias.n289 gnd 0.009185f
C5811 commonsourceibias.n290 gnd 0.010651f
C5812 commonsourceibias.n291 gnd 0.057546f
C5813 commonsourceibias.n292 gnd 0.010587f
C5814 commonsourceibias.n293 gnd 0.00772f
C5815 commonsourceibias.n294 gnd 0.00772f
C5816 commonsourceibias.n295 gnd 0.00772f
C5817 commonsourceibias.n296 gnd 0.010457f
C5818 commonsourceibias.n297 gnd 0.057546f
C5819 commonsourceibias.n298 gnd 0.010526f
C5820 commonsourceibias.n299 gnd 0.009515f
C5821 commonsourceibias.n300 gnd 0.00772f
C5822 commonsourceibias.n301 gnd 0.00772f
C5823 commonsourceibias.n302 gnd 0.007831f
C5824 commonsourceibias.n303 gnd 0.008096f
C5825 commonsourceibias.t2 gnd 0.155981f
C5826 commonsourceibias.n304 gnd 0.068855f
C5827 commonsourceibias.n305 gnd 0.076384f
C5828 commonsourceibias.t23 gnd 0.016658f
C5829 commonsourceibias.t3 gnd 0.016658f
C5830 commonsourceibias.n306 gnd 0.147197f
C5831 commonsourceibias.n307 gnd 0.12719f
C5832 commonsourceibias.t1 gnd 0.016658f
C5833 commonsourceibias.t39 gnd 0.016658f
C5834 commonsourceibias.n308 gnd 0.147197f
C5835 commonsourceibias.n309 gnd 0.067614f
C5836 commonsourceibias.t7 gnd 0.016658f
C5837 commonsourceibias.t29 gnd 0.016658f
C5838 commonsourceibias.n310 gnd 0.147197f
C5839 commonsourceibias.n311 gnd 0.056488f
C5840 commonsourceibias.n312 gnd 0.068401f
C5841 commonsourceibias.n313 gnd 0.055804f
C5842 commonsourceibias.n314 gnd 0.007683f
C5843 commonsourceibias.n315 gnd 0.010527f
C5844 commonsourceibias.n316 gnd 0.057546f
C5845 commonsourceibias.n317 gnd 0.010598f
C5846 commonsourceibias.t88 gnd 0.144227f
C5847 commonsourceibias.n318 gnd 0.057546f
C5848 commonsourceibias.n319 gnd 0.009442f
C5849 commonsourceibias.n320 gnd 0.00772f
C5850 commonsourceibias.n321 gnd 0.00772f
C5851 commonsourceibias.n322 gnd 0.00772f
C5852 commonsourceibias.n323 gnd 0.009185f
C5853 commonsourceibias.n324 gnd 0.010651f
C5854 commonsourceibias.n325 gnd 0.057546f
C5855 commonsourceibias.n326 gnd 0.010587f
C5856 commonsourceibias.n327 gnd 0.00772f
C5857 commonsourceibias.n328 gnd 0.00772f
C5858 commonsourceibias.n329 gnd 0.00772f
C5859 commonsourceibias.n330 gnd 0.010457f
C5860 commonsourceibias.n331 gnd 0.057546f
C5861 commonsourceibias.n332 gnd 0.010526f
C5862 commonsourceibias.n333 gnd 0.009515f
C5863 commonsourceibias.n334 gnd 0.00772f
C5864 commonsourceibias.n335 gnd 0.00772f
C5865 commonsourceibias.n336 gnd 0.007831f
C5866 commonsourceibias.n337 gnd 0.008096f
C5867 commonsourceibias.n338 gnd 0.068855f
C5868 commonsourceibias.n339 gnd 0.04456f
C5869 commonsourceibias.n340 gnd 0.010301f
C5870 commonsourceibias.t85 gnd 0.144227f
C5871 commonsourceibias.n341 gnd 0.057546f
C5872 commonsourceibias.n342 gnd 0.00772f
C5873 commonsourceibias.t93 gnd 0.144227f
C5874 commonsourceibias.n343 gnd 0.006245f
C5875 commonsourceibias.n344 gnd 0.00772f
C5876 commonsourceibias.t56 gnd 0.144227f
C5877 commonsourceibias.n345 gnd 0.007453f
C5878 commonsourceibias.n346 gnd 0.00772f
C5879 commonsourceibias.t89 gnd 0.144227f
C5880 commonsourceibias.n347 gnd 0.006235f
C5881 commonsourceibias.n348 gnd 0.00772f
C5882 commonsourceibias.t87 gnd 0.144227f
C5883 commonsourceibias.t74 gnd 0.144227f
C5884 commonsourceibias.n349 gnd 0.057546f
C5885 commonsourceibias.n350 gnd 0.00772f
C5886 commonsourceibias.t70 gnd 0.144227f
C5887 commonsourceibias.n351 gnd 0.057546f
C5888 commonsourceibias.n352 gnd 0.00772f
C5889 commonsourceibias.t82 gnd 0.144227f
C5890 commonsourceibias.n353 gnd 0.057546f
C5891 commonsourceibias.n354 gnd 0.038863f
C5892 commonsourceibias.t52 gnd 0.144227f
C5893 commonsourceibias.t65 gnd 0.162743f
C5894 commonsourceibias.n355 gnd 0.066782f
C5895 commonsourceibias.n356 gnd 0.069137f
C5896 commonsourceibias.n357 gnd 0.009515f
C5897 commonsourceibias.n358 gnd 0.010526f
C5898 commonsourceibias.n359 gnd 0.00772f
C5899 commonsourceibias.n360 gnd 0.00772f
C5900 commonsourceibias.n361 gnd 0.010457f
C5901 commonsourceibias.n362 gnd 0.006245f
C5902 commonsourceibias.n363 gnd 0.010587f
C5903 commonsourceibias.n364 gnd 0.00772f
C5904 commonsourceibias.n365 gnd 0.00772f
C5905 commonsourceibias.n366 gnd 0.010651f
C5906 commonsourceibias.n367 gnd 0.009185f
C5907 commonsourceibias.n368 gnd 0.007453f
C5908 commonsourceibias.n369 gnd 0.00772f
C5909 commonsourceibias.n370 gnd 0.00772f
C5910 commonsourceibias.n371 gnd 0.009442f
C5911 commonsourceibias.n372 gnd 0.010598f
C5912 commonsourceibias.n373 gnd 0.057546f
C5913 commonsourceibias.n374 gnd 0.010527f
C5914 commonsourceibias.n375 gnd 0.00772f
C5915 commonsourceibias.n376 gnd 0.00772f
C5916 commonsourceibias.n377 gnd 0.00772f
C5917 commonsourceibias.n378 gnd 0.010527f
C5918 commonsourceibias.n379 gnd 0.057546f
C5919 commonsourceibias.n380 gnd 0.010598f
C5920 commonsourceibias.t79 gnd 0.144227f
C5921 commonsourceibias.n381 gnd 0.057546f
C5922 commonsourceibias.n382 gnd 0.009442f
C5923 commonsourceibias.n383 gnd 0.00772f
C5924 commonsourceibias.n384 gnd 0.00772f
C5925 commonsourceibias.n385 gnd 0.00772f
C5926 commonsourceibias.n386 gnd 0.009185f
C5927 commonsourceibias.n387 gnd 0.010651f
C5928 commonsourceibias.n388 gnd 0.057546f
C5929 commonsourceibias.n389 gnd 0.010587f
C5930 commonsourceibias.n390 gnd 0.00772f
C5931 commonsourceibias.n391 gnd 0.00772f
C5932 commonsourceibias.n392 gnd 0.00772f
C5933 commonsourceibias.n393 gnd 0.010457f
C5934 commonsourceibias.n394 gnd 0.057546f
C5935 commonsourceibias.n395 gnd 0.010526f
C5936 commonsourceibias.n396 gnd 0.009515f
C5937 commonsourceibias.n397 gnd 0.00772f
C5938 commonsourceibias.n398 gnd 0.00772f
C5939 commonsourceibias.n399 gnd 0.007831f
C5940 commonsourceibias.n400 gnd 0.008096f
C5941 commonsourceibias.t73 gnd 0.155981f
C5942 commonsourceibias.n401 gnd 0.068855f
C5943 commonsourceibias.n402 gnd 0.023432f
C5944 commonsourceibias.n403 gnd 0.212991f
C5945 commonsourceibias.n404 gnd 4.01312f
.ends

