* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t31 plus.t0 drain_left.t5 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X1 a_n1886_n2088# a_n1886_n2088# a_n1886_n2088# a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=22.8 ps=103.6 w=6 l=0.15
X2 source.t0 minus.t0 drain_right.t15 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X3 drain_left.t10 plus.t1 source.t30 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X4 drain_left.t8 plus.t2 source.t29 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X5 drain_right.t14 minus.t1 source.t14 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X6 drain_right.t13 minus.t2 source.t2 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X7 source.t28 plus.t3 drain_left.t4 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X8 a_n1886_n2088# a_n1886_n2088# a_n1886_n2088# a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X9 a_n1886_n2088# a_n1886_n2088# a_n1886_n2088# a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X10 source.t9 minus.t3 drain_right.t12 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X11 a_n1886_n2088# a_n1886_n2088# a_n1886_n2088# a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X12 source.t11 minus.t4 drain_right.t11 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X13 source.t6 minus.t5 drain_right.t10 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X14 drain_right.t9 minus.t6 source.t15 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X15 drain_right.t8 minus.t7 source.t7 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X16 drain_right.t7 minus.t8 source.t10 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X17 source.t12 minus.t9 drain_right.t6 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X18 drain_right.t5 minus.t10 source.t4 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X19 drain_left.t13 plus.t4 source.t27 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X20 source.t26 plus.t5 drain_left.t9 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X21 drain_right.t4 minus.t11 source.t1 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X22 drain_right.t3 minus.t12 source.t3 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X23 source.t5 minus.t13 drain_right.t2 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X24 source.t13 minus.t14 drain_right.t1 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X25 source.t25 plus.t6 drain_left.t7 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X26 drain_left.t14 plus.t7 source.t24 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X27 source.t8 minus.t15 drain_right.t0 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X28 source.t23 plus.t8 drain_left.t0 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X29 source.t22 plus.t9 drain_left.t2 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X30 drain_left.t15 plus.t10 source.t21 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X31 drain_left.t12 plus.t11 source.t20 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X32 drain_left.t11 plus.t12 source.t19 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X33 source.t18 plus.t13 drain_left.t6 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X34 drain_left.t3 plus.t14 source.t17 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X35 source.t16 plus.t15 drain_left.t1 a_n1886_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
R0 plus.n5 plus.t5 1213.03
R1 plus.n21 plus.t4 1213.03
R2 plus.n28 plus.t1 1213.03
R3 plus.n44 plus.t13 1213.03
R4 plus.n6 plus.t12 1172.87
R5 plus.n3 plus.t9 1172.87
R6 plus.n12 plus.t7 1172.87
R7 plus.n14 plus.t15 1172.87
R8 plus.n1 plus.t11 1172.87
R9 plus.n20 plus.t8 1172.87
R10 plus.n29 plus.t3 1172.87
R11 plus.n26 plus.t10 1172.87
R12 plus.n35 plus.t0 1172.87
R13 plus.n37 plus.t2 1172.87
R14 plus.n24 plus.t6 1172.87
R15 plus.n43 plus.t14 1172.87
R16 plus.n5 plus.n4 161.489
R17 plus.n28 plus.n27 161.489
R18 plus.n7 plus.n4 161.3
R19 plus.n9 plus.n8 161.3
R20 plus.n11 plus.n10 161.3
R21 plus.n13 plus.n2 161.3
R22 plus.n16 plus.n15 161.3
R23 plus.n18 plus.n17 161.3
R24 plus.n19 plus.n0 161.3
R25 plus.n22 plus.n21 161.3
R26 plus.n30 plus.n27 161.3
R27 plus.n32 plus.n31 161.3
R28 plus.n34 plus.n33 161.3
R29 plus.n36 plus.n25 161.3
R30 plus.n39 plus.n38 161.3
R31 plus.n41 plus.n40 161.3
R32 plus.n42 plus.n23 161.3
R33 plus.n45 plus.n44 161.3
R34 plus.n8 plus.n7 73.0308
R35 plus.n19 plus.n18 73.0308
R36 plus.n42 plus.n41 73.0308
R37 plus.n31 plus.n30 73.0308
R38 plus.n11 plus.n3 69.3793
R39 plus.n15 plus.n1 69.3793
R40 plus.n38 plus.n24 69.3793
R41 plus.n34 plus.n26 69.3793
R42 plus.n6 plus.n5 54.7732
R43 plus.n21 plus.n20 54.7732
R44 plus.n44 plus.n43 54.7732
R45 plus.n29 plus.n28 54.7732
R46 plus.n13 plus.n12 47.4702
R47 plus.n14 plus.n13 47.4702
R48 plus.n37 plus.n36 47.4702
R49 plus.n36 plus.n35 47.4702
R50 plus plus.n45 27.8778
R51 plus.n12 plus.n11 25.5611
R52 plus.n15 plus.n14 25.5611
R53 plus.n38 plus.n37 25.5611
R54 plus.n35 plus.n34 25.5611
R55 plus.n7 plus.n6 18.2581
R56 plus.n20 plus.n19 18.2581
R57 plus.n43 plus.n42 18.2581
R58 plus.n30 plus.n29 18.2581
R59 plus plus.n22 9.8755
R60 plus.n8 plus.n3 3.65202
R61 plus.n18 plus.n1 3.65202
R62 plus.n41 plus.n24 3.65202
R63 plus.n31 plus.n26 3.65202
R64 plus.n9 plus.n4 0.189894
R65 plus.n10 plus.n9 0.189894
R66 plus.n10 plus.n2 0.189894
R67 plus.n16 plus.n2 0.189894
R68 plus.n17 plus.n16 0.189894
R69 plus.n17 plus.n0 0.189894
R70 plus.n22 plus.n0 0.189894
R71 plus.n45 plus.n23 0.189894
R72 plus.n40 plus.n23 0.189894
R73 plus.n40 plus.n39 0.189894
R74 plus.n39 plus.n25 0.189894
R75 plus.n33 plus.n25 0.189894
R76 plus.n33 plus.n32 0.189894
R77 plus.n32 plus.n27 0.189894
R78 drain_left.n9 drain_left.n7 67.7512
R79 drain_left.n5 drain_left.n3 67.751
R80 drain_left.n2 drain_left.n0 67.751
R81 drain_left.n11 drain_left.n10 67.1908
R82 drain_left.n9 drain_left.n8 67.1908
R83 drain_left.n13 drain_left.n12 67.1907
R84 drain_left.n5 drain_left.n4 67.1907
R85 drain_left.n2 drain_left.n1 67.1907
R86 drain_left drain_left.n6 26.4639
R87 drain_left drain_left.n13 6.21356
R88 drain_left.n3 drain_left.t4 5.0005
R89 drain_left.n3 drain_left.t10 5.0005
R90 drain_left.n4 drain_left.t5 5.0005
R91 drain_left.n4 drain_left.t15 5.0005
R92 drain_left.n1 drain_left.t7 5.0005
R93 drain_left.n1 drain_left.t8 5.0005
R94 drain_left.n0 drain_left.t6 5.0005
R95 drain_left.n0 drain_left.t3 5.0005
R96 drain_left.n12 drain_left.t0 5.0005
R97 drain_left.n12 drain_left.t13 5.0005
R98 drain_left.n10 drain_left.t1 5.0005
R99 drain_left.n10 drain_left.t12 5.0005
R100 drain_left.n8 drain_left.t2 5.0005
R101 drain_left.n8 drain_left.t14 5.0005
R102 drain_left.n7 drain_left.t9 5.0005
R103 drain_left.n7 drain_left.t11 5.0005
R104 drain_left.n11 drain_left.n9 0.560845
R105 drain_left.n13 drain_left.n11 0.560845
R106 drain_left.n6 drain_left.n5 0.225326
R107 drain_left.n6 drain_left.n2 0.225326
R108 source.n7 source.t26 55.512
R109 source.n8 source.t15 55.512
R110 source.n15 source.t13 55.512
R111 source.n0 source.t27 55.5119
R112 source.n31 source.t4 55.5119
R113 source.n24 source.t5 55.5119
R114 source.n23 source.t30 55.5119
R115 source.n16 source.t18 55.5119
R116 source.n2 source.n1 50.512
R117 source.n4 source.n3 50.512
R118 source.n6 source.n5 50.512
R119 source.n10 source.n9 50.512
R120 source.n12 source.n11 50.512
R121 source.n14 source.n13 50.512
R122 source.n30 source.n29 50.5119
R123 source.n28 source.n27 50.5119
R124 source.n26 source.n25 50.5119
R125 source.n22 source.n21 50.5119
R126 source.n20 source.n19 50.5119
R127 source.n18 source.n17 50.5119
R128 source.n16 source.n15 17.3026
R129 source.n32 source.n0 11.7595
R130 source.n32 source.n31 5.5436
R131 source.n29 source.t2 5.0005
R132 source.n29 source.t11 5.0005
R133 source.n27 source.t10 5.0005
R134 source.n27 source.t0 5.0005
R135 source.n25 source.t14 5.0005
R136 source.n25 source.t9 5.0005
R137 source.n21 source.t21 5.0005
R138 source.n21 source.t28 5.0005
R139 source.n19 source.t29 5.0005
R140 source.n19 source.t31 5.0005
R141 source.n17 source.t17 5.0005
R142 source.n17 source.t25 5.0005
R143 source.n1 source.t20 5.0005
R144 source.n1 source.t23 5.0005
R145 source.n3 source.t24 5.0005
R146 source.n3 source.t16 5.0005
R147 source.n5 source.t19 5.0005
R148 source.n5 source.t22 5.0005
R149 source.n9 source.t1 5.0005
R150 source.n9 source.t6 5.0005
R151 source.n11 source.t7 5.0005
R152 source.n11 source.t12 5.0005
R153 source.n13 source.t3 5.0005
R154 source.n13 source.t8 5.0005
R155 source.n15 source.n14 0.560845
R156 source.n14 source.n12 0.560845
R157 source.n12 source.n10 0.560845
R158 source.n10 source.n8 0.560845
R159 source.n7 source.n6 0.560845
R160 source.n6 source.n4 0.560845
R161 source.n4 source.n2 0.560845
R162 source.n2 source.n0 0.560845
R163 source.n18 source.n16 0.560845
R164 source.n20 source.n18 0.560845
R165 source.n22 source.n20 0.560845
R166 source.n23 source.n22 0.560845
R167 source.n26 source.n24 0.560845
R168 source.n28 source.n26 0.560845
R169 source.n30 source.n28 0.560845
R170 source.n31 source.n30 0.560845
R171 source.n8 source.n7 0.470328
R172 source.n24 source.n23 0.470328
R173 source source.n32 0.188
R174 minus.n21 minus.t14 1213.03
R175 minus.n5 minus.t6 1213.03
R176 minus.n44 minus.t10 1213.03
R177 minus.n28 minus.t13 1213.03
R178 minus.n20 minus.t12 1172.87
R179 minus.n1 minus.t15 1172.87
R180 minus.n14 minus.t7 1172.87
R181 minus.n12 minus.t9 1172.87
R182 minus.n3 minus.t11 1172.87
R183 minus.n6 minus.t5 1172.87
R184 minus.n43 minus.t4 1172.87
R185 minus.n24 minus.t2 1172.87
R186 minus.n37 minus.t0 1172.87
R187 minus.n35 minus.t8 1172.87
R188 minus.n26 minus.t3 1172.87
R189 minus.n29 minus.t1 1172.87
R190 minus.n5 minus.n4 161.489
R191 minus.n28 minus.n27 161.489
R192 minus.n22 minus.n21 161.3
R193 minus.n19 minus.n0 161.3
R194 minus.n18 minus.n17 161.3
R195 minus.n16 minus.n15 161.3
R196 minus.n13 minus.n2 161.3
R197 minus.n11 minus.n10 161.3
R198 minus.n9 minus.n8 161.3
R199 minus.n7 minus.n4 161.3
R200 minus.n45 minus.n44 161.3
R201 minus.n42 minus.n23 161.3
R202 minus.n41 minus.n40 161.3
R203 minus.n39 minus.n38 161.3
R204 minus.n36 minus.n25 161.3
R205 minus.n34 minus.n33 161.3
R206 minus.n32 minus.n31 161.3
R207 minus.n30 minus.n27 161.3
R208 minus.n19 minus.n18 73.0308
R209 minus.n8 minus.n7 73.0308
R210 minus.n31 minus.n30 73.0308
R211 minus.n42 minus.n41 73.0308
R212 minus.n15 minus.n1 69.3793
R213 minus.n11 minus.n3 69.3793
R214 minus.n34 minus.n26 69.3793
R215 minus.n38 minus.n24 69.3793
R216 minus.n21 minus.n20 54.7732
R217 minus.n6 minus.n5 54.7732
R218 minus.n29 minus.n28 54.7732
R219 minus.n44 minus.n43 54.7732
R220 minus.n14 minus.n13 47.4702
R221 minus.n13 minus.n12 47.4702
R222 minus.n36 minus.n35 47.4702
R223 minus.n37 minus.n36 47.4702
R224 minus.n46 minus.n22 31.724
R225 minus.n15 minus.n14 25.5611
R226 minus.n12 minus.n11 25.5611
R227 minus.n35 minus.n34 25.5611
R228 minus.n38 minus.n37 25.5611
R229 minus.n20 minus.n19 18.2581
R230 minus.n7 minus.n6 18.2581
R231 minus.n30 minus.n29 18.2581
R232 minus.n43 minus.n42 18.2581
R233 minus.n46 minus.n45 6.50429
R234 minus.n18 minus.n1 3.65202
R235 minus.n8 minus.n3 3.65202
R236 minus.n31 minus.n26 3.65202
R237 minus.n41 minus.n24 3.65202
R238 minus.n22 minus.n0 0.189894
R239 minus.n17 minus.n0 0.189894
R240 minus.n17 minus.n16 0.189894
R241 minus.n16 minus.n2 0.189894
R242 minus.n10 minus.n2 0.189894
R243 minus.n10 minus.n9 0.189894
R244 minus.n9 minus.n4 0.189894
R245 minus.n32 minus.n27 0.189894
R246 minus.n33 minus.n32 0.189894
R247 minus.n33 minus.n25 0.189894
R248 minus.n39 minus.n25 0.189894
R249 minus.n40 minus.n39 0.189894
R250 minus.n40 minus.n23 0.189894
R251 minus.n45 minus.n23 0.189894
R252 minus minus.n46 0.188
R253 drain_right.n9 drain_right.n7 67.751
R254 drain_right.n5 drain_right.n3 67.751
R255 drain_right.n2 drain_right.n0 67.751
R256 drain_right.n9 drain_right.n8 67.1908
R257 drain_right.n11 drain_right.n10 67.1908
R258 drain_right.n13 drain_right.n12 67.1908
R259 drain_right.n5 drain_right.n4 67.1907
R260 drain_right.n2 drain_right.n1 67.1907
R261 drain_right drain_right.n6 25.9106
R262 drain_right drain_right.n13 6.21356
R263 drain_right.n3 drain_right.t11 5.0005
R264 drain_right.n3 drain_right.t5 5.0005
R265 drain_right.n4 drain_right.t15 5.0005
R266 drain_right.n4 drain_right.t13 5.0005
R267 drain_right.n1 drain_right.t12 5.0005
R268 drain_right.n1 drain_right.t7 5.0005
R269 drain_right.n0 drain_right.t2 5.0005
R270 drain_right.n0 drain_right.t14 5.0005
R271 drain_right.n7 drain_right.t10 5.0005
R272 drain_right.n7 drain_right.t9 5.0005
R273 drain_right.n8 drain_right.t6 5.0005
R274 drain_right.n8 drain_right.t4 5.0005
R275 drain_right.n10 drain_right.t0 5.0005
R276 drain_right.n10 drain_right.t8 5.0005
R277 drain_right.n12 drain_right.t1 5.0005
R278 drain_right.n12 drain_right.t3 5.0005
R279 drain_right.n13 drain_right.n11 0.560845
R280 drain_right.n11 drain_right.n9 0.560845
R281 drain_right.n6 drain_right.n5 0.225326
R282 drain_right.n6 drain_right.n2 0.225326
C0 minus source 1.88403f
C1 drain_right plus 0.337321f
C2 drain_left source 17.0188f
C3 drain_right minus 2.03599f
C4 drain_right drain_left 0.96779f
C5 plus minus 4.38124f
C6 plus drain_left 2.21958f
C7 drain_left minus 0.170952f
C8 drain_right source 17.0191f
C9 plus source 1.89805f
C10 drain_right a_n1886_n2088# 4.91085f
C11 drain_left a_n1886_n2088# 5.19746f
C12 source a_n1886_n2088# 5.417755f
C13 minus a_n1886_n2088# 6.48188f
C14 plus a_n1886_n2088# 7.77649f
C15 drain_right.t2 a_n1886_n2088# 0.2012f
C16 drain_right.t14 a_n1886_n2088# 0.2012f
C17 drain_right.n0 a_n1886_n2088# 1.24711f
C18 drain_right.t12 a_n1886_n2088# 0.2012f
C19 drain_right.t7 a_n1886_n2088# 0.2012f
C20 drain_right.n1 a_n1886_n2088# 1.2443f
C21 drain_right.n2 a_n1886_n2088# 0.637981f
C22 drain_right.t11 a_n1886_n2088# 0.2012f
C23 drain_right.t5 a_n1886_n2088# 0.2012f
C24 drain_right.n3 a_n1886_n2088# 1.24711f
C25 drain_right.t15 a_n1886_n2088# 0.2012f
C26 drain_right.t13 a_n1886_n2088# 0.2012f
C27 drain_right.n4 a_n1886_n2088# 1.2443f
C28 drain_right.n5 a_n1886_n2088# 0.637981f
C29 drain_right.n6 a_n1886_n2088# 0.962524f
C30 drain_right.t10 a_n1886_n2088# 0.2012f
C31 drain_right.t9 a_n1886_n2088# 0.2012f
C32 drain_right.n7 a_n1886_n2088# 1.24711f
C33 drain_right.t6 a_n1886_n2088# 0.2012f
C34 drain_right.t4 a_n1886_n2088# 0.2012f
C35 drain_right.n8 a_n1886_n2088# 1.2443f
C36 drain_right.n9 a_n1886_n2088# 0.665367f
C37 drain_right.t0 a_n1886_n2088# 0.2012f
C38 drain_right.t8 a_n1886_n2088# 0.2012f
C39 drain_right.n10 a_n1886_n2088# 1.2443f
C40 drain_right.n11 a_n1886_n2088# 0.328445f
C41 drain_right.t1 a_n1886_n2088# 0.2012f
C42 drain_right.t3 a_n1886_n2088# 0.2012f
C43 drain_right.n12 a_n1886_n2088# 1.2443f
C44 drain_right.n13 a_n1886_n2088# 0.562333f
C45 minus.n0 a_n1886_n2088# 0.040873f
C46 minus.t14 a_n1886_n2088# 0.106548f
C47 minus.t12 a_n1886_n2088# 0.104809f
C48 minus.t15 a_n1886_n2088# 0.104809f
C49 minus.n1 a_n1886_n2088# 0.054409f
C50 minus.n2 a_n1886_n2088# 0.040873f
C51 minus.t7 a_n1886_n2088# 0.104809f
C52 minus.t9 a_n1886_n2088# 0.104809f
C53 minus.t11 a_n1886_n2088# 0.104809f
C54 minus.n3 a_n1886_n2088# 0.054409f
C55 minus.n4 a_n1886_n2088# 0.086732f
C56 minus.t5 a_n1886_n2088# 0.104809f
C57 minus.t6 a_n1886_n2088# 0.106548f
C58 minus.n5 a_n1886_n2088# 0.068173f
C59 minus.n6 a_n1886_n2088# 0.054409f
C60 minus.n7 a_n1886_n2088# 0.016709f
C61 minus.n8 a_n1886_n2088# 0.014189f
C62 minus.n9 a_n1886_n2088# 0.040873f
C63 minus.n10 a_n1886_n2088# 0.040873f
C64 minus.n11 a_n1886_n2088# 0.017339f
C65 minus.n12 a_n1886_n2088# 0.054409f
C66 minus.n13 a_n1886_n2088# 0.017339f
C67 minus.n14 a_n1886_n2088# 0.054409f
C68 minus.n15 a_n1886_n2088# 0.017339f
C69 minus.n16 a_n1886_n2088# 0.040873f
C70 minus.n17 a_n1886_n2088# 0.040873f
C71 minus.n18 a_n1886_n2088# 0.014189f
C72 minus.n19 a_n1886_n2088# 0.016709f
C73 minus.n20 a_n1886_n2088# 0.054409f
C74 minus.n21 a_n1886_n2088# 0.068119f
C75 minus.n22 a_n1886_n2088# 1.16833f
C76 minus.n23 a_n1886_n2088# 0.040873f
C77 minus.t4 a_n1886_n2088# 0.104809f
C78 minus.t2 a_n1886_n2088# 0.104809f
C79 minus.n24 a_n1886_n2088# 0.054409f
C80 minus.n25 a_n1886_n2088# 0.040873f
C81 minus.t0 a_n1886_n2088# 0.104809f
C82 minus.t8 a_n1886_n2088# 0.104809f
C83 minus.t3 a_n1886_n2088# 0.104809f
C84 minus.n26 a_n1886_n2088# 0.054409f
C85 minus.n27 a_n1886_n2088# 0.086732f
C86 minus.t1 a_n1886_n2088# 0.104809f
C87 minus.t13 a_n1886_n2088# 0.106548f
C88 minus.n28 a_n1886_n2088# 0.068173f
C89 minus.n29 a_n1886_n2088# 0.054409f
C90 minus.n30 a_n1886_n2088# 0.016709f
C91 minus.n31 a_n1886_n2088# 0.014189f
C92 minus.n32 a_n1886_n2088# 0.040873f
C93 minus.n33 a_n1886_n2088# 0.040873f
C94 minus.n34 a_n1886_n2088# 0.017339f
C95 minus.n35 a_n1886_n2088# 0.054409f
C96 minus.n36 a_n1886_n2088# 0.017339f
C97 minus.n37 a_n1886_n2088# 0.054409f
C98 minus.n38 a_n1886_n2088# 0.017339f
C99 minus.n39 a_n1886_n2088# 0.040873f
C100 minus.n40 a_n1886_n2088# 0.040873f
C101 minus.n41 a_n1886_n2088# 0.014189f
C102 minus.n42 a_n1886_n2088# 0.016709f
C103 minus.n43 a_n1886_n2088# 0.054409f
C104 minus.t10 a_n1886_n2088# 0.106548f
C105 minus.n44 a_n1886_n2088# 0.068119f
C106 minus.n45 a_n1886_n2088# 0.26763f
C107 minus.n46 a_n1886_n2088# 1.43624f
C108 source.t27 a_n1886_n2088# 1.14069f
C109 source.n0 a_n1886_n2088# 0.839181f
C110 source.t20 a_n1886_n2088# 0.162404f
C111 source.t23 a_n1886_n2088# 0.162404f
C112 source.n1 a_n1886_n2088# 0.945211f
C113 source.n2 a_n1886_n2088# 0.29355f
C114 source.t24 a_n1886_n2088# 0.162404f
C115 source.t16 a_n1886_n2088# 0.162404f
C116 source.n3 a_n1886_n2088# 0.945211f
C117 source.n4 a_n1886_n2088# 0.29355f
C118 source.t19 a_n1886_n2088# 0.162404f
C119 source.t22 a_n1886_n2088# 0.162404f
C120 source.n5 a_n1886_n2088# 0.945211f
C121 source.n6 a_n1886_n2088# 0.29355f
C122 source.t26 a_n1886_n2088# 1.1407f
C123 source.n7 a_n1886_n2088# 0.383795f
C124 source.t15 a_n1886_n2088# 1.1407f
C125 source.n8 a_n1886_n2088# 0.383795f
C126 source.t1 a_n1886_n2088# 0.162404f
C127 source.t6 a_n1886_n2088# 0.162404f
C128 source.n9 a_n1886_n2088# 0.945211f
C129 source.n10 a_n1886_n2088# 0.29355f
C130 source.t7 a_n1886_n2088# 0.162404f
C131 source.t12 a_n1886_n2088# 0.162404f
C132 source.n11 a_n1886_n2088# 0.945211f
C133 source.n12 a_n1886_n2088# 0.29355f
C134 source.t3 a_n1886_n2088# 0.162404f
C135 source.t8 a_n1886_n2088# 0.162404f
C136 source.n13 a_n1886_n2088# 0.945211f
C137 source.n14 a_n1886_n2088# 0.29355f
C138 source.t13 a_n1886_n2088# 1.1407f
C139 source.n15 a_n1886_n2088# 1.13057f
C140 source.t18 a_n1886_n2088# 1.14069f
C141 source.n16 a_n1886_n2088# 1.13058f
C142 source.t17 a_n1886_n2088# 0.162404f
C143 source.t25 a_n1886_n2088# 0.162404f
C144 source.n17 a_n1886_n2088# 0.945205f
C145 source.n18 a_n1886_n2088# 0.293556f
C146 source.t29 a_n1886_n2088# 0.162404f
C147 source.t31 a_n1886_n2088# 0.162404f
C148 source.n19 a_n1886_n2088# 0.945205f
C149 source.n20 a_n1886_n2088# 0.293556f
C150 source.t21 a_n1886_n2088# 0.162404f
C151 source.t28 a_n1886_n2088# 0.162404f
C152 source.n21 a_n1886_n2088# 0.945205f
C153 source.n22 a_n1886_n2088# 0.293556f
C154 source.t30 a_n1886_n2088# 1.14069f
C155 source.n23 a_n1886_n2088# 0.3838f
C156 source.t5 a_n1886_n2088# 1.14069f
C157 source.n24 a_n1886_n2088# 0.3838f
C158 source.t14 a_n1886_n2088# 0.162404f
C159 source.t9 a_n1886_n2088# 0.162404f
C160 source.n25 a_n1886_n2088# 0.945205f
C161 source.n26 a_n1886_n2088# 0.293556f
C162 source.t10 a_n1886_n2088# 0.162404f
C163 source.t0 a_n1886_n2088# 0.162404f
C164 source.n27 a_n1886_n2088# 0.945205f
C165 source.n28 a_n1886_n2088# 0.293556f
C166 source.t2 a_n1886_n2088# 0.162404f
C167 source.t11 a_n1886_n2088# 0.162404f
C168 source.n29 a_n1886_n2088# 0.945205f
C169 source.n30 a_n1886_n2088# 0.293556f
C170 source.t4 a_n1886_n2088# 1.14069f
C171 source.n31 a_n1886_n2088# 0.512418f
C172 source.n32 a_n1886_n2088# 0.925632f
C173 drain_left.t6 a_n1886_n2088# 0.202152f
C174 drain_left.t3 a_n1886_n2088# 0.202152f
C175 drain_left.n0 a_n1886_n2088# 1.25301f
C176 drain_left.t7 a_n1886_n2088# 0.202152f
C177 drain_left.t8 a_n1886_n2088# 0.202152f
C178 drain_left.n1 a_n1886_n2088# 1.25019f
C179 drain_left.n2 a_n1886_n2088# 0.641001f
C180 drain_left.t4 a_n1886_n2088# 0.202152f
C181 drain_left.t10 a_n1886_n2088# 0.202152f
C182 drain_left.n3 a_n1886_n2088# 1.25301f
C183 drain_left.t5 a_n1886_n2088# 0.202152f
C184 drain_left.t15 a_n1886_n2088# 0.202152f
C185 drain_left.n4 a_n1886_n2088# 1.25019f
C186 drain_left.n5 a_n1886_n2088# 0.641001f
C187 drain_left.n6 a_n1886_n2088# 1.02415f
C188 drain_left.t9 a_n1886_n2088# 0.202152f
C189 drain_left.t11 a_n1886_n2088# 0.202152f
C190 drain_left.n7 a_n1886_n2088# 1.25302f
C191 drain_left.t2 a_n1886_n2088# 0.202152f
C192 drain_left.t14 a_n1886_n2088# 0.202152f
C193 drain_left.n8 a_n1886_n2088# 1.25019f
C194 drain_left.n9 a_n1886_n2088# 0.668511f
C195 drain_left.t1 a_n1886_n2088# 0.202152f
C196 drain_left.t12 a_n1886_n2088# 0.202152f
C197 drain_left.n10 a_n1886_n2088# 1.25019f
C198 drain_left.n11 a_n1886_n2088# 0.33f
C199 drain_left.t0 a_n1886_n2088# 0.202152f
C200 drain_left.t13 a_n1886_n2088# 0.202152f
C201 drain_left.n12 a_n1886_n2088# 1.25019f
C202 drain_left.n13 a_n1886_n2088# 0.565f
C203 plus.n0 a_n1886_n2088# 0.042702f
C204 plus.t8 a_n1886_n2088# 0.109498f
C205 plus.t11 a_n1886_n2088# 0.109498f
C206 plus.n1 a_n1886_n2088# 0.056844f
C207 plus.n2 a_n1886_n2088# 0.042702f
C208 plus.t15 a_n1886_n2088# 0.109498f
C209 plus.t7 a_n1886_n2088# 0.109498f
C210 plus.t9 a_n1886_n2088# 0.109498f
C211 plus.n3 a_n1886_n2088# 0.056844f
C212 plus.n4 a_n1886_n2088# 0.090613f
C213 plus.t12 a_n1886_n2088# 0.109498f
C214 plus.t5 a_n1886_n2088# 0.111315f
C215 plus.n5 a_n1886_n2088# 0.071223f
C216 plus.n6 a_n1886_n2088# 0.056844f
C217 plus.n7 a_n1886_n2088# 0.017456f
C218 plus.n8 a_n1886_n2088# 0.014824f
C219 plus.n9 a_n1886_n2088# 0.042702f
C220 plus.n10 a_n1886_n2088# 0.042702f
C221 plus.n11 a_n1886_n2088# 0.018115f
C222 plus.n12 a_n1886_n2088# 0.056844f
C223 plus.n13 a_n1886_n2088# 0.018115f
C224 plus.n14 a_n1886_n2088# 0.056844f
C225 plus.n15 a_n1886_n2088# 0.018115f
C226 plus.n16 a_n1886_n2088# 0.042702f
C227 plus.n17 a_n1886_n2088# 0.042702f
C228 plus.n18 a_n1886_n2088# 0.014824f
C229 plus.n19 a_n1886_n2088# 0.017456f
C230 plus.n20 a_n1886_n2088# 0.056844f
C231 plus.t4 a_n1886_n2088# 0.111315f
C232 plus.n21 a_n1886_n2088# 0.071167f
C233 plus.n22 a_n1886_n2088# 0.366359f
C234 plus.n23 a_n1886_n2088# 0.042702f
C235 plus.t13 a_n1886_n2088# 0.111315f
C236 plus.t14 a_n1886_n2088# 0.109498f
C237 plus.t6 a_n1886_n2088# 0.109498f
C238 plus.n24 a_n1886_n2088# 0.056844f
C239 plus.n25 a_n1886_n2088# 0.042702f
C240 plus.t2 a_n1886_n2088# 0.109498f
C241 plus.t0 a_n1886_n2088# 0.109498f
C242 plus.t10 a_n1886_n2088# 0.109498f
C243 plus.n26 a_n1886_n2088# 0.056844f
C244 plus.n27 a_n1886_n2088# 0.090613f
C245 plus.t3 a_n1886_n2088# 0.109498f
C246 plus.t1 a_n1886_n2088# 0.111315f
C247 plus.n28 a_n1886_n2088# 0.071223f
C248 plus.n29 a_n1886_n2088# 0.056844f
C249 plus.n30 a_n1886_n2088# 0.017456f
C250 plus.n31 a_n1886_n2088# 0.014824f
C251 plus.n32 a_n1886_n2088# 0.042702f
C252 plus.n33 a_n1886_n2088# 0.042702f
C253 plus.n34 a_n1886_n2088# 0.018115f
C254 plus.n35 a_n1886_n2088# 0.056844f
C255 plus.n36 a_n1886_n2088# 0.018115f
C256 plus.n37 a_n1886_n2088# 0.056844f
C257 plus.n38 a_n1886_n2088# 0.018115f
C258 plus.n39 a_n1886_n2088# 0.042702f
C259 plus.n40 a_n1886_n2088# 0.042702f
C260 plus.n41 a_n1886_n2088# 0.014824f
C261 plus.n42 a_n1886_n2088# 0.017456f
C262 plus.n43 a_n1886_n2088# 0.056844f
C263 plus.n44 a_n1886_n2088# 0.071167f
C264 plus.n45 a_n1886_n2088# 1.10266f
.ends

