* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t47 plus.t0 drain_left.t2 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X1 drain_left.t0 plus.t1 source.t46 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X2 drain_right.t23 minus.t0 source.t6 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X3 drain_right.t22 minus.t1 source.t0 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X4 source.t45 plus.t2 drain_left.t1 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X5 source.t20 minus.t2 drain_right.t21 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X6 source.t44 plus.t3 drain_left.t23 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X7 drain_left.t3 plus.t4 source.t43 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X8 a_n2406_n1488# a_n2406_n1488# a_n2406_n1488# a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=11.4 ps=55.6 w=3 l=0.15
X9 drain_right.t20 minus.t3 source.t10 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X10 source.t14 minus.t4 drain_right.t19 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X11 drain_left.t4 plus.t5 source.t42 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X12 source.t8 minus.t5 drain_right.t18 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X13 a_n2406_n1488# a_n2406_n1488# a_n2406_n1488# a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X14 a_n2406_n1488# a_n2406_n1488# a_n2406_n1488# a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X15 source.t19 minus.t6 drain_right.t17 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X16 drain_right.t16 minus.t7 source.t23 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X17 source.t13 minus.t8 drain_right.t15 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X18 source.t41 plus.t6 drain_left.t5 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X19 drain_left.t6 plus.t7 source.t40 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X20 drain_right.t14 minus.t9 source.t15 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X21 drain_right.t13 minus.t10 source.t7 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X22 source.t12 minus.t11 drain_right.t12 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X23 source.t16 minus.t12 drain_right.t11 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X24 drain_left.t7 plus.t8 source.t39 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X25 drain_right.t10 minus.t13 source.t21 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X26 source.t38 plus.t9 drain_left.t8 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X27 drain_left.t9 plus.t10 source.t37 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X28 source.t36 plus.t11 drain_left.t10 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X29 drain_right.t9 minus.t14 source.t2 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X30 drain_right.t8 minus.t15 source.t9 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X31 source.t35 plus.t12 drain_left.t11 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X32 source.t11 minus.t16 drain_right.t7 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X33 source.t3 minus.t17 drain_right.t6 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X34 drain_left.t12 plus.t13 source.t34 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X35 source.t1 minus.t18 drain_right.t5 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X36 drain_right.t4 minus.t19 source.t5 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X37 drain_right.t3 minus.t20 source.t18 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X38 drain_left.t13 plus.t14 source.t33 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X39 source.t32 plus.t15 drain_left.t14 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X40 source.t31 plus.t16 drain_left.t15 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X41 drain_left.t16 plus.t17 source.t30 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X42 source.t17 minus.t21 drain_right.t2 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X43 source.t29 plus.t18 drain_left.t20 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X44 source.t28 plus.t19 drain_left.t21 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X45 drain_left.t17 plus.t20 source.t27 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X46 drain_left.t22 plus.t21 source.t26 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X47 a_n2406_n1488# a_n2406_n1488# a_n2406_n1488# a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X48 source.t22 minus.t22 drain_right.t1 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X49 drain_left.t18 plus.t22 source.t25 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X50 source.t24 plus.t23 drain_left.t19 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X51 drain_right.t0 minus.t23 source.t4 a_n2406_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
R0 plus.n6 plus.t11 738.337
R1 plus.n35 plus.t22 738.337
R2 plus.n45 plus.t4 738.337
R3 plus.n72 plus.t18 738.337
R4 plus.n7 plus.t21 690.867
R5 plus.n8 plus.t16 690.867
R6 plus.n14 plus.t13 690.867
R7 plus.n16 plus.t23 690.867
R8 plus.n17 plus.t20 690.867
R9 plus.n23 plus.t15 690.867
R10 plus.n25 plus.t10 690.867
R11 plus.n26 plus.t19 690.867
R12 plus.n32 plus.t14 690.867
R13 plus.n34 plus.t12 690.867
R14 plus.n47 plus.t2 690.867
R15 plus.n46 plus.t8 690.867
R16 plus.n53 plus.t6 690.867
R17 plus.n55 plus.t5 690.867
R18 plus.n43 plus.t0 690.867
R19 plus.n61 plus.t17 690.867
R20 plus.n63 plus.t9 690.867
R21 plus.n40 plus.t7 690.867
R22 plus.n69 plus.t3 690.867
R23 plus.n71 plus.t1 690.867
R24 plus.n10 plus.n6 161.489
R25 plus.n49 plus.n45 161.489
R26 plus.n10 plus.n9 161.3
R27 plus.n11 plus.n5 161.3
R28 plus.n13 plus.n12 161.3
R29 plus.n15 plus.n4 161.3
R30 plus.n19 plus.n18 161.3
R31 plus.n20 plus.n3 161.3
R32 plus.n22 plus.n21 161.3
R33 plus.n24 plus.n2 161.3
R34 plus.n28 plus.n27 161.3
R35 plus.n29 plus.n1 161.3
R36 plus.n31 plus.n30 161.3
R37 plus.n33 plus.n0 161.3
R38 plus.n36 plus.n35 161.3
R39 plus.n49 plus.n48 161.3
R40 plus.n50 plus.n44 161.3
R41 plus.n52 plus.n51 161.3
R42 plus.n54 plus.n42 161.3
R43 plus.n57 plus.n56 161.3
R44 plus.n58 plus.n41 161.3
R45 plus.n60 plus.n59 161.3
R46 plus.n62 plus.n39 161.3
R47 plus.n65 plus.n64 161.3
R48 plus.n66 plus.n38 161.3
R49 plus.n68 plus.n67 161.3
R50 plus.n70 plus.n37 161.3
R51 plus.n73 plus.n72 161.3
R52 plus.n13 plus.n5 73.0308
R53 plus.n22 plus.n3 73.0308
R54 plus.n31 plus.n1 73.0308
R55 plus.n68 plus.n38 73.0308
R56 plus.n60 plus.n41 73.0308
R57 plus.n52 plus.n44 73.0308
R58 plus.n9 plus.n8 69.3793
R59 plus.n33 plus.n32 69.3793
R60 plus.n70 plus.n69 69.3793
R61 plus.n48 plus.n46 69.3793
R62 plus.n18 plus.n17 62.0763
R63 plus.n24 plus.n23 62.0763
R64 plus.n62 plus.n61 62.0763
R65 plus.n56 plus.n43 62.0763
R66 plus.n15 plus.n14 54.7732
R67 plus.n27 plus.n26 54.7732
R68 plus.n64 plus.n40 54.7732
R69 plus.n54 plus.n53 54.7732
R70 plus.n7 plus.n6 47.4702
R71 plus.n35 plus.n34 47.4702
R72 plus.n72 plus.n71 47.4702
R73 plus.n47 plus.n45 47.4702
R74 plus.n16 plus.n15 40.1672
R75 plus.n27 plus.n25 40.1672
R76 plus.n64 plus.n63 40.1672
R77 plus.n55 plus.n54 40.1672
R78 plus.n18 plus.n16 32.8641
R79 plus.n25 plus.n24 32.8641
R80 plus.n63 plus.n62 32.8641
R81 plus.n56 plus.n55 32.8641
R82 plus plus.n73 28.7301
R83 plus.n9 plus.n7 25.5611
R84 plus.n34 plus.n33 25.5611
R85 plus.n71 plus.n70 25.5611
R86 plus.n48 plus.n47 25.5611
R87 plus.n14 plus.n13 18.2581
R88 plus.n26 plus.n1 18.2581
R89 plus.n40 plus.n38 18.2581
R90 plus.n53 plus.n52 18.2581
R91 plus.n17 plus.n3 10.955
R92 plus.n23 plus.n22 10.955
R93 plus.n61 plus.n60 10.955
R94 plus.n43 plus.n41 10.955
R95 plus plus.n36 8.75808
R96 plus.n8 plus.n5 3.65202
R97 plus.n32 plus.n31 3.65202
R98 plus.n69 plus.n68 3.65202
R99 plus.n46 plus.n44 3.65202
R100 plus.n11 plus.n10 0.189894
R101 plus.n12 plus.n11 0.189894
R102 plus.n12 plus.n4 0.189894
R103 plus.n19 plus.n4 0.189894
R104 plus.n20 plus.n19 0.189894
R105 plus.n21 plus.n20 0.189894
R106 plus.n21 plus.n2 0.189894
R107 plus.n28 plus.n2 0.189894
R108 plus.n29 plus.n28 0.189894
R109 plus.n30 plus.n29 0.189894
R110 plus.n30 plus.n0 0.189894
R111 plus.n36 plus.n0 0.189894
R112 plus.n73 plus.n37 0.189894
R113 plus.n67 plus.n37 0.189894
R114 plus.n67 plus.n66 0.189894
R115 plus.n66 plus.n65 0.189894
R116 plus.n65 plus.n39 0.189894
R117 plus.n59 plus.n39 0.189894
R118 plus.n59 plus.n58 0.189894
R119 plus.n58 plus.n57 0.189894
R120 plus.n57 plus.n42 0.189894
R121 plus.n51 plus.n42 0.189894
R122 plus.n51 plus.n50 0.189894
R123 plus.n50 plus.n49 0.189894
R124 drain_left.n13 drain_left.n11 80.3335
R125 drain_left.n7 drain_left.n5 80.3334
R126 drain_left.n2 drain_left.n0 80.3334
R127 drain_left.n21 drain_left.n20 79.7731
R128 drain_left.n19 drain_left.n18 79.7731
R129 drain_left.n17 drain_left.n16 79.7731
R130 drain_left.n15 drain_left.n14 79.7731
R131 drain_left.n13 drain_left.n12 79.7731
R132 drain_left.n7 drain_left.n6 79.773
R133 drain_left.n9 drain_left.n8 79.773
R134 drain_left.n4 drain_left.n3 79.773
R135 drain_left.n2 drain_left.n1 79.773
R136 drain_left drain_left.n10 25.8722
R137 drain_left.n5 drain_left.t1 10.0005
R138 drain_left.n5 drain_left.t3 10.0005
R139 drain_left.n6 drain_left.t5 10.0005
R140 drain_left.n6 drain_left.t7 10.0005
R141 drain_left.n8 drain_left.t2 10.0005
R142 drain_left.n8 drain_left.t4 10.0005
R143 drain_left.n3 drain_left.t8 10.0005
R144 drain_left.n3 drain_left.t16 10.0005
R145 drain_left.n1 drain_left.t23 10.0005
R146 drain_left.n1 drain_left.t6 10.0005
R147 drain_left.n0 drain_left.t20 10.0005
R148 drain_left.n0 drain_left.t0 10.0005
R149 drain_left.n20 drain_left.t11 10.0005
R150 drain_left.n20 drain_left.t18 10.0005
R151 drain_left.n18 drain_left.t21 10.0005
R152 drain_left.n18 drain_left.t13 10.0005
R153 drain_left.n16 drain_left.t14 10.0005
R154 drain_left.n16 drain_left.t9 10.0005
R155 drain_left.n14 drain_left.t19 10.0005
R156 drain_left.n14 drain_left.t17 10.0005
R157 drain_left.n12 drain_left.t15 10.0005
R158 drain_left.n12 drain_left.t12 10.0005
R159 drain_left.n11 drain_left.t10 10.0005
R160 drain_left.n11 drain_left.t22 10.0005
R161 drain_left drain_left.n21 6.21356
R162 drain_left.n9 drain_left.n7 0.560845
R163 drain_left.n4 drain_left.n2 0.560845
R164 drain_left.n15 drain_left.n13 0.560845
R165 drain_left.n17 drain_left.n15 0.560845
R166 drain_left.n19 drain_left.n17 0.560845
R167 drain_left.n21 drain_left.n19 0.560845
R168 drain_left.n10 drain_left.n9 0.225326
R169 drain_left.n10 drain_left.n4 0.225326
R170 source.n0 source.t25 73.0943
R171 source.n11 source.t36 73.0943
R172 source.n12 source.t15 73.0943
R173 source.n23 source.t3 73.0943
R174 source.n47 source.t4 73.0942
R175 source.n36 source.t19 73.0942
R176 source.n35 source.t43 73.0942
R177 source.n24 source.t29 73.0942
R178 source.n2 source.n1 63.0943
R179 source.n4 source.n3 63.0943
R180 source.n6 source.n5 63.0943
R181 source.n8 source.n7 63.0943
R182 source.n10 source.n9 63.0943
R183 source.n14 source.n13 63.0943
R184 source.n16 source.n15 63.0943
R185 source.n18 source.n17 63.0943
R186 source.n20 source.n19 63.0943
R187 source.n22 source.n21 63.0943
R188 source.n46 source.n45 63.0942
R189 source.n44 source.n43 63.0942
R190 source.n42 source.n41 63.0942
R191 source.n40 source.n39 63.0942
R192 source.n38 source.n37 63.0942
R193 source.n34 source.n33 63.0942
R194 source.n32 source.n31 63.0942
R195 source.n30 source.n29 63.0942
R196 source.n28 source.n27 63.0942
R197 source.n26 source.n25 63.0942
R198 source.n24 source.n23 15.0299
R199 source.n45 source.t23 10.0005
R200 source.n45 source.t14 10.0005
R201 source.n43 source.t6 10.0005
R202 source.n43 source.t16 10.0005
R203 source.n41 source.t10 10.0005
R204 source.n41 source.t20 10.0005
R205 source.n39 source.t5 10.0005
R206 source.n39 source.t8 10.0005
R207 source.n37 source.t0 10.0005
R208 source.n37 source.t22 10.0005
R209 source.n33 source.t39 10.0005
R210 source.n33 source.t45 10.0005
R211 source.n31 source.t42 10.0005
R212 source.n31 source.t41 10.0005
R213 source.n29 source.t30 10.0005
R214 source.n29 source.t47 10.0005
R215 source.n27 source.t40 10.0005
R216 source.n27 source.t38 10.0005
R217 source.n25 source.t46 10.0005
R218 source.n25 source.t44 10.0005
R219 source.n1 source.t33 10.0005
R220 source.n1 source.t35 10.0005
R221 source.n3 source.t37 10.0005
R222 source.n3 source.t28 10.0005
R223 source.n5 source.t27 10.0005
R224 source.n5 source.t32 10.0005
R225 source.n7 source.t34 10.0005
R226 source.n7 source.t24 10.0005
R227 source.n9 source.t26 10.0005
R228 source.n9 source.t31 10.0005
R229 source.n13 source.t2 10.0005
R230 source.n13 source.t13 10.0005
R231 source.n15 source.t7 10.0005
R232 source.n15 source.t12 10.0005
R233 source.n17 source.t9 10.0005
R234 source.n17 source.t1 10.0005
R235 source.n19 source.t21 10.0005
R236 source.n19 source.t11 10.0005
R237 source.n21 source.t18 10.0005
R238 source.n21 source.t17 10.0005
R239 source.n48 source.n0 9.48679
R240 source.n48 source.n47 5.5436
R241 source.n23 source.n22 0.560845
R242 source.n22 source.n20 0.560845
R243 source.n20 source.n18 0.560845
R244 source.n18 source.n16 0.560845
R245 source.n16 source.n14 0.560845
R246 source.n14 source.n12 0.560845
R247 source.n11 source.n10 0.560845
R248 source.n10 source.n8 0.560845
R249 source.n8 source.n6 0.560845
R250 source.n6 source.n4 0.560845
R251 source.n4 source.n2 0.560845
R252 source.n2 source.n0 0.560845
R253 source.n26 source.n24 0.560845
R254 source.n28 source.n26 0.560845
R255 source.n30 source.n28 0.560845
R256 source.n32 source.n30 0.560845
R257 source.n34 source.n32 0.560845
R258 source.n35 source.n34 0.560845
R259 source.n38 source.n36 0.560845
R260 source.n40 source.n38 0.560845
R261 source.n42 source.n40 0.560845
R262 source.n44 source.n42 0.560845
R263 source.n46 source.n44 0.560845
R264 source.n47 source.n46 0.560845
R265 source.n12 source.n11 0.470328
R266 source.n36 source.n35 0.470328
R267 source source.n48 0.188
R268 minus.n35 minus.t17 738.337
R269 minus.n8 minus.t9 738.337
R270 minus.n72 minus.t23 738.337
R271 minus.n43 minus.t6 738.337
R272 minus.n34 minus.t20 690.867
R273 minus.n32 minus.t21 690.867
R274 minus.n3 minus.t13 690.867
R275 minus.n26 minus.t16 690.867
R276 minus.n24 minus.t15 690.867
R277 minus.n6 minus.t18 690.867
R278 minus.n18 minus.t10 690.867
R279 minus.n16 minus.t11 690.867
R280 minus.n9 minus.t14 690.867
R281 minus.n10 minus.t8 690.867
R282 minus.n71 minus.t4 690.867
R283 minus.n69 minus.t7 690.867
R284 minus.n63 minus.t12 690.867
R285 minus.n62 minus.t0 690.867
R286 minus.n60 minus.t2 690.867
R287 minus.n54 minus.t3 690.867
R288 minus.n53 minus.t5 690.867
R289 minus.n51 minus.t19 690.867
R290 minus.n45 minus.t22 690.867
R291 minus.n44 minus.t1 690.867
R292 minus.n12 minus.n8 161.489
R293 minus.n47 minus.n43 161.489
R294 minus.n36 minus.n35 161.3
R295 minus.n33 minus.n0 161.3
R296 minus.n31 minus.n30 161.3
R297 minus.n29 minus.n1 161.3
R298 minus.n28 minus.n27 161.3
R299 minus.n25 minus.n2 161.3
R300 minus.n23 minus.n22 161.3
R301 minus.n21 minus.n4 161.3
R302 minus.n20 minus.n19 161.3
R303 minus.n17 minus.n5 161.3
R304 minus.n15 minus.n14 161.3
R305 minus.n13 minus.n7 161.3
R306 minus.n12 minus.n11 161.3
R307 minus.n73 minus.n72 161.3
R308 minus.n70 minus.n37 161.3
R309 minus.n68 minus.n67 161.3
R310 minus.n66 minus.n38 161.3
R311 minus.n65 minus.n64 161.3
R312 minus.n61 minus.n39 161.3
R313 minus.n59 minus.n58 161.3
R314 minus.n57 minus.n40 161.3
R315 minus.n56 minus.n55 161.3
R316 minus.n52 minus.n41 161.3
R317 minus.n50 minus.n49 161.3
R318 minus.n48 minus.n42 161.3
R319 minus.n47 minus.n46 161.3
R320 minus.n31 minus.n1 73.0308
R321 minus.n23 minus.n4 73.0308
R322 minus.n15 minus.n7 73.0308
R323 minus.n50 minus.n42 73.0308
R324 minus.n59 minus.n40 73.0308
R325 minus.n68 minus.n38 73.0308
R326 minus.n33 minus.n32 69.3793
R327 minus.n11 minus.n9 69.3793
R328 minus.n46 minus.n45 69.3793
R329 minus.n70 minus.n69 69.3793
R330 minus.n25 minus.n24 62.0763
R331 minus.n19 minus.n6 62.0763
R332 minus.n55 minus.n54 62.0763
R333 minus.n61 minus.n60 62.0763
R334 minus.n27 minus.n3 54.7732
R335 minus.n17 minus.n16 54.7732
R336 minus.n52 minus.n51 54.7732
R337 minus.n64 minus.n63 54.7732
R338 minus.n35 minus.n34 47.4702
R339 minus.n10 minus.n8 47.4702
R340 minus.n44 minus.n43 47.4702
R341 minus.n72 minus.n71 47.4702
R342 minus.n27 minus.n26 40.1672
R343 minus.n18 minus.n17 40.1672
R344 minus.n53 minus.n52 40.1672
R345 minus.n64 minus.n62 40.1672
R346 minus.n26 minus.n25 32.8641
R347 minus.n19 minus.n18 32.8641
R348 minus.n55 minus.n53 32.8641
R349 minus.n62 minus.n61 32.8641
R350 minus.n74 minus.n36 31.4399
R351 minus.n34 minus.n33 25.5611
R352 minus.n11 minus.n10 25.5611
R353 minus.n46 minus.n44 25.5611
R354 minus.n71 minus.n70 25.5611
R355 minus.n3 minus.n1 18.2581
R356 minus.n16 minus.n15 18.2581
R357 minus.n51 minus.n50 18.2581
R358 minus.n63 minus.n38 18.2581
R359 minus.n24 minus.n23 10.955
R360 minus.n6 minus.n4 10.955
R361 minus.n54 minus.n40 10.955
R362 minus.n60 minus.n59 10.955
R363 minus.n74 minus.n73 6.52323
R364 minus.n32 minus.n31 3.65202
R365 minus.n9 minus.n7 3.65202
R366 minus.n45 minus.n42 3.65202
R367 minus.n69 minus.n68 3.65202
R368 minus.n36 minus.n0 0.189894
R369 minus.n30 minus.n0 0.189894
R370 minus.n30 minus.n29 0.189894
R371 minus.n29 minus.n28 0.189894
R372 minus.n28 minus.n2 0.189894
R373 minus.n22 minus.n2 0.189894
R374 minus.n22 minus.n21 0.189894
R375 minus.n21 minus.n20 0.189894
R376 minus.n20 minus.n5 0.189894
R377 minus.n14 minus.n5 0.189894
R378 minus.n14 minus.n13 0.189894
R379 minus.n13 minus.n12 0.189894
R380 minus.n48 minus.n47 0.189894
R381 minus.n49 minus.n48 0.189894
R382 minus.n49 minus.n41 0.189894
R383 minus.n56 minus.n41 0.189894
R384 minus.n57 minus.n56 0.189894
R385 minus.n58 minus.n57 0.189894
R386 minus.n58 minus.n39 0.189894
R387 minus.n65 minus.n39 0.189894
R388 minus.n66 minus.n65 0.189894
R389 minus.n67 minus.n66 0.189894
R390 minus.n67 minus.n37 0.189894
R391 minus.n73 minus.n37 0.189894
R392 minus minus.n74 0.188
R393 drain_right.n13 drain_right.n11 80.3335
R394 drain_right.n7 drain_right.n5 80.3334
R395 drain_right.n2 drain_right.n0 80.3334
R396 drain_right.n13 drain_right.n12 79.7731
R397 drain_right.n15 drain_right.n14 79.7731
R398 drain_right.n17 drain_right.n16 79.7731
R399 drain_right.n19 drain_right.n18 79.7731
R400 drain_right.n21 drain_right.n20 79.7731
R401 drain_right.n7 drain_right.n6 79.773
R402 drain_right.n9 drain_right.n8 79.773
R403 drain_right.n4 drain_right.n3 79.773
R404 drain_right.n2 drain_right.n1 79.773
R405 drain_right drain_right.n10 25.3189
R406 drain_right.n5 drain_right.t19 10.0005
R407 drain_right.n5 drain_right.t0 10.0005
R408 drain_right.n6 drain_right.t11 10.0005
R409 drain_right.n6 drain_right.t16 10.0005
R410 drain_right.n8 drain_right.t21 10.0005
R411 drain_right.n8 drain_right.t23 10.0005
R412 drain_right.n3 drain_right.t18 10.0005
R413 drain_right.n3 drain_right.t20 10.0005
R414 drain_right.n1 drain_right.t1 10.0005
R415 drain_right.n1 drain_right.t4 10.0005
R416 drain_right.n0 drain_right.t17 10.0005
R417 drain_right.n0 drain_right.t22 10.0005
R418 drain_right.n11 drain_right.t15 10.0005
R419 drain_right.n11 drain_right.t14 10.0005
R420 drain_right.n12 drain_right.t12 10.0005
R421 drain_right.n12 drain_right.t9 10.0005
R422 drain_right.n14 drain_right.t5 10.0005
R423 drain_right.n14 drain_right.t13 10.0005
R424 drain_right.n16 drain_right.t7 10.0005
R425 drain_right.n16 drain_right.t8 10.0005
R426 drain_right.n18 drain_right.t2 10.0005
R427 drain_right.n18 drain_right.t10 10.0005
R428 drain_right.n20 drain_right.t6 10.0005
R429 drain_right.n20 drain_right.t3 10.0005
R430 drain_right drain_right.n21 6.21356
R431 drain_right.n9 drain_right.n7 0.560845
R432 drain_right.n4 drain_right.n2 0.560845
R433 drain_right.n21 drain_right.n19 0.560845
R434 drain_right.n19 drain_right.n17 0.560845
R435 drain_right.n17 drain_right.n15 0.560845
R436 drain_right.n15 drain_right.n13 0.560845
R437 drain_right.n10 drain_right.n9 0.225326
R438 drain_right.n10 drain_right.n4 0.225326
C0 drain_left plus 1.97368f
C1 plus drain_right 0.397886f
C2 drain_left drain_right 1.29455f
C3 plus minus 4.48207f
C4 drain_left minus 0.176743f
C5 drain_right minus 1.73594f
C6 plus source 1.86274f
C7 drain_left source 14.275201f
C8 drain_right source 14.2759f
C9 minus source 1.84874f
C10 drain_right a_n2406_n1488# 4.89066f
C11 drain_left a_n2406_n1488# 5.21728f
C12 source a_n2406_n1488# 4.040144f
C13 minus a_n2406_n1488# 8.177863f
C14 plus a_n2406_n1488# 8.941581f
C15 drain_right.t17 a_n2406_n1488# 0.090726f
C16 drain_right.t22 a_n2406_n1488# 0.090726f
C17 drain_right.n0 a_n2406_n1488# 0.495651f
C18 drain_right.t1 a_n2406_n1488# 0.090726f
C19 drain_right.t4 a_n2406_n1488# 0.090726f
C20 drain_right.n1 a_n2406_n1488# 0.493534f
C21 drain_right.n2 a_n2406_n1488# 0.594847f
C22 drain_right.t18 a_n2406_n1488# 0.090726f
C23 drain_right.t20 a_n2406_n1488# 0.090726f
C24 drain_right.n3 a_n2406_n1488# 0.493534f
C25 drain_right.n4 a_n2406_n1488# 0.268694f
C26 drain_right.t19 a_n2406_n1488# 0.090726f
C27 drain_right.t0 a_n2406_n1488# 0.090726f
C28 drain_right.n5 a_n2406_n1488# 0.495651f
C29 drain_right.t11 a_n2406_n1488# 0.090726f
C30 drain_right.t16 a_n2406_n1488# 0.090726f
C31 drain_right.n6 a_n2406_n1488# 0.493534f
C32 drain_right.n7 a_n2406_n1488# 0.594848f
C33 drain_right.t21 a_n2406_n1488# 0.090726f
C34 drain_right.t23 a_n2406_n1488# 0.090726f
C35 drain_right.n8 a_n2406_n1488# 0.493534f
C36 drain_right.n9 a_n2406_n1488# 0.268694f
C37 drain_right.n10 a_n2406_n1488# 0.856988f
C38 drain_right.t15 a_n2406_n1488# 0.090726f
C39 drain_right.t14 a_n2406_n1488# 0.090726f
C40 drain_right.n11 a_n2406_n1488# 0.495653f
C41 drain_right.t12 a_n2406_n1488# 0.090726f
C42 drain_right.t9 a_n2406_n1488# 0.090726f
C43 drain_right.n12 a_n2406_n1488# 0.493536f
C44 drain_right.n13 a_n2406_n1488# 0.594843f
C45 drain_right.t5 a_n2406_n1488# 0.090726f
C46 drain_right.t13 a_n2406_n1488# 0.090726f
C47 drain_right.n14 a_n2406_n1488# 0.493536f
C48 drain_right.n15 a_n2406_n1488# 0.293394f
C49 drain_right.t7 a_n2406_n1488# 0.090726f
C50 drain_right.t8 a_n2406_n1488# 0.090726f
C51 drain_right.n16 a_n2406_n1488# 0.493536f
C52 drain_right.n17 a_n2406_n1488# 0.293394f
C53 drain_right.t2 a_n2406_n1488# 0.090726f
C54 drain_right.t10 a_n2406_n1488# 0.090726f
C55 drain_right.n18 a_n2406_n1488# 0.493536f
C56 drain_right.n19 a_n2406_n1488# 0.293394f
C57 drain_right.t6 a_n2406_n1488# 0.090726f
C58 drain_right.t3 a_n2406_n1488# 0.090726f
C59 drain_right.n20 a_n2406_n1488# 0.493536f
C60 drain_right.n21 a_n2406_n1488# 0.504325f
C61 minus.n0 a_n2406_n1488# 0.02798f
C62 minus.t17 a_n2406_n1488# 0.038072f
C63 minus.t20 a_n2406_n1488# 0.036462f
C64 minus.t21 a_n2406_n1488# 0.036462f
C65 minus.n1 a_n2406_n1488# 0.011438f
C66 minus.n2 a_n2406_n1488# 0.02798f
C67 minus.t13 a_n2406_n1488# 0.036462f
C68 minus.n3 a_n2406_n1488# 0.025484f
C69 minus.t16 a_n2406_n1488# 0.036462f
C70 minus.t15 a_n2406_n1488# 0.036462f
C71 minus.n4 a_n2406_n1488# 0.010576f
C72 minus.n5 a_n2406_n1488# 0.02798f
C73 minus.t18 a_n2406_n1488# 0.036462f
C74 minus.n6 a_n2406_n1488# 0.025484f
C75 minus.t10 a_n2406_n1488# 0.036462f
C76 minus.t11 a_n2406_n1488# 0.036462f
C77 minus.n7 a_n2406_n1488# 0.009713f
C78 minus.t9 a_n2406_n1488# 0.038072f
C79 minus.n8 a_n2406_n1488# 0.03535f
C80 minus.t14 a_n2406_n1488# 0.036462f
C81 minus.n9 a_n2406_n1488# 0.025484f
C82 minus.t8 a_n2406_n1488# 0.036462f
C83 minus.n10 a_n2406_n1488# 0.025484f
C84 minus.n11 a_n2406_n1488# 0.011869f
C85 minus.n12 a_n2406_n1488# 0.061096f
C86 minus.n13 a_n2406_n1488# 0.02798f
C87 minus.n14 a_n2406_n1488# 0.02798f
C88 minus.n15 a_n2406_n1488# 0.011438f
C89 minus.n16 a_n2406_n1488# 0.025484f
C90 minus.n17 a_n2406_n1488# 0.011869f
C91 minus.n18 a_n2406_n1488# 0.025484f
C92 minus.n19 a_n2406_n1488# 0.011869f
C93 minus.n20 a_n2406_n1488# 0.02798f
C94 minus.n21 a_n2406_n1488# 0.02798f
C95 minus.n22 a_n2406_n1488# 0.02798f
C96 minus.n23 a_n2406_n1488# 0.010576f
C97 minus.n24 a_n2406_n1488# 0.025484f
C98 minus.n25 a_n2406_n1488# 0.011869f
C99 minus.n26 a_n2406_n1488# 0.025484f
C100 minus.n27 a_n2406_n1488# 0.011869f
C101 minus.n28 a_n2406_n1488# 0.02798f
C102 minus.n29 a_n2406_n1488# 0.02798f
C103 minus.n30 a_n2406_n1488# 0.02798f
C104 minus.n31 a_n2406_n1488# 0.009713f
C105 minus.n32 a_n2406_n1488# 0.025484f
C106 minus.n33 a_n2406_n1488# 0.011869f
C107 minus.n34 a_n2406_n1488# 0.025484f
C108 minus.n35 a_n2406_n1488# 0.035311f
C109 minus.n36 a_n2406_n1488# 0.788371f
C110 minus.n37 a_n2406_n1488# 0.02798f
C111 minus.t4 a_n2406_n1488# 0.036462f
C112 minus.t7 a_n2406_n1488# 0.036462f
C113 minus.n38 a_n2406_n1488# 0.011438f
C114 minus.n39 a_n2406_n1488# 0.02798f
C115 minus.t0 a_n2406_n1488# 0.036462f
C116 minus.t2 a_n2406_n1488# 0.036462f
C117 minus.n40 a_n2406_n1488# 0.010576f
C118 minus.n41 a_n2406_n1488# 0.02798f
C119 minus.t5 a_n2406_n1488# 0.036462f
C120 minus.t19 a_n2406_n1488# 0.036462f
C121 minus.n42 a_n2406_n1488# 0.009713f
C122 minus.t6 a_n2406_n1488# 0.038072f
C123 minus.n43 a_n2406_n1488# 0.03535f
C124 minus.t1 a_n2406_n1488# 0.036462f
C125 minus.n44 a_n2406_n1488# 0.025484f
C126 minus.t22 a_n2406_n1488# 0.036462f
C127 minus.n45 a_n2406_n1488# 0.025484f
C128 minus.n46 a_n2406_n1488# 0.011869f
C129 minus.n47 a_n2406_n1488# 0.061096f
C130 minus.n48 a_n2406_n1488# 0.02798f
C131 minus.n49 a_n2406_n1488# 0.02798f
C132 minus.n50 a_n2406_n1488# 0.011438f
C133 minus.n51 a_n2406_n1488# 0.025484f
C134 minus.n52 a_n2406_n1488# 0.011869f
C135 minus.n53 a_n2406_n1488# 0.025484f
C136 minus.t3 a_n2406_n1488# 0.036462f
C137 minus.n54 a_n2406_n1488# 0.025484f
C138 minus.n55 a_n2406_n1488# 0.011869f
C139 minus.n56 a_n2406_n1488# 0.02798f
C140 minus.n57 a_n2406_n1488# 0.02798f
C141 minus.n58 a_n2406_n1488# 0.02798f
C142 minus.n59 a_n2406_n1488# 0.010576f
C143 minus.n60 a_n2406_n1488# 0.025484f
C144 minus.n61 a_n2406_n1488# 0.011869f
C145 minus.n62 a_n2406_n1488# 0.025484f
C146 minus.t12 a_n2406_n1488# 0.036462f
C147 minus.n63 a_n2406_n1488# 0.025484f
C148 minus.n64 a_n2406_n1488# 0.011869f
C149 minus.n65 a_n2406_n1488# 0.02798f
C150 minus.n66 a_n2406_n1488# 0.02798f
C151 minus.n67 a_n2406_n1488# 0.02798f
C152 minus.n68 a_n2406_n1488# 0.009713f
C153 minus.n69 a_n2406_n1488# 0.025484f
C154 minus.n70 a_n2406_n1488# 0.011869f
C155 minus.n71 a_n2406_n1488# 0.025484f
C156 minus.t23 a_n2406_n1488# 0.038072f
C157 minus.n72 a_n2406_n1488# 0.035311f
C158 minus.n73 a_n2406_n1488# 0.184453f
C159 minus.n74 a_n2406_n1488# 0.969194f
C160 source.t25 a_n2406_n1488# 0.538322f
C161 source.n0 a_n2406_n1488# 0.710653f
C162 source.t33 a_n2406_n1488# 0.091399f
C163 source.t35 a_n2406_n1488# 0.091399f
C164 source.n1 a_n2406_n1488# 0.444638f
C165 source.n2 a_n2406_n1488# 0.31355f
C166 source.t37 a_n2406_n1488# 0.091399f
C167 source.t28 a_n2406_n1488# 0.091399f
C168 source.n3 a_n2406_n1488# 0.444638f
C169 source.n4 a_n2406_n1488# 0.31355f
C170 source.t27 a_n2406_n1488# 0.091399f
C171 source.t32 a_n2406_n1488# 0.091399f
C172 source.n5 a_n2406_n1488# 0.444638f
C173 source.n6 a_n2406_n1488# 0.31355f
C174 source.t34 a_n2406_n1488# 0.091399f
C175 source.t24 a_n2406_n1488# 0.091399f
C176 source.n7 a_n2406_n1488# 0.444638f
C177 source.n8 a_n2406_n1488# 0.31355f
C178 source.t26 a_n2406_n1488# 0.091399f
C179 source.t31 a_n2406_n1488# 0.091399f
C180 source.n9 a_n2406_n1488# 0.444638f
C181 source.n10 a_n2406_n1488# 0.31355f
C182 source.t36 a_n2406_n1488# 0.538322f
C183 source.n11 a_n2406_n1488# 0.376963f
C184 source.t15 a_n2406_n1488# 0.538322f
C185 source.n12 a_n2406_n1488# 0.376963f
C186 source.t2 a_n2406_n1488# 0.091399f
C187 source.t13 a_n2406_n1488# 0.091399f
C188 source.n13 a_n2406_n1488# 0.444638f
C189 source.n14 a_n2406_n1488# 0.31355f
C190 source.t7 a_n2406_n1488# 0.091399f
C191 source.t12 a_n2406_n1488# 0.091399f
C192 source.n15 a_n2406_n1488# 0.444638f
C193 source.n16 a_n2406_n1488# 0.31355f
C194 source.t9 a_n2406_n1488# 0.091399f
C195 source.t1 a_n2406_n1488# 0.091399f
C196 source.n17 a_n2406_n1488# 0.444638f
C197 source.n18 a_n2406_n1488# 0.31355f
C198 source.t21 a_n2406_n1488# 0.091399f
C199 source.t11 a_n2406_n1488# 0.091399f
C200 source.n19 a_n2406_n1488# 0.444638f
C201 source.n20 a_n2406_n1488# 0.31355f
C202 source.t18 a_n2406_n1488# 0.091399f
C203 source.t17 a_n2406_n1488# 0.091399f
C204 source.n21 a_n2406_n1488# 0.444638f
C205 source.n22 a_n2406_n1488# 0.31355f
C206 source.t3 a_n2406_n1488# 0.538322f
C207 source.n23 a_n2406_n1488# 0.976226f
C208 source.t29 a_n2406_n1488# 0.538319f
C209 source.n24 a_n2406_n1488# 0.976229f
C210 source.t46 a_n2406_n1488# 0.091399f
C211 source.t44 a_n2406_n1488# 0.091399f
C212 source.n25 a_n2406_n1488# 0.444635f
C213 source.n26 a_n2406_n1488# 0.313553f
C214 source.t40 a_n2406_n1488# 0.091399f
C215 source.t38 a_n2406_n1488# 0.091399f
C216 source.n27 a_n2406_n1488# 0.444635f
C217 source.n28 a_n2406_n1488# 0.313553f
C218 source.t30 a_n2406_n1488# 0.091399f
C219 source.t47 a_n2406_n1488# 0.091399f
C220 source.n29 a_n2406_n1488# 0.444635f
C221 source.n30 a_n2406_n1488# 0.313553f
C222 source.t42 a_n2406_n1488# 0.091399f
C223 source.t41 a_n2406_n1488# 0.091399f
C224 source.n31 a_n2406_n1488# 0.444635f
C225 source.n32 a_n2406_n1488# 0.313553f
C226 source.t39 a_n2406_n1488# 0.091399f
C227 source.t45 a_n2406_n1488# 0.091399f
C228 source.n33 a_n2406_n1488# 0.444635f
C229 source.n34 a_n2406_n1488# 0.313553f
C230 source.t43 a_n2406_n1488# 0.538319f
C231 source.n35 a_n2406_n1488# 0.376966f
C232 source.t19 a_n2406_n1488# 0.538319f
C233 source.n36 a_n2406_n1488# 0.376966f
C234 source.t0 a_n2406_n1488# 0.091399f
C235 source.t22 a_n2406_n1488# 0.091399f
C236 source.n37 a_n2406_n1488# 0.444635f
C237 source.n38 a_n2406_n1488# 0.313553f
C238 source.t5 a_n2406_n1488# 0.091399f
C239 source.t8 a_n2406_n1488# 0.091399f
C240 source.n39 a_n2406_n1488# 0.444635f
C241 source.n40 a_n2406_n1488# 0.313553f
C242 source.t10 a_n2406_n1488# 0.091399f
C243 source.t20 a_n2406_n1488# 0.091399f
C244 source.n41 a_n2406_n1488# 0.444635f
C245 source.n42 a_n2406_n1488# 0.313553f
C246 source.t6 a_n2406_n1488# 0.091399f
C247 source.t16 a_n2406_n1488# 0.091399f
C248 source.n43 a_n2406_n1488# 0.444635f
C249 source.n44 a_n2406_n1488# 0.313553f
C250 source.t23 a_n2406_n1488# 0.091399f
C251 source.t14 a_n2406_n1488# 0.091399f
C252 source.n45 a_n2406_n1488# 0.444635f
C253 source.n46 a_n2406_n1488# 0.313553f
C254 source.t4 a_n2406_n1488# 0.538319f
C255 source.n47 a_n2406_n1488# 0.521735f
C256 source.n48 a_n2406_n1488# 0.738166f
C257 drain_left.t20 a_n2406_n1488# 0.090103f
C258 drain_left.t0 a_n2406_n1488# 0.090103f
C259 drain_left.n0 a_n2406_n1488# 0.49225f
C260 drain_left.t23 a_n2406_n1488# 0.090103f
C261 drain_left.t6 a_n2406_n1488# 0.090103f
C262 drain_left.n1 a_n2406_n1488# 0.490147f
C263 drain_left.n2 a_n2406_n1488# 0.590766f
C264 drain_left.t8 a_n2406_n1488# 0.090103f
C265 drain_left.t16 a_n2406_n1488# 0.090103f
C266 drain_left.n3 a_n2406_n1488# 0.490147f
C267 drain_left.n4 a_n2406_n1488# 0.26685f
C268 drain_left.t1 a_n2406_n1488# 0.090103f
C269 drain_left.t3 a_n2406_n1488# 0.090103f
C270 drain_left.n5 a_n2406_n1488# 0.49225f
C271 drain_left.t5 a_n2406_n1488# 0.090103f
C272 drain_left.t7 a_n2406_n1488# 0.090103f
C273 drain_left.n6 a_n2406_n1488# 0.490147f
C274 drain_left.n7 a_n2406_n1488# 0.590766f
C275 drain_left.t2 a_n2406_n1488# 0.090103f
C276 drain_left.t4 a_n2406_n1488# 0.090103f
C277 drain_left.n8 a_n2406_n1488# 0.490147f
C278 drain_left.n9 a_n2406_n1488# 0.26685f
C279 drain_left.n10 a_n2406_n1488# 0.900471f
C280 drain_left.t10 a_n2406_n1488# 0.090103f
C281 drain_left.t22 a_n2406_n1488# 0.090103f
C282 drain_left.n11 a_n2406_n1488# 0.492252f
C283 drain_left.t15 a_n2406_n1488# 0.090103f
C284 drain_left.t12 a_n2406_n1488# 0.090103f
C285 drain_left.n12 a_n2406_n1488# 0.490149f
C286 drain_left.n13 a_n2406_n1488# 0.590761f
C287 drain_left.t19 a_n2406_n1488# 0.090103f
C288 drain_left.t17 a_n2406_n1488# 0.090103f
C289 drain_left.n14 a_n2406_n1488# 0.490149f
C290 drain_left.n15 a_n2406_n1488# 0.29138f
C291 drain_left.t14 a_n2406_n1488# 0.090103f
C292 drain_left.t9 a_n2406_n1488# 0.090103f
C293 drain_left.n16 a_n2406_n1488# 0.490149f
C294 drain_left.n17 a_n2406_n1488# 0.29138f
C295 drain_left.t21 a_n2406_n1488# 0.090103f
C296 drain_left.t13 a_n2406_n1488# 0.090103f
C297 drain_left.n18 a_n2406_n1488# 0.490149f
C298 drain_left.n19 a_n2406_n1488# 0.29138f
C299 drain_left.t11 a_n2406_n1488# 0.090103f
C300 drain_left.t18 a_n2406_n1488# 0.090103f
C301 drain_left.n20 a_n2406_n1488# 0.490149f
C302 drain_left.n21 a_n2406_n1488# 0.500864f
C303 plus.n0 a_n2406_n1488# 0.028336f
C304 plus.t12 a_n2406_n1488# 0.036926f
C305 plus.t14 a_n2406_n1488# 0.036926f
C306 plus.n1 a_n2406_n1488# 0.011584f
C307 plus.n2 a_n2406_n1488# 0.028336f
C308 plus.t10 a_n2406_n1488# 0.036926f
C309 plus.t15 a_n2406_n1488# 0.036926f
C310 plus.n3 a_n2406_n1488# 0.01071f
C311 plus.n4 a_n2406_n1488# 0.028336f
C312 plus.t23 a_n2406_n1488# 0.036926f
C313 plus.t13 a_n2406_n1488# 0.036926f
C314 plus.n5 a_n2406_n1488# 0.009837f
C315 plus.t11 a_n2406_n1488# 0.038557f
C316 plus.n6 a_n2406_n1488# 0.0358f
C317 plus.t21 a_n2406_n1488# 0.036926f
C318 plus.n7 a_n2406_n1488# 0.025809f
C319 plus.t16 a_n2406_n1488# 0.036926f
C320 plus.n8 a_n2406_n1488# 0.025809f
C321 plus.n9 a_n2406_n1488# 0.012021f
C322 plus.n10 a_n2406_n1488# 0.061874f
C323 plus.n11 a_n2406_n1488# 0.028336f
C324 plus.n12 a_n2406_n1488# 0.028336f
C325 plus.n13 a_n2406_n1488# 0.011584f
C326 plus.n14 a_n2406_n1488# 0.025809f
C327 plus.n15 a_n2406_n1488# 0.012021f
C328 plus.n16 a_n2406_n1488# 0.025809f
C329 plus.t20 a_n2406_n1488# 0.036926f
C330 plus.n17 a_n2406_n1488# 0.025809f
C331 plus.n18 a_n2406_n1488# 0.012021f
C332 plus.n19 a_n2406_n1488# 0.028336f
C333 plus.n20 a_n2406_n1488# 0.028336f
C334 plus.n21 a_n2406_n1488# 0.028336f
C335 plus.n22 a_n2406_n1488# 0.01071f
C336 plus.n23 a_n2406_n1488# 0.025809f
C337 plus.n24 a_n2406_n1488# 0.012021f
C338 plus.n25 a_n2406_n1488# 0.025809f
C339 plus.t19 a_n2406_n1488# 0.036926f
C340 plus.n26 a_n2406_n1488# 0.025809f
C341 plus.n27 a_n2406_n1488# 0.012021f
C342 plus.n28 a_n2406_n1488# 0.028336f
C343 plus.n29 a_n2406_n1488# 0.028336f
C344 plus.n30 a_n2406_n1488# 0.028336f
C345 plus.n31 a_n2406_n1488# 0.009837f
C346 plus.n32 a_n2406_n1488# 0.025809f
C347 plus.n33 a_n2406_n1488# 0.012021f
C348 plus.n34 a_n2406_n1488# 0.025809f
C349 plus.t22 a_n2406_n1488# 0.038557f
C350 plus.n35 a_n2406_n1488# 0.035761f
C351 plus.n36 a_n2406_n1488# 0.213297f
C352 plus.n37 a_n2406_n1488# 0.028336f
C353 plus.t18 a_n2406_n1488# 0.038557f
C354 plus.t1 a_n2406_n1488# 0.036926f
C355 plus.t3 a_n2406_n1488# 0.036926f
C356 plus.n38 a_n2406_n1488# 0.011584f
C357 plus.n39 a_n2406_n1488# 0.028336f
C358 plus.t7 a_n2406_n1488# 0.036926f
C359 plus.n40 a_n2406_n1488# 0.025809f
C360 plus.t9 a_n2406_n1488# 0.036926f
C361 plus.t17 a_n2406_n1488# 0.036926f
C362 plus.n41 a_n2406_n1488# 0.01071f
C363 plus.n42 a_n2406_n1488# 0.028336f
C364 plus.t0 a_n2406_n1488# 0.036926f
C365 plus.n43 a_n2406_n1488# 0.025809f
C366 plus.t5 a_n2406_n1488# 0.036926f
C367 plus.t6 a_n2406_n1488# 0.036926f
C368 plus.n44 a_n2406_n1488# 0.009837f
C369 plus.t4 a_n2406_n1488# 0.038557f
C370 plus.n45 a_n2406_n1488# 0.0358f
C371 plus.t8 a_n2406_n1488# 0.036926f
C372 plus.n46 a_n2406_n1488# 0.025809f
C373 plus.t2 a_n2406_n1488# 0.036926f
C374 plus.n47 a_n2406_n1488# 0.025809f
C375 plus.n48 a_n2406_n1488# 0.012021f
C376 plus.n49 a_n2406_n1488# 0.061874f
C377 plus.n50 a_n2406_n1488# 0.028336f
C378 plus.n51 a_n2406_n1488# 0.028336f
C379 plus.n52 a_n2406_n1488# 0.011584f
C380 plus.n53 a_n2406_n1488# 0.025809f
C381 plus.n54 a_n2406_n1488# 0.012021f
C382 plus.n55 a_n2406_n1488# 0.025809f
C383 plus.n56 a_n2406_n1488# 0.012021f
C384 plus.n57 a_n2406_n1488# 0.028336f
C385 plus.n58 a_n2406_n1488# 0.028336f
C386 plus.n59 a_n2406_n1488# 0.028336f
C387 plus.n60 a_n2406_n1488# 0.01071f
C388 plus.n61 a_n2406_n1488# 0.025809f
C389 plus.n62 a_n2406_n1488# 0.012021f
C390 plus.n63 a_n2406_n1488# 0.025809f
C391 plus.n64 a_n2406_n1488# 0.012021f
C392 plus.n65 a_n2406_n1488# 0.028336f
C393 plus.n66 a_n2406_n1488# 0.028336f
C394 plus.n67 a_n2406_n1488# 0.028336f
C395 plus.n68 a_n2406_n1488# 0.009837f
C396 plus.n69 a_n2406_n1488# 0.025809f
C397 plus.n70 a_n2406_n1488# 0.012021f
C398 plus.n71 a_n2406_n1488# 0.025809f
C399 plus.n72 a_n2406_n1488# 0.035761f
C400 plus.n73 a_n2406_n1488# 0.749436f
.ends

