* NGSPICE file created from opamp504.ext - technology: sky130A

.subckt opamp504 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n2804_13878.t29 a_n2982_13878.t33 a_n2982_13878.t34 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X1 CSoutput.t123 commonsourceibias.t80 gnd.t207 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X2 a_n2804_13878.t3 a_n2982_13878.t68 vdd.t249 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 vdd.t5 a_n8964_8799.t44 CSoutput.t2 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X4 gnd.t206 commonsourceibias.t81 CSoutput.t122 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X5 a_n8964_8799.t11 plus.t5 a_n2903_n3924.t20 gnd.t389 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X6 CSoutput.t121 commonsourceibias.t82 gnd.t205 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 CSoutput.t120 commonsourceibias.t83 gnd.t204 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 CSoutput.t3 a_n8964_8799.t45 vdd.t7 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X9 a_n2903_n3924.t19 plus.t6 a_n8964_8799.t0 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X10 gnd.t203 commonsourceibias.t84 CSoutput.t119 gnd.t124 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 CSoutput.t216 a_n2982_8322.t5 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X12 vdd.t181 a_n8964_8799.t46 CSoutput.t180 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X13 a_n2982_8322.t29 a_n2982_13878.t69 a_n8964_8799.t36 vdd.t246 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X14 CSoutput.t181 a_n8964_8799.t47 vdd.t183 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X15 vdd.t258 a_n8964_8799.t48 CSoutput.t198 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X16 vdd.t157 CSoutput.t217 output.t15 gnd.t373 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X17 CSoutput.t199 a_n8964_8799.t49 vdd.t259 vdd.t63 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X18 CSoutput.t118 commonsourceibias.t85 gnd.t197 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 gnd.t202 commonsourceibias.t86 CSoutput.t117 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 CSoutput.t116 commonsourceibias.t87 gnd.t198 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X21 gnd.t201 commonsourceibias.t88 CSoutput.t115 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X22 vdd.t50 a_n8964_8799.t50 CSoutput.t144 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X23 vdd.t52 a_n8964_8799.t51 CSoutput.t145 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X24 CSoutput.t114 commonsourceibias.t89 gnd.t200 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 CSoutput.t113 commonsourceibias.t90 gnd.t199 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 gnd.t196 commonsourceibias.t91 CSoutput.t112 gnd.t85 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 gnd.t340 gnd.t337 gnd.t339 gnd.t338 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X28 gnd.t336 gnd.t334 gnd.t335 gnd.t238 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X29 commonsourceibias.t13 commonsourceibias.t12 gnd.t195 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X30 a_n2982_13878.t16 minus.t5 a_n2903_n3924.t42 gnd.t388 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X31 CSoutput.t111 commonsourceibias.t92 gnd.t194 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 gnd.t333 gnd.t331 gnd.t332 gnd.t230 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X33 a_n8964_8799.t42 plus.t7 a_n2903_n3924.t18 gnd.t387 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X34 a_n8964_8799.t35 a_n2982_13878.t70 a_n2982_8322.t28 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X35 vdd.t170 a_n8964_8799.t52 CSoutput.t172 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X36 a_n2982_13878.t4 minus.t6 a_n2903_n3924.t25 gnd.t347 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X37 vdd.t172 a_n8964_8799.t53 CSoutput.t173 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X38 a_n8964_8799.t34 a_n2982_13878.t71 a_n2982_8322.t27 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X39 CSoutput.t110 commonsourceibias.t93 gnd.t193 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 gnd.t192 commonsourceibias.t94 CSoutput.t109 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X41 gnd.t330 gnd.t328 gnd.t329 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X42 CSoutput.t108 commonsourceibias.t95 gnd.t191 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 CSoutput.t107 commonsourceibias.t96 gnd.t190 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X44 CSoutput.t106 commonsourceibias.t97 gnd.t189 gnd.t87 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X45 a_n2903_n3924.t17 plus.t8 a_n8964_8799.t39 gnd.t364 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X46 a_n2903_n3924.t35 diffpairibias.t16 gnd.t369 gnd.t368 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X47 gnd.t188 commonsourceibias.t98 CSoutput.t105 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X48 a_n2903_n3924.t28 minus.t7 a_n2982_13878.t6 gnd.t353 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X49 CSoutput.t188 a_n8964_8799.t54 vdd.t190 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X50 gnd.t187 commonsourceibias.t99 CSoutput.t104 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 CSoutput.t103 commonsourceibias.t100 gnd.t186 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 vdd.t191 a_n8964_8799.t55 CSoutput.t189 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 CSoutput.t102 commonsourceibias.t101 gnd.t185 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X54 gnd.t175 commonsourceibias.t0 commonsourceibias.t1 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 CSoutput.t101 commonsourceibias.t102 gnd.t177 gnd.t87 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 gnd.t176 commonsourceibias.t103 CSoutput.t100 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X57 vdd.t266 a_n8964_8799.t56 CSoutput.t206 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X58 a_n2804_13878.t28 a_n2982_13878.t47 a_n2982_13878.t48 vdd.t203 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X59 CSoutput.t99 commonsourceibias.t104 gnd.t178 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X60 CSoutput.t98 commonsourceibias.t105 gnd.t184 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X61 gnd.t183 commonsourceibias.t106 CSoutput.t97 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X62 vdd.t158 CSoutput.t218 output.t14 gnd.t374 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X63 a_n2982_13878.t44 a_n2982_13878.t43 a_n2804_13878.t27 vdd.t216 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X64 CSoutput.t96 commonsourceibias.t107 gnd.t182 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X65 gnd.t181 commonsourceibias.t108 CSoutput.t95 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X66 CSoutput.t207 a_n8964_8799.t57 vdd.t267 vdd.t63 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X67 CSoutput.t219 a_n2982_8322.t4 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X68 vdd.t140 vdd.t138 vdd.t139 vdd.t115 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X69 gnd.t180 commonsourceibias.t2 commonsourceibias.t3 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 vdd.t272 a_n8964_8799.t58 CSoutput.t212 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 CSoutput.t94 commonsourceibias.t109 gnd.t179 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X72 a_n2903_n3924.t16 plus.t9 a_n8964_8799.t4 gnd.t351 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X73 vdd.t273 a_n8964_8799.t59 CSoutput.t213 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X74 gnd.t327 gnd.t325 gnd.t326 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X75 CSoutput.t93 commonsourceibias.t110 gnd.t174 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 plus.t4 gnd.t322 gnd.t324 gnd.t323 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X77 diffpairibias.t15 diffpairibias.t14 gnd.t399 gnd.t398 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X78 a_n2903_n3924.t15 plus.t10 a_n8964_8799.t43 gnd.t365 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X79 gnd.t321 gnd.t319 gnd.t320 gnd.t265 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X80 gnd.t173 commonsourceibias.t111 CSoutput.t92 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X81 a_n2982_13878.t36 a_n2982_13878.t35 a_n2804_13878.t26 vdd.t231 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X82 CSoutput.t91 commonsourceibias.t112 gnd.t172 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X83 CSoutput.t166 a_n8964_8799.t60 vdd.t162 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X84 CSoutput.t90 commonsourceibias.t113 gnd.t171 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 gnd.t170 commonsourceibias.t114 CSoutput.t89 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X86 a_n8964_8799.t33 a_n2982_13878.t72 a_n2982_8322.t26 vdd.t226 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X87 gnd.t169 commonsourceibias.t115 CSoutput.t88 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 vdd.t163 a_n8964_8799.t61 CSoutput.t167 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X89 CSoutput.t178 a_n8964_8799.t62 vdd.t178 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X90 gnd.t162 commonsourceibias.t116 CSoutput.t87 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 a_n2982_13878.t22 a_n2982_13878.t21 a_n2804_13878.t25 vdd.t247 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X92 vdd.t179 a_n8964_8799.t63 CSoutput.t179 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X93 vdd.t34 a_n8964_8799.t64 CSoutput.t134 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X94 a_n8964_8799.t28 a_n2982_13878.t73 a_n2982_8322.t25 vdd.t224 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X95 CSoutput.t86 commonsourceibias.t117 gnd.t163 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X96 diffpairibias.t13 diffpairibias.t12 gnd.t355 gnd.t354 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X97 CSoutput.t135 a_n8964_8799.t65 vdd.t35 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X98 gnd.t168 commonsourceibias.t34 commonsourceibias.t35 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X99 gnd.t167 commonsourceibias.t118 CSoutput.t85 gnd.t85 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X100 a_n8964_8799.t27 a_n2982_13878.t74 a_n2982_8322.t24 vdd.t239 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X101 CSoutput.t84 commonsourceibias.t119 gnd.t166 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X102 gnd.t165 commonsourceibias.t120 CSoutput.t83 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X103 CSoutput.t82 commonsourceibias.t121 gnd.t164 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 CSoutput.t81 commonsourceibias.t122 gnd.t161 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X105 a_n2982_8322.t23 a_n2982_13878.t75 a_n8964_8799.t30 vdd.t247 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X106 CSoutput.t80 commonsourceibias.t123 gnd.t160 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X107 gnd.t159 commonsourceibias.t124 CSoutput.t79 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 CSoutput.t162 a_n8964_8799.t66 vdd.t155 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X109 a_n2903_n3924.t0 minus.t8 a_n2982_13878.t0 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X110 gnd.t158 commonsourceibias.t78 commonsourceibias.t79 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X111 a_n2903_n3924.t14 plus.t11 a_n8964_8799.t6 gnd.t346 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X112 gnd.t157 commonsourceibias.t76 commonsourceibias.t77 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X113 CSoutput.t78 commonsourceibias.t125 gnd.t156 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X114 vdd.t173 CSoutput.t220 output.t13 gnd.t381 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X115 gnd.t318 gnd.t316 gnd.t317 gnd.t234 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X116 a_n8964_8799.t3 plus.t12 a_n2903_n3924.t13 gnd.t348 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X117 gnd.t315 gnd.t313 minus.t4 gnd.t314 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X118 output.t12 CSoutput.t221 vdd.t8 gnd.t3 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X119 CSoutput.t77 commonsourceibias.t126 gnd.t155 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 gnd.t154 commonsourceibias.t127 CSoutput.t76 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X121 vdd.t137 vdd.t135 vdd.t136 vdd.t111 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X122 a_n2903_n3924.t26 diffpairibias.t17 gnd.t350 gnd.t349 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X123 CSoutput.t222 a_n2982_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X124 vdd.t156 a_n8964_8799.t67 CSoutput.t163 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X125 gnd.t312 gnd.t310 gnd.t311 gnd.t226 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X126 vdd.t264 a_n8964_8799.t68 CSoutput.t204 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X127 a_n2982_13878.t46 a_n2982_13878.t45 a_n2804_13878.t24 vdd.t246 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X128 vdd.t265 a_n8964_8799.t69 CSoutput.t205 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X129 a_n2903_n3924.t12 plus.t13 a_n8964_8799.t2 gnd.t342 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X130 gnd.t153 commonsourceibias.t128 CSoutput.t75 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X131 gnd.t309 gnd.t306 gnd.t308 gnd.t307 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X132 a_n8964_8799.t29 a_n2982_13878.t76 a_n2982_8322.t22 vdd.t235 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X133 a_n2982_13878.t50 a_n2982_13878.t49 a_n2804_13878.t23 vdd.t198 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X134 gnd.t305 gnd.t303 gnd.t304 gnd.t226 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X135 gnd.t152 commonsourceibias.t129 CSoutput.t74 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X136 CSoutput.t73 commonsourceibias.t130 gnd.t149 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X137 commonsourceibias.t75 commonsourceibias.t74 gnd.t151 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 CSoutput.t210 a_n8964_8799.t70 vdd.t270 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X139 gnd.t150 commonsourceibias.t131 CSoutput.t72 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X140 gnd.t148 commonsourceibias.t132 CSoutput.t71 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X141 vdd.t134 vdd.t132 vdd.t133 vdd.t122 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X142 gnd.t147 commonsourceibias.t72 commonsourceibias.t73 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X143 CSoutput.t211 a_n8964_8799.t71 vdd.t271 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X144 gnd.t146 commonsourceibias.t133 CSoutput.t70 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X145 vdd.t131 vdd.t128 vdd.t130 vdd.t129 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X146 a_n2804_13878.t22 a_n2982_13878.t29 a_n2982_13878.t30 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X147 CSoutput.t154 a_n8964_8799.t72 vdd.t145 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X148 gnd.t302 gnd.t300 gnd.t301 gnd.t230 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X149 vdd.t147 a_n8964_8799.t73 CSoutput.t155 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X150 vdd.t245 a_n2982_13878.t77 a_n2982_8322.t37 vdd.t244 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X151 a_n2982_13878.t26 a_n2982_13878.t25 a_n2804_13878.t21 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X152 CSoutput.t69 commonsourceibias.t134 gnd.t123 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X153 a_n2982_8322.t36 a_n2982_13878.t78 vdd.t243 vdd.t242 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X154 CSoutput.t160 a_n8964_8799.t74 vdd.t153 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X155 gnd.t145 commonsourceibias.t135 CSoutput.t68 gnd.t85 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X156 a_n2903_n3924.t23 diffpairibias.t18 gnd.t345 gnd.t344 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X157 output.t11 CSoutput.t223 vdd.t9 gnd.t4 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X158 vdd.t10 CSoutput.t224 output.t10 gnd.t5 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X159 gnd.t144 commonsourceibias.t136 CSoutput.t67 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X160 gnd.t126 commonsourceibias.t6 commonsourceibias.t7 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 CSoutput.t66 commonsourceibias.t137 gnd.t143 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X162 gnd.t142 commonsourceibias.t138 CSoutput.t65 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X163 CSoutput.t64 commonsourceibias.t139 gnd.t141 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X164 CSoutput.t63 commonsourceibias.t140 gnd.t140 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X165 CSoutput.t62 commonsourceibias.t141 gnd.t139 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X166 vdd.t241 a_n2982_13878.t79 a_n2804_13878.t30 vdd.t240 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X167 vdd.t127 vdd.t125 vdd.t126 vdd.t111 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X168 vdd.t124 vdd.t121 vdd.t123 vdd.t122 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X169 vdd.t154 a_n8964_8799.t75 CSoutput.t161 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X170 vdd.t13 CSoutput.t225 output.t9 gnd.t208 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X171 gnd.t296 gnd.t294 gnd.t295 gnd.t226 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X172 a_n2804_13878.t20 a_n2982_13878.t23 a_n2982_13878.t24 vdd.t239 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X173 plus.t3 gnd.t297 gnd.t299 gnd.t298 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X174 vdd.t256 a_n8964_8799.t76 CSoutput.t196 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X175 a_n2982_8322.t21 a_n2982_13878.t80 a_n8964_8799.t32 vdd.t225 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X176 gnd.t293 gnd.t291 minus.t3 gnd.t292 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X177 a_n8964_8799.t9 plus.t14 a_n2903_n3924.t11 gnd.t386 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X178 vdd.t120 vdd.t118 vdd.t119 vdd.t88 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X179 a_n2982_13878.t11 minus.t9 a_n2903_n3924.t36 gnd.t372 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X180 vdd.t117 vdd.t114 vdd.t116 vdd.t115 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X181 a_n2982_8322.t35 a_n2982_13878.t81 vdd.t238 vdd.t237 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X182 a_n8964_8799.t31 a_n2982_13878.t82 a_n2982_8322.t20 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X183 a_n8964_8799.t5 plus.t15 a_n2903_n3924.t10 gnd.t360 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X184 CSoutput.t197 a_n8964_8799.t77 vdd.t257 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X185 diffpairibias.t11 diffpairibias.t10 gnd.t211 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X186 vdd.t252 a_n8964_8799.t78 CSoutput.t192 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X187 a_n2982_13878.t54 a_n2982_13878.t53 a_n2804_13878.t19 vdd.t219 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X188 CSoutput.t61 commonsourceibias.t142 gnd.t138 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 a_n8964_8799.t16 a_n2982_13878.t83 a_n2982_8322.t19 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X190 CSoutput.t193 a_n8964_8799.t79 vdd.t253 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X191 CSoutput.t132 a_n8964_8799.t80 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X192 commonsourceibias.t11 commonsourceibias.t10 gnd.t137 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 output.t8 CSoutput.t226 vdd.t14 gnd.t209 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X194 gnd.t122 commonsourceibias.t143 CSoutput.t60 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 a_n2804_13878.t18 a_n2982_13878.t37 a_n2982_13878.t38 vdd.t235 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X196 gnd.t125 commonsourceibias.t4 commonsourceibias.t5 gnd.t124 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X197 CSoutput.t59 commonsourceibias.t144 gnd.t136 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X198 vdd.t113 vdd.t110 vdd.t112 vdd.t111 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X199 vdd.t109 vdd.t107 vdd.t108 vdd.t84 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X200 vdd.t106 vdd.t104 vdd.t105 vdd.t70 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X201 CSoutput.t133 a_n8964_8799.t81 vdd.t32 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X202 gnd.t290 gnd.t288 minus.t2 gnd.t289 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X203 output.t7 CSoutput.t227 vdd.t11 gnd.t6 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X204 CSoutput.t58 commonsourceibias.t145 gnd.t135 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X205 vdd.t234 a_n2982_13878.t84 a_n2982_8322.t34 vdd.t233 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X206 a_n2804_13878.t17 a_n2982_13878.t41 a_n2982_13878.t42 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X207 vdd.t46 a_n8964_8799.t82 CSoutput.t142 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X208 vdd.t48 a_n8964_8799.t83 CSoutput.t143 vdd.t47 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X209 gnd.t134 commonsourceibias.t146 CSoutput.t57 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 gnd.t133 commonsourceibias.t147 CSoutput.t56 gnd.t124 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X211 a_n2982_13878.t66 minus.t10 a_n2903_n3924.t45 gnd.t389 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X212 a_n2903_n3924.t9 plus.t16 a_n8964_8799.t40 gnd.t343 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X213 a_n2982_13878.t28 a_n2982_13878.t27 a_n2804_13878.t16 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X214 gnd.t132 commonsourceibias.t148 CSoutput.t55 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 gnd.t131 commonsourceibias.t149 CSoutput.t54 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X216 commonsourceibias.t9 commonsourceibias.t8 gnd.t130 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X217 gnd.t128 commonsourceibias.t150 CSoutput.t53 gnd.t124 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 gnd.t287 gnd.t285 gnd.t286 gnd.t238 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X219 gnd.t127 commonsourceibias.t151 CSoutput.t52 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X220 vdd.t167 a_n8964_8799.t84 CSoutput.t170 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X221 CSoutput.t51 commonsourceibias.t152 gnd.t121 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X222 a_n2903_n3924.t37 diffpairibias.t19 gnd.t385 gnd.t384 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X223 gnd.t284 gnd.t281 gnd.t283 gnd.t282 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X224 a_n2903_n3924.t46 diffpairibias.t20 gnd.t403 gnd.t402 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X225 commonsourceibias.t31 commonsourceibias.t30 gnd.t120 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 a_n8964_8799.t37 plus.t17 a_n2903_n3924.t8 gnd.t352 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X227 vdd.t168 a_n8964_8799.t85 CSoutput.t171 vdd.t47 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X228 vdd.t159 a_n8964_8799.t86 CSoutput.t164 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 CSoutput.t165 a_n8964_8799.t87 vdd.t160 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X230 gnd.t280 gnd.t278 gnd.t279 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X231 vdd.t103 vdd.t101 vdd.t102 vdd.t88 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X232 CSoutput.t50 commonsourceibias.t153 gnd.t118 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X233 a_n8964_8799.t41 plus.t18 a_n2903_n3924.t7 gnd.t347 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X234 CSoutput.t49 commonsourceibias.t154 gnd.t117 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 a_n2804_13878.t15 a_n2982_13878.t63 a_n2982_13878.t64 vdd.t207 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X236 CSoutput.t186 a_n8964_8799.t88 vdd.t188 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X237 commonsourceibias.t29 commonsourceibias.t28 gnd.t116 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X238 gnd.t277 gnd.t274 gnd.t276 gnd.t275 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X239 a_n2982_8322.t18 a_n2982_13878.t85 a_n8964_8799.t15 vdd.t231 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X240 output.t18 outputibias.t8 gnd.t397 gnd.t396 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X241 CSoutput.t187 a_n8964_8799.t89 vdd.t189 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X242 CSoutput.t48 commonsourceibias.t155 gnd.t115 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 commonsourceibias.t27 commonsourceibias.t26 gnd.t113 gnd.t87 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X244 CSoutput.t47 commonsourceibias.t156 gnd.t112 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X245 outputibias.t7 outputibias.t6 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X246 gnd.t111 commonsourceibias.t46 commonsourceibias.t47 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X247 vdd.t12 CSoutput.t228 output.t6 gnd.t7 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X248 diffpairibias.t9 diffpairibias.t8 gnd.t391 gnd.t390 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X249 a_n2804_13878.t31 a_n2982_13878.t86 vdd.t230 vdd.t229 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X250 output.t19 outputibias.t9 gnd.t401 gnd.t400 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X251 a_n2982_13878.t7 minus.t11 a_n2903_n3924.t30 gnd.t341 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X252 vdd.t228 a_n2982_13878.t87 a_n2804_13878.t4 vdd.t227 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X253 CSoutput.t46 commonsourceibias.t157 gnd.t108 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 CSoutput.t45 commonsourceibias.t158 gnd.t109 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X255 CSoutput.t176 a_n8964_8799.t90 vdd.t176 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X256 CSoutput.t44 commonsourceibias.t159 gnd.t107 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X257 gnd.t106 commonsourceibias.t44 commonsourceibias.t45 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X258 a_n2903_n3924.t6 plus.t19 a_n8964_8799.t38 gnd.t353 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X259 vdd.t177 a_n8964_8799.t91 CSoutput.t177 vdd.t47 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X260 vdd.t26 a_n8964_8799.t92 CSoutput.t130 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X261 outputibias.t5 outputibias.t4 gnd.t215 gnd.t214 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X262 vdd.t28 a_n8964_8799.t93 CSoutput.t131 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X263 commonsourceibias.t37 commonsourceibias.t36 gnd.t99 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 gnd.t104 commonsourceibias.t160 CSoutput.t43 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X265 CSoutput.t0 a_n8964_8799.t94 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X266 a_n2804_13878.t14 a_n2982_13878.t57 a_n2982_13878.t58 vdd.t226 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X267 gnd.t103 commonsourceibias.t42 commonsourceibias.t43 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X268 gnd.t102 commonsourceibias.t161 CSoutput.t42 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 commonsourceibias.t41 commonsourceibias.t40 gnd.t101 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X270 vdd.t3 a_n8964_8799.t95 CSoutput.t1 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X271 gnd.t100 commonsourceibias.t38 commonsourceibias.t39 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X272 a_n2903_n3924.t31 minus.t12 a_n2982_13878.t8 gnd.t361 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X273 a_n2982_8322.t17 a_n2982_13878.t88 a_n8964_8799.t18 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X274 a_n2982_13878.t20 a_n2982_13878.t19 a_n2804_13878.t13 vdd.t225 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X275 CSoutput.t41 commonsourceibias.t162 gnd.t97 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X276 CSoutput.t174 a_n8964_8799.t96 vdd.t174 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X277 diffpairibias.t7 diffpairibias.t6 gnd.t376 gnd.t375 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X278 vdd.t175 a_n8964_8799.t97 CSoutput.t175 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X279 a_n2804_13878.t12 a_n2982_13878.t55 a_n2982_13878.t56 vdd.t224 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X280 commonsourceibias.t25 commonsourceibias.t24 gnd.t84 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X281 gnd.t273 gnd.t271 gnd.t272 gnd.t238 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X282 vdd.t223 a_n2982_13878.t89 a_n2982_8322.t33 vdd.t222 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X283 vdd.t142 a_n8964_8799.t98 CSoutput.t152 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X284 a_n2903_n3924.t33 minus.t13 a_n2982_13878.t10 gnd.t365 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X285 gnd.t267 gnd.t264 gnd.t266 gnd.t265 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X286 gnd.t96 commonsourceibias.t163 CSoutput.t40 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 gnd.t270 gnd.t268 plus.t2 gnd.t269 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X288 a_n2903_n3924.t21 minus.t14 a_n2982_13878.t1 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X289 CSoutput.t153 a_n8964_8799.t99 vdd.t144 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X290 minus.t1 gnd.t261 gnd.t263 gnd.t262 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X291 gnd.t95 commonsourceibias.t54 commonsourceibias.t55 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 CSoutput.t39 commonsourceibias.t164 gnd.t93 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X293 a_n2804_13878.t5 a_n2982_13878.t90 vdd.t221 vdd.t220 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X294 vdd.t100 vdd.t98 vdd.t99 vdd.t84 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X295 vdd.t254 a_n8964_8799.t100 CSoutput.t194 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X296 output.t5 CSoutput.t229 vdd.t40 gnd.t220 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X297 CSoutput.t195 a_n8964_8799.t101 vdd.t255 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X298 CSoutput.t190 a_n8964_8799.t102 vdd.t250 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X299 gnd.t92 commonsourceibias.t165 CSoutput.t38 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X300 vdd.t251 a_n8964_8799.t103 CSoutput.t191 vdd.t61 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 gnd.t260 gnd.t257 gnd.t259 gnd.t258 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X302 vdd.t97 vdd.t95 vdd.t96 vdd.t74 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X303 a_n2903_n3924.t34 diffpairibias.t21 gnd.t367 gnd.t366 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X304 a_n2982_8322.t16 a_n2982_13878.t91 a_n8964_8799.t17 vdd.t219 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X305 vdd.t218 a_n2982_13878.t92 a_n2982_8322.t32 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X306 CSoutput.t230 a_n2982_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X307 gnd.t91 commonsourceibias.t52 commonsourceibias.t53 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X308 a_n8964_8799.t10 plus.t20 a_n2903_n3924.t5 gnd.t388 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X309 outputibias.t3 outputibias.t2 gnd.t383 gnd.t382 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X310 a_n2982_13878.t14 minus.t15 a_n2903_n3924.t40 gnd.t387 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X311 vdd.t44 a_n8964_8799.t104 CSoutput.t140 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X312 a_n2903_n3924.t24 minus.t16 a_n2982_13878.t3 gnd.t346 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X313 output.t17 outputibias.t10 gnd.t378 gnd.t377 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X314 gnd.t89 commonsourceibias.t50 commonsourceibias.t51 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 vdd.t94 vdd.t91 vdd.t93 vdd.t92 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X316 CSoutput.t37 commonsourceibias.t166 gnd.t90 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X317 a_n2903_n3924.t41 minus.t17 a_n2982_13878.t15 gnd.t342 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X318 vdd.t45 a_n8964_8799.t105 CSoutput.t141 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 gnd.t256 gnd.t254 gnd.t255 gnd.t230 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X320 vdd.t36 CSoutput.t231 output.t4 gnd.t219 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X321 CSoutput.t168 a_n8964_8799.t106 vdd.t164 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 CSoutput.t36 commonsourceibias.t167 gnd.t88 gnd.t87 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X323 CSoutput.t169 a_n8964_8799.t107 vdd.t166 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X324 CSoutput.t184 a_n8964_8799.t108 vdd.t186 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 a_n2903_n3924.t32 minus.t18 a_n2982_13878.t9 gnd.t364 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X326 a_n2804_13878.t11 a_n2982_13878.t59 a_n2982_13878.t60 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X327 a_n2982_8322.t15 a_n2982_13878.t93 a_n8964_8799.t20 vdd.t216 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X328 diffpairibias.t5 diffpairibias.t4 gnd.t213 gnd.t212 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X329 CSoutput.t232 a_n2982_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X330 gnd.t253 gnd.t250 gnd.t252 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X331 CSoutput.t185 a_n8964_8799.t109 vdd.t187 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X332 CSoutput.t136 a_n8964_8799.t110 vdd.t38 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X333 gnd.t86 commonsourceibias.t48 commonsourceibias.t49 gnd.t85 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X334 output.t3 CSoutput.t233 vdd.t59 gnd.t358 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X335 vdd.t90 vdd.t87 vdd.t89 vdd.t88 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X336 vdd.t86 vdd.t83 vdd.t85 vdd.t84 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X337 CSoutput.t35 commonsourceibias.t168 gnd.t83 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X338 commonsourceibias.t23 commonsourceibias.t22 gnd.t81 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X339 gnd.t249 gnd.t247 plus.t1 gnd.t248 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X340 a_n2982_8322.t31 a_n2982_13878.t94 vdd.t215 vdd.t214 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X341 CSoutput.t137 a_n8964_8799.t111 vdd.t39 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X342 a_n2903_n3924.t44 minus.t19 a_n2982_13878.t65 gnd.t351 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X343 vdd.t268 a_n8964_8799.t112 CSoutput.t208 vdd.t61 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X344 gnd.t80 commonsourceibias.t169 CSoutput.t34 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X345 CSoutput.t209 a_n8964_8799.t113 vdd.t269 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X346 vdd.t213 a_n2982_13878.t95 a_n2804_13878.t2 vdd.t212 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X347 vdd.t62 a_n8964_8799.t114 CSoutput.t150 vdd.t61 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X348 CSoutput.t151 a_n8964_8799.t115 vdd.t64 vdd.t63 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X349 vdd.t262 a_n8964_8799.t116 CSoutput.t202 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X350 gnd.t79 commonsourceibias.t170 CSoutput.t33 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X351 gnd.t78 commonsourceibias.t171 CSoutput.t32 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X352 output.t2 CSoutput.t234 vdd.t60 gnd.t359 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X353 a_n2982_8322.t14 a_n2982_13878.t96 a_n8964_8799.t19 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X354 commonsourceibias.t21 commonsourceibias.t20 gnd.t77 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X355 a_n8964_8799.t26 a_n2982_13878.t97 a_n2982_8322.t13 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X356 a_n2804_13878.t1 a_n2982_13878.t98 vdd.t210 vdd.t209 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X357 gnd.t75 commonsourceibias.t172 CSoutput.t31 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X358 vdd.t82 vdd.t80 vdd.t81 vdd.t66 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X359 vdd.t263 a_n8964_8799.t117 CSoutput.t203 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X360 CSoutput.t182 a_n8964_8799.t118 vdd.t184 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X361 CSoutput.t183 a_n8964_8799.t119 vdd.t185 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X362 CSoutput.t148 a_n8964_8799.t120 vdd.t57 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X363 commonsourceibias.t19 commonsourceibias.t18 gnd.t74 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X364 a_n2982_13878.t18 a_n2982_13878.t17 a_n2804_13878.t10 vdd.t199 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X365 gnd.t246 gnd.t244 plus.t0 gnd.t245 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X366 a_n8964_8799.t25 a_n2982_13878.t99 a_n2982_8322.t12 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X367 a_n2903_n3924.t4 plus.t21 a_n8964_8799.t8 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X368 minus.t0 gnd.t241 gnd.t243 gnd.t242 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X369 output.t1 CSoutput.t235 vdd.t192 gnd.t394 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X370 a_n8964_8799.t14 a_n2982_13878.t100 a_n2982_8322.t11 vdd.t207 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X371 a_n2982_13878.t12 minus.t20 a_n2903_n3924.t38 gnd.t360 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X372 gnd.t240 gnd.t237 gnd.t239 gnd.t238 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X373 gnd.t72 commonsourceibias.t173 CSoutput.t30 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X374 a_n2982_8322.t10 a_n2982_13878.t101 a_n8964_8799.t13 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X375 commonsourceibias.t71 commonsourceibias.t70 gnd.t71 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X376 gnd.t69 commonsourceibias.t174 CSoutput.t29 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X377 gnd.t236 gnd.t233 gnd.t235 gnd.t234 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X378 a_n2982_13878.t67 minus.t21 a_n2903_n3924.t47 gnd.t348 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X379 CSoutput.t28 commonsourceibias.t175 gnd.t67 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X380 vdd.t58 a_n8964_8799.t121 CSoutput.t149 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X381 gnd.t66 commonsourceibias.t68 commonsourceibias.t69 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X382 CSoutput.t214 a_n8964_8799.t122 vdd.t274 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X383 CSoutput.t215 a_n8964_8799.t123 vdd.t275 vdd.t53 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X384 CSoutput.t146 a_n8964_8799.t124 vdd.t54 vdd.t53 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X385 a_n2804_13878.t9 a_n2982_13878.t51 a_n2982_13878.t52 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X386 outputibias.t1 outputibias.t0 gnd.t380 gnd.t379 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X387 vdd.t55 a_n8964_8799.t125 CSoutput.t147 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X388 gnd.t64 commonsourceibias.t66 commonsourceibias.t67 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X389 commonsourceibias.t65 commonsourceibias.t64 gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X390 gnd.t232 gnd.t229 gnd.t231 gnd.t230 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X391 gnd.t61 commonsourceibias.t176 CSoutput.t27 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X392 gnd.t60 commonsourceibias.t177 CSoutput.t26 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X393 a_n2903_n3924.t22 minus.t22 a_n2982_13878.t2 gnd.t343 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X394 a_n2903_n3924.t43 diffpairibias.t22 gnd.t393 gnd.t392 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X395 gnd.t59 commonsourceibias.t178 CSoutput.t25 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X396 vdd.t24 a_n8964_8799.t126 CSoutput.t128 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X397 CSoutput.t24 commonsourceibias.t179 gnd.t55 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X398 gnd.t57 commonsourceibias.t180 CSoutput.t23 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X399 CSoutput.t129 a_n8964_8799.t127 vdd.t25 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X400 CSoutput.t22 commonsourceibias.t181 gnd.t54 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X401 a_n2982_13878.t62 a_n2982_13878.t61 a_n2804_13878.t8 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X402 gnd.t228 gnd.t225 gnd.t227 gnd.t226 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X403 a_n8964_8799.t24 a_n2982_13878.t102 a_n2982_8322.t9 vdd.t203 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X404 vdd.t193 CSoutput.t236 output.t0 gnd.t395 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X405 vdd.t20 a_n8964_8799.t128 CSoutput.t126 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X406 CSoutput.t127 a_n8964_8799.t129 vdd.t22 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X407 vdd.t79 vdd.t77 vdd.t78 vdd.t74 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X408 CSoutput.t21 commonsourceibias.t182 gnd.t52 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X409 gnd.t49 commonsourceibias.t183 CSoutput.t20 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X410 commonsourceibias.t33 commonsourceibias.t32 gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X411 CSoutput.t19 commonsourceibias.t184 gnd.t51 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X412 CSoutput.t138 a_n8964_8799.t130 vdd.t41 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X413 gnd.t224 gnd.t221 gnd.t223 gnd.t222 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X414 diffpairibias.t3 diffpairibias.t2 gnd.t218 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X415 a_n2982_8322.t8 a_n2982_13878.t103 a_n8964_8799.t23 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X416 CSoutput.t18 commonsourceibias.t185 gnd.t45 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X417 gnd.t43 commonsourceibias.t186 CSoutput.t17 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X418 a_n2982_13878.t5 minus.t23 a_n2903_n3924.t27 gnd.t352 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X419 vdd.t42 a_n8964_8799.t131 CSoutput.t139 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X420 CSoutput.t156 a_n8964_8799.t132 vdd.t148 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X421 CSoutput.t157 a_n8964_8799.t133 vdd.t149 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X422 diffpairibias.t1 diffpairibias.t0 gnd.t371 gnd.t370 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X423 gnd.t42 commonsourceibias.t187 CSoutput.t16 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X424 CSoutput.t237 a_n2982_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X425 commonsourceibias.t61 commonsourceibias.t60 gnd.t40 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X426 gnd.t39 commonsourceibias.t188 CSoutput.t15 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X427 commonsourceibias.t17 commonsourceibias.t16 gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X428 CSoutput.t14 commonsourceibias.t189 gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X429 vdd.t201 a_n2982_13878.t104 a_n2804_13878.t0 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X430 CSoutput.t158 a_n8964_8799.t134 vdd.t150 vdd.t53 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X431 gnd.t34 commonsourceibias.t62 commonsourceibias.t63 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X432 vdd.t151 a_n8964_8799.t135 CSoutput.t159 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X433 gnd.t32 commonsourceibias.t58 commonsourceibias.t59 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X434 a_n8964_8799.t1 plus.t22 a_n2903_n3924.t3 gnd.t341 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X435 a_n2982_8322.t7 a_n2982_13878.t105 a_n8964_8799.t22 vdd.t199 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X436 gnd.t30 commonsourceibias.t190 CSoutput.t13 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X437 a_n2982_13878.t13 minus.t24 a_n2903_n3924.t39 gnd.t386 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X438 commonsourceibias.t57 commonsourceibias.t56 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X439 gnd.t26 commonsourceibias.t191 CSoutput.t12 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X440 gnd.t28 commonsourceibias.t192 CSoutput.t11 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X441 a_n8964_8799.t12 plus.t23 a_n2903_n3924.t2 gnd.t372 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X442 gnd.t22 commonsourceibias.t193 CSoutput.t10 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X443 a_n2982_8322.t6 a_n2982_13878.t106 a_n8964_8799.t21 vdd.t198 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X444 vdd.t260 a_n8964_8799.t136 CSoutput.t200 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X445 vdd.t261 a_n8964_8799.t137 CSoutput.t201 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X446 output.t16 outputibias.t11 gnd.t363 gnd.t362 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X447 CSoutput.t124 a_n8964_8799.t138 vdd.t16 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X448 gnd.t20 commonsourceibias.t194 CSoutput.t9 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X449 vdd.t76 vdd.t73 vdd.t75 vdd.t74 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X450 a_n2982_8322.t30 a_n2982_13878.t107 vdd.t197 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X451 gnd.t19 commonsourceibias.t195 CSoutput.t8 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X452 a_n2804_13878.t7 a_n2982_13878.t31 a_n2982_13878.t32 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X453 gnd.t17 commonsourceibias.t196 CSoutput.t7 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X454 CSoutput.t6 commonsourceibias.t197 gnd.t11 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X455 commonsourceibias.t15 commonsourceibias.t14 gnd.t13 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X456 CSoutput.t5 commonsourceibias.t198 gnd.t15 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X457 vdd.t72 vdd.t69 vdd.t71 vdd.t70 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X458 a_n2903_n3924.t1 plus.t24 a_n8964_8799.t7 gnd.t361 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X459 a_n2903_n3924.t29 diffpairibias.t23 gnd.t357 gnd.t356 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X460 vdd.t68 vdd.t65 vdd.t67 vdd.t66 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X461 CSoutput.t125 a_n8964_8799.t139 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X462 a_n2982_13878.t40 a_n2982_13878.t39 a_n2804_13878.t6 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X463 gnd.t9 commonsourceibias.t199 CSoutput.t4 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
R0 a_n2982_13878.n125 a_n2982_13878.t90 512.366
R1 a_n2982_13878.n115 a_n2982_13878.t79 512.366
R2 a_n2982_13878.n126 a_n2982_13878.t68 512.366
R3 a_n2982_13878.n123 a_n2982_13878.t98 512.366
R4 a_n2982_13878.n116 a_n2982_13878.t87 512.366
R5 a_n2982_13878.n124 a_n2982_13878.t86 512.366
R6 a_n2982_13878.n121 a_n2982_13878.t94 512.366
R7 a_n2982_13878.n117 a_n2982_13878.t77 512.366
R8 a_n2982_13878.n122 a_n2982_13878.t78 512.366
R9 a_n2982_13878.n119 a_n2982_13878.t81 512.366
R10 a_n2982_13878.n118 a_n2982_13878.t92 512.366
R11 a_n2982_13878.n120 a_n2982_13878.t107 512.366
R12 a_n2982_13878.n30 a_n2982_13878.t106 538.698
R13 a_n2982_13878.n134 a_n2982_13878.t83 512.366
R14 a_n2982_13878.n133 a_n2982_13878.t88 512.366
R15 a_n2982_13878.n86 a_n2982_13878.t76 512.366
R16 a_n2982_13878.n132 a_n2982_13878.t93 512.366
R17 a_n2982_13878.n131 a_n2982_13878.t102 512.366
R18 a_n2982_13878.n87 a_n2982_13878.t103 512.366
R19 a_n2982_13878.n130 a_n2982_13878.t70 512.366
R20 a_n2982_13878.n129 a_n2982_13878.t85 512.366
R21 a_n2982_13878.n88 a_n2982_13878.t73 512.366
R22 a_n2982_13878.n128 a_n2982_13878.t80 512.366
R23 a_n2982_13878.n49 a_n2982_13878.t31 532.5
R24 a_n2982_13878.n135 a_n2982_13878.t53 512.366
R25 a_n2982_13878.n83 a_n2982_13878.t51 512.366
R26 a_n2982_13878.n36 a_n2982_13878.t17 538.698
R27 a_n2982_13878.n151 a_n2982_13878.t23 512.366
R28 a_n2982_13878.n150 a_n2982_13878.t21 512.366
R29 a_n2982_13878.n84 a_n2982_13878.t63 512.366
R30 a_n2982_13878.n149 a_n2982_13878.t25 512.366
R31 a_n2982_13878.n148 a_n2982_13878.t57 512.366
R32 a_n2982_13878.n85 a_n2982_13878.t61 512.366
R33 a_n2982_13878.n147 a_n2982_13878.t59 512.366
R34 a_n2982_13878.n146 a_n2982_13878.t45 512.366
R35 a_n2982_13878.n18 a_n2982_13878.t49 538.698
R36 a_n2982_13878.n108 a_n2982_13878.t33 512.366
R37 a_n2982_13878.n97 a_n2982_13878.t39 512.366
R38 a_n2982_13878.n109 a_n2982_13878.t37 512.366
R39 a_n2982_13878.n96 a_n2982_13878.t43 512.366
R40 a_n2982_13878.n110 a_n2982_13878.t47 512.366
R41 a_n2982_13878.n111 a_n2982_13878.t27 512.366
R42 a_n2982_13878.n95 a_n2982_13878.t41 512.366
R43 a_n2982_13878.n112 a_n2982_13878.t35 512.366
R44 a_n2982_13878.n94 a_n2982_13878.t55 512.366
R45 a_n2982_13878.n113 a_n2982_13878.t19 512.366
R46 a_n2982_13878.n24 a_n2982_13878.t105 538.698
R47 a_n2982_13878.n102 a_n2982_13878.t74 512.366
R48 a_n2982_13878.n101 a_n2982_13878.t75 512.366
R49 a_n2982_13878.n103 a_n2982_13878.t100 512.366
R50 a_n2982_13878.n100 a_n2982_13878.t101 512.366
R51 a_n2982_13878.n104 a_n2982_13878.t72 512.366
R52 a_n2982_13878.n105 a_n2982_13878.t96 512.366
R53 a_n2982_13878.n99 a_n2982_13878.t97 512.366
R54 a_n2982_13878.n106 a_n2982_13878.t69 512.366
R55 a_n2982_13878.n98 a_n2982_13878.t82 512.366
R56 a_n2982_13878.n107 a_n2982_13878.t91 512.366
R57 a_n2982_13878.n4 a_n2982_13878.n81 70.1674
R58 a_n2982_13878.n6 a_n2982_13878.n79 70.1674
R59 a_n2982_13878.n8 a_n2982_13878.n77 70.1674
R60 a_n2982_13878.n11 a_n2982_13878.n75 70.1674
R61 a_n2982_13878.n57 a_n2982_13878.n25 70.5844
R62 a_n2982_13878.n48 a_n2982_13878.n31 74.73
R63 a_n2982_13878.n146 a_n2982_13878.n48 11.843
R64 a_n2982_13878.n47 a_n2982_13878.n32 80.4688
R65 a_n2982_13878.n47 a_n2982_13878.n147 0.365327
R66 a_n2982_13878.n33 a_n2982_13878.n46 75.0448
R67 a_n2982_13878.n45 a_n2982_13878.n33 70.1674
R68 a_n2982_13878.n149 a_n2982_13878.n45 20.9683
R69 a_n2982_13878.n35 a_n2982_13878.n44 70.3058
R70 a_n2982_13878.n44 a_n2982_13878.n84 20.6913
R71 a_n2982_13878.n43 a_n2982_13878.n35 75.3623
R72 a_n2982_13878.n150 a_n2982_13878.n43 10.5784
R73 a_n2982_13878.n34 a_n2982_13878.n36 44.7878
R74 a_n2982_13878.n82 a_n2982_13878.n83 20.9683
R75 a_n2982_13878.n49 a_n2982_13878.n31 70.5844
R76 a_n2982_13878.n31 a_n2982_13878.n82 70.1674
R77 a_n2982_13878.n25 a_n2982_13878.n56 70.1674
R78 a_n2982_13878.n56 a_n2982_13878.n88 20.9683
R79 a_n2982_13878.n55 a_n2982_13878.n26 74.73
R80 a_n2982_13878.n129 a_n2982_13878.n55 11.843
R81 a_n2982_13878.n54 a_n2982_13878.n26 80.4688
R82 a_n2982_13878.n54 a_n2982_13878.n130 0.365327
R83 a_n2982_13878.n27 a_n2982_13878.n53 75.0448
R84 a_n2982_13878.n52 a_n2982_13878.n27 70.1674
R85 a_n2982_13878.n132 a_n2982_13878.n52 20.9683
R86 a_n2982_13878.n29 a_n2982_13878.n51 70.3058
R87 a_n2982_13878.n51 a_n2982_13878.n86 20.6913
R88 a_n2982_13878.n50 a_n2982_13878.n29 75.3623
R89 a_n2982_13878.n133 a_n2982_13878.n50 10.5784
R90 a_n2982_13878.n28 a_n2982_13878.n30 44.7878
R91 a_n2982_13878.n14 a_n2982_13878.n73 70.5844
R92 a_n2982_13878.n20 a_n2982_13878.n65 70.5844
R93 a_n2982_13878.n64 a_n2982_13878.n20 70.1674
R94 a_n2982_13878.n64 a_n2982_13878.n98 20.9683
R95 a_n2982_13878.n19 a_n2982_13878.n63 74.73
R96 a_n2982_13878.n106 a_n2982_13878.n63 11.843
R97 a_n2982_13878.n62 a_n2982_13878.n19 80.4688
R98 a_n2982_13878.n62 a_n2982_13878.n99 0.365327
R99 a_n2982_13878.n21 a_n2982_13878.n61 75.0448
R100 a_n2982_13878.n60 a_n2982_13878.n21 70.1674
R101 a_n2982_13878.n60 a_n2982_13878.n100 20.9683
R102 a_n2982_13878.n22 a_n2982_13878.n59 70.3058
R103 a_n2982_13878.n103 a_n2982_13878.n59 20.6913
R104 a_n2982_13878.n58 a_n2982_13878.n22 75.3623
R105 a_n2982_13878.n58 a_n2982_13878.n101 10.5784
R106 a_n2982_13878.n24 a_n2982_13878.n23 44.7878
R107 a_n2982_13878.n72 a_n2982_13878.n14 70.1674
R108 a_n2982_13878.n72 a_n2982_13878.n94 20.9683
R109 a_n2982_13878.n13 a_n2982_13878.n71 74.73
R110 a_n2982_13878.n112 a_n2982_13878.n71 11.843
R111 a_n2982_13878.n70 a_n2982_13878.n13 80.4688
R112 a_n2982_13878.n70 a_n2982_13878.n95 0.365327
R113 a_n2982_13878.n15 a_n2982_13878.n69 75.0448
R114 a_n2982_13878.n68 a_n2982_13878.n15 70.1674
R115 a_n2982_13878.n68 a_n2982_13878.n96 20.9683
R116 a_n2982_13878.n16 a_n2982_13878.n67 70.3058
R117 a_n2982_13878.n109 a_n2982_13878.n67 20.6913
R118 a_n2982_13878.n66 a_n2982_13878.n16 75.3623
R119 a_n2982_13878.n66 a_n2982_13878.n97 10.5784
R120 a_n2982_13878.n18 a_n2982_13878.n17 44.7878
R121 a_n2982_13878.n120 a_n2982_13878.n75 20.9683
R122 a_n2982_13878.n74 a_n2982_13878.n12 75.0448
R123 a_n2982_13878.n74 a_n2982_13878.n118 11.2134
R124 a_n2982_13878.n12 a_n2982_13878.n119 161.3
R125 a_n2982_13878.n122 a_n2982_13878.n77 20.9683
R126 a_n2982_13878.n76 a_n2982_13878.n9 75.0448
R127 a_n2982_13878.n76 a_n2982_13878.n117 11.2134
R128 a_n2982_13878.n9 a_n2982_13878.n121 161.3
R129 a_n2982_13878.n124 a_n2982_13878.n79 20.9683
R130 a_n2982_13878.n78 a_n2982_13878.n7 75.0448
R131 a_n2982_13878.n78 a_n2982_13878.n116 11.2134
R132 a_n2982_13878.n7 a_n2982_13878.n123 161.3
R133 a_n2982_13878.n126 a_n2982_13878.n81 20.9683
R134 a_n2982_13878.n80 a_n2982_13878.n5 75.0448
R135 a_n2982_13878.n80 a_n2982_13878.n115 11.2134
R136 a_n2982_13878.n5 a_n2982_13878.n125 161.3
R137 a_n2982_13878.n3 a_n2982_13878.n144 81.4626
R138 a_n2982_13878.n1 a_n2982_13878.n139 81.4626
R139 a_n2982_13878.n0 a_n2982_13878.n136 81.4626
R140 a_n2982_13878.n3 a_n2982_13878.n145 80.9324
R141 a_n2982_13878.n3 a_n2982_13878.n143 80.9324
R142 a_n2982_13878.n2 a_n2982_13878.n142 80.9324
R143 a_n2982_13878.n2 a_n2982_13878.n141 80.9324
R144 a_n2982_13878.n1 a_n2982_13878.n140 80.9324
R145 a_n2982_13878.n1 a_n2982_13878.n138 80.9324
R146 a_n2982_13878.n0 a_n2982_13878.n137 80.9324
R147 a_n2982_13878.n42 a_n2982_13878.t32 74.6477
R148 a_n2982_13878.n37 a_n2982_13878.t50 74.6477
R149 a_n2982_13878.t18 a_n2982_13878.n41 74.2899
R150 a_n2982_13878.n39 a_n2982_13878.t30 74.2897
R151 a_n2982_13878.n42 a_n2982_13878.n153 70.6783
R152 a_n2982_13878.n42 a_n2982_13878.n154 70.6783
R153 a_n2982_13878.n40 a_n2982_13878.n155 70.6783
R154 a_n2982_13878.n40 a_n2982_13878.n156 70.6783
R155 a_n2982_13878.n41 a_n2982_13878.n157 70.6783
R156 a_n2982_13878.n39 a_n2982_13878.n93 70.6783
R157 a_n2982_13878.n38 a_n2982_13878.n92 70.6783
R158 a_n2982_13878.n38 a_n2982_13878.n91 70.6783
R159 a_n2982_13878.n37 a_n2982_13878.n90 70.6783
R160 a_n2982_13878.n37 a_n2982_13878.n89 70.6783
R161 a_n2982_13878.n125 a_n2982_13878.n115 48.2005
R162 a_n2982_13878.t95 a_n2982_13878.n81 533.335
R163 a_n2982_13878.n123 a_n2982_13878.n116 48.2005
R164 a_n2982_13878.t104 a_n2982_13878.n79 533.335
R165 a_n2982_13878.n121 a_n2982_13878.n117 48.2005
R166 a_n2982_13878.t89 a_n2982_13878.n77 533.335
R167 a_n2982_13878.n119 a_n2982_13878.n118 48.2005
R168 a_n2982_13878.t84 a_n2982_13878.n75 533.335
R169 a_n2982_13878.n134 a_n2982_13878.n133 48.2005
R170 a_n2982_13878.n52 a_n2982_13878.n131 20.9683
R171 a_n2982_13878.n130 a_n2982_13878.n87 48.2005
R172 a_n2982_13878.n128 a_n2982_13878.n56 20.9683
R173 a_n2982_13878.n135 a_n2982_13878.n82 20.9683
R174 a_n2982_13878.n151 a_n2982_13878.n150 48.2005
R175 a_n2982_13878.n45 a_n2982_13878.n148 20.9683
R176 a_n2982_13878.n147 a_n2982_13878.n85 48.2005
R177 a_n2982_13878.n108 a_n2982_13878.n97 48.2005
R178 a_n2982_13878.n110 a_n2982_13878.n68 20.9683
R179 a_n2982_13878.n111 a_n2982_13878.n95 48.2005
R180 a_n2982_13878.n113 a_n2982_13878.n72 20.9683
R181 a_n2982_13878.n102 a_n2982_13878.n101 48.2005
R182 a_n2982_13878.n104 a_n2982_13878.n60 20.9683
R183 a_n2982_13878.n105 a_n2982_13878.n99 48.2005
R184 a_n2982_13878.n107 a_n2982_13878.n64 20.9683
R185 a_n2982_13878.n132 a_n2982_13878.n51 21.4216
R186 a_n2982_13878.n149 a_n2982_13878.n44 21.4216
R187 a_n2982_13878.n96 a_n2982_13878.n67 21.4216
R188 a_n2982_13878.n100 a_n2982_13878.n59 21.4216
R189 a_n2982_13878.n57 a_n2982_13878.t99 532.5
R190 a_n2982_13878.t29 a_n2982_13878.n73 532.5
R191 a_n2982_13878.t71 a_n2982_13878.n65 532.5
R192 a_n2982_13878.n2 a_n2982_13878.n1 32.7898
R193 a_n2982_13878.n55 a_n2982_13878.n88 34.4824
R194 a_n2982_13878.n48 a_n2982_13878.n83 34.4824
R195 a_n2982_13878.n94 a_n2982_13878.n71 34.4824
R196 a_n2982_13878.n98 a_n2982_13878.n63 34.4824
R197 a_n2982_13878.n126 a_n2982_13878.n80 35.3134
R198 a_n2982_13878.n124 a_n2982_13878.n78 35.3134
R199 a_n2982_13878.n122 a_n2982_13878.n76 35.3134
R200 a_n2982_13878.n120 a_n2982_13878.n74 35.3134
R201 a_n2982_13878.n131 a_n2982_13878.n53 35.3134
R202 a_n2982_13878.n53 a_n2982_13878.n87 11.2134
R203 a_n2982_13878.n148 a_n2982_13878.n46 35.3134
R204 a_n2982_13878.n46 a_n2982_13878.n85 11.2134
R205 a_n2982_13878.n69 a_n2982_13878.n110 35.3134
R206 a_n2982_13878.n111 a_n2982_13878.n69 11.2134
R207 a_n2982_13878.n61 a_n2982_13878.n104 35.3134
R208 a_n2982_13878.n105 a_n2982_13878.n61 11.2134
R209 a_n2982_13878.n31 a_n2982_13878.n3 23.891
R210 a_n2982_13878.n50 a_n2982_13878.n86 36.139
R211 a_n2982_13878.n43 a_n2982_13878.n84 36.139
R212 a_n2982_13878.n109 a_n2982_13878.n66 36.139
R213 a_n2982_13878.n103 a_n2982_13878.n58 36.139
R214 a_n2982_13878.n23 a_n2982_13878.n10 13.9285
R215 a_n2982_13878.n25 a_n2982_13878.n127 13.724
R216 a_n2982_13878.n152 a_n2982_13878.n34 12.4191
R217 a_n2982_13878.n127 a_n2982_13878.n4 11.2486
R218 a_n2982_13878.n12 a_n2982_13878.n10 11.2486
R219 a_n2982_13878.n114 a_n2982_13878.n39 10.5745
R220 a_n2982_13878.n114 a_n2982_13878.n14 8.58383
R221 a_n2982_13878.n41 a_n2982_13878.n152 6.7311
R222 a_n2982_13878.n127 a_n2982_13878.n114 5.3452
R223 a_n2982_13878.n31 a_n2982_13878.n28 3.94368
R224 a_n2982_13878.n17 a_n2982_13878.n20 3.94368
R225 a_n2982_13878.n153 a_n2982_13878.t52 3.61217
R226 a_n2982_13878.n153 a_n2982_13878.t54 3.61217
R227 a_n2982_13878.n154 a_n2982_13878.t60 3.61217
R228 a_n2982_13878.n154 a_n2982_13878.t46 3.61217
R229 a_n2982_13878.n155 a_n2982_13878.t58 3.61217
R230 a_n2982_13878.n155 a_n2982_13878.t62 3.61217
R231 a_n2982_13878.n156 a_n2982_13878.t64 3.61217
R232 a_n2982_13878.n156 a_n2982_13878.t26 3.61217
R233 a_n2982_13878.n157 a_n2982_13878.t24 3.61217
R234 a_n2982_13878.n157 a_n2982_13878.t22 3.61217
R235 a_n2982_13878.n93 a_n2982_13878.t56 3.61217
R236 a_n2982_13878.n93 a_n2982_13878.t20 3.61217
R237 a_n2982_13878.n92 a_n2982_13878.t42 3.61217
R238 a_n2982_13878.n92 a_n2982_13878.t36 3.61217
R239 a_n2982_13878.n91 a_n2982_13878.t48 3.61217
R240 a_n2982_13878.n91 a_n2982_13878.t28 3.61217
R241 a_n2982_13878.n90 a_n2982_13878.t38 3.61217
R242 a_n2982_13878.n90 a_n2982_13878.t44 3.61217
R243 a_n2982_13878.n89 a_n2982_13878.t34 3.61217
R244 a_n2982_13878.n89 a_n2982_13878.t40 3.61217
R245 a_n2982_13878.n144 a_n2982_13878.t65 2.82907
R246 a_n2982_13878.n144 a_n2982_13878.t13 2.82907
R247 a_n2982_13878.n145 a_n2982_13878.t8 2.82907
R248 a_n2982_13878.n145 a_n2982_13878.t7 2.82907
R249 a_n2982_13878.n143 a_n2982_13878.t6 2.82907
R250 a_n2982_13878.n143 a_n2982_13878.t4 2.82907
R251 a_n2982_13878.n142 a_n2982_13878.t9 2.82907
R252 a_n2982_13878.n142 a_n2982_13878.t14 2.82907
R253 a_n2982_13878.n141 a_n2982_13878.t1 2.82907
R254 a_n2982_13878.n141 a_n2982_13878.t67 2.82907
R255 a_n2982_13878.n139 a_n2982_13878.t10 2.82907
R256 a_n2982_13878.n139 a_n2982_13878.t11 2.82907
R257 a_n2982_13878.n140 a_n2982_13878.t15 2.82907
R258 a_n2982_13878.n140 a_n2982_13878.t12 2.82907
R259 a_n2982_13878.n138 a_n2982_13878.t2 2.82907
R260 a_n2982_13878.n138 a_n2982_13878.t5 2.82907
R261 a_n2982_13878.n137 a_n2982_13878.t0 2.82907
R262 a_n2982_13878.n137 a_n2982_13878.t16 2.82907
R263 a_n2982_13878.n136 a_n2982_13878.t3 2.82907
R264 a_n2982_13878.n136 a_n2982_13878.t66 2.82907
R265 a_n2982_13878.n30 a_n2982_13878.n134 14.1668
R266 a_n2982_13878.n128 a_n2982_13878.n57 22.3251
R267 a_n2982_13878.n135 a_n2982_13878.n49 22.3251
R268 a_n2982_13878.n36 a_n2982_13878.n151 14.1668
R269 a_n2982_13878.n108 a_n2982_13878.n18 14.1668
R270 a_n2982_13878.n73 a_n2982_13878.n113 22.3251
R271 a_n2982_13878.n102 a_n2982_13878.n24 14.1668
R272 a_n2982_13878.n65 a_n2982_13878.n107 22.3251
R273 a_n2982_13878.n152 a_n2982_13878.n10 1.30542
R274 a_n2982_13878.n7 a_n2982_13878.n8 1.04595
R275 a_n2982_13878.n54 a_n2982_13878.n129 47.835
R276 a_n2982_13878.n47 a_n2982_13878.n146 47.835
R277 a_n2982_13878.n112 a_n2982_13878.n70 47.835
R278 a_n2982_13878.n106 a_n2982_13878.n62 47.835
R279 a_n2982_13878.n3 a_n2982_13878.n2 1.59102
R280 a_n2982_13878.n26 a_n2982_13878.n25 1.13686
R281 a_n2982_13878.n20 a_n2982_13878.n19 1.13686
R282 a_n2982_13878.n14 a_n2982_13878.n13 1.13686
R283 a_n2982_13878.n31 a_n2982_13878.n32 1.09898
R284 a_n2982_13878.n41 a_n2982_13878.n40 1.07378
R285 a_n2982_13878.n38 a_n2982_13878.n37 1.07378
R286 a_n2982_13878.n1 a_n2982_13878.n0 1.06084
R287 a_n2982_13878.n35 a_n2982_13878.n34 0.758076
R288 a_n2982_13878.n35 a_n2982_13878.n33 0.758076
R289 a_n2982_13878.n33 a_n2982_13878.n32 0.758076
R290 a_n2982_13878.n29 a_n2982_13878.n28 0.758076
R291 a_n2982_13878.n29 a_n2982_13878.n27 0.758076
R292 a_n2982_13878.n27 a_n2982_13878.n26 0.758076
R293 a_n2982_13878.n22 a_n2982_13878.n23 0.758076
R294 a_n2982_13878.n21 a_n2982_13878.n22 0.758076
R295 a_n2982_13878.n19 a_n2982_13878.n21 0.758076
R296 a_n2982_13878.n16 a_n2982_13878.n17 0.758076
R297 a_n2982_13878.n15 a_n2982_13878.n16 0.758076
R298 a_n2982_13878.n13 a_n2982_13878.n15 0.758076
R299 a_n2982_13878.n12 a_n2982_13878.n11 0.758076
R300 a_n2982_13878.n9 a_n2982_13878.n8 0.758076
R301 a_n2982_13878.n7 a_n2982_13878.n6 0.758076
R302 a_n2982_13878.n5 a_n2982_13878.n4 0.758076
R303 a_n2982_13878.n40 a_n2982_13878.n42 0.716017
R304 a_n2982_13878.n39 a_n2982_13878.n38 0.716017
R305 a_n2982_13878.n9 a_n2982_13878.n11 0.67853
R306 a_n2982_13878.n5 a_n2982_13878.n6 0.67853
R307 a_n2804_13878.n29 a_n2804_13878.n28 98.9632
R308 a_n2804_13878.n2 a_n2804_13878.n0 98.7517
R309 a_n2804_13878.n22 a_n2804_13878.n21 98.6055
R310 a_n2804_13878.n24 a_n2804_13878.n23 98.6055
R311 a_n2804_13878.n26 a_n2804_13878.n25 98.6055
R312 a_n2804_13878.n28 a_n2804_13878.n27 98.6055
R313 a_n2804_13878.n10 a_n2804_13878.n9 98.6055
R314 a_n2804_13878.n8 a_n2804_13878.n7 98.6055
R315 a_n2804_13878.n6 a_n2804_13878.n5 98.6055
R316 a_n2804_13878.n4 a_n2804_13878.n3 98.6055
R317 a_n2804_13878.n2 a_n2804_13878.n1 98.6055
R318 a_n2804_13878.n20 a_n2804_13878.n19 98.6054
R319 a_n2804_13878.n12 a_n2804_13878.t1 74.6477
R320 a_n2804_13878.n17 a_n2804_13878.t2 74.2899
R321 a_n2804_13878.n14 a_n2804_13878.t5 74.2899
R322 a_n2804_13878.n13 a_n2804_13878.t0 74.2899
R323 a_n2804_13878.n16 a_n2804_13878.n15 70.6783
R324 a_n2804_13878.n12 a_n2804_13878.n11 70.6783
R325 a_n2804_13878.n18 a_n2804_13878.n10 15.7159
R326 a_n2804_13878.n20 a_n2804_13878.n18 12.6495
R327 a_n2804_13878.n18 a_n2804_13878.n17 8.38735
R328 a_n2804_13878.n19 a_n2804_13878.t13 3.61217
R329 a_n2804_13878.n19 a_n2804_13878.t22 3.61217
R330 a_n2804_13878.n21 a_n2804_13878.t26 3.61217
R331 a_n2804_13878.n21 a_n2804_13878.t12 3.61217
R332 a_n2804_13878.n23 a_n2804_13878.t16 3.61217
R333 a_n2804_13878.n23 a_n2804_13878.t17 3.61217
R334 a_n2804_13878.n25 a_n2804_13878.t27 3.61217
R335 a_n2804_13878.n25 a_n2804_13878.t28 3.61217
R336 a_n2804_13878.n27 a_n2804_13878.t6 3.61217
R337 a_n2804_13878.n27 a_n2804_13878.t18 3.61217
R338 a_n2804_13878.n15 a_n2804_13878.t30 3.61217
R339 a_n2804_13878.n15 a_n2804_13878.t3 3.61217
R340 a_n2804_13878.n11 a_n2804_13878.t4 3.61217
R341 a_n2804_13878.n11 a_n2804_13878.t31 3.61217
R342 a_n2804_13878.n9 a_n2804_13878.t19 3.61217
R343 a_n2804_13878.n9 a_n2804_13878.t7 3.61217
R344 a_n2804_13878.n7 a_n2804_13878.t24 3.61217
R345 a_n2804_13878.n7 a_n2804_13878.t9 3.61217
R346 a_n2804_13878.n5 a_n2804_13878.t8 3.61217
R347 a_n2804_13878.n5 a_n2804_13878.t11 3.61217
R348 a_n2804_13878.n3 a_n2804_13878.t21 3.61217
R349 a_n2804_13878.n3 a_n2804_13878.t14 3.61217
R350 a_n2804_13878.n1 a_n2804_13878.t25 3.61217
R351 a_n2804_13878.n1 a_n2804_13878.t15 3.61217
R352 a_n2804_13878.n0 a_n2804_13878.t10 3.61217
R353 a_n2804_13878.n0 a_n2804_13878.t20 3.61217
R354 a_n2804_13878.n29 a_n2804_13878.t23 3.61217
R355 a_n2804_13878.t29 a_n2804_13878.n29 3.61217
R356 a_n2804_13878.n13 a_n2804_13878.n12 0.358259
R357 a_n2804_13878.n16 a_n2804_13878.n14 0.358259
R358 a_n2804_13878.n17 a_n2804_13878.n16 0.358259
R359 a_n2804_13878.n28 a_n2804_13878.n26 0.358259
R360 a_n2804_13878.n26 a_n2804_13878.n24 0.358259
R361 a_n2804_13878.n24 a_n2804_13878.n22 0.358259
R362 a_n2804_13878.n22 a_n2804_13878.n20 0.358259
R363 a_n2804_13878.n4 a_n2804_13878.n2 0.146627
R364 a_n2804_13878.n6 a_n2804_13878.n4 0.146627
R365 a_n2804_13878.n8 a_n2804_13878.n6 0.146627
R366 a_n2804_13878.n10 a_n2804_13878.n8 0.146627
R367 a_n2804_13878.n14 a_n2804_13878.n13 0.101793
R368 vdd.n315 vdd.n279 756.745
R369 vdd.n260 vdd.n224 756.745
R370 vdd.n217 vdd.n181 756.745
R371 vdd.n162 vdd.n126 756.745
R372 vdd.n120 vdd.n84 756.745
R373 vdd.n65 vdd.n29 756.745
R374 vdd.n2139 vdd.n2103 756.745
R375 vdd.n2194 vdd.n2158 756.745
R376 vdd.n2041 vdd.n2005 756.745
R377 vdd.n2096 vdd.n2060 756.745
R378 vdd.n1944 vdd.n1908 756.745
R379 vdd.n1999 vdd.n1963 756.745
R380 vdd.n1286 vdd.t69 640.208
R381 vdd.n981 vdd.t114 640.208
R382 vdd.n1290 vdd.t104 640.208
R383 vdd.n972 vdd.t138 640.208
R384 vdd.n867 vdd.t91 640.208
R385 vdd.n2740 vdd.t132 640.208
R386 vdd.n804 vdd.t80 640.208
R387 vdd.n2737 vdd.t121 640.208
R388 vdd.n768 vdd.t65 640.208
R389 vdd.n1042 vdd.t128 640.208
R390 vdd.n1603 vdd.t110 592.009
R391 vdd.n1759 vdd.t125 592.009
R392 vdd.n1795 vdd.t135 592.009
R393 vdd.n2279 vdd.t95 592.009
R394 vdd.n1219 vdd.t73 592.009
R395 vdd.n1179 vdd.t77 592.009
R396 vdd.n405 vdd.t107 592.009
R397 vdd.n419 vdd.t83 592.009
R398 vdd.n431 vdd.t98 592.009
R399 vdd.n723 vdd.t101 592.009
R400 vdd.n686 vdd.t118 592.009
R401 vdd.n3285 vdd.t87 592.009
R402 vdd.n316 vdd.n315 585
R403 vdd.n314 vdd.n281 585
R404 vdd.n313 vdd.n312 585
R405 vdd.n284 vdd.n282 585
R406 vdd.n307 vdd.n306 585
R407 vdd.n305 vdd.n304 585
R408 vdd.n288 vdd.n287 585
R409 vdd.n299 vdd.n298 585
R410 vdd.n297 vdd.n296 585
R411 vdd.n292 vdd.n291 585
R412 vdd.n261 vdd.n260 585
R413 vdd.n259 vdd.n226 585
R414 vdd.n258 vdd.n257 585
R415 vdd.n229 vdd.n227 585
R416 vdd.n252 vdd.n251 585
R417 vdd.n250 vdd.n249 585
R418 vdd.n233 vdd.n232 585
R419 vdd.n244 vdd.n243 585
R420 vdd.n242 vdd.n241 585
R421 vdd.n237 vdd.n236 585
R422 vdd.n218 vdd.n217 585
R423 vdd.n216 vdd.n183 585
R424 vdd.n215 vdd.n214 585
R425 vdd.n186 vdd.n184 585
R426 vdd.n209 vdd.n208 585
R427 vdd.n207 vdd.n206 585
R428 vdd.n190 vdd.n189 585
R429 vdd.n201 vdd.n200 585
R430 vdd.n199 vdd.n198 585
R431 vdd.n194 vdd.n193 585
R432 vdd.n163 vdd.n162 585
R433 vdd.n161 vdd.n128 585
R434 vdd.n160 vdd.n159 585
R435 vdd.n131 vdd.n129 585
R436 vdd.n154 vdd.n153 585
R437 vdd.n152 vdd.n151 585
R438 vdd.n135 vdd.n134 585
R439 vdd.n146 vdd.n145 585
R440 vdd.n144 vdd.n143 585
R441 vdd.n139 vdd.n138 585
R442 vdd.n121 vdd.n120 585
R443 vdd.n119 vdd.n86 585
R444 vdd.n118 vdd.n117 585
R445 vdd.n89 vdd.n87 585
R446 vdd.n112 vdd.n111 585
R447 vdd.n110 vdd.n109 585
R448 vdd.n93 vdd.n92 585
R449 vdd.n104 vdd.n103 585
R450 vdd.n102 vdd.n101 585
R451 vdd.n97 vdd.n96 585
R452 vdd.n66 vdd.n65 585
R453 vdd.n64 vdd.n31 585
R454 vdd.n63 vdd.n62 585
R455 vdd.n34 vdd.n32 585
R456 vdd.n57 vdd.n56 585
R457 vdd.n55 vdd.n54 585
R458 vdd.n38 vdd.n37 585
R459 vdd.n49 vdd.n48 585
R460 vdd.n47 vdd.n46 585
R461 vdd.n42 vdd.n41 585
R462 vdd.n2140 vdd.n2139 585
R463 vdd.n2138 vdd.n2105 585
R464 vdd.n2137 vdd.n2136 585
R465 vdd.n2108 vdd.n2106 585
R466 vdd.n2131 vdd.n2130 585
R467 vdd.n2129 vdd.n2128 585
R468 vdd.n2112 vdd.n2111 585
R469 vdd.n2123 vdd.n2122 585
R470 vdd.n2121 vdd.n2120 585
R471 vdd.n2116 vdd.n2115 585
R472 vdd.n2195 vdd.n2194 585
R473 vdd.n2193 vdd.n2160 585
R474 vdd.n2192 vdd.n2191 585
R475 vdd.n2163 vdd.n2161 585
R476 vdd.n2186 vdd.n2185 585
R477 vdd.n2184 vdd.n2183 585
R478 vdd.n2167 vdd.n2166 585
R479 vdd.n2178 vdd.n2177 585
R480 vdd.n2176 vdd.n2175 585
R481 vdd.n2171 vdd.n2170 585
R482 vdd.n2042 vdd.n2041 585
R483 vdd.n2040 vdd.n2007 585
R484 vdd.n2039 vdd.n2038 585
R485 vdd.n2010 vdd.n2008 585
R486 vdd.n2033 vdd.n2032 585
R487 vdd.n2031 vdd.n2030 585
R488 vdd.n2014 vdd.n2013 585
R489 vdd.n2025 vdd.n2024 585
R490 vdd.n2023 vdd.n2022 585
R491 vdd.n2018 vdd.n2017 585
R492 vdd.n2097 vdd.n2096 585
R493 vdd.n2095 vdd.n2062 585
R494 vdd.n2094 vdd.n2093 585
R495 vdd.n2065 vdd.n2063 585
R496 vdd.n2088 vdd.n2087 585
R497 vdd.n2086 vdd.n2085 585
R498 vdd.n2069 vdd.n2068 585
R499 vdd.n2080 vdd.n2079 585
R500 vdd.n2078 vdd.n2077 585
R501 vdd.n2073 vdd.n2072 585
R502 vdd.n1945 vdd.n1944 585
R503 vdd.n1943 vdd.n1910 585
R504 vdd.n1942 vdd.n1941 585
R505 vdd.n1913 vdd.n1911 585
R506 vdd.n1936 vdd.n1935 585
R507 vdd.n1934 vdd.n1933 585
R508 vdd.n1917 vdd.n1916 585
R509 vdd.n1928 vdd.n1927 585
R510 vdd.n1926 vdd.n1925 585
R511 vdd.n1921 vdd.n1920 585
R512 vdd.n2000 vdd.n1999 585
R513 vdd.n1998 vdd.n1965 585
R514 vdd.n1997 vdd.n1996 585
R515 vdd.n1968 vdd.n1966 585
R516 vdd.n1991 vdd.n1990 585
R517 vdd.n1989 vdd.n1988 585
R518 vdd.n1972 vdd.n1971 585
R519 vdd.n1983 vdd.n1982 585
R520 vdd.n1981 vdd.n1980 585
R521 vdd.n1976 vdd.n1975 585
R522 vdd.n445 vdd.n370 462.44
R523 vdd.n3523 vdd.n372 462.44
R524 vdd.n3418 vdd.n657 462.44
R525 vdd.n3416 vdd.n660 462.44
R526 vdd.n2274 vdd.n1502 462.44
R527 vdd.n2277 vdd.n2276 462.44
R528 vdd.n1830 vdd.n1600 462.44
R529 vdd.n1827 vdd.n1598 462.44
R530 vdd.n293 vdd.t57 329.043
R531 vdd.n238 vdd.t52 329.043
R532 vdd.n195 vdd.t148 329.043
R533 vdd.n140 vdd.t273 329.043
R534 vdd.n98 vdd.t160 329.043
R535 vdd.n43 vdd.t175 329.043
R536 vdd.n2117 vdd.t166 329.043
R537 vdd.n2172 vdd.t48 329.043
R538 vdd.n2019 vdd.t185 329.043
R539 vdd.n2074 vdd.t177 329.043
R540 vdd.n1922 vdd.t174 329.043
R541 vdd.n1977 vdd.t168 329.043
R542 vdd.n1603 vdd.t113 319.788
R543 vdd.n1759 vdd.t127 319.788
R544 vdd.n1795 vdd.t137 319.788
R545 vdd.n2279 vdd.t96 319.788
R546 vdd.n1219 vdd.t75 319.788
R547 vdd.n1179 vdd.t78 319.788
R548 vdd.n405 vdd.t108 319.788
R549 vdd.n419 vdd.t85 319.788
R550 vdd.n431 vdd.t99 319.788
R551 vdd.n723 vdd.t103 319.788
R552 vdd.n686 vdd.t120 319.788
R553 vdd.n3285 vdd.t90 319.788
R554 vdd.n1604 vdd.t112 303.69
R555 vdd.n1760 vdd.t126 303.69
R556 vdd.n1796 vdd.t136 303.69
R557 vdd.n2280 vdd.t97 303.69
R558 vdd.n1220 vdd.t76 303.69
R559 vdd.n1180 vdd.t79 303.69
R560 vdd.n406 vdd.t109 303.69
R561 vdd.n420 vdd.t86 303.69
R562 vdd.n432 vdd.t100 303.69
R563 vdd.n724 vdd.t102 303.69
R564 vdd.n687 vdd.t119 303.69
R565 vdd.n3286 vdd.t89 303.69
R566 vdd.n3007 vdd.n931 279.512
R567 vdd.n3247 vdd.n778 279.512
R568 vdd.n3184 vdd.n775 279.512
R569 vdd.n2939 vdd.n2938 279.512
R570 vdd.n2700 vdd.n969 279.512
R571 vdd.n2631 vdd.n2630 279.512
R572 vdd.n1326 vdd.n1325 279.512
R573 vdd.n2425 vdd.n1109 279.512
R574 vdd.n3163 vdd.n776 279.512
R575 vdd.n3250 vdd.n3249 279.512
R576 vdd.n2812 vdd.n2735 279.512
R577 vdd.n2743 vdd.n927 279.512
R578 vdd.n2628 vdd.n979 279.512
R579 vdd.n977 vdd.n951 279.512
R580 vdd.n1451 vdd.n1146 279.512
R581 vdd.n1251 vdd.n1104 279.512
R582 vdd.n2423 vdd.n1112 254.619
R583 vdd.n756 vdd.n658 254.619
R584 vdd.n3165 vdd.n776 185
R585 vdd.n3248 vdd.n776 185
R586 vdd.n3167 vdd.n3166 185
R587 vdd.n3166 vdd.n774 185
R588 vdd.n3168 vdd.n810 185
R589 vdd.n3178 vdd.n810 185
R590 vdd.n3169 vdd.n819 185
R591 vdd.n819 vdd.n817 185
R592 vdd.n3171 vdd.n3170 185
R593 vdd.n3172 vdd.n3171 185
R594 vdd.n3124 vdd.n818 185
R595 vdd.n818 vdd.n814 185
R596 vdd.n3123 vdd.n3122 185
R597 vdd.n3122 vdd.n3121 185
R598 vdd.n821 vdd.n820 185
R599 vdd.n822 vdd.n821 185
R600 vdd.n3114 vdd.n3113 185
R601 vdd.n3115 vdd.n3114 185
R602 vdd.n3112 vdd.n830 185
R603 vdd.n835 vdd.n830 185
R604 vdd.n3111 vdd.n3110 185
R605 vdd.n3110 vdd.n3109 185
R606 vdd.n832 vdd.n831 185
R607 vdd.n841 vdd.n832 185
R608 vdd.n3102 vdd.n3101 185
R609 vdd.n3103 vdd.n3102 185
R610 vdd.n3100 vdd.n842 185
R611 vdd.n848 vdd.n842 185
R612 vdd.n3099 vdd.n3098 185
R613 vdd.n3098 vdd.n3097 185
R614 vdd.n844 vdd.n843 185
R615 vdd.n845 vdd.n844 185
R616 vdd.n3090 vdd.n3089 185
R617 vdd.n3091 vdd.n3090 185
R618 vdd.n3088 vdd.n855 185
R619 vdd.n855 vdd.n852 185
R620 vdd.n3087 vdd.n3086 185
R621 vdd.n3086 vdd.n3085 185
R622 vdd.n857 vdd.n856 185
R623 vdd.n858 vdd.n857 185
R624 vdd.n3078 vdd.n3077 185
R625 vdd.n3079 vdd.n3078 185
R626 vdd.n3076 vdd.n866 185
R627 vdd.n872 vdd.n866 185
R628 vdd.n3075 vdd.n3074 185
R629 vdd.n3074 vdd.n3073 185
R630 vdd.n3064 vdd.n869 185
R631 vdd.n879 vdd.n869 185
R632 vdd.n3066 vdd.n3065 185
R633 vdd.n3067 vdd.n3066 185
R634 vdd.n3063 vdd.n880 185
R635 vdd.n880 vdd.n876 185
R636 vdd.n3062 vdd.n3061 185
R637 vdd.n3061 vdd.n3060 185
R638 vdd.n882 vdd.n881 185
R639 vdd.n883 vdd.n882 185
R640 vdd.n3053 vdd.n3052 185
R641 vdd.n3054 vdd.n3053 185
R642 vdd.n3051 vdd.n891 185
R643 vdd.n896 vdd.n891 185
R644 vdd.n3050 vdd.n3049 185
R645 vdd.n3049 vdd.n3048 185
R646 vdd.n893 vdd.n892 185
R647 vdd.n902 vdd.n893 185
R648 vdd.n3041 vdd.n3040 185
R649 vdd.n3042 vdd.n3041 185
R650 vdd.n3039 vdd.n903 185
R651 vdd.n2915 vdd.n903 185
R652 vdd.n3038 vdd.n3037 185
R653 vdd.n3037 vdd.n3036 185
R654 vdd.n905 vdd.n904 185
R655 vdd.n2921 vdd.n905 185
R656 vdd.n3029 vdd.n3028 185
R657 vdd.n3030 vdd.n3029 185
R658 vdd.n3027 vdd.n914 185
R659 vdd.n914 vdd.n911 185
R660 vdd.n3026 vdd.n3025 185
R661 vdd.n3025 vdd.n3024 185
R662 vdd.n916 vdd.n915 185
R663 vdd.n917 vdd.n916 185
R664 vdd.n3017 vdd.n3016 185
R665 vdd.n3018 vdd.n3017 185
R666 vdd.n3015 vdd.n925 185
R667 vdd.n2933 vdd.n925 185
R668 vdd.n3014 vdd.n3013 185
R669 vdd.n3013 vdd.n3012 185
R670 vdd.n927 vdd.n926 185
R671 vdd.n928 vdd.n927 185
R672 vdd.n2744 vdd.n2743 185
R673 vdd.n2746 vdd.n2745 185
R674 vdd.n2748 vdd.n2747 185
R675 vdd.n2750 vdd.n2749 185
R676 vdd.n2752 vdd.n2751 185
R677 vdd.n2754 vdd.n2753 185
R678 vdd.n2756 vdd.n2755 185
R679 vdd.n2758 vdd.n2757 185
R680 vdd.n2760 vdd.n2759 185
R681 vdd.n2762 vdd.n2761 185
R682 vdd.n2764 vdd.n2763 185
R683 vdd.n2766 vdd.n2765 185
R684 vdd.n2768 vdd.n2767 185
R685 vdd.n2770 vdd.n2769 185
R686 vdd.n2772 vdd.n2771 185
R687 vdd.n2774 vdd.n2773 185
R688 vdd.n2776 vdd.n2775 185
R689 vdd.n2778 vdd.n2777 185
R690 vdd.n2780 vdd.n2779 185
R691 vdd.n2782 vdd.n2781 185
R692 vdd.n2784 vdd.n2783 185
R693 vdd.n2786 vdd.n2785 185
R694 vdd.n2788 vdd.n2787 185
R695 vdd.n2790 vdd.n2789 185
R696 vdd.n2792 vdd.n2791 185
R697 vdd.n2794 vdd.n2793 185
R698 vdd.n2796 vdd.n2795 185
R699 vdd.n2798 vdd.n2797 185
R700 vdd.n2800 vdd.n2799 185
R701 vdd.n2802 vdd.n2801 185
R702 vdd.n2804 vdd.n2803 185
R703 vdd.n2806 vdd.n2805 185
R704 vdd.n2808 vdd.n2807 185
R705 vdd.n2810 vdd.n2809 185
R706 vdd.n2811 vdd.n2735 185
R707 vdd.n3005 vdd.n2735 185
R708 vdd.n3251 vdd.n3250 185
R709 vdd.n3252 vdd.n767 185
R710 vdd.n3254 vdd.n3253 185
R711 vdd.n3256 vdd.n765 185
R712 vdd.n3258 vdd.n3257 185
R713 vdd.n3259 vdd.n764 185
R714 vdd.n3261 vdd.n3260 185
R715 vdd.n3263 vdd.n762 185
R716 vdd.n3265 vdd.n3264 185
R717 vdd.n3266 vdd.n761 185
R718 vdd.n3268 vdd.n3267 185
R719 vdd.n3270 vdd.n759 185
R720 vdd.n3272 vdd.n3271 185
R721 vdd.n3273 vdd.n758 185
R722 vdd.n3275 vdd.n3274 185
R723 vdd.n3277 vdd.n757 185
R724 vdd.n3278 vdd.n754 185
R725 vdd.n3281 vdd.n3280 185
R726 vdd.n755 vdd.n753 185
R727 vdd.n3137 vdd.n3136 185
R728 vdd.n3139 vdd.n3138 185
R729 vdd.n3141 vdd.n3133 185
R730 vdd.n3143 vdd.n3142 185
R731 vdd.n3144 vdd.n3132 185
R732 vdd.n3146 vdd.n3145 185
R733 vdd.n3148 vdd.n3130 185
R734 vdd.n3150 vdd.n3149 185
R735 vdd.n3151 vdd.n3129 185
R736 vdd.n3153 vdd.n3152 185
R737 vdd.n3155 vdd.n3127 185
R738 vdd.n3157 vdd.n3156 185
R739 vdd.n3158 vdd.n3126 185
R740 vdd.n3160 vdd.n3159 185
R741 vdd.n3162 vdd.n3125 185
R742 vdd.n3164 vdd.n3163 185
R743 vdd.n3163 vdd.n756 185
R744 vdd.n3249 vdd.n771 185
R745 vdd.n3249 vdd.n3248 185
R746 vdd.n2866 vdd.n773 185
R747 vdd.n774 vdd.n773 185
R748 vdd.n2867 vdd.n809 185
R749 vdd.n3178 vdd.n809 185
R750 vdd.n2869 vdd.n2868 185
R751 vdd.n2868 vdd.n817 185
R752 vdd.n2870 vdd.n816 185
R753 vdd.n3172 vdd.n816 185
R754 vdd.n2872 vdd.n2871 185
R755 vdd.n2871 vdd.n814 185
R756 vdd.n2873 vdd.n824 185
R757 vdd.n3121 vdd.n824 185
R758 vdd.n2875 vdd.n2874 185
R759 vdd.n2874 vdd.n822 185
R760 vdd.n2876 vdd.n829 185
R761 vdd.n3115 vdd.n829 185
R762 vdd.n2878 vdd.n2877 185
R763 vdd.n2877 vdd.n835 185
R764 vdd.n2879 vdd.n834 185
R765 vdd.n3109 vdd.n834 185
R766 vdd.n2881 vdd.n2880 185
R767 vdd.n2880 vdd.n841 185
R768 vdd.n2882 vdd.n840 185
R769 vdd.n3103 vdd.n840 185
R770 vdd.n2884 vdd.n2883 185
R771 vdd.n2883 vdd.n848 185
R772 vdd.n2885 vdd.n847 185
R773 vdd.n3097 vdd.n847 185
R774 vdd.n2887 vdd.n2886 185
R775 vdd.n2886 vdd.n845 185
R776 vdd.n2888 vdd.n854 185
R777 vdd.n3091 vdd.n854 185
R778 vdd.n2890 vdd.n2889 185
R779 vdd.n2889 vdd.n852 185
R780 vdd.n2891 vdd.n860 185
R781 vdd.n3085 vdd.n860 185
R782 vdd.n2893 vdd.n2892 185
R783 vdd.n2892 vdd.n858 185
R784 vdd.n2894 vdd.n865 185
R785 vdd.n3079 vdd.n865 185
R786 vdd.n2896 vdd.n2895 185
R787 vdd.n2895 vdd.n872 185
R788 vdd.n2897 vdd.n871 185
R789 vdd.n3073 vdd.n871 185
R790 vdd.n2899 vdd.n2898 185
R791 vdd.n2898 vdd.n879 185
R792 vdd.n2900 vdd.n878 185
R793 vdd.n3067 vdd.n878 185
R794 vdd.n2902 vdd.n2901 185
R795 vdd.n2901 vdd.n876 185
R796 vdd.n2903 vdd.n885 185
R797 vdd.n3060 vdd.n885 185
R798 vdd.n2905 vdd.n2904 185
R799 vdd.n2904 vdd.n883 185
R800 vdd.n2906 vdd.n890 185
R801 vdd.n3054 vdd.n890 185
R802 vdd.n2908 vdd.n2907 185
R803 vdd.n2907 vdd.n896 185
R804 vdd.n2909 vdd.n895 185
R805 vdd.n3048 vdd.n895 185
R806 vdd.n2911 vdd.n2910 185
R807 vdd.n2910 vdd.n902 185
R808 vdd.n2912 vdd.n901 185
R809 vdd.n3042 vdd.n901 185
R810 vdd.n2914 vdd.n2913 185
R811 vdd.n2915 vdd.n2914 185
R812 vdd.n2815 vdd.n907 185
R813 vdd.n3036 vdd.n907 185
R814 vdd.n2923 vdd.n2922 185
R815 vdd.n2922 vdd.n2921 185
R816 vdd.n2924 vdd.n913 185
R817 vdd.n3030 vdd.n913 185
R818 vdd.n2926 vdd.n2925 185
R819 vdd.n2925 vdd.n911 185
R820 vdd.n2927 vdd.n919 185
R821 vdd.n3024 vdd.n919 185
R822 vdd.n2929 vdd.n2928 185
R823 vdd.n2928 vdd.n917 185
R824 vdd.n2930 vdd.n924 185
R825 vdd.n3018 vdd.n924 185
R826 vdd.n2932 vdd.n2931 185
R827 vdd.n2933 vdd.n2932 185
R828 vdd.n2814 vdd.n930 185
R829 vdd.n3012 vdd.n930 185
R830 vdd.n2813 vdd.n2812 185
R831 vdd.n2812 vdd.n928 185
R832 vdd.n2274 vdd.n2273 185
R833 vdd.n2275 vdd.n2274 185
R834 vdd.n1503 vdd.n1501 185
R835 vdd.n1501 vdd.n1500 185
R836 vdd.n2269 vdd.n2268 185
R837 vdd.n2268 vdd.n2267 185
R838 vdd.n1506 vdd.n1505 185
R839 vdd.n1507 vdd.n1506 185
R840 vdd.n2256 vdd.n2255 185
R841 vdd.n2257 vdd.n2256 185
R842 vdd.n1515 vdd.n1514 185
R843 vdd.n2248 vdd.n1514 185
R844 vdd.n2251 vdd.n2250 185
R845 vdd.n2250 vdd.n2249 185
R846 vdd.n1518 vdd.n1517 185
R847 vdd.n1524 vdd.n1518 185
R848 vdd.n2239 vdd.n2238 185
R849 vdd.n2240 vdd.n2239 185
R850 vdd.n1526 vdd.n1525 185
R851 vdd.n2231 vdd.n1525 185
R852 vdd.n2234 vdd.n2233 185
R853 vdd.n2233 vdd.n2232 185
R854 vdd.n1529 vdd.n1528 185
R855 vdd.n1530 vdd.n1529 185
R856 vdd.n2222 vdd.n2221 185
R857 vdd.n2223 vdd.n2222 185
R858 vdd.n1538 vdd.n1537 185
R859 vdd.n1537 vdd.n1536 185
R860 vdd.n2217 vdd.n2216 185
R861 vdd.n2216 vdd.n2215 185
R862 vdd.n1541 vdd.n1540 185
R863 vdd.n1547 vdd.n1541 185
R864 vdd.n2206 vdd.n2205 185
R865 vdd.n2207 vdd.n2206 185
R866 vdd.n1549 vdd.n1548 185
R867 vdd.n1903 vdd.n1548 185
R868 vdd.n1906 vdd.n1905 185
R869 vdd.n1905 vdd.n1904 185
R870 vdd.n1552 vdd.n1551 185
R871 vdd.n1559 vdd.n1552 185
R872 vdd.n1894 vdd.n1893 185
R873 vdd.n1895 vdd.n1894 185
R874 vdd.n1561 vdd.n1560 185
R875 vdd.n1560 vdd.n1558 185
R876 vdd.n1889 vdd.n1888 185
R877 vdd.n1888 vdd.n1887 185
R878 vdd.n1564 vdd.n1563 185
R879 vdd.n1565 vdd.n1564 185
R880 vdd.n1878 vdd.n1877 185
R881 vdd.n1879 vdd.n1878 185
R882 vdd.n1572 vdd.n1571 185
R883 vdd.n1870 vdd.n1571 185
R884 vdd.n1873 vdd.n1872 185
R885 vdd.n1872 vdd.n1871 185
R886 vdd.n1575 vdd.n1574 185
R887 vdd.n1581 vdd.n1575 185
R888 vdd.n1861 vdd.n1860 185
R889 vdd.n1862 vdd.n1861 185
R890 vdd.n1583 vdd.n1582 185
R891 vdd.n1853 vdd.n1582 185
R892 vdd.n1856 vdd.n1855 185
R893 vdd.n1855 vdd.n1854 185
R894 vdd.n1586 vdd.n1585 185
R895 vdd.n1587 vdd.n1586 185
R896 vdd.n1844 vdd.n1843 185
R897 vdd.n1845 vdd.n1844 185
R898 vdd.n1595 vdd.n1594 185
R899 vdd.n1594 vdd.n1593 185
R900 vdd.n1839 vdd.n1838 185
R901 vdd.n1838 vdd.n1837 185
R902 vdd.n1598 vdd.n1597 185
R903 vdd.n1599 vdd.n1598 185
R904 vdd.n1827 vdd.n1826 185
R905 vdd.n1825 vdd.n1638 185
R906 vdd.n1640 vdd.n1637 185
R907 vdd.n1829 vdd.n1637 185
R908 vdd.n1821 vdd.n1642 185
R909 vdd.n1820 vdd.n1643 185
R910 vdd.n1819 vdd.n1644 185
R911 vdd.n1647 vdd.n1645 185
R912 vdd.n1815 vdd.n1648 185
R913 vdd.n1814 vdd.n1649 185
R914 vdd.n1813 vdd.n1650 185
R915 vdd.n1653 vdd.n1651 185
R916 vdd.n1809 vdd.n1654 185
R917 vdd.n1808 vdd.n1655 185
R918 vdd.n1807 vdd.n1656 185
R919 vdd.n1659 vdd.n1657 185
R920 vdd.n1803 vdd.n1660 185
R921 vdd.n1802 vdd.n1661 185
R922 vdd.n1801 vdd.n1662 185
R923 vdd.n1793 vdd.n1663 185
R924 vdd.n1797 vdd.n1794 185
R925 vdd.n1792 vdd.n1665 185
R926 vdd.n1791 vdd.n1666 185
R927 vdd.n1669 vdd.n1667 185
R928 vdd.n1787 vdd.n1670 185
R929 vdd.n1786 vdd.n1671 185
R930 vdd.n1785 vdd.n1672 185
R931 vdd.n1675 vdd.n1673 185
R932 vdd.n1781 vdd.n1676 185
R933 vdd.n1780 vdd.n1677 185
R934 vdd.n1779 vdd.n1678 185
R935 vdd.n1681 vdd.n1679 185
R936 vdd.n1775 vdd.n1682 185
R937 vdd.n1774 vdd.n1683 185
R938 vdd.n1773 vdd.n1684 185
R939 vdd.n1687 vdd.n1685 185
R940 vdd.n1769 vdd.n1688 185
R941 vdd.n1768 vdd.n1689 185
R942 vdd.n1767 vdd.n1690 185
R943 vdd.n1693 vdd.n1691 185
R944 vdd.n1763 vdd.n1694 185
R945 vdd.n1762 vdd.n1695 185
R946 vdd.n1761 vdd.n1758 185
R947 vdd.n1698 vdd.n1696 185
R948 vdd.n1754 vdd.n1699 185
R949 vdd.n1753 vdd.n1700 185
R950 vdd.n1752 vdd.n1701 185
R951 vdd.n1704 vdd.n1702 185
R952 vdd.n1748 vdd.n1705 185
R953 vdd.n1747 vdd.n1706 185
R954 vdd.n1746 vdd.n1707 185
R955 vdd.n1710 vdd.n1708 185
R956 vdd.n1742 vdd.n1711 185
R957 vdd.n1741 vdd.n1712 185
R958 vdd.n1740 vdd.n1713 185
R959 vdd.n1716 vdd.n1714 185
R960 vdd.n1736 vdd.n1717 185
R961 vdd.n1735 vdd.n1718 185
R962 vdd.n1734 vdd.n1719 185
R963 vdd.n1722 vdd.n1720 185
R964 vdd.n1730 vdd.n1723 185
R965 vdd.n1729 vdd.n1724 185
R966 vdd.n1728 vdd.n1725 185
R967 vdd.n1726 vdd.n1606 185
R968 vdd.n1831 vdd.n1830 185
R969 vdd.n1830 vdd.n1829 185
R970 vdd.n2278 vdd.n2277 185
R971 vdd.n2282 vdd.n1496 185
R972 vdd.n1495 vdd.n1489 185
R973 vdd.n1493 vdd.n1492 185
R974 vdd.n1491 vdd.n1250 185
R975 vdd.n2286 vdd.n1247 185
R976 vdd.n2288 vdd.n2287 185
R977 vdd.n2290 vdd.n1245 185
R978 vdd.n2292 vdd.n2291 185
R979 vdd.n2293 vdd.n1240 185
R980 vdd.n2295 vdd.n2294 185
R981 vdd.n2297 vdd.n1238 185
R982 vdd.n2299 vdd.n2298 185
R983 vdd.n2300 vdd.n1233 185
R984 vdd.n2302 vdd.n2301 185
R985 vdd.n2304 vdd.n1231 185
R986 vdd.n2306 vdd.n2305 185
R987 vdd.n2307 vdd.n1227 185
R988 vdd.n2309 vdd.n2308 185
R989 vdd.n2311 vdd.n1224 185
R990 vdd.n2313 vdd.n2312 185
R991 vdd.n1225 vdd.n1218 185
R992 vdd.n2317 vdd.n1222 185
R993 vdd.n2318 vdd.n1214 185
R994 vdd.n2320 vdd.n2319 185
R995 vdd.n2322 vdd.n1212 185
R996 vdd.n2324 vdd.n2323 185
R997 vdd.n2325 vdd.n1207 185
R998 vdd.n2327 vdd.n2326 185
R999 vdd.n2329 vdd.n1205 185
R1000 vdd.n2331 vdd.n2330 185
R1001 vdd.n2332 vdd.n1200 185
R1002 vdd.n2334 vdd.n2333 185
R1003 vdd.n2336 vdd.n1198 185
R1004 vdd.n2338 vdd.n2337 185
R1005 vdd.n2339 vdd.n1193 185
R1006 vdd.n2341 vdd.n2340 185
R1007 vdd.n2343 vdd.n1191 185
R1008 vdd.n2345 vdd.n2344 185
R1009 vdd.n2346 vdd.n1187 185
R1010 vdd.n2348 vdd.n2347 185
R1011 vdd.n2350 vdd.n1184 185
R1012 vdd.n2352 vdd.n2351 185
R1013 vdd.n1185 vdd.n1178 185
R1014 vdd.n2356 vdd.n1182 185
R1015 vdd.n2357 vdd.n1174 185
R1016 vdd.n2359 vdd.n2358 185
R1017 vdd.n2361 vdd.n1172 185
R1018 vdd.n2363 vdd.n2362 185
R1019 vdd.n2364 vdd.n1167 185
R1020 vdd.n2366 vdd.n2365 185
R1021 vdd.n2368 vdd.n1165 185
R1022 vdd.n2370 vdd.n2369 185
R1023 vdd.n2371 vdd.n1160 185
R1024 vdd.n2373 vdd.n2372 185
R1025 vdd.n2375 vdd.n1158 185
R1026 vdd.n2377 vdd.n2376 185
R1027 vdd.n2378 vdd.n1156 185
R1028 vdd.n2380 vdd.n2379 185
R1029 vdd.n2383 vdd.n2382 185
R1030 vdd.n2385 vdd.n2384 185
R1031 vdd.n2387 vdd.n1154 185
R1032 vdd.n2389 vdd.n2388 185
R1033 vdd.n1502 vdd.n1153 185
R1034 vdd.n2276 vdd.n1499 185
R1035 vdd.n2276 vdd.n2275 185
R1036 vdd.n1510 vdd.n1498 185
R1037 vdd.n1500 vdd.n1498 185
R1038 vdd.n2266 vdd.n2265 185
R1039 vdd.n2267 vdd.n2266 185
R1040 vdd.n1509 vdd.n1508 185
R1041 vdd.n1508 vdd.n1507 185
R1042 vdd.n2259 vdd.n2258 185
R1043 vdd.n2258 vdd.n2257 185
R1044 vdd.n1513 vdd.n1512 185
R1045 vdd.n2248 vdd.n1513 185
R1046 vdd.n2247 vdd.n2246 185
R1047 vdd.n2249 vdd.n2247 185
R1048 vdd.n1520 vdd.n1519 185
R1049 vdd.n1524 vdd.n1519 185
R1050 vdd.n2242 vdd.n2241 185
R1051 vdd.n2241 vdd.n2240 185
R1052 vdd.n1523 vdd.n1522 185
R1053 vdd.n2231 vdd.n1523 185
R1054 vdd.n2230 vdd.n2229 185
R1055 vdd.n2232 vdd.n2230 185
R1056 vdd.n1532 vdd.n1531 185
R1057 vdd.n1531 vdd.n1530 185
R1058 vdd.n2225 vdd.n2224 185
R1059 vdd.n2224 vdd.n2223 185
R1060 vdd.n1535 vdd.n1534 185
R1061 vdd.n1536 vdd.n1535 185
R1062 vdd.n2214 vdd.n2213 185
R1063 vdd.n2215 vdd.n2214 185
R1064 vdd.n1543 vdd.n1542 185
R1065 vdd.n1547 vdd.n1542 185
R1066 vdd.n2209 vdd.n2208 185
R1067 vdd.n2208 vdd.n2207 185
R1068 vdd.n1546 vdd.n1545 185
R1069 vdd.n1903 vdd.n1546 185
R1070 vdd.n1902 vdd.n1901 185
R1071 vdd.n1904 vdd.n1902 185
R1072 vdd.n1554 vdd.n1553 185
R1073 vdd.n1559 vdd.n1553 185
R1074 vdd.n1897 vdd.n1896 185
R1075 vdd.n1896 vdd.n1895 185
R1076 vdd.n1557 vdd.n1556 185
R1077 vdd.n1558 vdd.n1557 185
R1078 vdd.n1886 vdd.n1885 185
R1079 vdd.n1887 vdd.n1886 185
R1080 vdd.n1567 vdd.n1566 185
R1081 vdd.n1566 vdd.n1565 185
R1082 vdd.n1881 vdd.n1880 185
R1083 vdd.n1880 vdd.n1879 185
R1084 vdd.n1570 vdd.n1569 185
R1085 vdd.n1870 vdd.n1570 185
R1086 vdd.n1869 vdd.n1868 185
R1087 vdd.n1871 vdd.n1869 185
R1088 vdd.n1577 vdd.n1576 185
R1089 vdd.n1581 vdd.n1576 185
R1090 vdd.n1864 vdd.n1863 185
R1091 vdd.n1863 vdd.n1862 185
R1092 vdd.n1580 vdd.n1579 185
R1093 vdd.n1853 vdd.n1580 185
R1094 vdd.n1852 vdd.n1851 185
R1095 vdd.n1854 vdd.n1852 185
R1096 vdd.n1589 vdd.n1588 185
R1097 vdd.n1588 vdd.n1587 185
R1098 vdd.n1847 vdd.n1846 185
R1099 vdd.n1846 vdd.n1845 185
R1100 vdd.n1592 vdd.n1591 185
R1101 vdd.n1593 vdd.n1592 185
R1102 vdd.n1836 vdd.n1835 185
R1103 vdd.n1837 vdd.n1836 185
R1104 vdd.n1601 vdd.n1600 185
R1105 vdd.n1600 vdd.n1599 185
R1106 vdd.n971 vdd.n969 185
R1107 vdd.n2629 vdd.n969 185
R1108 vdd.n2551 vdd.n989 185
R1109 vdd.n989 vdd.n976 185
R1110 vdd.n2553 vdd.n2552 185
R1111 vdd.n2554 vdd.n2553 185
R1112 vdd.n2550 vdd.n988 185
R1113 vdd.n1370 vdd.n988 185
R1114 vdd.n2549 vdd.n2548 185
R1115 vdd.n2548 vdd.n2547 185
R1116 vdd.n991 vdd.n990 185
R1117 vdd.n992 vdd.n991 185
R1118 vdd.n2538 vdd.n2537 185
R1119 vdd.n2539 vdd.n2538 185
R1120 vdd.n2536 vdd.n1002 185
R1121 vdd.n1002 vdd.n999 185
R1122 vdd.n2535 vdd.n2534 185
R1123 vdd.n2534 vdd.n2533 185
R1124 vdd.n1004 vdd.n1003 185
R1125 vdd.n1396 vdd.n1004 185
R1126 vdd.n2526 vdd.n2525 185
R1127 vdd.n2527 vdd.n2526 185
R1128 vdd.n2524 vdd.n1012 185
R1129 vdd.n1017 vdd.n1012 185
R1130 vdd.n2523 vdd.n2522 185
R1131 vdd.n2522 vdd.n2521 185
R1132 vdd.n1014 vdd.n1013 185
R1133 vdd.n1023 vdd.n1014 185
R1134 vdd.n2514 vdd.n2513 185
R1135 vdd.n2515 vdd.n2514 185
R1136 vdd.n2512 vdd.n1024 185
R1137 vdd.n1408 vdd.n1024 185
R1138 vdd.n2511 vdd.n2510 185
R1139 vdd.n2510 vdd.n2509 185
R1140 vdd.n1026 vdd.n1025 185
R1141 vdd.n1027 vdd.n1026 185
R1142 vdd.n2502 vdd.n2501 185
R1143 vdd.n2503 vdd.n2502 185
R1144 vdd.n2500 vdd.n1036 185
R1145 vdd.n1036 vdd.n1033 185
R1146 vdd.n2499 vdd.n2498 185
R1147 vdd.n2498 vdd.n2497 185
R1148 vdd.n1038 vdd.n1037 185
R1149 vdd.n1047 vdd.n1038 185
R1150 vdd.n2489 vdd.n2488 185
R1151 vdd.n2490 vdd.n2489 185
R1152 vdd.n2487 vdd.n1048 185
R1153 vdd.n1054 vdd.n1048 185
R1154 vdd.n2486 vdd.n2485 185
R1155 vdd.n2485 vdd.n2484 185
R1156 vdd.n1050 vdd.n1049 185
R1157 vdd.n1051 vdd.n1050 185
R1158 vdd.n2477 vdd.n2476 185
R1159 vdd.n2478 vdd.n2477 185
R1160 vdd.n2475 vdd.n1061 185
R1161 vdd.n1061 vdd.n1058 185
R1162 vdd.n2474 vdd.n2473 185
R1163 vdd.n2473 vdd.n2472 185
R1164 vdd.n1063 vdd.n1062 185
R1165 vdd.n1064 vdd.n1063 185
R1166 vdd.n2465 vdd.n2464 185
R1167 vdd.n2466 vdd.n2465 185
R1168 vdd.n2463 vdd.n1072 185
R1169 vdd.n1077 vdd.n1072 185
R1170 vdd.n2462 vdd.n2461 185
R1171 vdd.n2461 vdd.n2460 185
R1172 vdd.n1074 vdd.n1073 185
R1173 vdd.n1083 vdd.n1074 185
R1174 vdd.n2453 vdd.n2452 185
R1175 vdd.n2454 vdd.n2453 185
R1176 vdd.n2451 vdd.n1084 185
R1177 vdd.n1090 vdd.n1084 185
R1178 vdd.n2450 vdd.n2449 185
R1179 vdd.n2449 vdd.n2448 185
R1180 vdd.n1086 vdd.n1085 185
R1181 vdd.n1087 vdd.n1086 185
R1182 vdd.n2441 vdd.n2440 185
R1183 vdd.n2442 vdd.n2441 185
R1184 vdd.n2439 vdd.n1097 185
R1185 vdd.n1097 vdd.n1094 185
R1186 vdd.n2438 vdd.n2437 185
R1187 vdd.n2437 vdd.n2436 185
R1188 vdd.n1099 vdd.n1098 185
R1189 vdd.n1108 vdd.n1099 185
R1190 vdd.n2429 vdd.n2428 185
R1191 vdd.n2430 vdd.n2429 185
R1192 vdd.n2427 vdd.n1109 185
R1193 vdd.n1109 vdd.n1105 185
R1194 vdd.n2426 vdd.n2425 185
R1195 vdd.n1111 vdd.n1110 185
R1196 vdd.n2422 vdd.n2421 185
R1197 vdd.n2423 vdd.n2422 185
R1198 vdd.n2420 vdd.n1147 185
R1199 vdd.n2419 vdd.n2418 185
R1200 vdd.n2417 vdd.n2416 185
R1201 vdd.n2415 vdd.n2414 185
R1202 vdd.n2413 vdd.n2412 185
R1203 vdd.n2411 vdd.n2410 185
R1204 vdd.n2409 vdd.n2408 185
R1205 vdd.n2407 vdd.n2406 185
R1206 vdd.n2405 vdd.n2404 185
R1207 vdd.n2403 vdd.n2402 185
R1208 vdd.n2401 vdd.n2400 185
R1209 vdd.n2399 vdd.n2398 185
R1210 vdd.n2397 vdd.n2396 185
R1211 vdd.n2395 vdd.n2394 185
R1212 vdd.n2393 vdd.n2392 185
R1213 vdd.n1292 vdd.n1148 185
R1214 vdd.n1294 vdd.n1293 185
R1215 vdd.n1296 vdd.n1295 185
R1216 vdd.n1298 vdd.n1297 185
R1217 vdd.n1300 vdd.n1299 185
R1218 vdd.n1302 vdd.n1301 185
R1219 vdd.n1304 vdd.n1303 185
R1220 vdd.n1306 vdd.n1305 185
R1221 vdd.n1308 vdd.n1307 185
R1222 vdd.n1310 vdd.n1309 185
R1223 vdd.n1312 vdd.n1311 185
R1224 vdd.n1314 vdd.n1313 185
R1225 vdd.n1316 vdd.n1315 185
R1226 vdd.n1318 vdd.n1317 185
R1227 vdd.n1321 vdd.n1320 185
R1228 vdd.n1323 vdd.n1322 185
R1229 vdd.n1325 vdd.n1324 185
R1230 vdd.n2632 vdd.n2631 185
R1231 vdd.n2634 vdd.n2633 185
R1232 vdd.n2636 vdd.n2635 185
R1233 vdd.n2639 vdd.n2638 185
R1234 vdd.n2641 vdd.n2640 185
R1235 vdd.n2643 vdd.n2642 185
R1236 vdd.n2645 vdd.n2644 185
R1237 vdd.n2647 vdd.n2646 185
R1238 vdd.n2649 vdd.n2648 185
R1239 vdd.n2651 vdd.n2650 185
R1240 vdd.n2653 vdd.n2652 185
R1241 vdd.n2655 vdd.n2654 185
R1242 vdd.n2657 vdd.n2656 185
R1243 vdd.n2659 vdd.n2658 185
R1244 vdd.n2661 vdd.n2660 185
R1245 vdd.n2663 vdd.n2662 185
R1246 vdd.n2665 vdd.n2664 185
R1247 vdd.n2667 vdd.n2666 185
R1248 vdd.n2669 vdd.n2668 185
R1249 vdd.n2671 vdd.n2670 185
R1250 vdd.n2673 vdd.n2672 185
R1251 vdd.n2675 vdd.n2674 185
R1252 vdd.n2677 vdd.n2676 185
R1253 vdd.n2679 vdd.n2678 185
R1254 vdd.n2681 vdd.n2680 185
R1255 vdd.n2683 vdd.n2682 185
R1256 vdd.n2685 vdd.n2684 185
R1257 vdd.n2687 vdd.n2686 185
R1258 vdd.n2689 vdd.n2688 185
R1259 vdd.n2691 vdd.n2690 185
R1260 vdd.n2693 vdd.n2692 185
R1261 vdd.n2695 vdd.n2694 185
R1262 vdd.n2697 vdd.n2696 185
R1263 vdd.n2698 vdd.n970 185
R1264 vdd.n2700 vdd.n2699 185
R1265 vdd.n2701 vdd.n2700 185
R1266 vdd.n2630 vdd.n974 185
R1267 vdd.n2630 vdd.n2629 185
R1268 vdd.n1368 vdd.n975 185
R1269 vdd.n976 vdd.n975 185
R1270 vdd.n1369 vdd.n986 185
R1271 vdd.n2554 vdd.n986 185
R1272 vdd.n1372 vdd.n1371 185
R1273 vdd.n1371 vdd.n1370 185
R1274 vdd.n1373 vdd.n993 185
R1275 vdd.n2547 vdd.n993 185
R1276 vdd.n1375 vdd.n1374 185
R1277 vdd.n1374 vdd.n992 185
R1278 vdd.n1376 vdd.n1000 185
R1279 vdd.n2539 vdd.n1000 185
R1280 vdd.n1378 vdd.n1377 185
R1281 vdd.n1377 vdd.n999 185
R1282 vdd.n1379 vdd.n1005 185
R1283 vdd.n2533 vdd.n1005 185
R1284 vdd.n1398 vdd.n1397 185
R1285 vdd.n1397 vdd.n1396 185
R1286 vdd.n1399 vdd.n1010 185
R1287 vdd.n2527 vdd.n1010 185
R1288 vdd.n1401 vdd.n1400 185
R1289 vdd.n1400 vdd.n1017 185
R1290 vdd.n1402 vdd.n1015 185
R1291 vdd.n2521 vdd.n1015 185
R1292 vdd.n1404 vdd.n1403 185
R1293 vdd.n1403 vdd.n1023 185
R1294 vdd.n1405 vdd.n1021 185
R1295 vdd.n2515 vdd.n1021 185
R1296 vdd.n1407 vdd.n1406 185
R1297 vdd.n1408 vdd.n1407 185
R1298 vdd.n1367 vdd.n1028 185
R1299 vdd.n2509 vdd.n1028 185
R1300 vdd.n1366 vdd.n1365 185
R1301 vdd.n1365 vdd.n1027 185
R1302 vdd.n1364 vdd.n1034 185
R1303 vdd.n2503 vdd.n1034 185
R1304 vdd.n1363 vdd.n1362 185
R1305 vdd.n1362 vdd.n1033 185
R1306 vdd.n1361 vdd.n1039 185
R1307 vdd.n2497 vdd.n1039 185
R1308 vdd.n1360 vdd.n1359 185
R1309 vdd.n1359 vdd.n1047 185
R1310 vdd.n1358 vdd.n1045 185
R1311 vdd.n2490 vdd.n1045 185
R1312 vdd.n1357 vdd.n1356 185
R1313 vdd.n1356 vdd.n1054 185
R1314 vdd.n1355 vdd.n1052 185
R1315 vdd.n2484 vdd.n1052 185
R1316 vdd.n1354 vdd.n1353 185
R1317 vdd.n1353 vdd.n1051 185
R1318 vdd.n1352 vdd.n1059 185
R1319 vdd.n2478 vdd.n1059 185
R1320 vdd.n1351 vdd.n1350 185
R1321 vdd.n1350 vdd.n1058 185
R1322 vdd.n1349 vdd.n1065 185
R1323 vdd.n2472 vdd.n1065 185
R1324 vdd.n1348 vdd.n1347 185
R1325 vdd.n1347 vdd.n1064 185
R1326 vdd.n1346 vdd.n1070 185
R1327 vdd.n2466 vdd.n1070 185
R1328 vdd.n1345 vdd.n1344 185
R1329 vdd.n1344 vdd.n1077 185
R1330 vdd.n1343 vdd.n1075 185
R1331 vdd.n2460 vdd.n1075 185
R1332 vdd.n1342 vdd.n1341 185
R1333 vdd.n1341 vdd.n1083 185
R1334 vdd.n1340 vdd.n1081 185
R1335 vdd.n2454 vdd.n1081 185
R1336 vdd.n1339 vdd.n1338 185
R1337 vdd.n1338 vdd.n1090 185
R1338 vdd.n1337 vdd.n1088 185
R1339 vdd.n2448 vdd.n1088 185
R1340 vdd.n1336 vdd.n1335 185
R1341 vdd.n1335 vdd.n1087 185
R1342 vdd.n1334 vdd.n1095 185
R1343 vdd.n2442 vdd.n1095 185
R1344 vdd.n1333 vdd.n1332 185
R1345 vdd.n1332 vdd.n1094 185
R1346 vdd.n1331 vdd.n1100 185
R1347 vdd.n2436 vdd.n1100 185
R1348 vdd.n1330 vdd.n1329 185
R1349 vdd.n1329 vdd.n1108 185
R1350 vdd.n1328 vdd.n1106 185
R1351 vdd.n2430 vdd.n1106 185
R1352 vdd.n1327 vdd.n1326 185
R1353 vdd.n1326 vdd.n1105 185
R1354 vdd.n370 vdd.n369 185
R1355 vdd.n3526 vdd.n370 185
R1356 vdd.n3529 vdd.n3528 185
R1357 vdd.n3528 vdd.n3527 185
R1358 vdd.n3530 vdd.n364 185
R1359 vdd.n364 vdd.n363 185
R1360 vdd.n3532 vdd.n3531 185
R1361 vdd.n3533 vdd.n3532 185
R1362 vdd.n359 vdd.n358 185
R1363 vdd.n3534 vdd.n359 185
R1364 vdd.n3537 vdd.n3536 185
R1365 vdd.n3536 vdd.n3535 185
R1366 vdd.n3538 vdd.n353 185
R1367 vdd.n3508 vdd.n353 185
R1368 vdd.n3540 vdd.n3539 185
R1369 vdd.n3541 vdd.n3540 185
R1370 vdd.n348 vdd.n347 185
R1371 vdd.n3542 vdd.n348 185
R1372 vdd.n3545 vdd.n3544 185
R1373 vdd.n3544 vdd.n3543 185
R1374 vdd.n3546 vdd.n342 185
R1375 vdd.n349 vdd.n342 185
R1376 vdd.n3548 vdd.n3547 185
R1377 vdd.n3549 vdd.n3548 185
R1378 vdd.n338 vdd.n337 185
R1379 vdd.n3550 vdd.n338 185
R1380 vdd.n3553 vdd.n3552 185
R1381 vdd.n3552 vdd.n3551 185
R1382 vdd.n3554 vdd.n333 185
R1383 vdd.n333 vdd.n332 185
R1384 vdd.n3556 vdd.n3555 185
R1385 vdd.n3557 vdd.n3556 185
R1386 vdd.n327 vdd.n325 185
R1387 vdd.n3558 vdd.n327 185
R1388 vdd.n3561 vdd.n3560 185
R1389 vdd.n3560 vdd.n3559 185
R1390 vdd.n326 vdd.n324 185
R1391 vdd.n328 vdd.n326 185
R1392 vdd.n3484 vdd.n3483 185
R1393 vdd.n3485 vdd.n3484 185
R1394 vdd.n615 vdd.n614 185
R1395 vdd.n614 vdd.n613 185
R1396 vdd.n3479 vdd.n3478 185
R1397 vdd.n3478 vdd.n3477 185
R1398 vdd.n618 vdd.n617 185
R1399 vdd.n624 vdd.n618 185
R1400 vdd.n3465 vdd.n3464 185
R1401 vdd.n3466 vdd.n3465 185
R1402 vdd.n626 vdd.n625 185
R1403 vdd.n3457 vdd.n625 185
R1404 vdd.n3460 vdd.n3459 185
R1405 vdd.n3459 vdd.n3458 185
R1406 vdd.n629 vdd.n628 185
R1407 vdd.n636 vdd.n629 185
R1408 vdd.n3448 vdd.n3447 185
R1409 vdd.n3449 vdd.n3448 185
R1410 vdd.n638 vdd.n637 185
R1411 vdd.n637 vdd.n635 185
R1412 vdd.n3443 vdd.n3442 185
R1413 vdd.n3442 vdd.n3441 185
R1414 vdd.n641 vdd.n640 185
R1415 vdd.n642 vdd.n641 185
R1416 vdd.n3432 vdd.n3431 185
R1417 vdd.n3433 vdd.n3432 185
R1418 vdd.n650 vdd.n649 185
R1419 vdd.n649 vdd.n648 185
R1420 vdd.n3427 vdd.n3426 185
R1421 vdd.n3426 vdd.n3425 185
R1422 vdd.n653 vdd.n652 185
R1423 vdd.n659 vdd.n653 185
R1424 vdd.n3416 vdd.n3415 185
R1425 vdd.n3417 vdd.n3416 185
R1426 vdd.n3412 vdd.n660 185
R1427 vdd.n3411 vdd.n3410 185
R1428 vdd.n3408 vdd.n662 185
R1429 vdd.n3408 vdd.n658 185
R1430 vdd.n3407 vdd.n3406 185
R1431 vdd.n3405 vdd.n3404 185
R1432 vdd.n3403 vdd.n3402 185
R1433 vdd.n3401 vdd.n3400 185
R1434 vdd.n3399 vdd.n668 185
R1435 vdd.n3397 vdd.n3396 185
R1436 vdd.n3395 vdd.n669 185
R1437 vdd.n3394 vdd.n3393 185
R1438 vdd.n3391 vdd.n674 185
R1439 vdd.n3389 vdd.n3388 185
R1440 vdd.n3387 vdd.n675 185
R1441 vdd.n3386 vdd.n3385 185
R1442 vdd.n3383 vdd.n680 185
R1443 vdd.n3381 vdd.n3380 185
R1444 vdd.n3379 vdd.n681 185
R1445 vdd.n3378 vdd.n3377 185
R1446 vdd.n3375 vdd.n688 185
R1447 vdd.n3373 vdd.n3372 185
R1448 vdd.n3371 vdd.n689 185
R1449 vdd.n3370 vdd.n3369 185
R1450 vdd.n3367 vdd.n694 185
R1451 vdd.n3365 vdd.n3364 185
R1452 vdd.n3363 vdd.n695 185
R1453 vdd.n3362 vdd.n3361 185
R1454 vdd.n3359 vdd.n700 185
R1455 vdd.n3357 vdd.n3356 185
R1456 vdd.n3355 vdd.n701 185
R1457 vdd.n3354 vdd.n3353 185
R1458 vdd.n3351 vdd.n706 185
R1459 vdd.n3349 vdd.n3348 185
R1460 vdd.n3347 vdd.n707 185
R1461 vdd.n3346 vdd.n3345 185
R1462 vdd.n3343 vdd.n712 185
R1463 vdd.n3341 vdd.n3340 185
R1464 vdd.n3339 vdd.n713 185
R1465 vdd.n3338 vdd.n3337 185
R1466 vdd.n3335 vdd.n718 185
R1467 vdd.n3333 vdd.n3332 185
R1468 vdd.n3331 vdd.n719 185
R1469 vdd.n728 vdd.n722 185
R1470 vdd.n3327 vdd.n3326 185
R1471 vdd.n3324 vdd.n726 185
R1472 vdd.n3323 vdd.n3322 185
R1473 vdd.n3321 vdd.n3320 185
R1474 vdd.n3319 vdd.n732 185
R1475 vdd.n3317 vdd.n3316 185
R1476 vdd.n3315 vdd.n733 185
R1477 vdd.n3314 vdd.n3313 185
R1478 vdd.n3311 vdd.n738 185
R1479 vdd.n3309 vdd.n3308 185
R1480 vdd.n3307 vdd.n739 185
R1481 vdd.n3306 vdd.n3305 185
R1482 vdd.n3303 vdd.n744 185
R1483 vdd.n3301 vdd.n3300 185
R1484 vdd.n3299 vdd.n745 185
R1485 vdd.n3298 vdd.n3297 185
R1486 vdd.n3295 vdd.n3294 185
R1487 vdd.n3293 vdd.n3292 185
R1488 vdd.n3291 vdd.n3290 185
R1489 vdd.n3289 vdd.n3288 185
R1490 vdd.n3284 vdd.n657 185
R1491 vdd.n658 vdd.n657 185
R1492 vdd.n3523 vdd.n3522 185
R1493 vdd.n599 vdd.n404 185
R1494 vdd.n598 vdd.n597 185
R1495 vdd.n596 vdd.n595 185
R1496 vdd.n594 vdd.n409 185
R1497 vdd.n590 vdd.n589 185
R1498 vdd.n588 vdd.n587 185
R1499 vdd.n586 vdd.n585 185
R1500 vdd.n584 vdd.n411 185
R1501 vdd.n580 vdd.n579 185
R1502 vdd.n578 vdd.n577 185
R1503 vdd.n576 vdd.n575 185
R1504 vdd.n574 vdd.n413 185
R1505 vdd.n570 vdd.n569 185
R1506 vdd.n568 vdd.n567 185
R1507 vdd.n566 vdd.n565 185
R1508 vdd.n564 vdd.n415 185
R1509 vdd.n560 vdd.n559 185
R1510 vdd.n558 vdd.n557 185
R1511 vdd.n556 vdd.n555 185
R1512 vdd.n554 vdd.n417 185
R1513 vdd.n550 vdd.n549 185
R1514 vdd.n548 vdd.n547 185
R1515 vdd.n546 vdd.n545 185
R1516 vdd.n544 vdd.n421 185
R1517 vdd.n540 vdd.n539 185
R1518 vdd.n538 vdd.n537 185
R1519 vdd.n536 vdd.n535 185
R1520 vdd.n534 vdd.n423 185
R1521 vdd.n530 vdd.n529 185
R1522 vdd.n528 vdd.n527 185
R1523 vdd.n526 vdd.n525 185
R1524 vdd.n524 vdd.n425 185
R1525 vdd.n520 vdd.n519 185
R1526 vdd.n518 vdd.n517 185
R1527 vdd.n516 vdd.n515 185
R1528 vdd.n514 vdd.n427 185
R1529 vdd.n510 vdd.n509 185
R1530 vdd.n508 vdd.n507 185
R1531 vdd.n506 vdd.n505 185
R1532 vdd.n504 vdd.n429 185
R1533 vdd.n500 vdd.n499 185
R1534 vdd.n498 vdd.n497 185
R1535 vdd.n496 vdd.n495 185
R1536 vdd.n494 vdd.n433 185
R1537 vdd.n490 vdd.n489 185
R1538 vdd.n488 vdd.n487 185
R1539 vdd.n486 vdd.n485 185
R1540 vdd.n484 vdd.n435 185
R1541 vdd.n480 vdd.n479 185
R1542 vdd.n478 vdd.n477 185
R1543 vdd.n476 vdd.n475 185
R1544 vdd.n474 vdd.n437 185
R1545 vdd.n470 vdd.n469 185
R1546 vdd.n468 vdd.n467 185
R1547 vdd.n466 vdd.n465 185
R1548 vdd.n464 vdd.n439 185
R1549 vdd.n460 vdd.n459 185
R1550 vdd.n458 vdd.n457 185
R1551 vdd.n456 vdd.n455 185
R1552 vdd.n454 vdd.n441 185
R1553 vdd.n450 vdd.n449 185
R1554 vdd.n448 vdd.n447 185
R1555 vdd.n446 vdd.n445 185
R1556 vdd.n3519 vdd.n372 185
R1557 vdd.n3526 vdd.n372 185
R1558 vdd.n3518 vdd.n371 185
R1559 vdd.n3527 vdd.n371 185
R1560 vdd.n3517 vdd.n3516 185
R1561 vdd.n3516 vdd.n363 185
R1562 vdd.n602 vdd.n362 185
R1563 vdd.n3533 vdd.n362 185
R1564 vdd.n3512 vdd.n361 185
R1565 vdd.n3534 vdd.n361 185
R1566 vdd.n3511 vdd.n360 185
R1567 vdd.n3535 vdd.n360 185
R1568 vdd.n3510 vdd.n3509 185
R1569 vdd.n3509 vdd.n3508 185
R1570 vdd.n604 vdd.n352 185
R1571 vdd.n3541 vdd.n352 185
R1572 vdd.n3504 vdd.n351 185
R1573 vdd.n3542 vdd.n351 185
R1574 vdd.n3503 vdd.n350 185
R1575 vdd.n3543 vdd.n350 185
R1576 vdd.n3502 vdd.n3501 185
R1577 vdd.n3501 vdd.n349 185
R1578 vdd.n606 vdd.n341 185
R1579 vdd.n3549 vdd.n341 185
R1580 vdd.n3497 vdd.n340 185
R1581 vdd.n3550 vdd.n340 185
R1582 vdd.n3496 vdd.n339 185
R1583 vdd.n3551 vdd.n339 185
R1584 vdd.n3495 vdd.n3494 185
R1585 vdd.n3494 vdd.n332 185
R1586 vdd.n608 vdd.n331 185
R1587 vdd.n3557 vdd.n331 185
R1588 vdd.n3490 vdd.n330 185
R1589 vdd.n3558 vdd.n330 185
R1590 vdd.n3489 vdd.n329 185
R1591 vdd.n3559 vdd.n329 185
R1592 vdd.n3488 vdd.n3487 185
R1593 vdd.n3487 vdd.n328 185
R1594 vdd.n3486 vdd.n610 185
R1595 vdd.n3486 vdd.n3485 185
R1596 vdd.n3474 vdd.n612 185
R1597 vdd.n613 vdd.n612 185
R1598 vdd.n3476 vdd.n3475 185
R1599 vdd.n3477 vdd.n3476 185
R1600 vdd.n620 vdd.n619 185
R1601 vdd.n624 vdd.n619 185
R1602 vdd.n3468 vdd.n3467 185
R1603 vdd.n3467 vdd.n3466 185
R1604 vdd.n623 vdd.n622 185
R1605 vdd.n3457 vdd.n623 185
R1606 vdd.n3456 vdd.n3455 185
R1607 vdd.n3458 vdd.n3456 185
R1608 vdd.n631 vdd.n630 185
R1609 vdd.n636 vdd.n630 185
R1610 vdd.n3451 vdd.n3450 185
R1611 vdd.n3450 vdd.n3449 185
R1612 vdd.n634 vdd.n633 185
R1613 vdd.n635 vdd.n634 185
R1614 vdd.n3440 vdd.n3439 185
R1615 vdd.n3441 vdd.n3440 185
R1616 vdd.n644 vdd.n643 185
R1617 vdd.n643 vdd.n642 185
R1618 vdd.n3435 vdd.n3434 185
R1619 vdd.n3434 vdd.n3433 185
R1620 vdd.n647 vdd.n646 185
R1621 vdd.n648 vdd.n647 185
R1622 vdd.n3424 vdd.n3423 185
R1623 vdd.n3425 vdd.n3424 185
R1624 vdd.n655 vdd.n654 185
R1625 vdd.n659 vdd.n654 185
R1626 vdd.n3419 vdd.n3418 185
R1627 vdd.n3418 vdd.n3417 185
R1628 vdd.n3008 vdd.n3007 185
R1629 vdd.n933 vdd.n932 185
R1630 vdd.n3004 vdd.n3003 185
R1631 vdd.n3005 vdd.n3004 185
R1632 vdd.n3002 vdd.n2736 185
R1633 vdd.n3001 vdd.n3000 185
R1634 vdd.n2999 vdd.n2998 185
R1635 vdd.n2997 vdd.n2996 185
R1636 vdd.n2995 vdd.n2994 185
R1637 vdd.n2993 vdd.n2992 185
R1638 vdd.n2991 vdd.n2990 185
R1639 vdd.n2989 vdd.n2988 185
R1640 vdd.n2987 vdd.n2986 185
R1641 vdd.n2985 vdd.n2984 185
R1642 vdd.n2983 vdd.n2982 185
R1643 vdd.n2981 vdd.n2980 185
R1644 vdd.n2979 vdd.n2978 185
R1645 vdd.n2977 vdd.n2976 185
R1646 vdd.n2975 vdd.n2974 185
R1647 vdd.n2973 vdd.n2972 185
R1648 vdd.n2971 vdd.n2970 185
R1649 vdd.n2969 vdd.n2968 185
R1650 vdd.n2967 vdd.n2966 185
R1651 vdd.n2965 vdd.n2964 185
R1652 vdd.n2963 vdd.n2962 185
R1653 vdd.n2961 vdd.n2960 185
R1654 vdd.n2959 vdd.n2958 185
R1655 vdd.n2957 vdd.n2956 185
R1656 vdd.n2955 vdd.n2954 185
R1657 vdd.n2953 vdd.n2952 185
R1658 vdd.n2951 vdd.n2950 185
R1659 vdd.n2949 vdd.n2948 185
R1660 vdd.n2947 vdd.n2946 185
R1661 vdd.n2944 vdd.n2943 185
R1662 vdd.n2942 vdd.n2941 185
R1663 vdd.n2940 vdd.n2939 185
R1664 vdd.n3185 vdd.n3184 185
R1665 vdd.n3186 vdd.n803 185
R1666 vdd.n3188 vdd.n3187 185
R1667 vdd.n3190 vdd.n801 185
R1668 vdd.n3192 vdd.n3191 185
R1669 vdd.n3193 vdd.n800 185
R1670 vdd.n3195 vdd.n3194 185
R1671 vdd.n3197 vdd.n798 185
R1672 vdd.n3199 vdd.n3198 185
R1673 vdd.n3200 vdd.n797 185
R1674 vdd.n3202 vdd.n3201 185
R1675 vdd.n3204 vdd.n795 185
R1676 vdd.n3206 vdd.n3205 185
R1677 vdd.n3207 vdd.n794 185
R1678 vdd.n3209 vdd.n3208 185
R1679 vdd.n3211 vdd.n792 185
R1680 vdd.n3213 vdd.n3212 185
R1681 vdd.n3215 vdd.n791 185
R1682 vdd.n3217 vdd.n3216 185
R1683 vdd.n3219 vdd.n789 185
R1684 vdd.n3221 vdd.n3220 185
R1685 vdd.n3222 vdd.n788 185
R1686 vdd.n3224 vdd.n3223 185
R1687 vdd.n3226 vdd.n786 185
R1688 vdd.n3228 vdd.n3227 185
R1689 vdd.n3229 vdd.n785 185
R1690 vdd.n3231 vdd.n3230 185
R1691 vdd.n3233 vdd.n783 185
R1692 vdd.n3235 vdd.n3234 185
R1693 vdd.n3236 vdd.n782 185
R1694 vdd.n3238 vdd.n3237 185
R1695 vdd.n3240 vdd.n781 185
R1696 vdd.n3241 vdd.n780 185
R1697 vdd.n3244 vdd.n3243 185
R1698 vdd.n3245 vdd.n778 185
R1699 vdd.n778 vdd.n756 185
R1700 vdd.n3182 vdd.n775 185
R1701 vdd.n3248 vdd.n775 185
R1702 vdd.n3181 vdd.n3180 185
R1703 vdd.n3180 vdd.n774 185
R1704 vdd.n3179 vdd.n807 185
R1705 vdd.n3179 vdd.n3178 185
R1706 vdd.n2822 vdd.n808 185
R1707 vdd.n817 vdd.n808 185
R1708 vdd.n2823 vdd.n815 185
R1709 vdd.n3172 vdd.n815 185
R1710 vdd.n2825 vdd.n2824 185
R1711 vdd.n2824 vdd.n814 185
R1712 vdd.n2826 vdd.n823 185
R1713 vdd.n3121 vdd.n823 185
R1714 vdd.n2828 vdd.n2827 185
R1715 vdd.n2827 vdd.n822 185
R1716 vdd.n2829 vdd.n828 185
R1717 vdd.n3115 vdd.n828 185
R1718 vdd.n2831 vdd.n2830 185
R1719 vdd.n2830 vdd.n835 185
R1720 vdd.n2832 vdd.n833 185
R1721 vdd.n3109 vdd.n833 185
R1722 vdd.n2834 vdd.n2833 185
R1723 vdd.n2833 vdd.n841 185
R1724 vdd.n2835 vdd.n839 185
R1725 vdd.n3103 vdd.n839 185
R1726 vdd.n2837 vdd.n2836 185
R1727 vdd.n2836 vdd.n848 185
R1728 vdd.n2838 vdd.n846 185
R1729 vdd.n3097 vdd.n846 185
R1730 vdd.n2840 vdd.n2839 185
R1731 vdd.n2839 vdd.n845 185
R1732 vdd.n2841 vdd.n853 185
R1733 vdd.n3091 vdd.n853 185
R1734 vdd.n2843 vdd.n2842 185
R1735 vdd.n2842 vdd.n852 185
R1736 vdd.n2844 vdd.n859 185
R1737 vdd.n3085 vdd.n859 185
R1738 vdd.n2846 vdd.n2845 185
R1739 vdd.n2845 vdd.n858 185
R1740 vdd.n2847 vdd.n864 185
R1741 vdd.n3079 vdd.n864 185
R1742 vdd.n2849 vdd.n2848 185
R1743 vdd.n2848 vdd.n872 185
R1744 vdd.n2850 vdd.n870 185
R1745 vdd.n3073 vdd.n870 185
R1746 vdd.n2852 vdd.n2851 185
R1747 vdd.n2851 vdd.n879 185
R1748 vdd.n2853 vdd.n877 185
R1749 vdd.n3067 vdd.n877 185
R1750 vdd.n2855 vdd.n2854 185
R1751 vdd.n2854 vdd.n876 185
R1752 vdd.n2856 vdd.n884 185
R1753 vdd.n3060 vdd.n884 185
R1754 vdd.n2858 vdd.n2857 185
R1755 vdd.n2857 vdd.n883 185
R1756 vdd.n2859 vdd.n889 185
R1757 vdd.n3054 vdd.n889 185
R1758 vdd.n2861 vdd.n2860 185
R1759 vdd.n2860 vdd.n896 185
R1760 vdd.n2862 vdd.n894 185
R1761 vdd.n3048 vdd.n894 185
R1762 vdd.n2864 vdd.n2863 185
R1763 vdd.n2863 vdd.n902 185
R1764 vdd.n2865 vdd.n900 185
R1765 vdd.n3042 vdd.n900 185
R1766 vdd.n2917 vdd.n2916 185
R1767 vdd.n2916 vdd.n2915 185
R1768 vdd.n2918 vdd.n906 185
R1769 vdd.n3036 vdd.n906 185
R1770 vdd.n2920 vdd.n2919 185
R1771 vdd.n2921 vdd.n2920 185
R1772 vdd.n2821 vdd.n912 185
R1773 vdd.n3030 vdd.n912 185
R1774 vdd.n2820 vdd.n2819 185
R1775 vdd.n2819 vdd.n911 185
R1776 vdd.n2818 vdd.n918 185
R1777 vdd.n3024 vdd.n918 185
R1778 vdd.n2817 vdd.n2816 185
R1779 vdd.n2816 vdd.n917 185
R1780 vdd.n2739 vdd.n923 185
R1781 vdd.n3018 vdd.n923 185
R1782 vdd.n2935 vdd.n2934 185
R1783 vdd.n2934 vdd.n2933 185
R1784 vdd.n2936 vdd.n929 185
R1785 vdd.n3012 vdd.n929 185
R1786 vdd.n2938 vdd.n2937 185
R1787 vdd.n2938 vdd.n928 185
R1788 vdd.n3009 vdd.n931 185
R1789 vdd.n931 vdd.n928 185
R1790 vdd.n3011 vdd.n3010 185
R1791 vdd.n3012 vdd.n3011 185
R1792 vdd.n922 vdd.n921 185
R1793 vdd.n2933 vdd.n922 185
R1794 vdd.n3020 vdd.n3019 185
R1795 vdd.n3019 vdd.n3018 185
R1796 vdd.n3021 vdd.n920 185
R1797 vdd.n920 vdd.n917 185
R1798 vdd.n3023 vdd.n3022 185
R1799 vdd.n3024 vdd.n3023 185
R1800 vdd.n910 vdd.n909 185
R1801 vdd.n911 vdd.n910 185
R1802 vdd.n3032 vdd.n3031 185
R1803 vdd.n3031 vdd.n3030 185
R1804 vdd.n3033 vdd.n908 185
R1805 vdd.n2921 vdd.n908 185
R1806 vdd.n3035 vdd.n3034 185
R1807 vdd.n3036 vdd.n3035 185
R1808 vdd.n899 vdd.n898 185
R1809 vdd.n2915 vdd.n899 185
R1810 vdd.n3044 vdd.n3043 185
R1811 vdd.n3043 vdd.n3042 185
R1812 vdd.n3045 vdd.n897 185
R1813 vdd.n902 vdd.n897 185
R1814 vdd.n3047 vdd.n3046 185
R1815 vdd.n3048 vdd.n3047 185
R1816 vdd.n888 vdd.n887 185
R1817 vdd.n896 vdd.n888 185
R1818 vdd.n3056 vdd.n3055 185
R1819 vdd.n3055 vdd.n3054 185
R1820 vdd.n3057 vdd.n886 185
R1821 vdd.n886 vdd.n883 185
R1822 vdd.n3059 vdd.n3058 185
R1823 vdd.n3060 vdd.n3059 185
R1824 vdd.n875 vdd.n874 185
R1825 vdd.n876 vdd.n875 185
R1826 vdd.n3069 vdd.n3068 185
R1827 vdd.n3068 vdd.n3067 185
R1828 vdd.n3070 vdd.n873 185
R1829 vdd.n879 vdd.n873 185
R1830 vdd.n3072 vdd.n3071 185
R1831 vdd.n3073 vdd.n3072 185
R1832 vdd.n863 vdd.n862 185
R1833 vdd.n872 vdd.n863 185
R1834 vdd.n3081 vdd.n3080 185
R1835 vdd.n3080 vdd.n3079 185
R1836 vdd.n3082 vdd.n861 185
R1837 vdd.n861 vdd.n858 185
R1838 vdd.n3084 vdd.n3083 185
R1839 vdd.n3085 vdd.n3084 185
R1840 vdd.n851 vdd.n850 185
R1841 vdd.n852 vdd.n851 185
R1842 vdd.n3093 vdd.n3092 185
R1843 vdd.n3092 vdd.n3091 185
R1844 vdd.n3094 vdd.n849 185
R1845 vdd.n849 vdd.n845 185
R1846 vdd.n3096 vdd.n3095 185
R1847 vdd.n3097 vdd.n3096 185
R1848 vdd.n838 vdd.n837 185
R1849 vdd.n848 vdd.n838 185
R1850 vdd.n3105 vdd.n3104 185
R1851 vdd.n3104 vdd.n3103 185
R1852 vdd.n3106 vdd.n836 185
R1853 vdd.n841 vdd.n836 185
R1854 vdd.n3108 vdd.n3107 185
R1855 vdd.n3109 vdd.n3108 185
R1856 vdd.n827 vdd.n826 185
R1857 vdd.n835 vdd.n827 185
R1858 vdd.n3117 vdd.n3116 185
R1859 vdd.n3116 vdd.n3115 185
R1860 vdd.n3118 vdd.n825 185
R1861 vdd.n825 vdd.n822 185
R1862 vdd.n3120 vdd.n3119 185
R1863 vdd.n3121 vdd.n3120 185
R1864 vdd.n813 vdd.n812 185
R1865 vdd.n814 vdd.n813 185
R1866 vdd.n3174 vdd.n3173 185
R1867 vdd.n3173 vdd.n3172 185
R1868 vdd.n3175 vdd.n811 185
R1869 vdd.n817 vdd.n811 185
R1870 vdd.n3177 vdd.n3176 185
R1871 vdd.n3178 vdd.n3177 185
R1872 vdd.n779 vdd.n777 185
R1873 vdd.n777 vdd.n774 185
R1874 vdd.n3247 vdd.n3246 185
R1875 vdd.n3248 vdd.n3247 185
R1876 vdd.n2628 vdd.n2627 185
R1877 vdd.n2629 vdd.n2628 185
R1878 vdd.n980 vdd.n978 185
R1879 vdd.n978 vdd.n976 185
R1880 vdd.n2543 vdd.n987 185
R1881 vdd.n2554 vdd.n987 185
R1882 vdd.n2544 vdd.n996 185
R1883 vdd.n1370 vdd.n996 185
R1884 vdd.n2546 vdd.n2545 185
R1885 vdd.n2547 vdd.n2546 185
R1886 vdd.n2542 vdd.n995 185
R1887 vdd.n995 vdd.n992 185
R1888 vdd.n2541 vdd.n2540 185
R1889 vdd.n2540 vdd.n2539 185
R1890 vdd.n998 vdd.n997 185
R1891 vdd.n999 vdd.n998 185
R1892 vdd.n2532 vdd.n2531 185
R1893 vdd.n2533 vdd.n2532 185
R1894 vdd.n2530 vdd.n1007 185
R1895 vdd.n1396 vdd.n1007 185
R1896 vdd.n2529 vdd.n2528 185
R1897 vdd.n2528 vdd.n2527 185
R1898 vdd.n1009 vdd.n1008 185
R1899 vdd.n1017 vdd.n1009 185
R1900 vdd.n2520 vdd.n2519 185
R1901 vdd.n2521 vdd.n2520 185
R1902 vdd.n2518 vdd.n1018 185
R1903 vdd.n1023 vdd.n1018 185
R1904 vdd.n2517 vdd.n2516 185
R1905 vdd.n2516 vdd.n2515 185
R1906 vdd.n1020 vdd.n1019 185
R1907 vdd.n1408 vdd.n1020 185
R1908 vdd.n2508 vdd.n2507 185
R1909 vdd.n2509 vdd.n2508 185
R1910 vdd.n2506 vdd.n1030 185
R1911 vdd.n1030 vdd.n1027 185
R1912 vdd.n2505 vdd.n2504 185
R1913 vdd.n2504 vdd.n2503 185
R1914 vdd.n1032 vdd.n1031 185
R1915 vdd.n1033 vdd.n1032 185
R1916 vdd.n2496 vdd.n2495 185
R1917 vdd.n2497 vdd.n2496 185
R1918 vdd.n2493 vdd.n1041 185
R1919 vdd.n1047 vdd.n1041 185
R1920 vdd.n2492 vdd.n2491 185
R1921 vdd.n2491 vdd.n2490 185
R1922 vdd.n1044 vdd.n1043 185
R1923 vdd.n1054 vdd.n1044 185
R1924 vdd.n2483 vdd.n2482 185
R1925 vdd.n2484 vdd.n2483 185
R1926 vdd.n2481 vdd.n1055 185
R1927 vdd.n1055 vdd.n1051 185
R1928 vdd.n2480 vdd.n2479 185
R1929 vdd.n2479 vdd.n2478 185
R1930 vdd.n1057 vdd.n1056 185
R1931 vdd.n1058 vdd.n1057 185
R1932 vdd.n2471 vdd.n2470 185
R1933 vdd.n2472 vdd.n2471 185
R1934 vdd.n2469 vdd.n1067 185
R1935 vdd.n1067 vdd.n1064 185
R1936 vdd.n2468 vdd.n2467 185
R1937 vdd.n2467 vdd.n2466 185
R1938 vdd.n1069 vdd.n1068 185
R1939 vdd.n1077 vdd.n1069 185
R1940 vdd.n2459 vdd.n2458 185
R1941 vdd.n2460 vdd.n2459 185
R1942 vdd.n2457 vdd.n1078 185
R1943 vdd.n1083 vdd.n1078 185
R1944 vdd.n2456 vdd.n2455 185
R1945 vdd.n2455 vdd.n2454 185
R1946 vdd.n1080 vdd.n1079 185
R1947 vdd.n1090 vdd.n1080 185
R1948 vdd.n2447 vdd.n2446 185
R1949 vdd.n2448 vdd.n2447 185
R1950 vdd.n2445 vdd.n1091 185
R1951 vdd.n1091 vdd.n1087 185
R1952 vdd.n2444 vdd.n2443 185
R1953 vdd.n2443 vdd.n2442 185
R1954 vdd.n1093 vdd.n1092 185
R1955 vdd.n1094 vdd.n1093 185
R1956 vdd.n2435 vdd.n2434 185
R1957 vdd.n2436 vdd.n2435 185
R1958 vdd.n2433 vdd.n1102 185
R1959 vdd.n1108 vdd.n1102 185
R1960 vdd.n2432 vdd.n2431 185
R1961 vdd.n2431 vdd.n2430 185
R1962 vdd.n1104 vdd.n1103 185
R1963 vdd.n1105 vdd.n1104 185
R1964 vdd.n2559 vdd.n951 185
R1965 vdd.n2701 vdd.n951 185
R1966 vdd.n2561 vdd.n2560 185
R1967 vdd.n2563 vdd.n2562 185
R1968 vdd.n2565 vdd.n2564 185
R1969 vdd.n2567 vdd.n2566 185
R1970 vdd.n2569 vdd.n2568 185
R1971 vdd.n2571 vdd.n2570 185
R1972 vdd.n2573 vdd.n2572 185
R1973 vdd.n2575 vdd.n2574 185
R1974 vdd.n2577 vdd.n2576 185
R1975 vdd.n2579 vdd.n2578 185
R1976 vdd.n2581 vdd.n2580 185
R1977 vdd.n2583 vdd.n2582 185
R1978 vdd.n2585 vdd.n2584 185
R1979 vdd.n2587 vdd.n2586 185
R1980 vdd.n2589 vdd.n2588 185
R1981 vdd.n2591 vdd.n2590 185
R1982 vdd.n2593 vdd.n2592 185
R1983 vdd.n2595 vdd.n2594 185
R1984 vdd.n2597 vdd.n2596 185
R1985 vdd.n2599 vdd.n2598 185
R1986 vdd.n2601 vdd.n2600 185
R1987 vdd.n2603 vdd.n2602 185
R1988 vdd.n2605 vdd.n2604 185
R1989 vdd.n2607 vdd.n2606 185
R1990 vdd.n2609 vdd.n2608 185
R1991 vdd.n2611 vdd.n2610 185
R1992 vdd.n2613 vdd.n2612 185
R1993 vdd.n2615 vdd.n2614 185
R1994 vdd.n2617 vdd.n2616 185
R1995 vdd.n2619 vdd.n2618 185
R1996 vdd.n2621 vdd.n2620 185
R1997 vdd.n2623 vdd.n2622 185
R1998 vdd.n2625 vdd.n2624 185
R1999 vdd.n2626 vdd.n979 185
R2000 vdd.n2558 vdd.n977 185
R2001 vdd.n2629 vdd.n977 185
R2002 vdd.n2557 vdd.n2556 185
R2003 vdd.n2556 vdd.n976 185
R2004 vdd.n2555 vdd.n984 185
R2005 vdd.n2555 vdd.n2554 185
R2006 vdd.n1386 vdd.n985 185
R2007 vdd.n1370 vdd.n985 185
R2008 vdd.n1387 vdd.n994 185
R2009 vdd.n2547 vdd.n994 185
R2010 vdd.n1389 vdd.n1388 185
R2011 vdd.n1388 vdd.n992 185
R2012 vdd.n1390 vdd.n1001 185
R2013 vdd.n2539 vdd.n1001 185
R2014 vdd.n1392 vdd.n1391 185
R2015 vdd.n1391 vdd.n999 185
R2016 vdd.n1393 vdd.n1006 185
R2017 vdd.n2533 vdd.n1006 185
R2018 vdd.n1395 vdd.n1394 185
R2019 vdd.n1396 vdd.n1395 185
R2020 vdd.n1385 vdd.n1011 185
R2021 vdd.n2527 vdd.n1011 185
R2022 vdd.n1384 vdd.n1383 185
R2023 vdd.n1383 vdd.n1017 185
R2024 vdd.n1382 vdd.n1016 185
R2025 vdd.n2521 vdd.n1016 185
R2026 vdd.n1381 vdd.n1380 185
R2027 vdd.n1380 vdd.n1023 185
R2028 vdd.n1289 vdd.n1022 185
R2029 vdd.n2515 vdd.n1022 185
R2030 vdd.n1410 vdd.n1409 185
R2031 vdd.n1409 vdd.n1408 185
R2032 vdd.n1411 vdd.n1029 185
R2033 vdd.n2509 vdd.n1029 185
R2034 vdd.n1413 vdd.n1412 185
R2035 vdd.n1412 vdd.n1027 185
R2036 vdd.n1414 vdd.n1035 185
R2037 vdd.n2503 vdd.n1035 185
R2038 vdd.n1416 vdd.n1415 185
R2039 vdd.n1415 vdd.n1033 185
R2040 vdd.n1417 vdd.n1040 185
R2041 vdd.n2497 vdd.n1040 185
R2042 vdd.n1419 vdd.n1418 185
R2043 vdd.n1418 vdd.n1047 185
R2044 vdd.n1420 vdd.n1046 185
R2045 vdd.n2490 vdd.n1046 185
R2046 vdd.n1422 vdd.n1421 185
R2047 vdd.n1421 vdd.n1054 185
R2048 vdd.n1423 vdd.n1053 185
R2049 vdd.n2484 vdd.n1053 185
R2050 vdd.n1425 vdd.n1424 185
R2051 vdd.n1424 vdd.n1051 185
R2052 vdd.n1426 vdd.n1060 185
R2053 vdd.n2478 vdd.n1060 185
R2054 vdd.n1428 vdd.n1427 185
R2055 vdd.n1427 vdd.n1058 185
R2056 vdd.n1429 vdd.n1066 185
R2057 vdd.n2472 vdd.n1066 185
R2058 vdd.n1431 vdd.n1430 185
R2059 vdd.n1430 vdd.n1064 185
R2060 vdd.n1432 vdd.n1071 185
R2061 vdd.n2466 vdd.n1071 185
R2062 vdd.n1434 vdd.n1433 185
R2063 vdd.n1433 vdd.n1077 185
R2064 vdd.n1435 vdd.n1076 185
R2065 vdd.n2460 vdd.n1076 185
R2066 vdd.n1437 vdd.n1436 185
R2067 vdd.n1436 vdd.n1083 185
R2068 vdd.n1438 vdd.n1082 185
R2069 vdd.n2454 vdd.n1082 185
R2070 vdd.n1440 vdd.n1439 185
R2071 vdd.n1439 vdd.n1090 185
R2072 vdd.n1441 vdd.n1089 185
R2073 vdd.n2448 vdd.n1089 185
R2074 vdd.n1443 vdd.n1442 185
R2075 vdd.n1442 vdd.n1087 185
R2076 vdd.n1444 vdd.n1096 185
R2077 vdd.n2442 vdd.n1096 185
R2078 vdd.n1446 vdd.n1445 185
R2079 vdd.n1445 vdd.n1094 185
R2080 vdd.n1447 vdd.n1101 185
R2081 vdd.n2436 vdd.n1101 185
R2082 vdd.n1449 vdd.n1448 185
R2083 vdd.n1448 vdd.n1108 185
R2084 vdd.n1450 vdd.n1107 185
R2085 vdd.n2430 vdd.n1107 185
R2086 vdd.n1452 vdd.n1451 185
R2087 vdd.n1451 vdd.n1105 185
R2088 vdd.n1252 vdd.n1251 185
R2089 vdd.n1254 vdd.n1253 185
R2090 vdd.n1256 vdd.n1255 185
R2091 vdd.n1258 vdd.n1257 185
R2092 vdd.n1260 vdd.n1259 185
R2093 vdd.n1262 vdd.n1261 185
R2094 vdd.n1264 vdd.n1263 185
R2095 vdd.n1266 vdd.n1265 185
R2096 vdd.n1268 vdd.n1267 185
R2097 vdd.n1270 vdd.n1269 185
R2098 vdd.n1272 vdd.n1271 185
R2099 vdd.n1274 vdd.n1273 185
R2100 vdd.n1276 vdd.n1275 185
R2101 vdd.n1278 vdd.n1277 185
R2102 vdd.n1280 vdd.n1279 185
R2103 vdd.n1282 vdd.n1281 185
R2104 vdd.n1284 vdd.n1283 185
R2105 vdd.n1486 vdd.n1285 185
R2106 vdd.n1485 vdd.n1484 185
R2107 vdd.n1483 vdd.n1482 185
R2108 vdd.n1481 vdd.n1480 185
R2109 vdd.n1479 vdd.n1478 185
R2110 vdd.n1477 vdd.n1476 185
R2111 vdd.n1475 vdd.n1474 185
R2112 vdd.n1473 vdd.n1472 185
R2113 vdd.n1471 vdd.n1470 185
R2114 vdd.n1469 vdd.n1468 185
R2115 vdd.n1467 vdd.n1466 185
R2116 vdd.n1465 vdd.n1464 185
R2117 vdd.n1463 vdd.n1462 185
R2118 vdd.n1461 vdd.n1460 185
R2119 vdd.n1459 vdd.n1458 185
R2120 vdd.n1457 vdd.n1456 185
R2121 vdd.n1455 vdd.n1454 185
R2122 vdd.n1453 vdd.n1146 185
R2123 vdd.n2423 vdd.n1146 185
R2124 vdd.n315 vdd.n314 171.744
R2125 vdd.n314 vdd.n313 171.744
R2126 vdd.n313 vdd.n282 171.744
R2127 vdd.n306 vdd.n282 171.744
R2128 vdd.n306 vdd.n305 171.744
R2129 vdd.n305 vdd.n287 171.744
R2130 vdd.n298 vdd.n287 171.744
R2131 vdd.n298 vdd.n297 171.744
R2132 vdd.n297 vdd.n291 171.744
R2133 vdd.n260 vdd.n259 171.744
R2134 vdd.n259 vdd.n258 171.744
R2135 vdd.n258 vdd.n227 171.744
R2136 vdd.n251 vdd.n227 171.744
R2137 vdd.n251 vdd.n250 171.744
R2138 vdd.n250 vdd.n232 171.744
R2139 vdd.n243 vdd.n232 171.744
R2140 vdd.n243 vdd.n242 171.744
R2141 vdd.n242 vdd.n236 171.744
R2142 vdd.n217 vdd.n216 171.744
R2143 vdd.n216 vdd.n215 171.744
R2144 vdd.n215 vdd.n184 171.744
R2145 vdd.n208 vdd.n184 171.744
R2146 vdd.n208 vdd.n207 171.744
R2147 vdd.n207 vdd.n189 171.744
R2148 vdd.n200 vdd.n189 171.744
R2149 vdd.n200 vdd.n199 171.744
R2150 vdd.n199 vdd.n193 171.744
R2151 vdd.n162 vdd.n161 171.744
R2152 vdd.n161 vdd.n160 171.744
R2153 vdd.n160 vdd.n129 171.744
R2154 vdd.n153 vdd.n129 171.744
R2155 vdd.n153 vdd.n152 171.744
R2156 vdd.n152 vdd.n134 171.744
R2157 vdd.n145 vdd.n134 171.744
R2158 vdd.n145 vdd.n144 171.744
R2159 vdd.n144 vdd.n138 171.744
R2160 vdd.n120 vdd.n119 171.744
R2161 vdd.n119 vdd.n118 171.744
R2162 vdd.n118 vdd.n87 171.744
R2163 vdd.n111 vdd.n87 171.744
R2164 vdd.n111 vdd.n110 171.744
R2165 vdd.n110 vdd.n92 171.744
R2166 vdd.n103 vdd.n92 171.744
R2167 vdd.n103 vdd.n102 171.744
R2168 vdd.n102 vdd.n96 171.744
R2169 vdd.n65 vdd.n64 171.744
R2170 vdd.n64 vdd.n63 171.744
R2171 vdd.n63 vdd.n32 171.744
R2172 vdd.n56 vdd.n32 171.744
R2173 vdd.n56 vdd.n55 171.744
R2174 vdd.n55 vdd.n37 171.744
R2175 vdd.n48 vdd.n37 171.744
R2176 vdd.n48 vdd.n47 171.744
R2177 vdd.n47 vdd.n41 171.744
R2178 vdd.n2139 vdd.n2138 171.744
R2179 vdd.n2138 vdd.n2137 171.744
R2180 vdd.n2137 vdd.n2106 171.744
R2181 vdd.n2130 vdd.n2106 171.744
R2182 vdd.n2130 vdd.n2129 171.744
R2183 vdd.n2129 vdd.n2111 171.744
R2184 vdd.n2122 vdd.n2111 171.744
R2185 vdd.n2122 vdd.n2121 171.744
R2186 vdd.n2121 vdd.n2115 171.744
R2187 vdd.n2194 vdd.n2193 171.744
R2188 vdd.n2193 vdd.n2192 171.744
R2189 vdd.n2192 vdd.n2161 171.744
R2190 vdd.n2185 vdd.n2161 171.744
R2191 vdd.n2185 vdd.n2184 171.744
R2192 vdd.n2184 vdd.n2166 171.744
R2193 vdd.n2177 vdd.n2166 171.744
R2194 vdd.n2177 vdd.n2176 171.744
R2195 vdd.n2176 vdd.n2170 171.744
R2196 vdd.n2041 vdd.n2040 171.744
R2197 vdd.n2040 vdd.n2039 171.744
R2198 vdd.n2039 vdd.n2008 171.744
R2199 vdd.n2032 vdd.n2008 171.744
R2200 vdd.n2032 vdd.n2031 171.744
R2201 vdd.n2031 vdd.n2013 171.744
R2202 vdd.n2024 vdd.n2013 171.744
R2203 vdd.n2024 vdd.n2023 171.744
R2204 vdd.n2023 vdd.n2017 171.744
R2205 vdd.n2096 vdd.n2095 171.744
R2206 vdd.n2095 vdd.n2094 171.744
R2207 vdd.n2094 vdd.n2063 171.744
R2208 vdd.n2087 vdd.n2063 171.744
R2209 vdd.n2087 vdd.n2086 171.744
R2210 vdd.n2086 vdd.n2068 171.744
R2211 vdd.n2079 vdd.n2068 171.744
R2212 vdd.n2079 vdd.n2078 171.744
R2213 vdd.n2078 vdd.n2072 171.744
R2214 vdd.n1944 vdd.n1943 171.744
R2215 vdd.n1943 vdd.n1942 171.744
R2216 vdd.n1942 vdd.n1911 171.744
R2217 vdd.n1935 vdd.n1911 171.744
R2218 vdd.n1935 vdd.n1934 171.744
R2219 vdd.n1934 vdd.n1916 171.744
R2220 vdd.n1927 vdd.n1916 171.744
R2221 vdd.n1927 vdd.n1926 171.744
R2222 vdd.n1926 vdd.n1920 171.744
R2223 vdd.n1999 vdd.n1998 171.744
R2224 vdd.n1998 vdd.n1997 171.744
R2225 vdd.n1997 vdd.n1966 171.744
R2226 vdd.n1990 vdd.n1966 171.744
R2227 vdd.n1990 vdd.n1989 171.744
R2228 vdd.n1989 vdd.n1971 171.744
R2229 vdd.n1982 vdd.n1971 171.744
R2230 vdd.n1982 vdd.n1981 171.744
R2231 vdd.n1981 vdd.n1975 171.744
R2232 vdd.n449 vdd.n448 146.341
R2233 vdd.n455 vdd.n454 146.341
R2234 vdd.n459 vdd.n458 146.341
R2235 vdd.n465 vdd.n464 146.341
R2236 vdd.n469 vdd.n468 146.341
R2237 vdd.n475 vdd.n474 146.341
R2238 vdd.n479 vdd.n478 146.341
R2239 vdd.n485 vdd.n484 146.341
R2240 vdd.n489 vdd.n488 146.341
R2241 vdd.n495 vdd.n494 146.341
R2242 vdd.n499 vdd.n498 146.341
R2243 vdd.n505 vdd.n504 146.341
R2244 vdd.n509 vdd.n508 146.341
R2245 vdd.n515 vdd.n514 146.341
R2246 vdd.n519 vdd.n518 146.341
R2247 vdd.n525 vdd.n524 146.341
R2248 vdd.n529 vdd.n528 146.341
R2249 vdd.n535 vdd.n534 146.341
R2250 vdd.n539 vdd.n538 146.341
R2251 vdd.n545 vdd.n544 146.341
R2252 vdd.n549 vdd.n548 146.341
R2253 vdd.n555 vdd.n554 146.341
R2254 vdd.n559 vdd.n558 146.341
R2255 vdd.n565 vdd.n564 146.341
R2256 vdd.n569 vdd.n568 146.341
R2257 vdd.n575 vdd.n574 146.341
R2258 vdd.n579 vdd.n578 146.341
R2259 vdd.n585 vdd.n584 146.341
R2260 vdd.n589 vdd.n588 146.341
R2261 vdd.n595 vdd.n594 146.341
R2262 vdd.n597 vdd.n404 146.341
R2263 vdd.n3418 vdd.n654 146.341
R2264 vdd.n3424 vdd.n654 146.341
R2265 vdd.n3424 vdd.n647 146.341
R2266 vdd.n3434 vdd.n647 146.341
R2267 vdd.n3434 vdd.n643 146.341
R2268 vdd.n3440 vdd.n643 146.341
R2269 vdd.n3440 vdd.n634 146.341
R2270 vdd.n3450 vdd.n634 146.341
R2271 vdd.n3450 vdd.n630 146.341
R2272 vdd.n3456 vdd.n630 146.341
R2273 vdd.n3456 vdd.n623 146.341
R2274 vdd.n3467 vdd.n623 146.341
R2275 vdd.n3467 vdd.n619 146.341
R2276 vdd.n3476 vdd.n619 146.341
R2277 vdd.n3476 vdd.n612 146.341
R2278 vdd.n3486 vdd.n612 146.341
R2279 vdd.n3487 vdd.n3486 146.341
R2280 vdd.n3487 vdd.n329 146.341
R2281 vdd.n330 vdd.n329 146.341
R2282 vdd.n331 vdd.n330 146.341
R2283 vdd.n3494 vdd.n331 146.341
R2284 vdd.n3494 vdd.n339 146.341
R2285 vdd.n340 vdd.n339 146.341
R2286 vdd.n341 vdd.n340 146.341
R2287 vdd.n3501 vdd.n341 146.341
R2288 vdd.n3501 vdd.n350 146.341
R2289 vdd.n351 vdd.n350 146.341
R2290 vdd.n352 vdd.n351 146.341
R2291 vdd.n3509 vdd.n352 146.341
R2292 vdd.n3509 vdd.n360 146.341
R2293 vdd.n361 vdd.n360 146.341
R2294 vdd.n362 vdd.n361 146.341
R2295 vdd.n3516 vdd.n362 146.341
R2296 vdd.n3516 vdd.n371 146.341
R2297 vdd.n372 vdd.n371 146.341
R2298 vdd.n3410 vdd.n3408 146.341
R2299 vdd.n3408 vdd.n3407 146.341
R2300 vdd.n3404 vdd.n3403 146.341
R2301 vdd.n3400 vdd.n3399 146.341
R2302 vdd.n3397 vdd.n669 146.341
R2303 vdd.n3393 vdd.n3391 146.341
R2304 vdd.n3389 vdd.n675 146.341
R2305 vdd.n3385 vdd.n3383 146.341
R2306 vdd.n3381 vdd.n681 146.341
R2307 vdd.n3377 vdd.n3375 146.341
R2308 vdd.n3373 vdd.n689 146.341
R2309 vdd.n3369 vdd.n3367 146.341
R2310 vdd.n3365 vdd.n695 146.341
R2311 vdd.n3361 vdd.n3359 146.341
R2312 vdd.n3357 vdd.n701 146.341
R2313 vdd.n3353 vdd.n3351 146.341
R2314 vdd.n3349 vdd.n707 146.341
R2315 vdd.n3345 vdd.n3343 146.341
R2316 vdd.n3341 vdd.n713 146.341
R2317 vdd.n3337 vdd.n3335 146.341
R2318 vdd.n3333 vdd.n719 146.341
R2319 vdd.n3326 vdd.n728 146.341
R2320 vdd.n3324 vdd.n3323 146.341
R2321 vdd.n3320 vdd.n3319 146.341
R2322 vdd.n3317 vdd.n733 146.341
R2323 vdd.n3313 vdd.n3311 146.341
R2324 vdd.n3309 vdd.n739 146.341
R2325 vdd.n3305 vdd.n3303 146.341
R2326 vdd.n3301 vdd.n745 146.341
R2327 vdd.n3297 vdd.n3295 146.341
R2328 vdd.n3292 vdd.n3291 146.341
R2329 vdd.n3288 vdd.n657 146.341
R2330 vdd.n3416 vdd.n653 146.341
R2331 vdd.n3426 vdd.n653 146.341
R2332 vdd.n3426 vdd.n649 146.341
R2333 vdd.n3432 vdd.n649 146.341
R2334 vdd.n3432 vdd.n641 146.341
R2335 vdd.n3442 vdd.n641 146.341
R2336 vdd.n3442 vdd.n637 146.341
R2337 vdd.n3448 vdd.n637 146.341
R2338 vdd.n3448 vdd.n629 146.341
R2339 vdd.n3459 vdd.n629 146.341
R2340 vdd.n3459 vdd.n625 146.341
R2341 vdd.n3465 vdd.n625 146.341
R2342 vdd.n3465 vdd.n618 146.341
R2343 vdd.n3478 vdd.n618 146.341
R2344 vdd.n3478 vdd.n614 146.341
R2345 vdd.n3484 vdd.n614 146.341
R2346 vdd.n3484 vdd.n326 146.341
R2347 vdd.n3560 vdd.n326 146.341
R2348 vdd.n3560 vdd.n327 146.341
R2349 vdd.n3556 vdd.n327 146.341
R2350 vdd.n3556 vdd.n333 146.341
R2351 vdd.n3552 vdd.n333 146.341
R2352 vdd.n3552 vdd.n338 146.341
R2353 vdd.n3548 vdd.n338 146.341
R2354 vdd.n3548 vdd.n342 146.341
R2355 vdd.n3544 vdd.n342 146.341
R2356 vdd.n3544 vdd.n348 146.341
R2357 vdd.n3540 vdd.n348 146.341
R2358 vdd.n3540 vdd.n353 146.341
R2359 vdd.n3536 vdd.n353 146.341
R2360 vdd.n3536 vdd.n359 146.341
R2361 vdd.n3532 vdd.n359 146.341
R2362 vdd.n3532 vdd.n364 146.341
R2363 vdd.n3528 vdd.n364 146.341
R2364 vdd.n3528 vdd.n370 146.341
R2365 vdd.n2388 vdd.n2387 146.341
R2366 vdd.n2385 vdd.n2382 146.341
R2367 vdd.n2380 vdd.n1156 146.341
R2368 vdd.n2376 vdd.n2375 146.341
R2369 vdd.n2373 vdd.n1160 146.341
R2370 vdd.n2369 vdd.n2368 146.341
R2371 vdd.n2366 vdd.n1167 146.341
R2372 vdd.n2362 vdd.n2361 146.341
R2373 vdd.n2359 vdd.n1174 146.341
R2374 vdd.n1185 vdd.n1182 146.341
R2375 vdd.n2351 vdd.n2350 146.341
R2376 vdd.n2348 vdd.n1187 146.341
R2377 vdd.n2344 vdd.n2343 146.341
R2378 vdd.n2341 vdd.n1193 146.341
R2379 vdd.n2337 vdd.n2336 146.341
R2380 vdd.n2334 vdd.n1200 146.341
R2381 vdd.n2330 vdd.n2329 146.341
R2382 vdd.n2327 vdd.n1207 146.341
R2383 vdd.n2323 vdd.n2322 146.341
R2384 vdd.n2320 vdd.n1214 146.341
R2385 vdd.n1225 vdd.n1222 146.341
R2386 vdd.n2312 vdd.n2311 146.341
R2387 vdd.n2309 vdd.n1227 146.341
R2388 vdd.n2305 vdd.n2304 146.341
R2389 vdd.n2302 vdd.n1233 146.341
R2390 vdd.n2298 vdd.n2297 146.341
R2391 vdd.n2295 vdd.n1240 146.341
R2392 vdd.n2291 vdd.n2290 146.341
R2393 vdd.n2288 vdd.n1247 146.341
R2394 vdd.n1493 vdd.n1491 146.341
R2395 vdd.n1496 vdd.n1495 146.341
R2396 vdd.n1836 vdd.n1600 146.341
R2397 vdd.n1836 vdd.n1592 146.341
R2398 vdd.n1846 vdd.n1592 146.341
R2399 vdd.n1846 vdd.n1588 146.341
R2400 vdd.n1852 vdd.n1588 146.341
R2401 vdd.n1852 vdd.n1580 146.341
R2402 vdd.n1863 vdd.n1580 146.341
R2403 vdd.n1863 vdd.n1576 146.341
R2404 vdd.n1869 vdd.n1576 146.341
R2405 vdd.n1869 vdd.n1570 146.341
R2406 vdd.n1880 vdd.n1570 146.341
R2407 vdd.n1880 vdd.n1566 146.341
R2408 vdd.n1886 vdd.n1566 146.341
R2409 vdd.n1886 vdd.n1557 146.341
R2410 vdd.n1896 vdd.n1557 146.341
R2411 vdd.n1896 vdd.n1553 146.341
R2412 vdd.n1902 vdd.n1553 146.341
R2413 vdd.n1902 vdd.n1546 146.341
R2414 vdd.n2208 vdd.n1546 146.341
R2415 vdd.n2208 vdd.n1542 146.341
R2416 vdd.n2214 vdd.n1542 146.341
R2417 vdd.n2214 vdd.n1535 146.341
R2418 vdd.n2224 vdd.n1535 146.341
R2419 vdd.n2224 vdd.n1531 146.341
R2420 vdd.n2230 vdd.n1531 146.341
R2421 vdd.n2230 vdd.n1523 146.341
R2422 vdd.n2241 vdd.n1523 146.341
R2423 vdd.n2241 vdd.n1519 146.341
R2424 vdd.n2247 vdd.n1519 146.341
R2425 vdd.n2247 vdd.n1513 146.341
R2426 vdd.n2258 vdd.n1513 146.341
R2427 vdd.n2258 vdd.n1508 146.341
R2428 vdd.n2266 vdd.n1508 146.341
R2429 vdd.n2266 vdd.n1498 146.341
R2430 vdd.n2276 vdd.n1498 146.341
R2431 vdd.n1638 vdd.n1637 146.341
R2432 vdd.n1642 vdd.n1637 146.341
R2433 vdd.n1644 vdd.n1643 146.341
R2434 vdd.n1648 vdd.n1647 146.341
R2435 vdd.n1650 vdd.n1649 146.341
R2436 vdd.n1654 vdd.n1653 146.341
R2437 vdd.n1656 vdd.n1655 146.341
R2438 vdd.n1660 vdd.n1659 146.341
R2439 vdd.n1662 vdd.n1661 146.341
R2440 vdd.n1794 vdd.n1793 146.341
R2441 vdd.n1666 vdd.n1665 146.341
R2442 vdd.n1670 vdd.n1669 146.341
R2443 vdd.n1672 vdd.n1671 146.341
R2444 vdd.n1676 vdd.n1675 146.341
R2445 vdd.n1678 vdd.n1677 146.341
R2446 vdd.n1682 vdd.n1681 146.341
R2447 vdd.n1684 vdd.n1683 146.341
R2448 vdd.n1688 vdd.n1687 146.341
R2449 vdd.n1690 vdd.n1689 146.341
R2450 vdd.n1694 vdd.n1693 146.341
R2451 vdd.n1758 vdd.n1695 146.341
R2452 vdd.n1699 vdd.n1698 146.341
R2453 vdd.n1701 vdd.n1700 146.341
R2454 vdd.n1705 vdd.n1704 146.341
R2455 vdd.n1707 vdd.n1706 146.341
R2456 vdd.n1711 vdd.n1710 146.341
R2457 vdd.n1713 vdd.n1712 146.341
R2458 vdd.n1717 vdd.n1716 146.341
R2459 vdd.n1719 vdd.n1718 146.341
R2460 vdd.n1723 vdd.n1722 146.341
R2461 vdd.n1725 vdd.n1724 146.341
R2462 vdd.n1830 vdd.n1606 146.341
R2463 vdd.n1838 vdd.n1598 146.341
R2464 vdd.n1838 vdd.n1594 146.341
R2465 vdd.n1844 vdd.n1594 146.341
R2466 vdd.n1844 vdd.n1586 146.341
R2467 vdd.n1855 vdd.n1586 146.341
R2468 vdd.n1855 vdd.n1582 146.341
R2469 vdd.n1861 vdd.n1582 146.341
R2470 vdd.n1861 vdd.n1575 146.341
R2471 vdd.n1872 vdd.n1575 146.341
R2472 vdd.n1872 vdd.n1571 146.341
R2473 vdd.n1878 vdd.n1571 146.341
R2474 vdd.n1878 vdd.n1564 146.341
R2475 vdd.n1888 vdd.n1564 146.341
R2476 vdd.n1888 vdd.n1560 146.341
R2477 vdd.n1894 vdd.n1560 146.341
R2478 vdd.n1894 vdd.n1552 146.341
R2479 vdd.n1905 vdd.n1552 146.341
R2480 vdd.n1905 vdd.n1548 146.341
R2481 vdd.n2206 vdd.n1548 146.341
R2482 vdd.n2206 vdd.n1541 146.341
R2483 vdd.n2216 vdd.n1541 146.341
R2484 vdd.n2216 vdd.n1537 146.341
R2485 vdd.n2222 vdd.n1537 146.341
R2486 vdd.n2222 vdd.n1529 146.341
R2487 vdd.n2233 vdd.n1529 146.341
R2488 vdd.n2233 vdd.n1525 146.341
R2489 vdd.n2239 vdd.n1525 146.341
R2490 vdd.n2239 vdd.n1518 146.341
R2491 vdd.n2250 vdd.n1518 146.341
R2492 vdd.n2250 vdd.n1514 146.341
R2493 vdd.n2256 vdd.n1514 146.341
R2494 vdd.n2256 vdd.n1506 146.341
R2495 vdd.n2268 vdd.n1506 146.341
R2496 vdd.n2268 vdd.n1501 146.341
R2497 vdd.n2274 vdd.n1501 146.341
R2498 vdd.n1286 vdd.t72 127.284
R2499 vdd.n981 vdd.t116 127.284
R2500 vdd.n1290 vdd.t106 127.284
R2501 vdd.n972 vdd.t139 127.284
R2502 vdd.n867 vdd.t93 127.284
R2503 vdd.n867 vdd.t94 127.284
R2504 vdd.n2740 vdd.t134 127.284
R2505 vdd.n804 vdd.t81 127.284
R2506 vdd.n2737 vdd.t124 127.284
R2507 vdd.n768 vdd.t67 127.284
R2508 vdd.n1042 vdd.t130 127.284
R2509 vdd.n1042 vdd.t131 127.284
R2510 vdd.n22 vdd.n20 117.314
R2511 vdd.n17 vdd.n15 117.314
R2512 vdd.n27 vdd.n26 116.927
R2513 vdd.n24 vdd.n23 116.927
R2514 vdd.n22 vdd.n21 116.927
R2515 vdd.n17 vdd.n16 116.927
R2516 vdd.n19 vdd.n18 116.927
R2517 vdd.n27 vdd.n25 116.927
R2518 vdd.n1287 vdd.t71 111.188
R2519 vdd.n982 vdd.t117 111.188
R2520 vdd.n1291 vdd.t105 111.188
R2521 vdd.n973 vdd.t140 111.188
R2522 vdd.n2741 vdd.t133 111.188
R2523 vdd.n805 vdd.t82 111.188
R2524 vdd.n2738 vdd.t123 111.188
R2525 vdd.n769 vdd.t68 111.188
R2526 vdd.n3011 vdd.n931 99.5127
R2527 vdd.n3011 vdd.n922 99.5127
R2528 vdd.n3019 vdd.n922 99.5127
R2529 vdd.n3019 vdd.n920 99.5127
R2530 vdd.n3023 vdd.n920 99.5127
R2531 vdd.n3023 vdd.n910 99.5127
R2532 vdd.n3031 vdd.n910 99.5127
R2533 vdd.n3031 vdd.n908 99.5127
R2534 vdd.n3035 vdd.n908 99.5127
R2535 vdd.n3035 vdd.n899 99.5127
R2536 vdd.n3043 vdd.n899 99.5127
R2537 vdd.n3043 vdd.n897 99.5127
R2538 vdd.n3047 vdd.n897 99.5127
R2539 vdd.n3047 vdd.n888 99.5127
R2540 vdd.n3055 vdd.n888 99.5127
R2541 vdd.n3055 vdd.n886 99.5127
R2542 vdd.n3059 vdd.n886 99.5127
R2543 vdd.n3059 vdd.n875 99.5127
R2544 vdd.n3068 vdd.n875 99.5127
R2545 vdd.n3068 vdd.n873 99.5127
R2546 vdd.n3072 vdd.n873 99.5127
R2547 vdd.n3072 vdd.n863 99.5127
R2548 vdd.n3080 vdd.n863 99.5127
R2549 vdd.n3080 vdd.n861 99.5127
R2550 vdd.n3084 vdd.n861 99.5127
R2551 vdd.n3084 vdd.n851 99.5127
R2552 vdd.n3092 vdd.n851 99.5127
R2553 vdd.n3092 vdd.n849 99.5127
R2554 vdd.n3096 vdd.n849 99.5127
R2555 vdd.n3096 vdd.n838 99.5127
R2556 vdd.n3104 vdd.n838 99.5127
R2557 vdd.n3104 vdd.n836 99.5127
R2558 vdd.n3108 vdd.n836 99.5127
R2559 vdd.n3108 vdd.n827 99.5127
R2560 vdd.n3116 vdd.n827 99.5127
R2561 vdd.n3116 vdd.n825 99.5127
R2562 vdd.n3120 vdd.n825 99.5127
R2563 vdd.n3120 vdd.n813 99.5127
R2564 vdd.n3173 vdd.n813 99.5127
R2565 vdd.n3173 vdd.n811 99.5127
R2566 vdd.n3177 vdd.n811 99.5127
R2567 vdd.n3177 vdd.n777 99.5127
R2568 vdd.n3247 vdd.n777 99.5127
R2569 vdd.n3243 vdd.n778 99.5127
R2570 vdd.n3241 vdd.n3240 99.5127
R2571 vdd.n3238 vdd.n782 99.5127
R2572 vdd.n3234 vdd.n3233 99.5127
R2573 vdd.n3231 vdd.n785 99.5127
R2574 vdd.n3227 vdd.n3226 99.5127
R2575 vdd.n3224 vdd.n788 99.5127
R2576 vdd.n3220 vdd.n3219 99.5127
R2577 vdd.n3217 vdd.n791 99.5127
R2578 vdd.n3212 vdd.n3211 99.5127
R2579 vdd.n3209 vdd.n794 99.5127
R2580 vdd.n3205 vdd.n3204 99.5127
R2581 vdd.n3202 vdd.n797 99.5127
R2582 vdd.n3198 vdd.n3197 99.5127
R2583 vdd.n3195 vdd.n800 99.5127
R2584 vdd.n3191 vdd.n3190 99.5127
R2585 vdd.n3188 vdd.n803 99.5127
R2586 vdd.n2938 vdd.n929 99.5127
R2587 vdd.n2934 vdd.n929 99.5127
R2588 vdd.n2934 vdd.n923 99.5127
R2589 vdd.n2816 vdd.n923 99.5127
R2590 vdd.n2816 vdd.n918 99.5127
R2591 vdd.n2819 vdd.n918 99.5127
R2592 vdd.n2819 vdd.n912 99.5127
R2593 vdd.n2920 vdd.n912 99.5127
R2594 vdd.n2920 vdd.n906 99.5127
R2595 vdd.n2916 vdd.n906 99.5127
R2596 vdd.n2916 vdd.n900 99.5127
R2597 vdd.n2863 vdd.n900 99.5127
R2598 vdd.n2863 vdd.n894 99.5127
R2599 vdd.n2860 vdd.n894 99.5127
R2600 vdd.n2860 vdd.n889 99.5127
R2601 vdd.n2857 vdd.n889 99.5127
R2602 vdd.n2857 vdd.n884 99.5127
R2603 vdd.n2854 vdd.n884 99.5127
R2604 vdd.n2854 vdd.n877 99.5127
R2605 vdd.n2851 vdd.n877 99.5127
R2606 vdd.n2851 vdd.n870 99.5127
R2607 vdd.n2848 vdd.n870 99.5127
R2608 vdd.n2848 vdd.n864 99.5127
R2609 vdd.n2845 vdd.n864 99.5127
R2610 vdd.n2845 vdd.n859 99.5127
R2611 vdd.n2842 vdd.n859 99.5127
R2612 vdd.n2842 vdd.n853 99.5127
R2613 vdd.n2839 vdd.n853 99.5127
R2614 vdd.n2839 vdd.n846 99.5127
R2615 vdd.n2836 vdd.n846 99.5127
R2616 vdd.n2836 vdd.n839 99.5127
R2617 vdd.n2833 vdd.n839 99.5127
R2618 vdd.n2833 vdd.n833 99.5127
R2619 vdd.n2830 vdd.n833 99.5127
R2620 vdd.n2830 vdd.n828 99.5127
R2621 vdd.n2827 vdd.n828 99.5127
R2622 vdd.n2827 vdd.n823 99.5127
R2623 vdd.n2824 vdd.n823 99.5127
R2624 vdd.n2824 vdd.n815 99.5127
R2625 vdd.n815 vdd.n808 99.5127
R2626 vdd.n3179 vdd.n808 99.5127
R2627 vdd.n3180 vdd.n3179 99.5127
R2628 vdd.n3180 vdd.n775 99.5127
R2629 vdd.n3004 vdd.n933 99.5127
R2630 vdd.n3004 vdd.n2736 99.5127
R2631 vdd.n3000 vdd.n2999 99.5127
R2632 vdd.n2996 vdd.n2995 99.5127
R2633 vdd.n2992 vdd.n2991 99.5127
R2634 vdd.n2988 vdd.n2987 99.5127
R2635 vdd.n2984 vdd.n2983 99.5127
R2636 vdd.n2980 vdd.n2979 99.5127
R2637 vdd.n2976 vdd.n2975 99.5127
R2638 vdd.n2972 vdd.n2971 99.5127
R2639 vdd.n2968 vdd.n2967 99.5127
R2640 vdd.n2964 vdd.n2963 99.5127
R2641 vdd.n2960 vdd.n2959 99.5127
R2642 vdd.n2956 vdd.n2955 99.5127
R2643 vdd.n2952 vdd.n2951 99.5127
R2644 vdd.n2948 vdd.n2947 99.5127
R2645 vdd.n2943 vdd.n2942 99.5127
R2646 vdd.n2700 vdd.n970 99.5127
R2647 vdd.n2696 vdd.n2695 99.5127
R2648 vdd.n2692 vdd.n2691 99.5127
R2649 vdd.n2688 vdd.n2687 99.5127
R2650 vdd.n2684 vdd.n2683 99.5127
R2651 vdd.n2680 vdd.n2679 99.5127
R2652 vdd.n2676 vdd.n2675 99.5127
R2653 vdd.n2672 vdd.n2671 99.5127
R2654 vdd.n2668 vdd.n2667 99.5127
R2655 vdd.n2664 vdd.n2663 99.5127
R2656 vdd.n2660 vdd.n2659 99.5127
R2657 vdd.n2656 vdd.n2655 99.5127
R2658 vdd.n2652 vdd.n2651 99.5127
R2659 vdd.n2648 vdd.n2647 99.5127
R2660 vdd.n2644 vdd.n2643 99.5127
R2661 vdd.n2640 vdd.n2639 99.5127
R2662 vdd.n2635 vdd.n2634 99.5127
R2663 vdd.n1326 vdd.n1106 99.5127
R2664 vdd.n1329 vdd.n1106 99.5127
R2665 vdd.n1329 vdd.n1100 99.5127
R2666 vdd.n1332 vdd.n1100 99.5127
R2667 vdd.n1332 vdd.n1095 99.5127
R2668 vdd.n1335 vdd.n1095 99.5127
R2669 vdd.n1335 vdd.n1088 99.5127
R2670 vdd.n1338 vdd.n1088 99.5127
R2671 vdd.n1338 vdd.n1081 99.5127
R2672 vdd.n1341 vdd.n1081 99.5127
R2673 vdd.n1341 vdd.n1075 99.5127
R2674 vdd.n1344 vdd.n1075 99.5127
R2675 vdd.n1344 vdd.n1070 99.5127
R2676 vdd.n1347 vdd.n1070 99.5127
R2677 vdd.n1347 vdd.n1065 99.5127
R2678 vdd.n1350 vdd.n1065 99.5127
R2679 vdd.n1350 vdd.n1059 99.5127
R2680 vdd.n1353 vdd.n1059 99.5127
R2681 vdd.n1353 vdd.n1052 99.5127
R2682 vdd.n1356 vdd.n1052 99.5127
R2683 vdd.n1356 vdd.n1045 99.5127
R2684 vdd.n1359 vdd.n1045 99.5127
R2685 vdd.n1359 vdd.n1039 99.5127
R2686 vdd.n1362 vdd.n1039 99.5127
R2687 vdd.n1362 vdd.n1034 99.5127
R2688 vdd.n1365 vdd.n1034 99.5127
R2689 vdd.n1365 vdd.n1028 99.5127
R2690 vdd.n1407 vdd.n1028 99.5127
R2691 vdd.n1407 vdd.n1021 99.5127
R2692 vdd.n1403 vdd.n1021 99.5127
R2693 vdd.n1403 vdd.n1015 99.5127
R2694 vdd.n1400 vdd.n1015 99.5127
R2695 vdd.n1400 vdd.n1010 99.5127
R2696 vdd.n1397 vdd.n1010 99.5127
R2697 vdd.n1397 vdd.n1005 99.5127
R2698 vdd.n1377 vdd.n1005 99.5127
R2699 vdd.n1377 vdd.n1000 99.5127
R2700 vdd.n1374 vdd.n1000 99.5127
R2701 vdd.n1374 vdd.n993 99.5127
R2702 vdd.n1371 vdd.n993 99.5127
R2703 vdd.n1371 vdd.n986 99.5127
R2704 vdd.n986 vdd.n975 99.5127
R2705 vdd.n2630 vdd.n975 99.5127
R2706 vdd.n2422 vdd.n1111 99.5127
R2707 vdd.n2422 vdd.n1147 99.5127
R2708 vdd.n2418 vdd.n2417 99.5127
R2709 vdd.n2414 vdd.n2413 99.5127
R2710 vdd.n2410 vdd.n2409 99.5127
R2711 vdd.n2406 vdd.n2405 99.5127
R2712 vdd.n2402 vdd.n2401 99.5127
R2713 vdd.n2398 vdd.n2397 99.5127
R2714 vdd.n2394 vdd.n2393 99.5127
R2715 vdd.n1293 vdd.n1292 99.5127
R2716 vdd.n1297 vdd.n1296 99.5127
R2717 vdd.n1301 vdd.n1300 99.5127
R2718 vdd.n1305 vdd.n1304 99.5127
R2719 vdd.n1309 vdd.n1308 99.5127
R2720 vdd.n1313 vdd.n1312 99.5127
R2721 vdd.n1317 vdd.n1316 99.5127
R2722 vdd.n1322 vdd.n1321 99.5127
R2723 vdd.n2429 vdd.n1109 99.5127
R2724 vdd.n2429 vdd.n1099 99.5127
R2725 vdd.n2437 vdd.n1099 99.5127
R2726 vdd.n2437 vdd.n1097 99.5127
R2727 vdd.n2441 vdd.n1097 99.5127
R2728 vdd.n2441 vdd.n1086 99.5127
R2729 vdd.n2449 vdd.n1086 99.5127
R2730 vdd.n2449 vdd.n1084 99.5127
R2731 vdd.n2453 vdd.n1084 99.5127
R2732 vdd.n2453 vdd.n1074 99.5127
R2733 vdd.n2461 vdd.n1074 99.5127
R2734 vdd.n2461 vdd.n1072 99.5127
R2735 vdd.n2465 vdd.n1072 99.5127
R2736 vdd.n2465 vdd.n1063 99.5127
R2737 vdd.n2473 vdd.n1063 99.5127
R2738 vdd.n2473 vdd.n1061 99.5127
R2739 vdd.n2477 vdd.n1061 99.5127
R2740 vdd.n2477 vdd.n1050 99.5127
R2741 vdd.n2485 vdd.n1050 99.5127
R2742 vdd.n2485 vdd.n1048 99.5127
R2743 vdd.n2489 vdd.n1048 99.5127
R2744 vdd.n2489 vdd.n1038 99.5127
R2745 vdd.n2498 vdd.n1038 99.5127
R2746 vdd.n2498 vdd.n1036 99.5127
R2747 vdd.n2502 vdd.n1036 99.5127
R2748 vdd.n2502 vdd.n1026 99.5127
R2749 vdd.n2510 vdd.n1026 99.5127
R2750 vdd.n2510 vdd.n1024 99.5127
R2751 vdd.n2514 vdd.n1024 99.5127
R2752 vdd.n2514 vdd.n1014 99.5127
R2753 vdd.n2522 vdd.n1014 99.5127
R2754 vdd.n2522 vdd.n1012 99.5127
R2755 vdd.n2526 vdd.n1012 99.5127
R2756 vdd.n2526 vdd.n1004 99.5127
R2757 vdd.n2534 vdd.n1004 99.5127
R2758 vdd.n2534 vdd.n1002 99.5127
R2759 vdd.n2538 vdd.n1002 99.5127
R2760 vdd.n2538 vdd.n991 99.5127
R2761 vdd.n2548 vdd.n991 99.5127
R2762 vdd.n2548 vdd.n988 99.5127
R2763 vdd.n2553 vdd.n988 99.5127
R2764 vdd.n2553 vdd.n989 99.5127
R2765 vdd.n989 vdd.n969 99.5127
R2766 vdd.n3163 vdd.n3162 99.5127
R2767 vdd.n3160 vdd.n3126 99.5127
R2768 vdd.n3156 vdd.n3155 99.5127
R2769 vdd.n3153 vdd.n3129 99.5127
R2770 vdd.n3149 vdd.n3148 99.5127
R2771 vdd.n3146 vdd.n3132 99.5127
R2772 vdd.n3142 vdd.n3141 99.5127
R2773 vdd.n3139 vdd.n3136 99.5127
R2774 vdd.n3280 vdd.n755 99.5127
R2775 vdd.n3278 vdd.n3277 99.5127
R2776 vdd.n3275 vdd.n758 99.5127
R2777 vdd.n3271 vdd.n3270 99.5127
R2778 vdd.n3268 vdd.n761 99.5127
R2779 vdd.n3264 vdd.n3263 99.5127
R2780 vdd.n3261 vdd.n764 99.5127
R2781 vdd.n3257 vdd.n3256 99.5127
R2782 vdd.n3254 vdd.n767 99.5127
R2783 vdd.n2812 vdd.n930 99.5127
R2784 vdd.n2932 vdd.n930 99.5127
R2785 vdd.n2932 vdd.n924 99.5127
R2786 vdd.n2928 vdd.n924 99.5127
R2787 vdd.n2928 vdd.n919 99.5127
R2788 vdd.n2925 vdd.n919 99.5127
R2789 vdd.n2925 vdd.n913 99.5127
R2790 vdd.n2922 vdd.n913 99.5127
R2791 vdd.n2922 vdd.n907 99.5127
R2792 vdd.n2914 vdd.n907 99.5127
R2793 vdd.n2914 vdd.n901 99.5127
R2794 vdd.n2910 vdd.n901 99.5127
R2795 vdd.n2910 vdd.n895 99.5127
R2796 vdd.n2907 vdd.n895 99.5127
R2797 vdd.n2907 vdd.n890 99.5127
R2798 vdd.n2904 vdd.n890 99.5127
R2799 vdd.n2904 vdd.n885 99.5127
R2800 vdd.n2901 vdd.n885 99.5127
R2801 vdd.n2901 vdd.n878 99.5127
R2802 vdd.n2898 vdd.n878 99.5127
R2803 vdd.n2898 vdd.n871 99.5127
R2804 vdd.n2895 vdd.n871 99.5127
R2805 vdd.n2895 vdd.n865 99.5127
R2806 vdd.n2892 vdd.n865 99.5127
R2807 vdd.n2892 vdd.n860 99.5127
R2808 vdd.n2889 vdd.n860 99.5127
R2809 vdd.n2889 vdd.n854 99.5127
R2810 vdd.n2886 vdd.n854 99.5127
R2811 vdd.n2886 vdd.n847 99.5127
R2812 vdd.n2883 vdd.n847 99.5127
R2813 vdd.n2883 vdd.n840 99.5127
R2814 vdd.n2880 vdd.n840 99.5127
R2815 vdd.n2880 vdd.n834 99.5127
R2816 vdd.n2877 vdd.n834 99.5127
R2817 vdd.n2877 vdd.n829 99.5127
R2818 vdd.n2874 vdd.n829 99.5127
R2819 vdd.n2874 vdd.n824 99.5127
R2820 vdd.n2871 vdd.n824 99.5127
R2821 vdd.n2871 vdd.n816 99.5127
R2822 vdd.n2868 vdd.n816 99.5127
R2823 vdd.n2868 vdd.n809 99.5127
R2824 vdd.n809 vdd.n773 99.5127
R2825 vdd.n3249 vdd.n773 99.5127
R2826 vdd.n2747 vdd.n2746 99.5127
R2827 vdd.n2751 vdd.n2750 99.5127
R2828 vdd.n2755 vdd.n2754 99.5127
R2829 vdd.n2759 vdd.n2758 99.5127
R2830 vdd.n2763 vdd.n2762 99.5127
R2831 vdd.n2767 vdd.n2766 99.5127
R2832 vdd.n2771 vdd.n2770 99.5127
R2833 vdd.n2775 vdd.n2774 99.5127
R2834 vdd.n2779 vdd.n2778 99.5127
R2835 vdd.n2783 vdd.n2782 99.5127
R2836 vdd.n2787 vdd.n2786 99.5127
R2837 vdd.n2791 vdd.n2790 99.5127
R2838 vdd.n2795 vdd.n2794 99.5127
R2839 vdd.n2799 vdd.n2798 99.5127
R2840 vdd.n2803 vdd.n2802 99.5127
R2841 vdd.n2807 vdd.n2806 99.5127
R2842 vdd.n2809 vdd.n2735 99.5127
R2843 vdd.n3013 vdd.n927 99.5127
R2844 vdd.n3013 vdd.n925 99.5127
R2845 vdd.n3017 vdd.n925 99.5127
R2846 vdd.n3017 vdd.n916 99.5127
R2847 vdd.n3025 vdd.n916 99.5127
R2848 vdd.n3025 vdd.n914 99.5127
R2849 vdd.n3029 vdd.n914 99.5127
R2850 vdd.n3029 vdd.n905 99.5127
R2851 vdd.n3037 vdd.n905 99.5127
R2852 vdd.n3037 vdd.n903 99.5127
R2853 vdd.n3041 vdd.n903 99.5127
R2854 vdd.n3041 vdd.n893 99.5127
R2855 vdd.n3049 vdd.n893 99.5127
R2856 vdd.n3049 vdd.n891 99.5127
R2857 vdd.n3053 vdd.n891 99.5127
R2858 vdd.n3053 vdd.n882 99.5127
R2859 vdd.n3061 vdd.n882 99.5127
R2860 vdd.n3061 vdd.n880 99.5127
R2861 vdd.n3066 vdd.n880 99.5127
R2862 vdd.n3066 vdd.n869 99.5127
R2863 vdd.n3074 vdd.n869 99.5127
R2864 vdd.n3074 vdd.n866 99.5127
R2865 vdd.n3078 vdd.n866 99.5127
R2866 vdd.n3078 vdd.n857 99.5127
R2867 vdd.n3086 vdd.n857 99.5127
R2868 vdd.n3086 vdd.n855 99.5127
R2869 vdd.n3090 vdd.n855 99.5127
R2870 vdd.n3090 vdd.n844 99.5127
R2871 vdd.n3098 vdd.n844 99.5127
R2872 vdd.n3098 vdd.n842 99.5127
R2873 vdd.n3102 vdd.n842 99.5127
R2874 vdd.n3102 vdd.n832 99.5127
R2875 vdd.n3110 vdd.n832 99.5127
R2876 vdd.n3110 vdd.n830 99.5127
R2877 vdd.n3114 vdd.n830 99.5127
R2878 vdd.n3114 vdd.n821 99.5127
R2879 vdd.n3122 vdd.n821 99.5127
R2880 vdd.n3122 vdd.n818 99.5127
R2881 vdd.n3171 vdd.n818 99.5127
R2882 vdd.n3171 vdd.n819 99.5127
R2883 vdd.n819 vdd.n810 99.5127
R2884 vdd.n3166 vdd.n810 99.5127
R2885 vdd.n3166 vdd.n776 99.5127
R2886 vdd.n2624 vdd.n2623 99.5127
R2887 vdd.n2620 vdd.n2619 99.5127
R2888 vdd.n2616 vdd.n2615 99.5127
R2889 vdd.n2612 vdd.n2611 99.5127
R2890 vdd.n2608 vdd.n2607 99.5127
R2891 vdd.n2604 vdd.n2603 99.5127
R2892 vdd.n2600 vdd.n2599 99.5127
R2893 vdd.n2596 vdd.n2595 99.5127
R2894 vdd.n2592 vdd.n2591 99.5127
R2895 vdd.n2588 vdd.n2587 99.5127
R2896 vdd.n2584 vdd.n2583 99.5127
R2897 vdd.n2580 vdd.n2579 99.5127
R2898 vdd.n2576 vdd.n2575 99.5127
R2899 vdd.n2572 vdd.n2571 99.5127
R2900 vdd.n2568 vdd.n2567 99.5127
R2901 vdd.n2564 vdd.n2563 99.5127
R2902 vdd.n2560 vdd.n951 99.5127
R2903 vdd.n1451 vdd.n1107 99.5127
R2904 vdd.n1448 vdd.n1107 99.5127
R2905 vdd.n1448 vdd.n1101 99.5127
R2906 vdd.n1445 vdd.n1101 99.5127
R2907 vdd.n1445 vdd.n1096 99.5127
R2908 vdd.n1442 vdd.n1096 99.5127
R2909 vdd.n1442 vdd.n1089 99.5127
R2910 vdd.n1439 vdd.n1089 99.5127
R2911 vdd.n1439 vdd.n1082 99.5127
R2912 vdd.n1436 vdd.n1082 99.5127
R2913 vdd.n1436 vdd.n1076 99.5127
R2914 vdd.n1433 vdd.n1076 99.5127
R2915 vdd.n1433 vdd.n1071 99.5127
R2916 vdd.n1430 vdd.n1071 99.5127
R2917 vdd.n1430 vdd.n1066 99.5127
R2918 vdd.n1427 vdd.n1066 99.5127
R2919 vdd.n1427 vdd.n1060 99.5127
R2920 vdd.n1424 vdd.n1060 99.5127
R2921 vdd.n1424 vdd.n1053 99.5127
R2922 vdd.n1421 vdd.n1053 99.5127
R2923 vdd.n1421 vdd.n1046 99.5127
R2924 vdd.n1418 vdd.n1046 99.5127
R2925 vdd.n1418 vdd.n1040 99.5127
R2926 vdd.n1415 vdd.n1040 99.5127
R2927 vdd.n1415 vdd.n1035 99.5127
R2928 vdd.n1412 vdd.n1035 99.5127
R2929 vdd.n1412 vdd.n1029 99.5127
R2930 vdd.n1409 vdd.n1029 99.5127
R2931 vdd.n1409 vdd.n1022 99.5127
R2932 vdd.n1380 vdd.n1022 99.5127
R2933 vdd.n1380 vdd.n1016 99.5127
R2934 vdd.n1383 vdd.n1016 99.5127
R2935 vdd.n1383 vdd.n1011 99.5127
R2936 vdd.n1395 vdd.n1011 99.5127
R2937 vdd.n1395 vdd.n1006 99.5127
R2938 vdd.n1391 vdd.n1006 99.5127
R2939 vdd.n1391 vdd.n1001 99.5127
R2940 vdd.n1388 vdd.n1001 99.5127
R2941 vdd.n1388 vdd.n994 99.5127
R2942 vdd.n994 vdd.n985 99.5127
R2943 vdd.n2555 vdd.n985 99.5127
R2944 vdd.n2556 vdd.n2555 99.5127
R2945 vdd.n2556 vdd.n977 99.5127
R2946 vdd.n1255 vdd.n1254 99.5127
R2947 vdd.n1259 vdd.n1258 99.5127
R2948 vdd.n1263 vdd.n1262 99.5127
R2949 vdd.n1267 vdd.n1266 99.5127
R2950 vdd.n1271 vdd.n1270 99.5127
R2951 vdd.n1275 vdd.n1274 99.5127
R2952 vdd.n1279 vdd.n1278 99.5127
R2953 vdd.n1283 vdd.n1282 99.5127
R2954 vdd.n1484 vdd.n1285 99.5127
R2955 vdd.n1482 vdd.n1481 99.5127
R2956 vdd.n1478 vdd.n1477 99.5127
R2957 vdd.n1474 vdd.n1473 99.5127
R2958 vdd.n1470 vdd.n1469 99.5127
R2959 vdd.n1466 vdd.n1465 99.5127
R2960 vdd.n1462 vdd.n1461 99.5127
R2961 vdd.n1458 vdd.n1457 99.5127
R2962 vdd.n1454 vdd.n1146 99.5127
R2963 vdd.n2431 vdd.n1104 99.5127
R2964 vdd.n2431 vdd.n1102 99.5127
R2965 vdd.n2435 vdd.n1102 99.5127
R2966 vdd.n2435 vdd.n1093 99.5127
R2967 vdd.n2443 vdd.n1093 99.5127
R2968 vdd.n2443 vdd.n1091 99.5127
R2969 vdd.n2447 vdd.n1091 99.5127
R2970 vdd.n2447 vdd.n1080 99.5127
R2971 vdd.n2455 vdd.n1080 99.5127
R2972 vdd.n2455 vdd.n1078 99.5127
R2973 vdd.n2459 vdd.n1078 99.5127
R2974 vdd.n2459 vdd.n1069 99.5127
R2975 vdd.n2467 vdd.n1069 99.5127
R2976 vdd.n2467 vdd.n1067 99.5127
R2977 vdd.n2471 vdd.n1067 99.5127
R2978 vdd.n2471 vdd.n1057 99.5127
R2979 vdd.n2479 vdd.n1057 99.5127
R2980 vdd.n2479 vdd.n1055 99.5127
R2981 vdd.n2483 vdd.n1055 99.5127
R2982 vdd.n2483 vdd.n1044 99.5127
R2983 vdd.n2491 vdd.n1044 99.5127
R2984 vdd.n2491 vdd.n1041 99.5127
R2985 vdd.n2496 vdd.n1041 99.5127
R2986 vdd.n2496 vdd.n1032 99.5127
R2987 vdd.n2504 vdd.n1032 99.5127
R2988 vdd.n2504 vdd.n1030 99.5127
R2989 vdd.n2508 vdd.n1030 99.5127
R2990 vdd.n2508 vdd.n1020 99.5127
R2991 vdd.n2516 vdd.n1020 99.5127
R2992 vdd.n2516 vdd.n1018 99.5127
R2993 vdd.n2520 vdd.n1018 99.5127
R2994 vdd.n2520 vdd.n1009 99.5127
R2995 vdd.n2528 vdd.n1009 99.5127
R2996 vdd.n2528 vdd.n1007 99.5127
R2997 vdd.n2532 vdd.n1007 99.5127
R2998 vdd.n2532 vdd.n998 99.5127
R2999 vdd.n2540 vdd.n998 99.5127
R3000 vdd.n2540 vdd.n995 99.5127
R3001 vdd.n2546 vdd.n995 99.5127
R3002 vdd.n2546 vdd.n996 99.5127
R3003 vdd.n996 vdd.n987 99.5127
R3004 vdd.n987 vdd.n978 99.5127
R3005 vdd.n2628 vdd.n978 99.5127
R3006 vdd.n9 vdd.n7 98.9633
R3007 vdd.n2 vdd.n0 98.9633
R3008 vdd.n9 vdd.n8 98.6055
R3009 vdd.n11 vdd.n10 98.6055
R3010 vdd.n13 vdd.n12 98.6055
R3011 vdd.n6 vdd.n5 98.6055
R3012 vdd.n4 vdd.n3 98.6055
R3013 vdd.n2 vdd.n1 98.6055
R3014 vdd.t57 vdd.n291 85.8723
R3015 vdd.t52 vdd.n236 85.8723
R3016 vdd.t148 vdd.n193 85.8723
R3017 vdd.t273 vdd.n138 85.8723
R3018 vdd.t160 vdd.n96 85.8723
R3019 vdd.t175 vdd.n41 85.8723
R3020 vdd.t166 vdd.n2115 85.8723
R3021 vdd.t48 vdd.n2170 85.8723
R3022 vdd.t185 vdd.n2017 85.8723
R3023 vdd.t177 vdd.n2072 85.8723
R3024 vdd.t174 vdd.n1920 85.8723
R3025 vdd.t168 vdd.n1975 85.8723
R3026 vdd.n868 vdd.n867 78.546
R3027 vdd.n2494 vdd.n1042 78.546
R3028 vdd.n278 vdd.n277 75.1835
R3029 vdd.n276 vdd.n275 75.1835
R3030 vdd.n274 vdd.n273 75.1835
R3031 vdd.n272 vdd.n271 75.1835
R3032 vdd.n270 vdd.n269 75.1835
R3033 vdd.n268 vdd.n267 75.1835
R3034 vdd.n266 vdd.n265 75.1835
R3035 vdd.n180 vdd.n179 75.1835
R3036 vdd.n178 vdd.n177 75.1835
R3037 vdd.n176 vdd.n175 75.1835
R3038 vdd.n174 vdd.n173 75.1835
R3039 vdd.n172 vdd.n171 75.1835
R3040 vdd.n170 vdd.n169 75.1835
R3041 vdd.n168 vdd.n167 75.1835
R3042 vdd.n83 vdd.n82 75.1835
R3043 vdd.n81 vdd.n80 75.1835
R3044 vdd.n79 vdd.n78 75.1835
R3045 vdd.n77 vdd.n76 75.1835
R3046 vdd.n75 vdd.n74 75.1835
R3047 vdd.n73 vdd.n72 75.1835
R3048 vdd.n71 vdd.n70 75.1835
R3049 vdd.n2145 vdd.n2144 75.1835
R3050 vdd.n2147 vdd.n2146 75.1835
R3051 vdd.n2149 vdd.n2148 75.1835
R3052 vdd.n2151 vdd.n2150 75.1835
R3053 vdd.n2153 vdd.n2152 75.1835
R3054 vdd.n2155 vdd.n2154 75.1835
R3055 vdd.n2157 vdd.n2156 75.1835
R3056 vdd.n2047 vdd.n2046 75.1835
R3057 vdd.n2049 vdd.n2048 75.1835
R3058 vdd.n2051 vdd.n2050 75.1835
R3059 vdd.n2053 vdd.n2052 75.1835
R3060 vdd.n2055 vdd.n2054 75.1835
R3061 vdd.n2057 vdd.n2056 75.1835
R3062 vdd.n2059 vdd.n2058 75.1835
R3063 vdd.n1950 vdd.n1949 75.1835
R3064 vdd.n1952 vdd.n1951 75.1835
R3065 vdd.n1954 vdd.n1953 75.1835
R3066 vdd.n1956 vdd.n1955 75.1835
R3067 vdd.n1958 vdd.n1957 75.1835
R3068 vdd.n1960 vdd.n1959 75.1835
R3069 vdd.n1962 vdd.n1961 75.1835
R3070 vdd.n3005 vdd.n2718 72.8958
R3071 vdd.n3005 vdd.n2719 72.8958
R3072 vdd.n3005 vdd.n2720 72.8958
R3073 vdd.n3005 vdd.n2721 72.8958
R3074 vdd.n3005 vdd.n2722 72.8958
R3075 vdd.n3005 vdd.n2723 72.8958
R3076 vdd.n3005 vdd.n2724 72.8958
R3077 vdd.n3005 vdd.n2725 72.8958
R3078 vdd.n3005 vdd.n2726 72.8958
R3079 vdd.n3005 vdd.n2727 72.8958
R3080 vdd.n3005 vdd.n2728 72.8958
R3081 vdd.n3005 vdd.n2729 72.8958
R3082 vdd.n3005 vdd.n2730 72.8958
R3083 vdd.n3005 vdd.n2731 72.8958
R3084 vdd.n3005 vdd.n2732 72.8958
R3085 vdd.n3005 vdd.n2733 72.8958
R3086 vdd.n3005 vdd.n2734 72.8958
R3087 vdd.n772 vdd.n756 72.8958
R3088 vdd.n3255 vdd.n756 72.8958
R3089 vdd.n766 vdd.n756 72.8958
R3090 vdd.n3262 vdd.n756 72.8958
R3091 vdd.n763 vdd.n756 72.8958
R3092 vdd.n3269 vdd.n756 72.8958
R3093 vdd.n760 vdd.n756 72.8958
R3094 vdd.n3276 vdd.n756 72.8958
R3095 vdd.n3279 vdd.n756 72.8958
R3096 vdd.n3135 vdd.n756 72.8958
R3097 vdd.n3140 vdd.n756 72.8958
R3098 vdd.n3134 vdd.n756 72.8958
R3099 vdd.n3147 vdd.n756 72.8958
R3100 vdd.n3131 vdd.n756 72.8958
R3101 vdd.n3154 vdd.n756 72.8958
R3102 vdd.n3128 vdd.n756 72.8958
R3103 vdd.n3161 vdd.n756 72.8958
R3104 vdd.n2424 vdd.n2423 72.8958
R3105 vdd.n2423 vdd.n1113 72.8958
R3106 vdd.n2423 vdd.n1114 72.8958
R3107 vdd.n2423 vdd.n1115 72.8958
R3108 vdd.n2423 vdd.n1116 72.8958
R3109 vdd.n2423 vdd.n1117 72.8958
R3110 vdd.n2423 vdd.n1118 72.8958
R3111 vdd.n2423 vdd.n1119 72.8958
R3112 vdd.n2423 vdd.n1120 72.8958
R3113 vdd.n2423 vdd.n1121 72.8958
R3114 vdd.n2423 vdd.n1122 72.8958
R3115 vdd.n2423 vdd.n1123 72.8958
R3116 vdd.n2423 vdd.n1124 72.8958
R3117 vdd.n2423 vdd.n1125 72.8958
R3118 vdd.n2423 vdd.n1126 72.8958
R3119 vdd.n2423 vdd.n1127 72.8958
R3120 vdd.n2423 vdd.n1128 72.8958
R3121 vdd.n2701 vdd.n952 72.8958
R3122 vdd.n2701 vdd.n953 72.8958
R3123 vdd.n2701 vdd.n954 72.8958
R3124 vdd.n2701 vdd.n955 72.8958
R3125 vdd.n2701 vdd.n956 72.8958
R3126 vdd.n2701 vdd.n957 72.8958
R3127 vdd.n2701 vdd.n958 72.8958
R3128 vdd.n2701 vdd.n959 72.8958
R3129 vdd.n2701 vdd.n960 72.8958
R3130 vdd.n2701 vdd.n961 72.8958
R3131 vdd.n2701 vdd.n962 72.8958
R3132 vdd.n2701 vdd.n963 72.8958
R3133 vdd.n2701 vdd.n964 72.8958
R3134 vdd.n2701 vdd.n965 72.8958
R3135 vdd.n2701 vdd.n966 72.8958
R3136 vdd.n2701 vdd.n967 72.8958
R3137 vdd.n2701 vdd.n968 72.8958
R3138 vdd.n3006 vdd.n3005 72.8958
R3139 vdd.n3005 vdd.n2702 72.8958
R3140 vdd.n3005 vdd.n2703 72.8958
R3141 vdd.n3005 vdd.n2704 72.8958
R3142 vdd.n3005 vdd.n2705 72.8958
R3143 vdd.n3005 vdd.n2706 72.8958
R3144 vdd.n3005 vdd.n2707 72.8958
R3145 vdd.n3005 vdd.n2708 72.8958
R3146 vdd.n3005 vdd.n2709 72.8958
R3147 vdd.n3005 vdd.n2710 72.8958
R3148 vdd.n3005 vdd.n2711 72.8958
R3149 vdd.n3005 vdd.n2712 72.8958
R3150 vdd.n3005 vdd.n2713 72.8958
R3151 vdd.n3005 vdd.n2714 72.8958
R3152 vdd.n3005 vdd.n2715 72.8958
R3153 vdd.n3005 vdd.n2716 72.8958
R3154 vdd.n3005 vdd.n2717 72.8958
R3155 vdd.n3183 vdd.n756 72.8958
R3156 vdd.n3189 vdd.n756 72.8958
R3157 vdd.n802 vdd.n756 72.8958
R3158 vdd.n3196 vdd.n756 72.8958
R3159 vdd.n799 vdd.n756 72.8958
R3160 vdd.n3203 vdd.n756 72.8958
R3161 vdd.n796 vdd.n756 72.8958
R3162 vdd.n3210 vdd.n756 72.8958
R3163 vdd.n793 vdd.n756 72.8958
R3164 vdd.n3218 vdd.n756 72.8958
R3165 vdd.n790 vdd.n756 72.8958
R3166 vdd.n3225 vdd.n756 72.8958
R3167 vdd.n787 vdd.n756 72.8958
R3168 vdd.n3232 vdd.n756 72.8958
R3169 vdd.n784 vdd.n756 72.8958
R3170 vdd.n3239 vdd.n756 72.8958
R3171 vdd.n3242 vdd.n756 72.8958
R3172 vdd.n2701 vdd.n950 72.8958
R3173 vdd.n2701 vdd.n949 72.8958
R3174 vdd.n2701 vdd.n948 72.8958
R3175 vdd.n2701 vdd.n947 72.8958
R3176 vdd.n2701 vdd.n946 72.8958
R3177 vdd.n2701 vdd.n945 72.8958
R3178 vdd.n2701 vdd.n944 72.8958
R3179 vdd.n2701 vdd.n943 72.8958
R3180 vdd.n2701 vdd.n942 72.8958
R3181 vdd.n2701 vdd.n941 72.8958
R3182 vdd.n2701 vdd.n940 72.8958
R3183 vdd.n2701 vdd.n939 72.8958
R3184 vdd.n2701 vdd.n938 72.8958
R3185 vdd.n2701 vdd.n937 72.8958
R3186 vdd.n2701 vdd.n936 72.8958
R3187 vdd.n2701 vdd.n935 72.8958
R3188 vdd.n2701 vdd.n934 72.8958
R3189 vdd.n2423 vdd.n1129 72.8958
R3190 vdd.n2423 vdd.n1130 72.8958
R3191 vdd.n2423 vdd.n1131 72.8958
R3192 vdd.n2423 vdd.n1132 72.8958
R3193 vdd.n2423 vdd.n1133 72.8958
R3194 vdd.n2423 vdd.n1134 72.8958
R3195 vdd.n2423 vdd.n1135 72.8958
R3196 vdd.n2423 vdd.n1136 72.8958
R3197 vdd.n2423 vdd.n1137 72.8958
R3198 vdd.n2423 vdd.n1138 72.8958
R3199 vdd.n2423 vdd.n1139 72.8958
R3200 vdd.n2423 vdd.n1140 72.8958
R3201 vdd.n2423 vdd.n1141 72.8958
R3202 vdd.n2423 vdd.n1142 72.8958
R3203 vdd.n2423 vdd.n1143 72.8958
R3204 vdd.n2423 vdd.n1144 72.8958
R3205 vdd.n2423 vdd.n1145 72.8958
R3206 vdd.n1829 vdd.n1828 66.2847
R3207 vdd.n1829 vdd.n1607 66.2847
R3208 vdd.n1829 vdd.n1608 66.2847
R3209 vdd.n1829 vdd.n1609 66.2847
R3210 vdd.n1829 vdd.n1610 66.2847
R3211 vdd.n1829 vdd.n1611 66.2847
R3212 vdd.n1829 vdd.n1612 66.2847
R3213 vdd.n1829 vdd.n1613 66.2847
R3214 vdd.n1829 vdd.n1614 66.2847
R3215 vdd.n1829 vdd.n1615 66.2847
R3216 vdd.n1829 vdd.n1616 66.2847
R3217 vdd.n1829 vdd.n1617 66.2847
R3218 vdd.n1829 vdd.n1618 66.2847
R3219 vdd.n1829 vdd.n1619 66.2847
R3220 vdd.n1829 vdd.n1620 66.2847
R3221 vdd.n1829 vdd.n1621 66.2847
R3222 vdd.n1829 vdd.n1622 66.2847
R3223 vdd.n1829 vdd.n1623 66.2847
R3224 vdd.n1829 vdd.n1624 66.2847
R3225 vdd.n1829 vdd.n1625 66.2847
R3226 vdd.n1829 vdd.n1626 66.2847
R3227 vdd.n1829 vdd.n1627 66.2847
R3228 vdd.n1829 vdd.n1628 66.2847
R3229 vdd.n1829 vdd.n1629 66.2847
R3230 vdd.n1829 vdd.n1630 66.2847
R3231 vdd.n1829 vdd.n1631 66.2847
R3232 vdd.n1829 vdd.n1632 66.2847
R3233 vdd.n1829 vdd.n1633 66.2847
R3234 vdd.n1829 vdd.n1634 66.2847
R3235 vdd.n1829 vdd.n1635 66.2847
R3236 vdd.n1829 vdd.n1636 66.2847
R3237 vdd.n1497 vdd.n1112 66.2847
R3238 vdd.n1494 vdd.n1112 66.2847
R3239 vdd.n1490 vdd.n1112 66.2847
R3240 vdd.n2289 vdd.n1112 66.2847
R3241 vdd.n1246 vdd.n1112 66.2847
R3242 vdd.n2296 vdd.n1112 66.2847
R3243 vdd.n1239 vdd.n1112 66.2847
R3244 vdd.n2303 vdd.n1112 66.2847
R3245 vdd.n1232 vdd.n1112 66.2847
R3246 vdd.n2310 vdd.n1112 66.2847
R3247 vdd.n1226 vdd.n1112 66.2847
R3248 vdd.n1221 vdd.n1112 66.2847
R3249 vdd.n2321 vdd.n1112 66.2847
R3250 vdd.n1213 vdd.n1112 66.2847
R3251 vdd.n2328 vdd.n1112 66.2847
R3252 vdd.n1206 vdd.n1112 66.2847
R3253 vdd.n2335 vdd.n1112 66.2847
R3254 vdd.n1199 vdd.n1112 66.2847
R3255 vdd.n2342 vdd.n1112 66.2847
R3256 vdd.n1192 vdd.n1112 66.2847
R3257 vdd.n2349 vdd.n1112 66.2847
R3258 vdd.n1186 vdd.n1112 66.2847
R3259 vdd.n1181 vdd.n1112 66.2847
R3260 vdd.n2360 vdd.n1112 66.2847
R3261 vdd.n1173 vdd.n1112 66.2847
R3262 vdd.n2367 vdd.n1112 66.2847
R3263 vdd.n1166 vdd.n1112 66.2847
R3264 vdd.n2374 vdd.n1112 66.2847
R3265 vdd.n1159 vdd.n1112 66.2847
R3266 vdd.n2381 vdd.n1112 66.2847
R3267 vdd.n2386 vdd.n1112 66.2847
R3268 vdd.n1155 vdd.n1112 66.2847
R3269 vdd.n3409 vdd.n658 66.2847
R3270 vdd.n663 vdd.n658 66.2847
R3271 vdd.n666 vdd.n658 66.2847
R3272 vdd.n3398 vdd.n658 66.2847
R3273 vdd.n3392 vdd.n658 66.2847
R3274 vdd.n3390 vdd.n658 66.2847
R3275 vdd.n3384 vdd.n658 66.2847
R3276 vdd.n3382 vdd.n658 66.2847
R3277 vdd.n3376 vdd.n658 66.2847
R3278 vdd.n3374 vdd.n658 66.2847
R3279 vdd.n3368 vdd.n658 66.2847
R3280 vdd.n3366 vdd.n658 66.2847
R3281 vdd.n3360 vdd.n658 66.2847
R3282 vdd.n3358 vdd.n658 66.2847
R3283 vdd.n3352 vdd.n658 66.2847
R3284 vdd.n3350 vdd.n658 66.2847
R3285 vdd.n3344 vdd.n658 66.2847
R3286 vdd.n3342 vdd.n658 66.2847
R3287 vdd.n3336 vdd.n658 66.2847
R3288 vdd.n3334 vdd.n658 66.2847
R3289 vdd.n727 vdd.n658 66.2847
R3290 vdd.n3325 vdd.n658 66.2847
R3291 vdd.n729 vdd.n658 66.2847
R3292 vdd.n3318 vdd.n658 66.2847
R3293 vdd.n3312 vdd.n658 66.2847
R3294 vdd.n3310 vdd.n658 66.2847
R3295 vdd.n3304 vdd.n658 66.2847
R3296 vdd.n3302 vdd.n658 66.2847
R3297 vdd.n3296 vdd.n658 66.2847
R3298 vdd.n750 vdd.n658 66.2847
R3299 vdd.n752 vdd.n658 66.2847
R3300 vdd.n3525 vdd.n3524 66.2847
R3301 vdd.n3525 vdd.n403 66.2847
R3302 vdd.n3525 vdd.n402 66.2847
R3303 vdd.n3525 vdd.n401 66.2847
R3304 vdd.n3525 vdd.n400 66.2847
R3305 vdd.n3525 vdd.n399 66.2847
R3306 vdd.n3525 vdd.n398 66.2847
R3307 vdd.n3525 vdd.n397 66.2847
R3308 vdd.n3525 vdd.n396 66.2847
R3309 vdd.n3525 vdd.n395 66.2847
R3310 vdd.n3525 vdd.n394 66.2847
R3311 vdd.n3525 vdd.n393 66.2847
R3312 vdd.n3525 vdd.n392 66.2847
R3313 vdd.n3525 vdd.n391 66.2847
R3314 vdd.n3525 vdd.n390 66.2847
R3315 vdd.n3525 vdd.n389 66.2847
R3316 vdd.n3525 vdd.n388 66.2847
R3317 vdd.n3525 vdd.n387 66.2847
R3318 vdd.n3525 vdd.n386 66.2847
R3319 vdd.n3525 vdd.n385 66.2847
R3320 vdd.n3525 vdd.n384 66.2847
R3321 vdd.n3525 vdd.n383 66.2847
R3322 vdd.n3525 vdd.n382 66.2847
R3323 vdd.n3525 vdd.n381 66.2847
R3324 vdd.n3525 vdd.n380 66.2847
R3325 vdd.n3525 vdd.n379 66.2847
R3326 vdd.n3525 vdd.n378 66.2847
R3327 vdd.n3525 vdd.n377 66.2847
R3328 vdd.n3525 vdd.n376 66.2847
R3329 vdd.n3525 vdd.n375 66.2847
R3330 vdd.n3525 vdd.n374 66.2847
R3331 vdd.n3525 vdd.n373 66.2847
R3332 vdd.n448 vdd.n373 52.4337
R3333 vdd.n454 vdd.n374 52.4337
R3334 vdd.n458 vdd.n375 52.4337
R3335 vdd.n464 vdd.n376 52.4337
R3336 vdd.n468 vdd.n377 52.4337
R3337 vdd.n474 vdd.n378 52.4337
R3338 vdd.n478 vdd.n379 52.4337
R3339 vdd.n484 vdd.n380 52.4337
R3340 vdd.n488 vdd.n381 52.4337
R3341 vdd.n494 vdd.n382 52.4337
R3342 vdd.n498 vdd.n383 52.4337
R3343 vdd.n504 vdd.n384 52.4337
R3344 vdd.n508 vdd.n385 52.4337
R3345 vdd.n514 vdd.n386 52.4337
R3346 vdd.n518 vdd.n387 52.4337
R3347 vdd.n524 vdd.n388 52.4337
R3348 vdd.n528 vdd.n389 52.4337
R3349 vdd.n534 vdd.n390 52.4337
R3350 vdd.n538 vdd.n391 52.4337
R3351 vdd.n544 vdd.n392 52.4337
R3352 vdd.n548 vdd.n393 52.4337
R3353 vdd.n554 vdd.n394 52.4337
R3354 vdd.n558 vdd.n395 52.4337
R3355 vdd.n564 vdd.n396 52.4337
R3356 vdd.n568 vdd.n397 52.4337
R3357 vdd.n574 vdd.n398 52.4337
R3358 vdd.n578 vdd.n399 52.4337
R3359 vdd.n584 vdd.n400 52.4337
R3360 vdd.n588 vdd.n401 52.4337
R3361 vdd.n594 vdd.n402 52.4337
R3362 vdd.n597 vdd.n403 52.4337
R3363 vdd.n3524 vdd.n3523 52.4337
R3364 vdd.n3409 vdd.n660 52.4337
R3365 vdd.n3407 vdd.n663 52.4337
R3366 vdd.n3403 vdd.n666 52.4337
R3367 vdd.n3399 vdd.n3398 52.4337
R3368 vdd.n3392 vdd.n669 52.4337
R3369 vdd.n3391 vdd.n3390 52.4337
R3370 vdd.n3384 vdd.n675 52.4337
R3371 vdd.n3383 vdd.n3382 52.4337
R3372 vdd.n3376 vdd.n681 52.4337
R3373 vdd.n3375 vdd.n3374 52.4337
R3374 vdd.n3368 vdd.n689 52.4337
R3375 vdd.n3367 vdd.n3366 52.4337
R3376 vdd.n3360 vdd.n695 52.4337
R3377 vdd.n3359 vdd.n3358 52.4337
R3378 vdd.n3352 vdd.n701 52.4337
R3379 vdd.n3351 vdd.n3350 52.4337
R3380 vdd.n3344 vdd.n707 52.4337
R3381 vdd.n3343 vdd.n3342 52.4337
R3382 vdd.n3336 vdd.n713 52.4337
R3383 vdd.n3335 vdd.n3334 52.4337
R3384 vdd.n727 vdd.n719 52.4337
R3385 vdd.n3326 vdd.n3325 52.4337
R3386 vdd.n3323 vdd.n729 52.4337
R3387 vdd.n3319 vdd.n3318 52.4337
R3388 vdd.n3312 vdd.n733 52.4337
R3389 vdd.n3311 vdd.n3310 52.4337
R3390 vdd.n3304 vdd.n739 52.4337
R3391 vdd.n3303 vdd.n3302 52.4337
R3392 vdd.n3296 vdd.n745 52.4337
R3393 vdd.n3295 vdd.n750 52.4337
R3394 vdd.n3291 vdd.n752 52.4337
R3395 vdd.n2388 vdd.n1155 52.4337
R3396 vdd.n2386 vdd.n2385 52.4337
R3397 vdd.n2381 vdd.n2380 52.4337
R3398 vdd.n2376 vdd.n1159 52.4337
R3399 vdd.n2374 vdd.n2373 52.4337
R3400 vdd.n2369 vdd.n1166 52.4337
R3401 vdd.n2367 vdd.n2366 52.4337
R3402 vdd.n2362 vdd.n1173 52.4337
R3403 vdd.n2360 vdd.n2359 52.4337
R3404 vdd.n1182 vdd.n1181 52.4337
R3405 vdd.n2351 vdd.n1186 52.4337
R3406 vdd.n2349 vdd.n2348 52.4337
R3407 vdd.n2344 vdd.n1192 52.4337
R3408 vdd.n2342 vdd.n2341 52.4337
R3409 vdd.n2337 vdd.n1199 52.4337
R3410 vdd.n2335 vdd.n2334 52.4337
R3411 vdd.n2330 vdd.n1206 52.4337
R3412 vdd.n2328 vdd.n2327 52.4337
R3413 vdd.n2323 vdd.n1213 52.4337
R3414 vdd.n2321 vdd.n2320 52.4337
R3415 vdd.n1222 vdd.n1221 52.4337
R3416 vdd.n2312 vdd.n1226 52.4337
R3417 vdd.n2310 vdd.n2309 52.4337
R3418 vdd.n2305 vdd.n1232 52.4337
R3419 vdd.n2303 vdd.n2302 52.4337
R3420 vdd.n2298 vdd.n1239 52.4337
R3421 vdd.n2296 vdd.n2295 52.4337
R3422 vdd.n2291 vdd.n1246 52.4337
R3423 vdd.n2289 vdd.n2288 52.4337
R3424 vdd.n1491 vdd.n1490 52.4337
R3425 vdd.n1495 vdd.n1494 52.4337
R3426 vdd.n2277 vdd.n1497 52.4337
R3427 vdd.n1828 vdd.n1827 52.4337
R3428 vdd.n1642 vdd.n1607 52.4337
R3429 vdd.n1644 vdd.n1608 52.4337
R3430 vdd.n1648 vdd.n1609 52.4337
R3431 vdd.n1650 vdd.n1610 52.4337
R3432 vdd.n1654 vdd.n1611 52.4337
R3433 vdd.n1656 vdd.n1612 52.4337
R3434 vdd.n1660 vdd.n1613 52.4337
R3435 vdd.n1662 vdd.n1614 52.4337
R3436 vdd.n1794 vdd.n1615 52.4337
R3437 vdd.n1666 vdd.n1616 52.4337
R3438 vdd.n1670 vdd.n1617 52.4337
R3439 vdd.n1672 vdd.n1618 52.4337
R3440 vdd.n1676 vdd.n1619 52.4337
R3441 vdd.n1678 vdd.n1620 52.4337
R3442 vdd.n1682 vdd.n1621 52.4337
R3443 vdd.n1684 vdd.n1622 52.4337
R3444 vdd.n1688 vdd.n1623 52.4337
R3445 vdd.n1690 vdd.n1624 52.4337
R3446 vdd.n1694 vdd.n1625 52.4337
R3447 vdd.n1758 vdd.n1626 52.4337
R3448 vdd.n1699 vdd.n1627 52.4337
R3449 vdd.n1701 vdd.n1628 52.4337
R3450 vdd.n1705 vdd.n1629 52.4337
R3451 vdd.n1707 vdd.n1630 52.4337
R3452 vdd.n1711 vdd.n1631 52.4337
R3453 vdd.n1713 vdd.n1632 52.4337
R3454 vdd.n1717 vdd.n1633 52.4337
R3455 vdd.n1719 vdd.n1634 52.4337
R3456 vdd.n1723 vdd.n1635 52.4337
R3457 vdd.n1725 vdd.n1636 52.4337
R3458 vdd.n1828 vdd.n1638 52.4337
R3459 vdd.n1643 vdd.n1607 52.4337
R3460 vdd.n1647 vdd.n1608 52.4337
R3461 vdd.n1649 vdd.n1609 52.4337
R3462 vdd.n1653 vdd.n1610 52.4337
R3463 vdd.n1655 vdd.n1611 52.4337
R3464 vdd.n1659 vdd.n1612 52.4337
R3465 vdd.n1661 vdd.n1613 52.4337
R3466 vdd.n1793 vdd.n1614 52.4337
R3467 vdd.n1665 vdd.n1615 52.4337
R3468 vdd.n1669 vdd.n1616 52.4337
R3469 vdd.n1671 vdd.n1617 52.4337
R3470 vdd.n1675 vdd.n1618 52.4337
R3471 vdd.n1677 vdd.n1619 52.4337
R3472 vdd.n1681 vdd.n1620 52.4337
R3473 vdd.n1683 vdd.n1621 52.4337
R3474 vdd.n1687 vdd.n1622 52.4337
R3475 vdd.n1689 vdd.n1623 52.4337
R3476 vdd.n1693 vdd.n1624 52.4337
R3477 vdd.n1695 vdd.n1625 52.4337
R3478 vdd.n1698 vdd.n1626 52.4337
R3479 vdd.n1700 vdd.n1627 52.4337
R3480 vdd.n1704 vdd.n1628 52.4337
R3481 vdd.n1706 vdd.n1629 52.4337
R3482 vdd.n1710 vdd.n1630 52.4337
R3483 vdd.n1712 vdd.n1631 52.4337
R3484 vdd.n1716 vdd.n1632 52.4337
R3485 vdd.n1718 vdd.n1633 52.4337
R3486 vdd.n1722 vdd.n1634 52.4337
R3487 vdd.n1724 vdd.n1635 52.4337
R3488 vdd.n1636 vdd.n1606 52.4337
R3489 vdd.n1497 vdd.n1496 52.4337
R3490 vdd.n1494 vdd.n1493 52.4337
R3491 vdd.n1490 vdd.n1247 52.4337
R3492 vdd.n2290 vdd.n2289 52.4337
R3493 vdd.n1246 vdd.n1240 52.4337
R3494 vdd.n2297 vdd.n2296 52.4337
R3495 vdd.n1239 vdd.n1233 52.4337
R3496 vdd.n2304 vdd.n2303 52.4337
R3497 vdd.n1232 vdd.n1227 52.4337
R3498 vdd.n2311 vdd.n2310 52.4337
R3499 vdd.n1226 vdd.n1225 52.4337
R3500 vdd.n1221 vdd.n1214 52.4337
R3501 vdd.n2322 vdd.n2321 52.4337
R3502 vdd.n1213 vdd.n1207 52.4337
R3503 vdd.n2329 vdd.n2328 52.4337
R3504 vdd.n1206 vdd.n1200 52.4337
R3505 vdd.n2336 vdd.n2335 52.4337
R3506 vdd.n1199 vdd.n1193 52.4337
R3507 vdd.n2343 vdd.n2342 52.4337
R3508 vdd.n1192 vdd.n1187 52.4337
R3509 vdd.n2350 vdd.n2349 52.4337
R3510 vdd.n1186 vdd.n1185 52.4337
R3511 vdd.n1181 vdd.n1174 52.4337
R3512 vdd.n2361 vdd.n2360 52.4337
R3513 vdd.n1173 vdd.n1167 52.4337
R3514 vdd.n2368 vdd.n2367 52.4337
R3515 vdd.n1166 vdd.n1160 52.4337
R3516 vdd.n2375 vdd.n2374 52.4337
R3517 vdd.n1159 vdd.n1156 52.4337
R3518 vdd.n2382 vdd.n2381 52.4337
R3519 vdd.n2387 vdd.n2386 52.4337
R3520 vdd.n1502 vdd.n1155 52.4337
R3521 vdd.n3410 vdd.n3409 52.4337
R3522 vdd.n3404 vdd.n663 52.4337
R3523 vdd.n3400 vdd.n666 52.4337
R3524 vdd.n3398 vdd.n3397 52.4337
R3525 vdd.n3393 vdd.n3392 52.4337
R3526 vdd.n3390 vdd.n3389 52.4337
R3527 vdd.n3385 vdd.n3384 52.4337
R3528 vdd.n3382 vdd.n3381 52.4337
R3529 vdd.n3377 vdd.n3376 52.4337
R3530 vdd.n3374 vdd.n3373 52.4337
R3531 vdd.n3369 vdd.n3368 52.4337
R3532 vdd.n3366 vdd.n3365 52.4337
R3533 vdd.n3361 vdd.n3360 52.4337
R3534 vdd.n3358 vdd.n3357 52.4337
R3535 vdd.n3353 vdd.n3352 52.4337
R3536 vdd.n3350 vdd.n3349 52.4337
R3537 vdd.n3345 vdd.n3344 52.4337
R3538 vdd.n3342 vdd.n3341 52.4337
R3539 vdd.n3337 vdd.n3336 52.4337
R3540 vdd.n3334 vdd.n3333 52.4337
R3541 vdd.n728 vdd.n727 52.4337
R3542 vdd.n3325 vdd.n3324 52.4337
R3543 vdd.n3320 vdd.n729 52.4337
R3544 vdd.n3318 vdd.n3317 52.4337
R3545 vdd.n3313 vdd.n3312 52.4337
R3546 vdd.n3310 vdd.n3309 52.4337
R3547 vdd.n3305 vdd.n3304 52.4337
R3548 vdd.n3302 vdd.n3301 52.4337
R3549 vdd.n3297 vdd.n3296 52.4337
R3550 vdd.n3292 vdd.n750 52.4337
R3551 vdd.n3288 vdd.n752 52.4337
R3552 vdd.n3524 vdd.n404 52.4337
R3553 vdd.n595 vdd.n403 52.4337
R3554 vdd.n589 vdd.n402 52.4337
R3555 vdd.n585 vdd.n401 52.4337
R3556 vdd.n579 vdd.n400 52.4337
R3557 vdd.n575 vdd.n399 52.4337
R3558 vdd.n569 vdd.n398 52.4337
R3559 vdd.n565 vdd.n397 52.4337
R3560 vdd.n559 vdd.n396 52.4337
R3561 vdd.n555 vdd.n395 52.4337
R3562 vdd.n549 vdd.n394 52.4337
R3563 vdd.n545 vdd.n393 52.4337
R3564 vdd.n539 vdd.n392 52.4337
R3565 vdd.n535 vdd.n391 52.4337
R3566 vdd.n529 vdd.n390 52.4337
R3567 vdd.n525 vdd.n389 52.4337
R3568 vdd.n519 vdd.n388 52.4337
R3569 vdd.n515 vdd.n387 52.4337
R3570 vdd.n509 vdd.n386 52.4337
R3571 vdd.n505 vdd.n385 52.4337
R3572 vdd.n499 vdd.n384 52.4337
R3573 vdd.n495 vdd.n383 52.4337
R3574 vdd.n489 vdd.n382 52.4337
R3575 vdd.n485 vdd.n381 52.4337
R3576 vdd.n479 vdd.n380 52.4337
R3577 vdd.n475 vdd.n379 52.4337
R3578 vdd.n469 vdd.n378 52.4337
R3579 vdd.n465 vdd.n377 52.4337
R3580 vdd.n459 vdd.n376 52.4337
R3581 vdd.n455 vdd.n375 52.4337
R3582 vdd.n449 vdd.n374 52.4337
R3583 vdd.n445 vdd.n373 52.4337
R3584 vdd.t209 vdd.t222 51.4683
R3585 vdd.n266 vdd.n264 42.0461
R3586 vdd.n168 vdd.n166 42.0461
R3587 vdd.n71 vdd.n69 42.0461
R3588 vdd.n2145 vdd.n2143 42.0461
R3589 vdd.n2047 vdd.n2045 42.0461
R3590 vdd.n1950 vdd.n1948 42.0461
R3591 vdd.n320 vdd.n319 41.6884
R3592 vdd.n222 vdd.n221 41.6884
R3593 vdd.n125 vdd.n124 41.6884
R3594 vdd.n2199 vdd.n2198 41.6884
R3595 vdd.n2101 vdd.n2100 41.6884
R3596 vdd.n2004 vdd.n2003 41.6884
R3597 vdd.n1605 vdd.n1604 41.1157
R3598 vdd.n1761 vdd.n1760 41.1157
R3599 vdd.n1797 vdd.n1796 41.1157
R3600 vdd.n407 vdd.n406 41.1157
R3601 vdd.n547 vdd.n420 41.1157
R3602 vdd.n433 vdd.n432 41.1157
R3603 vdd.n3242 vdd.n3241 39.2114
R3604 vdd.n3239 vdd.n3238 39.2114
R3605 vdd.n3234 vdd.n784 39.2114
R3606 vdd.n3232 vdd.n3231 39.2114
R3607 vdd.n3227 vdd.n787 39.2114
R3608 vdd.n3225 vdd.n3224 39.2114
R3609 vdd.n3220 vdd.n790 39.2114
R3610 vdd.n3218 vdd.n3217 39.2114
R3611 vdd.n3212 vdd.n793 39.2114
R3612 vdd.n3210 vdd.n3209 39.2114
R3613 vdd.n3205 vdd.n796 39.2114
R3614 vdd.n3203 vdd.n3202 39.2114
R3615 vdd.n3198 vdd.n799 39.2114
R3616 vdd.n3196 vdd.n3195 39.2114
R3617 vdd.n3191 vdd.n802 39.2114
R3618 vdd.n3189 vdd.n3188 39.2114
R3619 vdd.n3184 vdd.n3183 39.2114
R3620 vdd.n3007 vdd.n3006 39.2114
R3621 vdd.n2736 vdd.n2702 39.2114
R3622 vdd.n2999 vdd.n2703 39.2114
R3623 vdd.n2995 vdd.n2704 39.2114
R3624 vdd.n2991 vdd.n2705 39.2114
R3625 vdd.n2987 vdd.n2706 39.2114
R3626 vdd.n2983 vdd.n2707 39.2114
R3627 vdd.n2979 vdd.n2708 39.2114
R3628 vdd.n2975 vdd.n2709 39.2114
R3629 vdd.n2971 vdd.n2710 39.2114
R3630 vdd.n2967 vdd.n2711 39.2114
R3631 vdd.n2963 vdd.n2712 39.2114
R3632 vdd.n2959 vdd.n2713 39.2114
R3633 vdd.n2955 vdd.n2714 39.2114
R3634 vdd.n2951 vdd.n2715 39.2114
R3635 vdd.n2947 vdd.n2716 39.2114
R3636 vdd.n2942 vdd.n2717 39.2114
R3637 vdd.n2696 vdd.n968 39.2114
R3638 vdd.n2692 vdd.n967 39.2114
R3639 vdd.n2688 vdd.n966 39.2114
R3640 vdd.n2684 vdd.n965 39.2114
R3641 vdd.n2680 vdd.n964 39.2114
R3642 vdd.n2676 vdd.n963 39.2114
R3643 vdd.n2672 vdd.n962 39.2114
R3644 vdd.n2668 vdd.n961 39.2114
R3645 vdd.n2664 vdd.n960 39.2114
R3646 vdd.n2660 vdd.n959 39.2114
R3647 vdd.n2656 vdd.n958 39.2114
R3648 vdd.n2652 vdd.n957 39.2114
R3649 vdd.n2648 vdd.n956 39.2114
R3650 vdd.n2644 vdd.n955 39.2114
R3651 vdd.n2640 vdd.n954 39.2114
R3652 vdd.n2635 vdd.n953 39.2114
R3653 vdd.n2631 vdd.n952 39.2114
R3654 vdd.n2425 vdd.n2424 39.2114
R3655 vdd.n1147 vdd.n1113 39.2114
R3656 vdd.n2417 vdd.n1114 39.2114
R3657 vdd.n2413 vdd.n1115 39.2114
R3658 vdd.n2409 vdd.n1116 39.2114
R3659 vdd.n2405 vdd.n1117 39.2114
R3660 vdd.n2401 vdd.n1118 39.2114
R3661 vdd.n2397 vdd.n1119 39.2114
R3662 vdd.n2393 vdd.n1120 39.2114
R3663 vdd.n1293 vdd.n1121 39.2114
R3664 vdd.n1297 vdd.n1122 39.2114
R3665 vdd.n1301 vdd.n1123 39.2114
R3666 vdd.n1305 vdd.n1124 39.2114
R3667 vdd.n1309 vdd.n1125 39.2114
R3668 vdd.n1313 vdd.n1126 39.2114
R3669 vdd.n1317 vdd.n1127 39.2114
R3670 vdd.n1322 vdd.n1128 39.2114
R3671 vdd.n3161 vdd.n3160 39.2114
R3672 vdd.n3156 vdd.n3128 39.2114
R3673 vdd.n3154 vdd.n3153 39.2114
R3674 vdd.n3149 vdd.n3131 39.2114
R3675 vdd.n3147 vdd.n3146 39.2114
R3676 vdd.n3142 vdd.n3134 39.2114
R3677 vdd.n3140 vdd.n3139 39.2114
R3678 vdd.n3135 vdd.n755 39.2114
R3679 vdd.n3279 vdd.n3278 39.2114
R3680 vdd.n3276 vdd.n3275 39.2114
R3681 vdd.n3271 vdd.n760 39.2114
R3682 vdd.n3269 vdd.n3268 39.2114
R3683 vdd.n3264 vdd.n763 39.2114
R3684 vdd.n3262 vdd.n3261 39.2114
R3685 vdd.n3257 vdd.n766 39.2114
R3686 vdd.n3255 vdd.n3254 39.2114
R3687 vdd.n3250 vdd.n772 39.2114
R3688 vdd.n2743 vdd.n2718 39.2114
R3689 vdd.n2747 vdd.n2719 39.2114
R3690 vdd.n2751 vdd.n2720 39.2114
R3691 vdd.n2755 vdd.n2721 39.2114
R3692 vdd.n2759 vdd.n2722 39.2114
R3693 vdd.n2763 vdd.n2723 39.2114
R3694 vdd.n2767 vdd.n2724 39.2114
R3695 vdd.n2771 vdd.n2725 39.2114
R3696 vdd.n2775 vdd.n2726 39.2114
R3697 vdd.n2779 vdd.n2727 39.2114
R3698 vdd.n2783 vdd.n2728 39.2114
R3699 vdd.n2787 vdd.n2729 39.2114
R3700 vdd.n2791 vdd.n2730 39.2114
R3701 vdd.n2795 vdd.n2731 39.2114
R3702 vdd.n2799 vdd.n2732 39.2114
R3703 vdd.n2803 vdd.n2733 39.2114
R3704 vdd.n2807 vdd.n2734 39.2114
R3705 vdd.n2746 vdd.n2718 39.2114
R3706 vdd.n2750 vdd.n2719 39.2114
R3707 vdd.n2754 vdd.n2720 39.2114
R3708 vdd.n2758 vdd.n2721 39.2114
R3709 vdd.n2762 vdd.n2722 39.2114
R3710 vdd.n2766 vdd.n2723 39.2114
R3711 vdd.n2770 vdd.n2724 39.2114
R3712 vdd.n2774 vdd.n2725 39.2114
R3713 vdd.n2778 vdd.n2726 39.2114
R3714 vdd.n2782 vdd.n2727 39.2114
R3715 vdd.n2786 vdd.n2728 39.2114
R3716 vdd.n2790 vdd.n2729 39.2114
R3717 vdd.n2794 vdd.n2730 39.2114
R3718 vdd.n2798 vdd.n2731 39.2114
R3719 vdd.n2802 vdd.n2732 39.2114
R3720 vdd.n2806 vdd.n2733 39.2114
R3721 vdd.n2809 vdd.n2734 39.2114
R3722 vdd.n772 vdd.n767 39.2114
R3723 vdd.n3256 vdd.n3255 39.2114
R3724 vdd.n766 vdd.n764 39.2114
R3725 vdd.n3263 vdd.n3262 39.2114
R3726 vdd.n763 vdd.n761 39.2114
R3727 vdd.n3270 vdd.n3269 39.2114
R3728 vdd.n760 vdd.n758 39.2114
R3729 vdd.n3277 vdd.n3276 39.2114
R3730 vdd.n3280 vdd.n3279 39.2114
R3731 vdd.n3136 vdd.n3135 39.2114
R3732 vdd.n3141 vdd.n3140 39.2114
R3733 vdd.n3134 vdd.n3132 39.2114
R3734 vdd.n3148 vdd.n3147 39.2114
R3735 vdd.n3131 vdd.n3129 39.2114
R3736 vdd.n3155 vdd.n3154 39.2114
R3737 vdd.n3128 vdd.n3126 39.2114
R3738 vdd.n3162 vdd.n3161 39.2114
R3739 vdd.n2424 vdd.n1111 39.2114
R3740 vdd.n2418 vdd.n1113 39.2114
R3741 vdd.n2414 vdd.n1114 39.2114
R3742 vdd.n2410 vdd.n1115 39.2114
R3743 vdd.n2406 vdd.n1116 39.2114
R3744 vdd.n2402 vdd.n1117 39.2114
R3745 vdd.n2398 vdd.n1118 39.2114
R3746 vdd.n2394 vdd.n1119 39.2114
R3747 vdd.n1292 vdd.n1120 39.2114
R3748 vdd.n1296 vdd.n1121 39.2114
R3749 vdd.n1300 vdd.n1122 39.2114
R3750 vdd.n1304 vdd.n1123 39.2114
R3751 vdd.n1308 vdd.n1124 39.2114
R3752 vdd.n1312 vdd.n1125 39.2114
R3753 vdd.n1316 vdd.n1126 39.2114
R3754 vdd.n1321 vdd.n1127 39.2114
R3755 vdd.n1325 vdd.n1128 39.2114
R3756 vdd.n2634 vdd.n952 39.2114
R3757 vdd.n2639 vdd.n953 39.2114
R3758 vdd.n2643 vdd.n954 39.2114
R3759 vdd.n2647 vdd.n955 39.2114
R3760 vdd.n2651 vdd.n956 39.2114
R3761 vdd.n2655 vdd.n957 39.2114
R3762 vdd.n2659 vdd.n958 39.2114
R3763 vdd.n2663 vdd.n959 39.2114
R3764 vdd.n2667 vdd.n960 39.2114
R3765 vdd.n2671 vdd.n961 39.2114
R3766 vdd.n2675 vdd.n962 39.2114
R3767 vdd.n2679 vdd.n963 39.2114
R3768 vdd.n2683 vdd.n964 39.2114
R3769 vdd.n2687 vdd.n965 39.2114
R3770 vdd.n2691 vdd.n966 39.2114
R3771 vdd.n2695 vdd.n967 39.2114
R3772 vdd.n970 vdd.n968 39.2114
R3773 vdd.n3006 vdd.n933 39.2114
R3774 vdd.n3000 vdd.n2702 39.2114
R3775 vdd.n2996 vdd.n2703 39.2114
R3776 vdd.n2992 vdd.n2704 39.2114
R3777 vdd.n2988 vdd.n2705 39.2114
R3778 vdd.n2984 vdd.n2706 39.2114
R3779 vdd.n2980 vdd.n2707 39.2114
R3780 vdd.n2976 vdd.n2708 39.2114
R3781 vdd.n2972 vdd.n2709 39.2114
R3782 vdd.n2968 vdd.n2710 39.2114
R3783 vdd.n2964 vdd.n2711 39.2114
R3784 vdd.n2960 vdd.n2712 39.2114
R3785 vdd.n2956 vdd.n2713 39.2114
R3786 vdd.n2952 vdd.n2714 39.2114
R3787 vdd.n2948 vdd.n2715 39.2114
R3788 vdd.n2943 vdd.n2716 39.2114
R3789 vdd.n2939 vdd.n2717 39.2114
R3790 vdd.n3183 vdd.n803 39.2114
R3791 vdd.n3190 vdd.n3189 39.2114
R3792 vdd.n802 vdd.n800 39.2114
R3793 vdd.n3197 vdd.n3196 39.2114
R3794 vdd.n799 vdd.n797 39.2114
R3795 vdd.n3204 vdd.n3203 39.2114
R3796 vdd.n796 vdd.n794 39.2114
R3797 vdd.n3211 vdd.n3210 39.2114
R3798 vdd.n793 vdd.n791 39.2114
R3799 vdd.n3219 vdd.n3218 39.2114
R3800 vdd.n790 vdd.n788 39.2114
R3801 vdd.n3226 vdd.n3225 39.2114
R3802 vdd.n787 vdd.n785 39.2114
R3803 vdd.n3233 vdd.n3232 39.2114
R3804 vdd.n784 vdd.n782 39.2114
R3805 vdd.n3240 vdd.n3239 39.2114
R3806 vdd.n3243 vdd.n3242 39.2114
R3807 vdd.n979 vdd.n934 39.2114
R3808 vdd.n2623 vdd.n935 39.2114
R3809 vdd.n2619 vdd.n936 39.2114
R3810 vdd.n2615 vdd.n937 39.2114
R3811 vdd.n2611 vdd.n938 39.2114
R3812 vdd.n2607 vdd.n939 39.2114
R3813 vdd.n2603 vdd.n940 39.2114
R3814 vdd.n2599 vdd.n941 39.2114
R3815 vdd.n2595 vdd.n942 39.2114
R3816 vdd.n2591 vdd.n943 39.2114
R3817 vdd.n2587 vdd.n944 39.2114
R3818 vdd.n2583 vdd.n945 39.2114
R3819 vdd.n2579 vdd.n946 39.2114
R3820 vdd.n2575 vdd.n947 39.2114
R3821 vdd.n2571 vdd.n948 39.2114
R3822 vdd.n2567 vdd.n949 39.2114
R3823 vdd.n2563 vdd.n950 39.2114
R3824 vdd.n1251 vdd.n1129 39.2114
R3825 vdd.n1255 vdd.n1130 39.2114
R3826 vdd.n1259 vdd.n1131 39.2114
R3827 vdd.n1263 vdd.n1132 39.2114
R3828 vdd.n1267 vdd.n1133 39.2114
R3829 vdd.n1271 vdd.n1134 39.2114
R3830 vdd.n1275 vdd.n1135 39.2114
R3831 vdd.n1279 vdd.n1136 39.2114
R3832 vdd.n1283 vdd.n1137 39.2114
R3833 vdd.n1484 vdd.n1138 39.2114
R3834 vdd.n1481 vdd.n1139 39.2114
R3835 vdd.n1477 vdd.n1140 39.2114
R3836 vdd.n1473 vdd.n1141 39.2114
R3837 vdd.n1469 vdd.n1142 39.2114
R3838 vdd.n1465 vdd.n1143 39.2114
R3839 vdd.n1461 vdd.n1144 39.2114
R3840 vdd.n1457 vdd.n1145 39.2114
R3841 vdd.n2560 vdd.n950 39.2114
R3842 vdd.n2564 vdd.n949 39.2114
R3843 vdd.n2568 vdd.n948 39.2114
R3844 vdd.n2572 vdd.n947 39.2114
R3845 vdd.n2576 vdd.n946 39.2114
R3846 vdd.n2580 vdd.n945 39.2114
R3847 vdd.n2584 vdd.n944 39.2114
R3848 vdd.n2588 vdd.n943 39.2114
R3849 vdd.n2592 vdd.n942 39.2114
R3850 vdd.n2596 vdd.n941 39.2114
R3851 vdd.n2600 vdd.n940 39.2114
R3852 vdd.n2604 vdd.n939 39.2114
R3853 vdd.n2608 vdd.n938 39.2114
R3854 vdd.n2612 vdd.n937 39.2114
R3855 vdd.n2616 vdd.n936 39.2114
R3856 vdd.n2620 vdd.n935 39.2114
R3857 vdd.n2624 vdd.n934 39.2114
R3858 vdd.n1254 vdd.n1129 39.2114
R3859 vdd.n1258 vdd.n1130 39.2114
R3860 vdd.n1262 vdd.n1131 39.2114
R3861 vdd.n1266 vdd.n1132 39.2114
R3862 vdd.n1270 vdd.n1133 39.2114
R3863 vdd.n1274 vdd.n1134 39.2114
R3864 vdd.n1278 vdd.n1135 39.2114
R3865 vdd.n1282 vdd.n1136 39.2114
R3866 vdd.n1285 vdd.n1137 39.2114
R3867 vdd.n1482 vdd.n1138 39.2114
R3868 vdd.n1478 vdd.n1139 39.2114
R3869 vdd.n1474 vdd.n1140 39.2114
R3870 vdd.n1470 vdd.n1141 39.2114
R3871 vdd.n1466 vdd.n1142 39.2114
R3872 vdd.n1462 vdd.n1143 39.2114
R3873 vdd.n1458 vdd.n1144 39.2114
R3874 vdd.n1454 vdd.n1145 39.2114
R3875 vdd.n2281 vdd.n2280 37.2369
R3876 vdd.n2317 vdd.n1220 37.2369
R3877 vdd.n2356 vdd.n1180 37.2369
R3878 vdd.n3331 vdd.n724 37.2369
R3879 vdd.n688 vdd.n687 37.2369
R3880 vdd.n3287 vdd.n3286 37.2369
R3881 vdd.n1288 vdd.n1287 30.449
R3882 vdd.n983 vdd.n982 30.449
R3883 vdd.n1319 vdd.n1291 30.449
R3884 vdd.n2637 vdd.n973 30.449
R3885 vdd.n2742 vdd.n2741 30.449
R3886 vdd.n806 vdd.n805 30.449
R3887 vdd.n2945 vdd.n2738 30.449
R3888 vdd.n770 vdd.n769 30.449
R3889 vdd.n2427 vdd.n2426 29.8151
R3890 vdd.n2699 vdd.n971 29.8151
R3891 vdd.n2632 vdd.n974 29.8151
R3892 vdd.n1327 vdd.n1324 29.8151
R3893 vdd.n2940 vdd.n2937 29.8151
R3894 vdd.n3185 vdd.n3182 29.8151
R3895 vdd.n3009 vdd.n3008 29.8151
R3896 vdd.n3246 vdd.n3245 29.8151
R3897 vdd.n3165 vdd.n3164 29.8151
R3898 vdd.n3251 vdd.n771 29.8151
R3899 vdd.n2813 vdd.n2811 29.8151
R3900 vdd.n2744 vdd.n926 29.8151
R3901 vdd.n1252 vdd.n1103 29.8151
R3902 vdd.n2627 vdd.n2626 29.8151
R3903 vdd.n2559 vdd.n2558 29.8151
R3904 vdd.n1453 vdd.n1452 29.8151
R3905 vdd.n1835 vdd.n1601 19.3944
R3906 vdd.n1835 vdd.n1591 19.3944
R3907 vdd.n1847 vdd.n1591 19.3944
R3908 vdd.n1847 vdd.n1589 19.3944
R3909 vdd.n1851 vdd.n1589 19.3944
R3910 vdd.n1851 vdd.n1579 19.3944
R3911 vdd.n1864 vdd.n1579 19.3944
R3912 vdd.n1864 vdd.n1577 19.3944
R3913 vdd.n1868 vdd.n1577 19.3944
R3914 vdd.n1868 vdd.n1569 19.3944
R3915 vdd.n1881 vdd.n1569 19.3944
R3916 vdd.n1881 vdd.n1567 19.3944
R3917 vdd.n1885 vdd.n1567 19.3944
R3918 vdd.n1885 vdd.n1556 19.3944
R3919 vdd.n1897 vdd.n1556 19.3944
R3920 vdd.n1897 vdd.n1554 19.3944
R3921 vdd.n1901 vdd.n1554 19.3944
R3922 vdd.n1901 vdd.n1545 19.3944
R3923 vdd.n2209 vdd.n1545 19.3944
R3924 vdd.n2209 vdd.n1543 19.3944
R3925 vdd.n2213 vdd.n1543 19.3944
R3926 vdd.n2213 vdd.n1534 19.3944
R3927 vdd.n2225 vdd.n1534 19.3944
R3928 vdd.n2225 vdd.n1532 19.3944
R3929 vdd.n2229 vdd.n1532 19.3944
R3930 vdd.n2229 vdd.n1522 19.3944
R3931 vdd.n2242 vdd.n1522 19.3944
R3932 vdd.n2242 vdd.n1520 19.3944
R3933 vdd.n2246 vdd.n1520 19.3944
R3934 vdd.n2246 vdd.n1512 19.3944
R3935 vdd.n2259 vdd.n1512 19.3944
R3936 vdd.n2259 vdd.n1509 19.3944
R3937 vdd.n2265 vdd.n1509 19.3944
R3938 vdd.n2265 vdd.n1510 19.3944
R3939 vdd.n1510 vdd.n1499 19.3944
R3940 vdd.n1754 vdd.n1696 19.3944
R3941 vdd.n1754 vdd.n1753 19.3944
R3942 vdd.n1753 vdd.n1752 19.3944
R3943 vdd.n1752 vdd.n1702 19.3944
R3944 vdd.n1748 vdd.n1702 19.3944
R3945 vdd.n1748 vdd.n1747 19.3944
R3946 vdd.n1747 vdd.n1746 19.3944
R3947 vdd.n1746 vdd.n1708 19.3944
R3948 vdd.n1742 vdd.n1708 19.3944
R3949 vdd.n1742 vdd.n1741 19.3944
R3950 vdd.n1741 vdd.n1740 19.3944
R3951 vdd.n1740 vdd.n1714 19.3944
R3952 vdd.n1736 vdd.n1714 19.3944
R3953 vdd.n1736 vdd.n1735 19.3944
R3954 vdd.n1735 vdd.n1734 19.3944
R3955 vdd.n1734 vdd.n1720 19.3944
R3956 vdd.n1730 vdd.n1720 19.3944
R3957 vdd.n1730 vdd.n1729 19.3944
R3958 vdd.n1729 vdd.n1728 19.3944
R3959 vdd.n1728 vdd.n1726 19.3944
R3960 vdd.n1792 vdd.n1791 19.3944
R3961 vdd.n1791 vdd.n1667 19.3944
R3962 vdd.n1787 vdd.n1667 19.3944
R3963 vdd.n1787 vdd.n1786 19.3944
R3964 vdd.n1786 vdd.n1785 19.3944
R3965 vdd.n1785 vdd.n1673 19.3944
R3966 vdd.n1781 vdd.n1673 19.3944
R3967 vdd.n1781 vdd.n1780 19.3944
R3968 vdd.n1780 vdd.n1779 19.3944
R3969 vdd.n1779 vdd.n1679 19.3944
R3970 vdd.n1775 vdd.n1679 19.3944
R3971 vdd.n1775 vdd.n1774 19.3944
R3972 vdd.n1774 vdd.n1773 19.3944
R3973 vdd.n1773 vdd.n1685 19.3944
R3974 vdd.n1769 vdd.n1685 19.3944
R3975 vdd.n1769 vdd.n1768 19.3944
R3976 vdd.n1768 vdd.n1767 19.3944
R3977 vdd.n1767 vdd.n1691 19.3944
R3978 vdd.n1763 vdd.n1691 19.3944
R3979 vdd.n1763 vdd.n1762 19.3944
R3980 vdd.n1826 vdd.n1825 19.3944
R3981 vdd.n1825 vdd.n1640 19.3944
R3982 vdd.n1821 vdd.n1640 19.3944
R3983 vdd.n1821 vdd.n1820 19.3944
R3984 vdd.n1820 vdd.n1819 19.3944
R3985 vdd.n1819 vdd.n1645 19.3944
R3986 vdd.n1815 vdd.n1645 19.3944
R3987 vdd.n1815 vdd.n1814 19.3944
R3988 vdd.n1814 vdd.n1813 19.3944
R3989 vdd.n1813 vdd.n1651 19.3944
R3990 vdd.n1809 vdd.n1651 19.3944
R3991 vdd.n1809 vdd.n1808 19.3944
R3992 vdd.n1808 vdd.n1807 19.3944
R3993 vdd.n1807 vdd.n1657 19.3944
R3994 vdd.n1803 vdd.n1657 19.3944
R3995 vdd.n1803 vdd.n1802 19.3944
R3996 vdd.n1802 vdd.n1801 19.3944
R3997 vdd.n1801 vdd.n1663 19.3944
R3998 vdd.n2313 vdd.n1218 19.3944
R3999 vdd.n2313 vdd.n1224 19.3944
R4000 vdd.n2308 vdd.n1224 19.3944
R4001 vdd.n2308 vdd.n2307 19.3944
R4002 vdd.n2307 vdd.n2306 19.3944
R4003 vdd.n2306 vdd.n1231 19.3944
R4004 vdd.n2301 vdd.n1231 19.3944
R4005 vdd.n2301 vdd.n2300 19.3944
R4006 vdd.n2300 vdd.n2299 19.3944
R4007 vdd.n2299 vdd.n1238 19.3944
R4008 vdd.n2294 vdd.n1238 19.3944
R4009 vdd.n2294 vdd.n2293 19.3944
R4010 vdd.n2293 vdd.n2292 19.3944
R4011 vdd.n2292 vdd.n1245 19.3944
R4012 vdd.n2287 vdd.n1245 19.3944
R4013 vdd.n2287 vdd.n2286 19.3944
R4014 vdd.n1492 vdd.n1250 19.3944
R4015 vdd.n2282 vdd.n1489 19.3944
R4016 vdd.n2352 vdd.n1178 19.3944
R4017 vdd.n2352 vdd.n1184 19.3944
R4018 vdd.n2347 vdd.n1184 19.3944
R4019 vdd.n2347 vdd.n2346 19.3944
R4020 vdd.n2346 vdd.n2345 19.3944
R4021 vdd.n2345 vdd.n1191 19.3944
R4022 vdd.n2340 vdd.n1191 19.3944
R4023 vdd.n2340 vdd.n2339 19.3944
R4024 vdd.n2339 vdd.n2338 19.3944
R4025 vdd.n2338 vdd.n1198 19.3944
R4026 vdd.n2333 vdd.n1198 19.3944
R4027 vdd.n2333 vdd.n2332 19.3944
R4028 vdd.n2332 vdd.n2331 19.3944
R4029 vdd.n2331 vdd.n1205 19.3944
R4030 vdd.n2326 vdd.n1205 19.3944
R4031 vdd.n2326 vdd.n2325 19.3944
R4032 vdd.n2325 vdd.n2324 19.3944
R4033 vdd.n2324 vdd.n1212 19.3944
R4034 vdd.n2319 vdd.n1212 19.3944
R4035 vdd.n2319 vdd.n2318 19.3944
R4036 vdd.n2389 vdd.n1153 19.3944
R4037 vdd.n2389 vdd.n1154 19.3944
R4038 vdd.n2384 vdd.n2383 19.3944
R4039 vdd.n2379 vdd.n2378 19.3944
R4040 vdd.n2378 vdd.n2377 19.3944
R4041 vdd.n2377 vdd.n1158 19.3944
R4042 vdd.n2372 vdd.n1158 19.3944
R4043 vdd.n2372 vdd.n2371 19.3944
R4044 vdd.n2371 vdd.n2370 19.3944
R4045 vdd.n2370 vdd.n1165 19.3944
R4046 vdd.n2365 vdd.n1165 19.3944
R4047 vdd.n2365 vdd.n2364 19.3944
R4048 vdd.n2364 vdd.n2363 19.3944
R4049 vdd.n2363 vdd.n1172 19.3944
R4050 vdd.n2358 vdd.n1172 19.3944
R4051 vdd.n2358 vdd.n2357 19.3944
R4052 vdd.n1839 vdd.n1597 19.3944
R4053 vdd.n1839 vdd.n1595 19.3944
R4054 vdd.n1843 vdd.n1595 19.3944
R4055 vdd.n1843 vdd.n1585 19.3944
R4056 vdd.n1856 vdd.n1585 19.3944
R4057 vdd.n1856 vdd.n1583 19.3944
R4058 vdd.n1860 vdd.n1583 19.3944
R4059 vdd.n1860 vdd.n1574 19.3944
R4060 vdd.n1873 vdd.n1574 19.3944
R4061 vdd.n1873 vdd.n1572 19.3944
R4062 vdd.n1877 vdd.n1572 19.3944
R4063 vdd.n1877 vdd.n1563 19.3944
R4064 vdd.n1889 vdd.n1563 19.3944
R4065 vdd.n1889 vdd.n1561 19.3944
R4066 vdd.n1893 vdd.n1561 19.3944
R4067 vdd.n1893 vdd.n1551 19.3944
R4068 vdd.n1906 vdd.n1551 19.3944
R4069 vdd.n1906 vdd.n1549 19.3944
R4070 vdd.n2205 vdd.n1549 19.3944
R4071 vdd.n2205 vdd.n1540 19.3944
R4072 vdd.n2217 vdd.n1540 19.3944
R4073 vdd.n2217 vdd.n1538 19.3944
R4074 vdd.n2221 vdd.n1538 19.3944
R4075 vdd.n2221 vdd.n1528 19.3944
R4076 vdd.n2234 vdd.n1528 19.3944
R4077 vdd.n2234 vdd.n1526 19.3944
R4078 vdd.n2238 vdd.n1526 19.3944
R4079 vdd.n2238 vdd.n1517 19.3944
R4080 vdd.n2251 vdd.n1517 19.3944
R4081 vdd.n2251 vdd.n1515 19.3944
R4082 vdd.n2255 vdd.n1515 19.3944
R4083 vdd.n2255 vdd.n1505 19.3944
R4084 vdd.n2269 vdd.n1505 19.3944
R4085 vdd.n2269 vdd.n1503 19.3944
R4086 vdd.n2273 vdd.n1503 19.3944
R4087 vdd.n3419 vdd.n655 19.3944
R4088 vdd.n3423 vdd.n655 19.3944
R4089 vdd.n3423 vdd.n646 19.3944
R4090 vdd.n3435 vdd.n646 19.3944
R4091 vdd.n3435 vdd.n644 19.3944
R4092 vdd.n3439 vdd.n644 19.3944
R4093 vdd.n3439 vdd.n633 19.3944
R4094 vdd.n3451 vdd.n633 19.3944
R4095 vdd.n3451 vdd.n631 19.3944
R4096 vdd.n3455 vdd.n631 19.3944
R4097 vdd.n3455 vdd.n622 19.3944
R4098 vdd.n3468 vdd.n622 19.3944
R4099 vdd.n3468 vdd.n620 19.3944
R4100 vdd.n3475 vdd.n620 19.3944
R4101 vdd.n3475 vdd.n3474 19.3944
R4102 vdd.n3474 vdd.n610 19.3944
R4103 vdd.n3488 vdd.n610 19.3944
R4104 vdd.n3489 vdd.n3488 19.3944
R4105 vdd.n3490 vdd.n3489 19.3944
R4106 vdd.n3490 vdd.n608 19.3944
R4107 vdd.n3495 vdd.n608 19.3944
R4108 vdd.n3496 vdd.n3495 19.3944
R4109 vdd.n3497 vdd.n3496 19.3944
R4110 vdd.n3497 vdd.n606 19.3944
R4111 vdd.n3502 vdd.n606 19.3944
R4112 vdd.n3503 vdd.n3502 19.3944
R4113 vdd.n3504 vdd.n3503 19.3944
R4114 vdd.n3504 vdd.n604 19.3944
R4115 vdd.n3510 vdd.n604 19.3944
R4116 vdd.n3511 vdd.n3510 19.3944
R4117 vdd.n3512 vdd.n3511 19.3944
R4118 vdd.n3512 vdd.n602 19.3944
R4119 vdd.n3517 vdd.n602 19.3944
R4120 vdd.n3518 vdd.n3517 19.3944
R4121 vdd.n3519 vdd.n3518 19.3944
R4122 vdd.n550 vdd.n417 19.3944
R4123 vdd.n556 vdd.n417 19.3944
R4124 vdd.n557 vdd.n556 19.3944
R4125 vdd.n560 vdd.n557 19.3944
R4126 vdd.n560 vdd.n415 19.3944
R4127 vdd.n566 vdd.n415 19.3944
R4128 vdd.n567 vdd.n566 19.3944
R4129 vdd.n570 vdd.n567 19.3944
R4130 vdd.n570 vdd.n413 19.3944
R4131 vdd.n576 vdd.n413 19.3944
R4132 vdd.n577 vdd.n576 19.3944
R4133 vdd.n580 vdd.n577 19.3944
R4134 vdd.n580 vdd.n411 19.3944
R4135 vdd.n586 vdd.n411 19.3944
R4136 vdd.n587 vdd.n586 19.3944
R4137 vdd.n590 vdd.n587 19.3944
R4138 vdd.n590 vdd.n409 19.3944
R4139 vdd.n596 vdd.n409 19.3944
R4140 vdd.n598 vdd.n596 19.3944
R4141 vdd.n599 vdd.n598 19.3944
R4142 vdd.n497 vdd.n496 19.3944
R4143 vdd.n500 vdd.n497 19.3944
R4144 vdd.n500 vdd.n429 19.3944
R4145 vdd.n506 vdd.n429 19.3944
R4146 vdd.n507 vdd.n506 19.3944
R4147 vdd.n510 vdd.n507 19.3944
R4148 vdd.n510 vdd.n427 19.3944
R4149 vdd.n516 vdd.n427 19.3944
R4150 vdd.n517 vdd.n516 19.3944
R4151 vdd.n520 vdd.n517 19.3944
R4152 vdd.n520 vdd.n425 19.3944
R4153 vdd.n526 vdd.n425 19.3944
R4154 vdd.n527 vdd.n526 19.3944
R4155 vdd.n530 vdd.n527 19.3944
R4156 vdd.n530 vdd.n423 19.3944
R4157 vdd.n536 vdd.n423 19.3944
R4158 vdd.n537 vdd.n536 19.3944
R4159 vdd.n540 vdd.n537 19.3944
R4160 vdd.n540 vdd.n421 19.3944
R4161 vdd.n546 vdd.n421 19.3944
R4162 vdd.n447 vdd.n446 19.3944
R4163 vdd.n450 vdd.n447 19.3944
R4164 vdd.n450 vdd.n441 19.3944
R4165 vdd.n456 vdd.n441 19.3944
R4166 vdd.n457 vdd.n456 19.3944
R4167 vdd.n460 vdd.n457 19.3944
R4168 vdd.n460 vdd.n439 19.3944
R4169 vdd.n466 vdd.n439 19.3944
R4170 vdd.n467 vdd.n466 19.3944
R4171 vdd.n470 vdd.n467 19.3944
R4172 vdd.n470 vdd.n437 19.3944
R4173 vdd.n476 vdd.n437 19.3944
R4174 vdd.n477 vdd.n476 19.3944
R4175 vdd.n480 vdd.n477 19.3944
R4176 vdd.n480 vdd.n435 19.3944
R4177 vdd.n486 vdd.n435 19.3944
R4178 vdd.n487 vdd.n486 19.3944
R4179 vdd.n490 vdd.n487 19.3944
R4180 vdd.n3415 vdd.n652 19.3944
R4181 vdd.n3427 vdd.n652 19.3944
R4182 vdd.n3427 vdd.n650 19.3944
R4183 vdd.n3431 vdd.n650 19.3944
R4184 vdd.n3431 vdd.n640 19.3944
R4185 vdd.n3443 vdd.n640 19.3944
R4186 vdd.n3443 vdd.n638 19.3944
R4187 vdd.n3447 vdd.n638 19.3944
R4188 vdd.n3447 vdd.n628 19.3944
R4189 vdd.n3460 vdd.n628 19.3944
R4190 vdd.n3460 vdd.n626 19.3944
R4191 vdd.n3464 vdd.n626 19.3944
R4192 vdd.n3464 vdd.n617 19.3944
R4193 vdd.n3479 vdd.n617 19.3944
R4194 vdd.n3479 vdd.n615 19.3944
R4195 vdd.n3483 vdd.n615 19.3944
R4196 vdd.n3483 vdd.n324 19.3944
R4197 vdd.n3561 vdd.n324 19.3944
R4198 vdd.n3561 vdd.n325 19.3944
R4199 vdd.n3555 vdd.n325 19.3944
R4200 vdd.n3555 vdd.n3554 19.3944
R4201 vdd.n3554 vdd.n3553 19.3944
R4202 vdd.n3553 vdd.n337 19.3944
R4203 vdd.n3547 vdd.n337 19.3944
R4204 vdd.n3547 vdd.n3546 19.3944
R4205 vdd.n3546 vdd.n3545 19.3944
R4206 vdd.n3545 vdd.n347 19.3944
R4207 vdd.n3539 vdd.n347 19.3944
R4208 vdd.n3539 vdd.n3538 19.3944
R4209 vdd.n3538 vdd.n3537 19.3944
R4210 vdd.n3537 vdd.n358 19.3944
R4211 vdd.n3531 vdd.n358 19.3944
R4212 vdd.n3531 vdd.n3530 19.3944
R4213 vdd.n3530 vdd.n3529 19.3944
R4214 vdd.n3529 vdd.n369 19.3944
R4215 vdd.n3372 vdd.n3371 19.3944
R4216 vdd.n3371 vdd.n3370 19.3944
R4217 vdd.n3370 vdd.n694 19.3944
R4218 vdd.n3364 vdd.n694 19.3944
R4219 vdd.n3364 vdd.n3363 19.3944
R4220 vdd.n3363 vdd.n3362 19.3944
R4221 vdd.n3362 vdd.n700 19.3944
R4222 vdd.n3356 vdd.n700 19.3944
R4223 vdd.n3356 vdd.n3355 19.3944
R4224 vdd.n3355 vdd.n3354 19.3944
R4225 vdd.n3354 vdd.n706 19.3944
R4226 vdd.n3348 vdd.n706 19.3944
R4227 vdd.n3348 vdd.n3347 19.3944
R4228 vdd.n3347 vdd.n3346 19.3944
R4229 vdd.n3346 vdd.n712 19.3944
R4230 vdd.n3340 vdd.n712 19.3944
R4231 vdd.n3340 vdd.n3339 19.3944
R4232 vdd.n3339 vdd.n3338 19.3944
R4233 vdd.n3338 vdd.n718 19.3944
R4234 vdd.n3332 vdd.n718 19.3944
R4235 vdd.n3412 vdd.n3411 19.3944
R4236 vdd.n3411 vdd.n662 19.3944
R4237 vdd.n3406 vdd.n3405 19.3944
R4238 vdd.n3402 vdd.n3401 19.3944
R4239 vdd.n3401 vdd.n668 19.3944
R4240 vdd.n3396 vdd.n668 19.3944
R4241 vdd.n3396 vdd.n3395 19.3944
R4242 vdd.n3395 vdd.n3394 19.3944
R4243 vdd.n3394 vdd.n674 19.3944
R4244 vdd.n3388 vdd.n674 19.3944
R4245 vdd.n3388 vdd.n3387 19.3944
R4246 vdd.n3387 vdd.n3386 19.3944
R4247 vdd.n3386 vdd.n680 19.3944
R4248 vdd.n3380 vdd.n680 19.3944
R4249 vdd.n3380 vdd.n3379 19.3944
R4250 vdd.n3379 vdd.n3378 19.3944
R4251 vdd.n3327 vdd.n722 19.3944
R4252 vdd.n3327 vdd.n726 19.3944
R4253 vdd.n3322 vdd.n726 19.3944
R4254 vdd.n3322 vdd.n3321 19.3944
R4255 vdd.n3321 vdd.n732 19.3944
R4256 vdd.n3316 vdd.n732 19.3944
R4257 vdd.n3316 vdd.n3315 19.3944
R4258 vdd.n3315 vdd.n3314 19.3944
R4259 vdd.n3314 vdd.n738 19.3944
R4260 vdd.n3308 vdd.n738 19.3944
R4261 vdd.n3308 vdd.n3307 19.3944
R4262 vdd.n3307 vdd.n3306 19.3944
R4263 vdd.n3306 vdd.n744 19.3944
R4264 vdd.n3300 vdd.n744 19.3944
R4265 vdd.n3300 vdd.n3299 19.3944
R4266 vdd.n3299 vdd.n3298 19.3944
R4267 vdd.n3294 vdd.n3293 19.3944
R4268 vdd.n3290 vdd.n3289 19.3944
R4269 vdd.n1761 vdd.n1696 19.0066
R4270 vdd.n2317 vdd.n1218 19.0066
R4271 vdd.n550 vdd.n547 19.0066
R4272 vdd.n3331 vdd.n722 19.0066
R4273 vdd.n1829 vdd.n1599 18.5924
R4274 vdd.n2275 vdd.n1112 18.5924
R4275 vdd.n3417 vdd.n658 18.5924
R4276 vdd.n3526 vdd.n3525 18.5924
R4277 vdd.n1287 vdd.n1286 16.0975
R4278 vdd.n982 vdd.n981 16.0975
R4279 vdd.n1604 vdd.n1603 16.0975
R4280 vdd.n1760 vdd.n1759 16.0975
R4281 vdd.n1796 vdd.n1795 16.0975
R4282 vdd.n2280 vdd.n2279 16.0975
R4283 vdd.n1220 vdd.n1219 16.0975
R4284 vdd.n1180 vdd.n1179 16.0975
R4285 vdd.n1291 vdd.n1290 16.0975
R4286 vdd.n973 vdd.n972 16.0975
R4287 vdd.n2741 vdd.n2740 16.0975
R4288 vdd.n406 vdd.n405 16.0975
R4289 vdd.n420 vdd.n419 16.0975
R4290 vdd.n432 vdd.n431 16.0975
R4291 vdd.n724 vdd.n723 16.0975
R4292 vdd.n687 vdd.n686 16.0975
R4293 vdd.n805 vdd.n804 16.0975
R4294 vdd.n2738 vdd.n2737 16.0975
R4295 vdd.n3286 vdd.n3285 16.0975
R4296 vdd.n769 vdd.n768 16.0975
R4297 vdd.t222 vdd.n2701 15.4182
R4298 vdd.n3005 vdd.t209 15.4182
R4299 vdd.n28 vdd.n27 14.7341
R4300 vdd.n316 vdd.n281 13.1884
R4301 vdd.n261 vdd.n226 13.1884
R4302 vdd.n218 vdd.n183 13.1884
R4303 vdd.n163 vdd.n128 13.1884
R4304 vdd.n121 vdd.n86 13.1884
R4305 vdd.n66 vdd.n31 13.1884
R4306 vdd.n2140 vdd.n2105 13.1884
R4307 vdd.n2195 vdd.n2160 13.1884
R4308 vdd.n2042 vdd.n2007 13.1884
R4309 vdd.n2097 vdd.n2062 13.1884
R4310 vdd.n1945 vdd.n1910 13.1884
R4311 vdd.n2000 vdd.n1965 13.1884
R4312 vdd.n2423 vdd.n1105 13.1509
R4313 vdd.n3248 vdd.n756 13.1509
R4314 vdd.n1797 vdd.n1792 12.9944
R4315 vdd.n1797 vdd.n1663 12.9944
R4316 vdd.n2356 vdd.n1178 12.9944
R4317 vdd.n2357 vdd.n2356 12.9944
R4318 vdd.n496 vdd.n433 12.9944
R4319 vdd.n490 vdd.n433 12.9944
R4320 vdd.n3372 vdd.n688 12.9944
R4321 vdd.n3378 vdd.n688 12.9944
R4322 vdd.n317 vdd.n279 12.8005
R4323 vdd.n312 vdd.n283 12.8005
R4324 vdd.n262 vdd.n224 12.8005
R4325 vdd.n257 vdd.n228 12.8005
R4326 vdd.n219 vdd.n181 12.8005
R4327 vdd.n214 vdd.n185 12.8005
R4328 vdd.n164 vdd.n126 12.8005
R4329 vdd.n159 vdd.n130 12.8005
R4330 vdd.n122 vdd.n84 12.8005
R4331 vdd.n117 vdd.n88 12.8005
R4332 vdd.n67 vdd.n29 12.8005
R4333 vdd.n62 vdd.n33 12.8005
R4334 vdd.n2141 vdd.n2103 12.8005
R4335 vdd.n2136 vdd.n2107 12.8005
R4336 vdd.n2196 vdd.n2158 12.8005
R4337 vdd.n2191 vdd.n2162 12.8005
R4338 vdd.n2043 vdd.n2005 12.8005
R4339 vdd.n2038 vdd.n2009 12.8005
R4340 vdd.n2098 vdd.n2060 12.8005
R4341 vdd.n2093 vdd.n2064 12.8005
R4342 vdd.n1946 vdd.n1908 12.8005
R4343 vdd.n1941 vdd.n1912 12.8005
R4344 vdd.n2001 vdd.n1963 12.8005
R4345 vdd.n1996 vdd.n1967 12.8005
R4346 vdd.n311 vdd.n284 12.0247
R4347 vdd.n256 vdd.n229 12.0247
R4348 vdd.n213 vdd.n186 12.0247
R4349 vdd.n158 vdd.n131 12.0247
R4350 vdd.n116 vdd.n89 12.0247
R4351 vdd.n61 vdd.n34 12.0247
R4352 vdd.n2135 vdd.n2108 12.0247
R4353 vdd.n2190 vdd.n2163 12.0247
R4354 vdd.n2037 vdd.n2010 12.0247
R4355 vdd.n2092 vdd.n2065 12.0247
R4356 vdd.n1940 vdd.n1913 12.0247
R4357 vdd.n1995 vdd.n1968 12.0247
R4358 vdd.n1837 vdd.n1599 11.337
R4359 vdd.n1845 vdd.n1593 11.337
R4360 vdd.n1845 vdd.n1587 11.337
R4361 vdd.n1854 vdd.n1587 11.337
R4362 vdd.n1862 vdd.n1581 11.337
R4363 vdd.n1871 vdd.n1870 11.337
R4364 vdd.n1887 vdd.n1565 11.337
R4365 vdd.n1895 vdd.n1558 11.337
R4366 vdd.n1904 vdd.n1903 11.337
R4367 vdd.n2207 vdd.n1547 11.337
R4368 vdd.n2223 vdd.n1536 11.337
R4369 vdd.n2232 vdd.n1530 11.337
R4370 vdd.n2240 vdd.n1524 11.337
R4371 vdd.n2249 vdd.n2248 11.337
R4372 vdd.n2257 vdd.n1507 11.337
R4373 vdd.n2267 vdd.n1507 11.337
R4374 vdd.n2275 vdd.n1500 11.337
R4375 vdd.n3417 vdd.n659 11.337
R4376 vdd.n3425 vdd.n648 11.337
R4377 vdd.n3433 vdd.n648 11.337
R4378 vdd.n3441 vdd.n642 11.337
R4379 vdd.n3449 vdd.n635 11.337
R4380 vdd.n3458 vdd.n3457 11.337
R4381 vdd.n3466 vdd.n624 11.337
R4382 vdd.n3485 vdd.n613 11.337
R4383 vdd.n3559 vdd.n328 11.337
R4384 vdd.n3557 vdd.n332 11.337
R4385 vdd.n3551 vdd.n3550 11.337
R4386 vdd.n3543 vdd.n349 11.337
R4387 vdd.n3542 vdd.n3541 11.337
R4388 vdd.n3535 vdd.n3534 11.337
R4389 vdd.n3534 vdd.n3533 11.337
R4390 vdd.n3533 vdd.n363 11.337
R4391 vdd.n3527 vdd.n3526 11.337
R4392 vdd.n308 vdd.n307 11.249
R4393 vdd.n253 vdd.n252 11.249
R4394 vdd.n210 vdd.n209 11.249
R4395 vdd.n155 vdd.n154 11.249
R4396 vdd.n113 vdd.n112 11.249
R4397 vdd.n58 vdd.n57 11.249
R4398 vdd.n2132 vdd.n2131 11.249
R4399 vdd.n2187 vdd.n2186 11.249
R4400 vdd.n2034 vdd.n2033 11.249
R4401 vdd.n2089 vdd.n2088 11.249
R4402 vdd.n1937 vdd.n1936 11.249
R4403 vdd.n1992 vdd.n1991 11.249
R4404 vdd.n2257 vdd.t165 10.7702
R4405 vdd.n3433 vdd.t51 10.7702
R4406 vdd.n293 vdd.n292 10.7238
R4407 vdd.n238 vdd.n237 10.7238
R4408 vdd.n195 vdd.n194 10.7238
R4409 vdd.n140 vdd.n139 10.7238
R4410 vdd.n98 vdd.n97 10.7238
R4411 vdd.n43 vdd.n42 10.7238
R4412 vdd.n2117 vdd.n2116 10.7238
R4413 vdd.n2172 vdd.n2171 10.7238
R4414 vdd.n2019 vdd.n2018 10.7238
R4415 vdd.n2074 vdd.n2073 10.7238
R4416 vdd.n1922 vdd.n1921 10.7238
R4417 vdd.n1977 vdd.n1976 10.7238
R4418 vdd.n2428 vdd.n2427 10.6151
R4419 vdd.n2428 vdd.n1098 10.6151
R4420 vdd.n2438 vdd.n1098 10.6151
R4421 vdd.n2439 vdd.n2438 10.6151
R4422 vdd.n2440 vdd.n2439 10.6151
R4423 vdd.n2440 vdd.n1085 10.6151
R4424 vdd.n2450 vdd.n1085 10.6151
R4425 vdd.n2451 vdd.n2450 10.6151
R4426 vdd.n2452 vdd.n2451 10.6151
R4427 vdd.n2452 vdd.n1073 10.6151
R4428 vdd.n2462 vdd.n1073 10.6151
R4429 vdd.n2463 vdd.n2462 10.6151
R4430 vdd.n2464 vdd.n2463 10.6151
R4431 vdd.n2464 vdd.n1062 10.6151
R4432 vdd.n2474 vdd.n1062 10.6151
R4433 vdd.n2475 vdd.n2474 10.6151
R4434 vdd.n2476 vdd.n2475 10.6151
R4435 vdd.n2476 vdd.n1049 10.6151
R4436 vdd.n2486 vdd.n1049 10.6151
R4437 vdd.n2487 vdd.n2486 10.6151
R4438 vdd.n2488 vdd.n2487 10.6151
R4439 vdd.n2488 vdd.n1037 10.6151
R4440 vdd.n2499 vdd.n1037 10.6151
R4441 vdd.n2500 vdd.n2499 10.6151
R4442 vdd.n2501 vdd.n2500 10.6151
R4443 vdd.n2501 vdd.n1025 10.6151
R4444 vdd.n2511 vdd.n1025 10.6151
R4445 vdd.n2512 vdd.n2511 10.6151
R4446 vdd.n2513 vdd.n2512 10.6151
R4447 vdd.n2513 vdd.n1013 10.6151
R4448 vdd.n2523 vdd.n1013 10.6151
R4449 vdd.n2524 vdd.n2523 10.6151
R4450 vdd.n2525 vdd.n2524 10.6151
R4451 vdd.n2525 vdd.n1003 10.6151
R4452 vdd.n2535 vdd.n1003 10.6151
R4453 vdd.n2536 vdd.n2535 10.6151
R4454 vdd.n2537 vdd.n2536 10.6151
R4455 vdd.n2537 vdd.n990 10.6151
R4456 vdd.n2549 vdd.n990 10.6151
R4457 vdd.n2550 vdd.n2549 10.6151
R4458 vdd.n2552 vdd.n2550 10.6151
R4459 vdd.n2552 vdd.n2551 10.6151
R4460 vdd.n2551 vdd.n971 10.6151
R4461 vdd.n2699 vdd.n2698 10.6151
R4462 vdd.n2698 vdd.n2697 10.6151
R4463 vdd.n2697 vdd.n2694 10.6151
R4464 vdd.n2694 vdd.n2693 10.6151
R4465 vdd.n2693 vdd.n2690 10.6151
R4466 vdd.n2690 vdd.n2689 10.6151
R4467 vdd.n2689 vdd.n2686 10.6151
R4468 vdd.n2686 vdd.n2685 10.6151
R4469 vdd.n2685 vdd.n2682 10.6151
R4470 vdd.n2682 vdd.n2681 10.6151
R4471 vdd.n2681 vdd.n2678 10.6151
R4472 vdd.n2678 vdd.n2677 10.6151
R4473 vdd.n2677 vdd.n2674 10.6151
R4474 vdd.n2674 vdd.n2673 10.6151
R4475 vdd.n2673 vdd.n2670 10.6151
R4476 vdd.n2670 vdd.n2669 10.6151
R4477 vdd.n2669 vdd.n2666 10.6151
R4478 vdd.n2666 vdd.n2665 10.6151
R4479 vdd.n2665 vdd.n2662 10.6151
R4480 vdd.n2662 vdd.n2661 10.6151
R4481 vdd.n2661 vdd.n2658 10.6151
R4482 vdd.n2658 vdd.n2657 10.6151
R4483 vdd.n2657 vdd.n2654 10.6151
R4484 vdd.n2654 vdd.n2653 10.6151
R4485 vdd.n2653 vdd.n2650 10.6151
R4486 vdd.n2650 vdd.n2649 10.6151
R4487 vdd.n2649 vdd.n2646 10.6151
R4488 vdd.n2646 vdd.n2645 10.6151
R4489 vdd.n2645 vdd.n2642 10.6151
R4490 vdd.n2642 vdd.n2641 10.6151
R4491 vdd.n2641 vdd.n2638 10.6151
R4492 vdd.n2636 vdd.n2633 10.6151
R4493 vdd.n2633 vdd.n2632 10.6151
R4494 vdd.n1328 vdd.n1327 10.6151
R4495 vdd.n1330 vdd.n1328 10.6151
R4496 vdd.n1331 vdd.n1330 10.6151
R4497 vdd.n1333 vdd.n1331 10.6151
R4498 vdd.n1334 vdd.n1333 10.6151
R4499 vdd.n1336 vdd.n1334 10.6151
R4500 vdd.n1337 vdd.n1336 10.6151
R4501 vdd.n1339 vdd.n1337 10.6151
R4502 vdd.n1340 vdd.n1339 10.6151
R4503 vdd.n1342 vdd.n1340 10.6151
R4504 vdd.n1343 vdd.n1342 10.6151
R4505 vdd.n1345 vdd.n1343 10.6151
R4506 vdd.n1346 vdd.n1345 10.6151
R4507 vdd.n1348 vdd.n1346 10.6151
R4508 vdd.n1349 vdd.n1348 10.6151
R4509 vdd.n1351 vdd.n1349 10.6151
R4510 vdd.n1352 vdd.n1351 10.6151
R4511 vdd.n1354 vdd.n1352 10.6151
R4512 vdd.n1355 vdd.n1354 10.6151
R4513 vdd.n1357 vdd.n1355 10.6151
R4514 vdd.n1358 vdd.n1357 10.6151
R4515 vdd.n1360 vdd.n1358 10.6151
R4516 vdd.n1361 vdd.n1360 10.6151
R4517 vdd.n1363 vdd.n1361 10.6151
R4518 vdd.n1364 vdd.n1363 10.6151
R4519 vdd.n1366 vdd.n1364 10.6151
R4520 vdd.n1367 vdd.n1366 10.6151
R4521 vdd.n1406 vdd.n1367 10.6151
R4522 vdd.n1406 vdd.n1405 10.6151
R4523 vdd.n1405 vdd.n1404 10.6151
R4524 vdd.n1404 vdd.n1402 10.6151
R4525 vdd.n1402 vdd.n1401 10.6151
R4526 vdd.n1401 vdd.n1399 10.6151
R4527 vdd.n1399 vdd.n1398 10.6151
R4528 vdd.n1398 vdd.n1379 10.6151
R4529 vdd.n1379 vdd.n1378 10.6151
R4530 vdd.n1378 vdd.n1376 10.6151
R4531 vdd.n1376 vdd.n1375 10.6151
R4532 vdd.n1375 vdd.n1373 10.6151
R4533 vdd.n1373 vdd.n1372 10.6151
R4534 vdd.n1372 vdd.n1369 10.6151
R4535 vdd.n1369 vdd.n1368 10.6151
R4536 vdd.n1368 vdd.n974 10.6151
R4537 vdd.n2426 vdd.n1110 10.6151
R4538 vdd.n2421 vdd.n1110 10.6151
R4539 vdd.n2421 vdd.n2420 10.6151
R4540 vdd.n2420 vdd.n2419 10.6151
R4541 vdd.n2419 vdd.n2416 10.6151
R4542 vdd.n2416 vdd.n2415 10.6151
R4543 vdd.n2415 vdd.n2412 10.6151
R4544 vdd.n2412 vdd.n2411 10.6151
R4545 vdd.n2411 vdd.n2408 10.6151
R4546 vdd.n2408 vdd.n2407 10.6151
R4547 vdd.n2407 vdd.n2404 10.6151
R4548 vdd.n2404 vdd.n2403 10.6151
R4549 vdd.n2403 vdd.n2400 10.6151
R4550 vdd.n2400 vdd.n2399 10.6151
R4551 vdd.n2399 vdd.n2396 10.6151
R4552 vdd.n2396 vdd.n2395 10.6151
R4553 vdd.n2395 vdd.n2392 10.6151
R4554 vdd.n2392 vdd.n1148 10.6151
R4555 vdd.n1294 vdd.n1148 10.6151
R4556 vdd.n1295 vdd.n1294 10.6151
R4557 vdd.n1298 vdd.n1295 10.6151
R4558 vdd.n1299 vdd.n1298 10.6151
R4559 vdd.n1302 vdd.n1299 10.6151
R4560 vdd.n1303 vdd.n1302 10.6151
R4561 vdd.n1306 vdd.n1303 10.6151
R4562 vdd.n1307 vdd.n1306 10.6151
R4563 vdd.n1310 vdd.n1307 10.6151
R4564 vdd.n1311 vdd.n1310 10.6151
R4565 vdd.n1314 vdd.n1311 10.6151
R4566 vdd.n1315 vdd.n1314 10.6151
R4567 vdd.n1318 vdd.n1315 10.6151
R4568 vdd.n1323 vdd.n1320 10.6151
R4569 vdd.n1324 vdd.n1323 10.6151
R4570 vdd.n2937 vdd.n2936 10.6151
R4571 vdd.n2936 vdd.n2935 10.6151
R4572 vdd.n2935 vdd.n2739 10.6151
R4573 vdd.n2817 vdd.n2739 10.6151
R4574 vdd.n2818 vdd.n2817 10.6151
R4575 vdd.n2820 vdd.n2818 10.6151
R4576 vdd.n2821 vdd.n2820 10.6151
R4577 vdd.n2919 vdd.n2821 10.6151
R4578 vdd.n2919 vdd.n2918 10.6151
R4579 vdd.n2918 vdd.n2917 10.6151
R4580 vdd.n2917 vdd.n2865 10.6151
R4581 vdd.n2865 vdd.n2864 10.6151
R4582 vdd.n2864 vdd.n2862 10.6151
R4583 vdd.n2862 vdd.n2861 10.6151
R4584 vdd.n2861 vdd.n2859 10.6151
R4585 vdd.n2859 vdd.n2858 10.6151
R4586 vdd.n2858 vdd.n2856 10.6151
R4587 vdd.n2856 vdd.n2855 10.6151
R4588 vdd.n2855 vdd.n2853 10.6151
R4589 vdd.n2853 vdd.n2852 10.6151
R4590 vdd.n2852 vdd.n2850 10.6151
R4591 vdd.n2850 vdd.n2849 10.6151
R4592 vdd.n2849 vdd.n2847 10.6151
R4593 vdd.n2847 vdd.n2846 10.6151
R4594 vdd.n2846 vdd.n2844 10.6151
R4595 vdd.n2844 vdd.n2843 10.6151
R4596 vdd.n2843 vdd.n2841 10.6151
R4597 vdd.n2841 vdd.n2840 10.6151
R4598 vdd.n2840 vdd.n2838 10.6151
R4599 vdd.n2838 vdd.n2837 10.6151
R4600 vdd.n2837 vdd.n2835 10.6151
R4601 vdd.n2835 vdd.n2834 10.6151
R4602 vdd.n2834 vdd.n2832 10.6151
R4603 vdd.n2832 vdd.n2831 10.6151
R4604 vdd.n2831 vdd.n2829 10.6151
R4605 vdd.n2829 vdd.n2828 10.6151
R4606 vdd.n2828 vdd.n2826 10.6151
R4607 vdd.n2826 vdd.n2825 10.6151
R4608 vdd.n2825 vdd.n2823 10.6151
R4609 vdd.n2823 vdd.n2822 10.6151
R4610 vdd.n2822 vdd.n807 10.6151
R4611 vdd.n3181 vdd.n807 10.6151
R4612 vdd.n3182 vdd.n3181 10.6151
R4613 vdd.n3008 vdd.n932 10.6151
R4614 vdd.n3003 vdd.n932 10.6151
R4615 vdd.n3003 vdd.n3002 10.6151
R4616 vdd.n3002 vdd.n3001 10.6151
R4617 vdd.n3001 vdd.n2998 10.6151
R4618 vdd.n2998 vdd.n2997 10.6151
R4619 vdd.n2997 vdd.n2994 10.6151
R4620 vdd.n2994 vdd.n2993 10.6151
R4621 vdd.n2993 vdd.n2990 10.6151
R4622 vdd.n2990 vdd.n2989 10.6151
R4623 vdd.n2989 vdd.n2986 10.6151
R4624 vdd.n2986 vdd.n2985 10.6151
R4625 vdd.n2985 vdd.n2982 10.6151
R4626 vdd.n2982 vdd.n2981 10.6151
R4627 vdd.n2981 vdd.n2978 10.6151
R4628 vdd.n2978 vdd.n2977 10.6151
R4629 vdd.n2977 vdd.n2974 10.6151
R4630 vdd.n2974 vdd.n2973 10.6151
R4631 vdd.n2973 vdd.n2970 10.6151
R4632 vdd.n2970 vdd.n2969 10.6151
R4633 vdd.n2969 vdd.n2966 10.6151
R4634 vdd.n2966 vdd.n2965 10.6151
R4635 vdd.n2965 vdd.n2962 10.6151
R4636 vdd.n2962 vdd.n2961 10.6151
R4637 vdd.n2961 vdd.n2958 10.6151
R4638 vdd.n2958 vdd.n2957 10.6151
R4639 vdd.n2957 vdd.n2954 10.6151
R4640 vdd.n2954 vdd.n2953 10.6151
R4641 vdd.n2953 vdd.n2950 10.6151
R4642 vdd.n2950 vdd.n2949 10.6151
R4643 vdd.n2949 vdd.n2946 10.6151
R4644 vdd.n2944 vdd.n2941 10.6151
R4645 vdd.n2941 vdd.n2940 10.6151
R4646 vdd.n3010 vdd.n3009 10.6151
R4647 vdd.n3010 vdd.n921 10.6151
R4648 vdd.n3020 vdd.n921 10.6151
R4649 vdd.n3021 vdd.n3020 10.6151
R4650 vdd.n3022 vdd.n3021 10.6151
R4651 vdd.n3022 vdd.n909 10.6151
R4652 vdd.n3032 vdd.n909 10.6151
R4653 vdd.n3033 vdd.n3032 10.6151
R4654 vdd.n3034 vdd.n3033 10.6151
R4655 vdd.n3034 vdd.n898 10.6151
R4656 vdd.n3044 vdd.n898 10.6151
R4657 vdd.n3045 vdd.n3044 10.6151
R4658 vdd.n3046 vdd.n3045 10.6151
R4659 vdd.n3046 vdd.n887 10.6151
R4660 vdd.n3056 vdd.n887 10.6151
R4661 vdd.n3057 vdd.n3056 10.6151
R4662 vdd.n3058 vdd.n3057 10.6151
R4663 vdd.n3058 vdd.n874 10.6151
R4664 vdd.n3069 vdd.n874 10.6151
R4665 vdd.n3070 vdd.n3069 10.6151
R4666 vdd.n3071 vdd.n3070 10.6151
R4667 vdd.n3071 vdd.n862 10.6151
R4668 vdd.n3081 vdd.n862 10.6151
R4669 vdd.n3082 vdd.n3081 10.6151
R4670 vdd.n3083 vdd.n3082 10.6151
R4671 vdd.n3083 vdd.n850 10.6151
R4672 vdd.n3093 vdd.n850 10.6151
R4673 vdd.n3094 vdd.n3093 10.6151
R4674 vdd.n3095 vdd.n3094 10.6151
R4675 vdd.n3095 vdd.n837 10.6151
R4676 vdd.n3105 vdd.n837 10.6151
R4677 vdd.n3106 vdd.n3105 10.6151
R4678 vdd.n3107 vdd.n3106 10.6151
R4679 vdd.n3107 vdd.n826 10.6151
R4680 vdd.n3117 vdd.n826 10.6151
R4681 vdd.n3118 vdd.n3117 10.6151
R4682 vdd.n3119 vdd.n3118 10.6151
R4683 vdd.n3119 vdd.n812 10.6151
R4684 vdd.n3174 vdd.n812 10.6151
R4685 vdd.n3175 vdd.n3174 10.6151
R4686 vdd.n3176 vdd.n3175 10.6151
R4687 vdd.n3176 vdd.n779 10.6151
R4688 vdd.n3246 vdd.n779 10.6151
R4689 vdd.n3245 vdd.n3244 10.6151
R4690 vdd.n3244 vdd.n780 10.6151
R4691 vdd.n781 vdd.n780 10.6151
R4692 vdd.n3237 vdd.n781 10.6151
R4693 vdd.n3237 vdd.n3236 10.6151
R4694 vdd.n3236 vdd.n3235 10.6151
R4695 vdd.n3235 vdd.n783 10.6151
R4696 vdd.n3230 vdd.n783 10.6151
R4697 vdd.n3230 vdd.n3229 10.6151
R4698 vdd.n3229 vdd.n3228 10.6151
R4699 vdd.n3228 vdd.n786 10.6151
R4700 vdd.n3223 vdd.n786 10.6151
R4701 vdd.n3223 vdd.n3222 10.6151
R4702 vdd.n3222 vdd.n3221 10.6151
R4703 vdd.n3221 vdd.n789 10.6151
R4704 vdd.n3216 vdd.n789 10.6151
R4705 vdd.n3216 vdd.n3215 10.6151
R4706 vdd.n3215 vdd.n3213 10.6151
R4707 vdd.n3213 vdd.n792 10.6151
R4708 vdd.n3208 vdd.n792 10.6151
R4709 vdd.n3208 vdd.n3207 10.6151
R4710 vdd.n3207 vdd.n3206 10.6151
R4711 vdd.n3206 vdd.n795 10.6151
R4712 vdd.n3201 vdd.n795 10.6151
R4713 vdd.n3201 vdd.n3200 10.6151
R4714 vdd.n3200 vdd.n3199 10.6151
R4715 vdd.n3199 vdd.n798 10.6151
R4716 vdd.n3194 vdd.n798 10.6151
R4717 vdd.n3194 vdd.n3193 10.6151
R4718 vdd.n3193 vdd.n3192 10.6151
R4719 vdd.n3192 vdd.n801 10.6151
R4720 vdd.n3187 vdd.n3186 10.6151
R4721 vdd.n3186 vdd.n3185 10.6151
R4722 vdd.n3164 vdd.n3125 10.6151
R4723 vdd.n3159 vdd.n3125 10.6151
R4724 vdd.n3159 vdd.n3158 10.6151
R4725 vdd.n3158 vdd.n3157 10.6151
R4726 vdd.n3157 vdd.n3127 10.6151
R4727 vdd.n3152 vdd.n3127 10.6151
R4728 vdd.n3152 vdd.n3151 10.6151
R4729 vdd.n3151 vdd.n3150 10.6151
R4730 vdd.n3150 vdd.n3130 10.6151
R4731 vdd.n3145 vdd.n3130 10.6151
R4732 vdd.n3145 vdd.n3144 10.6151
R4733 vdd.n3144 vdd.n3143 10.6151
R4734 vdd.n3143 vdd.n3133 10.6151
R4735 vdd.n3138 vdd.n3133 10.6151
R4736 vdd.n3138 vdd.n3137 10.6151
R4737 vdd.n3137 vdd.n753 10.6151
R4738 vdd.n3281 vdd.n753 10.6151
R4739 vdd.n3281 vdd.n754 10.6151
R4740 vdd.n757 vdd.n754 10.6151
R4741 vdd.n3274 vdd.n757 10.6151
R4742 vdd.n3274 vdd.n3273 10.6151
R4743 vdd.n3273 vdd.n3272 10.6151
R4744 vdd.n3272 vdd.n759 10.6151
R4745 vdd.n3267 vdd.n759 10.6151
R4746 vdd.n3267 vdd.n3266 10.6151
R4747 vdd.n3266 vdd.n3265 10.6151
R4748 vdd.n3265 vdd.n762 10.6151
R4749 vdd.n3260 vdd.n762 10.6151
R4750 vdd.n3260 vdd.n3259 10.6151
R4751 vdd.n3259 vdd.n3258 10.6151
R4752 vdd.n3258 vdd.n765 10.6151
R4753 vdd.n3253 vdd.n3252 10.6151
R4754 vdd.n3252 vdd.n3251 10.6151
R4755 vdd.n2814 vdd.n2813 10.6151
R4756 vdd.n2931 vdd.n2814 10.6151
R4757 vdd.n2931 vdd.n2930 10.6151
R4758 vdd.n2930 vdd.n2929 10.6151
R4759 vdd.n2929 vdd.n2927 10.6151
R4760 vdd.n2927 vdd.n2926 10.6151
R4761 vdd.n2926 vdd.n2924 10.6151
R4762 vdd.n2924 vdd.n2923 10.6151
R4763 vdd.n2923 vdd.n2815 10.6151
R4764 vdd.n2913 vdd.n2815 10.6151
R4765 vdd.n2913 vdd.n2912 10.6151
R4766 vdd.n2912 vdd.n2911 10.6151
R4767 vdd.n2911 vdd.n2909 10.6151
R4768 vdd.n2909 vdd.n2908 10.6151
R4769 vdd.n2908 vdd.n2906 10.6151
R4770 vdd.n2906 vdd.n2905 10.6151
R4771 vdd.n2905 vdd.n2903 10.6151
R4772 vdd.n2903 vdd.n2902 10.6151
R4773 vdd.n2902 vdd.n2900 10.6151
R4774 vdd.n2900 vdd.n2899 10.6151
R4775 vdd.n2899 vdd.n2897 10.6151
R4776 vdd.n2897 vdd.n2896 10.6151
R4777 vdd.n2896 vdd.n2894 10.6151
R4778 vdd.n2894 vdd.n2893 10.6151
R4779 vdd.n2893 vdd.n2891 10.6151
R4780 vdd.n2891 vdd.n2890 10.6151
R4781 vdd.n2890 vdd.n2888 10.6151
R4782 vdd.n2888 vdd.n2887 10.6151
R4783 vdd.n2887 vdd.n2885 10.6151
R4784 vdd.n2885 vdd.n2884 10.6151
R4785 vdd.n2884 vdd.n2882 10.6151
R4786 vdd.n2882 vdd.n2881 10.6151
R4787 vdd.n2881 vdd.n2879 10.6151
R4788 vdd.n2879 vdd.n2878 10.6151
R4789 vdd.n2878 vdd.n2876 10.6151
R4790 vdd.n2876 vdd.n2875 10.6151
R4791 vdd.n2875 vdd.n2873 10.6151
R4792 vdd.n2873 vdd.n2872 10.6151
R4793 vdd.n2872 vdd.n2870 10.6151
R4794 vdd.n2870 vdd.n2869 10.6151
R4795 vdd.n2869 vdd.n2867 10.6151
R4796 vdd.n2867 vdd.n2866 10.6151
R4797 vdd.n2866 vdd.n771 10.6151
R4798 vdd.n2745 vdd.n2744 10.6151
R4799 vdd.n2748 vdd.n2745 10.6151
R4800 vdd.n2749 vdd.n2748 10.6151
R4801 vdd.n2752 vdd.n2749 10.6151
R4802 vdd.n2753 vdd.n2752 10.6151
R4803 vdd.n2756 vdd.n2753 10.6151
R4804 vdd.n2757 vdd.n2756 10.6151
R4805 vdd.n2760 vdd.n2757 10.6151
R4806 vdd.n2761 vdd.n2760 10.6151
R4807 vdd.n2764 vdd.n2761 10.6151
R4808 vdd.n2765 vdd.n2764 10.6151
R4809 vdd.n2768 vdd.n2765 10.6151
R4810 vdd.n2769 vdd.n2768 10.6151
R4811 vdd.n2772 vdd.n2769 10.6151
R4812 vdd.n2773 vdd.n2772 10.6151
R4813 vdd.n2776 vdd.n2773 10.6151
R4814 vdd.n2777 vdd.n2776 10.6151
R4815 vdd.n2780 vdd.n2777 10.6151
R4816 vdd.n2781 vdd.n2780 10.6151
R4817 vdd.n2784 vdd.n2781 10.6151
R4818 vdd.n2785 vdd.n2784 10.6151
R4819 vdd.n2788 vdd.n2785 10.6151
R4820 vdd.n2789 vdd.n2788 10.6151
R4821 vdd.n2792 vdd.n2789 10.6151
R4822 vdd.n2793 vdd.n2792 10.6151
R4823 vdd.n2796 vdd.n2793 10.6151
R4824 vdd.n2797 vdd.n2796 10.6151
R4825 vdd.n2800 vdd.n2797 10.6151
R4826 vdd.n2801 vdd.n2800 10.6151
R4827 vdd.n2804 vdd.n2801 10.6151
R4828 vdd.n2805 vdd.n2804 10.6151
R4829 vdd.n2810 vdd.n2808 10.6151
R4830 vdd.n2811 vdd.n2810 10.6151
R4831 vdd.n3014 vdd.n926 10.6151
R4832 vdd.n3015 vdd.n3014 10.6151
R4833 vdd.n3016 vdd.n3015 10.6151
R4834 vdd.n3016 vdd.n915 10.6151
R4835 vdd.n3026 vdd.n915 10.6151
R4836 vdd.n3027 vdd.n3026 10.6151
R4837 vdd.n3028 vdd.n3027 10.6151
R4838 vdd.n3028 vdd.n904 10.6151
R4839 vdd.n3038 vdd.n904 10.6151
R4840 vdd.n3039 vdd.n3038 10.6151
R4841 vdd.n3040 vdd.n3039 10.6151
R4842 vdd.n3040 vdd.n892 10.6151
R4843 vdd.n3050 vdd.n892 10.6151
R4844 vdd.n3051 vdd.n3050 10.6151
R4845 vdd.n3052 vdd.n3051 10.6151
R4846 vdd.n3052 vdd.n881 10.6151
R4847 vdd.n3062 vdd.n881 10.6151
R4848 vdd.n3063 vdd.n3062 10.6151
R4849 vdd.n3065 vdd.n3063 10.6151
R4850 vdd.n3065 vdd.n3064 10.6151
R4851 vdd.n3076 vdd.n3075 10.6151
R4852 vdd.n3077 vdd.n3076 10.6151
R4853 vdd.n3077 vdd.n856 10.6151
R4854 vdd.n3087 vdd.n856 10.6151
R4855 vdd.n3088 vdd.n3087 10.6151
R4856 vdd.n3089 vdd.n3088 10.6151
R4857 vdd.n3089 vdd.n843 10.6151
R4858 vdd.n3099 vdd.n843 10.6151
R4859 vdd.n3100 vdd.n3099 10.6151
R4860 vdd.n3101 vdd.n3100 10.6151
R4861 vdd.n3101 vdd.n831 10.6151
R4862 vdd.n3111 vdd.n831 10.6151
R4863 vdd.n3112 vdd.n3111 10.6151
R4864 vdd.n3113 vdd.n3112 10.6151
R4865 vdd.n3113 vdd.n820 10.6151
R4866 vdd.n3123 vdd.n820 10.6151
R4867 vdd.n3124 vdd.n3123 10.6151
R4868 vdd.n3170 vdd.n3124 10.6151
R4869 vdd.n3170 vdd.n3169 10.6151
R4870 vdd.n3169 vdd.n3168 10.6151
R4871 vdd.n3168 vdd.n3167 10.6151
R4872 vdd.n3167 vdd.n3165 10.6151
R4873 vdd.n2432 vdd.n1103 10.6151
R4874 vdd.n2433 vdd.n2432 10.6151
R4875 vdd.n2434 vdd.n2433 10.6151
R4876 vdd.n2434 vdd.n1092 10.6151
R4877 vdd.n2444 vdd.n1092 10.6151
R4878 vdd.n2445 vdd.n2444 10.6151
R4879 vdd.n2446 vdd.n2445 10.6151
R4880 vdd.n2446 vdd.n1079 10.6151
R4881 vdd.n2456 vdd.n1079 10.6151
R4882 vdd.n2457 vdd.n2456 10.6151
R4883 vdd.n2458 vdd.n2457 10.6151
R4884 vdd.n2458 vdd.n1068 10.6151
R4885 vdd.n2468 vdd.n1068 10.6151
R4886 vdd.n2469 vdd.n2468 10.6151
R4887 vdd.n2470 vdd.n2469 10.6151
R4888 vdd.n2470 vdd.n1056 10.6151
R4889 vdd.n2480 vdd.n1056 10.6151
R4890 vdd.n2481 vdd.n2480 10.6151
R4891 vdd.n2482 vdd.n2481 10.6151
R4892 vdd.n2482 vdd.n1043 10.6151
R4893 vdd.n2492 vdd.n1043 10.6151
R4894 vdd.n2493 vdd.n2492 10.6151
R4895 vdd.n2495 vdd.n1031 10.6151
R4896 vdd.n2505 vdd.n1031 10.6151
R4897 vdd.n2506 vdd.n2505 10.6151
R4898 vdd.n2507 vdd.n2506 10.6151
R4899 vdd.n2507 vdd.n1019 10.6151
R4900 vdd.n2517 vdd.n1019 10.6151
R4901 vdd.n2518 vdd.n2517 10.6151
R4902 vdd.n2519 vdd.n2518 10.6151
R4903 vdd.n2519 vdd.n1008 10.6151
R4904 vdd.n2529 vdd.n1008 10.6151
R4905 vdd.n2530 vdd.n2529 10.6151
R4906 vdd.n2531 vdd.n2530 10.6151
R4907 vdd.n2531 vdd.n997 10.6151
R4908 vdd.n2541 vdd.n997 10.6151
R4909 vdd.n2542 vdd.n2541 10.6151
R4910 vdd.n2545 vdd.n2542 10.6151
R4911 vdd.n2545 vdd.n2544 10.6151
R4912 vdd.n2544 vdd.n2543 10.6151
R4913 vdd.n2543 vdd.n980 10.6151
R4914 vdd.n2627 vdd.n980 10.6151
R4915 vdd.n2626 vdd.n2625 10.6151
R4916 vdd.n2625 vdd.n2622 10.6151
R4917 vdd.n2622 vdd.n2621 10.6151
R4918 vdd.n2621 vdd.n2618 10.6151
R4919 vdd.n2618 vdd.n2617 10.6151
R4920 vdd.n2617 vdd.n2614 10.6151
R4921 vdd.n2614 vdd.n2613 10.6151
R4922 vdd.n2613 vdd.n2610 10.6151
R4923 vdd.n2610 vdd.n2609 10.6151
R4924 vdd.n2609 vdd.n2606 10.6151
R4925 vdd.n2606 vdd.n2605 10.6151
R4926 vdd.n2605 vdd.n2602 10.6151
R4927 vdd.n2602 vdd.n2601 10.6151
R4928 vdd.n2601 vdd.n2598 10.6151
R4929 vdd.n2598 vdd.n2597 10.6151
R4930 vdd.n2597 vdd.n2594 10.6151
R4931 vdd.n2594 vdd.n2593 10.6151
R4932 vdd.n2593 vdd.n2590 10.6151
R4933 vdd.n2590 vdd.n2589 10.6151
R4934 vdd.n2589 vdd.n2586 10.6151
R4935 vdd.n2586 vdd.n2585 10.6151
R4936 vdd.n2585 vdd.n2582 10.6151
R4937 vdd.n2582 vdd.n2581 10.6151
R4938 vdd.n2581 vdd.n2578 10.6151
R4939 vdd.n2578 vdd.n2577 10.6151
R4940 vdd.n2577 vdd.n2574 10.6151
R4941 vdd.n2574 vdd.n2573 10.6151
R4942 vdd.n2573 vdd.n2570 10.6151
R4943 vdd.n2570 vdd.n2569 10.6151
R4944 vdd.n2569 vdd.n2566 10.6151
R4945 vdd.n2566 vdd.n2565 10.6151
R4946 vdd.n2562 vdd.n2561 10.6151
R4947 vdd.n2561 vdd.n2559 10.6151
R4948 vdd.n1452 vdd.n1450 10.6151
R4949 vdd.n1450 vdd.n1449 10.6151
R4950 vdd.n1449 vdd.n1447 10.6151
R4951 vdd.n1447 vdd.n1446 10.6151
R4952 vdd.n1446 vdd.n1444 10.6151
R4953 vdd.n1444 vdd.n1443 10.6151
R4954 vdd.n1443 vdd.n1441 10.6151
R4955 vdd.n1441 vdd.n1440 10.6151
R4956 vdd.n1440 vdd.n1438 10.6151
R4957 vdd.n1438 vdd.n1437 10.6151
R4958 vdd.n1437 vdd.n1435 10.6151
R4959 vdd.n1435 vdd.n1434 10.6151
R4960 vdd.n1434 vdd.n1432 10.6151
R4961 vdd.n1432 vdd.n1431 10.6151
R4962 vdd.n1431 vdd.n1429 10.6151
R4963 vdd.n1429 vdd.n1428 10.6151
R4964 vdd.n1428 vdd.n1426 10.6151
R4965 vdd.n1426 vdd.n1425 10.6151
R4966 vdd.n1425 vdd.n1423 10.6151
R4967 vdd.n1423 vdd.n1422 10.6151
R4968 vdd.n1422 vdd.n1420 10.6151
R4969 vdd.n1420 vdd.n1419 10.6151
R4970 vdd.n1419 vdd.n1417 10.6151
R4971 vdd.n1417 vdd.n1416 10.6151
R4972 vdd.n1416 vdd.n1414 10.6151
R4973 vdd.n1414 vdd.n1413 10.6151
R4974 vdd.n1413 vdd.n1411 10.6151
R4975 vdd.n1411 vdd.n1410 10.6151
R4976 vdd.n1410 vdd.n1289 10.6151
R4977 vdd.n1381 vdd.n1289 10.6151
R4978 vdd.n1382 vdd.n1381 10.6151
R4979 vdd.n1384 vdd.n1382 10.6151
R4980 vdd.n1385 vdd.n1384 10.6151
R4981 vdd.n1394 vdd.n1385 10.6151
R4982 vdd.n1394 vdd.n1393 10.6151
R4983 vdd.n1393 vdd.n1392 10.6151
R4984 vdd.n1392 vdd.n1390 10.6151
R4985 vdd.n1390 vdd.n1389 10.6151
R4986 vdd.n1389 vdd.n1387 10.6151
R4987 vdd.n1387 vdd.n1386 10.6151
R4988 vdd.n1386 vdd.n984 10.6151
R4989 vdd.n2557 vdd.n984 10.6151
R4990 vdd.n2558 vdd.n2557 10.6151
R4991 vdd.n1253 vdd.n1252 10.6151
R4992 vdd.n1256 vdd.n1253 10.6151
R4993 vdd.n1257 vdd.n1256 10.6151
R4994 vdd.n1260 vdd.n1257 10.6151
R4995 vdd.n1261 vdd.n1260 10.6151
R4996 vdd.n1264 vdd.n1261 10.6151
R4997 vdd.n1265 vdd.n1264 10.6151
R4998 vdd.n1268 vdd.n1265 10.6151
R4999 vdd.n1269 vdd.n1268 10.6151
R5000 vdd.n1272 vdd.n1269 10.6151
R5001 vdd.n1273 vdd.n1272 10.6151
R5002 vdd.n1276 vdd.n1273 10.6151
R5003 vdd.n1277 vdd.n1276 10.6151
R5004 vdd.n1280 vdd.n1277 10.6151
R5005 vdd.n1281 vdd.n1280 10.6151
R5006 vdd.n1284 vdd.n1281 10.6151
R5007 vdd.n1486 vdd.n1284 10.6151
R5008 vdd.n1486 vdd.n1485 10.6151
R5009 vdd.n1485 vdd.n1483 10.6151
R5010 vdd.n1483 vdd.n1480 10.6151
R5011 vdd.n1480 vdd.n1479 10.6151
R5012 vdd.n1479 vdd.n1476 10.6151
R5013 vdd.n1476 vdd.n1475 10.6151
R5014 vdd.n1475 vdd.n1472 10.6151
R5015 vdd.n1472 vdd.n1471 10.6151
R5016 vdd.n1471 vdd.n1468 10.6151
R5017 vdd.n1468 vdd.n1467 10.6151
R5018 vdd.n1467 vdd.n1464 10.6151
R5019 vdd.n1464 vdd.n1463 10.6151
R5020 vdd.n1463 vdd.n1460 10.6151
R5021 vdd.n1460 vdd.n1459 10.6151
R5022 vdd.n1456 vdd.n1455 10.6151
R5023 vdd.n1455 vdd.n1453 10.6151
R5024 vdd.t19 vdd.n2231 10.5435
R5025 vdd.n636 vdd.t21 10.5435
R5026 vdd.n304 vdd.n286 10.4732
R5027 vdd.n249 vdd.n231 10.4732
R5028 vdd.n206 vdd.n188 10.4732
R5029 vdd.n151 vdd.n133 10.4732
R5030 vdd.n109 vdd.n91 10.4732
R5031 vdd.n54 vdd.n36 10.4732
R5032 vdd.n2128 vdd.n2110 10.4732
R5033 vdd.n2183 vdd.n2165 10.4732
R5034 vdd.n2030 vdd.n2012 10.4732
R5035 vdd.n2085 vdd.n2067 10.4732
R5036 vdd.n1933 vdd.n1915 10.4732
R5037 vdd.n1988 vdd.n1970 10.4732
R5038 vdd.n2215 vdd.t15 10.3167
R5039 vdd.n3477 vdd.t141 10.3167
R5040 vdd.t27 vdd.n1559 10.09
R5041 vdd.n2267 vdd.t74 10.09
R5042 vdd.n3425 vdd.t88 10.09
R5043 vdd.n3558 vdd.t0 10.09
R5044 vdd.n2392 vdd.n2391 9.98956
R5045 vdd.n3215 vdd.n3214 9.98956
R5046 vdd.n3282 vdd.n3281 9.98956
R5047 vdd.n2284 vdd.n1486 9.98956
R5048 vdd.n1879 vdd.t161 9.86327
R5049 vdd.n3549 vdd.t43 9.86327
R5050 vdd.n2629 vdd.t242 9.7499
R5051 vdd.t227 vdd.n928 9.7499
R5052 vdd.n303 vdd.n288 9.69747
R5053 vdd.n248 vdd.n233 9.69747
R5054 vdd.n205 vdd.n190 9.69747
R5055 vdd.n150 vdd.n135 9.69747
R5056 vdd.n108 vdd.n93 9.69747
R5057 vdd.n53 vdd.n38 9.69747
R5058 vdd.n2127 vdd.n2112 9.69747
R5059 vdd.n2182 vdd.n2167 9.69747
R5060 vdd.n2029 vdd.n2014 9.69747
R5061 vdd.n2084 vdd.n2069 9.69747
R5062 vdd.n1932 vdd.n1917 9.69747
R5063 vdd.n1987 vdd.n1972 9.69747
R5064 vdd.t47 vdd.n1853 9.63654
R5065 vdd.n3508 vdd.t56 9.63654
R5066 vdd.n319 vdd.n318 9.45567
R5067 vdd.n264 vdd.n263 9.45567
R5068 vdd.n221 vdd.n220 9.45567
R5069 vdd.n166 vdd.n165 9.45567
R5070 vdd.n124 vdd.n123 9.45567
R5071 vdd.n69 vdd.n68 9.45567
R5072 vdd.n2143 vdd.n2142 9.45567
R5073 vdd.n2198 vdd.n2197 9.45567
R5074 vdd.n2045 vdd.n2044 9.45567
R5075 vdd.n2100 vdd.n2099 9.45567
R5076 vdd.n1948 vdd.n1947 9.45567
R5077 vdd.n2003 vdd.n2002 9.45567
R5078 vdd.n2354 vdd.n1178 9.3005
R5079 vdd.n2353 vdd.n2352 9.3005
R5080 vdd.n1184 vdd.n1183 9.3005
R5081 vdd.n2347 vdd.n1188 9.3005
R5082 vdd.n2346 vdd.n1189 9.3005
R5083 vdd.n2345 vdd.n1190 9.3005
R5084 vdd.n1194 vdd.n1191 9.3005
R5085 vdd.n2340 vdd.n1195 9.3005
R5086 vdd.n2339 vdd.n1196 9.3005
R5087 vdd.n2338 vdd.n1197 9.3005
R5088 vdd.n1201 vdd.n1198 9.3005
R5089 vdd.n2333 vdd.n1202 9.3005
R5090 vdd.n2332 vdd.n1203 9.3005
R5091 vdd.n2331 vdd.n1204 9.3005
R5092 vdd.n1208 vdd.n1205 9.3005
R5093 vdd.n2326 vdd.n1209 9.3005
R5094 vdd.n2325 vdd.n1210 9.3005
R5095 vdd.n2324 vdd.n1211 9.3005
R5096 vdd.n1215 vdd.n1212 9.3005
R5097 vdd.n2319 vdd.n1216 9.3005
R5098 vdd.n2318 vdd.n1217 9.3005
R5099 vdd.n2317 vdd.n2316 9.3005
R5100 vdd.n2315 vdd.n1218 9.3005
R5101 vdd.n2314 vdd.n2313 9.3005
R5102 vdd.n1224 vdd.n1223 9.3005
R5103 vdd.n2308 vdd.n1228 9.3005
R5104 vdd.n2307 vdd.n1229 9.3005
R5105 vdd.n2306 vdd.n1230 9.3005
R5106 vdd.n1234 vdd.n1231 9.3005
R5107 vdd.n2301 vdd.n1235 9.3005
R5108 vdd.n2300 vdd.n1236 9.3005
R5109 vdd.n2299 vdd.n1237 9.3005
R5110 vdd.n1241 vdd.n1238 9.3005
R5111 vdd.n2294 vdd.n1242 9.3005
R5112 vdd.n2293 vdd.n1243 9.3005
R5113 vdd.n2292 vdd.n1244 9.3005
R5114 vdd.n1248 vdd.n1245 9.3005
R5115 vdd.n2287 vdd.n1249 9.3005
R5116 vdd.n2356 vdd.n2355 9.3005
R5117 vdd.n2378 vdd.n1149 9.3005
R5118 vdd.n2377 vdd.n1157 9.3005
R5119 vdd.n1161 vdd.n1158 9.3005
R5120 vdd.n2372 vdd.n1162 9.3005
R5121 vdd.n2371 vdd.n1163 9.3005
R5122 vdd.n2370 vdd.n1164 9.3005
R5123 vdd.n1168 vdd.n1165 9.3005
R5124 vdd.n2365 vdd.n1169 9.3005
R5125 vdd.n2364 vdd.n1170 9.3005
R5126 vdd.n2363 vdd.n1171 9.3005
R5127 vdd.n1175 vdd.n1172 9.3005
R5128 vdd.n2358 vdd.n1176 9.3005
R5129 vdd.n2357 vdd.n1177 9.3005
R5130 vdd.n2390 vdd.n2389 9.3005
R5131 vdd.n1153 vdd.n1152 9.3005
R5132 vdd.n2203 vdd.n1549 9.3005
R5133 vdd.n2205 vdd.n2204 9.3005
R5134 vdd.n1540 vdd.n1539 9.3005
R5135 vdd.n2218 vdd.n2217 9.3005
R5136 vdd.n2219 vdd.n1538 9.3005
R5137 vdd.n2221 vdd.n2220 9.3005
R5138 vdd.n1528 vdd.n1527 9.3005
R5139 vdd.n2235 vdd.n2234 9.3005
R5140 vdd.n2236 vdd.n1526 9.3005
R5141 vdd.n2238 vdd.n2237 9.3005
R5142 vdd.n1517 vdd.n1516 9.3005
R5143 vdd.n2252 vdd.n2251 9.3005
R5144 vdd.n2253 vdd.n1515 9.3005
R5145 vdd.n2255 vdd.n2254 9.3005
R5146 vdd.n1505 vdd.n1504 9.3005
R5147 vdd.n2270 vdd.n2269 9.3005
R5148 vdd.n2271 vdd.n1503 9.3005
R5149 vdd.n2273 vdd.n2272 9.3005
R5150 vdd.n295 vdd.n294 9.3005
R5151 vdd.n290 vdd.n289 9.3005
R5152 vdd.n301 vdd.n300 9.3005
R5153 vdd.n303 vdd.n302 9.3005
R5154 vdd.n286 vdd.n285 9.3005
R5155 vdd.n309 vdd.n308 9.3005
R5156 vdd.n311 vdd.n310 9.3005
R5157 vdd.n283 vdd.n280 9.3005
R5158 vdd.n318 vdd.n317 9.3005
R5159 vdd.n240 vdd.n239 9.3005
R5160 vdd.n235 vdd.n234 9.3005
R5161 vdd.n246 vdd.n245 9.3005
R5162 vdd.n248 vdd.n247 9.3005
R5163 vdd.n231 vdd.n230 9.3005
R5164 vdd.n254 vdd.n253 9.3005
R5165 vdd.n256 vdd.n255 9.3005
R5166 vdd.n228 vdd.n225 9.3005
R5167 vdd.n263 vdd.n262 9.3005
R5168 vdd.n197 vdd.n196 9.3005
R5169 vdd.n192 vdd.n191 9.3005
R5170 vdd.n203 vdd.n202 9.3005
R5171 vdd.n205 vdd.n204 9.3005
R5172 vdd.n188 vdd.n187 9.3005
R5173 vdd.n211 vdd.n210 9.3005
R5174 vdd.n213 vdd.n212 9.3005
R5175 vdd.n185 vdd.n182 9.3005
R5176 vdd.n220 vdd.n219 9.3005
R5177 vdd.n142 vdd.n141 9.3005
R5178 vdd.n137 vdd.n136 9.3005
R5179 vdd.n148 vdd.n147 9.3005
R5180 vdd.n150 vdd.n149 9.3005
R5181 vdd.n133 vdd.n132 9.3005
R5182 vdd.n156 vdd.n155 9.3005
R5183 vdd.n158 vdd.n157 9.3005
R5184 vdd.n130 vdd.n127 9.3005
R5185 vdd.n165 vdd.n164 9.3005
R5186 vdd.n100 vdd.n99 9.3005
R5187 vdd.n95 vdd.n94 9.3005
R5188 vdd.n106 vdd.n105 9.3005
R5189 vdd.n108 vdd.n107 9.3005
R5190 vdd.n91 vdd.n90 9.3005
R5191 vdd.n114 vdd.n113 9.3005
R5192 vdd.n116 vdd.n115 9.3005
R5193 vdd.n88 vdd.n85 9.3005
R5194 vdd.n123 vdd.n122 9.3005
R5195 vdd.n45 vdd.n44 9.3005
R5196 vdd.n40 vdd.n39 9.3005
R5197 vdd.n51 vdd.n50 9.3005
R5198 vdd.n53 vdd.n52 9.3005
R5199 vdd.n36 vdd.n35 9.3005
R5200 vdd.n59 vdd.n58 9.3005
R5201 vdd.n61 vdd.n60 9.3005
R5202 vdd.n33 vdd.n30 9.3005
R5203 vdd.n68 vdd.n67 9.3005
R5204 vdd.n3331 vdd.n3330 9.3005
R5205 vdd.n3332 vdd.n721 9.3005
R5206 vdd.n720 vdd.n718 9.3005
R5207 vdd.n3338 vdd.n717 9.3005
R5208 vdd.n3339 vdd.n716 9.3005
R5209 vdd.n3340 vdd.n715 9.3005
R5210 vdd.n714 vdd.n712 9.3005
R5211 vdd.n3346 vdd.n711 9.3005
R5212 vdd.n3347 vdd.n710 9.3005
R5213 vdd.n3348 vdd.n709 9.3005
R5214 vdd.n708 vdd.n706 9.3005
R5215 vdd.n3354 vdd.n705 9.3005
R5216 vdd.n3355 vdd.n704 9.3005
R5217 vdd.n3356 vdd.n703 9.3005
R5218 vdd.n702 vdd.n700 9.3005
R5219 vdd.n3362 vdd.n699 9.3005
R5220 vdd.n3363 vdd.n698 9.3005
R5221 vdd.n3364 vdd.n697 9.3005
R5222 vdd.n696 vdd.n694 9.3005
R5223 vdd.n3370 vdd.n693 9.3005
R5224 vdd.n3371 vdd.n692 9.3005
R5225 vdd.n3372 vdd.n691 9.3005
R5226 vdd.n690 vdd.n688 9.3005
R5227 vdd.n3378 vdd.n685 9.3005
R5228 vdd.n3379 vdd.n684 9.3005
R5229 vdd.n3380 vdd.n683 9.3005
R5230 vdd.n682 vdd.n680 9.3005
R5231 vdd.n3386 vdd.n679 9.3005
R5232 vdd.n3387 vdd.n678 9.3005
R5233 vdd.n3388 vdd.n677 9.3005
R5234 vdd.n676 vdd.n674 9.3005
R5235 vdd.n3394 vdd.n673 9.3005
R5236 vdd.n3395 vdd.n672 9.3005
R5237 vdd.n3396 vdd.n671 9.3005
R5238 vdd.n670 vdd.n668 9.3005
R5239 vdd.n3401 vdd.n667 9.3005
R5240 vdd.n3411 vdd.n661 9.3005
R5241 vdd.n3413 vdd.n3412 9.3005
R5242 vdd.n652 vdd.n651 9.3005
R5243 vdd.n3428 vdd.n3427 9.3005
R5244 vdd.n3429 vdd.n650 9.3005
R5245 vdd.n3431 vdd.n3430 9.3005
R5246 vdd.n640 vdd.n639 9.3005
R5247 vdd.n3444 vdd.n3443 9.3005
R5248 vdd.n3445 vdd.n638 9.3005
R5249 vdd.n3447 vdd.n3446 9.3005
R5250 vdd.n628 vdd.n627 9.3005
R5251 vdd.n3461 vdd.n3460 9.3005
R5252 vdd.n3462 vdd.n626 9.3005
R5253 vdd.n3464 vdd.n3463 9.3005
R5254 vdd.n617 vdd.n616 9.3005
R5255 vdd.n3480 vdd.n3479 9.3005
R5256 vdd.n3481 vdd.n615 9.3005
R5257 vdd.n3483 vdd.n3482 9.3005
R5258 vdd.n324 vdd.n322 9.3005
R5259 vdd.n3415 vdd.n3414 9.3005
R5260 vdd.n3562 vdd.n3561 9.3005
R5261 vdd.n325 vdd.n323 9.3005
R5262 vdd.n3555 vdd.n334 9.3005
R5263 vdd.n3554 vdd.n335 9.3005
R5264 vdd.n3553 vdd.n336 9.3005
R5265 vdd.n343 vdd.n337 9.3005
R5266 vdd.n3547 vdd.n344 9.3005
R5267 vdd.n3546 vdd.n345 9.3005
R5268 vdd.n3545 vdd.n346 9.3005
R5269 vdd.n354 vdd.n347 9.3005
R5270 vdd.n3539 vdd.n355 9.3005
R5271 vdd.n3538 vdd.n356 9.3005
R5272 vdd.n3537 vdd.n357 9.3005
R5273 vdd.n365 vdd.n358 9.3005
R5274 vdd.n3531 vdd.n366 9.3005
R5275 vdd.n3530 vdd.n367 9.3005
R5276 vdd.n3529 vdd.n368 9.3005
R5277 vdd.n443 vdd.n369 9.3005
R5278 vdd.n447 vdd.n442 9.3005
R5279 vdd.n451 vdd.n450 9.3005
R5280 vdd.n452 vdd.n441 9.3005
R5281 vdd.n456 vdd.n453 9.3005
R5282 vdd.n457 vdd.n440 9.3005
R5283 vdd.n461 vdd.n460 9.3005
R5284 vdd.n462 vdd.n439 9.3005
R5285 vdd.n466 vdd.n463 9.3005
R5286 vdd.n467 vdd.n438 9.3005
R5287 vdd.n471 vdd.n470 9.3005
R5288 vdd.n472 vdd.n437 9.3005
R5289 vdd.n476 vdd.n473 9.3005
R5290 vdd.n477 vdd.n436 9.3005
R5291 vdd.n481 vdd.n480 9.3005
R5292 vdd.n482 vdd.n435 9.3005
R5293 vdd.n486 vdd.n483 9.3005
R5294 vdd.n487 vdd.n434 9.3005
R5295 vdd.n491 vdd.n490 9.3005
R5296 vdd.n492 vdd.n433 9.3005
R5297 vdd.n496 vdd.n493 9.3005
R5298 vdd.n497 vdd.n430 9.3005
R5299 vdd.n501 vdd.n500 9.3005
R5300 vdd.n502 vdd.n429 9.3005
R5301 vdd.n506 vdd.n503 9.3005
R5302 vdd.n507 vdd.n428 9.3005
R5303 vdd.n511 vdd.n510 9.3005
R5304 vdd.n512 vdd.n427 9.3005
R5305 vdd.n516 vdd.n513 9.3005
R5306 vdd.n517 vdd.n426 9.3005
R5307 vdd.n521 vdd.n520 9.3005
R5308 vdd.n522 vdd.n425 9.3005
R5309 vdd.n526 vdd.n523 9.3005
R5310 vdd.n527 vdd.n424 9.3005
R5311 vdd.n531 vdd.n530 9.3005
R5312 vdd.n532 vdd.n423 9.3005
R5313 vdd.n536 vdd.n533 9.3005
R5314 vdd.n537 vdd.n422 9.3005
R5315 vdd.n541 vdd.n540 9.3005
R5316 vdd.n542 vdd.n421 9.3005
R5317 vdd.n546 vdd.n543 9.3005
R5318 vdd.n547 vdd.n418 9.3005
R5319 vdd.n551 vdd.n550 9.3005
R5320 vdd.n552 vdd.n417 9.3005
R5321 vdd.n556 vdd.n553 9.3005
R5322 vdd.n557 vdd.n416 9.3005
R5323 vdd.n561 vdd.n560 9.3005
R5324 vdd.n562 vdd.n415 9.3005
R5325 vdd.n566 vdd.n563 9.3005
R5326 vdd.n567 vdd.n414 9.3005
R5327 vdd.n571 vdd.n570 9.3005
R5328 vdd.n572 vdd.n413 9.3005
R5329 vdd.n576 vdd.n573 9.3005
R5330 vdd.n577 vdd.n412 9.3005
R5331 vdd.n581 vdd.n580 9.3005
R5332 vdd.n582 vdd.n411 9.3005
R5333 vdd.n586 vdd.n583 9.3005
R5334 vdd.n587 vdd.n410 9.3005
R5335 vdd.n591 vdd.n590 9.3005
R5336 vdd.n592 vdd.n409 9.3005
R5337 vdd.n596 vdd.n593 9.3005
R5338 vdd.n598 vdd.n408 9.3005
R5339 vdd.n600 vdd.n599 9.3005
R5340 vdd.n3522 vdd.n3521 9.3005
R5341 vdd.n446 vdd.n444 9.3005
R5342 vdd.n3421 vdd.n655 9.3005
R5343 vdd.n3423 vdd.n3422 9.3005
R5344 vdd.n646 vdd.n645 9.3005
R5345 vdd.n3436 vdd.n3435 9.3005
R5346 vdd.n3437 vdd.n644 9.3005
R5347 vdd.n3439 vdd.n3438 9.3005
R5348 vdd.n633 vdd.n632 9.3005
R5349 vdd.n3452 vdd.n3451 9.3005
R5350 vdd.n3453 vdd.n631 9.3005
R5351 vdd.n3455 vdd.n3454 9.3005
R5352 vdd.n622 vdd.n621 9.3005
R5353 vdd.n3469 vdd.n3468 9.3005
R5354 vdd.n3470 vdd.n620 9.3005
R5355 vdd.n3475 vdd.n3471 9.3005
R5356 vdd.n3474 vdd.n3473 9.3005
R5357 vdd.n3472 vdd.n610 9.3005
R5358 vdd.n3488 vdd.n611 9.3005
R5359 vdd.n3489 vdd.n609 9.3005
R5360 vdd.n3491 vdd.n3490 9.3005
R5361 vdd.n3492 vdd.n608 9.3005
R5362 vdd.n3495 vdd.n3493 9.3005
R5363 vdd.n3496 vdd.n607 9.3005
R5364 vdd.n3498 vdd.n3497 9.3005
R5365 vdd.n3499 vdd.n606 9.3005
R5366 vdd.n3502 vdd.n3500 9.3005
R5367 vdd.n3503 vdd.n605 9.3005
R5368 vdd.n3505 vdd.n3504 9.3005
R5369 vdd.n3506 vdd.n604 9.3005
R5370 vdd.n3510 vdd.n3507 9.3005
R5371 vdd.n3511 vdd.n603 9.3005
R5372 vdd.n3513 vdd.n3512 9.3005
R5373 vdd.n3514 vdd.n602 9.3005
R5374 vdd.n3517 vdd.n3515 9.3005
R5375 vdd.n3518 vdd.n601 9.3005
R5376 vdd.n3520 vdd.n3519 9.3005
R5377 vdd.n3420 vdd.n3419 9.3005
R5378 vdd.n3284 vdd.n656 9.3005
R5379 vdd.n3289 vdd.n3283 9.3005
R5380 vdd.n3299 vdd.n748 9.3005
R5381 vdd.n3300 vdd.n747 9.3005
R5382 vdd.n746 vdd.n744 9.3005
R5383 vdd.n3306 vdd.n743 9.3005
R5384 vdd.n3307 vdd.n742 9.3005
R5385 vdd.n3308 vdd.n741 9.3005
R5386 vdd.n740 vdd.n738 9.3005
R5387 vdd.n3314 vdd.n737 9.3005
R5388 vdd.n3315 vdd.n736 9.3005
R5389 vdd.n3316 vdd.n735 9.3005
R5390 vdd.n734 vdd.n732 9.3005
R5391 vdd.n3321 vdd.n731 9.3005
R5392 vdd.n3322 vdd.n730 9.3005
R5393 vdd.n726 vdd.n725 9.3005
R5394 vdd.n3328 vdd.n3327 9.3005
R5395 vdd.n3329 vdd.n722 9.3005
R5396 vdd.n2283 vdd.n2282 9.3005
R5397 vdd.n2278 vdd.n1488 9.3005
R5398 vdd.n1835 vdd.n1834 9.3005
R5399 vdd.n1591 vdd.n1590 9.3005
R5400 vdd.n1848 vdd.n1847 9.3005
R5401 vdd.n1849 vdd.n1589 9.3005
R5402 vdd.n1851 vdd.n1850 9.3005
R5403 vdd.n1579 vdd.n1578 9.3005
R5404 vdd.n1865 vdd.n1864 9.3005
R5405 vdd.n1866 vdd.n1577 9.3005
R5406 vdd.n1868 vdd.n1867 9.3005
R5407 vdd.n1569 vdd.n1568 9.3005
R5408 vdd.n1882 vdd.n1881 9.3005
R5409 vdd.n1883 vdd.n1567 9.3005
R5410 vdd.n1885 vdd.n1884 9.3005
R5411 vdd.n1556 vdd.n1555 9.3005
R5412 vdd.n1898 vdd.n1897 9.3005
R5413 vdd.n1899 vdd.n1554 9.3005
R5414 vdd.n1901 vdd.n1900 9.3005
R5415 vdd.n1545 vdd.n1544 9.3005
R5416 vdd.n2210 vdd.n2209 9.3005
R5417 vdd.n2211 vdd.n1543 9.3005
R5418 vdd.n2213 vdd.n2212 9.3005
R5419 vdd.n1534 vdd.n1533 9.3005
R5420 vdd.n2226 vdd.n2225 9.3005
R5421 vdd.n2227 vdd.n1532 9.3005
R5422 vdd.n2229 vdd.n2228 9.3005
R5423 vdd.n1522 vdd.n1521 9.3005
R5424 vdd.n2243 vdd.n2242 9.3005
R5425 vdd.n2244 vdd.n1520 9.3005
R5426 vdd.n2246 vdd.n2245 9.3005
R5427 vdd.n1512 vdd.n1511 9.3005
R5428 vdd.n2260 vdd.n2259 9.3005
R5429 vdd.n2261 vdd.n1509 9.3005
R5430 vdd.n2265 vdd.n2264 9.3005
R5431 vdd.n2263 vdd.n1510 9.3005
R5432 vdd.n2262 vdd.n1499 9.3005
R5433 vdd.n1833 vdd.n1601 9.3005
R5434 vdd.n1726 vdd.n1602 9.3005
R5435 vdd.n1728 vdd.n1727 9.3005
R5436 vdd.n1729 vdd.n1721 9.3005
R5437 vdd.n1731 vdd.n1730 9.3005
R5438 vdd.n1732 vdd.n1720 9.3005
R5439 vdd.n1734 vdd.n1733 9.3005
R5440 vdd.n1735 vdd.n1715 9.3005
R5441 vdd.n1737 vdd.n1736 9.3005
R5442 vdd.n1738 vdd.n1714 9.3005
R5443 vdd.n1740 vdd.n1739 9.3005
R5444 vdd.n1741 vdd.n1709 9.3005
R5445 vdd.n1743 vdd.n1742 9.3005
R5446 vdd.n1744 vdd.n1708 9.3005
R5447 vdd.n1746 vdd.n1745 9.3005
R5448 vdd.n1747 vdd.n1703 9.3005
R5449 vdd.n1749 vdd.n1748 9.3005
R5450 vdd.n1750 vdd.n1702 9.3005
R5451 vdd.n1752 vdd.n1751 9.3005
R5452 vdd.n1753 vdd.n1697 9.3005
R5453 vdd.n1755 vdd.n1754 9.3005
R5454 vdd.n1756 vdd.n1696 9.3005
R5455 vdd.n1761 vdd.n1757 9.3005
R5456 vdd.n1762 vdd.n1692 9.3005
R5457 vdd.n1764 vdd.n1763 9.3005
R5458 vdd.n1765 vdd.n1691 9.3005
R5459 vdd.n1767 vdd.n1766 9.3005
R5460 vdd.n1768 vdd.n1686 9.3005
R5461 vdd.n1770 vdd.n1769 9.3005
R5462 vdd.n1771 vdd.n1685 9.3005
R5463 vdd.n1773 vdd.n1772 9.3005
R5464 vdd.n1774 vdd.n1680 9.3005
R5465 vdd.n1776 vdd.n1775 9.3005
R5466 vdd.n1777 vdd.n1679 9.3005
R5467 vdd.n1779 vdd.n1778 9.3005
R5468 vdd.n1780 vdd.n1674 9.3005
R5469 vdd.n1782 vdd.n1781 9.3005
R5470 vdd.n1783 vdd.n1673 9.3005
R5471 vdd.n1785 vdd.n1784 9.3005
R5472 vdd.n1786 vdd.n1668 9.3005
R5473 vdd.n1788 vdd.n1787 9.3005
R5474 vdd.n1789 vdd.n1667 9.3005
R5475 vdd.n1791 vdd.n1790 9.3005
R5476 vdd.n1792 vdd.n1664 9.3005
R5477 vdd.n1798 vdd.n1797 9.3005
R5478 vdd.n1799 vdd.n1663 9.3005
R5479 vdd.n1801 vdd.n1800 9.3005
R5480 vdd.n1802 vdd.n1658 9.3005
R5481 vdd.n1804 vdd.n1803 9.3005
R5482 vdd.n1805 vdd.n1657 9.3005
R5483 vdd.n1807 vdd.n1806 9.3005
R5484 vdd.n1808 vdd.n1652 9.3005
R5485 vdd.n1810 vdd.n1809 9.3005
R5486 vdd.n1811 vdd.n1651 9.3005
R5487 vdd.n1813 vdd.n1812 9.3005
R5488 vdd.n1814 vdd.n1646 9.3005
R5489 vdd.n1816 vdd.n1815 9.3005
R5490 vdd.n1817 vdd.n1645 9.3005
R5491 vdd.n1819 vdd.n1818 9.3005
R5492 vdd.n1820 vdd.n1641 9.3005
R5493 vdd.n1822 vdd.n1821 9.3005
R5494 vdd.n1823 vdd.n1640 9.3005
R5495 vdd.n1825 vdd.n1824 9.3005
R5496 vdd.n1826 vdd.n1639 9.3005
R5497 vdd.n1832 vdd.n1831 9.3005
R5498 vdd.n1840 vdd.n1839 9.3005
R5499 vdd.n1841 vdd.n1595 9.3005
R5500 vdd.n1843 vdd.n1842 9.3005
R5501 vdd.n1585 vdd.n1584 9.3005
R5502 vdd.n1857 vdd.n1856 9.3005
R5503 vdd.n1858 vdd.n1583 9.3005
R5504 vdd.n1860 vdd.n1859 9.3005
R5505 vdd.n1574 vdd.n1573 9.3005
R5506 vdd.n1874 vdd.n1873 9.3005
R5507 vdd.n1875 vdd.n1572 9.3005
R5508 vdd.n1877 vdd.n1876 9.3005
R5509 vdd.n1563 vdd.n1562 9.3005
R5510 vdd.n1890 vdd.n1889 9.3005
R5511 vdd.n1891 vdd.n1561 9.3005
R5512 vdd.n1893 vdd.n1892 9.3005
R5513 vdd.n1551 vdd.n1550 9.3005
R5514 vdd.n1907 vdd.n1906 9.3005
R5515 vdd.n1597 vdd.n1596 9.3005
R5516 vdd.n2119 vdd.n2118 9.3005
R5517 vdd.n2114 vdd.n2113 9.3005
R5518 vdd.n2125 vdd.n2124 9.3005
R5519 vdd.n2127 vdd.n2126 9.3005
R5520 vdd.n2110 vdd.n2109 9.3005
R5521 vdd.n2133 vdd.n2132 9.3005
R5522 vdd.n2135 vdd.n2134 9.3005
R5523 vdd.n2107 vdd.n2104 9.3005
R5524 vdd.n2142 vdd.n2141 9.3005
R5525 vdd.n2174 vdd.n2173 9.3005
R5526 vdd.n2169 vdd.n2168 9.3005
R5527 vdd.n2180 vdd.n2179 9.3005
R5528 vdd.n2182 vdd.n2181 9.3005
R5529 vdd.n2165 vdd.n2164 9.3005
R5530 vdd.n2188 vdd.n2187 9.3005
R5531 vdd.n2190 vdd.n2189 9.3005
R5532 vdd.n2162 vdd.n2159 9.3005
R5533 vdd.n2197 vdd.n2196 9.3005
R5534 vdd.n2021 vdd.n2020 9.3005
R5535 vdd.n2016 vdd.n2015 9.3005
R5536 vdd.n2027 vdd.n2026 9.3005
R5537 vdd.n2029 vdd.n2028 9.3005
R5538 vdd.n2012 vdd.n2011 9.3005
R5539 vdd.n2035 vdd.n2034 9.3005
R5540 vdd.n2037 vdd.n2036 9.3005
R5541 vdd.n2009 vdd.n2006 9.3005
R5542 vdd.n2044 vdd.n2043 9.3005
R5543 vdd.n2076 vdd.n2075 9.3005
R5544 vdd.n2071 vdd.n2070 9.3005
R5545 vdd.n2082 vdd.n2081 9.3005
R5546 vdd.n2084 vdd.n2083 9.3005
R5547 vdd.n2067 vdd.n2066 9.3005
R5548 vdd.n2090 vdd.n2089 9.3005
R5549 vdd.n2092 vdd.n2091 9.3005
R5550 vdd.n2064 vdd.n2061 9.3005
R5551 vdd.n2099 vdd.n2098 9.3005
R5552 vdd.n1924 vdd.n1923 9.3005
R5553 vdd.n1919 vdd.n1918 9.3005
R5554 vdd.n1930 vdd.n1929 9.3005
R5555 vdd.n1932 vdd.n1931 9.3005
R5556 vdd.n1915 vdd.n1914 9.3005
R5557 vdd.n1938 vdd.n1937 9.3005
R5558 vdd.n1940 vdd.n1939 9.3005
R5559 vdd.n1912 vdd.n1909 9.3005
R5560 vdd.n1947 vdd.n1946 9.3005
R5561 vdd.n1979 vdd.n1978 9.3005
R5562 vdd.n1974 vdd.n1973 9.3005
R5563 vdd.n1985 vdd.n1984 9.3005
R5564 vdd.n1987 vdd.n1986 9.3005
R5565 vdd.n1970 vdd.n1969 9.3005
R5566 vdd.n1993 vdd.n1992 9.3005
R5567 vdd.n1995 vdd.n1994 9.3005
R5568 vdd.n1967 vdd.n1964 9.3005
R5569 vdd.n2002 vdd.n2001 9.3005
R5570 vdd.n1853 vdd.t182 9.18308
R5571 vdd.n3508 vdd.t49 9.18308
R5572 vdd.n1879 vdd.t61 8.95635
R5573 vdd.t6 vdd.n3549 8.95635
R5574 vdd.n300 vdd.n299 8.92171
R5575 vdd.n245 vdd.n244 8.92171
R5576 vdd.n202 vdd.n201 8.92171
R5577 vdd.n147 vdd.n146 8.92171
R5578 vdd.n105 vdd.n104 8.92171
R5579 vdd.n50 vdd.n49 8.92171
R5580 vdd.n2124 vdd.n2123 8.92171
R5581 vdd.n2179 vdd.n2178 8.92171
R5582 vdd.n2026 vdd.n2025 8.92171
R5583 vdd.n2081 vdd.n2080 8.92171
R5584 vdd.n1929 vdd.n1928 8.92171
R5585 vdd.n1984 vdd.n1983 8.92171
R5586 vdd.n223 vdd.n125 8.81535
R5587 vdd.n2102 vdd.n2004 8.81535
R5588 vdd.n1559 vdd.t143 8.72962
R5589 vdd.t169 vdd.n3558 8.72962
R5590 vdd.n2215 vdd.t2 8.50289
R5591 vdd.n3477 vdd.t53 8.50289
R5592 vdd.n28 vdd.n14 8.42249
R5593 vdd.n2231 vdd.t31 8.27616
R5594 vdd.t33 vdd.n636 8.27616
R5595 vdd.n3564 vdd.n3563 8.16225
R5596 vdd.n2202 vdd.n2201 8.16225
R5597 vdd.n296 vdd.n290 8.14595
R5598 vdd.n241 vdd.n235 8.14595
R5599 vdd.n198 vdd.n192 8.14595
R5600 vdd.n143 vdd.n137 8.14595
R5601 vdd.n101 vdd.n95 8.14595
R5602 vdd.n46 vdd.n40 8.14595
R5603 vdd.n2120 vdd.n2114 8.14595
R5604 vdd.n2175 vdd.n2169 8.14595
R5605 vdd.n2022 vdd.n2016 8.14595
R5606 vdd.n2077 vdd.n2071 8.14595
R5607 vdd.n1925 vdd.n1919 8.14595
R5608 vdd.n1980 vdd.n1974 8.14595
R5609 vdd.t111 vdd.n1593 7.8227
R5610 vdd.t84 vdd.n363 7.8227
R5611 vdd.n2430 vdd.n1105 7.70933
R5612 vdd.n2430 vdd.n1108 7.70933
R5613 vdd.n2436 vdd.n1094 7.70933
R5614 vdd.n2442 vdd.n1094 7.70933
R5615 vdd.n2442 vdd.n1087 7.70933
R5616 vdd.n2448 vdd.n1087 7.70933
R5617 vdd.n2448 vdd.n1090 7.70933
R5618 vdd.n2454 vdd.n1083 7.70933
R5619 vdd.n2460 vdd.n1077 7.70933
R5620 vdd.n2466 vdd.n1064 7.70933
R5621 vdd.n2472 vdd.n1064 7.70933
R5622 vdd.n2478 vdd.n1058 7.70933
R5623 vdd.n2484 vdd.n1051 7.70933
R5624 vdd.n2484 vdd.n1054 7.70933
R5625 vdd.n2490 vdd.n1047 7.70933
R5626 vdd.n2497 vdd.n1033 7.70933
R5627 vdd.n2503 vdd.n1033 7.70933
R5628 vdd.n2509 vdd.n1027 7.70933
R5629 vdd.n2515 vdd.n1023 7.70933
R5630 vdd.n2521 vdd.n1017 7.70933
R5631 vdd.n2539 vdd.n999 7.70933
R5632 vdd.n2539 vdd.n992 7.70933
R5633 vdd.n2547 vdd.n992 7.70933
R5634 vdd.n2629 vdd.n976 7.70933
R5635 vdd.n3012 vdd.n928 7.70933
R5636 vdd.n3024 vdd.n917 7.70933
R5637 vdd.n3024 vdd.n911 7.70933
R5638 vdd.n3030 vdd.n911 7.70933
R5639 vdd.n3042 vdd.n902 7.70933
R5640 vdd.n3048 vdd.n896 7.70933
R5641 vdd.n3060 vdd.n883 7.70933
R5642 vdd.n3067 vdd.n876 7.70933
R5643 vdd.n3067 vdd.n879 7.70933
R5644 vdd.n3073 vdd.n872 7.70933
R5645 vdd.n3079 vdd.n858 7.70933
R5646 vdd.n3085 vdd.n858 7.70933
R5647 vdd.n3091 vdd.n852 7.70933
R5648 vdd.n3097 vdd.n845 7.70933
R5649 vdd.n3097 vdd.n848 7.70933
R5650 vdd.n3103 vdd.n841 7.70933
R5651 vdd.n3109 vdd.n835 7.70933
R5652 vdd.n3115 vdd.n822 7.70933
R5653 vdd.n3121 vdd.n822 7.70933
R5654 vdd.n3121 vdd.n814 7.70933
R5655 vdd.n3172 vdd.n814 7.70933
R5656 vdd.n3172 vdd.n817 7.70933
R5657 vdd.n3178 vdd.n774 7.70933
R5658 vdd.n3248 vdd.n774 7.70933
R5659 vdd.n295 vdd.n292 7.3702
R5660 vdd.n240 vdd.n237 7.3702
R5661 vdd.n197 vdd.n194 7.3702
R5662 vdd.n142 vdd.n139 7.3702
R5663 vdd.n100 vdd.n97 7.3702
R5664 vdd.n45 vdd.n42 7.3702
R5665 vdd.n2119 vdd.n2116 7.3702
R5666 vdd.n2174 vdd.n2171 7.3702
R5667 vdd.n2021 vdd.n2018 7.3702
R5668 vdd.n2076 vdd.n2073 7.3702
R5669 vdd.n1924 vdd.n1921 7.3702
R5670 vdd.n1979 vdd.n1976 7.3702
R5671 vdd.n1077 vdd.t247 7.36923
R5672 vdd.n3103 vdd.t224 7.36923
R5673 vdd.n2454 vdd.t199 7.1425
R5674 vdd.n1396 vdd.t195 7.1425
R5675 vdd.n3036 vdd.t198 7.1425
R5676 vdd.n835 vdd.t208 7.1425
R5677 vdd.n1762 vdd.n1761 6.98232
R5678 vdd.n2318 vdd.n2317 6.98232
R5679 vdd.n547 vdd.n546 6.98232
R5680 vdd.n3332 vdd.n3331 6.98232
R5681 vdd.n2249 vdd.t4 6.91577
R5682 vdd.n3441 vdd.t63 6.91577
R5683 vdd.n1396 vdd.t196 6.80241
R5684 vdd.n3036 vdd.t240 6.80241
R5685 vdd.t37 vdd.n1530 6.68904
R5686 vdd.n3457 vdd.t171 6.68904
R5687 vdd.n2207 vdd.t23 6.46231
R5688 vdd.n2478 vdd.t206 6.46231
R5689 vdd.t211 vdd.n1027 6.46231
R5690 vdd.n3060 vdd.t216 6.46231
R5691 vdd.t232 vdd.n852 6.46231
R5692 vdd.n3485 vdd.t152 6.46231
R5693 vdd.n2554 vdd.t244 6.34895
R5694 vdd.n2933 vdd.t229 6.34895
R5695 vdd.n3564 vdd.n321 6.32949
R5696 vdd.n2201 vdd.n2200 6.32949
R5697 vdd.n3075 vdd.n868 6.2444
R5698 vdd.n2494 vdd.n2493 6.2444
R5699 vdd.t17 vdd.n1558 6.23558
R5700 vdd.t146 vdd.n332 6.23558
R5701 vdd.n1871 vdd.t180 6.00885
R5702 vdd.n3543 vdd.t29 6.00885
R5703 vdd.n2515 vdd.t237 5.89549
R5704 vdd.n896 vdd.t212 5.89549
R5705 vdd.n296 vdd.n295 5.81868
R5706 vdd.n241 vdd.n240 5.81868
R5707 vdd.n198 vdd.n197 5.81868
R5708 vdd.n143 vdd.n142 5.81868
R5709 vdd.n101 vdd.n100 5.81868
R5710 vdd.n46 vdd.n45 5.81868
R5711 vdd.n2120 vdd.n2119 5.81868
R5712 vdd.n2175 vdd.n2174 5.81868
R5713 vdd.n2022 vdd.n2021 5.81868
R5714 vdd.n2077 vdd.n2076 5.81868
R5715 vdd.n1925 vdd.n1924 5.81868
R5716 vdd.n1980 vdd.n1979 5.81868
R5717 vdd.n2637 vdd.n2636 5.77611
R5718 vdd.n1320 vdd.n1319 5.77611
R5719 vdd.n2945 vdd.n2944 5.77611
R5720 vdd.n3187 vdd.n806 5.77611
R5721 vdd.n3253 vdd.n770 5.77611
R5722 vdd.n2808 vdd.n2742 5.77611
R5723 vdd.n2562 vdd.n983 5.77611
R5724 vdd.n1456 vdd.n1288 5.77611
R5725 vdd.n1831 vdd.n1605 5.62474
R5726 vdd.n2281 vdd.n2278 5.62474
R5727 vdd.n3522 vdd.n407 5.62474
R5728 vdd.n3287 vdd.n3284 5.62474
R5729 vdd.n2490 vdd.t226 5.55539
R5730 vdd.n872 vdd.t202 5.55539
R5731 vdd.n1581 vdd.t180 5.32866
R5732 vdd.t29 vdd.n3542 5.32866
R5733 vdd.n1887 vdd.t17 5.10193
R5734 vdd.n3551 vdd.t146 5.10193
R5735 vdd.n299 vdd.n290 5.04292
R5736 vdd.n244 vdd.n235 5.04292
R5737 vdd.n201 vdd.n192 5.04292
R5738 vdd.n146 vdd.n137 5.04292
R5739 vdd.n104 vdd.n95 5.04292
R5740 vdd.n49 vdd.n40 5.04292
R5741 vdd.n2123 vdd.n2114 5.04292
R5742 vdd.n2178 vdd.n2169 5.04292
R5743 vdd.n2025 vdd.n2016 5.04292
R5744 vdd.n2080 vdd.n2071 5.04292
R5745 vdd.n1928 vdd.n1919 5.04292
R5746 vdd.n1983 vdd.n1974 5.04292
R5747 vdd.n1903 vdd.t23 4.8752
R5748 vdd.t205 vdd.t217 4.8752
R5749 vdd.t248 vdd.t194 4.8752
R5750 vdd.t152 vdd.n328 4.8752
R5751 vdd.n2638 vdd.n2637 4.83952
R5752 vdd.n1319 vdd.n1318 4.83952
R5753 vdd.n2946 vdd.n2945 4.83952
R5754 vdd.n806 vdd.n801 4.83952
R5755 vdd.n770 vdd.n765 4.83952
R5756 vdd.n2805 vdd.n2742 4.83952
R5757 vdd.n2565 vdd.n983 4.83952
R5758 vdd.n1459 vdd.n1288 4.83952
R5759 vdd.n1370 vdd.t214 4.76184
R5760 vdd.n3018 vdd.t200 4.76184
R5761 vdd.n2286 vdd.n2285 4.74817
R5762 vdd.n1492 vdd.n1487 4.74817
R5763 vdd.n1154 vdd.n1151 4.74817
R5764 vdd.n2379 vdd.n1150 4.74817
R5765 vdd.n2384 vdd.n1151 4.74817
R5766 vdd.n2383 vdd.n1150 4.74817
R5767 vdd.n664 vdd.n662 4.74817
R5768 vdd.n3402 vdd.n665 4.74817
R5769 vdd.n3405 vdd.n665 4.74817
R5770 vdd.n3406 vdd.n664 4.74817
R5771 vdd.n3294 vdd.n749 4.74817
R5772 vdd.n3290 vdd.n751 4.74817
R5773 vdd.n3293 vdd.n751 4.74817
R5774 vdd.n3298 vdd.n749 4.74817
R5775 vdd.n2285 vdd.n1250 4.74817
R5776 vdd.n1489 vdd.n1487 4.74817
R5777 vdd.n321 vdd.n320 4.7074
R5778 vdd.n223 vdd.n222 4.7074
R5779 vdd.n2200 vdd.n2199 4.7074
R5780 vdd.n2102 vdd.n2101 4.7074
R5781 vdd.n2223 vdd.t37 4.64847
R5782 vdd.t207 vdd.n1058 4.64847
R5783 vdd.n2509 vdd.t246 4.64847
R5784 vdd.t235 vdd.n883 4.64847
R5785 vdd.n3091 vdd.t231 4.64847
R5786 vdd.n3466 vdd.t171 4.64847
R5787 vdd.n1047 vdd.t129 4.53511
R5788 vdd.n3073 vdd.t92 4.53511
R5789 vdd.n1524 vdd.t4 4.42174
R5790 vdd.n2436 vdd.t70 4.42174
R5791 vdd.n1370 vdd.t115 4.42174
R5792 vdd.n3018 vdd.t122 4.42174
R5793 vdd.n817 vdd.t66 4.42174
R5794 vdd.t63 vdd.n635 4.42174
R5795 vdd.n3064 vdd.n868 4.37123
R5796 vdd.n2495 vdd.n2494 4.37123
R5797 vdd.n2533 vdd.t233 4.30838
R5798 vdd.n2921 vdd.t220 4.30838
R5799 vdd.n300 vdd.n288 4.26717
R5800 vdd.n245 vdd.n233 4.26717
R5801 vdd.n202 vdd.n190 4.26717
R5802 vdd.n147 vdd.n135 4.26717
R5803 vdd.n105 vdd.n93 4.26717
R5804 vdd.n50 vdd.n38 4.26717
R5805 vdd.n2124 vdd.n2112 4.26717
R5806 vdd.n2179 vdd.n2167 4.26717
R5807 vdd.n2026 vdd.n2014 4.26717
R5808 vdd.n2081 vdd.n2069 4.26717
R5809 vdd.n1929 vdd.n1917 4.26717
R5810 vdd.n1984 vdd.n1972 4.26717
R5811 vdd.n321 vdd.n223 4.10845
R5812 vdd.n2200 vdd.n2102 4.10845
R5813 vdd.n277 vdd.t30 4.06363
R5814 vdd.n277 vdd.t50 4.06363
R5815 vdd.n275 vdd.t149 4.06363
R5816 vdd.n275 vdd.t44 4.06363
R5817 vdd.n273 vdd.t250 4.06363
R5818 vdd.n273 vdd.t264 4.06363
R5819 vdd.n271 vdd.t155 4.06363
R5820 vdd.n271 vdd.t261 4.06363
R5821 vdd.n269 vdd.t275 4.06363
R5822 vdd.n269 vdd.t159 4.06363
R5823 vdd.n267 vdd.t35 4.06363
R5824 vdd.n267 vdd.t172 4.06363
R5825 vdd.n265 vdd.t259 4.06363
R5826 vdd.n265 vdd.t263 4.06363
R5827 vdd.n179 vdd.t188 4.06363
R5828 vdd.n179 vdd.t272 4.06363
R5829 vdd.n177 vdd.t7 4.06363
R5830 vdd.n177 vdd.t262 4.06363
R5831 vdd.n175 vdd.t39 4.06363
R5832 vdd.n175 vdd.t154 4.06363
R5833 vdd.n173 vdd.t153 4.06363
R5834 vdd.n173 vdd.t170 4.06363
R5835 vdd.n171 vdd.t150 4.06363
R5836 vdd.n171 vdd.t142 4.06363
R5837 vdd.n169 vdd.t271 4.06363
R5838 vdd.n169 vdd.t179 4.06363
R5839 vdd.n167 vdd.t267 4.06363
R5840 vdd.n167 vdd.t42 4.06363
R5841 vdd.n82 vdd.t255 4.06363
R5842 vdd.n82 vdd.t258 4.06363
R5843 vdd.n80 vdd.t269 4.06363
R5844 vdd.n80 vdd.t163 4.06363
R5845 vdd.n78 vdd.t1 4.06363
R5846 vdd.n78 vdd.t147 4.06363
R5847 vdd.n76 vdd.t164 4.06363
R5848 vdd.n76 vdd.t191 4.06363
R5849 vdd.n74 vdd.t54 4.06363
R5850 vdd.n74 vdd.t156 4.06363
R5851 vdd.n72 vdd.t22 4.06363
R5852 vdd.n72 vdd.t252 4.06363
R5853 vdd.n70 vdd.t64 4.06363
R5854 vdd.n70 vdd.t34 4.06363
R5855 vdd.n2144 vdd.t32 4.06363
R5856 vdd.n2144 vdd.t46 4.06363
R5857 vdd.n2146 vdd.t38 4.06363
R5858 vdd.n2146 vdd.t55 4.06363
R5859 vdd.n2148 vdd.t25 4.06363
R5860 vdd.n2148 vdd.t167 4.06363
R5861 vdd.n2150 vdd.t144 4.06363
R5862 vdd.n2150 vdd.t24 4.06363
R5863 vdd.n2152 vdd.t41 4.06363
R5864 vdd.n2152 vdd.t265 4.06363
R5865 vdd.n2154 vdd.t270 4.06363
R5866 vdd.n2154 vdd.t251 4.06363
R5867 vdd.n2156 vdd.t186 4.06363
R5868 vdd.n2156 vdd.t181 4.06363
R5869 vdd.n2046 vdd.t176 4.06363
R5870 vdd.n2046 vdd.t26 4.06363
R5871 vdd.n2048 vdd.t274 4.06363
R5872 vdd.n2048 vdd.t151 4.06363
R5873 vdd.n2050 vdd.t16 4.06363
R5874 vdd.n2050 vdd.t3 4.06363
R5875 vdd.n2052 vdd.t187 4.06363
R5876 vdd.n2052 vdd.t260 4.06363
R5877 vdd.n2054 vdd.t18 4.06363
R5878 vdd.n2054 vdd.t256 4.06363
R5879 vdd.n2056 vdd.t253 4.06363
R5880 vdd.n2056 vdd.t268 4.06363
R5881 vdd.n2058 vdd.t184 4.06363
R5882 vdd.n2058 vdd.t266 4.06363
R5883 vdd.n1949 vdd.t178 4.06363
R5884 vdd.n1949 vdd.t5 4.06363
R5885 vdd.n1951 vdd.t257 4.06363
R5886 vdd.n1951 vdd.t20 4.06363
R5887 vdd.n1953 vdd.t189 4.06363
R5888 vdd.n1953 vdd.t58 4.06363
R5889 vdd.n1955 vdd.t190 4.06363
R5890 vdd.n1955 vdd.t45 4.06363
R5891 vdd.n1957 vdd.t145 4.06363
R5892 vdd.n1957 vdd.t28 4.06363
R5893 vdd.n1959 vdd.t162 4.06363
R5894 vdd.n1959 vdd.t62 4.06363
R5895 vdd.n1961 vdd.t183 4.06363
R5896 vdd.n1961 vdd.t254 4.06363
R5897 vdd.n1083 vdd.t239 3.96828
R5898 vdd.n2527 vdd.t219 3.96828
R5899 vdd.n2915 vdd.t236 3.96828
R5900 vdd.n3109 vdd.t225 3.96828
R5901 vdd.n26 vdd.t40 3.9605
R5902 vdd.n26 vdd.t36 3.9605
R5903 vdd.n23 vdd.t59 3.9605
R5904 vdd.n23 vdd.t12 3.9605
R5905 vdd.n21 vdd.t11 3.9605
R5906 vdd.n21 vdd.t173 3.9605
R5907 vdd.n20 vdd.t192 3.9605
R5908 vdd.n20 vdd.t13 3.9605
R5909 vdd.n15 vdd.t14 3.9605
R5910 vdd.n15 vdd.t193 3.9605
R5911 vdd.n16 vdd.t60 3.9605
R5912 vdd.n16 vdd.t10 3.9605
R5913 vdd.n18 vdd.t8 3.9605
R5914 vdd.n18 vdd.t157 3.9605
R5915 vdd.n25 vdd.t9 3.9605
R5916 vdd.n25 vdd.t158 3.9605
R5917 vdd.n2460 vdd.t239 3.74155
R5918 vdd.n1017 vdd.t219 3.74155
R5919 vdd.n3042 vdd.t236 3.74155
R5920 vdd.n841 vdd.t225 3.74155
R5921 vdd.n7 vdd.t249 3.61217
R5922 vdd.n7 vdd.t213 3.61217
R5923 vdd.n8 vdd.t221 3.61217
R5924 vdd.n8 vdd.t241 3.61217
R5925 vdd.n10 vdd.t230 3.61217
R5926 vdd.n10 vdd.t201 3.61217
R5927 vdd.n12 vdd.t210 3.61217
R5928 vdd.n12 vdd.t228 3.61217
R5929 vdd.n5 vdd.t243 3.61217
R5930 vdd.n5 vdd.t223 3.61217
R5931 vdd.n3 vdd.t215 3.61217
R5932 vdd.n3 vdd.t245 3.61217
R5933 vdd.n1 vdd.t197 3.61217
R5934 vdd.n1 vdd.t234 3.61217
R5935 vdd.n0 vdd.t238 3.61217
R5936 vdd.n0 vdd.t218 3.61217
R5937 vdd.n1837 vdd.t111 3.51482
R5938 vdd.n3527 vdd.t84 3.51482
R5939 vdd.n304 vdd.n303 3.49141
R5940 vdd.n249 vdd.n248 3.49141
R5941 vdd.n206 vdd.n205 3.49141
R5942 vdd.n151 vdd.n150 3.49141
R5943 vdd.n109 vdd.n108 3.49141
R5944 vdd.n54 vdd.n53 3.49141
R5945 vdd.n2128 vdd.n2127 3.49141
R5946 vdd.n2183 vdd.n2182 3.49141
R5947 vdd.n2030 vdd.n2029 3.49141
R5948 vdd.n2085 vdd.n2084 3.49141
R5949 vdd.n1933 vdd.n1932 3.49141
R5950 vdd.n1988 vdd.n1987 3.49141
R5951 vdd.t233 vdd.n999 3.40145
R5952 vdd.n2701 vdd.t242 3.40145
R5953 vdd.n3005 vdd.t227 3.40145
R5954 vdd.n3030 vdd.t220 3.40145
R5955 vdd.n1108 vdd.t70 3.28809
R5956 vdd.n2554 vdd.t115 3.28809
R5957 vdd.n2933 vdd.t122 3.28809
R5958 vdd.n3178 vdd.t66 3.28809
R5959 vdd.n2240 vdd.t31 3.06136
R5960 vdd.n2472 vdd.t207 3.06136
R5961 vdd.n1408 vdd.t246 3.06136
R5962 vdd.n3054 vdd.t235 3.06136
R5963 vdd.t231 vdd.n845 3.06136
R5964 vdd.n3449 vdd.t33 3.06136
R5965 vdd.n2547 vdd.t214 2.94799
R5966 vdd.t200 vdd.n917 2.94799
R5967 vdd.t2 vdd.n1536 2.83463
R5968 vdd.n624 vdd.t53 2.83463
R5969 vdd.n307 vdd.n286 2.71565
R5970 vdd.n252 vdd.n231 2.71565
R5971 vdd.n209 vdd.n188 2.71565
R5972 vdd.n154 vdd.n133 2.71565
R5973 vdd.n112 vdd.n91 2.71565
R5974 vdd.n57 vdd.n36 2.71565
R5975 vdd.n2131 vdd.n2110 2.71565
R5976 vdd.n2186 vdd.n2165 2.71565
R5977 vdd.n2033 vdd.n2012 2.71565
R5978 vdd.n2088 vdd.n2067 2.71565
R5979 vdd.n1936 vdd.n1915 2.71565
R5980 vdd.n1991 vdd.n1970 2.71565
R5981 vdd.n1904 vdd.t143 2.6079
R5982 vdd.n3559 vdd.t169 2.6079
R5983 vdd.n2521 vdd.t217 2.49453
R5984 vdd.n902 vdd.t248 2.49453
R5985 vdd.n294 vdd.n293 2.4129
R5986 vdd.n239 vdd.n238 2.4129
R5987 vdd.n196 vdd.n195 2.4129
R5988 vdd.n141 vdd.n140 2.4129
R5989 vdd.n99 vdd.n98 2.4129
R5990 vdd.n44 vdd.n43 2.4129
R5991 vdd.n2118 vdd.n2117 2.4129
R5992 vdd.n2173 vdd.n2172 2.4129
R5993 vdd.n2020 vdd.n2019 2.4129
R5994 vdd.n2075 vdd.n2074 2.4129
R5995 vdd.n1923 vdd.n1922 2.4129
R5996 vdd.n1978 vdd.n1977 2.4129
R5997 vdd.t61 vdd.n1565 2.38117
R5998 vdd.n3550 vdd.t6 2.38117
R5999 vdd.n2391 vdd.n1151 2.27742
R6000 vdd.n2391 vdd.n1150 2.27742
R6001 vdd.n3214 vdd.n665 2.27742
R6002 vdd.n3214 vdd.n664 2.27742
R6003 vdd.n3282 vdd.n751 2.27742
R6004 vdd.n3282 vdd.n749 2.27742
R6005 vdd.n2285 vdd.n2284 2.27742
R6006 vdd.n2284 vdd.n1487 2.27742
R6007 vdd.n1862 vdd.t182 2.15444
R6008 vdd.n1054 vdd.t226 2.15444
R6009 vdd.n2497 vdd.t204 2.15444
R6010 vdd.n879 vdd.t203 2.15444
R6011 vdd.n3079 vdd.t202 2.15444
R6012 vdd.n3541 vdd.t49 2.15444
R6013 vdd.n308 vdd.n284 1.93989
R6014 vdd.n253 vdd.n229 1.93989
R6015 vdd.n210 vdd.n186 1.93989
R6016 vdd.n155 vdd.n131 1.93989
R6017 vdd.n113 vdd.n89 1.93989
R6018 vdd.n58 vdd.n34 1.93989
R6019 vdd.n2132 vdd.n2108 1.93989
R6020 vdd.n2187 vdd.n2163 1.93989
R6021 vdd.n2034 vdd.n2010 1.93989
R6022 vdd.n2089 vdd.n2065 1.93989
R6023 vdd.n1937 vdd.n1913 1.93989
R6024 vdd.n1992 vdd.n1968 1.93989
R6025 vdd.n1408 vdd.t237 1.81434
R6026 vdd.n3054 vdd.t212 1.81434
R6027 vdd.n1854 vdd.t47 1.70098
R6028 vdd.n3535 vdd.t56 1.70098
R6029 vdd.n1870 vdd.t161 1.47425
R6030 vdd.n349 vdd.t43 1.47425
R6031 vdd.t244 vdd.n976 1.36088
R6032 vdd.n3012 vdd.t229 1.36088
R6033 vdd.n1895 vdd.t27 1.24752
R6034 vdd.t74 vdd.n1500 1.24752
R6035 vdd.t206 vdd.n1051 1.24752
R6036 vdd.n2503 vdd.t211 1.24752
R6037 vdd.t216 vdd.n876 1.24752
R6038 vdd.n3085 vdd.t232 1.24752
R6039 vdd.n659 vdd.t88 1.24752
R6040 vdd.t0 vdd.n3557 1.24752
R6041 vdd.n2201 vdd.n28 1.16438
R6042 vdd.n319 vdd.n279 1.16414
R6043 vdd.n312 vdd.n311 1.16414
R6044 vdd.n264 vdd.n224 1.16414
R6045 vdd.n257 vdd.n256 1.16414
R6046 vdd.n221 vdd.n181 1.16414
R6047 vdd.n214 vdd.n213 1.16414
R6048 vdd.n166 vdd.n126 1.16414
R6049 vdd.n159 vdd.n158 1.16414
R6050 vdd.n124 vdd.n84 1.16414
R6051 vdd.n117 vdd.n116 1.16414
R6052 vdd.n69 vdd.n29 1.16414
R6053 vdd.n62 vdd.n61 1.16414
R6054 vdd.n2143 vdd.n2103 1.16414
R6055 vdd.n2136 vdd.n2135 1.16414
R6056 vdd.n2198 vdd.n2158 1.16414
R6057 vdd.n2191 vdd.n2190 1.16414
R6058 vdd.n2045 vdd.n2005 1.16414
R6059 vdd.n2038 vdd.n2037 1.16414
R6060 vdd.n2100 vdd.n2060 1.16414
R6061 vdd.n2093 vdd.n2092 1.16414
R6062 vdd.n1948 vdd.n1908 1.16414
R6063 vdd.n1941 vdd.n1940 1.16414
R6064 vdd.n2003 vdd.n1963 1.16414
R6065 vdd.n1996 vdd.n1995 1.16414
R6066 vdd vdd.n3564 1.15654
R6067 vdd.n1547 vdd.t15 1.02079
R6068 vdd.t129 vdd.t204 1.02079
R6069 vdd.t203 vdd.t92 1.02079
R6070 vdd.t141 vdd.n613 1.02079
R6071 vdd.n1726 vdd.n1605 0.970197
R6072 vdd.n2282 vdd.n2281 0.970197
R6073 vdd.n599 vdd.n407 0.970197
R6074 vdd.n3289 vdd.n3287 0.970197
R6075 vdd.n2527 vdd.t196 0.907421
R6076 vdd.n2915 vdd.t240 0.907421
R6077 vdd.n2232 vdd.t19 0.794056
R6078 vdd.n3458 vdd.t21 0.794056
R6079 vdd.n2248 vdd.t165 0.567326
R6080 vdd.n1090 vdd.t199 0.567326
R6081 vdd.n2533 vdd.t195 0.567326
R6082 vdd.n2921 vdd.t198 0.567326
R6083 vdd.n3115 vdd.t208 0.567326
R6084 vdd.t51 vdd.n642 0.567326
R6085 vdd.n2272 vdd.n1152 0.482207
R6086 vdd.n3414 vdd.n3413 0.482207
R6087 vdd.n444 vdd.n443 0.482207
R6088 vdd.n3521 vdd.n3520 0.482207
R6089 vdd.n3420 vdd.n656 0.482207
R6090 vdd.n2262 vdd.n1488 0.482207
R6091 vdd.n1833 vdd.n1832 0.482207
R6092 vdd.n1639 vdd.n1596 0.482207
R6093 vdd.n4 vdd.n2 0.459552
R6094 vdd.n11 vdd.n9 0.459552
R6095 vdd.n317 vdd.n316 0.388379
R6096 vdd.n283 vdd.n281 0.388379
R6097 vdd.n262 vdd.n261 0.388379
R6098 vdd.n228 vdd.n226 0.388379
R6099 vdd.n219 vdd.n218 0.388379
R6100 vdd.n185 vdd.n183 0.388379
R6101 vdd.n164 vdd.n163 0.388379
R6102 vdd.n130 vdd.n128 0.388379
R6103 vdd.n122 vdd.n121 0.388379
R6104 vdd.n88 vdd.n86 0.388379
R6105 vdd.n67 vdd.n66 0.388379
R6106 vdd.n33 vdd.n31 0.388379
R6107 vdd.n2141 vdd.n2140 0.388379
R6108 vdd.n2107 vdd.n2105 0.388379
R6109 vdd.n2196 vdd.n2195 0.388379
R6110 vdd.n2162 vdd.n2160 0.388379
R6111 vdd.n2043 vdd.n2042 0.388379
R6112 vdd.n2009 vdd.n2007 0.388379
R6113 vdd.n2098 vdd.n2097 0.388379
R6114 vdd.n2064 vdd.n2062 0.388379
R6115 vdd.n1946 vdd.n1945 0.388379
R6116 vdd.n1912 vdd.n1910 0.388379
R6117 vdd.n2001 vdd.n2000 0.388379
R6118 vdd.n1967 vdd.n1965 0.388379
R6119 vdd.n19 vdd.n17 0.387128
R6120 vdd.n24 vdd.n22 0.387128
R6121 vdd.n6 vdd.n4 0.358259
R6122 vdd.n13 vdd.n11 0.358259
R6123 vdd.n268 vdd.n266 0.358259
R6124 vdd.n270 vdd.n268 0.358259
R6125 vdd.n272 vdd.n270 0.358259
R6126 vdd.n274 vdd.n272 0.358259
R6127 vdd.n276 vdd.n274 0.358259
R6128 vdd.n278 vdd.n276 0.358259
R6129 vdd.n320 vdd.n278 0.358259
R6130 vdd.n170 vdd.n168 0.358259
R6131 vdd.n172 vdd.n170 0.358259
R6132 vdd.n174 vdd.n172 0.358259
R6133 vdd.n176 vdd.n174 0.358259
R6134 vdd.n178 vdd.n176 0.358259
R6135 vdd.n180 vdd.n178 0.358259
R6136 vdd.n222 vdd.n180 0.358259
R6137 vdd.n73 vdd.n71 0.358259
R6138 vdd.n75 vdd.n73 0.358259
R6139 vdd.n77 vdd.n75 0.358259
R6140 vdd.n79 vdd.n77 0.358259
R6141 vdd.n81 vdd.n79 0.358259
R6142 vdd.n83 vdd.n81 0.358259
R6143 vdd.n125 vdd.n83 0.358259
R6144 vdd.n2199 vdd.n2157 0.358259
R6145 vdd.n2157 vdd.n2155 0.358259
R6146 vdd.n2155 vdd.n2153 0.358259
R6147 vdd.n2153 vdd.n2151 0.358259
R6148 vdd.n2151 vdd.n2149 0.358259
R6149 vdd.n2149 vdd.n2147 0.358259
R6150 vdd.n2147 vdd.n2145 0.358259
R6151 vdd.n2101 vdd.n2059 0.358259
R6152 vdd.n2059 vdd.n2057 0.358259
R6153 vdd.n2057 vdd.n2055 0.358259
R6154 vdd.n2055 vdd.n2053 0.358259
R6155 vdd.n2053 vdd.n2051 0.358259
R6156 vdd.n2051 vdd.n2049 0.358259
R6157 vdd.n2049 vdd.n2047 0.358259
R6158 vdd.n2004 vdd.n1962 0.358259
R6159 vdd.n1962 vdd.n1960 0.358259
R6160 vdd.n1960 vdd.n1958 0.358259
R6161 vdd.n1958 vdd.n1956 0.358259
R6162 vdd.n1956 vdd.n1954 0.358259
R6163 vdd.n1954 vdd.n1952 0.358259
R6164 vdd.n1952 vdd.n1950 0.358259
R6165 vdd.n2466 vdd.t247 0.340595
R6166 vdd.n1023 vdd.t205 0.340595
R6167 vdd.n3048 vdd.t194 0.340595
R6168 vdd.n848 vdd.t224 0.340595
R6169 vdd.n14 vdd.n6 0.334552
R6170 vdd.n14 vdd.n13 0.334552
R6171 vdd.n27 vdd.n19 0.21707
R6172 vdd.n27 vdd.n24 0.21707
R6173 vdd.n318 vdd.n280 0.155672
R6174 vdd.n310 vdd.n280 0.155672
R6175 vdd.n310 vdd.n309 0.155672
R6176 vdd.n309 vdd.n285 0.155672
R6177 vdd.n302 vdd.n285 0.155672
R6178 vdd.n302 vdd.n301 0.155672
R6179 vdd.n301 vdd.n289 0.155672
R6180 vdd.n294 vdd.n289 0.155672
R6181 vdd.n263 vdd.n225 0.155672
R6182 vdd.n255 vdd.n225 0.155672
R6183 vdd.n255 vdd.n254 0.155672
R6184 vdd.n254 vdd.n230 0.155672
R6185 vdd.n247 vdd.n230 0.155672
R6186 vdd.n247 vdd.n246 0.155672
R6187 vdd.n246 vdd.n234 0.155672
R6188 vdd.n239 vdd.n234 0.155672
R6189 vdd.n220 vdd.n182 0.155672
R6190 vdd.n212 vdd.n182 0.155672
R6191 vdd.n212 vdd.n211 0.155672
R6192 vdd.n211 vdd.n187 0.155672
R6193 vdd.n204 vdd.n187 0.155672
R6194 vdd.n204 vdd.n203 0.155672
R6195 vdd.n203 vdd.n191 0.155672
R6196 vdd.n196 vdd.n191 0.155672
R6197 vdd.n165 vdd.n127 0.155672
R6198 vdd.n157 vdd.n127 0.155672
R6199 vdd.n157 vdd.n156 0.155672
R6200 vdd.n156 vdd.n132 0.155672
R6201 vdd.n149 vdd.n132 0.155672
R6202 vdd.n149 vdd.n148 0.155672
R6203 vdd.n148 vdd.n136 0.155672
R6204 vdd.n141 vdd.n136 0.155672
R6205 vdd.n123 vdd.n85 0.155672
R6206 vdd.n115 vdd.n85 0.155672
R6207 vdd.n115 vdd.n114 0.155672
R6208 vdd.n114 vdd.n90 0.155672
R6209 vdd.n107 vdd.n90 0.155672
R6210 vdd.n107 vdd.n106 0.155672
R6211 vdd.n106 vdd.n94 0.155672
R6212 vdd.n99 vdd.n94 0.155672
R6213 vdd.n68 vdd.n30 0.155672
R6214 vdd.n60 vdd.n30 0.155672
R6215 vdd.n60 vdd.n59 0.155672
R6216 vdd.n59 vdd.n35 0.155672
R6217 vdd.n52 vdd.n35 0.155672
R6218 vdd.n52 vdd.n51 0.155672
R6219 vdd.n51 vdd.n39 0.155672
R6220 vdd.n44 vdd.n39 0.155672
R6221 vdd.n2142 vdd.n2104 0.155672
R6222 vdd.n2134 vdd.n2104 0.155672
R6223 vdd.n2134 vdd.n2133 0.155672
R6224 vdd.n2133 vdd.n2109 0.155672
R6225 vdd.n2126 vdd.n2109 0.155672
R6226 vdd.n2126 vdd.n2125 0.155672
R6227 vdd.n2125 vdd.n2113 0.155672
R6228 vdd.n2118 vdd.n2113 0.155672
R6229 vdd.n2197 vdd.n2159 0.155672
R6230 vdd.n2189 vdd.n2159 0.155672
R6231 vdd.n2189 vdd.n2188 0.155672
R6232 vdd.n2188 vdd.n2164 0.155672
R6233 vdd.n2181 vdd.n2164 0.155672
R6234 vdd.n2181 vdd.n2180 0.155672
R6235 vdd.n2180 vdd.n2168 0.155672
R6236 vdd.n2173 vdd.n2168 0.155672
R6237 vdd.n2044 vdd.n2006 0.155672
R6238 vdd.n2036 vdd.n2006 0.155672
R6239 vdd.n2036 vdd.n2035 0.155672
R6240 vdd.n2035 vdd.n2011 0.155672
R6241 vdd.n2028 vdd.n2011 0.155672
R6242 vdd.n2028 vdd.n2027 0.155672
R6243 vdd.n2027 vdd.n2015 0.155672
R6244 vdd.n2020 vdd.n2015 0.155672
R6245 vdd.n2099 vdd.n2061 0.155672
R6246 vdd.n2091 vdd.n2061 0.155672
R6247 vdd.n2091 vdd.n2090 0.155672
R6248 vdd.n2090 vdd.n2066 0.155672
R6249 vdd.n2083 vdd.n2066 0.155672
R6250 vdd.n2083 vdd.n2082 0.155672
R6251 vdd.n2082 vdd.n2070 0.155672
R6252 vdd.n2075 vdd.n2070 0.155672
R6253 vdd.n1947 vdd.n1909 0.155672
R6254 vdd.n1939 vdd.n1909 0.155672
R6255 vdd.n1939 vdd.n1938 0.155672
R6256 vdd.n1938 vdd.n1914 0.155672
R6257 vdd.n1931 vdd.n1914 0.155672
R6258 vdd.n1931 vdd.n1930 0.155672
R6259 vdd.n1930 vdd.n1918 0.155672
R6260 vdd.n1923 vdd.n1918 0.155672
R6261 vdd.n2002 vdd.n1964 0.155672
R6262 vdd.n1994 vdd.n1964 0.155672
R6263 vdd.n1994 vdd.n1993 0.155672
R6264 vdd.n1993 vdd.n1969 0.155672
R6265 vdd.n1986 vdd.n1969 0.155672
R6266 vdd.n1986 vdd.n1985 0.155672
R6267 vdd.n1985 vdd.n1973 0.155672
R6268 vdd.n1978 vdd.n1973 0.155672
R6269 vdd.n1157 vdd.n1149 0.152939
R6270 vdd.n1161 vdd.n1157 0.152939
R6271 vdd.n1162 vdd.n1161 0.152939
R6272 vdd.n1163 vdd.n1162 0.152939
R6273 vdd.n1164 vdd.n1163 0.152939
R6274 vdd.n1168 vdd.n1164 0.152939
R6275 vdd.n1169 vdd.n1168 0.152939
R6276 vdd.n1170 vdd.n1169 0.152939
R6277 vdd.n1171 vdd.n1170 0.152939
R6278 vdd.n1175 vdd.n1171 0.152939
R6279 vdd.n1176 vdd.n1175 0.152939
R6280 vdd.n1177 vdd.n1176 0.152939
R6281 vdd.n2355 vdd.n1177 0.152939
R6282 vdd.n2355 vdd.n2354 0.152939
R6283 vdd.n2354 vdd.n2353 0.152939
R6284 vdd.n2353 vdd.n1183 0.152939
R6285 vdd.n1188 vdd.n1183 0.152939
R6286 vdd.n1189 vdd.n1188 0.152939
R6287 vdd.n1190 vdd.n1189 0.152939
R6288 vdd.n1194 vdd.n1190 0.152939
R6289 vdd.n1195 vdd.n1194 0.152939
R6290 vdd.n1196 vdd.n1195 0.152939
R6291 vdd.n1197 vdd.n1196 0.152939
R6292 vdd.n1201 vdd.n1197 0.152939
R6293 vdd.n1202 vdd.n1201 0.152939
R6294 vdd.n1203 vdd.n1202 0.152939
R6295 vdd.n1204 vdd.n1203 0.152939
R6296 vdd.n1208 vdd.n1204 0.152939
R6297 vdd.n1209 vdd.n1208 0.152939
R6298 vdd.n1210 vdd.n1209 0.152939
R6299 vdd.n1211 vdd.n1210 0.152939
R6300 vdd.n1215 vdd.n1211 0.152939
R6301 vdd.n1216 vdd.n1215 0.152939
R6302 vdd.n1217 vdd.n1216 0.152939
R6303 vdd.n2316 vdd.n1217 0.152939
R6304 vdd.n2316 vdd.n2315 0.152939
R6305 vdd.n2315 vdd.n2314 0.152939
R6306 vdd.n2314 vdd.n1223 0.152939
R6307 vdd.n1228 vdd.n1223 0.152939
R6308 vdd.n1229 vdd.n1228 0.152939
R6309 vdd.n1230 vdd.n1229 0.152939
R6310 vdd.n1234 vdd.n1230 0.152939
R6311 vdd.n1235 vdd.n1234 0.152939
R6312 vdd.n1236 vdd.n1235 0.152939
R6313 vdd.n1237 vdd.n1236 0.152939
R6314 vdd.n1241 vdd.n1237 0.152939
R6315 vdd.n1242 vdd.n1241 0.152939
R6316 vdd.n1243 vdd.n1242 0.152939
R6317 vdd.n1244 vdd.n1243 0.152939
R6318 vdd.n1248 vdd.n1244 0.152939
R6319 vdd.n1249 vdd.n1248 0.152939
R6320 vdd.n2390 vdd.n1152 0.152939
R6321 vdd.n2204 vdd.n2203 0.152939
R6322 vdd.n2204 vdd.n1539 0.152939
R6323 vdd.n2218 vdd.n1539 0.152939
R6324 vdd.n2219 vdd.n2218 0.152939
R6325 vdd.n2220 vdd.n2219 0.152939
R6326 vdd.n2220 vdd.n1527 0.152939
R6327 vdd.n2235 vdd.n1527 0.152939
R6328 vdd.n2236 vdd.n2235 0.152939
R6329 vdd.n2237 vdd.n2236 0.152939
R6330 vdd.n2237 vdd.n1516 0.152939
R6331 vdd.n2252 vdd.n1516 0.152939
R6332 vdd.n2253 vdd.n2252 0.152939
R6333 vdd.n2254 vdd.n2253 0.152939
R6334 vdd.n2254 vdd.n1504 0.152939
R6335 vdd.n2270 vdd.n1504 0.152939
R6336 vdd.n2271 vdd.n2270 0.152939
R6337 vdd.n2272 vdd.n2271 0.152939
R6338 vdd.n670 vdd.n667 0.152939
R6339 vdd.n671 vdd.n670 0.152939
R6340 vdd.n672 vdd.n671 0.152939
R6341 vdd.n673 vdd.n672 0.152939
R6342 vdd.n676 vdd.n673 0.152939
R6343 vdd.n677 vdd.n676 0.152939
R6344 vdd.n678 vdd.n677 0.152939
R6345 vdd.n679 vdd.n678 0.152939
R6346 vdd.n682 vdd.n679 0.152939
R6347 vdd.n683 vdd.n682 0.152939
R6348 vdd.n684 vdd.n683 0.152939
R6349 vdd.n685 vdd.n684 0.152939
R6350 vdd.n690 vdd.n685 0.152939
R6351 vdd.n691 vdd.n690 0.152939
R6352 vdd.n692 vdd.n691 0.152939
R6353 vdd.n693 vdd.n692 0.152939
R6354 vdd.n696 vdd.n693 0.152939
R6355 vdd.n697 vdd.n696 0.152939
R6356 vdd.n698 vdd.n697 0.152939
R6357 vdd.n699 vdd.n698 0.152939
R6358 vdd.n702 vdd.n699 0.152939
R6359 vdd.n703 vdd.n702 0.152939
R6360 vdd.n704 vdd.n703 0.152939
R6361 vdd.n705 vdd.n704 0.152939
R6362 vdd.n708 vdd.n705 0.152939
R6363 vdd.n709 vdd.n708 0.152939
R6364 vdd.n710 vdd.n709 0.152939
R6365 vdd.n711 vdd.n710 0.152939
R6366 vdd.n714 vdd.n711 0.152939
R6367 vdd.n715 vdd.n714 0.152939
R6368 vdd.n716 vdd.n715 0.152939
R6369 vdd.n717 vdd.n716 0.152939
R6370 vdd.n720 vdd.n717 0.152939
R6371 vdd.n721 vdd.n720 0.152939
R6372 vdd.n3330 vdd.n721 0.152939
R6373 vdd.n3330 vdd.n3329 0.152939
R6374 vdd.n3329 vdd.n3328 0.152939
R6375 vdd.n3328 vdd.n725 0.152939
R6376 vdd.n730 vdd.n725 0.152939
R6377 vdd.n731 vdd.n730 0.152939
R6378 vdd.n734 vdd.n731 0.152939
R6379 vdd.n735 vdd.n734 0.152939
R6380 vdd.n736 vdd.n735 0.152939
R6381 vdd.n737 vdd.n736 0.152939
R6382 vdd.n740 vdd.n737 0.152939
R6383 vdd.n741 vdd.n740 0.152939
R6384 vdd.n742 vdd.n741 0.152939
R6385 vdd.n743 vdd.n742 0.152939
R6386 vdd.n746 vdd.n743 0.152939
R6387 vdd.n747 vdd.n746 0.152939
R6388 vdd.n748 vdd.n747 0.152939
R6389 vdd.n3413 vdd.n661 0.152939
R6390 vdd.n3414 vdd.n651 0.152939
R6391 vdd.n3428 vdd.n651 0.152939
R6392 vdd.n3429 vdd.n3428 0.152939
R6393 vdd.n3430 vdd.n3429 0.152939
R6394 vdd.n3430 vdd.n639 0.152939
R6395 vdd.n3444 vdd.n639 0.152939
R6396 vdd.n3445 vdd.n3444 0.152939
R6397 vdd.n3446 vdd.n3445 0.152939
R6398 vdd.n3446 vdd.n627 0.152939
R6399 vdd.n3461 vdd.n627 0.152939
R6400 vdd.n3462 vdd.n3461 0.152939
R6401 vdd.n3463 vdd.n3462 0.152939
R6402 vdd.n3463 vdd.n616 0.152939
R6403 vdd.n3480 vdd.n616 0.152939
R6404 vdd.n3481 vdd.n3480 0.152939
R6405 vdd.n3482 vdd.n3481 0.152939
R6406 vdd.n3482 vdd.n322 0.152939
R6407 vdd.n3562 vdd.n323 0.152939
R6408 vdd.n334 vdd.n323 0.152939
R6409 vdd.n335 vdd.n334 0.152939
R6410 vdd.n336 vdd.n335 0.152939
R6411 vdd.n343 vdd.n336 0.152939
R6412 vdd.n344 vdd.n343 0.152939
R6413 vdd.n345 vdd.n344 0.152939
R6414 vdd.n346 vdd.n345 0.152939
R6415 vdd.n354 vdd.n346 0.152939
R6416 vdd.n355 vdd.n354 0.152939
R6417 vdd.n356 vdd.n355 0.152939
R6418 vdd.n357 vdd.n356 0.152939
R6419 vdd.n365 vdd.n357 0.152939
R6420 vdd.n366 vdd.n365 0.152939
R6421 vdd.n367 vdd.n366 0.152939
R6422 vdd.n368 vdd.n367 0.152939
R6423 vdd.n443 vdd.n368 0.152939
R6424 vdd.n444 vdd.n442 0.152939
R6425 vdd.n451 vdd.n442 0.152939
R6426 vdd.n452 vdd.n451 0.152939
R6427 vdd.n453 vdd.n452 0.152939
R6428 vdd.n453 vdd.n440 0.152939
R6429 vdd.n461 vdd.n440 0.152939
R6430 vdd.n462 vdd.n461 0.152939
R6431 vdd.n463 vdd.n462 0.152939
R6432 vdd.n463 vdd.n438 0.152939
R6433 vdd.n471 vdd.n438 0.152939
R6434 vdd.n472 vdd.n471 0.152939
R6435 vdd.n473 vdd.n472 0.152939
R6436 vdd.n473 vdd.n436 0.152939
R6437 vdd.n481 vdd.n436 0.152939
R6438 vdd.n482 vdd.n481 0.152939
R6439 vdd.n483 vdd.n482 0.152939
R6440 vdd.n483 vdd.n434 0.152939
R6441 vdd.n491 vdd.n434 0.152939
R6442 vdd.n492 vdd.n491 0.152939
R6443 vdd.n493 vdd.n492 0.152939
R6444 vdd.n493 vdd.n430 0.152939
R6445 vdd.n501 vdd.n430 0.152939
R6446 vdd.n502 vdd.n501 0.152939
R6447 vdd.n503 vdd.n502 0.152939
R6448 vdd.n503 vdd.n428 0.152939
R6449 vdd.n511 vdd.n428 0.152939
R6450 vdd.n512 vdd.n511 0.152939
R6451 vdd.n513 vdd.n512 0.152939
R6452 vdd.n513 vdd.n426 0.152939
R6453 vdd.n521 vdd.n426 0.152939
R6454 vdd.n522 vdd.n521 0.152939
R6455 vdd.n523 vdd.n522 0.152939
R6456 vdd.n523 vdd.n424 0.152939
R6457 vdd.n531 vdd.n424 0.152939
R6458 vdd.n532 vdd.n531 0.152939
R6459 vdd.n533 vdd.n532 0.152939
R6460 vdd.n533 vdd.n422 0.152939
R6461 vdd.n541 vdd.n422 0.152939
R6462 vdd.n542 vdd.n541 0.152939
R6463 vdd.n543 vdd.n542 0.152939
R6464 vdd.n543 vdd.n418 0.152939
R6465 vdd.n551 vdd.n418 0.152939
R6466 vdd.n552 vdd.n551 0.152939
R6467 vdd.n553 vdd.n552 0.152939
R6468 vdd.n553 vdd.n416 0.152939
R6469 vdd.n561 vdd.n416 0.152939
R6470 vdd.n562 vdd.n561 0.152939
R6471 vdd.n563 vdd.n562 0.152939
R6472 vdd.n563 vdd.n414 0.152939
R6473 vdd.n571 vdd.n414 0.152939
R6474 vdd.n572 vdd.n571 0.152939
R6475 vdd.n573 vdd.n572 0.152939
R6476 vdd.n573 vdd.n412 0.152939
R6477 vdd.n581 vdd.n412 0.152939
R6478 vdd.n582 vdd.n581 0.152939
R6479 vdd.n583 vdd.n582 0.152939
R6480 vdd.n583 vdd.n410 0.152939
R6481 vdd.n591 vdd.n410 0.152939
R6482 vdd.n592 vdd.n591 0.152939
R6483 vdd.n593 vdd.n592 0.152939
R6484 vdd.n593 vdd.n408 0.152939
R6485 vdd.n600 vdd.n408 0.152939
R6486 vdd.n3521 vdd.n600 0.152939
R6487 vdd.n3421 vdd.n3420 0.152939
R6488 vdd.n3422 vdd.n3421 0.152939
R6489 vdd.n3422 vdd.n645 0.152939
R6490 vdd.n3436 vdd.n645 0.152939
R6491 vdd.n3437 vdd.n3436 0.152939
R6492 vdd.n3438 vdd.n3437 0.152939
R6493 vdd.n3438 vdd.n632 0.152939
R6494 vdd.n3452 vdd.n632 0.152939
R6495 vdd.n3453 vdd.n3452 0.152939
R6496 vdd.n3454 vdd.n3453 0.152939
R6497 vdd.n3454 vdd.n621 0.152939
R6498 vdd.n3469 vdd.n621 0.152939
R6499 vdd.n3470 vdd.n3469 0.152939
R6500 vdd.n3471 vdd.n3470 0.152939
R6501 vdd.n3473 vdd.n3471 0.152939
R6502 vdd.n3473 vdd.n3472 0.152939
R6503 vdd.n3472 vdd.n611 0.152939
R6504 vdd.n611 vdd.n609 0.152939
R6505 vdd.n3491 vdd.n609 0.152939
R6506 vdd.n3492 vdd.n3491 0.152939
R6507 vdd.n3493 vdd.n3492 0.152939
R6508 vdd.n3493 vdd.n607 0.152939
R6509 vdd.n3498 vdd.n607 0.152939
R6510 vdd.n3499 vdd.n3498 0.152939
R6511 vdd.n3500 vdd.n3499 0.152939
R6512 vdd.n3500 vdd.n605 0.152939
R6513 vdd.n3505 vdd.n605 0.152939
R6514 vdd.n3506 vdd.n3505 0.152939
R6515 vdd.n3507 vdd.n3506 0.152939
R6516 vdd.n3507 vdd.n603 0.152939
R6517 vdd.n3513 vdd.n603 0.152939
R6518 vdd.n3514 vdd.n3513 0.152939
R6519 vdd.n3515 vdd.n3514 0.152939
R6520 vdd.n3515 vdd.n601 0.152939
R6521 vdd.n3520 vdd.n601 0.152939
R6522 vdd.n3283 vdd.n656 0.152939
R6523 vdd.n2283 vdd.n1488 0.152939
R6524 vdd.n1834 vdd.n1833 0.152939
R6525 vdd.n1834 vdd.n1590 0.152939
R6526 vdd.n1848 vdd.n1590 0.152939
R6527 vdd.n1849 vdd.n1848 0.152939
R6528 vdd.n1850 vdd.n1849 0.152939
R6529 vdd.n1850 vdd.n1578 0.152939
R6530 vdd.n1865 vdd.n1578 0.152939
R6531 vdd.n1866 vdd.n1865 0.152939
R6532 vdd.n1867 vdd.n1866 0.152939
R6533 vdd.n1867 vdd.n1568 0.152939
R6534 vdd.n1882 vdd.n1568 0.152939
R6535 vdd.n1883 vdd.n1882 0.152939
R6536 vdd.n1884 vdd.n1883 0.152939
R6537 vdd.n1884 vdd.n1555 0.152939
R6538 vdd.n1898 vdd.n1555 0.152939
R6539 vdd.n1899 vdd.n1898 0.152939
R6540 vdd.n1900 vdd.n1899 0.152939
R6541 vdd.n1900 vdd.n1544 0.152939
R6542 vdd.n2210 vdd.n1544 0.152939
R6543 vdd.n2211 vdd.n2210 0.152939
R6544 vdd.n2212 vdd.n2211 0.152939
R6545 vdd.n2212 vdd.n1533 0.152939
R6546 vdd.n2226 vdd.n1533 0.152939
R6547 vdd.n2227 vdd.n2226 0.152939
R6548 vdd.n2228 vdd.n2227 0.152939
R6549 vdd.n2228 vdd.n1521 0.152939
R6550 vdd.n2243 vdd.n1521 0.152939
R6551 vdd.n2244 vdd.n2243 0.152939
R6552 vdd.n2245 vdd.n2244 0.152939
R6553 vdd.n2245 vdd.n1511 0.152939
R6554 vdd.n2260 vdd.n1511 0.152939
R6555 vdd.n2261 vdd.n2260 0.152939
R6556 vdd.n2264 vdd.n2261 0.152939
R6557 vdd.n2264 vdd.n2263 0.152939
R6558 vdd.n2263 vdd.n2262 0.152939
R6559 vdd.n1824 vdd.n1639 0.152939
R6560 vdd.n1824 vdd.n1823 0.152939
R6561 vdd.n1823 vdd.n1822 0.152939
R6562 vdd.n1822 vdd.n1641 0.152939
R6563 vdd.n1818 vdd.n1641 0.152939
R6564 vdd.n1818 vdd.n1817 0.152939
R6565 vdd.n1817 vdd.n1816 0.152939
R6566 vdd.n1816 vdd.n1646 0.152939
R6567 vdd.n1812 vdd.n1646 0.152939
R6568 vdd.n1812 vdd.n1811 0.152939
R6569 vdd.n1811 vdd.n1810 0.152939
R6570 vdd.n1810 vdd.n1652 0.152939
R6571 vdd.n1806 vdd.n1652 0.152939
R6572 vdd.n1806 vdd.n1805 0.152939
R6573 vdd.n1805 vdd.n1804 0.152939
R6574 vdd.n1804 vdd.n1658 0.152939
R6575 vdd.n1800 vdd.n1658 0.152939
R6576 vdd.n1800 vdd.n1799 0.152939
R6577 vdd.n1799 vdd.n1798 0.152939
R6578 vdd.n1798 vdd.n1664 0.152939
R6579 vdd.n1790 vdd.n1664 0.152939
R6580 vdd.n1790 vdd.n1789 0.152939
R6581 vdd.n1789 vdd.n1788 0.152939
R6582 vdd.n1788 vdd.n1668 0.152939
R6583 vdd.n1784 vdd.n1668 0.152939
R6584 vdd.n1784 vdd.n1783 0.152939
R6585 vdd.n1783 vdd.n1782 0.152939
R6586 vdd.n1782 vdd.n1674 0.152939
R6587 vdd.n1778 vdd.n1674 0.152939
R6588 vdd.n1778 vdd.n1777 0.152939
R6589 vdd.n1777 vdd.n1776 0.152939
R6590 vdd.n1776 vdd.n1680 0.152939
R6591 vdd.n1772 vdd.n1680 0.152939
R6592 vdd.n1772 vdd.n1771 0.152939
R6593 vdd.n1771 vdd.n1770 0.152939
R6594 vdd.n1770 vdd.n1686 0.152939
R6595 vdd.n1766 vdd.n1686 0.152939
R6596 vdd.n1766 vdd.n1765 0.152939
R6597 vdd.n1765 vdd.n1764 0.152939
R6598 vdd.n1764 vdd.n1692 0.152939
R6599 vdd.n1757 vdd.n1692 0.152939
R6600 vdd.n1757 vdd.n1756 0.152939
R6601 vdd.n1756 vdd.n1755 0.152939
R6602 vdd.n1755 vdd.n1697 0.152939
R6603 vdd.n1751 vdd.n1697 0.152939
R6604 vdd.n1751 vdd.n1750 0.152939
R6605 vdd.n1750 vdd.n1749 0.152939
R6606 vdd.n1749 vdd.n1703 0.152939
R6607 vdd.n1745 vdd.n1703 0.152939
R6608 vdd.n1745 vdd.n1744 0.152939
R6609 vdd.n1744 vdd.n1743 0.152939
R6610 vdd.n1743 vdd.n1709 0.152939
R6611 vdd.n1739 vdd.n1709 0.152939
R6612 vdd.n1739 vdd.n1738 0.152939
R6613 vdd.n1738 vdd.n1737 0.152939
R6614 vdd.n1737 vdd.n1715 0.152939
R6615 vdd.n1733 vdd.n1715 0.152939
R6616 vdd.n1733 vdd.n1732 0.152939
R6617 vdd.n1732 vdd.n1731 0.152939
R6618 vdd.n1731 vdd.n1721 0.152939
R6619 vdd.n1727 vdd.n1721 0.152939
R6620 vdd.n1727 vdd.n1602 0.152939
R6621 vdd.n1832 vdd.n1602 0.152939
R6622 vdd.n1840 vdd.n1596 0.152939
R6623 vdd.n1841 vdd.n1840 0.152939
R6624 vdd.n1842 vdd.n1841 0.152939
R6625 vdd.n1842 vdd.n1584 0.152939
R6626 vdd.n1857 vdd.n1584 0.152939
R6627 vdd.n1858 vdd.n1857 0.152939
R6628 vdd.n1859 vdd.n1858 0.152939
R6629 vdd.n1859 vdd.n1573 0.152939
R6630 vdd.n1874 vdd.n1573 0.152939
R6631 vdd.n1875 vdd.n1874 0.152939
R6632 vdd.n1876 vdd.n1875 0.152939
R6633 vdd.n1876 vdd.n1562 0.152939
R6634 vdd.n1890 vdd.n1562 0.152939
R6635 vdd.n1891 vdd.n1890 0.152939
R6636 vdd.n1892 vdd.n1891 0.152939
R6637 vdd.n1892 vdd.n1550 0.152939
R6638 vdd.n1907 vdd.n1550 0.152939
R6639 vdd.n2391 vdd.n2390 0.110256
R6640 vdd.n3214 vdd.n661 0.110256
R6641 vdd.n3283 vdd.n3282 0.110256
R6642 vdd.n2284 vdd.n2283 0.110256
R6643 vdd.n2203 vdd.n2202 0.0695946
R6644 vdd.n3563 vdd.n322 0.0695946
R6645 vdd.n3563 vdd.n3562 0.0695946
R6646 vdd.n2202 vdd.n1907 0.0695946
R6647 vdd.n2391 vdd.n1149 0.0431829
R6648 vdd.n2284 vdd.n1249 0.0431829
R6649 vdd.n3214 vdd.n667 0.0431829
R6650 vdd.n3282 vdd.n748 0.0431829
R6651 vdd vdd.n28 0.00833333
R6652 commonsourceibias.n397 commonsourceibias.t184 222.032
R6653 commonsourceibias.n281 commonsourceibias.t134 222.032
R6654 commonsourceibias.n44 commonsourceibias.t22 222.032
R6655 commonsourceibias.n166 commonsourceibias.t140 222.032
R6656 commonsourceibias.n875 commonsourceibias.t191 222.032
R6657 commonsourceibias.n759 commonsourceibias.t98 222.032
R6658 commonsourceibias.n529 commonsourceibias.t76 222.032
R6659 commonsourceibias.n645 commonsourceibias.t177 222.032
R6660 commonsourceibias.n480 commonsourceibias.t183 207.983
R6661 commonsourceibias.n364 commonsourceibias.t88 207.983
R6662 commonsourceibias.n127 commonsourceibias.t66 207.983
R6663 commonsourceibias.n249 commonsourceibias.t151 207.983
R6664 commonsourceibias.n963 commonsourceibias.t101 207.983
R6665 commonsourceibias.n847 commonsourceibias.t189 207.983
R6666 commonsourceibias.n617 commonsourceibias.t40 207.983
R6667 commonsourceibias.n732 commonsourceibias.t112 207.983
R6668 commonsourceibias.n396 commonsourceibias.t150 168.701
R6669 commonsourceibias.n402 commonsourceibias.t155 168.701
R6670 commonsourceibias.n408 commonsourceibias.t199 168.701
R6671 commonsourceibias.n392 commonsourceibias.t175 168.701
R6672 commonsourceibias.n416 commonsourceibias.t165 168.701
R6673 commonsourceibias.n422 commonsourceibias.t96 168.701
R6674 commonsourceibias.n387 commonsourceibias.t187 168.701
R6675 commonsourceibias.n430 commonsourceibias.t168 168.701
R6676 commonsourceibias.n436 commonsourceibias.t172 168.701
R6677 commonsourceibias.n382 commonsourceibias.t80 168.701
R6678 commonsourceibias.n444 commonsourceibias.t173 168.701
R6679 commonsourceibias.n450 commonsourceibias.t182 168.701
R6680 commonsourceibias.n377 commonsourceibias.t149 168.701
R6681 commonsourceibias.n458 commonsourceibias.t110 168.701
R6682 commonsourceibias.n464 commonsourceibias.t194 168.701
R6683 commonsourceibias.n372 commonsourceibias.t157 168.701
R6684 commonsourceibias.n472 commonsourceibias.t163 168.701
R6685 commonsourceibias.n478 commonsourceibias.t92 168.701
R6686 commonsourceibias.n362 commonsourceibias.t198 168.701
R6687 commonsourceibias.n356 commonsourceibias.t186 168.701
R6688 commonsourceibias.n256 commonsourceibias.t95 168.701
R6689 commonsourceibias.n348 commonsourceibias.t196 168.701
R6690 commonsourceibias.n342 commonsourceibias.t105 168.701
R6691 commonsourceibias.n261 commonsourceibias.t94 168.701
R6692 commonsourceibias.n334 commonsourceibias.t197 168.701
R6693 commonsourceibias.n328 commonsourceibias.t115 168.701
R6694 commonsourceibias.n266 commonsourceibias.t141 168.701
R6695 commonsourceibias.n320 commonsourceibias.t195 168.701
R6696 commonsourceibias.n314 commonsourceibias.t113 168.701
R6697 commonsourceibias.n271 commonsourceibias.t138 168.701
R6698 commonsourceibias.n306 commonsourceibias.t130 168.701
R6699 commonsourceibias.n300 commonsourceibias.t114 168.701
R6700 commonsourceibias.n276 commonsourceibias.t139 168.701
R6701 commonsourceibias.n292 commonsourceibias.t129 168.701
R6702 commonsourceibias.n286 commonsourceibias.t125 168.701
R6703 commonsourceibias.n280 commonsourceibias.t147 168.701
R6704 commonsourceibias.n125 commonsourceibias.t10 168.701
R6705 commonsourceibias.n119 commonsourceibias.t58 168.701
R6706 commonsourceibias.n19 commonsourceibias.t64 168.701
R6707 commonsourceibias.n111 commonsourceibias.t2 168.701
R6708 commonsourceibias.n105 commonsourceibias.t70 168.701
R6709 commonsourceibias.n24 commonsourceibias.t54 168.701
R6710 commonsourceibias.n97 commonsourceibias.t60 168.701
R6711 commonsourceibias.n91 commonsourceibias.t68 168.701
R6712 commonsourceibias.n29 commonsourceibias.t30 168.701
R6713 commonsourceibias.n83 commonsourceibias.t50 168.701
R6714 commonsourceibias.n77 commonsourceibias.t24 168.701
R6715 commonsourceibias.n34 commonsourceibias.t78 168.701
R6716 commonsourceibias.n69 commonsourceibias.t18 168.701
R6717 commonsourceibias.n63 commonsourceibias.t6 168.701
R6718 commonsourceibias.n39 commonsourceibias.t14 168.701
R6719 commonsourceibias.n55 commonsourceibias.t42 168.701
R6720 commonsourceibias.n49 commonsourceibias.t28 168.701
R6721 commonsourceibias.n43 commonsourceibias.t4 168.701
R6722 commonsourceibias.n247 commonsourceibias.t83 168.701
R6723 commonsourceibias.n241 commonsourceibias.t161 168.701
R6724 commonsourceibias.n5 commonsourceibias.t152 168.701
R6725 commonsourceibias.n233 commonsourceibias.t171 168.701
R6726 commonsourceibias.n227 commonsourceibias.t145 168.701
R6727 commonsourceibias.n10 commonsourceibias.t124 168.701
R6728 commonsourceibias.n219 commonsourceibias.t158 168.701
R6729 commonsourceibias.n213 commonsourceibias.t148 168.701
R6730 commonsourceibias.n150 commonsourceibias.t93 168.701
R6731 commonsourceibias.n151 commonsourceibias.t131 168.701
R6732 commonsourceibias.n153 commonsourceibias.t117 168.701
R6733 commonsourceibias.n155 commonsourceibias.t176 168.701
R6734 commonsourceibias.n191 commonsourceibias.t144 168.701
R6735 commonsourceibias.n185 commonsourceibias.t190 168.701
R6736 commonsourceibias.n161 commonsourceibias.t164 168.701
R6737 commonsourceibias.n177 commonsourceibias.t111 168.701
R6738 commonsourceibias.n171 commonsourceibias.t100 168.701
R6739 commonsourceibias.n165 commonsourceibias.t84 168.701
R6740 commonsourceibias.n874 commonsourceibias.t156 168.701
R6741 commonsourceibias.n880 commonsourceibias.t146 168.701
R6742 commonsourceibias.n886 commonsourceibias.t126 168.701
R6743 commonsourceibias.n888 commonsourceibias.t91 168.701
R6744 commonsourceibias.n895 commonsourceibias.t181 168.701
R6745 commonsourceibias.n901 commonsourceibias.t136 168.701
R6746 commonsourceibias.n903 commonsourceibias.t107 168.701
R6747 commonsourceibias.n910 commonsourceibias.t192 168.701
R6748 commonsourceibias.n916 commonsourceibias.t167 168.701
R6749 commonsourceibias.n918 commonsourceibias.t127 168.701
R6750 commonsourceibias.n925 commonsourceibias.t87 168.701
R6751 commonsourceibias.n931 commonsourceibias.t99 168.701
R6752 commonsourceibias.n933 commonsourceibias.t137 168.701
R6753 commonsourceibias.n940 commonsourceibias.t143 168.701
R6754 commonsourceibias.n946 commonsourceibias.t122 168.701
R6755 commonsourceibias.n948 commonsourceibias.t170 168.701
R6756 commonsourceibias.n955 commonsourceibias.t153 168.701
R6757 commonsourceibias.n961 commonsourceibias.t133 168.701
R6758 commonsourceibias.n758 commonsourceibias.t123 168.701
R6759 commonsourceibias.n764 commonsourceibias.t132 168.701
R6760 commonsourceibias.n770 commonsourceibias.t104 168.701
R6761 commonsourceibias.n772 commonsourceibias.t118 168.701
R6762 commonsourceibias.n779 commonsourceibias.t85 168.701
R6763 commonsourceibias.n785 commonsourceibias.t106 168.701
R6764 commonsourceibias.n787 commonsourceibias.t119 168.701
R6765 commonsourceibias.n794 commonsourceibias.t86 168.701
R6766 commonsourceibias.n800 commonsourceibias.t97 168.701
R6767 commonsourceibias.n802 commonsourceibias.t120 168.701
R6768 commonsourceibias.n809 commonsourceibias.t89 168.701
R6769 commonsourceibias.n815 commonsourceibias.t178 168.701
R6770 commonsourceibias.n817 commonsourceibias.t121 168.701
R6771 commonsourceibias.n824 commonsourceibias.t81 168.701
R6772 commonsourceibias.n830 commonsourceibias.t179 168.701
R6773 commonsourceibias.n832 commonsourceibias.t193 168.701
R6774 commonsourceibias.n839 commonsourceibias.t82 168.701
R6775 commonsourceibias.n845 commonsourceibias.t180 168.701
R6776 commonsourceibias.n528 commonsourceibias.t16 168.701
R6777 commonsourceibias.n534 commonsourceibias.t62 168.701
R6778 commonsourceibias.n540 commonsourceibias.t74 168.701
R6779 commonsourceibias.n542 commonsourceibias.t48 168.701
R6780 commonsourceibias.n549 commonsourceibias.t12 168.701
R6781 commonsourceibias.n555 commonsourceibias.t46 168.701
R6782 commonsourceibias.n557 commonsourceibias.t56 168.701
R6783 commonsourceibias.n564 commonsourceibias.t72 168.701
R6784 commonsourceibias.n570 commonsourceibias.t26 168.701
R6785 commonsourceibias.n572 commonsourceibias.t34 168.701
R6786 commonsourceibias.n579 commonsourceibias.t36 168.701
R6787 commonsourceibias.n585 commonsourceibias.t52 168.701
R6788 commonsourceibias.n587 commonsourceibias.t8 168.701
R6789 commonsourceibias.n594 commonsourceibias.t44 168.701
R6790 commonsourceibias.n600 commonsourceibias.t32 168.701
R6791 commonsourceibias.n602 commonsourceibias.t38 168.701
R6792 commonsourceibias.n609 commonsourceibias.t20 168.701
R6793 commonsourceibias.n615 commonsourceibias.t0 168.701
R6794 commonsourceibias.n730 commonsourceibias.t169 168.701
R6795 commonsourceibias.n724 commonsourceibias.t142 168.701
R6796 commonsourceibias.n717 commonsourceibias.t116 168.701
R6797 commonsourceibias.n715 commonsourceibias.t154 168.701
R6798 commonsourceibias.n709 commonsourceibias.t108 168.701
R6799 commonsourceibias.n702 commonsourceibias.t90 168.701
R6800 commonsourceibias.n700 commonsourceibias.t128 168.701
R6801 commonsourceibias.n694 commonsourceibias.t109 168.701
R6802 commonsourceibias.n687 commonsourceibias.t174 168.701
R6803 commonsourceibias.n644 commonsourceibias.t159 168.701
R6804 commonsourceibias.n650 commonsourceibias.t160 168.701
R6805 commonsourceibias.n656 commonsourceibias.t185 168.701
R6806 commonsourceibias.n658 commonsourceibias.t135 168.701
R6807 commonsourceibias.n665 commonsourceibias.t166 168.701
R6808 commonsourceibias.n671 commonsourceibias.t103 168.701
R6809 commonsourceibias.n635 commonsourceibias.t162 168.701
R6810 commonsourceibias.n633 commonsourceibias.t188 168.701
R6811 commonsourceibias.n631 commonsourceibias.t102 168.701
R6812 commonsourceibias.n479 commonsourceibias.n367 161.3
R6813 commonsourceibias.n477 commonsourceibias.n476 161.3
R6814 commonsourceibias.n475 commonsourceibias.n368 161.3
R6815 commonsourceibias.n474 commonsourceibias.n473 161.3
R6816 commonsourceibias.n471 commonsourceibias.n369 161.3
R6817 commonsourceibias.n470 commonsourceibias.n469 161.3
R6818 commonsourceibias.n468 commonsourceibias.n370 161.3
R6819 commonsourceibias.n467 commonsourceibias.n466 161.3
R6820 commonsourceibias.n465 commonsourceibias.n371 161.3
R6821 commonsourceibias.n463 commonsourceibias.n462 161.3
R6822 commonsourceibias.n461 commonsourceibias.n373 161.3
R6823 commonsourceibias.n460 commonsourceibias.n459 161.3
R6824 commonsourceibias.n457 commonsourceibias.n374 161.3
R6825 commonsourceibias.n456 commonsourceibias.n455 161.3
R6826 commonsourceibias.n454 commonsourceibias.n375 161.3
R6827 commonsourceibias.n453 commonsourceibias.n452 161.3
R6828 commonsourceibias.n451 commonsourceibias.n376 161.3
R6829 commonsourceibias.n449 commonsourceibias.n448 161.3
R6830 commonsourceibias.n447 commonsourceibias.n378 161.3
R6831 commonsourceibias.n446 commonsourceibias.n445 161.3
R6832 commonsourceibias.n443 commonsourceibias.n379 161.3
R6833 commonsourceibias.n442 commonsourceibias.n441 161.3
R6834 commonsourceibias.n440 commonsourceibias.n380 161.3
R6835 commonsourceibias.n439 commonsourceibias.n438 161.3
R6836 commonsourceibias.n437 commonsourceibias.n381 161.3
R6837 commonsourceibias.n435 commonsourceibias.n434 161.3
R6838 commonsourceibias.n433 commonsourceibias.n383 161.3
R6839 commonsourceibias.n432 commonsourceibias.n431 161.3
R6840 commonsourceibias.n429 commonsourceibias.n384 161.3
R6841 commonsourceibias.n428 commonsourceibias.n427 161.3
R6842 commonsourceibias.n426 commonsourceibias.n385 161.3
R6843 commonsourceibias.n425 commonsourceibias.n424 161.3
R6844 commonsourceibias.n423 commonsourceibias.n386 161.3
R6845 commonsourceibias.n421 commonsourceibias.n420 161.3
R6846 commonsourceibias.n419 commonsourceibias.n388 161.3
R6847 commonsourceibias.n418 commonsourceibias.n417 161.3
R6848 commonsourceibias.n415 commonsourceibias.n389 161.3
R6849 commonsourceibias.n414 commonsourceibias.n413 161.3
R6850 commonsourceibias.n412 commonsourceibias.n390 161.3
R6851 commonsourceibias.n411 commonsourceibias.n410 161.3
R6852 commonsourceibias.n409 commonsourceibias.n391 161.3
R6853 commonsourceibias.n407 commonsourceibias.n406 161.3
R6854 commonsourceibias.n405 commonsourceibias.n393 161.3
R6855 commonsourceibias.n404 commonsourceibias.n403 161.3
R6856 commonsourceibias.n401 commonsourceibias.n394 161.3
R6857 commonsourceibias.n400 commonsourceibias.n399 161.3
R6858 commonsourceibias.n398 commonsourceibias.n395 161.3
R6859 commonsourceibias.n282 commonsourceibias.n279 161.3
R6860 commonsourceibias.n284 commonsourceibias.n283 161.3
R6861 commonsourceibias.n285 commonsourceibias.n278 161.3
R6862 commonsourceibias.n288 commonsourceibias.n287 161.3
R6863 commonsourceibias.n289 commonsourceibias.n277 161.3
R6864 commonsourceibias.n291 commonsourceibias.n290 161.3
R6865 commonsourceibias.n293 commonsourceibias.n275 161.3
R6866 commonsourceibias.n295 commonsourceibias.n294 161.3
R6867 commonsourceibias.n296 commonsourceibias.n274 161.3
R6868 commonsourceibias.n298 commonsourceibias.n297 161.3
R6869 commonsourceibias.n299 commonsourceibias.n273 161.3
R6870 commonsourceibias.n302 commonsourceibias.n301 161.3
R6871 commonsourceibias.n303 commonsourceibias.n272 161.3
R6872 commonsourceibias.n305 commonsourceibias.n304 161.3
R6873 commonsourceibias.n307 commonsourceibias.n270 161.3
R6874 commonsourceibias.n309 commonsourceibias.n308 161.3
R6875 commonsourceibias.n310 commonsourceibias.n269 161.3
R6876 commonsourceibias.n312 commonsourceibias.n311 161.3
R6877 commonsourceibias.n313 commonsourceibias.n268 161.3
R6878 commonsourceibias.n316 commonsourceibias.n315 161.3
R6879 commonsourceibias.n317 commonsourceibias.n267 161.3
R6880 commonsourceibias.n319 commonsourceibias.n318 161.3
R6881 commonsourceibias.n321 commonsourceibias.n265 161.3
R6882 commonsourceibias.n323 commonsourceibias.n322 161.3
R6883 commonsourceibias.n324 commonsourceibias.n264 161.3
R6884 commonsourceibias.n326 commonsourceibias.n325 161.3
R6885 commonsourceibias.n327 commonsourceibias.n263 161.3
R6886 commonsourceibias.n330 commonsourceibias.n329 161.3
R6887 commonsourceibias.n331 commonsourceibias.n262 161.3
R6888 commonsourceibias.n333 commonsourceibias.n332 161.3
R6889 commonsourceibias.n335 commonsourceibias.n260 161.3
R6890 commonsourceibias.n337 commonsourceibias.n336 161.3
R6891 commonsourceibias.n338 commonsourceibias.n259 161.3
R6892 commonsourceibias.n340 commonsourceibias.n339 161.3
R6893 commonsourceibias.n341 commonsourceibias.n258 161.3
R6894 commonsourceibias.n344 commonsourceibias.n343 161.3
R6895 commonsourceibias.n345 commonsourceibias.n257 161.3
R6896 commonsourceibias.n347 commonsourceibias.n346 161.3
R6897 commonsourceibias.n349 commonsourceibias.n255 161.3
R6898 commonsourceibias.n351 commonsourceibias.n350 161.3
R6899 commonsourceibias.n352 commonsourceibias.n254 161.3
R6900 commonsourceibias.n354 commonsourceibias.n353 161.3
R6901 commonsourceibias.n355 commonsourceibias.n253 161.3
R6902 commonsourceibias.n358 commonsourceibias.n357 161.3
R6903 commonsourceibias.n359 commonsourceibias.n252 161.3
R6904 commonsourceibias.n361 commonsourceibias.n360 161.3
R6905 commonsourceibias.n363 commonsourceibias.n251 161.3
R6906 commonsourceibias.n45 commonsourceibias.n42 161.3
R6907 commonsourceibias.n47 commonsourceibias.n46 161.3
R6908 commonsourceibias.n48 commonsourceibias.n41 161.3
R6909 commonsourceibias.n51 commonsourceibias.n50 161.3
R6910 commonsourceibias.n52 commonsourceibias.n40 161.3
R6911 commonsourceibias.n54 commonsourceibias.n53 161.3
R6912 commonsourceibias.n56 commonsourceibias.n38 161.3
R6913 commonsourceibias.n58 commonsourceibias.n57 161.3
R6914 commonsourceibias.n59 commonsourceibias.n37 161.3
R6915 commonsourceibias.n61 commonsourceibias.n60 161.3
R6916 commonsourceibias.n62 commonsourceibias.n36 161.3
R6917 commonsourceibias.n65 commonsourceibias.n64 161.3
R6918 commonsourceibias.n66 commonsourceibias.n35 161.3
R6919 commonsourceibias.n68 commonsourceibias.n67 161.3
R6920 commonsourceibias.n70 commonsourceibias.n33 161.3
R6921 commonsourceibias.n72 commonsourceibias.n71 161.3
R6922 commonsourceibias.n73 commonsourceibias.n32 161.3
R6923 commonsourceibias.n75 commonsourceibias.n74 161.3
R6924 commonsourceibias.n76 commonsourceibias.n31 161.3
R6925 commonsourceibias.n79 commonsourceibias.n78 161.3
R6926 commonsourceibias.n80 commonsourceibias.n30 161.3
R6927 commonsourceibias.n82 commonsourceibias.n81 161.3
R6928 commonsourceibias.n84 commonsourceibias.n28 161.3
R6929 commonsourceibias.n86 commonsourceibias.n85 161.3
R6930 commonsourceibias.n87 commonsourceibias.n27 161.3
R6931 commonsourceibias.n89 commonsourceibias.n88 161.3
R6932 commonsourceibias.n90 commonsourceibias.n26 161.3
R6933 commonsourceibias.n93 commonsourceibias.n92 161.3
R6934 commonsourceibias.n94 commonsourceibias.n25 161.3
R6935 commonsourceibias.n96 commonsourceibias.n95 161.3
R6936 commonsourceibias.n98 commonsourceibias.n23 161.3
R6937 commonsourceibias.n100 commonsourceibias.n99 161.3
R6938 commonsourceibias.n101 commonsourceibias.n22 161.3
R6939 commonsourceibias.n103 commonsourceibias.n102 161.3
R6940 commonsourceibias.n104 commonsourceibias.n21 161.3
R6941 commonsourceibias.n107 commonsourceibias.n106 161.3
R6942 commonsourceibias.n108 commonsourceibias.n20 161.3
R6943 commonsourceibias.n110 commonsourceibias.n109 161.3
R6944 commonsourceibias.n112 commonsourceibias.n18 161.3
R6945 commonsourceibias.n114 commonsourceibias.n113 161.3
R6946 commonsourceibias.n115 commonsourceibias.n17 161.3
R6947 commonsourceibias.n117 commonsourceibias.n116 161.3
R6948 commonsourceibias.n118 commonsourceibias.n16 161.3
R6949 commonsourceibias.n121 commonsourceibias.n120 161.3
R6950 commonsourceibias.n122 commonsourceibias.n15 161.3
R6951 commonsourceibias.n124 commonsourceibias.n123 161.3
R6952 commonsourceibias.n126 commonsourceibias.n14 161.3
R6953 commonsourceibias.n167 commonsourceibias.n164 161.3
R6954 commonsourceibias.n169 commonsourceibias.n168 161.3
R6955 commonsourceibias.n170 commonsourceibias.n163 161.3
R6956 commonsourceibias.n173 commonsourceibias.n172 161.3
R6957 commonsourceibias.n174 commonsourceibias.n162 161.3
R6958 commonsourceibias.n176 commonsourceibias.n175 161.3
R6959 commonsourceibias.n178 commonsourceibias.n160 161.3
R6960 commonsourceibias.n180 commonsourceibias.n179 161.3
R6961 commonsourceibias.n181 commonsourceibias.n159 161.3
R6962 commonsourceibias.n183 commonsourceibias.n182 161.3
R6963 commonsourceibias.n184 commonsourceibias.n158 161.3
R6964 commonsourceibias.n187 commonsourceibias.n186 161.3
R6965 commonsourceibias.n188 commonsourceibias.n157 161.3
R6966 commonsourceibias.n190 commonsourceibias.n189 161.3
R6967 commonsourceibias.n192 commonsourceibias.n156 161.3
R6968 commonsourceibias.n194 commonsourceibias.n193 161.3
R6969 commonsourceibias.n196 commonsourceibias.n195 161.3
R6970 commonsourceibias.n197 commonsourceibias.n154 161.3
R6971 commonsourceibias.n199 commonsourceibias.n198 161.3
R6972 commonsourceibias.n201 commonsourceibias.n200 161.3
R6973 commonsourceibias.n202 commonsourceibias.n152 161.3
R6974 commonsourceibias.n204 commonsourceibias.n203 161.3
R6975 commonsourceibias.n206 commonsourceibias.n205 161.3
R6976 commonsourceibias.n208 commonsourceibias.n207 161.3
R6977 commonsourceibias.n209 commonsourceibias.n13 161.3
R6978 commonsourceibias.n211 commonsourceibias.n210 161.3
R6979 commonsourceibias.n212 commonsourceibias.n12 161.3
R6980 commonsourceibias.n215 commonsourceibias.n214 161.3
R6981 commonsourceibias.n216 commonsourceibias.n11 161.3
R6982 commonsourceibias.n218 commonsourceibias.n217 161.3
R6983 commonsourceibias.n220 commonsourceibias.n9 161.3
R6984 commonsourceibias.n222 commonsourceibias.n221 161.3
R6985 commonsourceibias.n223 commonsourceibias.n8 161.3
R6986 commonsourceibias.n225 commonsourceibias.n224 161.3
R6987 commonsourceibias.n226 commonsourceibias.n7 161.3
R6988 commonsourceibias.n229 commonsourceibias.n228 161.3
R6989 commonsourceibias.n230 commonsourceibias.n6 161.3
R6990 commonsourceibias.n232 commonsourceibias.n231 161.3
R6991 commonsourceibias.n234 commonsourceibias.n4 161.3
R6992 commonsourceibias.n236 commonsourceibias.n235 161.3
R6993 commonsourceibias.n237 commonsourceibias.n3 161.3
R6994 commonsourceibias.n239 commonsourceibias.n238 161.3
R6995 commonsourceibias.n240 commonsourceibias.n2 161.3
R6996 commonsourceibias.n243 commonsourceibias.n242 161.3
R6997 commonsourceibias.n244 commonsourceibias.n1 161.3
R6998 commonsourceibias.n246 commonsourceibias.n245 161.3
R6999 commonsourceibias.n248 commonsourceibias.n0 161.3
R7000 commonsourceibias.n962 commonsourceibias.n850 161.3
R7001 commonsourceibias.n960 commonsourceibias.n959 161.3
R7002 commonsourceibias.n958 commonsourceibias.n851 161.3
R7003 commonsourceibias.n957 commonsourceibias.n956 161.3
R7004 commonsourceibias.n954 commonsourceibias.n852 161.3
R7005 commonsourceibias.n953 commonsourceibias.n952 161.3
R7006 commonsourceibias.n951 commonsourceibias.n853 161.3
R7007 commonsourceibias.n950 commonsourceibias.n949 161.3
R7008 commonsourceibias.n947 commonsourceibias.n854 161.3
R7009 commonsourceibias.n945 commonsourceibias.n944 161.3
R7010 commonsourceibias.n943 commonsourceibias.n855 161.3
R7011 commonsourceibias.n942 commonsourceibias.n941 161.3
R7012 commonsourceibias.n939 commonsourceibias.n856 161.3
R7013 commonsourceibias.n938 commonsourceibias.n937 161.3
R7014 commonsourceibias.n936 commonsourceibias.n857 161.3
R7015 commonsourceibias.n935 commonsourceibias.n934 161.3
R7016 commonsourceibias.n932 commonsourceibias.n858 161.3
R7017 commonsourceibias.n930 commonsourceibias.n929 161.3
R7018 commonsourceibias.n928 commonsourceibias.n859 161.3
R7019 commonsourceibias.n927 commonsourceibias.n926 161.3
R7020 commonsourceibias.n924 commonsourceibias.n860 161.3
R7021 commonsourceibias.n923 commonsourceibias.n922 161.3
R7022 commonsourceibias.n921 commonsourceibias.n861 161.3
R7023 commonsourceibias.n920 commonsourceibias.n919 161.3
R7024 commonsourceibias.n917 commonsourceibias.n862 161.3
R7025 commonsourceibias.n915 commonsourceibias.n914 161.3
R7026 commonsourceibias.n913 commonsourceibias.n863 161.3
R7027 commonsourceibias.n912 commonsourceibias.n911 161.3
R7028 commonsourceibias.n909 commonsourceibias.n864 161.3
R7029 commonsourceibias.n908 commonsourceibias.n907 161.3
R7030 commonsourceibias.n906 commonsourceibias.n865 161.3
R7031 commonsourceibias.n905 commonsourceibias.n904 161.3
R7032 commonsourceibias.n902 commonsourceibias.n866 161.3
R7033 commonsourceibias.n900 commonsourceibias.n899 161.3
R7034 commonsourceibias.n898 commonsourceibias.n867 161.3
R7035 commonsourceibias.n897 commonsourceibias.n896 161.3
R7036 commonsourceibias.n894 commonsourceibias.n868 161.3
R7037 commonsourceibias.n893 commonsourceibias.n892 161.3
R7038 commonsourceibias.n891 commonsourceibias.n869 161.3
R7039 commonsourceibias.n890 commonsourceibias.n889 161.3
R7040 commonsourceibias.n887 commonsourceibias.n870 161.3
R7041 commonsourceibias.n885 commonsourceibias.n884 161.3
R7042 commonsourceibias.n883 commonsourceibias.n871 161.3
R7043 commonsourceibias.n882 commonsourceibias.n881 161.3
R7044 commonsourceibias.n879 commonsourceibias.n872 161.3
R7045 commonsourceibias.n878 commonsourceibias.n877 161.3
R7046 commonsourceibias.n876 commonsourceibias.n873 161.3
R7047 commonsourceibias.n846 commonsourceibias.n734 161.3
R7048 commonsourceibias.n844 commonsourceibias.n843 161.3
R7049 commonsourceibias.n842 commonsourceibias.n735 161.3
R7050 commonsourceibias.n841 commonsourceibias.n840 161.3
R7051 commonsourceibias.n838 commonsourceibias.n736 161.3
R7052 commonsourceibias.n837 commonsourceibias.n836 161.3
R7053 commonsourceibias.n835 commonsourceibias.n737 161.3
R7054 commonsourceibias.n834 commonsourceibias.n833 161.3
R7055 commonsourceibias.n831 commonsourceibias.n738 161.3
R7056 commonsourceibias.n829 commonsourceibias.n828 161.3
R7057 commonsourceibias.n827 commonsourceibias.n739 161.3
R7058 commonsourceibias.n826 commonsourceibias.n825 161.3
R7059 commonsourceibias.n823 commonsourceibias.n740 161.3
R7060 commonsourceibias.n822 commonsourceibias.n821 161.3
R7061 commonsourceibias.n820 commonsourceibias.n741 161.3
R7062 commonsourceibias.n819 commonsourceibias.n818 161.3
R7063 commonsourceibias.n816 commonsourceibias.n742 161.3
R7064 commonsourceibias.n814 commonsourceibias.n813 161.3
R7065 commonsourceibias.n812 commonsourceibias.n743 161.3
R7066 commonsourceibias.n811 commonsourceibias.n810 161.3
R7067 commonsourceibias.n808 commonsourceibias.n744 161.3
R7068 commonsourceibias.n807 commonsourceibias.n806 161.3
R7069 commonsourceibias.n805 commonsourceibias.n745 161.3
R7070 commonsourceibias.n804 commonsourceibias.n803 161.3
R7071 commonsourceibias.n801 commonsourceibias.n746 161.3
R7072 commonsourceibias.n799 commonsourceibias.n798 161.3
R7073 commonsourceibias.n797 commonsourceibias.n747 161.3
R7074 commonsourceibias.n796 commonsourceibias.n795 161.3
R7075 commonsourceibias.n793 commonsourceibias.n748 161.3
R7076 commonsourceibias.n792 commonsourceibias.n791 161.3
R7077 commonsourceibias.n790 commonsourceibias.n749 161.3
R7078 commonsourceibias.n789 commonsourceibias.n788 161.3
R7079 commonsourceibias.n786 commonsourceibias.n750 161.3
R7080 commonsourceibias.n784 commonsourceibias.n783 161.3
R7081 commonsourceibias.n782 commonsourceibias.n751 161.3
R7082 commonsourceibias.n781 commonsourceibias.n780 161.3
R7083 commonsourceibias.n778 commonsourceibias.n752 161.3
R7084 commonsourceibias.n777 commonsourceibias.n776 161.3
R7085 commonsourceibias.n775 commonsourceibias.n753 161.3
R7086 commonsourceibias.n774 commonsourceibias.n773 161.3
R7087 commonsourceibias.n771 commonsourceibias.n754 161.3
R7088 commonsourceibias.n769 commonsourceibias.n768 161.3
R7089 commonsourceibias.n767 commonsourceibias.n755 161.3
R7090 commonsourceibias.n766 commonsourceibias.n765 161.3
R7091 commonsourceibias.n763 commonsourceibias.n756 161.3
R7092 commonsourceibias.n762 commonsourceibias.n761 161.3
R7093 commonsourceibias.n760 commonsourceibias.n757 161.3
R7094 commonsourceibias.n616 commonsourceibias.n504 161.3
R7095 commonsourceibias.n614 commonsourceibias.n613 161.3
R7096 commonsourceibias.n612 commonsourceibias.n505 161.3
R7097 commonsourceibias.n611 commonsourceibias.n610 161.3
R7098 commonsourceibias.n608 commonsourceibias.n506 161.3
R7099 commonsourceibias.n607 commonsourceibias.n606 161.3
R7100 commonsourceibias.n605 commonsourceibias.n507 161.3
R7101 commonsourceibias.n604 commonsourceibias.n603 161.3
R7102 commonsourceibias.n601 commonsourceibias.n508 161.3
R7103 commonsourceibias.n599 commonsourceibias.n598 161.3
R7104 commonsourceibias.n597 commonsourceibias.n509 161.3
R7105 commonsourceibias.n596 commonsourceibias.n595 161.3
R7106 commonsourceibias.n593 commonsourceibias.n510 161.3
R7107 commonsourceibias.n592 commonsourceibias.n591 161.3
R7108 commonsourceibias.n590 commonsourceibias.n511 161.3
R7109 commonsourceibias.n589 commonsourceibias.n588 161.3
R7110 commonsourceibias.n586 commonsourceibias.n512 161.3
R7111 commonsourceibias.n584 commonsourceibias.n583 161.3
R7112 commonsourceibias.n582 commonsourceibias.n513 161.3
R7113 commonsourceibias.n581 commonsourceibias.n580 161.3
R7114 commonsourceibias.n578 commonsourceibias.n514 161.3
R7115 commonsourceibias.n577 commonsourceibias.n576 161.3
R7116 commonsourceibias.n575 commonsourceibias.n515 161.3
R7117 commonsourceibias.n574 commonsourceibias.n573 161.3
R7118 commonsourceibias.n571 commonsourceibias.n516 161.3
R7119 commonsourceibias.n569 commonsourceibias.n568 161.3
R7120 commonsourceibias.n567 commonsourceibias.n517 161.3
R7121 commonsourceibias.n566 commonsourceibias.n565 161.3
R7122 commonsourceibias.n563 commonsourceibias.n518 161.3
R7123 commonsourceibias.n562 commonsourceibias.n561 161.3
R7124 commonsourceibias.n560 commonsourceibias.n519 161.3
R7125 commonsourceibias.n559 commonsourceibias.n558 161.3
R7126 commonsourceibias.n556 commonsourceibias.n520 161.3
R7127 commonsourceibias.n554 commonsourceibias.n553 161.3
R7128 commonsourceibias.n552 commonsourceibias.n521 161.3
R7129 commonsourceibias.n551 commonsourceibias.n550 161.3
R7130 commonsourceibias.n548 commonsourceibias.n522 161.3
R7131 commonsourceibias.n547 commonsourceibias.n546 161.3
R7132 commonsourceibias.n545 commonsourceibias.n523 161.3
R7133 commonsourceibias.n544 commonsourceibias.n543 161.3
R7134 commonsourceibias.n541 commonsourceibias.n524 161.3
R7135 commonsourceibias.n539 commonsourceibias.n538 161.3
R7136 commonsourceibias.n537 commonsourceibias.n525 161.3
R7137 commonsourceibias.n536 commonsourceibias.n535 161.3
R7138 commonsourceibias.n533 commonsourceibias.n526 161.3
R7139 commonsourceibias.n532 commonsourceibias.n531 161.3
R7140 commonsourceibias.n530 commonsourceibias.n527 161.3
R7141 commonsourceibias.n686 commonsourceibias.n685 161.3
R7142 commonsourceibias.n684 commonsourceibias.n683 161.3
R7143 commonsourceibias.n682 commonsourceibias.n632 161.3
R7144 commonsourceibias.n681 commonsourceibias.n680 161.3
R7145 commonsourceibias.n679 commonsourceibias.n678 161.3
R7146 commonsourceibias.n677 commonsourceibias.n634 161.3
R7147 commonsourceibias.n676 commonsourceibias.n675 161.3
R7148 commonsourceibias.n674 commonsourceibias.n673 161.3
R7149 commonsourceibias.n672 commonsourceibias.n636 161.3
R7150 commonsourceibias.n670 commonsourceibias.n669 161.3
R7151 commonsourceibias.n668 commonsourceibias.n637 161.3
R7152 commonsourceibias.n667 commonsourceibias.n666 161.3
R7153 commonsourceibias.n664 commonsourceibias.n638 161.3
R7154 commonsourceibias.n663 commonsourceibias.n662 161.3
R7155 commonsourceibias.n661 commonsourceibias.n639 161.3
R7156 commonsourceibias.n660 commonsourceibias.n659 161.3
R7157 commonsourceibias.n657 commonsourceibias.n640 161.3
R7158 commonsourceibias.n655 commonsourceibias.n654 161.3
R7159 commonsourceibias.n653 commonsourceibias.n641 161.3
R7160 commonsourceibias.n652 commonsourceibias.n651 161.3
R7161 commonsourceibias.n649 commonsourceibias.n642 161.3
R7162 commonsourceibias.n648 commonsourceibias.n647 161.3
R7163 commonsourceibias.n646 commonsourceibias.n643 161.3
R7164 commonsourceibias.n731 commonsourceibias.n483 161.3
R7165 commonsourceibias.n729 commonsourceibias.n728 161.3
R7166 commonsourceibias.n727 commonsourceibias.n484 161.3
R7167 commonsourceibias.n726 commonsourceibias.n725 161.3
R7168 commonsourceibias.n723 commonsourceibias.n485 161.3
R7169 commonsourceibias.n722 commonsourceibias.n721 161.3
R7170 commonsourceibias.n720 commonsourceibias.n486 161.3
R7171 commonsourceibias.n719 commonsourceibias.n718 161.3
R7172 commonsourceibias.n716 commonsourceibias.n487 161.3
R7173 commonsourceibias.n714 commonsourceibias.n713 161.3
R7174 commonsourceibias.n712 commonsourceibias.n488 161.3
R7175 commonsourceibias.n711 commonsourceibias.n710 161.3
R7176 commonsourceibias.n708 commonsourceibias.n489 161.3
R7177 commonsourceibias.n707 commonsourceibias.n706 161.3
R7178 commonsourceibias.n705 commonsourceibias.n490 161.3
R7179 commonsourceibias.n704 commonsourceibias.n703 161.3
R7180 commonsourceibias.n701 commonsourceibias.n491 161.3
R7181 commonsourceibias.n699 commonsourceibias.n698 161.3
R7182 commonsourceibias.n697 commonsourceibias.n492 161.3
R7183 commonsourceibias.n696 commonsourceibias.n695 161.3
R7184 commonsourceibias.n693 commonsourceibias.n493 161.3
R7185 commonsourceibias.n692 commonsourceibias.n691 161.3
R7186 commonsourceibias.n690 commonsourceibias.n494 161.3
R7187 commonsourceibias.n689 commonsourceibias.n688 161.3
R7188 commonsourceibias.n141 commonsourceibias.n139 81.5057
R7189 commonsourceibias.n497 commonsourceibias.n495 81.5057
R7190 commonsourceibias.n141 commonsourceibias.n140 80.9324
R7191 commonsourceibias.n143 commonsourceibias.n142 80.9324
R7192 commonsourceibias.n145 commonsourceibias.n144 80.9324
R7193 commonsourceibias.n147 commonsourceibias.n146 80.9324
R7194 commonsourceibias.n138 commonsourceibias.n137 80.9324
R7195 commonsourceibias.n136 commonsourceibias.n135 80.9324
R7196 commonsourceibias.n134 commonsourceibias.n133 80.9324
R7197 commonsourceibias.n132 commonsourceibias.n131 80.9324
R7198 commonsourceibias.n130 commonsourceibias.n129 80.9324
R7199 commonsourceibias.n620 commonsourceibias.n619 80.9324
R7200 commonsourceibias.n622 commonsourceibias.n621 80.9324
R7201 commonsourceibias.n624 commonsourceibias.n623 80.9324
R7202 commonsourceibias.n626 commonsourceibias.n625 80.9324
R7203 commonsourceibias.n628 commonsourceibias.n627 80.9324
R7204 commonsourceibias.n503 commonsourceibias.n502 80.9324
R7205 commonsourceibias.n501 commonsourceibias.n500 80.9324
R7206 commonsourceibias.n499 commonsourceibias.n498 80.9324
R7207 commonsourceibias.n497 commonsourceibias.n496 80.9324
R7208 commonsourceibias.n481 commonsourceibias.n480 80.6037
R7209 commonsourceibias.n365 commonsourceibias.n364 80.6037
R7210 commonsourceibias.n128 commonsourceibias.n127 80.6037
R7211 commonsourceibias.n250 commonsourceibias.n249 80.6037
R7212 commonsourceibias.n964 commonsourceibias.n963 80.6037
R7213 commonsourceibias.n848 commonsourceibias.n847 80.6037
R7214 commonsourceibias.n618 commonsourceibias.n617 80.6037
R7215 commonsourceibias.n733 commonsourceibias.n732 80.6037
R7216 commonsourceibias.n438 commonsourceibias.n437 56.5617
R7217 commonsourceibias.n452 commonsourceibias.n451 56.5617
R7218 commonsourceibias.n322 commonsourceibias.n321 56.5617
R7219 commonsourceibias.n308 commonsourceibias.n307 56.5617
R7220 commonsourceibias.n85 commonsourceibias.n84 56.5617
R7221 commonsourceibias.n71 commonsourceibias.n70 56.5617
R7222 commonsourceibias.n207 commonsourceibias.n206 56.5617
R7223 commonsourceibias.n193 commonsourceibias.n192 56.5617
R7224 commonsourceibias.n919 commonsourceibias.n917 56.5617
R7225 commonsourceibias.n934 commonsourceibias.n932 56.5617
R7226 commonsourceibias.n803 commonsourceibias.n801 56.5617
R7227 commonsourceibias.n818 commonsourceibias.n816 56.5617
R7228 commonsourceibias.n573 commonsourceibias.n571 56.5617
R7229 commonsourceibias.n588 commonsourceibias.n586 56.5617
R7230 commonsourceibias.n688 commonsourceibias.n686 56.5617
R7231 commonsourceibias.n410 commonsourceibias.n409 56.5617
R7232 commonsourceibias.n424 commonsourceibias.n423 56.5617
R7233 commonsourceibias.n466 commonsourceibias.n465 56.5617
R7234 commonsourceibias.n350 commonsourceibias.n349 56.5617
R7235 commonsourceibias.n336 commonsourceibias.n335 56.5617
R7236 commonsourceibias.n294 commonsourceibias.n293 56.5617
R7237 commonsourceibias.n113 commonsourceibias.n112 56.5617
R7238 commonsourceibias.n99 commonsourceibias.n98 56.5617
R7239 commonsourceibias.n57 commonsourceibias.n56 56.5617
R7240 commonsourceibias.n235 commonsourceibias.n234 56.5617
R7241 commonsourceibias.n221 commonsourceibias.n220 56.5617
R7242 commonsourceibias.n179 commonsourceibias.n178 56.5617
R7243 commonsourceibias.n889 commonsourceibias.n887 56.5617
R7244 commonsourceibias.n904 commonsourceibias.n902 56.5617
R7245 commonsourceibias.n949 commonsourceibias.n947 56.5617
R7246 commonsourceibias.n773 commonsourceibias.n771 56.5617
R7247 commonsourceibias.n788 commonsourceibias.n786 56.5617
R7248 commonsourceibias.n833 commonsourceibias.n831 56.5617
R7249 commonsourceibias.n543 commonsourceibias.n541 56.5617
R7250 commonsourceibias.n558 commonsourceibias.n556 56.5617
R7251 commonsourceibias.n603 commonsourceibias.n601 56.5617
R7252 commonsourceibias.n718 commonsourceibias.n716 56.5617
R7253 commonsourceibias.n703 commonsourceibias.n701 56.5617
R7254 commonsourceibias.n659 commonsourceibias.n657 56.5617
R7255 commonsourceibias.n673 commonsourceibias.n672 56.5617
R7256 commonsourceibias.n401 commonsourceibias.n400 51.2335
R7257 commonsourceibias.n473 commonsourceibias.n368 51.2335
R7258 commonsourceibias.n357 commonsourceibias.n252 51.2335
R7259 commonsourceibias.n285 commonsourceibias.n284 51.2335
R7260 commonsourceibias.n120 commonsourceibias.n15 51.2335
R7261 commonsourceibias.n48 commonsourceibias.n47 51.2335
R7262 commonsourceibias.n242 commonsourceibias.n1 51.2335
R7263 commonsourceibias.n170 commonsourceibias.n169 51.2335
R7264 commonsourceibias.n879 commonsourceibias.n878 51.2335
R7265 commonsourceibias.n956 commonsourceibias.n851 51.2335
R7266 commonsourceibias.n763 commonsourceibias.n762 51.2335
R7267 commonsourceibias.n840 commonsourceibias.n735 51.2335
R7268 commonsourceibias.n533 commonsourceibias.n532 51.2335
R7269 commonsourceibias.n610 commonsourceibias.n505 51.2335
R7270 commonsourceibias.n725 commonsourceibias.n484 51.2335
R7271 commonsourceibias.n649 commonsourceibias.n648 51.2335
R7272 commonsourceibias.n480 commonsourceibias.n479 50.9056
R7273 commonsourceibias.n364 commonsourceibias.n363 50.9056
R7274 commonsourceibias.n127 commonsourceibias.n126 50.9056
R7275 commonsourceibias.n249 commonsourceibias.n248 50.9056
R7276 commonsourceibias.n963 commonsourceibias.n962 50.9056
R7277 commonsourceibias.n847 commonsourceibias.n846 50.9056
R7278 commonsourceibias.n617 commonsourceibias.n616 50.9056
R7279 commonsourceibias.n732 commonsourceibias.n731 50.9056
R7280 commonsourceibias.n415 commonsourceibias.n414 50.2647
R7281 commonsourceibias.n459 commonsourceibias.n373 50.2647
R7282 commonsourceibias.n343 commonsourceibias.n257 50.2647
R7283 commonsourceibias.n299 commonsourceibias.n298 50.2647
R7284 commonsourceibias.n106 commonsourceibias.n20 50.2647
R7285 commonsourceibias.n62 commonsourceibias.n61 50.2647
R7286 commonsourceibias.n228 commonsourceibias.n6 50.2647
R7287 commonsourceibias.n184 commonsourceibias.n183 50.2647
R7288 commonsourceibias.n894 commonsourceibias.n893 50.2647
R7289 commonsourceibias.n941 commonsourceibias.n855 50.2647
R7290 commonsourceibias.n778 commonsourceibias.n777 50.2647
R7291 commonsourceibias.n825 commonsourceibias.n739 50.2647
R7292 commonsourceibias.n548 commonsourceibias.n547 50.2647
R7293 commonsourceibias.n595 commonsourceibias.n509 50.2647
R7294 commonsourceibias.n710 commonsourceibias.n488 50.2647
R7295 commonsourceibias.n664 commonsourceibias.n663 50.2647
R7296 commonsourceibias.n397 commonsourceibias.n396 49.9027
R7297 commonsourceibias.n281 commonsourceibias.n280 49.9027
R7298 commonsourceibias.n44 commonsourceibias.n43 49.9027
R7299 commonsourceibias.n166 commonsourceibias.n165 49.9027
R7300 commonsourceibias.n875 commonsourceibias.n874 49.9027
R7301 commonsourceibias.n759 commonsourceibias.n758 49.9027
R7302 commonsourceibias.n529 commonsourceibias.n528 49.9027
R7303 commonsourceibias.n645 commonsourceibias.n644 49.9027
R7304 commonsourceibias.n429 commonsourceibias.n428 49.296
R7305 commonsourceibias.n445 commonsourceibias.n378 49.296
R7306 commonsourceibias.n329 commonsourceibias.n262 49.296
R7307 commonsourceibias.n313 commonsourceibias.n312 49.296
R7308 commonsourceibias.n92 commonsourceibias.n25 49.296
R7309 commonsourceibias.n76 commonsourceibias.n75 49.296
R7310 commonsourceibias.n214 commonsourceibias.n11 49.296
R7311 commonsourceibias.n198 commonsourceibias.n197 49.296
R7312 commonsourceibias.n909 commonsourceibias.n908 49.296
R7313 commonsourceibias.n926 commonsourceibias.n859 49.296
R7314 commonsourceibias.n793 commonsourceibias.n792 49.296
R7315 commonsourceibias.n810 commonsourceibias.n743 49.296
R7316 commonsourceibias.n563 commonsourceibias.n562 49.296
R7317 commonsourceibias.n580 commonsourceibias.n513 49.296
R7318 commonsourceibias.n695 commonsourceibias.n492 49.296
R7319 commonsourceibias.n678 commonsourceibias.n677 49.296
R7320 commonsourceibias.n431 commonsourceibias.n383 48.3272
R7321 commonsourceibias.n443 commonsourceibias.n442 48.3272
R7322 commonsourceibias.n327 commonsourceibias.n326 48.3272
R7323 commonsourceibias.n315 commonsourceibias.n267 48.3272
R7324 commonsourceibias.n90 commonsourceibias.n89 48.3272
R7325 commonsourceibias.n78 commonsourceibias.n30 48.3272
R7326 commonsourceibias.n212 commonsourceibias.n211 48.3272
R7327 commonsourceibias.n202 commonsourceibias.n201 48.3272
R7328 commonsourceibias.n911 commonsourceibias.n863 48.3272
R7329 commonsourceibias.n924 commonsourceibias.n923 48.3272
R7330 commonsourceibias.n795 commonsourceibias.n747 48.3272
R7331 commonsourceibias.n808 commonsourceibias.n807 48.3272
R7332 commonsourceibias.n565 commonsourceibias.n517 48.3272
R7333 commonsourceibias.n578 commonsourceibias.n577 48.3272
R7334 commonsourceibias.n693 commonsourceibias.n692 48.3272
R7335 commonsourceibias.n682 commonsourceibias.n681 48.3272
R7336 commonsourceibias.n417 commonsourceibias.n388 47.3584
R7337 commonsourceibias.n457 commonsourceibias.n456 47.3584
R7338 commonsourceibias.n341 commonsourceibias.n340 47.3584
R7339 commonsourceibias.n301 commonsourceibias.n272 47.3584
R7340 commonsourceibias.n104 commonsourceibias.n103 47.3584
R7341 commonsourceibias.n64 commonsourceibias.n35 47.3584
R7342 commonsourceibias.n226 commonsourceibias.n225 47.3584
R7343 commonsourceibias.n186 commonsourceibias.n157 47.3584
R7344 commonsourceibias.n896 commonsourceibias.n867 47.3584
R7345 commonsourceibias.n939 commonsourceibias.n938 47.3584
R7346 commonsourceibias.n780 commonsourceibias.n751 47.3584
R7347 commonsourceibias.n823 commonsourceibias.n822 47.3584
R7348 commonsourceibias.n550 commonsourceibias.n521 47.3584
R7349 commonsourceibias.n593 commonsourceibias.n592 47.3584
R7350 commonsourceibias.n708 commonsourceibias.n707 47.3584
R7351 commonsourceibias.n666 commonsourceibias.n637 47.3584
R7352 commonsourceibias.n403 commonsourceibias.n393 46.3896
R7353 commonsourceibias.n471 commonsourceibias.n470 46.3896
R7354 commonsourceibias.n355 commonsourceibias.n354 46.3896
R7355 commonsourceibias.n287 commonsourceibias.n277 46.3896
R7356 commonsourceibias.n118 commonsourceibias.n117 46.3896
R7357 commonsourceibias.n50 commonsourceibias.n40 46.3896
R7358 commonsourceibias.n240 commonsourceibias.n239 46.3896
R7359 commonsourceibias.n172 commonsourceibias.n162 46.3896
R7360 commonsourceibias.n881 commonsourceibias.n871 46.3896
R7361 commonsourceibias.n954 commonsourceibias.n953 46.3896
R7362 commonsourceibias.n765 commonsourceibias.n755 46.3896
R7363 commonsourceibias.n838 commonsourceibias.n837 46.3896
R7364 commonsourceibias.n535 commonsourceibias.n525 46.3896
R7365 commonsourceibias.n608 commonsourceibias.n607 46.3896
R7366 commonsourceibias.n723 commonsourceibias.n722 46.3896
R7367 commonsourceibias.n651 commonsourceibias.n641 46.3896
R7368 commonsourceibias.n398 commonsourceibias.n397 44.7059
R7369 commonsourceibias.n876 commonsourceibias.n875 44.7059
R7370 commonsourceibias.n760 commonsourceibias.n759 44.7059
R7371 commonsourceibias.n530 commonsourceibias.n529 44.7059
R7372 commonsourceibias.n646 commonsourceibias.n645 44.7059
R7373 commonsourceibias.n282 commonsourceibias.n281 44.7059
R7374 commonsourceibias.n45 commonsourceibias.n44 44.7059
R7375 commonsourceibias.n167 commonsourceibias.n166 44.7059
R7376 commonsourceibias.n407 commonsourceibias.n393 34.7644
R7377 commonsourceibias.n470 commonsourceibias.n370 34.7644
R7378 commonsourceibias.n354 commonsourceibias.n254 34.7644
R7379 commonsourceibias.n291 commonsourceibias.n277 34.7644
R7380 commonsourceibias.n117 commonsourceibias.n17 34.7644
R7381 commonsourceibias.n54 commonsourceibias.n40 34.7644
R7382 commonsourceibias.n239 commonsourceibias.n3 34.7644
R7383 commonsourceibias.n176 commonsourceibias.n162 34.7644
R7384 commonsourceibias.n885 commonsourceibias.n871 34.7644
R7385 commonsourceibias.n953 commonsourceibias.n853 34.7644
R7386 commonsourceibias.n769 commonsourceibias.n755 34.7644
R7387 commonsourceibias.n837 commonsourceibias.n737 34.7644
R7388 commonsourceibias.n539 commonsourceibias.n525 34.7644
R7389 commonsourceibias.n607 commonsourceibias.n507 34.7644
R7390 commonsourceibias.n722 commonsourceibias.n486 34.7644
R7391 commonsourceibias.n655 commonsourceibias.n641 34.7644
R7392 commonsourceibias.n421 commonsourceibias.n388 33.7956
R7393 commonsourceibias.n456 commonsourceibias.n375 33.7956
R7394 commonsourceibias.n340 commonsourceibias.n259 33.7956
R7395 commonsourceibias.n305 commonsourceibias.n272 33.7956
R7396 commonsourceibias.n103 commonsourceibias.n22 33.7956
R7397 commonsourceibias.n68 commonsourceibias.n35 33.7956
R7398 commonsourceibias.n225 commonsourceibias.n8 33.7956
R7399 commonsourceibias.n190 commonsourceibias.n157 33.7956
R7400 commonsourceibias.n900 commonsourceibias.n867 33.7956
R7401 commonsourceibias.n938 commonsourceibias.n857 33.7956
R7402 commonsourceibias.n784 commonsourceibias.n751 33.7956
R7403 commonsourceibias.n822 commonsourceibias.n741 33.7956
R7404 commonsourceibias.n554 commonsourceibias.n521 33.7956
R7405 commonsourceibias.n592 commonsourceibias.n511 33.7956
R7406 commonsourceibias.n707 commonsourceibias.n490 33.7956
R7407 commonsourceibias.n670 commonsourceibias.n637 33.7956
R7408 commonsourceibias.n435 commonsourceibias.n383 32.8269
R7409 commonsourceibias.n442 commonsourceibias.n380 32.8269
R7410 commonsourceibias.n326 commonsourceibias.n264 32.8269
R7411 commonsourceibias.n319 commonsourceibias.n267 32.8269
R7412 commonsourceibias.n89 commonsourceibias.n27 32.8269
R7413 commonsourceibias.n82 commonsourceibias.n30 32.8269
R7414 commonsourceibias.n211 commonsourceibias.n13 32.8269
R7415 commonsourceibias.n203 commonsourceibias.n202 32.8269
R7416 commonsourceibias.n915 commonsourceibias.n863 32.8269
R7417 commonsourceibias.n923 commonsourceibias.n861 32.8269
R7418 commonsourceibias.n799 commonsourceibias.n747 32.8269
R7419 commonsourceibias.n807 commonsourceibias.n745 32.8269
R7420 commonsourceibias.n569 commonsourceibias.n517 32.8269
R7421 commonsourceibias.n577 commonsourceibias.n515 32.8269
R7422 commonsourceibias.n692 commonsourceibias.n494 32.8269
R7423 commonsourceibias.n683 commonsourceibias.n682 32.8269
R7424 commonsourceibias.n428 commonsourceibias.n385 31.8581
R7425 commonsourceibias.n449 commonsourceibias.n378 31.8581
R7426 commonsourceibias.n333 commonsourceibias.n262 31.8581
R7427 commonsourceibias.n312 commonsourceibias.n269 31.8581
R7428 commonsourceibias.n96 commonsourceibias.n25 31.8581
R7429 commonsourceibias.n75 commonsourceibias.n32 31.8581
R7430 commonsourceibias.n218 commonsourceibias.n11 31.8581
R7431 commonsourceibias.n197 commonsourceibias.n196 31.8581
R7432 commonsourceibias.n908 commonsourceibias.n865 31.8581
R7433 commonsourceibias.n930 commonsourceibias.n859 31.8581
R7434 commonsourceibias.n792 commonsourceibias.n749 31.8581
R7435 commonsourceibias.n814 commonsourceibias.n743 31.8581
R7436 commonsourceibias.n562 commonsourceibias.n519 31.8581
R7437 commonsourceibias.n584 commonsourceibias.n513 31.8581
R7438 commonsourceibias.n699 commonsourceibias.n492 31.8581
R7439 commonsourceibias.n677 commonsourceibias.n676 31.8581
R7440 commonsourceibias.n414 commonsourceibias.n390 30.8893
R7441 commonsourceibias.n463 commonsourceibias.n373 30.8893
R7442 commonsourceibias.n347 commonsourceibias.n257 30.8893
R7443 commonsourceibias.n298 commonsourceibias.n274 30.8893
R7444 commonsourceibias.n110 commonsourceibias.n20 30.8893
R7445 commonsourceibias.n61 commonsourceibias.n37 30.8893
R7446 commonsourceibias.n232 commonsourceibias.n6 30.8893
R7447 commonsourceibias.n183 commonsourceibias.n159 30.8893
R7448 commonsourceibias.n893 commonsourceibias.n869 30.8893
R7449 commonsourceibias.n945 commonsourceibias.n855 30.8893
R7450 commonsourceibias.n777 commonsourceibias.n753 30.8893
R7451 commonsourceibias.n829 commonsourceibias.n739 30.8893
R7452 commonsourceibias.n547 commonsourceibias.n523 30.8893
R7453 commonsourceibias.n599 commonsourceibias.n509 30.8893
R7454 commonsourceibias.n714 commonsourceibias.n488 30.8893
R7455 commonsourceibias.n663 commonsourceibias.n639 30.8893
R7456 commonsourceibias.n400 commonsourceibias.n395 29.9206
R7457 commonsourceibias.n477 commonsourceibias.n368 29.9206
R7458 commonsourceibias.n361 commonsourceibias.n252 29.9206
R7459 commonsourceibias.n284 commonsourceibias.n279 29.9206
R7460 commonsourceibias.n124 commonsourceibias.n15 29.9206
R7461 commonsourceibias.n47 commonsourceibias.n42 29.9206
R7462 commonsourceibias.n246 commonsourceibias.n1 29.9206
R7463 commonsourceibias.n169 commonsourceibias.n164 29.9206
R7464 commonsourceibias.n878 commonsourceibias.n873 29.9206
R7465 commonsourceibias.n960 commonsourceibias.n851 29.9206
R7466 commonsourceibias.n762 commonsourceibias.n757 29.9206
R7467 commonsourceibias.n844 commonsourceibias.n735 29.9206
R7468 commonsourceibias.n532 commonsourceibias.n527 29.9206
R7469 commonsourceibias.n614 commonsourceibias.n505 29.9206
R7470 commonsourceibias.n729 commonsourceibias.n484 29.9206
R7471 commonsourceibias.n648 commonsourceibias.n643 29.9206
R7472 commonsourceibias.n479 commonsourceibias.n478 21.8872
R7473 commonsourceibias.n363 commonsourceibias.n362 21.8872
R7474 commonsourceibias.n126 commonsourceibias.n125 21.8872
R7475 commonsourceibias.n248 commonsourceibias.n247 21.8872
R7476 commonsourceibias.n962 commonsourceibias.n961 21.8872
R7477 commonsourceibias.n846 commonsourceibias.n845 21.8872
R7478 commonsourceibias.n616 commonsourceibias.n615 21.8872
R7479 commonsourceibias.n731 commonsourceibias.n730 21.8872
R7480 commonsourceibias.n410 commonsourceibias.n392 21.3954
R7481 commonsourceibias.n465 commonsourceibias.n464 21.3954
R7482 commonsourceibias.n349 commonsourceibias.n348 21.3954
R7483 commonsourceibias.n294 commonsourceibias.n276 21.3954
R7484 commonsourceibias.n112 commonsourceibias.n111 21.3954
R7485 commonsourceibias.n57 commonsourceibias.n39 21.3954
R7486 commonsourceibias.n234 commonsourceibias.n233 21.3954
R7487 commonsourceibias.n179 commonsourceibias.n161 21.3954
R7488 commonsourceibias.n889 commonsourceibias.n888 21.3954
R7489 commonsourceibias.n947 commonsourceibias.n946 21.3954
R7490 commonsourceibias.n773 commonsourceibias.n772 21.3954
R7491 commonsourceibias.n831 commonsourceibias.n830 21.3954
R7492 commonsourceibias.n543 commonsourceibias.n542 21.3954
R7493 commonsourceibias.n601 commonsourceibias.n600 21.3954
R7494 commonsourceibias.n716 commonsourceibias.n715 21.3954
R7495 commonsourceibias.n659 commonsourceibias.n658 21.3954
R7496 commonsourceibias.n424 commonsourceibias.n387 20.9036
R7497 commonsourceibias.n451 commonsourceibias.n450 20.9036
R7498 commonsourceibias.n335 commonsourceibias.n334 20.9036
R7499 commonsourceibias.n308 commonsourceibias.n271 20.9036
R7500 commonsourceibias.n98 commonsourceibias.n97 20.9036
R7501 commonsourceibias.n71 commonsourceibias.n34 20.9036
R7502 commonsourceibias.n220 commonsourceibias.n219 20.9036
R7503 commonsourceibias.n193 commonsourceibias.n155 20.9036
R7504 commonsourceibias.n904 commonsourceibias.n903 20.9036
R7505 commonsourceibias.n932 commonsourceibias.n931 20.9036
R7506 commonsourceibias.n788 commonsourceibias.n787 20.9036
R7507 commonsourceibias.n816 commonsourceibias.n815 20.9036
R7508 commonsourceibias.n558 commonsourceibias.n557 20.9036
R7509 commonsourceibias.n586 commonsourceibias.n585 20.9036
R7510 commonsourceibias.n701 commonsourceibias.n700 20.9036
R7511 commonsourceibias.n673 commonsourceibias.n635 20.9036
R7512 commonsourceibias.n437 commonsourceibias.n436 20.4117
R7513 commonsourceibias.n438 commonsourceibias.n382 20.4117
R7514 commonsourceibias.n322 commonsourceibias.n266 20.4117
R7515 commonsourceibias.n321 commonsourceibias.n320 20.4117
R7516 commonsourceibias.n85 commonsourceibias.n29 20.4117
R7517 commonsourceibias.n84 commonsourceibias.n83 20.4117
R7518 commonsourceibias.n207 commonsourceibias.n150 20.4117
R7519 commonsourceibias.n206 commonsourceibias.n151 20.4117
R7520 commonsourceibias.n917 commonsourceibias.n916 20.4117
R7521 commonsourceibias.n919 commonsourceibias.n918 20.4117
R7522 commonsourceibias.n801 commonsourceibias.n800 20.4117
R7523 commonsourceibias.n803 commonsourceibias.n802 20.4117
R7524 commonsourceibias.n571 commonsourceibias.n570 20.4117
R7525 commonsourceibias.n573 commonsourceibias.n572 20.4117
R7526 commonsourceibias.n688 commonsourceibias.n687 20.4117
R7527 commonsourceibias.n686 commonsourceibias.n631 20.4117
R7528 commonsourceibias.n423 commonsourceibias.n422 19.9199
R7529 commonsourceibias.n452 commonsourceibias.n377 19.9199
R7530 commonsourceibias.n336 commonsourceibias.n261 19.9199
R7531 commonsourceibias.n307 commonsourceibias.n306 19.9199
R7532 commonsourceibias.n99 commonsourceibias.n24 19.9199
R7533 commonsourceibias.n70 commonsourceibias.n69 19.9199
R7534 commonsourceibias.n221 commonsourceibias.n10 19.9199
R7535 commonsourceibias.n192 commonsourceibias.n191 19.9199
R7536 commonsourceibias.n902 commonsourceibias.n901 19.9199
R7537 commonsourceibias.n934 commonsourceibias.n933 19.9199
R7538 commonsourceibias.n786 commonsourceibias.n785 19.9199
R7539 commonsourceibias.n818 commonsourceibias.n817 19.9199
R7540 commonsourceibias.n556 commonsourceibias.n555 19.9199
R7541 commonsourceibias.n588 commonsourceibias.n587 19.9199
R7542 commonsourceibias.n703 commonsourceibias.n702 19.9199
R7543 commonsourceibias.n672 commonsourceibias.n671 19.9199
R7544 commonsourceibias.n409 commonsourceibias.n408 19.4281
R7545 commonsourceibias.n466 commonsourceibias.n372 19.4281
R7546 commonsourceibias.n350 commonsourceibias.n256 19.4281
R7547 commonsourceibias.n293 commonsourceibias.n292 19.4281
R7548 commonsourceibias.n113 commonsourceibias.n19 19.4281
R7549 commonsourceibias.n56 commonsourceibias.n55 19.4281
R7550 commonsourceibias.n235 commonsourceibias.n5 19.4281
R7551 commonsourceibias.n178 commonsourceibias.n177 19.4281
R7552 commonsourceibias.n887 commonsourceibias.n886 19.4281
R7553 commonsourceibias.n949 commonsourceibias.n948 19.4281
R7554 commonsourceibias.n771 commonsourceibias.n770 19.4281
R7555 commonsourceibias.n833 commonsourceibias.n832 19.4281
R7556 commonsourceibias.n541 commonsourceibias.n540 19.4281
R7557 commonsourceibias.n603 commonsourceibias.n602 19.4281
R7558 commonsourceibias.n718 commonsourceibias.n717 19.4281
R7559 commonsourceibias.n657 commonsourceibias.n656 19.4281
R7560 commonsourceibias.n402 commonsourceibias.n401 13.526
R7561 commonsourceibias.n473 commonsourceibias.n472 13.526
R7562 commonsourceibias.n357 commonsourceibias.n356 13.526
R7563 commonsourceibias.n286 commonsourceibias.n285 13.526
R7564 commonsourceibias.n120 commonsourceibias.n119 13.526
R7565 commonsourceibias.n49 commonsourceibias.n48 13.526
R7566 commonsourceibias.n242 commonsourceibias.n241 13.526
R7567 commonsourceibias.n171 commonsourceibias.n170 13.526
R7568 commonsourceibias.n880 commonsourceibias.n879 13.526
R7569 commonsourceibias.n956 commonsourceibias.n955 13.526
R7570 commonsourceibias.n764 commonsourceibias.n763 13.526
R7571 commonsourceibias.n840 commonsourceibias.n839 13.526
R7572 commonsourceibias.n534 commonsourceibias.n533 13.526
R7573 commonsourceibias.n610 commonsourceibias.n609 13.526
R7574 commonsourceibias.n725 commonsourceibias.n724 13.526
R7575 commonsourceibias.n650 commonsourceibias.n649 13.526
R7576 commonsourceibias.n130 commonsourceibias.n128 13.2322
R7577 commonsourceibias.n620 commonsourceibias.n618 13.2322
R7578 commonsourceibias.n416 commonsourceibias.n415 13.0342
R7579 commonsourceibias.n459 commonsourceibias.n458 13.0342
R7580 commonsourceibias.n343 commonsourceibias.n342 13.0342
R7581 commonsourceibias.n300 commonsourceibias.n299 13.0342
R7582 commonsourceibias.n106 commonsourceibias.n105 13.0342
R7583 commonsourceibias.n63 commonsourceibias.n62 13.0342
R7584 commonsourceibias.n228 commonsourceibias.n227 13.0342
R7585 commonsourceibias.n185 commonsourceibias.n184 13.0342
R7586 commonsourceibias.n895 commonsourceibias.n894 13.0342
R7587 commonsourceibias.n941 commonsourceibias.n940 13.0342
R7588 commonsourceibias.n779 commonsourceibias.n778 13.0342
R7589 commonsourceibias.n825 commonsourceibias.n824 13.0342
R7590 commonsourceibias.n549 commonsourceibias.n548 13.0342
R7591 commonsourceibias.n595 commonsourceibias.n594 13.0342
R7592 commonsourceibias.n710 commonsourceibias.n709 13.0342
R7593 commonsourceibias.n665 commonsourceibias.n664 13.0342
R7594 commonsourceibias.n430 commonsourceibias.n429 12.5423
R7595 commonsourceibias.n445 commonsourceibias.n444 12.5423
R7596 commonsourceibias.n329 commonsourceibias.n328 12.5423
R7597 commonsourceibias.n314 commonsourceibias.n313 12.5423
R7598 commonsourceibias.n92 commonsourceibias.n91 12.5423
R7599 commonsourceibias.n77 commonsourceibias.n76 12.5423
R7600 commonsourceibias.n214 commonsourceibias.n213 12.5423
R7601 commonsourceibias.n198 commonsourceibias.n153 12.5423
R7602 commonsourceibias.n910 commonsourceibias.n909 12.5423
R7603 commonsourceibias.n926 commonsourceibias.n925 12.5423
R7604 commonsourceibias.n794 commonsourceibias.n793 12.5423
R7605 commonsourceibias.n810 commonsourceibias.n809 12.5423
R7606 commonsourceibias.n564 commonsourceibias.n563 12.5423
R7607 commonsourceibias.n580 commonsourceibias.n579 12.5423
R7608 commonsourceibias.n695 commonsourceibias.n694 12.5423
R7609 commonsourceibias.n678 commonsourceibias.n633 12.5423
R7610 commonsourceibias.n431 commonsourceibias.n430 12.0505
R7611 commonsourceibias.n444 commonsourceibias.n443 12.0505
R7612 commonsourceibias.n328 commonsourceibias.n327 12.0505
R7613 commonsourceibias.n315 commonsourceibias.n314 12.0505
R7614 commonsourceibias.n91 commonsourceibias.n90 12.0505
R7615 commonsourceibias.n78 commonsourceibias.n77 12.0505
R7616 commonsourceibias.n213 commonsourceibias.n212 12.0505
R7617 commonsourceibias.n201 commonsourceibias.n153 12.0505
R7618 commonsourceibias.n911 commonsourceibias.n910 12.0505
R7619 commonsourceibias.n925 commonsourceibias.n924 12.0505
R7620 commonsourceibias.n795 commonsourceibias.n794 12.0505
R7621 commonsourceibias.n809 commonsourceibias.n808 12.0505
R7622 commonsourceibias.n565 commonsourceibias.n564 12.0505
R7623 commonsourceibias.n579 commonsourceibias.n578 12.0505
R7624 commonsourceibias.n694 commonsourceibias.n693 12.0505
R7625 commonsourceibias.n681 commonsourceibias.n633 12.0505
R7626 commonsourceibias.n417 commonsourceibias.n416 11.5587
R7627 commonsourceibias.n458 commonsourceibias.n457 11.5587
R7628 commonsourceibias.n342 commonsourceibias.n341 11.5587
R7629 commonsourceibias.n301 commonsourceibias.n300 11.5587
R7630 commonsourceibias.n105 commonsourceibias.n104 11.5587
R7631 commonsourceibias.n64 commonsourceibias.n63 11.5587
R7632 commonsourceibias.n227 commonsourceibias.n226 11.5587
R7633 commonsourceibias.n186 commonsourceibias.n185 11.5587
R7634 commonsourceibias.n896 commonsourceibias.n895 11.5587
R7635 commonsourceibias.n940 commonsourceibias.n939 11.5587
R7636 commonsourceibias.n780 commonsourceibias.n779 11.5587
R7637 commonsourceibias.n824 commonsourceibias.n823 11.5587
R7638 commonsourceibias.n550 commonsourceibias.n549 11.5587
R7639 commonsourceibias.n594 commonsourceibias.n593 11.5587
R7640 commonsourceibias.n709 commonsourceibias.n708 11.5587
R7641 commonsourceibias.n666 commonsourceibias.n665 11.5587
R7642 commonsourceibias.n403 commonsourceibias.n402 11.0668
R7643 commonsourceibias.n472 commonsourceibias.n471 11.0668
R7644 commonsourceibias.n356 commonsourceibias.n355 11.0668
R7645 commonsourceibias.n287 commonsourceibias.n286 11.0668
R7646 commonsourceibias.n119 commonsourceibias.n118 11.0668
R7647 commonsourceibias.n50 commonsourceibias.n49 11.0668
R7648 commonsourceibias.n241 commonsourceibias.n240 11.0668
R7649 commonsourceibias.n172 commonsourceibias.n171 11.0668
R7650 commonsourceibias.n881 commonsourceibias.n880 11.0668
R7651 commonsourceibias.n955 commonsourceibias.n954 11.0668
R7652 commonsourceibias.n765 commonsourceibias.n764 11.0668
R7653 commonsourceibias.n839 commonsourceibias.n838 11.0668
R7654 commonsourceibias.n535 commonsourceibias.n534 11.0668
R7655 commonsourceibias.n609 commonsourceibias.n608 11.0668
R7656 commonsourceibias.n724 commonsourceibias.n723 11.0668
R7657 commonsourceibias.n651 commonsourceibias.n650 11.0668
R7658 commonsourceibias.n966 commonsourceibias.n482 10.122
R7659 commonsourceibias.n149 commonsourceibias.n148 9.50363
R7660 commonsourceibias.n630 commonsourceibias.n629 9.50363
R7661 commonsourceibias.n366 commonsourceibias.n250 8.76042
R7662 commonsourceibias.n849 commonsourceibias.n733 8.76042
R7663 commonsourceibias.n966 commonsourceibias.n965 8.46921
R7664 commonsourceibias.n408 commonsourceibias.n407 5.16479
R7665 commonsourceibias.n372 commonsourceibias.n370 5.16479
R7666 commonsourceibias.n256 commonsourceibias.n254 5.16479
R7667 commonsourceibias.n292 commonsourceibias.n291 5.16479
R7668 commonsourceibias.n19 commonsourceibias.n17 5.16479
R7669 commonsourceibias.n55 commonsourceibias.n54 5.16479
R7670 commonsourceibias.n5 commonsourceibias.n3 5.16479
R7671 commonsourceibias.n177 commonsourceibias.n176 5.16479
R7672 commonsourceibias.n886 commonsourceibias.n885 5.16479
R7673 commonsourceibias.n948 commonsourceibias.n853 5.16479
R7674 commonsourceibias.n770 commonsourceibias.n769 5.16479
R7675 commonsourceibias.n832 commonsourceibias.n737 5.16479
R7676 commonsourceibias.n540 commonsourceibias.n539 5.16479
R7677 commonsourceibias.n602 commonsourceibias.n507 5.16479
R7678 commonsourceibias.n717 commonsourceibias.n486 5.16479
R7679 commonsourceibias.n656 commonsourceibias.n655 5.16479
R7680 commonsourceibias.n482 commonsourceibias.n481 5.03125
R7681 commonsourceibias.n366 commonsourceibias.n365 5.03125
R7682 commonsourceibias.n965 commonsourceibias.n964 5.03125
R7683 commonsourceibias.n849 commonsourceibias.n848 5.03125
R7684 commonsourceibias.n422 commonsourceibias.n421 4.67295
R7685 commonsourceibias.n377 commonsourceibias.n375 4.67295
R7686 commonsourceibias.n261 commonsourceibias.n259 4.67295
R7687 commonsourceibias.n306 commonsourceibias.n305 4.67295
R7688 commonsourceibias.n24 commonsourceibias.n22 4.67295
R7689 commonsourceibias.n69 commonsourceibias.n68 4.67295
R7690 commonsourceibias.n10 commonsourceibias.n8 4.67295
R7691 commonsourceibias.n191 commonsourceibias.n190 4.67295
R7692 commonsourceibias.n901 commonsourceibias.n900 4.67295
R7693 commonsourceibias.n933 commonsourceibias.n857 4.67295
R7694 commonsourceibias.n785 commonsourceibias.n784 4.67295
R7695 commonsourceibias.n817 commonsourceibias.n741 4.67295
R7696 commonsourceibias.n555 commonsourceibias.n554 4.67295
R7697 commonsourceibias.n587 commonsourceibias.n511 4.67295
R7698 commonsourceibias.n702 commonsourceibias.n490 4.67295
R7699 commonsourceibias.n671 commonsourceibias.n670 4.67295
R7700 commonsourceibias commonsourceibias.n966 4.20978
R7701 commonsourceibias.n436 commonsourceibias.n435 4.18111
R7702 commonsourceibias.n382 commonsourceibias.n380 4.18111
R7703 commonsourceibias.n266 commonsourceibias.n264 4.18111
R7704 commonsourceibias.n320 commonsourceibias.n319 4.18111
R7705 commonsourceibias.n29 commonsourceibias.n27 4.18111
R7706 commonsourceibias.n83 commonsourceibias.n82 4.18111
R7707 commonsourceibias.n150 commonsourceibias.n13 4.18111
R7708 commonsourceibias.n203 commonsourceibias.n151 4.18111
R7709 commonsourceibias.n916 commonsourceibias.n915 4.18111
R7710 commonsourceibias.n918 commonsourceibias.n861 4.18111
R7711 commonsourceibias.n800 commonsourceibias.n799 4.18111
R7712 commonsourceibias.n802 commonsourceibias.n745 4.18111
R7713 commonsourceibias.n570 commonsourceibias.n569 4.18111
R7714 commonsourceibias.n572 commonsourceibias.n515 4.18111
R7715 commonsourceibias.n687 commonsourceibias.n494 4.18111
R7716 commonsourceibias.n683 commonsourceibias.n631 4.18111
R7717 commonsourceibias.n482 commonsourceibias.n366 3.72967
R7718 commonsourceibias.n965 commonsourceibias.n849 3.72967
R7719 commonsourceibias.n387 commonsourceibias.n385 3.68928
R7720 commonsourceibias.n450 commonsourceibias.n449 3.68928
R7721 commonsourceibias.n334 commonsourceibias.n333 3.68928
R7722 commonsourceibias.n271 commonsourceibias.n269 3.68928
R7723 commonsourceibias.n97 commonsourceibias.n96 3.68928
R7724 commonsourceibias.n34 commonsourceibias.n32 3.68928
R7725 commonsourceibias.n219 commonsourceibias.n218 3.68928
R7726 commonsourceibias.n196 commonsourceibias.n155 3.68928
R7727 commonsourceibias.n903 commonsourceibias.n865 3.68928
R7728 commonsourceibias.n931 commonsourceibias.n930 3.68928
R7729 commonsourceibias.n787 commonsourceibias.n749 3.68928
R7730 commonsourceibias.n815 commonsourceibias.n814 3.68928
R7731 commonsourceibias.n557 commonsourceibias.n519 3.68928
R7732 commonsourceibias.n585 commonsourceibias.n584 3.68928
R7733 commonsourceibias.n700 commonsourceibias.n699 3.68928
R7734 commonsourceibias.n676 commonsourceibias.n635 3.68928
R7735 commonsourceibias.n392 commonsourceibias.n390 3.19744
R7736 commonsourceibias.n464 commonsourceibias.n463 3.19744
R7737 commonsourceibias.n348 commonsourceibias.n347 3.19744
R7738 commonsourceibias.n276 commonsourceibias.n274 3.19744
R7739 commonsourceibias.n111 commonsourceibias.n110 3.19744
R7740 commonsourceibias.n39 commonsourceibias.n37 3.19744
R7741 commonsourceibias.n233 commonsourceibias.n232 3.19744
R7742 commonsourceibias.n161 commonsourceibias.n159 3.19744
R7743 commonsourceibias.n888 commonsourceibias.n869 3.19744
R7744 commonsourceibias.n946 commonsourceibias.n945 3.19744
R7745 commonsourceibias.n772 commonsourceibias.n753 3.19744
R7746 commonsourceibias.n830 commonsourceibias.n829 3.19744
R7747 commonsourceibias.n542 commonsourceibias.n523 3.19744
R7748 commonsourceibias.n600 commonsourceibias.n599 3.19744
R7749 commonsourceibias.n715 commonsourceibias.n714 3.19744
R7750 commonsourceibias.n658 commonsourceibias.n639 3.19744
R7751 commonsourceibias.n139 commonsourceibias.t5 2.82907
R7752 commonsourceibias.n139 commonsourceibias.t23 2.82907
R7753 commonsourceibias.n140 commonsourceibias.t43 2.82907
R7754 commonsourceibias.n140 commonsourceibias.t29 2.82907
R7755 commonsourceibias.n142 commonsourceibias.t7 2.82907
R7756 commonsourceibias.n142 commonsourceibias.t15 2.82907
R7757 commonsourceibias.n144 commonsourceibias.t79 2.82907
R7758 commonsourceibias.n144 commonsourceibias.t19 2.82907
R7759 commonsourceibias.n146 commonsourceibias.t51 2.82907
R7760 commonsourceibias.n146 commonsourceibias.t25 2.82907
R7761 commonsourceibias.n137 commonsourceibias.t69 2.82907
R7762 commonsourceibias.n137 commonsourceibias.t31 2.82907
R7763 commonsourceibias.n135 commonsourceibias.t55 2.82907
R7764 commonsourceibias.n135 commonsourceibias.t61 2.82907
R7765 commonsourceibias.n133 commonsourceibias.t3 2.82907
R7766 commonsourceibias.n133 commonsourceibias.t71 2.82907
R7767 commonsourceibias.n131 commonsourceibias.t59 2.82907
R7768 commonsourceibias.n131 commonsourceibias.t65 2.82907
R7769 commonsourceibias.n129 commonsourceibias.t67 2.82907
R7770 commonsourceibias.n129 commonsourceibias.t11 2.82907
R7771 commonsourceibias.n619 commonsourceibias.t1 2.82907
R7772 commonsourceibias.n619 commonsourceibias.t41 2.82907
R7773 commonsourceibias.n621 commonsourceibias.t39 2.82907
R7774 commonsourceibias.n621 commonsourceibias.t21 2.82907
R7775 commonsourceibias.n623 commonsourceibias.t45 2.82907
R7776 commonsourceibias.n623 commonsourceibias.t33 2.82907
R7777 commonsourceibias.n625 commonsourceibias.t53 2.82907
R7778 commonsourceibias.n625 commonsourceibias.t9 2.82907
R7779 commonsourceibias.n627 commonsourceibias.t35 2.82907
R7780 commonsourceibias.n627 commonsourceibias.t37 2.82907
R7781 commonsourceibias.n502 commonsourceibias.t73 2.82907
R7782 commonsourceibias.n502 commonsourceibias.t27 2.82907
R7783 commonsourceibias.n500 commonsourceibias.t47 2.82907
R7784 commonsourceibias.n500 commonsourceibias.t57 2.82907
R7785 commonsourceibias.n498 commonsourceibias.t49 2.82907
R7786 commonsourceibias.n498 commonsourceibias.t13 2.82907
R7787 commonsourceibias.n496 commonsourceibias.t63 2.82907
R7788 commonsourceibias.n496 commonsourceibias.t75 2.82907
R7789 commonsourceibias.n495 commonsourceibias.t77 2.82907
R7790 commonsourceibias.n495 commonsourceibias.t17 2.82907
R7791 commonsourceibias.n396 commonsourceibias.n395 2.7056
R7792 commonsourceibias.n478 commonsourceibias.n477 2.7056
R7793 commonsourceibias.n362 commonsourceibias.n361 2.7056
R7794 commonsourceibias.n280 commonsourceibias.n279 2.7056
R7795 commonsourceibias.n125 commonsourceibias.n124 2.7056
R7796 commonsourceibias.n43 commonsourceibias.n42 2.7056
R7797 commonsourceibias.n247 commonsourceibias.n246 2.7056
R7798 commonsourceibias.n165 commonsourceibias.n164 2.7056
R7799 commonsourceibias.n874 commonsourceibias.n873 2.7056
R7800 commonsourceibias.n961 commonsourceibias.n960 2.7056
R7801 commonsourceibias.n758 commonsourceibias.n757 2.7056
R7802 commonsourceibias.n845 commonsourceibias.n844 2.7056
R7803 commonsourceibias.n528 commonsourceibias.n527 2.7056
R7804 commonsourceibias.n615 commonsourceibias.n614 2.7056
R7805 commonsourceibias.n730 commonsourceibias.n729 2.7056
R7806 commonsourceibias.n644 commonsourceibias.n643 2.7056
R7807 commonsourceibias.n132 commonsourceibias.n130 0.573776
R7808 commonsourceibias.n134 commonsourceibias.n132 0.573776
R7809 commonsourceibias.n136 commonsourceibias.n134 0.573776
R7810 commonsourceibias.n138 commonsourceibias.n136 0.573776
R7811 commonsourceibias.n147 commonsourceibias.n145 0.573776
R7812 commonsourceibias.n145 commonsourceibias.n143 0.573776
R7813 commonsourceibias.n143 commonsourceibias.n141 0.573776
R7814 commonsourceibias.n499 commonsourceibias.n497 0.573776
R7815 commonsourceibias.n501 commonsourceibias.n499 0.573776
R7816 commonsourceibias.n503 commonsourceibias.n501 0.573776
R7817 commonsourceibias.n628 commonsourceibias.n626 0.573776
R7818 commonsourceibias.n626 commonsourceibias.n624 0.573776
R7819 commonsourceibias.n624 commonsourceibias.n622 0.573776
R7820 commonsourceibias.n622 commonsourceibias.n620 0.573776
R7821 commonsourceibias.n148 commonsourceibias.n138 0.287138
R7822 commonsourceibias.n148 commonsourceibias.n147 0.287138
R7823 commonsourceibias.n629 commonsourceibias.n503 0.287138
R7824 commonsourceibias.n629 commonsourceibias.n628 0.287138
R7825 commonsourceibias.n481 commonsourceibias.n367 0.285035
R7826 commonsourceibias.n365 commonsourceibias.n251 0.285035
R7827 commonsourceibias.n128 commonsourceibias.n14 0.285035
R7828 commonsourceibias.n250 commonsourceibias.n0 0.285035
R7829 commonsourceibias.n964 commonsourceibias.n850 0.285035
R7830 commonsourceibias.n848 commonsourceibias.n734 0.285035
R7831 commonsourceibias.n618 commonsourceibias.n504 0.285035
R7832 commonsourceibias.n733 commonsourceibias.n483 0.285035
R7833 commonsourceibias.n476 commonsourceibias.n367 0.189894
R7834 commonsourceibias.n476 commonsourceibias.n475 0.189894
R7835 commonsourceibias.n475 commonsourceibias.n474 0.189894
R7836 commonsourceibias.n474 commonsourceibias.n369 0.189894
R7837 commonsourceibias.n469 commonsourceibias.n369 0.189894
R7838 commonsourceibias.n469 commonsourceibias.n468 0.189894
R7839 commonsourceibias.n468 commonsourceibias.n467 0.189894
R7840 commonsourceibias.n467 commonsourceibias.n371 0.189894
R7841 commonsourceibias.n462 commonsourceibias.n371 0.189894
R7842 commonsourceibias.n462 commonsourceibias.n461 0.189894
R7843 commonsourceibias.n461 commonsourceibias.n460 0.189894
R7844 commonsourceibias.n460 commonsourceibias.n374 0.189894
R7845 commonsourceibias.n455 commonsourceibias.n374 0.189894
R7846 commonsourceibias.n455 commonsourceibias.n454 0.189894
R7847 commonsourceibias.n454 commonsourceibias.n453 0.189894
R7848 commonsourceibias.n453 commonsourceibias.n376 0.189894
R7849 commonsourceibias.n448 commonsourceibias.n376 0.189894
R7850 commonsourceibias.n448 commonsourceibias.n447 0.189894
R7851 commonsourceibias.n447 commonsourceibias.n446 0.189894
R7852 commonsourceibias.n446 commonsourceibias.n379 0.189894
R7853 commonsourceibias.n441 commonsourceibias.n379 0.189894
R7854 commonsourceibias.n441 commonsourceibias.n440 0.189894
R7855 commonsourceibias.n440 commonsourceibias.n439 0.189894
R7856 commonsourceibias.n439 commonsourceibias.n381 0.189894
R7857 commonsourceibias.n434 commonsourceibias.n381 0.189894
R7858 commonsourceibias.n434 commonsourceibias.n433 0.189894
R7859 commonsourceibias.n433 commonsourceibias.n432 0.189894
R7860 commonsourceibias.n432 commonsourceibias.n384 0.189894
R7861 commonsourceibias.n427 commonsourceibias.n384 0.189894
R7862 commonsourceibias.n427 commonsourceibias.n426 0.189894
R7863 commonsourceibias.n426 commonsourceibias.n425 0.189894
R7864 commonsourceibias.n425 commonsourceibias.n386 0.189894
R7865 commonsourceibias.n420 commonsourceibias.n386 0.189894
R7866 commonsourceibias.n420 commonsourceibias.n419 0.189894
R7867 commonsourceibias.n419 commonsourceibias.n418 0.189894
R7868 commonsourceibias.n418 commonsourceibias.n389 0.189894
R7869 commonsourceibias.n413 commonsourceibias.n389 0.189894
R7870 commonsourceibias.n413 commonsourceibias.n412 0.189894
R7871 commonsourceibias.n412 commonsourceibias.n411 0.189894
R7872 commonsourceibias.n411 commonsourceibias.n391 0.189894
R7873 commonsourceibias.n406 commonsourceibias.n391 0.189894
R7874 commonsourceibias.n406 commonsourceibias.n405 0.189894
R7875 commonsourceibias.n405 commonsourceibias.n404 0.189894
R7876 commonsourceibias.n404 commonsourceibias.n394 0.189894
R7877 commonsourceibias.n399 commonsourceibias.n394 0.189894
R7878 commonsourceibias.n399 commonsourceibias.n398 0.189894
R7879 commonsourceibias.n360 commonsourceibias.n251 0.189894
R7880 commonsourceibias.n360 commonsourceibias.n359 0.189894
R7881 commonsourceibias.n359 commonsourceibias.n358 0.189894
R7882 commonsourceibias.n358 commonsourceibias.n253 0.189894
R7883 commonsourceibias.n353 commonsourceibias.n253 0.189894
R7884 commonsourceibias.n353 commonsourceibias.n352 0.189894
R7885 commonsourceibias.n352 commonsourceibias.n351 0.189894
R7886 commonsourceibias.n351 commonsourceibias.n255 0.189894
R7887 commonsourceibias.n346 commonsourceibias.n255 0.189894
R7888 commonsourceibias.n346 commonsourceibias.n345 0.189894
R7889 commonsourceibias.n345 commonsourceibias.n344 0.189894
R7890 commonsourceibias.n344 commonsourceibias.n258 0.189894
R7891 commonsourceibias.n339 commonsourceibias.n258 0.189894
R7892 commonsourceibias.n339 commonsourceibias.n338 0.189894
R7893 commonsourceibias.n338 commonsourceibias.n337 0.189894
R7894 commonsourceibias.n337 commonsourceibias.n260 0.189894
R7895 commonsourceibias.n332 commonsourceibias.n260 0.189894
R7896 commonsourceibias.n332 commonsourceibias.n331 0.189894
R7897 commonsourceibias.n331 commonsourceibias.n330 0.189894
R7898 commonsourceibias.n330 commonsourceibias.n263 0.189894
R7899 commonsourceibias.n325 commonsourceibias.n263 0.189894
R7900 commonsourceibias.n325 commonsourceibias.n324 0.189894
R7901 commonsourceibias.n324 commonsourceibias.n323 0.189894
R7902 commonsourceibias.n323 commonsourceibias.n265 0.189894
R7903 commonsourceibias.n318 commonsourceibias.n265 0.189894
R7904 commonsourceibias.n318 commonsourceibias.n317 0.189894
R7905 commonsourceibias.n317 commonsourceibias.n316 0.189894
R7906 commonsourceibias.n316 commonsourceibias.n268 0.189894
R7907 commonsourceibias.n311 commonsourceibias.n268 0.189894
R7908 commonsourceibias.n311 commonsourceibias.n310 0.189894
R7909 commonsourceibias.n310 commonsourceibias.n309 0.189894
R7910 commonsourceibias.n309 commonsourceibias.n270 0.189894
R7911 commonsourceibias.n304 commonsourceibias.n270 0.189894
R7912 commonsourceibias.n304 commonsourceibias.n303 0.189894
R7913 commonsourceibias.n303 commonsourceibias.n302 0.189894
R7914 commonsourceibias.n302 commonsourceibias.n273 0.189894
R7915 commonsourceibias.n297 commonsourceibias.n273 0.189894
R7916 commonsourceibias.n297 commonsourceibias.n296 0.189894
R7917 commonsourceibias.n296 commonsourceibias.n295 0.189894
R7918 commonsourceibias.n295 commonsourceibias.n275 0.189894
R7919 commonsourceibias.n290 commonsourceibias.n275 0.189894
R7920 commonsourceibias.n290 commonsourceibias.n289 0.189894
R7921 commonsourceibias.n289 commonsourceibias.n288 0.189894
R7922 commonsourceibias.n288 commonsourceibias.n278 0.189894
R7923 commonsourceibias.n283 commonsourceibias.n278 0.189894
R7924 commonsourceibias.n283 commonsourceibias.n282 0.189894
R7925 commonsourceibias.n123 commonsourceibias.n14 0.189894
R7926 commonsourceibias.n123 commonsourceibias.n122 0.189894
R7927 commonsourceibias.n122 commonsourceibias.n121 0.189894
R7928 commonsourceibias.n121 commonsourceibias.n16 0.189894
R7929 commonsourceibias.n116 commonsourceibias.n16 0.189894
R7930 commonsourceibias.n116 commonsourceibias.n115 0.189894
R7931 commonsourceibias.n115 commonsourceibias.n114 0.189894
R7932 commonsourceibias.n114 commonsourceibias.n18 0.189894
R7933 commonsourceibias.n109 commonsourceibias.n18 0.189894
R7934 commonsourceibias.n109 commonsourceibias.n108 0.189894
R7935 commonsourceibias.n108 commonsourceibias.n107 0.189894
R7936 commonsourceibias.n107 commonsourceibias.n21 0.189894
R7937 commonsourceibias.n102 commonsourceibias.n21 0.189894
R7938 commonsourceibias.n102 commonsourceibias.n101 0.189894
R7939 commonsourceibias.n101 commonsourceibias.n100 0.189894
R7940 commonsourceibias.n100 commonsourceibias.n23 0.189894
R7941 commonsourceibias.n95 commonsourceibias.n23 0.189894
R7942 commonsourceibias.n95 commonsourceibias.n94 0.189894
R7943 commonsourceibias.n94 commonsourceibias.n93 0.189894
R7944 commonsourceibias.n93 commonsourceibias.n26 0.189894
R7945 commonsourceibias.n88 commonsourceibias.n26 0.189894
R7946 commonsourceibias.n88 commonsourceibias.n87 0.189894
R7947 commonsourceibias.n87 commonsourceibias.n86 0.189894
R7948 commonsourceibias.n86 commonsourceibias.n28 0.189894
R7949 commonsourceibias.n81 commonsourceibias.n28 0.189894
R7950 commonsourceibias.n81 commonsourceibias.n80 0.189894
R7951 commonsourceibias.n80 commonsourceibias.n79 0.189894
R7952 commonsourceibias.n79 commonsourceibias.n31 0.189894
R7953 commonsourceibias.n74 commonsourceibias.n31 0.189894
R7954 commonsourceibias.n74 commonsourceibias.n73 0.189894
R7955 commonsourceibias.n73 commonsourceibias.n72 0.189894
R7956 commonsourceibias.n72 commonsourceibias.n33 0.189894
R7957 commonsourceibias.n67 commonsourceibias.n33 0.189894
R7958 commonsourceibias.n67 commonsourceibias.n66 0.189894
R7959 commonsourceibias.n66 commonsourceibias.n65 0.189894
R7960 commonsourceibias.n65 commonsourceibias.n36 0.189894
R7961 commonsourceibias.n60 commonsourceibias.n36 0.189894
R7962 commonsourceibias.n60 commonsourceibias.n59 0.189894
R7963 commonsourceibias.n59 commonsourceibias.n58 0.189894
R7964 commonsourceibias.n58 commonsourceibias.n38 0.189894
R7965 commonsourceibias.n53 commonsourceibias.n38 0.189894
R7966 commonsourceibias.n53 commonsourceibias.n52 0.189894
R7967 commonsourceibias.n52 commonsourceibias.n51 0.189894
R7968 commonsourceibias.n51 commonsourceibias.n41 0.189894
R7969 commonsourceibias.n46 commonsourceibias.n41 0.189894
R7970 commonsourceibias.n46 commonsourceibias.n45 0.189894
R7971 commonsourceibias.n205 commonsourceibias.n204 0.189894
R7972 commonsourceibias.n204 commonsourceibias.n152 0.189894
R7973 commonsourceibias.n200 commonsourceibias.n152 0.189894
R7974 commonsourceibias.n200 commonsourceibias.n199 0.189894
R7975 commonsourceibias.n199 commonsourceibias.n154 0.189894
R7976 commonsourceibias.n195 commonsourceibias.n154 0.189894
R7977 commonsourceibias.n195 commonsourceibias.n194 0.189894
R7978 commonsourceibias.n194 commonsourceibias.n156 0.189894
R7979 commonsourceibias.n189 commonsourceibias.n156 0.189894
R7980 commonsourceibias.n189 commonsourceibias.n188 0.189894
R7981 commonsourceibias.n188 commonsourceibias.n187 0.189894
R7982 commonsourceibias.n187 commonsourceibias.n158 0.189894
R7983 commonsourceibias.n182 commonsourceibias.n158 0.189894
R7984 commonsourceibias.n182 commonsourceibias.n181 0.189894
R7985 commonsourceibias.n181 commonsourceibias.n180 0.189894
R7986 commonsourceibias.n180 commonsourceibias.n160 0.189894
R7987 commonsourceibias.n175 commonsourceibias.n160 0.189894
R7988 commonsourceibias.n175 commonsourceibias.n174 0.189894
R7989 commonsourceibias.n174 commonsourceibias.n173 0.189894
R7990 commonsourceibias.n173 commonsourceibias.n163 0.189894
R7991 commonsourceibias.n168 commonsourceibias.n163 0.189894
R7992 commonsourceibias.n168 commonsourceibias.n167 0.189894
R7993 commonsourceibias.n245 commonsourceibias.n0 0.189894
R7994 commonsourceibias.n245 commonsourceibias.n244 0.189894
R7995 commonsourceibias.n244 commonsourceibias.n243 0.189894
R7996 commonsourceibias.n243 commonsourceibias.n2 0.189894
R7997 commonsourceibias.n238 commonsourceibias.n2 0.189894
R7998 commonsourceibias.n238 commonsourceibias.n237 0.189894
R7999 commonsourceibias.n237 commonsourceibias.n236 0.189894
R8000 commonsourceibias.n236 commonsourceibias.n4 0.189894
R8001 commonsourceibias.n231 commonsourceibias.n4 0.189894
R8002 commonsourceibias.n231 commonsourceibias.n230 0.189894
R8003 commonsourceibias.n230 commonsourceibias.n229 0.189894
R8004 commonsourceibias.n229 commonsourceibias.n7 0.189894
R8005 commonsourceibias.n224 commonsourceibias.n7 0.189894
R8006 commonsourceibias.n224 commonsourceibias.n223 0.189894
R8007 commonsourceibias.n223 commonsourceibias.n222 0.189894
R8008 commonsourceibias.n222 commonsourceibias.n9 0.189894
R8009 commonsourceibias.n217 commonsourceibias.n9 0.189894
R8010 commonsourceibias.n217 commonsourceibias.n216 0.189894
R8011 commonsourceibias.n216 commonsourceibias.n215 0.189894
R8012 commonsourceibias.n215 commonsourceibias.n12 0.189894
R8013 commonsourceibias.n210 commonsourceibias.n12 0.189894
R8014 commonsourceibias.n210 commonsourceibias.n209 0.189894
R8015 commonsourceibias.n209 commonsourceibias.n208 0.189894
R8016 commonsourceibias.n877 commonsourceibias.n876 0.189894
R8017 commonsourceibias.n877 commonsourceibias.n872 0.189894
R8018 commonsourceibias.n882 commonsourceibias.n872 0.189894
R8019 commonsourceibias.n883 commonsourceibias.n882 0.189894
R8020 commonsourceibias.n884 commonsourceibias.n883 0.189894
R8021 commonsourceibias.n884 commonsourceibias.n870 0.189894
R8022 commonsourceibias.n890 commonsourceibias.n870 0.189894
R8023 commonsourceibias.n891 commonsourceibias.n890 0.189894
R8024 commonsourceibias.n892 commonsourceibias.n891 0.189894
R8025 commonsourceibias.n892 commonsourceibias.n868 0.189894
R8026 commonsourceibias.n897 commonsourceibias.n868 0.189894
R8027 commonsourceibias.n898 commonsourceibias.n897 0.189894
R8028 commonsourceibias.n899 commonsourceibias.n898 0.189894
R8029 commonsourceibias.n899 commonsourceibias.n866 0.189894
R8030 commonsourceibias.n905 commonsourceibias.n866 0.189894
R8031 commonsourceibias.n906 commonsourceibias.n905 0.189894
R8032 commonsourceibias.n907 commonsourceibias.n906 0.189894
R8033 commonsourceibias.n907 commonsourceibias.n864 0.189894
R8034 commonsourceibias.n912 commonsourceibias.n864 0.189894
R8035 commonsourceibias.n913 commonsourceibias.n912 0.189894
R8036 commonsourceibias.n914 commonsourceibias.n913 0.189894
R8037 commonsourceibias.n914 commonsourceibias.n862 0.189894
R8038 commonsourceibias.n920 commonsourceibias.n862 0.189894
R8039 commonsourceibias.n921 commonsourceibias.n920 0.189894
R8040 commonsourceibias.n922 commonsourceibias.n921 0.189894
R8041 commonsourceibias.n922 commonsourceibias.n860 0.189894
R8042 commonsourceibias.n927 commonsourceibias.n860 0.189894
R8043 commonsourceibias.n928 commonsourceibias.n927 0.189894
R8044 commonsourceibias.n929 commonsourceibias.n928 0.189894
R8045 commonsourceibias.n929 commonsourceibias.n858 0.189894
R8046 commonsourceibias.n935 commonsourceibias.n858 0.189894
R8047 commonsourceibias.n936 commonsourceibias.n935 0.189894
R8048 commonsourceibias.n937 commonsourceibias.n936 0.189894
R8049 commonsourceibias.n937 commonsourceibias.n856 0.189894
R8050 commonsourceibias.n942 commonsourceibias.n856 0.189894
R8051 commonsourceibias.n943 commonsourceibias.n942 0.189894
R8052 commonsourceibias.n944 commonsourceibias.n943 0.189894
R8053 commonsourceibias.n944 commonsourceibias.n854 0.189894
R8054 commonsourceibias.n950 commonsourceibias.n854 0.189894
R8055 commonsourceibias.n951 commonsourceibias.n950 0.189894
R8056 commonsourceibias.n952 commonsourceibias.n951 0.189894
R8057 commonsourceibias.n952 commonsourceibias.n852 0.189894
R8058 commonsourceibias.n957 commonsourceibias.n852 0.189894
R8059 commonsourceibias.n958 commonsourceibias.n957 0.189894
R8060 commonsourceibias.n959 commonsourceibias.n958 0.189894
R8061 commonsourceibias.n959 commonsourceibias.n850 0.189894
R8062 commonsourceibias.n761 commonsourceibias.n760 0.189894
R8063 commonsourceibias.n761 commonsourceibias.n756 0.189894
R8064 commonsourceibias.n766 commonsourceibias.n756 0.189894
R8065 commonsourceibias.n767 commonsourceibias.n766 0.189894
R8066 commonsourceibias.n768 commonsourceibias.n767 0.189894
R8067 commonsourceibias.n768 commonsourceibias.n754 0.189894
R8068 commonsourceibias.n774 commonsourceibias.n754 0.189894
R8069 commonsourceibias.n775 commonsourceibias.n774 0.189894
R8070 commonsourceibias.n776 commonsourceibias.n775 0.189894
R8071 commonsourceibias.n776 commonsourceibias.n752 0.189894
R8072 commonsourceibias.n781 commonsourceibias.n752 0.189894
R8073 commonsourceibias.n782 commonsourceibias.n781 0.189894
R8074 commonsourceibias.n783 commonsourceibias.n782 0.189894
R8075 commonsourceibias.n783 commonsourceibias.n750 0.189894
R8076 commonsourceibias.n789 commonsourceibias.n750 0.189894
R8077 commonsourceibias.n790 commonsourceibias.n789 0.189894
R8078 commonsourceibias.n791 commonsourceibias.n790 0.189894
R8079 commonsourceibias.n791 commonsourceibias.n748 0.189894
R8080 commonsourceibias.n796 commonsourceibias.n748 0.189894
R8081 commonsourceibias.n797 commonsourceibias.n796 0.189894
R8082 commonsourceibias.n798 commonsourceibias.n797 0.189894
R8083 commonsourceibias.n798 commonsourceibias.n746 0.189894
R8084 commonsourceibias.n804 commonsourceibias.n746 0.189894
R8085 commonsourceibias.n805 commonsourceibias.n804 0.189894
R8086 commonsourceibias.n806 commonsourceibias.n805 0.189894
R8087 commonsourceibias.n806 commonsourceibias.n744 0.189894
R8088 commonsourceibias.n811 commonsourceibias.n744 0.189894
R8089 commonsourceibias.n812 commonsourceibias.n811 0.189894
R8090 commonsourceibias.n813 commonsourceibias.n812 0.189894
R8091 commonsourceibias.n813 commonsourceibias.n742 0.189894
R8092 commonsourceibias.n819 commonsourceibias.n742 0.189894
R8093 commonsourceibias.n820 commonsourceibias.n819 0.189894
R8094 commonsourceibias.n821 commonsourceibias.n820 0.189894
R8095 commonsourceibias.n821 commonsourceibias.n740 0.189894
R8096 commonsourceibias.n826 commonsourceibias.n740 0.189894
R8097 commonsourceibias.n827 commonsourceibias.n826 0.189894
R8098 commonsourceibias.n828 commonsourceibias.n827 0.189894
R8099 commonsourceibias.n828 commonsourceibias.n738 0.189894
R8100 commonsourceibias.n834 commonsourceibias.n738 0.189894
R8101 commonsourceibias.n835 commonsourceibias.n834 0.189894
R8102 commonsourceibias.n836 commonsourceibias.n835 0.189894
R8103 commonsourceibias.n836 commonsourceibias.n736 0.189894
R8104 commonsourceibias.n841 commonsourceibias.n736 0.189894
R8105 commonsourceibias.n842 commonsourceibias.n841 0.189894
R8106 commonsourceibias.n843 commonsourceibias.n842 0.189894
R8107 commonsourceibias.n843 commonsourceibias.n734 0.189894
R8108 commonsourceibias.n531 commonsourceibias.n530 0.189894
R8109 commonsourceibias.n531 commonsourceibias.n526 0.189894
R8110 commonsourceibias.n536 commonsourceibias.n526 0.189894
R8111 commonsourceibias.n537 commonsourceibias.n536 0.189894
R8112 commonsourceibias.n538 commonsourceibias.n537 0.189894
R8113 commonsourceibias.n538 commonsourceibias.n524 0.189894
R8114 commonsourceibias.n544 commonsourceibias.n524 0.189894
R8115 commonsourceibias.n545 commonsourceibias.n544 0.189894
R8116 commonsourceibias.n546 commonsourceibias.n545 0.189894
R8117 commonsourceibias.n546 commonsourceibias.n522 0.189894
R8118 commonsourceibias.n551 commonsourceibias.n522 0.189894
R8119 commonsourceibias.n552 commonsourceibias.n551 0.189894
R8120 commonsourceibias.n553 commonsourceibias.n552 0.189894
R8121 commonsourceibias.n553 commonsourceibias.n520 0.189894
R8122 commonsourceibias.n559 commonsourceibias.n520 0.189894
R8123 commonsourceibias.n560 commonsourceibias.n559 0.189894
R8124 commonsourceibias.n561 commonsourceibias.n560 0.189894
R8125 commonsourceibias.n561 commonsourceibias.n518 0.189894
R8126 commonsourceibias.n566 commonsourceibias.n518 0.189894
R8127 commonsourceibias.n567 commonsourceibias.n566 0.189894
R8128 commonsourceibias.n568 commonsourceibias.n567 0.189894
R8129 commonsourceibias.n568 commonsourceibias.n516 0.189894
R8130 commonsourceibias.n574 commonsourceibias.n516 0.189894
R8131 commonsourceibias.n575 commonsourceibias.n574 0.189894
R8132 commonsourceibias.n576 commonsourceibias.n575 0.189894
R8133 commonsourceibias.n576 commonsourceibias.n514 0.189894
R8134 commonsourceibias.n581 commonsourceibias.n514 0.189894
R8135 commonsourceibias.n582 commonsourceibias.n581 0.189894
R8136 commonsourceibias.n583 commonsourceibias.n582 0.189894
R8137 commonsourceibias.n583 commonsourceibias.n512 0.189894
R8138 commonsourceibias.n589 commonsourceibias.n512 0.189894
R8139 commonsourceibias.n590 commonsourceibias.n589 0.189894
R8140 commonsourceibias.n591 commonsourceibias.n590 0.189894
R8141 commonsourceibias.n591 commonsourceibias.n510 0.189894
R8142 commonsourceibias.n596 commonsourceibias.n510 0.189894
R8143 commonsourceibias.n597 commonsourceibias.n596 0.189894
R8144 commonsourceibias.n598 commonsourceibias.n597 0.189894
R8145 commonsourceibias.n598 commonsourceibias.n508 0.189894
R8146 commonsourceibias.n604 commonsourceibias.n508 0.189894
R8147 commonsourceibias.n605 commonsourceibias.n604 0.189894
R8148 commonsourceibias.n606 commonsourceibias.n605 0.189894
R8149 commonsourceibias.n606 commonsourceibias.n506 0.189894
R8150 commonsourceibias.n611 commonsourceibias.n506 0.189894
R8151 commonsourceibias.n612 commonsourceibias.n611 0.189894
R8152 commonsourceibias.n613 commonsourceibias.n612 0.189894
R8153 commonsourceibias.n613 commonsourceibias.n504 0.189894
R8154 commonsourceibias.n647 commonsourceibias.n646 0.189894
R8155 commonsourceibias.n647 commonsourceibias.n642 0.189894
R8156 commonsourceibias.n652 commonsourceibias.n642 0.189894
R8157 commonsourceibias.n653 commonsourceibias.n652 0.189894
R8158 commonsourceibias.n654 commonsourceibias.n653 0.189894
R8159 commonsourceibias.n654 commonsourceibias.n640 0.189894
R8160 commonsourceibias.n660 commonsourceibias.n640 0.189894
R8161 commonsourceibias.n661 commonsourceibias.n660 0.189894
R8162 commonsourceibias.n662 commonsourceibias.n661 0.189894
R8163 commonsourceibias.n662 commonsourceibias.n638 0.189894
R8164 commonsourceibias.n667 commonsourceibias.n638 0.189894
R8165 commonsourceibias.n668 commonsourceibias.n667 0.189894
R8166 commonsourceibias.n669 commonsourceibias.n668 0.189894
R8167 commonsourceibias.n669 commonsourceibias.n636 0.189894
R8168 commonsourceibias.n674 commonsourceibias.n636 0.189894
R8169 commonsourceibias.n675 commonsourceibias.n674 0.189894
R8170 commonsourceibias.n675 commonsourceibias.n634 0.189894
R8171 commonsourceibias.n679 commonsourceibias.n634 0.189894
R8172 commonsourceibias.n680 commonsourceibias.n679 0.189894
R8173 commonsourceibias.n680 commonsourceibias.n632 0.189894
R8174 commonsourceibias.n684 commonsourceibias.n632 0.189894
R8175 commonsourceibias.n685 commonsourceibias.n684 0.189894
R8176 commonsourceibias.n690 commonsourceibias.n689 0.189894
R8177 commonsourceibias.n691 commonsourceibias.n690 0.189894
R8178 commonsourceibias.n691 commonsourceibias.n493 0.189894
R8179 commonsourceibias.n696 commonsourceibias.n493 0.189894
R8180 commonsourceibias.n697 commonsourceibias.n696 0.189894
R8181 commonsourceibias.n698 commonsourceibias.n697 0.189894
R8182 commonsourceibias.n698 commonsourceibias.n491 0.189894
R8183 commonsourceibias.n704 commonsourceibias.n491 0.189894
R8184 commonsourceibias.n705 commonsourceibias.n704 0.189894
R8185 commonsourceibias.n706 commonsourceibias.n705 0.189894
R8186 commonsourceibias.n706 commonsourceibias.n489 0.189894
R8187 commonsourceibias.n711 commonsourceibias.n489 0.189894
R8188 commonsourceibias.n712 commonsourceibias.n711 0.189894
R8189 commonsourceibias.n713 commonsourceibias.n712 0.189894
R8190 commonsourceibias.n713 commonsourceibias.n487 0.189894
R8191 commonsourceibias.n719 commonsourceibias.n487 0.189894
R8192 commonsourceibias.n720 commonsourceibias.n719 0.189894
R8193 commonsourceibias.n721 commonsourceibias.n720 0.189894
R8194 commonsourceibias.n721 commonsourceibias.n485 0.189894
R8195 commonsourceibias.n726 commonsourceibias.n485 0.189894
R8196 commonsourceibias.n727 commonsourceibias.n726 0.189894
R8197 commonsourceibias.n728 commonsourceibias.n727 0.189894
R8198 commonsourceibias.n728 commonsourceibias.n483 0.189894
R8199 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R8200 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R8201 commonsourceibias.n685 commonsourceibias.n630 0.0762576
R8202 commonsourceibias.n689 commonsourceibias.n630 0.0762576
R8203 gnd.n7496 gnd.n493 1564.47
R8204 gnd.n6792 gnd.n6745 939.716
R8205 gnd.n4493 gnd.n4492 771.183
R8206 gnd.n6201 gnd.n3010 771.183
R8207 gnd.n4773 gnd.n3926 771.183
R8208 gnd.n6203 gnd.n3005 771.183
R8209 gnd.n6807 gnd.n1006 766.379
R8210 gnd.n2354 gnd.n1003 766.379
R8211 gnd.n1625 gnd.n1528 766.379
R8212 gnd.n1621 gnd.n1526 766.379
R8213 gnd.n6791 gnd.n1000 756.769
R8214 gnd.n6802 gnd.n6801 756.769
R8215 gnd.n1718 gnd.n1435 756.769
R8216 gnd.n1716 gnd.n1438 756.769
R8217 gnd.n257 gnd.n246 751.963
R8218 gnd.n7795 gnd.n7794 751.963
R8219 gnd.n3186 gnd.n3074 751.963
R8220 gnd.n6012 gnd.n3188 751.963
R8221 gnd.n2766 gnd.n2754 751.963
R8222 gnd.n4766 gnd.n4765 751.963
R8223 gnd.n4164 gnd.n2393 751.963
R8224 gnd.n4120 gnd.n4119 751.963
R8225 gnd.n7004 gnd.n785 703.915
R8226 gnd.n7495 gnd.n494 703.915
R8227 gnd.n7709 gnd.n7707 703.915
R8228 gnd.n4230 gnd.n4223 703.915
R8229 gnd.n7974 gnd.n250 696.707
R8230 gnd.n7850 gnd.n7849 696.707
R8231 gnd.n6015 gnd.n6014 696.707
R8232 gnd.n6132 gnd.n3120 696.707
R8233 gnd.n6445 gnd.n2759 696.707
R8234 gnd.n4715 gnd.n3957 696.707
R8235 gnd.n6623 gnd.n2466 696.707
R8236 gnd.n6743 gnd.n2397 696.707
R8237 gnd.n7004 gnd.n7003 585
R8238 gnd.n7005 gnd.n7004 585
R8239 gnd.n7002 gnd.n787 585
R8240 gnd.n787 gnd.n786 585
R8241 gnd.n7001 gnd.n7000 585
R8242 gnd.n7000 gnd.n6999 585
R8243 gnd.n792 gnd.n791 585
R8244 gnd.n6998 gnd.n792 585
R8245 gnd.n6996 gnd.n6995 585
R8246 gnd.n6997 gnd.n6996 585
R8247 gnd.n6994 gnd.n794 585
R8248 gnd.n794 gnd.n793 585
R8249 gnd.n6993 gnd.n6992 585
R8250 gnd.n6992 gnd.n6991 585
R8251 gnd.n800 gnd.n799 585
R8252 gnd.n6990 gnd.n800 585
R8253 gnd.n6988 gnd.n6987 585
R8254 gnd.n6989 gnd.n6988 585
R8255 gnd.n6986 gnd.n802 585
R8256 gnd.n802 gnd.n801 585
R8257 gnd.n6985 gnd.n6984 585
R8258 gnd.n6984 gnd.n6983 585
R8259 gnd.n808 gnd.n807 585
R8260 gnd.n6982 gnd.n808 585
R8261 gnd.n6980 gnd.n6979 585
R8262 gnd.n6981 gnd.n6980 585
R8263 gnd.n6978 gnd.n810 585
R8264 gnd.n810 gnd.n809 585
R8265 gnd.n6977 gnd.n6976 585
R8266 gnd.n6976 gnd.n6975 585
R8267 gnd.n816 gnd.n815 585
R8268 gnd.n6974 gnd.n816 585
R8269 gnd.n6972 gnd.n6971 585
R8270 gnd.n6973 gnd.n6972 585
R8271 gnd.n6970 gnd.n818 585
R8272 gnd.n818 gnd.n817 585
R8273 gnd.n6969 gnd.n6968 585
R8274 gnd.n6968 gnd.n6967 585
R8275 gnd.n824 gnd.n823 585
R8276 gnd.n6966 gnd.n824 585
R8277 gnd.n6964 gnd.n6963 585
R8278 gnd.n6965 gnd.n6964 585
R8279 gnd.n6962 gnd.n826 585
R8280 gnd.n826 gnd.n825 585
R8281 gnd.n6961 gnd.n6960 585
R8282 gnd.n6960 gnd.n6959 585
R8283 gnd.n832 gnd.n831 585
R8284 gnd.n6958 gnd.n832 585
R8285 gnd.n6956 gnd.n6955 585
R8286 gnd.n6957 gnd.n6956 585
R8287 gnd.n6954 gnd.n834 585
R8288 gnd.n834 gnd.n833 585
R8289 gnd.n6953 gnd.n6952 585
R8290 gnd.n6952 gnd.n6951 585
R8291 gnd.n840 gnd.n839 585
R8292 gnd.n6950 gnd.n840 585
R8293 gnd.n6948 gnd.n6947 585
R8294 gnd.n6949 gnd.n6948 585
R8295 gnd.n6946 gnd.n842 585
R8296 gnd.n842 gnd.n841 585
R8297 gnd.n6945 gnd.n6944 585
R8298 gnd.n6944 gnd.n6943 585
R8299 gnd.n848 gnd.n847 585
R8300 gnd.n6942 gnd.n848 585
R8301 gnd.n6940 gnd.n6939 585
R8302 gnd.n6941 gnd.n6940 585
R8303 gnd.n6938 gnd.n850 585
R8304 gnd.n850 gnd.n849 585
R8305 gnd.n6937 gnd.n6936 585
R8306 gnd.n6936 gnd.n6935 585
R8307 gnd.n856 gnd.n855 585
R8308 gnd.n6934 gnd.n856 585
R8309 gnd.n6932 gnd.n6931 585
R8310 gnd.n6933 gnd.n6932 585
R8311 gnd.n6930 gnd.n858 585
R8312 gnd.n858 gnd.n857 585
R8313 gnd.n6929 gnd.n6928 585
R8314 gnd.n6928 gnd.n6927 585
R8315 gnd.n864 gnd.n863 585
R8316 gnd.n6926 gnd.n864 585
R8317 gnd.n6924 gnd.n6923 585
R8318 gnd.n6925 gnd.n6924 585
R8319 gnd.n6922 gnd.n866 585
R8320 gnd.n866 gnd.n865 585
R8321 gnd.n6921 gnd.n6920 585
R8322 gnd.n6920 gnd.n6919 585
R8323 gnd.n872 gnd.n871 585
R8324 gnd.n6918 gnd.n872 585
R8325 gnd.n6916 gnd.n6915 585
R8326 gnd.n6917 gnd.n6916 585
R8327 gnd.n6914 gnd.n874 585
R8328 gnd.n874 gnd.n873 585
R8329 gnd.n6913 gnd.n6912 585
R8330 gnd.n6912 gnd.n6911 585
R8331 gnd.n880 gnd.n879 585
R8332 gnd.n6910 gnd.n880 585
R8333 gnd.n6908 gnd.n6907 585
R8334 gnd.n6909 gnd.n6908 585
R8335 gnd.n6906 gnd.n882 585
R8336 gnd.n882 gnd.n881 585
R8337 gnd.n6905 gnd.n6904 585
R8338 gnd.n6904 gnd.n6903 585
R8339 gnd.n888 gnd.n887 585
R8340 gnd.n6902 gnd.n888 585
R8341 gnd.n6900 gnd.n6899 585
R8342 gnd.n6901 gnd.n6900 585
R8343 gnd.n6898 gnd.n890 585
R8344 gnd.n890 gnd.n889 585
R8345 gnd.n6897 gnd.n6896 585
R8346 gnd.n6896 gnd.n6895 585
R8347 gnd.n896 gnd.n895 585
R8348 gnd.n6894 gnd.n896 585
R8349 gnd.n6892 gnd.n6891 585
R8350 gnd.n6893 gnd.n6892 585
R8351 gnd.n6890 gnd.n898 585
R8352 gnd.n898 gnd.n897 585
R8353 gnd.n6889 gnd.n6888 585
R8354 gnd.n6888 gnd.n6887 585
R8355 gnd.n904 gnd.n903 585
R8356 gnd.n6886 gnd.n904 585
R8357 gnd.n6884 gnd.n6883 585
R8358 gnd.n6885 gnd.n6884 585
R8359 gnd.n6882 gnd.n906 585
R8360 gnd.n906 gnd.n905 585
R8361 gnd.n6881 gnd.n6880 585
R8362 gnd.n6880 gnd.n6879 585
R8363 gnd.n912 gnd.n911 585
R8364 gnd.n6878 gnd.n912 585
R8365 gnd.n6876 gnd.n6875 585
R8366 gnd.n6877 gnd.n6876 585
R8367 gnd.n6874 gnd.n914 585
R8368 gnd.n914 gnd.n913 585
R8369 gnd.n6873 gnd.n6872 585
R8370 gnd.n6872 gnd.n6871 585
R8371 gnd.n920 gnd.n919 585
R8372 gnd.n6870 gnd.n920 585
R8373 gnd.n6868 gnd.n6867 585
R8374 gnd.n6869 gnd.n6868 585
R8375 gnd.n6866 gnd.n922 585
R8376 gnd.n922 gnd.n921 585
R8377 gnd.n6865 gnd.n6864 585
R8378 gnd.n6864 gnd.n6863 585
R8379 gnd.n928 gnd.n927 585
R8380 gnd.n6862 gnd.n928 585
R8381 gnd.n6860 gnd.n6859 585
R8382 gnd.n6861 gnd.n6860 585
R8383 gnd.n6858 gnd.n930 585
R8384 gnd.n930 gnd.n929 585
R8385 gnd.n6857 gnd.n6856 585
R8386 gnd.n6856 gnd.n6855 585
R8387 gnd.n936 gnd.n935 585
R8388 gnd.n6854 gnd.n936 585
R8389 gnd.n6852 gnd.n6851 585
R8390 gnd.n6853 gnd.n6852 585
R8391 gnd.n6850 gnd.n938 585
R8392 gnd.n938 gnd.n937 585
R8393 gnd.n6849 gnd.n6848 585
R8394 gnd.n6848 gnd.n6847 585
R8395 gnd.n944 gnd.n943 585
R8396 gnd.n6846 gnd.n944 585
R8397 gnd.n6844 gnd.n6843 585
R8398 gnd.n6845 gnd.n6844 585
R8399 gnd.n6842 gnd.n946 585
R8400 gnd.n946 gnd.n945 585
R8401 gnd.n6841 gnd.n6840 585
R8402 gnd.n6840 gnd.n6839 585
R8403 gnd.n952 gnd.n951 585
R8404 gnd.n6838 gnd.n952 585
R8405 gnd.n785 gnd.n784 585
R8406 gnd.n7006 gnd.n785 585
R8407 gnd.n7009 gnd.n7008 585
R8408 gnd.n7008 gnd.n7007 585
R8409 gnd.n782 gnd.n781 585
R8410 gnd.n781 gnd.n780 585
R8411 gnd.n7014 gnd.n7013 585
R8412 gnd.n7015 gnd.n7014 585
R8413 gnd.n779 gnd.n778 585
R8414 gnd.n7016 gnd.n779 585
R8415 gnd.n7019 gnd.n7018 585
R8416 gnd.n7018 gnd.n7017 585
R8417 gnd.n776 gnd.n775 585
R8418 gnd.n775 gnd.n774 585
R8419 gnd.n7024 gnd.n7023 585
R8420 gnd.n7025 gnd.n7024 585
R8421 gnd.n773 gnd.n772 585
R8422 gnd.n7026 gnd.n773 585
R8423 gnd.n7029 gnd.n7028 585
R8424 gnd.n7028 gnd.n7027 585
R8425 gnd.n770 gnd.n769 585
R8426 gnd.n769 gnd.n768 585
R8427 gnd.n7034 gnd.n7033 585
R8428 gnd.n7035 gnd.n7034 585
R8429 gnd.n767 gnd.n766 585
R8430 gnd.n7036 gnd.n767 585
R8431 gnd.n7039 gnd.n7038 585
R8432 gnd.n7038 gnd.n7037 585
R8433 gnd.n764 gnd.n763 585
R8434 gnd.n763 gnd.n762 585
R8435 gnd.n7044 gnd.n7043 585
R8436 gnd.n7045 gnd.n7044 585
R8437 gnd.n761 gnd.n760 585
R8438 gnd.n7046 gnd.n761 585
R8439 gnd.n7049 gnd.n7048 585
R8440 gnd.n7048 gnd.n7047 585
R8441 gnd.n758 gnd.n757 585
R8442 gnd.n757 gnd.n756 585
R8443 gnd.n7054 gnd.n7053 585
R8444 gnd.n7055 gnd.n7054 585
R8445 gnd.n755 gnd.n754 585
R8446 gnd.n7056 gnd.n755 585
R8447 gnd.n7059 gnd.n7058 585
R8448 gnd.n7058 gnd.n7057 585
R8449 gnd.n752 gnd.n751 585
R8450 gnd.n751 gnd.n750 585
R8451 gnd.n7064 gnd.n7063 585
R8452 gnd.n7065 gnd.n7064 585
R8453 gnd.n749 gnd.n748 585
R8454 gnd.n7066 gnd.n749 585
R8455 gnd.n7069 gnd.n7068 585
R8456 gnd.n7068 gnd.n7067 585
R8457 gnd.n746 gnd.n745 585
R8458 gnd.n745 gnd.n744 585
R8459 gnd.n7074 gnd.n7073 585
R8460 gnd.n7075 gnd.n7074 585
R8461 gnd.n743 gnd.n742 585
R8462 gnd.n7076 gnd.n743 585
R8463 gnd.n7079 gnd.n7078 585
R8464 gnd.n7078 gnd.n7077 585
R8465 gnd.n740 gnd.n739 585
R8466 gnd.n739 gnd.n738 585
R8467 gnd.n7084 gnd.n7083 585
R8468 gnd.n7085 gnd.n7084 585
R8469 gnd.n737 gnd.n736 585
R8470 gnd.n7086 gnd.n737 585
R8471 gnd.n7089 gnd.n7088 585
R8472 gnd.n7088 gnd.n7087 585
R8473 gnd.n734 gnd.n733 585
R8474 gnd.n733 gnd.n732 585
R8475 gnd.n7094 gnd.n7093 585
R8476 gnd.n7095 gnd.n7094 585
R8477 gnd.n731 gnd.n730 585
R8478 gnd.n7096 gnd.n731 585
R8479 gnd.n7099 gnd.n7098 585
R8480 gnd.n7098 gnd.n7097 585
R8481 gnd.n728 gnd.n727 585
R8482 gnd.n727 gnd.n726 585
R8483 gnd.n7104 gnd.n7103 585
R8484 gnd.n7105 gnd.n7104 585
R8485 gnd.n725 gnd.n724 585
R8486 gnd.n7106 gnd.n725 585
R8487 gnd.n7109 gnd.n7108 585
R8488 gnd.n7108 gnd.n7107 585
R8489 gnd.n722 gnd.n721 585
R8490 gnd.n721 gnd.n720 585
R8491 gnd.n7114 gnd.n7113 585
R8492 gnd.n7115 gnd.n7114 585
R8493 gnd.n719 gnd.n718 585
R8494 gnd.n7116 gnd.n719 585
R8495 gnd.n7119 gnd.n7118 585
R8496 gnd.n7118 gnd.n7117 585
R8497 gnd.n716 gnd.n715 585
R8498 gnd.n715 gnd.n714 585
R8499 gnd.n7124 gnd.n7123 585
R8500 gnd.n7125 gnd.n7124 585
R8501 gnd.n713 gnd.n712 585
R8502 gnd.n7126 gnd.n713 585
R8503 gnd.n7129 gnd.n7128 585
R8504 gnd.n7128 gnd.n7127 585
R8505 gnd.n710 gnd.n709 585
R8506 gnd.n709 gnd.n708 585
R8507 gnd.n7134 gnd.n7133 585
R8508 gnd.n7135 gnd.n7134 585
R8509 gnd.n707 gnd.n706 585
R8510 gnd.n7136 gnd.n707 585
R8511 gnd.n7139 gnd.n7138 585
R8512 gnd.n7138 gnd.n7137 585
R8513 gnd.n704 gnd.n703 585
R8514 gnd.n703 gnd.n702 585
R8515 gnd.n7144 gnd.n7143 585
R8516 gnd.n7145 gnd.n7144 585
R8517 gnd.n701 gnd.n700 585
R8518 gnd.n7146 gnd.n701 585
R8519 gnd.n7149 gnd.n7148 585
R8520 gnd.n7148 gnd.n7147 585
R8521 gnd.n698 gnd.n697 585
R8522 gnd.n697 gnd.n696 585
R8523 gnd.n7154 gnd.n7153 585
R8524 gnd.n7155 gnd.n7154 585
R8525 gnd.n695 gnd.n694 585
R8526 gnd.n7156 gnd.n695 585
R8527 gnd.n7159 gnd.n7158 585
R8528 gnd.n7158 gnd.n7157 585
R8529 gnd.n692 gnd.n691 585
R8530 gnd.n691 gnd.n690 585
R8531 gnd.n7164 gnd.n7163 585
R8532 gnd.n7165 gnd.n7164 585
R8533 gnd.n689 gnd.n688 585
R8534 gnd.n7166 gnd.n689 585
R8535 gnd.n7169 gnd.n7168 585
R8536 gnd.n7168 gnd.n7167 585
R8537 gnd.n686 gnd.n685 585
R8538 gnd.n685 gnd.n684 585
R8539 gnd.n7174 gnd.n7173 585
R8540 gnd.n7175 gnd.n7174 585
R8541 gnd.n683 gnd.n682 585
R8542 gnd.n7176 gnd.n683 585
R8543 gnd.n7179 gnd.n7178 585
R8544 gnd.n7178 gnd.n7177 585
R8545 gnd.n680 gnd.n679 585
R8546 gnd.n679 gnd.n678 585
R8547 gnd.n7184 gnd.n7183 585
R8548 gnd.n7185 gnd.n7184 585
R8549 gnd.n677 gnd.n676 585
R8550 gnd.n7186 gnd.n677 585
R8551 gnd.n7189 gnd.n7188 585
R8552 gnd.n7188 gnd.n7187 585
R8553 gnd.n674 gnd.n673 585
R8554 gnd.n673 gnd.n672 585
R8555 gnd.n7194 gnd.n7193 585
R8556 gnd.n7195 gnd.n7194 585
R8557 gnd.n671 gnd.n670 585
R8558 gnd.n7196 gnd.n671 585
R8559 gnd.n7199 gnd.n7198 585
R8560 gnd.n7198 gnd.n7197 585
R8561 gnd.n668 gnd.n667 585
R8562 gnd.n667 gnd.n666 585
R8563 gnd.n7204 gnd.n7203 585
R8564 gnd.n7205 gnd.n7204 585
R8565 gnd.n665 gnd.n664 585
R8566 gnd.n7206 gnd.n665 585
R8567 gnd.n7209 gnd.n7208 585
R8568 gnd.n7208 gnd.n7207 585
R8569 gnd.n662 gnd.n661 585
R8570 gnd.n661 gnd.n660 585
R8571 gnd.n7214 gnd.n7213 585
R8572 gnd.n7215 gnd.n7214 585
R8573 gnd.n659 gnd.n658 585
R8574 gnd.n7216 gnd.n659 585
R8575 gnd.n7219 gnd.n7218 585
R8576 gnd.n7218 gnd.n7217 585
R8577 gnd.n656 gnd.n655 585
R8578 gnd.n655 gnd.n654 585
R8579 gnd.n7224 gnd.n7223 585
R8580 gnd.n7225 gnd.n7224 585
R8581 gnd.n653 gnd.n652 585
R8582 gnd.n7226 gnd.n653 585
R8583 gnd.n7229 gnd.n7228 585
R8584 gnd.n7228 gnd.n7227 585
R8585 gnd.n650 gnd.n649 585
R8586 gnd.n649 gnd.n648 585
R8587 gnd.n7234 gnd.n7233 585
R8588 gnd.n7235 gnd.n7234 585
R8589 gnd.n647 gnd.n646 585
R8590 gnd.n7236 gnd.n647 585
R8591 gnd.n7239 gnd.n7238 585
R8592 gnd.n7238 gnd.n7237 585
R8593 gnd.n644 gnd.n643 585
R8594 gnd.n643 gnd.n642 585
R8595 gnd.n7244 gnd.n7243 585
R8596 gnd.n7245 gnd.n7244 585
R8597 gnd.n641 gnd.n640 585
R8598 gnd.n7246 gnd.n641 585
R8599 gnd.n7249 gnd.n7248 585
R8600 gnd.n7248 gnd.n7247 585
R8601 gnd.n638 gnd.n637 585
R8602 gnd.n637 gnd.n636 585
R8603 gnd.n7254 gnd.n7253 585
R8604 gnd.n7255 gnd.n7254 585
R8605 gnd.n635 gnd.n634 585
R8606 gnd.n7256 gnd.n635 585
R8607 gnd.n7259 gnd.n7258 585
R8608 gnd.n7258 gnd.n7257 585
R8609 gnd.n632 gnd.n631 585
R8610 gnd.n631 gnd.n630 585
R8611 gnd.n7264 gnd.n7263 585
R8612 gnd.n7265 gnd.n7264 585
R8613 gnd.n629 gnd.n628 585
R8614 gnd.n7266 gnd.n629 585
R8615 gnd.n7269 gnd.n7268 585
R8616 gnd.n7268 gnd.n7267 585
R8617 gnd.n626 gnd.n625 585
R8618 gnd.n625 gnd.n624 585
R8619 gnd.n7274 gnd.n7273 585
R8620 gnd.n7275 gnd.n7274 585
R8621 gnd.n623 gnd.n622 585
R8622 gnd.n7276 gnd.n623 585
R8623 gnd.n7279 gnd.n7278 585
R8624 gnd.n7278 gnd.n7277 585
R8625 gnd.n620 gnd.n619 585
R8626 gnd.n619 gnd.n618 585
R8627 gnd.n7284 gnd.n7283 585
R8628 gnd.n7285 gnd.n7284 585
R8629 gnd.n617 gnd.n616 585
R8630 gnd.n7286 gnd.n617 585
R8631 gnd.n7289 gnd.n7288 585
R8632 gnd.n7288 gnd.n7287 585
R8633 gnd.n614 gnd.n613 585
R8634 gnd.n613 gnd.n612 585
R8635 gnd.n7294 gnd.n7293 585
R8636 gnd.n7295 gnd.n7294 585
R8637 gnd.n611 gnd.n610 585
R8638 gnd.n7296 gnd.n611 585
R8639 gnd.n7299 gnd.n7298 585
R8640 gnd.n7298 gnd.n7297 585
R8641 gnd.n608 gnd.n607 585
R8642 gnd.n607 gnd.n606 585
R8643 gnd.n7304 gnd.n7303 585
R8644 gnd.n7305 gnd.n7304 585
R8645 gnd.n605 gnd.n604 585
R8646 gnd.n7306 gnd.n605 585
R8647 gnd.n7309 gnd.n7308 585
R8648 gnd.n7308 gnd.n7307 585
R8649 gnd.n602 gnd.n601 585
R8650 gnd.n601 gnd.n600 585
R8651 gnd.n7314 gnd.n7313 585
R8652 gnd.n7315 gnd.n7314 585
R8653 gnd.n599 gnd.n598 585
R8654 gnd.n7316 gnd.n599 585
R8655 gnd.n7319 gnd.n7318 585
R8656 gnd.n7318 gnd.n7317 585
R8657 gnd.n596 gnd.n595 585
R8658 gnd.n595 gnd.n594 585
R8659 gnd.n7324 gnd.n7323 585
R8660 gnd.n7325 gnd.n7324 585
R8661 gnd.n593 gnd.n592 585
R8662 gnd.n7326 gnd.n593 585
R8663 gnd.n7329 gnd.n7328 585
R8664 gnd.n7328 gnd.n7327 585
R8665 gnd.n590 gnd.n589 585
R8666 gnd.n589 gnd.n588 585
R8667 gnd.n7334 gnd.n7333 585
R8668 gnd.n7335 gnd.n7334 585
R8669 gnd.n587 gnd.n586 585
R8670 gnd.n7336 gnd.n587 585
R8671 gnd.n7339 gnd.n7338 585
R8672 gnd.n7338 gnd.n7337 585
R8673 gnd.n584 gnd.n583 585
R8674 gnd.n583 gnd.n582 585
R8675 gnd.n7344 gnd.n7343 585
R8676 gnd.n7345 gnd.n7344 585
R8677 gnd.n581 gnd.n580 585
R8678 gnd.n7346 gnd.n581 585
R8679 gnd.n7349 gnd.n7348 585
R8680 gnd.n7348 gnd.n7347 585
R8681 gnd.n578 gnd.n577 585
R8682 gnd.n577 gnd.n576 585
R8683 gnd.n7354 gnd.n7353 585
R8684 gnd.n7355 gnd.n7354 585
R8685 gnd.n575 gnd.n574 585
R8686 gnd.n7356 gnd.n575 585
R8687 gnd.n7359 gnd.n7358 585
R8688 gnd.n7358 gnd.n7357 585
R8689 gnd.n572 gnd.n571 585
R8690 gnd.n571 gnd.n570 585
R8691 gnd.n7364 gnd.n7363 585
R8692 gnd.n7365 gnd.n7364 585
R8693 gnd.n569 gnd.n568 585
R8694 gnd.n7366 gnd.n569 585
R8695 gnd.n7369 gnd.n7368 585
R8696 gnd.n7368 gnd.n7367 585
R8697 gnd.n566 gnd.n565 585
R8698 gnd.n565 gnd.n564 585
R8699 gnd.n7374 gnd.n7373 585
R8700 gnd.n7375 gnd.n7374 585
R8701 gnd.n563 gnd.n562 585
R8702 gnd.n7376 gnd.n563 585
R8703 gnd.n7379 gnd.n7378 585
R8704 gnd.n7378 gnd.n7377 585
R8705 gnd.n560 gnd.n559 585
R8706 gnd.n559 gnd.n558 585
R8707 gnd.n7384 gnd.n7383 585
R8708 gnd.n7385 gnd.n7384 585
R8709 gnd.n557 gnd.n556 585
R8710 gnd.n7386 gnd.n557 585
R8711 gnd.n7389 gnd.n7388 585
R8712 gnd.n7388 gnd.n7387 585
R8713 gnd.n554 gnd.n553 585
R8714 gnd.n553 gnd.n552 585
R8715 gnd.n7394 gnd.n7393 585
R8716 gnd.n7395 gnd.n7394 585
R8717 gnd.n551 gnd.n550 585
R8718 gnd.n7396 gnd.n551 585
R8719 gnd.n7399 gnd.n7398 585
R8720 gnd.n7398 gnd.n7397 585
R8721 gnd.n548 gnd.n547 585
R8722 gnd.n547 gnd.n546 585
R8723 gnd.n7404 gnd.n7403 585
R8724 gnd.n7405 gnd.n7404 585
R8725 gnd.n545 gnd.n544 585
R8726 gnd.n7406 gnd.n545 585
R8727 gnd.n7409 gnd.n7408 585
R8728 gnd.n7408 gnd.n7407 585
R8729 gnd.n542 gnd.n541 585
R8730 gnd.n541 gnd.n540 585
R8731 gnd.n7414 gnd.n7413 585
R8732 gnd.n7415 gnd.n7414 585
R8733 gnd.n539 gnd.n538 585
R8734 gnd.n7416 gnd.n539 585
R8735 gnd.n7419 gnd.n7418 585
R8736 gnd.n7418 gnd.n7417 585
R8737 gnd.n536 gnd.n535 585
R8738 gnd.n535 gnd.n534 585
R8739 gnd.n7424 gnd.n7423 585
R8740 gnd.n7425 gnd.n7424 585
R8741 gnd.n533 gnd.n532 585
R8742 gnd.n7426 gnd.n533 585
R8743 gnd.n7429 gnd.n7428 585
R8744 gnd.n7428 gnd.n7427 585
R8745 gnd.n530 gnd.n529 585
R8746 gnd.n529 gnd.n528 585
R8747 gnd.n7434 gnd.n7433 585
R8748 gnd.n7435 gnd.n7434 585
R8749 gnd.n527 gnd.n526 585
R8750 gnd.n7436 gnd.n527 585
R8751 gnd.n7439 gnd.n7438 585
R8752 gnd.n7438 gnd.n7437 585
R8753 gnd.n524 gnd.n523 585
R8754 gnd.n523 gnd.n522 585
R8755 gnd.n7444 gnd.n7443 585
R8756 gnd.n7445 gnd.n7444 585
R8757 gnd.n521 gnd.n520 585
R8758 gnd.n7446 gnd.n521 585
R8759 gnd.n7449 gnd.n7448 585
R8760 gnd.n7448 gnd.n7447 585
R8761 gnd.n518 gnd.n517 585
R8762 gnd.n517 gnd.n516 585
R8763 gnd.n7454 gnd.n7453 585
R8764 gnd.n7455 gnd.n7454 585
R8765 gnd.n515 gnd.n514 585
R8766 gnd.n7456 gnd.n515 585
R8767 gnd.n7459 gnd.n7458 585
R8768 gnd.n7458 gnd.n7457 585
R8769 gnd.n512 gnd.n511 585
R8770 gnd.n511 gnd.n510 585
R8771 gnd.n7464 gnd.n7463 585
R8772 gnd.n7465 gnd.n7464 585
R8773 gnd.n509 gnd.n508 585
R8774 gnd.n7466 gnd.n509 585
R8775 gnd.n7469 gnd.n7468 585
R8776 gnd.n7468 gnd.n7467 585
R8777 gnd.n506 gnd.n505 585
R8778 gnd.n505 gnd.n504 585
R8779 gnd.n7474 gnd.n7473 585
R8780 gnd.n7475 gnd.n7474 585
R8781 gnd.n503 gnd.n502 585
R8782 gnd.n7476 gnd.n503 585
R8783 gnd.n7479 gnd.n7478 585
R8784 gnd.n7478 gnd.n7477 585
R8785 gnd.n500 gnd.n499 585
R8786 gnd.n499 gnd.n498 585
R8787 gnd.n7485 gnd.n7484 585
R8788 gnd.n7486 gnd.n7485 585
R8789 gnd.n497 gnd.n496 585
R8790 gnd.n7487 gnd.n497 585
R8791 gnd.n7490 gnd.n7489 585
R8792 gnd.n7489 gnd.n7488 585
R8793 gnd.n7491 gnd.n494 585
R8794 gnd.n494 gnd.n493 585
R8795 gnd.n369 gnd.n368 585
R8796 gnd.n7698 gnd.n368 585
R8797 gnd.n7701 gnd.n7700 585
R8798 gnd.n7700 gnd.n7699 585
R8799 gnd.n372 gnd.n371 585
R8800 gnd.n7697 gnd.n372 585
R8801 gnd.n7695 gnd.n7694 585
R8802 gnd.n7696 gnd.n7695 585
R8803 gnd.n375 gnd.n374 585
R8804 gnd.n374 gnd.n373 585
R8805 gnd.n7690 gnd.n7689 585
R8806 gnd.n7689 gnd.n7688 585
R8807 gnd.n378 gnd.n377 585
R8808 gnd.n7687 gnd.n378 585
R8809 gnd.n7685 gnd.n7684 585
R8810 gnd.n7686 gnd.n7685 585
R8811 gnd.n381 gnd.n380 585
R8812 gnd.n380 gnd.n379 585
R8813 gnd.n7680 gnd.n7679 585
R8814 gnd.n7679 gnd.n7678 585
R8815 gnd.n384 gnd.n383 585
R8816 gnd.n7677 gnd.n384 585
R8817 gnd.n7675 gnd.n7674 585
R8818 gnd.n7676 gnd.n7675 585
R8819 gnd.n387 gnd.n386 585
R8820 gnd.n386 gnd.n385 585
R8821 gnd.n7670 gnd.n7669 585
R8822 gnd.n7669 gnd.n7668 585
R8823 gnd.n390 gnd.n389 585
R8824 gnd.n7667 gnd.n390 585
R8825 gnd.n7665 gnd.n7664 585
R8826 gnd.n7666 gnd.n7665 585
R8827 gnd.n393 gnd.n392 585
R8828 gnd.n392 gnd.n391 585
R8829 gnd.n7660 gnd.n7659 585
R8830 gnd.n7659 gnd.n7658 585
R8831 gnd.n396 gnd.n395 585
R8832 gnd.n7657 gnd.n396 585
R8833 gnd.n7655 gnd.n7654 585
R8834 gnd.n7656 gnd.n7655 585
R8835 gnd.n399 gnd.n398 585
R8836 gnd.n398 gnd.n397 585
R8837 gnd.n7650 gnd.n7649 585
R8838 gnd.n7649 gnd.n7648 585
R8839 gnd.n402 gnd.n401 585
R8840 gnd.n7647 gnd.n402 585
R8841 gnd.n7645 gnd.n7644 585
R8842 gnd.n7646 gnd.n7645 585
R8843 gnd.n405 gnd.n404 585
R8844 gnd.n404 gnd.n403 585
R8845 gnd.n7640 gnd.n7639 585
R8846 gnd.n7639 gnd.n7638 585
R8847 gnd.n408 gnd.n407 585
R8848 gnd.n7637 gnd.n408 585
R8849 gnd.n7635 gnd.n7634 585
R8850 gnd.n7636 gnd.n7635 585
R8851 gnd.n411 gnd.n410 585
R8852 gnd.n410 gnd.n409 585
R8853 gnd.n7630 gnd.n7629 585
R8854 gnd.n7629 gnd.n7628 585
R8855 gnd.n414 gnd.n413 585
R8856 gnd.n7627 gnd.n414 585
R8857 gnd.n7625 gnd.n7624 585
R8858 gnd.n7626 gnd.n7625 585
R8859 gnd.n417 gnd.n416 585
R8860 gnd.n416 gnd.n415 585
R8861 gnd.n7620 gnd.n7619 585
R8862 gnd.n7619 gnd.n7618 585
R8863 gnd.n420 gnd.n419 585
R8864 gnd.n7617 gnd.n420 585
R8865 gnd.n7615 gnd.n7614 585
R8866 gnd.n7616 gnd.n7615 585
R8867 gnd.n423 gnd.n422 585
R8868 gnd.n422 gnd.n421 585
R8869 gnd.n7610 gnd.n7609 585
R8870 gnd.n7609 gnd.n7608 585
R8871 gnd.n426 gnd.n425 585
R8872 gnd.n7607 gnd.n426 585
R8873 gnd.n7605 gnd.n7604 585
R8874 gnd.n7606 gnd.n7605 585
R8875 gnd.n429 gnd.n428 585
R8876 gnd.n428 gnd.n427 585
R8877 gnd.n7600 gnd.n7599 585
R8878 gnd.n7599 gnd.n7598 585
R8879 gnd.n432 gnd.n431 585
R8880 gnd.n7597 gnd.n432 585
R8881 gnd.n7595 gnd.n7594 585
R8882 gnd.n7596 gnd.n7595 585
R8883 gnd.n435 gnd.n434 585
R8884 gnd.n434 gnd.n433 585
R8885 gnd.n7590 gnd.n7589 585
R8886 gnd.n7589 gnd.n7588 585
R8887 gnd.n438 gnd.n437 585
R8888 gnd.n7587 gnd.n438 585
R8889 gnd.n7585 gnd.n7584 585
R8890 gnd.n7586 gnd.n7585 585
R8891 gnd.n441 gnd.n440 585
R8892 gnd.n440 gnd.n439 585
R8893 gnd.n7580 gnd.n7579 585
R8894 gnd.n7579 gnd.n7578 585
R8895 gnd.n444 gnd.n443 585
R8896 gnd.n7577 gnd.n444 585
R8897 gnd.n7575 gnd.n7574 585
R8898 gnd.n7576 gnd.n7575 585
R8899 gnd.n447 gnd.n446 585
R8900 gnd.n446 gnd.n445 585
R8901 gnd.n7570 gnd.n7569 585
R8902 gnd.n7569 gnd.n7568 585
R8903 gnd.n450 gnd.n449 585
R8904 gnd.n7567 gnd.n450 585
R8905 gnd.n7565 gnd.n7564 585
R8906 gnd.n7566 gnd.n7565 585
R8907 gnd.n453 gnd.n452 585
R8908 gnd.n452 gnd.n451 585
R8909 gnd.n7560 gnd.n7559 585
R8910 gnd.n7559 gnd.n7558 585
R8911 gnd.n456 gnd.n455 585
R8912 gnd.n7557 gnd.n456 585
R8913 gnd.n7555 gnd.n7554 585
R8914 gnd.n7556 gnd.n7555 585
R8915 gnd.n459 gnd.n458 585
R8916 gnd.n458 gnd.n457 585
R8917 gnd.n7550 gnd.n7549 585
R8918 gnd.n7549 gnd.n7548 585
R8919 gnd.n462 gnd.n461 585
R8920 gnd.n7547 gnd.n462 585
R8921 gnd.n7545 gnd.n7544 585
R8922 gnd.n7546 gnd.n7545 585
R8923 gnd.n465 gnd.n464 585
R8924 gnd.n464 gnd.n463 585
R8925 gnd.n7540 gnd.n7539 585
R8926 gnd.n7539 gnd.n7538 585
R8927 gnd.n468 gnd.n467 585
R8928 gnd.n7537 gnd.n468 585
R8929 gnd.n7535 gnd.n7534 585
R8930 gnd.n7536 gnd.n7535 585
R8931 gnd.n471 gnd.n470 585
R8932 gnd.n470 gnd.n469 585
R8933 gnd.n7530 gnd.n7529 585
R8934 gnd.n7529 gnd.n7528 585
R8935 gnd.n474 gnd.n473 585
R8936 gnd.n7527 gnd.n474 585
R8937 gnd.n7525 gnd.n7524 585
R8938 gnd.n7526 gnd.n7525 585
R8939 gnd.n477 gnd.n476 585
R8940 gnd.n476 gnd.n475 585
R8941 gnd.n7520 gnd.n7519 585
R8942 gnd.n7519 gnd.n7518 585
R8943 gnd.n480 gnd.n479 585
R8944 gnd.n7517 gnd.n480 585
R8945 gnd.n7515 gnd.n7514 585
R8946 gnd.n7516 gnd.n7515 585
R8947 gnd.n483 gnd.n482 585
R8948 gnd.n482 gnd.n481 585
R8949 gnd.n7510 gnd.n7509 585
R8950 gnd.n7509 gnd.n7508 585
R8951 gnd.n486 gnd.n485 585
R8952 gnd.n7507 gnd.n486 585
R8953 gnd.n7505 gnd.n7504 585
R8954 gnd.n7506 gnd.n7505 585
R8955 gnd.n489 gnd.n488 585
R8956 gnd.n488 gnd.n487 585
R8957 gnd.n7500 gnd.n7499 585
R8958 gnd.n7499 gnd.n7498 585
R8959 gnd.n492 gnd.n491 585
R8960 gnd.n7497 gnd.n492 585
R8961 gnd.n7495 gnd.n7494 585
R8962 gnd.n7496 gnd.n7495 585
R8963 gnd.n2754 gnd.n2753 585
R8964 gnd.n4764 gnd.n2754 585
R8965 gnd.n6454 gnd.n6453 585
R8966 gnd.n6453 gnd.n6452 585
R8967 gnd.n6455 gnd.n2749 585
R8968 gnd.n4724 gnd.n2749 585
R8969 gnd.n6457 gnd.n6456 585
R8970 gnd.n6458 gnd.n6457 585
R8971 gnd.n2733 gnd.n2732 585
R8972 gnd.n4472 gnd.n2733 585
R8973 gnd.n6466 gnd.n6465 585
R8974 gnd.n6465 gnd.n6464 585
R8975 gnd.n6467 gnd.n2728 585
R8976 gnd.n4737 gnd.n2728 585
R8977 gnd.n6469 gnd.n6468 585
R8978 gnd.n6470 gnd.n6469 585
R8979 gnd.n2714 gnd.n2713 585
R8980 gnd.n4465 gnd.n2714 585
R8981 gnd.n6478 gnd.n6477 585
R8982 gnd.n6477 gnd.n6476 585
R8983 gnd.n6479 gnd.n2709 585
R8984 gnd.n4457 gnd.n2709 585
R8985 gnd.n6481 gnd.n6480 585
R8986 gnd.n6482 gnd.n6481 585
R8987 gnd.n2693 gnd.n2692 585
R8988 gnd.n4419 gnd.n2693 585
R8989 gnd.n6490 gnd.n6489 585
R8990 gnd.n6489 gnd.n6488 585
R8991 gnd.n6491 gnd.n2688 585
R8992 gnd.n4410 gnd.n2688 585
R8993 gnd.n6493 gnd.n6492 585
R8994 gnd.n6494 gnd.n6493 585
R8995 gnd.n2674 gnd.n2673 585
R8996 gnd.n4405 gnd.n2674 585
R8997 gnd.n6502 gnd.n6501 585
R8998 gnd.n6501 gnd.n6500 585
R8999 gnd.n6503 gnd.n2669 585
R9000 gnd.n4433 gnd.n2669 585
R9001 gnd.n6505 gnd.n6504 585
R9002 gnd.n6506 gnd.n6505 585
R9003 gnd.n2653 gnd.n2652 585
R9004 gnd.n4398 gnd.n2653 585
R9005 gnd.n6514 gnd.n6513 585
R9006 gnd.n6513 gnd.n6512 585
R9007 gnd.n6515 gnd.n2648 585
R9008 gnd.n4390 gnd.n2648 585
R9009 gnd.n6517 gnd.n6516 585
R9010 gnd.n6518 gnd.n6517 585
R9011 gnd.n2635 gnd.n2634 585
R9012 gnd.n4384 gnd.n2635 585
R9013 gnd.n6526 gnd.n6525 585
R9014 gnd.n6525 gnd.n6524 585
R9015 gnd.n6527 gnd.n2629 585
R9016 gnd.n4376 gnd.n2629 585
R9017 gnd.n6529 gnd.n6528 585
R9018 gnd.n6530 gnd.n6529 585
R9019 gnd.n2630 gnd.n2628 585
R9020 gnd.n4345 gnd.n2628 585
R9021 gnd.n4327 gnd.n4326 585
R9022 gnd.n4326 gnd.n4016 585
R9023 gnd.n4328 gnd.n4026 585
R9024 gnd.n4337 gnd.n4026 585
R9025 gnd.n4330 gnd.n4329 585
R9026 gnd.n4331 gnd.n4330 585
R9027 gnd.n4033 gnd.n4032 585
R9028 gnd.n4315 gnd.n4032 585
R9029 gnd.n4268 gnd.n4267 585
R9030 gnd.n4267 gnd.n4266 585
R9031 gnd.n2607 gnd.n2606 585
R9032 gnd.n4307 gnd.n2607 585
R9033 gnd.n6539 gnd.n6538 585
R9034 gnd.n6538 gnd.n6537 585
R9035 gnd.n6540 gnd.n2602 585
R9036 gnd.n4275 gnd.n2602 585
R9037 gnd.n6542 gnd.n6541 585
R9038 gnd.n6543 gnd.n6542 585
R9039 gnd.n2588 gnd.n2587 585
R9040 gnd.n4281 gnd.n2588 585
R9041 gnd.n6551 gnd.n6550 585
R9042 gnd.n6550 gnd.n6549 585
R9043 gnd.n6552 gnd.n2583 585
R9044 gnd.n4257 gnd.n2583 585
R9045 gnd.n6554 gnd.n6553 585
R9046 gnd.n6555 gnd.n6554 585
R9047 gnd.n2568 gnd.n2567 585
R9048 gnd.n4248 gnd.n2568 585
R9049 gnd.n6563 gnd.n6562 585
R9050 gnd.n6562 gnd.n6561 585
R9051 gnd.n6564 gnd.n2563 585
R9052 gnd.n4211 gnd.n2563 585
R9053 gnd.n6566 gnd.n6565 585
R9054 gnd.n6567 gnd.n6566 585
R9055 gnd.n2548 gnd.n2547 585
R9056 gnd.n4217 gnd.n2548 585
R9057 gnd.n6575 gnd.n6574 585
R9058 gnd.n6574 gnd.n6573 585
R9059 gnd.n6576 gnd.n2543 585
R9060 gnd.n4199 gnd.n2543 585
R9061 gnd.n6578 gnd.n6577 585
R9062 gnd.n6579 gnd.n6578 585
R9063 gnd.n2528 gnd.n2527 585
R9064 gnd.n2532 gnd.n2528 585
R9065 gnd.n6587 gnd.n6586 585
R9066 gnd.n6586 gnd.n6585 585
R9067 gnd.n6588 gnd.n2523 585
R9068 gnd.n2523 gnd.n2522 585
R9069 gnd.n6590 gnd.n6589 585
R9070 gnd.n6591 gnd.n6590 585
R9071 gnd.n2509 gnd.n2508 585
R9072 gnd.n2519 gnd.n2509 585
R9073 gnd.n6599 gnd.n6598 585
R9074 gnd.n6598 gnd.n6597 585
R9075 gnd.n6600 gnd.n2504 585
R9076 gnd.n2504 gnd.n2503 585
R9077 gnd.n6602 gnd.n6601 585
R9078 gnd.n6603 gnd.n6602 585
R9079 gnd.n2490 gnd.n2489 585
R9080 gnd.n2493 gnd.n2490 585
R9081 gnd.n6611 gnd.n6610 585
R9082 gnd.n6610 gnd.n6609 585
R9083 gnd.n6612 gnd.n2483 585
R9084 gnd.n2483 gnd.n2481 585
R9085 gnd.n6614 gnd.n6613 585
R9086 gnd.n6615 gnd.n6614 585
R9087 gnd.n2485 gnd.n2482 585
R9088 gnd.n2482 gnd.n2478 585
R9089 gnd.n2484 gnd.n2469 585
R9090 gnd.n6621 gnd.n2469 585
R9091 gnd.n4119 gnd.n2463 585
R9092 gnd.n4119 gnd.n2394 585
R9093 gnd.n4121 gnd.n4120 585
R9094 gnd.n4123 gnd.n4122 585
R9095 gnd.n4125 gnd.n4124 585
R9096 gnd.n4129 gnd.n4117 585
R9097 gnd.n4131 gnd.n4130 585
R9098 gnd.n4133 gnd.n4132 585
R9099 gnd.n4135 gnd.n4134 585
R9100 gnd.n4139 gnd.n4115 585
R9101 gnd.n4141 gnd.n4140 585
R9102 gnd.n4143 gnd.n4142 585
R9103 gnd.n4145 gnd.n4144 585
R9104 gnd.n4149 gnd.n4113 585
R9105 gnd.n4151 gnd.n4150 585
R9106 gnd.n4153 gnd.n4152 585
R9107 gnd.n4155 gnd.n4154 585
R9108 gnd.n4110 gnd.n4109 585
R9109 gnd.n4159 gnd.n4111 585
R9110 gnd.n4160 gnd.n4106 585
R9111 gnd.n4161 gnd.n2393 585
R9112 gnd.n6745 gnd.n2393 585
R9113 gnd.n4767 gnd.n4766 585
R9114 gnd.n4561 gnd.n3955 585
R9115 gnd.n4573 gnd.n4562 585
R9116 gnd.n4574 gnd.n4560 585
R9117 gnd.n4559 gnd.n4551 585
R9118 gnd.n4581 gnd.n4550 585
R9119 gnd.n4582 gnd.n4549 585
R9120 gnd.n4543 gnd.n4542 585
R9121 gnd.n4589 gnd.n4541 585
R9122 gnd.n4590 gnd.n4540 585
R9123 gnd.n4539 gnd.n4531 585
R9124 gnd.n4597 gnd.n4530 585
R9125 gnd.n4598 gnd.n4529 585
R9126 gnd.n4523 gnd.n4522 585
R9127 gnd.n4605 gnd.n4521 585
R9128 gnd.n4606 gnd.n4520 585
R9129 gnd.n4519 gnd.n4511 585
R9130 gnd.n4613 gnd.n4510 585
R9131 gnd.n4614 gnd.n2766 585
R9132 gnd.n6444 gnd.n2766 585
R9133 gnd.n4765 gnd.n3956 585
R9134 gnd.n4765 gnd.n4764 585
R9135 gnd.n4726 gnd.n2757 585
R9136 gnd.n6452 gnd.n2757 585
R9137 gnd.n4729 gnd.n4725 585
R9138 gnd.n4725 gnd.n4724 585
R9139 gnd.n4730 gnd.n2747 585
R9140 gnd.n6458 gnd.n2747 585
R9141 gnd.n4731 gnd.n3973 585
R9142 gnd.n4472 gnd.n3973 585
R9143 gnd.n3970 gnd.n2736 585
R9144 gnd.n6464 gnd.n2736 585
R9145 gnd.n4736 gnd.n4735 585
R9146 gnd.n4737 gnd.n4736 585
R9147 gnd.n3969 gnd.n2727 585
R9148 gnd.n6470 gnd.n2727 585
R9149 gnd.n4464 gnd.n4463 585
R9150 gnd.n4465 gnd.n4464 585
R9151 gnd.n3976 gnd.n2716 585
R9152 gnd.n6476 gnd.n2716 585
R9153 gnd.n4459 gnd.n4458 585
R9154 gnd.n4458 gnd.n4457 585
R9155 gnd.n3978 gnd.n2707 585
R9156 gnd.n6482 gnd.n2707 585
R9157 gnd.n4421 gnd.n4420 585
R9158 gnd.n4420 gnd.n4419 585
R9159 gnd.n3998 gnd.n2696 585
R9160 gnd.n6488 gnd.n2696 585
R9161 gnd.n4425 gnd.n3997 585
R9162 gnd.n4410 gnd.n3997 585
R9163 gnd.n4426 gnd.n2687 585
R9164 gnd.n6494 gnd.n2687 585
R9165 gnd.n4427 gnd.n3996 585
R9166 gnd.n4405 gnd.n3996 585
R9167 gnd.n3993 gnd.n2676 585
R9168 gnd.n6500 gnd.n2676 585
R9169 gnd.n4432 gnd.n4431 585
R9170 gnd.n4433 gnd.n4432 585
R9171 gnd.n3992 gnd.n2667 585
R9172 gnd.n6506 gnd.n2667 585
R9173 gnd.n4397 gnd.n4396 585
R9174 gnd.n4398 gnd.n4397 585
R9175 gnd.n4001 gnd.n2656 585
R9176 gnd.n6512 gnd.n2656 585
R9177 gnd.n4392 gnd.n4391 585
R9178 gnd.n4391 gnd.n4390 585
R9179 gnd.n4003 gnd.n2647 585
R9180 gnd.n6518 gnd.n2647 585
R9181 gnd.n4383 gnd.n4382 585
R9182 gnd.n4384 gnd.n4383 585
R9183 gnd.n4007 gnd.n2637 585
R9184 gnd.n6524 gnd.n2637 585
R9185 gnd.n4378 gnd.n4377 585
R9186 gnd.n4377 gnd.n4376 585
R9187 gnd.n4009 gnd.n2626 585
R9188 gnd.n6530 gnd.n2626 585
R9189 gnd.n4344 gnd.n4343 585
R9190 gnd.n4345 gnd.n4344 585
R9191 gnd.n4019 gnd.n4018 585
R9192 gnd.n4018 gnd.n4016 585
R9193 gnd.n4339 gnd.n4338 585
R9194 gnd.n4338 gnd.n4337 585
R9195 gnd.n4022 gnd.n4021 585
R9196 gnd.n4331 gnd.n4022 585
R9197 gnd.n4314 gnd.n4313 585
R9198 gnd.n4315 gnd.n4314 585
R9199 gnd.n4042 gnd.n4041 585
R9200 gnd.n4266 gnd.n4041 585
R9201 gnd.n4309 gnd.n4308 585
R9202 gnd.n4308 gnd.n4307 585
R9203 gnd.n4044 gnd.n2610 585
R9204 gnd.n6537 gnd.n2610 585
R9205 gnd.n4277 gnd.n4276 585
R9206 gnd.n4276 gnd.n4275 585
R9207 gnd.n4278 gnd.n2600 585
R9208 gnd.n6543 gnd.n2600 585
R9209 gnd.n4280 gnd.n4279 585
R9210 gnd.n4281 gnd.n4280 585
R9211 gnd.n4055 gnd.n2591 585
R9212 gnd.n6549 gnd.n2591 585
R9213 gnd.n4256 gnd.n4255 585
R9214 gnd.n4257 gnd.n4256 585
R9215 gnd.n4060 gnd.n2581 585
R9216 gnd.n6555 gnd.n2581 585
R9217 gnd.n4250 gnd.n4249 585
R9218 gnd.n4249 gnd.n4248 585
R9219 gnd.n4062 gnd.n2571 585
R9220 gnd.n6561 gnd.n2571 585
R9221 gnd.n4213 gnd.n4212 585
R9222 gnd.n4212 gnd.n4211 585
R9223 gnd.n4214 gnd.n2561 585
R9224 gnd.n6567 gnd.n2561 585
R9225 gnd.n4216 gnd.n4215 585
R9226 gnd.n4217 gnd.n4216 585
R9227 gnd.n4069 gnd.n2551 585
R9228 gnd.n6573 gnd.n2551 585
R9229 gnd.n4198 gnd.n4197 585
R9230 gnd.n4199 gnd.n4198 585
R9231 gnd.n4097 gnd.n2541 585
R9232 gnd.n6579 gnd.n2541 585
R9233 gnd.n4192 gnd.n4191 585
R9234 gnd.n4191 gnd.n2532 585
R9235 gnd.n4190 gnd.n2531 585
R9236 gnd.n6585 gnd.n2531 585
R9237 gnd.n4189 gnd.n4188 585
R9238 gnd.n4188 gnd.n2522 585
R9239 gnd.n4099 gnd.n2521 585
R9240 gnd.n6591 gnd.n2521 585
R9241 gnd.n4184 gnd.n4183 585
R9242 gnd.n4183 gnd.n2519 585
R9243 gnd.n4182 gnd.n2511 585
R9244 gnd.n6597 gnd.n2511 585
R9245 gnd.n4181 gnd.n4180 585
R9246 gnd.n4180 gnd.n2503 585
R9247 gnd.n4101 gnd.n2502 585
R9248 gnd.n6603 gnd.n2502 585
R9249 gnd.n4176 gnd.n4175 585
R9250 gnd.n4175 gnd.n2493 585
R9251 gnd.n4174 gnd.n2492 585
R9252 gnd.n6609 gnd.n2492 585
R9253 gnd.n4173 gnd.n4172 585
R9254 gnd.n4172 gnd.n2481 585
R9255 gnd.n4103 gnd.n2480 585
R9256 gnd.n6615 gnd.n2480 585
R9257 gnd.n4168 gnd.n4167 585
R9258 gnd.n4167 gnd.n2478 585
R9259 gnd.n4166 gnd.n2468 585
R9260 gnd.n6621 gnd.n2468 585
R9261 gnd.n4165 gnd.n4164 585
R9262 gnd.n4164 gnd.n2394 585
R9263 gnd.n6807 gnd.n6806 585
R9264 gnd.n6808 gnd.n6807 585
R9265 gnd.n1007 gnd.n1005 585
R9266 gnd.n1005 gnd.n1001 585
R9267 gnd.n987 gnd.n986 585
R9268 gnd.n2346 gnd.n987 585
R9269 gnd.n6818 gnd.n6817 585
R9270 gnd.n6817 gnd.n6816 585
R9271 gnd.n6819 gnd.n981 585
R9272 gnd.n2022 gnd.n981 585
R9273 gnd.n6821 gnd.n6820 585
R9274 gnd.n6822 gnd.n6821 585
R9275 gnd.n982 gnd.n980 585
R9276 gnd.n980 gnd.n976 585
R9277 gnd.n963 gnd.n962 585
R9278 gnd.n967 gnd.n963 585
R9279 gnd.n6832 gnd.n6831 585
R9280 gnd.n6831 gnd.n6830 585
R9281 gnd.n6833 gnd.n957 585
R9282 gnd.n2031 gnd.n957 585
R9283 gnd.n6835 gnd.n6834 585
R9284 gnd.n6836 gnd.n6835 585
R9285 gnd.n958 gnd.n956 585
R9286 gnd.n2035 gnd.n956 585
R9287 gnd.n2059 gnd.n2058 585
R9288 gnd.n2058 gnd.n2057 585
R9289 gnd.n1122 gnd.n1121 585
R9290 gnd.n2041 gnd.n1122 585
R9291 gnd.n2001 gnd.n1141 585
R9292 gnd.n1141 gnd.n1131 585
R9293 gnd.n2003 gnd.n2002 585
R9294 gnd.n2004 gnd.n2003 585
R9295 gnd.n1142 gnd.n1140 585
R9296 gnd.n1149 gnd.n1140 585
R9297 gnd.n1977 gnd.n1161 585
R9298 gnd.n1926 gnd.n1161 585
R9299 gnd.n1979 gnd.n1978 585
R9300 gnd.n1980 gnd.n1979 585
R9301 gnd.n1162 gnd.n1160 585
R9302 gnd.n1160 gnd.n1156 585
R9303 gnd.n1965 gnd.n1964 585
R9304 gnd.n1964 gnd.n1963 585
R9305 gnd.n1167 gnd.n1166 585
R9306 gnd.n1176 gnd.n1167 585
R9307 gnd.n1954 gnd.n1953 585
R9308 gnd.n1953 gnd.n1952 585
R9309 gnd.n1174 gnd.n1173 585
R9310 gnd.n1940 gnd.n1174 585
R9311 gnd.n1911 gnd.n1192 585
R9312 gnd.n1192 gnd.n1183 585
R9313 gnd.n1913 gnd.n1912 585
R9314 gnd.n1914 gnd.n1913 585
R9315 gnd.n1193 gnd.n1191 585
R9316 gnd.n1201 gnd.n1191 585
R9317 gnd.n1888 gnd.n1213 585
R9318 gnd.n1213 gnd.n1200 585
R9319 gnd.n1890 gnd.n1889 585
R9320 gnd.n1891 gnd.n1890 585
R9321 gnd.n1214 gnd.n1212 585
R9322 gnd.n1212 gnd.n1208 585
R9323 gnd.n1876 gnd.n1875 585
R9324 gnd.n1875 gnd.n1874 585
R9325 gnd.n1219 gnd.n1218 585
R9326 gnd.n1223 gnd.n1219 585
R9327 gnd.n1860 gnd.n1859 585
R9328 gnd.n1861 gnd.n1860 585
R9329 gnd.n1233 gnd.n1232 585
R9330 gnd.n1851 gnd.n1232 585
R9331 gnd.n1351 gnd.n1350 585
R9332 gnd.n1351 gnd.n1240 585
R9333 gnd.n1838 gnd.n1837 585
R9334 gnd.n1837 gnd.n1836 585
R9335 gnd.n1839 gnd.n1343 585
R9336 gnd.n1816 gnd.n1343 585
R9337 gnd.n1841 gnd.n1840 585
R9338 gnd.n1842 gnd.n1841 585
R9339 gnd.n1344 gnd.n1342 585
R9340 gnd.n1824 gnd.n1342 585
R9341 gnd.n1808 gnd.n1807 585
R9342 gnd.n1807 gnd.n1361 585
R9343 gnd.n1806 gnd.n1366 585
R9344 gnd.n1806 gnd.n1805 585
R9345 gnd.n1791 gnd.n1367 585
R9346 gnd.n1375 gnd.n1367 585
R9347 gnd.n1793 gnd.n1792 585
R9348 gnd.n1794 gnd.n1793 585
R9349 gnd.n1378 gnd.n1377 585
R9350 gnd.n1385 gnd.n1377 585
R9351 gnd.n1766 gnd.n1765 585
R9352 gnd.n1767 gnd.n1766 585
R9353 gnd.n1397 gnd.n1396 585
R9354 gnd.n1396 gnd.n1392 585
R9355 gnd.n1756 gnd.n1755 585
R9356 gnd.n1757 gnd.n1756 585
R9357 gnd.n1407 gnd.n1406 585
R9358 gnd.n1412 gnd.n1406 585
R9359 gnd.n1734 gnd.n1425 585
R9360 gnd.n1425 gnd.n1411 585
R9361 gnd.n1736 gnd.n1735 585
R9362 gnd.n1737 gnd.n1736 585
R9363 gnd.n1426 gnd.n1424 585
R9364 gnd.n1424 gnd.n1420 585
R9365 gnd.n1725 gnd.n1724 585
R9366 gnd.n1726 gnd.n1725 585
R9367 gnd.n1433 gnd.n1432 585
R9368 gnd.n1437 gnd.n1432 585
R9369 gnd.n1702 gnd.n1454 585
R9370 gnd.n1454 gnd.n1436 585
R9371 gnd.n1704 gnd.n1703 585
R9372 gnd.n1705 gnd.n1704 585
R9373 gnd.n1455 gnd.n1453 585
R9374 gnd.n1453 gnd.n1444 585
R9375 gnd.n1697 gnd.n1696 585
R9376 gnd.n1696 gnd.n1695 585
R9377 gnd.n1502 gnd.n1501 585
R9378 gnd.n1503 gnd.n1502 585
R9379 gnd.n1656 gnd.n1655 585
R9380 gnd.n1657 gnd.n1656 585
R9381 gnd.n1512 gnd.n1511 585
R9382 gnd.n1511 gnd.n1510 585
R9383 gnd.n1651 gnd.n1650 585
R9384 gnd.n1650 gnd.n1649 585
R9385 gnd.n1515 gnd.n1514 585
R9386 gnd.n1516 gnd.n1515 585
R9387 gnd.n1640 gnd.n1639 585
R9388 gnd.n1641 gnd.n1640 585
R9389 gnd.n1523 gnd.n1522 585
R9390 gnd.n1632 gnd.n1522 585
R9391 gnd.n1635 gnd.n1634 585
R9392 gnd.n1634 gnd.n1633 585
R9393 gnd.n1526 gnd.n1525 585
R9394 gnd.n1527 gnd.n1526 585
R9395 gnd.n1621 gnd.n1620 585
R9396 gnd.n1619 gnd.n1545 585
R9397 gnd.n1618 gnd.n1544 585
R9398 gnd.n1623 gnd.n1544 585
R9399 gnd.n1617 gnd.n1616 585
R9400 gnd.n1615 gnd.n1614 585
R9401 gnd.n1613 gnd.n1612 585
R9402 gnd.n1611 gnd.n1610 585
R9403 gnd.n1609 gnd.n1608 585
R9404 gnd.n1607 gnd.n1606 585
R9405 gnd.n1605 gnd.n1604 585
R9406 gnd.n1603 gnd.n1602 585
R9407 gnd.n1601 gnd.n1600 585
R9408 gnd.n1599 gnd.n1598 585
R9409 gnd.n1597 gnd.n1596 585
R9410 gnd.n1595 gnd.n1594 585
R9411 gnd.n1593 gnd.n1592 585
R9412 gnd.n1591 gnd.n1590 585
R9413 gnd.n1589 gnd.n1588 585
R9414 gnd.n1587 gnd.n1586 585
R9415 gnd.n1585 gnd.n1584 585
R9416 gnd.n1583 gnd.n1582 585
R9417 gnd.n1581 gnd.n1580 585
R9418 gnd.n1579 gnd.n1578 585
R9419 gnd.n1577 gnd.n1576 585
R9420 gnd.n1575 gnd.n1574 585
R9421 gnd.n1532 gnd.n1531 585
R9422 gnd.n1626 gnd.n1625 585
R9423 gnd.n2354 gnd.n2353 585
R9424 gnd.n1031 gnd.n1030 585
R9425 gnd.n1107 gnd.n1106 585
R9426 gnd.n1105 gnd.n1104 585
R9427 gnd.n1103 gnd.n1102 585
R9428 gnd.n1096 gnd.n1036 585
R9429 gnd.n1098 gnd.n1097 585
R9430 gnd.n1095 gnd.n1094 585
R9431 gnd.n1093 gnd.n1092 585
R9432 gnd.n1086 gnd.n1038 585
R9433 gnd.n1088 gnd.n1087 585
R9434 gnd.n1085 gnd.n1084 585
R9435 gnd.n1083 gnd.n1082 585
R9436 gnd.n1076 gnd.n1040 585
R9437 gnd.n1078 gnd.n1077 585
R9438 gnd.n1075 gnd.n1074 585
R9439 gnd.n1073 gnd.n1072 585
R9440 gnd.n1066 gnd.n1042 585
R9441 gnd.n1068 gnd.n1067 585
R9442 gnd.n1065 gnd.n1064 585
R9443 gnd.n1063 gnd.n1062 585
R9444 gnd.n1056 gnd.n1044 585
R9445 gnd.n1058 gnd.n1057 585
R9446 gnd.n1055 gnd.n1054 585
R9447 gnd.n1053 gnd.n1052 585
R9448 gnd.n1047 gnd.n1046 585
R9449 gnd.n1048 gnd.n1006 585
R9450 gnd.n6792 gnd.n1006 585
R9451 gnd.n2350 gnd.n1003 585
R9452 gnd.n6808 gnd.n1003 585
R9453 gnd.n2349 gnd.n2348 585
R9454 gnd.n2348 gnd.n1001 585
R9455 gnd.n2347 gnd.n1111 585
R9456 gnd.n2347 gnd.n2346 585
R9457 gnd.n2021 gnd.n989 585
R9458 gnd.n6816 gnd.n989 585
R9459 gnd.n2024 gnd.n2023 585
R9460 gnd.n2023 gnd.n2022 585
R9461 gnd.n2025 gnd.n978 585
R9462 gnd.n6822 gnd.n978 585
R9463 gnd.n2027 gnd.n2026 585
R9464 gnd.n2027 gnd.n976 585
R9465 gnd.n2029 gnd.n2028 585
R9466 gnd.n2028 gnd.n967 585
R9467 gnd.n2030 gnd.n965 585
R9468 gnd.n6830 gnd.n965 585
R9469 gnd.n2033 gnd.n2032 585
R9470 gnd.n2032 gnd.n2031 585
R9471 gnd.n2034 gnd.n954 585
R9472 gnd.n6836 gnd.n954 585
R9473 gnd.n2037 gnd.n2036 585
R9474 gnd.n2036 gnd.n2035 585
R9475 gnd.n2038 gnd.n1124 585
R9476 gnd.n2057 gnd.n1124 585
R9477 gnd.n2040 gnd.n2039 585
R9478 gnd.n2041 gnd.n2040 585
R9479 gnd.n1134 gnd.n1133 585
R9480 gnd.n1133 gnd.n1131 585
R9481 gnd.n2006 gnd.n2005 585
R9482 gnd.n2005 gnd.n2004 585
R9483 gnd.n1137 gnd.n1136 585
R9484 gnd.n1149 gnd.n1137 585
R9485 gnd.n1928 gnd.n1927 585
R9486 gnd.n1927 gnd.n1926 585
R9487 gnd.n1929 gnd.n1158 585
R9488 gnd.n1980 gnd.n1158 585
R9489 gnd.n1931 gnd.n1930 585
R9490 gnd.n1930 gnd.n1156 585
R9491 gnd.n1932 gnd.n1169 585
R9492 gnd.n1963 gnd.n1169 585
R9493 gnd.n1934 gnd.n1933 585
R9494 gnd.n1933 gnd.n1176 585
R9495 gnd.n1935 gnd.n1175 585
R9496 gnd.n1952 gnd.n1175 585
R9497 gnd.n1937 gnd.n1936 585
R9498 gnd.n1940 gnd.n1937 585
R9499 gnd.n1186 gnd.n1185 585
R9500 gnd.n1185 gnd.n1183 585
R9501 gnd.n1916 gnd.n1915 585
R9502 gnd.n1915 gnd.n1914 585
R9503 gnd.n1189 gnd.n1188 585
R9504 gnd.n1201 gnd.n1189 585
R9505 gnd.n1248 gnd.n1247 585
R9506 gnd.n1247 gnd.n1200 585
R9507 gnd.n1249 gnd.n1210 585
R9508 gnd.n1891 gnd.n1210 585
R9509 gnd.n1251 gnd.n1250 585
R9510 gnd.n1250 gnd.n1208 585
R9511 gnd.n1252 gnd.n1220 585
R9512 gnd.n1874 gnd.n1220 585
R9513 gnd.n1244 gnd.n1243 585
R9514 gnd.n1243 gnd.n1223 585
R9515 gnd.n1848 gnd.n1230 585
R9516 gnd.n1861 gnd.n1230 585
R9517 gnd.n1850 gnd.n1849 585
R9518 gnd.n1851 gnd.n1850 585
R9519 gnd.n1352 gnd.n1241 585
R9520 gnd.n1241 gnd.n1240 585
R9521 gnd.n1354 gnd.n1353 585
R9522 gnd.n1836 gnd.n1354 585
R9523 gnd.n1339 gnd.n1337 585
R9524 gnd.n1816 gnd.n1339 585
R9525 gnd.n1844 gnd.n1843 585
R9526 gnd.n1843 gnd.n1842 585
R9527 gnd.n1338 gnd.n1336 585
R9528 gnd.n1824 gnd.n1338 585
R9529 gnd.n1801 gnd.n1370 585
R9530 gnd.n1370 gnd.n1361 585
R9531 gnd.n1803 gnd.n1802 585
R9532 gnd.n1805 gnd.n1803 585
R9533 gnd.n1371 gnd.n1369 585
R9534 gnd.n1375 gnd.n1369 585
R9535 gnd.n1796 gnd.n1795 585
R9536 gnd.n1795 gnd.n1794 585
R9537 gnd.n1374 gnd.n1373 585
R9538 gnd.n1385 gnd.n1374 585
R9539 gnd.n1675 gnd.n1394 585
R9540 gnd.n1767 gnd.n1394 585
R9541 gnd.n1677 gnd.n1676 585
R9542 gnd.n1676 gnd.n1392 585
R9543 gnd.n1678 gnd.n1405 585
R9544 gnd.n1757 gnd.n1405 585
R9545 gnd.n1680 gnd.n1679 585
R9546 gnd.n1680 gnd.n1412 585
R9547 gnd.n1682 gnd.n1681 585
R9548 gnd.n1681 gnd.n1411 585
R9549 gnd.n1683 gnd.n1422 585
R9550 gnd.n1737 gnd.n1422 585
R9551 gnd.n1685 gnd.n1684 585
R9552 gnd.n1684 gnd.n1420 585
R9553 gnd.n1686 gnd.n1431 585
R9554 gnd.n1726 gnd.n1431 585
R9555 gnd.n1688 gnd.n1687 585
R9556 gnd.n1688 gnd.n1437 585
R9557 gnd.n1690 gnd.n1689 585
R9558 gnd.n1689 gnd.n1436 585
R9559 gnd.n1691 gnd.n1452 585
R9560 gnd.n1705 gnd.n1452 585
R9561 gnd.n1692 gnd.n1505 585
R9562 gnd.n1505 gnd.n1444 585
R9563 gnd.n1694 gnd.n1693 585
R9564 gnd.n1695 gnd.n1694 585
R9565 gnd.n1506 gnd.n1504 585
R9566 gnd.n1504 gnd.n1503 585
R9567 gnd.n1659 gnd.n1658 585
R9568 gnd.n1658 gnd.n1657 585
R9569 gnd.n1509 gnd.n1508 585
R9570 gnd.n1510 gnd.n1509 585
R9571 gnd.n1648 gnd.n1647 585
R9572 gnd.n1649 gnd.n1648 585
R9573 gnd.n1518 gnd.n1517 585
R9574 gnd.n1517 gnd.n1516 585
R9575 gnd.n1643 gnd.n1642 585
R9576 gnd.n1642 gnd.n1641 585
R9577 gnd.n1521 gnd.n1520 585
R9578 gnd.n1632 gnd.n1521 585
R9579 gnd.n1631 gnd.n1630 585
R9580 gnd.n1633 gnd.n1631 585
R9581 gnd.n1529 gnd.n1528 585
R9582 gnd.n1528 gnd.n1527 585
R9583 gnd.n246 gnd.n245 585
R9584 gnd.n249 gnd.n246 585
R9585 gnd.n7983 gnd.n7982 585
R9586 gnd.n7982 gnd.n7981 585
R9587 gnd.n7984 gnd.n241 585
R9588 gnd.n241 gnd.n240 585
R9589 gnd.n7986 gnd.n7985 585
R9590 gnd.n7987 gnd.n7986 585
R9591 gnd.n226 gnd.n225 585
R9592 gnd.n230 gnd.n226 585
R9593 gnd.n7995 gnd.n7994 585
R9594 gnd.n7994 gnd.n7993 585
R9595 gnd.n7996 gnd.n221 585
R9596 gnd.n227 gnd.n221 585
R9597 gnd.n7998 gnd.n7997 585
R9598 gnd.n7999 gnd.n7998 585
R9599 gnd.n208 gnd.n207 585
R9600 gnd.n211 gnd.n208 585
R9601 gnd.n8007 gnd.n8006 585
R9602 gnd.n8006 gnd.n8005 585
R9603 gnd.n8008 gnd.n203 585
R9604 gnd.n203 gnd.n202 585
R9605 gnd.n8010 gnd.n8009 585
R9606 gnd.n8011 gnd.n8010 585
R9607 gnd.n187 gnd.n186 585
R9608 gnd.n199 gnd.n187 585
R9609 gnd.n8019 gnd.n8018 585
R9610 gnd.n8018 gnd.n8017 585
R9611 gnd.n8020 gnd.n182 585
R9612 gnd.n188 gnd.n182 585
R9613 gnd.n8022 gnd.n8021 585
R9614 gnd.n8023 gnd.n8022 585
R9615 gnd.n168 gnd.n167 585
R9616 gnd.n7821 gnd.n168 585
R9617 gnd.n8031 gnd.n8030 585
R9618 gnd.n8030 gnd.n8029 585
R9619 gnd.n8032 gnd.n163 585
R9620 gnd.n7716 gnd.n163 585
R9621 gnd.n8034 gnd.n8033 585
R9622 gnd.n8035 gnd.n8034 585
R9623 gnd.n147 gnd.n146 585
R9624 gnd.n5872 gnd.n147 585
R9625 gnd.n8043 gnd.n8042 585
R9626 gnd.n8042 gnd.n8041 585
R9627 gnd.n8044 gnd.n142 585
R9628 gnd.n5878 gnd.n142 585
R9629 gnd.n8046 gnd.n8045 585
R9630 gnd.n8047 gnd.n8046 585
R9631 gnd.n129 gnd.n128 585
R9632 gnd.n5884 gnd.n129 585
R9633 gnd.n8055 gnd.n8054 585
R9634 gnd.n8054 gnd.n8053 585
R9635 gnd.n8056 gnd.n123 585
R9636 gnd.n5890 gnd.n123 585
R9637 gnd.n8058 gnd.n8057 585
R9638 gnd.n8059 gnd.n8058 585
R9639 gnd.n124 gnd.n122 585
R9640 gnd.n5829 gnd.n122 585
R9641 gnd.n5901 gnd.n5900 585
R9642 gnd.n5902 gnd.n5901 585
R9643 gnd.n3359 gnd.n104 585
R9644 gnd.n8067 gnd.n104 585
R9645 gnd.n5910 gnd.n5909 585
R9646 gnd.n5909 gnd.n5908 585
R9647 gnd.n5911 gnd.n3354 585
R9648 gnd.n3362 gnd.n3354 585
R9649 gnd.n5913 gnd.n5912 585
R9650 gnd.n5914 gnd.n5913 585
R9651 gnd.n3355 gnd.n3344 585
R9652 gnd.n5919 gnd.n3344 585
R9653 gnd.n5800 gnd.n5799 585
R9654 gnd.n5799 gnd.n3340 585
R9655 gnd.n5798 gnd.n5797 585
R9656 gnd.n5798 gnd.n3333 585
R9657 gnd.n3325 gnd.n3324 585
R9658 gnd.n5928 gnd.n3325 585
R9659 gnd.n5935 gnd.n5934 585
R9660 gnd.n5934 gnd.n5933 585
R9661 gnd.n5936 gnd.n3320 585
R9662 gnd.n5788 gnd.n3320 585
R9663 gnd.n5938 gnd.n5937 585
R9664 gnd.n5939 gnd.n5938 585
R9665 gnd.n3303 gnd.n3302 585
R9666 gnd.n5768 gnd.n3303 585
R9667 gnd.n5947 gnd.n5946 585
R9668 gnd.n5946 gnd.n5945 585
R9669 gnd.n5948 gnd.n3298 585
R9670 gnd.n5761 gnd.n3298 585
R9671 gnd.n5950 gnd.n5949 585
R9672 gnd.n5951 gnd.n5950 585
R9673 gnd.n3283 gnd.n3282 585
R9674 gnd.n5753 gnd.n3283 585
R9675 gnd.n5959 gnd.n5958 585
R9676 gnd.n5958 gnd.n5957 585
R9677 gnd.n5960 gnd.n3278 585
R9678 gnd.n5746 gnd.n3278 585
R9679 gnd.n5962 gnd.n5961 585
R9680 gnd.n5963 gnd.n5962 585
R9681 gnd.n3262 gnd.n3261 585
R9682 gnd.n5738 gnd.n3262 585
R9683 gnd.n5971 gnd.n5970 585
R9684 gnd.n5970 gnd.n5969 585
R9685 gnd.n5972 gnd.n3257 585
R9686 gnd.n5731 gnd.n3257 585
R9687 gnd.n5974 gnd.n5973 585
R9688 gnd.n5975 gnd.n5974 585
R9689 gnd.n3242 gnd.n3241 585
R9690 gnd.n5723 gnd.n3242 585
R9691 gnd.n5983 gnd.n5982 585
R9692 gnd.n5982 gnd.n5981 585
R9693 gnd.n5984 gnd.n3237 585
R9694 gnd.n5716 gnd.n3237 585
R9695 gnd.n5986 gnd.n5985 585
R9696 gnd.n5987 gnd.n5986 585
R9697 gnd.n3221 gnd.n3220 585
R9698 gnd.n5708 gnd.n3221 585
R9699 gnd.n5995 gnd.n5994 585
R9700 gnd.n5994 gnd.n5993 585
R9701 gnd.n5996 gnd.n3214 585
R9702 gnd.n5701 gnd.n3214 585
R9703 gnd.n5998 gnd.n5997 585
R9704 gnd.n5999 gnd.n5998 585
R9705 gnd.n3215 gnd.n3213 585
R9706 gnd.n5693 gnd.n3213 585
R9707 gnd.n3197 gnd.n3191 585
R9708 gnd.n6005 gnd.n3197 585
R9709 gnd.n6010 gnd.n3189 585
R9710 gnd.n5669 gnd.n3189 585
R9711 gnd.n6012 gnd.n6011 585
R9712 gnd.n6013 gnd.n6012 585
R9713 gnd.n3188 gnd.n3028 585
R9714 gnd.n6180 gnd.n3029 585
R9715 gnd.n6179 gnd.n3030 585
R9716 gnd.n3105 gnd.n3031 585
R9717 gnd.n6172 gnd.n3037 585
R9718 gnd.n6171 gnd.n3038 585
R9719 gnd.n3108 gnd.n3039 585
R9720 gnd.n6164 gnd.n3045 585
R9721 gnd.n6163 gnd.n3046 585
R9722 gnd.n3110 gnd.n3047 585
R9723 gnd.n6156 gnd.n3053 585
R9724 gnd.n6155 gnd.n3054 585
R9725 gnd.n3113 gnd.n3055 585
R9726 gnd.n6148 gnd.n3061 585
R9727 gnd.n6147 gnd.n3062 585
R9728 gnd.n3115 gnd.n3063 585
R9729 gnd.n6140 gnd.n3071 585
R9730 gnd.n6139 gnd.n6136 585
R9731 gnd.n3074 gnd.n3072 585
R9732 gnd.n6134 gnd.n3074 585
R9733 gnd.n7794 gnd.n7793 585
R9734 gnd.n7787 gnd.n7740 585
R9735 gnd.n7789 gnd.n7788 585
R9736 gnd.n7786 gnd.n7785 585
R9737 gnd.n7784 gnd.n7783 585
R9738 gnd.n7777 gnd.n7742 585
R9739 gnd.n7779 gnd.n7778 585
R9740 gnd.n7776 gnd.n7775 585
R9741 gnd.n7774 gnd.n7773 585
R9742 gnd.n7767 gnd.n7744 585
R9743 gnd.n7769 gnd.n7768 585
R9744 gnd.n7766 gnd.n7765 585
R9745 gnd.n7764 gnd.n7763 585
R9746 gnd.n7757 gnd.n7746 585
R9747 gnd.n7759 gnd.n7758 585
R9748 gnd.n7756 gnd.n7755 585
R9749 gnd.n7754 gnd.n7753 585
R9750 gnd.n7750 gnd.n7749 585
R9751 gnd.n7748 gnd.n257 585
R9752 gnd.n7973 gnd.n257 585
R9753 gnd.n7796 gnd.n7795 585
R9754 gnd.n7795 gnd.n249 585
R9755 gnd.n7797 gnd.n248 585
R9756 gnd.n7981 gnd.n248 585
R9757 gnd.n7799 gnd.n7798 585
R9758 gnd.n7798 gnd.n240 585
R9759 gnd.n7800 gnd.n239 585
R9760 gnd.n7987 gnd.n239 585
R9761 gnd.n7802 gnd.n7801 585
R9762 gnd.n7801 gnd.n230 585
R9763 gnd.n7803 gnd.n229 585
R9764 gnd.n7993 gnd.n229 585
R9765 gnd.n7805 gnd.n7804 585
R9766 gnd.n7804 gnd.n227 585
R9767 gnd.n7806 gnd.n220 585
R9768 gnd.n7999 gnd.n220 585
R9769 gnd.n7808 gnd.n7807 585
R9770 gnd.n7807 gnd.n211 585
R9771 gnd.n7809 gnd.n210 585
R9772 gnd.n8005 gnd.n210 585
R9773 gnd.n7811 gnd.n7810 585
R9774 gnd.n7810 gnd.n202 585
R9775 gnd.n7812 gnd.n201 585
R9776 gnd.n8011 gnd.n201 585
R9777 gnd.n7814 gnd.n7813 585
R9778 gnd.n7813 gnd.n199 585
R9779 gnd.n7815 gnd.n190 585
R9780 gnd.n8017 gnd.n190 585
R9781 gnd.n7817 gnd.n7816 585
R9782 gnd.n7816 gnd.n188 585
R9783 gnd.n7818 gnd.n181 585
R9784 gnd.n8023 gnd.n181 585
R9785 gnd.n7820 gnd.n7819 585
R9786 gnd.n7821 gnd.n7820 585
R9787 gnd.n357 gnd.n170 585
R9788 gnd.n8029 gnd.n170 585
R9789 gnd.n7718 gnd.n7717 585
R9790 gnd.n7717 gnd.n7716 585
R9791 gnd.n359 gnd.n161 585
R9792 gnd.n8035 gnd.n161 585
R9793 gnd.n5874 gnd.n5873 585
R9794 gnd.n5873 gnd.n5872 585
R9795 gnd.n5875 gnd.n150 585
R9796 gnd.n8041 gnd.n150 585
R9797 gnd.n5877 gnd.n5876 585
R9798 gnd.n5878 gnd.n5877 585
R9799 gnd.n5837 gnd.n141 585
R9800 gnd.n8047 gnd.n141 585
R9801 gnd.n5886 gnd.n5885 585
R9802 gnd.n5885 gnd.n5884 585
R9803 gnd.n5887 gnd.n131 585
R9804 gnd.n8053 gnd.n131 585
R9805 gnd.n5889 gnd.n5888 585
R9806 gnd.n5890 gnd.n5889 585
R9807 gnd.n5827 gnd.n120 585
R9808 gnd.n8059 gnd.n120 585
R9809 gnd.n5831 gnd.n5830 585
R9810 gnd.n5830 gnd.n5829 585
R9811 gnd.n100 gnd.n99 585
R9812 gnd.n5902 gnd.n100 585
R9813 gnd.n8069 gnd.n8068 585
R9814 gnd.n8068 gnd.n8067 585
R9815 gnd.n8070 gnd.n98 585
R9816 gnd.n5908 gnd.n98 585
R9817 gnd.n3361 gnd.n96 585
R9818 gnd.n3362 gnd.n3361 585
R9819 gnd.n5776 gnd.n3352 585
R9820 gnd.n5914 gnd.n3352 585
R9821 gnd.n5777 gnd.n3342 585
R9822 gnd.n5919 gnd.n3342 585
R9823 gnd.n5780 gnd.n5775 585
R9824 gnd.n5775 gnd.n3340 585
R9825 gnd.n5781 gnd.n5774 585
R9826 gnd.n5774 gnd.n3333 585
R9827 gnd.n5782 gnd.n3332 585
R9828 gnd.n5928 gnd.n3332 585
R9829 gnd.n3368 gnd.n3328 585
R9830 gnd.n5933 gnd.n3328 585
R9831 gnd.n5787 gnd.n5786 585
R9832 gnd.n5788 gnd.n5787 585
R9833 gnd.n3367 gnd.n3318 585
R9834 gnd.n5939 gnd.n3318 585
R9835 gnd.n5770 gnd.n5769 585
R9836 gnd.n5769 gnd.n5768 585
R9837 gnd.n3370 gnd.n3306 585
R9838 gnd.n5945 gnd.n3306 585
R9839 gnd.n5760 gnd.n5759 585
R9840 gnd.n5761 gnd.n5760 585
R9841 gnd.n3373 gnd.n3297 585
R9842 gnd.n5951 gnd.n3297 585
R9843 gnd.n5755 gnd.n5754 585
R9844 gnd.n5754 gnd.n5753 585
R9845 gnd.n3375 gnd.n3286 585
R9846 gnd.n5957 gnd.n3286 585
R9847 gnd.n5745 gnd.n5744 585
R9848 gnd.n5746 gnd.n5745 585
R9849 gnd.n3377 gnd.n3276 585
R9850 gnd.n5963 gnd.n3276 585
R9851 gnd.n5740 gnd.n5739 585
R9852 gnd.n5739 gnd.n5738 585
R9853 gnd.n3379 gnd.n3265 585
R9854 gnd.n5969 gnd.n3265 585
R9855 gnd.n5730 gnd.n5729 585
R9856 gnd.n5731 gnd.n5730 585
R9857 gnd.n3382 gnd.n3256 585
R9858 gnd.n5975 gnd.n3256 585
R9859 gnd.n5725 gnd.n5724 585
R9860 gnd.n5724 gnd.n5723 585
R9861 gnd.n3384 gnd.n3245 585
R9862 gnd.n5981 gnd.n3245 585
R9863 gnd.n5715 gnd.n5714 585
R9864 gnd.n5716 gnd.n5715 585
R9865 gnd.n3386 gnd.n3235 585
R9866 gnd.n5987 gnd.n3235 585
R9867 gnd.n5710 gnd.n5709 585
R9868 gnd.n5709 gnd.n5708 585
R9869 gnd.n3388 gnd.n3224 585
R9870 gnd.n5993 gnd.n3224 585
R9871 gnd.n5700 gnd.n5699 585
R9872 gnd.n5701 gnd.n5700 585
R9873 gnd.n3390 gnd.n3211 585
R9874 gnd.n5999 gnd.n3211 585
R9875 gnd.n5695 gnd.n5694 585
R9876 gnd.n5694 gnd.n5693 585
R9877 gnd.n5692 gnd.n3195 585
R9878 gnd.n6005 gnd.n3195 585
R9879 gnd.n5691 gnd.n3393 585
R9880 gnd.n5669 gnd.n3393 585
R9881 gnd.n3392 gnd.n3186 585
R9882 gnd.n6013 gnd.n3186 585
R9883 gnd.n1000 gnd.n999 585
R9884 gnd.n1004 gnd.n1000 585
R9885 gnd.n6811 gnd.n6810 585
R9886 gnd.n6810 gnd.n6809 585
R9887 gnd.n6812 gnd.n992 585
R9888 gnd.n2345 gnd.n992 585
R9889 gnd.n6814 gnd.n6813 585
R9890 gnd.n6815 gnd.n6814 585
R9891 gnd.n993 gnd.n991 585
R9892 gnd.n991 gnd.n988 585
R9893 gnd.n975 gnd.n974 585
R9894 gnd.n979 gnd.n975 585
R9895 gnd.n6825 gnd.n6824 585
R9896 gnd.n6824 gnd.n6823 585
R9897 gnd.n6826 gnd.n969 585
R9898 gnd.n1112 gnd.n969 585
R9899 gnd.n6828 gnd.n6827 585
R9900 gnd.n6829 gnd.n6828 585
R9901 gnd.n970 gnd.n968 585
R9902 gnd.n968 gnd.n964 585
R9903 gnd.n2052 gnd.n2051 585
R9904 gnd.n2051 gnd.n955 585
R9905 gnd.n2053 gnd.n1126 585
R9906 gnd.n1126 gnd.n953 585
R9907 gnd.n2055 gnd.n2054 585
R9908 gnd.n2056 gnd.n2055 585
R9909 gnd.n1127 gnd.n1125 585
R9910 gnd.n1125 gnd.n1123 585
R9911 gnd.n2044 gnd.n2043 585
R9912 gnd.n2043 gnd.n2042 585
R9913 gnd.n1130 gnd.n1129 585
R9914 gnd.n1139 gnd.n1130 585
R9915 gnd.n1988 gnd.n1151 585
R9916 gnd.n1151 gnd.n1138 585
R9917 gnd.n1990 gnd.n1989 585
R9918 gnd.n1991 gnd.n1990 585
R9919 gnd.n1152 gnd.n1150 585
R9920 gnd.n1159 gnd.n1150 585
R9921 gnd.n1983 gnd.n1982 585
R9922 gnd.n1982 gnd.n1981 585
R9923 gnd.n1155 gnd.n1154 585
R9924 gnd.n1962 gnd.n1155 585
R9925 gnd.n1948 gnd.n1178 585
R9926 gnd.n1178 gnd.n1168 585
R9927 gnd.n1950 gnd.n1949 585
R9928 gnd.n1951 gnd.n1950 585
R9929 gnd.n1179 gnd.n1177 585
R9930 gnd.n1939 gnd.n1177 585
R9931 gnd.n1943 gnd.n1942 585
R9932 gnd.n1942 gnd.n1941 585
R9933 gnd.n1182 gnd.n1181 585
R9934 gnd.n1905 gnd.n1182 585
R9935 gnd.n1899 gnd.n1203 585
R9936 gnd.n1203 gnd.n1190 585
R9937 gnd.n1901 gnd.n1900 585
R9938 gnd.n1902 gnd.n1901 585
R9939 gnd.n1204 gnd.n1202 585
R9940 gnd.n1211 gnd.n1202 585
R9941 gnd.n1894 gnd.n1893 585
R9942 gnd.n1893 gnd.n1892 585
R9943 gnd.n1207 gnd.n1206 585
R9944 gnd.n1873 gnd.n1207 585
R9945 gnd.n1869 gnd.n1868 585
R9946 gnd.n1870 gnd.n1869 585
R9947 gnd.n1225 gnd.n1224 585
R9948 gnd.n1231 gnd.n1224 585
R9949 gnd.n1864 gnd.n1863 585
R9950 gnd.n1863 gnd.n1862 585
R9951 gnd.n1228 gnd.n1227 585
R9952 gnd.n1852 gnd.n1228 585
R9953 gnd.n1834 gnd.n1833 585
R9954 gnd.n1835 gnd.n1834 585
R9955 gnd.n1356 gnd.n1355 585
R9956 gnd.n1817 gnd.n1355 585
R9957 gnd.n1829 gnd.n1828 585
R9958 gnd.n1828 gnd.n1341 585
R9959 gnd.n1827 gnd.n1358 585
R9960 gnd.n1827 gnd.n1340 585
R9961 gnd.n1826 gnd.n1360 585
R9962 gnd.n1826 gnd.n1825 585
R9963 gnd.n1778 gnd.n1359 585
R9964 gnd.n1804 gnd.n1359 585
R9965 gnd.n1780 gnd.n1779 585
R9966 gnd.n1779 gnd.n1368 585
R9967 gnd.n1781 gnd.n1387 585
R9968 gnd.n1387 gnd.n1376 585
R9969 gnd.n1783 gnd.n1782 585
R9970 gnd.n1784 gnd.n1783 585
R9971 gnd.n1388 gnd.n1386 585
R9972 gnd.n1395 gnd.n1386 585
R9973 gnd.n1770 gnd.n1769 585
R9974 gnd.n1769 gnd.n1768 585
R9975 gnd.n1391 gnd.n1390 585
R9976 gnd.n1758 gnd.n1391 585
R9977 gnd.n1745 gnd.n1415 585
R9978 gnd.n1415 gnd.n1414 585
R9979 gnd.n1747 gnd.n1746 585
R9980 gnd.n1748 gnd.n1747 585
R9981 gnd.n1416 gnd.n1413 585
R9982 gnd.n1423 gnd.n1413 585
R9983 gnd.n1740 gnd.n1739 585
R9984 gnd.n1739 gnd.n1738 585
R9985 gnd.n1419 gnd.n1418 585
R9986 gnd.n1727 gnd.n1419 585
R9987 gnd.n1714 gnd.n1440 585
R9988 gnd.n1440 gnd.n1439 585
R9989 gnd.n1716 gnd.n1715 585
R9990 gnd.n1717 gnd.n1716 585
R9991 gnd.n1710 gnd.n1438 585
R9992 gnd.n1709 gnd.n1708 585
R9993 gnd.n1443 gnd.n1442 585
R9994 gnd.n1706 gnd.n1443 585
R9995 gnd.n1465 gnd.n1464 585
R9996 gnd.n1468 gnd.n1467 585
R9997 gnd.n1466 gnd.n1461 585
R9998 gnd.n1473 gnd.n1472 585
R9999 gnd.n1475 gnd.n1474 585
R10000 gnd.n1478 gnd.n1477 585
R10001 gnd.n1476 gnd.n1459 585
R10002 gnd.n1483 gnd.n1482 585
R10003 gnd.n1485 gnd.n1484 585
R10004 gnd.n1488 gnd.n1487 585
R10005 gnd.n1486 gnd.n1457 585
R10006 gnd.n1493 gnd.n1492 585
R10007 gnd.n1497 gnd.n1494 585
R10008 gnd.n1498 gnd.n1435 585
R10009 gnd.n6801 gnd.n6800 585
R10010 gnd.n6794 gnd.n1014 585
R10011 gnd.n6796 gnd.n6795 585
R10012 gnd.n1017 gnd.n1016 585
R10013 gnd.n6766 gnd.n6765 585
R10014 gnd.n6768 gnd.n6767 585
R10015 gnd.n6770 gnd.n6769 585
R10016 gnd.n6772 gnd.n6771 585
R10017 gnd.n6774 gnd.n6773 585
R10018 gnd.n6776 gnd.n6775 585
R10019 gnd.n6778 gnd.n6777 585
R10020 gnd.n6780 gnd.n6779 585
R10021 gnd.n6782 gnd.n6781 585
R10022 gnd.n6785 gnd.n6784 585
R10023 gnd.n6783 gnd.n6755 585
R10024 gnd.n6789 gnd.n6752 585
R10025 gnd.n6791 gnd.n6790 585
R10026 gnd.n6792 gnd.n6791 585
R10027 gnd.n6803 gnd.n6802 585
R10028 gnd.n6802 gnd.n1004 585
R10029 gnd.n1010 gnd.n1002 585
R10030 gnd.n6809 gnd.n1002 585
R10031 gnd.n2344 gnd.n2343 585
R10032 gnd.n2345 gnd.n2344 585
R10033 gnd.n2338 gnd.n990 585
R10034 gnd.n6815 gnd.n990 585
R10035 gnd.n2337 gnd.n2336 585
R10036 gnd.n2336 gnd.n988 585
R10037 gnd.n2335 gnd.n2333 585
R10038 gnd.n2335 gnd.n979 585
R10039 gnd.n2075 gnd.n977 585
R10040 gnd.n6823 gnd.n977 585
R10041 gnd.n1114 gnd.n1113 585
R10042 gnd.n1113 gnd.n1112 585
R10043 gnd.n2069 gnd.n966 585
R10044 gnd.n6829 gnd.n966 585
R10045 gnd.n2068 gnd.n2067 585
R10046 gnd.n2067 gnd.n964 585
R10047 gnd.n2066 gnd.n1116 585
R10048 gnd.n2066 gnd.n955 585
R10049 gnd.n2065 gnd.n2064 585
R10050 gnd.n2065 gnd.n953 585
R10051 gnd.n1119 gnd.n1118 585
R10052 gnd.n2056 gnd.n1118 585
R10053 gnd.n1997 gnd.n1996 585
R10054 gnd.n1996 gnd.n1123 585
R10055 gnd.n1998 gnd.n1132 585
R10056 gnd.n2042 gnd.n1132 585
R10057 gnd.n1995 gnd.n1994 585
R10058 gnd.n1994 gnd.n1139 585
R10059 gnd.n1993 gnd.n1146 585
R10060 gnd.n1993 gnd.n1138 585
R10061 gnd.n1992 gnd.n1148 585
R10062 gnd.n1992 gnd.n1991 585
R10063 gnd.n1971 gnd.n1147 585
R10064 gnd.n1159 gnd.n1147 585
R10065 gnd.n1970 gnd.n1157 585
R10066 gnd.n1981 gnd.n1157 585
R10067 gnd.n1961 gnd.n1164 585
R10068 gnd.n1962 gnd.n1961 585
R10069 gnd.n1960 gnd.n1959 585
R10070 gnd.n1960 gnd.n1168 585
R10071 gnd.n1958 gnd.n1170 585
R10072 gnd.n1951 gnd.n1170 585
R10073 gnd.n1938 gnd.n1171 585
R10074 gnd.n1939 gnd.n1938 585
R10075 gnd.n1908 gnd.n1184 585
R10076 gnd.n1941 gnd.n1184 585
R10077 gnd.n1907 gnd.n1906 585
R10078 gnd.n1906 gnd.n1905 585
R10079 gnd.n1904 gnd.n1197 585
R10080 gnd.n1904 gnd.n1190 585
R10081 gnd.n1903 gnd.n1199 585
R10082 gnd.n1903 gnd.n1902 585
R10083 gnd.n1882 gnd.n1198 585
R10084 gnd.n1211 gnd.n1198 585
R10085 gnd.n1881 gnd.n1209 585
R10086 gnd.n1892 gnd.n1209 585
R10087 gnd.n1872 gnd.n1216 585
R10088 gnd.n1873 gnd.n1872 585
R10089 gnd.n1871 gnd.n1222 585
R10090 gnd.n1871 gnd.n1870 585
R10091 gnd.n1856 gnd.n1221 585
R10092 gnd.n1231 gnd.n1221 585
R10093 gnd.n1855 gnd.n1229 585
R10094 gnd.n1862 gnd.n1229 585
R10095 gnd.n1854 gnd.n1853 585
R10096 gnd.n1853 gnd.n1852 585
R10097 gnd.n1239 gnd.n1236 585
R10098 gnd.n1835 gnd.n1239 585
R10099 gnd.n1818 gnd.n1815 585
R10100 gnd.n1818 gnd.n1817 585
R10101 gnd.n1820 gnd.n1819 585
R10102 gnd.n1819 gnd.n1341 585
R10103 gnd.n1821 gnd.n1363 585
R10104 gnd.n1363 gnd.n1340 585
R10105 gnd.n1823 gnd.n1822 585
R10106 gnd.n1825 gnd.n1823 585
R10107 gnd.n1364 gnd.n1362 585
R10108 gnd.n1804 gnd.n1362 585
R10109 gnd.n1788 gnd.n1787 585
R10110 gnd.n1787 gnd.n1368 585
R10111 gnd.n1786 gnd.n1382 585
R10112 gnd.n1786 gnd.n1376 585
R10113 gnd.n1785 gnd.n1384 585
R10114 gnd.n1785 gnd.n1784 585
R10115 gnd.n1762 gnd.n1383 585
R10116 gnd.n1395 gnd.n1383 585
R10117 gnd.n1761 gnd.n1393 585
R10118 gnd.n1768 gnd.n1393 585
R10119 gnd.n1760 gnd.n1759 585
R10120 gnd.n1759 gnd.n1758 585
R10121 gnd.n1404 gnd.n1401 585
R10122 gnd.n1414 gnd.n1404 585
R10123 gnd.n1750 gnd.n1749 585
R10124 gnd.n1749 gnd.n1748 585
R10125 gnd.n1410 gnd.n1409 585
R10126 gnd.n1423 gnd.n1410 585
R10127 gnd.n1730 gnd.n1421 585
R10128 gnd.n1738 gnd.n1421 585
R10129 gnd.n1729 gnd.n1728 585
R10130 gnd.n1728 gnd.n1727 585
R10131 gnd.n1430 gnd.n1428 585
R10132 gnd.n1439 gnd.n1430 585
R10133 gnd.n1719 gnd.n1718 585
R10134 gnd.n1718 gnd.n1717 585
R10135 gnd.n5540 gnd.n5539 585
R10136 gnd.n5539 gnd.n3445 585
R10137 gnd.n5541 gnd.n3459 585
R10138 gnd.n3459 gnd.n3457 585
R10139 gnd.n5543 gnd.n5542 585
R10140 gnd.n5544 gnd.n5543 585
R10141 gnd.n3460 gnd.n3458 585
R10142 gnd.n5415 gnd.n3458 585
R10143 gnd.n3562 gnd.n3561 585
R10144 gnd.n3561 gnd.n3537 585
R10145 gnd.n5387 gnd.n3563 585
R10146 gnd.n5387 gnd.n5386 585
R10147 gnd.n5388 gnd.n3560 585
R10148 gnd.n5388 gnd.n3545 585
R10149 gnd.n5390 gnd.n5389 585
R10150 gnd.n5389 gnd.n3544 585
R10151 gnd.n5391 gnd.n3558 585
R10152 gnd.n5379 gnd.n3558 585
R10153 gnd.n5393 gnd.n5392 585
R10154 gnd.n5394 gnd.n5393 585
R10155 gnd.n3559 gnd.n3557 585
R10156 gnd.n3557 gnd.n3553 585
R10157 gnd.n5372 gnd.n5371 585
R10158 gnd.n5373 gnd.n5372 585
R10159 gnd.n5370 gnd.n3569 585
R10160 gnd.n3575 gnd.n3569 585
R10161 gnd.n5369 gnd.n5368 585
R10162 gnd.n5368 gnd.n5367 585
R10163 gnd.n3571 gnd.n3570 585
R10164 gnd.n3572 gnd.n3571 585
R10165 gnd.n5357 gnd.n5356 585
R10166 gnd.n5358 gnd.n5357 585
R10167 gnd.n5355 gnd.n3586 585
R10168 gnd.n3586 gnd.n3582 585
R10169 gnd.n5354 gnd.n5353 585
R10170 gnd.n5353 gnd.n5352 585
R10171 gnd.n3588 gnd.n3587 585
R10172 gnd.n3594 gnd.n3588 585
R10173 gnd.n5339 gnd.n5338 585
R10174 gnd.n5340 gnd.n5339 585
R10175 gnd.n5337 gnd.n3597 585
R10176 gnd.n3603 gnd.n3597 585
R10177 gnd.n5336 gnd.n5335 585
R10178 gnd.n5335 gnd.n5334 585
R10179 gnd.n3599 gnd.n3598 585
R10180 gnd.n3614 gnd.n3599 585
R10181 gnd.n5311 gnd.n3611 585
R10182 gnd.n5323 gnd.n3611 585
R10183 gnd.n5312 gnd.n3622 585
R10184 gnd.n3622 gnd.n3610 585
R10185 gnd.n5314 gnd.n5313 585
R10186 gnd.n5315 gnd.n5314 585
R10187 gnd.n5310 gnd.n3621 585
R10188 gnd.n5306 gnd.n3621 585
R10189 gnd.n5309 gnd.n5308 585
R10190 gnd.n5308 gnd.n5307 585
R10191 gnd.n3624 gnd.n3623 585
R10192 gnd.n3630 gnd.n3624 585
R10193 gnd.n5299 gnd.n5298 585
R10194 gnd.n5300 gnd.n5299 585
R10195 gnd.n5297 gnd.n3632 585
R10196 gnd.n3632 gnd.n3629 585
R10197 gnd.n5296 gnd.n5295 585
R10198 gnd.n5295 gnd.n5294 585
R10199 gnd.n3634 gnd.n3633 585
R10200 gnd.n3646 gnd.n3634 585
R10201 gnd.n5275 gnd.n5274 585
R10202 gnd.n5276 gnd.n5275 585
R10203 gnd.n5273 gnd.n3647 585
R10204 gnd.n5268 gnd.n3647 585
R10205 gnd.n5272 gnd.n5271 585
R10206 gnd.n5271 gnd.n5270 585
R10207 gnd.n3649 gnd.n3648 585
R10208 gnd.n3650 gnd.n3649 585
R10209 gnd.n5256 gnd.n5255 585
R10210 gnd.n5257 gnd.n5256 585
R10211 gnd.n5254 gnd.n3657 585
R10212 gnd.n5250 gnd.n3657 585
R10213 gnd.n5253 gnd.n5252 585
R10214 gnd.n5252 gnd.n5251 585
R10215 gnd.n3659 gnd.n3658 585
R10216 gnd.n5238 gnd.n3659 585
R10217 gnd.n5227 gnd.n3677 585
R10218 gnd.n3677 gnd.n3675 585
R10219 gnd.n5229 gnd.n5228 585
R10220 gnd.n5230 gnd.n5229 585
R10221 gnd.n5226 gnd.n3676 585
R10222 gnd.n3682 gnd.n3676 585
R10223 gnd.n5225 gnd.n5224 585
R10224 gnd.n5224 gnd.n5223 585
R10225 gnd.n3679 gnd.n3678 585
R10226 gnd.n5200 gnd.n3679 585
R10227 gnd.n5212 gnd.n5211 585
R10228 gnd.n5213 gnd.n5212 585
R10229 gnd.n5210 gnd.n3692 585
R10230 gnd.n3692 gnd.n3688 585
R10231 gnd.n5209 gnd.n5208 585
R10232 gnd.n5208 gnd.n5207 585
R10233 gnd.n3694 gnd.n3693 585
R10234 gnd.n3695 gnd.n3694 585
R10235 gnd.n5194 gnd.n5193 585
R10236 gnd.n5195 gnd.n5194 585
R10237 gnd.n5192 gnd.n3704 585
R10238 gnd.n5188 gnd.n3704 585
R10239 gnd.n5191 gnd.n5190 585
R10240 gnd.n5190 gnd.n5189 585
R10241 gnd.n3706 gnd.n3705 585
R10242 gnd.n3712 gnd.n3706 585
R10243 gnd.n5181 gnd.n5180 585
R10244 gnd.n5182 gnd.n5181 585
R10245 gnd.n5179 gnd.n3715 585
R10246 gnd.n3715 gnd.n3711 585
R10247 gnd.n5178 gnd.n5177 585
R10248 gnd.n5177 gnd.n5176 585
R10249 gnd.n3717 gnd.n3716 585
R10250 gnd.n3729 gnd.n3717 585
R10251 gnd.n5154 gnd.n5153 585
R10252 gnd.n5155 gnd.n5154 585
R10253 gnd.n5152 gnd.n3730 585
R10254 gnd.n5146 gnd.n3730 585
R10255 gnd.n5151 gnd.n5150 585
R10256 gnd.n5150 gnd.n5149 585
R10257 gnd.n3732 gnd.n3731 585
R10258 gnd.n3733 gnd.n3732 585
R10259 gnd.n5134 gnd.n5133 585
R10260 gnd.n5135 gnd.n5134 585
R10261 gnd.n5132 gnd.n3739 585
R10262 gnd.n5128 gnd.n3739 585
R10263 gnd.n5131 gnd.n5130 585
R10264 gnd.n5130 gnd.n5129 585
R10265 gnd.n3741 gnd.n3740 585
R10266 gnd.n5115 gnd.n3741 585
R10267 gnd.n5104 gnd.n3758 585
R10268 gnd.n3758 gnd.n3756 585
R10269 gnd.n5106 gnd.n5105 585
R10270 gnd.n5107 gnd.n5106 585
R10271 gnd.n5103 gnd.n3757 585
R10272 gnd.n3763 gnd.n3757 585
R10273 gnd.n5102 gnd.n5101 585
R10274 gnd.n5101 gnd.n5100 585
R10275 gnd.n3760 gnd.n3759 585
R10276 gnd.n5076 gnd.n3760 585
R10277 gnd.n5088 gnd.n5087 585
R10278 gnd.n5089 gnd.n5088 585
R10279 gnd.n5086 gnd.n3772 585
R10280 gnd.n3776 gnd.n3772 585
R10281 gnd.n5085 gnd.n5084 585
R10282 gnd.n5084 gnd.n5083 585
R10283 gnd.n3774 gnd.n3773 585
R10284 gnd.n3782 gnd.n3774 585
R10285 gnd.n5070 gnd.n5069 585
R10286 gnd.n5071 gnd.n5070 585
R10287 gnd.n5068 gnd.n3784 585
R10288 gnd.n5064 gnd.n3784 585
R10289 gnd.n5067 gnd.n5066 585
R10290 gnd.n5066 gnd.n5065 585
R10291 gnd.n3786 gnd.n3785 585
R10292 gnd.n3793 gnd.n3786 585
R10293 gnd.n5057 gnd.n5056 585
R10294 gnd.n5058 gnd.n5057 585
R10295 gnd.n5055 gnd.n3795 585
R10296 gnd.n3795 gnd.n3792 585
R10297 gnd.n5054 gnd.n5053 585
R10298 gnd.n5053 gnd.n5052 585
R10299 gnd.n3797 gnd.n3796 585
R10300 gnd.n3809 gnd.n3797 585
R10301 gnd.n5030 gnd.n5029 585
R10302 gnd.n5031 gnd.n5030 585
R10303 gnd.n5028 gnd.n3810 585
R10304 gnd.n5023 gnd.n3810 585
R10305 gnd.n5027 gnd.n5026 585
R10306 gnd.n5026 gnd.n5025 585
R10307 gnd.n3812 gnd.n3811 585
R10308 gnd.n5013 gnd.n3812 585
R10309 gnd.n5002 gnd.n5001 585
R10310 gnd.n5003 gnd.n5002 585
R10311 gnd.n5000 gnd.n3820 585
R10312 gnd.n3820 gnd.n3818 585
R10313 gnd.n4999 gnd.n4998 585
R10314 gnd.n4998 gnd.n4997 585
R10315 gnd.n3822 gnd.n3821 585
R10316 gnd.n3822 gnd.n2912 585
R10317 gnd.n4989 gnd.n4988 585
R10318 gnd.n4990 gnd.n4989 585
R10319 gnd.n4987 gnd.n4984 585
R10320 gnd.n4984 gnd.n4983 585
R10321 gnd.n4986 gnd.n4985 585
R10322 gnd.n4985 gnd.n2901 585
R10323 gnd.n2896 gnd.n2895 585
R10324 gnd.n6319 gnd.n2896 585
R10325 gnd.n6322 gnd.n6321 585
R10326 gnd.n6321 gnd.n6320 585
R10327 gnd.n6323 gnd.n2874 585
R10328 gnd.n3892 gnd.n2874 585
R10329 gnd.n6388 gnd.n6387 585
R10330 gnd.n6386 gnd.n2873 585
R10331 gnd.n6385 gnd.n2872 585
R10332 gnd.n6390 gnd.n2872 585
R10333 gnd.n6384 gnd.n6383 585
R10334 gnd.n6382 gnd.n6381 585
R10335 gnd.n6380 gnd.n6379 585
R10336 gnd.n6378 gnd.n6377 585
R10337 gnd.n6376 gnd.n6375 585
R10338 gnd.n6374 gnd.n6373 585
R10339 gnd.n6372 gnd.n6371 585
R10340 gnd.n6370 gnd.n6369 585
R10341 gnd.n6368 gnd.n6367 585
R10342 gnd.n6366 gnd.n6365 585
R10343 gnd.n6364 gnd.n6363 585
R10344 gnd.n6362 gnd.n6361 585
R10345 gnd.n6360 gnd.n6359 585
R10346 gnd.n6358 gnd.n6357 585
R10347 gnd.n6356 gnd.n6355 585
R10348 gnd.n6354 gnd.n6353 585
R10349 gnd.n6352 gnd.n6351 585
R10350 gnd.n6350 gnd.n6349 585
R10351 gnd.n6348 gnd.n6347 585
R10352 gnd.n6346 gnd.n6345 585
R10353 gnd.n6344 gnd.n6343 585
R10354 gnd.n6342 gnd.n6341 585
R10355 gnd.n6340 gnd.n6339 585
R10356 gnd.n6338 gnd.n6337 585
R10357 gnd.n6336 gnd.n6335 585
R10358 gnd.n6334 gnd.n6333 585
R10359 gnd.n6332 gnd.n6331 585
R10360 gnd.n6330 gnd.n6329 585
R10361 gnd.n6328 gnd.n2836 585
R10362 gnd.n6393 gnd.n6392 585
R10363 gnd.n2838 gnd.n2835 585
R10364 gnd.n3830 gnd.n3829 585
R10365 gnd.n3832 gnd.n3831 585
R10366 gnd.n3835 gnd.n3834 585
R10367 gnd.n3837 gnd.n3836 585
R10368 gnd.n3839 gnd.n3838 585
R10369 gnd.n3841 gnd.n3840 585
R10370 gnd.n3843 gnd.n3842 585
R10371 gnd.n3845 gnd.n3844 585
R10372 gnd.n3847 gnd.n3846 585
R10373 gnd.n3849 gnd.n3848 585
R10374 gnd.n3851 gnd.n3850 585
R10375 gnd.n3853 gnd.n3852 585
R10376 gnd.n3855 gnd.n3854 585
R10377 gnd.n3857 gnd.n3856 585
R10378 gnd.n3859 gnd.n3858 585
R10379 gnd.n3861 gnd.n3860 585
R10380 gnd.n3863 gnd.n3862 585
R10381 gnd.n3865 gnd.n3864 585
R10382 gnd.n3867 gnd.n3866 585
R10383 gnd.n3869 gnd.n3868 585
R10384 gnd.n3871 gnd.n3870 585
R10385 gnd.n3873 gnd.n3872 585
R10386 gnd.n3875 gnd.n3874 585
R10387 gnd.n3877 gnd.n3876 585
R10388 gnd.n3879 gnd.n3878 585
R10389 gnd.n3881 gnd.n3880 585
R10390 gnd.n3883 gnd.n3882 585
R10391 gnd.n3885 gnd.n3884 585
R10392 gnd.n3887 gnd.n3886 585
R10393 gnd.n3889 gnd.n3888 585
R10394 gnd.n3891 gnd.n3890 585
R10395 gnd.n5423 gnd.n5422 585
R10396 gnd.n5424 gnd.n3532 585
R10397 gnd.n5426 gnd.n5425 585
R10398 gnd.n5428 gnd.n3530 585
R10399 gnd.n5430 gnd.n5429 585
R10400 gnd.n5431 gnd.n3529 585
R10401 gnd.n5433 gnd.n5432 585
R10402 gnd.n5435 gnd.n3527 585
R10403 gnd.n5437 gnd.n5436 585
R10404 gnd.n5438 gnd.n3526 585
R10405 gnd.n5440 gnd.n5439 585
R10406 gnd.n5442 gnd.n3524 585
R10407 gnd.n5444 gnd.n5443 585
R10408 gnd.n5445 gnd.n3523 585
R10409 gnd.n5447 gnd.n5446 585
R10410 gnd.n5449 gnd.n3521 585
R10411 gnd.n5451 gnd.n5450 585
R10412 gnd.n5452 gnd.n3520 585
R10413 gnd.n5454 gnd.n5453 585
R10414 gnd.n5456 gnd.n3518 585
R10415 gnd.n5458 gnd.n5457 585
R10416 gnd.n5459 gnd.n3517 585
R10417 gnd.n5461 gnd.n5460 585
R10418 gnd.n5463 gnd.n3515 585
R10419 gnd.n5465 gnd.n5464 585
R10420 gnd.n5466 gnd.n3514 585
R10421 gnd.n5468 gnd.n5467 585
R10422 gnd.n5470 gnd.n3512 585
R10423 gnd.n5472 gnd.n5471 585
R10424 gnd.n5474 gnd.n3509 585
R10425 gnd.n5476 gnd.n5475 585
R10426 gnd.n5478 gnd.n3508 585
R10427 gnd.n5479 gnd.n3447 585
R10428 gnd.n5482 gnd.n3149 585
R10429 gnd.n5484 gnd.n5483 585
R10430 gnd.n5485 gnd.n3503 585
R10431 gnd.n5487 gnd.n5486 585
R10432 gnd.n5489 gnd.n3501 585
R10433 gnd.n5491 gnd.n5490 585
R10434 gnd.n5492 gnd.n3500 585
R10435 gnd.n5494 gnd.n5493 585
R10436 gnd.n5496 gnd.n3498 585
R10437 gnd.n5498 gnd.n5497 585
R10438 gnd.n5499 gnd.n3497 585
R10439 gnd.n5501 gnd.n5500 585
R10440 gnd.n5503 gnd.n3495 585
R10441 gnd.n5505 gnd.n5504 585
R10442 gnd.n5506 gnd.n3494 585
R10443 gnd.n5508 gnd.n5507 585
R10444 gnd.n5510 gnd.n3492 585
R10445 gnd.n5512 gnd.n5511 585
R10446 gnd.n5513 gnd.n3491 585
R10447 gnd.n5515 gnd.n5514 585
R10448 gnd.n5517 gnd.n3489 585
R10449 gnd.n5519 gnd.n5518 585
R10450 gnd.n5520 gnd.n3488 585
R10451 gnd.n5522 gnd.n5521 585
R10452 gnd.n5524 gnd.n3486 585
R10453 gnd.n5526 gnd.n5525 585
R10454 gnd.n5527 gnd.n3485 585
R10455 gnd.n5529 gnd.n5528 585
R10456 gnd.n5531 gnd.n3483 585
R10457 gnd.n5533 gnd.n5532 585
R10458 gnd.n5534 gnd.n3482 585
R10459 gnd.n5536 gnd.n5535 585
R10460 gnd.n5538 gnd.n3481 585
R10461 gnd.n5421 gnd.n3533 585
R10462 gnd.n5421 gnd.n3445 585
R10463 gnd.n5420 gnd.n5419 585
R10464 gnd.n5420 gnd.n3457 585
R10465 gnd.n5418 gnd.n3454 585
R10466 gnd.n5544 gnd.n3454 585
R10467 gnd.n5417 gnd.n5416 585
R10468 gnd.n5416 gnd.n5415 585
R10469 gnd.n3536 gnd.n3535 585
R10470 gnd.n3537 gnd.n3536 585
R10471 gnd.n5385 gnd.n5384 585
R10472 gnd.n5386 gnd.n5385 585
R10473 gnd.n5383 gnd.n3565 585
R10474 gnd.n3565 gnd.n3545 585
R10475 gnd.n5382 gnd.n5381 585
R10476 gnd.n5381 gnd.n3544 585
R10477 gnd.n5380 gnd.n5378 585
R10478 gnd.n5380 gnd.n5379 585
R10479 gnd.n5377 gnd.n3555 585
R10480 gnd.n5394 gnd.n3555 585
R10481 gnd.n5376 gnd.n5375 585
R10482 gnd.n5375 gnd.n3553 585
R10483 gnd.n5374 gnd.n3566 585
R10484 gnd.n5374 gnd.n5373 585
R10485 gnd.n5344 gnd.n3567 585
R10486 gnd.n3575 gnd.n3567 585
R10487 gnd.n5345 gnd.n3573 585
R10488 gnd.n5367 gnd.n3573 585
R10489 gnd.n5347 gnd.n5346 585
R10490 gnd.n5346 gnd.n3572 585
R10491 gnd.n5348 gnd.n3584 585
R10492 gnd.n5358 gnd.n3584 585
R10493 gnd.n5349 gnd.n3591 585
R10494 gnd.n3591 gnd.n3582 585
R10495 gnd.n5351 gnd.n5350 585
R10496 gnd.n5352 gnd.n5351 585
R10497 gnd.n5343 gnd.n3590 585
R10498 gnd.n3594 gnd.n3590 585
R10499 gnd.n5342 gnd.n5341 585
R10500 gnd.n5341 gnd.n5340 585
R10501 gnd.n3593 gnd.n3592 585
R10502 gnd.n3603 gnd.n3593 585
R10503 gnd.n5319 gnd.n3601 585
R10504 gnd.n5334 gnd.n3601 585
R10505 gnd.n5320 gnd.n3615 585
R10506 gnd.n3615 gnd.n3614 585
R10507 gnd.n5322 gnd.n5321 585
R10508 gnd.n5323 gnd.n5322 585
R10509 gnd.n5318 gnd.n3613 585
R10510 gnd.n3613 gnd.n3610 585
R10511 gnd.n5317 gnd.n5316 585
R10512 gnd.n5316 gnd.n5315 585
R10513 gnd.n3617 gnd.n3616 585
R10514 gnd.n5306 gnd.n3617 585
R10515 gnd.n5305 gnd.n5304 585
R10516 gnd.n5307 gnd.n5305 585
R10517 gnd.n5303 gnd.n3626 585
R10518 gnd.n3630 gnd.n3626 585
R10519 gnd.n5302 gnd.n5301 585
R10520 gnd.n5301 gnd.n5300 585
R10521 gnd.n3628 gnd.n3627 585
R10522 gnd.n3629 gnd.n3628 585
R10523 gnd.n5262 gnd.n3635 585
R10524 gnd.n5294 gnd.n3635 585
R10525 gnd.n5264 gnd.n5263 585
R10526 gnd.n5263 gnd.n3646 585
R10527 gnd.n5265 gnd.n3645 585
R10528 gnd.n5276 gnd.n3645 585
R10529 gnd.n5267 gnd.n5266 585
R10530 gnd.n5268 gnd.n5267 585
R10531 gnd.n5261 gnd.n3651 585
R10532 gnd.n5270 gnd.n3651 585
R10533 gnd.n5260 gnd.n5259 585
R10534 gnd.n5259 gnd.n3650 585
R10535 gnd.n5258 gnd.n3653 585
R10536 gnd.n5258 gnd.n5257 585
R10537 gnd.n5234 gnd.n3654 585
R10538 gnd.n5250 gnd.n3654 585
R10539 gnd.n5235 gnd.n3661 585
R10540 gnd.n5251 gnd.n3661 585
R10541 gnd.n5237 gnd.n5236 585
R10542 gnd.n5238 gnd.n5237 585
R10543 gnd.n5233 gnd.n3670 585
R10544 gnd.n3675 gnd.n3670 585
R10545 gnd.n5232 gnd.n5231 585
R10546 gnd.n5231 gnd.n5230 585
R10547 gnd.n3672 gnd.n3671 585
R10548 gnd.n3682 gnd.n3672 585
R10549 gnd.n5199 gnd.n3680 585
R10550 gnd.n5223 gnd.n3680 585
R10551 gnd.n5202 gnd.n5201 585
R10552 gnd.n5201 gnd.n5200 585
R10553 gnd.n5203 gnd.n3690 585
R10554 gnd.n5213 gnd.n3690 585
R10555 gnd.n5204 gnd.n3699 585
R10556 gnd.n3699 gnd.n3688 585
R10557 gnd.n5206 gnd.n5205 585
R10558 gnd.n5207 gnd.n5206 585
R10559 gnd.n5198 gnd.n3698 585
R10560 gnd.n3698 gnd.n3695 585
R10561 gnd.n5197 gnd.n5196 585
R10562 gnd.n5196 gnd.n5195 585
R10563 gnd.n3701 gnd.n3700 585
R10564 gnd.n5188 gnd.n3701 585
R10565 gnd.n5187 gnd.n5186 585
R10566 gnd.n5189 gnd.n5187 585
R10567 gnd.n5185 gnd.n3708 585
R10568 gnd.n3712 gnd.n3708 585
R10569 gnd.n5184 gnd.n5183 585
R10570 gnd.n5183 gnd.n5182 585
R10571 gnd.n3710 gnd.n3709 585
R10572 gnd.n3711 gnd.n3710 585
R10573 gnd.n5140 gnd.n3719 585
R10574 gnd.n5176 gnd.n3719 585
R10575 gnd.n5142 gnd.n5141 585
R10576 gnd.n5141 gnd.n3729 585
R10577 gnd.n5143 gnd.n3728 585
R10578 gnd.n5155 gnd.n3728 585
R10579 gnd.n5145 gnd.n5144 585
R10580 gnd.n5146 gnd.n5145 585
R10581 gnd.n5139 gnd.n3734 585
R10582 gnd.n5149 gnd.n3734 585
R10583 gnd.n5138 gnd.n5137 585
R10584 gnd.n5137 gnd.n3733 585
R10585 gnd.n5136 gnd.n3736 585
R10586 gnd.n5136 gnd.n5135 585
R10587 gnd.n5111 gnd.n3737 585
R10588 gnd.n5128 gnd.n3737 585
R10589 gnd.n5112 gnd.n3743 585
R10590 gnd.n5129 gnd.n3743 585
R10591 gnd.n5114 gnd.n5113 585
R10592 gnd.n5115 gnd.n5114 585
R10593 gnd.n5110 gnd.n3752 585
R10594 gnd.n3756 gnd.n3752 585
R10595 gnd.n5109 gnd.n5108 585
R10596 gnd.n5108 gnd.n5107 585
R10597 gnd.n3754 gnd.n3753 585
R10598 gnd.n3763 gnd.n3754 585
R10599 gnd.n5075 gnd.n3761 585
R10600 gnd.n5100 gnd.n3761 585
R10601 gnd.n5078 gnd.n5077 585
R10602 gnd.n5077 gnd.n5076 585
R10603 gnd.n5079 gnd.n3770 585
R10604 gnd.n5089 gnd.n3770 585
R10605 gnd.n5080 gnd.n3778 585
R10606 gnd.n3778 gnd.n3776 585
R10607 gnd.n5082 gnd.n5081 585
R10608 gnd.n5083 gnd.n5082 585
R10609 gnd.n5074 gnd.n3777 585
R10610 gnd.n3782 gnd.n3777 585
R10611 gnd.n5073 gnd.n5072 585
R10612 gnd.n5072 gnd.n5071 585
R10613 gnd.n3780 gnd.n3779 585
R10614 gnd.n5064 gnd.n3780 585
R10615 gnd.n5063 gnd.n5062 585
R10616 gnd.n5065 gnd.n5063 585
R10617 gnd.n5061 gnd.n3789 585
R10618 gnd.n3793 gnd.n3789 585
R10619 gnd.n5060 gnd.n5059 585
R10620 gnd.n5059 gnd.n5058 585
R10621 gnd.n3791 gnd.n3790 585
R10622 gnd.n3792 gnd.n3791 585
R10623 gnd.n5017 gnd.n3799 585
R10624 gnd.n5052 gnd.n3799 585
R10625 gnd.n5019 gnd.n5018 585
R10626 gnd.n5018 gnd.n3809 585
R10627 gnd.n5020 gnd.n3808 585
R10628 gnd.n5031 gnd.n3808 585
R10629 gnd.n5022 gnd.n5021 585
R10630 gnd.n5023 gnd.n5022 585
R10631 gnd.n5016 gnd.n3813 585
R10632 gnd.n5025 gnd.n3813 585
R10633 gnd.n5015 gnd.n5014 585
R10634 gnd.n5014 gnd.n5013 585
R10635 gnd.n3816 gnd.n3815 585
R10636 gnd.n5003 gnd.n3816 585
R10637 gnd.n4994 gnd.n3825 585
R10638 gnd.n3825 gnd.n3818 585
R10639 gnd.n4996 gnd.n4995 585
R10640 gnd.n4997 gnd.n4996 585
R10641 gnd.n4993 gnd.n3824 585
R10642 gnd.n3824 gnd.n2912 585
R10643 gnd.n4992 gnd.n4991 585
R10644 gnd.n4991 gnd.n4990 585
R10645 gnd.n3899 gnd.n3826 585
R10646 gnd.n4983 gnd.n3899 585
R10647 gnd.n3898 gnd.n3897 585
R10648 gnd.n3898 gnd.n2901 585
R10649 gnd.n3896 gnd.n2899 585
R10650 gnd.n6319 gnd.n2899 585
R10651 gnd.n3895 gnd.n2898 585
R10652 gnd.n6320 gnd.n2898 585
R10653 gnd.n3894 gnd.n3893 585
R10654 gnd.n3893 gnd.n3892 585
R10655 gnd.n6449 gnd.n2759 585
R10656 gnd.n4764 gnd.n2759 585
R10657 gnd.n6451 gnd.n6450 585
R10658 gnd.n6452 gnd.n6451 585
R10659 gnd.n2744 gnd.n2743 585
R10660 gnd.n4724 gnd.n2744 585
R10661 gnd.n6460 gnd.n6459 585
R10662 gnd.n6459 gnd.n6458 585
R10663 gnd.n6461 gnd.n2738 585
R10664 gnd.n4472 gnd.n2738 585
R10665 gnd.n6463 gnd.n6462 585
R10666 gnd.n6464 gnd.n6463 585
R10667 gnd.n2724 gnd.n2723 585
R10668 gnd.n4737 gnd.n2724 585
R10669 gnd.n6472 gnd.n6471 585
R10670 gnd.n6471 gnd.n6470 585
R10671 gnd.n6473 gnd.n2718 585
R10672 gnd.n4465 gnd.n2718 585
R10673 gnd.n6475 gnd.n6474 585
R10674 gnd.n6476 gnd.n6475 585
R10675 gnd.n2704 gnd.n2703 585
R10676 gnd.n4457 gnd.n2704 585
R10677 gnd.n6484 gnd.n6483 585
R10678 gnd.n6483 gnd.n6482 585
R10679 gnd.n6485 gnd.n2698 585
R10680 gnd.n4419 gnd.n2698 585
R10681 gnd.n6487 gnd.n6486 585
R10682 gnd.n6488 gnd.n6487 585
R10683 gnd.n2684 gnd.n2683 585
R10684 gnd.n4410 gnd.n2684 585
R10685 gnd.n6496 gnd.n6495 585
R10686 gnd.n6495 gnd.n6494 585
R10687 gnd.n6497 gnd.n2678 585
R10688 gnd.n4405 gnd.n2678 585
R10689 gnd.n6499 gnd.n6498 585
R10690 gnd.n6500 gnd.n6499 585
R10691 gnd.n2664 gnd.n2663 585
R10692 gnd.n4433 gnd.n2664 585
R10693 gnd.n6508 gnd.n6507 585
R10694 gnd.n6507 gnd.n6506 585
R10695 gnd.n6509 gnd.n2658 585
R10696 gnd.n4398 gnd.n2658 585
R10697 gnd.n6511 gnd.n6510 585
R10698 gnd.n6512 gnd.n6511 585
R10699 gnd.n2644 gnd.n2643 585
R10700 gnd.n4390 gnd.n2644 585
R10701 gnd.n6520 gnd.n6519 585
R10702 gnd.n6519 gnd.n6518 585
R10703 gnd.n6521 gnd.n2639 585
R10704 gnd.n4384 gnd.n2639 585
R10705 gnd.n6523 gnd.n6522 585
R10706 gnd.n6524 gnd.n6523 585
R10707 gnd.n2623 gnd.n2621 585
R10708 gnd.n4376 gnd.n2623 585
R10709 gnd.n6532 gnd.n6531 585
R10710 gnd.n6531 gnd.n6530 585
R10711 gnd.n2622 gnd.n2620 585
R10712 gnd.n4345 gnd.n2622 585
R10713 gnd.n4334 gnd.n4333 585
R10714 gnd.n4333 gnd.n4016 585
R10715 gnd.n4336 gnd.n4335 585
R10716 gnd.n4337 gnd.n4336 585
R10717 gnd.n4332 gnd.n4029 585
R10718 gnd.n4332 gnd.n4331 585
R10719 gnd.n4028 gnd.n4027 585
R10720 gnd.n4315 gnd.n4027 585
R10721 gnd.n4265 gnd.n4264 585
R10722 gnd.n4266 gnd.n4265 585
R10723 gnd.n2614 gnd.n2612 585
R10724 gnd.n4307 gnd.n2612 585
R10725 gnd.n6536 gnd.n6535 585
R10726 gnd.n6537 gnd.n6536 585
R10727 gnd.n2613 gnd.n2597 585
R10728 gnd.n4275 gnd.n2597 585
R10729 gnd.n6545 gnd.n6544 585
R10730 gnd.n6544 gnd.n6543 585
R10731 gnd.n6546 gnd.n2592 585
R10732 gnd.n4281 gnd.n2592 585
R10733 gnd.n6548 gnd.n6547 585
R10734 gnd.n6549 gnd.n6548 585
R10735 gnd.n2579 gnd.n2578 585
R10736 gnd.n4257 gnd.n2579 585
R10737 gnd.n6557 gnd.n6556 585
R10738 gnd.n6556 gnd.n6555 585
R10739 gnd.n6558 gnd.n2573 585
R10740 gnd.n4248 gnd.n2573 585
R10741 gnd.n6560 gnd.n6559 585
R10742 gnd.n6561 gnd.n6560 585
R10743 gnd.n2558 gnd.n2557 585
R10744 gnd.n4211 gnd.n2558 585
R10745 gnd.n6569 gnd.n6568 585
R10746 gnd.n6568 gnd.n6567 585
R10747 gnd.n6570 gnd.n2552 585
R10748 gnd.n4217 gnd.n2552 585
R10749 gnd.n6572 gnd.n6571 585
R10750 gnd.n6573 gnd.n6572 585
R10751 gnd.n2539 gnd.n2538 585
R10752 gnd.n4199 gnd.n2539 585
R10753 gnd.n6581 gnd.n6580 585
R10754 gnd.n6580 gnd.n6579 585
R10755 gnd.n6582 gnd.n2533 585
R10756 gnd.n2533 gnd.n2532 585
R10757 gnd.n6584 gnd.n6583 585
R10758 gnd.n6585 gnd.n6584 585
R10759 gnd.n2518 gnd.n2517 585
R10760 gnd.n2522 gnd.n2518 585
R10761 gnd.n6593 gnd.n6592 585
R10762 gnd.n6592 gnd.n6591 585
R10763 gnd.n6594 gnd.n2512 585
R10764 gnd.n2519 gnd.n2512 585
R10765 gnd.n6596 gnd.n6595 585
R10766 gnd.n6597 gnd.n6596 585
R10767 gnd.n2500 gnd.n2499 585
R10768 gnd.n2503 gnd.n2500 585
R10769 gnd.n6605 gnd.n6604 585
R10770 gnd.n6604 gnd.n6603 585
R10771 gnd.n6606 gnd.n2494 585
R10772 gnd.n2494 gnd.n2493 585
R10773 gnd.n6608 gnd.n6607 585
R10774 gnd.n6609 gnd.n6608 585
R10775 gnd.n2477 gnd.n2476 585
R10776 gnd.n2481 gnd.n2477 585
R10777 gnd.n6617 gnd.n6616 585
R10778 gnd.n6616 gnd.n6615 585
R10779 gnd.n6618 gnd.n2470 585
R10780 gnd.n2478 gnd.n2470 585
R10781 gnd.n6620 gnd.n6619 585
R10782 gnd.n6621 gnd.n6620 585
R10783 gnd.n2471 gnd.n2397 585
R10784 gnd.n2397 gnd.n2394 585
R10785 gnd.n6743 gnd.n6742 585
R10786 gnd.n6741 gnd.n2396 585
R10787 gnd.n6740 gnd.n2395 585
R10788 gnd.n6745 gnd.n2395 585
R10789 gnd.n6739 gnd.n6738 585
R10790 gnd.n6737 gnd.n6736 585
R10791 gnd.n6735 gnd.n6734 585
R10792 gnd.n6733 gnd.n6732 585
R10793 gnd.n6731 gnd.n6730 585
R10794 gnd.n6729 gnd.n6728 585
R10795 gnd.n6727 gnd.n6726 585
R10796 gnd.n6725 gnd.n6724 585
R10797 gnd.n6723 gnd.n6722 585
R10798 gnd.n6721 gnd.n6720 585
R10799 gnd.n6719 gnd.n6718 585
R10800 gnd.n6717 gnd.n6716 585
R10801 gnd.n6715 gnd.n6714 585
R10802 gnd.n6713 gnd.n6712 585
R10803 gnd.n6711 gnd.n6710 585
R10804 gnd.n6708 gnd.n6707 585
R10805 gnd.n6706 gnd.n6705 585
R10806 gnd.n6704 gnd.n6703 585
R10807 gnd.n6702 gnd.n6701 585
R10808 gnd.n6700 gnd.n6699 585
R10809 gnd.n6698 gnd.n6697 585
R10810 gnd.n6696 gnd.n6695 585
R10811 gnd.n6694 gnd.n6693 585
R10812 gnd.n6692 gnd.n6691 585
R10813 gnd.n6690 gnd.n6689 585
R10814 gnd.n6688 gnd.n6687 585
R10815 gnd.n6686 gnd.n6685 585
R10816 gnd.n6684 gnd.n6683 585
R10817 gnd.n6682 gnd.n6681 585
R10818 gnd.n6680 gnd.n6679 585
R10819 gnd.n6678 gnd.n6677 585
R10820 gnd.n6676 gnd.n6675 585
R10821 gnd.n6674 gnd.n6673 585
R10822 gnd.n6672 gnd.n6671 585
R10823 gnd.n6670 gnd.n6669 585
R10824 gnd.n6668 gnd.n6667 585
R10825 gnd.n6666 gnd.n6665 585
R10826 gnd.n6664 gnd.n6663 585
R10827 gnd.n6662 gnd.n6661 585
R10828 gnd.n6660 gnd.n6659 585
R10829 gnd.n6658 gnd.n6657 585
R10830 gnd.n6656 gnd.n6655 585
R10831 gnd.n6654 gnd.n6653 585
R10832 gnd.n6652 gnd.n6651 585
R10833 gnd.n6650 gnd.n6649 585
R10834 gnd.n6648 gnd.n6647 585
R10835 gnd.n6646 gnd.n6645 585
R10836 gnd.n6644 gnd.n6643 585
R10837 gnd.n6642 gnd.n6641 585
R10838 gnd.n6640 gnd.n6639 585
R10839 gnd.n6638 gnd.n6637 585
R10840 gnd.n6636 gnd.n6635 585
R10841 gnd.n6634 gnd.n6633 585
R10842 gnd.n6632 gnd.n6631 585
R10843 gnd.n6630 gnd.n6629 585
R10844 gnd.n2466 gnd.n2459 585
R10845 gnd.n4716 gnd.n4715 585
R10846 gnd.n4714 gnd.n4625 585
R10847 gnd.n4713 gnd.n4712 585
R10848 gnd.n4706 gnd.n4626 585
R10849 gnd.n4708 gnd.n4707 585
R10850 gnd.n4705 gnd.n4704 585
R10851 gnd.n4703 gnd.n4702 585
R10852 gnd.n4696 gnd.n4628 585
R10853 gnd.n4698 gnd.n4697 585
R10854 gnd.n4695 gnd.n4694 585
R10855 gnd.n4693 gnd.n4692 585
R10856 gnd.n4686 gnd.n4630 585
R10857 gnd.n4688 gnd.n4687 585
R10858 gnd.n4685 gnd.n4684 585
R10859 gnd.n4683 gnd.n4682 585
R10860 gnd.n4676 gnd.n4632 585
R10861 gnd.n4678 gnd.n4677 585
R10862 gnd.n4675 gnd.n4674 585
R10863 gnd.n4673 gnd.n4672 585
R10864 gnd.n4666 gnd.n4634 585
R10865 gnd.n4668 gnd.n4667 585
R10866 gnd.n4665 gnd.n4638 585
R10867 gnd.n4664 gnd.n4663 585
R10868 gnd.n4657 gnd.n4639 585
R10869 gnd.n4659 gnd.n4658 585
R10870 gnd.n4656 gnd.n4655 585
R10871 gnd.n4654 gnd.n4653 585
R10872 gnd.n4647 gnd.n4641 585
R10873 gnd.n4649 gnd.n4648 585
R10874 gnd.n4646 gnd.n4645 585
R10875 gnd.n4644 gnd.n2832 585
R10876 gnd.n6396 gnd.n6395 585
R10877 gnd.n6398 gnd.n6397 585
R10878 gnd.n6400 gnd.n6399 585
R10879 gnd.n6402 gnd.n6401 585
R10880 gnd.n6404 gnd.n6403 585
R10881 gnd.n6406 gnd.n6405 585
R10882 gnd.n6408 gnd.n6407 585
R10883 gnd.n6410 gnd.n6409 585
R10884 gnd.n6413 gnd.n6412 585
R10885 gnd.n6415 gnd.n6414 585
R10886 gnd.n6417 gnd.n6416 585
R10887 gnd.n6419 gnd.n6418 585
R10888 gnd.n6421 gnd.n6420 585
R10889 gnd.n6423 gnd.n6422 585
R10890 gnd.n6425 gnd.n6424 585
R10891 gnd.n6427 gnd.n6426 585
R10892 gnd.n6429 gnd.n6428 585
R10893 gnd.n6431 gnd.n6430 585
R10894 gnd.n6433 gnd.n6432 585
R10895 gnd.n6435 gnd.n6434 585
R10896 gnd.n6437 gnd.n6436 585
R10897 gnd.n6439 gnd.n6438 585
R10898 gnd.n6440 gnd.n2805 585
R10899 gnd.n6442 gnd.n6441 585
R10900 gnd.n2764 gnd.n2763 585
R10901 gnd.n6446 gnd.n6445 585
R10902 gnd.n6445 gnd.n6444 585
R10903 gnd.n4720 gnd.n3957 585
R10904 gnd.n4764 gnd.n3957 585
R10905 gnd.n4721 gnd.n2756 585
R10906 gnd.n6452 gnd.n2756 585
R10907 gnd.n4723 gnd.n4722 585
R10908 gnd.n4724 gnd.n4723 585
R10909 gnd.n4475 gnd.n2746 585
R10910 gnd.n6458 gnd.n2746 585
R10911 gnd.n4474 gnd.n4473 585
R10912 gnd.n4473 gnd.n4472 585
R10913 gnd.n4470 gnd.n2735 585
R10914 gnd.n6464 gnd.n2735 585
R10915 gnd.n4469 gnd.n3968 585
R10916 gnd.n4737 gnd.n3968 585
R10917 gnd.n4468 gnd.n2726 585
R10918 gnd.n6470 gnd.n2726 585
R10919 gnd.n4467 gnd.n4466 585
R10920 gnd.n4466 gnd.n4465 585
R10921 gnd.n3974 gnd.n2715 585
R10922 gnd.n6476 gnd.n2715 585
R10923 gnd.n4415 gnd.n3979 585
R10924 gnd.n4457 gnd.n3979 585
R10925 gnd.n4416 gnd.n2706 585
R10926 gnd.n6482 gnd.n2706 585
R10927 gnd.n4418 gnd.n4417 585
R10928 gnd.n4419 gnd.n4418 585
R10929 gnd.n4413 gnd.n2695 585
R10930 gnd.n6488 gnd.n2695 585
R10931 gnd.n4412 gnd.n4411 585
R10932 gnd.n4411 gnd.n4410 585
R10933 gnd.n4408 gnd.n2686 585
R10934 gnd.n6494 gnd.n2686 585
R10935 gnd.n4407 gnd.n4406 585
R10936 gnd.n4406 gnd.n4405 585
R10937 gnd.n4403 gnd.n2675 585
R10938 gnd.n6500 gnd.n2675 585
R10939 gnd.n4402 gnd.n3991 585
R10940 gnd.n4433 gnd.n3991 585
R10941 gnd.n4401 gnd.n2666 585
R10942 gnd.n6506 gnd.n2666 585
R10943 gnd.n4400 gnd.n4399 585
R10944 gnd.n4399 gnd.n4398 585
R10945 gnd.n3999 gnd.n2655 585
R10946 gnd.n6512 gnd.n2655 585
R10947 gnd.n4389 gnd.n4388 585
R10948 gnd.n4390 gnd.n4389 585
R10949 gnd.n4387 gnd.n2646 585
R10950 gnd.n6518 gnd.n2646 585
R10951 gnd.n4386 gnd.n4385 585
R10952 gnd.n4385 gnd.n4384 585
R10953 gnd.n4005 gnd.n2636 585
R10954 gnd.n6524 gnd.n2636 585
R10955 gnd.n4320 gnd.n4010 585
R10956 gnd.n4376 gnd.n4010 585
R10957 gnd.n4321 gnd.n2625 585
R10958 gnd.n6530 gnd.n2625 585
R10959 gnd.n4322 gnd.n4017 585
R10960 gnd.n4345 gnd.n4017 585
R10961 gnd.n4324 gnd.n4323 585
R10962 gnd.n4323 gnd.n4016 585
R10963 gnd.n4319 gnd.n4024 585
R10964 gnd.n4337 gnd.n4024 585
R10965 gnd.n4318 gnd.n4031 585
R10966 gnd.n4331 gnd.n4031 585
R10967 gnd.n4317 gnd.n4316 585
R10968 gnd.n4316 gnd.n4315 585
R10969 gnd.n4039 gnd.n4037 585
R10970 gnd.n4266 gnd.n4039 585
R10971 gnd.n4271 gnd.n4045 585
R10972 gnd.n4307 gnd.n4045 585
R10973 gnd.n4272 gnd.n2609 585
R10974 gnd.n6537 gnd.n2609 585
R10975 gnd.n4274 gnd.n4273 585
R10976 gnd.n4275 gnd.n4274 585
R10977 gnd.n4263 gnd.n2599 585
R10978 gnd.n6543 gnd.n2599 585
R10979 gnd.n4262 gnd.n4054 585
R10980 gnd.n4281 gnd.n4054 585
R10981 gnd.n4260 gnd.n2590 585
R10982 gnd.n6549 gnd.n2590 585
R10983 gnd.n4259 gnd.n4258 585
R10984 gnd.n4258 gnd.n4257 585
R10985 gnd.n4059 gnd.n2580 585
R10986 gnd.n6555 gnd.n2580 585
R10987 gnd.n4207 gnd.n4063 585
R10988 gnd.n4248 gnd.n4063 585
R10989 gnd.n4208 gnd.n2570 585
R10990 gnd.n6561 gnd.n2570 585
R10991 gnd.n4210 gnd.n4209 585
R10992 gnd.n4211 gnd.n4210 585
R10993 gnd.n4205 gnd.n2560 585
R10994 gnd.n6567 gnd.n2560 585
R10995 gnd.n4204 gnd.n4068 585
R10996 gnd.n4217 gnd.n4068 585
R10997 gnd.n4202 gnd.n2550 585
R10998 gnd.n6573 gnd.n2550 585
R10999 gnd.n4201 gnd.n4200 585
R11000 gnd.n4200 gnd.n4199 585
R11001 gnd.n4096 gnd.n2540 585
R11002 gnd.n6579 gnd.n2540 585
R11003 gnd.n4095 gnd.n4094 585
R11004 gnd.n4094 gnd.n2532 585
R11005 gnd.n4092 gnd.n2530 585
R11006 gnd.n6585 gnd.n2530 585
R11007 gnd.n4091 gnd.n4090 585
R11008 gnd.n4090 gnd.n2522 585
R11009 gnd.n4089 gnd.n2520 585
R11010 gnd.n6591 gnd.n2520 585
R11011 gnd.n4088 gnd.n4087 585
R11012 gnd.n4087 gnd.n2519 585
R11013 gnd.n4085 gnd.n2510 585
R11014 gnd.n6597 gnd.n2510 585
R11015 gnd.n4084 gnd.n4083 585
R11016 gnd.n4083 gnd.n2503 585
R11017 gnd.n4082 gnd.n2501 585
R11018 gnd.n6603 gnd.n2501 585
R11019 gnd.n4081 gnd.n4080 585
R11020 gnd.n4080 gnd.n2493 585
R11021 gnd.n4078 gnd.n2491 585
R11022 gnd.n6609 gnd.n2491 585
R11023 gnd.n4077 gnd.n4076 585
R11024 gnd.n4076 gnd.n2481 585
R11025 gnd.n4075 gnd.n2479 585
R11026 gnd.n6615 gnd.n2479 585
R11027 gnd.n4074 gnd.n2467 585
R11028 gnd.n2478 gnd.n2467 585
R11029 gnd.n6622 gnd.n2465 585
R11030 gnd.n6622 gnd.n6621 585
R11031 gnd.n6624 gnd.n6623 585
R11032 gnd.n6623 gnd.n2394 585
R11033 gnd.n7978 gnd.n250 585
R11034 gnd.n250 gnd.n249 585
R11035 gnd.n7980 gnd.n7979 585
R11036 gnd.n7981 gnd.n7980 585
R11037 gnd.n237 gnd.n236 585
R11038 gnd.n240 gnd.n237 585
R11039 gnd.n7989 gnd.n7988 585
R11040 gnd.n7988 gnd.n7987 585
R11041 gnd.n7990 gnd.n231 585
R11042 gnd.n231 gnd.n230 585
R11043 gnd.n7992 gnd.n7991 585
R11044 gnd.n7993 gnd.n7992 585
R11045 gnd.n218 gnd.n217 585
R11046 gnd.n227 gnd.n218 585
R11047 gnd.n8001 gnd.n8000 585
R11048 gnd.n8000 gnd.n7999 585
R11049 gnd.n8002 gnd.n212 585
R11050 gnd.n212 gnd.n211 585
R11051 gnd.n8004 gnd.n8003 585
R11052 gnd.n8005 gnd.n8004 585
R11053 gnd.n198 gnd.n197 585
R11054 gnd.n202 gnd.n198 585
R11055 gnd.n8013 gnd.n8012 585
R11056 gnd.n8012 gnd.n8011 585
R11057 gnd.n8014 gnd.n192 585
R11058 gnd.n199 gnd.n192 585
R11059 gnd.n8016 gnd.n8015 585
R11060 gnd.n8017 gnd.n8016 585
R11061 gnd.n178 gnd.n177 585
R11062 gnd.n188 gnd.n178 585
R11063 gnd.n8025 gnd.n8024 585
R11064 gnd.n8024 gnd.n8023 585
R11065 gnd.n8026 gnd.n172 585
R11066 gnd.n7821 gnd.n172 585
R11067 gnd.n8028 gnd.n8027 585
R11068 gnd.n8029 gnd.n8028 585
R11069 gnd.n158 gnd.n157 585
R11070 gnd.n7716 gnd.n158 585
R11071 gnd.n8037 gnd.n8036 585
R11072 gnd.n8036 gnd.n8035 585
R11073 gnd.n8038 gnd.n152 585
R11074 gnd.n5872 gnd.n152 585
R11075 gnd.n8040 gnd.n8039 585
R11076 gnd.n8041 gnd.n8040 585
R11077 gnd.n138 gnd.n137 585
R11078 gnd.n5878 gnd.n138 585
R11079 gnd.n8049 gnd.n8048 585
R11080 gnd.n8048 gnd.n8047 585
R11081 gnd.n8050 gnd.n133 585
R11082 gnd.n5884 gnd.n133 585
R11083 gnd.n8052 gnd.n8051 585
R11084 gnd.n8053 gnd.n8052 585
R11085 gnd.n117 gnd.n115 585
R11086 gnd.n5890 gnd.n117 585
R11087 gnd.n8061 gnd.n8060 585
R11088 gnd.n8060 gnd.n8059 585
R11089 gnd.n116 gnd.n108 585
R11090 gnd.n5829 gnd.n116 585
R11091 gnd.n8064 gnd.n106 585
R11092 gnd.n5902 gnd.n106 585
R11093 gnd.n8066 gnd.n8065 585
R11094 gnd.n8067 gnd.n8066 585
R11095 gnd.n3348 gnd.n105 585
R11096 gnd.n5908 gnd.n105 585
R11097 gnd.n3350 gnd.n3349 585
R11098 gnd.n3362 gnd.n3350 585
R11099 gnd.n5916 gnd.n5915 585
R11100 gnd.n5915 gnd.n5914 585
R11101 gnd.n5918 gnd.n5917 585
R11102 gnd.n5919 gnd.n5918 585
R11103 gnd.n3347 gnd.n3346 585
R11104 gnd.n3347 gnd.n3340 585
R11105 gnd.n3345 gnd.n3330 585
R11106 gnd.n3333 gnd.n3330 585
R11107 gnd.n5930 gnd.n5929 585
R11108 gnd.n5929 gnd.n5928 585
R11109 gnd.n5932 gnd.n5931 585
R11110 gnd.n5933 gnd.n5932 585
R11111 gnd.n3315 gnd.n3314 585
R11112 gnd.n5788 gnd.n3315 585
R11113 gnd.n5941 gnd.n5940 585
R11114 gnd.n5940 gnd.n5939 585
R11115 gnd.n5942 gnd.n3308 585
R11116 gnd.n5768 gnd.n3308 585
R11117 gnd.n5944 gnd.n5943 585
R11118 gnd.n5945 gnd.n5944 585
R11119 gnd.n3294 gnd.n3293 585
R11120 gnd.n5761 gnd.n3294 585
R11121 gnd.n5953 gnd.n5952 585
R11122 gnd.n5952 gnd.n5951 585
R11123 gnd.n5954 gnd.n3288 585
R11124 gnd.n5753 gnd.n3288 585
R11125 gnd.n5956 gnd.n5955 585
R11126 gnd.n5957 gnd.n5956 585
R11127 gnd.n3273 gnd.n3272 585
R11128 gnd.n5746 gnd.n3273 585
R11129 gnd.n5965 gnd.n5964 585
R11130 gnd.n5964 gnd.n5963 585
R11131 gnd.n5966 gnd.n3267 585
R11132 gnd.n5738 gnd.n3267 585
R11133 gnd.n5968 gnd.n5967 585
R11134 gnd.n5969 gnd.n5968 585
R11135 gnd.n3253 gnd.n3252 585
R11136 gnd.n5731 gnd.n3253 585
R11137 gnd.n5977 gnd.n5976 585
R11138 gnd.n5976 gnd.n5975 585
R11139 gnd.n5978 gnd.n3247 585
R11140 gnd.n5723 gnd.n3247 585
R11141 gnd.n5980 gnd.n5979 585
R11142 gnd.n5981 gnd.n5980 585
R11143 gnd.n3232 gnd.n3231 585
R11144 gnd.n5716 gnd.n3232 585
R11145 gnd.n5989 gnd.n5988 585
R11146 gnd.n5988 gnd.n5987 585
R11147 gnd.n5990 gnd.n3226 585
R11148 gnd.n5708 gnd.n3226 585
R11149 gnd.n5992 gnd.n5991 585
R11150 gnd.n5993 gnd.n5992 585
R11151 gnd.n3208 gnd.n3207 585
R11152 gnd.n5701 gnd.n3208 585
R11153 gnd.n6001 gnd.n6000 585
R11154 gnd.n6000 gnd.n5999 585
R11155 gnd.n6002 gnd.n3199 585
R11156 gnd.n5693 gnd.n3199 585
R11157 gnd.n6004 gnd.n6003 585
R11158 gnd.n6005 gnd.n6004 585
R11159 gnd.n3200 gnd.n3198 585
R11160 gnd.n5669 gnd.n3198 585
R11161 gnd.n3201 gnd.n3120 585
R11162 gnd.n6013 gnd.n3120 585
R11163 gnd.n6132 gnd.n6131 585
R11164 gnd.n6130 gnd.n3119 585
R11165 gnd.n6129 gnd.n3118 585
R11166 gnd.n6134 gnd.n3118 585
R11167 gnd.n6128 gnd.n6127 585
R11168 gnd.n6126 gnd.n6125 585
R11169 gnd.n6124 gnd.n6123 585
R11170 gnd.n6122 gnd.n6121 585
R11171 gnd.n6120 gnd.n6119 585
R11172 gnd.n6118 gnd.n6117 585
R11173 gnd.n6116 gnd.n6115 585
R11174 gnd.n6114 gnd.n6113 585
R11175 gnd.n6112 gnd.n6111 585
R11176 gnd.n6110 gnd.n6109 585
R11177 gnd.n6108 gnd.n6107 585
R11178 gnd.n6106 gnd.n6105 585
R11179 gnd.n6104 gnd.n6103 585
R11180 gnd.n6102 gnd.n6101 585
R11181 gnd.n6100 gnd.n6099 585
R11182 gnd.n6097 gnd.n6096 585
R11183 gnd.n6095 gnd.n6094 585
R11184 gnd.n6093 gnd.n6092 585
R11185 gnd.n6091 gnd.n6090 585
R11186 gnd.n6089 gnd.n6088 585
R11187 gnd.n6087 gnd.n6086 585
R11188 gnd.n6085 gnd.n6084 585
R11189 gnd.n6083 gnd.n6082 585
R11190 gnd.n6080 gnd.n6079 585
R11191 gnd.n6078 gnd.n6077 585
R11192 gnd.n6076 gnd.n6075 585
R11193 gnd.n6074 gnd.n6073 585
R11194 gnd.n6072 gnd.n6071 585
R11195 gnd.n6070 gnd.n6069 585
R11196 gnd.n6068 gnd.n6067 585
R11197 gnd.n6066 gnd.n6065 585
R11198 gnd.n6064 gnd.n6063 585
R11199 gnd.n6062 gnd.n6061 585
R11200 gnd.n6060 gnd.n6059 585
R11201 gnd.n6058 gnd.n6057 585
R11202 gnd.n6056 gnd.n6055 585
R11203 gnd.n6054 gnd.n6053 585
R11204 gnd.n6052 gnd.n6051 585
R11205 gnd.n6050 gnd.n6049 585
R11206 gnd.n6048 gnd.n6047 585
R11207 gnd.n6046 gnd.n6045 585
R11208 gnd.n6044 gnd.n6043 585
R11209 gnd.n6042 gnd.n6041 585
R11210 gnd.n6040 gnd.n6039 585
R11211 gnd.n6038 gnd.n6037 585
R11212 gnd.n6036 gnd.n6035 585
R11213 gnd.n6034 gnd.n6033 585
R11214 gnd.n6032 gnd.n6031 585
R11215 gnd.n6030 gnd.n6029 585
R11216 gnd.n6028 gnd.n6027 585
R11217 gnd.n6026 gnd.n6025 585
R11218 gnd.n6024 gnd.n6023 585
R11219 gnd.n6022 gnd.n6021 585
R11220 gnd.n6016 gnd.n6015 585
R11221 gnd.n7849 gnd.n351 585
R11222 gnd.n7857 gnd.n7856 585
R11223 gnd.n7859 gnd.n7858 585
R11224 gnd.n7861 gnd.n7860 585
R11225 gnd.n7863 gnd.n7862 585
R11226 gnd.n7865 gnd.n7864 585
R11227 gnd.n7867 gnd.n7866 585
R11228 gnd.n7869 gnd.n7868 585
R11229 gnd.n7871 gnd.n7870 585
R11230 gnd.n7873 gnd.n7872 585
R11231 gnd.n7875 gnd.n7874 585
R11232 gnd.n7877 gnd.n7876 585
R11233 gnd.n7879 gnd.n7878 585
R11234 gnd.n7881 gnd.n7880 585
R11235 gnd.n7883 gnd.n7882 585
R11236 gnd.n7885 gnd.n7884 585
R11237 gnd.n7887 gnd.n7886 585
R11238 gnd.n7889 gnd.n7888 585
R11239 gnd.n7891 gnd.n7890 585
R11240 gnd.n7894 gnd.n7893 585
R11241 gnd.n7892 gnd.n331 585
R11242 gnd.n7899 gnd.n7898 585
R11243 gnd.n7901 gnd.n7900 585
R11244 gnd.n7903 gnd.n7902 585
R11245 gnd.n7905 gnd.n7904 585
R11246 gnd.n7907 gnd.n7906 585
R11247 gnd.n7909 gnd.n7908 585
R11248 gnd.n7911 gnd.n7910 585
R11249 gnd.n7913 gnd.n7912 585
R11250 gnd.n7915 gnd.n7914 585
R11251 gnd.n7917 gnd.n7916 585
R11252 gnd.n7919 gnd.n7918 585
R11253 gnd.n7921 gnd.n7920 585
R11254 gnd.n7923 gnd.n7922 585
R11255 gnd.n7925 gnd.n7924 585
R11256 gnd.n7927 gnd.n7926 585
R11257 gnd.n7929 gnd.n7928 585
R11258 gnd.n7931 gnd.n7930 585
R11259 gnd.n7933 gnd.n7932 585
R11260 gnd.n7935 gnd.n7934 585
R11261 gnd.n7937 gnd.n7936 585
R11262 gnd.n7942 gnd.n7941 585
R11263 gnd.n7944 gnd.n7943 585
R11264 gnd.n7946 gnd.n7945 585
R11265 gnd.n7948 gnd.n7947 585
R11266 gnd.n7950 gnd.n7949 585
R11267 gnd.n7952 gnd.n7951 585
R11268 gnd.n7954 gnd.n7953 585
R11269 gnd.n7956 gnd.n7955 585
R11270 gnd.n7958 gnd.n7957 585
R11271 gnd.n7960 gnd.n7959 585
R11272 gnd.n7962 gnd.n7961 585
R11273 gnd.n7964 gnd.n7963 585
R11274 gnd.n7966 gnd.n7965 585
R11275 gnd.n7968 gnd.n7967 585
R11276 gnd.n7969 gnd.n295 585
R11277 gnd.n7971 gnd.n7970 585
R11278 gnd.n255 gnd.n254 585
R11279 gnd.n7975 gnd.n7974 585
R11280 gnd.n7974 gnd.n7973 585
R11281 gnd.n7851 gnd.n7850 585
R11282 gnd.n7850 gnd.n249 585
R11283 gnd.n7848 gnd.n247 585
R11284 gnd.n7981 gnd.n247 585
R11285 gnd.n7847 gnd.n7846 585
R11286 gnd.n7846 gnd.n240 585
R11287 gnd.n7845 gnd.n238 585
R11288 gnd.n7987 gnd.n238 585
R11289 gnd.n7844 gnd.n7843 585
R11290 gnd.n7843 gnd.n230 585
R11291 gnd.n7841 gnd.n228 585
R11292 gnd.n7993 gnd.n228 585
R11293 gnd.n7840 gnd.n7839 585
R11294 gnd.n7839 gnd.n227 585
R11295 gnd.n7838 gnd.n219 585
R11296 gnd.n7999 gnd.n219 585
R11297 gnd.n7837 gnd.n7836 585
R11298 gnd.n7836 gnd.n211 585
R11299 gnd.n7834 gnd.n209 585
R11300 gnd.n8005 gnd.n209 585
R11301 gnd.n7833 gnd.n7832 585
R11302 gnd.n7832 gnd.n202 585
R11303 gnd.n7831 gnd.n200 585
R11304 gnd.n8011 gnd.n200 585
R11305 gnd.n7830 gnd.n7829 585
R11306 gnd.n7829 gnd.n199 585
R11307 gnd.n7827 gnd.n189 585
R11308 gnd.n8017 gnd.n189 585
R11309 gnd.n7826 gnd.n7825 585
R11310 gnd.n7825 gnd.n188 585
R11311 gnd.n7824 gnd.n180 585
R11312 gnd.n8023 gnd.n180 585
R11313 gnd.n7823 gnd.n7822 585
R11314 gnd.n7822 gnd.n7821 585
R11315 gnd.n355 gnd.n169 585
R11316 gnd.n8029 gnd.n169 585
R11317 gnd.n5868 gnd.n360 585
R11318 gnd.n7716 gnd.n360 585
R11319 gnd.n5869 gnd.n160 585
R11320 gnd.n8035 gnd.n160 585
R11321 gnd.n5871 gnd.n5870 585
R11322 gnd.n5872 gnd.n5871 585
R11323 gnd.n5842 gnd.n149 585
R11324 gnd.n8041 gnd.n149 585
R11325 gnd.n5880 gnd.n5879 585
R11326 gnd.n5879 gnd.n5878 585
R11327 gnd.n5881 gnd.n140 585
R11328 gnd.n8047 gnd.n140 585
R11329 gnd.n5883 gnd.n5882 585
R11330 gnd.n5884 gnd.n5883 585
R11331 gnd.n5840 gnd.n130 585
R11332 gnd.n8053 gnd.n130 585
R11333 gnd.n5839 gnd.n5826 585
R11334 gnd.n5890 gnd.n5826 585
R11335 gnd.n5838 gnd.n119 585
R11336 gnd.n8059 gnd.n119 585
R11337 gnd.n5810 gnd.n5809 585
R11338 gnd.n5829 gnd.n5810 585
R11339 gnd.n5904 gnd.n5903 585
R11340 gnd.n5903 gnd.n5902 585
R11341 gnd.n5905 gnd.n102 585
R11342 gnd.n8067 gnd.n102 585
R11343 gnd.n5907 gnd.n5906 585
R11344 gnd.n5908 gnd.n5907 585
R11345 gnd.n5805 gnd.n3363 585
R11346 gnd.n3363 gnd.n3362 585
R11347 gnd.n5804 gnd.n3351 585
R11348 gnd.n5914 gnd.n3351 585
R11349 gnd.n5803 gnd.n3341 585
R11350 gnd.n5919 gnd.n3341 585
R11351 gnd.n5793 gnd.n3364 585
R11352 gnd.n5793 gnd.n3340 585
R11353 gnd.n5795 gnd.n5794 585
R11354 gnd.n5794 gnd.n3333 585
R11355 gnd.n5792 gnd.n3331 585
R11356 gnd.n5928 gnd.n3331 585
R11357 gnd.n5791 gnd.n3327 585
R11358 gnd.n5933 gnd.n3327 585
R11359 gnd.n5790 gnd.n5789 585
R11360 gnd.n5789 gnd.n5788 585
R11361 gnd.n3366 gnd.n3317 585
R11362 gnd.n5939 gnd.n3317 585
R11363 gnd.n5767 gnd.n5766 585
R11364 gnd.n5768 gnd.n5767 585
R11365 gnd.n5764 gnd.n3305 585
R11366 gnd.n5945 gnd.n3305 585
R11367 gnd.n5763 gnd.n5762 585
R11368 gnd.n5762 gnd.n5761 585
R11369 gnd.n3371 gnd.n3296 585
R11370 gnd.n5951 gnd.n3296 585
R11371 gnd.n5752 gnd.n5751 585
R11372 gnd.n5753 gnd.n5752 585
R11373 gnd.n5749 gnd.n3285 585
R11374 gnd.n5957 gnd.n3285 585
R11375 gnd.n5748 gnd.n5747 585
R11376 gnd.n5747 gnd.n5746 585
R11377 gnd.n3376 gnd.n3275 585
R11378 gnd.n5963 gnd.n3275 585
R11379 gnd.n5737 gnd.n5736 585
R11380 gnd.n5738 gnd.n5737 585
R11381 gnd.n5734 gnd.n3264 585
R11382 gnd.n5969 gnd.n3264 585
R11383 gnd.n5733 gnd.n5732 585
R11384 gnd.n5732 gnd.n5731 585
R11385 gnd.n3380 gnd.n3255 585
R11386 gnd.n5975 gnd.n3255 585
R11387 gnd.n5722 gnd.n5721 585
R11388 gnd.n5723 gnd.n5722 585
R11389 gnd.n5719 gnd.n3244 585
R11390 gnd.n5981 gnd.n3244 585
R11391 gnd.n5718 gnd.n5717 585
R11392 gnd.n5717 gnd.n5716 585
R11393 gnd.n3385 gnd.n3234 585
R11394 gnd.n5987 gnd.n3234 585
R11395 gnd.n5707 gnd.n5706 585
R11396 gnd.n5708 gnd.n5707 585
R11397 gnd.n5704 gnd.n3223 585
R11398 gnd.n5993 gnd.n3223 585
R11399 gnd.n5703 gnd.n5702 585
R11400 gnd.n5702 gnd.n5701 585
R11401 gnd.n3389 gnd.n3210 585
R11402 gnd.n5999 gnd.n3210 585
R11403 gnd.n3194 gnd.n3193 585
R11404 gnd.n5693 gnd.n3194 585
R11405 gnd.n6007 gnd.n6006 585
R11406 gnd.n6006 gnd.n6005 585
R11407 gnd.n6008 gnd.n3183 585
R11408 gnd.n5669 gnd.n3183 585
R11409 gnd.n6014 gnd.n3184 585
R11410 gnd.n6014 gnd.n6013 585
R11411 gnd.n4225 gnd.n4223 585
R11412 gnd.n4223 gnd.n2529 585
R11413 gnd.n7707 gnd.n7706 585
R11414 gnd.n7707 gnd.n191 585
R11415 gnd.n7709 gnd.n367 585
R11416 gnd.n7709 gnd.n7708 585
R11417 gnd.n7711 gnd.n7710 585
R11418 gnd.n7710 gnd.n179 585
R11419 gnd.n7712 gnd.n362 585
R11420 gnd.n362 gnd.n171 585
R11421 gnd.n7714 gnd.n7713 585
R11422 gnd.n7715 gnd.n7714 585
R11423 gnd.n363 gnd.n361 585
R11424 gnd.n361 gnd.n162 585
R11425 gnd.n5856 gnd.n5855 585
R11426 gnd.n5856 gnd.n159 585
R11427 gnd.n5858 gnd.n5857 585
R11428 gnd.n5857 gnd.n151 585
R11429 gnd.n5859 gnd.n5844 585
R11430 gnd.n5844 gnd.n148 585
R11431 gnd.n5861 gnd.n5860 585
R11432 gnd.n5862 gnd.n5861 585
R11433 gnd.n5845 gnd.n5843 585
R11434 gnd.n5843 gnd.n139 585
R11435 gnd.n5847 gnd.n5825 585
R11436 gnd.n5825 gnd.n132 585
R11437 gnd.n5892 gnd.n5824 585
R11438 gnd.n5892 gnd.n5891 585
R11439 gnd.n5894 gnd.n5893 585
R11440 gnd.n5893 gnd.n121 585
R11441 gnd.n5895 gnd.n5812 585
R11442 gnd.n5812 gnd.n118 585
R11443 gnd.n5898 gnd.n5897 585
R11444 gnd.n5899 gnd.n5898 585
R11445 gnd.n5822 gnd.n5811 585
R11446 gnd.n5811 gnd.n103 585
R11447 gnd.n5820 gnd.n5819 585
R11448 gnd.n5819 gnd.n101 585
R11449 gnd.n5818 gnd.n5813 585
R11450 gnd.n5818 gnd.n3360 585
R11451 gnd.n5817 gnd.n5816 585
R11452 gnd.n5817 gnd.n3353 585
R11453 gnd.n5814 gnd.n3338 585
R11454 gnd.n3343 gnd.n3338 585
R11455 gnd.n5922 gnd.n5921 585
R11456 gnd.n5921 gnd.n5920 585
R11457 gnd.n5923 gnd.n3335 585
R11458 gnd.n3339 gnd.n3335 585
R11459 gnd.n5926 gnd.n5925 585
R11460 gnd.n5927 gnd.n5926 585
R11461 gnd.n3336 gnd.n3334 585
R11462 gnd.n3334 gnd.n3329 585
R11463 gnd.n5634 gnd.n5633 585
R11464 gnd.n5633 gnd.n3326 585
R11465 gnd.n5635 gnd.n5627 585
R11466 gnd.n5627 gnd.n3319 585
R11467 gnd.n5637 gnd.n5636 585
R11468 gnd.n5637 gnd.n3316 585
R11469 gnd.n5638 gnd.n5626 585
R11470 gnd.n5638 gnd.n3307 585
R11471 gnd.n5640 gnd.n5639 585
R11472 gnd.n5639 gnd.n3304 585
R11473 gnd.n5641 gnd.n5621 585
R11474 gnd.n5621 gnd.n3372 585
R11475 gnd.n5643 gnd.n5642 585
R11476 gnd.n5643 gnd.n3295 585
R11477 gnd.n5644 gnd.n5620 585
R11478 gnd.n5644 gnd.n3287 585
R11479 gnd.n5646 gnd.n5645 585
R11480 gnd.n5645 gnd.n3284 585
R11481 gnd.n5647 gnd.n5615 585
R11482 gnd.n5615 gnd.n3277 585
R11483 gnd.n5649 gnd.n5648 585
R11484 gnd.n5649 gnd.n3274 585
R11485 gnd.n5650 gnd.n5614 585
R11486 gnd.n5650 gnd.n3266 585
R11487 gnd.n5652 gnd.n5651 585
R11488 gnd.n5651 gnd.n3263 585
R11489 gnd.n5653 gnd.n5609 585
R11490 gnd.n5609 gnd.n3381 585
R11491 gnd.n5655 gnd.n5654 585
R11492 gnd.n5655 gnd.n3254 585
R11493 gnd.n5656 gnd.n5608 585
R11494 gnd.n5656 gnd.n3246 585
R11495 gnd.n5658 gnd.n5657 585
R11496 gnd.n5657 gnd.n3243 585
R11497 gnd.n5659 gnd.n5603 585
R11498 gnd.n5603 gnd.n3236 585
R11499 gnd.n5661 gnd.n5660 585
R11500 gnd.n5661 gnd.n3233 585
R11501 gnd.n5662 gnd.n5602 585
R11502 gnd.n5662 gnd.n3225 585
R11503 gnd.n5664 gnd.n5663 585
R11504 gnd.n5663 gnd.n3222 585
R11505 gnd.n5665 gnd.n5597 585
R11506 gnd.n5597 gnd.n3212 585
R11507 gnd.n5667 gnd.n5666 585
R11508 gnd.n5667 gnd.n3209 585
R11509 gnd.n5668 gnd.n5596 585
R11510 gnd.n5668 gnd.n3196 585
R11511 gnd.n5672 gnd.n5671 585
R11512 gnd.n5671 gnd.n5670 585
R11513 gnd.n5673 gnd.n5591 585
R11514 gnd.n5591 gnd.n3187 585
R11515 gnd.n5675 gnd.n5674 585
R11516 gnd.n5675 gnd.n3185 585
R11517 gnd.n5676 gnd.n5590 585
R11518 gnd.n5676 gnd.n3117 585
R11519 gnd.n5678 gnd.n5677 585
R11520 gnd.n5677 gnd.n3075 585
R11521 gnd.n5679 gnd.n3422 585
R11522 gnd.n3422 gnd.n3420 585
R11523 gnd.n5681 gnd.n5680 585
R11524 gnd.n5682 gnd.n5681 585
R11525 gnd.n3423 gnd.n3421 585
R11526 gnd.n3421 gnd.n3008 585
R11527 gnd.n5584 gnd.n3007 585
R11528 gnd.n6202 gnd.n3007 585
R11529 gnd.n5583 gnd.n5582 585
R11530 gnd.n5582 gnd.n3006 585
R11531 gnd.n5581 gnd.n3425 585
R11532 gnd.n5581 gnd.n5580 585
R11533 gnd.n5569 gnd.n3426 585
R11534 gnd.n3427 gnd.n3426 585
R11535 gnd.n5571 gnd.n5570 585
R11536 gnd.n5572 gnd.n5571 585
R11537 gnd.n3436 gnd.n3435 585
R11538 gnd.n3435 gnd.n3434 585
R11539 gnd.n5563 gnd.n5562 585
R11540 gnd.n5562 gnd.n5561 585
R11541 gnd.n3439 gnd.n3438 585
R11542 gnd.n3446 gnd.n3439 585
R11543 gnd.n5552 gnd.n5551 585
R11544 gnd.n5553 gnd.n5552 585
R11545 gnd.n3449 gnd.n3448 585
R11546 gnd.n3456 gnd.n3448 585
R11547 gnd.n5547 gnd.n5546 585
R11548 gnd.n5546 gnd.n5545 585
R11549 gnd.n3452 gnd.n3451 585
R11550 gnd.n5414 gnd.n3452 585
R11551 gnd.n5402 gnd.n3548 585
R11552 gnd.n3564 gnd.n3548 585
R11553 gnd.n5404 gnd.n5403 585
R11554 gnd.n5405 gnd.n5404 585
R11555 gnd.n3549 gnd.n3547 585
R11556 gnd.n3556 gnd.n3547 585
R11557 gnd.n5397 gnd.n5396 585
R11558 gnd.n5396 gnd.n5395 585
R11559 gnd.n3552 gnd.n3551 585
R11560 gnd.n3568 gnd.n3552 585
R11561 gnd.n5365 gnd.n5364 585
R11562 gnd.n5366 gnd.n5365 585
R11563 gnd.n3578 gnd.n3577 585
R11564 gnd.n3585 gnd.n3577 585
R11565 gnd.n5360 gnd.n5359 585
R11566 gnd.n5359 gnd.t365 585
R11567 gnd.n3581 gnd.n3580 585
R11568 gnd.n3589 gnd.n3581 585
R11569 gnd.n5330 gnd.n3605 585
R11570 gnd.n3605 gnd.n3596 585
R11571 gnd.n5332 gnd.n5331 585
R11572 gnd.n5333 gnd.n5332 585
R11573 gnd.n3606 gnd.n3604 585
R11574 gnd.n3604 gnd.n3600 585
R11575 gnd.n5325 gnd.n5324 585
R11576 gnd.n5324 gnd.n5323 585
R11577 gnd.n3609 gnd.n3608 585
R11578 gnd.n3620 gnd.n3609 585
R11579 gnd.n5287 gnd.n5286 585
R11580 gnd.n5287 gnd.n3618 585
R11581 gnd.n5289 gnd.n5288 585
R11582 gnd.n5288 gnd.n3625 585
R11583 gnd.n5290 gnd.n3639 585
R11584 gnd.n3639 gnd.n3631 585
R11585 gnd.n5292 gnd.n5291 585
R11586 gnd.n5293 gnd.n5292 585
R11587 gnd.n3640 gnd.n3638 585
R11588 gnd.n4876 gnd.n3638 585
R11589 gnd.n5279 gnd.n5278 585
R11590 gnd.n5278 gnd.n5277 585
R11591 gnd.n3643 gnd.n3642 585
R11592 gnd.n5269 gnd.n3643 585
R11593 gnd.n5246 gnd.n3664 585
R11594 gnd.n3664 gnd.n3656 585
R11595 gnd.n5248 gnd.n5247 585
R11596 gnd.n5249 gnd.n5248 585
R11597 gnd.n3665 gnd.n3663 585
R11598 gnd.n3663 gnd.n3660 585
R11599 gnd.n5241 gnd.n5240 585
R11600 gnd.n5240 gnd.n5239 585
R11601 gnd.n3668 gnd.n3667 585
R11602 gnd.n3674 gnd.n3668 585
R11603 gnd.n5221 gnd.n5220 585
R11604 gnd.n5222 gnd.n5221 585
R11605 gnd.n3684 gnd.n3683 585
R11606 gnd.n3691 gnd.n3683 585
R11607 gnd.n5216 gnd.n5215 585
R11608 gnd.n5215 gnd.n5214 585
R11609 gnd.n3687 gnd.n3686 585
R11610 gnd.n5207 gnd.n3687 585
R11611 gnd.n5168 gnd.n5167 585
R11612 gnd.n5168 gnd.n3703 585
R11613 gnd.n5169 gnd.n5164 585
R11614 gnd.n5169 gnd.n3702 585
R11615 gnd.n5171 gnd.n5170 585
R11616 gnd.n5170 gnd.n3707 585
R11617 gnd.n5172 gnd.n3722 585
R11618 gnd.n3722 gnd.n3714 585
R11619 gnd.n5174 gnd.n5173 585
R11620 gnd.n5175 gnd.n5174 585
R11621 gnd.n3723 gnd.n3721 585
R11622 gnd.n3721 gnd.n3718 585
R11623 gnd.n5158 gnd.n5157 585
R11624 gnd.n5157 gnd.n5156 585
R11625 gnd.n3726 gnd.n3725 585
R11626 gnd.n5148 gnd.n3726 585
R11627 gnd.n5124 gnd.n3746 585
R11628 gnd.n3746 gnd.n3738 585
R11629 gnd.n5126 gnd.n5125 585
R11630 gnd.n5127 gnd.n5126 585
R11631 gnd.n3747 gnd.n3745 585
R11632 gnd.n3745 gnd.n3742 585
R11633 gnd.n5119 gnd.n5118 585
R11634 gnd.n5118 gnd.n5117 585
R11635 gnd.n3750 gnd.n3749 585
R11636 gnd.n3755 gnd.n3750 585
R11637 gnd.n5098 gnd.n5097 585
R11638 gnd.n5099 gnd.n5098 585
R11639 gnd.n3765 gnd.n3764 585
R11640 gnd.n3771 gnd.n3764 585
R11641 gnd.n5093 gnd.n5092 585
R11642 gnd.n5092 gnd.n5091 585
R11643 gnd.n3768 gnd.n3767 585
R11644 gnd.n5083 gnd.n3768 585
R11645 gnd.n5045 gnd.n5044 585
R11646 gnd.n5045 gnd.n3783 585
R11647 gnd.n5046 gnd.n5041 585
R11648 gnd.n5046 gnd.n3781 585
R11649 gnd.n5048 gnd.n5047 585
R11650 gnd.n5047 gnd.n3788 585
R11651 gnd.n5049 gnd.n3802 585
R11652 gnd.n3802 gnd.n3794 585
R11653 gnd.n5051 gnd.n5050 585
R11654 gnd.t348 gnd.n5051 585
R11655 gnd.n3803 gnd.n3801 585
R11656 gnd.n3801 gnd.n3798 585
R11657 gnd.n5035 gnd.n5034 585
R11658 gnd.n5034 gnd.n5033 585
R11659 gnd.n3806 gnd.n3805 585
R11660 gnd.n5024 gnd.n3806 585
R11661 gnd.n5011 gnd.n5010 585
R11662 gnd.n5012 gnd.n5011 585
R11663 gnd.n5006 gnd.n5005 585
R11664 gnd.n5005 gnd.n5004 585
R11665 gnd.n2910 gnd.n2909 585
R11666 gnd.n3823 gnd.n2910 585
R11667 gnd.n6314 gnd.n6313 585
R11668 gnd.n6313 gnd.n6312 585
R11669 gnd.n6315 gnd.n2904 585
R11670 gnd.n4982 gnd.n2904 585
R11671 gnd.n6317 gnd.n6316 585
R11672 gnd.n6318 gnd.n6317 585
R11673 gnd.n2905 gnd.n2903 585
R11674 gnd.n2903 gnd.n2897 585
R11675 gnd.n4819 gnd.n4818 585
R11676 gnd.n4819 gnd.n2871 585
R11677 gnd.n4821 gnd.n4820 585
R11678 gnd.n4820 gnd.n2839 585
R11679 gnd.n4822 gnd.n3913 585
R11680 gnd.n3913 gnd.n3910 585
R11681 gnd.n4824 gnd.n4823 585
R11682 gnd.n4825 gnd.n4824 585
R11683 gnd.n3914 gnd.n3912 585
R11684 gnd.n3912 gnd.n3909 585
R11685 gnd.n4810 gnd.n4809 585
R11686 gnd.n4809 gnd.n4808 585
R11687 gnd.n3917 gnd.n3916 585
R11688 gnd.n3918 gnd.n3917 585
R11689 gnd.n4782 gnd.n4781 585
R11690 gnd.n4783 gnd.n4782 585
R11691 gnd.n3930 gnd.n3929 585
R11692 gnd.n3929 gnd.n3927 585
R11693 gnd.n4777 gnd.n4776 585
R11694 gnd.n4776 gnd.n4775 585
R11695 gnd.n3933 gnd.n3932 585
R11696 gnd.n4774 gnd.n3933 585
R11697 gnd.n4757 gnd.n4756 585
R11698 gnd.n4757 gnd.n3934 585
R11699 gnd.n4759 gnd.n4758 585
R11700 gnd.n4758 gnd.n2776 585
R11701 gnd.n4760 gnd.n3959 585
R11702 gnd.n3959 gnd.n2765 585
R11703 gnd.n4762 gnd.n4761 585
R11704 gnd.n4763 gnd.n4762 585
R11705 gnd.n3960 gnd.n3958 585
R11706 gnd.n3958 gnd.n2758 585
R11707 gnd.n4749 gnd.n4748 585
R11708 gnd.n4748 gnd.n2755 585
R11709 gnd.n4747 gnd.n3962 585
R11710 gnd.n4747 gnd.n2748 585
R11711 gnd.n4746 gnd.n4745 585
R11712 gnd.n4746 gnd.n2745 585
R11713 gnd.n3964 gnd.n3963 585
R11714 gnd.n3963 gnd.n2737 585
R11715 gnd.n4741 gnd.n4740 585
R11716 gnd.n4740 gnd.n2734 585
R11717 gnd.n4739 gnd.n3966 585
R11718 gnd.n4739 gnd.n4738 585
R11719 gnd.n4452 gnd.n3967 585
R11720 gnd.n3967 gnd.n2725 585
R11721 gnd.n4453 gnd.n3981 585
R11722 gnd.n3981 gnd.n2717 585
R11723 gnd.n4455 gnd.n4454 585
R11724 gnd.n4456 gnd.n4455 585
R11725 gnd.n3982 gnd.n3980 585
R11726 gnd.n3980 gnd.n2708 585
R11727 gnd.n4446 gnd.n4445 585
R11728 gnd.n4445 gnd.n2705 585
R11729 gnd.n4444 gnd.n3984 585
R11730 gnd.n4444 gnd.n2697 585
R11731 gnd.n4443 gnd.n4442 585
R11732 gnd.n4443 gnd.n2694 585
R11733 gnd.n3986 gnd.n3985 585
R11734 gnd.n4409 gnd.n3985 585
R11735 gnd.n4438 gnd.n4437 585
R11736 gnd.n4437 gnd.n2685 585
R11737 gnd.n4436 gnd.n3988 585
R11738 gnd.n4436 gnd.n2677 585
R11739 gnd.n4435 gnd.n3990 585
R11740 gnd.n4435 gnd.n4434 585
R11741 gnd.n4363 gnd.n3989 585
R11742 gnd.n3989 gnd.n2668 585
R11743 gnd.n4365 gnd.n4364 585
R11744 gnd.n4364 gnd.n2665 585
R11745 gnd.n4366 gnd.n4356 585
R11746 gnd.n4356 gnd.n2657 585
R11747 gnd.n4368 gnd.n4367 585
R11748 gnd.n4368 gnd.n2654 585
R11749 gnd.n4369 gnd.n4355 585
R11750 gnd.n4369 gnd.n4004 585
R11751 gnd.n4371 gnd.n4370 585
R11752 gnd.n4370 gnd.n2645 585
R11753 gnd.n4372 gnd.n4012 585
R11754 gnd.n4012 gnd.n2638 585
R11755 gnd.n4374 gnd.n4373 585
R11756 gnd.n4375 gnd.n4374 585
R11757 gnd.n4350 gnd.n4011 585
R11758 gnd.n4011 gnd.n2627 585
R11759 gnd.n4349 gnd.n4348 585
R11760 gnd.n4348 gnd.n2624 585
R11761 gnd.n4347 gnd.n4015 585
R11762 gnd.n4347 gnd.n4346 585
R11763 gnd.n4296 gnd.n4014 585
R11764 gnd.n4025 gnd.n4014 585
R11765 gnd.n4299 gnd.n4298 585
R11766 gnd.n4299 gnd.n4023 585
R11767 gnd.n4301 gnd.n4300 585
R11768 gnd.n4300 gnd.n4030 585
R11769 gnd.n4303 gnd.n4047 585
R11770 gnd.n4047 gnd.n4040 585
R11771 gnd.n4305 gnd.n4304 585
R11772 gnd.n4306 gnd.n4305 585
R11773 gnd.n4294 gnd.n4046 585
R11774 gnd.n4046 gnd.n2611 585
R11775 gnd.n4293 gnd.n4292 585
R11776 gnd.n4292 gnd.n2608 585
R11777 gnd.n4291 gnd.n4290 585
R11778 gnd.n4291 gnd.n2601 585
R11779 gnd.n4289 gnd.n4049 585
R11780 gnd.n4049 gnd.n2598 585
R11781 gnd.n4283 gnd.n4050 585
R11782 gnd.n4283 gnd.n4282 585
R11783 gnd.n4285 gnd.n4284 585
R11784 gnd.n4284 gnd.n2589 585
R11785 gnd.n4053 gnd.n4052 585
R11786 gnd.n4053 gnd.n2582 585
R11787 gnd.n4246 gnd.n4245 585
R11788 gnd.n4247 gnd.n4246 585
R11789 gnd.n4065 gnd.n4064 585
R11790 gnd.n4064 gnd.n2572 585
R11791 gnd.n4241 gnd.n4240 585
R11792 gnd.n4240 gnd.n2569 585
R11793 gnd.n4239 gnd.n4067 585
R11794 gnd.n4239 gnd.n2562 585
R11795 gnd.n4238 gnd.n4237 585
R11796 gnd.n4238 gnd.n2559 585
R11797 gnd.n4220 gnd.n4219 585
R11798 gnd.n4219 gnd.n4218 585
R11799 gnd.n4233 gnd.n4232 585
R11800 gnd.n4232 gnd.n2549 585
R11801 gnd.n4231 gnd.n4222 585
R11802 gnd.n4231 gnd.n2542 585
R11803 gnd.n4230 gnd.n4228 585
R11804 gnd.n4230 gnd.n4229 585
R11805 gnd.n6201 gnd.n6200 585
R11806 gnd.n6202 gnd.n6201 585
R11807 gnd.n3011 gnd.n3009 585
R11808 gnd.n3009 gnd.n3006 585
R11809 gnd.n5579 gnd.n5578 585
R11810 gnd.n5580 gnd.n5579 585
R11811 gnd.n3429 gnd.n3428 585
R11812 gnd.n3428 gnd.n3427 585
R11813 gnd.n5574 gnd.n5573 585
R11814 gnd.n5573 gnd.n5572 585
R11815 gnd.n3432 gnd.n3431 585
R11816 gnd.n3434 gnd.n3432 585
R11817 gnd.n5560 gnd.n5559 585
R11818 gnd.n5561 gnd.n5560 585
R11819 gnd.n3441 gnd.n3440 585
R11820 gnd.n3446 gnd.n3440 585
R11821 gnd.n5555 gnd.n5554 585
R11822 gnd.n5554 gnd.n5553 585
R11823 gnd.n3444 gnd.n3443 585
R11824 gnd.n3456 gnd.n3444 585
R11825 gnd.n3540 gnd.n3453 585
R11826 gnd.n5545 gnd.n3453 585
R11827 gnd.n5413 gnd.n5412 585
R11828 gnd.n5414 gnd.n5413 585
R11829 gnd.n3539 gnd.n3538 585
R11830 gnd.n3564 gnd.n3538 585
R11831 gnd.n5407 gnd.n5406 585
R11832 gnd.n5406 gnd.n5405 585
R11833 gnd.n3543 gnd.n3542 585
R11834 gnd.n3556 gnd.n3543 585
R11835 gnd.n4896 gnd.n3554 585
R11836 gnd.n5395 gnd.n3554 585
R11837 gnd.n4897 gnd.n4894 585
R11838 gnd.n4894 gnd.n3568 585
R11839 gnd.n4898 gnd.n3574 585
R11840 gnd.n5366 gnd.n3574 585
R11841 gnd.n4892 gnd.n4891 585
R11842 gnd.n4891 gnd.n3585 585
R11843 gnd.n4902 gnd.n3583 585
R11844 gnd.t365 gnd.n3583 585
R11845 gnd.n4903 gnd.n4890 585
R11846 gnd.n4890 gnd.n3589 585
R11847 gnd.n4904 gnd.n4889 585
R11848 gnd.n4889 gnd.n3596 585
R11849 gnd.n4887 gnd.n3602 585
R11850 gnd.n5333 gnd.n3602 585
R11851 gnd.n4908 gnd.n4886 585
R11852 gnd.n4886 gnd.n3600 585
R11853 gnd.n4909 gnd.n3612 585
R11854 gnd.n5323 gnd.n3612 585
R11855 gnd.n4910 gnd.n4885 585
R11856 gnd.n4885 gnd.n3620 585
R11857 gnd.n4884 gnd.n4882 585
R11858 gnd.n4884 gnd.n3618 585
R11859 gnd.n4914 gnd.n4881 585
R11860 gnd.n4881 gnd.n3625 585
R11861 gnd.n4915 gnd.n4880 585
R11862 gnd.n4880 gnd.n3631 585
R11863 gnd.n4916 gnd.n3636 585
R11864 gnd.n5293 gnd.n3636 585
R11865 gnd.n4878 gnd.n4877 585
R11866 gnd.n4877 gnd.n4876 585
R11867 gnd.n4920 gnd.n3644 585
R11868 gnd.n5277 gnd.n3644 585
R11869 gnd.n4921 gnd.n3652 585
R11870 gnd.n5269 gnd.n3652 585
R11871 gnd.n4922 gnd.n4875 585
R11872 gnd.n4875 gnd.n3656 585
R11873 gnd.n4873 gnd.n3662 585
R11874 gnd.n5249 gnd.n3662 585
R11875 gnd.n4926 gnd.n4872 585
R11876 gnd.n4872 gnd.n3660 585
R11877 gnd.n4927 gnd.n3669 585
R11878 gnd.n5239 gnd.n3669 585
R11879 gnd.n4928 gnd.n4871 585
R11880 gnd.n4871 gnd.n3674 585
R11881 gnd.n4869 gnd.n3681 585
R11882 gnd.n5222 gnd.n3681 585
R11883 gnd.n4932 gnd.n4868 585
R11884 gnd.n4868 gnd.n3691 585
R11885 gnd.n4933 gnd.n3689 585
R11886 gnd.n5214 gnd.n3689 585
R11887 gnd.n4934 gnd.n3696 585
R11888 gnd.n5207 gnd.n3696 585
R11889 gnd.n4866 gnd.n4865 585
R11890 gnd.n4865 gnd.n3703 585
R11891 gnd.n4938 gnd.n4864 585
R11892 gnd.n4864 gnd.n3702 585
R11893 gnd.n4939 gnd.n4863 585
R11894 gnd.n4863 gnd.n3707 585
R11895 gnd.n4940 gnd.n4862 585
R11896 gnd.n4862 gnd.n3714 585
R11897 gnd.n4860 gnd.n3720 585
R11898 gnd.n5175 gnd.n3720 585
R11899 gnd.n4944 gnd.n4859 585
R11900 gnd.n4859 gnd.n3718 585
R11901 gnd.n4945 gnd.n3727 585
R11902 gnd.n5156 gnd.n3727 585
R11903 gnd.n4946 gnd.n3735 585
R11904 gnd.n5148 gnd.n3735 585
R11905 gnd.n4857 gnd.n4856 585
R11906 gnd.n4856 gnd.n3738 585
R11907 gnd.n4950 gnd.n3744 585
R11908 gnd.n5127 gnd.n3744 585
R11909 gnd.n4951 gnd.n4855 585
R11910 gnd.n4855 gnd.n3742 585
R11911 gnd.n4952 gnd.n3751 585
R11912 gnd.n5117 gnd.n3751 585
R11913 gnd.n4853 gnd.n4852 585
R11914 gnd.n4852 gnd.n3755 585
R11915 gnd.n4956 gnd.n3762 585
R11916 gnd.n5099 gnd.n3762 585
R11917 gnd.n4957 gnd.n4851 585
R11918 gnd.n4851 gnd.n3771 585
R11919 gnd.n4958 gnd.n3769 585
R11920 gnd.n5091 gnd.n3769 585
R11921 gnd.n4849 gnd.n3775 585
R11922 gnd.n5083 gnd.n3775 585
R11923 gnd.n4962 gnd.n4848 585
R11924 gnd.n4848 gnd.n3783 585
R11925 gnd.n4963 gnd.n4847 585
R11926 gnd.n4847 gnd.n3781 585
R11927 gnd.n4964 gnd.n4846 585
R11928 gnd.n4846 gnd.n3788 585
R11929 gnd.n4845 gnd.n4843 585
R11930 gnd.n4845 gnd.n3794 585
R11931 gnd.n4968 gnd.n3800 585
R11932 gnd.t348 gnd.n3800 585
R11933 gnd.n4969 gnd.n4842 585
R11934 gnd.n4842 gnd.n3798 585
R11935 gnd.n4970 gnd.n3807 585
R11936 gnd.n5033 gnd.n3807 585
R11937 gnd.n4840 gnd.n3814 585
R11938 gnd.n5024 gnd.n3814 585
R11939 gnd.n4974 gnd.n3817 585
R11940 gnd.n5012 gnd.n3817 585
R11941 gnd.n4975 gnd.n3819 585
R11942 gnd.n5004 gnd.n3819 585
R11943 gnd.n4976 gnd.n4839 585
R11944 gnd.n4839 gnd.n3823 585
R11945 gnd.n3901 gnd.n2911 585
R11946 gnd.n6312 gnd.n2911 585
R11947 gnd.n4981 gnd.n4980 585
R11948 gnd.n4982 gnd.n4981 585
R11949 gnd.n3900 gnd.n2900 585
R11950 gnd.n6318 gnd.n2900 585
R11951 gnd.n4835 gnd.n4834 585
R11952 gnd.n4834 gnd.n2897 585
R11953 gnd.n4833 gnd.n3903 585
R11954 gnd.n4833 gnd.n2871 585
R11955 gnd.n4832 gnd.n4831 585
R11956 gnd.n4832 gnd.n2839 585
R11957 gnd.n3905 gnd.n3904 585
R11958 gnd.n3910 gnd.n3904 585
R11959 gnd.n4827 gnd.n4826 585
R11960 gnd.n4826 gnd.n4825 585
R11961 gnd.n3908 gnd.n3907 585
R11962 gnd.n3909 gnd.n3908 585
R11963 gnd.n4486 gnd.n3919 585
R11964 gnd.n4808 gnd.n3919 585
R11965 gnd.n4487 gnd.n4485 585
R11966 gnd.n4485 gnd.n3918 585
R11967 gnd.n4483 gnd.n3928 585
R11968 gnd.n4783 gnd.n3928 585
R11969 gnd.n4492 gnd.n4491 585
R11970 gnd.n4492 gnd.n3927 585
R11971 gnd.n4494 gnd.n4493 585
R11972 gnd.n4496 gnd.n4495 585
R11973 gnd.n4498 gnd.n4497 585
R11974 gnd.n4479 gnd.n4478 585
R11975 gnd.n4502 gnd.n4480 585
R11976 gnd.n4504 gnd.n4503 585
R11977 gnd.n4619 gnd.n4505 585
R11978 gnd.n4618 gnd.n4506 585
R11979 gnd.n4617 gnd.n4507 585
R11980 gnd.n4513 gnd.n4508 585
R11981 gnd.n4610 gnd.n4514 585
R11982 gnd.n4609 gnd.n4515 585
R11983 gnd.n4517 gnd.n4516 585
R11984 gnd.n4602 gnd.n4525 585
R11985 gnd.n4601 gnd.n4526 585
R11986 gnd.n4533 gnd.n4527 585
R11987 gnd.n4594 gnd.n4534 585
R11988 gnd.n4593 gnd.n4535 585
R11989 gnd.n4537 gnd.n4536 585
R11990 gnd.n4586 gnd.n4545 585
R11991 gnd.n4585 gnd.n4546 585
R11992 gnd.n4553 gnd.n4547 585
R11993 gnd.n4578 gnd.n4554 585
R11994 gnd.n4577 gnd.n4555 585
R11995 gnd.n4557 gnd.n4556 585
R11996 gnd.n4570 gnd.n4567 585
R11997 gnd.n4569 gnd.n4568 585
R11998 gnd.n3950 gnd.n3949 585
R11999 gnd.n4773 gnd.n4772 585
R12000 gnd.n4774 gnd.n4773 585
R12001 gnd.n6204 gnd.n6203 585
R12002 gnd.n6203 gnd.n6202 585
R12003 gnd.n3004 gnd.n3002 585
R12004 gnd.n3006 gnd.n3004 585
R12005 gnd.n6208 gnd.n3001 585
R12006 gnd.n5580 gnd.n3001 585
R12007 gnd.n6209 gnd.n3000 585
R12008 gnd.n3427 gnd.n3000 585
R12009 gnd.n6210 gnd.n2999 585
R12010 gnd.n5572 gnd.n2999 585
R12011 gnd.n3433 gnd.n2997 585
R12012 gnd.n3434 gnd.n3433 585
R12013 gnd.n6214 gnd.n2996 585
R12014 gnd.n5561 gnd.n2996 585
R12015 gnd.n6215 gnd.n2995 585
R12016 gnd.n3446 gnd.n2995 585
R12017 gnd.n6216 gnd.n2994 585
R12018 gnd.n5553 gnd.n2994 585
R12019 gnd.n3455 gnd.n2992 585
R12020 gnd.n3456 gnd.n3455 585
R12021 gnd.n6220 gnd.n2991 585
R12022 gnd.n5545 gnd.n2991 585
R12023 gnd.n6221 gnd.n2990 585
R12024 gnd.n5414 gnd.n2990 585
R12025 gnd.n6222 gnd.n2989 585
R12026 gnd.n3564 gnd.n2989 585
R12027 gnd.n3546 gnd.n2987 585
R12028 gnd.n5405 gnd.n3546 585
R12029 gnd.n6226 gnd.n2986 585
R12030 gnd.n3556 gnd.n2986 585
R12031 gnd.n6227 gnd.n2985 585
R12032 gnd.n5395 gnd.n2985 585
R12033 gnd.n6228 gnd.n2984 585
R12034 gnd.n3568 gnd.n2984 585
R12035 gnd.n3576 gnd.n2982 585
R12036 gnd.n5366 gnd.n3576 585
R12037 gnd.n6232 gnd.n2981 585
R12038 gnd.n3585 gnd.n2981 585
R12039 gnd.n6233 gnd.n2980 585
R12040 gnd.t365 gnd.n2980 585
R12041 gnd.n6234 gnd.n2979 585
R12042 gnd.n3589 gnd.n2979 585
R12043 gnd.n3595 gnd.n2977 585
R12044 gnd.n3596 gnd.n3595 585
R12045 gnd.n6238 gnd.n2976 585
R12046 gnd.n5333 gnd.n2976 585
R12047 gnd.n6239 gnd.n2975 585
R12048 gnd.n3600 gnd.n2975 585
R12049 gnd.n6240 gnd.n2974 585
R12050 gnd.n5323 gnd.n2974 585
R12051 gnd.n3619 gnd.n2972 585
R12052 gnd.n3620 gnd.n3619 585
R12053 gnd.n6244 gnd.n2971 585
R12054 gnd.n3618 gnd.n2971 585
R12055 gnd.n6245 gnd.n2970 585
R12056 gnd.n3625 gnd.n2970 585
R12057 gnd.n6246 gnd.n2969 585
R12058 gnd.n3631 gnd.n2969 585
R12059 gnd.n3637 gnd.n2967 585
R12060 gnd.n5293 gnd.n3637 585
R12061 gnd.n6250 gnd.n2966 585
R12062 gnd.n4876 gnd.n2966 585
R12063 gnd.n6251 gnd.n2965 585
R12064 gnd.n5277 gnd.n2965 585
R12065 gnd.n6252 gnd.n2964 585
R12066 gnd.n5269 gnd.n2964 585
R12067 gnd.n3655 gnd.n2962 585
R12068 gnd.n3656 gnd.n3655 585
R12069 gnd.n6256 gnd.n2961 585
R12070 gnd.n5249 gnd.n2961 585
R12071 gnd.n6257 gnd.n2960 585
R12072 gnd.n3660 gnd.n2960 585
R12073 gnd.n6258 gnd.n2959 585
R12074 gnd.n5239 gnd.n2959 585
R12075 gnd.n3673 gnd.n2957 585
R12076 gnd.n3674 gnd.n3673 585
R12077 gnd.n6262 gnd.n2956 585
R12078 gnd.n5222 gnd.n2956 585
R12079 gnd.n6263 gnd.n2955 585
R12080 gnd.n3691 gnd.n2955 585
R12081 gnd.n6264 gnd.n2954 585
R12082 gnd.n5214 gnd.n2954 585
R12083 gnd.n3697 gnd.n2952 585
R12084 gnd.n5207 gnd.n3697 585
R12085 gnd.n6268 gnd.n2951 585
R12086 gnd.n3703 gnd.n2951 585
R12087 gnd.n6269 gnd.n2950 585
R12088 gnd.n3702 gnd.n2950 585
R12089 gnd.n6270 gnd.n2949 585
R12090 gnd.n3707 gnd.n2949 585
R12091 gnd.n3713 gnd.n2947 585
R12092 gnd.n3714 gnd.n3713 585
R12093 gnd.n6274 gnd.n2946 585
R12094 gnd.n5175 gnd.n2946 585
R12095 gnd.n6275 gnd.n2945 585
R12096 gnd.n3718 gnd.n2945 585
R12097 gnd.n6276 gnd.n2944 585
R12098 gnd.n5156 gnd.n2944 585
R12099 gnd.n5147 gnd.n2942 585
R12100 gnd.n5148 gnd.n5147 585
R12101 gnd.n6280 gnd.n2941 585
R12102 gnd.n3738 gnd.n2941 585
R12103 gnd.n6281 gnd.n2940 585
R12104 gnd.n5127 gnd.n2940 585
R12105 gnd.n6282 gnd.n2939 585
R12106 gnd.n3742 gnd.n2939 585
R12107 gnd.n5116 gnd.n2937 585
R12108 gnd.n5117 gnd.n5116 585
R12109 gnd.n6286 gnd.n2936 585
R12110 gnd.n3755 gnd.n2936 585
R12111 gnd.n6287 gnd.n2935 585
R12112 gnd.n5099 gnd.n2935 585
R12113 gnd.n6288 gnd.n2934 585
R12114 gnd.n3771 gnd.n2934 585
R12115 gnd.n5090 gnd.n2932 585
R12116 gnd.n5091 gnd.n5090 585
R12117 gnd.n6292 gnd.n2931 585
R12118 gnd.n5083 gnd.n2931 585
R12119 gnd.n6293 gnd.n2930 585
R12120 gnd.n3783 gnd.n2930 585
R12121 gnd.n6294 gnd.n2929 585
R12122 gnd.n3781 gnd.n2929 585
R12123 gnd.n3787 gnd.n2927 585
R12124 gnd.n3788 gnd.n3787 585
R12125 gnd.n6298 gnd.n2926 585
R12126 gnd.n3794 gnd.n2926 585
R12127 gnd.n6299 gnd.n2925 585
R12128 gnd.t348 gnd.n2925 585
R12129 gnd.n6300 gnd.n2924 585
R12130 gnd.n3798 gnd.n2924 585
R12131 gnd.n5032 gnd.n2922 585
R12132 gnd.n5033 gnd.n5032 585
R12133 gnd.n6304 gnd.n2921 585
R12134 gnd.n5024 gnd.n2921 585
R12135 gnd.n6305 gnd.n2920 585
R12136 gnd.n5012 gnd.n2920 585
R12137 gnd.n6306 gnd.n2919 585
R12138 gnd.n5004 gnd.n2919 585
R12139 gnd.n2916 gnd.n2914 585
R12140 gnd.n3823 gnd.n2914 585
R12141 gnd.n6311 gnd.n6310 585
R12142 gnd.n6312 gnd.n6311 585
R12143 gnd.n2915 gnd.n2913 585
R12144 gnd.n4982 gnd.n2913 585
R12145 gnd.n4795 gnd.n2902 585
R12146 gnd.n6318 gnd.n2902 585
R12147 gnd.n4796 gnd.n4794 585
R12148 gnd.n4794 gnd.n2897 585
R12149 gnd.n4793 gnd.n4791 585
R12150 gnd.n4793 gnd.n2871 585
R12151 gnd.n4800 gnd.n4790 585
R12152 gnd.n4790 gnd.n2839 585
R12153 gnd.n4801 gnd.n4789 585
R12154 gnd.n4789 gnd.n3910 585
R12155 gnd.n4802 gnd.n3911 585
R12156 gnd.n4825 gnd.n3911 585
R12157 gnd.n3923 gnd.n3921 585
R12158 gnd.n3921 gnd.n3909 585
R12159 gnd.n4807 gnd.n4806 585
R12160 gnd.n4808 gnd.n4807 585
R12161 gnd.n3922 gnd.n3920 585
R12162 gnd.n3920 gnd.n3918 585
R12163 gnd.n4785 gnd.n4784 585
R12164 gnd.n4784 gnd.n4783 585
R12165 gnd.n3926 gnd.n3925 585
R12166 gnd.n3927 gnd.n3926 585
R12167 gnd.n6143 gnd.n3066 585
R12168 gnd.n6144 gnd.n3065 585
R12169 gnd.n3415 gnd.n3059 585
R12170 gnd.n6151 gnd.n3058 585
R12171 gnd.n6152 gnd.n3057 585
R12172 gnd.n3412 gnd.n3051 585
R12173 gnd.n6159 gnd.n3050 585
R12174 gnd.n6160 gnd.n3049 585
R12175 gnd.n3410 gnd.n3043 585
R12176 gnd.n6167 gnd.n3042 585
R12177 gnd.n6168 gnd.n3041 585
R12178 gnd.n3407 gnd.n3035 585
R12179 gnd.n6175 gnd.n3034 585
R12180 gnd.n6176 gnd.n3033 585
R12181 gnd.n3405 gnd.n3026 585
R12182 gnd.n6183 gnd.n3025 585
R12183 gnd.n6184 gnd.n3024 585
R12184 gnd.n3402 gnd.n3021 585
R12185 gnd.n6189 gnd.n3020 585
R12186 gnd.n6190 gnd.n3019 585
R12187 gnd.n6191 gnd.n3018 585
R12188 gnd.n3399 gnd.n3016 585
R12189 gnd.n6195 gnd.n3015 585
R12190 gnd.n6196 gnd.n3014 585
R12191 gnd.n6197 gnd.n3010 585
R12192 gnd.n5685 gnd.n3005 585
R12193 gnd.n5682 gnd.n3005 585
R12194 gnd.n5686 gnd.n5684 585
R12195 gnd.n3397 gnd.n3396 585
R12196 gnd.n3418 gnd.n3417 585
R12197 gnd.n5539 gnd.n5538 468.476
R12198 gnd.n5422 gnd.n5421 468.476
R12199 gnd.n3893 gnd.n3891 468.476
R12200 gnd.n6388 gnd.n2874 468.476
R12201 gnd.n7006 gnd.n7005 452.659
R12202 gnd.n3827 gnd.t316 389.64
R12203 gnd.n3510 gnd.t264 389.64
R12204 gnd.n6325 gnd.t233 389.64
R12205 gnd.n3504 gnd.t319 389.64
R12206 gnd.n4564 gnd.t281 371.625
R12207 gnd.n6137 gnd.t310 371.625
R12208 gnd.n3953 gnd.t328 371.625
R12209 gnd.n3139 gnd.t303 371.625
R12210 gnd.n3162 gnd.t294 371.625
R12211 gnd.n6017 gnd.t225 371.625
R12212 gnd.n352 gnd.t334 371.625
R12213 gnd.n332 gnd.t237 371.625
R12214 gnd.n7938 gnd.t271 371.625
R12215 gnd.n7738 gnd.t285 371.625
R12216 gnd.n2416 gnd.t300 371.625
R12217 gnd.n2438 gnd.t229 371.625
R12218 gnd.n2460 gnd.t254 371.625
R12219 gnd.n4107 gnd.t331 371.625
R12220 gnd.n2822 gnd.t325 371.625
R12221 gnd.n4623 gnd.t250 371.625
R12222 gnd.n4636 gnd.t278 371.625
R12223 gnd.n3067 gnd.t257 371.625
R12224 gnd.n1495 gnd.t274 323.425
R12225 gnd.n1012 gnd.t306 323.425
R12226 gnd.n2324 gnd.n2298 289.615
R12227 gnd.n2292 gnd.n2266 289.615
R12228 gnd.n2260 gnd.n2234 289.615
R12229 gnd.n2229 gnd.n2203 289.615
R12230 gnd.n2197 gnd.n2171 289.615
R12231 gnd.n2165 gnd.n2139 289.615
R12232 gnd.n2133 gnd.n2107 289.615
R12233 gnd.n2102 gnd.n2076 289.615
R12234 gnd.n1569 gnd.t221 279.217
R12235 gnd.n1033 gnd.t337 279.217
R12236 gnd.n2881 gnd.t246 260.649
R12237 gnd.n3472 gnd.t290 260.649
R12238 gnd.n6390 gnd.n6389 256.663
R12239 gnd.n6390 gnd.n2840 256.663
R12240 gnd.n6390 gnd.n2841 256.663
R12241 gnd.n6390 gnd.n2842 256.663
R12242 gnd.n6390 gnd.n2843 256.663
R12243 gnd.n6390 gnd.n2844 256.663
R12244 gnd.n6390 gnd.n2845 256.663
R12245 gnd.n6390 gnd.n2846 256.663
R12246 gnd.n6390 gnd.n2847 256.663
R12247 gnd.n6390 gnd.n2848 256.663
R12248 gnd.n6390 gnd.n2849 256.663
R12249 gnd.n6390 gnd.n2850 256.663
R12250 gnd.n6390 gnd.n2851 256.663
R12251 gnd.n6390 gnd.n2852 256.663
R12252 gnd.n6390 gnd.n2853 256.663
R12253 gnd.n6390 gnd.n2854 256.663
R12254 gnd.n6393 gnd.n2837 256.663
R12255 gnd.n6391 gnd.n6390 256.663
R12256 gnd.n6390 gnd.n2855 256.663
R12257 gnd.n6390 gnd.n2856 256.663
R12258 gnd.n6390 gnd.n2857 256.663
R12259 gnd.n6390 gnd.n2858 256.663
R12260 gnd.n6390 gnd.n2859 256.663
R12261 gnd.n6390 gnd.n2860 256.663
R12262 gnd.n6390 gnd.n2861 256.663
R12263 gnd.n6390 gnd.n2862 256.663
R12264 gnd.n6390 gnd.n2863 256.663
R12265 gnd.n6390 gnd.n2864 256.663
R12266 gnd.n6390 gnd.n2865 256.663
R12267 gnd.n6390 gnd.n2866 256.663
R12268 gnd.n6390 gnd.n2867 256.663
R12269 gnd.n6390 gnd.n2868 256.663
R12270 gnd.n6390 gnd.n2869 256.663
R12271 gnd.n6390 gnd.n2870 256.663
R12272 gnd.n3534 gnd.n3447 256.663
R12273 gnd.n5427 gnd.n3447 256.663
R12274 gnd.n3531 gnd.n3447 256.663
R12275 gnd.n5434 gnd.n3447 256.663
R12276 gnd.n3528 gnd.n3447 256.663
R12277 gnd.n5441 gnd.n3447 256.663
R12278 gnd.n3525 gnd.n3447 256.663
R12279 gnd.n5448 gnd.n3447 256.663
R12280 gnd.n3522 gnd.n3447 256.663
R12281 gnd.n5455 gnd.n3447 256.663
R12282 gnd.n3519 gnd.n3447 256.663
R12283 gnd.n5462 gnd.n3447 256.663
R12284 gnd.n3516 gnd.n3447 256.663
R12285 gnd.n5469 gnd.n3447 256.663
R12286 gnd.n3513 gnd.n3447 256.663
R12287 gnd.n5477 gnd.n3447 256.663
R12288 gnd.n5480 gnd.n3149 256.663
R12289 gnd.n5481 gnd.n3447 256.663
R12290 gnd.n3507 gnd.n3447 256.663
R12291 gnd.n5488 gnd.n3447 256.663
R12292 gnd.n3502 gnd.n3447 256.663
R12293 gnd.n5495 gnd.n3447 256.663
R12294 gnd.n3499 gnd.n3447 256.663
R12295 gnd.n5502 gnd.n3447 256.663
R12296 gnd.n3496 gnd.n3447 256.663
R12297 gnd.n5509 gnd.n3447 256.663
R12298 gnd.n3493 gnd.n3447 256.663
R12299 gnd.n5516 gnd.n3447 256.663
R12300 gnd.n3490 gnd.n3447 256.663
R12301 gnd.n5523 gnd.n3447 256.663
R12302 gnd.n3487 gnd.n3447 256.663
R12303 gnd.n5530 gnd.n3447 256.663
R12304 gnd.n3484 gnd.n3447 256.663
R12305 gnd.n5537 gnd.n3447 256.663
R12306 gnd.n6745 gnd.n2384 242.672
R12307 gnd.n6745 gnd.n2385 242.672
R12308 gnd.n6745 gnd.n2386 242.672
R12309 gnd.n6745 gnd.n2387 242.672
R12310 gnd.n6745 gnd.n2388 242.672
R12311 gnd.n6745 gnd.n2389 242.672
R12312 gnd.n6745 gnd.n2390 242.672
R12313 gnd.n6745 gnd.n2391 242.672
R12314 gnd.n6745 gnd.n2392 242.672
R12315 gnd.n6444 gnd.n2775 242.672
R12316 gnd.n6444 gnd.n2774 242.672
R12317 gnd.n6444 gnd.n2773 242.672
R12318 gnd.n6444 gnd.n2772 242.672
R12319 gnd.n6444 gnd.n2771 242.672
R12320 gnd.n6444 gnd.n2770 242.672
R12321 gnd.n6444 gnd.n2769 242.672
R12322 gnd.n6444 gnd.n2768 242.672
R12323 gnd.n6444 gnd.n2767 242.672
R12324 gnd.n1623 gnd.n1622 242.672
R12325 gnd.n1623 gnd.n1533 242.672
R12326 gnd.n1623 gnd.n1534 242.672
R12327 gnd.n1623 gnd.n1535 242.672
R12328 gnd.n1623 gnd.n1536 242.672
R12329 gnd.n1623 gnd.n1537 242.672
R12330 gnd.n1623 gnd.n1538 242.672
R12331 gnd.n1623 gnd.n1539 242.672
R12332 gnd.n1623 gnd.n1540 242.672
R12333 gnd.n1623 gnd.n1541 242.672
R12334 gnd.n1623 gnd.n1542 242.672
R12335 gnd.n1623 gnd.n1543 242.672
R12336 gnd.n1624 gnd.n1623 242.672
R12337 gnd.n6792 gnd.n2355 242.672
R12338 gnd.n6792 gnd.n1029 242.672
R12339 gnd.n6792 gnd.n1028 242.672
R12340 gnd.n6792 gnd.n1027 242.672
R12341 gnd.n6792 gnd.n1026 242.672
R12342 gnd.n6792 gnd.n1025 242.672
R12343 gnd.n6792 gnd.n1024 242.672
R12344 gnd.n6792 gnd.n1023 242.672
R12345 gnd.n6792 gnd.n1022 242.672
R12346 gnd.n6792 gnd.n1021 242.672
R12347 gnd.n6792 gnd.n1020 242.672
R12348 gnd.n6792 gnd.n1019 242.672
R12349 gnd.n6792 gnd.n1018 242.672
R12350 gnd.n6134 gnd.n3104 242.672
R12351 gnd.n6134 gnd.n3106 242.672
R12352 gnd.n6134 gnd.n3107 242.672
R12353 gnd.n6134 gnd.n3109 242.672
R12354 gnd.n6134 gnd.n3111 242.672
R12355 gnd.n6134 gnd.n3112 242.672
R12356 gnd.n6134 gnd.n3114 242.672
R12357 gnd.n6134 gnd.n3116 242.672
R12358 gnd.n6135 gnd.n6134 242.672
R12359 gnd.n7973 gnd.n266 242.672
R12360 gnd.n7973 gnd.n265 242.672
R12361 gnd.n7973 gnd.n264 242.672
R12362 gnd.n7973 gnd.n263 242.672
R12363 gnd.n7973 gnd.n262 242.672
R12364 gnd.n7973 gnd.n261 242.672
R12365 gnd.n7973 gnd.n260 242.672
R12366 gnd.n7973 gnd.n259 242.672
R12367 gnd.n7973 gnd.n258 242.672
R12368 gnd.n1707 gnd.n1706 242.672
R12369 gnd.n1706 gnd.n1445 242.672
R12370 gnd.n1706 gnd.n1446 242.672
R12371 gnd.n1706 gnd.n1447 242.672
R12372 gnd.n1706 gnd.n1448 242.672
R12373 gnd.n1706 gnd.n1449 242.672
R12374 gnd.n1706 gnd.n1450 242.672
R12375 gnd.n1706 gnd.n1451 242.672
R12376 gnd.n6792 gnd.n1011 242.672
R12377 gnd.n6793 gnd.n6792 242.672
R12378 gnd.n6792 gnd.n6746 242.672
R12379 gnd.n6792 gnd.n6747 242.672
R12380 gnd.n6792 gnd.n6748 242.672
R12381 gnd.n6792 gnd.n6749 242.672
R12382 gnd.n6792 gnd.n6750 242.672
R12383 gnd.n6792 gnd.n6751 242.672
R12384 gnd.n6745 gnd.n6744 242.672
R12385 gnd.n6745 gnd.n2356 242.672
R12386 gnd.n6745 gnd.n2357 242.672
R12387 gnd.n6745 gnd.n2358 242.672
R12388 gnd.n6745 gnd.n2359 242.672
R12389 gnd.n6745 gnd.n2360 242.672
R12390 gnd.n6745 gnd.n2361 242.672
R12391 gnd.n6745 gnd.n2362 242.672
R12392 gnd.n6745 gnd.n2363 242.672
R12393 gnd.n6745 gnd.n2364 242.672
R12394 gnd.n6745 gnd.n2365 242.672
R12395 gnd.n6745 gnd.n2366 242.672
R12396 gnd.n6745 gnd.n2367 242.672
R12397 gnd.n6745 gnd.n2368 242.672
R12398 gnd.n6745 gnd.n2369 242.672
R12399 gnd.n6745 gnd.n2370 242.672
R12400 gnd.n6745 gnd.n2371 242.672
R12401 gnd.n6745 gnd.n2372 242.672
R12402 gnd.n6745 gnd.n2373 242.672
R12403 gnd.n6745 gnd.n2374 242.672
R12404 gnd.n6745 gnd.n2375 242.672
R12405 gnd.n6745 gnd.n2376 242.672
R12406 gnd.n6745 gnd.n2377 242.672
R12407 gnd.n6745 gnd.n2378 242.672
R12408 gnd.n6745 gnd.n2379 242.672
R12409 gnd.n6745 gnd.n2380 242.672
R12410 gnd.n6745 gnd.n2381 242.672
R12411 gnd.n6745 gnd.n2382 242.672
R12412 gnd.n6745 gnd.n2383 242.672
R12413 gnd.n6444 gnd.n2777 242.672
R12414 gnd.n6444 gnd.n2778 242.672
R12415 gnd.n6444 gnd.n2779 242.672
R12416 gnd.n6444 gnd.n2780 242.672
R12417 gnd.n6444 gnd.n2781 242.672
R12418 gnd.n6444 gnd.n2782 242.672
R12419 gnd.n6444 gnd.n2783 242.672
R12420 gnd.n6444 gnd.n2784 242.672
R12421 gnd.n6444 gnd.n2785 242.672
R12422 gnd.n6444 gnd.n2786 242.672
R12423 gnd.n6444 gnd.n2787 242.672
R12424 gnd.n6444 gnd.n2788 242.672
R12425 gnd.n6444 gnd.n2789 242.672
R12426 gnd.n6444 gnd.n2790 242.672
R12427 gnd.n6444 gnd.n2791 242.672
R12428 gnd.n6444 gnd.n2792 242.672
R12429 gnd.n6394 gnd.n2833 242.672
R12430 gnd.n6444 gnd.n2793 242.672
R12431 gnd.n6444 gnd.n2794 242.672
R12432 gnd.n6444 gnd.n2795 242.672
R12433 gnd.n6444 gnd.n2796 242.672
R12434 gnd.n6444 gnd.n2797 242.672
R12435 gnd.n6444 gnd.n2798 242.672
R12436 gnd.n6444 gnd.n2799 242.672
R12437 gnd.n6444 gnd.n2800 242.672
R12438 gnd.n6444 gnd.n2801 242.672
R12439 gnd.n6444 gnd.n2802 242.672
R12440 gnd.n6444 gnd.n2803 242.672
R12441 gnd.n6444 gnd.n2804 242.672
R12442 gnd.n6444 gnd.n6443 242.672
R12443 gnd.n6134 gnd.n6133 242.672
R12444 gnd.n6134 gnd.n3076 242.672
R12445 gnd.n6134 gnd.n3077 242.672
R12446 gnd.n6134 gnd.n3078 242.672
R12447 gnd.n6134 gnd.n3079 242.672
R12448 gnd.n6134 gnd.n3080 242.672
R12449 gnd.n6134 gnd.n3081 242.672
R12450 gnd.n6134 gnd.n3082 242.672
R12451 gnd.n6134 gnd.n3083 242.672
R12452 gnd.n6134 gnd.n3084 242.672
R12453 gnd.n6134 gnd.n3085 242.672
R12454 gnd.n6134 gnd.n3086 242.672
R12455 gnd.n6134 gnd.n3087 242.672
R12456 gnd.n6081 gnd.n3150 242.672
R12457 gnd.n6134 gnd.n3088 242.672
R12458 gnd.n6134 gnd.n3089 242.672
R12459 gnd.n6134 gnd.n3090 242.672
R12460 gnd.n6134 gnd.n3091 242.672
R12461 gnd.n6134 gnd.n3092 242.672
R12462 gnd.n6134 gnd.n3093 242.672
R12463 gnd.n6134 gnd.n3094 242.672
R12464 gnd.n6134 gnd.n3095 242.672
R12465 gnd.n6134 gnd.n3096 242.672
R12466 gnd.n6134 gnd.n3097 242.672
R12467 gnd.n6134 gnd.n3098 242.672
R12468 gnd.n6134 gnd.n3099 242.672
R12469 gnd.n6134 gnd.n3100 242.672
R12470 gnd.n6134 gnd.n3101 242.672
R12471 gnd.n6134 gnd.n3102 242.672
R12472 gnd.n6134 gnd.n3103 242.672
R12473 gnd.n7973 gnd.n267 242.672
R12474 gnd.n7973 gnd.n268 242.672
R12475 gnd.n7973 gnd.n269 242.672
R12476 gnd.n7973 gnd.n270 242.672
R12477 gnd.n7973 gnd.n271 242.672
R12478 gnd.n7973 gnd.n272 242.672
R12479 gnd.n7973 gnd.n273 242.672
R12480 gnd.n7973 gnd.n274 242.672
R12481 gnd.n7973 gnd.n275 242.672
R12482 gnd.n7973 gnd.n276 242.672
R12483 gnd.n7973 gnd.n277 242.672
R12484 gnd.n7973 gnd.n278 242.672
R12485 gnd.n7973 gnd.n279 242.672
R12486 gnd.n7973 gnd.n280 242.672
R12487 gnd.n7973 gnd.n281 242.672
R12488 gnd.n7973 gnd.n282 242.672
R12489 gnd.n7973 gnd.n283 242.672
R12490 gnd.n7973 gnd.n284 242.672
R12491 gnd.n7973 gnd.n285 242.672
R12492 gnd.n7973 gnd.n286 242.672
R12493 gnd.n7973 gnd.n287 242.672
R12494 gnd.n7973 gnd.n288 242.672
R12495 gnd.n7973 gnd.n289 242.672
R12496 gnd.n7973 gnd.n290 242.672
R12497 gnd.n7973 gnd.n291 242.672
R12498 gnd.n7973 gnd.n292 242.672
R12499 gnd.n7973 gnd.n293 242.672
R12500 gnd.n7973 gnd.n294 242.672
R12501 gnd.n7973 gnd.n7972 242.672
R12502 gnd.n4774 gnd.n3935 242.672
R12503 gnd.n4774 gnd.n3936 242.672
R12504 gnd.n4774 gnd.n3937 242.672
R12505 gnd.n4774 gnd.n3938 242.672
R12506 gnd.n4774 gnd.n3939 242.672
R12507 gnd.n4774 gnd.n3940 242.672
R12508 gnd.n4774 gnd.n3941 242.672
R12509 gnd.n4774 gnd.n3942 242.672
R12510 gnd.n4774 gnd.n3943 242.672
R12511 gnd.n4774 gnd.n3944 242.672
R12512 gnd.n4774 gnd.n3945 242.672
R12513 gnd.n4774 gnd.n3946 242.672
R12514 gnd.n4774 gnd.n3947 242.672
R12515 gnd.n4774 gnd.n3948 242.672
R12516 gnd.n5682 gnd.n3419 242.672
R12517 gnd.n5682 gnd.n3416 242.672
R12518 gnd.n5682 gnd.n3414 242.672
R12519 gnd.n5682 gnd.n3413 242.672
R12520 gnd.n5682 gnd.n3411 242.672
R12521 gnd.n5682 gnd.n3409 242.672
R12522 gnd.n5682 gnd.n3408 242.672
R12523 gnd.n5682 gnd.n3406 242.672
R12524 gnd.n5682 gnd.n3404 242.672
R12525 gnd.n5682 gnd.n3403 242.672
R12526 gnd.n5682 gnd.n3401 242.672
R12527 gnd.n5682 gnd.n3400 242.672
R12528 gnd.n5682 gnd.n3398 242.672
R12529 gnd.n5683 gnd.n5682 242.672
R12530 gnd.n7974 gnd.n255 240.244
R12531 gnd.n7971 gnd.n295 240.244
R12532 gnd.n7967 gnd.n7966 240.244
R12533 gnd.n7963 gnd.n7962 240.244
R12534 gnd.n7959 gnd.n7958 240.244
R12535 gnd.n7955 gnd.n7954 240.244
R12536 gnd.n7951 gnd.n7950 240.244
R12537 gnd.n7947 gnd.n7946 240.244
R12538 gnd.n7943 gnd.n7942 240.244
R12539 gnd.n7936 gnd.n7935 240.244
R12540 gnd.n7932 gnd.n7931 240.244
R12541 gnd.n7928 gnd.n7927 240.244
R12542 gnd.n7924 gnd.n7923 240.244
R12543 gnd.n7920 gnd.n7919 240.244
R12544 gnd.n7916 gnd.n7915 240.244
R12545 gnd.n7912 gnd.n7911 240.244
R12546 gnd.n7908 gnd.n7907 240.244
R12547 gnd.n7904 gnd.n7903 240.244
R12548 gnd.n7900 gnd.n7899 240.244
R12549 gnd.n7893 gnd.n7892 240.244
R12550 gnd.n7890 gnd.n7889 240.244
R12551 gnd.n7886 gnd.n7885 240.244
R12552 gnd.n7882 gnd.n7881 240.244
R12553 gnd.n7878 gnd.n7877 240.244
R12554 gnd.n7874 gnd.n7873 240.244
R12555 gnd.n7870 gnd.n7869 240.244
R12556 gnd.n7866 gnd.n7865 240.244
R12557 gnd.n7862 gnd.n7861 240.244
R12558 gnd.n7858 gnd.n7857 240.244
R12559 gnd.n6014 gnd.n3183 240.244
R12560 gnd.n6006 gnd.n3183 240.244
R12561 gnd.n6006 gnd.n3194 240.244
R12562 gnd.n3210 gnd.n3194 240.244
R12563 gnd.n5702 gnd.n3210 240.244
R12564 gnd.n5702 gnd.n3223 240.244
R12565 gnd.n5707 gnd.n3223 240.244
R12566 gnd.n5707 gnd.n3234 240.244
R12567 gnd.n5717 gnd.n3234 240.244
R12568 gnd.n5717 gnd.n3244 240.244
R12569 gnd.n5722 gnd.n3244 240.244
R12570 gnd.n5722 gnd.n3255 240.244
R12571 gnd.n5732 gnd.n3255 240.244
R12572 gnd.n5732 gnd.n3264 240.244
R12573 gnd.n5737 gnd.n3264 240.244
R12574 gnd.n5737 gnd.n3275 240.244
R12575 gnd.n5747 gnd.n3275 240.244
R12576 gnd.n5747 gnd.n3285 240.244
R12577 gnd.n5752 gnd.n3285 240.244
R12578 gnd.n5752 gnd.n3296 240.244
R12579 gnd.n5762 gnd.n3296 240.244
R12580 gnd.n5762 gnd.n3305 240.244
R12581 gnd.n5767 gnd.n3305 240.244
R12582 gnd.n5767 gnd.n3317 240.244
R12583 gnd.n5789 gnd.n3317 240.244
R12584 gnd.n5789 gnd.n3327 240.244
R12585 gnd.n3331 gnd.n3327 240.244
R12586 gnd.n5794 gnd.n3331 240.244
R12587 gnd.n5794 gnd.n5793 240.244
R12588 gnd.n5793 gnd.n3341 240.244
R12589 gnd.n3351 gnd.n3341 240.244
R12590 gnd.n3363 gnd.n3351 240.244
R12591 gnd.n5907 gnd.n3363 240.244
R12592 gnd.n5907 gnd.n102 240.244
R12593 gnd.n5903 gnd.n102 240.244
R12594 gnd.n5903 gnd.n5810 240.244
R12595 gnd.n5810 gnd.n119 240.244
R12596 gnd.n5826 gnd.n119 240.244
R12597 gnd.n5826 gnd.n130 240.244
R12598 gnd.n5883 gnd.n130 240.244
R12599 gnd.n5883 gnd.n140 240.244
R12600 gnd.n5879 gnd.n140 240.244
R12601 gnd.n5879 gnd.n149 240.244
R12602 gnd.n5871 gnd.n149 240.244
R12603 gnd.n5871 gnd.n160 240.244
R12604 gnd.n360 gnd.n160 240.244
R12605 gnd.n360 gnd.n169 240.244
R12606 gnd.n7822 gnd.n169 240.244
R12607 gnd.n7822 gnd.n180 240.244
R12608 gnd.n7825 gnd.n180 240.244
R12609 gnd.n7825 gnd.n189 240.244
R12610 gnd.n7829 gnd.n189 240.244
R12611 gnd.n7829 gnd.n200 240.244
R12612 gnd.n7832 gnd.n200 240.244
R12613 gnd.n7832 gnd.n209 240.244
R12614 gnd.n7836 gnd.n209 240.244
R12615 gnd.n7836 gnd.n219 240.244
R12616 gnd.n7839 gnd.n219 240.244
R12617 gnd.n7839 gnd.n228 240.244
R12618 gnd.n7843 gnd.n228 240.244
R12619 gnd.n7843 gnd.n238 240.244
R12620 gnd.n7846 gnd.n238 240.244
R12621 gnd.n7846 gnd.n247 240.244
R12622 gnd.n7850 gnd.n247 240.244
R12623 gnd.n3119 gnd.n3118 240.244
R12624 gnd.n6127 gnd.n3118 240.244
R12625 gnd.n6125 gnd.n6124 240.244
R12626 gnd.n6121 gnd.n6120 240.244
R12627 gnd.n6117 gnd.n6116 240.244
R12628 gnd.n6113 gnd.n6112 240.244
R12629 gnd.n6109 gnd.n6108 240.244
R12630 gnd.n6105 gnd.n6104 240.244
R12631 gnd.n6101 gnd.n6100 240.244
R12632 gnd.n6096 gnd.n6095 240.244
R12633 gnd.n6092 gnd.n6091 240.244
R12634 gnd.n6088 gnd.n6087 240.244
R12635 gnd.n6084 gnd.n6083 240.244
R12636 gnd.n6079 gnd.n6078 240.244
R12637 gnd.n6075 gnd.n6074 240.244
R12638 gnd.n6071 gnd.n6070 240.244
R12639 gnd.n6067 gnd.n6066 240.244
R12640 gnd.n6063 gnd.n6062 240.244
R12641 gnd.n6059 gnd.n6058 240.244
R12642 gnd.n6055 gnd.n6054 240.244
R12643 gnd.n6051 gnd.n6050 240.244
R12644 gnd.n6047 gnd.n6046 240.244
R12645 gnd.n6043 gnd.n6042 240.244
R12646 gnd.n6039 gnd.n6038 240.244
R12647 gnd.n6035 gnd.n6034 240.244
R12648 gnd.n6031 gnd.n6030 240.244
R12649 gnd.n6027 gnd.n6026 240.244
R12650 gnd.n6023 gnd.n6022 240.244
R12651 gnd.n3198 gnd.n3120 240.244
R12652 gnd.n6004 gnd.n3198 240.244
R12653 gnd.n6004 gnd.n3199 240.244
R12654 gnd.n6000 gnd.n3199 240.244
R12655 gnd.n6000 gnd.n3208 240.244
R12656 gnd.n5992 gnd.n3208 240.244
R12657 gnd.n5992 gnd.n3226 240.244
R12658 gnd.n5988 gnd.n3226 240.244
R12659 gnd.n5988 gnd.n3232 240.244
R12660 gnd.n5980 gnd.n3232 240.244
R12661 gnd.n5980 gnd.n3247 240.244
R12662 gnd.n5976 gnd.n3247 240.244
R12663 gnd.n5976 gnd.n3253 240.244
R12664 gnd.n5968 gnd.n3253 240.244
R12665 gnd.n5968 gnd.n3267 240.244
R12666 gnd.n5964 gnd.n3267 240.244
R12667 gnd.n5964 gnd.n3273 240.244
R12668 gnd.n5956 gnd.n3273 240.244
R12669 gnd.n5956 gnd.n3288 240.244
R12670 gnd.n5952 gnd.n3288 240.244
R12671 gnd.n5952 gnd.n3294 240.244
R12672 gnd.n5944 gnd.n3294 240.244
R12673 gnd.n5944 gnd.n3308 240.244
R12674 gnd.n5940 gnd.n3308 240.244
R12675 gnd.n5940 gnd.n3315 240.244
R12676 gnd.n5932 gnd.n3315 240.244
R12677 gnd.n5932 gnd.n5929 240.244
R12678 gnd.n5929 gnd.n3330 240.244
R12679 gnd.n3347 gnd.n3330 240.244
R12680 gnd.n5918 gnd.n3347 240.244
R12681 gnd.n5918 gnd.n5915 240.244
R12682 gnd.n5915 gnd.n3350 240.244
R12683 gnd.n3350 gnd.n105 240.244
R12684 gnd.n8066 gnd.n105 240.244
R12685 gnd.n8066 gnd.n106 240.244
R12686 gnd.n116 gnd.n106 240.244
R12687 gnd.n8060 gnd.n116 240.244
R12688 gnd.n8060 gnd.n117 240.244
R12689 gnd.n8052 gnd.n117 240.244
R12690 gnd.n8052 gnd.n133 240.244
R12691 gnd.n8048 gnd.n133 240.244
R12692 gnd.n8048 gnd.n138 240.244
R12693 gnd.n8040 gnd.n138 240.244
R12694 gnd.n8040 gnd.n152 240.244
R12695 gnd.n8036 gnd.n152 240.244
R12696 gnd.n8036 gnd.n158 240.244
R12697 gnd.n8028 gnd.n158 240.244
R12698 gnd.n8028 gnd.n172 240.244
R12699 gnd.n8024 gnd.n172 240.244
R12700 gnd.n8024 gnd.n178 240.244
R12701 gnd.n8016 gnd.n178 240.244
R12702 gnd.n8016 gnd.n192 240.244
R12703 gnd.n8012 gnd.n192 240.244
R12704 gnd.n8012 gnd.n198 240.244
R12705 gnd.n8004 gnd.n198 240.244
R12706 gnd.n8004 gnd.n212 240.244
R12707 gnd.n8000 gnd.n212 240.244
R12708 gnd.n8000 gnd.n218 240.244
R12709 gnd.n7992 gnd.n218 240.244
R12710 gnd.n7992 gnd.n231 240.244
R12711 gnd.n7988 gnd.n231 240.244
R12712 gnd.n7988 gnd.n237 240.244
R12713 gnd.n7980 gnd.n237 240.244
R12714 gnd.n7980 gnd.n250 240.244
R12715 gnd.n6445 gnd.n2764 240.244
R12716 gnd.n6442 gnd.n2805 240.244
R12717 gnd.n6438 gnd.n6437 240.244
R12718 gnd.n6434 gnd.n6433 240.244
R12719 gnd.n6430 gnd.n6429 240.244
R12720 gnd.n6426 gnd.n6425 240.244
R12721 gnd.n6422 gnd.n6421 240.244
R12722 gnd.n6418 gnd.n6417 240.244
R12723 gnd.n6414 gnd.n6413 240.244
R12724 gnd.n6409 gnd.n6408 240.244
R12725 gnd.n6405 gnd.n6404 240.244
R12726 gnd.n6401 gnd.n6400 240.244
R12727 gnd.n6397 gnd.n6396 240.244
R12728 gnd.n4645 gnd.n4644 240.244
R12729 gnd.n4648 gnd.n4647 240.244
R12730 gnd.n4655 gnd.n4654 240.244
R12731 gnd.n4658 gnd.n4657 240.244
R12732 gnd.n4663 gnd.n4638 240.244
R12733 gnd.n4667 gnd.n4666 240.244
R12734 gnd.n4674 gnd.n4673 240.244
R12735 gnd.n4677 gnd.n4676 240.244
R12736 gnd.n4684 gnd.n4683 240.244
R12737 gnd.n4687 gnd.n4686 240.244
R12738 gnd.n4694 gnd.n4693 240.244
R12739 gnd.n4697 gnd.n4696 240.244
R12740 gnd.n4704 gnd.n4703 240.244
R12741 gnd.n4707 gnd.n4706 240.244
R12742 gnd.n4712 gnd.n4625 240.244
R12743 gnd.n6623 gnd.n6622 240.244
R12744 gnd.n6622 gnd.n2467 240.244
R12745 gnd.n2479 gnd.n2467 240.244
R12746 gnd.n4076 gnd.n2479 240.244
R12747 gnd.n4076 gnd.n2491 240.244
R12748 gnd.n4080 gnd.n2491 240.244
R12749 gnd.n4080 gnd.n2501 240.244
R12750 gnd.n4083 gnd.n2501 240.244
R12751 gnd.n4083 gnd.n2510 240.244
R12752 gnd.n4087 gnd.n2510 240.244
R12753 gnd.n4087 gnd.n2520 240.244
R12754 gnd.n4090 gnd.n2520 240.244
R12755 gnd.n4090 gnd.n2530 240.244
R12756 gnd.n4094 gnd.n2530 240.244
R12757 gnd.n4094 gnd.n2540 240.244
R12758 gnd.n4200 gnd.n2540 240.244
R12759 gnd.n4200 gnd.n2550 240.244
R12760 gnd.n4068 gnd.n2550 240.244
R12761 gnd.n4068 gnd.n2560 240.244
R12762 gnd.n4210 gnd.n2560 240.244
R12763 gnd.n4210 gnd.n2570 240.244
R12764 gnd.n4063 gnd.n2570 240.244
R12765 gnd.n4063 gnd.n2580 240.244
R12766 gnd.n4258 gnd.n2580 240.244
R12767 gnd.n4258 gnd.n2590 240.244
R12768 gnd.n4054 gnd.n2590 240.244
R12769 gnd.n4054 gnd.n2599 240.244
R12770 gnd.n4274 gnd.n2599 240.244
R12771 gnd.n4274 gnd.n2609 240.244
R12772 gnd.n4045 gnd.n2609 240.244
R12773 gnd.n4045 gnd.n4039 240.244
R12774 gnd.n4316 gnd.n4039 240.244
R12775 gnd.n4316 gnd.n4031 240.244
R12776 gnd.n4031 gnd.n4024 240.244
R12777 gnd.n4323 gnd.n4024 240.244
R12778 gnd.n4323 gnd.n4017 240.244
R12779 gnd.n4017 gnd.n2625 240.244
R12780 gnd.n4010 gnd.n2625 240.244
R12781 gnd.n4010 gnd.n2636 240.244
R12782 gnd.n4385 gnd.n2636 240.244
R12783 gnd.n4385 gnd.n2646 240.244
R12784 gnd.n4389 gnd.n2646 240.244
R12785 gnd.n4389 gnd.n2655 240.244
R12786 gnd.n4399 gnd.n2655 240.244
R12787 gnd.n4399 gnd.n2666 240.244
R12788 gnd.n3991 gnd.n2666 240.244
R12789 gnd.n3991 gnd.n2675 240.244
R12790 gnd.n4406 gnd.n2675 240.244
R12791 gnd.n4406 gnd.n2686 240.244
R12792 gnd.n4411 gnd.n2686 240.244
R12793 gnd.n4411 gnd.n2695 240.244
R12794 gnd.n4418 gnd.n2695 240.244
R12795 gnd.n4418 gnd.n2706 240.244
R12796 gnd.n3979 gnd.n2706 240.244
R12797 gnd.n3979 gnd.n2715 240.244
R12798 gnd.n4466 gnd.n2715 240.244
R12799 gnd.n4466 gnd.n2726 240.244
R12800 gnd.n3968 gnd.n2726 240.244
R12801 gnd.n3968 gnd.n2735 240.244
R12802 gnd.n4473 gnd.n2735 240.244
R12803 gnd.n4473 gnd.n2746 240.244
R12804 gnd.n4723 gnd.n2746 240.244
R12805 gnd.n4723 gnd.n2756 240.244
R12806 gnd.n3957 gnd.n2756 240.244
R12807 gnd.n2396 gnd.n2395 240.244
R12808 gnd.n6738 gnd.n2395 240.244
R12809 gnd.n6736 gnd.n6735 240.244
R12810 gnd.n6732 gnd.n6731 240.244
R12811 gnd.n6728 gnd.n6727 240.244
R12812 gnd.n6724 gnd.n6723 240.244
R12813 gnd.n6720 gnd.n6719 240.244
R12814 gnd.n6716 gnd.n6715 240.244
R12815 gnd.n6712 gnd.n6711 240.244
R12816 gnd.n6707 gnd.n6706 240.244
R12817 gnd.n6703 gnd.n6702 240.244
R12818 gnd.n6699 gnd.n6698 240.244
R12819 gnd.n6695 gnd.n6694 240.244
R12820 gnd.n6691 gnd.n6690 240.244
R12821 gnd.n6687 gnd.n6686 240.244
R12822 gnd.n6683 gnd.n6682 240.244
R12823 gnd.n6679 gnd.n6678 240.244
R12824 gnd.n6675 gnd.n6674 240.244
R12825 gnd.n6671 gnd.n6670 240.244
R12826 gnd.n6667 gnd.n6666 240.244
R12827 gnd.n6663 gnd.n6662 240.244
R12828 gnd.n6659 gnd.n6658 240.244
R12829 gnd.n6655 gnd.n6654 240.244
R12830 gnd.n6651 gnd.n6650 240.244
R12831 gnd.n6647 gnd.n6646 240.244
R12832 gnd.n6643 gnd.n6642 240.244
R12833 gnd.n6639 gnd.n6638 240.244
R12834 gnd.n6635 gnd.n6634 240.244
R12835 gnd.n6631 gnd.n6630 240.244
R12836 gnd.n6620 gnd.n2397 240.244
R12837 gnd.n6620 gnd.n2470 240.244
R12838 gnd.n6616 gnd.n2470 240.244
R12839 gnd.n6616 gnd.n2477 240.244
R12840 gnd.n6608 gnd.n2477 240.244
R12841 gnd.n6608 gnd.n2494 240.244
R12842 gnd.n6604 gnd.n2494 240.244
R12843 gnd.n6604 gnd.n2500 240.244
R12844 gnd.n6596 gnd.n2500 240.244
R12845 gnd.n6596 gnd.n2512 240.244
R12846 gnd.n6592 gnd.n2512 240.244
R12847 gnd.n6592 gnd.n2518 240.244
R12848 gnd.n6584 gnd.n2518 240.244
R12849 gnd.n6584 gnd.n2533 240.244
R12850 gnd.n6580 gnd.n2533 240.244
R12851 gnd.n6580 gnd.n2539 240.244
R12852 gnd.n6572 gnd.n2539 240.244
R12853 gnd.n6572 gnd.n2552 240.244
R12854 gnd.n6568 gnd.n2552 240.244
R12855 gnd.n6568 gnd.n2558 240.244
R12856 gnd.n6560 gnd.n2558 240.244
R12857 gnd.n6560 gnd.n2573 240.244
R12858 gnd.n6556 gnd.n2573 240.244
R12859 gnd.n6556 gnd.n2579 240.244
R12860 gnd.n6548 gnd.n2579 240.244
R12861 gnd.n6548 gnd.n2592 240.244
R12862 gnd.n6544 gnd.n2592 240.244
R12863 gnd.n6544 gnd.n2597 240.244
R12864 gnd.n6536 gnd.n2597 240.244
R12865 gnd.n6536 gnd.n2612 240.244
R12866 gnd.n4265 gnd.n2612 240.244
R12867 gnd.n4265 gnd.n4027 240.244
R12868 gnd.n4332 gnd.n4027 240.244
R12869 gnd.n4336 gnd.n4332 240.244
R12870 gnd.n4336 gnd.n4333 240.244
R12871 gnd.n4333 gnd.n2622 240.244
R12872 gnd.n6531 gnd.n2622 240.244
R12873 gnd.n6531 gnd.n2623 240.244
R12874 gnd.n6523 gnd.n2623 240.244
R12875 gnd.n6523 gnd.n2639 240.244
R12876 gnd.n6519 gnd.n2639 240.244
R12877 gnd.n6519 gnd.n2644 240.244
R12878 gnd.n6511 gnd.n2644 240.244
R12879 gnd.n6511 gnd.n2658 240.244
R12880 gnd.n6507 gnd.n2658 240.244
R12881 gnd.n6507 gnd.n2664 240.244
R12882 gnd.n6499 gnd.n2664 240.244
R12883 gnd.n6499 gnd.n2678 240.244
R12884 gnd.n6495 gnd.n2678 240.244
R12885 gnd.n6495 gnd.n2684 240.244
R12886 gnd.n6487 gnd.n2684 240.244
R12887 gnd.n6487 gnd.n2698 240.244
R12888 gnd.n6483 gnd.n2698 240.244
R12889 gnd.n6483 gnd.n2704 240.244
R12890 gnd.n6475 gnd.n2704 240.244
R12891 gnd.n6475 gnd.n2718 240.244
R12892 gnd.n6471 gnd.n2718 240.244
R12893 gnd.n6471 gnd.n2724 240.244
R12894 gnd.n6463 gnd.n2724 240.244
R12895 gnd.n6463 gnd.n2738 240.244
R12896 gnd.n6459 gnd.n2738 240.244
R12897 gnd.n6459 gnd.n2744 240.244
R12898 gnd.n6451 gnd.n2744 240.244
R12899 gnd.n6451 gnd.n2759 240.244
R12900 gnd.n6791 gnd.n6752 240.244
R12901 gnd.n6784 gnd.n6783 240.244
R12902 gnd.n6781 gnd.n6780 240.244
R12903 gnd.n6777 gnd.n6776 240.244
R12904 gnd.n6773 gnd.n6772 240.244
R12905 gnd.n6769 gnd.n6768 240.244
R12906 gnd.n6765 gnd.n1017 240.244
R12907 gnd.n6795 gnd.n6794 240.244
R12908 gnd.n1718 gnd.n1430 240.244
R12909 gnd.n1728 gnd.n1430 240.244
R12910 gnd.n1728 gnd.n1421 240.244
R12911 gnd.n1421 gnd.n1410 240.244
R12912 gnd.n1749 gnd.n1410 240.244
R12913 gnd.n1749 gnd.n1404 240.244
R12914 gnd.n1759 gnd.n1404 240.244
R12915 gnd.n1759 gnd.n1393 240.244
R12916 gnd.n1393 gnd.n1383 240.244
R12917 gnd.n1785 gnd.n1383 240.244
R12918 gnd.n1786 gnd.n1785 240.244
R12919 gnd.n1787 gnd.n1786 240.244
R12920 gnd.n1787 gnd.n1362 240.244
R12921 gnd.n1823 gnd.n1362 240.244
R12922 gnd.n1823 gnd.n1363 240.244
R12923 gnd.n1819 gnd.n1363 240.244
R12924 gnd.n1819 gnd.n1818 240.244
R12925 gnd.n1818 gnd.n1239 240.244
R12926 gnd.n1853 gnd.n1239 240.244
R12927 gnd.n1853 gnd.n1229 240.244
R12928 gnd.n1229 gnd.n1221 240.244
R12929 gnd.n1871 gnd.n1221 240.244
R12930 gnd.n1872 gnd.n1871 240.244
R12931 gnd.n1872 gnd.n1209 240.244
R12932 gnd.n1209 gnd.n1198 240.244
R12933 gnd.n1903 gnd.n1198 240.244
R12934 gnd.n1904 gnd.n1903 240.244
R12935 gnd.n1906 gnd.n1904 240.244
R12936 gnd.n1906 gnd.n1184 240.244
R12937 gnd.n1938 gnd.n1184 240.244
R12938 gnd.n1938 gnd.n1170 240.244
R12939 gnd.n1960 gnd.n1170 240.244
R12940 gnd.n1961 gnd.n1960 240.244
R12941 gnd.n1961 gnd.n1157 240.244
R12942 gnd.n1157 gnd.n1147 240.244
R12943 gnd.n1992 gnd.n1147 240.244
R12944 gnd.n1993 gnd.n1992 240.244
R12945 gnd.n1994 gnd.n1993 240.244
R12946 gnd.n1994 gnd.n1132 240.244
R12947 gnd.n1996 gnd.n1132 240.244
R12948 gnd.n1996 gnd.n1118 240.244
R12949 gnd.n2065 gnd.n1118 240.244
R12950 gnd.n2066 gnd.n2065 240.244
R12951 gnd.n2067 gnd.n2066 240.244
R12952 gnd.n2067 gnd.n966 240.244
R12953 gnd.n1113 gnd.n966 240.244
R12954 gnd.n1113 gnd.n977 240.244
R12955 gnd.n2335 gnd.n977 240.244
R12956 gnd.n2336 gnd.n2335 240.244
R12957 gnd.n2336 gnd.n990 240.244
R12958 gnd.n2344 gnd.n990 240.244
R12959 gnd.n2344 gnd.n1002 240.244
R12960 gnd.n6802 gnd.n1002 240.244
R12961 gnd.n1708 gnd.n1443 240.244
R12962 gnd.n1464 gnd.n1443 240.244
R12963 gnd.n1467 gnd.n1466 240.244
R12964 gnd.n1474 gnd.n1473 240.244
R12965 gnd.n1477 gnd.n1476 240.244
R12966 gnd.n1484 gnd.n1483 240.244
R12967 gnd.n1487 gnd.n1486 240.244
R12968 gnd.n1494 gnd.n1493 240.244
R12969 gnd.n1716 gnd.n1440 240.244
R12970 gnd.n1440 gnd.n1419 240.244
R12971 gnd.n1739 gnd.n1419 240.244
R12972 gnd.n1739 gnd.n1413 240.244
R12973 gnd.n1747 gnd.n1413 240.244
R12974 gnd.n1747 gnd.n1415 240.244
R12975 gnd.n1415 gnd.n1391 240.244
R12976 gnd.n1769 gnd.n1391 240.244
R12977 gnd.n1769 gnd.n1386 240.244
R12978 gnd.n1783 gnd.n1386 240.244
R12979 gnd.n1783 gnd.n1387 240.244
R12980 gnd.n1779 gnd.n1387 240.244
R12981 gnd.n1779 gnd.n1359 240.244
R12982 gnd.n1826 gnd.n1359 240.244
R12983 gnd.n1827 gnd.n1826 240.244
R12984 gnd.n1828 gnd.n1827 240.244
R12985 gnd.n1828 gnd.n1355 240.244
R12986 gnd.n1834 gnd.n1355 240.244
R12987 gnd.n1834 gnd.n1228 240.244
R12988 gnd.n1863 gnd.n1228 240.244
R12989 gnd.n1863 gnd.n1224 240.244
R12990 gnd.n1869 gnd.n1224 240.244
R12991 gnd.n1869 gnd.n1207 240.244
R12992 gnd.n1893 gnd.n1207 240.244
R12993 gnd.n1893 gnd.n1202 240.244
R12994 gnd.n1901 gnd.n1202 240.244
R12995 gnd.n1901 gnd.n1203 240.244
R12996 gnd.n1203 gnd.n1182 240.244
R12997 gnd.n1942 gnd.n1182 240.244
R12998 gnd.n1942 gnd.n1177 240.244
R12999 gnd.n1950 gnd.n1177 240.244
R13000 gnd.n1950 gnd.n1178 240.244
R13001 gnd.n1178 gnd.n1155 240.244
R13002 gnd.n1982 gnd.n1155 240.244
R13003 gnd.n1982 gnd.n1150 240.244
R13004 gnd.n1990 gnd.n1150 240.244
R13005 gnd.n1990 gnd.n1151 240.244
R13006 gnd.n1151 gnd.n1130 240.244
R13007 gnd.n2043 gnd.n1130 240.244
R13008 gnd.n2043 gnd.n1125 240.244
R13009 gnd.n2055 gnd.n1125 240.244
R13010 gnd.n2055 gnd.n1126 240.244
R13011 gnd.n2051 gnd.n1126 240.244
R13012 gnd.n2051 gnd.n968 240.244
R13013 gnd.n6828 gnd.n968 240.244
R13014 gnd.n6828 gnd.n969 240.244
R13015 gnd.n6824 gnd.n969 240.244
R13016 gnd.n6824 gnd.n975 240.244
R13017 gnd.n991 gnd.n975 240.244
R13018 gnd.n6814 gnd.n991 240.244
R13019 gnd.n6814 gnd.n992 240.244
R13020 gnd.n6810 gnd.n992 240.244
R13021 gnd.n6810 gnd.n1000 240.244
R13022 gnd.n7749 gnd.n257 240.244
R13023 gnd.n7755 gnd.n7754 240.244
R13024 gnd.n7758 gnd.n7757 240.244
R13025 gnd.n7765 gnd.n7764 240.244
R13026 gnd.n7768 gnd.n7767 240.244
R13027 gnd.n7775 gnd.n7774 240.244
R13028 gnd.n7778 gnd.n7777 240.244
R13029 gnd.n7785 gnd.n7784 240.244
R13030 gnd.n7788 gnd.n7787 240.244
R13031 gnd.n3393 gnd.n3186 240.244
R13032 gnd.n3393 gnd.n3195 240.244
R13033 gnd.n5694 gnd.n3195 240.244
R13034 gnd.n5694 gnd.n3211 240.244
R13035 gnd.n5700 gnd.n3211 240.244
R13036 gnd.n5700 gnd.n3224 240.244
R13037 gnd.n5709 gnd.n3224 240.244
R13038 gnd.n5709 gnd.n3235 240.244
R13039 gnd.n5715 gnd.n3235 240.244
R13040 gnd.n5715 gnd.n3245 240.244
R13041 gnd.n5724 gnd.n3245 240.244
R13042 gnd.n5724 gnd.n3256 240.244
R13043 gnd.n5730 gnd.n3256 240.244
R13044 gnd.n5730 gnd.n3265 240.244
R13045 gnd.n5739 gnd.n3265 240.244
R13046 gnd.n5739 gnd.n3276 240.244
R13047 gnd.n5745 gnd.n3276 240.244
R13048 gnd.n5745 gnd.n3286 240.244
R13049 gnd.n5754 gnd.n3286 240.244
R13050 gnd.n5754 gnd.n3297 240.244
R13051 gnd.n5760 gnd.n3297 240.244
R13052 gnd.n5760 gnd.n3306 240.244
R13053 gnd.n5769 gnd.n3306 240.244
R13054 gnd.n5769 gnd.n3318 240.244
R13055 gnd.n5787 gnd.n3318 240.244
R13056 gnd.n5787 gnd.n3328 240.244
R13057 gnd.n3332 gnd.n3328 240.244
R13058 gnd.n5774 gnd.n3332 240.244
R13059 gnd.n5775 gnd.n5774 240.244
R13060 gnd.n5775 gnd.n3342 240.244
R13061 gnd.n3352 gnd.n3342 240.244
R13062 gnd.n3361 gnd.n3352 240.244
R13063 gnd.n3361 gnd.n98 240.244
R13064 gnd.n8068 gnd.n98 240.244
R13065 gnd.n8068 gnd.n100 240.244
R13066 gnd.n5830 gnd.n100 240.244
R13067 gnd.n5830 gnd.n120 240.244
R13068 gnd.n5889 gnd.n120 240.244
R13069 gnd.n5889 gnd.n131 240.244
R13070 gnd.n5885 gnd.n131 240.244
R13071 gnd.n5885 gnd.n141 240.244
R13072 gnd.n5877 gnd.n141 240.244
R13073 gnd.n5877 gnd.n150 240.244
R13074 gnd.n5873 gnd.n150 240.244
R13075 gnd.n5873 gnd.n161 240.244
R13076 gnd.n7717 gnd.n161 240.244
R13077 gnd.n7717 gnd.n170 240.244
R13078 gnd.n7820 gnd.n170 240.244
R13079 gnd.n7820 gnd.n181 240.244
R13080 gnd.n7816 gnd.n181 240.244
R13081 gnd.n7816 gnd.n190 240.244
R13082 gnd.n7813 gnd.n190 240.244
R13083 gnd.n7813 gnd.n201 240.244
R13084 gnd.n7810 gnd.n201 240.244
R13085 gnd.n7810 gnd.n210 240.244
R13086 gnd.n7807 gnd.n210 240.244
R13087 gnd.n7807 gnd.n220 240.244
R13088 gnd.n7804 gnd.n220 240.244
R13089 gnd.n7804 gnd.n229 240.244
R13090 gnd.n7801 gnd.n229 240.244
R13091 gnd.n7801 gnd.n239 240.244
R13092 gnd.n7798 gnd.n239 240.244
R13093 gnd.n7798 gnd.n248 240.244
R13094 gnd.n7795 gnd.n248 240.244
R13095 gnd.n3030 gnd.n3029 240.244
R13096 gnd.n3105 gnd.n3037 240.244
R13097 gnd.n3108 gnd.n3038 240.244
R13098 gnd.n3046 gnd.n3045 240.244
R13099 gnd.n3110 gnd.n3053 240.244
R13100 gnd.n3113 gnd.n3054 240.244
R13101 gnd.n3062 gnd.n3061 240.244
R13102 gnd.n3115 gnd.n3071 240.244
R13103 gnd.n6136 gnd.n3074 240.244
R13104 gnd.n6012 gnd.n3189 240.244
R13105 gnd.n3197 gnd.n3189 240.244
R13106 gnd.n3213 gnd.n3197 240.244
R13107 gnd.n5998 gnd.n3213 240.244
R13108 gnd.n5998 gnd.n3214 240.244
R13109 gnd.n5994 gnd.n3214 240.244
R13110 gnd.n5994 gnd.n3221 240.244
R13111 gnd.n5986 gnd.n3221 240.244
R13112 gnd.n5986 gnd.n3237 240.244
R13113 gnd.n5982 gnd.n3237 240.244
R13114 gnd.n5982 gnd.n3242 240.244
R13115 gnd.n5974 gnd.n3242 240.244
R13116 gnd.n5974 gnd.n3257 240.244
R13117 gnd.n5970 gnd.n3257 240.244
R13118 gnd.n5970 gnd.n3262 240.244
R13119 gnd.n5962 gnd.n3262 240.244
R13120 gnd.n5962 gnd.n3278 240.244
R13121 gnd.n5958 gnd.n3278 240.244
R13122 gnd.n5958 gnd.n3283 240.244
R13123 gnd.n5950 gnd.n3283 240.244
R13124 gnd.n5950 gnd.n3298 240.244
R13125 gnd.n5946 gnd.n3298 240.244
R13126 gnd.n5946 gnd.n3303 240.244
R13127 gnd.n5938 gnd.n3303 240.244
R13128 gnd.n5938 gnd.n3320 240.244
R13129 gnd.n5934 gnd.n3320 240.244
R13130 gnd.n5934 gnd.n3325 240.244
R13131 gnd.n5798 gnd.n3325 240.244
R13132 gnd.n5799 gnd.n5798 240.244
R13133 gnd.n5799 gnd.n3344 240.244
R13134 gnd.n5913 gnd.n3344 240.244
R13135 gnd.n5913 gnd.n3354 240.244
R13136 gnd.n5909 gnd.n3354 240.244
R13137 gnd.n5909 gnd.n104 240.244
R13138 gnd.n5901 gnd.n104 240.244
R13139 gnd.n5901 gnd.n122 240.244
R13140 gnd.n8058 gnd.n122 240.244
R13141 gnd.n8058 gnd.n123 240.244
R13142 gnd.n8054 gnd.n123 240.244
R13143 gnd.n8054 gnd.n129 240.244
R13144 gnd.n8046 gnd.n129 240.244
R13145 gnd.n8046 gnd.n142 240.244
R13146 gnd.n8042 gnd.n142 240.244
R13147 gnd.n8042 gnd.n147 240.244
R13148 gnd.n8034 gnd.n147 240.244
R13149 gnd.n8034 gnd.n163 240.244
R13150 gnd.n8030 gnd.n163 240.244
R13151 gnd.n8030 gnd.n168 240.244
R13152 gnd.n8022 gnd.n168 240.244
R13153 gnd.n8022 gnd.n182 240.244
R13154 gnd.n8018 gnd.n182 240.244
R13155 gnd.n8018 gnd.n187 240.244
R13156 gnd.n8010 gnd.n187 240.244
R13157 gnd.n8010 gnd.n203 240.244
R13158 gnd.n8006 gnd.n203 240.244
R13159 gnd.n8006 gnd.n208 240.244
R13160 gnd.n7998 gnd.n208 240.244
R13161 gnd.n7998 gnd.n221 240.244
R13162 gnd.n7994 gnd.n221 240.244
R13163 gnd.n7994 gnd.n226 240.244
R13164 gnd.n7986 gnd.n226 240.244
R13165 gnd.n7986 gnd.n241 240.244
R13166 gnd.n7982 gnd.n241 240.244
R13167 gnd.n7982 gnd.n246 240.244
R13168 gnd.n1046 gnd.n1006 240.244
R13169 gnd.n1054 gnd.n1053 240.244
R13170 gnd.n1057 gnd.n1056 240.244
R13171 gnd.n1064 gnd.n1063 240.244
R13172 gnd.n1067 gnd.n1066 240.244
R13173 gnd.n1074 gnd.n1073 240.244
R13174 gnd.n1077 gnd.n1076 240.244
R13175 gnd.n1084 gnd.n1083 240.244
R13176 gnd.n1087 gnd.n1086 240.244
R13177 gnd.n1094 gnd.n1093 240.244
R13178 gnd.n1097 gnd.n1096 240.244
R13179 gnd.n1104 gnd.n1103 240.244
R13180 gnd.n1106 gnd.n1030 240.244
R13181 gnd.n1631 gnd.n1528 240.244
R13182 gnd.n1631 gnd.n1521 240.244
R13183 gnd.n1642 gnd.n1521 240.244
R13184 gnd.n1642 gnd.n1517 240.244
R13185 gnd.n1648 gnd.n1517 240.244
R13186 gnd.n1648 gnd.n1509 240.244
R13187 gnd.n1658 gnd.n1509 240.244
R13188 gnd.n1658 gnd.n1504 240.244
R13189 gnd.n1694 gnd.n1504 240.244
R13190 gnd.n1694 gnd.n1505 240.244
R13191 gnd.n1505 gnd.n1452 240.244
R13192 gnd.n1689 gnd.n1452 240.244
R13193 gnd.n1689 gnd.n1688 240.244
R13194 gnd.n1688 gnd.n1431 240.244
R13195 gnd.n1684 gnd.n1431 240.244
R13196 gnd.n1684 gnd.n1422 240.244
R13197 gnd.n1681 gnd.n1422 240.244
R13198 gnd.n1681 gnd.n1680 240.244
R13199 gnd.n1680 gnd.n1405 240.244
R13200 gnd.n1676 gnd.n1405 240.244
R13201 gnd.n1676 gnd.n1394 240.244
R13202 gnd.n1394 gnd.n1374 240.244
R13203 gnd.n1795 gnd.n1374 240.244
R13204 gnd.n1795 gnd.n1369 240.244
R13205 gnd.n1803 gnd.n1369 240.244
R13206 gnd.n1803 gnd.n1370 240.244
R13207 gnd.n1370 gnd.n1338 240.244
R13208 gnd.n1843 gnd.n1338 240.244
R13209 gnd.n1843 gnd.n1339 240.244
R13210 gnd.n1354 gnd.n1339 240.244
R13211 gnd.n1354 gnd.n1241 240.244
R13212 gnd.n1850 gnd.n1241 240.244
R13213 gnd.n1850 gnd.n1230 240.244
R13214 gnd.n1243 gnd.n1230 240.244
R13215 gnd.n1243 gnd.n1220 240.244
R13216 gnd.n1250 gnd.n1220 240.244
R13217 gnd.n1250 gnd.n1210 240.244
R13218 gnd.n1247 gnd.n1210 240.244
R13219 gnd.n1247 gnd.n1189 240.244
R13220 gnd.n1915 gnd.n1189 240.244
R13221 gnd.n1915 gnd.n1185 240.244
R13222 gnd.n1937 gnd.n1185 240.244
R13223 gnd.n1937 gnd.n1175 240.244
R13224 gnd.n1933 gnd.n1175 240.244
R13225 gnd.n1933 gnd.n1169 240.244
R13226 gnd.n1930 gnd.n1169 240.244
R13227 gnd.n1930 gnd.n1158 240.244
R13228 gnd.n1927 gnd.n1158 240.244
R13229 gnd.n1927 gnd.n1137 240.244
R13230 gnd.n2005 gnd.n1137 240.244
R13231 gnd.n2005 gnd.n1133 240.244
R13232 gnd.n2040 gnd.n1133 240.244
R13233 gnd.n2040 gnd.n1124 240.244
R13234 gnd.n2036 gnd.n1124 240.244
R13235 gnd.n2036 gnd.n954 240.244
R13236 gnd.n2032 gnd.n954 240.244
R13237 gnd.n2032 gnd.n965 240.244
R13238 gnd.n2028 gnd.n965 240.244
R13239 gnd.n2028 gnd.n2027 240.244
R13240 gnd.n2027 gnd.n978 240.244
R13241 gnd.n2023 gnd.n978 240.244
R13242 gnd.n2023 gnd.n989 240.244
R13243 gnd.n2347 gnd.n989 240.244
R13244 gnd.n2348 gnd.n2347 240.244
R13245 gnd.n2348 gnd.n1003 240.244
R13246 gnd.n1545 gnd.n1544 240.244
R13247 gnd.n1616 gnd.n1544 240.244
R13248 gnd.n1614 gnd.n1613 240.244
R13249 gnd.n1610 gnd.n1609 240.244
R13250 gnd.n1606 gnd.n1605 240.244
R13251 gnd.n1602 gnd.n1601 240.244
R13252 gnd.n1598 gnd.n1597 240.244
R13253 gnd.n1594 gnd.n1593 240.244
R13254 gnd.n1590 gnd.n1589 240.244
R13255 gnd.n1586 gnd.n1585 240.244
R13256 gnd.n1582 gnd.n1581 240.244
R13257 gnd.n1578 gnd.n1577 240.244
R13258 gnd.n1574 gnd.n1532 240.244
R13259 gnd.n1634 gnd.n1526 240.244
R13260 gnd.n1634 gnd.n1522 240.244
R13261 gnd.n1640 gnd.n1522 240.244
R13262 gnd.n1640 gnd.n1515 240.244
R13263 gnd.n1650 gnd.n1515 240.244
R13264 gnd.n1650 gnd.n1511 240.244
R13265 gnd.n1656 gnd.n1511 240.244
R13266 gnd.n1656 gnd.n1502 240.244
R13267 gnd.n1696 gnd.n1502 240.244
R13268 gnd.n1696 gnd.n1453 240.244
R13269 gnd.n1704 gnd.n1453 240.244
R13270 gnd.n1704 gnd.n1454 240.244
R13271 gnd.n1454 gnd.n1432 240.244
R13272 gnd.n1725 gnd.n1432 240.244
R13273 gnd.n1725 gnd.n1424 240.244
R13274 gnd.n1736 gnd.n1424 240.244
R13275 gnd.n1736 gnd.n1425 240.244
R13276 gnd.n1425 gnd.n1406 240.244
R13277 gnd.n1756 gnd.n1406 240.244
R13278 gnd.n1756 gnd.n1396 240.244
R13279 gnd.n1766 gnd.n1396 240.244
R13280 gnd.n1766 gnd.n1377 240.244
R13281 gnd.n1793 gnd.n1377 240.244
R13282 gnd.n1793 gnd.n1367 240.244
R13283 gnd.n1806 gnd.n1367 240.244
R13284 gnd.n1807 gnd.n1806 240.244
R13285 gnd.n1807 gnd.n1342 240.244
R13286 gnd.n1841 gnd.n1342 240.244
R13287 gnd.n1841 gnd.n1343 240.244
R13288 gnd.n1837 gnd.n1343 240.244
R13289 gnd.n1837 gnd.n1351 240.244
R13290 gnd.n1351 gnd.n1232 240.244
R13291 gnd.n1860 gnd.n1232 240.244
R13292 gnd.n1860 gnd.n1219 240.244
R13293 gnd.n1875 gnd.n1219 240.244
R13294 gnd.n1875 gnd.n1212 240.244
R13295 gnd.n1890 gnd.n1212 240.244
R13296 gnd.n1890 gnd.n1213 240.244
R13297 gnd.n1213 gnd.n1191 240.244
R13298 gnd.n1913 gnd.n1191 240.244
R13299 gnd.n1913 gnd.n1192 240.244
R13300 gnd.n1192 gnd.n1174 240.244
R13301 gnd.n1953 gnd.n1174 240.244
R13302 gnd.n1953 gnd.n1167 240.244
R13303 gnd.n1964 gnd.n1167 240.244
R13304 gnd.n1964 gnd.n1160 240.244
R13305 gnd.n1979 gnd.n1160 240.244
R13306 gnd.n1979 gnd.n1161 240.244
R13307 gnd.n1161 gnd.n1140 240.244
R13308 gnd.n2003 gnd.n1140 240.244
R13309 gnd.n2003 gnd.n1141 240.244
R13310 gnd.n1141 gnd.n1122 240.244
R13311 gnd.n2058 gnd.n1122 240.244
R13312 gnd.n2058 gnd.n956 240.244
R13313 gnd.n6835 gnd.n956 240.244
R13314 gnd.n6835 gnd.n957 240.244
R13315 gnd.n6831 gnd.n957 240.244
R13316 gnd.n6831 gnd.n963 240.244
R13317 gnd.n980 gnd.n963 240.244
R13318 gnd.n6821 gnd.n980 240.244
R13319 gnd.n6821 gnd.n981 240.244
R13320 gnd.n6817 gnd.n981 240.244
R13321 gnd.n6817 gnd.n987 240.244
R13322 gnd.n1005 gnd.n987 240.244
R13323 gnd.n6807 gnd.n1005 240.244
R13324 gnd.n4510 gnd.n2766 240.244
R13325 gnd.n4520 gnd.n4519 240.244
R13326 gnd.n4522 gnd.n4521 240.244
R13327 gnd.n4530 gnd.n4529 240.244
R13328 gnd.n4540 gnd.n4539 240.244
R13329 gnd.n4542 gnd.n4541 240.244
R13330 gnd.n4550 gnd.n4549 240.244
R13331 gnd.n4560 gnd.n4559 240.244
R13332 gnd.n4562 gnd.n4561 240.244
R13333 gnd.n4164 gnd.n2468 240.244
R13334 gnd.n4167 gnd.n2468 240.244
R13335 gnd.n4167 gnd.n2480 240.244
R13336 gnd.n4172 gnd.n2480 240.244
R13337 gnd.n4172 gnd.n2492 240.244
R13338 gnd.n4175 gnd.n2492 240.244
R13339 gnd.n4175 gnd.n2502 240.244
R13340 gnd.n4180 gnd.n2502 240.244
R13341 gnd.n4180 gnd.n2511 240.244
R13342 gnd.n4183 gnd.n2511 240.244
R13343 gnd.n4183 gnd.n2521 240.244
R13344 gnd.n4188 gnd.n2521 240.244
R13345 gnd.n4188 gnd.n2531 240.244
R13346 gnd.n4191 gnd.n2531 240.244
R13347 gnd.n4191 gnd.n2541 240.244
R13348 gnd.n4198 gnd.n2541 240.244
R13349 gnd.n4198 gnd.n2551 240.244
R13350 gnd.n4216 gnd.n2551 240.244
R13351 gnd.n4216 gnd.n2561 240.244
R13352 gnd.n4212 gnd.n2561 240.244
R13353 gnd.n4212 gnd.n2571 240.244
R13354 gnd.n4249 gnd.n2571 240.244
R13355 gnd.n4249 gnd.n2581 240.244
R13356 gnd.n4256 gnd.n2581 240.244
R13357 gnd.n4256 gnd.n2591 240.244
R13358 gnd.n4280 gnd.n2591 240.244
R13359 gnd.n4280 gnd.n2600 240.244
R13360 gnd.n4276 gnd.n2600 240.244
R13361 gnd.n4276 gnd.n2610 240.244
R13362 gnd.n4308 gnd.n2610 240.244
R13363 gnd.n4308 gnd.n4041 240.244
R13364 gnd.n4314 gnd.n4041 240.244
R13365 gnd.n4314 gnd.n4022 240.244
R13366 gnd.n4338 gnd.n4022 240.244
R13367 gnd.n4338 gnd.n4018 240.244
R13368 gnd.n4344 gnd.n4018 240.244
R13369 gnd.n4344 gnd.n2626 240.244
R13370 gnd.n4377 gnd.n2626 240.244
R13371 gnd.n4377 gnd.n2637 240.244
R13372 gnd.n4383 gnd.n2637 240.244
R13373 gnd.n4383 gnd.n2647 240.244
R13374 gnd.n4391 gnd.n2647 240.244
R13375 gnd.n4391 gnd.n2656 240.244
R13376 gnd.n4397 gnd.n2656 240.244
R13377 gnd.n4397 gnd.n2667 240.244
R13378 gnd.n4432 gnd.n2667 240.244
R13379 gnd.n4432 gnd.n2676 240.244
R13380 gnd.n3996 gnd.n2676 240.244
R13381 gnd.n3996 gnd.n2687 240.244
R13382 gnd.n3997 gnd.n2687 240.244
R13383 gnd.n3997 gnd.n2696 240.244
R13384 gnd.n4420 gnd.n2696 240.244
R13385 gnd.n4420 gnd.n2707 240.244
R13386 gnd.n4458 gnd.n2707 240.244
R13387 gnd.n4458 gnd.n2716 240.244
R13388 gnd.n4464 gnd.n2716 240.244
R13389 gnd.n4464 gnd.n2727 240.244
R13390 gnd.n4736 gnd.n2727 240.244
R13391 gnd.n4736 gnd.n2736 240.244
R13392 gnd.n3973 gnd.n2736 240.244
R13393 gnd.n3973 gnd.n2747 240.244
R13394 gnd.n4725 gnd.n2747 240.244
R13395 gnd.n4725 gnd.n2757 240.244
R13396 gnd.n4765 gnd.n2757 240.244
R13397 gnd.n4124 gnd.n4123 240.244
R13398 gnd.n4130 gnd.n4129 240.244
R13399 gnd.n4134 gnd.n4133 240.244
R13400 gnd.n4140 gnd.n4139 240.244
R13401 gnd.n4144 gnd.n4143 240.244
R13402 gnd.n4150 gnd.n4149 240.244
R13403 gnd.n4154 gnd.n4153 240.244
R13404 gnd.n4111 gnd.n4110 240.244
R13405 gnd.n4106 gnd.n2393 240.244
R13406 gnd.n4119 gnd.n2469 240.244
R13407 gnd.n2482 gnd.n2469 240.244
R13408 gnd.n6614 gnd.n2482 240.244
R13409 gnd.n6614 gnd.n2483 240.244
R13410 gnd.n6610 gnd.n2483 240.244
R13411 gnd.n6610 gnd.n2490 240.244
R13412 gnd.n6602 gnd.n2490 240.244
R13413 gnd.n6602 gnd.n2504 240.244
R13414 gnd.n6598 gnd.n2504 240.244
R13415 gnd.n6598 gnd.n2509 240.244
R13416 gnd.n6590 gnd.n2509 240.244
R13417 gnd.n6590 gnd.n2523 240.244
R13418 gnd.n6586 gnd.n2523 240.244
R13419 gnd.n6586 gnd.n2528 240.244
R13420 gnd.n6578 gnd.n2528 240.244
R13421 gnd.n6578 gnd.n2543 240.244
R13422 gnd.n6574 gnd.n2543 240.244
R13423 gnd.n6574 gnd.n2548 240.244
R13424 gnd.n6566 gnd.n2548 240.244
R13425 gnd.n6566 gnd.n2563 240.244
R13426 gnd.n6562 gnd.n2563 240.244
R13427 gnd.n6562 gnd.n2568 240.244
R13428 gnd.n6554 gnd.n2568 240.244
R13429 gnd.n6554 gnd.n2583 240.244
R13430 gnd.n6550 gnd.n2583 240.244
R13431 gnd.n6550 gnd.n2588 240.244
R13432 gnd.n6542 gnd.n2588 240.244
R13433 gnd.n6542 gnd.n2602 240.244
R13434 gnd.n6538 gnd.n2602 240.244
R13435 gnd.n6538 gnd.n2607 240.244
R13436 gnd.n4267 gnd.n2607 240.244
R13437 gnd.n4267 gnd.n4032 240.244
R13438 gnd.n4330 gnd.n4032 240.244
R13439 gnd.n4330 gnd.n4026 240.244
R13440 gnd.n4326 gnd.n4026 240.244
R13441 gnd.n4326 gnd.n2628 240.244
R13442 gnd.n6529 gnd.n2628 240.244
R13443 gnd.n6529 gnd.n2629 240.244
R13444 gnd.n6525 gnd.n2629 240.244
R13445 gnd.n6525 gnd.n2635 240.244
R13446 gnd.n6517 gnd.n2635 240.244
R13447 gnd.n6517 gnd.n2648 240.244
R13448 gnd.n6513 gnd.n2648 240.244
R13449 gnd.n6513 gnd.n2653 240.244
R13450 gnd.n6505 gnd.n2653 240.244
R13451 gnd.n6505 gnd.n2669 240.244
R13452 gnd.n6501 gnd.n2669 240.244
R13453 gnd.n6501 gnd.n2674 240.244
R13454 gnd.n6493 gnd.n2674 240.244
R13455 gnd.n6493 gnd.n2688 240.244
R13456 gnd.n6489 gnd.n2688 240.244
R13457 gnd.n6489 gnd.n2693 240.244
R13458 gnd.n6481 gnd.n2693 240.244
R13459 gnd.n6481 gnd.n2709 240.244
R13460 gnd.n6477 gnd.n2709 240.244
R13461 gnd.n6477 gnd.n2714 240.244
R13462 gnd.n6469 gnd.n2714 240.244
R13463 gnd.n6469 gnd.n2728 240.244
R13464 gnd.n6465 gnd.n2728 240.244
R13465 gnd.n6465 gnd.n2733 240.244
R13466 gnd.n6457 gnd.n2733 240.244
R13467 gnd.n6457 gnd.n2749 240.244
R13468 gnd.n6453 gnd.n2749 240.244
R13469 gnd.n6453 gnd.n2754 240.244
R13470 gnd.n7008 gnd.n785 240.244
R13471 gnd.n7008 gnd.n781 240.244
R13472 gnd.n7014 gnd.n781 240.244
R13473 gnd.n7014 gnd.n779 240.244
R13474 gnd.n7018 gnd.n779 240.244
R13475 gnd.n7018 gnd.n775 240.244
R13476 gnd.n7024 gnd.n775 240.244
R13477 gnd.n7024 gnd.n773 240.244
R13478 gnd.n7028 gnd.n773 240.244
R13479 gnd.n7028 gnd.n769 240.244
R13480 gnd.n7034 gnd.n769 240.244
R13481 gnd.n7034 gnd.n767 240.244
R13482 gnd.n7038 gnd.n767 240.244
R13483 gnd.n7038 gnd.n763 240.244
R13484 gnd.n7044 gnd.n763 240.244
R13485 gnd.n7044 gnd.n761 240.244
R13486 gnd.n7048 gnd.n761 240.244
R13487 gnd.n7048 gnd.n757 240.244
R13488 gnd.n7054 gnd.n757 240.244
R13489 gnd.n7054 gnd.n755 240.244
R13490 gnd.n7058 gnd.n755 240.244
R13491 gnd.n7058 gnd.n751 240.244
R13492 gnd.n7064 gnd.n751 240.244
R13493 gnd.n7064 gnd.n749 240.244
R13494 gnd.n7068 gnd.n749 240.244
R13495 gnd.n7068 gnd.n745 240.244
R13496 gnd.n7074 gnd.n745 240.244
R13497 gnd.n7074 gnd.n743 240.244
R13498 gnd.n7078 gnd.n743 240.244
R13499 gnd.n7078 gnd.n739 240.244
R13500 gnd.n7084 gnd.n739 240.244
R13501 gnd.n7084 gnd.n737 240.244
R13502 gnd.n7088 gnd.n737 240.244
R13503 gnd.n7088 gnd.n733 240.244
R13504 gnd.n7094 gnd.n733 240.244
R13505 gnd.n7094 gnd.n731 240.244
R13506 gnd.n7098 gnd.n731 240.244
R13507 gnd.n7098 gnd.n727 240.244
R13508 gnd.n7104 gnd.n727 240.244
R13509 gnd.n7104 gnd.n725 240.244
R13510 gnd.n7108 gnd.n725 240.244
R13511 gnd.n7108 gnd.n721 240.244
R13512 gnd.n7114 gnd.n721 240.244
R13513 gnd.n7114 gnd.n719 240.244
R13514 gnd.n7118 gnd.n719 240.244
R13515 gnd.n7118 gnd.n715 240.244
R13516 gnd.n7124 gnd.n715 240.244
R13517 gnd.n7124 gnd.n713 240.244
R13518 gnd.n7128 gnd.n713 240.244
R13519 gnd.n7128 gnd.n709 240.244
R13520 gnd.n7134 gnd.n709 240.244
R13521 gnd.n7134 gnd.n707 240.244
R13522 gnd.n7138 gnd.n707 240.244
R13523 gnd.n7138 gnd.n703 240.244
R13524 gnd.n7144 gnd.n703 240.244
R13525 gnd.n7144 gnd.n701 240.244
R13526 gnd.n7148 gnd.n701 240.244
R13527 gnd.n7148 gnd.n697 240.244
R13528 gnd.n7154 gnd.n697 240.244
R13529 gnd.n7154 gnd.n695 240.244
R13530 gnd.n7158 gnd.n695 240.244
R13531 gnd.n7158 gnd.n691 240.244
R13532 gnd.n7164 gnd.n691 240.244
R13533 gnd.n7164 gnd.n689 240.244
R13534 gnd.n7168 gnd.n689 240.244
R13535 gnd.n7168 gnd.n685 240.244
R13536 gnd.n7174 gnd.n685 240.244
R13537 gnd.n7174 gnd.n683 240.244
R13538 gnd.n7178 gnd.n683 240.244
R13539 gnd.n7178 gnd.n679 240.244
R13540 gnd.n7184 gnd.n679 240.244
R13541 gnd.n7184 gnd.n677 240.244
R13542 gnd.n7188 gnd.n677 240.244
R13543 gnd.n7188 gnd.n673 240.244
R13544 gnd.n7194 gnd.n673 240.244
R13545 gnd.n7194 gnd.n671 240.244
R13546 gnd.n7198 gnd.n671 240.244
R13547 gnd.n7198 gnd.n667 240.244
R13548 gnd.n7204 gnd.n667 240.244
R13549 gnd.n7204 gnd.n665 240.244
R13550 gnd.n7208 gnd.n665 240.244
R13551 gnd.n7208 gnd.n661 240.244
R13552 gnd.n7214 gnd.n661 240.244
R13553 gnd.n7214 gnd.n659 240.244
R13554 gnd.n7218 gnd.n659 240.244
R13555 gnd.n7218 gnd.n655 240.244
R13556 gnd.n7224 gnd.n655 240.244
R13557 gnd.n7224 gnd.n653 240.244
R13558 gnd.n7228 gnd.n653 240.244
R13559 gnd.n7228 gnd.n649 240.244
R13560 gnd.n7234 gnd.n649 240.244
R13561 gnd.n7234 gnd.n647 240.244
R13562 gnd.n7238 gnd.n647 240.244
R13563 gnd.n7238 gnd.n643 240.244
R13564 gnd.n7244 gnd.n643 240.244
R13565 gnd.n7244 gnd.n641 240.244
R13566 gnd.n7248 gnd.n641 240.244
R13567 gnd.n7248 gnd.n637 240.244
R13568 gnd.n7254 gnd.n637 240.244
R13569 gnd.n7254 gnd.n635 240.244
R13570 gnd.n7258 gnd.n635 240.244
R13571 gnd.n7258 gnd.n631 240.244
R13572 gnd.n7264 gnd.n631 240.244
R13573 gnd.n7264 gnd.n629 240.244
R13574 gnd.n7268 gnd.n629 240.244
R13575 gnd.n7268 gnd.n625 240.244
R13576 gnd.n7274 gnd.n625 240.244
R13577 gnd.n7274 gnd.n623 240.244
R13578 gnd.n7278 gnd.n623 240.244
R13579 gnd.n7278 gnd.n619 240.244
R13580 gnd.n7284 gnd.n619 240.244
R13581 gnd.n7284 gnd.n617 240.244
R13582 gnd.n7288 gnd.n617 240.244
R13583 gnd.n7288 gnd.n613 240.244
R13584 gnd.n7294 gnd.n613 240.244
R13585 gnd.n7294 gnd.n611 240.244
R13586 gnd.n7298 gnd.n611 240.244
R13587 gnd.n7298 gnd.n607 240.244
R13588 gnd.n7304 gnd.n607 240.244
R13589 gnd.n7304 gnd.n605 240.244
R13590 gnd.n7308 gnd.n605 240.244
R13591 gnd.n7308 gnd.n601 240.244
R13592 gnd.n7314 gnd.n601 240.244
R13593 gnd.n7314 gnd.n599 240.244
R13594 gnd.n7318 gnd.n599 240.244
R13595 gnd.n7318 gnd.n595 240.244
R13596 gnd.n7324 gnd.n595 240.244
R13597 gnd.n7324 gnd.n593 240.244
R13598 gnd.n7328 gnd.n593 240.244
R13599 gnd.n7328 gnd.n589 240.244
R13600 gnd.n7334 gnd.n589 240.244
R13601 gnd.n7334 gnd.n587 240.244
R13602 gnd.n7338 gnd.n587 240.244
R13603 gnd.n7338 gnd.n583 240.244
R13604 gnd.n7344 gnd.n583 240.244
R13605 gnd.n7344 gnd.n581 240.244
R13606 gnd.n7348 gnd.n581 240.244
R13607 gnd.n7348 gnd.n577 240.244
R13608 gnd.n7354 gnd.n577 240.244
R13609 gnd.n7354 gnd.n575 240.244
R13610 gnd.n7358 gnd.n575 240.244
R13611 gnd.n7358 gnd.n571 240.244
R13612 gnd.n7364 gnd.n571 240.244
R13613 gnd.n7364 gnd.n569 240.244
R13614 gnd.n7368 gnd.n569 240.244
R13615 gnd.n7368 gnd.n565 240.244
R13616 gnd.n7374 gnd.n565 240.244
R13617 gnd.n7374 gnd.n563 240.244
R13618 gnd.n7378 gnd.n563 240.244
R13619 gnd.n7378 gnd.n559 240.244
R13620 gnd.n7384 gnd.n559 240.244
R13621 gnd.n7384 gnd.n557 240.244
R13622 gnd.n7388 gnd.n557 240.244
R13623 gnd.n7388 gnd.n553 240.244
R13624 gnd.n7394 gnd.n553 240.244
R13625 gnd.n7394 gnd.n551 240.244
R13626 gnd.n7398 gnd.n551 240.244
R13627 gnd.n7398 gnd.n547 240.244
R13628 gnd.n7404 gnd.n547 240.244
R13629 gnd.n7404 gnd.n545 240.244
R13630 gnd.n7408 gnd.n545 240.244
R13631 gnd.n7408 gnd.n541 240.244
R13632 gnd.n7414 gnd.n541 240.244
R13633 gnd.n7414 gnd.n539 240.244
R13634 gnd.n7418 gnd.n539 240.244
R13635 gnd.n7418 gnd.n535 240.244
R13636 gnd.n7424 gnd.n535 240.244
R13637 gnd.n7424 gnd.n533 240.244
R13638 gnd.n7428 gnd.n533 240.244
R13639 gnd.n7428 gnd.n529 240.244
R13640 gnd.n7434 gnd.n529 240.244
R13641 gnd.n7434 gnd.n527 240.244
R13642 gnd.n7438 gnd.n527 240.244
R13643 gnd.n7438 gnd.n523 240.244
R13644 gnd.n7444 gnd.n523 240.244
R13645 gnd.n7444 gnd.n521 240.244
R13646 gnd.n7448 gnd.n521 240.244
R13647 gnd.n7448 gnd.n517 240.244
R13648 gnd.n7454 gnd.n517 240.244
R13649 gnd.n7454 gnd.n515 240.244
R13650 gnd.n7458 gnd.n515 240.244
R13651 gnd.n7458 gnd.n511 240.244
R13652 gnd.n7464 gnd.n511 240.244
R13653 gnd.n7464 gnd.n509 240.244
R13654 gnd.n7468 gnd.n509 240.244
R13655 gnd.n7468 gnd.n505 240.244
R13656 gnd.n7474 gnd.n505 240.244
R13657 gnd.n7474 gnd.n503 240.244
R13658 gnd.n7478 gnd.n503 240.244
R13659 gnd.n7478 gnd.n499 240.244
R13660 gnd.n7485 gnd.n499 240.244
R13661 gnd.n7485 gnd.n497 240.244
R13662 gnd.n7489 gnd.n497 240.244
R13663 gnd.n7489 gnd.n494 240.244
R13664 gnd.n7495 gnd.n492 240.244
R13665 gnd.n7499 gnd.n492 240.244
R13666 gnd.n7499 gnd.n488 240.244
R13667 gnd.n7505 gnd.n488 240.244
R13668 gnd.n7505 gnd.n486 240.244
R13669 gnd.n7509 gnd.n486 240.244
R13670 gnd.n7509 gnd.n482 240.244
R13671 gnd.n7515 gnd.n482 240.244
R13672 gnd.n7515 gnd.n480 240.244
R13673 gnd.n7519 gnd.n480 240.244
R13674 gnd.n7519 gnd.n476 240.244
R13675 gnd.n7525 gnd.n476 240.244
R13676 gnd.n7525 gnd.n474 240.244
R13677 gnd.n7529 gnd.n474 240.244
R13678 gnd.n7529 gnd.n470 240.244
R13679 gnd.n7535 gnd.n470 240.244
R13680 gnd.n7535 gnd.n468 240.244
R13681 gnd.n7539 gnd.n468 240.244
R13682 gnd.n7539 gnd.n464 240.244
R13683 gnd.n7545 gnd.n464 240.244
R13684 gnd.n7545 gnd.n462 240.244
R13685 gnd.n7549 gnd.n462 240.244
R13686 gnd.n7549 gnd.n458 240.244
R13687 gnd.n7555 gnd.n458 240.244
R13688 gnd.n7555 gnd.n456 240.244
R13689 gnd.n7559 gnd.n456 240.244
R13690 gnd.n7559 gnd.n452 240.244
R13691 gnd.n7565 gnd.n452 240.244
R13692 gnd.n7565 gnd.n450 240.244
R13693 gnd.n7569 gnd.n450 240.244
R13694 gnd.n7569 gnd.n446 240.244
R13695 gnd.n7575 gnd.n446 240.244
R13696 gnd.n7575 gnd.n444 240.244
R13697 gnd.n7579 gnd.n444 240.244
R13698 gnd.n7579 gnd.n440 240.244
R13699 gnd.n7585 gnd.n440 240.244
R13700 gnd.n7585 gnd.n438 240.244
R13701 gnd.n7589 gnd.n438 240.244
R13702 gnd.n7589 gnd.n434 240.244
R13703 gnd.n7595 gnd.n434 240.244
R13704 gnd.n7595 gnd.n432 240.244
R13705 gnd.n7599 gnd.n432 240.244
R13706 gnd.n7599 gnd.n428 240.244
R13707 gnd.n7605 gnd.n428 240.244
R13708 gnd.n7605 gnd.n426 240.244
R13709 gnd.n7609 gnd.n426 240.244
R13710 gnd.n7609 gnd.n422 240.244
R13711 gnd.n7615 gnd.n422 240.244
R13712 gnd.n7615 gnd.n420 240.244
R13713 gnd.n7619 gnd.n420 240.244
R13714 gnd.n7619 gnd.n416 240.244
R13715 gnd.n7625 gnd.n416 240.244
R13716 gnd.n7625 gnd.n414 240.244
R13717 gnd.n7629 gnd.n414 240.244
R13718 gnd.n7629 gnd.n410 240.244
R13719 gnd.n7635 gnd.n410 240.244
R13720 gnd.n7635 gnd.n408 240.244
R13721 gnd.n7639 gnd.n408 240.244
R13722 gnd.n7639 gnd.n404 240.244
R13723 gnd.n7645 gnd.n404 240.244
R13724 gnd.n7645 gnd.n402 240.244
R13725 gnd.n7649 gnd.n402 240.244
R13726 gnd.n7649 gnd.n398 240.244
R13727 gnd.n7655 gnd.n398 240.244
R13728 gnd.n7655 gnd.n396 240.244
R13729 gnd.n7659 gnd.n396 240.244
R13730 gnd.n7659 gnd.n392 240.244
R13731 gnd.n7665 gnd.n392 240.244
R13732 gnd.n7665 gnd.n390 240.244
R13733 gnd.n7669 gnd.n390 240.244
R13734 gnd.n7669 gnd.n386 240.244
R13735 gnd.n7675 gnd.n386 240.244
R13736 gnd.n7675 gnd.n384 240.244
R13737 gnd.n7679 gnd.n384 240.244
R13738 gnd.n7679 gnd.n380 240.244
R13739 gnd.n7685 gnd.n380 240.244
R13740 gnd.n7685 gnd.n378 240.244
R13741 gnd.n7689 gnd.n378 240.244
R13742 gnd.n7689 gnd.n374 240.244
R13743 gnd.n7695 gnd.n374 240.244
R13744 gnd.n7695 gnd.n372 240.244
R13745 gnd.n7700 gnd.n372 240.244
R13746 gnd.n7700 gnd.n368 240.244
R13747 gnd.n7707 gnd.n368 240.244
R13748 gnd.n4231 gnd.n4230 240.244
R13749 gnd.n4232 gnd.n4231 240.244
R13750 gnd.n4232 gnd.n4219 240.244
R13751 gnd.n4238 gnd.n4219 240.244
R13752 gnd.n4239 gnd.n4238 240.244
R13753 gnd.n4240 gnd.n4239 240.244
R13754 gnd.n4240 gnd.n4064 240.244
R13755 gnd.n4246 gnd.n4064 240.244
R13756 gnd.n4246 gnd.n4053 240.244
R13757 gnd.n4284 gnd.n4053 240.244
R13758 gnd.n4284 gnd.n4283 240.244
R13759 gnd.n4283 gnd.n4049 240.244
R13760 gnd.n4291 gnd.n4049 240.244
R13761 gnd.n4292 gnd.n4291 240.244
R13762 gnd.n4292 gnd.n4046 240.244
R13763 gnd.n4305 gnd.n4046 240.244
R13764 gnd.n4305 gnd.n4047 240.244
R13765 gnd.n4300 gnd.n4047 240.244
R13766 gnd.n4300 gnd.n4299 240.244
R13767 gnd.n4299 gnd.n4014 240.244
R13768 gnd.n4347 gnd.n4014 240.244
R13769 gnd.n4348 gnd.n4347 240.244
R13770 gnd.n4348 gnd.n4011 240.244
R13771 gnd.n4374 gnd.n4011 240.244
R13772 gnd.n4374 gnd.n4012 240.244
R13773 gnd.n4370 gnd.n4012 240.244
R13774 gnd.n4370 gnd.n4369 240.244
R13775 gnd.n4369 gnd.n4368 240.244
R13776 gnd.n4368 gnd.n4356 240.244
R13777 gnd.n4364 gnd.n4356 240.244
R13778 gnd.n4364 gnd.n3989 240.244
R13779 gnd.n4435 gnd.n3989 240.244
R13780 gnd.n4436 gnd.n4435 240.244
R13781 gnd.n4437 gnd.n4436 240.244
R13782 gnd.n4437 gnd.n3985 240.244
R13783 gnd.n4443 gnd.n3985 240.244
R13784 gnd.n4444 gnd.n4443 240.244
R13785 gnd.n4445 gnd.n4444 240.244
R13786 gnd.n4445 gnd.n3980 240.244
R13787 gnd.n4455 gnd.n3980 240.244
R13788 gnd.n4455 gnd.n3981 240.244
R13789 gnd.n3981 gnd.n3967 240.244
R13790 gnd.n4739 gnd.n3967 240.244
R13791 gnd.n4740 gnd.n4739 240.244
R13792 gnd.n4740 gnd.n3963 240.244
R13793 gnd.n4746 gnd.n3963 240.244
R13794 gnd.n4747 gnd.n4746 240.244
R13795 gnd.n4748 gnd.n4747 240.244
R13796 gnd.n4748 gnd.n3958 240.244
R13797 gnd.n4762 gnd.n3958 240.244
R13798 gnd.n4762 gnd.n3959 240.244
R13799 gnd.n4758 gnd.n3959 240.244
R13800 gnd.n4758 gnd.n4757 240.244
R13801 gnd.n4757 gnd.n3933 240.244
R13802 gnd.n4776 gnd.n3933 240.244
R13803 gnd.n4776 gnd.n3929 240.244
R13804 gnd.n4782 gnd.n3929 240.244
R13805 gnd.n4782 gnd.n3917 240.244
R13806 gnd.n4809 gnd.n3917 240.244
R13807 gnd.n4809 gnd.n3912 240.244
R13808 gnd.n4824 gnd.n3912 240.244
R13809 gnd.n4824 gnd.n3913 240.244
R13810 gnd.n4820 gnd.n3913 240.244
R13811 gnd.n4820 gnd.n4819 240.244
R13812 gnd.n4819 gnd.n2903 240.244
R13813 gnd.n6317 gnd.n2903 240.244
R13814 gnd.n6317 gnd.n2904 240.244
R13815 gnd.n6313 gnd.n2904 240.244
R13816 gnd.n6313 gnd.n2910 240.244
R13817 gnd.n5005 gnd.n2910 240.244
R13818 gnd.n5011 gnd.n5005 240.244
R13819 gnd.n5011 gnd.n3806 240.244
R13820 gnd.n5034 gnd.n3806 240.244
R13821 gnd.n5034 gnd.n3801 240.244
R13822 gnd.n5051 gnd.n3801 240.244
R13823 gnd.n5051 gnd.n3802 240.244
R13824 gnd.n5047 gnd.n3802 240.244
R13825 gnd.n5047 gnd.n5046 240.244
R13826 gnd.n5046 gnd.n5045 240.244
R13827 gnd.n5045 gnd.n3768 240.244
R13828 gnd.n5092 gnd.n3768 240.244
R13829 gnd.n5092 gnd.n3764 240.244
R13830 gnd.n5098 gnd.n3764 240.244
R13831 gnd.n5098 gnd.n3750 240.244
R13832 gnd.n5118 gnd.n3750 240.244
R13833 gnd.n5118 gnd.n3745 240.244
R13834 gnd.n5126 gnd.n3745 240.244
R13835 gnd.n5126 gnd.n3746 240.244
R13836 gnd.n3746 gnd.n3726 240.244
R13837 gnd.n5157 gnd.n3726 240.244
R13838 gnd.n5157 gnd.n3721 240.244
R13839 gnd.n5174 gnd.n3721 240.244
R13840 gnd.n5174 gnd.n3722 240.244
R13841 gnd.n5170 gnd.n3722 240.244
R13842 gnd.n5170 gnd.n5169 240.244
R13843 gnd.n5169 gnd.n5168 240.244
R13844 gnd.n5168 gnd.n3687 240.244
R13845 gnd.n5215 gnd.n3687 240.244
R13846 gnd.n5215 gnd.n3683 240.244
R13847 gnd.n5221 gnd.n3683 240.244
R13848 gnd.n5221 gnd.n3668 240.244
R13849 gnd.n5240 gnd.n3668 240.244
R13850 gnd.n5240 gnd.n3663 240.244
R13851 gnd.n5248 gnd.n3663 240.244
R13852 gnd.n5248 gnd.n3664 240.244
R13853 gnd.n3664 gnd.n3643 240.244
R13854 gnd.n5278 gnd.n3643 240.244
R13855 gnd.n5278 gnd.n3638 240.244
R13856 gnd.n5292 gnd.n3638 240.244
R13857 gnd.n5292 gnd.n3639 240.244
R13858 gnd.n5288 gnd.n3639 240.244
R13859 gnd.n5288 gnd.n5287 240.244
R13860 gnd.n5287 gnd.n3609 240.244
R13861 gnd.n5324 gnd.n3609 240.244
R13862 gnd.n5324 gnd.n3604 240.244
R13863 gnd.n5332 gnd.n3604 240.244
R13864 gnd.n5332 gnd.n3605 240.244
R13865 gnd.n3605 gnd.n3581 240.244
R13866 gnd.n5359 gnd.n3581 240.244
R13867 gnd.n5359 gnd.n3577 240.244
R13868 gnd.n5365 gnd.n3577 240.244
R13869 gnd.n5365 gnd.n3552 240.244
R13870 gnd.n5396 gnd.n3552 240.244
R13871 gnd.n5396 gnd.n3547 240.244
R13872 gnd.n5404 gnd.n3547 240.244
R13873 gnd.n5404 gnd.n3548 240.244
R13874 gnd.n3548 gnd.n3452 240.244
R13875 gnd.n5546 gnd.n3452 240.244
R13876 gnd.n5546 gnd.n3448 240.244
R13877 gnd.n5552 gnd.n3448 240.244
R13878 gnd.n5552 gnd.n3439 240.244
R13879 gnd.n5562 gnd.n3439 240.244
R13880 gnd.n5562 gnd.n3435 240.244
R13881 gnd.n5571 gnd.n3435 240.244
R13882 gnd.n5571 gnd.n3426 240.244
R13883 gnd.n5581 gnd.n3426 240.244
R13884 gnd.n5582 gnd.n5581 240.244
R13885 gnd.n5582 gnd.n3007 240.244
R13886 gnd.n3421 gnd.n3007 240.244
R13887 gnd.n5681 gnd.n3421 240.244
R13888 gnd.n5681 gnd.n3422 240.244
R13889 gnd.n5677 gnd.n3422 240.244
R13890 gnd.n5677 gnd.n5676 240.244
R13891 gnd.n5676 gnd.n5675 240.244
R13892 gnd.n5675 gnd.n5591 240.244
R13893 gnd.n5671 gnd.n5591 240.244
R13894 gnd.n5671 gnd.n5668 240.244
R13895 gnd.n5668 gnd.n5667 240.244
R13896 gnd.n5667 gnd.n5597 240.244
R13897 gnd.n5663 gnd.n5597 240.244
R13898 gnd.n5663 gnd.n5662 240.244
R13899 gnd.n5662 gnd.n5661 240.244
R13900 gnd.n5661 gnd.n5603 240.244
R13901 gnd.n5657 gnd.n5603 240.244
R13902 gnd.n5657 gnd.n5656 240.244
R13903 gnd.n5656 gnd.n5655 240.244
R13904 gnd.n5655 gnd.n5609 240.244
R13905 gnd.n5651 gnd.n5609 240.244
R13906 gnd.n5651 gnd.n5650 240.244
R13907 gnd.n5650 gnd.n5649 240.244
R13908 gnd.n5649 gnd.n5615 240.244
R13909 gnd.n5645 gnd.n5615 240.244
R13910 gnd.n5645 gnd.n5644 240.244
R13911 gnd.n5644 gnd.n5643 240.244
R13912 gnd.n5643 gnd.n5621 240.244
R13913 gnd.n5639 gnd.n5621 240.244
R13914 gnd.n5639 gnd.n5638 240.244
R13915 gnd.n5638 gnd.n5637 240.244
R13916 gnd.n5637 gnd.n5627 240.244
R13917 gnd.n5633 gnd.n5627 240.244
R13918 gnd.n5633 gnd.n3334 240.244
R13919 gnd.n5926 gnd.n3334 240.244
R13920 gnd.n5926 gnd.n3335 240.244
R13921 gnd.n5921 gnd.n3335 240.244
R13922 gnd.n5921 gnd.n3338 240.244
R13923 gnd.n5817 gnd.n3338 240.244
R13924 gnd.n5818 gnd.n5817 240.244
R13925 gnd.n5819 gnd.n5818 240.244
R13926 gnd.n5819 gnd.n5811 240.244
R13927 gnd.n5898 gnd.n5811 240.244
R13928 gnd.n5898 gnd.n5812 240.244
R13929 gnd.n5893 gnd.n5812 240.244
R13930 gnd.n5893 gnd.n5892 240.244
R13931 gnd.n5892 gnd.n5825 240.244
R13932 gnd.n5843 gnd.n5825 240.244
R13933 gnd.n5861 gnd.n5843 240.244
R13934 gnd.n5861 gnd.n5844 240.244
R13935 gnd.n5857 gnd.n5844 240.244
R13936 gnd.n5857 gnd.n5856 240.244
R13937 gnd.n5856 gnd.n361 240.244
R13938 gnd.n7714 gnd.n361 240.244
R13939 gnd.n7714 gnd.n362 240.244
R13940 gnd.n7710 gnd.n362 240.244
R13941 gnd.n7710 gnd.n7709 240.244
R13942 gnd.n7004 gnd.n787 240.244
R13943 gnd.n7000 gnd.n787 240.244
R13944 gnd.n7000 gnd.n792 240.244
R13945 gnd.n6996 gnd.n792 240.244
R13946 gnd.n6996 gnd.n794 240.244
R13947 gnd.n6992 gnd.n794 240.244
R13948 gnd.n6992 gnd.n800 240.244
R13949 gnd.n6988 gnd.n800 240.244
R13950 gnd.n6988 gnd.n802 240.244
R13951 gnd.n6984 gnd.n802 240.244
R13952 gnd.n6984 gnd.n808 240.244
R13953 gnd.n6980 gnd.n808 240.244
R13954 gnd.n6980 gnd.n810 240.244
R13955 gnd.n6976 gnd.n810 240.244
R13956 gnd.n6976 gnd.n816 240.244
R13957 gnd.n6972 gnd.n816 240.244
R13958 gnd.n6972 gnd.n818 240.244
R13959 gnd.n6968 gnd.n818 240.244
R13960 gnd.n6968 gnd.n824 240.244
R13961 gnd.n6964 gnd.n824 240.244
R13962 gnd.n6964 gnd.n826 240.244
R13963 gnd.n6960 gnd.n826 240.244
R13964 gnd.n6960 gnd.n832 240.244
R13965 gnd.n6956 gnd.n832 240.244
R13966 gnd.n6956 gnd.n834 240.244
R13967 gnd.n6952 gnd.n834 240.244
R13968 gnd.n6952 gnd.n840 240.244
R13969 gnd.n6948 gnd.n840 240.244
R13970 gnd.n6948 gnd.n842 240.244
R13971 gnd.n6944 gnd.n842 240.244
R13972 gnd.n6944 gnd.n848 240.244
R13973 gnd.n6940 gnd.n848 240.244
R13974 gnd.n6940 gnd.n850 240.244
R13975 gnd.n6936 gnd.n850 240.244
R13976 gnd.n6936 gnd.n856 240.244
R13977 gnd.n6932 gnd.n856 240.244
R13978 gnd.n6932 gnd.n858 240.244
R13979 gnd.n6928 gnd.n858 240.244
R13980 gnd.n6928 gnd.n864 240.244
R13981 gnd.n6924 gnd.n864 240.244
R13982 gnd.n6924 gnd.n866 240.244
R13983 gnd.n6920 gnd.n866 240.244
R13984 gnd.n6920 gnd.n872 240.244
R13985 gnd.n6916 gnd.n872 240.244
R13986 gnd.n6916 gnd.n874 240.244
R13987 gnd.n6912 gnd.n874 240.244
R13988 gnd.n6912 gnd.n880 240.244
R13989 gnd.n6908 gnd.n880 240.244
R13990 gnd.n6908 gnd.n882 240.244
R13991 gnd.n6904 gnd.n882 240.244
R13992 gnd.n6904 gnd.n888 240.244
R13993 gnd.n6900 gnd.n888 240.244
R13994 gnd.n6900 gnd.n890 240.244
R13995 gnd.n6896 gnd.n890 240.244
R13996 gnd.n6896 gnd.n896 240.244
R13997 gnd.n6892 gnd.n896 240.244
R13998 gnd.n6892 gnd.n898 240.244
R13999 gnd.n6888 gnd.n898 240.244
R14000 gnd.n6888 gnd.n904 240.244
R14001 gnd.n6884 gnd.n904 240.244
R14002 gnd.n6884 gnd.n906 240.244
R14003 gnd.n6880 gnd.n906 240.244
R14004 gnd.n6880 gnd.n912 240.244
R14005 gnd.n6876 gnd.n912 240.244
R14006 gnd.n6876 gnd.n914 240.244
R14007 gnd.n6872 gnd.n914 240.244
R14008 gnd.n6872 gnd.n920 240.244
R14009 gnd.n6868 gnd.n920 240.244
R14010 gnd.n6868 gnd.n922 240.244
R14011 gnd.n6864 gnd.n922 240.244
R14012 gnd.n6864 gnd.n928 240.244
R14013 gnd.n6860 gnd.n928 240.244
R14014 gnd.n6860 gnd.n930 240.244
R14015 gnd.n6856 gnd.n930 240.244
R14016 gnd.n6856 gnd.n936 240.244
R14017 gnd.n6852 gnd.n936 240.244
R14018 gnd.n6852 gnd.n938 240.244
R14019 gnd.n6848 gnd.n938 240.244
R14020 gnd.n6848 gnd.n944 240.244
R14021 gnd.n6844 gnd.n944 240.244
R14022 gnd.n6844 gnd.n946 240.244
R14023 gnd.n6840 gnd.n946 240.244
R14024 gnd.n6840 gnd.n952 240.244
R14025 gnd.n4223 gnd.n952 240.244
R14026 gnd.n4492 gnd.n3928 240.244
R14027 gnd.n4485 gnd.n3928 240.244
R14028 gnd.n4485 gnd.n3919 240.244
R14029 gnd.n3919 gnd.n3908 240.244
R14030 gnd.n4826 gnd.n3908 240.244
R14031 gnd.n4826 gnd.n3904 240.244
R14032 gnd.n4832 gnd.n3904 240.244
R14033 gnd.n4833 gnd.n4832 240.244
R14034 gnd.n4834 gnd.n4833 240.244
R14035 gnd.n4834 gnd.n2900 240.244
R14036 gnd.n4981 gnd.n2900 240.244
R14037 gnd.n4981 gnd.n2911 240.244
R14038 gnd.n4839 gnd.n2911 240.244
R14039 gnd.n4839 gnd.n3819 240.244
R14040 gnd.n3819 gnd.n3817 240.244
R14041 gnd.n3817 gnd.n3814 240.244
R14042 gnd.n3814 gnd.n3807 240.244
R14043 gnd.n4842 gnd.n3807 240.244
R14044 gnd.n4842 gnd.n3800 240.244
R14045 gnd.n4845 gnd.n3800 240.244
R14046 gnd.n4846 gnd.n4845 240.244
R14047 gnd.n4847 gnd.n4846 240.244
R14048 gnd.n4848 gnd.n4847 240.244
R14049 gnd.n4848 gnd.n3775 240.244
R14050 gnd.n3775 gnd.n3769 240.244
R14051 gnd.n4851 gnd.n3769 240.244
R14052 gnd.n4851 gnd.n3762 240.244
R14053 gnd.n4852 gnd.n3762 240.244
R14054 gnd.n4852 gnd.n3751 240.244
R14055 gnd.n4855 gnd.n3751 240.244
R14056 gnd.n4855 gnd.n3744 240.244
R14057 gnd.n4856 gnd.n3744 240.244
R14058 gnd.n4856 gnd.n3735 240.244
R14059 gnd.n3735 gnd.n3727 240.244
R14060 gnd.n4859 gnd.n3727 240.244
R14061 gnd.n4859 gnd.n3720 240.244
R14062 gnd.n4862 gnd.n3720 240.244
R14063 gnd.n4863 gnd.n4862 240.244
R14064 gnd.n4864 gnd.n4863 240.244
R14065 gnd.n4865 gnd.n4864 240.244
R14066 gnd.n4865 gnd.n3696 240.244
R14067 gnd.n3696 gnd.n3689 240.244
R14068 gnd.n4868 gnd.n3689 240.244
R14069 gnd.n4868 gnd.n3681 240.244
R14070 gnd.n4871 gnd.n3681 240.244
R14071 gnd.n4871 gnd.n3669 240.244
R14072 gnd.n4872 gnd.n3669 240.244
R14073 gnd.n4872 gnd.n3662 240.244
R14074 gnd.n4875 gnd.n3662 240.244
R14075 gnd.n4875 gnd.n3652 240.244
R14076 gnd.n3652 gnd.n3644 240.244
R14077 gnd.n4877 gnd.n3644 240.244
R14078 gnd.n4877 gnd.n3636 240.244
R14079 gnd.n4880 gnd.n3636 240.244
R14080 gnd.n4881 gnd.n4880 240.244
R14081 gnd.n4884 gnd.n4881 240.244
R14082 gnd.n4885 gnd.n4884 240.244
R14083 gnd.n4885 gnd.n3612 240.244
R14084 gnd.n4886 gnd.n3612 240.244
R14085 gnd.n4886 gnd.n3602 240.244
R14086 gnd.n4889 gnd.n3602 240.244
R14087 gnd.n4890 gnd.n4889 240.244
R14088 gnd.n4890 gnd.n3583 240.244
R14089 gnd.n4891 gnd.n3583 240.244
R14090 gnd.n4891 gnd.n3574 240.244
R14091 gnd.n4894 gnd.n3574 240.244
R14092 gnd.n4894 gnd.n3554 240.244
R14093 gnd.n3554 gnd.n3543 240.244
R14094 gnd.n5406 gnd.n3543 240.244
R14095 gnd.n5406 gnd.n3538 240.244
R14096 gnd.n5413 gnd.n3538 240.244
R14097 gnd.n5413 gnd.n3453 240.244
R14098 gnd.n3453 gnd.n3444 240.244
R14099 gnd.n5554 gnd.n3444 240.244
R14100 gnd.n5554 gnd.n3440 240.244
R14101 gnd.n5560 gnd.n3440 240.244
R14102 gnd.n5560 gnd.n3432 240.244
R14103 gnd.n5573 gnd.n3432 240.244
R14104 gnd.n5573 gnd.n3428 240.244
R14105 gnd.n5579 gnd.n3428 240.244
R14106 gnd.n5579 gnd.n3009 240.244
R14107 gnd.n6201 gnd.n3009 240.244
R14108 gnd.n4497 gnd.n4496 240.244
R14109 gnd.n4480 gnd.n4479 240.244
R14110 gnd.n4505 gnd.n4504 240.244
R14111 gnd.n4507 gnd.n4506 240.244
R14112 gnd.n4514 gnd.n4513 240.244
R14113 gnd.n4516 gnd.n4515 240.244
R14114 gnd.n4526 gnd.n4525 240.244
R14115 gnd.n4534 gnd.n4533 240.244
R14116 gnd.n4536 gnd.n4535 240.244
R14117 gnd.n4546 gnd.n4545 240.244
R14118 gnd.n4554 gnd.n4553 240.244
R14119 gnd.n4556 gnd.n4555 240.244
R14120 gnd.n4568 gnd.n4567 240.244
R14121 gnd.n4773 gnd.n3949 240.244
R14122 gnd.n4784 gnd.n3926 240.244
R14123 gnd.n4784 gnd.n3920 240.244
R14124 gnd.n4807 gnd.n3920 240.244
R14125 gnd.n4807 gnd.n3921 240.244
R14126 gnd.n3921 gnd.n3911 240.244
R14127 gnd.n4789 gnd.n3911 240.244
R14128 gnd.n4790 gnd.n4789 240.244
R14129 gnd.n4793 gnd.n4790 240.244
R14130 gnd.n4794 gnd.n4793 240.244
R14131 gnd.n4794 gnd.n2902 240.244
R14132 gnd.n2913 gnd.n2902 240.244
R14133 gnd.n6311 gnd.n2913 240.244
R14134 gnd.n6311 gnd.n2914 240.244
R14135 gnd.n2919 gnd.n2914 240.244
R14136 gnd.n2920 gnd.n2919 240.244
R14137 gnd.n2921 gnd.n2920 240.244
R14138 gnd.n5032 gnd.n2921 240.244
R14139 gnd.n5032 gnd.n2924 240.244
R14140 gnd.n2925 gnd.n2924 240.244
R14141 gnd.n2926 gnd.n2925 240.244
R14142 gnd.n3787 gnd.n2926 240.244
R14143 gnd.n3787 gnd.n2929 240.244
R14144 gnd.n2930 gnd.n2929 240.244
R14145 gnd.n2931 gnd.n2930 240.244
R14146 gnd.n5090 gnd.n2931 240.244
R14147 gnd.n5090 gnd.n2934 240.244
R14148 gnd.n2935 gnd.n2934 240.244
R14149 gnd.n2936 gnd.n2935 240.244
R14150 gnd.n5116 gnd.n2936 240.244
R14151 gnd.n5116 gnd.n2939 240.244
R14152 gnd.n2940 gnd.n2939 240.244
R14153 gnd.n2941 gnd.n2940 240.244
R14154 gnd.n5147 gnd.n2941 240.244
R14155 gnd.n5147 gnd.n2944 240.244
R14156 gnd.n2945 gnd.n2944 240.244
R14157 gnd.n2946 gnd.n2945 240.244
R14158 gnd.n3713 gnd.n2946 240.244
R14159 gnd.n3713 gnd.n2949 240.244
R14160 gnd.n2950 gnd.n2949 240.244
R14161 gnd.n2951 gnd.n2950 240.244
R14162 gnd.n3697 gnd.n2951 240.244
R14163 gnd.n3697 gnd.n2954 240.244
R14164 gnd.n2955 gnd.n2954 240.244
R14165 gnd.n2956 gnd.n2955 240.244
R14166 gnd.n3673 gnd.n2956 240.244
R14167 gnd.n3673 gnd.n2959 240.244
R14168 gnd.n2960 gnd.n2959 240.244
R14169 gnd.n2961 gnd.n2960 240.244
R14170 gnd.n3655 gnd.n2961 240.244
R14171 gnd.n3655 gnd.n2964 240.244
R14172 gnd.n2965 gnd.n2964 240.244
R14173 gnd.n2966 gnd.n2965 240.244
R14174 gnd.n3637 gnd.n2966 240.244
R14175 gnd.n3637 gnd.n2969 240.244
R14176 gnd.n2970 gnd.n2969 240.244
R14177 gnd.n2971 gnd.n2970 240.244
R14178 gnd.n3619 gnd.n2971 240.244
R14179 gnd.n3619 gnd.n2974 240.244
R14180 gnd.n2975 gnd.n2974 240.244
R14181 gnd.n2976 gnd.n2975 240.244
R14182 gnd.n3595 gnd.n2976 240.244
R14183 gnd.n3595 gnd.n2979 240.244
R14184 gnd.n2980 gnd.n2979 240.244
R14185 gnd.n2981 gnd.n2980 240.244
R14186 gnd.n3576 gnd.n2981 240.244
R14187 gnd.n3576 gnd.n2984 240.244
R14188 gnd.n2985 gnd.n2984 240.244
R14189 gnd.n2986 gnd.n2985 240.244
R14190 gnd.n3546 gnd.n2986 240.244
R14191 gnd.n3546 gnd.n2989 240.244
R14192 gnd.n2990 gnd.n2989 240.244
R14193 gnd.n2991 gnd.n2990 240.244
R14194 gnd.n3455 gnd.n2991 240.244
R14195 gnd.n3455 gnd.n2994 240.244
R14196 gnd.n2995 gnd.n2994 240.244
R14197 gnd.n2996 gnd.n2995 240.244
R14198 gnd.n3433 gnd.n2996 240.244
R14199 gnd.n3433 gnd.n2999 240.244
R14200 gnd.n3000 gnd.n2999 240.244
R14201 gnd.n3001 gnd.n3000 240.244
R14202 gnd.n3004 gnd.n3001 240.244
R14203 gnd.n6203 gnd.n3004 240.244
R14204 gnd.n3015 gnd.n3014 240.244
R14205 gnd.n3399 gnd.n3018 240.244
R14206 gnd.n3020 gnd.n3019 240.244
R14207 gnd.n3402 gnd.n3024 240.244
R14208 gnd.n3405 gnd.n3025 240.244
R14209 gnd.n3034 gnd.n3033 240.244
R14210 gnd.n3407 gnd.n3041 240.244
R14211 gnd.n3410 gnd.n3042 240.244
R14212 gnd.n3050 gnd.n3049 240.244
R14213 gnd.n3412 gnd.n3057 240.244
R14214 gnd.n3415 gnd.n3058 240.244
R14215 gnd.n3066 gnd.n3065 240.244
R14216 gnd.n3418 gnd.n3397 240.244
R14217 gnd.n5684 gnd.n3005 240.244
R14218 gnd.n2881 gnd.n2880 240.132
R14219 gnd.n3472 gnd.n3471 240.132
R14220 gnd.n7007 gnd.n7006 225.874
R14221 gnd.n7007 gnd.n780 225.874
R14222 gnd.n7015 gnd.n780 225.874
R14223 gnd.n7016 gnd.n7015 225.874
R14224 gnd.n7017 gnd.n7016 225.874
R14225 gnd.n7017 gnd.n774 225.874
R14226 gnd.n7025 gnd.n774 225.874
R14227 gnd.n7026 gnd.n7025 225.874
R14228 gnd.n7027 gnd.n7026 225.874
R14229 gnd.n7027 gnd.n768 225.874
R14230 gnd.n7035 gnd.n768 225.874
R14231 gnd.n7036 gnd.n7035 225.874
R14232 gnd.n7037 gnd.n7036 225.874
R14233 gnd.n7037 gnd.n762 225.874
R14234 gnd.n7045 gnd.n762 225.874
R14235 gnd.n7046 gnd.n7045 225.874
R14236 gnd.n7047 gnd.n7046 225.874
R14237 gnd.n7047 gnd.n756 225.874
R14238 gnd.n7055 gnd.n756 225.874
R14239 gnd.n7056 gnd.n7055 225.874
R14240 gnd.n7057 gnd.n7056 225.874
R14241 gnd.n7057 gnd.n750 225.874
R14242 gnd.n7065 gnd.n750 225.874
R14243 gnd.n7066 gnd.n7065 225.874
R14244 gnd.n7067 gnd.n7066 225.874
R14245 gnd.n7067 gnd.n744 225.874
R14246 gnd.n7075 gnd.n744 225.874
R14247 gnd.n7076 gnd.n7075 225.874
R14248 gnd.n7077 gnd.n7076 225.874
R14249 gnd.n7077 gnd.n738 225.874
R14250 gnd.n7085 gnd.n738 225.874
R14251 gnd.n7086 gnd.n7085 225.874
R14252 gnd.n7087 gnd.n7086 225.874
R14253 gnd.n7087 gnd.n732 225.874
R14254 gnd.n7095 gnd.n732 225.874
R14255 gnd.n7096 gnd.n7095 225.874
R14256 gnd.n7097 gnd.n7096 225.874
R14257 gnd.n7097 gnd.n726 225.874
R14258 gnd.n7105 gnd.n726 225.874
R14259 gnd.n7106 gnd.n7105 225.874
R14260 gnd.n7107 gnd.n7106 225.874
R14261 gnd.n7107 gnd.n720 225.874
R14262 gnd.n7115 gnd.n720 225.874
R14263 gnd.n7116 gnd.n7115 225.874
R14264 gnd.n7117 gnd.n7116 225.874
R14265 gnd.n7117 gnd.n714 225.874
R14266 gnd.n7125 gnd.n714 225.874
R14267 gnd.n7126 gnd.n7125 225.874
R14268 gnd.n7127 gnd.n7126 225.874
R14269 gnd.n7127 gnd.n708 225.874
R14270 gnd.n7135 gnd.n708 225.874
R14271 gnd.n7136 gnd.n7135 225.874
R14272 gnd.n7137 gnd.n7136 225.874
R14273 gnd.n7137 gnd.n702 225.874
R14274 gnd.n7145 gnd.n702 225.874
R14275 gnd.n7146 gnd.n7145 225.874
R14276 gnd.n7147 gnd.n7146 225.874
R14277 gnd.n7147 gnd.n696 225.874
R14278 gnd.n7155 gnd.n696 225.874
R14279 gnd.n7156 gnd.n7155 225.874
R14280 gnd.n7157 gnd.n7156 225.874
R14281 gnd.n7157 gnd.n690 225.874
R14282 gnd.n7165 gnd.n690 225.874
R14283 gnd.n7166 gnd.n7165 225.874
R14284 gnd.n7167 gnd.n7166 225.874
R14285 gnd.n7167 gnd.n684 225.874
R14286 gnd.n7175 gnd.n684 225.874
R14287 gnd.n7176 gnd.n7175 225.874
R14288 gnd.n7177 gnd.n7176 225.874
R14289 gnd.n7177 gnd.n678 225.874
R14290 gnd.n7185 gnd.n678 225.874
R14291 gnd.n7186 gnd.n7185 225.874
R14292 gnd.n7187 gnd.n7186 225.874
R14293 gnd.n7187 gnd.n672 225.874
R14294 gnd.n7195 gnd.n672 225.874
R14295 gnd.n7196 gnd.n7195 225.874
R14296 gnd.n7197 gnd.n7196 225.874
R14297 gnd.n7197 gnd.n666 225.874
R14298 gnd.n7205 gnd.n666 225.874
R14299 gnd.n7206 gnd.n7205 225.874
R14300 gnd.n7207 gnd.n7206 225.874
R14301 gnd.n7207 gnd.n660 225.874
R14302 gnd.n7215 gnd.n660 225.874
R14303 gnd.n7216 gnd.n7215 225.874
R14304 gnd.n7217 gnd.n7216 225.874
R14305 gnd.n7217 gnd.n654 225.874
R14306 gnd.n7225 gnd.n654 225.874
R14307 gnd.n7226 gnd.n7225 225.874
R14308 gnd.n7227 gnd.n7226 225.874
R14309 gnd.n7227 gnd.n648 225.874
R14310 gnd.n7235 gnd.n648 225.874
R14311 gnd.n7236 gnd.n7235 225.874
R14312 gnd.n7237 gnd.n7236 225.874
R14313 gnd.n7237 gnd.n642 225.874
R14314 gnd.n7245 gnd.n642 225.874
R14315 gnd.n7246 gnd.n7245 225.874
R14316 gnd.n7247 gnd.n7246 225.874
R14317 gnd.n7247 gnd.n636 225.874
R14318 gnd.n7255 gnd.n636 225.874
R14319 gnd.n7256 gnd.n7255 225.874
R14320 gnd.n7257 gnd.n7256 225.874
R14321 gnd.n7257 gnd.n630 225.874
R14322 gnd.n7265 gnd.n630 225.874
R14323 gnd.n7266 gnd.n7265 225.874
R14324 gnd.n7267 gnd.n7266 225.874
R14325 gnd.n7267 gnd.n624 225.874
R14326 gnd.n7275 gnd.n624 225.874
R14327 gnd.n7276 gnd.n7275 225.874
R14328 gnd.n7277 gnd.n7276 225.874
R14329 gnd.n7277 gnd.n618 225.874
R14330 gnd.n7285 gnd.n618 225.874
R14331 gnd.n7286 gnd.n7285 225.874
R14332 gnd.n7287 gnd.n7286 225.874
R14333 gnd.n7287 gnd.n612 225.874
R14334 gnd.n7295 gnd.n612 225.874
R14335 gnd.n7296 gnd.n7295 225.874
R14336 gnd.n7297 gnd.n7296 225.874
R14337 gnd.n7297 gnd.n606 225.874
R14338 gnd.n7305 gnd.n606 225.874
R14339 gnd.n7306 gnd.n7305 225.874
R14340 gnd.n7307 gnd.n7306 225.874
R14341 gnd.n7307 gnd.n600 225.874
R14342 gnd.n7315 gnd.n600 225.874
R14343 gnd.n7316 gnd.n7315 225.874
R14344 gnd.n7317 gnd.n7316 225.874
R14345 gnd.n7317 gnd.n594 225.874
R14346 gnd.n7325 gnd.n594 225.874
R14347 gnd.n7326 gnd.n7325 225.874
R14348 gnd.n7327 gnd.n7326 225.874
R14349 gnd.n7327 gnd.n588 225.874
R14350 gnd.n7335 gnd.n588 225.874
R14351 gnd.n7336 gnd.n7335 225.874
R14352 gnd.n7337 gnd.n7336 225.874
R14353 gnd.n7337 gnd.n582 225.874
R14354 gnd.n7345 gnd.n582 225.874
R14355 gnd.n7346 gnd.n7345 225.874
R14356 gnd.n7347 gnd.n7346 225.874
R14357 gnd.n7347 gnd.n576 225.874
R14358 gnd.n7355 gnd.n576 225.874
R14359 gnd.n7356 gnd.n7355 225.874
R14360 gnd.n7357 gnd.n7356 225.874
R14361 gnd.n7357 gnd.n570 225.874
R14362 gnd.n7365 gnd.n570 225.874
R14363 gnd.n7366 gnd.n7365 225.874
R14364 gnd.n7367 gnd.n7366 225.874
R14365 gnd.n7367 gnd.n564 225.874
R14366 gnd.n7375 gnd.n564 225.874
R14367 gnd.n7376 gnd.n7375 225.874
R14368 gnd.n7377 gnd.n7376 225.874
R14369 gnd.n7377 gnd.n558 225.874
R14370 gnd.n7385 gnd.n558 225.874
R14371 gnd.n7386 gnd.n7385 225.874
R14372 gnd.n7387 gnd.n7386 225.874
R14373 gnd.n7387 gnd.n552 225.874
R14374 gnd.n7395 gnd.n552 225.874
R14375 gnd.n7396 gnd.n7395 225.874
R14376 gnd.n7397 gnd.n7396 225.874
R14377 gnd.n7397 gnd.n546 225.874
R14378 gnd.n7405 gnd.n546 225.874
R14379 gnd.n7406 gnd.n7405 225.874
R14380 gnd.n7407 gnd.n7406 225.874
R14381 gnd.n7407 gnd.n540 225.874
R14382 gnd.n7415 gnd.n540 225.874
R14383 gnd.n7416 gnd.n7415 225.874
R14384 gnd.n7417 gnd.n7416 225.874
R14385 gnd.n7417 gnd.n534 225.874
R14386 gnd.n7425 gnd.n534 225.874
R14387 gnd.n7426 gnd.n7425 225.874
R14388 gnd.n7427 gnd.n7426 225.874
R14389 gnd.n7427 gnd.n528 225.874
R14390 gnd.n7435 gnd.n528 225.874
R14391 gnd.n7436 gnd.n7435 225.874
R14392 gnd.n7437 gnd.n7436 225.874
R14393 gnd.n7437 gnd.n522 225.874
R14394 gnd.n7445 gnd.n522 225.874
R14395 gnd.n7446 gnd.n7445 225.874
R14396 gnd.n7447 gnd.n7446 225.874
R14397 gnd.n7447 gnd.n516 225.874
R14398 gnd.n7455 gnd.n516 225.874
R14399 gnd.n7456 gnd.n7455 225.874
R14400 gnd.n7457 gnd.n7456 225.874
R14401 gnd.n7457 gnd.n510 225.874
R14402 gnd.n7465 gnd.n510 225.874
R14403 gnd.n7466 gnd.n7465 225.874
R14404 gnd.n7467 gnd.n7466 225.874
R14405 gnd.n7467 gnd.n504 225.874
R14406 gnd.n7475 gnd.n504 225.874
R14407 gnd.n7476 gnd.n7475 225.874
R14408 gnd.n7477 gnd.n7476 225.874
R14409 gnd.n7477 gnd.n498 225.874
R14410 gnd.n7486 gnd.n498 225.874
R14411 gnd.n7487 gnd.n7486 225.874
R14412 gnd.n7488 gnd.n7487 225.874
R14413 gnd.n7488 gnd.n493 225.874
R14414 gnd.n1569 gnd.t224 224.174
R14415 gnd.n1033 gnd.t339 224.174
R14416 gnd.n3150 gnd.n3087 199.319
R14417 gnd.n3150 gnd.n3088 199.319
R14418 gnd.n2833 gnd.n2793 199.319
R14419 gnd.n2833 gnd.n2792 199.319
R14420 gnd.n2882 gnd.n2879 186.49
R14421 gnd.n3473 gnd.n3470 186.49
R14422 gnd.n2325 gnd.n2324 185
R14423 gnd.n2323 gnd.n2322 185
R14424 gnd.n2302 gnd.n2301 185
R14425 gnd.n2317 gnd.n2316 185
R14426 gnd.n2315 gnd.n2314 185
R14427 gnd.n2306 gnd.n2305 185
R14428 gnd.n2309 gnd.n2308 185
R14429 gnd.n2293 gnd.n2292 185
R14430 gnd.n2291 gnd.n2290 185
R14431 gnd.n2270 gnd.n2269 185
R14432 gnd.n2285 gnd.n2284 185
R14433 gnd.n2283 gnd.n2282 185
R14434 gnd.n2274 gnd.n2273 185
R14435 gnd.n2277 gnd.n2276 185
R14436 gnd.n2261 gnd.n2260 185
R14437 gnd.n2259 gnd.n2258 185
R14438 gnd.n2238 gnd.n2237 185
R14439 gnd.n2253 gnd.n2252 185
R14440 gnd.n2251 gnd.n2250 185
R14441 gnd.n2242 gnd.n2241 185
R14442 gnd.n2245 gnd.n2244 185
R14443 gnd.n2230 gnd.n2229 185
R14444 gnd.n2228 gnd.n2227 185
R14445 gnd.n2207 gnd.n2206 185
R14446 gnd.n2222 gnd.n2221 185
R14447 gnd.n2220 gnd.n2219 185
R14448 gnd.n2211 gnd.n2210 185
R14449 gnd.n2214 gnd.n2213 185
R14450 gnd.n2198 gnd.n2197 185
R14451 gnd.n2196 gnd.n2195 185
R14452 gnd.n2175 gnd.n2174 185
R14453 gnd.n2190 gnd.n2189 185
R14454 gnd.n2188 gnd.n2187 185
R14455 gnd.n2179 gnd.n2178 185
R14456 gnd.n2182 gnd.n2181 185
R14457 gnd.n2166 gnd.n2165 185
R14458 gnd.n2164 gnd.n2163 185
R14459 gnd.n2143 gnd.n2142 185
R14460 gnd.n2158 gnd.n2157 185
R14461 gnd.n2156 gnd.n2155 185
R14462 gnd.n2147 gnd.n2146 185
R14463 gnd.n2150 gnd.n2149 185
R14464 gnd.n2134 gnd.n2133 185
R14465 gnd.n2132 gnd.n2131 185
R14466 gnd.n2111 gnd.n2110 185
R14467 gnd.n2126 gnd.n2125 185
R14468 gnd.n2124 gnd.n2123 185
R14469 gnd.n2115 gnd.n2114 185
R14470 gnd.n2118 gnd.n2117 185
R14471 gnd.n2103 gnd.n2102 185
R14472 gnd.n2101 gnd.n2100 185
R14473 gnd.n2080 gnd.n2079 185
R14474 gnd.n2095 gnd.n2094 185
R14475 gnd.n2093 gnd.n2092 185
R14476 gnd.n2084 gnd.n2083 185
R14477 gnd.n2087 gnd.n2086 185
R14478 gnd.n1570 gnd.t223 178.987
R14479 gnd.n1034 gnd.t340 178.987
R14480 gnd.n1 gnd.t367 170.774
R14481 gnd.n7 gnd.t345 170.103
R14482 gnd.n6 gnd.t393 170.103
R14483 gnd.n5 gnd.t403 170.103
R14484 gnd.n4 gnd.t357 170.103
R14485 gnd.n3 gnd.t385 170.103
R14486 gnd.n2 gnd.t369 170.103
R14487 gnd.n1 gnd.t350 170.103
R14488 gnd.n5536 gnd.n3482 163.367
R14489 gnd.n5532 gnd.n5531 163.367
R14490 gnd.n5529 gnd.n3485 163.367
R14491 gnd.n5525 gnd.n5524 163.367
R14492 gnd.n5522 gnd.n3488 163.367
R14493 gnd.n5518 gnd.n5517 163.367
R14494 gnd.n5515 gnd.n3491 163.367
R14495 gnd.n5511 gnd.n5510 163.367
R14496 gnd.n5508 gnd.n3494 163.367
R14497 gnd.n5504 gnd.n5503 163.367
R14498 gnd.n5501 gnd.n3497 163.367
R14499 gnd.n5497 gnd.n5496 163.367
R14500 gnd.n5494 gnd.n3500 163.367
R14501 gnd.n5490 gnd.n5489 163.367
R14502 gnd.n5487 gnd.n3503 163.367
R14503 gnd.n5483 gnd.n5482 163.367
R14504 gnd.n5479 gnd.n5478 163.367
R14505 gnd.n5476 gnd.n3509 163.367
R14506 gnd.n5471 gnd.n5470 163.367
R14507 gnd.n5468 gnd.n3514 163.367
R14508 gnd.n5464 gnd.n5463 163.367
R14509 gnd.n5461 gnd.n3517 163.367
R14510 gnd.n5457 gnd.n5456 163.367
R14511 gnd.n5454 gnd.n3520 163.367
R14512 gnd.n5450 gnd.n5449 163.367
R14513 gnd.n5447 gnd.n3523 163.367
R14514 gnd.n5443 gnd.n5442 163.367
R14515 gnd.n5440 gnd.n3526 163.367
R14516 gnd.n5436 gnd.n5435 163.367
R14517 gnd.n5433 gnd.n3529 163.367
R14518 gnd.n5429 gnd.n5428 163.367
R14519 gnd.n5426 gnd.n3532 163.367
R14520 gnd.n3893 gnd.n2898 163.367
R14521 gnd.n2899 gnd.n2898 163.367
R14522 gnd.n3898 gnd.n2899 163.367
R14523 gnd.n3899 gnd.n3898 163.367
R14524 gnd.n4991 gnd.n3899 163.367
R14525 gnd.n4991 gnd.n3824 163.367
R14526 gnd.n4996 gnd.n3824 163.367
R14527 gnd.n4996 gnd.n3825 163.367
R14528 gnd.n3825 gnd.n3816 163.367
R14529 gnd.n5014 gnd.n3816 163.367
R14530 gnd.n5014 gnd.n3813 163.367
R14531 gnd.n5022 gnd.n3813 163.367
R14532 gnd.n5022 gnd.n3808 163.367
R14533 gnd.n5018 gnd.n3808 163.367
R14534 gnd.n5018 gnd.n3799 163.367
R14535 gnd.n3799 gnd.n3791 163.367
R14536 gnd.n5059 gnd.n3791 163.367
R14537 gnd.n5059 gnd.n3789 163.367
R14538 gnd.n5063 gnd.n3789 163.367
R14539 gnd.n5063 gnd.n3780 163.367
R14540 gnd.n5072 gnd.n3780 163.367
R14541 gnd.n5072 gnd.n3777 163.367
R14542 gnd.n5082 gnd.n3777 163.367
R14543 gnd.n5082 gnd.n3778 163.367
R14544 gnd.n3778 gnd.n3770 163.367
R14545 gnd.n5077 gnd.n3770 163.367
R14546 gnd.n5077 gnd.n3761 163.367
R14547 gnd.n3761 gnd.n3754 163.367
R14548 gnd.n5108 gnd.n3754 163.367
R14549 gnd.n5108 gnd.n3752 163.367
R14550 gnd.n5114 gnd.n3752 163.367
R14551 gnd.n5114 gnd.n3743 163.367
R14552 gnd.n3743 gnd.n3737 163.367
R14553 gnd.n5136 gnd.n3737 163.367
R14554 gnd.n5137 gnd.n5136 163.367
R14555 gnd.n5137 gnd.n3734 163.367
R14556 gnd.n5145 gnd.n3734 163.367
R14557 gnd.n5145 gnd.n3728 163.367
R14558 gnd.n5141 gnd.n3728 163.367
R14559 gnd.n5141 gnd.n3719 163.367
R14560 gnd.n3719 gnd.n3710 163.367
R14561 gnd.n5183 gnd.n3710 163.367
R14562 gnd.n5183 gnd.n3708 163.367
R14563 gnd.n5187 gnd.n3708 163.367
R14564 gnd.n5187 gnd.n3701 163.367
R14565 gnd.n5196 gnd.n3701 163.367
R14566 gnd.n5196 gnd.n3698 163.367
R14567 gnd.n5206 gnd.n3698 163.367
R14568 gnd.n5206 gnd.n3699 163.367
R14569 gnd.n3699 gnd.n3690 163.367
R14570 gnd.n5201 gnd.n3690 163.367
R14571 gnd.n5201 gnd.n3680 163.367
R14572 gnd.n3680 gnd.n3672 163.367
R14573 gnd.n5231 gnd.n3672 163.367
R14574 gnd.n5231 gnd.n3670 163.367
R14575 gnd.n5237 gnd.n3670 163.367
R14576 gnd.n5237 gnd.n3661 163.367
R14577 gnd.n3661 gnd.n3654 163.367
R14578 gnd.n5258 gnd.n3654 163.367
R14579 gnd.n5259 gnd.n5258 163.367
R14580 gnd.n5259 gnd.n3651 163.367
R14581 gnd.n5267 gnd.n3651 163.367
R14582 gnd.n5267 gnd.n3645 163.367
R14583 gnd.n5263 gnd.n3645 163.367
R14584 gnd.n5263 gnd.n3635 163.367
R14585 gnd.n3635 gnd.n3628 163.367
R14586 gnd.n5301 gnd.n3628 163.367
R14587 gnd.n5301 gnd.n3626 163.367
R14588 gnd.n5305 gnd.n3626 163.367
R14589 gnd.n5305 gnd.n3617 163.367
R14590 gnd.n5316 gnd.n3617 163.367
R14591 gnd.n5316 gnd.n3613 163.367
R14592 gnd.n5322 gnd.n3613 163.367
R14593 gnd.n5322 gnd.n3615 163.367
R14594 gnd.n3615 gnd.n3601 163.367
R14595 gnd.n3601 gnd.n3593 163.367
R14596 gnd.n5341 gnd.n3593 163.367
R14597 gnd.n5341 gnd.n3590 163.367
R14598 gnd.n5351 gnd.n3590 163.367
R14599 gnd.n5351 gnd.n3591 163.367
R14600 gnd.n3591 gnd.n3584 163.367
R14601 gnd.n5346 gnd.n3584 163.367
R14602 gnd.n5346 gnd.n3573 163.367
R14603 gnd.n3573 gnd.n3567 163.367
R14604 gnd.n5374 gnd.n3567 163.367
R14605 gnd.n5375 gnd.n5374 163.367
R14606 gnd.n5375 gnd.n3555 163.367
R14607 gnd.n5380 gnd.n3555 163.367
R14608 gnd.n5381 gnd.n5380 163.367
R14609 gnd.n5381 gnd.n3565 163.367
R14610 gnd.n5385 gnd.n3565 163.367
R14611 gnd.n5385 gnd.n3536 163.367
R14612 gnd.n5416 gnd.n3536 163.367
R14613 gnd.n5416 gnd.n3454 163.367
R14614 gnd.n5420 gnd.n3454 163.367
R14615 gnd.n5421 gnd.n5420 163.367
R14616 gnd.n2873 gnd.n2872 163.367
R14617 gnd.n6383 gnd.n2872 163.367
R14618 gnd.n6381 gnd.n6380 163.367
R14619 gnd.n6377 gnd.n6376 163.367
R14620 gnd.n6373 gnd.n6372 163.367
R14621 gnd.n6369 gnd.n6368 163.367
R14622 gnd.n6365 gnd.n6364 163.367
R14623 gnd.n6361 gnd.n6360 163.367
R14624 gnd.n6357 gnd.n6356 163.367
R14625 gnd.n6353 gnd.n6352 163.367
R14626 gnd.n6349 gnd.n6348 163.367
R14627 gnd.n6345 gnd.n6344 163.367
R14628 gnd.n6341 gnd.n6340 163.367
R14629 gnd.n6337 gnd.n6336 163.367
R14630 gnd.n6333 gnd.n6332 163.367
R14631 gnd.n6329 gnd.n6328 163.367
R14632 gnd.n6392 gnd.n2838 163.367
R14633 gnd.n3831 gnd.n3830 163.367
R14634 gnd.n3836 gnd.n3835 163.367
R14635 gnd.n3840 gnd.n3839 163.367
R14636 gnd.n3844 gnd.n3843 163.367
R14637 gnd.n3848 gnd.n3847 163.367
R14638 gnd.n3852 gnd.n3851 163.367
R14639 gnd.n3856 gnd.n3855 163.367
R14640 gnd.n3860 gnd.n3859 163.367
R14641 gnd.n3864 gnd.n3863 163.367
R14642 gnd.n3868 gnd.n3867 163.367
R14643 gnd.n3872 gnd.n3871 163.367
R14644 gnd.n3876 gnd.n3875 163.367
R14645 gnd.n3880 gnd.n3879 163.367
R14646 gnd.n3884 gnd.n3883 163.367
R14647 gnd.n3888 gnd.n3887 163.367
R14648 gnd.n6321 gnd.n2874 163.367
R14649 gnd.n6321 gnd.n2896 163.367
R14650 gnd.n4985 gnd.n2896 163.367
R14651 gnd.n4985 gnd.n4984 163.367
R14652 gnd.n4989 gnd.n4984 163.367
R14653 gnd.n4989 gnd.n3822 163.367
R14654 gnd.n4998 gnd.n3822 163.367
R14655 gnd.n4998 gnd.n3820 163.367
R14656 gnd.n5002 gnd.n3820 163.367
R14657 gnd.n5002 gnd.n3812 163.367
R14658 gnd.n5026 gnd.n3812 163.367
R14659 gnd.n5026 gnd.n3810 163.367
R14660 gnd.n5030 gnd.n3810 163.367
R14661 gnd.n5030 gnd.n3797 163.367
R14662 gnd.n5053 gnd.n3797 163.367
R14663 gnd.n5053 gnd.n3795 163.367
R14664 gnd.n5057 gnd.n3795 163.367
R14665 gnd.n5057 gnd.n3786 163.367
R14666 gnd.n5066 gnd.n3786 163.367
R14667 gnd.n5066 gnd.n3784 163.367
R14668 gnd.n5070 gnd.n3784 163.367
R14669 gnd.n5070 gnd.n3774 163.367
R14670 gnd.n5084 gnd.n3774 163.367
R14671 gnd.n5084 gnd.n3772 163.367
R14672 gnd.n5088 gnd.n3772 163.367
R14673 gnd.n5088 gnd.n3760 163.367
R14674 gnd.n5101 gnd.n3760 163.367
R14675 gnd.n5101 gnd.n3757 163.367
R14676 gnd.n5106 gnd.n3757 163.367
R14677 gnd.n5106 gnd.n3758 163.367
R14678 gnd.n3758 gnd.n3741 163.367
R14679 gnd.n5130 gnd.n3741 163.367
R14680 gnd.n5130 gnd.n3739 163.367
R14681 gnd.n5134 gnd.n3739 163.367
R14682 gnd.n5134 gnd.n3732 163.367
R14683 gnd.n5150 gnd.n3732 163.367
R14684 gnd.n5150 gnd.n3730 163.367
R14685 gnd.n5154 gnd.n3730 163.367
R14686 gnd.n5154 gnd.n3717 163.367
R14687 gnd.n5177 gnd.n3717 163.367
R14688 gnd.n5177 gnd.n3715 163.367
R14689 gnd.n5181 gnd.n3715 163.367
R14690 gnd.n5181 gnd.n3706 163.367
R14691 gnd.n5190 gnd.n3706 163.367
R14692 gnd.n5190 gnd.n3704 163.367
R14693 gnd.n5194 gnd.n3704 163.367
R14694 gnd.n5194 gnd.n3694 163.367
R14695 gnd.n5208 gnd.n3694 163.367
R14696 gnd.n5208 gnd.n3692 163.367
R14697 gnd.n5212 gnd.n3692 163.367
R14698 gnd.n5212 gnd.n3679 163.367
R14699 gnd.n5224 gnd.n3679 163.367
R14700 gnd.n5224 gnd.n3676 163.367
R14701 gnd.n5229 gnd.n3676 163.367
R14702 gnd.n5229 gnd.n3677 163.367
R14703 gnd.n3677 gnd.n3659 163.367
R14704 gnd.n5252 gnd.n3659 163.367
R14705 gnd.n5252 gnd.n3657 163.367
R14706 gnd.n5256 gnd.n3657 163.367
R14707 gnd.n5256 gnd.n3649 163.367
R14708 gnd.n5271 gnd.n3649 163.367
R14709 gnd.n5271 gnd.n3647 163.367
R14710 gnd.n5275 gnd.n3647 163.367
R14711 gnd.n5275 gnd.n3634 163.367
R14712 gnd.n5295 gnd.n3634 163.367
R14713 gnd.n5295 gnd.n3632 163.367
R14714 gnd.n5299 gnd.n3632 163.367
R14715 gnd.n5299 gnd.n3624 163.367
R14716 gnd.n5308 gnd.n3624 163.367
R14717 gnd.n5308 gnd.n3621 163.367
R14718 gnd.n5314 gnd.n3621 163.367
R14719 gnd.n5314 gnd.n3622 163.367
R14720 gnd.n3622 gnd.n3611 163.367
R14721 gnd.n3611 gnd.n3599 163.367
R14722 gnd.n5335 gnd.n3599 163.367
R14723 gnd.n5335 gnd.n3597 163.367
R14724 gnd.n5339 gnd.n3597 163.367
R14725 gnd.n5339 gnd.n3588 163.367
R14726 gnd.n5353 gnd.n3588 163.367
R14727 gnd.n5353 gnd.n3586 163.367
R14728 gnd.n5357 gnd.n3586 163.367
R14729 gnd.n5357 gnd.n3571 163.367
R14730 gnd.n5368 gnd.n3571 163.367
R14731 gnd.n5368 gnd.n3569 163.367
R14732 gnd.n5372 gnd.n3569 163.367
R14733 gnd.n5372 gnd.n3557 163.367
R14734 gnd.n5393 gnd.n3557 163.367
R14735 gnd.n5393 gnd.n3558 163.367
R14736 gnd.n5389 gnd.n3558 163.367
R14737 gnd.n5389 gnd.n5388 163.367
R14738 gnd.n5388 gnd.n5387 163.367
R14739 gnd.n5387 gnd.n3561 163.367
R14740 gnd.n3561 gnd.n3458 163.367
R14741 gnd.n5543 gnd.n3458 163.367
R14742 gnd.n5543 gnd.n3459 163.367
R14743 gnd.n5539 gnd.n3459 163.367
R14744 gnd.n3479 gnd.n3478 156.462
R14745 gnd.n2265 gnd.n2233 153.042
R14746 gnd.n2329 gnd.n2328 152.079
R14747 gnd.n2297 gnd.n2296 152.079
R14748 gnd.n2265 gnd.n2264 152.079
R14749 gnd.n2887 gnd.n2886 152
R14750 gnd.n2888 gnd.n2877 152
R14751 gnd.n2890 gnd.n2889 152
R14752 gnd.n2892 gnd.n2875 152
R14753 gnd.n2894 gnd.n2893 152
R14754 gnd.n3477 gnd.n3461 152
R14755 gnd.n3469 gnd.n3462 152
R14756 gnd.n3468 gnd.n3467 152
R14757 gnd.n3466 gnd.n3463 152
R14758 gnd.n3464 gnd.t288 150.546
R14759 gnd.n7497 gnd.n7496 150.119
R14760 gnd.n7498 gnd.n7497 150.119
R14761 gnd.n7498 gnd.n487 150.119
R14762 gnd.n7506 gnd.n487 150.119
R14763 gnd.n7507 gnd.n7506 150.119
R14764 gnd.n7508 gnd.n7507 150.119
R14765 gnd.n7508 gnd.n481 150.119
R14766 gnd.n7516 gnd.n481 150.119
R14767 gnd.n7517 gnd.n7516 150.119
R14768 gnd.n7518 gnd.n7517 150.119
R14769 gnd.n7518 gnd.n475 150.119
R14770 gnd.n7526 gnd.n475 150.119
R14771 gnd.n7527 gnd.n7526 150.119
R14772 gnd.n7528 gnd.n7527 150.119
R14773 gnd.n7528 gnd.n469 150.119
R14774 gnd.n7536 gnd.n469 150.119
R14775 gnd.n7537 gnd.n7536 150.119
R14776 gnd.n7538 gnd.n7537 150.119
R14777 gnd.n7538 gnd.n463 150.119
R14778 gnd.n7546 gnd.n463 150.119
R14779 gnd.n7547 gnd.n7546 150.119
R14780 gnd.n7548 gnd.n7547 150.119
R14781 gnd.n7548 gnd.n457 150.119
R14782 gnd.n7556 gnd.n457 150.119
R14783 gnd.n7557 gnd.n7556 150.119
R14784 gnd.n7558 gnd.n7557 150.119
R14785 gnd.n7558 gnd.n451 150.119
R14786 gnd.n7566 gnd.n451 150.119
R14787 gnd.n7567 gnd.n7566 150.119
R14788 gnd.n7568 gnd.n7567 150.119
R14789 gnd.n7568 gnd.n445 150.119
R14790 gnd.n7576 gnd.n445 150.119
R14791 gnd.n7577 gnd.n7576 150.119
R14792 gnd.n7578 gnd.n7577 150.119
R14793 gnd.n7578 gnd.n439 150.119
R14794 gnd.n7586 gnd.n439 150.119
R14795 gnd.n7587 gnd.n7586 150.119
R14796 gnd.n7588 gnd.n7587 150.119
R14797 gnd.n7588 gnd.n433 150.119
R14798 gnd.n7596 gnd.n433 150.119
R14799 gnd.n7597 gnd.n7596 150.119
R14800 gnd.n7598 gnd.n7597 150.119
R14801 gnd.n7598 gnd.n427 150.119
R14802 gnd.n7606 gnd.n427 150.119
R14803 gnd.n7607 gnd.n7606 150.119
R14804 gnd.n7608 gnd.n7607 150.119
R14805 gnd.n7608 gnd.n421 150.119
R14806 gnd.n7616 gnd.n421 150.119
R14807 gnd.n7617 gnd.n7616 150.119
R14808 gnd.n7618 gnd.n7617 150.119
R14809 gnd.n7618 gnd.n415 150.119
R14810 gnd.n7626 gnd.n415 150.119
R14811 gnd.n7627 gnd.n7626 150.119
R14812 gnd.n7628 gnd.n7627 150.119
R14813 gnd.n7628 gnd.n409 150.119
R14814 gnd.n7636 gnd.n409 150.119
R14815 gnd.n7637 gnd.n7636 150.119
R14816 gnd.n7638 gnd.n7637 150.119
R14817 gnd.n7638 gnd.n403 150.119
R14818 gnd.n7646 gnd.n403 150.119
R14819 gnd.n7647 gnd.n7646 150.119
R14820 gnd.n7648 gnd.n7647 150.119
R14821 gnd.n7648 gnd.n397 150.119
R14822 gnd.n7656 gnd.n397 150.119
R14823 gnd.n7657 gnd.n7656 150.119
R14824 gnd.n7658 gnd.n7657 150.119
R14825 gnd.n7658 gnd.n391 150.119
R14826 gnd.n7666 gnd.n391 150.119
R14827 gnd.n7667 gnd.n7666 150.119
R14828 gnd.n7668 gnd.n7667 150.119
R14829 gnd.n7668 gnd.n385 150.119
R14830 gnd.n7676 gnd.n385 150.119
R14831 gnd.n7677 gnd.n7676 150.119
R14832 gnd.n7678 gnd.n7677 150.119
R14833 gnd.n7678 gnd.n379 150.119
R14834 gnd.n7686 gnd.n379 150.119
R14835 gnd.n7687 gnd.n7686 150.119
R14836 gnd.n7688 gnd.n7687 150.119
R14837 gnd.n7688 gnd.n373 150.119
R14838 gnd.n7696 gnd.n373 150.119
R14839 gnd.n7697 gnd.n7696 150.119
R14840 gnd.n7699 gnd.n7697 150.119
R14841 gnd.n7699 gnd.n7698 150.119
R14842 gnd.t397 gnd.n2307 147.661
R14843 gnd.t378 gnd.n2275 147.661
R14844 gnd.t363 gnd.n2243 147.661
R14845 gnd.t401 gnd.n2212 147.661
R14846 gnd.t1 gnd.n2180 147.661
R14847 gnd.t380 gnd.n2148 147.661
R14848 gnd.t383 gnd.n2116 147.661
R14849 gnd.t215 gnd.n2085 147.661
R14850 gnd.n5481 gnd.n5480 143.351
R14851 gnd.n2854 gnd.n2837 143.351
R14852 gnd.n6391 gnd.n2837 143.351
R14853 gnd.n2884 gnd.t247 130.484
R14854 gnd.n2893 gnd.t244 126.766
R14855 gnd.n2891 gnd.t297 126.766
R14856 gnd.n2877 gnd.t268 126.766
R14857 gnd.n2885 gnd.t322 126.766
R14858 gnd.n3465 gnd.t261 126.766
R14859 gnd.n3467 gnd.t291 126.766
R14860 gnd.n3476 gnd.t241 126.766
R14861 gnd.n3478 gnd.t313 126.766
R14862 gnd.n2324 gnd.n2323 104.615
R14863 gnd.n2323 gnd.n2301 104.615
R14864 gnd.n2316 gnd.n2301 104.615
R14865 gnd.n2316 gnd.n2315 104.615
R14866 gnd.n2315 gnd.n2305 104.615
R14867 gnd.n2308 gnd.n2305 104.615
R14868 gnd.n2292 gnd.n2291 104.615
R14869 gnd.n2291 gnd.n2269 104.615
R14870 gnd.n2284 gnd.n2269 104.615
R14871 gnd.n2284 gnd.n2283 104.615
R14872 gnd.n2283 gnd.n2273 104.615
R14873 gnd.n2276 gnd.n2273 104.615
R14874 gnd.n2260 gnd.n2259 104.615
R14875 gnd.n2259 gnd.n2237 104.615
R14876 gnd.n2252 gnd.n2237 104.615
R14877 gnd.n2252 gnd.n2251 104.615
R14878 gnd.n2251 gnd.n2241 104.615
R14879 gnd.n2244 gnd.n2241 104.615
R14880 gnd.n2229 gnd.n2228 104.615
R14881 gnd.n2228 gnd.n2206 104.615
R14882 gnd.n2221 gnd.n2206 104.615
R14883 gnd.n2221 gnd.n2220 104.615
R14884 gnd.n2220 gnd.n2210 104.615
R14885 gnd.n2213 gnd.n2210 104.615
R14886 gnd.n2197 gnd.n2196 104.615
R14887 gnd.n2196 gnd.n2174 104.615
R14888 gnd.n2189 gnd.n2174 104.615
R14889 gnd.n2189 gnd.n2188 104.615
R14890 gnd.n2188 gnd.n2178 104.615
R14891 gnd.n2181 gnd.n2178 104.615
R14892 gnd.n2165 gnd.n2164 104.615
R14893 gnd.n2164 gnd.n2142 104.615
R14894 gnd.n2157 gnd.n2142 104.615
R14895 gnd.n2157 gnd.n2156 104.615
R14896 gnd.n2156 gnd.n2146 104.615
R14897 gnd.n2149 gnd.n2146 104.615
R14898 gnd.n2133 gnd.n2132 104.615
R14899 gnd.n2132 gnd.n2110 104.615
R14900 gnd.n2125 gnd.n2110 104.615
R14901 gnd.n2125 gnd.n2124 104.615
R14902 gnd.n2124 gnd.n2114 104.615
R14903 gnd.n2117 gnd.n2114 104.615
R14904 gnd.n2102 gnd.n2101 104.615
R14905 gnd.n2101 gnd.n2079 104.615
R14906 gnd.n2094 gnd.n2079 104.615
R14907 gnd.n2094 gnd.n2093 104.615
R14908 gnd.n2093 gnd.n2083 104.615
R14909 gnd.n2086 gnd.n2083 104.615
R14910 gnd.n1495 gnd.t277 100.632
R14911 gnd.n1012 gnd.t308 100.632
R14912 gnd.n7972 gnd.n7971 99.6594
R14913 gnd.n7967 gnd.n294 99.6594
R14914 gnd.n7963 gnd.n293 99.6594
R14915 gnd.n7959 gnd.n292 99.6594
R14916 gnd.n7955 gnd.n291 99.6594
R14917 gnd.n7951 gnd.n290 99.6594
R14918 gnd.n7947 gnd.n289 99.6594
R14919 gnd.n7943 gnd.n288 99.6594
R14920 gnd.n7936 gnd.n287 99.6594
R14921 gnd.n7932 gnd.n286 99.6594
R14922 gnd.n7928 gnd.n285 99.6594
R14923 gnd.n7924 gnd.n284 99.6594
R14924 gnd.n7920 gnd.n283 99.6594
R14925 gnd.n7916 gnd.n282 99.6594
R14926 gnd.n7912 gnd.n281 99.6594
R14927 gnd.n7908 gnd.n280 99.6594
R14928 gnd.n7904 gnd.n279 99.6594
R14929 gnd.n7900 gnd.n278 99.6594
R14930 gnd.n7892 gnd.n277 99.6594
R14931 gnd.n7890 gnd.n276 99.6594
R14932 gnd.n7886 gnd.n275 99.6594
R14933 gnd.n7882 gnd.n274 99.6594
R14934 gnd.n7878 gnd.n273 99.6594
R14935 gnd.n7874 gnd.n272 99.6594
R14936 gnd.n7870 gnd.n271 99.6594
R14937 gnd.n7866 gnd.n270 99.6594
R14938 gnd.n7862 gnd.n269 99.6594
R14939 gnd.n7858 gnd.n268 99.6594
R14940 gnd.n7849 gnd.n267 99.6594
R14941 gnd.n6133 gnd.n6132 99.6594
R14942 gnd.n6127 gnd.n3076 99.6594
R14943 gnd.n6124 gnd.n3077 99.6594
R14944 gnd.n6120 gnd.n3078 99.6594
R14945 gnd.n6116 gnd.n3079 99.6594
R14946 gnd.n6112 gnd.n3080 99.6594
R14947 gnd.n6108 gnd.n3081 99.6594
R14948 gnd.n6104 gnd.n3082 99.6594
R14949 gnd.n6100 gnd.n3083 99.6594
R14950 gnd.n6095 gnd.n3084 99.6594
R14951 gnd.n6091 gnd.n3085 99.6594
R14952 gnd.n6087 gnd.n3086 99.6594
R14953 gnd.n6083 gnd.n3087 99.6594
R14954 gnd.n6078 gnd.n3089 99.6594
R14955 gnd.n6074 gnd.n3090 99.6594
R14956 gnd.n6070 gnd.n3091 99.6594
R14957 gnd.n6066 gnd.n3092 99.6594
R14958 gnd.n6062 gnd.n3093 99.6594
R14959 gnd.n6058 gnd.n3094 99.6594
R14960 gnd.n6054 gnd.n3095 99.6594
R14961 gnd.n6050 gnd.n3096 99.6594
R14962 gnd.n6046 gnd.n3097 99.6594
R14963 gnd.n6042 gnd.n3098 99.6594
R14964 gnd.n6038 gnd.n3099 99.6594
R14965 gnd.n6034 gnd.n3100 99.6594
R14966 gnd.n6030 gnd.n3101 99.6594
R14967 gnd.n6026 gnd.n3102 99.6594
R14968 gnd.n6022 gnd.n3103 99.6594
R14969 gnd.n6443 gnd.n6442 99.6594
R14970 gnd.n6438 gnd.n2804 99.6594
R14971 gnd.n6434 gnd.n2803 99.6594
R14972 gnd.n6430 gnd.n2802 99.6594
R14973 gnd.n6426 gnd.n2801 99.6594
R14974 gnd.n6422 gnd.n2800 99.6594
R14975 gnd.n6418 gnd.n2799 99.6594
R14976 gnd.n6414 gnd.n2798 99.6594
R14977 gnd.n6409 gnd.n2797 99.6594
R14978 gnd.n6405 gnd.n2796 99.6594
R14979 gnd.n6401 gnd.n2795 99.6594
R14980 gnd.n6397 gnd.n2794 99.6594
R14981 gnd.n4644 gnd.n2792 99.6594
R14982 gnd.n4648 gnd.n2791 99.6594
R14983 gnd.n4654 gnd.n2790 99.6594
R14984 gnd.n4658 gnd.n2789 99.6594
R14985 gnd.n4663 gnd.n2788 99.6594
R14986 gnd.n4667 gnd.n2787 99.6594
R14987 gnd.n4673 gnd.n2786 99.6594
R14988 gnd.n4677 gnd.n2785 99.6594
R14989 gnd.n4683 gnd.n2784 99.6594
R14990 gnd.n4687 gnd.n2783 99.6594
R14991 gnd.n4693 gnd.n2782 99.6594
R14992 gnd.n4697 gnd.n2781 99.6594
R14993 gnd.n4703 gnd.n2780 99.6594
R14994 gnd.n4707 gnd.n2779 99.6594
R14995 gnd.n4712 gnd.n2778 99.6594
R14996 gnd.n4715 gnd.n2777 99.6594
R14997 gnd.n6744 gnd.n6743 99.6594
R14998 gnd.n6738 gnd.n2356 99.6594
R14999 gnd.n6735 gnd.n2357 99.6594
R15000 gnd.n6731 gnd.n2358 99.6594
R15001 gnd.n6727 gnd.n2359 99.6594
R15002 gnd.n6723 gnd.n2360 99.6594
R15003 gnd.n6719 gnd.n2361 99.6594
R15004 gnd.n6715 gnd.n2362 99.6594
R15005 gnd.n6711 gnd.n2363 99.6594
R15006 gnd.n6706 gnd.n2364 99.6594
R15007 gnd.n6702 gnd.n2365 99.6594
R15008 gnd.n6698 gnd.n2366 99.6594
R15009 gnd.n6694 gnd.n2367 99.6594
R15010 gnd.n6690 gnd.n2368 99.6594
R15011 gnd.n6686 gnd.n2369 99.6594
R15012 gnd.n6682 gnd.n2370 99.6594
R15013 gnd.n6678 gnd.n2371 99.6594
R15014 gnd.n6674 gnd.n2372 99.6594
R15015 gnd.n6670 gnd.n2373 99.6594
R15016 gnd.n6666 gnd.n2374 99.6594
R15017 gnd.n6662 gnd.n2375 99.6594
R15018 gnd.n6658 gnd.n2376 99.6594
R15019 gnd.n6654 gnd.n2377 99.6594
R15020 gnd.n6650 gnd.n2378 99.6594
R15021 gnd.n6646 gnd.n2379 99.6594
R15022 gnd.n6642 gnd.n2380 99.6594
R15023 gnd.n6638 gnd.n2381 99.6594
R15024 gnd.n6634 gnd.n2382 99.6594
R15025 gnd.n6630 gnd.n2383 99.6594
R15026 gnd.n6783 gnd.n6751 99.6594
R15027 gnd.n6781 gnd.n6750 99.6594
R15028 gnd.n6777 gnd.n6749 99.6594
R15029 gnd.n6773 gnd.n6748 99.6594
R15030 gnd.n6769 gnd.n6747 99.6594
R15031 gnd.n6765 gnd.n6746 99.6594
R15032 gnd.n6795 gnd.n6793 99.6594
R15033 gnd.n6801 gnd.n1011 99.6594
R15034 gnd.n1707 gnd.n1438 99.6594
R15035 gnd.n1464 gnd.n1445 99.6594
R15036 gnd.n1466 gnd.n1446 99.6594
R15037 gnd.n1474 gnd.n1447 99.6594
R15038 gnd.n1476 gnd.n1448 99.6594
R15039 gnd.n1484 gnd.n1449 99.6594
R15040 gnd.n1486 gnd.n1450 99.6594
R15041 gnd.n1494 gnd.n1451 99.6594
R15042 gnd.n7754 gnd.n258 99.6594
R15043 gnd.n7758 gnd.n259 99.6594
R15044 gnd.n7764 gnd.n260 99.6594
R15045 gnd.n7768 gnd.n261 99.6594
R15046 gnd.n7774 gnd.n262 99.6594
R15047 gnd.n7778 gnd.n263 99.6594
R15048 gnd.n7784 gnd.n264 99.6594
R15049 gnd.n7788 gnd.n265 99.6594
R15050 gnd.n7794 gnd.n266 99.6594
R15051 gnd.n3188 gnd.n3104 99.6594
R15052 gnd.n3106 gnd.n3030 99.6594
R15053 gnd.n3107 gnd.n3037 99.6594
R15054 gnd.n3109 gnd.n3108 99.6594
R15055 gnd.n3111 gnd.n3046 99.6594
R15056 gnd.n3112 gnd.n3053 99.6594
R15057 gnd.n3114 gnd.n3113 99.6594
R15058 gnd.n3116 gnd.n3062 99.6594
R15059 gnd.n6135 gnd.n3071 99.6594
R15060 gnd.n1053 gnd.n1018 99.6594
R15061 gnd.n1057 gnd.n1019 99.6594
R15062 gnd.n1063 gnd.n1020 99.6594
R15063 gnd.n1067 gnd.n1021 99.6594
R15064 gnd.n1073 gnd.n1022 99.6594
R15065 gnd.n1077 gnd.n1023 99.6594
R15066 gnd.n1083 gnd.n1024 99.6594
R15067 gnd.n1087 gnd.n1025 99.6594
R15068 gnd.n1093 gnd.n1026 99.6594
R15069 gnd.n1097 gnd.n1027 99.6594
R15070 gnd.n1103 gnd.n1028 99.6594
R15071 gnd.n1106 gnd.n1029 99.6594
R15072 gnd.n2355 gnd.n2354 99.6594
R15073 gnd.n1622 gnd.n1621 99.6594
R15074 gnd.n1616 gnd.n1533 99.6594
R15075 gnd.n1613 gnd.n1534 99.6594
R15076 gnd.n1609 gnd.n1535 99.6594
R15077 gnd.n1605 gnd.n1536 99.6594
R15078 gnd.n1601 gnd.n1537 99.6594
R15079 gnd.n1597 gnd.n1538 99.6594
R15080 gnd.n1593 gnd.n1539 99.6594
R15081 gnd.n1589 gnd.n1540 99.6594
R15082 gnd.n1585 gnd.n1541 99.6594
R15083 gnd.n1581 gnd.n1542 99.6594
R15084 gnd.n1577 gnd.n1543 99.6594
R15085 gnd.n1624 gnd.n1532 99.6594
R15086 gnd.n4519 gnd.n2767 99.6594
R15087 gnd.n4521 gnd.n2768 99.6594
R15088 gnd.n4529 gnd.n2769 99.6594
R15089 gnd.n4539 gnd.n2770 99.6594
R15090 gnd.n4541 gnd.n2771 99.6594
R15091 gnd.n4549 gnd.n2772 99.6594
R15092 gnd.n4559 gnd.n2773 99.6594
R15093 gnd.n4562 gnd.n2774 99.6594
R15094 gnd.n4766 gnd.n2775 99.6594
R15095 gnd.n4120 gnd.n2384 99.6594
R15096 gnd.n4124 gnd.n2385 99.6594
R15097 gnd.n4130 gnd.n2386 99.6594
R15098 gnd.n4134 gnd.n2387 99.6594
R15099 gnd.n4140 gnd.n2388 99.6594
R15100 gnd.n4144 gnd.n2389 99.6594
R15101 gnd.n4150 gnd.n2390 99.6594
R15102 gnd.n4154 gnd.n2391 99.6594
R15103 gnd.n4111 gnd.n2392 99.6594
R15104 gnd.n4123 gnd.n2384 99.6594
R15105 gnd.n4129 gnd.n2385 99.6594
R15106 gnd.n4133 gnd.n2386 99.6594
R15107 gnd.n4139 gnd.n2387 99.6594
R15108 gnd.n4143 gnd.n2388 99.6594
R15109 gnd.n4149 gnd.n2389 99.6594
R15110 gnd.n4153 gnd.n2390 99.6594
R15111 gnd.n4110 gnd.n2391 99.6594
R15112 gnd.n4106 gnd.n2392 99.6594
R15113 gnd.n4561 gnd.n2775 99.6594
R15114 gnd.n4560 gnd.n2774 99.6594
R15115 gnd.n4550 gnd.n2773 99.6594
R15116 gnd.n4542 gnd.n2772 99.6594
R15117 gnd.n4540 gnd.n2771 99.6594
R15118 gnd.n4530 gnd.n2770 99.6594
R15119 gnd.n4522 gnd.n2769 99.6594
R15120 gnd.n4520 gnd.n2768 99.6594
R15121 gnd.n4510 gnd.n2767 99.6594
R15122 gnd.n1622 gnd.n1545 99.6594
R15123 gnd.n1614 gnd.n1533 99.6594
R15124 gnd.n1610 gnd.n1534 99.6594
R15125 gnd.n1606 gnd.n1535 99.6594
R15126 gnd.n1602 gnd.n1536 99.6594
R15127 gnd.n1598 gnd.n1537 99.6594
R15128 gnd.n1594 gnd.n1538 99.6594
R15129 gnd.n1590 gnd.n1539 99.6594
R15130 gnd.n1586 gnd.n1540 99.6594
R15131 gnd.n1582 gnd.n1541 99.6594
R15132 gnd.n1578 gnd.n1542 99.6594
R15133 gnd.n1574 gnd.n1543 99.6594
R15134 gnd.n1625 gnd.n1624 99.6594
R15135 gnd.n2355 gnd.n1030 99.6594
R15136 gnd.n1104 gnd.n1029 99.6594
R15137 gnd.n1096 gnd.n1028 99.6594
R15138 gnd.n1094 gnd.n1027 99.6594
R15139 gnd.n1086 gnd.n1026 99.6594
R15140 gnd.n1084 gnd.n1025 99.6594
R15141 gnd.n1076 gnd.n1024 99.6594
R15142 gnd.n1074 gnd.n1023 99.6594
R15143 gnd.n1066 gnd.n1022 99.6594
R15144 gnd.n1064 gnd.n1021 99.6594
R15145 gnd.n1056 gnd.n1020 99.6594
R15146 gnd.n1054 gnd.n1019 99.6594
R15147 gnd.n1046 gnd.n1018 99.6594
R15148 gnd.n3104 gnd.n3029 99.6594
R15149 gnd.n3106 gnd.n3105 99.6594
R15150 gnd.n3107 gnd.n3038 99.6594
R15151 gnd.n3109 gnd.n3045 99.6594
R15152 gnd.n3111 gnd.n3110 99.6594
R15153 gnd.n3112 gnd.n3054 99.6594
R15154 gnd.n3114 gnd.n3061 99.6594
R15155 gnd.n3116 gnd.n3115 99.6594
R15156 gnd.n6136 gnd.n6135 99.6594
R15157 gnd.n7787 gnd.n266 99.6594
R15158 gnd.n7785 gnd.n265 99.6594
R15159 gnd.n7777 gnd.n264 99.6594
R15160 gnd.n7775 gnd.n263 99.6594
R15161 gnd.n7767 gnd.n262 99.6594
R15162 gnd.n7765 gnd.n261 99.6594
R15163 gnd.n7757 gnd.n260 99.6594
R15164 gnd.n7755 gnd.n259 99.6594
R15165 gnd.n7749 gnd.n258 99.6594
R15166 gnd.n1708 gnd.n1707 99.6594
R15167 gnd.n1467 gnd.n1445 99.6594
R15168 gnd.n1473 gnd.n1446 99.6594
R15169 gnd.n1477 gnd.n1447 99.6594
R15170 gnd.n1483 gnd.n1448 99.6594
R15171 gnd.n1487 gnd.n1449 99.6594
R15172 gnd.n1493 gnd.n1450 99.6594
R15173 gnd.n1451 gnd.n1435 99.6594
R15174 gnd.n6794 gnd.n1011 99.6594
R15175 gnd.n6793 gnd.n1017 99.6594
R15176 gnd.n6768 gnd.n6746 99.6594
R15177 gnd.n6772 gnd.n6747 99.6594
R15178 gnd.n6776 gnd.n6748 99.6594
R15179 gnd.n6780 gnd.n6749 99.6594
R15180 gnd.n6784 gnd.n6750 99.6594
R15181 gnd.n6752 gnd.n6751 99.6594
R15182 gnd.n6744 gnd.n2396 99.6594
R15183 gnd.n6736 gnd.n2356 99.6594
R15184 gnd.n6732 gnd.n2357 99.6594
R15185 gnd.n6728 gnd.n2358 99.6594
R15186 gnd.n6724 gnd.n2359 99.6594
R15187 gnd.n6720 gnd.n2360 99.6594
R15188 gnd.n6716 gnd.n2361 99.6594
R15189 gnd.n6712 gnd.n2362 99.6594
R15190 gnd.n6707 gnd.n2363 99.6594
R15191 gnd.n6703 gnd.n2364 99.6594
R15192 gnd.n6699 gnd.n2365 99.6594
R15193 gnd.n6695 gnd.n2366 99.6594
R15194 gnd.n6691 gnd.n2367 99.6594
R15195 gnd.n6687 gnd.n2368 99.6594
R15196 gnd.n6683 gnd.n2369 99.6594
R15197 gnd.n6679 gnd.n2370 99.6594
R15198 gnd.n6675 gnd.n2371 99.6594
R15199 gnd.n6671 gnd.n2372 99.6594
R15200 gnd.n6667 gnd.n2373 99.6594
R15201 gnd.n6663 gnd.n2374 99.6594
R15202 gnd.n6659 gnd.n2375 99.6594
R15203 gnd.n6655 gnd.n2376 99.6594
R15204 gnd.n6651 gnd.n2377 99.6594
R15205 gnd.n6647 gnd.n2378 99.6594
R15206 gnd.n6643 gnd.n2379 99.6594
R15207 gnd.n6639 gnd.n2380 99.6594
R15208 gnd.n6635 gnd.n2381 99.6594
R15209 gnd.n6631 gnd.n2382 99.6594
R15210 gnd.n2466 gnd.n2383 99.6594
R15211 gnd.n4625 gnd.n2777 99.6594
R15212 gnd.n4706 gnd.n2778 99.6594
R15213 gnd.n4704 gnd.n2779 99.6594
R15214 gnd.n4696 gnd.n2780 99.6594
R15215 gnd.n4694 gnd.n2781 99.6594
R15216 gnd.n4686 gnd.n2782 99.6594
R15217 gnd.n4684 gnd.n2783 99.6594
R15218 gnd.n4676 gnd.n2784 99.6594
R15219 gnd.n4674 gnd.n2785 99.6594
R15220 gnd.n4666 gnd.n2786 99.6594
R15221 gnd.n4638 gnd.n2787 99.6594
R15222 gnd.n4657 gnd.n2788 99.6594
R15223 gnd.n4655 gnd.n2789 99.6594
R15224 gnd.n4647 gnd.n2790 99.6594
R15225 gnd.n4645 gnd.n2791 99.6594
R15226 gnd.n6396 gnd.n2793 99.6594
R15227 gnd.n6400 gnd.n2794 99.6594
R15228 gnd.n6404 gnd.n2795 99.6594
R15229 gnd.n6408 gnd.n2796 99.6594
R15230 gnd.n6413 gnd.n2797 99.6594
R15231 gnd.n6417 gnd.n2798 99.6594
R15232 gnd.n6421 gnd.n2799 99.6594
R15233 gnd.n6425 gnd.n2800 99.6594
R15234 gnd.n6429 gnd.n2801 99.6594
R15235 gnd.n6433 gnd.n2802 99.6594
R15236 gnd.n6437 gnd.n2803 99.6594
R15237 gnd.n2805 gnd.n2804 99.6594
R15238 gnd.n6443 gnd.n2764 99.6594
R15239 gnd.n6133 gnd.n3119 99.6594
R15240 gnd.n6125 gnd.n3076 99.6594
R15241 gnd.n6121 gnd.n3077 99.6594
R15242 gnd.n6117 gnd.n3078 99.6594
R15243 gnd.n6113 gnd.n3079 99.6594
R15244 gnd.n6109 gnd.n3080 99.6594
R15245 gnd.n6105 gnd.n3081 99.6594
R15246 gnd.n6101 gnd.n3082 99.6594
R15247 gnd.n6096 gnd.n3083 99.6594
R15248 gnd.n6092 gnd.n3084 99.6594
R15249 gnd.n6088 gnd.n3085 99.6594
R15250 gnd.n6084 gnd.n3086 99.6594
R15251 gnd.n6079 gnd.n3088 99.6594
R15252 gnd.n6075 gnd.n3089 99.6594
R15253 gnd.n6071 gnd.n3090 99.6594
R15254 gnd.n6067 gnd.n3091 99.6594
R15255 gnd.n6063 gnd.n3092 99.6594
R15256 gnd.n6059 gnd.n3093 99.6594
R15257 gnd.n6055 gnd.n3094 99.6594
R15258 gnd.n6051 gnd.n3095 99.6594
R15259 gnd.n6047 gnd.n3096 99.6594
R15260 gnd.n6043 gnd.n3097 99.6594
R15261 gnd.n6039 gnd.n3098 99.6594
R15262 gnd.n6035 gnd.n3099 99.6594
R15263 gnd.n6031 gnd.n3100 99.6594
R15264 gnd.n6027 gnd.n3101 99.6594
R15265 gnd.n6023 gnd.n3102 99.6594
R15266 gnd.n6015 gnd.n3103 99.6594
R15267 gnd.n7857 gnd.n267 99.6594
R15268 gnd.n7861 gnd.n268 99.6594
R15269 gnd.n7865 gnd.n269 99.6594
R15270 gnd.n7869 gnd.n270 99.6594
R15271 gnd.n7873 gnd.n271 99.6594
R15272 gnd.n7877 gnd.n272 99.6594
R15273 gnd.n7881 gnd.n273 99.6594
R15274 gnd.n7885 gnd.n274 99.6594
R15275 gnd.n7889 gnd.n275 99.6594
R15276 gnd.n7893 gnd.n276 99.6594
R15277 gnd.n7899 gnd.n277 99.6594
R15278 gnd.n7903 gnd.n278 99.6594
R15279 gnd.n7907 gnd.n279 99.6594
R15280 gnd.n7911 gnd.n280 99.6594
R15281 gnd.n7915 gnd.n281 99.6594
R15282 gnd.n7919 gnd.n282 99.6594
R15283 gnd.n7923 gnd.n283 99.6594
R15284 gnd.n7927 gnd.n284 99.6594
R15285 gnd.n7931 gnd.n285 99.6594
R15286 gnd.n7935 gnd.n286 99.6594
R15287 gnd.n7942 gnd.n287 99.6594
R15288 gnd.n7946 gnd.n288 99.6594
R15289 gnd.n7950 gnd.n289 99.6594
R15290 gnd.n7954 gnd.n290 99.6594
R15291 gnd.n7958 gnd.n291 99.6594
R15292 gnd.n7962 gnd.n292 99.6594
R15293 gnd.n7966 gnd.n293 99.6594
R15294 gnd.n295 gnd.n294 99.6594
R15295 gnd.n7972 gnd.n255 99.6594
R15296 gnd.n4493 gnd.n3935 99.6594
R15297 gnd.n4497 gnd.n3936 99.6594
R15298 gnd.n4480 gnd.n3937 99.6594
R15299 gnd.n4505 gnd.n3938 99.6594
R15300 gnd.n4507 gnd.n3939 99.6594
R15301 gnd.n4514 gnd.n3940 99.6594
R15302 gnd.n4516 gnd.n3941 99.6594
R15303 gnd.n4526 gnd.n3942 99.6594
R15304 gnd.n4534 gnd.n3943 99.6594
R15305 gnd.n4536 gnd.n3944 99.6594
R15306 gnd.n4546 gnd.n3945 99.6594
R15307 gnd.n4554 gnd.n3946 99.6594
R15308 gnd.n4556 gnd.n3947 99.6594
R15309 gnd.n4568 gnd.n3948 99.6594
R15310 gnd.n4496 gnd.n3935 99.6594
R15311 gnd.n4479 gnd.n3936 99.6594
R15312 gnd.n4504 gnd.n3937 99.6594
R15313 gnd.n4506 gnd.n3938 99.6594
R15314 gnd.n4513 gnd.n3939 99.6594
R15315 gnd.n4515 gnd.n3940 99.6594
R15316 gnd.n4525 gnd.n3941 99.6594
R15317 gnd.n4533 gnd.n3942 99.6594
R15318 gnd.n4535 gnd.n3943 99.6594
R15319 gnd.n4545 gnd.n3944 99.6594
R15320 gnd.n4553 gnd.n3945 99.6594
R15321 gnd.n4555 gnd.n3946 99.6594
R15322 gnd.n4567 gnd.n3947 99.6594
R15323 gnd.n3949 gnd.n3948 99.6594
R15324 gnd.n3398 gnd.n3010 99.6594
R15325 gnd.n3400 gnd.n3015 99.6594
R15326 gnd.n3401 gnd.n3018 99.6594
R15327 gnd.n3403 gnd.n3020 99.6594
R15328 gnd.n3404 gnd.n3024 99.6594
R15329 gnd.n3406 gnd.n3405 99.6594
R15330 gnd.n3408 gnd.n3034 99.6594
R15331 gnd.n3409 gnd.n3041 99.6594
R15332 gnd.n3411 gnd.n3410 99.6594
R15333 gnd.n3413 gnd.n3050 99.6594
R15334 gnd.n3414 gnd.n3057 99.6594
R15335 gnd.n3416 gnd.n3415 99.6594
R15336 gnd.n3419 gnd.n3066 99.6594
R15337 gnd.n5683 gnd.n3397 99.6594
R15338 gnd.n3416 gnd.n3065 99.6594
R15339 gnd.n3414 gnd.n3058 99.6594
R15340 gnd.n3413 gnd.n3412 99.6594
R15341 gnd.n3411 gnd.n3049 99.6594
R15342 gnd.n3409 gnd.n3042 99.6594
R15343 gnd.n3408 gnd.n3407 99.6594
R15344 gnd.n3406 gnd.n3033 99.6594
R15345 gnd.n3404 gnd.n3025 99.6594
R15346 gnd.n3403 gnd.n3402 99.6594
R15347 gnd.n3401 gnd.n3019 99.6594
R15348 gnd.n3400 gnd.n3399 99.6594
R15349 gnd.n3398 gnd.n3014 99.6594
R15350 gnd.n5684 gnd.n5683 99.6594
R15351 gnd.n3419 gnd.n3418 99.6594
R15352 gnd.n4564 gnd.t284 98.63
R15353 gnd.n6137 gnd.t312 98.63
R15354 gnd.n3953 gnd.t329 98.63
R15355 gnd.n3139 gnd.t305 98.63
R15356 gnd.n3162 gnd.t296 98.63
R15357 gnd.n6017 gnd.t228 98.63
R15358 gnd.n352 gnd.t335 98.63
R15359 gnd.n332 gnd.t239 98.63
R15360 gnd.n7938 gnd.t272 98.63
R15361 gnd.n7738 gnd.t286 98.63
R15362 gnd.n2416 gnd.t302 98.63
R15363 gnd.n2438 gnd.t232 98.63
R15364 gnd.n2460 gnd.t256 98.63
R15365 gnd.n4107 gnd.t333 98.63
R15366 gnd.n2822 gnd.t326 98.63
R15367 gnd.n4623 gnd.t252 98.63
R15368 gnd.n4636 gnd.t279 98.63
R15369 gnd.n3067 gnd.t259 98.63
R15370 gnd.n3827 gnd.t318 96.6984
R15371 gnd.n3510 gnd.t266 96.6984
R15372 gnd.n6325 gnd.t236 96.6906
R15373 gnd.n3504 gnd.t320 96.6906
R15374 gnd.n7698 gnd.n256 90.0721
R15375 gnd.n2884 gnd.n2883 81.8399
R15376 gnd.n6081 gnd.n3149 77.1205
R15377 gnd.n6394 gnd.n6393 77.1205
R15378 gnd.n1496 gnd.t276 74.8376
R15379 gnd.n1013 gnd.t309 74.8376
R15380 gnd.n3828 gnd.t317 72.8438
R15381 gnd.n3511 gnd.t267 72.8438
R15382 gnd.n2885 gnd.n2878 72.8411
R15383 gnd.n2891 gnd.n2876 72.8411
R15384 gnd.n3476 gnd.n3475 72.8411
R15385 gnd.n4565 gnd.t283 72.836
R15386 gnd.n6326 gnd.t235 72.836
R15387 gnd.n3505 gnd.t321 72.836
R15388 gnd.n6138 gnd.t311 72.836
R15389 gnd.n3954 gnd.t330 72.836
R15390 gnd.n3140 gnd.t304 72.836
R15391 gnd.n3163 gnd.t295 72.836
R15392 gnd.n6018 gnd.t227 72.836
R15393 gnd.n353 gnd.t336 72.836
R15394 gnd.n333 gnd.t240 72.836
R15395 gnd.n7939 gnd.t273 72.836
R15396 gnd.n7739 gnd.t287 72.836
R15397 gnd.n2417 gnd.t301 72.836
R15398 gnd.n2439 gnd.t231 72.836
R15399 gnd.n2461 gnd.t255 72.836
R15400 gnd.n4108 gnd.t332 72.836
R15401 gnd.n2823 gnd.t327 72.836
R15402 gnd.n4624 gnd.t253 72.836
R15403 gnd.n4637 gnd.t280 72.836
R15404 gnd.n3068 gnd.t260 72.836
R15405 gnd.n5537 gnd.n5536 71.676
R15406 gnd.n5532 gnd.n3484 71.676
R15407 gnd.n5530 gnd.n5529 71.676
R15408 gnd.n5525 gnd.n3487 71.676
R15409 gnd.n5523 gnd.n5522 71.676
R15410 gnd.n5518 gnd.n3490 71.676
R15411 gnd.n5516 gnd.n5515 71.676
R15412 gnd.n5511 gnd.n3493 71.676
R15413 gnd.n5509 gnd.n5508 71.676
R15414 gnd.n5504 gnd.n3496 71.676
R15415 gnd.n5502 gnd.n5501 71.676
R15416 gnd.n5497 gnd.n3499 71.676
R15417 gnd.n5495 gnd.n5494 71.676
R15418 gnd.n5490 gnd.n3502 71.676
R15419 gnd.n5488 gnd.n5487 71.676
R15420 gnd.n5483 gnd.n3507 71.676
R15421 gnd.n5480 gnd.n5479 71.676
R15422 gnd.n5477 gnd.n5476 71.676
R15423 gnd.n5471 gnd.n3513 71.676
R15424 gnd.n5469 gnd.n5468 71.676
R15425 gnd.n5464 gnd.n3516 71.676
R15426 gnd.n5462 gnd.n5461 71.676
R15427 gnd.n5457 gnd.n3519 71.676
R15428 gnd.n5455 gnd.n5454 71.676
R15429 gnd.n5450 gnd.n3522 71.676
R15430 gnd.n5448 gnd.n5447 71.676
R15431 gnd.n5443 gnd.n3525 71.676
R15432 gnd.n5441 gnd.n5440 71.676
R15433 gnd.n5436 gnd.n3528 71.676
R15434 gnd.n5434 gnd.n5433 71.676
R15435 gnd.n5429 gnd.n3531 71.676
R15436 gnd.n5427 gnd.n5426 71.676
R15437 gnd.n5422 gnd.n3534 71.676
R15438 gnd.n6389 gnd.n6388 71.676
R15439 gnd.n6383 gnd.n2840 71.676
R15440 gnd.n6380 gnd.n2841 71.676
R15441 gnd.n6376 gnd.n2842 71.676
R15442 gnd.n6372 gnd.n2843 71.676
R15443 gnd.n6368 gnd.n2844 71.676
R15444 gnd.n6364 gnd.n2845 71.676
R15445 gnd.n6360 gnd.n2846 71.676
R15446 gnd.n6356 gnd.n2847 71.676
R15447 gnd.n6352 gnd.n2848 71.676
R15448 gnd.n6348 gnd.n2849 71.676
R15449 gnd.n6344 gnd.n2850 71.676
R15450 gnd.n6340 gnd.n2851 71.676
R15451 gnd.n6336 gnd.n2852 71.676
R15452 gnd.n6332 gnd.n2853 71.676
R15453 gnd.n6328 gnd.n2854 71.676
R15454 gnd.n2855 gnd.n2838 71.676
R15455 gnd.n3831 gnd.n2856 71.676
R15456 gnd.n3836 gnd.n2857 71.676
R15457 gnd.n3840 gnd.n2858 71.676
R15458 gnd.n3844 gnd.n2859 71.676
R15459 gnd.n3848 gnd.n2860 71.676
R15460 gnd.n3852 gnd.n2861 71.676
R15461 gnd.n3856 gnd.n2862 71.676
R15462 gnd.n3860 gnd.n2863 71.676
R15463 gnd.n3864 gnd.n2864 71.676
R15464 gnd.n3868 gnd.n2865 71.676
R15465 gnd.n3872 gnd.n2866 71.676
R15466 gnd.n3876 gnd.n2867 71.676
R15467 gnd.n3880 gnd.n2868 71.676
R15468 gnd.n3884 gnd.n2869 71.676
R15469 gnd.n3888 gnd.n2870 71.676
R15470 gnd.n6389 gnd.n2873 71.676
R15471 gnd.n6381 gnd.n2840 71.676
R15472 gnd.n6377 gnd.n2841 71.676
R15473 gnd.n6373 gnd.n2842 71.676
R15474 gnd.n6369 gnd.n2843 71.676
R15475 gnd.n6365 gnd.n2844 71.676
R15476 gnd.n6361 gnd.n2845 71.676
R15477 gnd.n6357 gnd.n2846 71.676
R15478 gnd.n6353 gnd.n2847 71.676
R15479 gnd.n6349 gnd.n2848 71.676
R15480 gnd.n6345 gnd.n2849 71.676
R15481 gnd.n6341 gnd.n2850 71.676
R15482 gnd.n6337 gnd.n2851 71.676
R15483 gnd.n6333 gnd.n2852 71.676
R15484 gnd.n6329 gnd.n2853 71.676
R15485 gnd.n6392 gnd.n6391 71.676
R15486 gnd.n3830 gnd.n2855 71.676
R15487 gnd.n3835 gnd.n2856 71.676
R15488 gnd.n3839 gnd.n2857 71.676
R15489 gnd.n3843 gnd.n2858 71.676
R15490 gnd.n3847 gnd.n2859 71.676
R15491 gnd.n3851 gnd.n2860 71.676
R15492 gnd.n3855 gnd.n2861 71.676
R15493 gnd.n3859 gnd.n2862 71.676
R15494 gnd.n3863 gnd.n2863 71.676
R15495 gnd.n3867 gnd.n2864 71.676
R15496 gnd.n3871 gnd.n2865 71.676
R15497 gnd.n3875 gnd.n2866 71.676
R15498 gnd.n3879 gnd.n2867 71.676
R15499 gnd.n3883 gnd.n2868 71.676
R15500 gnd.n3887 gnd.n2869 71.676
R15501 gnd.n3891 gnd.n2870 71.676
R15502 gnd.n3534 gnd.n3532 71.676
R15503 gnd.n5428 gnd.n5427 71.676
R15504 gnd.n3531 gnd.n3529 71.676
R15505 gnd.n5435 gnd.n5434 71.676
R15506 gnd.n3528 gnd.n3526 71.676
R15507 gnd.n5442 gnd.n5441 71.676
R15508 gnd.n3525 gnd.n3523 71.676
R15509 gnd.n5449 gnd.n5448 71.676
R15510 gnd.n3522 gnd.n3520 71.676
R15511 gnd.n5456 gnd.n5455 71.676
R15512 gnd.n3519 gnd.n3517 71.676
R15513 gnd.n5463 gnd.n5462 71.676
R15514 gnd.n3516 gnd.n3514 71.676
R15515 gnd.n5470 gnd.n5469 71.676
R15516 gnd.n3513 gnd.n3509 71.676
R15517 gnd.n5478 gnd.n5477 71.676
R15518 gnd.n5482 gnd.n5481 71.676
R15519 gnd.n3507 gnd.n3503 71.676
R15520 gnd.n5489 gnd.n5488 71.676
R15521 gnd.n3502 gnd.n3500 71.676
R15522 gnd.n5496 gnd.n5495 71.676
R15523 gnd.n3499 gnd.n3497 71.676
R15524 gnd.n5503 gnd.n5502 71.676
R15525 gnd.n3496 gnd.n3494 71.676
R15526 gnd.n5510 gnd.n5509 71.676
R15527 gnd.n3493 gnd.n3491 71.676
R15528 gnd.n5517 gnd.n5516 71.676
R15529 gnd.n3490 gnd.n3488 71.676
R15530 gnd.n5524 gnd.n5523 71.676
R15531 gnd.n3487 gnd.n3485 71.676
R15532 gnd.n5531 gnd.n5530 71.676
R15533 gnd.n3484 gnd.n3482 71.676
R15534 gnd.n5538 gnd.n5537 71.676
R15535 gnd.n8 gnd.t399 69.1507
R15536 gnd.n14 gnd.t371 68.4792
R15537 gnd.n13 gnd.t391 68.4792
R15538 gnd.n12 gnd.t211 68.4792
R15539 gnd.n11 gnd.t376 68.4792
R15540 gnd.n10 gnd.t218 68.4792
R15541 gnd.n9 gnd.t355 68.4792
R15542 gnd.n8 gnd.t213 68.4792
R15543 gnd.n1623 gnd.n1527 64.369
R15544 gnd.n3833 gnd.n3828 59.5399
R15545 gnd.n5473 gnd.n3511 59.5399
R15546 gnd.n6327 gnd.n6326 59.5399
R15547 gnd.n3506 gnd.n3505 59.5399
R15548 gnd.n6324 gnd.n2894 59.1804
R15549 gnd.n6792 gnd.n1004 57.3586
R15550 gnd.n1314 gnd.t101 56.407
R15551 gnd.n1255 gnd.t185 56.407
R15552 gnd.n1274 gnd.t36 56.407
R15553 gnd.n1294 gnd.t172 56.407
R15554 gnd.n76 gnd.t64 56.407
R15555 gnd.n17 gnd.t49 56.407
R15556 gnd.n36 gnd.t201 56.407
R15557 gnd.n56 gnd.t127 56.407
R15558 gnd.n1331 gnd.t157 55.8337
R15559 gnd.n1272 gnd.t26 55.8337
R15560 gnd.n1291 gnd.t188 55.8337
R15561 gnd.n1311 gnd.t60 55.8337
R15562 gnd.n93 gnd.t81 55.8337
R15563 gnd.n34 gnd.t51 55.8337
R15564 gnd.n53 gnd.t123 55.8337
R15565 gnd.n73 gnd.t140 55.8337
R15566 gnd.n2882 gnd.n2881 54.358
R15567 gnd.n3473 gnd.n3472 54.358
R15568 gnd.n1314 gnd.n1313 53.0052
R15569 gnd.n1316 gnd.n1315 53.0052
R15570 gnd.n1318 gnd.n1317 53.0052
R15571 gnd.n1320 gnd.n1319 53.0052
R15572 gnd.n1322 gnd.n1321 53.0052
R15573 gnd.n1324 gnd.n1323 53.0052
R15574 gnd.n1326 gnd.n1325 53.0052
R15575 gnd.n1328 gnd.n1327 53.0052
R15576 gnd.n1330 gnd.n1329 53.0052
R15577 gnd.n1255 gnd.n1254 53.0052
R15578 gnd.n1257 gnd.n1256 53.0052
R15579 gnd.n1259 gnd.n1258 53.0052
R15580 gnd.n1261 gnd.n1260 53.0052
R15581 gnd.n1263 gnd.n1262 53.0052
R15582 gnd.n1265 gnd.n1264 53.0052
R15583 gnd.n1267 gnd.n1266 53.0052
R15584 gnd.n1269 gnd.n1268 53.0052
R15585 gnd.n1271 gnd.n1270 53.0052
R15586 gnd.n1274 gnd.n1273 53.0052
R15587 gnd.n1276 gnd.n1275 53.0052
R15588 gnd.n1278 gnd.n1277 53.0052
R15589 gnd.n1280 gnd.n1279 53.0052
R15590 gnd.n1282 gnd.n1281 53.0052
R15591 gnd.n1284 gnd.n1283 53.0052
R15592 gnd.n1286 gnd.n1285 53.0052
R15593 gnd.n1288 gnd.n1287 53.0052
R15594 gnd.n1290 gnd.n1289 53.0052
R15595 gnd.n1294 gnd.n1293 53.0052
R15596 gnd.n1296 gnd.n1295 53.0052
R15597 gnd.n1298 gnd.n1297 53.0052
R15598 gnd.n1300 gnd.n1299 53.0052
R15599 gnd.n1302 gnd.n1301 53.0052
R15600 gnd.n1304 gnd.n1303 53.0052
R15601 gnd.n1306 gnd.n1305 53.0052
R15602 gnd.n1308 gnd.n1307 53.0052
R15603 gnd.n1310 gnd.n1309 53.0052
R15604 gnd.n92 gnd.n91 53.0052
R15605 gnd.n90 gnd.n89 53.0052
R15606 gnd.n88 gnd.n87 53.0052
R15607 gnd.n86 gnd.n85 53.0052
R15608 gnd.n84 gnd.n83 53.0052
R15609 gnd.n82 gnd.n81 53.0052
R15610 gnd.n80 gnd.n79 53.0052
R15611 gnd.n78 gnd.n77 53.0052
R15612 gnd.n76 gnd.n75 53.0052
R15613 gnd.n33 gnd.n32 53.0052
R15614 gnd.n31 gnd.n30 53.0052
R15615 gnd.n29 gnd.n28 53.0052
R15616 gnd.n27 gnd.n26 53.0052
R15617 gnd.n25 gnd.n24 53.0052
R15618 gnd.n23 gnd.n22 53.0052
R15619 gnd.n21 gnd.n20 53.0052
R15620 gnd.n19 gnd.n18 53.0052
R15621 gnd.n17 gnd.n16 53.0052
R15622 gnd.n52 gnd.n51 53.0052
R15623 gnd.n50 gnd.n49 53.0052
R15624 gnd.n48 gnd.n47 53.0052
R15625 gnd.n46 gnd.n45 53.0052
R15626 gnd.n44 gnd.n43 53.0052
R15627 gnd.n42 gnd.n41 53.0052
R15628 gnd.n40 gnd.n39 53.0052
R15629 gnd.n38 gnd.n37 53.0052
R15630 gnd.n36 gnd.n35 53.0052
R15631 gnd.n72 gnd.n71 53.0052
R15632 gnd.n70 gnd.n69 53.0052
R15633 gnd.n68 gnd.n67 53.0052
R15634 gnd.n66 gnd.n65 53.0052
R15635 gnd.n64 gnd.n63 53.0052
R15636 gnd.n62 gnd.n61 53.0052
R15637 gnd.n60 gnd.n59 53.0052
R15638 gnd.n58 gnd.n57 53.0052
R15639 gnd.n56 gnd.n55 53.0052
R15640 gnd.n3464 gnd.n3463 52.4801
R15641 gnd.n2308 gnd.t397 52.3082
R15642 gnd.n2276 gnd.t378 52.3082
R15643 gnd.n2244 gnd.t363 52.3082
R15644 gnd.n2213 gnd.t401 52.3082
R15645 gnd.n2181 gnd.t1 52.3082
R15646 gnd.n2149 gnd.t380 52.3082
R15647 gnd.n2117 gnd.t383 52.3082
R15648 gnd.n2086 gnd.t215 52.3082
R15649 gnd.n6745 gnd.n2394 51.6227
R15650 gnd.n2138 gnd.n2106 51.4173
R15651 gnd.n2202 gnd.n2201 50.455
R15652 gnd.n2170 gnd.n2169 50.455
R15653 gnd.n2138 gnd.n2137 50.455
R15654 gnd.n1570 gnd.n1569 45.1884
R15655 gnd.n1034 gnd.n1033 45.1884
R15656 gnd.n3480 gnd.n3479 44.3322
R15657 gnd.n2885 gnd.n2884 44.3189
R15658 gnd.n4566 gnd.n4565 42.2793
R15659 gnd.n6139 gnd.n6138 42.2793
R15660 gnd.n1571 gnd.n1570 42.2793
R15661 gnd.n1035 gnd.n1034 42.2793
R15662 gnd.n1497 gnd.n1496 42.2793
R15663 gnd.n1014 gnd.n1013 42.2793
R15664 gnd.n3955 gnd.n3954 42.2793
R15665 gnd.n6098 gnd.n3140 42.2793
R15666 gnd.n6061 gnd.n3163 42.2793
R15667 gnd.n6021 gnd.n6018 42.2793
R15668 gnd.n7856 gnd.n353 42.2793
R15669 gnd.n7898 gnd.n333 42.2793
R15670 gnd.n7940 gnd.n7939 42.2793
R15671 gnd.n7740 gnd.n7739 42.2793
R15672 gnd.n6709 gnd.n2417 42.2793
R15673 gnd.n6669 gnd.n2439 42.2793
R15674 gnd.n6629 gnd.n2461 42.2793
R15675 gnd.n4160 gnd.n4108 42.2793
R15676 gnd.n6411 gnd.n2823 42.2793
R15677 gnd.n4714 gnd.n4624 42.2793
R15678 gnd.n4665 gnd.n4637 42.2793
R15679 gnd.n3069 gnd.n3068 42.2793
R15680 gnd.n2883 gnd.n2882 41.6274
R15681 gnd.n3474 gnd.n3473 41.6274
R15682 gnd.n2892 gnd.n2891 40.8975
R15683 gnd.n3477 gnd.n3476 40.8975
R15684 gnd.n7005 gnd.n786 38.268
R15685 gnd.n6999 gnd.n786 38.268
R15686 gnd.n6999 gnd.n6998 38.268
R15687 gnd.n6998 gnd.n6997 38.268
R15688 gnd.n6997 gnd.n793 38.268
R15689 gnd.n6991 gnd.n793 38.268
R15690 gnd.n6991 gnd.n6990 38.268
R15691 gnd.n6990 gnd.n6989 38.268
R15692 gnd.n6989 gnd.n801 38.268
R15693 gnd.n6983 gnd.n801 38.268
R15694 gnd.n6983 gnd.n6982 38.268
R15695 gnd.n6982 gnd.n6981 38.268
R15696 gnd.n6981 gnd.n809 38.268
R15697 gnd.n6975 gnd.n809 38.268
R15698 gnd.n6975 gnd.n6974 38.268
R15699 gnd.n6974 gnd.n6973 38.268
R15700 gnd.n6973 gnd.n817 38.268
R15701 gnd.n6967 gnd.n817 38.268
R15702 gnd.n6967 gnd.n6966 38.268
R15703 gnd.n6966 gnd.n6965 38.268
R15704 gnd.n6965 gnd.n825 38.268
R15705 gnd.n6959 gnd.n825 38.268
R15706 gnd.n6959 gnd.n6958 38.268
R15707 gnd.n6958 gnd.n6957 38.268
R15708 gnd.n6957 gnd.n833 38.268
R15709 gnd.n6951 gnd.n833 38.268
R15710 gnd.n6951 gnd.n6950 38.268
R15711 gnd.n6950 gnd.n6949 38.268
R15712 gnd.n6949 gnd.n841 38.268
R15713 gnd.n6943 gnd.n841 38.268
R15714 gnd.n6943 gnd.n6942 38.268
R15715 gnd.n6942 gnd.n6941 38.268
R15716 gnd.n6941 gnd.n849 38.268
R15717 gnd.n6935 gnd.n849 38.268
R15718 gnd.n6935 gnd.n6934 38.268
R15719 gnd.n6934 gnd.n6933 38.268
R15720 gnd.n6933 gnd.n857 38.268
R15721 gnd.n6927 gnd.n857 38.268
R15722 gnd.n6927 gnd.n6926 38.268
R15723 gnd.n6926 gnd.n6925 38.268
R15724 gnd.n6925 gnd.n865 38.268
R15725 gnd.n6919 gnd.n865 38.268
R15726 gnd.n6919 gnd.n6918 38.268
R15727 gnd.n6918 gnd.n6917 38.268
R15728 gnd.n6917 gnd.n873 38.268
R15729 gnd.n6911 gnd.n873 38.268
R15730 gnd.n6911 gnd.n6910 38.268
R15731 gnd.n6910 gnd.n6909 38.268
R15732 gnd.n6909 gnd.n881 38.268
R15733 gnd.n6903 gnd.n881 38.268
R15734 gnd.n6903 gnd.n6902 38.268
R15735 gnd.n6902 gnd.n6901 38.268
R15736 gnd.n6901 gnd.n889 38.268
R15737 gnd.n6895 gnd.n889 38.268
R15738 gnd.n6895 gnd.n6894 38.268
R15739 gnd.n6894 gnd.n6893 38.268
R15740 gnd.n6893 gnd.n897 38.268
R15741 gnd.n6887 gnd.n897 38.268
R15742 gnd.n6887 gnd.n6886 38.268
R15743 gnd.n6886 gnd.n6885 38.268
R15744 gnd.n6885 gnd.n905 38.268
R15745 gnd.n6879 gnd.n905 38.268
R15746 gnd.n6879 gnd.n6878 38.268
R15747 gnd.n6878 gnd.n6877 38.268
R15748 gnd.n6877 gnd.n913 38.268
R15749 gnd.n6871 gnd.n913 38.268
R15750 gnd.n6871 gnd.n6870 38.268
R15751 gnd.n6870 gnd.n6869 38.268
R15752 gnd.n6869 gnd.n921 38.268
R15753 gnd.n6863 gnd.n921 38.268
R15754 gnd.n6863 gnd.n6862 38.268
R15755 gnd.n6862 gnd.n6861 38.268
R15756 gnd.n6861 gnd.n929 38.268
R15757 gnd.n6855 gnd.n929 38.268
R15758 gnd.n6855 gnd.n6854 38.268
R15759 gnd.n6854 gnd.n6853 38.268
R15760 gnd.n6853 gnd.n937 38.268
R15761 gnd.n6847 gnd.n937 38.268
R15762 gnd.n6847 gnd.n6846 38.268
R15763 gnd.n6846 gnd.n6845 38.268
R15764 gnd.n6845 gnd.n945 38.268
R15765 gnd.n6839 gnd.n945 38.268
R15766 gnd.n6839 gnd.n6838 38.268
R15767 gnd.n7973 gnd.n256 35.69
R15768 gnd.n2891 gnd.n2890 35.055
R15769 gnd.n2886 gnd.n2885 35.055
R15770 gnd.n3466 gnd.n3465 35.055
R15771 gnd.n3476 gnd.n3462 35.055
R15772 gnd.n1633 gnd.n1527 31.8661
R15773 gnd.n1633 gnd.n1632 31.8661
R15774 gnd.n1641 gnd.n1516 31.8661
R15775 gnd.n1649 gnd.n1516 31.8661
R15776 gnd.n1649 gnd.n1510 31.8661
R15777 gnd.n1657 gnd.n1510 31.8661
R15778 gnd.n1657 gnd.n1503 31.8661
R15779 gnd.n1695 gnd.n1503 31.8661
R15780 gnd.n1705 gnd.n1436 31.8661
R15781 gnd.n6621 gnd.n2394 31.8661
R15782 gnd.n6615 gnd.n2478 31.8661
R15783 gnd.n6615 gnd.n2481 31.8661
R15784 gnd.n6609 gnd.n2481 31.8661
R15785 gnd.n6609 gnd.n2493 31.8661
R15786 gnd.n6603 gnd.n2503 31.8661
R15787 gnd.n6597 gnd.n2503 31.8661
R15788 gnd.n6591 gnd.n2519 31.8661
R15789 gnd.n6591 gnd.n2522 31.8661
R15790 gnd.n6585 gnd.n2532 31.8661
R15791 gnd.n4763 gnd.n2765 31.8661
R15792 gnd.n3934 gnd.n2776 31.8661
R15793 gnd.n4774 gnd.n3934 31.8661
R15794 gnd.n4775 gnd.n4774 31.8661
R15795 gnd.n4775 gnd.n3927 31.8661
R15796 gnd.n4783 gnd.n3927 31.8661
R15797 gnd.n4808 gnd.n3918 31.8661
R15798 gnd.n4808 gnd.n3909 31.8661
R15799 gnd.n4825 gnd.n3909 31.8661
R15800 gnd.n4825 gnd.n3910 31.8661
R15801 gnd.n5561 gnd.n3434 31.8661
R15802 gnd.n5572 gnd.n3434 31.8661
R15803 gnd.n5572 gnd.n3427 31.8661
R15804 gnd.n5580 gnd.n3427 31.8661
R15805 gnd.n6202 gnd.n3006 31.8661
R15806 gnd.n6202 gnd.n3008 31.8661
R15807 gnd.n5682 gnd.n3008 31.8661
R15808 gnd.n5682 gnd.n3420 31.8661
R15809 gnd.n3420 gnd.n3075 31.8661
R15810 gnd.n3185 gnd.n3117 31.8661
R15811 gnd.n8017 gnd.n188 31.8661
R15812 gnd.n8011 gnd.n199 31.8661
R15813 gnd.n8011 gnd.n202 31.8661
R15814 gnd.n8005 gnd.n211 31.8661
R15815 gnd.n7999 gnd.n211 31.8661
R15816 gnd.n7993 gnd.n227 31.8661
R15817 gnd.n7993 gnd.n230 31.8661
R15818 gnd.n7987 gnd.n230 31.8661
R15819 gnd.n7987 gnd.n240 31.8661
R15820 gnd.n7981 gnd.n249 31.8661
R15821 gnd.n5423 gnd.n3533 30.4395
R15822 gnd.n3894 gnd.n3890 30.4395
R15823 gnd.n6621 gnd.t230 28.3609
R15824 gnd.n7981 gnd.t238 28.3609
R15825 gnd.n6444 gnd.n2776 27.4049
R15826 gnd.n6134 gnd.n3075 27.4049
R15827 gnd.n6390 gnd.n2871 25.8116
R15828 gnd.n5553 gnd.n3447 25.8116
R15829 gnd.n4565 gnd.n4564 25.7944
R15830 gnd.n6138 gnd.n6137 25.7944
R15831 gnd.n1496 gnd.n1495 25.7944
R15832 gnd.n1013 gnd.n1012 25.7944
R15833 gnd.n3954 gnd.n3953 25.7944
R15834 gnd.n3140 gnd.n3139 25.7944
R15835 gnd.n3163 gnd.n3162 25.7944
R15836 gnd.n6018 gnd.n6017 25.7944
R15837 gnd.n353 gnd.n352 25.7944
R15838 gnd.n333 gnd.n332 25.7944
R15839 gnd.n7939 gnd.n7938 25.7944
R15840 gnd.n7739 gnd.n7738 25.7944
R15841 gnd.n2417 gnd.n2416 25.7944
R15842 gnd.n2439 gnd.n2438 25.7944
R15843 gnd.n2461 gnd.n2460 25.7944
R15844 gnd.n4108 gnd.n4107 25.7944
R15845 gnd.n2823 gnd.n2822 25.7944
R15846 gnd.n4624 gnd.n4623 25.7944
R15847 gnd.n4637 gnd.n4636 25.7944
R15848 gnd.n3068 gnd.n3067 25.7944
R15849 gnd.n1717 gnd.n1437 24.8557
R15850 gnd.n1727 gnd.n1420 24.8557
R15851 gnd.n1423 gnd.n1411 24.8557
R15852 gnd.n1748 gnd.n1412 24.8557
R15853 gnd.n1758 gnd.n1392 24.8557
R15854 gnd.n1768 gnd.n1767 24.8557
R15855 gnd.n1376 gnd.n1375 24.8557
R15856 gnd.n1805 gnd.n1368 24.8557
R15857 gnd.n1804 gnd.n1361 24.8557
R15858 gnd.n1842 gnd.n1340 24.8557
R15859 gnd.n1816 gnd.n1341 24.8557
R15860 gnd.n1835 gnd.n1240 24.8557
R15861 gnd.n1852 gnd.n1851 24.8557
R15862 gnd.n1862 gnd.n1861 24.8557
R15863 gnd.n1231 gnd.n1223 24.8557
R15864 gnd.n1892 gnd.n1891 24.8557
R15865 gnd.n1902 gnd.n1201 24.8557
R15866 gnd.n1914 gnd.n1190 24.8557
R15867 gnd.n1905 gnd.n1183 24.8557
R15868 gnd.n1941 gnd.n1940 24.8557
R15869 gnd.n1951 gnd.n1176 24.8557
R15870 gnd.n1963 gnd.n1168 24.8557
R15871 gnd.n1981 gnd.n1980 24.8557
R15872 gnd.n1926 gnd.n1159 24.8557
R15873 gnd.n1991 gnd.n1149 24.8557
R15874 gnd.n2004 gnd.n1138 24.8557
R15875 gnd.n2042 gnd.n2041 24.8557
R15876 gnd.n2057 gnd.n1123 24.8557
R15877 gnd.n6830 gnd.n964 24.8557
R15878 gnd.n6829 gnd.n967 24.8557
R15879 gnd.n6823 gnd.n6822 24.8557
R15880 gnd.n2022 gnd.n979 24.8557
R15881 gnd.n6816 gnd.n988 24.8557
R15882 gnd.n6809 gnd.n6808 24.8557
R15883 gnd.n3828 gnd.n3827 23.855
R15884 gnd.n3511 gnd.n3510 23.855
R15885 gnd.n6326 gnd.n6325 23.855
R15886 gnd.n3505 gnd.n3504 23.855
R15887 gnd.n1738 gnd.t214 23.2624
R15888 gnd.t25 gnd.n2493 23.2624
R15889 gnd.n227 gnd.t50 23.2624
R15890 gnd.n6838 gnd.n6837 22.961
R15891 gnd.n1439 gnd.t275 22.6251
R15892 gnd.n2529 gnd.t33 22.3064
R15893 gnd.t114 gnd.n191 22.3064
R15894 gnd.n6320 gnd.n6319 21.6691
R15895 gnd.n5031 gnd.n3809 21.6691
R15896 gnd.n5058 gnd.n3792 21.6691
R15897 gnd.n5083 gnd.n3776 21.6691
R15898 gnd.n5107 gnd.n3756 21.6691
R15899 gnd.n5129 gnd.n5128 21.6691
R15900 gnd.n5149 gnd.n3733 21.6691
R15901 gnd.n5155 gnd.n3729 21.6691
R15902 gnd.n5182 gnd.n3711 21.6691
R15903 gnd.n5207 gnd.n3695 21.6691
R15904 gnd.n5207 gnd.n3688 21.6691
R15905 gnd.n5230 gnd.n3675 21.6691
R15906 gnd.n5251 gnd.n5250 21.6691
R15907 gnd.n5270 gnd.n3650 21.6691
R15908 gnd.n5276 gnd.n3646 21.6691
R15909 gnd.n5300 gnd.n3629 21.6691
R15910 gnd.n5323 gnd.n3610 21.6691
R15911 gnd.n5352 gnd.n3582 21.6691
R15912 gnd.n5367 gnd.n3572 21.6691
R15913 gnd.n5386 gnd.n3537 21.6691
R15914 gnd.n5544 gnd.n3457 21.6691
R15915 gnd.t400 gnd.n1444 21.3504
R15916 gnd.n2035 gnd.t5 20.7131
R15917 gnd.t366 gnd.n2839 20.7131
R15918 gnd.n3446 gnd.t370 20.7131
R15919 gnd.n3892 gnd.n2897 20.3945
R15920 gnd.t323 gnd.n3818 20.3945
R15921 gnd.n5071 gnd.n3781 20.3945
R15922 gnd.n5089 gnd.n3771 20.3945
R15923 gnd.n5195 gnd.n3702 20.3945
R15924 gnd.n5213 gnd.n3691 20.3945
R15925 gnd.n5315 gnd.n3618 20.3945
R15926 gnd.n5334 gnd.n5333 20.3945
R15927 gnd.t3 gnd.n1156 20.0758
R15928 gnd.n2880 gnd.t299 19.8005
R15929 gnd.n2880 gnd.t270 19.8005
R15930 gnd.n2879 gnd.t324 19.8005
R15931 gnd.n2879 gnd.t249 19.8005
R15932 gnd.n3471 gnd.t263 19.8005
R15933 gnd.n3471 gnd.t293 19.8005
R15934 gnd.n3470 gnd.t243 19.8005
R15935 gnd.n3470 gnd.t315 19.8005
R15936 gnd.n2876 gnd.n2875 19.5087
R15937 gnd.n2889 gnd.n2876 19.5087
R15938 gnd.n2887 gnd.n2878 19.5087
R15939 gnd.n3475 gnd.n3469 19.5087
R15940 gnd.t374 gnd.n1200 19.4385
R15941 gnd.n2519 gnd.t37 19.4385
R15942 gnd.t124 gnd.n202 19.4385
R15943 gnd.n4785 gnd.n3925 19.3944
R15944 gnd.n4785 gnd.n3922 19.3944
R15945 gnd.n4806 gnd.n3922 19.3944
R15946 gnd.n4806 gnd.n3923 19.3944
R15947 gnd.n4802 gnd.n3923 19.3944
R15948 gnd.n4802 gnd.n4801 19.3944
R15949 gnd.n4801 gnd.n4800 19.3944
R15950 gnd.n4800 gnd.n4791 19.3944
R15951 gnd.n4796 gnd.n4791 19.3944
R15952 gnd.n4796 gnd.n4795 19.3944
R15953 gnd.n4795 gnd.n2915 19.3944
R15954 gnd.n6310 gnd.n2915 19.3944
R15955 gnd.n6310 gnd.n2916 19.3944
R15956 gnd.n6306 gnd.n2916 19.3944
R15957 gnd.n6306 gnd.n6305 19.3944
R15958 gnd.n6305 gnd.n6304 19.3944
R15959 gnd.n6304 gnd.n2922 19.3944
R15960 gnd.n6300 gnd.n2922 19.3944
R15961 gnd.n6300 gnd.n6299 19.3944
R15962 gnd.n6299 gnd.n6298 19.3944
R15963 gnd.n6298 gnd.n2927 19.3944
R15964 gnd.n6294 gnd.n2927 19.3944
R15965 gnd.n6294 gnd.n6293 19.3944
R15966 gnd.n6293 gnd.n6292 19.3944
R15967 gnd.n6292 gnd.n2932 19.3944
R15968 gnd.n6288 gnd.n2932 19.3944
R15969 gnd.n6288 gnd.n6287 19.3944
R15970 gnd.n6287 gnd.n6286 19.3944
R15971 gnd.n6286 gnd.n2937 19.3944
R15972 gnd.n6282 gnd.n2937 19.3944
R15973 gnd.n6282 gnd.n6281 19.3944
R15974 gnd.n6281 gnd.n6280 19.3944
R15975 gnd.n6280 gnd.n2942 19.3944
R15976 gnd.n6276 gnd.n2942 19.3944
R15977 gnd.n6276 gnd.n6275 19.3944
R15978 gnd.n6275 gnd.n6274 19.3944
R15979 gnd.n6274 gnd.n2947 19.3944
R15980 gnd.n6270 gnd.n2947 19.3944
R15981 gnd.n6270 gnd.n6269 19.3944
R15982 gnd.n6269 gnd.n6268 19.3944
R15983 gnd.n6268 gnd.n2952 19.3944
R15984 gnd.n6264 gnd.n2952 19.3944
R15985 gnd.n6264 gnd.n6263 19.3944
R15986 gnd.n6263 gnd.n6262 19.3944
R15987 gnd.n6262 gnd.n2957 19.3944
R15988 gnd.n6258 gnd.n2957 19.3944
R15989 gnd.n6258 gnd.n6257 19.3944
R15990 gnd.n6257 gnd.n6256 19.3944
R15991 gnd.n6256 gnd.n2962 19.3944
R15992 gnd.n6252 gnd.n2962 19.3944
R15993 gnd.n6252 gnd.n6251 19.3944
R15994 gnd.n6251 gnd.n6250 19.3944
R15995 gnd.n6250 gnd.n2967 19.3944
R15996 gnd.n6246 gnd.n2967 19.3944
R15997 gnd.n6246 gnd.n6245 19.3944
R15998 gnd.n6245 gnd.n6244 19.3944
R15999 gnd.n6244 gnd.n2972 19.3944
R16000 gnd.n6240 gnd.n2972 19.3944
R16001 gnd.n6240 gnd.n6239 19.3944
R16002 gnd.n6239 gnd.n6238 19.3944
R16003 gnd.n6238 gnd.n2977 19.3944
R16004 gnd.n6234 gnd.n2977 19.3944
R16005 gnd.n6234 gnd.n6233 19.3944
R16006 gnd.n6233 gnd.n6232 19.3944
R16007 gnd.n6232 gnd.n2982 19.3944
R16008 gnd.n6228 gnd.n2982 19.3944
R16009 gnd.n6228 gnd.n6227 19.3944
R16010 gnd.n6227 gnd.n6226 19.3944
R16011 gnd.n6226 gnd.n2987 19.3944
R16012 gnd.n6222 gnd.n2987 19.3944
R16013 gnd.n6222 gnd.n6221 19.3944
R16014 gnd.n6221 gnd.n6220 19.3944
R16015 gnd.n6220 gnd.n2992 19.3944
R16016 gnd.n6216 gnd.n2992 19.3944
R16017 gnd.n6216 gnd.n6215 19.3944
R16018 gnd.n6215 gnd.n6214 19.3944
R16019 gnd.n6214 gnd.n2997 19.3944
R16020 gnd.n6210 gnd.n2997 19.3944
R16021 gnd.n6210 gnd.n6209 19.3944
R16022 gnd.n6209 gnd.n6208 19.3944
R16023 gnd.n6208 gnd.n3002 19.3944
R16024 gnd.n6204 gnd.n3002 19.3944
R16025 gnd.n4570 gnd.n4569 19.3944
R16026 gnd.n4569 gnd.n3950 19.3944
R16027 gnd.n4772 gnd.n3950 19.3944
R16028 gnd.n4495 gnd.n4494 19.3944
R16029 gnd.n4498 gnd.n4495 19.3944
R16030 gnd.n4498 gnd.n4478 19.3944
R16031 gnd.n4502 gnd.n4478 19.3944
R16032 gnd.n4503 gnd.n4502 19.3944
R16033 gnd.n4619 gnd.n4503 19.3944
R16034 gnd.n4619 gnd.n4618 19.3944
R16035 gnd.n4618 gnd.n4617 19.3944
R16036 gnd.n4617 gnd.n4508 19.3944
R16037 gnd.n4610 gnd.n4508 19.3944
R16038 gnd.n4610 gnd.n4609 19.3944
R16039 gnd.n4609 gnd.n4517 19.3944
R16040 gnd.n4602 gnd.n4517 19.3944
R16041 gnd.n4602 gnd.n4601 19.3944
R16042 gnd.n4601 gnd.n4527 19.3944
R16043 gnd.n4594 gnd.n4527 19.3944
R16044 gnd.n4594 gnd.n4593 19.3944
R16045 gnd.n4593 gnd.n4537 19.3944
R16046 gnd.n4586 gnd.n4537 19.3944
R16047 gnd.n4586 gnd.n4585 19.3944
R16048 gnd.n4585 gnd.n4547 19.3944
R16049 gnd.n4578 gnd.n4547 19.3944
R16050 gnd.n4578 gnd.n4577 19.3944
R16051 gnd.n4577 gnd.n4557 19.3944
R16052 gnd.n6180 gnd.n3028 19.3944
R16053 gnd.n6180 gnd.n6179 19.3944
R16054 gnd.n6179 gnd.n3031 19.3944
R16055 gnd.n6172 gnd.n3031 19.3944
R16056 gnd.n6172 gnd.n6171 19.3944
R16057 gnd.n6171 gnd.n3039 19.3944
R16058 gnd.n6164 gnd.n3039 19.3944
R16059 gnd.n6164 gnd.n6163 19.3944
R16060 gnd.n6163 gnd.n3047 19.3944
R16061 gnd.n6156 gnd.n3047 19.3944
R16062 gnd.n6156 gnd.n6155 19.3944
R16063 gnd.n6155 gnd.n3055 19.3944
R16064 gnd.n6148 gnd.n3055 19.3944
R16065 gnd.n6148 gnd.n6147 19.3944
R16066 gnd.n6147 gnd.n3063 19.3944
R16067 gnd.n6140 gnd.n3063 19.3944
R16068 gnd.n1620 gnd.n1619 19.3944
R16069 gnd.n1619 gnd.n1618 19.3944
R16070 gnd.n1618 gnd.n1617 19.3944
R16071 gnd.n1617 gnd.n1615 19.3944
R16072 gnd.n1615 gnd.n1612 19.3944
R16073 gnd.n1612 gnd.n1611 19.3944
R16074 gnd.n1611 gnd.n1608 19.3944
R16075 gnd.n1608 gnd.n1607 19.3944
R16076 gnd.n1607 gnd.n1604 19.3944
R16077 gnd.n1604 gnd.n1603 19.3944
R16078 gnd.n1603 gnd.n1600 19.3944
R16079 gnd.n1600 gnd.n1599 19.3944
R16080 gnd.n1599 gnd.n1596 19.3944
R16081 gnd.n1596 gnd.n1595 19.3944
R16082 gnd.n1595 gnd.n1592 19.3944
R16083 gnd.n1592 gnd.n1591 19.3944
R16084 gnd.n1591 gnd.n1588 19.3944
R16085 gnd.n1588 gnd.n1587 19.3944
R16086 gnd.n1587 gnd.n1584 19.3944
R16087 gnd.n1584 gnd.n1583 19.3944
R16088 gnd.n1583 gnd.n1580 19.3944
R16089 gnd.n1580 gnd.n1579 19.3944
R16090 gnd.n1576 gnd.n1575 19.3944
R16091 gnd.n1575 gnd.n1531 19.3944
R16092 gnd.n1626 gnd.n1531 19.3944
R16093 gnd.n1107 gnd.n1105 19.3944
R16094 gnd.n1107 gnd.n1031 19.3944
R16095 gnd.n2353 gnd.n1031 19.3944
R16096 gnd.n1048 gnd.n1047 19.3944
R16097 gnd.n1052 gnd.n1047 19.3944
R16098 gnd.n1055 gnd.n1052 19.3944
R16099 gnd.n1058 gnd.n1055 19.3944
R16100 gnd.n1058 gnd.n1044 19.3944
R16101 gnd.n1062 gnd.n1044 19.3944
R16102 gnd.n1065 gnd.n1062 19.3944
R16103 gnd.n1068 gnd.n1065 19.3944
R16104 gnd.n1068 gnd.n1042 19.3944
R16105 gnd.n1072 gnd.n1042 19.3944
R16106 gnd.n1075 gnd.n1072 19.3944
R16107 gnd.n1078 gnd.n1075 19.3944
R16108 gnd.n1078 gnd.n1040 19.3944
R16109 gnd.n1082 gnd.n1040 19.3944
R16110 gnd.n1085 gnd.n1082 19.3944
R16111 gnd.n1088 gnd.n1085 19.3944
R16112 gnd.n1088 gnd.n1038 19.3944
R16113 gnd.n1092 gnd.n1038 19.3944
R16114 gnd.n1095 gnd.n1092 19.3944
R16115 gnd.n1098 gnd.n1095 19.3944
R16116 gnd.n1098 gnd.n1036 19.3944
R16117 gnd.n1102 gnd.n1036 19.3944
R16118 gnd.n1719 gnd.n1428 19.3944
R16119 gnd.n1729 gnd.n1428 19.3944
R16120 gnd.n1730 gnd.n1729 19.3944
R16121 gnd.n1730 gnd.n1409 19.3944
R16122 gnd.n1750 gnd.n1409 19.3944
R16123 gnd.n1750 gnd.n1401 19.3944
R16124 gnd.n1760 gnd.n1401 19.3944
R16125 gnd.n1761 gnd.n1760 19.3944
R16126 gnd.n1762 gnd.n1761 19.3944
R16127 gnd.n1762 gnd.n1384 19.3944
R16128 gnd.n1384 gnd.n1382 19.3944
R16129 gnd.n1788 gnd.n1382 19.3944
R16130 gnd.n1788 gnd.n1364 19.3944
R16131 gnd.n1822 gnd.n1364 19.3944
R16132 gnd.n1822 gnd.n1821 19.3944
R16133 gnd.n1821 gnd.n1820 19.3944
R16134 gnd.n1820 gnd.n1815 19.3944
R16135 gnd.n1815 gnd.n1236 19.3944
R16136 gnd.n1854 gnd.n1236 19.3944
R16137 gnd.n1855 gnd.n1854 19.3944
R16138 gnd.n1856 gnd.n1855 19.3944
R16139 gnd.n1856 gnd.n1222 19.3944
R16140 gnd.n1222 gnd.n1216 19.3944
R16141 gnd.n1881 gnd.n1216 19.3944
R16142 gnd.n1882 gnd.n1881 19.3944
R16143 gnd.n1882 gnd.n1199 19.3944
R16144 gnd.n1199 gnd.n1197 19.3944
R16145 gnd.n1907 gnd.n1197 19.3944
R16146 gnd.n1908 gnd.n1907 19.3944
R16147 gnd.n1908 gnd.n1171 19.3944
R16148 gnd.n1958 gnd.n1171 19.3944
R16149 gnd.n1959 gnd.n1958 19.3944
R16150 gnd.n1959 gnd.n1164 19.3944
R16151 gnd.n1970 gnd.n1164 19.3944
R16152 gnd.n1971 gnd.n1970 19.3944
R16153 gnd.n1971 gnd.n1148 19.3944
R16154 gnd.n1148 gnd.n1146 19.3944
R16155 gnd.n1995 gnd.n1146 19.3944
R16156 gnd.n1998 gnd.n1995 19.3944
R16157 gnd.n1998 gnd.n1997 19.3944
R16158 gnd.n1997 gnd.n1119 19.3944
R16159 gnd.n2064 gnd.n1119 19.3944
R16160 gnd.n2064 gnd.n1116 19.3944
R16161 gnd.n2068 gnd.n1116 19.3944
R16162 gnd.n2069 gnd.n2068 19.3944
R16163 gnd.n2069 gnd.n1114 19.3944
R16164 gnd.n2075 gnd.n1114 19.3944
R16165 gnd.n2333 gnd.n2075 19.3944
R16166 gnd.n2337 gnd.n2333 19.3944
R16167 gnd.n2338 gnd.n2337 19.3944
R16168 gnd.n2343 gnd.n2338 19.3944
R16169 gnd.n2343 gnd.n1010 19.3944
R16170 gnd.n6803 gnd.n1010 19.3944
R16171 gnd.n1710 gnd.n1709 19.3944
R16172 gnd.n1709 gnd.n1442 19.3944
R16173 gnd.n1465 gnd.n1442 19.3944
R16174 gnd.n1468 gnd.n1465 19.3944
R16175 gnd.n1468 gnd.n1461 19.3944
R16176 gnd.n1472 gnd.n1461 19.3944
R16177 gnd.n1475 gnd.n1472 19.3944
R16178 gnd.n1478 gnd.n1475 19.3944
R16179 gnd.n1478 gnd.n1459 19.3944
R16180 gnd.n1482 gnd.n1459 19.3944
R16181 gnd.n1485 gnd.n1482 19.3944
R16182 gnd.n1488 gnd.n1485 19.3944
R16183 gnd.n1488 gnd.n1457 19.3944
R16184 gnd.n1492 gnd.n1457 19.3944
R16185 gnd.n1715 gnd.n1714 19.3944
R16186 gnd.n1714 gnd.n1418 19.3944
R16187 gnd.n1740 gnd.n1418 19.3944
R16188 gnd.n1740 gnd.n1416 19.3944
R16189 gnd.n1746 gnd.n1416 19.3944
R16190 gnd.n1746 gnd.n1745 19.3944
R16191 gnd.n1745 gnd.n1390 19.3944
R16192 gnd.n1770 gnd.n1390 19.3944
R16193 gnd.n1770 gnd.n1388 19.3944
R16194 gnd.n1782 gnd.n1388 19.3944
R16195 gnd.n1782 gnd.n1781 19.3944
R16196 gnd.n1781 gnd.n1780 19.3944
R16197 gnd.n1780 gnd.n1778 19.3944
R16198 gnd.n1778 gnd.n1360 19.3944
R16199 gnd.n1360 gnd.n1358 19.3944
R16200 gnd.n1829 gnd.n1358 19.3944
R16201 gnd.n1829 gnd.n1356 19.3944
R16202 gnd.n1833 gnd.n1356 19.3944
R16203 gnd.n1833 gnd.n1227 19.3944
R16204 gnd.n1864 gnd.n1227 19.3944
R16205 gnd.n1864 gnd.n1225 19.3944
R16206 gnd.n1868 gnd.n1225 19.3944
R16207 gnd.n1868 gnd.n1206 19.3944
R16208 gnd.n1894 gnd.n1206 19.3944
R16209 gnd.n1894 gnd.n1204 19.3944
R16210 gnd.n1900 gnd.n1204 19.3944
R16211 gnd.n1900 gnd.n1899 19.3944
R16212 gnd.n1899 gnd.n1181 19.3944
R16213 gnd.n1943 gnd.n1181 19.3944
R16214 gnd.n1943 gnd.n1179 19.3944
R16215 gnd.n1949 gnd.n1179 19.3944
R16216 gnd.n1949 gnd.n1948 19.3944
R16217 gnd.n1948 gnd.n1154 19.3944
R16218 gnd.n1983 gnd.n1154 19.3944
R16219 gnd.n1983 gnd.n1152 19.3944
R16220 gnd.n1989 gnd.n1152 19.3944
R16221 gnd.n1989 gnd.n1988 19.3944
R16222 gnd.n1988 gnd.n1129 19.3944
R16223 gnd.n2044 gnd.n1129 19.3944
R16224 gnd.n2044 gnd.n1127 19.3944
R16225 gnd.n2054 gnd.n1127 19.3944
R16226 gnd.n2054 gnd.n2053 19.3944
R16227 gnd.n2053 gnd.n2052 19.3944
R16228 gnd.n2052 gnd.n970 19.3944
R16229 gnd.n6827 gnd.n970 19.3944
R16230 gnd.n6827 gnd.n6826 19.3944
R16231 gnd.n6826 gnd.n6825 19.3944
R16232 gnd.n6825 gnd.n974 19.3944
R16233 gnd.n993 gnd.n974 19.3944
R16234 gnd.n6813 gnd.n993 19.3944
R16235 gnd.n6813 gnd.n6812 19.3944
R16236 gnd.n6812 gnd.n6811 19.3944
R16237 gnd.n6811 gnd.n999 19.3944
R16238 gnd.n6790 gnd.n6789 19.3944
R16239 gnd.n6789 gnd.n6755 19.3944
R16240 gnd.n6785 gnd.n6755 19.3944
R16241 gnd.n6785 gnd.n6782 19.3944
R16242 gnd.n6782 gnd.n6779 19.3944
R16243 gnd.n6779 gnd.n6778 19.3944
R16244 gnd.n6778 gnd.n6775 19.3944
R16245 gnd.n6775 gnd.n6774 19.3944
R16246 gnd.n6774 gnd.n6771 19.3944
R16247 gnd.n6771 gnd.n6770 19.3944
R16248 gnd.n6770 gnd.n6767 19.3944
R16249 gnd.n6767 gnd.n6766 19.3944
R16250 gnd.n6766 gnd.n1016 19.3944
R16251 gnd.n6796 gnd.n1016 19.3944
R16252 gnd.n1630 gnd.n1529 19.3944
R16253 gnd.n1630 gnd.n1520 19.3944
R16254 gnd.n1643 gnd.n1520 19.3944
R16255 gnd.n1643 gnd.n1518 19.3944
R16256 gnd.n1647 gnd.n1518 19.3944
R16257 gnd.n1647 gnd.n1508 19.3944
R16258 gnd.n1659 gnd.n1508 19.3944
R16259 gnd.n1659 gnd.n1506 19.3944
R16260 gnd.n1693 gnd.n1506 19.3944
R16261 gnd.n1693 gnd.n1692 19.3944
R16262 gnd.n1692 gnd.n1691 19.3944
R16263 gnd.n1691 gnd.n1690 19.3944
R16264 gnd.n1690 gnd.n1687 19.3944
R16265 gnd.n1687 gnd.n1686 19.3944
R16266 gnd.n1686 gnd.n1685 19.3944
R16267 gnd.n1685 gnd.n1683 19.3944
R16268 gnd.n1683 gnd.n1682 19.3944
R16269 gnd.n1682 gnd.n1679 19.3944
R16270 gnd.n1679 gnd.n1678 19.3944
R16271 gnd.n1678 gnd.n1677 19.3944
R16272 gnd.n1677 gnd.n1675 19.3944
R16273 gnd.n1675 gnd.n1373 19.3944
R16274 gnd.n1796 gnd.n1373 19.3944
R16275 gnd.n1796 gnd.n1371 19.3944
R16276 gnd.n1802 gnd.n1371 19.3944
R16277 gnd.n1802 gnd.n1801 19.3944
R16278 gnd.n1801 gnd.n1336 19.3944
R16279 gnd.n1844 gnd.n1336 19.3944
R16280 gnd.n1844 gnd.n1337 19.3944
R16281 gnd.n1353 gnd.n1352 19.3944
R16282 gnd.n1849 gnd.n1848 19.3944
R16283 gnd.n1252 gnd.n1244 19.3944
R16284 gnd.n1251 gnd.n1249 19.3944
R16285 gnd.n1249 gnd.n1248 19.3944
R16286 gnd.n1248 gnd.n1188 19.3944
R16287 gnd.n1916 gnd.n1188 19.3944
R16288 gnd.n1916 gnd.n1186 19.3944
R16289 gnd.n1936 gnd.n1186 19.3944
R16290 gnd.n1936 gnd.n1935 19.3944
R16291 gnd.n1935 gnd.n1934 19.3944
R16292 gnd.n1934 gnd.n1932 19.3944
R16293 gnd.n1932 gnd.n1931 19.3944
R16294 gnd.n1931 gnd.n1929 19.3944
R16295 gnd.n1929 gnd.n1928 19.3944
R16296 gnd.n1928 gnd.n1136 19.3944
R16297 gnd.n2006 gnd.n1136 19.3944
R16298 gnd.n2006 gnd.n1134 19.3944
R16299 gnd.n2039 gnd.n1134 19.3944
R16300 gnd.n2039 gnd.n2038 19.3944
R16301 gnd.n2038 gnd.n2037 19.3944
R16302 gnd.n2037 gnd.n2034 19.3944
R16303 gnd.n2034 gnd.n2033 19.3944
R16304 gnd.n2033 gnd.n2030 19.3944
R16305 gnd.n2030 gnd.n2029 19.3944
R16306 gnd.n2029 gnd.n2026 19.3944
R16307 gnd.n2026 gnd.n2025 19.3944
R16308 gnd.n2025 gnd.n2024 19.3944
R16309 gnd.n2024 gnd.n2021 19.3944
R16310 gnd.n2021 gnd.n1111 19.3944
R16311 gnd.n2349 gnd.n1111 19.3944
R16312 gnd.n2350 gnd.n2349 19.3944
R16313 gnd.n1635 gnd.n1525 19.3944
R16314 gnd.n1635 gnd.n1523 19.3944
R16315 gnd.n1639 gnd.n1523 19.3944
R16316 gnd.n1639 gnd.n1514 19.3944
R16317 gnd.n1651 gnd.n1514 19.3944
R16318 gnd.n1651 gnd.n1512 19.3944
R16319 gnd.n1655 gnd.n1512 19.3944
R16320 gnd.n1655 gnd.n1501 19.3944
R16321 gnd.n1697 gnd.n1501 19.3944
R16322 gnd.n1697 gnd.n1455 19.3944
R16323 gnd.n1703 gnd.n1455 19.3944
R16324 gnd.n1703 gnd.n1702 19.3944
R16325 gnd.n1702 gnd.n1433 19.3944
R16326 gnd.n1724 gnd.n1433 19.3944
R16327 gnd.n1724 gnd.n1426 19.3944
R16328 gnd.n1735 gnd.n1426 19.3944
R16329 gnd.n1735 gnd.n1734 19.3944
R16330 gnd.n1734 gnd.n1407 19.3944
R16331 gnd.n1755 gnd.n1407 19.3944
R16332 gnd.n1755 gnd.n1397 19.3944
R16333 gnd.n1765 gnd.n1397 19.3944
R16334 gnd.n1765 gnd.n1378 19.3944
R16335 gnd.n1792 gnd.n1378 19.3944
R16336 gnd.n1792 gnd.n1791 19.3944
R16337 gnd.n1791 gnd.n1366 19.3944
R16338 gnd.n1808 gnd.n1366 19.3944
R16339 gnd.n1808 gnd.n1344 19.3944
R16340 gnd.n1840 gnd.n1344 19.3944
R16341 gnd.n1840 gnd.n1839 19.3944
R16342 gnd.n1839 gnd.n1838 19.3944
R16343 gnd.n1838 gnd.n1350 19.3944
R16344 gnd.n1350 gnd.n1233 19.3944
R16345 gnd.n1859 gnd.n1233 19.3944
R16346 gnd.n1859 gnd.n1218 19.3944
R16347 gnd.n1876 gnd.n1218 19.3944
R16348 gnd.n1876 gnd.n1214 19.3944
R16349 gnd.n1889 gnd.n1214 19.3944
R16350 gnd.n1889 gnd.n1888 19.3944
R16351 gnd.n1888 gnd.n1193 19.3944
R16352 gnd.n1912 gnd.n1193 19.3944
R16353 gnd.n1912 gnd.n1911 19.3944
R16354 gnd.n1911 gnd.n1173 19.3944
R16355 gnd.n1954 gnd.n1173 19.3944
R16356 gnd.n1954 gnd.n1166 19.3944
R16357 gnd.n1965 gnd.n1166 19.3944
R16358 gnd.n1965 gnd.n1162 19.3944
R16359 gnd.n1978 gnd.n1162 19.3944
R16360 gnd.n1978 gnd.n1977 19.3944
R16361 gnd.n1977 gnd.n1142 19.3944
R16362 gnd.n2002 gnd.n1142 19.3944
R16363 gnd.n2002 gnd.n2001 19.3944
R16364 gnd.n2001 gnd.n1121 19.3944
R16365 gnd.n2059 gnd.n1121 19.3944
R16366 gnd.n2059 gnd.n958 19.3944
R16367 gnd.n6834 gnd.n958 19.3944
R16368 gnd.n6834 gnd.n6833 19.3944
R16369 gnd.n6833 gnd.n6832 19.3944
R16370 gnd.n6832 gnd.n962 19.3944
R16371 gnd.n982 gnd.n962 19.3944
R16372 gnd.n6820 gnd.n982 19.3944
R16373 gnd.n6820 gnd.n6819 19.3944
R16374 gnd.n6819 gnd.n6818 19.3944
R16375 gnd.n6818 gnd.n986 19.3944
R16376 gnd.n1007 gnd.n986 19.3944
R16377 gnd.n6806 gnd.n1007 19.3944
R16378 gnd.n4614 gnd.n4613 19.3944
R16379 gnd.n4613 gnd.n4511 19.3944
R16380 gnd.n4606 gnd.n4511 19.3944
R16381 gnd.n4606 gnd.n4605 19.3944
R16382 gnd.n4605 gnd.n4523 19.3944
R16383 gnd.n4598 gnd.n4523 19.3944
R16384 gnd.n4598 gnd.n4597 19.3944
R16385 gnd.n4597 gnd.n4531 19.3944
R16386 gnd.n4590 gnd.n4531 19.3944
R16387 gnd.n4590 gnd.n4589 19.3944
R16388 gnd.n4589 gnd.n4543 19.3944
R16389 gnd.n4582 gnd.n4543 19.3944
R16390 gnd.n4582 gnd.n4581 19.3944
R16391 gnd.n4581 gnd.n4551 19.3944
R16392 gnd.n4574 gnd.n4551 19.3944
R16393 gnd.n4574 gnd.n4573 19.3944
R16394 gnd.n7494 gnd.n491 19.3944
R16395 gnd.n7500 gnd.n491 19.3944
R16396 gnd.n7500 gnd.n489 19.3944
R16397 gnd.n7504 gnd.n489 19.3944
R16398 gnd.n7504 gnd.n485 19.3944
R16399 gnd.n7510 gnd.n485 19.3944
R16400 gnd.n7510 gnd.n483 19.3944
R16401 gnd.n7514 gnd.n483 19.3944
R16402 gnd.n7514 gnd.n479 19.3944
R16403 gnd.n7520 gnd.n479 19.3944
R16404 gnd.n7520 gnd.n477 19.3944
R16405 gnd.n7524 gnd.n477 19.3944
R16406 gnd.n7524 gnd.n473 19.3944
R16407 gnd.n7530 gnd.n473 19.3944
R16408 gnd.n7530 gnd.n471 19.3944
R16409 gnd.n7534 gnd.n471 19.3944
R16410 gnd.n7534 gnd.n467 19.3944
R16411 gnd.n7540 gnd.n467 19.3944
R16412 gnd.n7540 gnd.n465 19.3944
R16413 gnd.n7544 gnd.n465 19.3944
R16414 gnd.n7544 gnd.n461 19.3944
R16415 gnd.n7550 gnd.n461 19.3944
R16416 gnd.n7550 gnd.n459 19.3944
R16417 gnd.n7554 gnd.n459 19.3944
R16418 gnd.n7554 gnd.n455 19.3944
R16419 gnd.n7560 gnd.n455 19.3944
R16420 gnd.n7560 gnd.n453 19.3944
R16421 gnd.n7564 gnd.n453 19.3944
R16422 gnd.n7564 gnd.n449 19.3944
R16423 gnd.n7570 gnd.n449 19.3944
R16424 gnd.n7570 gnd.n447 19.3944
R16425 gnd.n7574 gnd.n447 19.3944
R16426 gnd.n7574 gnd.n443 19.3944
R16427 gnd.n7580 gnd.n443 19.3944
R16428 gnd.n7580 gnd.n441 19.3944
R16429 gnd.n7584 gnd.n441 19.3944
R16430 gnd.n7584 gnd.n437 19.3944
R16431 gnd.n7590 gnd.n437 19.3944
R16432 gnd.n7590 gnd.n435 19.3944
R16433 gnd.n7594 gnd.n435 19.3944
R16434 gnd.n7594 gnd.n431 19.3944
R16435 gnd.n7600 gnd.n431 19.3944
R16436 gnd.n7600 gnd.n429 19.3944
R16437 gnd.n7604 gnd.n429 19.3944
R16438 gnd.n7604 gnd.n425 19.3944
R16439 gnd.n7610 gnd.n425 19.3944
R16440 gnd.n7610 gnd.n423 19.3944
R16441 gnd.n7614 gnd.n423 19.3944
R16442 gnd.n7614 gnd.n419 19.3944
R16443 gnd.n7620 gnd.n419 19.3944
R16444 gnd.n7620 gnd.n417 19.3944
R16445 gnd.n7624 gnd.n417 19.3944
R16446 gnd.n7624 gnd.n413 19.3944
R16447 gnd.n7630 gnd.n413 19.3944
R16448 gnd.n7630 gnd.n411 19.3944
R16449 gnd.n7634 gnd.n411 19.3944
R16450 gnd.n7634 gnd.n407 19.3944
R16451 gnd.n7640 gnd.n407 19.3944
R16452 gnd.n7640 gnd.n405 19.3944
R16453 gnd.n7644 gnd.n405 19.3944
R16454 gnd.n7644 gnd.n401 19.3944
R16455 gnd.n7650 gnd.n401 19.3944
R16456 gnd.n7650 gnd.n399 19.3944
R16457 gnd.n7654 gnd.n399 19.3944
R16458 gnd.n7654 gnd.n395 19.3944
R16459 gnd.n7660 gnd.n395 19.3944
R16460 gnd.n7660 gnd.n393 19.3944
R16461 gnd.n7664 gnd.n393 19.3944
R16462 gnd.n7664 gnd.n389 19.3944
R16463 gnd.n7670 gnd.n389 19.3944
R16464 gnd.n7670 gnd.n387 19.3944
R16465 gnd.n7674 gnd.n387 19.3944
R16466 gnd.n7674 gnd.n383 19.3944
R16467 gnd.n7680 gnd.n383 19.3944
R16468 gnd.n7680 gnd.n381 19.3944
R16469 gnd.n7684 gnd.n381 19.3944
R16470 gnd.n7684 gnd.n377 19.3944
R16471 gnd.n7690 gnd.n377 19.3944
R16472 gnd.n7690 gnd.n375 19.3944
R16473 gnd.n7694 gnd.n375 19.3944
R16474 gnd.n7694 gnd.n371 19.3944
R16475 gnd.n7701 gnd.n371 19.3944
R16476 gnd.n7701 gnd.n369 19.3944
R16477 gnd.n7706 gnd.n369 19.3944
R16478 gnd.n7009 gnd.n784 19.3944
R16479 gnd.n7009 gnd.n782 19.3944
R16480 gnd.n7013 gnd.n782 19.3944
R16481 gnd.n7013 gnd.n778 19.3944
R16482 gnd.n7019 gnd.n778 19.3944
R16483 gnd.n7019 gnd.n776 19.3944
R16484 gnd.n7023 gnd.n776 19.3944
R16485 gnd.n7023 gnd.n772 19.3944
R16486 gnd.n7029 gnd.n772 19.3944
R16487 gnd.n7029 gnd.n770 19.3944
R16488 gnd.n7033 gnd.n770 19.3944
R16489 gnd.n7033 gnd.n766 19.3944
R16490 gnd.n7039 gnd.n766 19.3944
R16491 gnd.n7039 gnd.n764 19.3944
R16492 gnd.n7043 gnd.n764 19.3944
R16493 gnd.n7043 gnd.n760 19.3944
R16494 gnd.n7049 gnd.n760 19.3944
R16495 gnd.n7049 gnd.n758 19.3944
R16496 gnd.n7053 gnd.n758 19.3944
R16497 gnd.n7053 gnd.n754 19.3944
R16498 gnd.n7059 gnd.n754 19.3944
R16499 gnd.n7059 gnd.n752 19.3944
R16500 gnd.n7063 gnd.n752 19.3944
R16501 gnd.n7063 gnd.n748 19.3944
R16502 gnd.n7069 gnd.n748 19.3944
R16503 gnd.n7069 gnd.n746 19.3944
R16504 gnd.n7073 gnd.n746 19.3944
R16505 gnd.n7073 gnd.n742 19.3944
R16506 gnd.n7079 gnd.n742 19.3944
R16507 gnd.n7079 gnd.n740 19.3944
R16508 gnd.n7083 gnd.n740 19.3944
R16509 gnd.n7083 gnd.n736 19.3944
R16510 gnd.n7089 gnd.n736 19.3944
R16511 gnd.n7089 gnd.n734 19.3944
R16512 gnd.n7093 gnd.n734 19.3944
R16513 gnd.n7093 gnd.n730 19.3944
R16514 gnd.n7099 gnd.n730 19.3944
R16515 gnd.n7099 gnd.n728 19.3944
R16516 gnd.n7103 gnd.n728 19.3944
R16517 gnd.n7103 gnd.n724 19.3944
R16518 gnd.n7109 gnd.n724 19.3944
R16519 gnd.n7109 gnd.n722 19.3944
R16520 gnd.n7113 gnd.n722 19.3944
R16521 gnd.n7113 gnd.n718 19.3944
R16522 gnd.n7119 gnd.n718 19.3944
R16523 gnd.n7119 gnd.n716 19.3944
R16524 gnd.n7123 gnd.n716 19.3944
R16525 gnd.n7123 gnd.n712 19.3944
R16526 gnd.n7129 gnd.n712 19.3944
R16527 gnd.n7129 gnd.n710 19.3944
R16528 gnd.n7133 gnd.n710 19.3944
R16529 gnd.n7133 gnd.n706 19.3944
R16530 gnd.n7139 gnd.n706 19.3944
R16531 gnd.n7139 gnd.n704 19.3944
R16532 gnd.n7143 gnd.n704 19.3944
R16533 gnd.n7143 gnd.n700 19.3944
R16534 gnd.n7149 gnd.n700 19.3944
R16535 gnd.n7149 gnd.n698 19.3944
R16536 gnd.n7153 gnd.n698 19.3944
R16537 gnd.n7153 gnd.n694 19.3944
R16538 gnd.n7159 gnd.n694 19.3944
R16539 gnd.n7159 gnd.n692 19.3944
R16540 gnd.n7163 gnd.n692 19.3944
R16541 gnd.n7163 gnd.n688 19.3944
R16542 gnd.n7169 gnd.n688 19.3944
R16543 gnd.n7169 gnd.n686 19.3944
R16544 gnd.n7173 gnd.n686 19.3944
R16545 gnd.n7173 gnd.n682 19.3944
R16546 gnd.n7179 gnd.n682 19.3944
R16547 gnd.n7179 gnd.n680 19.3944
R16548 gnd.n7183 gnd.n680 19.3944
R16549 gnd.n7183 gnd.n676 19.3944
R16550 gnd.n7189 gnd.n676 19.3944
R16551 gnd.n7189 gnd.n674 19.3944
R16552 gnd.n7193 gnd.n674 19.3944
R16553 gnd.n7193 gnd.n670 19.3944
R16554 gnd.n7199 gnd.n670 19.3944
R16555 gnd.n7199 gnd.n668 19.3944
R16556 gnd.n7203 gnd.n668 19.3944
R16557 gnd.n7203 gnd.n664 19.3944
R16558 gnd.n7209 gnd.n664 19.3944
R16559 gnd.n7209 gnd.n662 19.3944
R16560 gnd.n7213 gnd.n662 19.3944
R16561 gnd.n7213 gnd.n658 19.3944
R16562 gnd.n7219 gnd.n658 19.3944
R16563 gnd.n7219 gnd.n656 19.3944
R16564 gnd.n7223 gnd.n656 19.3944
R16565 gnd.n7223 gnd.n652 19.3944
R16566 gnd.n7229 gnd.n652 19.3944
R16567 gnd.n7229 gnd.n650 19.3944
R16568 gnd.n7233 gnd.n650 19.3944
R16569 gnd.n7233 gnd.n646 19.3944
R16570 gnd.n7239 gnd.n646 19.3944
R16571 gnd.n7239 gnd.n644 19.3944
R16572 gnd.n7243 gnd.n644 19.3944
R16573 gnd.n7243 gnd.n640 19.3944
R16574 gnd.n7249 gnd.n640 19.3944
R16575 gnd.n7249 gnd.n638 19.3944
R16576 gnd.n7253 gnd.n638 19.3944
R16577 gnd.n7253 gnd.n634 19.3944
R16578 gnd.n7259 gnd.n634 19.3944
R16579 gnd.n7259 gnd.n632 19.3944
R16580 gnd.n7263 gnd.n632 19.3944
R16581 gnd.n7263 gnd.n628 19.3944
R16582 gnd.n7269 gnd.n628 19.3944
R16583 gnd.n7269 gnd.n626 19.3944
R16584 gnd.n7273 gnd.n626 19.3944
R16585 gnd.n7273 gnd.n622 19.3944
R16586 gnd.n7279 gnd.n622 19.3944
R16587 gnd.n7279 gnd.n620 19.3944
R16588 gnd.n7283 gnd.n620 19.3944
R16589 gnd.n7283 gnd.n616 19.3944
R16590 gnd.n7289 gnd.n616 19.3944
R16591 gnd.n7289 gnd.n614 19.3944
R16592 gnd.n7293 gnd.n614 19.3944
R16593 gnd.n7293 gnd.n610 19.3944
R16594 gnd.n7299 gnd.n610 19.3944
R16595 gnd.n7299 gnd.n608 19.3944
R16596 gnd.n7303 gnd.n608 19.3944
R16597 gnd.n7303 gnd.n604 19.3944
R16598 gnd.n7309 gnd.n604 19.3944
R16599 gnd.n7309 gnd.n602 19.3944
R16600 gnd.n7313 gnd.n602 19.3944
R16601 gnd.n7313 gnd.n598 19.3944
R16602 gnd.n7319 gnd.n598 19.3944
R16603 gnd.n7319 gnd.n596 19.3944
R16604 gnd.n7323 gnd.n596 19.3944
R16605 gnd.n7323 gnd.n592 19.3944
R16606 gnd.n7329 gnd.n592 19.3944
R16607 gnd.n7329 gnd.n590 19.3944
R16608 gnd.n7333 gnd.n590 19.3944
R16609 gnd.n7333 gnd.n586 19.3944
R16610 gnd.n7339 gnd.n586 19.3944
R16611 gnd.n7339 gnd.n584 19.3944
R16612 gnd.n7343 gnd.n584 19.3944
R16613 gnd.n7343 gnd.n580 19.3944
R16614 gnd.n7349 gnd.n580 19.3944
R16615 gnd.n7349 gnd.n578 19.3944
R16616 gnd.n7353 gnd.n578 19.3944
R16617 gnd.n7353 gnd.n574 19.3944
R16618 gnd.n7359 gnd.n574 19.3944
R16619 gnd.n7359 gnd.n572 19.3944
R16620 gnd.n7363 gnd.n572 19.3944
R16621 gnd.n7363 gnd.n568 19.3944
R16622 gnd.n7369 gnd.n568 19.3944
R16623 gnd.n7369 gnd.n566 19.3944
R16624 gnd.n7373 gnd.n566 19.3944
R16625 gnd.n7373 gnd.n562 19.3944
R16626 gnd.n7379 gnd.n562 19.3944
R16627 gnd.n7379 gnd.n560 19.3944
R16628 gnd.n7383 gnd.n560 19.3944
R16629 gnd.n7383 gnd.n556 19.3944
R16630 gnd.n7389 gnd.n556 19.3944
R16631 gnd.n7389 gnd.n554 19.3944
R16632 gnd.n7393 gnd.n554 19.3944
R16633 gnd.n7393 gnd.n550 19.3944
R16634 gnd.n7399 gnd.n550 19.3944
R16635 gnd.n7399 gnd.n548 19.3944
R16636 gnd.n7403 gnd.n548 19.3944
R16637 gnd.n7403 gnd.n544 19.3944
R16638 gnd.n7409 gnd.n544 19.3944
R16639 gnd.n7409 gnd.n542 19.3944
R16640 gnd.n7413 gnd.n542 19.3944
R16641 gnd.n7413 gnd.n538 19.3944
R16642 gnd.n7419 gnd.n538 19.3944
R16643 gnd.n7419 gnd.n536 19.3944
R16644 gnd.n7423 gnd.n536 19.3944
R16645 gnd.n7423 gnd.n532 19.3944
R16646 gnd.n7429 gnd.n532 19.3944
R16647 gnd.n7429 gnd.n530 19.3944
R16648 gnd.n7433 gnd.n530 19.3944
R16649 gnd.n7433 gnd.n526 19.3944
R16650 gnd.n7439 gnd.n526 19.3944
R16651 gnd.n7439 gnd.n524 19.3944
R16652 gnd.n7443 gnd.n524 19.3944
R16653 gnd.n7443 gnd.n520 19.3944
R16654 gnd.n7449 gnd.n520 19.3944
R16655 gnd.n7449 gnd.n518 19.3944
R16656 gnd.n7453 gnd.n518 19.3944
R16657 gnd.n7453 gnd.n514 19.3944
R16658 gnd.n7459 gnd.n514 19.3944
R16659 gnd.n7459 gnd.n512 19.3944
R16660 gnd.n7463 gnd.n512 19.3944
R16661 gnd.n7463 gnd.n508 19.3944
R16662 gnd.n7469 gnd.n508 19.3944
R16663 gnd.n7469 gnd.n506 19.3944
R16664 gnd.n7473 gnd.n506 19.3944
R16665 gnd.n7473 gnd.n502 19.3944
R16666 gnd.n7479 gnd.n502 19.3944
R16667 gnd.n7479 gnd.n500 19.3944
R16668 gnd.n7484 gnd.n500 19.3944
R16669 gnd.n7484 gnd.n496 19.3944
R16670 gnd.n7490 gnd.n496 19.3944
R16671 gnd.n7491 gnd.n7490 19.3944
R16672 gnd.n6131 gnd.n6130 19.3944
R16673 gnd.n6130 gnd.n6129 19.3944
R16674 gnd.n6129 gnd.n6128 19.3944
R16675 gnd.n6128 gnd.n6126 19.3944
R16676 gnd.n6126 gnd.n6123 19.3944
R16677 gnd.n6123 gnd.n6122 19.3944
R16678 gnd.n6122 gnd.n6119 19.3944
R16679 gnd.n6119 gnd.n6118 19.3944
R16680 gnd.n6118 gnd.n6115 19.3944
R16681 gnd.n6115 gnd.n6114 19.3944
R16682 gnd.n6114 gnd.n6111 19.3944
R16683 gnd.n6111 gnd.n6110 19.3944
R16684 gnd.n6110 gnd.n6107 19.3944
R16685 gnd.n6107 gnd.n6106 19.3944
R16686 gnd.n6106 gnd.n6103 19.3944
R16687 gnd.n6103 gnd.n6102 19.3944
R16688 gnd.n6102 gnd.n6099 19.3944
R16689 gnd.n6097 gnd.n6094 19.3944
R16690 gnd.n6094 gnd.n6093 19.3944
R16691 gnd.n6093 gnd.n6090 19.3944
R16692 gnd.n6090 gnd.n6089 19.3944
R16693 gnd.n6089 gnd.n6086 19.3944
R16694 gnd.n6086 gnd.n6085 19.3944
R16695 gnd.n6085 gnd.n6082 19.3944
R16696 gnd.n6080 gnd.n6077 19.3944
R16697 gnd.n6077 gnd.n6076 19.3944
R16698 gnd.n6076 gnd.n6073 19.3944
R16699 gnd.n6073 gnd.n6072 19.3944
R16700 gnd.n6072 gnd.n6069 19.3944
R16701 gnd.n6069 gnd.n6068 19.3944
R16702 gnd.n6068 gnd.n6065 19.3944
R16703 gnd.n6065 gnd.n6064 19.3944
R16704 gnd.n6060 gnd.n6057 19.3944
R16705 gnd.n6057 gnd.n6056 19.3944
R16706 gnd.n6056 gnd.n6053 19.3944
R16707 gnd.n6053 gnd.n6052 19.3944
R16708 gnd.n6052 gnd.n6049 19.3944
R16709 gnd.n6049 gnd.n6048 19.3944
R16710 gnd.n6048 gnd.n6045 19.3944
R16711 gnd.n6045 gnd.n6044 19.3944
R16712 gnd.n6044 gnd.n6041 19.3944
R16713 gnd.n6041 gnd.n6040 19.3944
R16714 gnd.n6040 gnd.n6037 19.3944
R16715 gnd.n6037 gnd.n6036 19.3944
R16716 gnd.n6036 gnd.n6033 19.3944
R16717 gnd.n6033 gnd.n6032 19.3944
R16718 gnd.n6032 gnd.n6029 19.3944
R16719 gnd.n6029 gnd.n6028 19.3944
R16720 gnd.n6028 gnd.n6025 19.3944
R16721 gnd.n6025 gnd.n6024 19.3944
R16722 gnd.n6008 gnd.n3184 19.3944
R16723 gnd.n6008 gnd.n6007 19.3944
R16724 gnd.n6007 gnd.n3193 19.3944
R16725 gnd.n3389 gnd.n3193 19.3944
R16726 gnd.n5703 gnd.n3389 19.3944
R16727 gnd.n5704 gnd.n5703 19.3944
R16728 gnd.n5706 gnd.n5704 19.3944
R16729 gnd.n5706 gnd.n3385 19.3944
R16730 gnd.n5718 gnd.n3385 19.3944
R16731 gnd.n5719 gnd.n5718 19.3944
R16732 gnd.n5721 gnd.n5719 19.3944
R16733 gnd.n5721 gnd.n3380 19.3944
R16734 gnd.n5733 gnd.n3380 19.3944
R16735 gnd.n5734 gnd.n5733 19.3944
R16736 gnd.n5736 gnd.n5734 19.3944
R16737 gnd.n5736 gnd.n3376 19.3944
R16738 gnd.n5748 gnd.n3376 19.3944
R16739 gnd.n5749 gnd.n5748 19.3944
R16740 gnd.n5751 gnd.n5749 19.3944
R16741 gnd.n5751 gnd.n3371 19.3944
R16742 gnd.n5763 gnd.n3371 19.3944
R16743 gnd.n5764 gnd.n5763 19.3944
R16744 gnd.n5766 gnd.n5764 19.3944
R16745 gnd.n5766 gnd.n3366 19.3944
R16746 gnd.n5790 gnd.n3366 19.3944
R16747 gnd.n5791 gnd.n5790 19.3944
R16748 gnd.n5792 gnd.n5791 19.3944
R16749 gnd.n5795 gnd.n5792 19.3944
R16750 gnd.n5795 gnd.n3364 19.3944
R16751 gnd.n5803 gnd.n3364 19.3944
R16752 gnd.n5804 gnd.n5803 19.3944
R16753 gnd.n5805 gnd.n5804 19.3944
R16754 gnd.n5906 gnd.n5805 19.3944
R16755 gnd.n5906 gnd.n5905 19.3944
R16756 gnd.n5905 gnd.n5904 19.3944
R16757 gnd.n5904 gnd.n5809 19.3944
R16758 gnd.n5838 gnd.n5809 19.3944
R16759 gnd.n5839 gnd.n5838 19.3944
R16760 gnd.n5840 gnd.n5839 19.3944
R16761 gnd.n5882 gnd.n5840 19.3944
R16762 gnd.n5882 gnd.n5881 19.3944
R16763 gnd.n5881 gnd.n5880 19.3944
R16764 gnd.n5880 gnd.n5842 19.3944
R16765 gnd.n5870 gnd.n5842 19.3944
R16766 gnd.n5870 gnd.n5869 19.3944
R16767 gnd.n5869 gnd.n5868 19.3944
R16768 gnd.n5868 gnd.n355 19.3944
R16769 gnd.n7823 gnd.n355 19.3944
R16770 gnd.n7824 gnd.n7823 19.3944
R16771 gnd.n7826 gnd.n7824 19.3944
R16772 gnd.n7827 gnd.n7826 19.3944
R16773 gnd.n7830 gnd.n7827 19.3944
R16774 gnd.n7831 gnd.n7830 19.3944
R16775 gnd.n7833 gnd.n7831 19.3944
R16776 gnd.n7834 gnd.n7833 19.3944
R16777 gnd.n7837 gnd.n7834 19.3944
R16778 gnd.n7838 gnd.n7837 19.3944
R16779 gnd.n7840 gnd.n7838 19.3944
R16780 gnd.n7841 gnd.n7840 19.3944
R16781 gnd.n7844 gnd.n7841 19.3944
R16782 gnd.n7845 gnd.n7844 19.3944
R16783 gnd.n7847 gnd.n7845 19.3944
R16784 gnd.n7848 gnd.n7847 19.3944
R16785 gnd.n7851 gnd.n7848 19.3944
R16786 gnd.n6011 gnd.n6010 19.3944
R16787 gnd.n6010 gnd.n3191 19.3944
R16788 gnd.n3215 gnd.n3191 19.3944
R16789 gnd.n5997 gnd.n3215 19.3944
R16790 gnd.n5997 gnd.n5996 19.3944
R16791 gnd.n5996 gnd.n5995 19.3944
R16792 gnd.n5995 gnd.n3220 19.3944
R16793 gnd.n5985 gnd.n3220 19.3944
R16794 gnd.n5985 gnd.n5984 19.3944
R16795 gnd.n5984 gnd.n5983 19.3944
R16796 gnd.n5983 gnd.n3241 19.3944
R16797 gnd.n5973 gnd.n3241 19.3944
R16798 gnd.n5973 gnd.n5972 19.3944
R16799 gnd.n5972 gnd.n5971 19.3944
R16800 gnd.n5971 gnd.n3261 19.3944
R16801 gnd.n5961 gnd.n3261 19.3944
R16802 gnd.n5961 gnd.n5960 19.3944
R16803 gnd.n5960 gnd.n5959 19.3944
R16804 gnd.n5959 gnd.n3282 19.3944
R16805 gnd.n5949 gnd.n3282 19.3944
R16806 gnd.n5949 gnd.n5948 19.3944
R16807 gnd.n5948 gnd.n5947 19.3944
R16808 gnd.n5947 gnd.n3302 19.3944
R16809 gnd.n5937 gnd.n3302 19.3944
R16810 gnd.n5937 gnd.n5936 19.3944
R16811 gnd.n5936 gnd.n5935 19.3944
R16812 gnd.n5935 gnd.n3324 19.3944
R16813 gnd.n5797 gnd.n3324 19.3944
R16814 gnd.n5800 gnd.n5797 19.3944
R16815 gnd.n5800 gnd.n3355 19.3944
R16816 gnd.n5912 gnd.n3355 19.3944
R16817 gnd.n5912 gnd.n5911 19.3944
R16818 gnd.n5911 gnd.n5910 19.3944
R16819 gnd.n5910 gnd.n3359 19.3944
R16820 gnd.n5900 gnd.n3359 19.3944
R16821 gnd.n5900 gnd.n124 19.3944
R16822 gnd.n8057 gnd.n124 19.3944
R16823 gnd.n8057 gnd.n8056 19.3944
R16824 gnd.n8056 gnd.n8055 19.3944
R16825 gnd.n8055 gnd.n128 19.3944
R16826 gnd.n8045 gnd.n128 19.3944
R16827 gnd.n8045 gnd.n8044 19.3944
R16828 gnd.n8044 gnd.n8043 19.3944
R16829 gnd.n8043 gnd.n146 19.3944
R16830 gnd.n8033 gnd.n146 19.3944
R16831 gnd.n8033 gnd.n8032 19.3944
R16832 gnd.n8032 gnd.n8031 19.3944
R16833 gnd.n8031 gnd.n167 19.3944
R16834 gnd.n8021 gnd.n167 19.3944
R16835 gnd.n8021 gnd.n8020 19.3944
R16836 gnd.n8020 gnd.n8019 19.3944
R16837 gnd.n8019 gnd.n186 19.3944
R16838 gnd.n8009 gnd.n186 19.3944
R16839 gnd.n8009 gnd.n8008 19.3944
R16840 gnd.n8008 gnd.n8007 19.3944
R16841 gnd.n8007 gnd.n207 19.3944
R16842 gnd.n7997 gnd.n207 19.3944
R16843 gnd.n7997 gnd.n7996 19.3944
R16844 gnd.n7996 gnd.n7995 19.3944
R16845 gnd.n7995 gnd.n225 19.3944
R16846 gnd.n7985 gnd.n225 19.3944
R16847 gnd.n7985 gnd.n7984 19.3944
R16848 gnd.n7984 gnd.n7983 19.3944
R16849 gnd.n7983 gnd.n245 19.3944
R16850 gnd.n7894 gnd.n331 19.3944
R16851 gnd.n7894 gnd.n7891 19.3944
R16852 gnd.n7891 gnd.n7888 19.3944
R16853 gnd.n7888 gnd.n7887 19.3944
R16854 gnd.n7887 gnd.n7884 19.3944
R16855 gnd.n7884 gnd.n7883 19.3944
R16856 gnd.n7883 gnd.n7880 19.3944
R16857 gnd.n7880 gnd.n7879 19.3944
R16858 gnd.n7879 gnd.n7876 19.3944
R16859 gnd.n7876 gnd.n7875 19.3944
R16860 gnd.n7875 gnd.n7872 19.3944
R16861 gnd.n7872 gnd.n7871 19.3944
R16862 gnd.n7871 gnd.n7868 19.3944
R16863 gnd.n7868 gnd.n7867 19.3944
R16864 gnd.n7867 gnd.n7864 19.3944
R16865 gnd.n7864 gnd.n7863 19.3944
R16866 gnd.n7863 gnd.n7860 19.3944
R16867 gnd.n7860 gnd.n7859 19.3944
R16868 gnd.n7937 gnd.n7934 19.3944
R16869 gnd.n7934 gnd.n7933 19.3944
R16870 gnd.n7933 gnd.n7930 19.3944
R16871 gnd.n7930 gnd.n7929 19.3944
R16872 gnd.n7929 gnd.n7926 19.3944
R16873 gnd.n7926 gnd.n7925 19.3944
R16874 gnd.n7925 gnd.n7922 19.3944
R16875 gnd.n7922 gnd.n7921 19.3944
R16876 gnd.n7921 gnd.n7918 19.3944
R16877 gnd.n7918 gnd.n7917 19.3944
R16878 gnd.n7917 gnd.n7914 19.3944
R16879 gnd.n7914 gnd.n7913 19.3944
R16880 gnd.n7913 gnd.n7910 19.3944
R16881 gnd.n7910 gnd.n7909 19.3944
R16882 gnd.n7909 gnd.n7906 19.3944
R16883 gnd.n7906 gnd.n7905 19.3944
R16884 gnd.n7905 gnd.n7902 19.3944
R16885 gnd.n7902 gnd.n7901 19.3944
R16886 gnd.n7975 gnd.n254 19.3944
R16887 gnd.n7970 gnd.n254 19.3944
R16888 gnd.n7970 gnd.n7969 19.3944
R16889 gnd.n7969 gnd.n7968 19.3944
R16890 gnd.n7968 gnd.n7965 19.3944
R16891 gnd.n7965 gnd.n7964 19.3944
R16892 gnd.n7964 gnd.n7961 19.3944
R16893 gnd.n7961 gnd.n7960 19.3944
R16894 gnd.n7960 gnd.n7957 19.3944
R16895 gnd.n7957 gnd.n7956 19.3944
R16896 gnd.n7956 gnd.n7953 19.3944
R16897 gnd.n7953 gnd.n7952 19.3944
R16898 gnd.n7952 gnd.n7949 19.3944
R16899 gnd.n7949 gnd.n7948 19.3944
R16900 gnd.n7948 gnd.n7945 19.3944
R16901 gnd.n7945 gnd.n7944 19.3944
R16902 gnd.n7944 gnd.n7941 19.3944
R16903 gnd.n7750 gnd.n7748 19.3944
R16904 gnd.n7753 gnd.n7750 19.3944
R16905 gnd.n7756 gnd.n7753 19.3944
R16906 gnd.n7759 gnd.n7756 19.3944
R16907 gnd.n7759 gnd.n7746 19.3944
R16908 gnd.n7763 gnd.n7746 19.3944
R16909 gnd.n7766 gnd.n7763 19.3944
R16910 gnd.n7769 gnd.n7766 19.3944
R16911 gnd.n7769 gnd.n7744 19.3944
R16912 gnd.n7773 gnd.n7744 19.3944
R16913 gnd.n7776 gnd.n7773 19.3944
R16914 gnd.n7779 gnd.n7776 19.3944
R16915 gnd.n7779 gnd.n7742 19.3944
R16916 gnd.n7783 gnd.n7742 19.3944
R16917 gnd.n7786 gnd.n7783 19.3944
R16918 gnd.n7789 gnd.n7786 19.3944
R16919 gnd.n5691 gnd.n3392 19.3944
R16920 gnd.n5692 gnd.n5691 19.3944
R16921 gnd.n5695 gnd.n5692 19.3944
R16922 gnd.n5695 gnd.n3390 19.3944
R16923 gnd.n5699 gnd.n3390 19.3944
R16924 gnd.n5699 gnd.n3388 19.3944
R16925 gnd.n5710 gnd.n3388 19.3944
R16926 gnd.n5710 gnd.n3386 19.3944
R16927 gnd.n5714 gnd.n3386 19.3944
R16928 gnd.n5714 gnd.n3384 19.3944
R16929 gnd.n5725 gnd.n3384 19.3944
R16930 gnd.n5725 gnd.n3382 19.3944
R16931 gnd.n5729 gnd.n3382 19.3944
R16932 gnd.n5729 gnd.n3379 19.3944
R16933 gnd.n5740 gnd.n3379 19.3944
R16934 gnd.n5740 gnd.n3377 19.3944
R16935 gnd.n5744 gnd.n3377 19.3944
R16936 gnd.n5744 gnd.n3375 19.3944
R16937 gnd.n5755 gnd.n3375 19.3944
R16938 gnd.n5755 gnd.n3373 19.3944
R16939 gnd.n5759 gnd.n3373 19.3944
R16940 gnd.n5759 gnd.n3370 19.3944
R16941 gnd.n5770 gnd.n3370 19.3944
R16942 gnd.n5770 gnd.n3367 19.3944
R16943 gnd.n5786 gnd.n3367 19.3944
R16944 gnd.n5786 gnd.n3368 19.3944
R16945 gnd.n5782 gnd.n3368 19.3944
R16946 gnd.n5782 gnd.n5781 19.3944
R16947 gnd.n5781 gnd.n5780 19.3944
R16948 gnd.n5780 gnd.n5777 19.3944
R16949 gnd.n5777 gnd.n5776 19.3944
R16950 gnd.n5776 gnd.n96 19.3944
R16951 gnd.n8070 gnd.n96 19.3944
R16952 gnd.n8070 gnd.n8069 19.3944
R16953 gnd.n8069 gnd.n99 19.3944
R16954 gnd.n5831 gnd.n99 19.3944
R16955 gnd.n5831 gnd.n5827 19.3944
R16956 gnd.n5888 gnd.n5827 19.3944
R16957 gnd.n5888 gnd.n5887 19.3944
R16958 gnd.n5887 gnd.n5886 19.3944
R16959 gnd.n5886 gnd.n5837 19.3944
R16960 gnd.n5876 gnd.n5837 19.3944
R16961 gnd.n5876 gnd.n5875 19.3944
R16962 gnd.n5875 gnd.n5874 19.3944
R16963 gnd.n5874 gnd.n359 19.3944
R16964 gnd.n7718 gnd.n359 19.3944
R16965 gnd.n7718 gnd.n357 19.3944
R16966 gnd.n7819 gnd.n357 19.3944
R16967 gnd.n7819 gnd.n7818 19.3944
R16968 gnd.n7818 gnd.n7817 19.3944
R16969 gnd.n7817 gnd.n7815 19.3944
R16970 gnd.n7815 gnd.n7814 19.3944
R16971 gnd.n7814 gnd.n7812 19.3944
R16972 gnd.n7812 gnd.n7811 19.3944
R16973 gnd.n7811 gnd.n7809 19.3944
R16974 gnd.n7809 gnd.n7808 19.3944
R16975 gnd.n7808 gnd.n7806 19.3944
R16976 gnd.n7806 gnd.n7805 19.3944
R16977 gnd.n7805 gnd.n7803 19.3944
R16978 gnd.n7803 gnd.n7802 19.3944
R16979 gnd.n7802 gnd.n7800 19.3944
R16980 gnd.n7800 gnd.n7799 19.3944
R16981 gnd.n7799 gnd.n7797 19.3944
R16982 gnd.n7797 gnd.n7796 19.3944
R16983 gnd.n3201 gnd.n3200 19.3944
R16984 gnd.n6003 gnd.n3200 19.3944
R16985 gnd.n6003 gnd.n6002 19.3944
R16986 gnd.n6002 gnd.n6001 19.3944
R16987 gnd.n6001 gnd.n3207 19.3944
R16988 gnd.n5991 gnd.n3207 19.3944
R16989 gnd.n5991 gnd.n5990 19.3944
R16990 gnd.n5990 gnd.n5989 19.3944
R16991 gnd.n5989 gnd.n3231 19.3944
R16992 gnd.n5979 gnd.n3231 19.3944
R16993 gnd.n5979 gnd.n5978 19.3944
R16994 gnd.n5978 gnd.n5977 19.3944
R16995 gnd.n5977 gnd.n3252 19.3944
R16996 gnd.n5967 gnd.n3252 19.3944
R16997 gnd.n5967 gnd.n5966 19.3944
R16998 gnd.n5966 gnd.n5965 19.3944
R16999 gnd.n5965 gnd.n3272 19.3944
R17000 gnd.n5955 gnd.n3272 19.3944
R17001 gnd.n5955 gnd.n5954 19.3944
R17002 gnd.n5954 gnd.n5953 19.3944
R17003 gnd.n5953 gnd.n3293 19.3944
R17004 gnd.n5943 gnd.n3293 19.3944
R17005 gnd.n5943 gnd.n5942 19.3944
R17006 gnd.n5942 gnd.n5941 19.3944
R17007 gnd.n5941 gnd.n3314 19.3944
R17008 gnd.n5931 gnd.n3314 19.3944
R17009 gnd.n5931 gnd.n5930 19.3944
R17010 gnd.n3346 gnd.n3345 19.3944
R17011 gnd.n5917 gnd.n5916 19.3944
R17012 gnd.n3349 gnd.n3348 19.3944
R17013 gnd.n8065 gnd.n8064 19.3944
R17014 gnd.n8061 gnd.n108 19.3944
R17015 gnd.n8061 gnd.n115 19.3944
R17016 gnd.n8051 gnd.n115 19.3944
R17017 gnd.n8051 gnd.n8050 19.3944
R17018 gnd.n8050 gnd.n8049 19.3944
R17019 gnd.n8049 gnd.n137 19.3944
R17020 gnd.n8039 gnd.n137 19.3944
R17021 gnd.n8039 gnd.n8038 19.3944
R17022 gnd.n8038 gnd.n8037 19.3944
R17023 gnd.n8037 gnd.n157 19.3944
R17024 gnd.n8027 gnd.n157 19.3944
R17025 gnd.n8027 gnd.n8026 19.3944
R17026 gnd.n8026 gnd.n8025 19.3944
R17027 gnd.n8025 gnd.n177 19.3944
R17028 gnd.n8015 gnd.n177 19.3944
R17029 gnd.n8015 gnd.n8014 19.3944
R17030 gnd.n8014 gnd.n8013 19.3944
R17031 gnd.n8013 gnd.n197 19.3944
R17032 gnd.n8003 gnd.n197 19.3944
R17033 gnd.n8003 gnd.n8002 19.3944
R17034 gnd.n8002 gnd.n8001 19.3944
R17035 gnd.n8001 gnd.n217 19.3944
R17036 gnd.n7991 gnd.n217 19.3944
R17037 gnd.n7991 gnd.n7990 19.3944
R17038 gnd.n7990 gnd.n7989 19.3944
R17039 gnd.n7989 gnd.n236 19.3944
R17040 gnd.n7979 gnd.n236 19.3944
R17041 gnd.n7979 gnd.n7978 19.3944
R17042 gnd.n4228 gnd.n4222 19.3944
R17043 gnd.n4233 gnd.n4222 19.3944
R17044 gnd.n4233 gnd.n4220 19.3944
R17045 gnd.n4237 gnd.n4220 19.3944
R17046 gnd.n4237 gnd.n4067 19.3944
R17047 gnd.n4241 gnd.n4067 19.3944
R17048 gnd.n4241 gnd.n4065 19.3944
R17049 gnd.n4245 gnd.n4065 19.3944
R17050 gnd.n4245 gnd.n4052 19.3944
R17051 gnd.n4285 gnd.n4052 19.3944
R17052 gnd.n4285 gnd.n4050 19.3944
R17053 gnd.n4289 gnd.n4050 19.3944
R17054 gnd.n4290 gnd.n4289 19.3944
R17055 gnd.n4294 gnd.n4293 19.3944
R17056 gnd.n4304 gnd.n4303 19.3944
R17057 gnd.n4301 gnd.n4298 19.3944
R17058 gnd.n4296 gnd.n4015 19.3944
R17059 gnd.n4350 gnd.n4349 19.3944
R17060 gnd.n4373 gnd.n4350 19.3944
R17061 gnd.n4373 gnd.n4372 19.3944
R17062 gnd.n4372 gnd.n4371 19.3944
R17063 gnd.n4371 gnd.n4355 19.3944
R17064 gnd.n4367 gnd.n4355 19.3944
R17065 gnd.n4367 gnd.n4366 19.3944
R17066 gnd.n4366 gnd.n4365 19.3944
R17067 gnd.n4365 gnd.n4363 19.3944
R17068 gnd.n4363 gnd.n3990 19.3944
R17069 gnd.n3990 gnd.n3988 19.3944
R17070 gnd.n4438 gnd.n3988 19.3944
R17071 gnd.n4438 gnd.n3986 19.3944
R17072 gnd.n4442 gnd.n3986 19.3944
R17073 gnd.n4442 gnd.n3984 19.3944
R17074 gnd.n4446 gnd.n3984 19.3944
R17075 gnd.n4446 gnd.n3982 19.3944
R17076 gnd.n4454 gnd.n3982 19.3944
R17077 gnd.n4454 gnd.n4453 19.3944
R17078 gnd.n4453 gnd.n4452 19.3944
R17079 gnd.n4452 gnd.n3966 19.3944
R17080 gnd.n4741 gnd.n3966 19.3944
R17081 gnd.n4741 gnd.n3964 19.3944
R17082 gnd.n4745 gnd.n3964 19.3944
R17083 gnd.n4745 gnd.n3962 19.3944
R17084 gnd.n4749 gnd.n3962 19.3944
R17085 gnd.n4749 gnd.n3960 19.3944
R17086 gnd.n4761 gnd.n3960 19.3944
R17087 gnd.n4761 gnd.n4760 19.3944
R17088 gnd.n4760 gnd.n4759 19.3944
R17089 gnd.n4759 gnd.n4756 19.3944
R17090 gnd.n4756 gnd.n3932 19.3944
R17091 gnd.n4777 gnd.n3932 19.3944
R17092 gnd.n4777 gnd.n3930 19.3944
R17093 gnd.n4781 gnd.n3930 19.3944
R17094 gnd.n4781 gnd.n3916 19.3944
R17095 gnd.n4810 gnd.n3916 19.3944
R17096 gnd.n4810 gnd.n3914 19.3944
R17097 gnd.n4823 gnd.n3914 19.3944
R17098 gnd.n4823 gnd.n4822 19.3944
R17099 gnd.n4822 gnd.n4821 19.3944
R17100 gnd.n4821 gnd.n4818 19.3944
R17101 gnd.n4818 gnd.n2905 19.3944
R17102 gnd.n6316 gnd.n2905 19.3944
R17103 gnd.n6316 gnd.n6315 19.3944
R17104 gnd.n6315 gnd.n6314 19.3944
R17105 gnd.n6314 gnd.n2909 19.3944
R17106 gnd.n5006 gnd.n2909 19.3944
R17107 gnd.n5010 gnd.n5006 19.3944
R17108 gnd.n5010 gnd.n3805 19.3944
R17109 gnd.n5035 gnd.n3805 19.3944
R17110 gnd.n5035 gnd.n3803 19.3944
R17111 gnd.n5050 gnd.n3803 19.3944
R17112 gnd.n5050 gnd.n5049 19.3944
R17113 gnd.n5049 gnd.n5048 19.3944
R17114 gnd.n5048 gnd.n5041 19.3944
R17115 gnd.n5044 gnd.n5041 19.3944
R17116 gnd.n5044 gnd.n3767 19.3944
R17117 gnd.n5093 gnd.n3767 19.3944
R17118 gnd.n5093 gnd.n3765 19.3944
R17119 gnd.n5097 gnd.n3765 19.3944
R17120 gnd.n5097 gnd.n3749 19.3944
R17121 gnd.n5119 gnd.n3749 19.3944
R17122 gnd.n5119 gnd.n3747 19.3944
R17123 gnd.n5125 gnd.n3747 19.3944
R17124 gnd.n5125 gnd.n5124 19.3944
R17125 gnd.n5124 gnd.n3725 19.3944
R17126 gnd.n5158 gnd.n3725 19.3944
R17127 gnd.n5158 gnd.n3723 19.3944
R17128 gnd.n5173 gnd.n3723 19.3944
R17129 gnd.n5173 gnd.n5172 19.3944
R17130 gnd.n5172 gnd.n5171 19.3944
R17131 gnd.n5171 gnd.n5164 19.3944
R17132 gnd.n5167 gnd.n5164 19.3944
R17133 gnd.n5167 gnd.n3686 19.3944
R17134 gnd.n5216 gnd.n3686 19.3944
R17135 gnd.n5216 gnd.n3684 19.3944
R17136 gnd.n5220 gnd.n3684 19.3944
R17137 gnd.n5220 gnd.n3667 19.3944
R17138 gnd.n5241 gnd.n3667 19.3944
R17139 gnd.n5241 gnd.n3665 19.3944
R17140 gnd.n5247 gnd.n3665 19.3944
R17141 gnd.n5247 gnd.n5246 19.3944
R17142 gnd.n5246 gnd.n3642 19.3944
R17143 gnd.n5279 gnd.n3642 19.3944
R17144 gnd.n5279 gnd.n3640 19.3944
R17145 gnd.n5291 gnd.n3640 19.3944
R17146 gnd.n5291 gnd.n5290 19.3944
R17147 gnd.n5290 gnd.n5289 19.3944
R17148 gnd.n5289 gnd.n5286 19.3944
R17149 gnd.n5286 gnd.n3608 19.3944
R17150 gnd.n5325 gnd.n3608 19.3944
R17151 gnd.n5325 gnd.n3606 19.3944
R17152 gnd.n5331 gnd.n3606 19.3944
R17153 gnd.n5331 gnd.n5330 19.3944
R17154 gnd.n5330 gnd.n3580 19.3944
R17155 gnd.n5360 gnd.n3580 19.3944
R17156 gnd.n5360 gnd.n3578 19.3944
R17157 gnd.n5364 gnd.n3578 19.3944
R17158 gnd.n5364 gnd.n3551 19.3944
R17159 gnd.n5397 gnd.n3551 19.3944
R17160 gnd.n5397 gnd.n3549 19.3944
R17161 gnd.n5403 gnd.n3549 19.3944
R17162 gnd.n5403 gnd.n5402 19.3944
R17163 gnd.n5402 gnd.n3451 19.3944
R17164 gnd.n5547 gnd.n3451 19.3944
R17165 gnd.n5547 gnd.n3449 19.3944
R17166 gnd.n5551 gnd.n3449 19.3944
R17167 gnd.n5551 gnd.n3438 19.3944
R17168 gnd.n5563 gnd.n3438 19.3944
R17169 gnd.n5563 gnd.n3436 19.3944
R17170 gnd.n5570 gnd.n3436 19.3944
R17171 gnd.n5570 gnd.n5569 19.3944
R17172 gnd.n5569 gnd.n3425 19.3944
R17173 gnd.n5583 gnd.n3425 19.3944
R17174 gnd.n5584 gnd.n5583 19.3944
R17175 gnd.n5584 gnd.n3423 19.3944
R17176 gnd.n5680 gnd.n3423 19.3944
R17177 gnd.n5680 gnd.n5679 19.3944
R17178 gnd.n5679 gnd.n5678 19.3944
R17179 gnd.n5678 gnd.n5590 19.3944
R17180 gnd.n5674 gnd.n5590 19.3944
R17181 gnd.n5674 gnd.n5673 19.3944
R17182 gnd.n5673 gnd.n5672 19.3944
R17183 gnd.n5672 gnd.n5596 19.3944
R17184 gnd.n5666 gnd.n5596 19.3944
R17185 gnd.n5666 gnd.n5665 19.3944
R17186 gnd.n5665 gnd.n5664 19.3944
R17187 gnd.n5664 gnd.n5602 19.3944
R17188 gnd.n5660 gnd.n5602 19.3944
R17189 gnd.n5660 gnd.n5659 19.3944
R17190 gnd.n5659 gnd.n5658 19.3944
R17191 gnd.n5658 gnd.n5608 19.3944
R17192 gnd.n5654 gnd.n5608 19.3944
R17193 gnd.n5654 gnd.n5653 19.3944
R17194 gnd.n5653 gnd.n5652 19.3944
R17195 gnd.n5652 gnd.n5614 19.3944
R17196 gnd.n5648 gnd.n5614 19.3944
R17197 gnd.n5648 gnd.n5647 19.3944
R17198 gnd.n5647 gnd.n5646 19.3944
R17199 gnd.n5646 gnd.n5620 19.3944
R17200 gnd.n5642 gnd.n5620 19.3944
R17201 gnd.n5642 gnd.n5641 19.3944
R17202 gnd.n5641 gnd.n5640 19.3944
R17203 gnd.n5640 gnd.n5626 19.3944
R17204 gnd.n5636 gnd.n5626 19.3944
R17205 gnd.n5636 gnd.n5635 19.3944
R17206 gnd.n5635 gnd.n5634 19.3944
R17207 gnd.n5634 gnd.n3336 19.3944
R17208 gnd.n5925 gnd.n3336 19.3944
R17209 gnd.n5923 gnd.n5922 19.3944
R17210 gnd.n5816 gnd.n5814 19.3944
R17211 gnd.n5820 gnd.n5813 19.3944
R17212 gnd.n5897 gnd.n5822 19.3944
R17213 gnd.n5895 gnd.n5894 19.3944
R17214 gnd.n5894 gnd.n5824 19.3944
R17215 gnd.n5847 gnd.n5824 19.3944
R17216 gnd.n5847 gnd.n5845 19.3944
R17217 gnd.n5860 gnd.n5845 19.3944
R17218 gnd.n5860 gnd.n5859 19.3944
R17219 gnd.n5859 gnd.n5858 19.3944
R17220 gnd.n5858 gnd.n5855 19.3944
R17221 gnd.n5855 gnd.n363 19.3944
R17222 gnd.n7713 gnd.n363 19.3944
R17223 gnd.n7713 gnd.n7712 19.3944
R17224 gnd.n7712 gnd.n7711 19.3944
R17225 gnd.n7711 gnd.n367 19.3944
R17226 gnd.n6742 gnd.n6741 19.3944
R17227 gnd.n6741 gnd.n6740 19.3944
R17228 gnd.n6740 gnd.n6739 19.3944
R17229 gnd.n6739 gnd.n6737 19.3944
R17230 gnd.n6737 gnd.n6734 19.3944
R17231 gnd.n6734 gnd.n6733 19.3944
R17232 gnd.n6733 gnd.n6730 19.3944
R17233 gnd.n6730 gnd.n6729 19.3944
R17234 gnd.n6729 gnd.n6726 19.3944
R17235 gnd.n6726 gnd.n6725 19.3944
R17236 gnd.n6725 gnd.n6722 19.3944
R17237 gnd.n6722 gnd.n6721 19.3944
R17238 gnd.n6721 gnd.n6718 19.3944
R17239 gnd.n6718 gnd.n6717 19.3944
R17240 gnd.n6717 gnd.n6714 19.3944
R17241 gnd.n6714 gnd.n6713 19.3944
R17242 gnd.n6713 gnd.n6710 19.3944
R17243 gnd.n6708 gnd.n6705 19.3944
R17244 gnd.n6705 gnd.n6704 19.3944
R17245 gnd.n6704 gnd.n6701 19.3944
R17246 gnd.n6701 gnd.n6700 19.3944
R17247 gnd.n6700 gnd.n6697 19.3944
R17248 gnd.n6697 gnd.n6696 19.3944
R17249 gnd.n6696 gnd.n6693 19.3944
R17250 gnd.n6693 gnd.n6692 19.3944
R17251 gnd.n6692 gnd.n6689 19.3944
R17252 gnd.n6689 gnd.n6688 19.3944
R17253 gnd.n6688 gnd.n6685 19.3944
R17254 gnd.n6685 gnd.n6684 19.3944
R17255 gnd.n6684 gnd.n6681 19.3944
R17256 gnd.n6681 gnd.n6680 19.3944
R17257 gnd.n6680 gnd.n6677 19.3944
R17258 gnd.n6677 gnd.n6676 19.3944
R17259 gnd.n6676 gnd.n6673 19.3944
R17260 gnd.n6673 gnd.n6672 19.3944
R17261 gnd.n6668 gnd.n6665 19.3944
R17262 gnd.n6665 gnd.n6664 19.3944
R17263 gnd.n6664 gnd.n6661 19.3944
R17264 gnd.n6661 gnd.n6660 19.3944
R17265 gnd.n6660 gnd.n6657 19.3944
R17266 gnd.n6657 gnd.n6656 19.3944
R17267 gnd.n6656 gnd.n6653 19.3944
R17268 gnd.n6653 gnd.n6652 19.3944
R17269 gnd.n6652 gnd.n6649 19.3944
R17270 gnd.n6649 gnd.n6648 19.3944
R17271 gnd.n6648 gnd.n6645 19.3944
R17272 gnd.n6645 gnd.n6644 19.3944
R17273 gnd.n6644 gnd.n6641 19.3944
R17274 gnd.n6641 gnd.n6640 19.3944
R17275 gnd.n6640 gnd.n6637 19.3944
R17276 gnd.n6637 gnd.n6636 19.3944
R17277 gnd.n6636 gnd.n6633 19.3944
R17278 gnd.n6633 gnd.n6632 19.3944
R17279 gnd.n4122 gnd.n4121 19.3944
R17280 gnd.n4125 gnd.n4122 19.3944
R17281 gnd.n4125 gnd.n4117 19.3944
R17282 gnd.n4131 gnd.n4117 19.3944
R17283 gnd.n4132 gnd.n4131 19.3944
R17284 gnd.n4135 gnd.n4132 19.3944
R17285 gnd.n4135 gnd.n4115 19.3944
R17286 gnd.n4141 gnd.n4115 19.3944
R17287 gnd.n4142 gnd.n4141 19.3944
R17288 gnd.n4145 gnd.n4142 19.3944
R17289 gnd.n4145 gnd.n4113 19.3944
R17290 gnd.n4151 gnd.n4113 19.3944
R17291 gnd.n4152 gnd.n4151 19.3944
R17292 gnd.n4155 gnd.n4152 19.3944
R17293 gnd.n4155 gnd.n4109 19.3944
R17294 gnd.n4159 gnd.n4109 19.3944
R17295 gnd.n4166 gnd.n4165 19.3944
R17296 gnd.n4168 gnd.n4166 19.3944
R17297 gnd.n4168 gnd.n4103 19.3944
R17298 gnd.n4173 gnd.n4103 19.3944
R17299 gnd.n4174 gnd.n4173 19.3944
R17300 gnd.n4176 gnd.n4174 19.3944
R17301 gnd.n4176 gnd.n4101 19.3944
R17302 gnd.n4181 gnd.n4101 19.3944
R17303 gnd.n4182 gnd.n4181 19.3944
R17304 gnd.n4184 gnd.n4182 19.3944
R17305 gnd.n4184 gnd.n4099 19.3944
R17306 gnd.n4189 gnd.n4099 19.3944
R17307 gnd.n4190 gnd.n4189 19.3944
R17308 gnd.n4192 gnd.n4190 19.3944
R17309 gnd.n4192 gnd.n4097 19.3944
R17310 gnd.n4197 gnd.n4097 19.3944
R17311 gnd.n4197 gnd.n4069 19.3944
R17312 gnd.n4215 gnd.n4069 19.3944
R17313 gnd.n4215 gnd.n4214 19.3944
R17314 gnd.n4214 gnd.n4213 19.3944
R17315 gnd.n4213 gnd.n4062 19.3944
R17316 gnd.n4250 gnd.n4062 19.3944
R17317 gnd.n4250 gnd.n4060 19.3944
R17318 gnd.n4255 gnd.n4060 19.3944
R17319 gnd.n4255 gnd.n4055 19.3944
R17320 gnd.n4279 gnd.n4055 19.3944
R17321 gnd.n4279 gnd.n4278 19.3944
R17322 gnd.n4278 gnd.n4277 19.3944
R17323 gnd.n4277 gnd.n4044 19.3944
R17324 gnd.n4309 gnd.n4044 19.3944
R17325 gnd.n4309 gnd.n4042 19.3944
R17326 gnd.n4313 gnd.n4042 19.3944
R17327 gnd.n4313 gnd.n4021 19.3944
R17328 gnd.n4339 gnd.n4021 19.3944
R17329 gnd.n4339 gnd.n4019 19.3944
R17330 gnd.n4343 gnd.n4019 19.3944
R17331 gnd.n4343 gnd.n4009 19.3944
R17332 gnd.n4378 gnd.n4009 19.3944
R17333 gnd.n4378 gnd.n4007 19.3944
R17334 gnd.n4382 gnd.n4007 19.3944
R17335 gnd.n4382 gnd.n4003 19.3944
R17336 gnd.n4392 gnd.n4003 19.3944
R17337 gnd.n4392 gnd.n4001 19.3944
R17338 gnd.n4396 gnd.n4001 19.3944
R17339 gnd.n4396 gnd.n3992 19.3944
R17340 gnd.n4431 gnd.n3992 19.3944
R17341 gnd.n4431 gnd.n3993 19.3944
R17342 gnd.n4427 gnd.n3993 19.3944
R17343 gnd.n4427 gnd.n4426 19.3944
R17344 gnd.n4426 gnd.n4425 19.3944
R17345 gnd.n4425 gnd.n3998 19.3944
R17346 gnd.n4421 gnd.n3998 19.3944
R17347 gnd.n4421 gnd.n3978 19.3944
R17348 gnd.n4459 gnd.n3978 19.3944
R17349 gnd.n4459 gnd.n3976 19.3944
R17350 gnd.n4463 gnd.n3976 19.3944
R17351 gnd.n4463 gnd.n3969 19.3944
R17352 gnd.n4735 gnd.n3969 19.3944
R17353 gnd.n4735 gnd.n3970 19.3944
R17354 gnd.n4731 gnd.n3970 19.3944
R17355 gnd.n4731 gnd.n4730 19.3944
R17356 gnd.n4730 gnd.n4729 19.3944
R17357 gnd.n4729 gnd.n4726 19.3944
R17358 gnd.n4726 gnd.n3956 19.3944
R17359 gnd.n6624 gnd.n2465 19.3944
R17360 gnd.n4074 gnd.n2465 19.3944
R17361 gnd.n4075 gnd.n4074 19.3944
R17362 gnd.n4077 gnd.n4075 19.3944
R17363 gnd.n4078 gnd.n4077 19.3944
R17364 gnd.n4081 gnd.n4078 19.3944
R17365 gnd.n4082 gnd.n4081 19.3944
R17366 gnd.n4084 gnd.n4082 19.3944
R17367 gnd.n4085 gnd.n4084 19.3944
R17368 gnd.n4088 gnd.n4085 19.3944
R17369 gnd.n4089 gnd.n4088 19.3944
R17370 gnd.n4091 gnd.n4089 19.3944
R17371 gnd.n4092 gnd.n4091 19.3944
R17372 gnd.n4095 gnd.n4092 19.3944
R17373 gnd.n4096 gnd.n4095 19.3944
R17374 gnd.n4201 gnd.n4096 19.3944
R17375 gnd.n4202 gnd.n4201 19.3944
R17376 gnd.n4204 gnd.n4202 19.3944
R17377 gnd.n4205 gnd.n4204 19.3944
R17378 gnd.n4209 gnd.n4205 19.3944
R17379 gnd.n4209 gnd.n4208 19.3944
R17380 gnd.n4208 gnd.n4207 19.3944
R17381 gnd.n4207 gnd.n4059 19.3944
R17382 gnd.n4259 gnd.n4059 19.3944
R17383 gnd.n4260 gnd.n4259 19.3944
R17384 gnd.n4262 gnd.n4260 19.3944
R17385 gnd.n4263 gnd.n4262 19.3944
R17386 gnd.n4273 gnd.n4263 19.3944
R17387 gnd.n4273 gnd.n4272 19.3944
R17388 gnd.n4272 gnd.n4271 19.3944
R17389 gnd.n4271 gnd.n4037 19.3944
R17390 gnd.n4317 gnd.n4037 19.3944
R17391 gnd.n4318 gnd.n4317 19.3944
R17392 gnd.n4319 gnd.n4318 19.3944
R17393 gnd.n4324 gnd.n4319 19.3944
R17394 gnd.n4324 gnd.n4322 19.3944
R17395 gnd.n4322 gnd.n4321 19.3944
R17396 gnd.n4321 gnd.n4320 19.3944
R17397 gnd.n4320 gnd.n4005 19.3944
R17398 gnd.n4386 gnd.n4005 19.3944
R17399 gnd.n4387 gnd.n4386 19.3944
R17400 gnd.n4388 gnd.n4387 19.3944
R17401 gnd.n4388 gnd.n3999 19.3944
R17402 gnd.n4400 gnd.n3999 19.3944
R17403 gnd.n4401 gnd.n4400 19.3944
R17404 gnd.n4402 gnd.n4401 19.3944
R17405 gnd.n4403 gnd.n4402 19.3944
R17406 gnd.n4407 gnd.n4403 19.3944
R17407 gnd.n4408 gnd.n4407 19.3944
R17408 gnd.n4412 gnd.n4408 19.3944
R17409 gnd.n4413 gnd.n4412 19.3944
R17410 gnd.n4417 gnd.n4413 19.3944
R17411 gnd.n4417 gnd.n4416 19.3944
R17412 gnd.n4416 gnd.n4415 19.3944
R17413 gnd.n4415 gnd.n3974 19.3944
R17414 gnd.n4467 gnd.n3974 19.3944
R17415 gnd.n4468 gnd.n4467 19.3944
R17416 gnd.n4469 gnd.n4468 19.3944
R17417 gnd.n4470 gnd.n4469 19.3944
R17418 gnd.n4474 gnd.n4470 19.3944
R17419 gnd.n4475 gnd.n4474 19.3944
R17420 gnd.n4722 gnd.n4475 19.3944
R17421 gnd.n4722 gnd.n4721 19.3944
R17422 gnd.n4721 gnd.n4720 19.3944
R17423 gnd.n2484 gnd.n2463 19.3944
R17424 gnd.n2485 gnd.n2484 19.3944
R17425 gnd.n6613 gnd.n2485 19.3944
R17426 gnd.n6613 gnd.n6612 19.3944
R17427 gnd.n6612 gnd.n6611 19.3944
R17428 gnd.n6611 gnd.n2489 19.3944
R17429 gnd.n6601 gnd.n2489 19.3944
R17430 gnd.n6601 gnd.n6600 19.3944
R17431 gnd.n6600 gnd.n6599 19.3944
R17432 gnd.n6599 gnd.n2508 19.3944
R17433 gnd.n6589 gnd.n2508 19.3944
R17434 gnd.n6589 gnd.n6588 19.3944
R17435 gnd.n6588 gnd.n6587 19.3944
R17436 gnd.n6587 gnd.n2527 19.3944
R17437 gnd.n6577 gnd.n2527 19.3944
R17438 gnd.n6577 gnd.n6576 19.3944
R17439 gnd.n6576 gnd.n6575 19.3944
R17440 gnd.n6575 gnd.n2547 19.3944
R17441 gnd.n6565 gnd.n2547 19.3944
R17442 gnd.n6565 gnd.n6564 19.3944
R17443 gnd.n6564 gnd.n6563 19.3944
R17444 gnd.n6563 gnd.n2567 19.3944
R17445 gnd.n6553 gnd.n2567 19.3944
R17446 gnd.n6553 gnd.n6552 19.3944
R17447 gnd.n6552 gnd.n6551 19.3944
R17448 gnd.n6551 gnd.n2587 19.3944
R17449 gnd.n6541 gnd.n2587 19.3944
R17450 gnd.n6541 gnd.n6540 19.3944
R17451 gnd.n6540 gnd.n6539 19.3944
R17452 gnd.n6539 gnd.n2606 19.3944
R17453 gnd.n4268 gnd.n2606 19.3944
R17454 gnd.n4268 gnd.n4033 19.3944
R17455 gnd.n4329 gnd.n4033 19.3944
R17456 gnd.n4329 gnd.n4328 19.3944
R17457 gnd.n4328 gnd.n4327 19.3944
R17458 gnd.n4327 gnd.n2630 19.3944
R17459 gnd.n6528 gnd.n2630 19.3944
R17460 gnd.n6528 gnd.n6527 19.3944
R17461 gnd.n6527 gnd.n6526 19.3944
R17462 gnd.n6526 gnd.n2634 19.3944
R17463 gnd.n6516 gnd.n2634 19.3944
R17464 gnd.n6516 gnd.n6515 19.3944
R17465 gnd.n6515 gnd.n6514 19.3944
R17466 gnd.n6514 gnd.n2652 19.3944
R17467 gnd.n6504 gnd.n2652 19.3944
R17468 gnd.n6504 gnd.n6503 19.3944
R17469 gnd.n6503 gnd.n6502 19.3944
R17470 gnd.n6502 gnd.n2673 19.3944
R17471 gnd.n6492 gnd.n2673 19.3944
R17472 gnd.n6492 gnd.n6491 19.3944
R17473 gnd.n6491 gnd.n6490 19.3944
R17474 gnd.n6490 gnd.n2692 19.3944
R17475 gnd.n6480 gnd.n2692 19.3944
R17476 gnd.n6480 gnd.n6479 19.3944
R17477 gnd.n6479 gnd.n6478 19.3944
R17478 gnd.n6478 gnd.n2713 19.3944
R17479 gnd.n6468 gnd.n2713 19.3944
R17480 gnd.n6468 gnd.n6467 19.3944
R17481 gnd.n6467 gnd.n6466 19.3944
R17482 gnd.n6466 gnd.n2732 19.3944
R17483 gnd.n6456 gnd.n2732 19.3944
R17484 gnd.n6456 gnd.n6455 19.3944
R17485 gnd.n6455 gnd.n6454 19.3944
R17486 gnd.n6454 gnd.n2753 19.3944
R17487 gnd.n6446 gnd.n2763 19.3944
R17488 gnd.n6441 gnd.n2763 19.3944
R17489 gnd.n6441 gnd.n6440 19.3944
R17490 gnd.n6440 gnd.n6439 19.3944
R17491 gnd.n6439 gnd.n6436 19.3944
R17492 gnd.n6436 gnd.n6435 19.3944
R17493 gnd.n6435 gnd.n6432 19.3944
R17494 gnd.n6432 gnd.n6431 19.3944
R17495 gnd.n6431 gnd.n6428 19.3944
R17496 gnd.n6428 gnd.n6427 19.3944
R17497 gnd.n6427 gnd.n6424 19.3944
R17498 gnd.n6424 gnd.n6423 19.3944
R17499 gnd.n6423 gnd.n6420 19.3944
R17500 gnd.n6420 gnd.n6419 19.3944
R17501 gnd.n6419 gnd.n6416 19.3944
R17502 gnd.n6416 gnd.n6415 19.3944
R17503 gnd.n6415 gnd.n6412 19.3944
R17504 gnd.n4668 gnd.n4634 19.3944
R17505 gnd.n4672 gnd.n4634 19.3944
R17506 gnd.n4675 gnd.n4672 19.3944
R17507 gnd.n4678 gnd.n4675 19.3944
R17508 gnd.n4678 gnd.n4632 19.3944
R17509 gnd.n4682 gnd.n4632 19.3944
R17510 gnd.n4685 gnd.n4682 19.3944
R17511 gnd.n4688 gnd.n4685 19.3944
R17512 gnd.n4688 gnd.n4630 19.3944
R17513 gnd.n4692 gnd.n4630 19.3944
R17514 gnd.n4695 gnd.n4692 19.3944
R17515 gnd.n4698 gnd.n4695 19.3944
R17516 gnd.n4698 gnd.n4628 19.3944
R17517 gnd.n4702 gnd.n4628 19.3944
R17518 gnd.n4705 gnd.n4702 19.3944
R17519 gnd.n4708 gnd.n4705 19.3944
R17520 gnd.n4708 gnd.n4626 19.3944
R17521 gnd.n4713 gnd.n4626 19.3944
R17522 gnd.n4646 gnd.n2832 19.3944
R17523 gnd.n4649 gnd.n4646 19.3944
R17524 gnd.n4649 gnd.n4641 19.3944
R17525 gnd.n4653 gnd.n4641 19.3944
R17526 gnd.n4656 gnd.n4653 19.3944
R17527 gnd.n4659 gnd.n4656 19.3944
R17528 gnd.n4659 gnd.n4639 19.3944
R17529 gnd.n4664 gnd.n4639 19.3944
R17530 gnd.n6410 gnd.n6407 19.3944
R17531 gnd.n6407 gnd.n6406 19.3944
R17532 gnd.n6406 gnd.n6403 19.3944
R17533 gnd.n6403 gnd.n6402 19.3944
R17534 gnd.n6402 gnd.n6399 19.3944
R17535 gnd.n6399 gnd.n6398 19.3944
R17536 gnd.n6398 gnd.n6395 19.3944
R17537 gnd.n6619 gnd.n2471 19.3944
R17538 gnd.n6619 gnd.n6618 19.3944
R17539 gnd.n6618 gnd.n6617 19.3944
R17540 gnd.n6617 gnd.n2476 19.3944
R17541 gnd.n6607 gnd.n2476 19.3944
R17542 gnd.n6607 gnd.n6606 19.3944
R17543 gnd.n6606 gnd.n6605 19.3944
R17544 gnd.n6605 gnd.n2499 19.3944
R17545 gnd.n6595 gnd.n2499 19.3944
R17546 gnd.n6595 gnd.n6594 19.3944
R17547 gnd.n6594 gnd.n6593 19.3944
R17548 gnd.n6593 gnd.n2517 19.3944
R17549 gnd.n6583 gnd.n2517 19.3944
R17550 gnd.n6583 gnd.n6582 19.3944
R17551 gnd.n6582 gnd.n6581 19.3944
R17552 gnd.n6581 gnd.n2538 19.3944
R17553 gnd.n6571 gnd.n2538 19.3944
R17554 gnd.n6571 gnd.n6570 19.3944
R17555 gnd.n6570 gnd.n6569 19.3944
R17556 gnd.n6569 gnd.n2557 19.3944
R17557 gnd.n6559 gnd.n2557 19.3944
R17558 gnd.n6559 gnd.n6558 19.3944
R17559 gnd.n6558 gnd.n6557 19.3944
R17560 gnd.n6557 gnd.n2578 19.3944
R17561 gnd.n6547 gnd.n2578 19.3944
R17562 gnd.n6547 gnd.n6546 19.3944
R17563 gnd.n6546 gnd.n6545 19.3944
R17564 gnd.n6535 gnd.n2613 19.3944
R17565 gnd.n4264 gnd.n2614 19.3944
R17566 gnd.n4029 gnd.n4028 19.3944
R17567 gnd.n4335 gnd.n4334 19.3944
R17568 gnd.n6532 gnd.n2620 19.3944
R17569 gnd.n6532 gnd.n2621 19.3944
R17570 gnd.n6522 gnd.n2621 19.3944
R17571 gnd.n6522 gnd.n6521 19.3944
R17572 gnd.n6521 gnd.n6520 19.3944
R17573 gnd.n6520 gnd.n2643 19.3944
R17574 gnd.n6510 gnd.n2643 19.3944
R17575 gnd.n6510 gnd.n6509 19.3944
R17576 gnd.n6509 gnd.n6508 19.3944
R17577 gnd.n6508 gnd.n2663 19.3944
R17578 gnd.n6498 gnd.n2663 19.3944
R17579 gnd.n6498 gnd.n6497 19.3944
R17580 gnd.n6497 gnd.n6496 19.3944
R17581 gnd.n6496 gnd.n2683 19.3944
R17582 gnd.n6486 gnd.n2683 19.3944
R17583 gnd.n6486 gnd.n6485 19.3944
R17584 gnd.n6485 gnd.n6484 19.3944
R17585 gnd.n6484 gnd.n2703 19.3944
R17586 gnd.n6474 gnd.n2703 19.3944
R17587 gnd.n6474 gnd.n6473 19.3944
R17588 gnd.n6473 gnd.n6472 19.3944
R17589 gnd.n6472 gnd.n2723 19.3944
R17590 gnd.n6462 gnd.n2723 19.3944
R17591 gnd.n6462 gnd.n6461 19.3944
R17592 gnd.n6461 gnd.n6460 19.3944
R17593 gnd.n6460 gnd.n2743 19.3944
R17594 gnd.n6450 gnd.n2743 19.3944
R17595 gnd.n6450 gnd.n6449 19.3944
R17596 gnd.n7003 gnd.n7002 19.3944
R17597 gnd.n7002 gnd.n7001 19.3944
R17598 gnd.n7001 gnd.n791 19.3944
R17599 gnd.n6995 gnd.n791 19.3944
R17600 gnd.n6995 gnd.n6994 19.3944
R17601 gnd.n6994 gnd.n6993 19.3944
R17602 gnd.n6993 gnd.n799 19.3944
R17603 gnd.n6987 gnd.n799 19.3944
R17604 gnd.n6987 gnd.n6986 19.3944
R17605 gnd.n6986 gnd.n6985 19.3944
R17606 gnd.n6985 gnd.n807 19.3944
R17607 gnd.n6979 gnd.n807 19.3944
R17608 gnd.n6979 gnd.n6978 19.3944
R17609 gnd.n6978 gnd.n6977 19.3944
R17610 gnd.n6977 gnd.n815 19.3944
R17611 gnd.n6971 gnd.n815 19.3944
R17612 gnd.n6971 gnd.n6970 19.3944
R17613 gnd.n6970 gnd.n6969 19.3944
R17614 gnd.n6969 gnd.n823 19.3944
R17615 gnd.n6963 gnd.n823 19.3944
R17616 gnd.n6963 gnd.n6962 19.3944
R17617 gnd.n6962 gnd.n6961 19.3944
R17618 gnd.n6961 gnd.n831 19.3944
R17619 gnd.n6955 gnd.n831 19.3944
R17620 gnd.n6955 gnd.n6954 19.3944
R17621 gnd.n6954 gnd.n6953 19.3944
R17622 gnd.n6953 gnd.n839 19.3944
R17623 gnd.n6947 gnd.n839 19.3944
R17624 gnd.n6947 gnd.n6946 19.3944
R17625 gnd.n6946 gnd.n6945 19.3944
R17626 gnd.n6945 gnd.n847 19.3944
R17627 gnd.n6939 gnd.n847 19.3944
R17628 gnd.n6939 gnd.n6938 19.3944
R17629 gnd.n6938 gnd.n6937 19.3944
R17630 gnd.n6937 gnd.n855 19.3944
R17631 gnd.n6931 gnd.n855 19.3944
R17632 gnd.n6931 gnd.n6930 19.3944
R17633 gnd.n6930 gnd.n6929 19.3944
R17634 gnd.n6929 gnd.n863 19.3944
R17635 gnd.n6923 gnd.n863 19.3944
R17636 gnd.n6923 gnd.n6922 19.3944
R17637 gnd.n6922 gnd.n6921 19.3944
R17638 gnd.n6921 gnd.n871 19.3944
R17639 gnd.n6915 gnd.n871 19.3944
R17640 gnd.n6915 gnd.n6914 19.3944
R17641 gnd.n6914 gnd.n6913 19.3944
R17642 gnd.n6913 gnd.n879 19.3944
R17643 gnd.n6907 gnd.n879 19.3944
R17644 gnd.n6907 gnd.n6906 19.3944
R17645 gnd.n6906 gnd.n6905 19.3944
R17646 gnd.n6905 gnd.n887 19.3944
R17647 gnd.n6899 gnd.n887 19.3944
R17648 gnd.n6899 gnd.n6898 19.3944
R17649 gnd.n6898 gnd.n6897 19.3944
R17650 gnd.n6897 gnd.n895 19.3944
R17651 gnd.n6891 gnd.n895 19.3944
R17652 gnd.n6891 gnd.n6890 19.3944
R17653 gnd.n6890 gnd.n6889 19.3944
R17654 gnd.n6889 gnd.n903 19.3944
R17655 gnd.n6883 gnd.n903 19.3944
R17656 gnd.n6883 gnd.n6882 19.3944
R17657 gnd.n6882 gnd.n6881 19.3944
R17658 gnd.n6881 gnd.n911 19.3944
R17659 gnd.n6875 gnd.n911 19.3944
R17660 gnd.n6875 gnd.n6874 19.3944
R17661 gnd.n6874 gnd.n6873 19.3944
R17662 gnd.n6873 gnd.n919 19.3944
R17663 gnd.n6867 gnd.n919 19.3944
R17664 gnd.n6867 gnd.n6866 19.3944
R17665 gnd.n6866 gnd.n6865 19.3944
R17666 gnd.n6865 gnd.n927 19.3944
R17667 gnd.n6859 gnd.n927 19.3944
R17668 gnd.n6859 gnd.n6858 19.3944
R17669 gnd.n6858 gnd.n6857 19.3944
R17670 gnd.n6857 gnd.n935 19.3944
R17671 gnd.n6851 gnd.n935 19.3944
R17672 gnd.n6851 gnd.n6850 19.3944
R17673 gnd.n6850 gnd.n6849 19.3944
R17674 gnd.n6849 gnd.n943 19.3944
R17675 gnd.n6843 gnd.n943 19.3944
R17676 gnd.n6843 gnd.n6842 19.3944
R17677 gnd.n6842 gnd.n6841 19.3944
R17678 gnd.n6841 gnd.n951 19.3944
R17679 gnd.n4225 gnd.n951 19.3944
R17680 gnd.n4491 gnd.n4483 19.3944
R17681 gnd.n4487 gnd.n4483 19.3944
R17682 gnd.n4487 gnd.n4486 19.3944
R17683 gnd.n4486 gnd.n3907 19.3944
R17684 gnd.n4827 gnd.n3907 19.3944
R17685 gnd.n4827 gnd.n3905 19.3944
R17686 gnd.n4831 gnd.n3905 19.3944
R17687 gnd.n4831 gnd.n3903 19.3944
R17688 gnd.n4835 gnd.n3903 19.3944
R17689 gnd.n4835 gnd.n3900 19.3944
R17690 gnd.n4980 gnd.n3900 19.3944
R17691 gnd.n4980 gnd.n3901 19.3944
R17692 gnd.n4976 gnd.n3901 19.3944
R17693 gnd.n4976 gnd.n4975 19.3944
R17694 gnd.n4975 gnd.n4974 19.3944
R17695 gnd.n4974 gnd.n4840 19.3944
R17696 gnd.n4970 gnd.n4840 19.3944
R17697 gnd.n4970 gnd.n4969 19.3944
R17698 gnd.n4969 gnd.n4968 19.3944
R17699 gnd.n4968 gnd.n4843 19.3944
R17700 gnd.n4964 gnd.n4843 19.3944
R17701 gnd.n4964 gnd.n4963 19.3944
R17702 gnd.n4963 gnd.n4962 19.3944
R17703 gnd.n4962 gnd.n4849 19.3944
R17704 gnd.n4958 gnd.n4849 19.3944
R17705 gnd.n4958 gnd.n4957 19.3944
R17706 gnd.n4957 gnd.n4956 19.3944
R17707 gnd.n4956 gnd.n4853 19.3944
R17708 gnd.n4952 gnd.n4853 19.3944
R17709 gnd.n4952 gnd.n4951 19.3944
R17710 gnd.n4951 gnd.n4950 19.3944
R17711 gnd.n4950 gnd.n4857 19.3944
R17712 gnd.n4946 gnd.n4857 19.3944
R17713 gnd.n4946 gnd.n4945 19.3944
R17714 gnd.n4945 gnd.n4944 19.3944
R17715 gnd.n4944 gnd.n4860 19.3944
R17716 gnd.n4940 gnd.n4860 19.3944
R17717 gnd.n4940 gnd.n4939 19.3944
R17718 gnd.n4939 gnd.n4938 19.3944
R17719 gnd.n4938 gnd.n4866 19.3944
R17720 gnd.n4934 gnd.n4866 19.3944
R17721 gnd.n4934 gnd.n4933 19.3944
R17722 gnd.n4933 gnd.n4932 19.3944
R17723 gnd.n4932 gnd.n4869 19.3944
R17724 gnd.n4928 gnd.n4869 19.3944
R17725 gnd.n4928 gnd.n4927 19.3944
R17726 gnd.n4927 gnd.n4926 19.3944
R17727 gnd.n4926 gnd.n4873 19.3944
R17728 gnd.n4922 gnd.n4873 19.3944
R17729 gnd.n4922 gnd.n4921 19.3944
R17730 gnd.n4921 gnd.n4920 19.3944
R17731 gnd.n4920 gnd.n4878 19.3944
R17732 gnd.n4916 gnd.n4878 19.3944
R17733 gnd.n4916 gnd.n4915 19.3944
R17734 gnd.n4915 gnd.n4914 19.3944
R17735 gnd.n4914 gnd.n4882 19.3944
R17736 gnd.n4910 gnd.n4882 19.3944
R17737 gnd.n4910 gnd.n4909 19.3944
R17738 gnd.n4909 gnd.n4908 19.3944
R17739 gnd.n4908 gnd.n4887 19.3944
R17740 gnd.n4904 gnd.n4887 19.3944
R17741 gnd.n4904 gnd.n4903 19.3944
R17742 gnd.n4903 gnd.n4902 19.3944
R17743 gnd.n4902 gnd.n4892 19.3944
R17744 gnd.n4898 gnd.n4892 19.3944
R17745 gnd.n4898 gnd.n4897 19.3944
R17746 gnd.n4897 gnd.n4896 19.3944
R17747 gnd.n4896 gnd.n3542 19.3944
R17748 gnd.n5407 gnd.n3542 19.3944
R17749 gnd.n5407 gnd.n3539 19.3944
R17750 gnd.n5412 gnd.n3539 19.3944
R17751 gnd.n5412 gnd.n3540 19.3944
R17752 gnd.n3540 gnd.n3443 19.3944
R17753 gnd.n5555 gnd.n3443 19.3944
R17754 gnd.n5555 gnd.n3441 19.3944
R17755 gnd.n5559 gnd.n3441 19.3944
R17756 gnd.n5559 gnd.n3431 19.3944
R17757 gnd.n5574 gnd.n3431 19.3944
R17758 gnd.n5574 gnd.n3429 19.3944
R17759 gnd.n5578 gnd.n3429 19.3944
R17760 gnd.n5578 gnd.n3011 19.3944
R17761 gnd.n6200 gnd.n3011 19.3944
R17762 gnd.n6197 gnd.n6196 19.3944
R17763 gnd.n6196 gnd.n6195 19.3944
R17764 gnd.n6195 gnd.n3016 19.3944
R17765 gnd.n6191 gnd.n3016 19.3944
R17766 gnd.n6191 gnd.n6190 19.3944
R17767 gnd.n6190 gnd.n6189 19.3944
R17768 gnd.n6189 gnd.n3021 19.3944
R17769 gnd.n6184 gnd.n3021 19.3944
R17770 gnd.n6184 gnd.n6183 19.3944
R17771 gnd.n6183 gnd.n3026 19.3944
R17772 gnd.n6176 gnd.n3026 19.3944
R17773 gnd.n6176 gnd.n6175 19.3944
R17774 gnd.n6175 gnd.n3035 19.3944
R17775 gnd.n6168 gnd.n3035 19.3944
R17776 gnd.n6168 gnd.n6167 19.3944
R17777 gnd.n6167 gnd.n3043 19.3944
R17778 gnd.n6160 gnd.n3043 19.3944
R17779 gnd.n6160 gnd.n6159 19.3944
R17780 gnd.n6159 gnd.n3051 19.3944
R17781 gnd.n6152 gnd.n3051 19.3944
R17782 gnd.n6152 gnd.n6151 19.3944
R17783 gnd.n6151 gnd.n3059 19.3944
R17784 gnd.n6144 gnd.n3059 19.3944
R17785 gnd.n6144 gnd.n6143 19.3944
R17786 gnd.n3417 gnd.n3396 19.3944
R17787 gnd.n5686 gnd.n3396 19.3944
R17788 gnd.n5686 gnd.n5685 19.3944
R17789 gnd.n3782 gnd.t387 19.1199
R17790 gnd.n3763 gnd.n3755 19.1199
R17791 gnd.n3714 gnd.n3712 19.1199
R17792 gnd.n3682 gnd.n3674 19.1199
R17793 gnd.n3631 gnd.n3630 19.1199
R17794 gnd.n3614 gnd.t342 19.1199
R17795 gnd.n1836 gnd.t358 18.8012
R17796 gnd.n1873 gnd.t377 18.8012
R17797 gnd.n1706 gnd.n1705 18.4825
R17798 gnd.n6837 gnd.n953 18.4825
R17799 gnd.n6082 gnd.n6081 18.4247
R17800 gnd.n6395 gnd.n6394 18.4247
R17801 gnd.n6324 gnd.n6323 18.2639
R17802 gnd.n5540 gnd.n3480 18.2639
R17803 gnd.n6140 gnd.n6139 18.2308
R17804 gnd.n4573 gnd.n3955 18.2308
R17805 gnd.n7789 gnd.n7740 18.2308
R17806 gnd.n4160 gnd.n4159 18.2308
R17807 gnd.t208 gnd.n1385 18.1639
R17808 gnd.t398 gnd.n2901 18.1639
R17809 gnd.n5415 gnd.t344 18.1639
R17810 gnd.n3823 gnd.n2912 17.8452
R17811 gnd.n5052 gnd.n3798 17.8452
R17812 gnd.n5176 gnd.n3718 17.8452
R17813 gnd.n5238 gnd.n3660 17.8452
R17814 gnd.n5358 gnd.n3585 17.8452
R17815 gnd.t289 gnd.n3544 17.8452
R17816 gnd.n5405 gnd.n3545 17.8452
R17817 gnd.n1414 gnd.t394 17.5266
R17818 gnd.t354 gnd.n3742 17.5266
R17819 gnd.n4876 gnd.t402 17.5266
R17820 gnd.n1825 gnd.t381 16.8893
R17821 gnd.n6064 gnd.n6061 16.6793
R17822 gnd.n7901 gnd.n7898 16.6793
R17823 gnd.n6672 gnd.n6669 16.6793
R17824 gnd.n4665 gnd.n4664 16.6793
R17825 gnd.n4199 gnd.n2542 16.5706
R17826 gnd.n6573 gnd.n2549 16.5706
R17827 gnd.n4218 gnd.n4217 16.5706
R17828 gnd.n6567 gnd.n2559 16.5706
R17829 gnd.n4211 gnd.n2562 16.5706
R17830 gnd.n6561 gnd.n2569 16.5706
R17831 gnd.n4248 gnd.n2572 16.5706
R17832 gnd.n4257 gnd.n2582 16.5706
R17833 gnd.n6549 gnd.n2589 16.5706
R17834 gnd.n4282 gnd.n4281 16.5706
R17835 gnd.n6543 gnd.n2598 16.5706
R17836 gnd.n4275 gnd.n2601 16.5706
R17837 gnd.n6537 gnd.n2608 16.5706
R17838 gnd.n4307 gnd.n2611 16.5706
R17839 gnd.n4315 gnd.n4040 16.5706
R17840 gnd.n4331 gnd.n4030 16.5706
R17841 gnd.n4337 gnd.n4023 16.5706
R17842 gnd.n4025 gnd.n4016 16.5706
R17843 gnd.n6530 gnd.n2624 16.5706
R17844 gnd.n4376 gnd.n2627 16.5706
R17845 gnd.n4384 gnd.n2638 16.5706
R17846 gnd.n6518 gnd.n2645 16.5706
R17847 gnd.n4390 gnd.n4004 16.5706
R17848 gnd.n6512 gnd.n2654 16.5706
R17849 gnd.n6506 gnd.n2665 16.5706
R17850 gnd.n4433 gnd.n2668 16.5706
R17851 gnd.n4405 gnd.n2677 16.5706
R17852 gnd.n6494 gnd.n2685 16.5706
R17853 gnd.n4410 gnd.n4409 16.5706
R17854 gnd.n6488 gnd.n2694 16.5706
R17855 gnd.n6482 gnd.n2705 16.5706
R17856 gnd.n4457 gnd.n2708 16.5706
R17857 gnd.n4465 gnd.n2717 16.5706
R17858 gnd.n6470 gnd.n2725 16.5706
R17859 gnd.n4738 gnd.n4737 16.5706
R17860 gnd.n6464 gnd.n2734 16.5706
R17861 gnd.n4472 gnd.n2737 16.5706
R17862 gnd.n6458 gnd.n2745 16.5706
R17863 gnd.n4724 gnd.n2748 16.5706
R17864 gnd.n6452 gnd.n2755 16.5706
R17865 gnd.n4764 gnd.n2758 16.5706
R17866 gnd.n5024 gnd.n5023 16.5706
R17867 gnd.n5135 gnd.n3738 16.5706
R17868 gnd.n5148 gnd.n5146 16.5706
R17869 gnd.n5257 gnd.n3656 16.5706
R17870 gnd.n5269 gnd.n5268 16.5706
R17871 gnd.n3575 gnd.n3568 16.5706
R17872 gnd.n5395 gnd.n5394 16.5706
R17873 gnd.n6013 gnd.n3187 16.5706
R17874 gnd.n5670 gnd.n5669 16.5706
R17875 gnd.n6005 gnd.n3196 16.5706
R17876 gnd.n5693 gnd.n3209 16.5706
R17877 gnd.n5999 gnd.n3212 16.5706
R17878 gnd.n5701 gnd.n3222 16.5706
R17879 gnd.n5993 gnd.n3225 16.5706
R17880 gnd.n5708 gnd.n3233 16.5706
R17881 gnd.n5987 gnd.n3236 16.5706
R17882 gnd.n5981 gnd.n3246 16.5706
R17883 gnd.n5723 gnd.n3254 16.5706
R17884 gnd.n5731 gnd.n3263 16.5706
R17885 gnd.n5969 gnd.n3266 16.5706
R17886 gnd.n5738 gnd.n3274 16.5706
R17887 gnd.n5963 gnd.n3277 16.5706
R17888 gnd.n5957 gnd.n3287 16.5706
R17889 gnd.n5753 gnd.n3295 16.5706
R17890 gnd.n5761 gnd.n3304 16.5706
R17891 gnd.n5945 gnd.n3307 16.5706
R17892 gnd.n5768 gnd.n3316 16.5706
R17893 gnd.n5939 gnd.n3319 16.5706
R17894 gnd.n5933 gnd.n3329 16.5706
R17895 gnd.n5928 gnd.n5927 16.5706
R17896 gnd.n5920 gnd.n3340 16.5706
R17897 gnd.n5919 gnd.n3343 16.5706
R17898 gnd.n5914 gnd.n3353 16.5706
R17899 gnd.n3362 gnd.n3360 16.5706
R17900 gnd.n8067 gnd.n103 16.5706
R17901 gnd.n5902 gnd.n5899 16.5706
R17902 gnd.n5829 gnd.n118 16.5706
R17903 gnd.n8059 gnd.n121 16.5706
R17904 gnd.n5891 gnd.n5890 16.5706
R17905 gnd.n8053 gnd.n132 16.5706
R17906 gnd.n5884 gnd.n139 16.5706
R17907 gnd.n5878 gnd.n148 16.5706
R17908 gnd.n8041 gnd.n151 16.5706
R17909 gnd.n5872 gnd.n159 16.5706
R17910 gnd.n8035 gnd.n162 16.5706
R17911 gnd.n7716 gnd.n7715 16.5706
R17912 gnd.n8029 gnd.n171 16.5706
R17913 gnd.n7821 gnd.n179 16.5706
R17914 gnd.n1641 gnd.t222 16.2519
R17915 gnd.n1870 gnd.t4 16.2519
R17916 gnd.n4346 gnd.t98 16.2519
R17917 gnd.n4783 gnd.t282 16.2519
R17918 gnd.t258 gnd.n3006 16.2519
R17919 gnd.n3339 gnd.t65 16.2519
R17920 gnd.t364 gnd.n5064 15.9333
R17921 gnd.n3603 gnd.t360 15.9333
R17922 gnd.n256 gnd.n249 15.9333
R17923 gnd.n2309 gnd.n2307 15.6674
R17924 gnd.n2277 gnd.n2275 15.6674
R17925 gnd.n2245 gnd.n2243 15.6674
R17926 gnd.n2214 gnd.n2212 15.6674
R17927 gnd.n2182 gnd.n2180 15.6674
R17928 gnd.n2150 gnd.n2148 15.6674
R17929 gnd.n2118 gnd.n2116 15.6674
R17930 gnd.n2087 gnd.n2085 15.6674
R17931 gnd.n1632 gnd.t222 15.6146
R17932 gnd.n2346 gnd.t338 15.6146
R17933 gnd.t307 gnd.n1001 15.6146
R17934 gnd.t105 gnd.n2657 15.6146
R17935 gnd.t282 gnd.n3918 15.6146
R17936 gnd.n5580 gnd.t258 15.6146
R17937 gnd.n3372 gnd.t70 15.6146
R17938 gnd.n6021 gnd.n6016 15.3217
R17939 gnd.n7856 gnd.n351 15.3217
R17940 gnd.n6629 gnd.n2459 15.3217
R17941 gnd.n4716 gnd.n4714 15.3217
R17942 gnd.n4229 gnd.n2532 15.296
R17943 gnd.n6579 gnd.n2542 15.296
R17944 gnd.n4199 gnd.n2549 15.296
R17945 gnd.n4217 gnd.n2559 15.296
R17946 gnd.n6567 gnd.n2562 15.296
R17947 gnd.n6561 gnd.n2572 15.296
R17948 gnd.n4248 gnd.n4247 15.296
R17949 gnd.n6555 gnd.n2582 15.296
R17950 gnd.n4257 gnd.n2589 15.296
R17951 gnd.n4281 gnd.n2598 15.296
R17952 gnd.n6543 gnd.n2601 15.296
R17953 gnd.n6537 gnd.n2611 15.296
R17954 gnd.n4307 gnd.n4306 15.296
R17955 gnd.n4266 gnd.n4040 15.296
R17956 gnd.n4315 gnd.n4030 15.296
R17957 gnd.n4337 gnd.n4025 15.296
R17958 gnd.n4346 gnd.n4016 15.296
R17959 gnd.n4345 gnd.n2624 15.296
R17960 gnd.n6530 gnd.n2627 15.296
R17961 gnd.n4376 gnd.n4375 15.296
R17962 gnd.n6524 gnd.n2638 15.296
R17963 gnd.n4384 gnd.n2645 15.296
R17964 gnd.n4390 gnd.n2654 15.296
R17965 gnd.n6512 gnd.n2657 15.296
R17966 gnd.n4398 gnd.n2665 15.296
R17967 gnd.n6506 gnd.n2668 15.296
R17968 gnd.n4434 gnd.n4433 15.296
R17969 gnd.n6500 gnd.n2677 15.296
R17970 gnd.n4405 gnd.n2685 15.296
R17971 gnd.n4410 gnd.n2694 15.296
R17972 gnd.n6488 gnd.n2697 15.296
R17973 gnd.n4419 gnd.n2705 15.296
R17974 gnd.n6482 gnd.n2708 15.296
R17975 gnd.n4457 gnd.n4456 15.296
R17976 gnd.n6476 gnd.n2717 15.296
R17977 gnd.n4465 gnd.n2725 15.296
R17978 gnd.n4737 gnd.n2734 15.296
R17979 gnd.n6464 gnd.n2737 15.296
R17980 gnd.n4472 gnd.n2745 15.296
R17981 gnd.n6458 gnd.n2748 15.296
R17982 gnd.n6452 gnd.n2758 15.296
R17983 gnd.n4764 gnd.n4763 15.296
R17984 gnd.n5004 gnd.n5003 15.296
R17985 gnd.n5394 gnd.n3556 15.296
R17986 gnd.n6013 gnd.n3185 15.296
R17987 gnd.n5669 gnd.n3187 15.296
R17988 gnd.n5693 gnd.n3196 15.296
R17989 gnd.n5999 gnd.n3209 15.296
R17990 gnd.n5701 gnd.n3212 15.296
R17991 gnd.n5993 gnd.n3222 15.296
R17992 gnd.n5987 gnd.n3233 15.296
R17993 gnd.n5716 gnd.n3236 15.296
R17994 gnd.n5981 gnd.n3243 15.296
R17995 gnd.n5723 gnd.n3246 15.296
R17996 gnd.n5975 gnd.n3254 15.296
R17997 gnd.n5731 gnd.n3381 15.296
R17998 gnd.n5969 gnd.n3263 15.296
R17999 gnd.n5963 gnd.n3274 15.296
R18000 gnd.n5746 gnd.n3277 15.296
R18001 gnd.n5957 gnd.n3284 15.296
R18002 gnd.n5753 gnd.n3287 15.296
R18003 gnd.n5951 gnd.n3295 15.296
R18004 gnd.n5761 gnd.n3372 15.296
R18005 gnd.n5945 gnd.n3304 15.296
R18006 gnd.n5939 gnd.n3316 15.296
R18007 gnd.n5788 gnd.n3319 15.296
R18008 gnd.n5933 gnd.n3326 15.296
R18009 gnd.n5928 gnd.n3329 15.296
R18010 gnd.n5927 gnd.n3333 15.296
R18011 gnd.n3340 gnd.n3339 15.296
R18012 gnd.n5920 gnd.n5919 15.296
R18013 gnd.n3362 gnd.n3353 15.296
R18014 gnd.n5908 gnd.n3360 15.296
R18015 gnd.n8067 gnd.n101 15.296
R18016 gnd.n5902 gnd.n103 15.296
R18017 gnd.n8059 gnd.n118 15.296
R18018 gnd.n5890 gnd.n121 15.296
R18019 gnd.n5884 gnd.n132 15.296
R18020 gnd.n8047 gnd.n139 15.296
R18021 gnd.n5878 gnd.n5862 15.296
R18022 gnd.n8041 gnd.n148 15.296
R18023 gnd.n8035 gnd.n159 15.296
R18024 gnd.n7716 gnd.n162 15.296
R18025 gnd.n7821 gnd.n171 15.296
R18026 gnd.n8023 gnd.n179 15.296
R18027 gnd.n7708 gnd.n188 15.296
R18028 gnd.n3465 gnd.n3464 15.0827
R18029 gnd.n2883 gnd.n2878 15.0481
R18030 gnd.n3475 gnd.n3474 15.0481
R18031 gnd.n1139 gnd.t359 14.9773
R18032 gnd.t27 gnd.n2608 14.9773
R18033 gnd.t76 gnd.n2697 14.9773
R18034 gnd.n3381 gnd.t31 14.9773
R18035 gnd.n5899 gnd.t82 14.9773
R18036 gnd.n5033 gnd.t2 14.6587
R18037 gnd.n5366 gnd.t372 14.6587
R18038 gnd.t0 gnd.n955 14.34
R18039 gnd.n1112 gnd.t395 14.34
R18040 gnd.t53 gnd.n2569 14.34
R18041 gnd.t29 gnd.n151 14.34
R18042 gnd.n6312 gnd.n2912 14.0214
R18043 gnd.n5052 gnd.t348 14.0214
R18044 gnd.n5117 gnd.n5115 14.0214
R18045 gnd.n5176 gnd.n5175 14.0214
R18046 gnd.n5239 gnd.n5238 14.0214
R18047 gnd.n5294 gnd.n5293 14.0214
R18048 gnd.t365 gnd.n5358 14.0214
R18049 gnd.n1794 gnd.t362 13.7027
R18050 gnd.n5013 gnd.t349 13.7027
R18051 gnd.t390 gnd.n3553 13.7027
R18052 gnd.n1498 gnd.n1497 13.5763
R18053 gnd.n6800 gnd.n1014 13.5763
R18054 gnd.n1706 gnd.n1444 13.384
R18055 gnd.n4983 gnd.t269 13.384
R18056 gnd.t262 gnd.n3545 13.384
R18057 gnd.n2894 gnd.n2875 13.1884
R18058 gnd.n2889 gnd.n2888 13.1884
R18059 gnd.n2888 gnd.n2887 13.1884
R18060 gnd.n3468 gnd.n3463 13.1884
R18061 gnd.n3469 gnd.n3468 13.1884
R18062 gnd.n2890 gnd.n2877 13.146
R18063 gnd.n2886 gnd.n2877 13.146
R18064 gnd.n3467 gnd.n3466 13.146
R18065 gnd.n3467 gnd.n3462 13.146
R18066 gnd.n2310 gnd.n2306 12.8005
R18067 gnd.n2278 gnd.n2274 12.8005
R18068 gnd.n2246 gnd.n2242 12.8005
R18069 gnd.n2215 gnd.n2211 12.8005
R18070 gnd.n2183 gnd.n2179 12.8005
R18071 gnd.n2151 gnd.n2147 12.8005
R18072 gnd.n2119 gnd.n2115 12.8005
R18073 gnd.n2088 gnd.n2084 12.8005
R18074 gnd.n6318 gnd.n2901 12.7467
R18075 gnd.n3793 gnd.n3788 12.7467
R18076 gnd.n5099 gnd.n3763 12.7467
R18077 gnd.n3712 gnd.n3707 12.7467
R18078 gnd.n5189 gnd.t386 12.7467
R18079 gnd.n5223 gnd.t346 12.7467
R18080 gnd.n5222 gnd.n3682 12.7467
R18081 gnd.n3630 gnd.n3625 12.7467
R18082 gnd.n3596 gnd.n3594 12.7467
R18083 gnd.n6597 gnd.t37 12.4281
R18084 gnd.n6476 gnd.t56 12.4281
R18085 gnd.t212 gnd.n3793 12.4281
R18086 gnd.n3594 gnd.t392 12.4281
R18087 gnd.n5716 gnd.t14 12.4281
R18088 gnd.n8005 gnd.t124 12.4281
R18089 gnd.n1497 gnd.n1492 12.4126
R18090 gnd.n6796 gnd.n1014 12.4126
R18091 gnd.n6387 gnd.n6324 12.1761
R18092 gnd.n3481 gnd.n3480 12.1761
R18093 gnd.n2314 gnd.n2313 12.0247
R18094 gnd.n2282 gnd.n2281 12.0247
R18095 gnd.n2250 gnd.n2249 12.0247
R18096 gnd.n2219 gnd.n2218 12.0247
R18097 gnd.n2187 gnd.n2186 12.0247
R18098 gnd.n2155 gnd.n2154 12.0247
R18099 gnd.n2123 gnd.n2122 12.0247
R18100 gnd.n2092 gnd.n2091 12.0247
R18101 gnd.n6573 gnd.t85 11.7908
R18102 gnd.n6500 gnd.t46 11.7908
R18103 gnd.t251 gnd.n2755 11.7908
R18104 gnd.n5670 gnd.t226 11.7908
R18105 gnd.n5746 gnd.t16 11.7908
R18106 gnd.n8029 gnd.t12 11.7908
R18107 gnd.n5071 gnd.n3783 11.4721
R18108 gnd.n5091 gnd.n5089 11.4721
R18109 gnd.n5195 gnd.n3703 11.4721
R18110 gnd.n5214 gnd.n5213 11.4721
R18111 gnd.n5315 gnd.n3620 11.4721
R18112 gnd.n5334 gnd.n3600 11.4721
R18113 gnd.n5545 gnd.t292 11.4721
R18114 gnd.n5553 gnd.n3445 11.4721
R18115 gnd.n2317 gnd.n2304 11.249
R18116 gnd.n2285 gnd.n2272 11.249
R18117 gnd.n2253 gnd.n2240 11.249
R18118 gnd.n2222 gnd.n2209 11.249
R18119 gnd.n2190 gnd.n2177 11.249
R18120 gnd.n2158 gnd.n2145 11.249
R18121 gnd.n2126 gnd.n2113 11.249
R18122 gnd.n2095 gnd.n2082 11.249
R18123 gnd.n1784 gnd.t362 11.1535
R18124 gnd.n6549 gnd.t23 11.1535
R18125 gnd.n6524 gnd.t58 11.1535
R18126 gnd.n3910 gnd.t366 11.1535
R18127 gnd.n5561 gnd.t370 11.1535
R18128 gnd.n5788 gnd.t10 11.1535
R18129 gnd.n8053 gnd.t41 11.1535
R18130 gnd.n5003 gnd.t248 10.8348
R18131 gnd.n5076 gnd.t353 10.8348
R18132 gnd.n5100 gnd.t353 10.8348
R18133 gnd.n5307 gnd.t352 10.8348
R18134 gnd.t352 gnd.n5306 10.8348
R18135 gnd.t242 gnd.n3445 10.8348
R18136 gnd.n6024 gnd.n6021 10.6672
R18137 gnd.n7859 gnd.n7856 10.6672
R18138 gnd.n6632 gnd.n6629 10.6672
R18139 gnd.n4714 gnd.n4713 10.6672
R18140 gnd.n5475 gnd.n3508 10.6151
R18141 gnd.n5475 gnd.n5474 10.6151
R18142 gnd.n5472 gnd.n3512 10.6151
R18143 gnd.n5467 gnd.n3512 10.6151
R18144 gnd.n5467 gnd.n5466 10.6151
R18145 gnd.n5466 gnd.n5465 10.6151
R18146 gnd.n5465 gnd.n3515 10.6151
R18147 gnd.n5460 gnd.n3515 10.6151
R18148 gnd.n5460 gnd.n5459 10.6151
R18149 gnd.n5459 gnd.n5458 10.6151
R18150 gnd.n5458 gnd.n3518 10.6151
R18151 gnd.n5453 gnd.n3518 10.6151
R18152 gnd.n5453 gnd.n5452 10.6151
R18153 gnd.n5452 gnd.n5451 10.6151
R18154 gnd.n5451 gnd.n3521 10.6151
R18155 gnd.n5446 gnd.n3521 10.6151
R18156 gnd.n5446 gnd.n5445 10.6151
R18157 gnd.n5445 gnd.n5444 10.6151
R18158 gnd.n5444 gnd.n3524 10.6151
R18159 gnd.n5439 gnd.n3524 10.6151
R18160 gnd.n5439 gnd.n5438 10.6151
R18161 gnd.n5438 gnd.n5437 10.6151
R18162 gnd.n5437 gnd.n3527 10.6151
R18163 gnd.n5432 gnd.n3527 10.6151
R18164 gnd.n5432 gnd.n5431 10.6151
R18165 gnd.n5431 gnd.n5430 10.6151
R18166 gnd.n5430 gnd.n3530 10.6151
R18167 gnd.n5425 gnd.n3530 10.6151
R18168 gnd.n5425 gnd.n5424 10.6151
R18169 gnd.n5424 gnd.n5423 10.6151
R18170 gnd.n3895 gnd.n3894 10.6151
R18171 gnd.n3896 gnd.n3895 10.6151
R18172 gnd.n3897 gnd.n3896 10.6151
R18173 gnd.n3897 gnd.n3826 10.6151
R18174 gnd.n4992 gnd.n3826 10.6151
R18175 gnd.n4993 gnd.n4992 10.6151
R18176 gnd.n4995 gnd.n4993 10.6151
R18177 gnd.n4995 gnd.n4994 10.6151
R18178 gnd.n4994 gnd.n3815 10.6151
R18179 gnd.n5015 gnd.n3815 10.6151
R18180 gnd.n5016 gnd.n5015 10.6151
R18181 gnd.n5021 gnd.n5016 10.6151
R18182 gnd.n5021 gnd.n5020 10.6151
R18183 gnd.n5020 gnd.n5019 10.6151
R18184 gnd.n5019 gnd.n5017 10.6151
R18185 gnd.n5017 gnd.n3790 10.6151
R18186 gnd.n5060 gnd.n3790 10.6151
R18187 gnd.n5061 gnd.n5060 10.6151
R18188 gnd.n5062 gnd.n5061 10.6151
R18189 gnd.n5062 gnd.n3779 10.6151
R18190 gnd.n5073 gnd.n3779 10.6151
R18191 gnd.n5074 gnd.n5073 10.6151
R18192 gnd.n5081 gnd.n5074 10.6151
R18193 gnd.n5081 gnd.n5080 10.6151
R18194 gnd.n5080 gnd.n5079 10.6151
R18195 gnd.n5079 gnd.n5078 10.6151
R18196 gnd.n5078 gnd.n5075 10.6151
R18197 gnd.n5075 gnd.n3753 10.6151
R18198 gnd.n5109 gnd.n3753 10.6151
R18199 gnd.n5110 gnd.n5109 10.6151
R18200 gnd.n5113 gnd.n5110 10.6151
R18201 gnd.n5113 gnd.n5112 10.6151
R18202 gnd.n5112 gnd.n5111 10.6151
R18203 gnd.n5111 gnd.n3736 10.6151
R18204 gnd.n5138 gnd.n3736 10.6151
R18205 gnd.n5139 gnd.n5138 10.6151
R18206 gnd.n5144 gnd.n5139 10.6151
R18207 gnd.n5144 gnd.n5143 10.6151
R18208 gnd.n5143 gnd.n5142 10.6151
R18209 gnd.n5142 gnd.n5140 10.6151
R18210 gnd.n5140 gnd.n3709 10.6151
R18211 gnd.n5184 gnd.n3709 10.6151
R18212 gnd.n5185 gnd.n5184 10.6151
R18213 gnd.n5186 gnd.n5185 10.6151
R18214 gnd.n5186 gnd.n3700 10.6151
R18215 gnd.n5197 gnd.n3700 10.6151
R18216 gnd.n5198 gnd.n5197 10.6151
R18217 gnd.n5205 gnd.n5198 10.6151
R18218 gnd.n5205 gnd.n5204 10.6151
R18219 gnd.n5204 gnd.n5203 10.6151
R18220 gnd.n5203 gnd.n5202 10.6151
R18221 gnd.n5202 gnd.n5199 10.6151
R18222 gnd.n5199 gnd.n3671 10.6151
R18223 gnd.n5232 gnd.n3671 10.6151
R18224 gnd.n5233 gnd.n5232 10.6151
R18225 gnd.n5236 gnd.n5233 10.6151
R18226 gnd.n5236 gnd.n5235 10.6151
R18227 gnd.n5235 gnd.n5234 10.6151
R18228 gnd.n5234 gnd.n3653 10.6151
R18229 gnd.n5260 gnd.n3653 10.6151
R18230 gnd.n5261 gnd.n5260 10.6151
R18231 gnd.n5266 gnd.n5261 10.6151
R18232 gnd.n5266 gnd.n5265 10.6151
R18233 gnd.n5265 gnd.n5264 10.6151
R18234 gnd.n5264 gnd.n5262 10.6151
R18235 gnd.n5262 gnd.n3627 10.6151
R18236 gnd.n5302 gnd.n3627 10.6151
R18237 gnd.n5303 gnd.n5302 10.6151
R18238 gnd.n5304 gnd.n5303 10.6151
R18239 gnd.n5304 gnd.n3616 10.6151
R18240 gnd.n5317 gnd.n3616 10.6151
R18241 gnd.n5318 gnd.n5317 10.6151
R18242 gnd.n5321 gnd.n5318 10.6151
R18243 gnd.n5321 gnd.n5320 10.6151
R18244 gnd.n5320 gnd.n5319 10.6151
R18245 gnd.n5319 gnd.n3592 10.6151
R18246 gnd.n5342 gnd.n3592 10.6151
R18247 gnd.n5343 gnd.n5342 10.6151
R18248 gnd.n5350 gnd.n5343 10.6151
R18249 gnd.n5350 gnd.n5349 10.6151
R18250 gnd.n5349 gnd.n5348 10.6151
R18251 gnd.n5348 gnd.n5347 10.6151
R18252 gnd.n5347 gnd.n5345 10.6151
R18253 gnd.n5345 gnd.n5344 10.6151
R18254 gnd.n5344 gnd.n3566 10.6151
R18255 gnd.n5376 gnd.n3566 10.6151
R18256 gnd.n5377 gnd.n5376 10.6151
R18257 gnd.n5378 gnd.n5377 10.6151
R18258 gnd.n5382 gnd.n5378 10.6151
R18259 gnd.n5383 gnd.n5382 10.6151
R18260 gnd.n5384 gnd.n5383 10.6151
R18261 gnd.n5384 gnd.n3535 10.6151
R18262 gnd.n5417 gnd.n3535 10.6151
R18263 gnd.n5418 gnd.n5417 10.6151
R18264 gnd.n5419 gnd.n5418 10.6151
R18265 gnd.n5419 gnd.n3533 10.6151
R18266 gnd.n3829 gnd.n2835 10.6151
R18267 gnd.n3832 gnd.n3829 10.6151
R18268 gnd.n3837 gnd.n3834 10.6151
R18269 gnd.n3838 gnd.n3837 10.6151
R18270 gnd.n3841 gnd.n3838 10.6151
R18271 gnd.n3842 gnd.n3841 10.6151
R18272 gnd.n3845 gnd.n3842 10.6151
R18273 gnd.n3846 gnd.n3845 10.6151
R18274 gnd.n3849 gnd.n3846 10.6151
R18275 gnd.n3850 gnd.n3849 10.6151
R18276 gnd.n3853 gnd.n3850 10.6151
R18277 gnd.n3854 gnd.n3853 10.6151
R18278 gnd.n3857 gnd.n3854 10.6151
R18279 gnd.n3858 gnd.n3857 10.6151
R18280 gnd.n3861 gnd.n3858 10.6151
R18281 gnd.n3862 gnd.n3861 10.6151
R18282 gnd.n3865 gnd.n3862 10.6151
R18283 gnd.n3866 gnd.n3865 10.6151
R18284 gnd.n3869 gnd.n3866 10.6151
R18285 gnd.n3870 gnd.n3869 10.6151
R18286 gnd.n3873 gnd.n3870 10.6151
R18287 gnd.n3874 gnd.n3873 10.6151
R18288 gnd.n3877 gnd.n3874 10.6151
R18289 gnd.n3878 gnd.n3877 10.6151
R18290 gnd.n3881 gnd.n3878 10.6151
R18291 gnd.n3882 gnd.n3881 10.6151
R18292 gnd.n3885 gnd.n3882 10.6151
R18293 gnd.n3886 gnd.n3885 10.6151
R18294 gnd.n3889 gnd.n3886 10.6151
R18295 gnd.n3890 gnd.n3889 10.6151
R18296 gnd.n6387 gnd.n6386 10.6151
R18297 gnd.n6386 gnd.n6385 10.6151
R18298 gnd.n6385 gnd.n6384 10.6151
R18299 gnd.n6384 gnd.n6382 10.6151
R18300 gnd.n6382 gnd.n6379 10.6151
R18301 gnd.n6379 gnd.n6378 10.6151
R18302 gnd.n6378 gnd.n6375 10.6151
R18303 gnd.n6375 gnd.n6374 10.6151
R18304 gnd.n6374 gnd.n6371 10.6151
R18305 gnd.n6371 gnd.n6370 10.6151
R18306 gnd.n6370 gnd.n6367 10.6151
R18307 gnd.n6367 gnd.n6366 10.6151
R18308 gnd.n6366 gnd.n6363 10.6151
R18309 gnd.n6363 gnd.n6362 10.6151
R18310 gnd.n6362 gnd.n6359 10.6151
R18311 gnd.n6359 gnd.n6358 10.6151
R18312 gnd.n6358 gnd.n6355 10.6151
R18313 gnd.n6355 gnd.n6354 10.6151
R18314 gnd.n6354 gnd.n6351 10.6151
R18315 gnd.n6351 gnd.n6350 10.6151
R18316 gnd.n6350 gnd.n6347 10.6151
R18317 gnd.n6347 gnd.n6346 10.6151
R18318 gnd.n6346 gnd.n6343 10.6151
R18319 gnd.n6343 gnd.n6342 10.6151
R18320 gnd.n6342 gnd.n6339 10.6151
R18321 gnd.n6339 gnd.n6338 10.6151
R18322 gnd.n6338 gnd.n6335 10.6151
R18323 gnd.n6335 gnd.n6334 10.6151
R18324 gnd.n6331 gnd.n6330 10.6151
R18325 gnd.n6330 gnd.n2836 10.6151
R18326 gnd.n5535 gnd.n3481 10.6151
R18327 gnd.n5535 gnd.n5534 10.6151
R18328 gnd.n5534 gnd.n5533 10.6151
R18329 gnd.n5533 gnd.n3483 10.6151
R18330 gnd.n5528 gnd.n3483 10.6151
R18331 gnd.n5528 gnd.n5527 10.6151
R18332 gnd.n5527 gnd.n5526 10.6151
R18333 gnd.n5526 gnd.n3486 10.6151
R18334 gnd.n5521 gnd.n3486 10.6151
R18335 gnd.n5521 gnd.n5520 10.6151
R18336 gnd.n5520 gnd.n5519 10.6151
R18337 gnd.n5519 gnd.n3489 10.6151
R18338 gnd.n5514 gnd.n3489 10.6151
R18339 gnd.n5514 gnd.n5513 10.6151
R18340 gnd.n5513 gnd.n5512 10.6151
R18341 gnd.n5512 gnd.n3492 10.6151
R18342 gnd.n5507 gnd.n3492 10.6151
R18343 gnd.n5507 gnd.n5506 10.6151
R18344 gnd.n5506 gnd.n5505 10.6151
R18345 gnd.n5505 gnd.n3495 10.6151
R18346 gnd.n5500 gnd.n3495 10.6151
R18347 gnd.n5500 gnd.n5499 10.6151
R18348 gnd.n5499 gnd.n5498 10.6151
R18349 gnd.n5498 gnd.n3498 10.6151
R18350 gnd.n5493 gnd.n3498 10.6151
R18351 gnd.n5493 gnd.n5492 10.6151
R18352 gnd.n5492 gnd.n5491 10.6151
R18353 gnd.n5491 gnd.n3501 10.6151
R18354 gnd.n5486 gnd.n5485 10.6151
R18355 gnd.n5485 gnd.n5484 10.6151
R18356 gnd.n6323 gnd.n6322 10.6151
R18357 gnd.n6322 gnd.n2895 10.6151
R18358 gnd.n4986 gnd.n2895 10.6151
R18359 gnd.n4987 gnd.n4986 10.6151
R18360 gnd.n4988 gnd.n4987 10.6151
R18361 gnd.n4988 gnd.n3821 10.6151
R18362 gnd.n4999 gnd.n3821 10.6151
R18363 gnd.n5000 gnd.n4999 10.6151
R18364 gnd.n5001 gnd.n5000 10.6151
R18365 gnd.n5001 gnd.n3811 10.6151
R18366 gnd.n5027 gnd.n3811 10.6151
R18367 gnd.n5028 gnd.n5027 10.6151
R18368 gnd.n5029 gnd.n5028 10.6151
R18369 gnd.n5029 gnd.n3796 10.6151
R18370 gnd.n5054 gnd.n3796 10.6151
R18371 gnd.n5055 gnd.n5054 10.6151
R18372 gnd.n5056 gnd.n5055 10.6151
R18373 gnd.n5056 gnd.n3785 10.6151
R18374 gnd.n5067 gnd.n3785 10.6151
R18375 gnd.n5068 gnd.n5067 10.6151
R18376 gnd.n5069 gnd.n5068 10.6151
R18377 gnd.n5069 gnd.n3773 10.6151
R18378 gnd.n5085 gnd.n3773 10.6151
R18379 gnd.n5086 gnd.n5085 10.6151
R18380 gnd.n5087 gnd.n5086 10.6151
R18381 gnd.n5087 gnd.n3759 10.6151
R18382 gnd.n5102 gnd.n3759 10.6151
R18383 gnd.n5103 gnd.n5102 10.6151
R18384 gnd.n5105 gnd.n5103 10.6151
R18385 gnd.n5105 gnd.n5104 10.6151
R18386 gnd.n5104 gnd.n3740 10.6151
R18387 gnd.n5131 gnd.n3740 10.6151
R18388 gnd.n5132 gnd.n5131 10.6151
R18389 gnd.n5133 gnd.n5132 10.6151
R18390 gnd.n5133 gnd.n3731 10.6151
R18391 gnd.n5151 gnd.n3731 10.6151
R18392 gnd.n5152 gnd.n5151 10.6151
R18393 gnd.n5153 gnd.n5152 10.6151
R18394 gnd.n5153 gnd.n3716 10.6151
R18395 gnd.n5178 gnd.n3716 10.6151
R18396 gnd.n5179 gnd.n5178 10.6151
R18397 gnd.n5180 gnd.n5179 10.6151
R18398 gnd.n5180 gnd.n3705 10.6151
R18399 gnd.n5191 gnd.n3705 10.6151
R18400 gnd.n5192 gnd.n5191 10.6151
R18401 gnd.n5193 gnd.n5192 10.6151
R18402 gnd.n5193 gnd.n3693 10.6151
R18403 gnd.n5209 gnd.n3693 10.6151
R18404 gnd.n5210 gnd.n5209 10.6151
R18405 gnd.n5211 gnd.n5210 10.6151
R18406 gnd.n5211 gnd.n3678 10.6151
R18407 gnd.n5225 gnd.n3678 10.6151
R18408 gnd.n5226 gnd.n5225 10.6151
R18409 gnd.n5228 gnd.n5226 10.6151
R18410 gnd.n5228 gnd.n5227 10.6151
R18411 gnd.n5227 gnd.n3658 10.6151
R18412 gnd.n5253 gnd.n3658 10.6151
R18413 gnd.n5254 gnd.n5253 10.6151
R18414 gnd.n5255 gnd.n5254 10.6151
R18415 gnd.n5255 gnd.n3648 10.6151
R18416 gnd.n5272 gnd.n3648 10.6151
R18417 gnd.n5273 gnd.n5272 10.6151
R18418 gnd.n5274 gnd.n5273 10.6151
R18419 gnd.n5274 gnd.n3633 10.6151
R18420 gnd.n5296 gnd.n3633 10.6151
R18421 gnd.n5297 gnd.n5296 10.6151
R18422 gnd.n5298 gnd.n5297 10.6151
R18423 gnd.n5298 gnd.n3623 10.6151
R18424 gnd.n5309 gnd.n3623 10.6151
R18425 gnd.n5310 gnd.n5309 10.6151
R18426 gnd.n5313 gnd.n5310 10.6151
R18427 gnd.n5313 gnd.n5312 10.6151
R18428 gnd.n5312 gnd.n5311 10.6151
R18429 gnd.n5311 gnd.n3598 10.6151
R18430 gnd.n5336 gnd.n3598 10.6151
R18431 gnd.n5337 gnd.n5336 10.6151
R18432 gnd.n5338 gnd.n5337 10.6151
R18433 gnd.n5338 gnd.n3587 10.6151
R18434 gnd.n5354 gnd.n3587 10.6151
R18435 gnd.n5355 gnd.n5354 10.6151
R18436 gnd.n5356 gnd.n5355 10.6151
R18437 gnd.n5356 gnd.n3570 10.6151
R18438 gnd.n5369 gnd.n3570 10.6151
R18439 gnd.n5370 gnd.n5369 10.6151
R18440 gnd.n5371 gnd.n5370 10.6151
R18441 gnd.n5371 gnd.n3559 10.6151
R18442 gnd.n5392 gnd.n3559 10.6151
R18443 gnd.n5392 gnd.n5391 10.6151
R18444 gnd.n5391 gnd.n5390 10.6151
R18445 gnd.n5390 gnd.n3560 10.6151
R18446 gnd.n3563 gnd.n3560 10.6151
R18447 gnd.n3563 gnd.n3562 10.6151
R18448 gnd.n3562 gnd.n3460 10.6151
R18449 gnd.n5542 gnd.n3460 10.6151
R18450 gnd.n5542 gnd.n5541 10.6151
R18451 gnd.n5541 gnd.n5540 10.6151
R18452 gnd.n1695 gnd.t400 10.5161
R18453 gnd.n2031 gnd.t0 10.5161
R18454 gnd.t395 gnd.n976 10.5161
R18455 gnd.n4266 gnd.t87 10.5161
R18456 gnd.n4331 gnd.t68 10.5161
R18457 gnd.n5914 gnd.t119 10.5161
R18458 gnd.n5908 gnd.t18 10.5161
R18459 gnd.n2318 gnd.n2302 10.4732
R18460 gnd.n2286 gnd.n2270 10.4732
R18461 gnd.n2254 gnd.n2238 10.4732
R18462 gnd.n2223 gnd.n2207 10.4732
R18463 gnd.n2191 gnd.n2175 10.4732
R18464 gnd.n2159 gnd.n2143 10.4732
R18465 gnd.n2127 gnd.n2111 10.4732
R18466 gnd.n2096 gnd.n2080 10.4732
R18467 gnd.n3783 gnd.n3782 10.1975
R18468 gnd.n3703 gnd.n3695 10.1975
R18469 gnd.n5214 gnd.n3688 10.1975
R18470 gnd.n3614 gnd.n3600 10.1975
R18471 gnd.t359 gnd.n1131 9.87883
R18472 gnd.n6555 gnd.t110 9.87883
R18473 gnd.n6518 gnd.t129 9.87883
R18474 gnd.n5768 gnd.t94 9.87883
R18475 gnd.n8047 gnd.t73 9.87883
R18476 gnd.n2322 gnd.n2321 9.69747
R18477 gnd.n2290 gnd.n2289 9.69747
R18478 gnd.n2258 gnd.n2257 9.69747
R18479 gnd.n2227 gnd.n2226 9.69747
R18480 gnd.n2195 gnd.n2194 9.69747
R18481 gnd.n2163 gnd.n2162 9.69747
R18482 gnd.n2131 gnd.n2130 9.69747
R18483 gnd.n2100 gnd.n2099 9.69747
R18484 gnd.n5127 gnd.t361 9.56018
R18485 gnd.n5277 gnd.t388 9.56018
R18486 gnd.n3456 gnd.t242 9.56018
R18487 gnd.n2328 gnd.n2327 9.45567
R18488 gnd.n2296 gnd.n2295 9.45567
R18489 gnd.n2264 gnd.n2263 9.45567
R18490 gnd.n2233 gnd.n2232 9.45567
R18491 gnd.n2201 gnd.n2200 9.45567
R18492 gnd.n2169 gnd.n2168 9.45567
R18493 gnd.n2137 gnd.n2136 9.45567
R18494 gnd.n2106 gnd.n2105 9.45567
R18495 gnd.n6061 gnd.n6060 9.30959
R18496 gnd.n7898 gnd.n331 9.30959
R18497 gnd.n6669 gnd.n6668 9.30959
R18498 gnd.n4668 gnd.n4665 9.30959
R18499 gnd.n2327 gnd.n2326 9.3005
R18500 gnd.n2300 gnd.n2299 9.3005
R18501 gnd.n2321 gnd.n2320 9.3005
R18502 gnd.n2319 gnd.n2318 9.3005
R18503 gnd.n2304 gnd.n2303 9.3005
R18504 gnd.n2313 gnd.n2312 9.3005
R18505 gnd.n2311 gnd.n2310 9.3005
R18506 gnd.n2295 gnd.n2294 9.3005
R18507 gnd.n2268 gnd.n2267 9.3005
R18508 gnd.n2289 gnd.n2288 9.3005
R18509 gnd.n2287 gnd.n2286 9.3005
R18510 gnd.n2272 gnd.n2271 9.3005
R18511 gnd.n2281 gnd.n2280 9.3005
R18512 gnd.n2279 gnd.n2278 9.3005
R18513 gnd.n2263 gnd.n2262 9.3005
R18514 gnd.n2236 gnd.n2235 9.3005
R18515 gnd.n2257 gnd.n2256 9.3005
R18516 gnd.n2255 gnd.n2254 9.3005
R18517 gnd.n2240 gnd.n2239 9.3005
R18518 gnd.n2249 gnd.n2248 9.3005
R18519 gnd.n2247 gnd.n2246 9.3005
R18520 gnd.n2232 gnd.n2231 9.3005
R18521 gnd.n2205 gnd.n2204 9.3005
R18522 gnd.n2226 gnd.n2225 9.3005
R18523 gnd.n2224 gnd.n2223 9.3005
R18524 gnd.n2209 gnd.n2208 9.3005
R18525 gnd.n2218 gnd.n2217 9.3005
R18526 gnd.n2216 gnd.n2215 9.3005
R18527 gnd.n2200 gnd.n2199 9.3005
R18528 gnd.n2173 gnd.n2172 9.3005
R18529 gnd.n2194 gnd.n2193 9.3005
R18530 gnd.n2192 gnd.n2191 9.3005
R18531 gnd.n2177 gnd.n2176 9.3005
R18532 gnd.n2186 gnd.n2185 9.3005
R18533 gnd.n2184 gnd.n2183 9.3005
R18534 gnd.n2168 gnd.n2167 9.3005
R18535 gnd.n2141 gnd.n2140 9.3005
R18536 gnd.n2162 gnd.n2161 9.3005
R18537 gnd.n2160 gnd.n2159 9.3005
R18538 gnd.n2145 gnd.n2144 9.3005
R18539 gnd.n2154 gnd.n2153 9.3005
R18540 gnd.n2152 gnd.n2151 9.3005
R18541 gnd.n2136 gnd.n2135 9.3005
R18542 gnd.n2109 gnd.n2108 9.3005
R18543 gnd.n2130 gnd.n2129 9.3005
R18544 gnd.n2128 gnd.n2127 9.3005
R18545 gnd.n2113 gnd.n2112 9.3005
R18546 gnd.n2122 gnd.n2121 9.3005
R18547 gnd.n2120 gnd.n2119 9.3005
R18548 gnd.n2105 gnd.n2104 9.3005
R18549 gnd.n2078 gnd.n2077 9.3005
R18550 gnd.n2099 gnd.n2098 9.3005
R18551 gnd.n2097 gnd.n2096 9.3005
R18552 gnd.n2082 gnd.n2081 9.3005
R18553 gnd.n2091 gnd.n2090 9.3005
R18554 gnd.n2089 gnd.n2088 9.3005
R18555 gnd.n6789 gnd.n6788 9.3005
R18556 gnd.n6787 gnd.n6755 9.3005
R18557 gnd.n6786 gnd.n6785 9.3005
R18558 gnd.n6782 gnd.n6756 9.3005
R18559 gnd.n6779 gnd.n6757 9.3005
R18560 gnd.n6778 gnd.n6758 9.3005
R18561 gnd.n6775 gnd.n6759 9.3005
R18562 gnd.n6774 gnd.n6760 9.3005
R18563 gnd.n6771 gnd.n6761 9.3005
R18564 gnd.n6770 gnd.n6762 9.3005
R18565 gnd.n6767 gnd.n6763 9.3005
R18566 gnd.n6766 gnd.n6764 9.3005
R18567 gnd.n1016 gnd.n1015 9.3005
R18568 gnd.n6797 gnd.n6796 9.3005
R18569 gnd.n6798 gnd.n1014 9.3005
R18570 gnd.n6800 gnd.n6799 9.3005
R18571 gnd.n6790 gnd.n6754 9.3005
R18572 gnd.n1714 gnd.n1713 9.3005
R18573 gnd.n1418 gnd.n1417 9.3005
R18574 gnd.n1741 gnd.n1740 9.3005
R18575 gnd.n1742 gnd.n1416 9.3005
R18576 gnd.n1746 gnd.n1743 9.3005
R18577 gnd.n1745 gnd.n1744 9.3005
R18578 gnd.n1390 gnd.n1389 9.3005
R18579 gnd.n1771 gnd.n1770 9.3005
R18580 gnd.n1772 gnd.n1388 9.3005
R18581 gnd.n1782 gnd.n1773 9.3005
R18582 gnd.n1781 gnd.n1774 9.3005
R18583 gnd.n1780 gnd.n1775 9.3005
R18584 gnd.n1778 gnd.n1777 9.3005
R18585 gnd.n1776 gnd.n1360 9.3005
R18586 gnd.n1358 gnd.n1357 9.3005
R18587 gnd.n1830 gnd.n1829 9.3005
R18588 gnd.n1831 gnd.n1356 9.3005
R18589 gnd.n1833 gnd.n1832 9.3005
R18590 gnd.n1227 gnd.n1226 9.3005
R18591 gnd.n1865 gnd.n1864 9.3005
R18592 gnd.n1866 gnd.n1225 9.3005
R18593 gnd.n1868 gnd.n1867 9.3005
R18594 gnd.n1206 gnd.n1205 9.3005
R18595 gnd.n1895 gnd.n1894 9.3005
R18596 gnd.n1896 gnd.n1204 9.3005
R18597 gnd.n1900 gnd.n1897 9.3005
R18598 gnd.n1899 gnd.n1898 9.3005
R18599 gnd.n1181 gnd.n1180 9.3005
R18600 gnd.n1944 gnd.n1943 9.3005
R18601 gnd.n1945 gnd.n1179 9.3005
R18602 gnd.n1949 gnd.n1946 9.3005
R18603 gnd.n1948 gnd.n1947 9.3005
R18604 gnd.n1154 gnd.n1153 9.3005
R18605 gnd.n1984 gnd.n1983 9.3005
R18606 gnd.n1985 gnd.n1152 9.3005
R18607 gnd.n1989 gnd.n1986 9.3005
R18608 gnd.n1988 gnd.n1987 9.3005
R18609 gnd.n1129 gnd.n1128 9.3005
R18610 gnd.n2045 gnd.n2044 9.3005
R18611 gnd.n2046 gnd.n1127 9.3005
R18612 gnd.n2054 gnd.n2047 9.3005
R18613 gnd.n2053 gnd.n2048 9.3005
R18614 gnd.n2052 gnd.n2050 9.3005
R18615 gnd.n2049 gnd.n970 9.3005
R18616 gnd.n6827 gnd.n971 9.3005
R18617 gnd.n6826 gnd.n972 9.3005
R18618 gnd.n6825 gnd.n973 9.3005
R18619 gnd.n994 gnd.n974 9.3005
R18620 gnd.n995 gnd.n993 9.3005
R18621 gnd.n6813 gnd.n996 9.3005
R18622 gnd.n6812 gnd.n997 9.3005
R18623 gnd.n6811 gnd.n998 9.3005
R18624 gnd.n6753 gnd.n999 9.3005
R18625 gnd.n1715 gnd.n1712 9.3005
R18626 gnd.n1497 gnd.n1456 9.3005
R18627 gnd.n1492 gnd.n1491 9.3005
R18628 gnd.n1490 gnd.n1457 9.3005
R18629 gnd.n1489 gnd.n1488 9.3005
R18630 gnd.n1485 gnd.n1458 9.3005
R18631 gnd.n1482 gnd.n1481 9.3005
R18632 gnd.n1480 gnd.n1459 9.3005
R18633 gnd.n1479 gnd.n1478 9.3005
R18634 gnd.n1475 gnd.n1460 9.3005
R18635 gnd.n1472 gnd.n1471 9.3005
R18636 gnd.n1470 gnd.n1461 9.3005
R18637 gnd.n1469 gnd.n1468 9.3005
R18638 gnd.n1465 gnd.n1463 9.3005
R18639 gnd.n1462 gnd.n1442 9.3005
R18640 gnd.n1709 gnd.n1441 9.3005
R18641 gnd.n1711 gnd.n1710 9.3005
R18642 gnd.n1499 gnd.n1498 9.3005
R18643 gnd.n1722 gnd.n1428 9.3005
R18644 gnd.n1729 gnd.n1429 9.3005
R18645 gnd.n1731 gnd.n1730 9.3005
R18646 gnd.n1732 gnd.n1409 9.3005
R18647 gnd.n1751 gnd.n1750 9.3005
R18648 gnd.n1753 gnd.n1401 9.3005
R18649 gnd.n1760 gnd.n1403 9.3005
R18650 gnd.n1761 gnd.n1398 9.3005
R18651 gnd.n1763 gnd.n1762 9.3005
R18652 gnd.n1399 gnd.n1384 9.3005
R18653 gnd.n1382 gnd.n1380 9.3005
R18654 gnd.n1789 gnd.n1788 9.3005
R18655 gnd.n1365 gnd.n1364 9.3005
R18656 gnd.n1822 gnd.n1810 9.3005
R18657 gnd.n1821 gnd.n1812 9.3005
R18658 gnd.n1820 gnd.n1813 9.3005
R18659 gnd.n1815 gnd.n1814 9.3005
R18660 gnd.n1348 gnd.n1236 9.3005
R18661 gnd.n1854 gnd.n1238 9.3005
R18662 gnd.n1855 gnd.n1234 9.3005
R18663 gnd.n1857 gnd.n1856 9.3005
R18664 gnd.n1222 gnd.n1217 9.3005
R18665 gnd.n1878 gnd.n1216 9.3005
R18666 gnd.n1881 gnd.n1880 9.3005
R18667 gnd.n1883 gnd.n1882 9.3005
R18668 gnd.n1886 gnd.n1199 9.3005
R18669 gnd.n1884 gnd.n1197 9.3005
R18670 gnd.n1907 gnd.n1195 9.3005
R18671 gnd.n1909 gnd.n1908 9.3005
R18672 gnd.n1172 gnd.n1171 9.3005
R18673 gnd.n1958 gnd.n1957 9.3005
R18674 gnd.n1959 gnd.n1165 9.3005
R18675 gnd.n1967 gnd.n1164 9.3005
R18676 gnd.n1970 gnd.n1969 9.3005
R18677 gnd.n1972 gnd.n1971 9.3005
R18678 gnd.n1975 gnd.n1148 9.3005
R18679 gnd.n1973 gnd.n1146 9.3005
R18680 gnd.n1995 gnd.n1144 9.3005
R18681 gnd.n1999 gnd.n1998 9.3005
R18682 gnd.n1997 gnd.n1120 9.3005
R18683 gnd.n2061 gnd.n1119 9.3005
R18684 gnd.n2064 gnd.n2063 9.3005
R18685 gnd.n1116 gnd.n1115 9.3005
R18686 gnd.n2068 gnd.n1117 9.3005
R18687 gnd.n2070 gnd.n2069 9.3005
R18688 gnd.n2072 gnd.n1114 9.3005
R18689 gnd.n2075 gnd.n2074 9.3005
R18690 gnd.n2333 gnd.n2332 9.3005
R18691 gnd.n2337 gnd.n2334 9.3005
R18692 gnd.n2339 gnd.n2338 9.3005
R18693 gnd.n2343 gnd.n2342 9.3005
R18694 gnd.n1010 gnd.n1008 9.3005
R18695 gnd.n6804 gnd.n6803 9.3005
R18696 gnd.n1720 gnd.n1719 9.3005
R18697 gnd.n1050 gnd.n1047 9.3005
R18698 gnd.n1052 gnd.n1051 9.3005
R18699 gnd.n1055 gnd.n1045 9.3005
R18700 gnd.n1059 gnd.n1058 9.3005
R18701 gnd.n1060 gnd.n1044 9.3005
R18702 gnd.n1062 gnd.n1061 9.3005
R18703 gnd.n1065 gnd.n1043 9.3005
R18704 gnd.n1069 gnd.n1068 9.3005
R18705 gnd.n1070 gnd.n1042 9.3005
R18706 gnd.n1072 gnd.n1071 9.3005
R18707 gnd.n1075 gnd.n1041 9.3005
R18708 gnd.n1079 gnd.n1078 9.3005
R18709 gnd.n1080 gnd.n1040 9.3005
R18710 gnd.n1082 gnd.n1081 9.3005
R18711 gnd.n1085 gnd.n1039 9.3005
R18712 gnd.n1089 gnd.n1088 9.3005
R18713 gnd.n1090 gnd.n1038 9.3005
R18714 gnd.n1092 gnd.n1091 9.3005
R18715 gnd.n1095 gnd.n1037 9.3005
R18716 gnd.n1099 gnd.n1098 9.3005
R18717 gnd.n1100 gnd.n1036 9.3005
R18718 gnd.n1102 gnd.n1101 9.3005
R18719 gnd.n1105 gnd.n1032 9.3005
R18720 gnd.n1108 gnd.n1107 9.3005
R18721 gnd.n1109 gnd.n1031 9.3005
R18722 gnd.n2353 gnd.n2352 9.3005
R18723 gnd.n1049 gnd.n1048 9.3005
R18724 gnd.n1249 gnd.n1245 9.3005
R18725 gnd.n1248 gnd.n1246 9.3005
R18726 gnd.n1188 gnd.n1187 9.3005
R18727 gnd.n1917 gnd.n1916 9.3005
R18728 gnd.n1918 gnd.n1186 9.3005
R18729 gnd.n1936 gnd.n1919 9.3005
R18730 gnd.n1935 gnd.n1920 9.3005
R18731 gnd.n1934 gnd.n1921 9.3005
R18732 gnd.n1932 gnd.n1922 9.3005
R18733 gnd.n1931 gnd.n1923 9.3005
R18734 gnd.n1929 gnd.n1924 9.3005
R18735 gnd.n1928 gnd.n1925 9.3005
R18736 gnd.n1136 gnd.n1135 9.3005
R18737 gnd.n2007 gnd.n2006 9.3005
R18738 gnd.n2008 gnd.n1134 9.3005
R18739 gnd.n2039 gnd.n2009 9.3005
R18740 gnd.n2038 gnd.n2010 9.3005
R18741 gnd.n2037 gnd.n2011 9.3005
R18742 gnd.n2034 gnd.n2012 9.3005
R18743 gnd.n2033 gnd.n2013 9.3005
R18744 gnd.n2030 gnd.n2014 9.3005
R18745 gnd.n2029 gnd.n2015 9.3005
R18746 gnd.n2026 gnd.n2016 9.3005
R18747 gnd.n2025 gnd.n2017 9.3005
R18748 gnd.n2024 gnd.n2018 9.3005
R18749 gnd.n2021 gnd.n2020 9.3005
R18750 gnd.n2019 gnd.n1111 9.3005
R18751 gnd.n2349 gnd.n1110 9.3005
R18752 gnd.n2351 gnd.n2350 9.3005
R18753 gnd.n1630 gnd.n1629 9.3005
R18754 gnd.n1520 gnd.n1519 9.3005
R18755 gnd.n1644 gnd.n1643 9.3005
R18756 gnd.n1645 gnd.n1518 9.3005
R18757 gnd.n1647 gnd.n1646 9.3005
R18758 gnd.n1508 gnd.n1507 9.3005
R18759 gnd.n1660 gnd.n1659 9.3005
R18760 gnd.n1661 gnd.n1506 9.3005
R18761 gnd.n1693 gnd.n1662 9.3005
R18762 gnd.n1692 gnd.n1663 9.3005
R18763 gnd.n1691 gnd.n1664 9.3005
R18764 gnd.n1690 gnd.n1665 9.3005
R18765 gnd.n1687 gnd.n1666 9.3005
R18766 gnd.n1686 gnd.n1667 9.3005
R18767 gnd.n1685 gnd.n1668 9.3005
R18768 gnd.n1683 gnd.n1669 9.3005
R18769 gnd.n1682 gnd.n1670 9.3005
R18770 gnd.n1679 gnd.n1671 9.3005
R18771 gnd.n1678 gnd.n1672 9.3005
R18772 gnd.n1677 gnd.n1673 9.3005
R18773 gnd.n1675 gnd.n1674 9.3005
R18774 gnd.n1373 gnd.n1372 9.3005
R18775 gnd.n1797 gnd.n1796 9.3005
R18776 gnd.n1798 gnd.n1371 9.3005
R18777 gnd.n1802 gnd.n1799 9.3005
R18778 gnd.n1801 gnd.n1800 9.3005
R18779 gnd.n1336 gnd.n1335 9.3005
R18780 gnd.n1845 gnd.n1844 9.3005
R18781 gnd.n1628 gnd.n1529 9.3005
R18782 gnd.n1531 gnd.n1530 9.3005
R18783 gnd.n1575 gnd.n1573 9.3005
R18784 gnd.n1576 gnd.n1572 9.3005
R18785 gnd.n1579 gnd.n1568 9.3005
R18786 gnd.n1580 gnd.n1567 9.3005
R18787 gnd.n1583 gnd.n1566 9.3005
R18788 gnd.n1584 gnd.n1565 9.3005
R18789 gnd.n1587 gnd.n1564 9.3005
R18790 gnd.n1588 gnd.n1563 9.3005
R18791 gnd.n1591 gnd.n1562 9.3005
R18792 gnd.n1592 gnd.n1561 9.3005
R18793 gnd.n1595 gnd.n1560 9.3005
R18794 gnd.n1596 gnd.n1559 9.3005
R18795 gnd.n1599 gnd.n1558 9.3005
R18796 gnd.n1600 gnd.n1557 9.3005
R18797 gnd.n1603 gnd.n1556 9.3005
R18798 gnd.n1604 gnd.n1555 9.3005
R18799 gnd.n1607 gnd.n1554 9.3005
R18800 gnd.n1608 gnd.n1553 9.3005
R18801 gnd.n1611 gnd.n1552 9.3005
R18802 gnd.n1612 gnd.n1551 9.3005
R18803 gnd.n1615 gnd.n1550 9.3005
R18804 gnd.n1617 gnd.n1549 9.3005
R18805 gnd.n1618 gnd.n1548 9.3005
R18806 gnd.n1619 gnd.n1547 9.3005
R18807 gnd.n1620 gnd.n1546 9.3005
R18808 gnd.n1627 gnd.n1626 9.3005
R18809 gnd.n1636 gnd.n1635 9.3005
R18810 gnd.n1637 gnd.n1523 9.3005
R18811 gnd.n1639 gnd.n1638 9.3005
R18812 gnd.n1514 gnd.n1513 9.3005
R18813 gnd.n1652 gnd.n1651 9.3005
R18814 gnd.n1653 gnd.n1512 9.3005
R18815 gnd.n1655 gnd.n1654 9.3005
R18816 gnd.n1501 gnd.n1500 9.3005
R18817 gnd.n1698 gnd.n1697 9.3005
R18818 gnd.n1699 gnd.n1455 9.3005
R18819 gnd.n1703 gnd.n1701 9.3005
R18820 gnd.n1702 gnd.n1434 9.3005
R18821 gnd.n1721 gnd.n1433 9.3005
R18822 gnd.n1724 gnd.n1723 9.3005
R18823 gnd.n1427 gnd.n1426 9.3005
R18824 gnd.n1735 gnd.n1733 9.3005
R18825 gnd.n1734 gnd.n1408 9.3005
R18826 gnd.n1752 gnd.n1407 9.3005
R18827 gnd.n1755 gnd.n1754 9.3005
R18828 gnd.n1402 gnd.n1397 9.3005
R18829 gnd.n1765 gnd.n1764 9.3005
R18830 gnd.n1400 gnd.n1378 9.3005
R18831 gnd.n1792 gnd.n1379 9.3005
R18832 gnd.n1791 gnd.n1790 9.3005
R18833 gnd.n1381 gnd.n1366 9.3005
R18834 gnd.n1809 gnd.n1808 9.3005
R18835 gnd.n1811 gnd.n1344 9.3005
R18836 gnd.n1840 gnd.n1345 9.3005
R18837 gnd.n1839 gnd.n1346 9.3005
R18838 gnd.n1838 gnd.n1347 9.3005
R18839 gnd.n1350 gnd.n1349 9.3005
R18840 gnd.n1237 gnd.n1233 9.3005
R18841 gnd.n1859 gnd.n1858 9.3005
R18842 gnd.n1235 gnd.n1218 9.3005
R18843 gnd.n1877 gnd.n1876 9.3005
R18844 gnd.n1879 gnd.n1214 9.3005
R18845 gnd.n1889 gnd.n1215 9.3005
R18846 gnd.n1888 gnd.n1887 9.3005
R18847 gnd.n1885 gnd.n1193 9.3005
R18848 gnd.n1912 gnd.n1194 9.3005
R18849 gnd.n1911 gnd.n1910 9.3005
R18850 gnd.n1196 gnd.n1173 9.3005
R18851 gnd.n1955 gnd.n1954 9.3005
R18852 gnd.n1956 gnd.n1166 9.3005
R18853 gnd.n1966 gnd.n1965 9.3005
R18854 gnd.n1968 gnd.n1162 9.3005
R18855 gnd.n1978 gnd.n1163 9.3005
R18856 gnd.n1977 gnd.n1976 9.3005
R18857 gnd.n1974 gnd.n1142 9.3005
R18858 gnd.n2002 gnd.n1143 9.3005
R18859 gnd.n2001 gnd.n2000 9.3005
R18860 gnd.n1145 gnd.n1121 9.3005
R18861 gnd.n2060 gnd.n2059 9.3005
R18862 gnd.n2062 gnd.n958 9.3005
R18863 gnd.n6834 gnd.n959 9.3005
R18864 gnd.n6833 gnd.n960 9.3005
R18865 gnd.n6832 gnd.n961 9.3005
R18866 gnd.n2071 gnd.n962 9.3005
R18867 gnd.n2073 gnd.n982 9.3005
R18868 gnd.n6820 gnd.n983 9.3005
R18869 gnd.n6819 gnd.n984 9.3005
R18870 gnd.n6818 gnd.n985 9.3005
R18871 gnd.n2340 gnd.n986 9.3005
R18872 gnd.n2341 gnd.n1007 9.3005
R18873 gnd.n6806 gnd.n6805 9.3005
R18874 gnd.n1525 gnd.n1524 9.3005
R18875 gnd.n784 gnd.n783 9.3005
R18876 gnd.n7010 gnd.n7009 9.3005
R18877 gnd.n7011 gnd.n782 9.3005
R18878 gnd.n7013 gnd.n7012 9.3005
R18879 gnd.n778 gnd.n777 9.3005
R18880 gnd.n7020 gnd.n7019 9.3005
R18881 gnd.n7021 gnd.n776 9.3005
R18882 gnd.n7023 gnd.n7022 9.3005
R18883 gnd.n772 gnd.n771 9.3005
R18884 gnd.n7030 gnd.n7029 9.3005
R18885 gnd.n7031 gnd.n770 9.3005
R18886 gnd.n7033 gnd.n7032 9.3005
R18887 gnd.n766 gnd.n765 9.3005
R18888 gnd.n7040 gnd.n7039 9.3005
R18889 gnd.n7041 gnd.n764 9.3005
R18890 gnd.n7043 gnd.n7042 9.3005
R18891 gnd.n760 gnd.n759 9.3005
R18892 gnd.n7050 gnd.n7049 9.3005
R18893 gnd.n7051 gnd.n758 9.3005
R18894 gnd.n7053 gnd.n7052 9.3005
R18895 gnd.n754 gnd.n753 9.3005
R18896 gnd.n7060 gnd.n7059 9.3005
R18897 gnd.n7061 gnd.n752 9.3005
R18898 gnd.n7063 gnd.n7062 9.3005
R18899 gnd.n748 gnd.n747 9.3005
R18900 gnd.n7070 gnd.n7069 9.3005
R18901 gnd.n7071 gnd.n746 9.3005
R18902 gnd.n7073 gnd.n7072 9.3005
R18903 gnd.n742 gnd.n741 9.3005
R18904 gnd.n7080 gnd.n7079 9.3005
R18905 gnd.n7081 gnd.n740 9.3005
R18906 gnd.n7083 gnd.n7082 9.3005
R18907 gnd.n736 gnd.n735 9.3005
R18908 gnd.n7090 gnd.n7089 9.3005
R18909 gnd.n7091 gnd.n734 9.3005
R18910 gnd.n7093 gnd.n7092 9.3005
R18911 gnd.n730 gnd.n729 9.3005
R18912 gnd.n7100 gnd.n7099 9.3005
R18913 gnd.n7101 gnd.n728 9.3005
R18914 gnd.n7103 gnd.n7102 9.3005
R18915 gnd.n724 gnd.n723 9.3005
R18916 gnd.n7110 gnd.n7109 9.3005
R18917 gnd.n7111 gnd.n722 9.3005
R18918 gnd.n7113 gnd.n7112 9.3005
R18919 gnd.n718 gnd.n717 9.3005
R18920 gnd.n7120 gnd.n7119 9.3005
R18921 gnd.n7121 gnd.n716 9.3005
R18922 gnd.n7123 gnd.n7122 9.3005
R18923 gnd.n712 gnd.n711 9.3005
R18924 gnd.n7130 gnd.n7129 9.3005
R18925 gnd.n7131 gnd.n710 9.3005
R18926 gnd.n7133 gnd.n7132 9.3005
R18927 gnd.n706 gnd.n705 9.3005
R18928 gnd.n7140 gnd.n7139 9.3005
R18929 gnd.n7141 gnd.n704 9.3005
R18930 gnd.n7143 gnd.n7142 9.3005
R18931 gnd.n700 gnd.n699 9.3005
R18932 gnd.n7150 gnd.n7149 9.3005
R18933 gnd.n7151 gnd.n698 9.3005
R18934 gnd.n7153 gnd.n7152 9.3005
R18935 gnd.n694 gnd.n693 9.3005
R18936 gnd.n7160 gnd.n7159 9.3005
R18937 gnd.n7161 gnd.n692 9.3005
R18938 gnd.n7163 gnd.n7162 9.3005
R18939 gnd.n688 gnd.n687 9.3005
R18940 gnd.n7170 gnd.n7169 9.3005
R18941 gnd.n7171 gnd.n686 9.3005
R18942 gnd.n7173 gnd.n7172 9.3005
R18943 gnd.n682 gnd.n681 9.3005
R18944 gnd.n7180 gnd.n7179 9.3005
R18945 gnd.n7181 gnd.n680 9.3005
R18946 gnd.n7183 gnd.n7182 9.3005
R18947 gnd.n676 gnd.n675 9.3005
R18948 gnd.n7190 gnd.n7189 9.3005
R18949 gnd.n7191 gnd.n674 9.3005
R18950 gnd.n7193 gnd.n7192 9.3005
R18951 gnd.n670 gnd.n669 9.3005
R18952 gnd.n7200 gnd.n7199 9.3005
R18953 gnd.n7201 gnd.n668 9.3005
R18954 gnd.n7203 gnd.n7202 9.3005
R18955 gnd.n664 gnd.n663 9.3005
R18956 gnd.n7210 gnd.n7209 9.3005
R18957 gnd.n7211 gnd.n662 9.3005
R18958 gnd.n7213 gnd.n7212 9.3005
R18959 gnd.n658 gnd.n657 9.3005
R18960 gnd.n7220 gnd.n7219 9.3005
R18961 gnd.n7221 gnd.n656 9.3005
R18962 gnd.n7223 gnd.n7222 9.3005
R18963 gnd.n652 gnd.n651 9.3005
R18964 gnd.n7230 gnd.n7229 9.3005
R18965 gnd.n7231 gnd.n650 9.3005
R18966 gnd.n7233 gnd.n7232 9.3005
R18967 gnd.n646 gnd.n645 9.3005
R18968 gnd.n7240 gnd.n7239 9.3005
R18969 gnd.n7241 gnd.n644 9.3005
R18970 gnd.n7243 gnd.n7242 9.3005
R18971 gnd.n640 gnd.n639 9.3005
R18972 gnd.n7250 gnd.n7249 9.3005
R18973 gnd.n7251 gnd.n638 9.3005
R18974 gnd.n7253 gnd.n7252 9.3005
R18975 gnd.n634 gnd.n633 9.3005
R18976 gnd.n7260 gnd.n7259 9.3005
R18977 gnd.n7261 gnd.n632 9.3005
R18978 gnd.n7263 gnd.n7262 9.3005
R18979 gnd.n628 gnd.n627 9.3005
R18980 gnd.n7270 gnd.n7269 9.3005
R18981 gnd.n7271 gnd.n626 9.3005
R18982 gnd.n7273 gnd.n7272 9.3005
R18983 gnd.n622 gnd.n621 9.3005
R18984 gnd.n7280 gnd.n7279 9.3005
R18985 gnd.n7281 gnd.n620 9.3005
R18986 gnd.n7283 gnd.n7282 9.3005
R18987 gnd.n616 gnd.n615 9.3005
R18988 gnd.n7290 gnd.n7289 9.3005
R18989 gnd.n7291 gnd.n614 9.3005
R18990 gnd.n7293 gnd.n7292 9.3005
R18991 gnd.n610 gnd.n609 9.3005
R18992 gnd.n7300 gnd.n7299 9.3005
R18993 gnd.n7301 gnd.n608 9.3005
R18994 gnd.n7303 gnd.n7302 9.3005
R18995 gnd.n604 gnd.n603 9.3005
R18996 gnd.n7310 gnd.n7309 9.3005
R18997 gnd.n7311 gnd.n602 9.3005
R18998 gnd.n7313 gnd.n7312 9.3005
R18999 gnd.n598 gnd.n597 9.3005
R19000 gnd.n7320 gnd.n7319 9.3005
R19001 gnd.n7321 gnd.n596 9.3005
R19002 gnd.n7323 gnd.n7322 9.3005
R19003 gnd.n592 gnd.n591 9.3005
R19004 gnd.n7330 gnd.n7329 9.3005
R19005 gnd.n7331 gnd.n590 9.3005
R19006 gnd.n7333 gnd.n7332 9.3005
R19007 gnd.n586 gnd.n585 9.3005
R19008 gnd.n7340 gnd.n7339 9.3005
R19009 gnd.n7341 gnd.n584 9.3005
R19010 gnd.n7343 gnd.n7342 9.3005
R19011 gnd.n580 gnd.n579 9.3005
R19012 gnd.n7350 gnd.n7349 9.3005
R19013 gnd.n7351 gnd.n578 9.3005
R19014 gnd.n7353 gnd.n7352 9.3005
R19015 gnd.n574 gnd.n573 9.3005
R19016 gnd.n7360 gnd.n7359 9.3005
R19017 gnd.n7361 gnd.n572 9.3005
R19018 gnd.n7363 gnd.n7362 9.3005
R19019 gnd.n568 gnd.n567 9.3005
R19020 gnd.n7370 gnd.n7369 9.3005
R19021 gnd.n7371 gnd.n566 9.3005
R19022 gnd.n7373 gnd.n7372 9.3005
R19023 gnd.n562 gnd.n561 9.3005
R19024 gnd.n7380 gnd.n7379 9.3005
R19025 gnd.n7381 gnd.n560 9.3005
R19026 gnd.n7383 gnd.n7382 9.3005
R19027 gnd.n556 gnd.n555 9.3005
R19028 gnd.n7390 gnd.n7389 9.3005
R19029 gnd.n7391 gnd.n554 9.3005
R19030 gnd.n7393 gnd.n7392 9.3005
R19031 gnd.n550 gnd.n549 9.3005
R19032 gnd.n7400 gnd.n7399 9.3005
R19033 gnd.n7401 gnd.n548 9.3005
R19034 gnd.n7403 gnd.n7402 9.3005
R19035 gnd.n544 gnd.n543 9.3005
R19036 gnd.n7410 gnd.n7409 9.3005
R19037 gnd.n7411 gnd.n542 9.3005
R19038 gnd.n7413 gnd.n7412 9.3005
R19039 gnd.n538 gnd.n537 9.3005
R19040 gnd.n7420 gnd.n7419 9.3005
R19041 gnd.n7421 gnd.n536 9.3005
R19042 gnd.n7423 gnd.n7422 9.3005
R19043 gnd.n532 gnd.n531 9.3005
R19044 gnd.n7430 gnd.n7429 9.3005
R19045 gnd.n7431 gnd.n530 9.3005
R19046 gnd.n7433 gnd.n7432 9.3005
R19047 gnd.n526 gnd.n525 9.3005
R19048 gnd.n7440 gnd.n7439 9.3005
R19049 gnd.n7441 gnd.n524 9.3005
R19050 gnd.n7443 gnd.n7442 9.3005
R19051 gnd.n520 gnd.n519 9.3005
R19052 gnd.n7450 gnd.n7449 9.3005
R19053 gnd.n7451 gnd.n518 9.3005
R19054 gnd.n7453 gnd.n7452 9.3005
R19055 gnd.n514 gnd.n513 9.3005
R19056 gnd.n7460 gnd.n7459 9.3005
R19057 gnd.n7461 gnd.n512 9.3005
R19058 gnd.n7463 gnd.n7462 9.3005
R19059 gnd.n508 gnd.n507 9.3005
R19060 gnd.n7470 gnd.n7469 9.3005
R19061 gnd.n7471 gnd.n506 9.3005
R19062 gnd.n7473 gnd.n7472 9.3005
R19063 gnd.n502 gnd.n501 9.3005
R19064 gnd.n7480 gnd.n7479 9.3005
R19065 gnd.n7481 gnd.n500 9.3005
R19066 gnd.n7484 gnd.n7483 9.3005
R19067 gnd.n7482 gnd.n496 9.3005
R19068 gnd.n7490 gnd.n495 9.3005
R19069 gnd.n7492 gnd.n7491 9.3005
R19070 gnd.n491 gnd.n490 9.3005
R19071 gnd.n7501 gnd.n7500 9.3005
R19072 gnd.n7502 gnd.n489 9.3005
R19073 gnd.n7504 gnd.n7503 9.3005
R19074 gnd.n485 gnd.n484 9.3005
R19075 gnd.n7511 gnd.n7510 9.3005
R19076 gnd.n7512 gnd.n483 9.3005
R19077 gnd.n7514 gnd.n7513 9.3005
R19078 gnd.n479 gnd.n478 9.3005
R19079 gnd.n7521 gnd.n7520 9.3005
R19080 gnd.n7522 gnd.n477 9.3005
R19081 gnd.n7524 gnd.n7523 9.3005
R19082 gnd.n473 gnd.n472 9.3005
R19083 gnd.n7531 gnd.n7530 9.3005
R19084 gnd.n7532 gnd.n471 9.3005
R19085 gnd.n7534 gnd.n7533 9.3005
R19086 gnd.n467 gnd.n466 9.3005
R19087 gnd.n7541 gnd.n7540 9.3005
R19088 gnd.n7542 gnd.n465 9.3005
R19089 gnd.n7544 gnd.n7543 9.3005
R19090 gnd.n461 gnd.n460 9.3005
R19091 gnd.n7551 gnd.n7550 9.3005
R19092 gnd.n7552 gnd.n459 9.3005
R19093 gnd.n7554 gnd.n7553 9.3005
R19094 gnd.n455 gnd.n454 9.3005
R19095 gnd.n7561 gnd.n7560 9.3005
R19096 gnd.n7562 gnd.n453 9.3005
R19097 gnd.n7564 gnd.n7563 9.3005
R19098 gnd.n449 gnd.n448 9.3005
R19099 gnd.n7571 gnd.n7570 9.3005
R19100 gnd.n7572 gnd.n447 9.3005
R19101 gnd.n7574 gnd.n7573 9.3005
R19102 gnd.n443 gnd.n442 9.3005
R19103 gnd.n7581 gnd.n7580 9.3005
R19104 gnd.n7582 gnd.n441 9.3005
R19105 gnd.n7584 gnd.n7583 9.3005
R19106 gnd.n437 gnd.n436 9.3005
R19107 gnd.n7591 gnd.n7590 9.3005
R19108 gnd.n7592 gnd.n435 9.3005
R19109 gnd.n7594 gnd.n7593 9.3005
R19110 gnd.n431 gnd.n430 9.3005
R19111 gnd.n7601 gnd.n7600 9.3005
R19112 gnd.n7602 gnd.n429 9.3005
R19113 gnd.n7604 gnd.n7603 9.3005
R19114 gnd.n425 gnd.n424 9.3005
R19115 gnd.n7611 gnd.n7610 9.3005
R19116 gnd.n7612 gnd.n423 9.3005
R19117 gnd.n7614 gnd.n7613 9.3005
R19118 gnd.n419 gnd.n418 9.3005
R19119 gnd.n7621 gnd.n7620 9.3005
R19120 gnd.n7622 gnd.n417 9.3005
R19121 gnd.n7624 gnd.n7623 9.3005
R19122 gnd.n413 gnd.n412 9.3005
R19123 gnd.n7631 gnd.n7630 9.3005
R19124 gnd.n7632 gnd.n411 9.3005
R19125 gnd.n7634 gnd.n7633 9.3005
R19126 gnd.n407 gnd.n406 9.3005
R19127 gnd.n7641 gnd.n7640 9.3005
R19128 gnd.n7642 gnd.n405 9.3005
R19129 gnd.n7644 gnd.n7643 9.3005
R19130 gnd.n401 gnd.n400 9.3005
R19131 gnd.n7651 gnd.n7650 9.3005
R19132 gnd.n7652 gnd.n399 9.3005
R19133 gnd.n7654 gnd.n7653 9.3005
R19134 gnd.n395 gnd.n394 9.3005
R19135 gnd.n7661 gnd.n7660 9.3005
R19136 gnd.n7662 gnd.n393 9.3005
R19137 gnd.n7664 gnd.n7663 9.3005
R19138 gnd.n389 gnd.n388 9.3005
R19139 gnd.n7671 gnd.n7670 9.3005
R19140 gnd.n7672 gnd.n387 9.3005
R19141 gnd.n7674 gnd.n7673 9.3005
R19142 gnd.n383 gnd.n382 9.3005
R19143 gnd.n7681 gnd.n7680 9.3005
R19144 gnd.n7682 gnd.n381 9.3005
R19145 gnd.n7684 gnd.n7683 9.3005
R19146 gnd.n377 gnd.n376 9.3005
R19147 gnd.n7691 gnd.n7690 9.3005
R19148 gnd.n7692 gnd.n375 9.3005
R19149 gnd.n7694 gnd.n7693 9.3005
R19150 gnd.n371 gnd.n370 9.3005
R19151 gnd.n7702 gnd.n7701 9.3005
R19152 gnd.n7703 gnd.n369 9.3005
R19153 gnd.n7706 gnd.n7705 9.3005
R19154 gnd.n7494 gnd.n7493 9.3005
R19155 gnd.n8071 gnd.n8070 9.3005
R19156 gnd.n8069 gnd.n97 9.3005
R19157 gnd.n5828 gnd.n99 9.3005
R19158 gnd.n5832 gnd.n5831 9.3005
R19159 gnd.n5833 gnd.n5827 9.3005
R19160 gnd.n5888 gnd.n5834 9.3005
R19161 gnd.n5887 gnd.n5835 9.3005
R19162 gnd.n5886 gnd.n5836 9.3005
R19163 gnd.n5863 gnd.n5837 9.3005
R19164 gnd.n5876 gnd.n5864 9.3005
R19165 gnd.n5875 gnd.n5865 9.3005
R19166 gnd.n5874 gnd.n5866 9.3005
R19167 gnd.n359 gnd.n358 9.3005
R19168 gnd.n7719 gnd.n7718 9.3005
R19169 gnd.n7720 gnd.n357 9.3005
R19170 gnd.n7819 gnd.n7721 9.3005
R19171 gnd.n7818 gnd.n7722 9.3005
R19172 gnd.n7817 gnd.n7723 9.3005
R19173 gnd.n7815 gnd.n7724 9.3005
R19174 gnd.n7814 gnd.n7725 9.3005
R19175 gnd.n7812 gnd.n7726 9.3005
R19176 gnd.n7811 gnd.n7727 9.3005
R19177 gnd.n7809 gnd.n7728 9.3005
R19178 gnd.n7808 gnd.n7729 9.3005
R19179 gnd.n7806 gnd.n7730 9.3005
R19180 gnd.n7805 gnd.n7731 9.3005
R19181 gnd.n7803 gnd.n7732 9.3005
R19182 gnd.n7802 gnd.n7733 9.3005
R19183 gnd.n7800 gnd.n7734 9.3005
R19184 gnd.n7799 gnd.n7735 9.3005
R19185 gnd.n7797 gnd.n7736 9.3005
R19186 gnd.n7796 gnd.n7737 9.3005
R19187 gnd.n7751 gnd.n7750 9.3005
R19188 gnd.n7753 gnd.n7752 9.3005
R19189 gnd.n7756 gnd.n7747 9.3005
R19190 gnd.n7760 gnd.n7759 9.3005
R19191 gnd.n7761 gnd.n7746 9.3005
R19192 gnd.n7763 gnd.n7762 9.3005
R19193 gnd.n7766 gnd.n7745 9.3005
R19194 gnd.n7770 gnd.n7769 9.3005
R19195 gnd.n7771 gnd.n7744 9.3005
R19196 gnd.n7773 gnd.n7772 9.3005
R19197 gnd.n7776 gnd.n7743 9.3005
R19198 gnd.n7780 gnd.n7779 9.3005
R19199 gnd.n7781 gnd.n7742 9.3005
R19200 gnd.n7783 gnd.n7782 9.3005
R19201 gnd.n7786 gnd.n7741 9.3005
R19202 gnd.n7790 gnd.n7789 9.3005
R19203 gnd.n7791 gnd.n7740 9.3005
R19204 gnd.n7793 gnd.n7792 9.3005
R19205 gnd.n7748 gnd.n354 9.3005
R19206 gnd.n254 gnd.n253 9.3005
R19207 gnd.n7970 gnd.n296 9.3005
R19208 gnd.n7969 gnd.n297 9.3005
R19209 gnd.n7968 gnd.n298 9.3005
R19210 gnd.n7965 gnd.n299 9.3005
R19211 gnd.n7964 gnd.n300 9.3005
R19212 gnd.n7961 gnd.n301 9.3005
R19213 gnd.n7960 gnd.n302 9.3005
R19214 gnd.n7957 gnd.n303 9.3005
R19215 gnd.n7956 gnd.n304 9.3005
R19216 gnd.n7953 gnd.n305 9.3005
R19217 gnd.n7952 gnd.n306 9.3005
R19218 gnd.n7949 gnd.n307 9.3005
R19219 gnd.n7948 gnd.n308 9.3005
R19220 gnd.n7945 gnd.n309 9.3005
R19221 gnd.n7944 gnd.n310 9.3005
R19222 gnd.n7941 gnd.n311 9.3005
R19223 gnd.n7937 gnd.n312 9.3005
R19224 gnd.n7934 gnd.n313 9.3005
R19225 gnd.n7933 gnd.n314 9.3005
R19226 gnd.n7930 gnd.n315 9.3005
R19227 gnd.n7929 gnd.n316 9.3005
R19228 gnd.n7926 gnd.n317 9.3005
R19229 gnd.n7925 gnd.n318 9.3005
R19230 gnd.n7922 gnd.n319 9.3005
R19231 gnd.n7921 gnd.n320 9.3005
R19232 gnd.n7918 gnd.n321 9.3005
R19233 gnd.n7917 gnd.n322 9.3005
R19234 gnd.n7914 gnd.n323 9.3005
R19235 gnd.n7913 gnd.n324 9.3005
R19236 gnd.n7910 gnd.n325 9.3005
R19237 gnd.n7909 gnd.n326 9.3005
R19238 gnd.n7906 gnd.n327 9.3005
R19239 gnd.n7905 gnd.n328 9.3005
R19240 gnd.n7902 gnd.n329 9.3005
R19241 gnd.n7901 gnd.n330 9.3005
R19242 gnd.n7898 gnd.n7897 9.3005
R19243 gnd.n7896 gnd.n331 9.3005
R19244 gnd.n7895 gnd.n7894 9.3005
R19245 gnd.n7891 gnd.n334 9.3005
R19246 gnd.n7888 gnd.n335 9.3005
R19247 gnd.n7887 gnd.n336 9.3005
R19248 gnd.n7884 gnd.n337 9.3005
R19249 gnd.n7883 gnd.n338 9.3005
R19250 gnd.n7880 gnd.n339 9.3005
R19251 gnd.n7879 gnd.n340 9.3005
R19252 gnd.n7876 gnd.n341 9.3005
R19253 gnd.n7875 gnd.n342 9.3005
R19254 gnd.n7872 gnd.n343 9.3005
R19255 gnd.n7871 gnd.n344 9.3005
R19256 gnd.n7868 gnd.n345 9.3005
R19257 gnd.n7867 gnd.n346 9.3005
R19258 gnd.n7864 gnd.n347 9.3005
R19259 gnd.n7863 gnd.n348 9.3005
R19260 gnd.n7860 gnd.n349 9.3005
R19261 gnd.n7859 gnd.n350 9.3005
R19262 gnd.n7856 gnd.n7855 9.3005
R19263 gnd.n7854 gnd.n351 9.3005
R19264 gnd.n7976 gnd.n7975 9.3005
R19265 gnd.n6010 gnd.n6009 9.3005
R19266 gnd.n3192 gnd.n3191 9.3005
R19267 gnd.n3216 gnd.n3215 9.3005
R19268 gnd.n5997 gnd.n3217 9.3005
R19269 gnd.n5996 gnd.n3218 9.3005
R19270 gnd.n5995 gnd.n3219 9.3005
R19271 gnd.n5705 gnd.n3220 9.3005
R19272 gnd.n5985 gnd.n3238 9.3005
R19273 gnd.n5984 gnd.n3239 9.3005
R19274 gnd.n5983 gnd.n3240 9.3005
R19275 gnd.n5720 gnd.n3241 9.3005
R19276 gnd.n5973 gnd.n3258 9.3005
R19277 gnd.n5972 gnd.n3259 9.3005
R19278 gnd.n5971 gnd.n3260 9.3005
R19279 gnd.n5735 gnd.n3261 9.3005
R19280 gnd.n5961 gnd.n3279 9.3005
R19281 gnd.n5960 gnd.n3280 9.3005
R19282 gnd.n5959 gnd.n3281 9.3005
R19283 gnd.n5750 gnd.n3282 9.3005
R19284 gnd.n5949 gnd.n3299 9.3005
R19285 gnd.n5948 gnd.n3300 9.3005
R19286 gnd.n5947 gnd.n3301 9.3005
R19287 gnd.n5765 gnd.n3302 9.3005
R19288 gnd.n5937 gnd.n3321 9.3005
R19289 gnd.n5936 gnd.n3322 9.3005
R19290 gnd.n5935 gnd.n3323 9.3005
R19291 gnd.n3365 gnd.n3324 9.3005
R19292 gnd.n5797 gnd.n5796 9.3005
R19293 gnd.n5801 gnd.n5800 9.3005
R19294 gnd.n5802 gnd.n3355 9.3005
R19295 gnd.n5912 gnd.n3356 9.3005
R19296 gnd.n5911 gnd.n3357 9.3005
R19297 gnd.n5910 gnd.n3358 9.3005
R19298 gnd.n5806 gnd.n3359 9.3005
R19299 gnd.n5900 gnd.n5807 9.3005
R19300 gnd.n5808 gnd.n124 9.3005
R19301 gnd.n8057 gnd.n125 9.3005
R19302 gnd.n8056 gnd.n126 9.3005
R19303 gnd.n8055 gnd.n127 9.3005
R19304 gnd.n5841 gnd.n128 9.3005
R19305 gnd.n8045 gnd.n143 9.3005
R19306 gnd.n8044 gnd.n144 9.3005
R19307 gnd.n8043 gnd.n145 9.3005
R19308 gnd.n5867 gnd.n146 9.3005
R19309 gnd.n8033 gnd.n164 9.3005
R19310 gnd.n8032 gnd.n165 9.3005
R19311 gnd.n8031 gnd.n166 9.3005
R19312 gnd.n356 gnd.n167 9.3005
R19313 gnd.n8021 gnd.n183 9.3005
R19314 gnd.n8020 gnd.n184 9.3005
R19315 gnd.n8019 gnd.n185 9.3005
R19316 gnd.n7828 gnd.n186 9.3005
R19317 gnd.n8009 gnd.n204 9.3005
R19318 gnd.n8008 gnd.n205 9.3005
R19319 gnd.n8007 gnd.n206 9.3005
R19320 gnd.n7835 gnd.n207 9.3005
R19321 gnd.n7997 gnd.n222 9.3005
R19322 gnd.n7996 gnd.n223 9.3005
R19323 gnd.n7995 gnd.n224 9.3005
R19324 gnd.n7842 gnd.n225 9.3005
R19325 gnd.n7985 gnd.n242 9.3005
R19326 gnd.n7984 gnd.n243 9.3005
R19327 gnd.n7983 gnd.n244 9.3005
R19328 gnd.n7852 gnd.n245 9.3005
R19329 gnd.n6011 gnd.n3190 9.3005
R19330 gnd.n6009 gnd.n6008 9.3005
R19331 gnd.n6007 gnd.n3192 9.3005
R19332 gnd.n3216 gnd.n3193 9.3005
R19333 gnd.n3389 gnd.n3217 9.3005
R19334 gnd.n5703 gnd.n3218 9.3005
R19335 gnd.n5704 gnd.n3219 9.3005
R19336 gnd.n5706 gnd.n5705 9.3005
R19337 gnd.n3385 gnd.n3238 9.3005
R19338 gnd.n5718 gnd.n3239 9.3005
R19339 gnd.n5719 gnd.n3240 9.3005
R19340 gnd.n5721 gnd.n5720 9.3005
R19341 gnd.n3380 gnd.n3258 9.3005
R19342 gnd.n5733 gnd.n3259 9.3005
R19343 gnd.n5734 gnd.n3260 9.3005
R19344 gnd.n5736 gnd.n5735 9.3005
R19345 gnd.n3376 gnd.n3279 9.3005
R19346 gnd.n5748 gnd.n3280 9.3005
R19347 gnd.n5749 gnd.n3281 9.3005
R19348 gnd.n5751 gnd.n5750 9.3005
R19349 gnd.n3371 gnd.n3299 9.3005
R19350 gnd.n5763 gnd.n3300 9.3005
R19351 gnd.n5764 gnd.n3301 9.3005
R19352 gnd.n5766 gnd.n5765 9.3005
R19353 gnd.n3366 gnd.n3321 9.3005
R19354 gnd.n5790 gnd.n3322 9.3005
R19355 gnd.n5791 gnd.n3323 9.3005
R19356 gnd.n5792 gnd.n3365 9.3005
R19357 gnd.n5796 gnd.n5795 9.3005
R19358 gnd.n5801 gnd.n3364 9.3005
R19359 gnd.n5803 gnd.n5802 9.3005
R19360 gnd.n5804 gnd.n3356 9.3005
R19361 gnd.n5805 gnd.n3357 9.3005
R19362 gnd.n5906 gnd.n3358 9.3005
R19363 gnd.n5905 gnd.n5806 9.3005
R19364 gnd.n5904 gnd.n5807 9.3005
R19365 gnd.n5809 gnd.n5808 9.3005
R19366 gnd.n5838 gnd.n125 9.3005
R19367 gnd.n5839 gnd.n126 9.3005
R19368 gnd.n5840 gnd.n127 9.3005
R19369 gnd.n5882 gnd.n5841 9.3005
R19370 gnd.n5881 gnd.n143 9.3005
R19371 gnd.n5880 gnd.n144 9.3005
R19372 gnd.n5842 gnd.n145 9.3005
R19373 gnd.n5870 gnd.n5867 9.3005
R19374 gnd.n5869 gnd.n164 9.3005
R19375 gnd.n5868 gnd.n165 9.3005
R19376 gnd.n355 gnd.n166 9.3005
R19377 gnd.n7823 gnd.n356 9.3005
R19378 gnd.n7824 gnd.n183 9.3005
R19379 gnd.n7826 gnd.n184 9.3005
R19380 gnd.n7827 gnd.n185 9.3005
R19381 gnd.n7830 gnd.n7828 9.3005
R19382 gnd.n7831 gnd.n204 9.3005
R19383 gnd.n7833 gnd.n205 9.3005
R19384 gnd.n7834 gnd.n206 9.3005
R19385 gnd.n7837 gnd.n7835 9.3005
R19386 gnd.n7838 gnd.n222 9.3005
R19387 gnd.n7840 gnd.n223 9.3005
R19388 gnd.n7841 gnd.n224 9.3005
R19389 gnd.n7844 gnd.n7842 9.3005
R19390 gnd.n7845 gnd.n242 9.3005
R19391 gnd.n7847 gnd.n243 9.3005
R19392 gnd.n7848 gnd.n244 9.3005
R19393 gnd.n7852 gnd.n7851 9.3005
R19394 gnd.n3190 gnd.n3184 9.3005
R19395 gnd.n6021 gnd.n6020 9.3005
R19396 gnd.n6024 gnd.n3182 9.3005
R19397 gnd.n6025 gnd.n3181 9.3005
R19398 gnd.n6028 gnd.n3180 9.3005
R19399 gnd.n6029 gnd.n3179 9.3005
R19400 gnd.n6032 gnd.n3178 9.3005
R19401 gnd.n6033 gnd.n3177 9.3005
R19402 gnd.n6036 gnd.n3176 9.3005
R19403 gnd.n6037 gnd.n3175 9.3005
R19404 gnd.n6040 gnd.n3174 9.3005
R19405 gnd.n6041 gnd.n3173 9.3005
R19406 gnd.n6044 gnd.n3172 9.3005
R19407 gnd.n6045 gnd.n3171 9.3005
R19408 gnd.n6048 gnd.n3170 9.3005
R19409 gnd.n6049 gnd.n3169 9.3005
R19410 gnd.n6052 gnd.n3168 9.3005
R19411 gnd.n6053 gnd.n3167 9.3005
R19412 gnd.n6056 gnd.n3166 9.3005
R19413 gnd.n6057 gnd.n3165 9.3005
R19414 gnd.n6060 gnd.n3164 9.3005
R19415 gnd.n6064 gnd.n3160 9.3005
R19416 gnd.n6065 gnd.n3159 9.3005
R19417 gnd.n6068 gnd.n3158 9.3005
R19418 gnd.n6069 gnd.n3157 9.3005
R19419 gnd.n6072 gnd.n3156 9.3005
R19420 gnd.n6073 gnd.n3155 9.3005
R19421 gnd.n6076 gnd.n3154 9.3005
R19422 gnd.n6077 gnd.n3153 9.3005
R19423 gnd.n6080 gnd.n3152 9.3005
R19424 gnd.n6082 gnd.n3148 9.3005
R19425 gnd.n6085 gnd.n3147 9.3005
R19426 gnd.n6086 gnd.n3146 9.3005
R19427 gnd.n6089 gnd.n3145 9.3005
R19428 gnd.n6090 gnd.n3144 9.3005
R19429 gnd.n6093 gnd.n3143 9.3005
R19430 gnd.n6094 gnd.n3142 9.3005
R19431 gnd.n6097 gnd.n3141 9.3005
R19432 gnd.n6099 gnd.n3138 9.3005
R19433 gnd.n6102 gnd.n3137 9.3005
R19434 gnd.n6103 gnd.n3136 9.3005
R19435 gnd.n6106 gnd.n3135 9.3005
R19436 gnd.n6107 gnd.n3134 9.3005
R19437 gnd.n6110 gnd.n3133 9.3005
R19438 gnd.n6111 gnd.n3132 9.3005
R19439 gnd.n6114 gnd.n3131 9.3005
R19440 gnd.n6115 gnd.n3130 9.3005
R19441 gnd.n6118 gnd.n3129 9.3005
R19442 gnd.n6119 gnd.n3128 9.3005
R19443 gnd.n6122 gnd.n3127 9.3005
R19444 gnd.n6123 gnd.n3126 9.3005
R19445 gnd.n6126 gnd.n3125 9.3005
R19446 gnd.n6128 gnd.n3124 9.3005
R19447 gnd.n6129 gnd.n3123 9.3005
R19448 gnd.n6130 gnd.n3122 9.3005
R19449 gnd.n6131 gnd.n3121 9.3005
R19450 gnd.n6061 gnd.n3161 9.3005
R19451 gnd.n6019 gnd.n6016 9.3005
R19452 gnd.n3203 gnd.n3200 9.3005
R19453 gnd.n6003 gnd.n3204 9.3005
R19454 gnd.n6002 gnd.n3205 9.3005
R19455 gnd.n6001 gnd.n3206 9.3005
R19456 gnd.n3227 gnd.n3207 9.3005
R19457 gnd.n5991 gnd.n3228 9.3005
R19458 gnd.n5990 gnd.n3229 9.3005
R19459 gnd.n5989 gnd.n3230 9.3005
R19460 gnd.n3248 gnd.n3231 9.3005
R19461 gnd.n5979 gnd.n3249 9.3005
R19462 gnd.n5978 gnd.n3250 9.3005
R19463 gnd.n5977 gnd.n3251 9.3005
R19464 gnd.n3268 gnd.n3252 9.3005
R19465 gnd.n5967 gnd.n3269 9.3005
R19466 gnd.n5966 gnd.n3270 9.3005
R19467 gnd.n5965 gnd.n3271 9.3005
R19468 gnd.n3289 gnd.n3272 9.3005
R19469 gnd.n5955 gnd.n3290 9.3005
R19470 gnd.n5954 gnd.n3291 9.3005
R19471 gnd.n5953 gnd.n3292 9.3005
R19472 gnd.n3309 gnd.n3293 9.3005
R19473 gnd.n5943 gnd.n3310 9.3005
R19474 gnd.n5942 gnd.n3311 9.3005
R19475 gnd.n5941 gnd.n3312 9.3005
R19476 gnd.n3314 gnd.n3313 9.3005
R19477 gnd.n5931 gnd.n110 9.3005
R19478 gnd.n115 gnd.n109 9.3005
R19479 gnd.n8051 gnd.n134 9.3005
R19480 gnd.n8050 gnd.n135 9.3005
R19481 gnd.n8049 gnd.n136 9.3005
R19482 gnd.n153 gnd.n137 9.3005
R19483 gnd.n8039 gnd.n154 9.3005
R19484 gnd.n8038 gnd.n155 9.3005
R19485 gnd.n8037 gnd.n156 9.3005
R19486 gnd.n173 gnd.n157 9.3005
R19487 gnd.n8027 gnd.n174 9.3005
R19488 gnd.n8026 gnd.n175 9.3005
R19489 gnd.n8025 gnd.n176 9.3005
R19490 gnd.n193 gnd.n177 9.3005
R19491 gnd.n8015 gnd.n194 9.3005
R19492 gnd.n8014 gnd.n195 9.3005
R19493 gnd.n8013 gnd.n196 9.3005
R19494 gnd.n213 gnd.n197 9.3005
R19495 gnd.n8003 gnd.n214 9.3005
R19496 gnd.n8002 gnd.n215 9.3005
R19497 gnd.n8001 gnd.n216 9.3005
R19498 gnd.n232 gnd.n217 9.3005
R19499 gnd.n7991 gnd.n233 9.3005
R19500 gnd.n7990 gnd.n234 9.3005
R19501 gnd.n7989 gnd.n235 9.3005
R19502 gnd.n251 gnd.n236 9.3005
R19503 gnd.n7979 gnd.n252 9.3005
R19504 gnd.n7978 gnd.n7977 9.3005
R19505 gnd.n3202 gnd.n3201 9.3005
R19506 gnd.n8062 gnd.n8061 9.3005
R19507 gnd.n4351 gnd.n4350 9.3005
R19508 gnd.n4373 gnd.n4352 9.3005
R19509 gnd.n4372 gnd.n4353 9.3005
R19510 gnd.n4371 gnd.n4354 9.3005
R19511 gnd.n4357 gnd.n4355 9.3005
R19512 gnd.n4367 gnd.n4358 9.3005
R19513 gnd.n4366 gnd.n4359 9.3005
R19514 gnd.n4365 gnd.n4360 9.3005
R19515 gnd.n4363 gnd.n4362 9.3005
R19516 gnd.n4361 gnd.n3990 9.3005
R19517 gnd.n3988 gnd.n3987 9.3005
R19518 gnd.n4439 gnd.n4438 9.3005
R19519 gnd.n4440 gnd.n3986 9.3005
R19520 gnd.n4442 gnd.n4441 9.3005
R19521 gnd.n3984 gnd.n3983 9.3005
R19522 gnd.n4447 gnd.n4446 9.3005
R19523 gnd.n4448 gnd.n3982 9.3005
R19524 gnd.n4454 gnd.n4449 9.3005
R19525 gnd.n4453 gnd.n4450 9.3005
R19526 gnd.n4452 gnd.n4451 9.3005
R19527 gnd.n3966 gnd.n3965 9.3005
R19528 gnd.n4742 gnd.n4741 9.3005
R19529 gnd.n4743 gnd.n3964 9.3005
R19530 gnd.n4745 gnd.n4744 9.3005
R19531 gnd.n3962 gnd.n3961 9.3005
R19532 gnd.n4750 gnd.n4749 9.3005
R19533 gnd.n4751 gnd.n3960 9.3005
R19534 gnd.n4761 gnd.n4752 9.3005
R19535 gnd.n4760 gnd.n4753 9.3005
R19536 gnd.n4759 gnd.n4754 9.3005
R19537 gnd.n4756 gnd.n4755 9.3005
R19538 gnd.n3932 gnd.n3931 9.3005
R19539 gnd.n4778 gnd.n4777 9.3005
R19540 gnd.n4779 gnd.n3930 9.3005
R19541 gnd.n4781 gnd.n4780 9.3005
R19542 gnd.n3916 gnd.n3915 9.3005
R19543 gnd.n4811 gnd.n4810 9.3005
R19544 gnd.n4812 gnd.n3914 9.3005
R19545 gnd.n4823 gnd.n4813 9.3005
R19546 gnd.n4822 gnd.n4814 9.3005
R19547 gnd.n4821 gnd.n4815 9.3005
R19548 gnd.n4818 gnd.n4817 9.3005
R19549 gnd.n4816 gnd.n2905 9.3005
R19550 gnd.n6316 gnd.n2906 9.3005
R19551 gnd.n6315 gnd.n2907 9.3005
R19552 gnd.n6314 gnd.n2908 9.3005
R19553 gnd.n5007 gnd.n2909 9.3005
R19554 gnd.n5008 gnd.n5006 9.3005
R19555 gnd.n5010 gnd.n5009 9.3005
R19556 gnd.n3805 gnd.n3804 9.3005
R19557 gnd.n5036 gnd.n5035 9.3005
R19558 gnd.n5037 gnd.n3803 9.3005
R19559 gnd.n5050 gnd.n5038 9.3005
R19560 gnd.n5049 gnd.n5039 9.3005
R19561 gnd.n5048 gnd.n5040 9.3005
R19562 gnd.n5042 gnd.n5041 9.3005
R19563 gnd.n5044 gnd.n5043 9.3005
R19564 gnd.n3767 gnd.n3766 9.3005
R19565 gnd.n5094 gnd.n5093 9.3005
R19566 gnd.n5095 gnd.n3765 9.3005
R19567 gnd.n5097 gnd.n5096 9.3005
R19568 gnd.n3749 gnd.n3748 9.3005
R19569 gnd.n5120 gnd.n5119 9.3005
R19570 gnd.n5121 gnd.n3747 9.3005
R19571 gnd.n5125 gnd.n5122 9.3005
R19572 gnd.n5124 gnd.n5123 9.3005
R19573 gnd.n3725 gnd.n3724 9.3005
R19574 gnd.n5159 gnd.n5158 9.3005
R19575 gnd.n5160 gnd.n3723 9.3005
R19576 gnd.n5173 gnd.n5161 9.3005
R19577 gnd.n5172 gnd.n5162 9.3005
R19578 gnd.n5171 gnd.n5163 9.3005
R19579 gnd.n5165 gnd.n5164 9.3005
R19580 gnd.n5167 gnd.n5166 9.3005
R19581 gnd.n3686 gnd.n3685 9.3005
R19582 gnd.n5217 gnd.n5216 9.3005
R19583 gnd.n5218 gnd.n3684 9.3005
R19584 gnd.n5220 gnd.n5219 9.3005
R19585 gnd.n3667 gnd.n3666 9.3005
R19586 gnd.n5242 gnd.n5241 9.3005
R19587 gnd.n5243 gnd.n3665 9.3005
R19588 gnd.n5247 gnd.n5244 9.3005
R19589 gnd.n5246 gnd.n5245 9.3005
R19590 gnd.n3642 gnd.n3641 9.3005
R19591 gnd.n5280 gnd.n5279 9.3005
R19592 gnd.n5281 gnd.n3640 9.3005
R19593 gnd.n5291 gnd.n5282 9.3005
R19594 gnd.n5290 gnd.n5283 9.3005
R19595 gnd.n5289 gnd.n5284 9.3005
R19596 gnd.n5286 gnd.n5285 9.3005
R19597 gnd.n3608 gnd.n3607 9.3005
R19598 gnd.n5326 gnd.n5325 9.3005
R19599 gnd.n5327 gnd.n3606 9.3005
R19600 gnd.n5331 gnd.n5328 9.3005
R19601 gnd.n5330 gnd.n5329 9.3005
R19602 gnd.n3580 gnd.n3579 9.3005
R19603 gnd.n5361 gnd.n5360 9.3005
R19604 gnd.n5362 gnd.n3578 9.3005
R19605 gnd.n5364 gnd.n5363 9.3005
R19606 gnd.n3551 gnd.n3550 9.3005
R19607 gnd.n5398 gnd.n5397 9.3005
R19608 gnd.n5399 gnd.n3549 9.3005
R19609 gnd.n5403 gnd.n5400 9.3005
R19610 gnd.n5402 gnd.n5401 9.3005
R19611 gnd.n3451 gnd.n3450 9.3005
R19612 gnd.n5548 gnd.n5547 9.3005
R19613 gnd.n5549 gnd.n3449 9.3005
R19614 gnd.n5551 gnd.n5550 9.3005
R19615 gnd.n3438 gnd.n3437 9.3005
R19616 gnd.n5564 gnd.n5563 9.3005
R19617 gnd.n5565 gnd.n3436 9.3005
R19618 gnd.n5570 gnd.n5566 9.3005
R19619 gnd.n5569 gnd.n5568 9.3005
R19620 gnd.n5567 gnd.n3425 9.3005
R19621 gnd.n5583 gnd.n3424 9.3005
R19622 gnd.n5585 gnd.n5584 9.3005
R19623 gnd.n5586 gnd.n3423 9.3005
R19624 gnd.n5680 gnd.n5587 9.3005
R19625 gnd.n5679 gnd.n5588 9.3005
R19626 gnd.n5678 gnd.n5589 9.3005
R19627 gnd.n5592 gnd.n5590 9.3005
R19628 gnd.n5674 gnd.n5593 9.3005
R19629 gnd.n5673 gnd.n5594 9.3005
R19630 gnd.n5672 gnd.n5595 9.3005
R19631 gnd.n5598 gnd.n5596 9.3005
R19632 gnd.n5666 gnd.n5599 9.3005
R19633 gnd.n5665 gnd.n5600 9.3005
R19634 gnd.n5664 gnd.n5601 9.3005
R19635 gnd.n5604 gnd.n5602 9.3005
R19636 gnd.n5660 gnd.n5605 9.3005
R19637 gnd.n5659 gnd.n5606 9.3005
R19638 gnd.n5658 gnd.n5607 9.3005
R19639 gnd.n5610 gnd.n5608 9.3005
R19640 gnd.n5654 gnd.n5611 9.3005
R19641 gnd.n5653 gnd.n5612 9.3005
R19642 gnd.n5652 gnd.n5613 9.3005
R19643 gnd.n5616 gnd.n5614 9.3005
R19644 gnd.n5648 gnd.n5617 9.3005
R19645 gnd.n5647 gnd.n5618 9.3005
R19646 gnd.n5646 gnd.n5619 9.3005
R19647 gnd.n5622 gnd.n5620 9.3005
R19648 gnd.n5642 gnd.n5623 9.3005
R19649 gnd.n5641 gnd.n5624 9.3005
R19650 gnd.n5640 gnd.n5625 9.3005
R19651 gnd.n5628 gnd.n5626 9.3005
R19652 gnd.n5636 gnd.n5629 9.3005
R19653 gnd.n5635 gnd.n5630 9.3005
R19654 gnd.n5634 gnd.n5632 9.3005
R19655 gnd.n5631 gnd.n3336 9.3005
R19656 gnd.n5894 gnd.n5823 9.3005
R19657 gnd.n5846 gnd.n5824 9.3005
R19658 gnd.n5848 gnd.n5847 9.3005
R19659 gnd.n5849 gnd.n5845 9.3005
R19660 gnd.n5860 gnd.n5850 9.3005
R19661 gnd.n5859 gnd.n5851 9.3005
R19662 gnd.n5858 gnd.n5852 9.3005
R19663 gnd.n5855 gnd.n5854 9.3005
R19664 gnd.n5853 gnd.n363 9.3005
R19665 gnd.n7713 gnd.n364 9.3005
R19666 gnd.n7712 gnd.n365 9.3005
R19667 gnd.n7711 gnd.n366 9.3005
R19668 gnd.n7704 gnd.n367 9.3005
R19669 gnd.n4313 gnd.n4312 9.3005
R19670 gnd.n4166 gnd.n4104 9.3005
R19671 gnd.n4169 gnd.n4168 9.3005
R19672 gnd.n4170 gnd.n4103 9.3005
R19673 gnd.n4173 gnd.n4171 9.3005
R19674 gnd.n4174 gnd.n4102 9.3005
R19675 gnd.n4177 gnd.n4176 9.3005
R19676 gnd.n4178 gnd.n4101 9.3005
R19677 gnd.n4181 gnd.n4179 9.3005
R19678 gnd.n4182 gnd.n4100 9.3005
R19679 gnd.n4185 gnd.n4184 9.3005
R19680 gnd.n4186 gnd.n4099 9.3005
R19681 gnd.n4189 gnd.n4187 9.3005
R19682 gnd.n4190 gnd.n4098 9.3005
R19683 gnd.n4193 gnd.n4192 9.3005
R19684 gnd.n4194 gnd.n4097 9.3005
R19685 gnd.n4197 gnd.n4196 9.3005
R19686 gnd.n4195 gnd.n4069 9.3005
R19687 gnd.n4215 gnd.n4070 9.3005
R19688 gnd.n4214 gnd.n4071 9.3005
R19689 gnd.n4213 gnd.n4072 9.3005
R19690 gnd.n4062 gnd.n4061 9.3005
R19691 gnd.n4251 gnd.n4250 9.3005
R19692 gnd.n4252 gnd.n4060 9.3005
R19693 gnd.n4255 gnd.n4254 9.3005
R19694 gnd.n4253 gnd.n4055 9.3005
R19695 gnd.n4279 gnd.n4056 9.3005
R19696 gnd.n4278 gnd.n4057 9.3005
R19697 gnd.n4277 gnd.n4058 9.3005
R19698 gnd.n4044 gnd.n4043 9.3005
R19699 gnd.n4310 gnd.n4309 9.3005
R19700 gnd.n4311 gnd.n4042 9.3005
R19701 gnd.n4165 gnd.n4163 9.3005
R19702 gnd.n4159 gnd.n4158 9.3005
R19703 gnd.n4157 gnd.n4109 9.3005
R19704 gnd.n4156 gnd.n4155 9.3005
R19705 gnd.n4152 gnd.n4112 9.3005
R19706 gnd.n4151 gnd.n4148 9.3005
R19707 gnd.n4147 gnd.n4113 9.3005
R19708 gnd.n4146 gnd.n4145 9.3005
R19709 gnd.n4142 gnd.n4114 9.3005
R19710 gnd.n4141 gnd.n4138 9.3005
R19711 gnd.n4137 gnd.n4115 9.3005
R19712 gnd.n4136 gnd.n4135 9.3005
R19713 gnd.n4132 gnd.n4116 9.3005
R19714 gnd.n4131 gnd.n4128 9.3005
R19715 gnd.n4127 gnd.n4117 9.3005
R19716 gnd.n4126 gnd.n4125 9.3005
R19717 gnd.n4122 gnd.n4118 9.3005
R19718 gnd.n4121 gnd.n2462 9.3005
R19719 gnd.n4160 gnd.n4105 9.3005
R19720 gnd.n4162 gnd.n4161 9.3005
R19721 gnd.n6395 gnd.n2831 9.3005
R19722 gnd.n6398 gnd.n2830 9.3005
R19723 gnd.n6399 gnd.n2829 9.3005
R19724 gnd.n6402 gnd.n2828 9.3005
R19725 gnd.n6403 gnd.n2827 9.3005
R19726 gnd.n6406 gnd.n2826 9.3005
R19727 gnd.n6407 gnd.n2825 9.3005
R19728 gnd.n6410 gnd.n2824 9.3005
R19729 gnd.n6412 gnd.n2821 9.3005
R19730 gnd.n6415 gnd.n2820 9.3005
R19731 gnd.n6416 gnd.n2819 9.3005
R19732 gnd.n6419 gnd.n2818 9.3005
R19733 gnd.n6420 gnd.n2817 9.3005
R19734 gnd.n6423 gnd.n2816 9.3005
R19735 gnd.n6424 gnd.n2815 9.3005
R19736 gnd.n6427 gnd.n2814 9.3005
R19737 gnd.n6428 gnd.n2813 9.3005
R19738 gnd.n6431 gnd.n2812 9.3005
R19739 gnd.n6432 gnd.n2811 9.3005
R19740 gnd.n6435 gnd.n2810 9.3005
R19741 gnd.n6436 gnd.n2809 9.3005
R19742 gnd.n6439 gnd.n2808 9.3005
R19743 gnd.n6440 gnd.n2807 9.3005
R19744 gnd.n6441 gnd.n2806 9.3005
R19745 gnd.n2763 gnd.n2762 9.3005
R19746 gnd.n6447 gnd.n6446 9.3005
R19747 gnd.n4646 gnd.n4643 9.3005
R19748 gnd.n4650 gnd.n4649 9.3005
R19749 gnd.n4651 gnd.n4641 9.3005
R19750 gnd.n4653 gnd.n4652 9.3005
R19751 gnd.n4656 gnd.n4640 9.3005
R19752 gnd.n4660 gnd.n4659 9.3005
R19753 gnd.n4661 gnd.n4639 9.3005
R19754 gnd.n4664 gnd.n4662 9.3005
R19755 gnd.n4665 gnd.n4635 9.3005
R19756 gnd.n4669 gnd.n4668 9.3005
R19757 gnd.n4670 gnd.n4634 9.3005
R19758 gnd.n4672 gnd.n4671 9.3005
R19759 gnd.n4675 gnd.n4633 9.3005
R19760 gnd.n4679 gnd.n4678 9.3005
R19761 gnd.n4680 gnd.n4632 9.3005
R19762 gnd.n4682 gnd.n4681 9.3005
R19763 gnd.n4685 gnd.n4631 9.3005
R19764 gnd.n4689 gnd.n4688 9.3005
R19765 gnd.n4690 gnd.n4630 9.3005
R19766 gnd.n4692 gnd.n4691 9.3005
R19767 gnd.n4695 gnd.n4629 9.3005
R19768 gnd.n4699 gnd.n4698 9.3005
R19769 gnd.n4700 gnd.n4628 9.3005
R19770 gnd.n4702 gnd.n4701 9.3005
R19771 gnd.n4705 gnd.n4627 9.3005
R19772 gnd.n4709 gnd.n4708 9.3005
R19773 gnd.n4710 gnd.n4626 9.3005
R19774 gnd.n4713 gnd.n4711 9.3005
R19775 gnd.n4714 gnd.n4622 9.3005
R19776 gnd.n4717 gnd.n4716 9.3005
R19777 gnd.n4642 gnd.n2832 9.3005
R19778 gnd.n2484 gnd.n2464 9.3005
R19779 gnd.n4073 gnd.n2485 9.3005
R19780 gnd.n6613 gnd.n2486 9.3005
R19781 gnd.n6612 gnd.n2487 9.3005
R19782 gnd.n6611 gnd.n2488 9.3005
R19783 gnd.n4079 gnd.n2489 9.3005
R19784 gnd.n6601 gnd.n2505 9.3005
R19785 gnd.n6600 gnd.n2506 9.3005
R19786 gnd.n6599 gnd.n2507 9.3005
R19787 gnd.n4086 gnd.n2508 9.3005
R19788 gnd.n6589 gnd.n2524 9.3005
R19789 gnd.n6588 gnd.n2525 9.3005
R19790 gnd.n6587 gnd.n2526 9.3005
R19791 gnd.n4093 gnd.n2527 9.3005
R19792 gnd.n6577 gnd.n2544 9.3005
R19793 gnd.n6576 gnd.n2545 9.3005
R19794 gnd.n6575 gnd.n2546 9.3005
R19795 gnd.n4203 gnd.n2547 9.3005
R19796 gnd.n6565 gnd.n2564 9.3005
R19797 gnd.n6564 gnd.n2565 9.3005
R19798 gnd.n6563 gnd.n2566 9.3005
R19799 gnd.n4206 gnd.n2567 9.3005
R19800 gnd.n6553 gnd.n2584 9.3005
R19801 gnd.n6552 gnd.n2585 9.3005
R19802 gnd.n6551 gnd.n2586 9.3005
R19803 gnd.n4261 gnd.n2587 9.3005
R19804 gnd.n6541 gnd.n2603 9.3005
R19805 gnd.n6540 gnd.n2604 9.3005
R19806 gnd.n6539 gnd.n2605 9.3005
R19807 gnd.n4270 gnd.n2606 9.3005
R19808 gnd.n4269 gnd.n4268 9.3005
R19809 gnd.n4038 gnd.n4033 9.3005
R19810 gnd.n4329 gnd.n4034 9.3005
R19811 gnd.n4328 gnd.n4035 9.3005
R19812 gnd.n4327 gnd.n4325 9.3005
R19813 gnd.n4036 gnd.n2630 9.3005
R19814 gnd.n6528 gnd.n2631 9.3005
R19815 gnd.n6527 gnd.n2632 9.3005
R19816 gnd.n6526 gnd.n2633 9.3005
R19817 gnd.n4006 gnd.n2634 9.3005
R19818 gnd.n6516 gnd.n2649 9.3005
R19819 gnd.n6515 gnd.n2650 9.3005
R19820 gnd.n6514 gnd.n2651 9.3005
R19821 gnd.n4000 gnd.n2652 9.3005
R19822 gnd.n6504 gnd.n2670 9.3005
R19823 gnd.n6503 gnd.n2671 9.3005
R19824 gnd.n6502 gnd.n2672 9.3005
R19825 gnd.n4404 gnd.n2673 9.3005
R19826 gnd.n6492 gnd.n2689 9.3005
R19827 gnd.n6491 gnd.n2690 9.3005
R19828 gnd.n6490 gnd.n2691 9.3005
R19829 gnd.n4414 gnd.n2692 9.3005
R19830 gnd.n6480 gnd.n2710 9.3005
R19831 gnd.n6479 gnd.n2711 9.3005
R19832 gnd.n6478 gnd.n2712 9.3005
R19833 gnd.n3975 gnd.n2713 9.3005
R19834 gnd.n6468 gnd.n2729 9.3005
R19835 gnd.n6467 gnd.n2730 9.3005
R19836 gnd.n6466 gnd.n2731 9.3005
R19837 gnd.n4471 gnd.n2732 9.3005
R19838 gnd.n6456 gnd.n2750 9.3005
R19839 gnd.n6455 gnd.n2751 9.3005
R19840 gnd.n6454 gnd.n2752 9.3005
R19841 gnd.n4719 gnd.n2753 9.3005
R19842 gnd.n6625 gnd.n2463 9.3005
R19843 gnd.n2465 gnd.n2464 9.3005
R19844 gnd.n4074 gnd.n4073 9.3005
R19845 gnd.n4075 gnd.n2486 9.3005
R19846 gnd.n4077 gnd.n2487 9.3005
R19847 gnd.n4078 gnd.n2488 9.3005
R19848 gnd.n4081 gnd.n4079 9.3005
R19849 gnd.n4082 gnd.n2505 9.3005
R19850 gnd.n4084 gnd.n2506 9.3005
R19851 gnd.n4085 gnd.n2507 9.3005
R19852 gnd.n4088 gnd.n4086 9.3005
R19853 gnd.n4089 gnd.n2524 9.3005
R19854 gnd.n4091 gnd.n2525 9.3005
R19855 gnd.n4092 gnd.n2526 9.3005
R19856 gnd.n4095 gnd.n4093 9.3005
R19857 gnd.n4096 gnd.n2544 9.3005
R19858 gnd.n4201 gnd.n2545 9.3005
R19859 gnd.n4202 gnd.n2546 9.3005
R19860 gnd.n4204 gnd.n4203 9.3005
R19861 gnd.n4205 gnd.n2564 9.3005
R19862 gnd.n4209 gnd.n2565 9.3005
R19863 gnd.n4208 gnd.n2566 9.3005
R19864 gnd.n4207 gnd.n4206 9.3005
R19865 gnd.n4059 gnd.n2584 9.3005
R19866 gnd.n4259 gnd.n2585 9.3005
R19867 gnd.n4260 gnd.n2586 9.3005
R19868 gnd.n4262 gnd.n4261 9.3005
R19869 gnd.n4263 gnd.n2603 9.3005
R19870 gnd.n4273 gnd.n2604 9.3005
R19871 gnd.n4272 gnd.n2605 9.3005
R19872 gnd.n4271 gnd.n4270 9.3005
R19873 gnd.n4269 gnd.n4037 9.3005
R19874 gnd.n4317 gnd.n4038 9.3005
R19875 gnd.n4318 gnd.n4034 9.3005
R19876 gnd.n4319 gnd.n4035 9.3005
R19877 gnd.n4325 gnd.n4324 9.3005
R19878 gnd.n4322 gnd.n4036 9.3005
R19879 gnd.n4321 gnd.n2631 9.3005
R19880 gnd.n4320 gnd.n2632 9.3005
R19881 gnd.n4005 gnd.n2633 9.3005
R19882 gnd.n4386 gnd.n4006 9.3005
R19883 gnd.n4387 gnd.n2649 9.3005
R19884 gnd.n4388 gnd.n2650 9.3005
R19885 gnd.n3999 gnd.n2651 9.3005
R19886 gnd.n4400 gnd.n4000 9.3005
R19887 gnd.n4401 gnd.n2670 9.3005
R19888 gnd.n4402 gnd.n2671 9.3005
R19889 gnd.n4403 gnd.n2672 9.3005
R19890 gnd.n4407 gnd.n4404 9.3005
R19891 gnd.n4408 gnd.n2689 9.3005
R19892 gnd.n4412 gnd.n2690 9.3005
R19893 gnd.n4413 gnd.n2691 9.3005
R19894 gnd.n4417 gnd.n4414 9.3005
R19895 gnd.n4416 gnd.n2710 9.3005
R19896 gnd.n4415 gnd.n2711 9.3005
R19897 gnd.n3974 gnd.n2712 9.3005
R19898 gnd.n4467 gnd.n3975 9.3005
R19899 gnd.n4468 gnd.n2729 9.3005
R19900 gnd.n4469 gnd.n2730 9.3005
R19901 gnd.n4470 gnd.n2731 9.3005
R19902 gnd.n4474 gnd.n4471 9.3005
R19903 gnd.n4475 gnd.n2750 9.3005
R19904 gnd.n4722 gnd.n2751 9.3005
R19905 gnd.n4721 gnd.n2752 9.3005
R19906 gnd.n4720 gnd.n4719 9.3005
R19907 gnd.n6625 gnd.n6624 9.3005
R19908 gnd.n6629 gnd.n6628 9.3005
R19909 gnd.n6632 gnd.n2458 9.3005
R19910 gnd.n6633 gnd.n2457 9.3005
R19911 gnd.n6636 gnd.n2456 9.3005
R19912 gnd.n6637 gnd.n2455 9.3005
R19913 gnd.n6640 gnd.n2454 9.3005
R19914 gnd.n6641 gnd.n2453 9.3005
R19915 gnd.n6644 gnd.n2452 9.3005
R19916 gnd.n6645 gnd.n2451 9.3005
R19917 gnd.n6648 gnd.n2450 9.3005
R19918 gnd.n6649 gnd.n2449 9.3005
R19919 gnd.n6652 gnd.n2448 9.3005
R19920 gnd.n6653 gnd.n2447 9.3005
R19921 gnd.n6656 gnd.n2446 9.3005
R19922 gnd.n6657 gnd.n2445 9.3005
R19923 gnd.n6660 gnd.n2444 9.3005
R19924 gnd.n6661 gnd.n2443 9.3005
R19925 gnd.n6664 gnd.n2442 9.3005
R19926 gnd.n6665 gnd.n2441 9.3005
R19927 gnd.n6668 gnd.n2440 9.3005
R19928 gnd.n6672 gnd.n2436 9.3005
R19929 gnd.n6673 gnd.n2435 9.3005
R19930 gnd.n6676 gnd.n2434 9.3005
R19931 gnd.n6677 gnd.n2433 9.3005
R19932 gnd.n6680 gnd.n2432 9.3005
R19933 gnd.n6681 gnd.n2431 9.3005
R19934 gnd.n6684 gnd.n2430 9.3005
R19935 gnd.n6685 gnd.n2429 9.3005
R19936 gnd.n6688 gnd.n2428 9.3005
R19937 gnd.n6689 gnd.n2427 9.3005
R19938 gnd.n6692 gnd.n2426 9.3005
R19939 gnd.n6693 gnd.n2425 9.3005
R19940 gnd.n6696 gnd.n2424 9.3005
R19941 gnd.n6697 gnd.n2423 9.3005
R19942 gnd.n6700 gnd.n2422 9.3005
R19943 gnd.n6701 gnd.n2421 9.3005
R19944 gnd.n6704 gnd.n2420 9.3005
R19945 gnd.n6705 gnd.n2419 9.3005
R19946 gnd.n6708 gnd.n2418 9.3005
R19947 gnd.n6710 gnd.n2415 9.3005
R19948 gnd.n6713 gnd.n2414 9.3005
R19949 gnd.n6714 gnd.n2413 9.3005
R19950 gnd.n6717 gnd.n2412 9.3005
R19951 gnd.n6718 gnd.n2411 9.3005
R19952 gnd.n6721 gnd.n2410 9.3005
R19953 gnd.n6722 gnd.n2409 9.3005
R19954 gnd.n6725 gnd.n2408 9.3005
R19955 gnd.n6726 gnd.n2407 9.3005
R19956 gnd.n6729 gnd.n2406 9.3005
R19957 gnd.n6730 gnd.n2405 9.3005
R19958 gnd.n6733 gnd.n2404 9.3005
R19959 gnd.n6734 gnd.n2403 9.3005
R19960 gnd.n6737 gnd.n2402 9.3005
R19961 gnd.n6739 gnd.n2401 9.3005
R19962 gnd.n6740 gnd.n2400 9.3005
R19963 gnd.n6741 gnd.n2399 9.3005
R19964 gnd.n6742 gnd.n2398 9.3005
R19965 gnd.n6669 gnd.n2437 9.3005
R19966 gnd.n6627 gnd.n2459 9.3005
R19967 gnd.n6619 gnd.n2473 9.3005
R19968 gnd.n6618 gnd.n2474 9.3005
R19969 gnd.n6617 gnd.n2475 9.3005
R19970 gnd.n2495 gnd.n2476 9.3005
R19971 gnd.n6607 gnd.n2496 9.3005
R19972 gnd.n6606 gnd.n2497 9.3005
R19973 gnd.n6605 gnd.n2498 9.3005
R19974 gnd.n2513 gnd.n2499 9.3005
R19975 gnd.n6595 gnd.n2514 9.3005
R19976 gnd.n6594 gnd.n2515 9.3005
R19977 gnd.n6593 gnd.n2516 9.3005
R19978 gnd.n2534 gnd.n2517 9.3005
R19979 gnd.n6583 gnd.n2535 9.3005
R19980 gnd.n6582 gnd.n2536 9.3005
R19981 gnd.n6581 gnd.n2537 9.3005
R19982 gnd.n2553 gnd.n2538 9.3005
R19983 gnd.n6571 gnd.n2554 9.3005
R19984 gnd.n6570 gnd.n2555 9.3005
R19985 gnd.n6569 gnd.n2556 9.3005
R19986 gnd.n2574 gnd.n2557 9.3005
R19987 gnd.n6559 gnd.n2575 9.3005
R19988 gnd.n6558 gnd.n2576 9.3005
R19989 gnd.n6557 gnd.n2577 9.3005
R19990 gnd.n2593 gnd.n2578 9.3005
R19991 gnd.n6547 gnd.n2594 9.3005
R19992 gnd.n6546 gnd.n2595 9.3005
R19993 gnd.n2621 gnd.n2615 9.3005
R19994 gnd.n6522 gnd.n2640 9.3005
R19995 gnd.n6521 gnd.n2641 9.3005
R19996 gnd.n6520 gnd.n2642 9.3005
R19997 gnd.n2659 gnd.n2643 9.3005
R19998 gnd.n6510 gnd.n2660 9.3005
R19999 gnd.n6509 gnd.n2661 9.3005
R20000 gnd.n6508 gnd.n2662 9.3005
R20001 gnd.n2679 gnd.n2663 9.3005
R20002 gnd.n6498 gnd.n2680 9.3005
R20003 gnd.n6497 gnd.n2681 9.3005
R20004 gnd.n6496 gnd.n2682 9.3005
R20005 gnd.n2699 gnd.n2683 9.3005
R20006 gnd.n6486 gnd.n2700 9.3005
R20007 gnd.n6485 gnd.n2701 9.3005
R20008 gnd.n6484 gnd.n2702 9.3005
R20009 gnd.n2719 gnd.n2703 9.3005
R20010 gnd.n6474 gnd.n2720 9.3005
R20011 gnd.n6473 gnd.n2721 9.3005
R20012 gnd.n6472 gnd.n2722 9.3005
R20013 gnd.n2739 gnd.n2723 9.3005
R20014 gnd.n6462 gnd.n2740 9.3005
R20015 gnd.n6461 gnd.n2741 9.3005
R20016 gnd.n6460 gnd.n2742 9.3005
R20017 gnd.n2760 gnd.n2743 9.3005
R20018 gnd.n6450 gnd.n2761 9.3005
R20019 gnd.n6449 gnd.n6448 9.3005
R20020 gnd.n2472 gnd.n2471 9.3005
R20021 gnd.n6533 gnd.n6532 9.3005
R20022 gnd.n4222 gnd.n4221 9.3005
R20023 gnd.n4234 gnd.n4233 9.3005
R20024 gnd.n4235 gnd.n4220 9.3005
R20025 gnd.n4237 gnd.n4236 9.3005
R20026 gnd.n4067 gnd.n4066 9.3005
R20027 gnd.n4242 gnd.n4241 9.3005
R20028 gnd.n4243 gnd.n4065 9.3005
R20029 gnd.n4245 gnd.n4244 9.3005
R20030 gnd.n4052 gnd.n4051 9.3005
R20031 gnd.n4286 gnd.n4285 9.3005
R20032 gnd.n4287 gnd.n4050 9.3005
R20033 gnd.n4289 gnd.n4288 9.3005
R20034 gnd.n4228 gnd.n4227 9.3005
R20035 gnd.n4224 gnd.n951 9.3005
R20036 gnd.n6841 gnd.n950 9.3005
R20037 gnd.n6842 gnd.n949 9.3005
R20038 gnd.n6843 gnd.n948 9.3005
R20039 gnd.n947 gnd.n943 9.3005
R20040 gnd.n6849 gnd.n942 9.3005
R20041 gnd.n6850 gnd.n941 9.3005
R20042 gnd.n6851 gnd.n940 9.3005
R20043 gnd.n939 gnd.n935 9.3005
R20044 gnd.n6857 gnd.n934 9.3005
R20045 gnd.n6858 gnd.n933 9.3005
R20046 gnd.n6859 gnd.n932 9.3005
R20047 gnd.n931 gnd.n927 9.3005
R20048 gnd.n6865 gnd.n926 9.3005
R20049 gnd.n6866 gnd.n925 9.3005
R20050 gnd.n6867 gnd.n924 9.3005
R20051 gnd.n923 gnd.n919 9.3005
R20052 gnd.n6873 gnd.n918 9.3005
R20053 gnd.n6874 gnd.n917 9.3005
R20054 gnd.n6875 gnd.n916 9.3005
R20055 gnd.n915 gnd.n911 9.3005
R20056 gnd.n6881 gnd.n910 9.3005
R20057 gnd.n6882 gnd.n909 9.3005
R20058 gnd.n6883 gnd.n908 9.3005
R20059 gnd.n907 gnd.n903 9.3005
R20060 gnd.n6889 gnd.n902 9.3005
R20061 gnd.n6890 gnd.n901 9.3005
R20062 gnd.n6891 gnd.n900 9.3005
R20063 gnd.n899 gnd.n895 9.3005
R20064 gnd.n6897 gnd.n894 9.3005
R20065 gnd.n6898 gnd.n893 9.3005
R20066 gnd.n6899 gnd.n892 9.3005
R20067 gnd.n891 gnd.n887 9.3005
R20068 gnd.n6905 gnd.n886 9.3005
R20069 gnd.n6906 gnd.n885 9.3005
R20070 gnd.n6907 gnd.n884 9.3005
R20071 gnd.n883 gnd.n879 9.3005
R20072 gnd.n6913 gnd.n878 9.3005
R20073 gnd.n6914 gnd.n877 9.3005
R20074 gnd.n6915 gnd.n876 9.3005
R20075 gnd.n875 gnd.n871 9.3005
R20076 gnd.n6921 gnd.n870 9.3005
R20077 gnd.n6922 gnd.n869 9.3005
R20078 gnd.n6923 gnd.n868 9.3005
R20079 gnd.n867 gnd.n863 9.3005
R20080 gnd.n6929 gnd.n862 9.3005
R20081 gnd.n6930 gnd.n861 9.3005
R20082 gnd.n6931 gnd.n860 9.3005
R20083 gnd.n859 gnd.n855 9.3005
R20084 gnd.n6937 gnd.n854 9.3005
R20085 gnd.n6938 gnd.n853 9.3005
R20086 gnd.n6939 gnd.n852 9.3005
R20087 gnd.n851 gnd.n847 9.3005
R20088 gnd.n6945 gnd.n846 9.3005
R20089 gnd.n6946 gnd.n845 9.3005
R20090 gnd.n6947 gnd.n844 9.3005
R20091 gnd.n843 gnd.n839 9.3005
R20092 gnd.n6953 gnd.n838 9.3005
R20093 gnd.n6954 gnd.n837 9.3005
R20094 gnd.n6955 gnd.n836 9.3005
R20095 gnd.n835 gnd.n831 9.3005
R20096 gnd.n6961 gnd.n830 9.3005
R20097 gnd.n6962 gnd.n829 9.3005
R20098 gnd.n6963 gnd.n828 9.3005
R20099 gnd.n827 gnd.n823 9.3005
R20100 gnd.n6969 gnd.n822 9.3005
R20101 gnd.n6970 gnd.n821 9.3005
R20102 gnd.n6971 gnd.n820 9.3005
R20103 gnd.n819 gnd.n815 9.3005
R20104 gnd.n6977 gnd.n814 9.3005
R20105 gnd.n6978 gnd.n813 9.3005
R20106 gnd.n6979 gnd.n812 9.3005
R20107 gnd.n811 gnd.n807 9.3005
R20108 gnd.n6985 gnd.n806 9.3005
R20109 gnd.n6986 gnd.n805 9.3005
R20110 gnd.n6987 gnd.n804 9.3005
R20111 gnd.n803 gnd.n799 9.3005
R20112 gnd.n6993 gnd.n798 9.3005
R20113 gnd.n6994 gnd.n797 9.3005
R20114 gnd.n6995 gnd.n796 9.3005
R20115 gnd.n795 gnd.n791 9.3005
R20116 gnd.n7001 gnd.n790 9.3005
R20117 gnd.n7002 gnd.n789 9.3005
R20118 gnd.n7003 gnd.n788 9.3005
R20119 gnd.n4226 gnd.n4225 9.3005
R20120 gnd.n5685 gnd.n3003 9.3005
R20121 gnd.n4786 gnd.n4785 9.3005
R20122 gnd.n4787 gnd.n3922 9.3005
R20123 gnd.n4806 gnd.n4805 9.3005
R20124 gnd.n4804 gnd.n3923 9.3005
R20125 gnd.n4803 gnd.n4802 9.3005
R20126 gnd.n4801 gnd.n4788 9.3005
R20127 gnd.n4800 gnd.n4799 9.3005
R20128 gnd.n4798 gnd.n4791 9.3005
R20129 gnd.n4797 gnd.n4796 9.3005
R20130 gnd.n4795 gnd.n4792 9.3005
R20131 gnd.n2917 gnd.n2915 9.3005
R20132 gnd.n6310 gnd.n6309 9.3005
R20133 gnd.n6308 gnd.n2916 9.3005
R20134 gnd.n6307 gnd.n6306 9.3005
R20135 gnd.n6305 gnd.n2918 9.3005
R20136 gnd.n6304 gnd.n6303 9.3005
R20137 gnd.n6302 gnd.n2922 9.3005
R20138 gnd.n6301 gnd.n6300 9.3005
R20139 gnd.n6299 gnd.n2923 9.3005
R20140 gnd.n6298 gnd.n6297 9.3005
R20141 gnd.n6296 gnd.n2927 9.3005
R20142 gnd.n6295 gnd.n6294 9.3005
R20143 gnd.n6293 gnd.n2928 9.3005
R20144 gnd.n6292 gnd.n6291 9.3005
R20145 gnd.n6290 gnd.n2932 9.3005
R20146 gnd.n6289 gnd.n6288 9.3005
R20147 gnd.n6287 gnd.n2933 9.3005
R20148 gnd.n6286 gnd.n6285 9.3005
R20149 gnd.n6284 gnd.n2937 9.3005
R20150 gnd.n6283 gnd.n6282 9.3005
R20151 gnd.n6281 gnd.n2938 9.3005
R20152 gnd.n6280 gnd.n6279 9.3005
R20153 gnd.n6278 gnd.n2942 9.3005
R20154 gnd.n6277 gnd.n6276 9.3005
R20155 gnd.n6275 gnd.n2943 9.3005
R20156 gnd.n6274 gnd.n6273 9.3005
R20157 gnd.n6272 gnd.n2947 9.3005
R20158 gnd.n6271 gnd.n6270 9.3005
R20159 gnd.n6269 gnd.n2948 9.3005
R20160 gnd.n6268 gnd.n6267 9.3005
R20161 gnd.n6266 gnd.n2952 9.3005
R20162 gnd.n6265 gnd.n6264 9.3005
R20163 gnd.n6263 gnd.n2953 9.3005
R20164 gnd.n6262 gnd.n6261 9.3005
R20165 gnd.n6260 gnd.n2957 9.3005
R20166 gnd.n6259 gnd.n6258 9.3005
R20167 gnd.n6257 gnd.n2958 9.3005
R20168 gnd.n6256 gnd.n6255 9.3005
R20169 gnd.n6254 gnd.n2962 9.3005
R20170 gnd.n6253 gnd.n6252 9.3005
R20171 gnd.n6251 gnd.n2963 9.3005
R20172 gnd.n6250 gnd.n6249 9.3005
R20173 gnd.n6248 gnd.n2967 9.3005
R20174 gnd.n6247 gnd.n6246 9.3005
R20175 gnd.n6245 gnd.n2968 9.3005
R20176 gnd.n6244 gnd.n6243 9.3005
R20177 gnd.n6242 gnd.n2972 9.3005
R20178 gnd.n6241 gnd.n6240 9.3005
R20179 gnd.n6239 gnd.n2973 9.3005
R20180 gnd.n6238 gnd.n6237 9.3005
R20181 gnd.n6236 gnd.n2977 9.3005
R20182 gnd.n6235 gnd.n6234 9.3005
R20183 gnd.n6233 gnd.n2978 9.3005
R20184 gnd.n6232 gnd.n6231 9.3005
R20185 gnd.n6230 gnd.n2982 9.3005
R20186 gnd.n6229 gnd.n6228 9.3005
R20187 gnd.n6227 gnd.n2983 9.3005
R20188 gnd.n6226 gnd.n6225 9.3005
R20189 gnd.n6224 gnd.n2987 9.3005
R20190 gnd.n6223 gnd.n6222 9.3005
R20191 gnd.n6221 gnd.n2988 9.3005
R20192 gnd.n6220 gnd.n6219 9.3005
R20193 gnd.n6218 gnd.n2992 9.3005
R20194 gnd.n6217 gnd.n6216 9.3005
R20195 gnd.n6215 gnd.n2993 9.3005
R20196 gnd.n6214 gnd.n6213 9.3005
R20197 gnd.n6212 gnd.n2997 9.3005
R20198 gnd.n6211 gnd.n6210 9.3005
R20199 gnd.n6209 gnd.n2998 9.3005
R20200 gnd.n6208 gnd.n6207 9.3005
R20201 gnd.n6206 gnd.n3002 9.3005
R20202 gnd.n6205 gnd.n6204 9.3005
R20203 gnd.n3925 gnd.n3924 9.3005
R20204 gnd.n4772 gnd.n4771 9.3005
R20205 gnd.n4021 gnd.n4020 9.3005
R20206 gnd.n4340 gnd.n4339 9.3005
R20207 gnd.n4341 gnd.n4019 9.3005
R20208 gnd.n4343 gnd.n4342 9.3005
R20209 gnd.n4009 gnd.n4008 9.3005
R20210 gnd.n4379 gnd.n4378 9.3005
R20211 gnd.n4380 gnd.n4007 9.3005
R20212 gnd.n4382 gnd.n4381 9.3005
R20213 gnd.n4003 gnd.n4002 9.3005
R20214 gnd.n4393 gnd.n4392 9.3005
R20215 gnd.n4394 gnd.n4001 9.3005
R20216 gnd.n4396 gnd.n4395 9.3005
R20217 gnd.n3994 gnd.n3992 9.3005
R20218 gnd.n4431 gnd.n4430 9.3005
R20219 gnd.n4429 gnd.n3993 9.3005
R20220 gnd.n4428 gnd.n4427 9.3005
R20221 gnd.n4426 gnd.n3995 9.3005
R20222 gnd.n4425 gnd.n4424 9.3005
R20223 gnd.n4423 gnd.n3998 9.3005
R20224 gnd.n4422 gnd.n4421 9.3005
R20225 gnd.n3978 gnd.n3977 9.3005
R20226 gnd.n4460 gnd.n4459 9.3005
R20227 gnd.n4461 gnd.n3976 9.3005
R20228 gnd.n4463 gnd.n4462 9.3005
R20229 gnd.n3971 gnd.n3969 9.3005
R20230 gnd.n4735 gnd.n4734 9.3005
R20231 gnd.n4733 gnd.n3970 9.3005
R20232 gnd.n4732 gnd.n4731 9.3005
R20233 gnd.n4730 gnd.n3972 9.3005
R20234 gnd.n4729 gnd.n4728 9.3005
R20235 gnd.n4727 gnd.n4726 9.3005
R20236 gnd.n3956 gnd.n3951 9.3005
R20237 gnd.n4613 gnd.n4612 9.3005
R20238 gnd.n4512 gnd.n4511 9.3005
R20239 gnd.n4607 gnd.n4606 9.3005
R20240 gnd.n4605 gnd.n4604 9.3005
R20241 gnd.n4524 gnd.n4523 9.3005
R20242 gnd.n4599 gnd.n4598 9.3005
R20243 gnd.n4597 gnd.n4596 9.3005
R20244 gnd.n4532 gnd.n4531 9.3005
R20245 gnd.n4591 gnd.n4590 9.3005
R20246 gnd.n4589 gnd.n4588 9.3005
R20247 gnd.n4544 gnd.n4543 9.3005
R20248 gnd.n4583 gnd.n4582 9.3005
R20249 gnd.n4581 gnd.n4580 9.3005
R20250 gnd.n4552 gnd.n4551 9.3005
R20251 gnd.n4575 gnd.n4574 9.3005
R20252 gnd.n4573 gnd.n4572 9.3005
R20253 gnd.n4563 gnd.n3955 9.3005
R20254 gnd.n4768 gnd.n4767 9.3005
R20255 gnd.n4615 gnd.n4614 9.3005
R20256 gnd.n4769 gnd.n3950 9.3005
R20257 gnd.n4569 gnd.n3952 9.3005
R20258 gnd.n4571 gnd.n4570 9.3005
R20259 gnd.n4558 gnd.n4557 9.3005
R20260 gnd.n4577 gnd.n4576 9.3005
R20261 gnd.n4579 gnd.n4578 9.3005
R20262 gnd.n4548 gnd.n4547 9.3005
R20263 gnd.n4585 gnd.n4584 9.3005
R20264 gnd.n4587 gnd.n4586 9.3005
R20265 gnd.n4538 gnd.n4537 9.3005
R20266 gnd.n4593 gnd.n4592 9.3005
R20267 gnd.n4595 gnd.n4594 9.3005
R20268 gnd.n4528 gnd.n4527 9.3005
R20269 gnd.n4601 gnd.n4600 9.3005
R20270 gnd.n4603 gnd.n4602 9.3005
R20271 gnd.n4518 gnd.n4517 9.3005
R20272 gnd.n4609 gnd.n4608 9.3005
R20273 gnd.n4611 gnd.n4610 9.3005
R20274 gnd.n4509 gnd.n4508 9.3005
R20275 gnd.n4617 gnd.n4616 9.3005
R20276 gnd.n4618 gnd.n4476 9.3005
R20277 gnd.n4620 gnd.n4619 9.3005
R20278 gnd.n4503 gnd.n4477 9.3005
R20279 gnd.n4502 gnd.n4501 9.3005
R20280 gnd.n4500 gnd.n4478 9.3005
R20281 gnd.n4499 gnd.n4498 9.3005
R20282 gnd.n4495 gnd.n4481 9.3005
R20283 gnd.n4494 gnd.n4482 9.3005
R20284 gnd.n4489 gnd.n4483 9.3005
R20285 gnd.n4488 gnd.n4487 9.3005
R20286 gnd.n4486 gnd.n4484 9.3005
R20287 gnd.n3907 gnd.n3906 9.3005
R20288 gnd.n4828 gnd.n4827 9.3005
R20289 gnd.n4829 gnd.n3905 9.3005
R20290 gnd.n4831 gnd.n4830 9.3005
R20291 gnd.n3903 gnd.n3902 9.3005
R20292 gnd.n4836 gnd.n4835 9.3005
R20293 gnd.n4837 gnd.n3900 9.3005
R20294 gnd.n4980 gnd.n4979 9.3005
R20295 gnd.n4978 gnd.n3901 9.3005
R20296 gnd.n4977 gnd.n4976 9.3005
R20297 gnd.n4975 gnd.n4838 9.3005
R20298 gnd.n4974 gnd.n4973 9.3005
R20299 gnd.n4972 gnd.n4840 9.3005
R20300 gnd.n4971 gnd.n4970 9.3005
R20301 gnd.n4969 gnd.n4841 9.3005
R20302 gnd.n4968 gnd.n4967 9.3005
R20303 gnd.n4966 gnd.n4843 9.3005
R20304 gnd.n4965 gnd.n4964 9.3005
R20305 gnd.n4963 gnd.n4844 9.3005
R20306 gnd.n4962 gnd.n4961 9.3005
R20307 gnd.n4960 gnd.n4849 9.3005
R20308 gnd.n4959 gnd.n4958 9.3005
R20309 gnd.n4957 gnd.n4850 9.3005
R20310 gnd.n4956 gnd.n4955 9.3005
R20311 gnd.n4954 gnd.n4853 9.3005
R20312 gnd.n4953 gnd.n4952 9.3005
R20313 gnd.n4951 gnd.n4854 9.3005
R20314 gnd.n4950 gnd.n4949 9.3005
R20315 gnd.n4948 gnd.n4857 9.3005
R20316 gnd.n4947 gnd.n4946 9.3005
R20317 gnd.n4945 gnd.n4858 9.3005
R20318 gnd.n4944 gnd.n4943 9.3005
R20319 gnd.n4942 gnd.n4860 9.3005
R20320 gnd.n4941 gnd.n4940 9.3005
R20321 gnd.n4939 gnd.n4861 9.3005
R20322 gnd.n4938 gnd.n4937 9.3005
R20323 gnd.n4936 gnd.n4866 9.3005
R20324 gnd.n4935 gnd.n4934 9.3005
R20325 gnd.n4933 gnd.n4867 9.3005
R20326 gnd.n4932 gnd.n4931 9.3005
R20327 gnd.n4930 gnd.n4869 9.3005
R20328 gnd.n4929 gnd.n4928 9.3005
R20329 gnd.n4927 gnd.n4870 9.3005
R20330 gnd.n4926 gnd.n4925 9.3005
R20331 gnd.n4924 gnd.n4873 9.3005
R20332 gnd.n4923 gnd.n4922 9.3005
R20333 gnd.n4921 gnd.n4874 9.3005
R20334 gnd.n4920 gnd.n4919 9.3005
R20335 gnd.n4918 gnd.n4878 9.3005
R20336 gnd.n4917 gnd.n4916 9.3005
R20337 gnd.n4915 gnd.n4879 9.3005
R20338 gnd.n4914 gnd.n4913 9.3005
R20339 gnd.n4912 gnd.n4882 9.3005
R20340 gnd.n4911 gnd.n4910 9.3005
R20341 gnd.n4909 gnd.n4883 9.3005
R20342 gnd.n4908 gnd.n4907 9.3005
R20343 gnd.n4906 gnd.n4887 9.3005
R20344 gnd.n4905 gnd.n4904 9.3005
R20345 gnd.n4903 gnd.n4888 9.3005
R20346 gnd.n4902 gnd.n4901 9.3005
R20347 gnd.n4900 gnd.n4892 9.3005
R20348 gnd.n4899 gnd.n4898 9.3005
R20349 gnd.n4897 gnd.n4893 9.3005
R20350 gnd.n4896 gnd.n4895 9.3005
R20351 gnd.n3542 gnd.n3541 9.3005
R20352 gnd.n5408 gnd.n5407 9.3005
R20353 gnd.n5409 gnd.n3539 9.3005
R20354 gnd.n5412 gnd.n5411 9.3005
R20355 gnd.n5410 gnd.n3540 9.3005
R20356 gnd.n3443 gnd.n3442 9.3005
R20357 gnd.n5556 gnd.n5555 9.3005
R20358 gnd.n5557 gnd.n3441 9.3005
R20359 gnd.n5559 gnd.n5558 9.3005
R20360 gnd.n3431 gnd.n3430 9.3005
R20361 gnd.n5575 gnd.n5574 9.3005
R20362 gnd.n5576 gnd.n3429 9.3005
R20363 gnd.n5578 gnd.n5577 9.3005
R20364 gnd.n3012 gnd.n3011 9.3005
R20365 gnd.n6200 gnd.n6199 9.3005
R20366 gnd.n4491 gnd.n4490 9.3005
R20367 gnd.n6196 gnd.n3013 9.3005
R20368 gnd.n6195 gnd.n6194 9.3005
R20369 gnd.n6193 gnd.n3016 9.3005
R20370 gnd.n6192 gnd.n6191 9.3005
R20371 gnd.n6190 gnd.n3017 9.3005
R20372 gnd.n6189 gnd.n6188 9.3005
R20373 gnd.n6198 gnd.n6197 9.3005
R20374 gnd.n6141 gnd.n6140 9.3005
R20375 gnd.n3064 gnd.n3063 9.3005
R20376 gnd.n6147 gnd.n6146 9.3005
R20377 gnd.n6149 gnd.n6148 9.3005
R20378 gnd.n3056 gnd.n3055 9.3005
R20379 gnd.n6155 gnd.n6154 9.3005
R20380 gnd.n6157 gnd.n6156 9.3005
R20381 gnd.n3048 gnd.n3047 9.3005
R20382 gnd.n6163 gnd.n6162 9.3005
R20383 gnd.n6165 gnd.n6164 9.3005
R20384 gnd.n3040 gnd.n3039 9.3005
R20385 gnd.n6171 gnd.n6170 9.3005
R20386 gnd.n6173 gnd.n6172 9.3005
R20387 gnd.n3032 gnd.n3031 9.3005
R20388 gnd.n6179 gnd.n6178 9.3005
R20389 gnd.n6181 gnd.n6180 9.3005
R20390 gnd.n3028 gnd.n3023 9.3005
R20391 gnd.n6139 gnd.n3073 9.3005
R20392 gnd.n3394 gnd.n3072 9.3005
R20393 gnd.n6186 gnd.n3021 9.3005
R20394 gnd.n6185 gnd.n6184 9.3005
R20395 gnd.n6183 gnd.n6182 9.3005
R20396 gnd.n3027 gnd.n3026 9.3005
R20397 gnd.n6177 gnd.n6176 9.3005
R20398 gnd.n6175 gnd.n6174 9.3005
R20399 gnd.n3036 gnd.n3035 9.3005
R20400 gnd.n6169 gnd.n6168 9.3005
R20401 gnd.n6167 gnd.n6166 9.3005
R20402 gnd.n3044 gnd.n3043 9.3005
R20403 gnd.n6161 gnd.n6160 9.3005
R20404 gnd.n6159 gnd.n6158 9.3005
R20405 gnd.n3052 gnd.n3051 9.3005
R20406 gnd.n6153 gnd.n6152 9.3005
R20407 gnd.n6151 gnd.n6150 9.3005
R20408 gnd.n3060 gnd.n3059 9.3005
R20409 gnd.n6145 gnd.n6144 9.3005
R20410 gnd.n6143 gnd.n6142 9.3005
R20411 gnd.n3417 gnd.n3070 9.3005
R20412 gnd.n3396 gnd.n3395 9.3005
R20413 gnd.n5687 gnd.n5686 9.3005
R20414 gnd.n5691 gnd.n5690 9.3005
R20415 gnd.n5692 gnd.n3391 9.3005
R20416 gnd.n5696 gnd.n5695 9.3005
R20417 gnd.n5697 gnd.n3390 9.3005
R20418 gnd.n5699 gnd.n5698 9.3005
R20419 gnd.n3388 gnd.n3387 9.3005
R20420 gnd.n5711 gnd.n5710 9.3005
R20421 gnd.n5712 gnd.n3386 9.3005
R20422 gnd.n5714 gnd.n5713 9.3005
R20423 gnd.n3384 gnd.n3383 9.3005
R20424 gnd.n5726 gnd.n5725 9.3005
R20425 gnd.n5727 gnd.n3382 9.3005
R20426 gnd.n5729 gnd.n5728 9.3005
R20427 gnd.n3379 gnd.n3378 9.3005
R20428 gnd.n5741 gnd.n5740 9.3005
R20429 gnd.n5742 gnd.n3377 9.3005
R20430 gnd.n5744 gnd.n5743 9.3005
R20431 gnd.n3375 gnd.n3374 9.3005
R20432 gnd.n5756 gnd.n5755 9.3005
R20433 gnd.n5757 gnd.n3373 9.3005
R20434 gnd.n5759 gnd.n5758 9.3005
R20435 gnd.n3370 gnd.n3369 9.3005
R20436 gnd.n5771 gnd.n5770 9.3005
R20437 gnd.n5772 gnd.n3367 9.3005
R20438 gnd.n5786 gnd.n5785 9.3005
R20439 gnd.n5784 gnd.n3368 9.3005
R20440 gnd.n5783 gnd.n5782 9.3005
R20441 gnd.n5781 gnd.n5773 9.3005
R20442 gnd.n5780 gnd.n5779 9.3005
R20443 gnd.n5778 gnd.n5777 9.3005
R20444 gnd.n5776 gnd.n95 9.3005
R20445 gnd.n5689 gnd.n3392 9.3005
R20446 gnd.n8072 gnd.n96 9.3005
R20447 gnd.n1952 gnd.t219 9.24152
R20448 gnd.n6815 gnd.t338 9.24152
R20449 gnd.n2345 gnd.t307 9.24152
R20450 gnd.n6579 gnd.t44 9.24152
R20451 gnd.n6494 gnd.t21 9.24152
R20452 gnd.n5738 gnd.t62 9.24152
R20453 gnd.n8023 gnd.t8 9.24152
R20454 gnd.t379 gnd.t219 8.92286
R20455 gnd.n5065 gnd.n3788 8.92286
R20456 gnd.n5100 gnd.n5099 8.92286
R20457 gnd.n5189 gnd.n3707 8.92286
R20458 gnd.n5223 gnd.n5222 8.92286
R20459 gnd.n5307 gnd.n3625 8.92286
R20460 gnd.n5340 gnd.n3596 8.92286
R20461 gnd.n5545 gnd.n5544 8.92286
R20462 gnd.n2325 gnd.n2300 8.92171
R20463 gnd.n2293 gnd.n2268 8.92171
R20464 gnd.n2261 gnd.n2236 8.92171
R20465 gnd.n2230 gnd.n2205 8.92171
R20466 gnd.n2198 gnd.n2173 8.92171
R20467 gnd.n2166 gnd.n2141 8.92171
R20468 gnd.n2134 gnd.n2109 8.92171
R20469 gnd.n2103 gnd.n2078 8.92171
R20470 gnd.n3479 gnd.n3461 8.72777
R20471 gnd.n1874 gnd.t4 8.60421
R20472 gnd.n6603 gnd.t25 8.60421
R20473 gnd.n6470 gnd.t35 8.60421
R20474 gnd.t217 gnd.n5188 8.60421
R20475 gnd.n5200 gnd.t356 8.60421
R20476 gnd.n5708 gnd.t48 8.60421
R20477 gnd.n7999 gnd.t50 8.60421
R20478 gnd.n1292 gnd.n1272 8.43656
R20479 gnd.n54 gnd.n34 8.43656
R20480 gnd.n4990 gnd.t269 8.28555
R20481 gnd.n2326 gnd.n2298 8.14595
R20482 gnd.n2294 gnd.n2266 8.14595
R20483 gnd.n2262 gnd.n2234 8.14595
R20484 gnd.n2231 gnd.n2203 8.14595
R20485 gnd.n2199 gnd.n2171 8.14595
R20486 gnd.n2167 gnd.n2139 8.14595
R20487 gnd.n2135 gnd.n2107 8.14595
R20488 gnd.n2104 gnd.n2076 8.14595
R20489 gnd.n4312 gnd.n0 8.10675
R20490 gnd.n8073 gnd.n8072 8.10675
R20491 gnd.n2331 gnd.n2330 7.97301
R20492 gnd.t381 gnd.n1824 7.9669
R20493 gnd.n6585 gnd.n2529 7.9669
R20494 gnd.n5025 gnd.t349 7.9669
R20495 gnd.n5373 gnd.t390 7.9669
R20496 gnd.n8017 gnd.n191 7.9669
R20497 gnd.n8073 gnd.n94 7.95236
R20498 gnd.n6139 gnd.n3072 7.75808
R20499 gnd.n4767 gnd.n3955 7.75808
R20500 gnd.n7793 gnd.n7740 7.75808
R20501 gnd.n4161 gnd.n4160 7.75808
R20502 gnd.t348 gnd.n3792 7.64824
R20503 gnd.n5146 gnd.t341 7.64824
R20504 gnd.n5156 gnd.t341 7.64824
R20505 gnd.n5249 gnd.t216 7.64824
R20506 gnd.n5257 gnd.t216 7.64824
R20507 gnd.t365 gnd.n3582 7.64824
R20508 gnd.n1333 gnd.n1332 7.53171
R20509 gnd.n1757 gnd.t394 7.32958
R20510 gnd.n4229 gnd.t44 7.32958
R20511 gnd.n7708 gnd.t8 7.32958
R20512 gnd.n2893 gnd.n2892 7.30353
R20513 gnd.n3478 gnd.n3477 7.30353
R20514 gnd.n1717 gnd.n1436 7.01093
R20515 gnd.n1439 gnd.n1437 7.01093
R20516 gnd.n1727 gnd.n1726 7.01093
R20517 gnd.n1738 gnd.n1420 7.01093
R20518 gnd.n1737 gnd.n1423 7.01093
R20519 gnd.n1748 gnd.n1411 7.01093
R20520 gnd.n1414 gnd.n1412 7.01093
R20521 gnd.n1758 gnd.n1757 7.01093
R20522 gnd.n1768 gnd.n1392 7.01093
R20523 gnd.n1767 gnd.n1395 7.01093
R20524 gnd.n1784 gnd.n1385 7.01093
R20525 gnd.n1794 gnd.n1376 7.01093
R20526 gnd.n1805 gnd.n1804 7.01093
R20527 gnd.n1825 gnd.n1361 7.01093
R20528 gnd.n1824 gnd.n1340 7.01093
R20529 gnd.n1842 gnd.n1341 7.01093
R20530 gnd.n1836 gnd.n1835 7.01093
R20531 gnd.n1852 gnd.n1240 7.01093
R20532 gnd.n1861 gnd.n1231 7.01093
R20533 gnd.n1870 gnd.n1223 7.01093
R20534 gnd.n1874 gnd.n1873 7.01093
R20535 gnd.n1892 gnd.n1208 7.01093
R20536 gnd.n1891 gnd.n1211 7.01093
R20537 gnd.n1902 gnd.n1200 7.01093
R20538 gnd.n1201 gnd.n1190 7.01093
R20539 gnd.n1941 gnd.n1183 7.01093
R20540 gnd.n1940 gnd.n1939 7.01093
R20541 gnd.n1952 gnd.n1951 7.01093
R20542 gnd.n1176 gnd.n1168 7.01093
R20543 gnd.n1963 gnd.n1962 7.01093
R20544 gnd.n1981 gnd.n1156 7.01093
R20545 gnd.n1980 gnd.n1159 7.01093
R20546 gnd.n2004 gnd.n1139 7.01093
R20547 gnd.n2042 gnd.n1131 7.01093
R20548 gnd.n2041 gnd.n1123 7.01093
R20549 gnd.n2057 gnd.n2056 7.01093
R20550 gnd.n2035 gnd.n953 7.01093
R20551 gnd.n6836 gnd.n955 7.01093
R20552 gnd.n6830 gnd.n6829 7.01093
R20553 gnd.n1112 gnd.n967 7.01093
R20554 gnd.n6823 gnd.n976 7.01093
R20555 gnd.n6822 gnd.n979 7.01093
R20556 gnd.n2022 gnd.n988 7.01093
R20557 gnd.n6816 gnd.n6815 7.01093
R20558 gnd.n2346 gnd.n2345 7.01093
R20559 gnd.n6809 gnd.n1001 7.01093
R20560 gnd.n6808 gnd.n1004 7.01093
R20561 gnd.n5175 gnd.t351 7.01093
R20562 gnd.n5239 gnd.t389 7.01093
R20563 gnd.n1395 gnd.t208 6.69227
R20564 gnd.n1939 gnd.t379 6.69227
R20565 gnd.t209 gnd.n964 6.69227
R20566 gnd.n4247 gnd.t110 6.69227
R20567 gnd.n4738 gnd.t35 6.69227
R20568 gnd.n3794 gnd.t212 6.69227
R20569 gnd.t392 gnd.n3589 6.69227
R20570 gnd.t48 gnd.n3225 6.69227
R20571 gnd.n5862 gnd.t73 6.69227
R20572 gnd.n5474 gnd.n5473 6.5566
R20573 gnd.n3833 gnd.n3832 6.5566
R20574 gnd.n6331 gnd.n6327 6.5566
R20575 gnd.n5486 gnd.n3506 6.5566
R20576 gnd.n6837 gnd.n6836 6.37362
R20577 gnd.n5004 gnd.n3818 6.37362
R20578 gnd.n5033 gnd.n5031 6.37362
R20579 gnd.n5128 gnd.n5127 6.37362
R20580 gnd.n5277 gnd.n5276 6.37362
R20581 gnd.n5367 gnd.n5366 6.37362
R20582 gnd.n5379 gnd.n3556 6.37362
R20583 gnd.n4570 gnd.n4566 6.20656
R20584 gnd.n3417 gnd.n3069 6.20656
R20585 gnd.t382 gnd.n1816 6.05496
R20586 gnd.n1817 gnd.t358 6.05496
R20587 gnd.t377 gnd.n1208 6.05496
R20588 gnd.n1991 gnd.t373 6.05496
R20589 gnd.n4306 gnd.t87 6.05496
R20590 gnd.n4409 gnd.t21 6.05496
R20591 gnd.n6390 gnd.n2839 6.05496
R20592 gnd.t62 gnd.n3266 6.05496
R20593 gnd.t18 gnd.n101 6.05496
R20594 gnd.n2328 gnd.n2298 5.81868
R20595 gnd.n2296 gnd.n2266 5.81868
R20596 gnd.n2264 gnd.n2234 5.81868
R20597 gnd.n2233 gnd.n2203 5.81868
R20598 gnd.n2201 gnd.n2171 5.81868
R20599 gnd.n2169 gnd.n2139 5.81868
R20600 gnd.n2137 gnd.n2107 5.81868
R20601 gnd.n2106 gnd.n2076 5.81868
R20602 gnd.t245 gnd.n2871 5.73631
R20603 gnd.n3892 gnd.t245 5.73631
R20604 gnd.n5012 gnd.t248 5.73631
R20605 gnd.n5065 gnd.t364 5.73631
R20606 gnd.n5135 gnd.t361 5.73631
R20607 gnd.n5268 gnd.t388 5.73631
R20608 gnd.n5340 gnd.t360 5.73631
R20609 gnd.n3508 gnd.n3149 5.62001
R20610 gnd.n6393 gnd.n2835 5.62001
R20611 gnd.n6393 gnd.n2836 5.62001
R20612 gnd.n5484 gnd.n3149 5.62001
R20613 gnd.n1576 gnd.n1571 5.4308
R20614 gnd.n1105 gnd.n1035 5.4308
R20615 gnd.n1211 gnd.t374 5.41765
R20616 gnd.n1905 gnd.t220 5.41765
R20617 gnd.t396 gnd.n1138 5.41765
R20618 gnd.n4375 gnd.t58 5.41765
R20619 gnd.n4004 gnd.t129 5.41765
R20620 gnd.n5091 gnd.t368 5.41765
R20621 gnd.n3620 gnd.t210 5.41765
R20622 gnd.t94 gnd.n3307 5.41765
R20623 gnd.t10 gnd.n3326 5.41765
R20624 gnd.t298 gnd.n6318 5.09899
R20625 gnd.n5013 gnd.n5012 5.09899
R20626 gnd.n5025 gnd.n5024 5.09899
R20627 gnd.n5117 gnd.t347 5.09899
R20628 gnd.n3738 gnd.n3733 5.09899
R20629 gnd.n5149 gnd.n5148 5.09899
R20630 gnd.n3656 gnd.n3650 5.09899
R20631 gnd.n5270 gnd.n5269 5.09899
R20632 gnd.n5293 gnd.t343 5.09899
R20633 gnd.n5373 gnd.n3568 5.09899
R20634 gnd.n5395 gnd.n3553 5.09899
R20635 gnd.n2326 gnd.n2325 5.04292
R20636 gnd.n2294 gnd.n2293 5.04292
R20637 gnd.n2262 gnd.n2261 5.04292
R20638 gnd.n2231 gnd.n2230 5.04292
R20639 gnd.n2199 gnd.n2198 5.04292
R20640 gnd.n2167 gnd.n2166 5.04292
R20641 gnd.n2135 gnd.n2134 5.04292
R20642 gnd.n2104 gnd.n2103 5.04292
R20643 gnd.n1862 gnd.t7 4.78034
R20644 gnd.n1962 gnd.t3 4.78034
R20645 gnd.t68 gnd.n4023 4.78034
R20646 gnd.n4434 gnd.t46 4.78034
R20647 gnd.n3776 gnd.t368 4.78034
R20648 gnd.t210 gnd.n3610 4.78034
R20649 gnd.n3447 gnd.t314 4.78034
R20650 gnd.t16 gnd.n3284 4.78034
R20651 gnd.t119 gnd.n3343 4.78034
R20652 gnd.n1337 gnd.n1334 4.74817
R20653 gnd.n1849 gnd.n1242 4.74817
R20654 gnd.n1847 gnd.n1244 4.74817
R20655 gnd.n1253 gnd.n1251 4.74817
R20656 gnd.n1353 gnd.n1334 4.74817
R20657 gnd.n1352 gnd.n1242 4.74817
R20658 gnd.n1848 gnd.n1847 4.74817
R20659 gnd.n1253 gnd.n1252 4.74817
R20660 gnd.n3345 gnd.n114 4.74817
R20661 gnd.n5917 gnd.n113 4.74817
R20662 gnd.n3349 gnd.n112 4.74817
R20663 gnd.n8065 gnd.n107 4.74817
R20664 gnd.n8063 gnd.n108 4.74817
R20665 gnd.n5930 gnd.n114 4.74817
R20666 gnd.n3346 gnd.n113 4.74817
R20667 gnd.n5916 gnd.n112 4.74817
R20668 gnd.n3348 gnd.n107 4.74817
R20669 gnd.n8064 gnd.n8063 4.74817
R20670 gnd.n4290 gnd.n4048 4.74817
R20671 gnd.n4304 gnd.n4295 4.74817
R20672 gnd.n4302 gnd.n4301 4.74817
R20673 gnd.n4297 gnd.n4296 4.74817
R20674 gnd.n4349 gnd.n4013 4.74817
R20675 gnd.n5924 gnd.n5923 4.74817
R20676 gnd.n5814 gnd.n3337 4.74817
R20677 gnd.n5815 gnd.n5813 4.74817
R20678 gnd.n5822 gnd.n5821 4.74817
R20679 gnd.n5896 gnd.n5895 4.74817
R20680 gnd.n5925 gnd.n5924 4.74817
R20681 gnd.n5922 gnd.n3337 4.74817
R20682 gnd.n5816 gnd.n5815 4.74817
R20683 gnd.n5821 gnd.n5820 4.74817
R20684 gnd.n5897 gnd.n5896 4.74817
R20685 gnd.n2613 gnd.n2596 4.74817
R20686 gnd.n6534 gnd.n2614 4.74817
R20687 gnd.n4028 gnd.n2619 4.74817
R20688 gnd.n4335 gnd.n2618 4.74817
R20689 gnd.n2620 gnd.n2617 4.74817
R20690 gnd.n6545 gnd.n2596 4.74817
R20691 gnd.n6535 gnd.n6534 4.74817
R20692 gnd.n4264 gnd.n2619 4.74817
R20693 gnd.n4029 gnd.n2618 4.74817
R20694 gnd.n4334 gnd.n2617 4.74817
R20695 gnd.n4293 gnd.n4048 4.74817
R20696 gnd.n4295 gnd.n4294 4.74817
R20697 gnd.n4303 gnd.n4302 4.74817
R20698 gnd.n4298 gnd.n4297 4.74817
R20699 gnd.n4015 gnd.n4013 4.74817
R20700 gnd.n1332 gnd.n1331 4.74296
R20701 gnd.n94 gnd.n93 4.74296
R20702 gnd.n1292 gnd.n1291 4.7074
R20703 gnd.n1312 gnd.n1311 4.7074
R20704 gnd.n54 gnd.n53 4.7074
R20705 gnd.n74 gnd.n73 4.7074
R20706 gnd.n1332 gnd.n1312 4.65959
R20707 gnd.n94 gnd.n74 4.65959
R20708 gnd.n6081 gnd.n3151 4.6132
R20709 gnd.n6394 gnd.n2834 4.6132
R20710 gnd.n6444 gnd.n2765 4.46168
R20711 gnd.n4990 gnd.t234 4.46168
R20712 gnd.n5386 gnd.t265 4.46168
R20713 gnd.n6134 gnd.n3117 4.46168
R20714 gnd.n3474 gnd.n3461 4.46111
R20715 gnd.n2311 gnd.n2307 4.38594
R20716 gnd.n2279 gnd.n2275 4.38594
R20717 gnd.n2247 gnd.n2243 4.38594
R20718 gnd.n2216 gnd.n2212 4.38594
R20719 gnd.n2184 gnd.n2180 4.38594
R20720 gnd.n2152 gnd.n2148 4.38594
R20721 gnd.n2120 gnd.n2116 4.38594
R20722 gnd.n2089 gnd.n2085 4.38594
R20723 gnd.n2322 gnd.n2300 4.26717
R20724 gnd.n2290 gnd.n2268 4.26717
R20725 gnd.n2258 gnd.n2236 4.26717
R20726 gnd.n2227 gnd.n2205 4.26717
R20727 gnd.n2195 gnd.n2173 4.26717
R20728 gnd.n2163 gnd.n2141 4.26717
R20729 gnd.n2131 gnd.n2109 4.26717
R20730 gnd.n2100 gnd.n2078 4.26717
R20731 gnd.t6 gnd.n1368 4.14303
R20732 gnd.n2056 gnd.t5 4.14303
R20733 gnd.n4282 gnd.t23 4.14303
R20734 gnd.n4456 gnd.t56 4.14303
R20735 gnd.t384 gnd.n5155 4.14303
R20736 gnd.n5250 gnd.t375 4.14303
R20737 gnd.t14 gnd.n3243 4.14303
R20738 gnd.n5891 gnd.t41 4.14303
R20739 gnd.n2330 gnd.n2329 4.08274
R20740 gnd.n5473 gnd.n5472 4.05904
R20741 gnd.n3834 gnd.n3833 4.05904
R20742 gnd.n6334 gnd.n6327 4.05904
R20743 gnd.n3506 gnd.n3501 4.05904
R20744 gnd.n15 gnd.n7 3.99943
R20745 gnd.n6319 gnd.t298 3.82437
R20746 gnd.n4997 gnd.n3823 3.82437
R20747 gnd.n3809 gnd.n3798 3.82437
R20748 gnd.n5129 gnd.n3742 3.82437
R20749 gnd.n3729 gnd.n3718 3.82437
R20750 gnd.n5251 gnd.n3660 3.82437
R20751 gnd.n4876 gnd.n3646 3.82437
R20752 gnd.n3585 gnd.n3572 3.82437
R20753 gnd.n5379 gnd.t289 3.82437
R20754 gnd.n5405 gnd.n3544 3.82437
R20755 gnd.n1846 gnd.n1333 3.81325
R20756 gnd.n1312 gnd.n1292 3.72967
R20757 gnd.n74 gnd.n54 3.72967
R20758 gnd.n2330 gnd.n2202 3.70378
R20759 gnd.n15 gnd.n14 3.60163
R20760 gnd.n2478 gnd.t230 3.50571
R20761 gnd.n4218 gnd.t85 3.50571
R20762 gnd.n4724 gnd.t251 3.50571
R20763 gnd.n6005 gnd.t226 3.50571
R20764 gnd.n7715 gnd.t12 3.50571
R20765 gnd.t238 gnd.n240 3.50571
R20766 gnd.n2321 gnd.n2302 3.49141
R20767 gnd.n2289 gnd.n2270 3.49141
R20768 gnd.n2257 gnd.n2238 3.49141
R20769 gnd.n2226 gnd.n2207 3.49141
R20770 gnd.n2194 gnd.n2175 3.49141
R20771 gnd.n2162 gnd.n2143 3.49141
R20772 gnd.n2130 gnd.n2111 3.49141
R20773 gnd.n2099 gnd.n2080 3.49141
R20774 gnd.n6099 gnd.n6098 3.29747
R20775 gnd.n6098 gnd.n6097 3.29747
R20776 gnd.n7940 gnd.n7937 3.29747
R20777 gnd.n7941 gnd.n7940 3.29747
R20778 gnd.n6710 gnd.n6709 3.29747
R20779 gnd.n6709 gnd.n6708 3.29747
R20780 gnd.n6412 gnd.n6411 3.29747
R20781 gnd.n6411 gnd.n6410 3.29747
R20782 gnd.n6312 gnd.t234 3.18706
R20783 gnd.t265 gnd.n3564 3.18706
R20784 gnd.n1375 gnd.t6 2.8684
R20785 gnd.n1313 gnd.t77 2.82907
R20786 gnd.n1313 gnd.t175 2.82907
R20787 gnd.n1315 gnd.t47 2.82907
R20788 gnd.n1315 gnd.t100 2.82907
R20789 gnd.n1317 gnd.t130 2.82907
R20790 gnd.n1317 gnd.t106 2.82907
R20791 gnd.n1319 gnd.t99 2.82907
R20792 gnd.n1319 gnd.t91 2.82907
R20793 gnd.n1321 gnd.t113 2.82907
R20794 gnd.n1321 gnd.t168 2.82907
R20795 gnd.n1323 gnd.t24 2.82907
R20796 gnd.n1323 gnd.t147 2.82907
R20797 gnd.n1325 gnd.t195 2.82907
R20798 gnd.n1325 gnd.t111 2.82907
R20799 gnd.n1327 gnd.t151 2.82907
R20800 gnd.n1327 gnd.t86 2.82907
R20801 gnd.n1329 gnd.t38 2.82907
R20802 gnd.n1329 gnd.t34 2.82907
R20803 gnd.n1254 gnd.t118 2.82907
R20804 gnd.n1254 gnd.t146 2.82907
R20805 gnd.n1256 gnd.t161 2.82907
R20806 gnd.n1256 gnd.t79 2.82907
R20807 gnd.n1258 gnd.t143 2.82907
R20808 gnd.n1258 gnd.t122 2.82907
R20809 gnd.n1260 gnd.t198 2.82907
R20810 gnd.n1260 gnd.t187 2.82907
R20811 gnd.n1262 gnd.t88 2.82907
R20812 gnd.n1262 gnd.t154 2.82907
R20813 gnd.n1264 gnd.t182 2.82907
R20814 gnd.n1264 gnd.t28 2.82907
R20815 gnd.n1266 gnd.t54 2.82907
R20816 gnd.n1266 gnd.t144 2.82907
R20817 gnd.n1268 gnd.t155 2.82907
R20818 gnd.n1268 gnd.t196 2.82907
R20819 gnd.n1270 gnd.t112 2.82907
R20820 gnd.n1270 gnd.t134 2.82907
R20821 gnd.n1273 gnd.t205 2.82907
R20822 gnd.n1273 gnd.t57 2.82907
R20823 gnd.n1275 gnd.t55 2.82907
R20824 gnd.n1275 gnd.t22 2.82907
R20825 gnd.n1277 gnd.t164 2.82907
R20826 gnd.n1277 gnd.t206 2.82907
R20827 gnd.n1279 gnd.t200 2.82907
R20828 gnd.n1279 gnd.t59 2.82907
R20829 gnd.n1281 gnd.t189 2.82907
R20830 gnd.n1281 gnd.t165 2.82907
R20831 gnd.n1283 gnd.t166 2.82907
R20832 gnd.n1283 gnd.t202 2.82907
R20833 gnd.n1285 gnd.t197 2.82907
R20834 gnd.n1285 gnd.t183 2.82907
R20835 gnd.n1287 gnd.t178 2.82907
R20836 gnd.n1287 gnd.t167 2.82907
R20837 gnd.n1289 gnd.t160 2.82907
R20838 gnd.n1289 gnd.t148 2.82907
R20839 gnd.n1293 gnd.t138 2.82907
R20840 gnd.n1293 gnd.t80 2.82907
R20841 gnd.n1295 gnd.t117 2.82907
R20842 gnd.n1295 gnd.t162 2.82907
R20843 gnd.n1297 gnd.t199 2.82907
R20844 gnd.n1297 gnd.t181 2.82907
R20845 gnd.n1299 gnd.t179 2.82907
R20846 gnd.n1299 gnd.t153 2.82907
R20847 gnd.n1301 gnd.t177 2.82907
R20848 gnd.n1301 gnd.t69 2.82907
R20849 gnd.n1303 gnd.t97 2.82907
R20850 gnd.n1303 gnd.t39 2.82907
R20851 gnd.n1305 gnd.t90 2.82907
R20852 gnd.n1305 gnd.t176 2.82907
R20853 gnd.n1307 gnd.t45 2.82907
R20854 gnd.n1307 gnd.t145 2.82907
R20855 gnd.n1309 gnd.t107 2.82907
R20856 gnd.n1309 gnd.t104 2.82907
R20857 gnd.n91 gnd.t116 2.82907
R20858 gnd.n91 gnd.t125 2.82907
R20859 gnd.n89 gnd.t13 2.82907
R20860 gnd.n89 gnd.t103 2.82907
R20861 gnd.n87 gnd.t74 2.82907
R20862 gnd.n87 gnd.t126 2.82907
R20863 gnd.n85 gnd.t84 2.82907
R20864 gnd.n85 gnd.t158 2.82907
R20865 gnd.n83 gnd.t120 2.82907
R20866 gnd.n83 gnd.t89 2.82907
R20867 gnd.n81 gnd.t40 2.82907
R20868 gnd.n81 gnd.t66 2.82907
R20869 gnd.n79 gnd.t71 2.82907
R20870 gnd.n79 gnd.t95 2.82907
R20871 gnd.n77 gnd.t63 2.82907
R20872 gnd.n77 gnd.t180 2.82907
R20873 gnd.n75 gnd.t137 2.82907
R20874 gnd.n75 gnd.t32 2.82907
R20875 gnd.n32 gnd.t115 2.82907
R20876 gnd.n32 gnd.t128 2.82907
R20877 gnd.n30 gnd.t67 2.82907
R20878 gnd.n30 gnd.t9 2.82907
R20879 gnd.n28 gnd.t190 2.82907
R20880 gnd.n28 gnd.t92 2.82907
R20881 gnd.n26 gnd.t83 2.82907
R20882 gnd.n26 gnd.t42 2.82907
R20883 gnd.n24 gnd.t207 2.82907
R20884 gnd.n24 gnd.t75 2.82907
R20885 gnd.n22 gnd.t52 2.82907
R20886 gnd.n22 gnd.t72 2.82907
R20887 gnd.n20 gnd.t174 2.82907
R20888 gnd.n20 gnd.t131 2.82907
R20889 gnd.n18 gnd.t108 2.82907
R20890 gnd.n18 gnd.t20 2.82907
R20891 gnd.n16 gnd.t194 2.82907
R20892 gnd.n16 gnd.t96 2.82907
R20893 gnd.n51 gnd.t156 2.82907
R20894 gnd.n51 gnd.t133 2.82907
R20895 gnd.n49 gnd.t141 2.82907
R20896 gnd.n49 gnd.t152 2.82907
R20897 gnd.n47 gnd.t149 2.82907
R20898 gnd.n47 gnd.t170 2.82907
R20899 gnd.n45 gnd.t171 2.82907
R20900 gnd.n45 gnd.t142 2.82907
R20901 gnd.n43 gnd.t139 2.82907
R20902 gnd.n43 gnd.t19 2.82907
R20903 gnd.n41 gnd.t11 2.82907
R20904 gnd.n41 gnd.t169 2.82907
R20905 gnd.n39 gnd.t184 2.82907
R20906 gnd.n39 gnd.t192 2.82907
R20907 gnd.n37 gnd.t191 2.82907
R20908 gnd.n37 gnd.t17 2.82907
R20909 gnd.n35 gnd.t15 2.82907
R20910 gnd.n35 gnd.t43 2.82907
R20911 gnd.n71 gnd.t186 2.82907
R20912 gnd.n71 gnd.t203 2.82907
R20913 gnd.n69 gnd.t93 2.82907
R20914 gnd.n69 gnd.t173 2.82907
R20915 gnd.n67 gnd.t136 2.82907
R20916 gnd.n67 gnd.t30 2.82907
R20917 gnd.n65 gnd.t163 2.82907
R20918 gnd.n65 gnd.t61 2.82907
R20919 gnd.n63 gnd.t193 2.82907
R20920 gnd.n63 gnd.t150 2.82907
R20921 gnd.n61 gnd.t109 2.82907
R20922 gnd.n61 gnd.t132 2.82907
R20923 gnd.n59 gnd.t135 2.82907
R20924 gnd.n59 gnd.t159 2.82907
R20925 gnd.n57 gnd.t121 2.82907
R20926 gnd.n57 gnd.t78 2.82907
R20927 gnd.n55 gnd.t204 2.82907
R20928 gnd.n55 gnd.t102 2.82907
R20929 gnd.n2318 gnd.n2317 2.71565
R20930 gnd.n2286 gnd.n2285 2.71565
R20931 gnd.n2254 gnd.n2253 2.71565
R20932 gnd.n2223 gnd.n2222 2.71565
R20933 gnd.n2191 gnd.n2190 2.71565
R20934 gnd.n2159 gnd.n2158 2.71565
R20935 gnd.n2127 gnd.n2126 2.71565
R20936 gnd.n2096 gnd.n2095 2.71565
R20937 gnd.n4983 gnd.n4982 2.54975
R20938 gnd.n5058 gnd.n3794 2.54975
R20939 gnd.n5083 gnd.t387 2.54975
R20940 gnd.n5107 gnd.n3755 2.54975
R20941 gnd.n3756 gnd.t347 2.54975
R20942 gnd.n5182 gnd.n3714 2.54975
R20943 gnd.n5230 gnd.n3674 2.54975
R20944 gnd.t343 gnd.n3629 2.54975
R20945 gnd.n5300 gnd.n3631 2.54975
R20946 gnd.n5323 gnd.t342 2.54975
R20947 gnd.n5352 gnd.n3589 2.54975
R20948 gnd.n5414 gnd.n3537 2.54975
R20949 gnd.n1846 gnd.n1334 2.27742
R20950 gnd.n1846 gnd.n1242 2.27742
R20951 gnd.n1847 gnd.n1846 2.27742
R20952 gnd.n1846 gnd.n1253 2.27742
R20953 gnd.n8062 gnd.n114 2.27742
R20954 gnd.n8062 gnd.n113 2.27742
R20955 gnd.n8062 gnd.n112 2.27742
R20956 gnd.n8062 gnd.n107 2.27742
R20957 gnd.n8063 gnd.n8062 2.27742
R20958 gnd.n5924 gnd.n111 2.27742
R20959 gnd.n3337 gnd.n111 2.27742
R20960 gnd.n5815 gnd.n111 2.27742
R20961 gnd.n5821 gnd.n111 2.27742
R20962 gnd.n5896 gnd.n111 2.27742
R20963 gnd.n6533 gnd.n2596 2.27742
R20964 gnd.n6534 gnd.n6533 2.27742
R20965 gnd.n6533 gnd.n2619 2.27742
R20966 gnd.n6533 gnd.n2618 2.27742
R20967 gnd.n6533 gnd.n2617 2.27742
R20968 gnd.n4048 gnd.n2616 2.27742
R20969 gnd.n4295 gnd.n2616 2.27742
R20970 gnd.n4302 gnd.n2616 2.27742
R20971 gnd.n4297 gnd.n2616 2.27742
R20972 gnd.n4013 gnd.n2616 2.27742
R20973 gnd.n1726 gnd.t275 2.23109
R20974 gnd.n1851 gnd.t7 2.23109
R20975 gnd.n5156 gnd.t384 2.23109
R20976 gnd.t375 gnd.n5249 2.23109
R20977 gnd.n2314 gnd.n2304 1.93989
R20978 gnd.n2282 gnd.n2272 1.93989
R20979 gnd.n2250 gnd.n2240 1.93989
R20980 gnd.n2219 gnd.n2209 1.93989
R20981 gnd.n2187 gnd.n2177 1.93989
R20982 gnd.n2155 gnd.n2145 1.93989
R20983 gnd.n2123 gnd.n2113 1.93989
R20984 gnd.n2092 gnd.n2082 1.93989
R20985 gnd.t214 gnd.n1737 1.59378
R20986 gnd.n1914 gnd.t220 1.59378
R20987 gnd.n1149 gnd.t396 1.59378
R20988 gnd.t33 gnd.n2522 1.59378
R20989 gnd.n4419 gnd.t76 1.59378
R20990 gnd.n5975 gnd.t31 1.59378
R20991 gnd.n199 gnd.t114 1.59378
R20992 gnd.n6320 gnd.n2897 1.27512
R20993 gnd.n4997 gnd.t323 1.27512
R20994 gnd.n5064 gnd.n3781 1.27512
R20995 gnd.n5076 gnd.n3771 1.27512
R20996 gnd.n5188 gnd.n3702 1.27512
R20997 gnd.n5200 gnd.n3691 1.27512
R20998 gnd.n5306 gnd.n3618 1.27512
R20999 gnd.n5333 gnd.n3603 1.27512
R21000 gnd.n5415 gnd.t292 1.27512
R21001 gnd.n3457 gnd.n3456 1.27512
R21002 gnd.t314 gnd.n3446 1.27512
R21003 gnd.n1579 gnd.n1571 1.16414
R21004 gnd.n1102 gnd.n1035 1.16414
R21005 gnd.n2313 gnd.n2306 1.16414
R21006 gnd.n2281 gnd.n2274 1.16414
R21007 gnd.n2249 gnd.n2242 1.16414
R21008 gnd.n2218 gnd.n2211 1.16414
R21009 gnd.n2186 gnd.n2179 1.16414
R21010 gnd.n2154 gnd.n2147 1.16414
R21011 gnd.n2122 gnd.n2115 1.16414
R21012 gnd.n2091 gnd.n2084 1.16414
R21013 gnd.n6081 gnd.n6080 0.970197
R21014 gnd.n6394 gnd.n2832 0.970197
R21015 gnd.n2297 gnd.n2265 0.962709
R21016 gnd.n2329 gnd.n2297 0.962709
R21017 gnd.n2170 gnd.n2138 0.962709
R21018 gnd.n2202 gnd.n2170 0.962709
R21019 gnd.n1817 gnd.t382 0.956468
R21020 gnd.n1926 gnd.t373 0.956468
R21021 gnd.n4211 gnd.t53 0.956468
R21022 gnd.n4398 gnd.t105 0.956468
R21023 gnd.n4982 gnd.t398 0.956468
R21024 gnd.t344 gnd.n5414 0.956468
R21025 gnd.n5951 gnd.t70 0.956468
R21026 gnd.n5872 gnd.t29 0.956468
R21027 gnd.n2 gnd.n1 0.672012
R21028 gnd.n3 gnd.n2 0.672012
R21029 gnd.n4 gnd.n3 0.672012
R21030 gnd.n5 gnd.n4 0.672012
R21031 gnd.n6 gnd.n5 0.672012
R21032 gnd.n7 gnd.n6 0.672012
R21033 gnd.n9 gnd.n8 0.672012
R21034 gnd.n10 gnd.n9 0.672012
R21035 gnd.n11 gnd.n10 0.672012
R21036 gnd.n12 gnd.n11 0.672012
R21037 gnd.n13 gnd.n12 0.672012
R21038 gnd.n14 gnd.n13 0.672012
R21039 gnd.n5023 gnd.t2 0.637812
R21040 gnd.t351 gnd.n3711 0.637812
R21041 gnd.n3675 gnd.t389 0.637812
R21042 gnd.t372 gnd.n3575 0.637812
R21043 gnd.n3564 gnd.t262 0.637812
R21044 gnd.n8074 gnd.n8073 0.63688
R21045 gnd gnd.n0 0.634843
R21046 gnd.n1331 gnd.n1330 0.573776
R21047 gnd.n1330 gnd.n1328 0.573776
R21048 gnd.n1328 gnd.n1326 0.573776
R21049 gnd.n1326 gnd.n1324 0.573776
R21050 gnd.n1324 gnd.n1322 0.573776
R21051 gnd.n1322 gnd.n1320 0.573776
R21052 gnd.n1320 gnd.n1318 0.573776
R21053 gnd.n1318 gnd.n1316 0.573776
R21054 gnd.n1316 gnd.n1314 0.573776
R21055 gnd.n1272 gnd.n1271 0.573776
R21056 gnd.n1271 gnd.n1269 0.573776
R21057 gnd.n1269 gnd.n1267 0.573776
R21058 gnd.n1267 gnd.n1265 0.573776
R21059 gnd.n1265 gnd.n1263 0.573776
R21060 gnd.n1263 gnd.n1261 0.573776
R21061 gnd.n1261 gnd.n1259 0.573776
R21062 gnd.n1259 gnd.n1257 0.573776
R21063 gnd.n1257 gnd.n1255 0.573776
R21064 gnd.n1291 gnd.n1290 0.573776
R21065 gnd.n1290 gnd.n1288 0.573776
R21066 gnd.n1288 gnd.n1286 0.573776
R21067 gnd.n1286 gnd.n1284 0.573776
R21068 gnd.n1284 gnd.n1282 0.573776
R21069 gnd.n1282 gnd.n1280 0.573776
R21070 gnd.n1280 gnd.n1278 0.573776
R21071 gnd.n1278 gnd.n1276 0.573776
R21072 gnd.n1276 gnd.n1274 0.573776
R21073 gnd.n1311 gnd.n1310 0.573776
R21074 gnd.n1310 gnd.n1308 0.573776
R21075 gnd.n1308 gnd.n1306 0.573776
R21076 gnd.n1306 gnd.n1304 0.573776
R21077 gnd.n1304 gnd.n1302 0.573776
R21078 gnd.n1302 gnd.n1300 0.573776
R21079 gnd.n1300 gnd.n1298 0.573776
R21080 gnd.n1298 gnd.n1296 0.573776
R21081 gnd.n1296 gnd.n1294 0.573776
R21082 gnd.n78 gnd.n76 0.573776
R21083 gnd.n80 gnd.n78 0.573776
R21084 gnd.n82 gnd.n80 0.573776
R21085 gnd.n84 gnd.n82 0.573776
R21086 gnd.n86 gnd.n84 0.573776
R21087 gnd.n88 gnd.n86 0.573776
R21088 gnd.n90 gnd.n88 0.573776
R21089 gnd.n92 gnd.n90 0.573776
R21090 gnd.n93 gnd.n92 0.573776
R21091 gnd.n19 gnd.n17 0.573776
R21092 gnd.n21 gnd.n19 0.573776
R21093 gnd.n23 gnd.n21 0.573776
R21094 gnd.n25 gnd.n23 0.573776
R21095 gnd.n27 gnd.n25 0.573776
R21096 gnd.n29 gnd.n27 0.573776
R21097 gnd.n31 gnd.n29 0.573776
R21098 gnd.n33 gnd.n31 0.573776
R21099 gnd.n34 gnd.n33 0.573776
R21100 gnd.n38 gnd.n36 0.573776
R21101 gnd.n40 gnd.n38 0.573776
R21102 gnd.n42 gnd.n40 0.573776
R21103 gnd.n44 gnd.n42 0.573776
R21104 gnd.n46 gnd.n44 0.573776
R21105 gnd.n48 gnd.n46 0.573776
R21106 gnd.n50 gnd.n48 0.573776
R21107 gnd.n52 gnd.n50 0.573776
R21108 gnd.n53 gnd.n52 0.573776
R21109 gnd.n58 gnd.n56 0.573776
R21110 gnd.n60 gnd.n58 0.573776
R21111 gnd.n62 gnd.n60 0.573776
R21112 gnd.n64 gnd.n62 0.573776
R21113 gnd.n66 gnd.n64 0.573776
R21114 gnd.n68 gnd.n66 0.573776
R21115 gnd.n70 gnd.n68 0.573776
R21116 gnd.n72 gnd.n70 0.573776
R21117 gnd.n73 gnd.n72 0.573776
R21118 gnd.n6205 gnd.n3003 0.489829
R21119 gnd.n4771 gnd.n3924 0.489829
R21120 gnd.n4490 gnd.n4482 0.489829
R21121 gnd.n6199 gnd.n6198 0.489829
R21122 gnd.n2352 gnd.n2351 0.486781
R21123 gnd.n1628 gnd.n1627 0.48678
R21124 gnd.n6754 gnd.n6753 0.480683
R21125 gnd.n1712 gnd.n1711 0.480683
R21126 gnd.n7792 gnd.n7737 0.477634
R21127 gnd.n4163 gnd.n4162 0.477634
R21128 gnd.n788 gnd.n783 0.447146
R21129 gnd.n7493 gnd.n7492 0.447146
R21130 gnd.n7705 gnd.n7704 0.447146
R21131 gnd.n4227 gnd.n4226 0.447146
R21132 gnd.n7977 gnd.n7976 0.442573
R21133 gnd.n3202 gnd.n3121 0.442573
R21134 gnd.n6448 gnd.n6447 0.442573
R21135 gnd.n2472 gnd.n2398 0.442573
R21136 gnd.n8062 gnd.n111 0.4255
R21137 gnd.n6533 gnd.n2616 0.4255
R21138 gnd.n4566 gnd.n4557 0.388379
R21139 gnd.n2310 gnd.n2309 0.388379
R21140 gnd.n2278 gnd.n2277 0.388379
R21141 gnd.n2246 gnd.n2245 0.388379
R21142 gnd.n2215 gnd.n2214 0.388379
R21143 gnd.n2183 gnd.n2182 0.388379
R21144 gnd.n2151 gnd.n2150 0.388379
R21145 gnd.n2119 gnd.n2118 0.388379
R21146 gnd.n2088 gnd.n2087 0.388379
R21147 gnd.n6143 gnd.n3069 0.388379
R21148 gnd.n8074 gnd.n15 0.374463
R21149 gnd.n2031 gnd.t209 0.319156
R21150 gnd.n4275 gnd.t27 0.319156
R21151 gnd.t98 gnd.n4345 0.319156
R21152 gnd.n5115 gnd.t354 0.319156
R21153 gnd.t386 gnd.t217 0.319156
R21154 gnd.t356 gnd.t346 0.319156
R21155 gnd.n5294 gnd.t402 0.319156
R21156 gnd.t65 gnd.n3333 0.319156
R21157 gnd.n5829 gnd.t82 0.319156
R21158 gnd.n1546 gnd.n1524 0.311721
R21159 gnd gnd.n8074 0.295112
R21160 gnd.n7853 gnd.n354 0.293183
R21161 gnd.n6626 gnd.n2462 0.293183
R21162 gnd.n6799 gnd.n1009 0.268793
R21163 gnd.n7854 gnd.n7853 0.258122
R21164 gnd.n6019 gnd.n3022 0.258122
R21165 gnd.n4718 gnd.n4717 0.258122
R21166 gnd.n6627 gnd.n6626 0.258122
R21167 gnd.n4770 gnd.n3951 0.247451
R21168 gnd.n5689 gnd.n5688 0.247451
R21169 gnd.n1049 gnd.n1009 0.241354
R21170 gnd.n3151 gnd.n3148 0.229039
R21171 gnd.n3152 gnd.n3151 0.229039
R21172 gnd.n2834 gnd.n2831 0.229039
R21173 gnd.n4642 gnd.n2834 0.229039
R21174 gnd.n1333 gnd.n0 0.210825
R21175 gnd.n1700 gnd.n1499 0.206293
R21176 gnd.n2327 gnd.n2299 0.155672
R21177 gnd.n2320 gnd.n2299 0.155672
R21178 gnd.n2320 gnd.n2319 0.155672
R21179 gnd.n2319 gnd.n2303 0.155672
R21180 gnd.n2312 gnd.n2303 0.155672
R21181 gnd.n2312 gnd.n2311 0.155672
R21182 gnd.n2295 gnd.n2267 0.155672
R21183 gnd.n2288 gnd.n2267 0.155672
R21184 gnd.n2288 gnd.n2287 0.155672
R21185 gnd.n2287 gnd.n2271 0.155672
R21186 gnd.n2280 gnd.n2271 0.155672
R21187 gnd.n2280 gnd.n2279 0.155672
R21188 gnd.n2263 gnd.n2235 0.155672
R21189 gnd.n2256 gnd.n2235 0.155672
R21190 gnd.n2256 gnd.n2255 0.155672
R21191 gnd.n2255 gnd.n2239 0.155672
R21192 gnd.n2248 gnd.n2239 0.155672
R21193 gnd.n2248 gnd.n2247 0.155672
R21194 gnd.n2232 gnd.n2204 0.155672
R21195 gnd.n2225 gnd.n2204 0.155672
R21196 gnd.n2225 gnd.n2224 0.155672
R21197 gnd.n2224 gnd.n2208 0.155672
R21198 gnd.n2217 gnd.n2208 0.155672
R21199 gnd.n2217 gnd.n2216 0.155672
R21200 gnd.n2200 gnd.n2172 0.155672
R21201 gnd.n2193 gnd.n2172 0.155672
R21202 gnd.n2193 gnd.n2192 0.155672
R21203 gnd.n2192 gnd.n2176 0.155672
R21204 gnd.n2185 gnd.n2176 0.155672
R21205 gnd.n2185 gnd.n2184 0.155672
R21206 gnd.n2168 gnd.n2140 0.155672
R21207 gnd.n2161 gnd.n2140 0.155672
R21208 gnd.n2161 gnd.n2160 0.155672
R21209 gnd.n2160 gnd.n2144 0.155672
R21210 gnd.n2153 gnd.n2144 0.155672
R21211 gnd.n2153 gnd.n2152 0.155672
R21212 gnd.n2136 gnd.n2108 0.155672
R21213 gnd.n2129 gnd.n2108 0.155672
R21214 gnd.n2129 gnd.n2128 0.155672
R21215 gnd.n2128 gnd.n2112 0.155672
R21216 gnd.n2121 gnd.n2112 0.155672
R21217 gnd.n2121 gnd.n2120 0.155672
R21218 gnd.n2105 gnd.n2077 0.155672
R21219 gnd.n2098 gnd.n2077 0.155672
R21220 gnd.n2098 gnd.n2097 0.155672
R21221 gnd.n2097 gnd.n2081 0.155672
R21222 gnd.n2090 gnd.n2081 0.155672
R21223 gnd.n2090 gnd.n2089 0.155672
R21224 gnd.n6788 gnd.n6754 0.152939
R21225 gnd.n6788 gnd.n6787 0.152939
R21226 gnd.n6787 gnd.n6786 0.152939
R21227 gnd.n6786 gnd.n6756 0.152939
R21228 gnd.n6757 gnd.n6756 0.152939
R21229 gnd.n6758 gnd.n6757 0.152939
R21230 gnd.n6759 gnd.n6758 0.152939
R21231 gnd.n6760 gnd.n6759 0.152939
R21232 gnd.n6761 gnd.n6760 0.152939
R21233 gnd.n6762 gnd.n6761 0.152939
R21234 gnd.n6763 gnd.n6762 0.152939
R21235 gnd.n6764 gnd.n6763 0.152939
R21236 gnd.n6764 gnd.n1015 0.152939
R21237 gnd.n6797 gnd.n1015 0.152939
R21238 gnd.n6798 gnd.n6797 0.152939
R21239 gnd.n6799 gnd.n6798 0.152939
R21240 gnd.n1713 gnd.n1712 0.152939
R21241 gnd.n1713 gnd.n1417 0.152939
R21242 gnd.n1741 gnd.n1417 0.152939
R21243 gnd.n1742 gnd.n1741 0.152939
R21244 gnd.n1743 gnd.n1742 0.152939
R21245 gnd.n1744 gnd.n1743 0.152939
R21246 gnd.n1744 gnd.n1389 0.152939
R21247 gnd.n1771 gnd.n1389 0.152939
R21248 gnd.n1772 gnd.n1771 0.152939
R21249 gnd.n1773 gnd.n1772 0.152939
R21250 gnd.n1774 gnd.n1773 0.152939
R21251 gnd.n1775 gnd.n1774 0.152939
R21252 gnd.n1777 gnd.n1775 0.152939
R21253 gnd.n1777 gnd.n1776 0.152939
R21254 gnd.n1776 gnd.n1357 0.152939
R21255 gnd.n1830 gnd.n1357 0.152939
R21256 gnd.n1831 gnd.n1830 0.152939
R21257 gnd.n1832 gnd.n1831 0.152939
R21258 gnd.n1832 gnd.n1226 0.152939
R21259 gnd.n1865 gnd.n1226 0.152939
R21260 gnd.n1866 gnd.n1865 0.152939
R21261 gnd.n1867 gnd.n1866 0.152939
R21262 gnd.n1867 gnd.n1205 0.152939
R21263 gnd.n1895 gnd.n1205 0.152939
R21264 gnd.n1896 gnd.n1895 0.152939
R21265 gnd.n1897 gnd.n1896 0.152939
R21266 gnd.n1898 gnd.n1897 0.152939
R21267 gnd.n1898 gnd.n1180 0.152939
R21268 gnd.n1944 gnd.n1180 0.152939
R21269 gnd.n1945 gnd.n1944 0.152939
R21270 gnd.n1946 gnd.n1945 0.152939
R21271 gnd.n1947 gnd.n1946 0.152939
R21272 gnd.n1947 gnd.n1153 0.152939
R21273 gnd.n1984 gnd.n1153 0.152939
R21274 gnd.n1985 gnd.n1984 0.152939
R21275 gnd.n1986 gnd.n1985 0.152939
R21276 gnd.n1987 gnd.n1986 0.152939
R21277 gnd.n1987 gnd.n1128 0.152939
R21278 gnd.n2045 gnd.n1128 0.152939
R21279 gnd.n2046 gnd.n2045 0.152939
R21280 gnd.n2047 gnd.n2046 0.152939
R21281 gnd.n2048 gnd.n2047 0.152939
R21282 gnd.n2050 gnd.n2048 0.152939
R21283 gnd.n2050 gnd.n2049 0.152939
R21284 gnd.n2049 gnd.n971 0.152939
R21285 gnd.n972 gnd.n971 0.152939
R21286 gnd.n973 gnd.n972 0.152939
R21287 gnd.n994 gnd.n973 0.152939
R21288 gnd.n995 gnd.n994 0.152939
R21289 gnd.n996 gnd.n995 0.152939
R21290 gnd.n997 gnd.n996 0.152939
R21291 gnd.n998 gnd.n997 0.152939
R21292 gnd.n6753 gnd.n998 0.152939
R21293 gnd.n1711 gnd.n1441 0.152939
R21294 gnd.n1462 gnd.n1441 0.152939
R21295 gnd.n1463 gnd.n1462 0.152939
R21296 gnd.n1469 gnd.n1463 0.152939
R21297 gnd.n1470 gnd.n1469 0.152939
R21298 gnd.n1471 gnd.n1470 0.152939
R21299 gnd.n1471 gnd.n1460 0.152939
R21300 gnd.n1479 gnd.n1460 0.152939
R21301 gnd.n1480 gnd.n1479 0.152939
R21302 gnd.n1481 gnd.n1480 0.152939
R21303 gnd.n1481 gnd.n1458 0.152939
R21304 gnd.n1489 gnd.n1458 0.152939
R21305 gnd.n1490 gnd.n1489 0.152939
R21306 gnd.n1491 gnd.n1490 0.152939
R21307 gnd.n1491 gnd.n1456 0.152939
R21308 gnd.n1499 gnd.n1456 0.152939
R21309 gnd.n1050 gnd.n1049 0.152939
R21310 gnd.n1051 gnd.n1050 0.152939
R21311 gnd.n1051 gnd.n1045 0.152939
R21312 gnd.n1059 gnd.n1045 0.152939
R21313 gnd.n1060 gnd.n1059 0.152939
R21314 gnd.n1061 gnd.n1060 0.152939
R21315 gnd.n1061 gnd.n1043 0.152939
R21316 gnd.n1069 gnd.n1043 0.152939
R21317 gnd.n1070 gnd.n1069 0.152939
R21318 gnd.n1071 gnd.n1070 0.152939
R21319 gnd.n1071 gnd.n1041 0.152939
R21320 gnd.n1079 gnd.n1041 0.152939
R21321 gnd.n1080 gnd.n1079 0.152939
R21322 gnd.n1081 gnd.n1080 0.152939
R21323 gnd.n1081 gnd.n1039 0.152939
R21324 gnd.n1089 gnd.n1039 0.152939
R21325 gnd.n1090 gnd.n1089 0.152939
R21326 gnd.n1091 gnd.n1090 0.152939
R21327 gnd.n1091 gnd.n1037 0.152939
R21328 gnd.n1099 gnd.n1037 0.152939
R21329 gnd.n1100 gnd.n1099 0.152939
R21330 gnd.n1101 gnd.n1100 0.152939
R21331 gnd.n1101 gnd.n1032 0.152939
R21332 gnd.n1108 gnd.n1032 0.152939
R21333 gnd.n1109 gnd.n1108 0.152939
R21334 gnd.n2352 gnd.n1109 0.152939
R21335 gnd.n1246 gnd.n1245 0.152939
R21336 gnd.n1246 gnd.n1187 0.152939
R21337 gnd.n1917 gnd.n1187 0.152939
R21338 gnd.n1918 gnd.n1917 0.152939
R21339 gnd.n1919 gnd.n1918 0.152939
R21340 gnd.n1920 gnd.n1919 0.152939
R21341 gnd.n1921 gnd.n1920 0.152939
R21342 gnd.n1922 gnd.n1921 0.152939
R21343 gnd.n1923 gnd.n1922 0.152939
R21344 gnd.n1924 gnd.n1923 0.152939
R21345 gnd.n1925 gnd.n1924 0.152939
R21346 gnd.n1925 gnd.n1135 0.152939
R21347 gnd.n2007 gnd.n1135 0.152939
R21348 gnd.n2008 gnd.n2007 0.152939
R21349 gnd.n2009 gnd.n2008 0.152939
R21350 gnd.n2010 gnd.n2009 0.152939
R21351 gnd.n2011 gnd.n2010 0.152939
R21352 gnd.n2012 gnd.n2011 0.152939
R21353 gnd.n2013 gnd.n2012 0.152939
R21354 gnd.n2014 gnd.n2013 0.152939
R21355 gnd.n2015 gnd.n2014 0.152939
R21356 gnd.n2016 gnd.n2015 0.152939
R21357 gnd.n2017 gnd.n2016 0.152939
R21358 gnd.n2018 gnd.n2017 0.152939
R21359 gnd.n2020 gnd.n2018 0.152939
R21360 gnd.n2020 gnd.n2019 0.152939
R21361 gnd.n2019 gnd.n1110 0.152939
R21362 gnd.n2351 gnd.n1110 0.152939
R21363 gnd.n1629 gnd.n1628 0.152939
R21364 gnd.n1629 gnd.n1519 0.152939
R21365 gnd.n1644 gnd.n1519 0.152939
R21366 gnd.n1645 gnd.n1644 0.152939
R21367 gnd.n1646 gnd.n1645 0.152939
R21368 gnd.n1646 gnd.n1507 0.152939
R21369 gnd.n1660 gnd.n1507 0.152939
R21370 gnd.n1661 gnd.n1660 0.152939
R21371 gnd.n1662 gnd.n1661 0.152939
R21372 gnd.n1663 gnd.n1662 0.152939
R21373 gnd.n1664 gnd.n1663 0.152939
R21374 gnd.n1665 gnd.n1664 0.152939
R21375 gnd.n1666 gnd.n1665 0.152939
R21376 gnd.n1667 gnd.n1666 0.152939
R21377 gnd.n1668 gnd.n1667 0.152939
R21378 gnd.n1669 gnd.n1668 0.152939
R21379 gnd.n1670 gnd.n1669 0.152939
R21380 gnd.n1671 gnd.n1670 0.152939
R21381 gnd.n1672 gnd.n1671 0.152939
R21382 gnd.n1673 gnd.n1672 0.152939
R21383 gnd.n1674 gnd.n1673 0.152939
R21384 gnd.n1674 gnd.n1372 0.152939
R21385 gnd.n1797 gnd.n1372 0.152939
R21386 gnd.n1798 gnd.n1797 0.152939
R21387 gnd.n1799 gnd.n1798 0.152939
R21388 gnd.n1800 gnd.n1799 0.152939
R21389 gnd.n1800 gnd.n1335 0.152939
R21390 gnd.n1845 gnd.n1335 0.152939
R21391 gnd.n1547 gnd.n1546 0.152939
R21392 gnd.n1548 gnd.n1547 0.152939
R21393 gnd.n1549 gnd.n1548 0.152939
R21394 gnd.n1550 gnd.n1549 0.152939
R21395 gnd.n1551 gnd.n1550 0.152939
R21396 gnd.n1552 gnd.n1551 0.152939
R21397 gnd.n1553 gnd.n1552 0.152939
R21398 gnd.n1554 gnd.n1553 0.152939
R21399 gnd.n1555 gnd.n1554 0.152939
R21400 gnd.n1556 gnd.n1555 0.152939
R21401 gnd.n1557 gnd.n1556 0.152939
R21402 gnd.n1558 gnd.n1557 0.152939
R21403 gnd.n1559 gnd.n1558 0.152939
R21404 gnd.n1560 gnd.n1559 0.152939
R21405 gnd.n1561 gnd.n1560 0.152939
R21406 gnd.n1562 gnd.n1561 0.152939
R21407 gnd.n1563 gnd.n1562 0.152939
R21408 gnd.n1564 gnd.n1563 0.152939
R21409 gnd.n1565 gnd.n1564 0.152939
R21410 gnd.n1566 gnd.n1565 0.152939
R21411 gnd.n1567 gnd.n1566 0.152939
R21412 gnd.n1568 gnd.n1567 0.152939
R21413 gnd.n1572 gnd.n1568 0.152939
R21414 gnd.n1573 gnd.n1572 0.152939
R21415 gnd.n1573 gnd.n1530 0.152939
R21416 gnd.n1627 gnd.n1530 0.152939
R21417 gnd.n7010 gnd.n783 0.152939
R21418 gnd.n7011 gnd.n7010 0.152939
R21419 gnd.n7012 gnd.n7011 0.152939
R21420 gnd.n7012 gnd.n777 0.152939
R21421 gnd.n7020 gnd.n777 0.152939
R21422 gnd.n7021 gnd.n7020 0.152939
R21423 gnd.n7022 gnd.n7021 0.152939
R21424 gnd.n7022 gnd.n771 0.152939
R21425 gnd.n7030 gnd.n771 0.152939
R21426 gnd.n7031 gnd.n7030 0.152939
R21427 gnd.n7032 gnd.n7031 0.152939
R21428 gnd.n7032 gnd.n765 0.152939
R21429 gnd.n7040 gnd.n765 0.152939
R21430 gnd.n7041 gnd.n7040 0.152939
R21431 gnd.n7042 gnd.n7041 0.152939
R21432 gnd.n7042 gnd.n759 0.152939
R21433 gnd.n7050 gnd.n759 0.152939
R21434 gnd.n7051 gnd.n7050 0.152939
R21435 gnd.n7052 gnd.n7051 0.152939
R21436 gnd.n7052 gnd.n753 0.152939
R21437 gnd.n7060 gnd.n753 0.152939
R21438 gnd.n7061 gnd.n7060 0.152939
R21439 gnd.n7062 gnd.n7061 0.152939
R21440 gnd.n7062 gnd.n747 0.152939
R21441 gnd.n7070 gnd.n747 0.152939
R21442 gnd.n7071 gnd.n7070 0.152939
R21443 gnd.n7072 gnd.n7071 0.152939
R21444 gnd.n7072 gnd.n741 0.152939
R21445 gnd.n7080 gnd.n741 0.152939
R21446 gnd.n7081 gnd.n7080 0.152939
R21447 gnd.n7082 gnd.n7081 0.152939
R21448 gnd.n7082 gnd.n735 0.152939
R21449 gnd.n7090 gnd.n735 0.152939
R21450 gnd.n7091 gnd.n7090 0.152939
R21451 gnd.n7092 gnd.n7091 0.152939
R21452 gnd.n7092 gnd.n729 0.152939
R21453 gnd.n7100 gnd.n729 0.152939
R21454 gnd.n7101 gnd.n7100 0.152939
R21455 gnd.n7102 gnd.n7101 0.152939
R21456 gnd.n7102 gnd.n723 0.152939
R21457 gnd.n7110 gnd.n723 0.152939
R21458 gnd.n7111 gnd.n7110 0.152939
R21459 gnd.n7112 gnd.n7111 0.152939
R21460 gnd.n7112 gnd.n717 0.152939
R21461 gnd.n7120 gnd.n717 0.152939
R21462 gnd.n7121 gnd.n7120 0.152939
R21463 gnd.n7122 gnd.n7121 0.152939
R21464 gnd.n7122 gnd.n711 0.152939
R21465 gnd.n7130 gnd.n711 0.152939
R21466 gnd.n7131 gnd.n7130 0.152939
R21467 gnd.n7132 gnd.n7131 0.152939
R21468 gnd.n7132 gnd.n705 0.152939
R21469 gnd.n7140 gnd.n705 0.152939
R21470 gnd.n7141 gnd.n7140 0.152939
R21471 gnd.n7142 gnd.n7141 0.152939
R21472 gnd.n7142 gnd.n699 0.152939
R21473 gnd.n7150 gnd.n699 0.152939
R21474 gnd.n7151 gnd.n7150 0.152939
R21475 gnd.n7152 gnd.n7151 0.152939
R21476 gnd.n7152 gnd.n693 0.152939
R21477 gnd.n7160 gnd.n693 0.152939
R21478 gnd.n7161 gnd.n7160 0.152939
R21479 gnd.n7162 gnd.n7161 0.152939
R21480 gnd.n7162 gnd.n687 0.152939
R21481 gnd.n7170 gnd.n687 0.152939
R21482 gnd.n7171 gnd.n7170 0.152939
R21483 gnd.n7172 gnd.n7171 0.152939
R21484 gnd.n7172 gnd.n681 0.152939
R21485 gnd.n7180 gnd.n681 0.152939
R21486 gnd.n7181 gnd.n7180 0.152939
R21487 gnd.n7182 gnd.n7181 0.152939
R21488 gnd.n7182 gnd.n675 0.152939
R21489 gnd.n7190 gnd.n675 0.152939
R21490 gnd.n7191 gnd.n7190 0.152939
R21491 gnd.n7192 gnd.n7191 0.152939
R21492 gnd.n7192 gnd.n669 0.152939
R21493 gnd.n7200 gnd.n669 0.152939
R21494 gnd.n7201 gnd.n7200 0.152939
R21495 gnd.n7202 gnd.n7201 0.152939
R21496 gnd.n7202 gnd.n663 0.152939
R21497 gnd.n7210 gnd.n663 0.152939
R21498 gnd.n7211 gnd.n7210 0.152939
R21499 gnd.n7212 gnd.n7211 0.152939
R21500 gnd.n7212 gnd.n657 0.152939
R21501 gnd.n7220 gnd.n657 0.152939
R21502 gnd.n7221 gnd.n7220 0.152939
R21503 gnd.n7222 gnd.n7221 0.152939
R21504 gnd.n7222 gnd.n651 0.152939
R21505 gnd.n7230 gnd.n651 0.152939
R21506 gnd.n7231 gnd.n7230 0.152939
R21507 gnd.n7232 gnd.n7231 0.152939
R21508 gnd.n7232 gnd.n645 0.152939
R21509 gnd.n7240 gnd.n645 0.152939
R21510 gnd.n7241 gnd.n7240 0.152939
R21511 gnd.n7242 gnd.n7241 0.152939
R21512 gnd.n7242 gnd.n639 0.152939
R21513 gnd.n7250 gnd.n639 0.152939
R21514 gnd.n7251 gnd.n7250 0.152939
R21515 gnd.n7252 gnd.n7251 0.152939
R21516 gnd.n7252 gnd.n633 0.152939
R21517 gnd.n7260 gnd.n633 0.152939
R21518 gnd.n7261 gnd.n7260 0.152939
R21519 gnd.n7262 gnd.n7261 0.152939
R21520 gnd.n7262 gnd.n627 0.152939
R21521 gnd.n7270 gnd.n627 0.152939
R21522 gnd.n7271 gnd.n7270 0.152939
R21523 gnd.n7272 gnd.n7271 0.152939
R21524 gnd.n7272 gnd.n621 0.152939
R21525 gnd.n7280 gnd.n621 0.152939
R21526 gnd.n7281 gnd.n7280 0.152939
R21527 gnd.n7282 gnd.n7281 0.152939
R21528 gnd.n7282 gnd.n615 0.152939
R21529 gnd.n7290 gnd.n615 0.152939
R21530 gnd.n7291 gnd.n7290 0.152939
R21531 gnd.n7292 gnd.n7291 0.152939
R21532 gnd.n7292 gnd.n609 0.152939
R21533 gnd.n7300 gnd.n609 0.152939
R21534 gnd.n7301 gnd.n7300 0.152939
R21535 gnd.n7302 gnd.n7301 0.152939
R21536 gnd.n7302 gnd.n603 0.152939
R21537 gnd.n7310 gnd.n603 0.152939
R21538 gnd.n7311 gnd.n7310 0.152939
R21539 gnd.n7312 gnd.n7311 0.152939
R21540 gnd.n7312 gnd.n597 0.152939
R21541 gnd.n7320 gnd.n597 0.152939
R21542 gnd.n7321 gnd.n7320 0.152939
R21543 gnd.n7322 gnd.n7321 0.152939
R21544 gnd.n7322 gnd.n591 0.152939
R21545 gnd.n7330 gnd.n591 0.152939
R21546 gnd.n7331 gnd.n7330 0.152939
R21547 gnd.n7332 gnd.n7331 0.152939
R21548 gnd.n7332 gnd.n585 0.152939
R21549 gnd.n7340 gnd.n585 0.152939
R21550 gnd.n7341 gnd.n7340 0.152939
R21551 gnd.n7342 gnd.n7341 0.152939
R21552 gnd.n7342 gnd.n579 0.152939
R21553 gnd.n7350 gnd.n579 0.152939
R21554 gnd.n7351 gnd.n7350 0.152939
R21555 gnd.n7352 gnd.n7351 0.152939
R21556 gnd.n7352 gnd.n573 0.152939
R21557 gnd.n7360 gnd.n573 0.152939
R21558 gnd.n7361 gnd.n7360 0.152939
R21559 gnd.n7362 gnd.n7361 0.152939
R21560 gnd.n7362 gnd.n567 0.152939
R21561 gnd.n7370 gnd.n567 0.152939
R21562 gnd.n7371 gnd.n7370 0.152939
R21563 gnd.n7372 gnd.n7371 0.152939
R21564 gnd.n7372 gnd.n561 0.152939
R21565 gnd.n7380 gnd.n561 0.152939
R21566 gnd.n7381 gnd.n7380 0.152939
R21567 gnd.n7382 gnd.n7381 0.152939
R21568 gnd.n7382 gnd.n555 0.152939
R21569 gnd.n7390 gnd.n555 0.152939
R21570 gnd.n7391 gnd.n7390 0.152939
R21571 gnd.n7392 gnd.n7391 0.152939
R21572 gnd.n7392 gnd.n549 0.152939
R21573 gnd.n7400 gnd.n549 0.152939
R21574 gnd.n7401 gnd.n7400 0.152939
R21575 gnd.n7402 gnd.n7401 0.152939
R21576 gnd.n7402 gnd.n543 0.152939
R21577 gnd.n7410 gnd.n543 0.152939
R21578 gnd.n7411 gnd.n7410 0.152939
R21579 gnd.n7412 gnd.n7411 0.152939
R21580 gnd.n7412 gnd.n537 0.152939
R21581 gnd.n7420 gnd.n537 0.152939
R21582 gnd.n7421 gnd.n7420 0.152939
R21583 gnd.n7422 gnd.n7421 0.152939
R21584 gnd.n7422 gnd.n531 0.152939
R21585 gnd.n7430 gnd.n531 0.152939
R21586 gnd.n7431 gnd.n7430 0.152939
R21587 gnd.n7432 gnd.n7431 0.152939
R21588 gnd.n7432 gnd.n525 0.152939
R21589 gnd.n7440 gnd.n525 0.152939
R21590 gnd.n7441 gnd.n7440 0.152939
R21591 gnd.n7442 gnd.n7441 0.152939
R21592 gnd.n7442 gnd.n519 0.152939
R21593 gnd.n7450 gnd.n519 0.152939
R21594 gnd.n7451 gnd.n7450 0.152939
R21595 gnd.n7452 gnd.n7451 0.152939
R21596 gnd.n7452 gnd.n513 0.152939
R21597 gnd.n7460 gnd.n513 0.152939
R21598 gnd.n7461 gnd.n7460 0.152939
R21599 gnd.n7462 gnd.n7461 0.152939
R21600 gnd.n7462 gnd.n507 0.152939
R21601 gnd.n7470 gnd.n507 0.152939
R21602 gnd.n7471 gnd.n7470 0.152939
R21603 gnd.n7472 gnd.n7471 0.152939
R21604 gnd.n7472 gnd.n501 0.152939
R21605 gnd.n7480 gnd.n501 0.152939
R21606 gnd.n7481 gnd.n7480 0.152939
R21607 gnd.n7483 gnd.n7481 0.152939
R21608 gnd.n7483 gnd.n7482 0.152939
R21609 gnd.n7482 gnd.n495 0.152939
R21610 gnd.n7492 gnd.n495 0.152939
R21611 gnd.n7493 gnd.n490 0.152939
R21612 gnd.n7501 gnd.n490 0.152939
R21613 gnd.n7502 gnd.n7501 0.152939
R21614 gnd.n7503 gnd.n7502 0.152939
R21615 gnd.n7503 gnd.n484 0.152939
R21616 gnd.n7511 gnd.n484 0.152939
R21617 gnd.n7512 gnd.n7511 0.152939
R21618 gnd.n7513 gnd.n7512 0.152939
R21619 gnd.n7513 gnd.n478 0.152939
R21620 gnd.n7521 gnd.n478 0.152939
R21621 gnd.n7522 gnd.n7521 0.152939
R21622 gnd.n7523 gnd.n7522 0.152939
R21623 gnd.n7523 gnd.n472 0.152939
R21624 gnd.n7531 gnd.n472 0.152939
R21625 gnd.n7532 gnd.n7531 0.152939
R21626 gnd.n7533 gnd.n7532 0.152939
R21627 gnd.n7533 gnd.n466 0.152939
R21628 gnd.n7541 gnd.n466 0.152939
R21629 gnd.n7542 gnd.n7541 0.152939
R21630 gnd.n7543 gnd.n7542 0.152939
R21631 gnd.n7543 gnd.n460 0.152939
R21632 gnd.n7551 gnd.n460 0.152939
R21633 gnd.n7552 gnd.n7551 0.152939
R21634 gnd.n7553 gnd.n7552 0.152939
R21635 gnd.n7553 gnd.n454 0.152939
R21636 gnd.n7561 gnd.n454 0.152939
R21637 gnd.n7562 gnd.n7561 0.152939
R21638 gnd.n7563 gnd.n7562 0.152939
R21639 gnd.n7563 gnd.n448 0.152939
R21640 gnd.n7571 gnd.n448 0.152939
R21641 gnd.n7572 gnd.n7571 0.152939
R21642 gnd.n7573 gnd.n7572 0.152939
R21643 gnd.n7573 gnd.n442 0.152939
R21644 gnd.n7581 gnd.n442 0.152939
R21645 gnd.n7582 gnd.n7581 0.152939
R21646 gnd.n7583 gnd.n7582 0.152939
R21647 gnd.n7583 gnd.n436 0.152939
R21648 gnd.n7591 gnd.n436 0.152939
R21649 gnd.n7592 gnd.n7591 0.152939
R21650 gnd.n7593 gnd.n7592 0.152939
R21651 gnd.n7593 gnd.n430 0.152939
R21652 gnd.n7601 gnd.n430 0.152939
R21653 gnd.n7602 gnd.n7601 0.152939
R21654 gnd.n7603 gnd.n7602 0.152939
R21655 gnd.n7603 gnd.n424 0.152939
R21656 gnd.n7611 gnd.n424 0.152939
R21657 gnd.n7612 gnd.n7611 0.152939
R21658 gnd.n7613 gnd.n7612 0.152939
R21659 gnd.n7613 gnd.n418 0.152939
R21660 gnd.n7621 gnd.n418 0.152939
R21661 gnd.n7622 gnd.n7621 0.152939
R21662 gnd.n7623 gnd.n7622 0.152939
R21663 gnd.n7623 gnd.n412 0.152939
R21664 gnd.n7631 gnd.n412 0.152939
R21665 gnd.n7632 gnd.n7631 0.152939
R21666 gnd.n7633 gnd.n7632 0.152939
R21667 gnd.n7633 gnd.n406 0.152939
R21668 gnd.n7641 gnd.n406 0.152939
R21669 gnd.n7642 gnd.n7641 0.152939
R21670 gnd.n7643 gnd.n7642 0.152939
R21671 gnd.n7643 gnd.n400 0.152939
R21672 gnd.n7651 gnd.n400 0.152939
R21673 gnd.n7652 gnd.n7651 0.152939
R21674 gnd.n7653 gnd.n7652 0.152939
R21675 gnd.n7653 gnd.n394 0.152939
R21676 gnd.n7661 gnd.n394 0.152939
R21677 gnd.n7662 gnd.n7661 0.152939
R21678 gnd.n7663 gnd.n7662 0.152939
R21679 gnd.n7663 gnd.n388 0.152939
R21680 gnd.n7671 gnd.n388 0.152939
R21681 gnd.n7672 gnd.n7671 0.152939
R21682 gnd.n7673 gnd.n7672 0.152939
R21683 gnd.n7673 gnd.n382 0.152939
R21684 gnd.n7681 gnd.n382 0.152939
R21685 gnd.n7682 gnd.n7681 0.152939
R21686 gnd.n7683 gnd.n7682 0.152939
R21687 gnd.n7683 gnd.n376 0.152939
R21688 gnd.n7691 gnd.n376 0.152939
R21689 gnd.n7692 gnd.n7691 0.152939
R21690 gnd.n7693 gnd.n7692 0.152939
R21691 gnd.n7693 gnd.n370 0.152939
R21692 gnd.n7702 gnd.n370 0.152939
R21693 gnd.n7703 gnd.n7702 0.152939
R21694 gnd.n7705 gnd.n7703 0.152939
R21695 gnd.n5846 gnd.n5823 0.152939
R21696 gnd.n5848 gnd.n5846 0.152939
R21697 gnd.n5849 gnd.n5848 0.152939
R21698 gnd.n5850 gnd.n5849 0.152939
R21699 gnd.n5851 gnd.n5850 0.152939
R21700 gnd.n5852 gnd.n5851 0.152939
R21701 gnd.n5854 gnd.n5852 0.152939
R21702 gnd.n5854 gnd.n5853 0.152939
R21703 gnd.n5853 gnd.n364 0.152939
R21704 gnd.n365 gnd.n364 0.152939
R21705 gnd.n366 gnd.n365 0.152939
R21706 gnd.n7704 gnd.n366 0.152939
R21707 gnd.n8062 gnd.n109 0.152939
R21708 gnd.n134 gnd.n109 0.152939
R21709 gnd.n135 gnd.n134 0.152939
R21710 gnd.n136 gnd.n135 0.152939
R21711 gnd.n153 gnd.n136 0.152939
R21712 gnd.n154 gnd.n153 0.152939
R21713 gnd.n155 gnd.n154 0.152939
R21714 gnd.n156 gnd.n155 0.152939
R21715 gnd.n173 gnd.n156 0.152939
R21716 gnd.n174 gnd.n173 0.152939
R21717 gnd.n175 gnd.n174 0.152939
R21718 gnd.n176 gnd.n175 0.152939
R21719 gnd.n193 gnd.n176 0.152939
R21720 gnd.n194 gnd.n193 0.152939
R21721 gnd.n195 gnd.n194 0.152939
R21722 gnd.n196 gnd.n195 0.152939
R21723 gnd.n213 gnd.n196 0.152939
R21724 gnd.n214 gnd.n213 0.152939
R21725 gnd.n215 gnd.n214 0.152939
R21726 gnd.n216 gnd.n215 0.152939
R21727 gnd.n232 gnd.n216 0.152939
R21728 gnd.n233 gnd.n232 0.152939
R21729 gnd.n234 gnd.n233 0.152939
R21730 gnd.n235 gnd.n234 0.152939
R21731 gnd.n251 gnd.n235 0.152939
R21732 gnd.n252 gnd.n251 0.152939
R21733 gnd.n7977 gnd.n252 0.152939
R21734 gnd.n8071 gnd.n97 0.152939
R21735 gnd.n5828 gnd.n97 0.152939
R21736 gnd.n5832 gnd.n5828 0.152939
R21737 gnd.n5833 gnd.n5832 0.152939
R21738 gnd.n5834 gnd.n5833 0.152939
R21739 gnd.n5835 gnd.n5834 0.152939
R21740 gnd.n5836 gnd.n5835 0.152939
R21741 gnd.n5863 gnd.n5836 0.152939
R21742 gnd.n5864 gnd.n5863 0.152939
R21743 gnd.n5865 gnd.n5864 0.152939
R21744 gnd.n5866 gnd.n5865 0.152939
R21745 gnd.n5866 gnd.n358 0.152939
R21746 gnd.n7719 gnd.n358 0.152939
R21747 gnd.n7720 gnd.n7719 0.152939
R21748 gnd.n7721 gnd.n7720 0.152939
R21749 gnd.n7722 gnd.n7721 0.152939
R21750 gnd.n7723 gnd.n7722 0.152939
R21751 gnd.n7724 gnd.n7723 0.152939
R21752 gnd.n7725 gnd.n7724 0.152939
R21753 gnd.n7726 gnd.n7725 0.152939
R21754 gnd.n7727 gnd.n7726 0.152939
R21755 gnd.n7728 gnd.n7727 0.152939
R21756 gnd.n7729 gnd.n7728 0.152939
R21757 gnd.n7730 gnd.n7729 0.152939
R21758 gnd.n7731 gnd.n7730 0.152939
R21759 gnd.n7732 gnd.n7731 0.152939
R21760 gnd.n7733 gnd.n7732 0.152939
R21761 gnd.n7734 gnd.n7733 0.152939
R21762 gnd.n7735 gnd.n7734 0.152939
R21763 gnd.n7736 gnd.n7735 0.152939
R21764 gnd.n7737 gnd.n7736 0.152939
R21765 gnd.n7751 gnd.n354 0.152939
R21766 gnd.n7752 gnd.n7751 0.152939
R21767 gnd.n7752 gnd.n7747 0.152939
R21768 gnd.n7760 gnd.n7747 0.152939
R21769 gnd.n7761 gnd.n7760 0.152939
R21770 gnd.n7762 gnd.n7761 0.152939
R21771 gnd.n7762 gnd.n7745 0.152939
R21772 gnd.n7770 gnd.n7745 0.152939
R21773 gnd.n7771 gnd.n7770 0.152939
R21774 gnd.n7772 gnd.n7771 0.152939
R21775 gnd.n7772 gnd.n7743 0.152939
R21776 gnd.n7780 gnd.n7743 0.152939
R21777 gnd.n7781 gnd.n7780 0.152939
R21778 gnd.n7782 gnd.n7781 0.152939
R21779 gnd.n7782 gnd.n7741 0.152939
R21780 gnd.n7790 gnd.n7741 0.152939
R21781 gnd.n7791 gnd.n7790 0.152939
R21782 gnd.n7792 gnd.n7791 0.152939
R21783 gnd.n7976 gnd.n253 0.152939
R21784 gnd.n296 gnd.n253 0.152939
R21785 gnd.n297 gnd.n296 0.152939
R21786 gnd.n298 gnd.n297 0.152939
R21787 gnd.n299 gnd.n298 0.152939
R21788 gnd.n300 gnd.n299 0.152939
R21789 gnd.n301 gnd.n300 0.152939
R21790 gnd.n302 gnd.n301 0.152939
R21791 gnd.n303 gnd.n302 0.152939
R21792 gnd.n304 gnd.n303 0.152939
R21793 gnd.n305 gnd.n304 0.152939
R21794 gnd.n306 gnd.n305 0.152939
R21795 gnd.n307 gnd.n306 0.152939
R21796 gnd.n308 gnd.n307 0.152939
R21797 gnd.n309 gnd.n308 0.152939
R21798 gnd.n310 gnd.n309 0.152939
R21799 gnd.n311 gnd.n310 0.152939
R21800 gnd.n312 gnd.n311 0.152939
R21801 gnd.n313 gnd.n312 0.152939
R21802 gnd.n314 gnd.n313 0.152939
R21803 gnd.n315 gnd.n314 0.152939
R21804 gnd.n316 gnd.n315 0.152939
R21805 gnd.n317 gnd.n316 0.152939
R21806 gnd.n318 gnd.n317 0.152939
R21807 gnd.n319 gnd.n318 0.152939
R21808 gnd.n320 gnd.n319 0.152939
R21809 gnd.n321 gnd.n320 0.152939
R21810 gnd.n322 gnd.n321 0.152939
R21811 gnd.n323 gnd.n322 0.152939
R21812 gnd.n324 gnd.n323 0.152939
R21813 gnd.n325 gnd.n324 0.152939
R21814 gnd.n326 gnd.n325 0.152939
R21815 gnd.n327 gnd.n326 0.152939
R21816 gnd.n328 gnd.n327 0.152939
R21817 gnd.n329 gnd.n328 0.152939
R21818 gnd.n330 gnd.n329 0.152939
R21819 gnd.n7897 gnd.n330 0.152939
R21820 gnd.n7897 gnd.n7896 0.152939
R21821 gnd.n7896 gnd.n7895 0.152939
R21822 gnd.n7895 gnd.n334 0.152939
R21823 gnd.n335 gnd.n334 0.152939
R21824 gnd.n336 gnd.n335 0.152939
R21825 gnd.n337 gnd.n336 0.152939
R21826 gnd.n338 gnd.n337 0.152939
R21827 gnd.n339 gnd.n338 0.152939
R21828 gnd.n340 gnd.n339 0.152939
R21829 gnd.n341 gnd.n340 0.152939
R21830 gnd.n342 gnd.n341 0.152939
R21831 gnd.n343 gnd.n342 0.152939
R21832 gnd.n344 gnd.n343 0.152939
R21833 gnd.n345 gnd.n344 0.152939
R21834 gnd.n346 gnd.n345 0.152939
R21835 gnd.n347 gnd.n346 0.152939
R21836 gnd.n348 gnd.n347 0.152939
R21837 gnd.n349 gnd.n348 0.152939
R21838 gnd.n350 gnd.n349 0.152939
R21839 gnd.n7855 gnd.n350 0.152939
R21840 gnd.n7855 gnd.n7854 0.152939
R21841 gnd.n3122 gnd.n3121 0.152939
R21842 gnd.n3123 gnd.n3122 0.152939
R21843 gnd.n3124 gnd.n3123 0.152939
R21844 gnd.n3125 gnd.n3124 0.152939
R21845 gnd.n3126 gnd.n3125 0.152939
R21846 gnd.n3127 gnd.n3126 0.152939
R21847 gnd.n3128 gnd.n3127 0.152939
R21848 gnd.n3129 gnd.n3128 0.152939
R21849 gnd.n3130 gnd.n3129 0.152939
R21850 gnd.n3131 gnd.n3130 0.152939
R21851 gnd.n3132 gnd.n3131 0.152939
R21852 gnd.n3133 gnd.n3132 0.152939
R21853 gnd.n3134 gnd.n3133 0.152939
R21854 gnd.n3135 gnd.n3134 0.152939
R21855 gnd.n3136 gnd.n3135 0.152939
R21856 gnd.n3137 gnd.n3136 0.152939
R21857 gnd.n3138 gnd.n3137 0.152939
R21858 gnd.n3141 gnd.n3138 0.152939
R21859 gnd.n3142 gnd.n3141 0.152939
R21860 gnd.n3143 gnd.n3142 0.152939
R21861 gnd.n3144 gnd.n3143 0.152939
R21862 gnd.n3145 gnd.n3144 0.152939
R21863 gnd.n3146 gnd.n3145 0.152939
R21864 gnd.n3147 gnd.n3146 0.152939
R21865 gnd.n3148 gnd.n3147 0.152939
R21866 gnd.n3153 gnd.n3152 0.152939
R21867 gnd.n3154 gnd.n3153 0.152939
R21868 gnd.n3155 gnd.n3154 0.152939
R21869 gnd.n3156 gnd.n3155 0.152939
R21870 gnd.n3157 gnd.n3156 0.152939
R21871 gnd.n3158 gnd.n3157 0.152939
R21872 gnd.n3159 gnd.n3158 0.152939
R21873 gnd.n3160 gnd.n3159 0.152939
R21874 gnd.n3161 gnd.n3160 0.152939
R21875 gnd.n3164 gnd.n3161 0.152939
R21876 gnd.n3165 gnd.n3164 0.152939
R21877 gnd.n3166 gnd.n3165 0.152939
R21878 gnd.n3167 gnd.n3166 0.152939
R21879 gnd.n3168 gnd.n3167 0.152939
R21880 gnd.n3169 gnd.n3168 0.152939
R21881 gnd.n3170 gnd.n3169 0.152939
R21882 gnd.n3171 gnd.n3170 0.152939
R21883 gnd.n3172 gnd.n3171 0.152939
R21884 gnd.n3173 gnd.n3172 0.152939
R21885 gnd.n3174 gnd.n3173 0.152939
R21886 gnd.n3175 gnd.n3174 0.152939
R21887 gnd.n3176 gnd.n3175 0.152939
R21888 gnd.n3177 gnd.n3176 0.152939
R21889 gnd.n3178 gnd.n3177 0.152939
R21890 gnd.n3179 gnd.n3178 0.152939
R21891 gnd.n3180 gnd.n3179 0.152939
R21892 gnd.n3181 gnd.n3180 0.152939
R21893 gnd.n3182 gnd.n3181 0.152939
R21894 gnd.n6020 gnd.n3182 0.152939
R21895 gnd.n6020 gnd.n6019 0.152939
R21896 gnd.n3203 gnd.n3202 0.152939
R21897 gnd.n3204 gnd.n3203 0.152939
R21898 gnd.n3205 gnd.n3204 0.152939
R21899 gnd.n3206 gnd.n3205 0.152939
R21900 gnd.n3227 gnd.n3206 0.152939
R21901 gnd.n3228 gnd.n3227 0.152939
R21902 gnd.n3229 gnd.n3228 0.152939
R21903 gnd.n3230 gnd.n3229 0.152939
R21904 gnd.n3248 gnd.n3230 0.152939
R21905 gnd.n3249 gnd.n3248 0.152939
R21906 gnd.n3250 gnd.n3249 0.152939
R21907 gnd.n3251 gnd.n3250 0.152939
R21908 gnd.n3268 gnd.n3251 0.152939
R21909 gnd.n3269 gnd.n3268 0.152939
R21910 gnd.n3270 gnd.n3269 0.152939
R21911 gnd.n3271 gnd.n3270 0.152939
R21912 gnd.n3289 gnd.n3271 0.152939
R21913 gnd.n3290 gnd.n3289 0.152939
R21914 gnd.n3291 gnd.n3290 0.152939
R21915 gnd.n3292 gnd.n3291 0.152939
R21916 gnd.n3309 gnd.n3292 0.152939
R21917 gnd.n3310 gnd.n3309 0.152939
R21918 gnd.n3311 gnd.n3310 0.152939
R21919 gnd.n3312 gnd.n3311 0.152939
R21920 gnd.n3313 gnd.n3312 0.152939
R21921 gnd.n3313 gnd.n110 0.152939
R21922 gnd.n8062 gnd.n110 0.152939
R21923 gnd.n4352 gnd.n4351 0.152939
R21924 gnd.n4353 gnd.n4352 0.152939
R21925 gnd.n4354 gnd.n4353 0.152939
R21926 gnd.n4357 gnd.n4354 0.152939
R21927 gnd.n4358 gnd.n4357 0.152939
R21928 gnd.n4359 gnd.n4358 0.152939
R21929 gnd.n4360 gnd.n4359 0.152939
R21930 gnd.n4362 gnd.n4360 0.152939
R21931 gnd.n4362 gnd.n4361 0.152939
R21932 gnd.n4361 gnd.n3987 0.152939
R21933 gnd.n4439 gnd.n3987 0.152939
R21934 gnd.n4440 gnd.n4439 0.152939
R21935 gnd.n4441 gnd.n4440 0.152939
R21936 gnd.n4441 gnd.n3983 0.152939
R21937 gnd.n4447 gnd.n3983 0.152939
R21938 gnd.n4448 gnd.n4447 0.152939
R21939 gnd.n4449 gnd.n4448 0.152939
R21940 gnd.n4450 gnd.n4449 0.152939
R21941 gnd.n4451 gnd.n4450 0.152939
R21942 gnd.n4451 gnd.n3965 0.152939
R21943 gnd.n4742 gnd.n3965 0.152939
R21944 gnd.n4743 gnd.n4742 0.152939
R21945 gnd.n4744 gnd.n4743 0.152939
R21946 gnd.n4744 gnd.n3961 0.152939
R21947 gnd.n4750 gnd.n3961 0.152939
R21948 gnd.n4751 gnd.n4750 0.152939
R21949 gnd.n4752 gnd.n4751 0.152939
R21950 gnd.n4753 gnd.n4752 0.152939
R21951 gnd.n4754 gnd.n4753 0.152939
R21952 gnd.n4755 gnd.n4754 0.152939
R21953 gnd.n4755 gnd.n3931 0.152939
R21954 gnd.n4778 gnd.n3931 0.152939
R21955 gnd.n4779 gnd.n4778 0.152939
R21956 gnd.n4780 gnd.n4779 0.152939
R21957 gnd.n4780 gnd.n3915 0.152939
R21958 gnd.n4811 gnd.n3915 0.152939
R21959 gnd.n4812 gnd.n4811 0.152939
R21960 gnd.n4813 gnd.n4812 0.152939
R21961 gnd.n4814 gnd.n4813 0.152939
R21962 gnd.n4815 gnd.n4814 0.152939
R21963 gnd.n4817 gnd.n4815 0.152939
R21964 gnd.n4817 gnd.n4816 0.152939
R21965 gnd.n4816 gnd.n2906 0.152939
R21966 gnd.n2907 gnd.n2906 0.152939
R21967 gnd.n2908 gnd.n2907 0.152939
R21968 gnd.n5007 gnd.n2908 0.152939
R21969 gnd.n5008 gnd.n5007 0.152939
R21970 gnd.n5009 gnd.n5008 0.152939
R21971 gnd.n5009 gnd.n3804 0.152939
R21972 gnd.n5036 gnd.n3804 0.152939
R21973 gnd.n5037 gnd.n5036 0.152939
R21974 gnd.n5038 gnd.n5037 0.152939
R21975 gnd.n5039 gnd.n5038 0.152939
R21976 gnd.n5040 gnd.n5039 0.152939
R21977 gnd.n5042 gnd.n5040 0.152939
R21978 gnd.n5043 gnd.n5042 0.152939
R21979 gnd.n5043 gnd.n3766 0.152939
R21980 gnd.n5094 gnd.n3766 0.152939
R21981 gnd.n5095 gnd.n5094 0.152939
R21982 gnd.n5096 gnd.n5095 0.152939
R21983 gnd.n5096 gnd.n3748 0.152939
R21984 gnd.n5120 gnd.n3748 0.152939
R21985 gnd.n5121 gnd.n5120 0.152939
R21986 gnd.n5122 gnd.n5121 0.152939
R21987 gnd.n5123 gnd.n5122 0.152939
R21988 gnd.n5123 gnd.n3724 0.152939
R21989 gnd.n5159 gnd.n3724 0.152939
R21990 gnd.n5160 gnd.n5159 0.152939
R21991 gnd.n5161 gnd.n5160 0.152939
R21992 gnd.n5162 gnd.n5161 0.152939
R21993 gnd.n5163 gnd.n5162 0.152939
R21994 gnd.n5165 gnd.n5163 0.152939
R21995 gnd.n5166 gnd.n5165 0.152939
R21996 gnd.n5166 gnd.n3685 0.152939
R21997 gnd.n5217 gnd.n3685 0.152939
R21998 gnd.n5218 gnd.n5217 0.152939
R21999 gnd.n5219 gnd.n5218 0.152939
R22000 gnd.n5219 gnd.n3666 0.152939
R22001 gnd.n5242 gnd.n3666 0.152939
R22002 gnd.n5243 gnd.n5242 0.152939
R22003 gnd.n5244 gnd.n5243 0.152939
R22004 gnd.n5245 gnd.n5244 0.152939
R22005 gnd.n5245 gnd.n3641 0.152939
R22006 gnd.n5280 gnd.n3641 0.152939
R22007 gnd.n5281 gnd.n5280 0.152939
R22008 gnd.n5282 gnd.n5281 0.152939
R22009 gnd.n5283 gnd.n5282 0.152939
R22010 gnd.n5284 gnd.n5283 0.152939
R22011 gnd.n5285 gnd.n5284 0.152939
R22012 gnd.n5285 gnd.n3607 0.152939
R22013 gnd.n5326 gnd.n3607 0.152939
R22014 gnd.n5327 gnd.n5326 0.152939
R22015 gnd.n5328 gnd.n5327 0.152939
R22016 gnd.n5329 gnd.n5328 0.152939
R22017 gnd.n5329 gnd.n3579 0.152939
R22018 gnd.n5361 gnd.n3579 0.152939
R22019 gnd.n5362 gnd.n5361 0.152939
R22020 gnd.n5363 gnd.n5362 0.152939
R22021 gnd.n5363 gnd.n3550 0.152939
R22022 gnd.n5398 gnd.n3550 0.152939
R22023 gnd.n5399 gnd.n5398 0.152939
R22024 gnd.n5400 gnd.n5399 0.152939
R22025 gnd.n5401 gnd.n5400 0.152939
R22026 gnd.n5401 gnd.n3450 0.152939
R22027 gnd.n5548 gnd.n3450 0.152939
R22028 gnd.n5549 gnd.n5548 0.152939
R22029 gnd.n5550 gnd.n5549 0.152939
R22030 gnd.n5550 gnd.n3437 0.152939
R22031 gnd.n5564 gnd.n3437 0.152939
R22032 gnd.n5565 gnd.n5564 0.152939
R22033 gnd.n5566 gnd.n5565 0.152939
R22034 gnd.n5568 gnd.n5566 0.152939
R22035 gnd.n5568 gnd.n5567 0.152939
R22036 gnd.n5567 gnd.n3424 0.152939
R22037 gnd.n5585 gnd.n3424 0.152939
R22038 gnd.n5586 gnd.n5585 0.152939
R22039 gnd.n5587 gnd.n5586 0.152939
R22040 gnd.n5588 gnd.n5587 0.152939
R22041 gnd.n5589 gnd.n5588 0.152939
R22042 gnd.n5592 gnd.n5589 0.152939
R22043 gnd.n5593 gnd.n5592 0.152939
R22044 gnd.n5594 gnd.n5593 0.152939
R22045 gnd.n5595 gnd.n5594 0.152939
R22046 gnd.n5598 gnd.n5595 0.152939
R22047 gnd.n5599 gnd.n5598 0.152939
R22048 gnd.n5600 gnd.n5599 0.152939
R22049 gnd.n5601 gnd.n5600 0.152939
R22050 gnd.n5604 gnd.n5601 0.152939
R22051 gnd.n5605 gnd.n5604 0.152939
R22052 gnd.n5606 gnd.n5605 0.152939
R22053 gnd.n5607 gnd.n5606 0.152939
R22054 gnd.n5610 gnd.n5607 0.152939
R22055 gnd.n5611 gnd.n5610 0.152939
R22056 gnd.n5612 gnd.n5611 0.152939
R22057 gnd.n5613 gnd.n5612 0.152939
R22058 gnd.n5616 gnd.n5613 0.152939
R22059 gnd.n5617 gnd.n5616 0.152939
R22060 gnd.n5618 gnd.n5617 0.152939
R22061 gnd.n5619 gnd.n5618 0.152939
R22062 gnd.n5622 gnd.n5619 0.152939
R22063 gnd.n5623 gnd.n5622 0.152939
R22064 gnd.n5624 gnd.n5623 0.152939
R22065 gnd.n5625 gnd.n5624 0.152939
R22066 gnd.n5628 gnd.n5625 0.152939
R22067 gnd.n5629 gnd.n5628 0.152939
R22068 gnd.n5630 gnd.n5629 0.152939
R22069 gnd.n5632 gnd.n5630 0.152939
R22070 gnd.n5632 gnd.n5631 0.152939
R22071 gnd.n4163 gnd.n4104 0.152939
R22072 gnd.n4169 gnd.n4104 0.152939
R22073 gnd.n4170 gnd.n4169 0.152939
R22074 gnd.n4171 gnd.n4170 0.152939
R22075 gnd.n4171 gnd.n4102 0.152939
R22076 gnd.n4177 gnd.n4102 0.152939
R22077 gnd.n4178 gnd.n4177 0.152939
R22078 gnd.n4179 gnd.n4178 0.152939
R22079 gnd.n4179 gnd.n4100 0.152939
R22080 gnd.n4185 gnd.n4100 0.152939
R22081 gnd.n4186 gnd.n4185 0.152939
R22082 gnd.n4187 gnd.n4186 0.152939
R22083 gnd.n4187 gnd.n4098 0.152939
R22084 gnd.n4193 gnd.n4098 0.152939
R22085 gnd.n4194 gnd.n4193 0.152939
R22086 gnd.n4196 gnd.n4194 0.152939
R22087 gnd.n4196 gnd.n4195 0.152939
R22088 gnd.n4195 gnd.n4070 0.152939
R22089 gnd.n4071 gnd.n4070 0.152939
R22090 gnd.n4072 gnd.n4071 0.152939
R22091 gnd.n4072 gnd.n4061 0.152939
R22092 gnd.n4251 gnd.n4061 0.152939
R22093 gnd.n4252 gnd.n4251 0.152939
R22094 gnd.n4254 gnd.n4252 0.152939
R22095 gnd.n4254 gnd.n4253 0.152939
R22096 gnd.n4253 gnd.n4056 0.152939
R22097 gnd.n4057 gnd.n4056 0.152939
R22098 gnd.n4058 gnd.n4057 0.152939
R22099 gnd.n4058 gnd.n4043 0.152939
R22100 gnd.n4310 gnd.n4043 0.152939
R22101 gnd.n4311 gnd.n4310 0.152939
R22102 gnd.n4118 gnd.n2462 0.152939
R22103 gnd.n4126 gnd.n4118 0.152939
R22104 gnd.n4127 gnd.n4126 0.152939
R22105 gnd.n4128 gnd.n4127 0.152939
R22106 gnd.n4128 gnd.n4116 0.152939
R22107 gnd.n4136 gnd.n4116 0.152939
R22108 gnd.n4137 gnd.n4136 0.152939
R22109 gnd.n4138 gnd.n4137 0.152939
R22110 gnd.n4138 gnd.n4114 0.152939
R22111 gnd.n4146 gnd.n4114 0.152939
R22112 gnd.n4147 gnd.n4146 0.152939
R22113 gnd.n4148 gnd.n4147 0.152939
R22114 gnd.n4148 gnd.n4112 0.152939
R22115 gnd.n4156 gnd.n4112 0.152939
R22116 gnd.n4157 gnd.n4156 0.152939
R22117 gnd.n4158 gnd.n4157 0.152939
R22118 gnd.n4158 gnd.n4105 0.152939
R22119 gnd.n4162 gnd.n4105 0.152939
R22120 gnd.n6533 gnd.n2615 0.152939
R22121 gnd.n2640 gnd.n2615 0.152939
R22122 gnd.n2641 gnd.n2640 0.152939
R22123 gnd.n2642 gnd.n2641 0.152939
R22124 gnd.n2659 gnd.n2642 0.152939
R22125 gnd.n2660 gnd.n2659 0.152939
R22126 gnd.n2661 gnd.n2660 0.152939
R22127 gnd.n2662 gnd.n2661 0.152939
R22128 gnd.n2679 gnd.n2662 0.152939
R22129 gnd.n2680 gnd.n2679 0.152939
R22130 gnd.n2681 gnd.n2680 0.152939
R22131 gnd.n2682 gnd.n2681 0.152939
R22132 gnd.n2699 gnd.n2682 0.152939
R22133 gnd.n2700 gnd.n2699 0.152939
R22134 gnd.n2701 gnd.n2700 0.152939
R22135 gnd.n2702 gnd.n2701 0.152939
R22136 gnd.n2719 gnd.n2702 0.152939
R22137 gnd.n2720 gnd.n2719 0.152939
R22138 gnd.n2721 gnd.n2720 0.152939
R22139 gnd.n2722 gnd.n2721 0.152939
R22140 gnd.n2739 gnd.n2722 0.152939
R22141 gnd.n2740 gnd.n2739 0.152939
R22142 gnd.n2741 gnd.n2740 0.152939
R22143 gnd.n2742 gnd.n2741 0.152939
R22144 gnd.n2760 gnd.n2742 0.152939
R22145 gnd.n2761 gnd.n2760 0.152939
R22146 gnd.n6448 gnd.n2761 0.152939
R22147 gnd.n6447 gnd.n2762 0.152939
R22148 gnd.n2806 gnd.n2762 0.152939
R22149 gnd.n2807 gnd.n2806 0.152939
R22150 gnd.n2808 gnd.n2807 0.152939
R22151 gnd.n2809 gnd.n2808 0.152939
R22152 gnd.n2810 gnd.n2809 0.152939
R22153 gnd.n2811 gnd.n2810 0.152939
R22154 gnd.n2812 gnd.n2811 0.152939
R22155 gnd.n2813 gnd.n2812 0.152939
R22156 gnd.n2814 gnd.n2813 0.152939
R22157 gnd.n2815 gnd.n2814 0.152939
R22158 gnd.n2816 gnd.n2815 0.152939
R22159 gnd.n2817 gnd.n2816 0.152939
R22160 gnd.n2818 gnd.n2817 0.152939
R22161 gnd.n2819 gnd.n2818 0.152939
R22162 gnd.n2820 gnd.n2819 0.152939
R22163 gnd.n2821 gnd.n2820 0.152939
R22164 gnd.n2824 gnd.n2821 0.152939
R22165 gnd.n2825 gnd.n2824 0.152939
R22166 gnd.n2826 gnd.n2825 0.152939
R22167 gnd.n2827 gnd.n2826 0.152939
R22168 gnd.n2828 gnd.n2827 0.152939
R22169 gnd.n2829 gnd.n2828 0.152939
R22170 gnd.n2830 gnd.n2829 0.152939
R22171 gnd.n2831 gnd.n2830 0.152939
R22172 gnd.n4643 gnd.n4642 0.152939
R22173 gnd.n4650 gnd.n4643 0.152939
R22174 gnd.n4651 gnd.n4650 0.152939
R22175 gnd.n4652 gnd.n4651 0.152939
R22176 gnd.n4652 gnd.n4640 0.152939
R22177 gnd.n4660 gnd.n4640 0.152939
R22178 gnd.n4661 gnd.n4660 0.152939
R22179 gnd.n4662 gnd.n4661 0.152939
R22180 gnd.n4662 gnd.n4635 0.152939
R22181 gnd.n4669 gnd.n4635 0.152939
R22182 gnd.n4670 gnd.n4669 0.152939
R22183 gnd.n4671 gnd.n4670 0.152939
R22184 gnd.n4671 gnd.n4633 0.152939
R22185 gnd.n4679 gnd.n4633 0.152939
R22186 gnd.n4680 gnd.n4679 0.152939
R22187 gnd.n4681 gnd.n4680 0.152939
R22188 gnd.n4681 gnd.n4631 0.152939
R22189 gnd.n4689 gnd.n4631 0.152939
R22190 gnd.n4690 gnd.n4689 0.152939
R22191 gnd.n4691 gnd.n4690 0.152939
R22192 gnd.n4691 gnd.n4629 0.152939
R22193 gnd.n4699 gnd.n4629 0.152939
R22194 gnd.n4700 gnd.n4699 0.152939
R22195 gnd.n4701 gnd.n4700 0.152939
R22196 gnd.n4701 gnd.n4627 0.152939
R22197 gnd.n4709 gnd.n4627 0.152939
R22198 gnd.n4710 gnd.n4709 0.152939
R22199 gnd.n4711 gnd.n4710 0.152939
R22200 gnd.n4711 gnd.n4622 0.152939
R22201 gnd.n4717 gnd.n4622 0.152939
R22202 gnd.n2399 gnd.n2398 0.152939
R22203 gnd.n2400 gnd.n2399 0.152939
R22204 gnd.n2401 gnd.n2400 0.152939
R22205 gnd.n2402 gnd.n2401 0.152939
R22206 gnd.n2403 gnd.n2402 0.152939
R22207 gnd.n2404 gnd.n2403 0.152939
R22208 gnd.n2405 gnd.n2404 0.152939
R22209 gnd.n2406 gnd.n2405 0.152939
R22210 gnd.n2407 gnd.n2406 0.152939
R22211 gnd.n2408 gnd.n2407 0.152939
R22212 gnd.n2409 gnd.n2408 0.152939
R22213 gnd.n2410 gnd.n2409 0.152939
R22214 gnd.n2411 gnd.n2410 0.152939
R22215 gnd.n2412 gnd.n2411 0.152939
R22216 gnd.n2413 gnd.n2412 0.152939
R22217 gnd.n2414 gnd.n2413 0.152939
R22218 gnd.n2415 gnd.n2414 0.152939
R22219 gnd.n2418 gnd.n2415 0.152939
R22220 gnd.n2419 gnd.n2418 0.152939
R22221 gnd.n2420 gnd.n2419 0.152939
R22222 gnd.n2421 gnd.n2420 0.152939
R22223 gnd.n2422 gnd.n2421 0.152939
R22224 gnd.n2423 gnd.n2422 0.152939
R22225 gnd.n2424 gnd.n2423 0.152939
R22226 gnd.n2425 gnd.n2424 0.152939
R22227 gnd.n2426 gnd.n2425 0.152939
R22228 gnd.n2427 gnd.n2426 0.152939
R22229 gnd.n2428 gnd.n2427 0.152939
R22230 gnd.n2429 gnd.n2428 0.152939
R22231 gnd.n2430 gnd.n2429 0.152939
R22232 gnd.n2431 gnd.n2430 0.152939
R22233 gnd.n2432 gnd.n2431 0.152939
R22234 gnd.n2433 gnd.n2432 0.152939
R22235 gnd.n2434 gnd.n2433 0.152939
R22236 gnd.n2435 gnd.n2434 0.152939
R22237 gnd.n2436 gnd.n2435 0.152939
R22238 gnd.n2437 gnd.n2436 0.152939
R22239 gnd.n2440 gnd.n2437 0.152939
R22240 gnd.n2441 gnd.n2440 0.152939
R22241 gnd.n2442 gnd.n2441 0.152939
R22242 gnd.n2443 gnd.n2442 0.152939
R22243 gnd.n2444 gnd.n2443 0.152939
R22244 gnd.n2445 gnd.n2444 0.152939
R22245 gnd.n2446 gnd.n2445 0.152939
R22246 gnd.n2447 gnd.n2446 0.152939
R22247 gnd.n2448 gnd.n2447 0.152939
R22248 gnd.n2449 gnd.n2448 0.152939
R22249 gnd.n2450 gnd.n2449 0.152939
R22250 gnd.n2451 gnd.n2450 0.152939
R22251 gnd.n2452 gnd.n2451 0.152939
R22252 gnd.n2453 gnd.n2452 0.152939
R22253 gnd.n2454 gnd.n2453 0.152939
R22254 gnd.n2455 gnd.n2454 0.152939
R22255 gnd.n2456 gnd.n2455 0.152939
R22256 gnd.n2457 gnd.n2456 0.152939
R22257 gnd.n2458 gnd.n2457 0.152939
R22258 gnd.n6628 gnd.n2458 0.152939
R22259 gnd.n6628 gnd.n6627 0.152939
R22260 gnd.n2473 gnd.n2472 0.152939
R22261 gnd.n2474 gnd.n2473 0.152939
R22262 gnd.n2475 gnd.n2474 0.152939
R22263 gnd.n2495 gnd.n2475 0.152939
R22264 gnd.n2496 gnd.n2495 0.152939
R22265 gnd.n2497 gnd.n2496 0.152939
R22266 gnd.n2498 gnd.n2497 0.152939
R22267 gnd.n2513 gnd.n2498 0.152939
R22268 gnd.n2514 gnd.n2513 0.152939
R22269 gnd.n2515 gnd.n2514 0.152939
R22270 gnd.n2516 gnd.n2515 0.152939
R22271 gnd.n2534 gnd.n2516 0.152939
R22272 gnd.n2535 gnd.n2534 0.152939
R22273 gnd.n2536 gnd.n2535 0.152939
R22274 gnd.n2537 gnd.n2536 0.152939
R22275 gnd.n2553 gnd.n2537 0.152939
R22276 gnd.n2554 gnd.n2553 0.152939
R22277 gnd.n2555 gnd.n2554 0.152939
R22278 gnd.n2556 gnd.n2555 0.152939
R22279 gnd.n2574 gnd.n2556 0.152939
R22280 gnd.n2575 gnd.n2574 0.152939
R22281 gnd.n2576 gnd.n2575 0.152939
R22282 gnd.n2577 gnd.n2576 0.152939
R22283 gnd.n2593 gnd.n2577 0.152939
R22284 gnd.n2594 gnd.n2593 0.152939
R22285 gnd.n2595 gnd.n2594 0.152939
R22286 gnd.n6533 gnd.n2595 0.152939
R22287 gnd.n4227 gnd.n4221 0.152939
R22288 gnd.n4234 gnd.n4221 0.152939
R22289 gnd.n4235 gnd.n4234 0.152939
R22290 gnd.n4236 gnd.n4235 0.152939
R22291 gnd.n4236 gnd.n4066 0.152939
R22292 gnd.n4242 gnd.n4066 0.152939
R22293 gnd.n4243 gnd.n4242 0.152939
R22294 gnd.n4244 gnd.n4243 0.152939
R22295 gnd.n4244 gnd.n4051 0.152939
R22296 gnd.n4286 gnd.n4051 0.152939
R22297 gnd.n4287 gnd.n4286 0.152939
R22298 gnd.n4288 gnd.n4287 0.152939
R22299 gnd.n789 gnd.n788 0.152939
R22300 gnd.n790 gnd.n789 0.152939
R22301 gnd.n795 gnd.n790 0.152939
R22302 gnd.n796 gnd.n795 0.152939
R22303 gnd.n797 gnd.n796 0.152939
R22304 gnd.n798 gnd.n797 0.152939
R22305 gnd.n803 gnd.n798 0.152939
R22306 gnd.n804 gnd.n803 0.152939
R22307 gnd.n805 gnd.n804 0.152939
R22308 gnd.n806 gnd.n805 0.152939
R22309 gnd.n811 gnd.n806 0.152939
R22310 gnd.n812 gnd.n811 0.152939
R22311 gnd.n813 gnd.n812 0.152939
R22312 gnd.n814 gnd.n813 0.152939
R22313 gnd.n819 gnd.n814 0.152939
R22314 gnd.n820 gnd.n819 0.152939
R22315 gnd.n821 gnd.n820 0.152939
R22316 gnd.n822 gnd.n821 0.152939
R22317 gnd.n827 gnd.n822 0.152939
R22318 gnd.n828 gnd.n827 0.152939
R22319 gnd.n829 gnd.n828 0.152939
R22320 gnd.n830 gnd.n829 0.152939
R22321 gnd.n835 gnd.n830 0.152939
R22322 gnd.n836 gnd.n835 0.152939
R22323 gnd.n837 gnd.n836 0.152939
R22324 gnd.n838 gnd.n837 0.152939
R22325 gnd.n843 gnd.n838 0.152939
R22326 gnd.n844 gnd.n843 0.152939
R22327 gnd.n845 gnd.n844 0.152939
R22328 gnd.n846 gnd.n845 0.152939
R22329 gnd.n851 gnd.n846 0.152939
R22330 gnd.n852 gnd.n851 0.152939
R22331 gnd.n853 gnd.n852 0.152939
R22332 gnd.n854 gnd.n853 0.152939
R22333 gnd.n859 gnd.n854 0.152939
R22334 gnd.n860 gnd.n859 0.152939
R22335 gnd.n861 gnd.n860 0.152939
R22336 gnd.n862 gnd.n861 0.152939
R22337 gnd.n867 gnd.n862 0.152939
R22338 gnd.n868 gnd.n867 0.152939
R22339 gnd.n869 gnd.n868 0.152939
R22340 gnd.n870 gnd.n869 0.152939
R22341 gnd.n875 gnd.n870 0.152939
R22342 gnd.n876 gnd.n875 0.152939
R22343 gnd.n877 gnd.n876 0.152939
R22344 gnd.n878 gnd.n877 0.152939
R22345 gnd.n883 gnd.n878 0.152939
R22346 gnd.n884 gnd.n883 0.152939
R22347 gnd.n885 gnd.n884 0.152939
R22348 gnd.n886 gnd.n885 0.152939
R22349 gnd.n891 gnd.n886 0.152939
R22350 gnd.n892 gnd.n891 0.152939
R22351 gnd.n893 gnd.n892 0.152939
R22352 gnd.n894 gnd.n893 0.152939
R22353 gnd.n899 gnd.n894 0.152939
R22354 gnd.n900 gnd.n899 0.152939
R22355 gnd.n901 gnd.n900 0.152939
R22356 gnd.n902 gnd.n901 0.152939
R22357 gnd.n907 gnd.n902 0.152939
R22358 gnd.n908 gnd.n907 0.152939
R22359 gnd.n909 gnd.n908 0.152939
R22360 gnd.n910 gnd.n909 0.152939
R22361 gnd.n915 gnd.n910 0.152939
R22362 gnd.n916 gnd.n915 0.152939
R22363 gnd.n917 gnd.n916 0.152939
R22364 gnd.n918 gnd.n917 0.152939
R22365 gnd.n923 gnd.n918 0.152939
R22366 gnd.n924 gnd.n923 0.152939
R22367 gnd.n925 gnd.n924 0.152939
R22368 gnd.n926 gnd.n925 0.152939
R22369 gnd.n931 gnd.n926 0.152939
R22370 gnd.n932 gnd.n931 0.152939
R22371 gnd.n933 gnd.n932 0.152939
R22372 gnd.n934 gnd.n933 0.152939
R22373 gnd.n939 gnd.n934 0.152939
R22374 gnd.n940 gnd.n939 0.152939
R22375 gnd.n941 gnd.n940 0.152939
R22376 gnd.n942 gnd.n941 0.152939
R22377 gnd.n947 gnd.n942 0.152939
R22378 gnd.n948 gnd.n947 0.152939
R22379 gnd.n949 gnd.n948 0.152939
R22380 gnd.n950 gnd.n949 0.152939
R22381 gnd.n4224 gnd.n950 0.152939
R22382 gnd.n4226 gnd.n4224 0.152939
R22383 gnd.n4786 gnd.n3924 0.152939
R22384 gnd.n4787 gnd.n4786 0.152939
R22385 gnd.n4805 gnd.n4787 0.152939
R22386 gnd.n4805 gnd.n4804 0.152939
R22387 gnd.n4804 gnd.n4803 0.152939
R22388 gnd.n4803 gnd.n4788 0.152939
R22389 gnd.n4799 gnd.n4788 0.152939
R22390 gnd.n4799 gnd.n4798 0.152939
R22391 gnd.n4798 gnd.n4797 0.152939
R22392 gnd.n4797 gnd.n4792 0.152939
R22393 gnd.n4792 gnd.n2917 0.152939
R22394 gnd.n6309 gnd.n2917 0.152939
R22395 gnd.n6309 gnd.n6308 0.152939
R22396 gnd.n6308 gnd.n6307 0.152939
R22397 gnd.n6307 gnd.n2918 0.152939
R22398 gnd.n6303 gnd.n2918 0.152939
R22399 gnd.n6303 gnd.n6302 0.152939
R22400 gnd.n6302 gnd.n6301 0.152939
R22401 gnd.n6301 gnd.n2923 0.152939
R22402 gnd.n6297 gnd.n2923 0.152939
R22403 gnd.n6297 gnd.n6296 0.152939
R22404 gnd.n6296 gnd.n6295 0.152939
R22405 gnd.n6295 gnd.n2928 0.152939
R22406 gnd.n6291 gnd.n2928 0.152939
R22407 gnd.n6291 gnd.n6290 0.152939
R22408 gnd.n6290 gnd.n6289 0.152939
R22409 gnd.n6289 gnd.n2933 0.152939
R22410 gnd.n6285 gnd.n2933 0.152939
R22411 gnd.n6285 gnd.n6284 0.152939
R22412 gnd.n6284 gnd.n6283 0.152939
R22413 gnd.n6283 gnd.n2938 0.152939
R22414 gnd.n6279 gnd.n2938 0.152939
R22415 gnd.n6279 gnd.n6278 0.152939
R22416 gnd.n6278 gnd.n6277 0.152939
R22417 gnd.n6277 gnd.n2943 0.152939
R22418 gnd.n6273 gnd.n2943 0.152939
R22419 gnd.n6273 gnd.n6272 0.152939
R22420 gnd.n6272 gnd.n6271 0.152939
R22421 gnd.n6271 gnd.n2948 0.152939
R22422 gnd.n6267 gnd.n2948 0.152939
R22423 gnd.n6267 gnd.n6266 0.152939
R22424 gnd.n6266 gnd.n6265 0.152939
R22425 gnd.n6265 gnd.n2953 0.152939
R22426 gnd.n6261 gnd.n2953 0.152939
R22427 gnd.n6261 gnd.n6260 0.152939
R22428 gnd.n6260 gnd.n6259 0.152939
R22429 gnd.n6259 gnd.n2958 0.152939
R22430 gnd.n6255 gnd.n2958 0.152939
R22431 gnd.n6255 gnd.n6254 0.152939
R22432 gnd.n6254 gnd.n6253 0.152939
R22433 gnd.n6253 gnd.n2963 0.152939
R22434 gnd.n6249 gnd.n2963 0.152939
R22435 gnd.n6249 gnd.n6248 0.152939
R22436 gnd.n6248 gnd.n6247 0.152939
R22437 gnd.n6247 gnd.n2968 0.152939
R22438 gnd.n6243 gnd.n2968 0.152939
R22439 gnd.n6243 gnd.n6242 0.152939
R22440 gnd.n6242 gnd.n6241 0.152939
R22441 gnd.n6241 gnd.n2973 0.152939
R22442 gnd.n6237 gnd.n2973 0.152939
R22443 gnd.n6237 gnd.n6236 0.152939
R22444 gnd.n6236 gnd.n6235 0.152939
R22445 gnd.n6235 gnd.n2978 0.152939
R22446 gnd.n6231 gnd.n2978 0.152939
R22447 gnd.n6231 gnd.n6230 0.152939
R22448 gnd.n6230 gnd.n6229 0.152939
R22449 gnd.n6229 gnd.n2983 0.152939
R22450 gnd.n6225 gnd.n2983 0.152939
R22451 gnd.n6225 gnd.n6224 0.152939
R22452 gnd.n6224 gnd.n6223 0.152939
R22453 gnd.n6223 gnd.n2988 0.152939
R22454 gnd.n6219 gnd.n2988 0.152939
R22455 gnd.n6219 gnd.n6218 0.152939
R22456 gnd.n6218 gnd.n6217 0.152939
R22457 gnd.n6217 gnd.n2993 0.152939
R22458 gnd.n6213 gnd.n2993 0.152939
R22459 gnd.n6213 gnd.n6212 0.152939
R22460 gnd.n6212 gnd.n6211 0.152939
R22461 gnd.n6211 gnd.n2998 0.152939
R22462 gnd.n6207 gnd.n2998 0.152939
R22463 gnd.n6207 gnd.n6206 0.152939
R22464 gnd.n6206 gnd.n6205 0.152939
R22465 gnd.n4340 gnd.n4020 0.152939
R22466 gnd.n4341 gnd.n4340 0.152939
R22467 gnd.n4342 gnd.n4341 0.152939
R22468 gnd.n4342 gnd.n4008 0.152939
R22469 gnd.n4379 gnd.n4008 0.152939
R22470 gnd.n4380 gnd.n4379 0.152939
R22471 gnd.n4381 gnd.n4380 0.152939
R22472 gnd.n4381 gnd.n4002 0.152939
R22473 gnd.n4393 gnd.n4002 0.152939
R22474 gnd.n4394 gnd.n4393 0.152939
R22475 gnd.n4395 gnd.n4394 0.152939
R22476 gnd.n4395 gnd.n3994 0.152939
R22477 gnd.n4430 gnd.n3994 0.152939
R22478 gnd.n4430 gnd.n4429 0.152939
R22479 gnd.n4429 gnd.n4428 0.152939
R22480 gnd.n4428 gnd.n3995 0.152939
R22481 gnd.n4424 gnd.n3995 0.152939
R22482 gnd.n4424 gnd.n4423 0.152939
R22483 gnd.n4423 gnd.n4422 0.152939
R22484 gnd.n4422 gnd.n3977 0.152939
R22485 gnd.n4460 gnd.n3977 0.152939
R22486 gnd.n4461 gnd.n4460 0.152939
R22487 gnd.n4462 gnd.n4461 0.152939
R22488 gnd.n4462 gnd.n3971 0.152939
R22489 gnd.n4734 gnd.n3971 0.152939
R22490 gnd.n4734 gnd.n4733 0.152939
R22491 gnd.n4733 gnd.n4732 0.152939
R22492 gnd.n4732 gnd.n3972 0.152939
R22493 gnd.n4728 gnd.n3972 0.152939
R22494 gnd.n4728 gnd.n4727 0.152939
R22495 gnd.n4727 gnd.n3951 0.152939
R22496 gnd.n4482 gnd.n4481 0.152939
R22497 gnd.n4499 gnd.n4481 0.152939
R22498 gnd.n4500 gnd.n4499 0.152939
R22499 gnd.n4501 gnd.n4500 0.152939
R22500 gnd.n4501 gnd.n4477 0.152939
R22501 gnd.n4620 gnd.n4477 0.152939
R22502 gnd.n4490 gnd.n4489 0.152939
R22503 gnd.n4489 gnd.n4488 0.152939
R22504 gnd.n4488 gnd.n4484 0.152939
R22505 gnd.n4484 gnd.n3906 0.152939
R22506 gnd.n4828 gnd.n3906 0.152939
R22507 gnd.n4829 gnd.n4828 0.152939
R22508 gnd.n4830 gnd.n4829 0.152939
R22509 gnd.n4830 gnd.n3902 0.152939
R22510 gnd.n4836 gnd.n3902 0.152939
R22511 gnd.n4837 gnd.n4836 0.152939
R22512 gnd.n4979 gnd.n4837 0.152939
R22513 gnd.n4979 gnd.n4978 0.152939
R22514 gnd.n4978 gnd.n4977 0.152939
R22515 gnd.n4977 gnd.n4838 0.152939
R22516 gnd.n4973 gnd.n4838 0.152939
R22517 gnd.n4973 gnd.n4972 0.152939
R22518 gnd.n4972 gnd.n4971 0.152939
R22519 gnd.n4971 gnd.n4841 0.152939
R22520 gnd.n4967 gnd.n4841 0.152939
R22521 gnd.n4967 gnd.n4966 0.152939
R22522 gnd.n4966 gnd.n4965 0.152939
R22523 gnd.n4965 gnd.n4844 0.152939
R22524 gnd.n4961 gnd.n4844 0.152939
R22525 gnd.n4961 gnd.n4960 0.152939
R22526 gnd.n4960 gnd.n4959 0.152939
R22527 gnd.n4959 gnd.n4850 0.152939
R22528 gnd.n4955 gnd.n4850 0.152939
R22529 gnd.n4955 gnd.n4954 0.152939
R22530 gnd.n4954 gnd.n4953 0.152939
R22531 gnd.n4953 gnd.n4854 0.152939
R22532 gnd.n4949 gnd.n4854 0.152939
R22533 gnd.n4949 gnd.n4948 0.152939
R22534 gnd.n4948 gnd.n4947 0.152939
R22535 gnd.n4947 gnd.n4858 0.152939
R22536 gnd.n4943 gnd.n4858 0.152939
R22537 gnd.n4943 gnd.n4942 0.152939
R22538 gnd.n4942 gnd.n4941 0.152939
R22539 gnd.n4941 gnd.n4861 0.152939
R22540 gnd.n4937 gnd.n4861 0.152939
R22541 gnd.n4937 gnd.n4936 0.152939
R22542 gnd.n4936 gnd.n4935 0.152939
R22543 gnd.n4935 gnd.n4867 0.152939
R22544 gnd.n4931 gnd.n4867 0.152939
R22545 gnd.n4931 gnd.n4930 0.152939
R22546 gnd.n4930 gnd.n4929 0.152939
R22547 gnd.n4929 gnd.n4870 0.152939
R22548 gnd.n4925 gnd.n4870 0.152939
R22549 gnd.n4925 gnd.n4924 0.152939
R22550 gnd.n4924 gnd.n4923 0.152939
R22551 gnd.n4923 gnd.n4874 0.152939
R22552 gnd.n4919 gnd.n4874 0.152939
R22553 gnd.n4919 gnd.n4918 0.152939
R22554 gnd.n4918 gnd.n4917 0.152939
R22555 gnd.n4917 gnd.n4879 0.152939
R22556 gnd.n4913 gnd.n4879 0.152939
R22557 gnd.n4913 gnd.n4912 0.152939
R22558 gnd.n4912 gnd.n4911 0.152939
R22559 gnd.n4911 gnd.n4883 0.152939
R22560 gnd.n4907 gnd.n4883 0.152939
R22561 gnd.n4907 gnd.n4906 0.152939
R22562 gnd.n4906 gnd.n4905 0.152939
R22563 gnd.n4905 gnd.n4888 0.152939
R22564 gnd.n4901 gnd.n4888 0.152939
R22565 gnd.n4901 gnd.n4900 0.152939
R22566 gnd.n4900 gnd.n4899 0.152939
R22567 gnd.n4899 gnd.n4893 0.152939
R22568 gnd.n4895 gnd.n4893 0.152939
R22569 gnd.n4895 gnd.n3541 0.152939
R22570 gnd.n5408 gnd.n3541 0.152939
R22571 gnd.n5409 gnd.n5408 0.152939
R22572 gnd.n5411 gnd.n5409 0.152939
R22573 gnd.n5411 gnd.n5410 0.152939
R22574 gnd.n5410 gnd.n3442 0.152939
R22575 gnd.n5556 gnd.n3442 0.152939
R22576 gnd.n5557 gnd.n5556 0.152939
R22577 gnd.n5558 gnd.n5557 0.152939
R22578 gnd.n5558 gnd.n3430 0.152939
R22579 gnd.n5575 gnd.n3430 0.152939
R22580 gnd.n5576 gnd.n5575 0.152939
R22581 gnd.n5577 gnd.n5576 0.152939
R22582 gnd.n5577 gnd.n3012 0.152939
R22583 gnd.n6199 gnd.n3012 0.152939
R22584 gnd.n6198 gnd.n3013 0.152939
R22585 gnd.n6194 gnd.n3013 0.152939
R22586 gnd.n6194 gnd.n6193 0.152939
R22587 gnd.n6193 gnd.n6192 0.152939
R22588 gnd.n6192 gnd.n3017 0.152939
R22589 gnd.n6188 gnd.n3017 0.152939
R22590 gnd.n5690 gnd.n5689 0.152939
R22591 gnd.n5690 gnd.n3391 0.152939
R22592 gnd.n5696 gnd.n3391 0.152939
R22593 gnd.n5697 gnd.n5696 0.152939
R22594 gnd.n5698 gnd.n5697 0.152939
R22595 gnd.n5698 gnd.n3387 0.152939
R22596 gnd.n5711 gnd.n3387 0.152939
R22597 gnd.n5712 gnd.n5711 0.152939
R22598 gnd.n5713 gnd.n5712 0.152939
R22599 gnd.n5713 gnd.n3383 0.152939
R22600 gnd.n5726 gnd.n3383 0.152939
R22601 gnd.n5727 gnd.n5726 0.152939
R22602 gnd.n5728 gnd.n5727 0.152939
R22603 gnd.n5728 gnd.n3378 0.152939
R22604 gnd.n5741 gnd.n3378 0.152939
R22605 gnd.n5742 gnd.n5741 0.152939
R22606 gnd.n5743 gnd.n5742 0.152939
R22607 gnd.n5743 gnd.n3374 0.152939
R22608 gnd.n5756 gnd.n3374 0.152939
R22609 gnd.n5757 gnd.n5756 0.152939
R22610 gnd.n5758 gnd.n5757 0.152939
R22611 gnd.n5758 gnd.n3369 0.152939
R22612 gnd.n5771 gnd.n3369 0.152939
R22613 gnd.n5772 gnd.n5771 0.152939
R22614 gnd.n5785 gnd.n5772 0.152939
R22615 gnd.n5785 gnd.n5784 0.152939
R22616 gnd.n5784 gnd.n5783 0.152939
R22617 gnd.n5783 gnd.n5773 0.152939
R22618 gnd.n5779 gnd.n5773 0.152939
R22619 gnd.n5779 gnd.n5778 0.152939
R22620 gnd.n5778 gnd.n95 0.152939
R22621 gnd.n8072 gnd.n8071 0.145814
R22622 gnd.n4312 gnd.n4311 0.145814
R22623 gnd.n4312 gnd.n4020 0.145814
R22624 gnd.n8072 gnd.n95 0.145814
R22625 gnd.n4621 gnd.n4620 0.128549
R22626 gnd.n6188 gnd.n6187 0.128549
R22627 gnd.n5823 gnd.n111 0.0797683
R22628 gnd.n4288 gnd.n2616 0.0797683
R22629 gnd.n1846 gnd.n1245 0.0767195
R22630 gnd.n1846 gnd.n1845 0.0767195
R22631 gnd.n4351 gnd.n2616 0.0736707
R22632 gnd.n5631 gnd.n111 0.0736707
R22633 gnd.n4718 gnd.n4621 0.063
R22634 gnd.n6187 gnd.n3022 0.063
R22635 gnd.n6804 gnd.n1009 0.0477147
R22636 gnd.n1636 gnd.n1524 0.0442063
R22637 gnd.n1637 gnd.n1636 0.0442063
R22638 gnd.n1638 gnd.n1637 0.0442063
R22639 gnd.n1638 gnd.n1513 0.0442063
R22640 gnd.n1652 gnd.n1513 0.0442063
R22641 gnd.n1653 gnd.n1652 0.0442063
R22642 gnd.n1654 gnd.n1653 0.0442063
R22643 gnd.n1654 gnd.n1500 0.0442063
R22644 gnd.n1698 gnd.n1500 0.0442063
R22645 gnd.n1699 gnd.n1698 0.0442063
R22646 gnd.n3190 gnd.n3022 0.0416005
R22647 gnd.n7853 gnd.n7852 0.0416005
R22648 gnd.n6626 gnd.n6625 0.0416005
R22649 gnd.n4719 gnd.n4718 0.0416005
R22650 gnd.n1701 gnd.n1434 0.0344674
R22651 gnd.n6009 gnd.n3190 0.0344674
R22652 gnd.n6009 gnd.n3192 0.0344674
R22653 gnd.n3216 gnd.n3192 0.0344674
R22654 gnd.n3217 gnd.n3216 0.0344674
R22655 gnd.n3218 gnd.n3217 0.0344674
R22656 gnd.n3219 gnd.n3218 0.0344674
R22657 gnd.n5705 gnd.n3219 0.0344674
R22658 gnd.n5705 gnd.n3238 0.0344674
R22659 gnd.n3239 gnd.n3238 0.0344674
R22660 gnd.n3240 gnd.n3239 0.0344674
R22661 gnd.n5720 gnd.n3240 0.0344674
R22662 gnd.n5720 gnd.n3258 0.0344674
R22663 gnd.n3259 gnd.n3258 0.0344674
R22664 gnd.n3260 gnd.n3259 0.0344674
R22665 gnd.n5735 gnd.n3260 0.0344674
R22666 gnd.n5735 gnd.n3279 0.0344674
R22667 gnd.n3280 gnd.n3279 0.0344674
R22668 gnd.n3281 gnd.n3280 0.0344674
R22669 gnd.n5750 gnd.n3281 0.0344674
R22670 gnd.n5750 gnd.n3299 0.0344674
R22671 gnd.n3300 gnd.n3299 0.0344674
R22672 gnd.n3301 gnd.n3300 0.0344674
R22673 gnd.n5765 gnd.n3301 0.0344674
R22674 gnd.n5765 gnd.n3321 0.0344674
R22675 gnd.n3322 gnd.n3321 0.0344674
R22676 gnd.n3323 gnd.n3322 0.0344674
R22677 gnd.n3365 gnd.n3323 0.0344674
R22678 gnd.n5796 gnd.n3365 0.0344674
R22679 gnd.n5801 gnd.n5796 0.0344674
R22680 gnd.n5802 gnd.n5801 0.0344674
R22681 gnd.n5802 gnd.n3356 0.0344674
R22682 gnd.n3357 gnd.n3356 0.0344674
R22683 gnd.n3358 gnd.n3357 0.0344674
R22684 gnd.n5806 gnd.n3358 0.0344674
R22685 gnd.n5807 gnd.n5806 0.0344674
R22686 gnd.n5808 gnd.n5807 0.0344674
R22687 gnd.n5808 gnd.n125 0.0344674
R22688 gnd.n126 gnd.n125 0.0344674
R22689 gnd.n127 gnd.n126 0.0344674
R22690 gnd.n5841 gnd.n127 0.0344674
R22691 gnd.n5841 gnd.n143 0.0344674
R22692 gnd.n144 gnd.n143 0.0344674
R22693 gnd.n145 gnd.n144 0.0344674
R22694 gnd.n5867 gnd.n145 0.0344674
R22695 gnd.n5867 gnd.n164 0.0344674
R22696 gnd.n165 gnd.n164 0.0344674
R22697 gnd.n166 gnd.n165 0.0344674
R22698 gnd.n356 gnd.n166 0.0344674
R22699 gnd.n356 gnd.n183 0.0344674
R22700 gnd.n184 gnd.n183 0.0344674
R22701 gnd.n185 gnd.n184 0.0344674
R22702 gnd.n7828 gnd.n185 0.0344674
R22703 gnd.n7828 gnd.n204 0.0344674
R22704 gnd.n205 gnd.n204 0.0344674
R22705 gnd.n206 gnd.n205 0.0344674
R22706 gnd.n7835 gnd.n206 0.0344674
R22707 gnd.n7835 gnd.n222 0.0344674
R22708 gnd.n223 gnd.n222 0.0344674
R22709 gnd.n224 gnd.n223 0.0344674
R22710 gnd.n7842 gnd.n224 0.0344674
R22711 gnd.n7842 gnd.n242 0.0344674
R22712 gnd.n243 gnd.n242 0.0344674
R22713 gnd.n244 gnd.n243 0.0344674
R22714 gnd.n7852 gnd.n244 0.0344674
R22715 gnd.n6625 gnd.n2464 0.0344674
R22716 gnd.n4073 gnd.n2464 0.0344674
R22717 gnd.n4073 gnd.n2486 0.0344674
R22718 gnd.n2487 gnd.n2486 0.0344674
R22719 gnd.n2488 gnd.n2487 0.0344674
R22720 gnd.n4079 gnd.n2488 0.0344674
R22721 gnd.n4079 gnd.n2505 0.0344674
R22722 gnd.n2506 gnd.n2505 0.0344674
R22723 gnd.n2507 gnd.n2506 0.0344674
R22724 gnd.n4086 gnd.n2507 0.0344674
R22725 gnd.n4086 gnd.n2524 0.0344674
R22726 gnd.n2525 gnd.n2524 0.0344674
R22727 gnd.n2526 gnd.n2525 0.0344674
R22728 gnd.n4093 gnd.n2526 0.0344674
R22729 gnd.n4093 gnd.n2544 0.0344674
R22730 gnd.n2545 gnd.n2544 0.0344674
R22731 gnd.n2546 gnd.n2545 0.0344674
R22732 gnd.n4203 gnd.n2546 0.0344674
R22733 gnd.n4203 gnd.n2564 0.0344674
R22734 gnd.n2565 gnd.n2564 0.0344674
R22735 gnd.n2566 gnd.n2565 0.0344674
R22736 gnd.n4206 gnd.n2566 0.0344674
R22737 gnd.n4206 gnd.n2584 0.0344674
R22738 gnd.n2585 gnd.n2584 0.0344674
R22739 gnd.n2586 gnd.n2585 0.0344674
R22740 gnd.n4261 gnd.n2586 0.0344674
R22741 gnd.n4261 gnd.n2603 0.0344674
R22742 gnd.n2604 gnd.n2603 0.0344674
R22743 gnd.n2605 gnd.n2604 0.0344674
R22744 gnd.n4270 gnd.n2605 0.0344674
R22745 gnd.n4270 gnd.n4269 0.0344674
R22746 gnd.n4269 gnd.n4038 0.0344674
R22747 gnd.n4038 gnd.n4034 0.0344674
R22748 gnd.n4035 gnd.n4034 0.0344674
R22749 gnd.n4325 gnd.n4035 0.0344674
R22750 gnd.n4325 gnd.n4036 0.0344674
R22751 gnd.n4036 gnd.n2631 0.0344674
R22752 gnd.n2632 gnd.n2631 0.0344674
R22753 gnd.n2633 gnd.n2632 0.0344674
R22754 gnd.n4006 gnd.n2633 0.0344674
R22755 gnd.n4006 gnd.n2649 0.0344674
R22756 gnd.n2650 gnd.n2649 0.0344674
R22757 gnd.n2651 gnd.n2650 0.0344674
R22758 gnd.n4000 gnd.n2651 0.0344674
R22759 gnd.n4000 gnd.n2670 0.0344674
R22760 gnd.n2671 gnd.n2670 0.0344674
R22761 gnd.n2672 gnd.n2671 0.0344674
R22762 gnd.n4404 gnd.n2672 0.0344674
R22763 gnd.n4404 gnd.n2689 0.0344674
R22764 gnd.n2690 gnd.n2689 0.0344674
R22765 gnd.n2691 gnd.n2690 0.0344674
R22766 gnd.n4414 gnd.n2691 0.0344674
R22767 gnd.n4414 gnd.n2710 0.0344674
R22768 gnd.n2711 gnd.n2710 0.0344674
R22769 gnd.n2712 gnd.n2711 0.0344674
R22770 gnd.n3975 gnd.n2712 0.0344674
R22771 gnd.n3975 gnd.n2729 0.0344674
R22772 gnd.n2730 gnd.n2729 0.0344674
R22773 gnd.n2731 gnd.n2730 0.0344674
R22774 gnd.n4471 gnd.n2731 0.0344674
R22775 gnd.n4471 gnd.n2750 0.0344674
R22776 gnd.n2751 gnd.n2750 0.0344674
R22777 gnd.n2752 gnd.n2751 0.0344674
R22778 gnd.n4719 gnd.n2752 0.0344674
R22779 gnd.n4616 gnd.n4476 0.0344674
R22780 gnd.n6186 gnd.n6185 0.0344674
R22781 gnd.n4770 gnd.n4769 0.029712
R22782 gnd.n5688 gnd.n5687 0.029712
R22783 gnd.n1721 gnd.n1720 0.0269946
R22784 gnd.n1723 gnd.n1722 0.0269946
R22785 gnd.n1429 gnd.n1427 0.0269946
R22786 gnd.n1733 gnd.n1731 0.0269946
R22787 gnd.n1732 gnd.n1408 0.0269946
R22788 gnd.n1752 gnd.n1751 0.0269946
R22789 gnd.n1754 gnd.n1753 0.0269946
R22790 gnd.n1403 gnd.n1402 0.0269946
R22791 gnd.n1764 gnd.n1398 0.0269946
R22792 gnd.n1763 gnd.n1400 0.0269946
R22793 gnd.n1399 gnd.n1379 0.0269946
R22794 gnd.n1790 gnd.n1380 0.0269946
R22795 gnd.n1789 gnd.n1381 0.0269946
R22796 gnd.n1809 gnd.n1365 0.0269946
R22797 gnd.n1811 gnd.n1810 0.0269946
R22798 gnd.n1812 gnd.n1345 0.0269946
R22799 gnd.n1813 gnd.n1346 0.0269946
R22800 gnd.n1814 gnd.n1347 0.0269946
R22801 gnd.n1349 gnd.n1348 0.0269946
R22802 gnd.n1238 gnd.n1237 0.0269946
R22803 gnd.n1858 gnd.n1234 0.0269946
R22804 gnd.n1857 gnd.n1235 0.0269946
R22805 gnd.n1877 gnd.n1217 0.0269946
R22806 gnd.n1879 gnd.n1878 0.0269946
R22807 gnd.n1880 gnd.n1215 0.0269946
R22808 gnd.n1887 gnd.n1883 0.0269946
R22809 gnd.n1886 gnd.n1885 0.0269946
R22810 gnd.n1884 gnd.n1194 0.0269946
R22811 gnd.n1910 gnd.n1195 0.0269946
R22812 gnd.n1909 gnd.n1196 0.0269946
R22813 gnd.n1955 gnd.n1172 0.0269946
R22814 gnd.n1957 gnd.n1956 0.0269946
R22815 gnd.n1966 gnd.n1165 0.0269946
R22816 gnd.n1968 gnd.n1967 0.0269946
R22817 gnd.n1969 gnd.n1163 0.0269946
R22818 gnd.n1976 gnd.n1972 0.0269946
R22819 gnd.n1975 gnd.n1974 0.0269946
R22820 gnd.n1973 gnd.n1143 0.0269946
R22821 gnd.n2000 gnd.n1144 0.0269946
R22822 gnd.n1999 gnd.n1145 0.0269946
R22823 gnd.n2060 gnd.n1120 0.0269946
R22824 gnd.n2062 gnd.n2061 0.0269946
R22825 gnd.n2063 gnd.n959 0.0269946
R22826 gnd.n1115 gnd.n960 0.0269946
R22827 gnd.n1117 gnd.n961 0.0269946
R22828 gnd.n2071 gnd.n2070 0.0269946
R22829 gnd.n2073 gnd.n2072 0.0269946
R22830 gnd.n2074 gnd.n983 0.0269946
R22831 gnd.n2334 gnd.n985 0.0269946
R22832 gnd.n2340 gnd.n2339 0.0269946
R22833 gnd.n2342 gnd.n2341 0.0269946
R22834 gnd.n6805 gnd.n1008 0.0269946
R22835 gnd.n4615 gnd.n4509 0.0225788
R22836 gnd.n4612 gnd.n4611 0.0225788
R22837 gnd.n4608 gnd.n4512 0.0225788
R22838 gnd.n4607 gnd.n4518 0.0225788
R22839 gnd.n4604 gnd.n4603 0.0225788
R22840 gnd.n4600 gnd.n4524 0.0225788
R22841 gnd.n4599 gnd.n4528 0.0225788
R22842 gnd.n4596 gnd.n4595 0.0225788
R22843 gnd.n4592 gnd.n4532 0.0225788
R22844 gnd.n4591 gnd.n4538 0.0225788
R22845 gnd.n4588 gnd.n4587 0.0225788
R22846 gnd.n4584 gnd.n4544 0.0225788
R22847 gnd.n4583 gnd.n4548 0.0225788
R22848 gnd.n4580 gnd.n4579 0.0225788
R22849 gnd.n4576 gnd.n4552 0.0225788
R22850 gnd.n4575 gnd.n4558 0.0225788
R22851 gnd.n4572 gnd.n4571 0.0225788
R22852 gnd.n4563 gnd.n3952 0.0225788
R22853 gnd.n4769 gnd.n4768 0.0225788
R22854 gnd.n6182 gnd.n3023 0.0225788
R22855 gnd.n6181 gnd.n3027 0.0225788
R22856 gnd.n6178 gnd.n6177 0.0225788
R22857 gnd.n6174 gnd.n3032 0.0225788
R22858 gnd.n6173 gnd.n3036 0.0225788
R22859 gnd.n6170 gnd.n6169 0.0225788
R22860 gnd.n6166 gnd.n3040 0.0225788
R22861 gnd.n6165 gnd.n3044 0.0225788
R22862 gnd.n6162 gnd.n6161 0.0225788
R22863 gnd.n6158 gnd.n3048 0.0225788
R22864 gnd.n6157 gnd.n3052 0.0225788
R22865 gnd.n6154 gnd.n6153 0.0225788
R22866 gnd.n6150 gnd.n3056 0.0225788
R22867 gnd.n6149 gnd.n3060 0.0225788
R22868 gnd.n6146 gnd.n6145 0.0225788
R22869 gnd.n6142 gnd.n3064 0.0225788
R22870 gnd.n6141 gnd.n3070 0.0225788
R22871 gnd.n3395 gnd.n3073 0.0225788
R22872 gnd.n5687 gnd.n3394 0.0225788
R22873 gnd.n5688 gnd.n3003 0.0218415
R22874 gnd.n4771 gnd.n4770 0.0218415
R22875 gnd.n1701 gnd.n1700 0.0202011
R22876 gnd.n1700 gnd.n1699 0.0148637
R22877 gnd.n2332 gnd.n2331 0.0144266
R22878 gnd.n2331 gnd.n984 0.0130679
R22879 gnd.n4616 gnd.n4615 0.0123886
R22880 gnd.n4612 gnd.n4509 0.0123886
R22881 gnd.n4611 gnd.n4512 0.0123886
R22882 gnd.n4608 gnd.n4607 0.0123886
R22883 gnd.n4604 gnd.n4518 0.0123886
R22884 gnd.n4603 gnd.n4524 0.0123886
R22885 gnd.n4600 gnd.n4599 0.0123886
R22886 gnd.n4596 gnd.n4528 0.0123886
R22887 gnd.n4595 gnd.n4532 0.0123886
R22888 gnd.n4592 gnd.n4591 0.0123886
R22889 gnd.n4588 gnd.n4538 0.0123886
R22890 gnd.n4587 gnd.n4544 0.0123886
R22891 gnd.n4584 gnd.n4583 0.0123886
R22892 gnd.n4580 gnd.n4548 0.0123886
R22893 gnd.n4579 gnd.n4552 0.0123886
R22894 gnd.n4576 gnd.n4575 0.0123886
R22895 gnd.n4572 gnd.n4558 0.0123886
R22896 gnd.n4571 gnd.n4563 0.0123886
R22897 gnd.n4768 gnd.n3952 0.0123886
R22898 gnd.n6185 gnd.n3023 0.0123886
R22899 gnd.n6182 gnd.n6181 0.0123886
R22900 gnd.n6178 gnd.n3027 0.0123886
R22901 gnd.n6177 gnd.n3032 0.0123886
R22902 gnd.n6174 gnd.n6173 0.0123886
R22903 gnd.n6170 gnd.n3036 0.0123886
R22904 gnd.n6169 gnd.n3040 0.0123886
R22905 gnd.n6166 gnd.n6165 0.0123886
R22906 gnd.n6162 gnd.n3044 0.0123886
R22907 gnd.n6161 gnd.n3048 0.0123886
R22908 gnd.n6158 gnd.n6157 0.0123886
R22909 gnd.n6154 gnd.n3052 0.0123886
R22910 gnd.n6153 gnd.n3056 0.0123886
R22911 gnd.n6150 gnd.n6149 0.0123886
R22912 gnd.n6146 gnd.n3060 0.0123886
R22913 gnd.n6145 gnd.n3064 0.0123886
R22914 gnd.n6142 gnd.n6141 0.0123886
R22915 gnd.n3073 gnd.n3070 0.0123886
R22916 gnd.n3395 gnd.n3394 0.0123886
R22917 gnd.n1720 gnd.n1434 0.00797283
R22918 gnd.n1722 gnd.n1721 0.00797283
R22919 gnd.n1723 gnd.n1429 0.00797283
R22920 gnd.n1731 gnd.n1427 0.00797283
R22921 gnd.n1733 gnd.n1732 0.00797283
R22922 gnd.n1751 gnd.n1408 0.00797283
R22923 gnd.n1753 gnd.n1752 0.00797283
R22924 gnd.n1754 gnd.n1403 0.00797283
R22925 gnd.n1402 gnd.n1398 0.00797283
R22926 gnd.n1764 gnd.n1763 0.00797283
R22927 gnd.n1400 gnd.n1399 0.00797283
R22928 gnd.n1380 gnd.n1379 0.00797283
R22929 gnd.n1790 gnd.n1789 0.00797283
R22930 gnd.n1381 gnd.n1365 0.00797283
R22931 gnd.n1810 gnd.n1809 0.00797283
R22932 gnd.n1812 gnd.n1811 0.00797283
R22933 gnd.n1813 gnd.n1345 0.00797283
R22934 gnd.n1814 gnd.n1346 0.00797283
R22935 gnd.n1348 gnd.n1347 0.00797283
R22936 gnd.n1349 gnd.n1238 0.00797283
R22937 gnd.n1237 gnd.n1234 0.00797283
R22938 gnd.n1858 gnd.n1857 0.00797283
R22939 gnd.n1235 gnd.n1217 0.00797283
R22940 gnd.n1878 gnd.n1877 0.00797283
R22941 gnd.n1880 gnd.n1879 0.00797283
R22942 gnd.n1883 gnd.n1215 0.00797283
R22943 gnd.n1887 gnd.n1886 0.00797283
R22944 gnd.n1885 gnd.n1884 0.00797283
R22945 gnd.n1195 gnd.n1194 0.00797283
R22946 gnd.n1910 gnd.n1909 0.00797283
R22947 gnd.n1196 gnd.n1172 0.00797283
R22948 gnd.n1957 gnd.n1955 0.00797283
R22949 gnd.n1956 gnd.n1165 0.00797283
R22950 gnd.n1967 gnd.n1966 0.00797283
R22951 gnd.n1969 gnd.n1968 0.00797283
R22952 gnd.n1972 gnd.n1163 0.00797283
R22953 gnd.n1976 gnd.n1975 0.00797283
R22954 gnd.n1974 gnd.n1973 0.00797283
R22955 gnd.n1144 gnd.n1143 0.00797283
R22956 gnd.n2000 gnd.n1999 0.00797283
R22957 gnd.n1145 gnd.n1120 0.00797283
R22958 gnd.n2061 gnd.n2060 0.00797283
R22959 gnd.n2063 gnd.n2062 0.00797283
R22960 gnd.n1115 gnd.n959 0.00797283
R22961 gnd.n1117 gnd.n960 0.00797283
R22962 gnd.n2070 gnd.n961 0.00797283
R22963 gnd.n2072 gnd.n2071 0.00797283
R22964 gnd.n2074 gnd.n2073 0.00797283
R22965 gnd.n2332 gnd.n983 0.00797283
R22966 gnd.n2334 gnd.n984 0.00797283
R22967 gnd.n2339 gnd.n985 0.00797283
R22968 gnd.n2342 gnd.n2340 0.00797283
R22969 gnd.n2341 gnd.n1008 0.00797283
R22970 gnd.n6805 gnd.n6804 0.00797283
R22971 gnd.n4621 gnd.n4476 0.00593478
R22972 gnd.n6187 gnd.n6186 0.00593478
R22973 CSoutput.n19 CSoutput.t235 184.661
R22974 CSoutput.n78 CSoutput.n77 165.8
R22975 CSoutput.n76 CSoutput.n0 165.8
R22976 CSoutput.n75 CSoutput.n74 165.8
R22977 CSoutput.n73 CSoutput.n72 165.8
R22978 CSoutput.n71 CSoutput.n2 165.8
R22979 CSoutput.n69 CSoutput.n68 165.8
R22980 CSoutput.n67 CSoutput.n3 165.8
R22981 CSoutput.n66 CSoutput.n65 165.8
R22982 CSoutput.n63 CSoutput.n4 165.8
R22983 CSoutput.n61 CSoutput.n60 165.8
R22984 CSoutput.n59 CSoutput.n5 165.8
R22985 CSoutput.n58 CSoutput.n57 165.8
R22986 CSoutput.n55 CSoutput.n6 165.8
R22987 CSoutput.n54 CSoutput.n53 165.8
R22988 CSoutput.n52 CSoutput.n51 165.8
R22989 CSoutput.n50 CSoutput.n8 165.8
R22990 CSoutput.n48 CSoutput.n47 165.8
R22991 CSoutput.n46 CSoutput.n9 165.8
R22992 CSoutput.n45 CSoutput.n44 165.8
R22993 CSoutput.n42 CSoutput.n10 165.8
R22994 CSoutput.n41 CSoutput.n40 165.8
R22995 CSoutput.n39 CSoutput.n38 165.8
R22996 CSoutput.n37 CSoutput.n12 165.8
R22997 CSoutput.n35 CSoutput.n34 165.8
R22998 CSoutput.n33 CSoutput.n13 165.8
R22999 CSoutput.n32 CSoutput.n31 165.8
R23000 CSoutput.n29 CSoutput.n14 165.8
R23001 CSoutput.n28 CSoutput.n27 165.8
R23002 CSoutput.n26 CSoutput.n25 165.8
R23003 CSoutput.n24 CSoutput.n16 165.8
R23004 CSoutput.n22 CSoutput.n21 165.8
R23005 CSoutput.n20 CSoutput.n17 165.8
R23006 CSoutput.n77 CSoutput.t236 162.194
R23007 CSoutput.n18 CSoutput.t225 120.501
R23008 CSoutput.n23 CSoutput.t227 120.501
R23009 CSoutput.n15 CSoutput.t220 120.501
R23010 CSoutput.n30 CSoutput.t233 120.501
R23011 CSoutput.n36 CSoutput.t228 120.501
R23012 CSoutput.n11 CSoutput.t223 120.501
R23013 CSoutput.n43 CSoutput.t218 120.501
R23014 CSoutput.n49 CSoutput.t229 120.501
R23015 CSoutput.n7 CSoutput.t231 120.501
R23016 CSoutput.n56 CSoutput.t221 120.501
R23017 CSoutput.n62 CSoutput.t217 120.501
R23018 CSoutput.n64 CSoutput.t234 120.501
R23019 CSoutput.n70 CSoutput.t224 120.501
R23020 CSoutput.n1 CSoutput.t226 120.501
R23021 CSoutput.n310 CSoutput.n308 103.469
R23022 CSoutput.n294 CSoutput.n292 103.469
R23023 CSoutput.n279 CSoutput.n277 103.469
R23024 CSoutput.n112 CSoutput.n110 103.469
R23025 CSoutput.n96 CSoutput.n94 103.469
R23026 CSoutput.n81 CSoutput.n79 103.469
R23027 CSoutput.n320 CSoutput.n319 103.111
R23028 CSoutput.n318 CSoutput.n317 103.111
R23029 CSoutput.n316 CSoutput.n315 103.111
R23030 CSoutput.n314 CSoutput.n313 103.111
R23031 CSoutput.n312 CSoutput.n311 103.111
R23032 CSoutput.n310 CSoutput.n309 103.111
R23033 CSoutput.n306 CSoutput.n305 103.111
R23034 CSoutput.n304 CSoutput.n303 103.111
R23035 CSoutput.n302 CSoutput.n301 103.111
R23036 CSoutput.n300 CSoutput.n299 103.111
R23037 CSoutput.n298 CSoutput.n297 103.111
R23038 CSoutput.n296 CSoutput.n295 103.111
R23039 CSoutput.n294 CSoutput.n293 103.111
R23040 CSoutput.n291 CSoutput.n290 103.111
R23041 CSoutput.n289 CSoutput.n288 103.111
R23042 CSoutput.n287 CSoutput.n286 103.111
R23043 CSoutput.n285 CSoutput.n284 103.111
R23044 CSoutput.n283 CSoutput.n282 103.111
R23045 CSoutput.n281 CSoutput.n280 103.111
R23046 CSoutput.n279 CSoutput.n278 103.111
R23047 CSoutput.n112 CSoutput.n111 103.111
R23048 CSoutput.n114 CSoutput.n113 103.111
R23049 CSoutput.n116 CSoutput.n115 103.111
R23050 CSoutput.n118 CSoutput.n117 103.111
R23051 CSoutput.n120 CSoutput.n119 103.111
R23052 CSoutput.n122 CSoutput.n121 103.111
R23053 CSoutput.n124 CSoutput.n123 103.111
R23054 CSoutput.n96 CSoutput.n95 103.111
R23055 CSoutput.n98 CSoutput.n97 103.111
R23056 CSoutput.n100 CSoutput.n99 103.111
R23057 CSoutput.n102 CSoutput.n101 103.111
R23058 CSoutput.n104 CSoutput.n103 103.111
R23059 CSoutput.n106 CSoutput.n105 103.111
R23060 CSoutput.n108 CSoutput.n107 103.111
R23061 CSoutput.n81 CSoutput.n80 103.111
R23062 CSoutput.n83 CSoutput.n82 103.111
R23063 CSoutput.n85 CSoutput.n84 103.111
R23064 CSoutput.n87 CSoutput.n86 103.111
R23065 CSoutput.n89 CSoutput.n88 103.111
R23066 CSoutput.n91 CSoutput.n90 103.111
R23067 CSoutput.n93 CSoutput.n92 103.111
R23068 CSoutput.n322 CSoutput.n321 103.111
R23069 CSoutput.n366 CSoutput.n364 81.5057
R23070 CSoutput.n346 CSoutput.n344 81.5057
R23071 CSoutput.n327 CSoutput.n325 81.5057
R23072 CSoutput.n426 CSoutput.n424 81.5057
R23073 CSoutput.n406 CSoutput.n404 81.5057
R23074 CSoutput.n387 CSoutput.n385 81.5057
R23075 CSoutput.n382 CSoutput.n381 80.9324
R23076 CSoutput.n380 CSoutput.n379 80.9324
R23077 CSoutput.n378 CSoutput.n377 80.9324
R23078 CSoutput.n376 CSoutput.n375 80.9324
R23079 CSoutput.n374 CSoutput.n373 80.9324
R23080 CSoutput.n372 CSoutput.n371 80.9324
R23081 CSoutput.n370 CSoutput.n369 80.9324
R23082 CSoutput.n368 CSoutput.n367 80.9324
R23083 CSoutput.n366 CSoutput.n365 80.9324
R23084 CSoutput.n362 CSoutput.n361 80.9324
R23085 CSoutput.n360 CSoutput.n359 80.9324
R23086 CSoutput.n358 CSoutput.n357 80.9324
R23087 CSoutput.n356 CSoutput.n355 80.9324
R23088 CSoutput.n354 CSoutput.n353 80.9324
R23089 CSoutput.n352 CSoutput.n351 80.9324
R23090 CSoutput.n350 CSoutput.n349 80.9324
R23091 CSoutput.n348 CSoutput.n347 80.9324
R23092 CSoutput.n346 CSoutput.n345 80.9324
R23093 CSoutput.n343 CSoutput.n342 80.9324
R23094 CSoutput.n341 CSoutput.n340 80.9324
R23095 CSoutput.n339 CSoutput.n338 80.9324
R23096 CSoutput.n337 CSoutput.n336 80.9324
R23097 CSoutput.n335 CSoutput.n334 80.9324
R23098 CSoutput.n333 CSoutput.n332 80.9324
R23099 CSoutput.n331 CSoutput.n330 80.9324
R23100 CSoutput.n329 CSoutput.n328 80.9324
R23101 CSoutput.n327 CSoutput.n326 80.9324
R23102 CSoutput.n426 CSoutput.n425 80.9324
R23103 CSoutput.n428 CSoutput.n427 80.9324
R23104 CSoutput.n430 CSoutput.n429 80.9324
R23105 CSoutput.n432 CSoutput.n431 80.9324
R23106 CSoutput.n434 CSoutput.n433 80.9324
R23107 CSoutput.n436 CSoutput.n435 80.9324
R23108 CSoutput.n438 CSoutput.n437 80.9324
R23109 CSoutput.n440 CSoutput.n439 80.9324
R23110 CSoutput.n442 CSoutput.n441 80.9324
R23111 CSoutput.n406 CSoutput.n405 80.9324
R23112 CSoutput.n408 CSoutput.n407 80.9324
R23113 CSoutput.n410 CSoutput.n409 80.9324
R23114 CSoutput.n412 CSoutput.n411 80.9324
R23115 CSoutput.n414 CSoutput.n413 80.9324
R23116 CSoutput.n416 CSoutput.n415 80.9324
R23117 CSoutput.n418 CSoutput.n417 80.9324
R23118 CSoutput.n420 CSoutput.n419 80.9324
R23119 CSoutput.n422 CSoutput.n421 80.9324
R23120 CSoutput.n387 CSoutput.n386 80.9324
R23121 CSoutput.n389 CSoutput.n388 80.9324
R23122 CSoutput.n391 CSoutput.n390 80.9324
R23123 CSoutput.n393 CSoutput.n392 80.9324
R23124 CSoutput.n395 CSoutput.n394 80.9324
R23125 CSoutput.n397 CSoutput.n396 80.9324
R23126 CSoutput.n399 CSoutput.n398 80.9324
R23127 CSoutput.n401 CSoutput.n400 80.9324
R23128 CSoutput.n403 CSoutput.n402 80.9324
R23129 CSoutput.n25 CSoutput.n24 48.1486
R23130 CSoutput.n69 CSoutput.n3 48.1486
R23131 CSoutput.n38 CSoutput.n37 48.1486
R23132 CSoutput.n42 CSoutput.n41 48.1486
R23133 CSoutput.n51 CSoutput.n50 48.1486
R23134 CSoutput.n55 CSoutput.n54 48.1486
R23135 CSoutput.n22 CSoutput.n17 46.462
R23136 CSoutput.n72 CSoutput.n71 46.462
R23137 CSoutput.n20 CSoutput.n19 44.9055
R23138 CSoutput.n29 CSoutput.n28 43.7635
R23139 CSoutput.n65 CSoutput.n63 43.7635
R23140 CSoutput.n35 CSoutput.n13 41.7396
R23141 CSoutput.n57 CSoutput.n5 41.7396
R23142 CSoutput.n44 CSoutput.n9 37.0171
R23143 CSoutput.n48 CSoutput.n9 37.0171
R23144 CSoutput.n76 CSoutput.n75 34.9932
R23145 CSoutput.n31 CSoutput.n13 32.2947
R23146 CSoutput.n61 CSoutput.n5 32.2947
R23147 CSoutput.n30 CSoutput.n29 29.6014
R23148 CSoutput.n63 CSoutput.n62 29.6014
R23149 CSoutput.n19 CSoutput.n18 28.4085
R23150 CSoutput.n18 CSoutput.n17 25.1176
R23151 CSoutput.n72 CSoutput.n1 25.1176
R23152 CSoutput.n43 CSoutput.n42 22.0922
R23153 CSoutput.n50 CSoutput.n49 22.0922
R23154 CSoutput.n77 CSoutput.n76 21.8586
R23155 CSoutput.n37 CSoutput.n36 18.9681
R23156 CSoutput.n56 CSoutput.n55 18.9681
R23157 CSoutput.n25 CSoutput.n15 17.6292
R23158 CSoutput.n64 CSoutput.n3 17.6292
R23159 CSoutput.n24 CSoutput.n23 15.844
R23160 CSoutput.n70 CSoutput.n69 15.844
R23161 CSoutput.n38 CSoutput.n11 14.5051
R23162 CSoutput.n54 CSoutput.n7 14.5051
R23163 CSoutput.n445 CSoutput.n78 11.4982
R23164 CSoutput.n41 CSoutput.n11 11.3811
R23165 CSoutput.n51 CSoutput.n7 11.3811
R23166 CSoutput.n23 CSoutput.n22 10.0422
R23167 CSoutput.n71 CSoutput.n70 10.0422
R23168 CSoutput.n307 CSoutput.n291 9.25285
R23169 CSoutput.n109 CSoutput.n93 9.25285
R23170 CSoutput.n363 CSoutput.n343 8.98182
R23171 CSoutput.n423 CSoutput.n403 8.98182
R23172 CSoutput.n384 CSoutput.n324 8.74155
R23173 CSoutput.n28 CSoutput.n15 8.25698
R23174 CSoutput.n65 CSoutput.n64 8.25698
R23175 CSoutput.n324 CSoutput.n323 7.12641
R23176 CSoutput.n126 CSoutput.n125 7.12641
R23177 CSoutput.n36 CSoutput.n35 6.91809
R23178 CSoutput.n57 CSoutput.n56 6.91809
R23179 CSoutput.n384 CSoutput.n383 6.02792
R23180 CSoutput.n444 CSoutput.n443 6.02792
R23181 CSoutput.n383 CSoutput.n382 5.25266
R23182 CSoutput.n363 CSoutput.n362 5.25266
R23183 CSoutput.n443 CSoutput.n442 5.25266
R23184 CSoutput.n423 CSoutput.n422 5.25266
R23185 CSoutput.n445 CSoutput.n126 5.14911
R23186 CSoutput.n323 CSoutput.n322 5.1449
R23187 CSoutput.n307 CSoutput.n306 5.1449
R23188 CSoutput.n125 CSoutput.n124 5.1449
R23189 CSoutput.n109 CSoutput.n108 5.1449
R23190 CSoutput.n217 CSoutput.n170 4.5005
R23191 CSoutput.n186 CSoutput.n170 4.5005
R23192 CSoutput.n181 CSoutput.n165 4.5005
R23193 CSoutput.n181 CSoutput.n167 4.5005
R23194 CSoutput.n181 CSoutput.n164 4.5005
R23195 CSoutput.n181 CSoutput.n168 4.5005
R23196 CSoutput.n181 CSoutput.n163 4.5005
R23197 CSoutput.n181 CSoutput.t237 4.5005
R23198 CSoutput.n181 CSoutput.n162 4.5005
R23199 CSoutput.n181 CSoutput.n169 4.5005
R23200 CSoutput.n181 CSoutput.n170 4.5005
R23201 CSoutput.n179 CSoutput.n165 4.5005
R23202 CSoutput.n179 CSoutput.n167 4.5005
R23203 CSoutput.n179 CSoutput.n164 4.5005
R23204 CSoutput.n179 CSoutput.n168 4.5005
R23205 CSoutput.n179 CSoutput.n163 4.5005
R23206 CSoutput.n179 CSoutput.t237 4.5005
R23207 CSoutput.n179 CSoutput.n162 4.5005
R23208 CSoutput.n179 CSoutput.n169 4.5005
R23209 CSoutput.n179 CSoutput.n170 4.5005
R23210 CSoutput.n178 CSoutput.n165 4.5005
R23211 CSoutput.n178 CSoutput.n167 4.5005
R23212 CSoutput.n178 CSoutput.n164 4.5005
R23213 CSoutput.n178 CSoutput.n168 4.5005
R23214 CSoutput.n178 CSoutput.n163 4.5005
R23215 CSoutput.n178 CSoutput.t237 4.5005
R23216 CSoutput.n178 CSoutput.n162 4.5005
R23217 CSoutput.n178 CSoutput.n169 4.5005
R23218 CSoutput.n178 CSoutput.n170 4.5005
R23219 CSoutput.n263 CSoutput.n165 4.5005
R23220 CSoutput.n263 CSoutput.n167 4.5005
R23221 CSoutput.n263 CSoutput.n164 4.5005
R23222 CSoutput.n263 CSoutput.n168 4.5005
R23223 CSoutput.n263 CSoutput.n163 4.5005
R23224 CSoutput.n263 CSoutput.t237 4.5005
R23225 CSoutput.n263 CSoutput.n162 4.5005
R23226 CSoutput.n263 CSoutput.n169 4.5005
R23227 CSoutput.n263 CSoutput.n170 4.5005
R23228 CSoutput.n261 CSoutput.n165 4.5005
R23229 CSoutput.n261 CSoutput.n167 4.5005
R23230 CSoutput.n261 CSoutput.n164 4.5005
R23231 CSoutput.n261 CSoutput.n168 4.5005
R23232 CSoutput.n261 CSoutput.n163 4.5005
R23233 CSoutput.n261 CSoutput.t237 4.5005
R23234 CSoutput.n261 CSoutput.n162 4.5005
R23235 CSoutput.n261 CSoutput.n169 4.5005
R23236 CSoutput.n259 CSoutput.n165 4.5005
R23237 CSoutput.n259 CSoutput.n167 4.5005
R23238 CSoutput.n259 CSoutput.n164 4.5005
R23239 CSoutput.n259 CSoutput.n168 4.5005
R23240 CSoutput.n259 CSoutput.n163 4.5005
R23241 CSoutput.n259 CSoutput.t237 4.5005
R23242 CSoutput.n259 CSoutput.n162 4.5005
R23243 CSoutput.n259 CSoutput.n169 4.5005
R23244 CSoutput.n189 CSoutput.n165 4.5005
R23245 CSoutput.n189 CSoutput.n167 4.5005
R23246 CSoutput.n189 CSoutput.n164 4.5005
R23247 CSoutput.n189 CSoutput.n168 4.5005
R23248 CSoutput.n189 CSoutput.n163 4.5005
R23249 CSoutput.n189 CSoutput.t237 4.5005
R23250 CSoutput.n189 CSoutput.n162 4.5005
R23251 CSoutput.n189 CSoutput.n169 4.5005
R23252 CSoutput.n189 CSoutput.n170 4.5005
R23253 CSoutput.n188 CSoutput.n165 4.5005
R23254 CSoutput.n188 CSoutput.n167 4.5005
R23255 CSoutput.n188 CSoutput.n164 4.5005
R23256 CSoutput.n188 CSoutput.n168 4.5005
R23257 CSoutput.n188 CSoutput.n163 4.5005
R23258 CSoutput.n188 CSoutput.t237 4.5005
R23259 CSoutput.n188 CSoutput.n162 4.5005
R23260 CSoutput.n188 CSoutput.n169 4.5005
R23261 CSoutput.n188 CSoutput.n170 4.5005
R23262 CSoutput.n192 CSoutput.n165 4.5005
R23263 CSoutput.n192 CSoutput.n167 4.5005
R23264 CSoutput.n192 CSoutput.n164 4.5005
R23265 CSoutput.n192 CSoutput.n168 4.5005
R23266 CSoutput.n192 CSoutput.n163 4.5005
R23267 CSoutput.n192 CSoutput.t237 4.5005
R23268 CSoutput.n192 CSoutput.n162 4.5005
R23269 CSoutput.n192 CSoutput.n169 4.5005
R23270 CSoutput.n192 CSoutput.n170 4.5005
R23271 CSoutput.n191 CSoutput.n165 4.5005
R23272 CSoutput.n191 CSoutput.n167 4.5005
R23273 CSoutput.n191 CSoutput.n164 4.5005
R23274 CSoutput.n191 CSoutput.n168 4.5005
R23275 CSoutput.n191 CSoutput.n163 4.5005
R23276 CSoutput.n191 CSoutput.t237 4.5005
R23277 CSoutput.n191 CSoutput.n162 4.5005
R23278 CSoutput.n191 CSoutput.n169 4.5005
R23279 CSoutput.n191 CSoutput.n170 4.5005
R23280 CSoutput.n174 CSoutput.n165 4.5005
R23281 CSoutput.n174 CSoutput.n167 4.5005
R23282 CSoutput.n174 CSoutput.n164 4.5005
R23283 CSoutput.n174 CSoutput.n168 4.5005
R23284 CSoutput.n174 CSoutput.n163 4.5005
R23285 CSoutput.n174 CSoutput.t237 4.5005
R23286 CSoutput.n174 CSoutput.n162 4.5005
R23287 CSoutput.n174 CSoutput.n169 4.5005
R23288 CSoutput.n174 CSoutput.n170 4.5005
R23289 CSoutput.n266 CSoutput.n165 4.5005
R23290 CSoutput.n266 CSoutput.n167 4.5005
R23291 CSoutput.n266 CSoutput.n164 4.5005
R23292 CSoutput.n266 CSoutput.n168 4.5005
R23293 CSoutput.n266 CSoutput.n163 4.5005
R23294 CSoutput.n266 CSoutput.t237 4.5005
R23295 CSoutput.n266 CSoutput.n162 4.5005
R23296 CSoutput.n266 CSoutput.n169 4.5005
R23297 CSoutput.n266 CSoutput.n170 4.5005
R23298 CSoutput.n253 CSoutput.n224 4.5005
R23299 CSoutput.n253 CSoutput.n230 4.5005
R23300 CSoutput.n211 CSoutput.n200 4.5005
R23301 CSoutput.n211 CSoutput.n202 4.5005
R23302 CSoutput.n211 CSoutput.n199 4.5005
R23303 CSoutput.n211 CSoutput.n203 4.5005
R23304 CSoutput.n211 CSoutput.n198 4.5005
R23305 CSoutput.n211 CSoutput.t232 4.5005
R23306 CSoutput.n211 CSoutput.n197 4.5005
R23307 CSoutput.n211 CSoutput.n204 4.5005
R23308 CSoutput.n253 CSoutput.n211 4.5005
R23309 CSoutput.n232 CSoutput.n200 4.5005
R23310 CSoutput.n232 CSoutput.n202 4.5005
R23311 CSoutput.n232 CSoutput.n199 4.5005
R23312 CSoutput.n232 CSoutput.n203 4.5005
R23313 CSoutput.n232 CSoutput.n198 4.5005
R23314 CSoutput.n232 CSoutput.t232 4.5005
R23315 CSoutput.n232 CSoutput.n197 4.5005
R23316 CSoutput.n232 CSoutput.n204 4.5005
R23317 CSoutput.n253 CSoutput.n232 4.5005
R23318 CSoutput.n210 CSoutput.n200 4.5005
R23319 CSoutput.n210 CSoutput.n202 4.5005
R23320 CSoutput.n210 CSoutput.n199 4.5005
R23321 CSoutput.n210 CSoutput.n203 4.5005
R23322 CSoutput.n210 CSoutput.n198 4.5005
R23323 CSoutput.n210 CSoutput.t232 4.5005
R23324 CSoutput.n210 CSoutput.n197 4.5005
R23325 CSoutput.n210 CSoutput.n204 4.5005
R23326 CSoutput.n253 CSoutput.n210 4.5005
R23327 CSoutput.n234 CSoutput.n200 4.5005
R23328 CSoutput.n234 CSoutput.n202 4.5005
R23329 CSoutput.n234 CSoutput.n199 4.5005
R23330 CSoutput.n234 CSoutput.n203 4.5005
R23331 CSoutput.n234 CSoutput.n198 4.5005
R23332 CSoutput.n234 CSoutput.t232 4.5005
R23333 CSoutput.n234 CSoutput.n197 4.5005
R23334 CSoutput.n234 CSoutput.n204 4.5005
R23335 CSoutput.n253 CSoutput.n234 4.5005
R23336 CSoutput.n200 CSoutput.n195 4.5005
R23337 CSoutput.n202 CSoutput.n195 4.5005
R23338 CSoutput.n199 CSoutput.n195 4.5005
R23339 CSoutput.n203 CSoutput.n195 4.5005
R23340 CSoutput.n198 CSoutput.n195 4.5005
R23341 CSoutput.t232 CSoutput.n195 4.5005
R23342 CSoutput.n197 CSoutput.n195 4.5005
R23343 CSoutput.n204 CSoutput.n195 4.5005
R23344 CSoutput.n256 CSoutput.n200 4.5005
R23345 CSoutput.n256 CSoutput.n202 4.5005
R23346 CSoutput.n256 CSoutput.n199 4.5005
R23347 CSoutput.n256 CSoutput.n203 4.5005
R23348 CSoutput.n256 CSoutput.n198 4.5005
R23349 CSoutput.n256 CSoutput.t232 4.5005
R23350 CSoutput.n256 CSoutput.n197 4.5005
R23351 CSoutput.n256 CSoutput.n204 4.5005
R23352 CSoutput.n254 CSoutput.n200 4.5005
R23353 CSoutput.n254 CSoutput.n202 4.5005
R23354 CSoutput.n254 CSoutput.n199 4.5005
R23355 CSoutput.n254 CSoutput.n203 4.5005
R23356 CSoutput.n254 CSoutput.n198 4.5005
R23357 CSoutput.n254 CSoutput.t232 4.5005
R23358 CSoutput.n254 CSoutput.n197 4.5005
R23359 CSoutput.n254 CSoutput.n204 4.5005
R23360 CSoutput.n254 CSoutput.n253 4.5005
R23361 CSoutput.n236 CSoutput.n200 4.5005
R23362 CSoutput.n236 CSoutput.n202 4.5005
R23363 CSoutput.n236 CSoutput.n199 4.5005
R23364 CSoutput.n236 CSoutput.n203 4.5005
R23365 CSoutput.n236 CSoutput.n198 4.5005
R23366 CSoutput.n236 CSoutput.t232 4.5005
R23367 CSoutput.n236 CSoutput.n197 4.5005
R23368 CSoutput.n236 CSoutput.n204 4.5005
R23369 CSoutput.n253 CSoutput.n236 4.5005
R23370 CSoutput.n208 CSoutput.n200 4.5005
R23371 CSoutput.n208 CSoutput.n202 4.5005
R23372 CSoutput.n208 CSoutput.n199 4.5005
R23373 CSoutput.n208 CSoutput.n203 4.5005
R23374 CSoutput.n208 CSoutput.n198 4.5005
R23375 CSoutput.n208 CSoutput.t232 4.5005
R23376 CSoutput.n208 CSoutput.n197 4.5005
R23377 CSoutput.n208 CSoutput.n204 4.5005
R23378 CSoutput.n253 CSoutput.n208 4.5005
R23379 CSoutput.n238 CSoutput.n200 4.5005
R23380 CSoutput.n238 CSoutput.n202 4.5005
R23381 CSoutput.n238 CSoutput.n199 4.5005
R23382 CSoutput.n238 CSoutput.n203 4.5005
R23383 CSoutput.n238 CSoutput.n198 4.5005
R23384 CSoutput.n238 CSoutput.t232 4.5005
R23385 CSoutput.n238 CSoutput.n197 4.5005
R23386 CSoutput.n238 CSoutput.n204 4.5005
R23387 CSoutput.n253 CSoutput.n238 4.5005
R23388 CSoutput.n207 CSoutput.n200 4.5005
R23389 CSoutput.n207 CSoutput.n202 4.5005
R23390 CSoutput.n207 CSoutput.n199 4.5005
R23391 CSoutput.n207 CSoutput.n203 4.5005
R23392 CSoutput.n207 CSoutput.n198 4.5005
R23393 CSoutput.n207 CSoutput.t232 4.5005
R23394 CSoutput.n207 CSoutput.n197 4.5005
R23395 CSoutput.n207 CSoutput.n204 4.5005
R23396 CSoutput.n253 CSoutput.n207 4.5005
R23397 CSoutput.n252 CSoutput.n200 4.5005
R23398 CSoutput.n252 CSoutput.n202 4.5005
R23399 CSoutput.n252 CSoutput.n199 4.5005
R23400 CSoutput.n252 CSoutput.n203 4.5005
R23401 CSoutput.n252 CSoutput.n198 4.5005
R23402 CSoutput.n252 CSoutput.t232 4.5005
R23403 CSoutput.n252 CSoutput.n197 4.5005
R23404 CSoutput.n252 CSoutput.n204 4.5005
R23405 CSoutput.n253 CSoutput.n252 4.5005
R23406 CSoutput.n251 CSoutput.n136 4.5005
R23407 CSoutput.n152 CSoutput.n136 4.5005
R23408 CSoutput.n147 CSoutput.n131 4.5005
R23409 CSoutput.n147 CSoutput.n133 4.5005
R23410 CSoutput.n147 CSoutput.n130 4.5005
R23411 CSoutput.n147 CSoutput.n134 4.5005
R23412 CSoutput.n147 CSoutput.n129 4.5005
R23413 CSoutput.n147 CSoutput.t230 4.5005
R23414 CSoutput.n147 CSoutput.n128 4.5005
R23415 CSoutput.n147 CSoutput.n135 4.5005
R23416 CSoutput.n147 CSoutput.n136 4.5005
R23417 CSoutput.n145 CSoutput.n131 4.5005
R23418 CSoutput.n145 CSoutput.n133 4.5005
R23419 CSoutput.n145 CSoutput.n130 4.5005
R23420 CSoutput.n145 CSoutput.n134 4.5005
R23421 CSoutput.n145 CSoutput.n129 4.5005
R23422 CSoutput.n145 CSoutput.t230 4.5005
R23423 CSoutput.n145 CSoutput.n128 4.5005
R23424 CSoutput.n145 CSoutput.n135 4.5005
R23425 CSoutput.n145 CSoutput.n136 4.5005
R23426 CSoutput.n144 CSoutput.n131 4.5005
R23427 CSoutput.n144 CSoutput.n133 4.5005
R23428 CSoutput.n144 CSoutput.n130 4.5005
R23429 CSoutput.n144 CSoutput.n134 4.5005
R23430 CSoutput.n144 CSoutput.n129 4.5005
R23431 CSoutput.n144 CSoutput.t230 4.5005
R23432 CSoutput.n144 CSoutput.n128 4.5005
R23433 CSoutput.n144 CSoutput.n135 4.5005
R23434 CSoutput.n144 CSoutput.n136 4.5005
R23435 CSoutput.n273 CSoutput.n131 4.5005
R23436 CSoutput.n273 CSoutput.n133 4.5005
R23437 CSoutput.n273 CSoutput.n130 4.5005
R23438 CSoutput.n273 CSoutput.n134 4.5005
R23439 CSoutput.n273 CSoutput.n129 4.5005
R23440 CSoutput.n273 CSoutput.t230 4.5005
R23441 CSoutput.n273 CSoutput.n128 4.5005
R23442 CSoutput.n273 CSoutput.n135 4.5005
R23443 CSoutput.n273 CSoutput.n136 4.5005
R23444 CSoutput.n271 CSoutput.n131 4.5005
R23445 CSoutput.n271 CSoutput.n133 4.5005
R23446 CSoutput.n271 CSoutput.n130 4.5005
R23447 CSoutput.n271 CSoutput.n134 4.5005
R23448 CSoutput.n271 CSoutput.n129 4.5005
R23449 CSoutput.n271 CSoutput.t230 4.5005
R23450 CSoutput.n271 CSoutput.n128 4.5005
R23451 CSoutput.n271 CSoutput.n135 4.5005
R23452 CSoutput.n269 CSoutput.n131 4.5005
R23453 CSoutput.n269 CSoutput.n133 4.5005
R23454 CSoutput.n269 CSoutput.n130 4.5005
R23455 CSoutput.n269 CSoutput.n134 4.5005
R23456 CSoutput.n269 CSoutput.n129 4.5005
R23457 CSoutput.n269 CSoutput.t230 4.5005
R23458 CSoutput.n269 CSoutput.n128 4.5005
R23459 CSoutput.n269 CSoutput.n135 4.5005
R23460 CSoutput.n155 CSoutput.n131 4.5005
R23461 CSoutput.n155 CSoutput.n133 4.5005
R23462 CSoutput.n155 CSoutput.n130 4.5005
R23463 CSoutput.n155 CSoutput.n134 4.5005
R23464 CSoutput.n155 CSoutput.n129 4.5005
R23465 CSoutput.n155 CSoutput.t230 4.5005
R23466 CSoutput.n155 CSoutput.n128 4.5005
R23467 CSoutput.n155 CSoutput.n135 4.5005
R23468 CSoutput.n155 CSoutput.n136 4.5005
R23469 CSoutput.n154 CSoutput.n131 4.5005
R23470 CSoutput.n154 CSoutput.n133 4.5005
R23471 CSoutput.n154 CSoutput.n130 4.5005
R23472 CSoutput.n154 CSoutput.n134 4.5005
R23473 CSoutput.n154 CSoutput.n129 4.5005
R23474 CSoutput.n154 CSoutput.t230 4.5005
R23475 CSoutput.n154 CSoutput.n128 4.5005
R23476 CSoutput.n154 CSoutput.n135 4.5005
R23477 CSoutput.n154 CSoutput.n136 4.5005
R23478 CSoutput.n158 CSoutput.n131 4.5005
R23479 CSoutput.n158 CSoutput.n133 4.5005
R23480 CSoutput.n158 CSoutput.n130 4.5005
R23481 CSoutput.n158 CSoutput.n134 4.5005
R23482 CSoutput.n158 CSoutput.n129 4.5005
R23483 CSoutput.n158 CSoutput.t230 4.5005
R23484 CSoutput.n158 CSoutput.n128 4.5005
R23485 CSoutput.n158 CSoutput.n135 4.5005
R23486 CSoutput.n158 CSoutput.n136 4.5005
R23487 CSoutput.n157 CSoutput.n131 4.5005
R23488 CSoutput.n157 CSoutput.n133 4.5005
R23489 CSoutput.n157 CSoutput.n130 4.5005
R23490 CSoutput.n157 CSoutput.n134 4.5005
R23491 CSoutput.n157 CSoutput.n129 4.5005
R23492 CSoutput.n157 CSoutput.t230 4.5005
R23493 CSoutput.n157 CSoutput.n128 4.5005
R23494 CSoutput.n157 CSoutput.n135 4.5005
R23495 CSoutput.n157 CSoutput.n136 4.5005
R23496 CSoutput.n140 CSoutput.n131 4.5005
R23497 CSoutput.n140 CSoutput.n133 4.5005
R23498 CSoutput.n140 CSoutput.n130 4.5005
R23499 CSoutput.n140 CSoutput.n134 4.5005
R23500 CSoutput.n140 CSoutput.n129 4.5005
R23501 CSoutput.n140 CSoutput.t230 4.5005
R23502 CSoutput.n140 CSoutput.n128 4.5005
R23503 CSoutput.n140 CSoutput.n135 4.5005
R23504 CSoutput.n140 CSoutput.n136 4.5005
R23505 CSoutput.n276 CSoutput.n131 4.5005
R23506 CSoutput.n276 CSoutput.n133 4.5005
R23507 CSoutput.n276 CSoutput.n130 4.5005
R23508 CSoutput.n276 CSoutput.n134 4.5005
R23509 CSoutput.n276 CSoutput.n129 4.5005
R23510 CSoutput.n276 CSoutput.t230 4.5005
R23511 CSoutput.n276 CSoutput.n128 4.5005
R23512 CSoutput.n276 CSoutput.n135 4.5005
R23513 CSoutput.n276 CSoutput.n136 4.5005
R23514 CSoutput.n323 CSoutput.n307 4.10845
R23515 CSoutput.n125 CSoutput.n109 4.10845
R23516 CSoutput.n321 CSoutput.t144 4.06363
R23517 CSoutput.n321 CSoutput.t148 4.06363
R23518 CSoutput.n319 CSoutput.t140 4.06363
R23519 CSoutput.n319 CSoutput.t132 4.06363
R23520 CSoutput.n317 CSoutput.t204 4.06363
R23521 CSoutput.n317 CSoutput.t157 4.06363
R23522 CSoutput.n315 CSoutput.t201 4.06363
R23523 CSoutput.n315 CSoutput.t190 4.06363
R23524 CSoutput.n313 CSoutput.t164 4.06363
R23525 CSoutput.n313 CSoutput.t162 4.06363
R23526 CSoutput.n311 CSoutput.t173 4.06363
R23527 CSoutput.n311 CSoutput.t215 4.06363
R23528 CSoutput.n309 CSoutput.t203 4.06363
R23529 CSoutput.n309 CSoutput.t135 4.06363
R23530 CSoutput.n308 CSoutput.t145 4.06363
R23531 CSoutput.n308 CSoutput.t199 4.06363
R23532 CSoutput.n305 CSoutput.t212 4.06363
R23533 CSoutput.n305 CSoutput.t156 4.06363
R23534 CSoutput.n303 CSoutput.t202 4.06363
R23535 CSoutput.n303 CSoutput.t186 4.06363
R23536 CSoutput.n301 CSoutput.t161 4.06363
R23537 CSoutput.n301 CSoutput.t3 4.06363
R23538 CSoutput.n299 CSoutput.t172 4.06363
R23539 CSoutput.n299 CSoutput.t137 4.06363
R23540 CSoutput.n297 CSoutput.t152 4.06363
R23541 CSoutput.n297 CSoutput.t160 4.06363
R23542 CSoutput.n295 CSoutput.t179 4.06363
R23543 CSoutput.n295 CSoutput.t158 4.06363
R23544 CSoutput.n293 CSoutput.t139 4.06363
R23545 CSoutput.n293 CSoutput.t211 4.06363
R23546 CSoutput.n292 CSoutput.t213 4.06363
R23547 CSoutput.n292 CSoutput.t207 4.06363
R23548 CSoutput.n290 CSoutput.t198 4.06363
R23549 CSoutput.n290 CSoutput.t165 4.06363
R23550 CSoutput.n288 CSoutput.t167 4.06363
R23551 CSoutput.n288 CSoutput.t195 4.06363
R23552 CSoutput.n286 CSoutput.t155 4.06363
R23553 CSoutput.n286 CSoutput.t209 4.06363
R23554 CSoutput.n284 CSoutput.t189 4.06363
R23555 CSoutput.n284 CSoutput.t0 4.06363
R23556 CSoutput.n282 CSoutput.t163 4.06363
R23557 CSoutput.n282 CSoutput.t168 4.06363
R23558 CSoutput.n280 CSoutput.t192 4.06363
R23559 CSoutput.n280 CSoutput.t146 4.06363
R23560 CSoutput.n278 CSoutput.t134 4.06363
R23561 CSoutput.n278 CSoutput.t127 4.06363
R23562 CSoutput.n277 CSoutput.t175 4.06363
R23563 CSoutput.n277 CSoutput.t151 4.06363
R23564 CSoutput.n110 CSoutput.t142 4.06363
R23565 CSoutput.n110 CSoutput.t169 4.06363
R23566 CSoutput.n111 CSoutput.t147 4.06363
R23567 CSoutput.n111 CSoutput.t133 4.06363
R23568 CSoutput.n113 CSoutput.t170 4.06363
R23569 CSoutput.n113 CSoutput.t136 4.06363
R23570 CSoutput.n115 CSoutput.t128 4.06363
R23571 CSoutput.n115 CSoutput.t129 4.06363
R23572 CSoutput.n117 CSoutput.t205 4.06363
R23573 CSoutput.n117 CSoutput.t153 4.06363
R23574 CSoutput.n119 CSoutput.t191 4.06363
R23575 CSoutput.n119 CSoutput.t138 4.06363
R23576 CSoutput.n121 CSoutput.t180 4.06363
R23577 CSoutput.n121 CSoutput.t210 4.06363
R23578 CSoutput.n123 CSoutput.t143 4.06363
R23579 CSoutput.n123 CSoutput.t184 4.06363
R23580 CSoutput.n94 CSoutput.t130 4.06363
R23581 CSoutput.n94 CSoutput.t183 4.06363
R23582 CSoutput.n95 CSoutput.t159 4.06363
R23583 CSoutput.n95 CSoutput.t176 4.06363
R23584 CSoutput.n97 CSoutput.t1 4.06363
R23585 CSoutput.n97 CSoutput.t214 4.06363
R23586 CSoutput.n99 CSoutput.t200 4.06363
R23587 CSoutput.n99 CSoutput.t124 4.06363
R23588 CSoutput.n101 CSoutput.t196 4.06363
R23589 CSoutput.n101 CSoutput.t185 4.06363
R23590 CSoutput.n103 CSoutput.t208 4.06363
R23591 CSoutput.n103 CSoutput.t125 4.06363
R23592 CSoutput.n105 CSoutput.t206 4.06363
R23593 CSoutput.n105 CSoutput.t193 4.06363
R23594 CSoutput.n107 CSoutput.t177 4.06363
R23595 CSoutput.n107 CSoutput.t182 4.06363
R23596 CSoutput.n79 CSoutput.t2 4.06363
R23597 CSoutput.n79 CSoutput.t174 4.06363
R23598 CSoutput.n80 CSoutput.t126 4.06363
R23599 CSoutput.n80 CSoutput.t178 4.06363
R23600 CSoutput.n82 CSoutput.t149 4.06363
R23601 CSoutput.n82 CSoutput.t197 4.06363
R23602 CSoutput.n84 CSoutput.t141 4.06363
R23603 CSoutput.n84 CSoutput.t187 4.06363
R23604 CSoutput.n86 CSoutput.t131 4.06363
R23605 CSoutput.n86 CSoutput.t188 4.06363
R23606 CSoutput.n88 CSoutput.t150 4.06363
R23607 CSoutput.n88 CSoutput.t154 4.06363
R23608 CSoutput.n90 CSoutput.t194 4.06363
R23609 CSoutput.n90 CSoutput.t166 4.06363
R23610 CSoutput.n92 CSoutput.t171 4.06363
R23611 CSoutput.n92 CSoutput.t181 4.06363
R23612 CSoutput.n44 CSoutput.n43 3.79402
R23613 CSoutput.n49 CSoutput.n48 3.79402
R23614 CSoutput.n383 CSoutput.n363 3.72967
R23615 CSoutput.n443 CSoutput.n423 3.72967
R23616 CSoutput.n445 CSoutput.n444 3.57343
R23617 CSoutput.n444 CSoutput.n384 3.42304
R23618 CSoutput.n324 CSoutput.n126 2.99158
R23619 CSoutput.n381 CSoutput.t53 2.82907
R23620 CSoutput.n381 CSoutput.t19 2.82907
R23621 CSoutput.n379 CSoutput.t4 2.82907
R23622 CSoutput.n379 CSoutput.t48 2.82907
R23623 CSoutput.n377 CSoutput.t38 2.82907
R23624 CSoutput.n377 CSoutput.t28 2.82907
R23625 CSoutput.n375 CSoutput.t16 2.82907
R23626 CSoutput.n375 CSoutput.t107 2.82907
R23627 CSoutput.n373 CSoutput.t31 2.82907
R23628 CSoutput.n373 CSoutput.t35 2.82907
R23629 CSoutput.n371 CSoutput.t30 2.82907
R23630 CSoutput.n371 CSoutput.t123 2.82907
R23631 CSoutput.n369 CSoutput.t54 2.82907
R23632 CSoutput.n369 CSoutput.t21 2.82907
R23633 CSoutput.n367 CSoutput.t9 2.82907
R23634 CSoutput.n367 CSoutput.t93 2.82907
R23635 CSoutput.n365 CSoutput.t40 2.82907
R23636 CSoutput.n365 CSoutput.t46 2.82907
R23637 CSoutput.n364 CSoutput.t20 2.82907
R23638 CSoutput.n364 CSoutput.t111 2.82907
R23639 CSoutput.n361 CSoutput.t56 2.82907
R23640 CSoutput.n361 CSoutput.t69 2.82907
R23641 CSoutput.n359 CSoutput.t74 2.82907
R23642 CSoutput.n359 CSoutput.t78 2.82907
R23643 CSoutput.n357 CSoutput.t89 2.82907
R23644 CSoutput.n357 CSoutput.t64 2.82907
R23645 CSoutput.n355 CSoutput.t65 2.82907
R23646 CSoutput.n355 CSoutput.t73 2.82907
R23647 CSoutput.n353 CSoutput.t8 2.82907
R23648 CSoutput.n353 CSoutput.t90 2.82907
R23649 CSoutput.n351 CSoutput.t88 2.82907
R23650 CSoutput.n351 CSoutput.t62 2.82907
R23651 CSoutput.n349 CSoutput.t109 2.82907
R23652 CSoutput.n349 CSoutput.t6 2.82907
R23653 CSoutput.n347 CSoutput.t7 2.82907
R23654 CSoutput.n347 CSoutput.t98 2.82907
R23655 CSoutput.n345 CSoutput.t17 2.82907
R23656 CSoutput.n345 CSoutput.t108 2.82907
R23657 CSoutput.n344 CSoutput.t115 2.82907
R23658 CSoutput.n344 CSoutput.t5 2.82907
R23659 CSoutput.n342 CSoutput.t119 2.82907
R23660 CSoutput.n342 CSoutput.t63 2.82907
R23661 CSoutput.n340 CSoutput.t92 2.82907
R23662 CSoutput.n340 CSoutput.t103 2.82907
R23663 CSoutput.n338 CSoutput.t13 2.82907
R23664 CSoutput.n338 CSoutput.t39 2.82907
R23665 CSoutput.n336 CSoutput.t27 2.82907
R23666 CSoutput.n336 CSoutput.t59 2.82907
R23667 CSoutput.n334 CSoutput.t72 2.82907
R23668 CSoutput.n334 CSoutput.t86 2.82907
R23669 CSoutput.n332 CSoutput.t55 2.82907
R23670 CSoutput.n332 CSoutput.t110 2.82907
R23671 CSoutput.n330 CSoutput.t79 2.82907
R23672 CSoutput.n330 CSoutput.t45 2.82907
R23673 CSoutput.n328 CSoutput.t32 2.82907
R23674 CSoutput.n328 CSoutput.t58 2.82907
R23675 CSoutput.n326 CSoutput.t42 2.82907
R23676 CSoutput.n326 CSoutput.t51 2.82907
R23677 CSoutput.n325 CSoutput.t52 2.82907
R23678 CSoutput.n325 CSoutput.t120 2.82907
R23679 CSoutput.n424 CSoutput.t70 2.82907
R23680 CSoutput.n424 CSoutput.t102 2.82907
R23681 CSoutput.n425 CSoutput.t33 2.82907
R23682 CSoutput.n425 CSoutput.t50 2.82907
R23683 CSoutput.n427 CSoutput.t60 2.82907
R23684 CSoutput.n427 CSoutput.t81 2.82907
R23685 CSoutput.n429 CSoutput.t104 2.82907
R23686 CSoutput.n429 CSoutput.t66 2.82907
R23687 CSoutput.n431 CSoutput.t76 2.82907
R23688 CSoutput.n431 CSoutput.t116 2.82907
R23689 CSoutput.n433 CSoutput.t11 2.82907
R23690 CSoutput.n433 CSoutput.t36 2.82907
R23691 CSoutput.n435 CSoutput.t67 2.82907
R23692 CSoutput.n435 CSoutput.t96 2.82907
R23693 CSoutput.n437 CSoutput.t112 2.82907
R23694 CSoutput.n437 CSoutput.t22 2.82907
R23695 CSoutput.n439 CSoutput.t57 2.82907
R23696 CSoutput.n439 CSoutput.t77 2.82907
R23697 CSoutput.n441 CSoutput.t12 2.82907
R23698 CSoutput.n441 CSoutput.t47 2.82907
R23699 CSoutput.n404 CSoutput.t23 2.82907
R23700 CSoutput.n404 CSoutput.t14 2.82907
R23701 CSoutput.n405 CSoutput.t10 2.82907
R23702 CSoutput.n405 CSoutput.t121 2.82907
R23703 CSoutput.n407 CSoutput.t122 2.82907
R23704 CSoutput.n407 CSoutput.t24 2.82907
R23705 CSoutput.n409 CSoutput.t25 2.82907
R23706 CSoutput.n409 CSoutput.t82 2.82907
R23707 CSoutput.n411 CSoutput.t83 2.82907
R23708 CSoutput.n411 CSoutput.t114 2.82907
R23709 CSoutput.n413 CSoutput.t117 2.82907
R23710 CSoutput.n413 CSoutput.t106 2.82907
R23711 CSoutput.n415 CSoutput.t97 2.82907
R23712 CSoutput.n415 CSoutput.t84 2.82907
R23713 CSoutput.n417 CSoutput.t85 2.82907
R23714 CSoutput.n417 CSoutput.t118 2.82907
R23715 CSoutput.n419 CSoutput.t71 2.82907
R23716 CSoutput.n419 CSoutput.t99 2.82907
R23717 CSoutput.n421 CSoutput.t105 2.82907
R23718 CSoutput.n421 CSoutput.t80 2.82907
R23719 CSoutput.n385 CSoutput.t34 2.82907
R23720 CSoutput.n385 CSoutput.t91 2.82907
R23721 CSoutput.n386 CSoutput.t87 2.82907
R23722 CSoutput.n386 CSoutput.t61 2.82907
R23723 CSoutput.n388 CSoutput.t95 2.82907
R23724 CSoutput.n388 CSoutput.t49 2.82907
R23725 CSoutput.n390 CSoutput.t75 2.82907
R23726 CSoutput.n390 CSoutput.t113 2.82907
R23727 CSoutput.n392 CSoutput.t29 2.82907
R23728 CSoutput.n392 CSoutput.t94 2.82907
R23729 CSoutput.n394 CSoutput.t15 2.82907
R23730 CSoutput.n394 CSoutput.t101 2.82907
R23731 CSoutput.n396 CSoutput.t100 2.82907
R23732 CSoutput.n396 CSoutput.t41 2.82907
R23733 CSoutput.n398 CSoutput.t68 2.82907
R23734 CSoutput.n398 CSoutput.t37 2.82907
R23735 CSoutput.n400 CSoutput.t43 2.82907
R23736 CSoutput.n400 CSoutput.t18 2.82907
R23737 CSoutput.n402 CSoutput.t26 2.82907
R23738 CSoutput.n402 CSoutput.t44 2.82907
R23739 CSoutput.n75 CSoutput.n1 2.45513
R23740 CSoutput.n217 CSoutput.n215 2.251
R23741 CSoutput.n217 CSoutput.n214 2.251
R23742 CSoutput.n217 CSoutput.n213 2.251
R23743 CSoutput.n217 CSoutput.n212 2.251
R23744 CSoutput.n186 CSoutput.n185 2.251
R23745 CSoutput.n186 CSoutput.n184 2.251
R23746 CSoutput.n186 CSoutput.n183 2.251
R23747 CSoutput.n186 CSoutput.n182 2.251
R23748 CSoutput.n259 CSoutput.n258 2.251
R23749 CSoutput.n224 CSoutput.n222 2.251
R23750 CSoutput.n224 CSoutput.n221 2.251
R23751 CSoutput.n224 CSoutput.n220 2.251
R23752 CSoutput.n242 CSoutput.n224 2.251
R23753 CSoutput.n230 CSoutput.n229 2.251
R23754 CSoutput.n230 CSoutput.n228 2.251
R23755 CSoutput.n230 CSoutput.n227 2.251
R23756 CSoutput.n230 CSoutput.n226 2.251
R23757 CSoutput.n256 CSoutput.n196 2.251
R23758 CSoutput.n251 CSoutput.n249 2.251
R23759 CSoutput.n251 CSoutput.n248 2.251
R23760 CSoutput.n251 CSoutput.n247 2.251
R23761 CSoutput.n251 CSoutput.n246 2.251
R23762 CSoutput.n152 CSoutput.n151 2.251
R23763 CSoutput.n152 CSoutput.n150 2.251
R23764 CSoutput.n152 CSoutput.n149 2.251
R23765 CSoutput.n152 CSoutput.n148 2.251
R23766 CSoutput.n269 CSoutput.n268 2.251
R23767 CSoutput.n186 CSoutput.n166 2.2505
R23768 CSoutput.n181 CSoutput.n166 2.2505
R23769 CSoutput.n179 CSoutput.n166 2.2505
R23770 CSoutput.n178 CSoutput.n166 2.2505
R23771 CSoutput.n263 CSoutput.n166 2.2505
R23772 CSoutput.n261 CSoutput.n166 2.2505
R23773 CSoutput.n259 CSoutput.n166 2.2505
R23774 CSoutput.n189 CSoutput.n166 2.2505
R23775 CSoutput.n188 CSoutput.n166 2.2505
R23776 CSoutput.n192 CSoutput.n166 2.2505
R23777 CSoutput.n191 CSoutput.n166 2.2505
R23778 CSoutput.n174 CSoutput.n166 2.2505
R23779 CSoutput.n266 CSoutput.n166 2.2505
R23780 CSoutput.n266 CSoutput.n265 2.2505
R23781 CSoutput.n230 CSoutput.n201 2.2505
R23782 CSoutput.n211 CSoutput.n201 2.2505
R23783 CSoutput.n232 CSoutput.n201 2.2505
R23784 CSoutput.n210 CSoutput.n201 2.2505
R23785 CSoutput.n234 CSoutput.n201 2.2505
R23786 CSoutput.n201 CSoutput.n195 2.2505
R23787 CSoutput.n256 CSoutput.n201 2.2505
R23788 CSoutput.n254 CSoutput.n201 2.2505
R23789 CSoutput.n236 CSoutput.n201 2.2505
R23790 CSoutput.n208 CSoutput.n201 2.2505
R23791 CSoutput.n238 CSoutput.n201 2.2505
R23792 CSoutput.n207 CSoutput.n201 2.2505
R23793 CSoutput.n252 CSoutput.n201 2.2505
R23794 CSoutput.n252 CSoutput.n205 2.2505
R23795 CSoutput.n152 CSoutput.n132 2.2505
R23796 CSoutput.n147 CSoutput.n132 2.2505
R23797 CSoutput.n145 CSoutput.n132 2.2505
R23798 CSoutput.n144 CSoutput.n132 2.2505
R23799 CSoutput.n273 CSoutput.n132 2.2505
R23800 CSoutput.n271 CSoutput.n132 2.2505
R23801 CSoutput.n269 CSoutput.n132 2.2505
R23802 CSoutput.n155 CSoutput.n132 2.2505
R23803 CSoutput.n154 CSoutput.n132 2.2505
R23804 CSoutput.n158 CSoutput.n132 2.2505
R23805 CSoutput.n157 CSoutput.n132 2.2505
R23806 CSoutput.n140 CSoutput.n132 2.2505
R23807 CSoutput.n276 CSoutput.n132 2.2505
R23808 CSoutput.n276 CSoutput.n275 2.2505
R23809 CSoutput.n194 CSoutput.n187 2.25024
R23810 CSoutput.n194 CSoutput.n180 2.25024
R23811 CSoutput.n262 CSoutput.n194 2.25024
R23812 CSoutput.n194 CSoutput.n190 2.25024
R23813 CSoutput.n194 CSoutput.n193 2.25024
R23814 CSoutput.n194 CSoutput.n161 2.25024
R23815 CSoutput.n244 CSoutput.n241 2.25024
R23816 CSoutput.n244 CSoutput.n240 2.25024
R23817 CSoutput.n244 CSoutput.n239 2.25024
R23818 CSoutput.n244 CSoutput.n206 2.25024
R23819 CSoutput.n244 CSoutput.n243 2.25024
R23820 CSoutput.n245 CSoutput.n244 2.25024
R23821 CSoutput.n160 CSoutput.n153 2.25024
R23822 CSoutput.n160 CSoutput.n146 2.25024
R23823 CSoutput.n272 CSoutput.n160 2.25024
R23824 CSoutput.n160 CSoutput.n156 2.25024
R23825 CSoutput.n160 CSoutput.n159 2.25024
R23826 CSoutput.n160 CSoutput.n127 2.25024
R23827 CSoutput.n261 CSoutput.n171 1.50111
R23828 CSoutput.n209 CSoutput.n195 1.50111
R23829 CSoutput.n271 CSoutput.n137 1.50111
R23830 CSoutput.n217 CSoutput.n216 1.501
R23831 CSoutput.n224 CSoutput.n223 1.501
R23832 CSoutput.n251 CSoutput.n250 1.501
R23833 CSoutput.n265 CSoutput.n176 1.12536
R23834 CSoutput.n265 CSoutput.n177 1.12536
R23835 CSoutput.n265 CSoutput.n264 1.12536
R23836 CSoutput.n225 CSoutput.n205 1.12536
R23837 CSoutput.n231 CSoutput.n205 1.12536
R23838 CSoutput.n233 CSoutput.n205 1.12536
R23839 CSoutput.n275 CSoutput.n142 1.12536
R23840 CSoutput.n275 CSoutput.n143 1.12536
R23841 CSoutput.n275 CSoutput.n274 1.12536
R23842 CSoutput.n265 CSoutput.n172 1.12536
R23843 CSoutput.n265 CSoutput.n173 1.12536
R23844 CSoutput.n265 CSoutput.n175 1.12536
R23845 CSoutput.n255 CSoutput.n205 1.12536
R23846 CSoutput.n235 CSoutput.n205 1.12536
R23847 CSoutput.n237 CSoutput.n205 1.12536
R23848 CSoutput.n275 CSoutput.n138 1.12536
R23849 CSoutput.n275 CSoutput.n139 1.12536
R23850 CSoutput.n275 CSoutput.n141 1.12536
R23851 CSoutput.n31 CSoutput.n30 0.669944
R23852 CSoutput.n62 CSoutput.n61 0.669944
R23853 CSoutput.n368 CSoutput.n366 0.573776
R23854 CSoutput.n370 CSoutput.n368 0.573776
R23855 CSoutput.n372 CSoutput.n370 0.573776
R23856 CSoutput.n374 CSoutput.n372 0.573776
R23857 CSoutput.n376 CSoutput.n374 0.573776
R23858 CSoutput.n378 CSoutput.n376 0.573776
R23859 CSoutput.n380 CSoutput.n378 0.573776
R23860 CSoutput.n382 CSoutput.n380 0.573776
R23861 CSoutput.n348 CSoutput.n346 0.573776
R23862 CSoutput.n350 CSoutput.n348 0.573776
R23863 CSoutput.n352 CSoutput.n350 0.573776
R23864 CSoutput.n354 CSoutput.n352 0.573776
R23865 CSoutput.n356 CSoutput.n354 0.573776
R23866 CSoutput.n358 CSoutput.n356 0.573776
R23867 CSoutput.n360 CSoutput.n358 0.573776
R23868 CSoutput.n362 CSoutput.n360 0.573776
R23869 CSoutput.n329 CSoutput.n327 0.573776
R23870 CSoutput.n331 CSoutput.n329 0.573776
R23871 CSoutput.n333 CSoutput.n331 0.573776
R23872 CSoutput.n335 CSoutput.n333 0.573776
R23873 CSoutput.n337 CSoutput.n335 0.573776
R23874 CSoutput.n339 CSoutput.n337 0.573776
R23875 CSoutput.n341 CSoutput.n339 0.573776
R23876 CSoutput.n343 CSoutput.n341 0.573776
R23877 CSoutput.n442 CSoutput.n440 0.573776
R23878 CSoutput.n440 CSoutput.n438 0.573776
R23879 CSoutput.n438 CSoutput.n436 0.573776
R23880 CSoutput.n436 CSoutput.n434 0.573776
R23881 CSoutput.n434 CSoutput.n432 0.573776
R23882 CSoutput.n432 CSoutput.n430 0.573776
R23883 CSoutput.n430 CSoutput.n428 0.573776
R23884 CSoutput.n428 CSoutput.n426 0.573776
R23885 CSoutput.n422 CSoutput.n420 0.573776
R23886 CSoutput.n420 CSoutput.n418 0.573776
R23887 CSoutput.n418 CSoutput.n416 0.573776
R23888 CSoutput.n416 CSoutput.n414 0.573776
R23889 CSoutput.n414 CSoutput.n412 0.573776
R23890 CSoutput.n412 CSoutput.n410 0.573776
R23891 CSoutput.n410 CSoutput.n408 0.573776
R23892 CSoutput.n408 CSoutput.n406 0.573776
R23893 CSoutput.n403 CSoutput.n401 0.573776
R23894 CSoutput.n401 CSoutput.n399 0.573776
R23895 CSoutput.n399 CSoutput.n397 0.573776
R23896 CSoutput.n397 CSoutput.n395 0.573776
R23897 CSoutput.n395 CSoutput.n393 0.573776
R23898 CSoutput.n393 CSoutput.n391 0.573776
R23899 CSoutput.n391 CSoutput.n389 0.573776
R23900 CSoutput.n389 CSoutput.n387 0.573776
R23901 CSoutput.n445 CSoutput.n276 0.53442
R23902 CSoutput.n312 CSoutput.n310 0.358259
R23903 CSoutput.n314 CSoutput.n312 0.358259
R23904 CSoutput.n316 CSoutput.n314 0.358259
R23905 CSoutput.n318 CSoutput.n316 0.358259
R23906 CSoutput.n320 CSoutput.n318 0.358259
R23907 CSoutput.n322 CSoutput.n320 0.358259
R23908 CSoutput.n296 CSoutput.n294 0.358259
R23909 CSoutput.n298 CSoutput.n296 0.358259
R23910 CSoutput.n300 CSoutput.n298 0.358259
R23911 CSoutput.n302 CSoutput.n300 0.358259
R23912 CSoutput.n304 CSoutput.n302 0.358259
R23913 CSoutput.n306 CSoutput.n304 0.358259
R23914 CSoutput.n281 CSoutput.n279 0.358259
R23915 CSoutput.n283 CSoutput.n281 0.358259
R23916 CSoutput.n285 CSoutput.n283 0.358259
R23917 CSoutput.n287 CSoutput.n285 0.358259
R23918 CSoutput.n289 CSoutput.n287 0.358259
R23919 CSoutput.n291 CSoutput.n289 0.358259
R23920 CSoutput.n124 CSoutput.n122 0.358259
R23921 CSoutput.n122 CSoutput.n120 0.358259
R23922 CSoutput.n120 CSoutput.n118 0.358259
R23923 CSoutput.n118 CSoutput.n116 0.358259
R23924 CSoutput.n116 CSoutput.n114 0.358259
R23925 CSoutput.n114 CSoutput.n112 0.358259
R23926 CSoutput.n108 CSoutput.n106 0.358259
R23927 CSoutput.n106 CSoutput.n104 0.358259
R23928 CSoutput.n104 CSoutput.n102 0.358259
R23929 CSoutput.n102 CSoutput.n100 0.358259
R23930 CSoutput.n100 CSoutput.n98 0.358259
R23931 CSoutput.n98 CSoutput.n96 0.358259
R23932 CSoutput.n93 CSoutput.n91 0.358259
R23933 CSoutput.n91 CSoutput.n89 0.358259
R23934 CSoutput.n89 CSoutput.n87 0.358259
R23935 CSoutput.n87 CSoutput.n85 0.358259
R23936 CSoutput.n85 CSoutput.n83 0.358259
R23937 CSoutput.n83 CSoutput.n81 0.358259
R23938 CSoutput.n21 CSoutput.n20 0.169105
R23939 CSoutput.n21 CSoutput.n16 0.169105
R23940 CSoutput.n26 CSoutput.n16 0.169105
R23941 CSoutput.n27 CSoutput.n26 0.169105
R23942 CSoutput.n27 CSoutput.n14 0.169105
R23943 CSoutput.n32 CSoutput.n14 0.169105
R23944 CSoutput.n33 CSoutput.n32 0.169105
R23945 CSoutput.n34 CSoutput.n33 0.169105
R23946 CSoutput.n34 CSoutput.n12 0.169105
R23947 CSoutput.n39 CSoutput.n12 0.169105
R23948 CSoutput.n40 CSoutput.n39 0.169105
R23949 CSoutput.n40 CSoutput.n10 0.169105
R23950 CSoutput.n45 CSoutput.n10 0.169105
R23951 CSoutput.n46 CSoutput.n45 0.169105
R23952 CSoutput.n47 CSoutput.n46 0.169105
R23953 CSoutput.n47 CSoutput.n8 0.169105
R23954 CSoutput.n52 CSoutput.n8 0.169105
R23955 CSoutput.n53 CSoutput.n52 0.169105
R23956 CSoutput.n53 CSoutput.n6 0.169105
R23957 CSoutput.n58 CSoutput.n6 0.169105
R23958 CSoutput.n59 CSoutput.n58 0.169105
R23959 CSoutput.n60 CSoutput.n59 0.169105
R23960 CSoutput.n60 CSoutput.n4 0.169105
R23961 CSoutput.n66 CSoutput.n4 0.169105
R23962 CSoutput.n67 CSoutput.n66 0.169105
R23963 CSoutput.n68 CSoutput.n67 0.169105
R23964 CSoutput.n68 CSoutput.n2 0.169105
R23965 CSoutput.n73 CSoutput.n2 0.169105
R23966 CSoutput.n74 CSoutput.n73 0.169105
R23967 CSoutput.n74 CSoutput.n0 0.169105
R23968 CSoutput.n78 CSoutput.n0 0.169105
R23969 CSoutput.n219 CSoutput.n218 0.0910737
R23970 CSoutput.n270 CSoutput.n267 0.0723685
R23971 CSoutput.n224 CSoutput.n219 0.0522944
R23972 CSoutput.n267 CSoutput.n266 0.0499135
R23973 CSoutput.n218 CSoutput.n217 0.0499135
R23974 CSoutput.n252 CSoutput.n251 0.0464294
R23975 CSoutput.n260 CSoutput.n257 0.0391444
R23976 CSoutput.n219 CSoutput.t216 0.023435
R23977 CSoutput.n267 CSoutput.t219 0.02262
R23978 CSoutput.n218 CSoutput.t222 0.02262
R23979 CSoutput CSoutput.n445 0.0052
R23980 CSoutput.n189 CSoutput.n172 0.00365111
R23981 CSoutput.n192 CSoutput.n173 0.00365111
R23982 CSoutput.n175 CSoutput.n174 0.00365111
R23983 CSoutput.n217 CSoutput.n176 0.00365111
R23984 CSoutput.n181 CSoutput.n177 0.00365111
R23985 CSoutput.n264 CSoutput.n178 0.00365111
R23986 CSoutput.n255 CSoutput.n254 0.00365111
R23987 CSoutput.n235 CSoutput.n208 0.00365111
R23988 CSoutput.n237 CSoutput.n207 0.00365111
R23989 CSoutput.n225 CSoutput.n224 0.00365111
R23990 CSoutput.n231 CSoutput.n211 0.00365111
R23991 CSoutput.n233 CSoutput.n210 0.00365111
R23992 CSoutput.n155 CSoutput.n138 0.00365111
R23993 CSoutput.n158 CSoutput.n139 0.00365111
R23994 CSoutput.n141 CSoutput.n140 0.00365111
R23995 CSoutput.n251 CSoutput.n142 0.00365111
R23996 CSoutput.n147 CSoutput.n143 0.00365111
R23997 CSoutput.n274 CSoutput.n144 0.00365111
R23998 CSoutput.n186 CSoutput.n176 0.00340054
R23999 CSoutput.n179 CSoutput.n177 0.00340054
R24000 CSoutput.n264 CSoutput.n263 0.00340054
R24001 CSoutput.n259 CSoutput.n172 0.00340054
R24002 CSoutput.n188 CSoutput.n173 0.00340054
R24003 CSoutput.n191 CSoutput.n175 0.00340054
R24004 CSoutput.n230 CSoutput.n225 0.00340054
R24005 CSoutput.n232 CSoutput.n231 0.00340054
R24006 CSoutput.n234 CSoutput.n233 0.00340054
R24007 CSoutput.n256 CSoutput.n255 0.00340054
R24008 CSoutput.n236 CSoutput.n235 0.00340054
R24009 CSoutput.n238 CSoutput.n237 0.00340054
R24010 CSoutput.n152 CSoutput.n142 0.00340054
R24011 CSoutput.n145 CSoutput.n143 0.00340054
R24012 CSoutput.n274 CSoutput.n273 0.00340054
R24013 CSoutput.n269 CSoutput.n138 0.00340054
R24014 CSoutput.n154 CSoutput.n139 0.00340054
R24015 CSoutput.n157 CSoutput.n141 0.00340054
R24016 CSoutput.n187 CSoutput.n181 0.00252698
R24017 CSoutput.n180 CSoutput.n178 0.00252698
R24018 CSoutput.n262 CSoutput.n261 0.00252698
R24019 CSoutput.n190 CSoutput.n188 0.00252698
R24020 CSoutput.n193 CSoutput.n191 0.00252698
R24021 CSoutput.n266 CSoutput.n161 0.00252698
R24022 CSoutput.n187 CSoutput.n186 0.00252698
R24023 CSoutput.n180 CSoutput.n179 0.00252698
R24024 CSoutput.n263 CSoutput.n262 0.00252698
R24025 CSoutput.n190 CSoutput.n189 0.00252698
R24026 CSoutput.n193 CSoutput.n192 0.00252698
R24027 CSoutput.n174 CSoutput.n161 0.00252698
R24028 CSoutput.n241 CSoutput.n211 0.00252698
R24029 CSoutput.n240 CSoutput.n210 0.00252698
R24030 CSoutput.n239 CSoutput.n195 0.00252698
R24031 CSoutput.n236 CSoutput.n206 0.00252698
R24032 CSoutput.n243 CSoutput.n238 0.00252698
R24033 CSoutput.n252 CSoutput.n245 0.00252698
R24034 CSoutput.n241 CSoutput.n230 0.00252698
R24035 CSoutput.n240 CSoutput.n232 0.00252698
R24036 CSoutput.n239 CSoutput.n234 0.00252698
R24037 CSoutput.n254 CSoutput.n206 0.00252698
R24038 CSoutput.n243 CSoutput.n208 0.00252698
R24039 CSoutput.n245 CSoutput.n207 0.00252698
R24040 CSoutput.n153 CSoutput.n147 0.00252698
R24041 CSoutput.n146 CSoutput.n144 0.00252698
R24042 CSoutput.n272 CSoutput.n271 0.00252698
R24043 CSoutput.n156 CSoutput.n154 0.00252698
R24044 CSoutput.n159 CSoutput.n157 0.00252698
R24045 CSoutput.n276 CSoutput.n127 0.00252698
R24046 CSoutput.n153 CSoutput.n152 0.00252698
R24047 CSoutput.n146 CSoutput.n145 0.00252698
R24048 CSoutput.n273 CSoutput.n272 0.00252698
R24049 CSoutput.n156 CSoutput.n155 0.00252698
R24050 CSoutput.n159 CSoutput.n158 0.00252698
R24051 CSoutput.n140 CSoutput.n127 0.00252698
R24052 CSoutput.n261 CSoutput.n260 0.0020275
R24053 CSoutput.n260 CSoutput.n259 0.0020275
R24054 CSoutput.n257 CSoutput.n195 0.0020275
R24055 CSoutput.n257 CSoutput.n256 0.0020275
R24056 CSoutput.n271 CSoutput.n270 0.0020275
R24057 CSoutput.n270 CSoutput.n269 0.0020275
R24058 CSoutput.n171 CSoutput.n170 0.00166668
R24059 CSoutput.n253 CSoutput.n209 0.00166668
R24060 CSoutput.n137 CSoutput.n136 0.00166668
R24061 CSoutput.n275 CSoutput.n137 0.00133328
R24062 CSoutput.n209 CSoutput.n205 0.00133328
R24063 CSoutput.n265 CSoutput.n171 0.00133328
R24064 CSoutput.n268 CSoutput.n160 0.001
R24065 CSoutput.n246 CSoutput.n160 0.001
R24066 CSoutput.n148 CSoutput.n128 0.001
R24067 CSoutput.n247 CSoutput.n128 0.001
R24068 CSoutput.n149 CSoutput.n129 0.001
R24069 CSoutput.n248 CSoutput.n129 0.001
R24070 CSoutput.n150 CSoutput.n130 0.001
R24071 CSoutput.n249 CSoutput.n130 0.001
R24072 CSoutput.n151 CSoutput.n131 0.001
R24073 CSoutput.n250 CSoutput.n131 0.001
R24074 CSoutput.n244 CSoutput.n196 0.001
R24075 CSoutput.n244 CSoutput.n242 0.001
R24076 CSoutput.n226 CSoutput.n197 0.001
R24077 CSoutput.n220 CSoutput.n197 0.001
R24078 CSoutput.n227 CSoutput.n198 0.001
R24079 CSoutput.n221 CSoutput.n198 0.001
R24080 CSoutput.n228 CSoutput.n199 0.001
R24081 CSoutput.n222 CSoutput.n199 0.001
R24082 CSoutput.n229 CSoutput.n200 0.001
R24083 CSoutput.n223 CSoutput.n200 0.001
R24084 CSoutput.n258 CSoutput.n194 0.001
R24085 CSoutput.n212 CSoutput.n194 0.001
R24086 CSoutput.n182 CSoutput.n162 0.001
R24087 CSoutput.n213 CSoutput.n162 0.001
R24088 CSoutput.n183 CSoutput.n163 0.001
R24089 CSoutput.n214 CSoutput.n163 0.001
R24090 CSoutput.n184 CSoutput.n164 0.001
R24091 CSoutput.n215 CSoutput.n164 0.001
R24092 CSoutput.n185 CSoutput.n165 0.001
R24093 CSoutput.n216 CSoutput.n165 0.001
R24094 CSoutput.n216 CSoutput.n166 0.001
R24095 CSoutput.n215 CSoutput.n167 0.001
R24096 CSoutput.n214 CSoutput.n168 0.001
R24097 CSoutput.n213 CSoutput.t237 0.001
R24098 CSoutput.n212 CSoutput.n169 0.001
R24099 CSoutput.n185 CSoutput.n167 0.001
R24100 CSoutput.n184 CSoutput.n168 0.001
R24101 CSoutput.n183 CSoutput.t237 0.001
R24102 CSoutput.n182 CSoutput.n169 0.001
R24103 CSoutput.n258 CSoutput.n170 0.001
R24104 CSoutput.n223 CSoutput.n201 0.001
R24105 CSoutput.n222 CSoutput.n202 0.001
R24106 CSoutput.n221 CSoutput.n203 0.001
R24107 CSoutput.n220 CSoutput.t232 0.001
R24108 CSoutput.n242 CSoutput.n204 0.001
R24109 CSoutput.n229 CSoutput.n202 0.001
R24110 CSoutput.n228 CSoutput.n203 0.001
R24111 CSoutput.n227 CSoutput.t232 0.001
R24112 CSoutput.n226 CSoutput.n204 0.001
R24113 CSoutput.n253 CSoutput.n196 0.001
R24114 CSoutput.n250 CSoutput.n132 0.001
R24115 CSoutput.n249 CSoutput.n133 0.001
R24116 CSoutput.n248 CSoutput.n134 0.001
R24117 CSoutput.n247 CSoutput.t230 0.001
R24118 CSoutput.n246 CSoutput.n135 0.001
R24119 CSoutput.n151 CSoutput.n133 0.001
R24120 CSoutput.n150 CSoutput.n134 0.001
R24121 CSoutput.n149 CSoutput.t230 0.001
R24122 CSoutput.n148 CSoutput.n135 0.001
R24123 CSoutput.n268 CSoutput.n136 0.001
R24124 a_n8964_8799.n183 a_n8964_8799.t120 485.149
R24125 a_n8964_8799.n199 a_n8964_8799.t132 485.149
R24126 a_n8964_8799.n216 a_n8964_8799.t87 485.149
R24127 a_n8964_8799.n132 a_n8964_8799.t83 485.149
R24128 a_n8964_8799.n148 a_n8964_8799.t91 485.149
R24129 a_n8964_8799.n165 a_n8964_8799.t85 485.149
R24130 a_n8964_8799.n193 a_n8964_8799.t51 464.166
R24131 a_n8964_8799.n192 a_n8964_8799.t49 464.166
R24132 a_n8964_8799.n178 a_n8964_8799.t117 464.166
R24133 a_n8964_8799.n191 a_n8964_8799.t65 464.166
R24134 a_n8964_8799.n190 a_n8964_8799.t53 464.166
R24135 a_n8964_8799.n179 a_n8964_8799.t123 464.166
R24136 a_n8964_8799.n189 a_n8964_8799.t86 464.166
R24137 a_n8964_8799.n188 a_n8964_8799.t66 464.166
R24138 a_n8964_8799.n180 a_n8964_8799.t137 464.166
R24139 a_n8964_8799.n187 a_n8964_8799.t102 464.166
R24140 a_n8964_8799.n186 a_n8964_8799.t68 464.166
R24141 a_n8964_8799.n181 a_n8964_8799.t133 464.166
R24142 a_n8964_8799.n185 a_n8964_8799.t104 464.166
R24143 a_n8964_8799.n184 a_n8964_8799.t80 464.166
R24144 a_n8964_8799.n182 a_n8964_8799.t50 464.166
R24145 a_n8964_8799.n209 a_n8964_8799.t59 464.166
R24146 a_n8964_8799.n208 a_n8964_8799.t57 464.166
R24147 a_n8964_8799.n194 a_n8964_8799.t131 464.166
R24148 a_n8964_8799.n207 a_n8964_8799.t71 464.166
R24149 a_n8964_8799.n206 a_n8964_8799.t63 464.166
R24150 a_n8964_8799.n195 a_n8964_8799.t134 464.166
R24151 a_n8964_8799.n205 a_n8964_8799.t98 464.166
R24152 a_n8964_8799.n204 a_n8964_8799.t74 464.166
R24153 a_n8964_8799.n196 a_n8964_8799.t52 464.166
R24154 a_n8964_8799.n203 a_n8964_8799.t111 464.166
R24155 a_n8964_8799.n202 a_n8964_8799.t75 464.166
R24156 a_n8964_8799.n197 a_n8964_8799.t45 464.166
R24157 a_n8964_8799.n201 a_n8964_8799.t116 464.166
R24158 a_n8964_8799.n200 a_n8964_8799.t88 464.166
R24159 a_n8964_8799.n198 a_n8964_8799.t58 464.166
R24160 a_n8964_8799.n226 a_n8964_8799.t97 464.166
R24161 a_n8964_8799.n225 a_n8964_8799.t115 464.166
R24162 a_n8964_8799.n211 a_n8964_8799.t64 464.166
R24163 a_n8964_8799.n224 a_n8964_8799.t129 464.166
R24164 a_n8964_8799.n223 a_n8964_8799.t78 464.166
R24165 a_n8964_8799.n212 a_n8964_8799.t124 464.166
R24166 a_n8964_8799.n222 a_n8964_8799.t67 464.166
R24167 a_n8964_8799.n221 a_n8964_8799.t106 464.166
R24168 a_n8964_8799.n213 a_n8964_8799.t55 464.166
R24169 a_n8964_8799.n220 a_n8964_8799.t94 464.166
R24170 a_n8964_8799.n219 a_n8964_8799.t73 464.166
R24171 a_n8964_8799.n214 a_n8964_8799.t113 464.166
R24172 a_n8964_8799.n218 a_n8964_8799.t61 464.166
R24173 a_n8964_8799.n217 a_n8964_8799.t101 464.166
R24174 a_n8964_8799.n215 a_n8964_8799.t48 464.166
R24175 a_n8964_8799.n131 a_n8964_8799.t108 464.166
R24176 a_n8964_8799.n134 a_n8964_8799.t46 464.166
R24177 a_n8964_8799.n130 a_n8964_8799.t70 464.166
R24178 a_n8964_8799.n135 a_n8964_8799.t103 464.166
R24179 a_n8964_8799.n136 a_n8964_8799.t130 464.166
R24180 a_n8964_8799.n137 a_n8964_8799.t69 464.166
R24181 a_n8964_8799.n138 a_n8964_8799.t99 464.166
R24182 a_n8964_8799.n129 a_n8964_8799.t126 464.166
R24183 a_n8964_8799.n139 a_n8964_8799.t127 464.166
R24184 a_n8964_8799.n140 a_n8964_8799.t84 464.166
R24185 a_n8964_8799.n141 a_n8964_8799.t110 464.166
R24186 a_n8964_8799.n142 a_n8964_8799.t125 464.166
R24187 a_n8964_8799.n128 a_n8964_8799.t81 464.166
R24188 a_n8964_8799.n143 a_n8964_8799.t82 464.166
R24189 a_n8964_8799.n147 a_n8964_8799.t118 464.166
R24190 a_n8964_8799.n150 a_n8964_8799.t56 464.166
R24191 a_n8964_8799.n146 a_n8964_8799.t79 464.166
R24192 a_n8964_8799.n151 a_n8964_8799.t112 464.166
R24193 a_n8964_8799.n152 a_n8964_8799.t139 464.166
R24194 a_n8964_8799.n153 a_n8964_8799.t76 464.166
R24195 a_n8964_8799.n154 a_n8964_8799.t109 464.166
R24196 a_n8964_8799.n145 a_n8964_8799.t136 464.166
R24197 a_n8964_8799.n155 a_n8964_8799.t138 464.166
R24198 a_n8964_8799.n156 a_n8964_8799.t95 464.166
R24199 a_n8964_8799.n157 a_n8964_8799.t122 464.166
R24200 a_n8964_8799.n158 a_n8964_8799.t135 464.166
R24201 a_n8964_8799.n144 a_n8964_8799.t90 464.166
R24202 a_n8964_8799.n159 a_n8964_8799.t92 464.166
R24203 a_n8964_8799.n164 a_n8964_8799.t47 464.166
R24204 a_n8964_8799.n167 a_n8964_8799.t100 464.166
R24205 a_n8964_8799.n163 a_n8964_8799.t60 464.166
R24206 a_n8964_8799.n168 a_n8964_8799.t114 464.166
R24207 a_n8964_8799.n169 a_n8964_8799.t72 464.166
R24208 a_n8964_8799.n170 a_n8964_8799.t93 464.166
R24209 a_n8964_8799.n171 a_n8964_8799.t54 464.166
R24210 a_n8964_8799.n162 a_n8964_8799.t105 464.166
R24211 a_n8964_8799.n172 a_n8964_8799.t89 464.166
R24212 a_n8964_8799.n173 a_n8964_8799.t121 464.166
R24213 a_n8964_8799.n174 a_n8964_8799.t77 464.166
R24214 a_n8964_8799.n175 a_n8964_8799.t128 464.166
R24215 a_n8964_8799.n161 a_n8964_8799.t62 464.166
R24216 a_n8964_8799.n176 a_n8964_8799.t44 464.166
R24217 a_n8964_8799.n56 a_n8964_8799.n34 74.4178
R24218 a_n8964_8799.n184 a_n8964_8799.n56 12.4674
R24219 a_n8964_8799.n55 a_n8964_8799.n34 80.107
R24220 a_n8964_8799.n55 a_n8964_8799.n185 1.08907
R24221 a_n8964_8799.n35 a_n8964_8799.n54 75.3623
R24222 a_n8964_8799.n53 a_n8964_8799.n35 70.3058
R24223 a_n8964_8799.n37 a_n8964_8799.n52 70.1674
R24224 a_n8964_8799.n52 a_n8964_8799.n180 20.9683
R24225 a_n8964_8799.n51 a_n8964_8799.n37 75.0448
R24226 a_n8964_8799.n188 a_n8964_8799.n51 11.2134
R24227 a_n8964_8799.n50 a_n8964_8799.n36 80.4688
R24228 a_n8964_8799.n36 a_n8964_8799.n49 74.73
R24229 a_n8964_8799.n48 a_n8964_8799.n38 70.1674
R24230 a_n8964_8799.n191 a_n8964_8799.n48 20.9683
R24231 a_n8964_8799.n38 a_n8964_8799.n47 70.5844
R24232 a_n8964_8799.n47 a_n8964_8799.n178 20.1342
R24233 a_n8964_8799.n46 a_n8964_8799.n39 75.6825
R24234 a_n8964_8799.n192 a_n8964_8799.n46 9.93802
R24235 a_n8964_8799.n39 a_n8964_8799.n193 161.3
R24236 a_n8964_8799.n67 a_n8964_8799.n28 74.4178
R24237 a_n8964_8799.n200 a_n8964_8799.n67 12.4674
R24238 a_n8964_8799.n66 a_n8964_8799.n28 80.107
R24239 a_n8964_8799.n66 a_n8964_8799.n201 1.08907
R24240 a_n8964_8799.n29 a_n8964_8799.n65 75.3623
R24241 a_n8964_8799.n64 a_n8964_8799.n29 70.3058
R24242 a_n8964_8799.n31 a_n8964_8799.n63 70.1674
R24243 a_n8964_8799.n63 a_n8964_8799.n196 20.9683
R24244 a_n8964_8799.n62 a_n8964_8799.n31 75.0448
R24245 a_n8964_8799.n204 a_n8964_8799.n62 11.2134
R24246 a_n8964_8799.n61 a_n8964_8799.n30 80.4688
R24247 a_n8964_8799.n30 a_n8964_8799.n60 74.73
R24248 a_n8964_8799.n59 a_n8964_8799.n32 70.1674
R24249 a_n8964_8799.n207 a_n8964_8799.n59 20.9683
R24250 a_n8964_8799.n32 a_n8964_8799.n58 70.5844
R24251 a_n8964_8799.n58 a_n8964_8799.n194 20.1342
R24252 a_n8964_8799.n57 a_n8964_8799.n33 75.6825
R24253 a_n8964_8799.n208 a_n8964_8799.n57 9.93802
R24254 a_n8964_8799.n33 a_n8964_8799.n209 161.3
R24255 a_n8964_8799.n78 a_n8964_8799.n22 74.4178
R24256 a_n8964_8799.n217 a_n8964_8799.n78 12.4674
R24257 a_n8964_8799.n77 a_n8964_8799.n22 80.107
R24258 a_n8964_8799.n77 a_n8964_8799.n218 1.08907
R24259 a_n8964_8799.n23 a_n8964_8799.n76 75.3623
R24260 a_n8964_8799.n75 a_n8964_8799.n23 70.3058
R24261 a_n8964_8799.n25 a_n8964_8799.n74 70.1674
R24262 a_n8964_8799.n74 a_n8964_8799.n213 20.9683
R24263 a_n8964_8799.n73 a_n8964_8799.n25 75.0448
R24264 a_n8964_8799.n221 a_n8964_8799.n73 11.2134
R24265 a_n8964_8799.n72 a_n8964_8799.n24 80.4688
R24266 a_n8964_8799.n24 a_n8964_8799.n71 74.73
R24267 a_n8964_8799.n70 a_n8964_8799.n26 70.1674
R24268 a_n8964_8799.n224 a_n8964_8799.n70 20.9683
R24269 a_n8964_8799.n26 a_n8964_8799.n69 70.5844
R24270 a_n8964_8799.n69 a_n8964_8799.n211 20.1342
R24271 a_n8964_8799.n68 a_n8964_8799.n27 75.6825
R24272 a_n8964_8799.n225 a_n8964_8799.n68 9.93802
R24273 a_n8964_8799.n27 a_n8964_8799.n226 161.3
R24274 a_n8964_8799.n17 a_n8964_8799.n89 70.1674
R24275 a_n8964_8799.n143 a_n8964_8799.n89 20.9683
R24276 a_n8964_8799.n88 a_n8964_8799.n17 74.4178
R24277 a_n8964_8799.n88 a_n8964_8799.n128 12.4674
R24278 a_n8964_8799.n16 a_n8964_8799.n87 80.107
R24279 a_n8964_8799.n142 a_n8964_8799.n87 1.08907
R24280 a_n8964_8799.n86 a_n8964_8799.n16 75.3623
R24281 a_n8964_8799.n18 a_n8964_8799.n85 70.3058
R24282 a_n8964_8799.n84 a_n8964_8799.n18 70.1674
R24283 a_n8964_8799.n84 a_n8964_8799.n129 20.9683
R24284 a_n8964_8799.n19 a_n8964_8799.n83 75.0448
R24285 a_n8964_8799.n138 a_n8964_8799.n83 11.2134
R24286 a_n8964_8799.n82 a_n8964_8799.n19 80.4688
R24287 a_n8964_8799.n20 a_n8964_8799.n81 74.73
R24288 a_n8964_8799.n80 a_n8964_8799.n20 70.1674
R24289 a_n8964_8799.n80 a_n8964_8799.n130 20.9683
R24290 a_n8964_8799.n21 a_n8964_8799.n79 70.5844
R24291 a_n8964_8799.n134 a_n8964_8799.n79 20.1342
R24292 a_n8964_8799.n133 a_n8964_8799.n21 161.3
R24293 a_n8964_8799.n11 a_n8964_8799.n100 70.1674
R24294 a_n8964_8799.n159 a_n8964_8799.n100 20.9683
R24295 a_n8964_8799.n99 a_n8964_8799.n11 74.4178
R24296 a_n8964_8799.n99 a_n8964_8799.n144 12.4674
R24297 a_n8964_8799.n10 a_n8964_8799.n98 80.107
R24298 a_n8964_8799.n158 a_n8964_8799.n98 1.08907
R24299 a_n8964_8799.n97 a_n8964_8799.n10 75.3623
R24300 a_n8964_8799.n12 a_n8964_8799.n96 70.3058
R24301 a_n8964_8799.n95 a_n8964_8799.n12 70.1674
R24302 a_n8964_8799.n95 a_n8964_8799.n145 20.9683
R24303 a_n8964_8799.n13 a_n8964_8799.n94 75.0448
R24304 a_n8964_8799.n154 a_n8964_8799.n94 11.2134
R24305 a_n8964_8799.n93 a_n8964_8799.n13 80.4688
R24306 a_n8964_8799.n14 a_n8964_8799.n92 74.73
R24307 a_n8964_8799.n91 a_n8964_8799.n14 70.1674
R24308 a_n8964_8799.n91 a_n8964_8799.n146 20.9683
R24309 a_n8964_8799.n15 a_n8964_8799.n90 70.5844
R24310 a_n8964_8799.n150 a_n8964_8799.n90 20.1342
R24311 a_n8964_8799.n149 a_n8964_8799.n15 161.3
R24312 a_n8964_8799.n5 a_n8964_8799.n111 70.1674
R24313 a_n8964_8799.n176 a_n8964_8799.n111 20.9683
R24314 a_n8964_8799.n110 a_n8964_8799.n5 74.4178
R24315 a_n8964_8799.n110 a_n8964_8799.n161 12.4674
R24316 a_n8964_8799.n4 a_n8964_8799.n109 80.107
R24317 a_n8964_8799.n175 a_n8964_8799.n109 1.08907
R24318 a_n8964_8799.n108 a_n8964_8799.n4 75.3623
R24319 a_n8964_8799.n6 a_n8964_8799.n107 70.3058
R24320 a_n8964_8799.n106 a_n8964_8799.n6 70.1674
R24321 a_n8964_8799.n106 a_n8964_8799.n162 20.9683
R24322 a_n8964_8799.n7 a_n8964_8799.n105 75.0448
R24323 a_n8964_8799.n171 a_n8964_8799.n105 11.2134
R24324 a_n8964_8799.n104 a_n8964_8799.n7 80.4688
R24325 a_n8964_8799.n8 a_n8964_8799.n103 74.73
R24326 a_n8964_8799.n102 a_n8964_8799.n8 70.1674
R24327 a_n8964_8799.n102 a_n8964_8799.n163 20.9683
R24328 a_n8964_8799.n9 a_n8964_8799.n101 70.5844
R24329 a_n8964_8799.n167 a_n8964_8799.n101 20.1342
R24330 a_n8964_8799.n166 a_n8964_8799.n9 161.3
R24331 a_n8964_8799.n40 a_n8964_8799.n112 98.9633
R24332 a_n8964_8799.n43 a_n8964_8799.n233 98.9631
R24333 a_n8964_8799.n43 a_n8964_8799.n234 98.6055
R24334 a_n8964_8799.n43 a_n8964_8799.n235 98.6055
R24335 a_n8964_8799.n45 a_n8964_8799.n232 98.6055
R24336 a_n8964_8799.n44 a_n8964_8799.n231 98.6055
R24337 a_n8964_8799.n42 a_n8964_8799.n117 98.6055
R24338 a_n8964_8799.n42 a_n8964_8799.n116 98.6055
R24339 a_n8964_8799.n41 a_n8964_8799.n115 98.6055
R24340 a_n8964_8799.n41 a_n8964_8799.n114 98.6055
R24341 a_n8964_8799.n40 a_n8964_8799.n113 98.6055
R24342 a_n8964_8799.n236 a_n8964_8799.n45 98.6054
R24343 a_n8964_8799.n3 a_n8964_8799.n118 81.4626
R24344 a_n8964_8799.n1 a_n8964_8799.n124 81.4626
R24345 a_n8964_8799.n0 a_n8964_8799.n121 81.4626
R24346 a_n8964_8799.n2 a_n8964_8799.n126 80.9324
R24347 a_n8964_8799.n2 a_n8964_8799.n127 80.9324
R24348 a_n8964_8799.n3 a_n8964_8799.n120 80.9324
R24349 a_n8964_8799.n3 a_n8964_8799.n119 80.9324
R24350 a_n8964_8799.n1 a_n8964_8799.n125 80.9324
R24351 a_n8964_8799.n1 a_n8964_8799.n123 80.9324
R24352 a_n8964_8799.n0 a_n8964_8799.n122 80.9324
R24353 a_n8964_8799.n34 a_n8964_8799.n183 70.4033
R24354 a_n8964_8799.n28 a_n8964_8799.n199 70.4033
R24355 a_n8964_8799.n22 a_n8964_8799.n216 70.4033
R24356 a_n8964_8799.n21 a_n8964_8799.n132 70.4033
R24357 a_n8964_8799.n15 a_n8964_8799.n148 70.4033
R24358 a_n8964_8799.n9 a_n8964_8799.n165 70.4033
R24359 a_n8964_8799.n193 a_n8964_8799.n192 48.2005
R24360 a_n8964_8799.n48 a_n8964_8799.n190 20.9683
R24361 a_n8964_8799.n189 a_n8964_8799.n188 48.2005
R24362 a_n8964_8799.n187 a_n8964_8799.n52 20.9683
R24363 a_n8964_8799.n185 a_n8964_8799.n181 48.2005
R24364 a_n8964_8799.n209 a_n8964_8799.n208 48.2005
R24365 a_n8964_8799.n59 a_n8964_8799.n206 20.9683
R24366 a_n8964_8799.n205 a_n8964_8799.n204 48.2005
R24367 a_n8964_8799.n203 a_n8964_8799.n63 20.9683
R24368 a_n8964_8799.n201 a_n8964_8799.n197 48.2005
R24369 a_n8964_8799.n226 a_n8964_8799.n225 48.2005
R24370 a_n8964_8799.n70 a_n8964_8799.n223 20.9683
R24371 a_n8964_8799.n222 a_n8964_8799.n221 48.2005
R24372 a_n8964_8799.n220 a_n8964_8799.n74 20.9683
R24373 a_n8964_8799.n218 a_n8964_8799.n214 48.2005
R24374 a_n8964_8799.n135 a_n8964_8799.n80 20.9683
R24375 a_n8964_8799.n138 a_n8964_8799.n137 48.2005
R24376 a_n8964_8799.n139 a_n8964_8799.n84 20.9683
R24377 a_n8964_8799.n142 a_n8964_8799.n141 48.2005
R24378 a_n8964_8799.t107 a_n8964_8799.n89 485.135
R24379 a_n8964_8799.n151 a_n8964_8799.n91 20.9683
R24380 a_n8964_8799.n154 a_n8964_8799.n153 48.2005
R24381 a_n8964_8799.n155 a_n8964_8799.n95 20.9683
R24382 a_n8964_8799.n158 a_n8964_8799.n157 48.2005
R24383 a_n8964_8799.t119 a_n8964_8799.n100 485.135
R24384 a_n8964_8799.n168 a_n8964_8799.n102 20.9683
R24385 a_n8964_8799.n171 a_n8964_8799.n170 48.2005
R24386 a_n8964_8799.n172 a_n8964_8799.n106 20.9683
R24387 a_n8964_8799.n175 a_n8964_8799.n174 48.2005
R24388 a_n8964_8799.t96 a_n8964_8799.n111 485.135
R24389 a_n8964_8799.n50 a_n8964_8799.n179 47.835
R24390 a_n8964_8799.n53 a_n8964_8799.n186 20.6913
R24391 a_n8964_8799.n61 a_n8964_8799.n195 47.835
R24392 a_n8964_8799.n64 a_n8964_8799.n202 20.6913
R24393 a_n8964_8799.n72 a_n8964_8799.n212 47.835
R24394 a_n8964_8799.n75 a_n8964_8799.n219 20.6913
R24395 a_n8964_8799.n136 a_n8964_8799.n82 47.835
R24396 a_n8964_8799.n140 a_n8964_8799.n85 20.6913
R24397 a_n8964_8799.n152 a_n8964_8799.n93 47.835
R24398 a_n8964_8799.n156 a_n8964_8799.n96 20.6913
R24399 a_n8964_8799.n169 a_n8964_8799.n104 47.835
R24400 a_n8964_8799.n173 a_n8964_8799.n107 20.6913
R24401 a_n8964_8799.n191 a_n8964_8799.n47 22.3251
R24402 a_n8964_8799.n207 a_n8964_8799.n58 22.3251
R24403 a_n8964_8799.n224 a_n8964_8799.n69 22.3251
R24404 a_n8964_8799.n130 a_n8964_8799.n79 22.3251
R24405 a_n8964_8799.n146 a_n8964_8799.n90 22.3251
R24406 a_n8964_8799.n163 a_n8964_8799.n101 22.3251
R24407 a_n8964_8799.n44 a_n8964_8799.n230 34.1489
R24408 a_n8964_8799.n2 a_n8964_8799.n1 33.5285
R24409 a_n8964_8799.n56 a_n8964_8799.n182 33.6462
R24410 a_n8964_8799.n67 a_n8964_8799.n198 33.6462
R24411 a_n8964_8799.n78 a_n8964_8799.n215 33.6462
R24412 a_n8964_8799.n134 a_n8964_8799.n133 27.0217
R24413 a_n8964_8799.n143 a_n8964_8799.n88 33.6462
R24414 a_n8964_8799.n150 a_n8964_8799.n149 27.0217
R24415 a_n8964_8799.n159 a_n8964_8799.n99 33.6462
R24416 a_n8964_8799.n167 a_n8964_8799.n166 27.0217
R24417 a_n8964_8799.n176 a_n8964_8799.n110 33.6462
R24418 a_n8964_8799.n49 a_n8964_8799.n179 11.843
R24419 a_n8964_8799.n186 a_n8964_8799.n54 36.139
R24420 a_n8964_8799.n60 a_n8964_8799.n195 11.843
R24421 a_n8964_8799.n202 a_n8964_8799.n65 36.139
R24422 a_n8964_8799.n71 a_n8964_8799.n212 11.843
R24423 a_n8964_8799.n219 a_n8964_8799.n76 36.139
R24424 a_n8964_8799.n136 a_n8964_8799.n81 11.843
R24425 a_n8964_8799.n140 a_n8964_8799.n86 36.139
R24426 a_n8964_8799.n152 a_n8964_8799.n92 11.843
R24427 a_n8964_8799.n156 a_n8964_8799.n97 36.139
R24428 a_n8964_8799.n169 a_n8964_8799.n103 11.843
R24429 a_n8964_8799.n173 a_n8964_8799.n108 36.139
R24430 a_n8964_8799.n51 a_n8964_8799.n180 35.3134
R24431 a_n8964_8799.n62 a_n8964_8799.n196 35.3134
R24432 a_n8964_8799.n73 a_n8964_8799.n213 35.3134
R24433 a_n8964_8799.n129 a_n8964_8799.n83 35.3134
R24434 a_n8964_8799.n145 a_n8964_8799.n94 35.3134
R24435 a_n8964_8799.n162 a_n8964_8799.n105 35.3134
R24436 a_n8964_8799.n190 a_n8964_8799.n49 34.4824
R24437 a_n8964_8799.n54 a_n8964_8799.n181 10.5784
R24438 a_n8964_8799.n206 a_n8964_8799.n60 34.4824
R24439 a_n8964_8799.n65 a_n8964_8799.n197 10.5784
R24440 a_n8964_8799.n223 a_n8964_8799.n71 34.4824
R24441 a_n8964_8799.n76 a_n8964_8799.n214 10.5784
R24442 a_n8964_8799.n81 a_n8964_8799.n135 34.4824
R24443 a_n8964_8799.n141 a_n8964_8799.n86 10.5784
R24444 a_n8964_8799.n92 a_n8964_8799.n151 34.4824
R24445 a_n8964_8799.n157 a_n8964_8799.n97 10.5784
R24446 a_n8964_8799.n103 a_n8964_8799.n168 34.4824
R24447 a_n8964_8799.n174 a_n8964_8799.n108 10.5784
R24448 a_n8964_8799.n46 a_n8964_8799.n178 36.9592
R24449 a_n8964_8799.n57 a_n8964_8799.n194 36.9592
R24450 a_n8964_8799.n68 a_n8964_8799.n211 36.9592
R24451 a_n8964_8799.n133 a_n8964_8799.n131 21.1793
R24452 a_n8964_8799.n149 a_n8964_8799.n147 21.1793
R24453 a_n8964_8799.n166 a_n8964_8799.n164 21.1793
R24454 a_n8964_8799.n183 a_n8964_8799.n182 20.9576
R24455 a_n8964_8799.n199 a_n8964_8799.n198 20.9576
R24456 a_n8964_8799.n216 a_n8964_8799.n215 20.9576
R24457 a_n8964_8799.n132 a_n8964_8799.n131 20.9576
R24458 a_n8964_8799.n148 a_n8964_8799.n147 20.9576
R24459 a_n8964_8799.n165 a_n8964_8799.n164 20.9576
R24460 a_n8964_8799.n230 a_n8964_8799.n42 20.7404
R24461 a_n8964_8799.n229 a_n8964_8799.n3 12.3339
R24462 a_n8964_8799.n230 a_n8964_8799.n229 11.4887
R24463 a_n8964_8799.n210 a_n8964_8799.n39 9.07815
R24464 a_n8964_8799.n160 a_n8964_8799.n17 9.07815
R24465 a_n8964_8799.n228 a_n8964_8799.n177 7.21326
R24466 a_n8964_8799.n228 a_n8964_8799.n227 6.79371
R24467 a_n8964_8799.n210 a_n8964_8799.n33 4.9702
R24468 a_n8964_8799.n227 a_n8964_8799.n27 4.9702
R24469 a_n8964_8799.n160 a_n8964_8799.n11 4.9702
R24470 a_n8964_8799.n177 a_n8964_8799.n5 4.9702
R24471 a_n8964_8799.n227 a_n8964_8799.n210 4.10845
R24472 a_n8964_8799.n177 a_n8964_8799.n160 4.10845
R24473 a_n8964_8799.n233 a_n8964_8799.t17 3.61217
R24474 a_n8964_8799.n233 a_n8964_8799.t34 3.61217
R24475 a_n8964_8799.n234 a_n8964_8799.t36 3.61217
R24476 a_n8964_8799.n234 a_n8964_8799.t31 3.61217
R24477 a_n8964_8799.n235 a_n8964_8799.t19 3.61217
R24478 a_n8964_8799.n235 a_n8964_8799.t26 3.61217
R24479 a_n8964_8799.n232 a_n8964_8799.t30 3.61217
R24480 a_n8964_8799.n232 a_n8964_8799.t14 3.61217
R24481 a_n8964_8799.n231 a_n8964_8799.t22 3.61217
R24482 a_n8964_8799.n231 a_n8964_8799.t27 3.61217
R24483 a_n8964_8799.n117 a_n8964_8799.t32 3.61217
R24484 a_n8964_8799.n117 a_n8964_8799.t25 3.61217
R24485 a_n8964_8799.n116 a_n8964_8799.t15 3.61217
R24486 a_n8964_8799.n116 a_n8964_8799.t28 3.61217
R24487 a_n8964_8799.n115 a_n8964_8799.t23 3.61217
R24488 a_n8964_8799.n115 a_n8964_8799.t35 3.61217
R24489 a_n8964_8799.n114 a_n8964_8799.t20 3.61217
R24490 a_n8964_8799.n114 a_n8964_8799.t24 3.61217
R24491 a_n8964_8799.n113 a_n8964_8799.t18 3.61217
R24492 a_n8964_8799.n113 a_n8964_8799.t29 3.61217
R24493 a_n8964_8799.n112 a_n8964_8799.t21 3.61217
R24494 a_n8964_8799.n112 a_n8964_8799.t16 3.61217
R24495 a_n8964_8799.t13 a_n8964_8799.n236 3.61217
R24496 a_n8964_8799.n236 a_n8964_8799.t33 3.61217
R24497 a_n8964_8799.n229 a_n8964_8799.n228 3.4105
R24498 a_n8964_8799.n126 a_n8964_8799.t43 2.82907
R24499 a_n8964_8799.n126 a_n8964_8799.t12 2.82907
R24500 a_n8964_8799.n127 a_n8964_8799.t2 2.82907
R24501 a_n8964_8799.n127 a_n8964_8799.t5 2.82907
R24502 a_n8964_8799.n120 a_n8964_8799.t40 2.82907
R24503 a_n8964_8799.n120 a_n8964_8799.t37 2.82907
R24504 a_n8964_8799.n119 a_n8964_8799.t8 2.82907
R24505 a_n8964_8799.n119 a_n8964_8799.t10 2.82907
R24506 a_n8964_8799.n118 a_n8964_8799.t6 2.82907
R24507 a_n8964_8799.n118 a_n8964_8799.t11 2.82907
R24508 a_n8964_8799.n124 a_n8964_8799.t4 2.82907
R24509 a_n8964_8799.n124 a_n8964_8799.t9 2.82907
R24510 a_n8964_8799.n125 a_n8964_8799.t7 2.82907
R24511 a_n8964_8799.n125 a_n8964_8799.t1 2.82907
R24512 a_n8964_8799.n123 a_n8964_8799.t38 2.82907
R24513 a_n8964_8799.n123 a_n8964_8799.t41 2.82907
R24514 a_n8964_8799.n122 a_n8964_8799.t39 2.82907
R24515 a_n8964_8799.n122 a_n8964_8799.t42 2.82907
R24516 a_n8964_8799.n121 a_n8964_8799.t0 2.82907
R24517 a_n8964_8799.n121 a_n8964_8799.t3 2.82907
R24518 a_n8964_8799.n55 a_n8964_8799.n184 47.0982
R24519 a_n8964_8799.n66 a_n8964_8799.n200 47.0982
R24520 a_n8964_8799.n77 a_n8964_8799.n217 47.0982
R24521 a_n8964_8799.n128 a_n8964_8799.n87 47.0982
R24522 a_n8964_8799.n144 a_n8964_8799.n98 47.0982
R24523 a_n8964_8799.n161 a_n8964_8799.n109 47.0982
R24524 a_n8964_8799.n50 a_n8964_8799.n189 0.365327
R24525 a_n8964_8799.n187 a_n8964_8799.n53 21.4216
R24526 a_n8964_8799.n61 a_n8964_8799.n205 0.365327
R24527 a_n8964_8799.n203 a_n8964_8799.n64 21.4216
R24528 a_n8964_8799.n72 a_n8964_8799.n222 0.365327
R24529 a_n8964_8799.n220 a_n8964_8799.n75 21.4216
R24530 a_n8964_8799.n137 a_n8964_8799.n82 0.365327
R24531 a_n8964_8799.n85 a_n8964_8799.n139 21.4216
R24532 a_n8964_8799.n153 a_n8964_8799.n93 0.365327
R24533 a_n8964_8799.n96 a_n8964_8799.n155 21.4216
R24534 a_n8964_8799.n170 a_n8964_8799.n104 0.365327
R24535 a_n8964_8799.n107 a_n8964_8799.n172 21.4216
R24536 a_n8964_8799.n3 a_n8964_8799.n2 1.59102
R24537 a_n8964_8799.n35 a_n8964_8799.n34 1.13686
R24538 a_n8964_8799.n29 a_n8964_8799.n28 1.13686
R24539 a_n8964_8799.n23 a_n8964_8799.n22 1.13686
R24540 a_n8964_8799.n17 a_n8964_8799.n16 1.13686
R24541 a_n8964_8799.n11 a_n8964_8799.n10 1.13686
R24542 a_n8964_8799.n5 a_n8964_8799.n4 1.13686
R24543 a_n8964_8799.n1 a_n8964_8799.n0 1.06084
R24544 a_n8964_8799.n39 a_n8964_8799.n38 0.758076
R24545 a_n8964_8799.n36 a_n8964_8799.n38 0.758076
R24546 a_n8964_8799.n37 a_n8964_8799.n36 0.758076
R24547 a_n8964_8799.n37 a_n8964_8799.n35 0.758076
R24548 a_n8964_8799.n33 a_n8964_8799.n32 0.758076
R24549 a_n8964_8799.n30 a_n8964_8799.n32 0.758076
R24550 a_n8964_8799.n31 a_n8964_8799.n30 0.758076
R24551 a_n8964_8799.n31 a_n8964_8799.n29 0.758076
R24552 a_n8964_8799.n27 a_n8964_8799.n26 0.758076
R24553 a_n8964_8799.n24 a_n8964_8799.n26 0.758076
R24554 a_n8964_8799.n25 a_n8964_8799.n24 0.758076
R24555 a_n8964_8799.n25 a_n8964_8799.n23 0.758076
R24556 a_n8964_8799.n20 a_n8964_8799.n21 0.758076
R24557 a_n8964_8799.n19 a_n8964_8799.n20 0.758076
R24558 a_n8964_8799.n18 a_n8964_8799.n19 0.758076
R24559 a_n8964_8799.n16 a_n8964_8799.n18 0.758076
R24560 a_n8964_8799.n14 a_n8964_8799.n15 0.758076
R24561 a_n8964_8799.n13 a_n8964_8799.n14 0.758076
R24562 a_n8964_8799.n12 a_n8964_8799.n13 0.758076
R24563 a_n8964_8799.n10 a_n8964_8799.n12 0.758076
R24564 a_n8964_8799.n8 a_n8964_8799.n9 0.758076
R24565 a_n8964_8799.n7 a_n8964_8799.n8 0.758076
R24566 a_n8964_8799.n6 a_n8964_8799.n7 0.758076
R24567 a_n8964_8799.n4 a_n8964_8799.n6 0.758076
R24568 a_n8964_8799.n45 a_n8964_8799.n43 0.716017
R24569 a_n8964_8799.n45 a_n8964_8799.n44 0.716017
R24570 a_n8964_8799.n42 a_n8964_8799.n41 0.716017
R24571 a_n8964_8799.n41 a_n8964_8799.n40 0.716017
R24572 plus.n61 plus.t11 251.488
R24573 plus.n12 plus.t14 251.488
R24574 plus.n100 plus.t1 243.97
R24575 plus.n96 plus.t23 231.093
R24576 plus.n47 plus.t6 231.093
R24577 plus.n100 plus.n99 223.454
R24578 plus.n102 plus.n101 223.454
R24579 plus.n60 plus.t5 187.445
R24580 plus.n65 plus.t21 187.445
R24581 plus.n71 plus.t20 187.445
R24582 plus.n56 plus.t16 187.445
R24583 plus.n54 plus.t17 187.445
R24584 plus.n83 plus.t13 187.445
R24585 plus.n89 plus.t15 187.445
R24586 plus.n50 plus.t10 187.445
R24587 plus.n1 plus.t12 187.445
R24588 plus.n40 plus.t8 187.445
R24589 plus.n34 plus.t7 187.445
R24590 plus.n5 plus.t19 187.445
R24591 plus.n7 plus.t18 187.445
R24592 plus.n22 plus.t24 187.445
R24593 plus.n16 plus.t22 187.445
R24594 plus.n11 plus.t9 187.445
R24595 plus.n97 plus.n96 161.3
R24596 plus.n95 plus.n49 161.3
R24597 plus.n94 plus.n93 161.3
R24598 plus.n92 plus.n91 161.3
R24599 plus.n90 plus.n51 161.3
R24600 plus.n88 plus.n87 161.3
R24601 plus.n86 plus.n52 161.3
R24602 plus.n85 plus.n84 161.3
R24603 plus.n82 plus.n53 161.3
R24604 plus.n81 plus.n80 161.3
R24605 plus.n79 plus.n78 161.3
R24606 plus.n77 plus.n55 161.3
R24607 plus.n76 plus.n75 161.3
R24608 plus.n74 plus.n73 161.3
R24609 plus.n72 plus.n57 161.3
R24610 plus.n70 plus.n69 161.3
R24611 plus.n68 plus.n58 161.3
R24612 plus.n67 plus.n66 161.3
R24613 plus.n64 plus.n59 161.3
R24614 plus.n63 plus.n62 161.3
R24615 plus.n14 plus.n13 161.3
R24616 plus.n15 plus.n10 161.3
R24617 plus.n18 plus.n17 161.3
R24618 plus.n19 plus.n9 161.3
R24619 plus.n21 plus.n20 161.3
R24620 plus.n23 plus.n8 161.3
R24621 plus.n25 plus.n24 161.3
R24622 plus.n27 plus.n26 161.3
R24623 plus.n28 plus.n6 161.3
R24624 plus.n30 plus.n29 161.3
R24625 plus.n32 plus.n31 161.3
R24626 plus.n33 plus.n4 161.3
R24627 plus.n36 plus.n35 161.3
R24628 plus.n37 plus.n3 161.3
R24629 plus.n39 plus.n38 161.3
R24630 plus.n41 plus.n2 161.3
R24631 plus.n43 plus.n42 161.3
R24632 plus.n45 plus.n44 161.3
R24633 plus.n46 plus.n0 161.3
R24634 plus.n48 plus.n47 161.3
R24635 plus.n64 plus.n63 56.5617
R24636 plus.n91 plus.n90 56.5617
R24637 plus.n42 plus.n41 56.5617
R24638 plus.n15 plus.n14 56.5617
R24639 plus.n73 plus.n72 56.5617
R24640 plus.n82 plus.n81 56.5617
R24641 plus.n33 plus.n32 56.5617
R24642 plus.n24 plus.n23 56.5617
R24643 plus.n95 plus.n94 48.3272
R24644 plus.n46 plus.n45 48.3272
R24645 plus.n70 plus.n58 44.4521
R24646 plus.n84 plus.n52 44.4521
R24647 plus.n35 plus.n3 44.4521
R24648 plus.n21 plus.n9 44.4521
R24649 plus.n62 plus.n61 43.0014
R24650 plus.n13 plus.n12 43.0014
R24651 plus.n77 plus.n76 40.577
R24652 plus.n78 plus.n77 40.577
R24653 plus.n29 plus.n28 40.577
R24654 plus.n28 plus.n27 40.577
R24655 plus.n61 plus.n60 39.4345
R24656 plus.n12 plus.n11 39.4345
R24657 plus.n66 plus.n58 36.702
R24658 plus.n88 plus.n52 36.702
R24659 plus.n39 plus.n3 36.702
R24660 plus.n17 plus.n9 36.702
R24661 plus.n98 plus.n97 33.3471
R24662 plus.n65 plus.n64 20.9036
R24663 plus.n90 plus.n89 20.9036
R24664 plus.n41 plus.n40 20.9036
R24665 plus.n16 plus.n15 20.9036
R24666 plus.n99 plus.t2 19.8005
R24667 plus.n99 plus.t4 19.8005
R24668 plus.n101 plus.t0 19.8005
R24669 plus.n101 plus.t3 19.8005
R24670 plus.n73 plus.n56 18.9362
R24671 plus.n81 plus.n54 18.9362
R24672 plus.n32 plus.n5 18.9362
R24673 plus.n24 plus.n7 18.9362
R24674 plus.n72 plus.n71 16.9689
R24675 plus.n83 plus.n82 16.9689
R24676 plus.n34 plus.n33 16.9689
R24677 plus.n23 plus.n22 16.9689
R24678 plus.n63 plus.n60 15.0015
R24679 plus.n91 plus.n50 15.0015
R24680 plus.n42 plus.n1 15.0015
R24681 plus.n14 plus.n11 15.0015
R24682 plus plus.n103 14.9146
R24683 plus.n96 plus.n95 12.4157
R24684 plus.n47 plus.n46 12.4157
R24685 plus.n98 plus.n48 11.9418
R24686 plus.n94 plus.n50 9.59132
R24687 plus.n45 plus.n1 9.59132
R24688 plus.n71 plus.n70 7.62397
R24689 plus.n84 plus.n83 7.62397
R24690 plus.n35 plus.n34 7.62397
R24691 plus.n22 plus.n21 7.62397
R24692 plus.n76 plus.n56 5.65662
R24693 plus.n78 plus.n54 5.65662
R24694 plus.n29 plus.n5 5.65662
R24695 plus.n27 plus.n7 5.65662
R24696 plus.n103 plus.n102 5.40567
R24697 plus.n66 plus.n65 3.68928
R24698 plus.n89 plus.n88 3.68928
R24699 plus.n40 plus.n39 3.68928
R24700 plus.n17 plus.n16 3.68928
R24701 plus.n103 plus.n98 1.188
R24702 plus.n102 plus.n100 0.716017
R24703 plus.n62 plus.n59 0.189894
R24704 plus.n67 plus.n59 0.189894
R24705 plus.n68 plus.n67 0.189894
R24706 plus.n69 plus.n68 0.189894
R24707 plus.n69 plus.n57 0.189894
R24708 plus.n74 plus.n57 0.189894
R24709 plus.n75 plus.n74 0.189894
R24710 plus.n75 plus.n55 0.189894
R24711 plus.n79 plus.n55 0.189894
R24712 plus.n80 plus.n79 0.189894
R24713 plus.n80 plus.n53 0.189894
R24714 plus.n85 plus.n53 0.189894
R24715 plus.n86 plus.n85 0.189894
R24716 plus.n87 plus.n86 0.189894
R24717 plus.n87 plus.n51 0.189894
R24718 plus.n92 plus.n51 0.189894
R24719 plus.n93 plus.n92 0.189894
R24720 plus.n93 plus.n49 0.189894
R24721 plus.n97 plus.n49 0.189894
R24722 plus.n48 plus.n0 0.189894
R24723 plus.n44 plus.n0 0.189894
R24724 plus.n44 plus.n43 0.189894
R24725 plus.n43 plus.n2 0.189894
R24726 plus.n38 plus.n2 0.189894
R24727 plus.n38 plus.n37 0.189894
R24728 plus.n37 plus.n36 0.189894
R24729 plus.n36 plus.n4 0.189894
R24730 plus.n31 plus.n4 0.189894
R24731 plus.n31 plus.n30 0.189894
R24732 plus.n30 plus.n6 0.189894
R24733 plus.n26 plus.n6 0.189894
R24734 plus.n26 plus.n25 0.189894
R24735 plus.n25 plus.n8 0.189894
R24736 plus.n20 plus.n8 0.189894
R24737 plus.n20 plus.n19 0.189894
R24738 plus.n19 plus.n18 0.189894
R24739 plus.n18 plus.n10 0.189894
R24740 plus.n13 plus.n10 0.189894
R24741 a_n2903_n3924.n18 a_n2903_n3924.t34 214.624
R24742 a_n2903_n3924.n1 a_n2903_n3924.t23 214.321
R24743 a_n2903_n3924.n12 a_n2903_n3924.t43 214.321
R24744 a_n2903_n3924.n13 a_n2903_n3924.t46 214.321
R24745 a_n2903_n3924.n14 a_n2903_n3924.t29 214.321
R24746 a_n2903_n3924.n15 a_n2903_n3924.t37 214.321
R24747 a_n2903_n3924.n16 a_n2903_n3924.t35 214.321
R24748 a_n2903_n3924.n17 a_n2903_n3924.t26 214.321
R24749 a_n2903_n3924.n0 a_n2903_n3924.t14 55.8337
R24750 a_n2903_n3924.n2 a_n2903_n3924.t39 55.8337
R24751 a_n2903_n3924.n11 a_n2903_n3924.t21 55.8337
R24752 a_n2903_n3924.n41 a_n2903_n3924.t2 55.8335
R24753 a_n2903_n3924.n39 a_n2903_n3924.t36 55.8335
R24754 a_n2903_n3924.n30 a_n2903_n3924.t24 55.8335
R24755 a_n2903_n3924.n29 a_n2903_n3924.t11 55.8335
R24756 a_n2903_n3924.n20 a_n2903_n3924.t19 55.8335
R24757 a_n2903_n3924.n43 a_n2903_n3924.n42 53.0052
R24758 a_n2903_n3924.n45 a_n2903_n3924.n44 53.0052
R24759 a_n2903_n3924.n47 a_n2903_n3924.n46 53.0052
R24760 a_n2903_n3924.n4 a_n2903_n3924.n3 53.0052
R24761 a_n2903_n3924.n6 a_n2903_n3924.n5 53.0052
R24762 a_n2903_n3924.n8 a_n2903_n3924.n7 53.0052
R24763 a_n2903_n3924.n10 a_n2903_n3924.n9 53.0052
R24764 a_n2903_n3924.n38 a_n2903_n3924.n37 53.0051
R24765 a_n2903_n3924.n36 a_n2903_n3924.n35 53.0051
R24766 a_n2903_n3924.n34 a_n2903_n3924.n33 53.0051
R24767 a_n2903_n3924.n32 a_n2903_n3924.n31 53.0051
R24768 a_n2903_n3924.n28 a_n2903_n3924.n27 53.0051
R24769 a_n2903_n3924.n26 a_n2903_n3924.n25 53.0051
R24770 a_n2903_n3924.n24 a_n2903_n3924.n23 53.0051
R24771 a_n2903_n3924.n22 a_n2903_n3924.n21 53.0051
R24772 a_n2903_n3924.n49 a_n2903_n3924.n48 53.0051
R24773 a_n2903_n3924.n19 a_n2903_n3924.n11 12.2417
R24774 a_n2903_n3924.n41 a_n2903_n3924.n40 12.2417
R24775 a_n2903_n3924.n20 a_n2903_n3924.n19 5.16214
R24776 a_n2903_n3924.n40 a_n2903_n3924.n39 5.16214
R24777 a_n2903_n3924.n42 a_n2903_n3924.t10 2.82907
R24778 a_n2903_n3924.n42 a_n2903_n3924.t15 2.82907
R24779 a_n2903_n3924.n44 a_n2903_n3924.t8 2.82907
R24780 a_n2903_n3924.n44 a_n2903_n3924.t12 2.82907
R24781 a_n2903_n3924.n46 a_n2903_n3924.t5 2.82907
R24782 a_n2903_n3924.n46 a_n2903_n3924.t9 2.82907
R24783 a_n2903_n3924.n3 a_n2903_n3924.t30 2.82907
R24784 a_n2903_n3924.n3 a_n2903_n3924.t44 2.82907
R24785 a_n2903_n3924.n5 a_n2903_n3924.t25 2.82907
R24786 a_n2903_n3924.n5 a_n2903_n3924.t31 2.82907
R24787 a_n2903_n3924.n7 a_n2903_n3924.t40 2.82907
R24788 a_n2903_n3924.n7 a_n2903_n3924.t28 2.82907
R24789 a_n2903_n3924.n9 a_n2903_n3924.t47 2.82907
R24790 a_n2903_n3924.n9 a_n2903_n3924.t32 2.82907
R24791 a_n2903_n3924.n37 a_n2903_n3924.t38 2.82907
R24792 a_n2903_n3924.n37 a_n2903_n3924.t33 2.82907
R24793 a_n2903_n3924.n35 a_n2903_n3924.t27 2.82907
R24794 a_n2903_n3924.n35 a_n2903_n3924.t41 2.82907
R24795 a_n2903_n3924.n33 a_n2903_n3924.t42 2.82907
R24796 a_n2903_n3924.n33 a_n2903_n3924.t22 2.82907
R24797 a_n2903_n3924.n31 a_n2903_n3924.t45 2.82907
R24798 a_n2903_n3924.n31 a_n2903_n3924.t0 2.82907
R24799 a_n2903_n3924.n27 a_n2903_n3924.t3 2.82907
R24800 a_n2903_n3924.n27 a_n2903_n3924.t16 2.82907
R24801 a_n2903_n3924.n25 a_n2903_n3924.t7 2.82907
R24802 a_n2903_n3924.n25 a_n2903_n3924.t1 2.82907
R24803 a_n2903_n3924.n23 a_n2903_n3924.t18 2.82907
R24804 a_n2903_n3924.n23 a_n2903_n3924.t6 2.82907
R24805 a_n2903_n3924.n21 a_n2903_n3924.t13 2.82907
R24806 a_n2903_n3924.n21 a_n2903_n3924.t17 2.82907
R24807 a_n2903_n3924.t20 a_n2903_n3924.n49 2.82907
R24808 a_n2903_n3924.n49 a_n2903_n3924.t4 2.82907
R24809 a_n2903_n3924.n40 a_n2903_n3924.n1 2.18441
R24810 a_n2903_n3924.n19 a_n2903_n3924.n18 1.95694
R24811 a_n2903_n3924.n17 a_n2903_n3924.n16 0.672012
R24812 a_n2903_n3924.n16 a_n2903_n3924.n15 0.672012
R24813 a_n2903_n3924.n15 a_n2903_n3924.n14 0.672012
R24814 a_n2903_n3924.n14 a_n2903_n3924.n13 0.672012
R24815 a_n2903_n3924.n13 a_n2903_n3924.n12 0.672012
R24816 a_n2903_n3924.n12 a_n2903_n3924.n1 0.672012
R24817 a_n2903_n3924.n22 a_n2903_n3924.n20 0.530672
R24818 a_n2903_n3924.n24 a_n2903_n3924.n22 0.530672
R24819 a_n2903_n3924.n26 a_n2903_n3924.n24 0.530672
R24820 a_n2903_n3924.n28 a_n2903_n3924.n26 0.530672
R24821 a_n2903_n3924.n29 a_n2903_n3924.n28 0.530672
R24822 a_n2903_n3924.n32 a_n2903_n3924.n30 0.530672
R24823 a_n2903_n3924.n34 a_n2903_n3924.n32 0.530672
R24824 a_n2903_n3924.n36 a_n2903_n3924.n34 0.530672
R24825 a_n2903_n3924.n38 a_n2903_n3924.n36 0.530672
R24826 a_n2903_n3924.n39 a_n2903_n3924.n38 0.530672
R24827 a_n2903_n3924.n11 a_n2903_n3924.n10 0.530672
R24828 a_n2903_n3924.n10 a_n2903_n3924.n8 0.530672
R24829 a_n2903_n3924.n8 a_n2903_n3924.n6 0.530672
R24830 a_n2903_n3924.n6 a_n2903_n3924.n4 0.530672
R24831 a_n2903_n3924.n4 a_n2903_n3924.n2 0.530672
R24832 a_n2903_n3924.n48 a_n2903_n3924.n0 0.530672
R24833 a_n2903_n3924.n48 a_n2903_n3924.n47 0.530672
R24834 a_n2903_n3924.n47 a_n2903_n3924.n45 0.530672
R24835 a_n2903_n3924.n45 a_n2903_n3924.n43 0.530672
R24836 a_n2903_n3924.n43 a_n2903_n3924.n41 0.530672
R24837 a_n2903_n3924.n18 a_n2903_n3924.n17 0.370413
R24838 a_n2903_n3924.n30 a_n2903_n3924.n29 0.235414
R24839 a_n2903_n3924.n2 a_n2903_n3924.n0 0.235414
R24840 a_n2982_8322.n12 a_n2982_8322.t33 74.6477
R24841 a_n2982_8322.n1 a_n2982_8322.t12 74.6477
R24842 a_n2982_8322.n28 a_n2982_8322.t27 74.6474
R24843 a_n2982_8322.n20 a_n2982_8322.t7 74.2899
R24844 a_n2982_8322.n13 a_n2982_8322.t31 74.2899
R24845 a_n2982_8322.n14 a_n2982_8322.t34 74.2899
R24846 a_n2982_8322.n17 a_n2982_8322.t35 74.2899
R24847 a_n2982_8322.n10 a_n2982_8322.t6 74.2899
R24848 a_n2982_8322.n28 a_n2982_8322.n27 70.6783
R24849 a_n2982_8322.n26 a_n2982_8322.n25 70.6783
R24850 a_n2982_8322.n24 a_n2982_8322.n23 70.6783
R24851 a_n2982_8322.n22 a_n2982_8322.n21 70.6783
R24852 a_n2982_8322.n12 a_n2982_8322.n11 70.6783
R24853 a_n2982_8322.n16 a_n2982_8322.n15 70.6783
R24854 a_n2982_8322.n1 a_n2982_8322.n0 70.6783
R24855 a_n2982_8322.n3 a_n2982_8322.n2 70.6783
R24856 a_n2982_8322.n5 a_n2982_8322.n4 70.6783
R24857 a_n2982_8322.n7 a_n2982_8322.n6 70.6783
R24858 a_n2982_8322.n9 a_n2982_8322.n8 70.6783
R24859 a_n2982_8322.n30 a_n2982_8322.n29 70.6782
R24860 a_n2982_8322.n18 a_n2982_8322.n10 24.9022
R24861 a_n2982_8322.n19 a_n2982_8322.t5 9.81851
R24862 a_n2982_8322.n18 a_n2982_8322.n17 8.38735
R24863 a_n2982_8322.n20 a_n2982_8322.n19 6.90998
R24864 a_n2982_8322.n19 a_n2982_8322.n18 5.3452
R24865 a_n2982_8322.n27 a_n2982_8322.t20 3.61217
R24866 a_n2982_8322.n27 a_n2982_8322.t16 3.61217
R24867 a_n2982_8322.n25 a_n2982_8322.t26 3.61217
R24868 a_n2982_8322.n25 a_n2982_8322.t14 3.61217
R24869 a_n2982_8322.n23 a_n2982_8322.t11 3.61217
R24870 a_n2982_8322.n23 a_n2982_8322.t10 3.61217
R24871 a_n2982_8322.n21 a_n2982_8322.t24 3.61217
R24872 a_n2982_8322.n21 a_n2982_8322.t23 3.61217
R24873 a_n2982_8322.n11 a_n2982_8322.t37 3.61217
R24874 a_n2982_8322.n11 a_n2982_8322.t36 3.61217
R24875 a_n2982_8322.n15 a_n2982_8322.t32 3.61217
R24876 a_n2982_8322.n15 a_n2982_8322.t30 3.61217
R24877 a_n2982_8322.n0 a_n2982_8322.t25 3.61217
R24878 a_n2982_8322.n0 a_n2982_8322.t21 3.61217
R24879 a_n2982_8322.n2 a_n2982_8322.t28 3.61217
R24880 a_n2982_8322.n2 a_n2982_8322.t18 3.61217
R24881 a_n2982_8322.n4 a_n2982_8322.t9 3.61217
R24882 a_n2982_8322.n4 a_n2982_8322.t8 3.61217
R24883 a_n2982_8322.n6 a_n2982_8322.t22 3.61217
R24884 a_n2982_8322.n6 a_n2982_8322.t15 3.61217
R24885 a_n2982_8322.n8 a_n2982_8322.t19 3.61217
R24886 a_n2982_8322.n8 a_n2982_8322.t17 3.61217
R24887 a_n2982_8322.n30 a_n2982_8322.t13 3.61217
R24888 a_n2982_8322.t29 a_n2982_8322.n30 3.61217
R24889 a_n2982_8322.n17 a_n2982_8322.n16 0.358259
R24890 a_n2982_8322.n16 a_n2982_8322.n14 0.358259
R24891 a_n2982_8322.n13 a_n2982_8322.n12 0.358259
R24892 a_n2982_8322.n10 a_n2982_8322.n9 0.358259
R24893 a_n2982_8322.n9 a_n2982_8322.n7 0.358259
R24894 a_n2982_8322.n7 a_n2982_8322.n5 0.358259
R24895 a_n2982_8322.n5 a_n2982_8322.n3 0.358259
R24896 a_n2982_8322.n3 a_n2982_8322.n1 0.358259
R24897 a_n2982_8322.n22 a_n2982_8322.n20 0.358259
R24898 a_n2982_8322.n24 a_n2982_8322.n22 0.358259
R24899 a_n2982_8322.n26 a_n2982_8322.n24 0.358259
R24900 a_n2982_8322.n29 a_n2982_8322.n26 0.358259
R24901 a_n2982_8322.n29 a_n2982_8322.n28 0.358259
R24902 a_n2982_8322.n14 a_n2982_8322.n13 0.101793
R24903 a_n2982_8322.t4 a_n2982_8322.t2 0.0788333
R24904 a_n2982_8322.t0 a_n2982_8322.t1 0.0788333
R24905 a_n2982_8322.t5 a_n2982_8322.t3 0.0788333
R24906 a_n2982_8322.t0 a_n2982_8322.t4 0.0318333
R24907 a_n2982_8322.t5 a_n2982_8322.t1 0.0318333
R24908 a_n2982_8322.t2 a_n2982_8322.t1 0.0318333
R24909 a_n2982_8322.t3 a_n2982_8322.t0 0.0318333
R24910 output.n41 output.n15 289.615
R24911 output.n72 output.n46 289.615
R24912 output.n104 output.n78 289.615
R24913 output.n136 output.n110 289.615
R24914 output.n77 output.n45 197.26
R24915 output.n77 output.n76 196.298
R24916 output.n109 output.n108 196.298
R24917 output.n141 output.n140 196.298
R24918 output.n42 output.n41 185
R24919 output.n40 output.n39 185
R24920 output.n19 output.n18 185
R24921 output.n34 output.n33 185
R24922 output.n32 output.n31 185
R24923 output.n23 output.n22 185
R24924 output.n26 output.n25 185
R24925 output.n73 output.n72 185
R24926 output.n71 output.n70 185
R24927 output.n50 output.n49 185
R24928 output.n65 output.n64 185
R24929 output.n63 output.n62 185
R24930 output.n54 output.n53 185
R24931 output.n57 output.n56 185
R24932 output.n105 output.n104 185
R24933 output.n103 output.n102 185
R24934 output.n82 output.n81 185
R24935 output.n97 output.n96 185
R24936 output.n95 output.n94 185
R24937 output.n86 output.n85 185
R24938 output.n89 output.n88 185
R24939 output.n137 output.n136 185
R24940 output.n135 output.n134 185
R24941 output.n114 output.n113 185
R24942 output.n129 output.n128 185
R24943 output.n127 output.n126 185
R24944 output.n118 output.n117 185
R24945 output.n121 output.n120 185
R24946 output.t18 output.n24 147.661
R24947 output.t17 output.n55 147.661
R24948 output.t16 output.n87 147.661
R24949 output.t19 output.n119 147.661
R24950 output.n41 output.n40 104.615
R24951 output.n40 output.n18 104.615
R24952 output.n33 output.n18 104.615
R24953 output.n33 output.n32 104.615
R24954 output.n32 output.n22 104.615
R24955 output.n25 output.n22 104.615
R24956 output.n72 output.n71 104.615
R24957 output.n71 output.n49 104.615
R24958 output.n64 output.n49 104.615
R24959 output.n64 output.n63 104.615
R24960 output.n63 output.n53 104.615
R24961 output.n56 output.n53 104.615
R24962 output.n104 output.n103 104.615
R24963 output.n103 output.n81 104.615
R24964 output.n96 output.n81 104.615
R24965 output.n96 output.n95 104.615
R24966 output.n95 output.n85 104.615
R24967 output.n88 output.n85 104.615
R24968 output.n136 output.n135 104.615
R24969 output.n135 output.n113 104.615
R24970 output.n128 output.n113 104.615
R24971 output.n128 output.n127 104.615
R24972 output.n127 output.n117 104.615
R24973 output.n120 output.n117 104.615
R24974 output.n1 output.t0 77.056
R24975 output.n14 output.t1 76.6694
R24976 output.n1 output.n0 72.7095
R24977 output.n3 output.n2 72.7095
R24978 output.n5 output.n4 72.7095
R24979 output.n7 output.n6 72.7095
R24980 output.n9 output.n8 72.7095
R24981 output.n11 output.n10 72.7095
R24982 output.n13 output.n12 72.7095
R24983 output.n25 output.t18 52.3082
R24984 output.n56 output.t17 52.3082
R24985 output.n88 output.t16 52.3082
R24986 output.n120 output.t19 52.3082
R24987 output.n26 output.n24 15.6674
R24988 output.n57 output.n55 15.6674
R24989 output.n89 output.n87 15.6674
R24990 output.n121 output.n119 15.6674
R24991 output.n27 output.n23 12.8005
R24992 output.n58 output.n54 12.8005
R24993 output.n90 output.n86 12.8005
R24994 output.n122 output.n118 12.8005
R24995 output.n31 output.n30 12.0247
R24996 output.n62 output.n61 12.0247
R24997 output.n94 output.n93 12.0247
R24998 output.n126 output.n125 12.0247
R24999 output.n34 output.n21 11.249
R25000 output.n65 output.n52 11.249
R25001 output.n97 output.n84 11.249
R25002 output.n129 output.n116 11.249
R25003 output.n35 output.n19 10.4732
R25004 output.n66 output.n50 10.4732
R25005 output.n98 output.n82 10.4732
R25006 output.n130 output.n114 10.4732
R25007 output.n39 output.n38 9.69747
R25008 output.n70 output.n69 9.69747
R25009 output.n102 output.n101 9.69747
R25010 output.n134 output.n133 9.69747
R25011 output.n45 output.n44 9.45567
R25012 output.n76 output.n75 9.45567
R25013 output.n108 output.n107 9.45567
R25014 output.n140 output.n139 9.45567
R25015 output.n44 output.n43 9.3005
R25016 output.n17 output.n16 9.3005
R25017 output.n38 output.n37 9.3005
R25018 output.n36 output.n35 9.3005
R25019 output.n21 output.n20 9.3005
R25020 output.n30 output.n29 9.3005
R25021 output.n28 output.n27 9.3005
R25022 output.n75 output.n74 9.3005
R25023 output.n48 output.n47 9.3005
R25024 output.n69 output.n68 9.3005
R25025 output.n67 output.n66 9.3005
R25026 output.n52 output.n51 9.3005
R25027 output.n61 output.n60 9.3005
R25028 output.n59 output.n58 9.3005
R25029 output.n107 output.n106 9.3005
R25030 output.n80 output.n79 9.3005
R25031 output.n101 output.n100 9.3005
R25032 output.n99 output.n98 9.3005
R25033 output.n84 output.n83 9.3005
R25034 output.n93 output.n92 9.3005
R25035 output.n91 output.n90 9.3005
R25036 output.n139 output.n138 9.3005
R25037 output.n112 output.n111 9.3005
R25038 output.n133 output.n132 9.3005
R25039 output.n131 output.n130 9.3005
R25040 output.n116 output.n115 9.3005
R25041 output.n125 output.n124 9.3005
R25042 output.n123 output.n122 9.3005
R25043 output.n42 output.n17 8.92171
R25044 output.n73 output.n48 8.92171
R25045 output.n105 output.n80 8.92171
R25046 output.n137 output.n112 8.92171
R25047 output output.n141 8.15037
R25048 output.n43 output.n15 8.14595
R25049 output.n74 output.n46 8.14595
R25050 output.n106 output.n78 8.14595
R25051 output.n138 output.n110 8.14595
R25052 output.n45 output.n15 5.81868
R25053 output.n76 output.n46 5.81868
R25054 output.n108 output.n78 5.81868
R25055 output.n140 output.n110 5.81868
R25056 output.n43 output.n42 5.04292
R25057 output.n74 output.n73 5.04292
R25058 output.n106 output.n105 5.04292
R25059 output.n138 output.n137 5.04292
R25060 output.n28 output.n24 4.38594
R25061 output.n59 output.n55 4.38594
R25062 output.n91 output.n87 4.38594
R25063 output.n123 output.n119 4.38594
R25064 output.n39 output.n17 4.26717
R25065 output.n70 output.n48 4.26717
R25066 output.n102 output.n80 4.26717
R25067 output.n134 output.n112 4.26717
R25068 output.n0 output.t10 3.9605
R25069 output.n0 output.t8 3.9605
R25070 output.n2 output.t15 3.9605
R25071 output.n2 output.t2 3.9605
R25072 output.n4 output.t4 3.9605
R25073 output.n4 output.t12 3.9605
R25074 output.n6 output.t14 3.9605
R25075 output.n6 output.t5 3.9605
R25076 output.n8 output.t6 3.9605
R25077 output.n8 output.t11 3.9605
R25078 output.n10 output.t13 3.9605
R25079 output.n10 output.t3 3.9605
R25080 output.n12 output.t9 3.9605
R25081 output.n12 output.t7 3.9605
R25082 output.n38 output.n19 3.49141
R25083 output.n69 output.n50 3.49141
R25084 output.n101 output.n82 3.49141
R25085 output.n133 output.n114 3.49141
R25086 output.n35 output.n34 2.71565
R25087 output.n66 output.n65 2.71565
R25088 output.n98 output.n97 2.71565
R25089 output.n130 output.n129 2.71565
R25090 output.n31 output.n21 1.93989
R25091 output.n62 output.n52 1.93989
R25092 output.n94 output.n84 1.93989
R25093 output.n126 output.n116 1.93989
R25094 output.n30 output.n23 1.16414
R25095 output.n61 output.n54 1.16414
R25096 output.n93 output.n86 1.16414
R25097 output.n125 output.n118 1.16414
R25098 output.n141 output.n109 0.962709
R25099 output.n109 output.n77 0.962709
R25100 output.n27 output.n26 0.388379
R25101 output.n58 output.n57 0.388379
R25102 output.n90 output.n89 0.388379
R25103 output.n122 output.n121 0.388379
R25104 output.n14 output.n13 0.387128
R25105 output.n13 output.n11 0.387128
R25106 output.n11 output.n9 0.387128
R25107 output.n9 output.n7 0.387128
R25108 output.n7 output.n5 0.387128
R25109 output.n5 output.n3 0.387128
R25110 output.n3 output.n1 0.387128
R25111 output.n44 output.n16 0.155672
R25112 output.n37 output.n16 0.155672
R25113 output.n37 output.n36 0.155672
R25114 output.n36 output.n20 0.155672
R25115 output.n29 output.n20 0.155672
R25116 output.n29 output.n28 0.155672
R25117 output.n75 output.n47 0.155672
R25118 output.n68 output.n47 0.155672
R25119 output.n68 output.n67 0.155672
R25120 output.n67 output.n51 0.155672
R25121 output.n60 output.n51 0.155672
R25122 output.n60 output.n59 0.155672
R25123 output.n107 output.n79 0.155672
R25124 output.n100 output.n79 0.155672
R25125 output.n100 output.n99 0.155672
R25126 output.n99 output.n83 0.155672
R25127 output.n92 output.n83 0.155672
R25128 output.n92 output.n91 0.155672
R25129 output.n139 output.n111 0.155672
R25130 output.n132 output.n111 0.155672
R25131 output.n132 output.n131 0.155672
R25132 output.n131 output.n115 0.155672
R25133 output.n124 output.n115 0.155672
R25134 output.n124 output.n123 0.155672
R25135 output output.n14 0.126227
R25136 minus.n61 minus.t24 251.488
R25137 minus.n12 minus.t16 251.488
R25138 minus.n102 minus.t4 243.255
R25139 minus.n96 minus.t14 231.093
R25140 minus.n47 minus.t9 231.093
R25141 minus.n101 minus.n99 224.169
R25142 minus.n101 minus.n100 223.454
R25143 minus.n50 minus.t21 187.445
R25144 minus.n89 minus.t18 187.445
R25145 minus.n83 minus.t15 187.445
R25146 minus.n54 minus.t7 187.445
R25147 minus.n56 minus.t6 187.445
R25148 minus.n71 minus.t12 187.445
R25149 minus.n65 minus.t11 187.445
R25150 minus.n60 minus.t19 187.445
R25151 minus.n11 minus.t10 187.445
R25152 minus.n16 minus.t8 187.445
R25153 minus.n22 minus.t5 187.445
R25154 minus.n7 minus.t22 187.445
R25155 minus.n5 minus.t23 187.445
R25156 minus.n34 minus.t17 187.445
R25157 minus.n40 minus.t20 187.445
R25158 minus.n1 minus.t13 187.445
R25159 minus.n63 minus.n62 161.3
R25160 minus.n64 minus.n59 161.3
R25161 minus.n67 minus.n66 161.3
R25162 minus.n68 minus.n58 161.3
R25163 minus.n70 minus.n69 161.3
R25164 minus.n72 minus.n57 161.3
R25165 minus.n74 minus.n73 161.3
R25166 minus.n76 minus.n75 161.3
R25167 minus.n77 minus.n55 161.3
R25168 minus.n79 minus.n78 161.3
R25169 minus.n81 minus.n80 161.3
R25170 minus.n82 minus.n53 161.3
R25171 minus.n85 minus.n84 161.3
R25172 minus.n86 minus.n52 161.3
R25173 minus.n88 minus.n87 161.3
R25174 minus.n90 minus.n51 161.3
R25175 minus.n92 minus.n91 161.3
R25176 minus.n94 minus.n93 161.3
R25177 minus.n95 minus.n49 161.3
R25178 minus.n97 minus.n96 161.3
R25179 minus.n48 minus.n47 161.3
R25180 minus.n46 minus.n0 161.3
R25181 minus.n45 minus.n44 161.3
R25182 minus.n43 minus.n42 161.3
R25183 minus.n41 minus.n2 161.3
R25184 minus.n39 minus.n38 161.3
R25185 minus.n37 minus.n3 161.3
R25186 minus.n36 minus.n35 161.3
R25187 minus.n33 minus.n4 161.3
R25188 minus.n32 minus.n31 161.3
R25189 minus.n30 minus.n29 161.3
R25190 minus.n28 minus.n6 161.3
R25191 minus.n27 minus.n26 161.3
R25192 minus.n25 minus.n24 161.3
R25193 minus.n23 minus.n8 161.3
R25194 minus.n21 minus.n20 161.3
R25195 minus.n19 minus.n9 161.3
R25196 minus.n18 minus.n17 161.3
R25197 minus.n15 minus.n10 161.3
R25198 minus.n14 minus.n13 161.3
R25199 minus.n91 minus.n90 56.5617
R25200 minus.n64 minus.n63 56.5617
R25201 minus.n15 minus.n14 56.5617
R25202 minus.n42 minus.n41 56.5617
R25203 minus.n82 minus.n81 56.5617
R25204 minus.n73 minus.n72 56.5617
R25205 minus.n24 minus.n23 56.5617
R25206 minus.n33 minus.n32 56.5617
R25207 minus.n95 minus.n94 48.3272
R25208 minus.n46 minus.n45 48.3272
R25209 minus.n84 minus.n52 44.4521
R25210 minus.n70 minus.n58 44.4521
R25211 minus.n21 minus.n9 44.4521
R25212 minus.n35 minus.n3 44.4521
R25213 minus.n13 minus.n12 43.0014
R25214 minus.n62 minus.n61 43.0014
R25215 minus.n78 minus.n77 40.577
R25216 minus.n77 minus.n76 40.577
R25217 minus.n28 minus.n27 40.577
R25218 minus.n29 minus.n28 40.577
R25219 minus.n61 minus.n60 39.4345
R25220 minus.n12 minus.n11 39.4345
R25221 minus.n88 minus.n52 36.702
R25222 minus.n66 minus.n58 36.702
R25223 minus.n17 minus.n9 36.702
R25224 minus.n39 minus.n3 36.702
R25225 minus.n98 minus.n97 33.563
R25226 minus.n90 minus.n89 20.9036
R25227 minus.n65 minus.n64 20.9036
R25228 minus.n16 minus.n15 20.9036
R25229 minus.n41 minus.n40 20.9036
R25230 minus.n100 minus.t3 19.8005
R25231 minus.n100 minus.t0 19.8005
R25232 minus.n99 minus.t2 19.8005
R25233 minus.n99 minus.t1 19.8005
R25234 minus.n81 minus.n54 18.9362
R25235 minus.n73 minus.n56 18.9362
R25236 minus.n24 minus.n7 18.9362
R25237 minus.n32 minus.n5 18.9362
R25238 minus.n83 minus.n82 16.9689
R25239 minus.n72 minus.n71 16.9689
R25240 minus.n23 minus.n22 16.9689
R25241 minus.n34 minus.n33 16.9689
R25242 minus.n91 minus.n50 15.0015
R25243 minus.n63 minus.n60 15.0015
R25244 minus.n14 minus.n11 15.0015
R25245 minus.n42 minus.n1 15.0015
R25246 minus.n96 minus.n95 12.4157
R25247 minus.n47 minus.n46 12.4157
R25248 minus.n98 minus.n48 12.1577
R25249 minus minus.n103 11.7349
R25250 minus.n94 minus.n50 9.59132
R25251 minus.n45 minus.n1 9.59132
R25252 minus.n84 minus.n83 7.62397
R25253 minus.n71 minus.n70 7.62397
R25254 minus.n22 minus.n21 7.62397
R25255 minus.n35 minus.n34 7.62397
R25256 minus.n78 minus.n54 5.65662
R25257 minus.n76 minus.n56 5.65662
R25258 minus.n27 minus.n7 5.65662
R25259 minus.n29 minus.n5 5.65662
R25260 minus.n103 minus.n102 4.80222
R25261 minus.n89 minus.n88 3.68928
R25262 minus.n66 minus.n65 3.68928
R25263 minus.n17 minus.n16 3.68928
R25264 minus.n40 minus.n39 3.68928
R25265 minus.n103 minus.n98 0.972091
R25266 minus.n102 minus.n101 0.716017
R25267 minus.n97 minus.n49 0.189894
R25268 minus.n93 minus.n49 0.189894
R25269 minus.n93 minus.n92 0.189894
R25270 minus.n92 minus.n51 0.189894
R25271 minus.n87 minus.n51 0.189894
R25272 minus.n87 minus.n86 0.189894
R25273 minus.n86 minus.n85 0.189894
R25274 minus.n85 minus.n53 0.189894
R25275 minus.n80 minus.n53 0.189894
R25276 minus.n80 minus.n79 0.189894
R25277 minus.n79 minus.n55 0.189894
R25278 minus.n75 minus.n55 0.189894
R25279 minus.n75 minus.n74 0.189894
R25280 minus.n74 minus.n57 0.189894
R25281 minus.n69 minus.n57 0.189894
R25282 minus.n69 minus.n68 0.189894
R25283 minus.n68 minus.n67 0.189894
R25284 minus.n67 minus.n59 0.189894
R25285 minus.n62 minus.n59 0.189894
R25286 minus.n13 minus.n10 0.189894
R25287 minus.n18 minus.n10 0.189894
R25288 minus.n19 minus.n18 0.189894
R25289 minus.n20 minus.n19 0.189894
R25290 minus.n20 minus.n8 0.189894
R25291 minus.n25 minus.n8 0.189894
R25292 minus.n26 minus.n25 0.189894
R25293 minus.n26 minus.n6 0.189894
R25294 minus.n30 minus.n6 0.189894
R25295 minus.n31 minus.n30 0.189894
R25296 minus.n31 minus.n4 0.189894
R25297 minus.n36 minus.n4 0.189894
R25298 minus.n37 minus.n36 0.189894
R25299 minus.n38 minus.n37 0.189894
R25300 minus.n38 minus.n2 0.189894
R25301 minus.n43 minus.n2 0.189894
R25302 minus.n44 minus.n43 0.189894
R25303 minus.n44 minus.n0 0.189894
R25304 minus.n48 minus.n0 0.189894
R25305 diffpairibias.n0 diffpairibias.t18 436.822
R25306 diffpairibias.n21 diffpairibias.t19 435.479
R25307 diffpairibias.n20 diffpairibias.t16 435.479
R25308 diffpairibias.n19 diffpairibias.t17 435.479
R25309 diffpairibias.n18 diffpairibias.t21 435.479
R25310 diffpairibias.n0 diffpairibias.t22 435.479
R25311 diffpairibias.n1 diffpairibias.t20 435.479
R25312 diffpairibias.n2 diffpairibias.t23 435.479
R25313 diffpairibias.n10 diffpairibias.t0 377.536
R25314 diffpairibias.n10 diffpairibias.t8 376.193
R25315 diffpairibias.n11 diffpairibias.t10 376.193
R25316 diffpairibias.n12 diffpairibias.t6 376.193
R25317 diffpairibias.n13 diffpairibias.t2 376.193
R25318 diffpairibias.n14 diffpairibias.t12 376.193
R25319 diffpairibias.n15 diffpairibias.t4 376.193
R25320 diffpairibias.n16 diffpairibias.t14 376.193
R25321 diffpairibias.n3 diffpairibias.t1 113.368
R25322 diffpairibias.n3 diffpairibias.t9 112.698
R25323 diffpairibias.n4 diffpairibias.t11 112.698
R25324 diffpairibias.n5 diffpairibias.t7 112.698
R25325 diffpairibias.n6 diffpairibias.t3 112.698
R25326 diffpairibias.n7 diffpairibias.t13 112.698
R25327 diffpairibias.n8 diffpairibias.t5 112.698
R25328 diffpairibias.n9 diffpairibias.t15 112.698
R25329 diffpairibias.n17 diffpairibias.n16 4.77242
R25330 diffpairibias.n17 diffpairibias.n9 4.30807
R25331 diffpairibias.n18 diffpairibias.n17 4.13945
R25332 diffpairibias.n16 diffpairibias.n15 1.34352
R25333 diffpairibias.n15 diffpairibias.n14 1.34352
R25334 diffpairibias.n14 diffpairibias.n13 1.34352
R25335 diffpairibias.n13 diffpairibias.n12 1.34352
R25336 diffpairibias.n12 diffpairibias.n11 1.34352
R25337 diffpairibias.n11 diffpairibias.n10 1.34352
R25338 diffpairibias.n2 diffpairibias.n1 1.34352
R25339 diffpairibias.n1 diffpairibias.n0 1.34352
R25340 diffpairibias.n19 diffpairibias.n18 1.34352
R25341 diffpairibias.n20 diffpairibias.n19 1.34352
R25342 diffpairibias.n21 diffpairibias.n20 1.34352
R25343 diffpairibias.n22 diffpairibias.n21 0.862419
R25344 diffpairibias diffpairibias.n22 0.684875
R25345 diffpairibias.n9 diffpairibias.n8 0.672012
R25346 diffpairibias.n8 diffpairibias.n7 0.672012
R25347 diffpairibias.n7 diffpairibias.n6 0.672012
R25348 diffpairibias.n6 diffpairibias.n5 0.672012
R25349 diffpairibias.n5 diffpairibias.n4 0.672012
R25350 diffpairibias.n4 diffpairibias.n3 0.672012
R25351 diffpairibias.n22 diffpairibias.n2 0.190907
R25352 outputibias.n27 outputibias.n1 289.615
R25353 outputibias.n58 outputibias.n32 289.615
R25354 outputibias.n90 outputibias.n64 289.615
R25355 outputibias.n122 outputibias.n96 289.615
R25356 outputibias.n28 outputibias.n27 185
R25357 outputibias.n26 outputibias.n25 185
R25358 outputibias.n5 outputibias.n4 185
R25359 outputibias.n20 outputibias.n19 185
R25360 outputibias.n18 outputibias.n17 185
R25361 outputibias.n9 outputibias.n8 185
R25362 outputibias.n12 outputibias.n11 185
R25363 outputibias.n59 outputibias.n58 185
R25364 outputibias.n57 outputibias.n56 185
R25365 outputibias.n36 outputibias.n35 185
R25366 outputibias.n51 outputibias.n50 185
R25367 outputibias.n49 outputibias.n48 185
R25368 outputibias.n40 outputibias.n39 185
R25369 outputibias.n43 outputibias.n42 185
R25370 outputibias.n91 outputibias.n90 185
R25371 outputibias.n89 outputibias.n88 185
R25372 outputibias.n68 outputibias.n67 185
R25373 outputibias.n83 outputibias.n82 185
R25374 outputibias.n81 outputibias.n80 185
R25375 outputibias.n72 outputibias.n71 185
R25376 outputibias.n75 outputibias.n74 185
R25377 outputibias.n123 outputibias.n122 185
R25378 outputibias.n121 outputibias.n120 185
R25379 outputibias.n100 outputibias.n99 185
R25380 outputibias.n115 outputibias.n114 185
R25381 outputibias.n113 outputibias.n112 185
R25382 outputibias.n104 outputibias.n103 185
R25383 outputibias.n107 outputibias.n106 185
R25384 outputibias.n0 outputibias.t8 178.945
R25385 outputibias.n133 outputibias.t11 177.018
R25386 outputibias.n132 outputibias.t9 177.018
R25387 outputibias.n0 outputibias.t10 177.018
R25388 outputibias.t7 outputibias.n10 147.661
R25389 outputibias.t1 outputibias.n41 147.661
R25390 outputibias.t3 outputibias.n73 147.661
R25391 outputibias.t5 outputibias.n105 147.661
R25392 outputibias.n128 outputibias.t6 132.363
R25393 outputibias.n128 outputibias.t0 130.436
R25394 outputibias.n129 outputibias.t2 130.436
R25395 outputibias.n130 outputibias.t4 130.436
R25396 outputibias.n27 outputibias.n26 104.615
R25397 outputibias.n26 outputibias.n4 104.615
R25398 outputibias.n19 outputibias.n4 104.615
R25399 outputibias.n19 outputibias.n18 104.615
R25400 outputibias.n18 outputibias.n8 104.615
R25401 outputibias.n11 outputibias.n8 104.615
R25402 outputibias.n58 outputibias.n57 104.615
R25403 outputibias.n57 outputibias.n35 104.615
R25404 outputibias.n50 outputibias.n35 104.615
R25405 outputibias.n50 outputibias.n49 104.615
R25406 outputibias.n49 outputibias.n39 104.615
R25407 outputibias.n42 outputibias.n39 104.615
R25408 outputibias.n90 outputibias.n89 104.615
R25409 outputibias.n89 outputibias.n67 104.615
R25410 outputibias.n82 outputibias.n67 104.615
R25411 outputibias.n82 outputibias.n81 104.615
R25412 outputibias.n81 outputibias.n71 104.615
R25413 outputibias.n74 outputibias.n71 104.615
R25414 outputibias.n122 outputibias.n121 104.615
R25415 outputibias.n121 outputibias.n99 104.615
R25416 outputibias.n114 outputibias.n99 104.615
R25417 outputibias.n114 outputibias.n113 104.615
R25418 outputibias.n113 outputibias.n103 104.615
R25419 outputibias.n106 outputibias.n103 104.615
R25420 outputibias.n63 outputibias.n31 95.6354
R25421 outputibias.n63 outputibias.n62 94.6732
R25422 outputibias.n95 outputibias.n94 94.6732
R25423 outputibias.n127 outputibias.n126 94.6732
R25424 outputibias.n11 outputibias.t7 52.3082
R25425 outputibias.n42 outputibias.t1 52.3082
R25426 outputibias.n74 outputibias.t3 52.3082
R25427 outputibias.n106 outputibias.t5 52.3082
R25428 outputibias.n12 outputibias.n10 15.6674
R25429 outputibias.n43 outputibias.n41 15.6674
R25430 outputibias.n75 outputibias.n73 15.6674
R25431 outputibias.n107 outputibias.n105 15.6674
R25432 outputibias.n13 outputibias.n9 12.8005
R25433 outputibias.n44 outputibias.n40 12.8005
R25434 outputibias.n76 outputibias.n72 12.8005
R25435 outputibias.n108 outputibias.n104 12.8005
R25436 outputibias.n17 outputibias.n16 12.0247
R25437 outputibias.n48 outputibias.n47 12.0247
R25438 outputibias.n80 outputibias.n79 12.0247
R25439 outputibias.n112 outputibias.n111 12.0247
R25440 outputibias.n20 outputibias.n7 11.249
R25441 outputibias.n51 outputibias.n38 11.249
R25442 outputibias.n83 outputibias.n70 11.249
R25443 outputibias.n115 outputibias.n102 11.249
R25444 outputibias.n21 outputibias.n5 10.4732
R25445 outputibias.n52 outputibias.n36 10.4732
R25446 outputibias.n84 outputibias.n68 10.4732
R25447 outputibias.n116 outputibias.n100 10.4732
R25448 outputibias.n25 outputibias.n24 9.69747
R25449 outputibias.n56 outputibias.n55 9.69747
R25450 outputibias.n88 outputibias.n87 9.69747
R25451 outputibias.n120 outputibias.n119 9.69747
R25452 outputibias.n31 outputibias.n30 9.45567
R25453 outputibias.n62 outputibias.n61 9.45567
R25454 outputibias.n94 outputibias.n93 9.45567
R25455 outputibias.n126 outputibias.n125 9.45567
R25456 outputibias.n30 outputibias.n29 9.3005
R25457 outputibias.n3 outputibias.n2 9.3005
R25458 outputibias.n24 outputibias.n23 9.3005
R25459 outputibias.n22 outputibias.n21 9.3005
R25460 outputibias.n7 outputibias.n6 9.3005
R25461 outputibias.n16 outputibias.n15 9.3005
R25462 outputibias.n14 outputibias.n13 9.3005
R25463 outputibias.n61 outputibias.n60 9.3005
R25464 outputibias.n34 outputibias.n33 9.3005
R25465 outputibias.n55 outputibias.n54 9.3005
R25466 outputibias.n53 outputibias.n52 9.3005
R25467 outputibias.n38 outputibias.n37 9.3005
R25468 outputibias.n47 outputibias.n46 9.3005
R25469 outputibias.n45 outputibias.n44 9.3005
R25470 outputibias.n93 outputibias.n92 9.3005
R25471 outputibias.n66 outputibias.n65 9.3005
R25472 outputibias.n87 outputibias.n86 9.3005
R25473 outputibias.n85 outputibias.n84 9.3005
R25474 outputibias.n70 outputibias.n69 9.3005
R25475 outputibias.n79 outputibias.n78 9.3005
R25476 outputibias.n77 outputibias.n76 9.3005
R25477 outputibias.n125 outputibias.n124 9.3005
R25478 outputibias.n98 outputibias.n97 9.3005
R25479 outputibias.n119 outputibias.n118 9.3005
R25480 outputibias.n117 outputibias.n116 9.3005
R25481 outputibias.n102 outputibias.n101 9.3005
R25482 outputibias.n111 outputibias.n110 9.3005
R25483 outputibias.n109 outputibias.n108 9.3005
R25484 outputibias.n28 outputibias.n3 8.92171
R25485 outputibias.n59 outputibias.n34 8.92171
R25486 outputibias.n91 outputibias.n66 8.92171
R25487 outputibias.n123 outputibias.n98 8.92171
R25488 outputibias.n29 outputibias.n1 8.14595
R25489 outputibias.n60 outputibias.n32 8.14595
R25490 outputibias.n92 outputibias.n64 8.14595
R25491 outputibias.n124 outputibias.n96 8.14595
R25492 outputibias.n31 outputibias.n1 5.81868
R25493 outputibias.n62 outputibias.n32 5.81868
R25494 outputibias.n94 outputibias.n64 5.81868
R25495 outputibias.n126 outputibias.n96 5.81868
R25496 outputibias.n131 outputibias.n130 5.20947
R25497 outputibias.n29 outputibias.n28 5.04292
R25498 outputibias.n60 outputibias.n59 5.04292
R25499 outputibias.n92 outputibias.n91 5.04292
R25500 outputibias.n124 outputibias.n123 5.04292
R25501 outputibias.n131 outputibias.n127 4.42209
R25502 outputibias.n14 outputibias.n10 4.38594
R25503 outputibias.n45 outputibias.n41 4.38594
R25504 outputibias.n77 outputibias.n73 4.38594
R25505 outputibias.n109 outputibias.n105 4.38594
R25506 outputibias.n132 outputibias.n131 4.28454
R25507 outputibias.n25 outputibias.n3 4.26717
R25508 outputibias.n56 outputibias.n34 4.26717
R25509 outputibias.n88 outputibias.n66 4.26717
R25510 outputibias.n120 outputibias.n98 4.26717
R25511 outputibias.n24 outputibias.n5 3.49141
R25512 outputibias.n55 outputibias.n36 3.49141
R25513 outputibias.n87 outputibias.n68 3.49141
R25514 outputibias.n119 outputibias.n100 3.49141
R25515 outputibias.n21 outputibias.n20 2.71565
R25516 outputibias.n52 outputibias.n51 2.71565
R25517 outputibias.n84 outputibias.n83 2.71565
R25518 outputibias.n116 outputibias.n115 2.71565
R25519 outputibias.n17 outputibias.n7 1.93989
R25520 outputibias.n48 outputibias.n38 1.93989
R25521 outputibias.n80 outputibias.n70 1.93989
R25522 outputibias.n112 outputibias.n102 1.93989
R25523 outputibias.n130 outputibias.n129 1.9266
R25524 outputibias.n129 outputibias.n128 1.9266
R25525 outputibias.n133 outputibias.n132 1.92658
R25526 outputibias.n134 outputibias.n133 1.29913
R25527 outputibias.n16 outputibias.n9 1.16414
R25528 outputibias.n47 outputibias.n40 1.16414
R25529 outputibias.n79 outputibias.n72 1.16414
R25530 outputibias.n111 outputibias.n104 1.16414
R25531 outputibias.n127 outputibias.n95 0.962709
R25532 outputibias.n95 outputibias.n63 0.962709
R25533 outputibias.n13 outputibias.n12 0.388379
R25534 outputibias.n44 outputibias.n43 0.388379
R25535 outputibias.n76 outputibias.n75 0.388379
R25536 outputibias.n108 outputibias.n107 0.388379
R25537 outputibias.n134 outputibias.n0 0.337251
R25538 outputibias outputibias.n134 0.302375
R25539 outputibias.n30 outputibias.n2 0.155672
R25540 outputibias.n23 outputibias.n2 0.155672
R25541 outputibias.n23 outputibias.n22 0.155672
R25542 outputibias.n22 outputibias.n6 0.155672
R25543 outputibias.n15 outputibias.n6 0.155672
R25544 outputibias.n15 outputibias.n14 0.155672
R25545 outputibias.n61 outputibias.n33 0.155672
R25546 outputibias.n54 outputibias.n33 0.155672
R25547 outputibias.n54 outputibias.n53 0.155672
R25548 outputibias.n53 outputibias.n37 0.155672
R25549 outputibias.n46 outputibias.n37 0.155672
R25550 outputibias.n46 outputibias.n45 0.155672
R25551 outputibias.n93 outputibias.n65 0.155672
R25552 outputibias.n86 outputibias.n65 0.155672
R25553 outputibias.n86 outputibias.n85 0.155672
R25554 outputibias.n85 outputibias.n69 0.155672
R25555 outputibias.n78 outputibias.n69 0.155672
R25556 outputibias.n78 outputibias.n77 0.155672
R25557 outputibias.n125 outputibias.n97 0.155672
R25558 outputibias.n118 outputibias.n97 0.155672
R25559 outputibias.n118 outputibias.n117 0.155672
R25560 outputibias.n117 outputibias.n101 0.155672
R25561 outputibias.n110 outputibias.n101 0.155672
R25562 outputibias.n110 outputibias.n109 0.155672
C0 commonsourceibias outputibias 0.003832f
C1 plus diffpairibias 4.13e-19
C2 vdd commonsourceibias 0.004218f
C3 CSoutput plus 0.895742f
C4 commonsourceibias diffpairibias 0.06482f
C5 CSoutput commonsourceibias 66.33679f
C6 minus plus 9.99291f
C7 minus commonsourceibias 0.462932f
C8 plus commonsourceibias 0.417773f
C9 output outputibias 2.34152f
C10 vdd output 7.23429f
C11 CSoutput output 6.13881f
C12 CSoutput outputibias 0.032386f
C13 vdd CSoutput 0.117233p
C14 minus diffpairibias 5.12e-19
C15 commonsourceibias output 0.006808f
C16 CSoutput minus 2.92497f
C17 vdd plus 0.095754f
C18 diffpairibias gnd 48.98024f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.22223p
C22 plus gnd 36.411797f
C23 minus gnd 29.63035f
C24 CSoutput gnd 0.143055p
C25 vdd gnd 0.511372p
C26 outputibias.t10 gnd 0.11477f
C27 outputibias.t8 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t7 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t1 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t3 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t5 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t4 gnd 0.108319f
C161 outputibias.t2 gnd 0.108319f
C162 outputibias.t0 gnd 0.108319f
C163 outputibias.t6 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t9 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t11 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 diffpairibias.t18 gnd 0.087401f
C174 diffpairibias.t22 gnd 0.087239f
C175 diffpairibias.n0 gnd 0.102784f
C176 diffpairibias.t20 gnd 0.087239f
C177 diffpairibias.n1 gnd 0.050171f
C178 diffpairibias.t23 gnd 0.087239f
C179 diffpairibias.n2 gnd 0.039841f
C180 diffpairibias.t1 gnd 0.083757f
C181 diffpairibias.t9 gnd 0.083392f
C182 diffpairibias.n3 gnd 0.131682f
C183 diffpairibias.t11 gnd 0.083392f
C184 diffpairibias.n4 gnd 0.07027f
C185 diffpairibias.t7 gnd 0.083392f
C186 diffpairibias.n5 gnd 0.07027f
C187 diffpairibias.t3 gnd 0.083392f
C188 diffpairibias.n6 gnd 0.07027f
C189 diffpairibias.t13 gnd 0.083392f
C190 diffpairibias.n7 gnd 0.07027f
C191 diffpairibias.t5 gnd 0.083392f
C192 diffpairibias.n8 gnd 0.07027f
C193 diffpairibias.t15 gnd 0.083392f
C194 diffpairibias.n9 gnd 0.099771f
C195 diffpairibias.t0 gnd 0.08427f
C196 diffpairibias.t8 gnd 0.084123f
C197 diffpairibias.n10 gnd 0.091784f
C198 diffpairibias.t10 gnd 0.084123f
C199 diffpairibias.n11 gnd 0.050681f
C200 diffpairibias.t6 gnd 0.084123f
C201 diffpairibias.n12 gnd 0.050681f
C202 diffpairibias.t2 gnd 0.084123f
C203 diffpairibias.n13 gnd 0.050681f
C204 diffpairibias.t12 gnd 0.084123f
C205 diffpairibias.n14 gnd 0.050681f
C206 diffpairibias.t4 gnd 0.084123f
C207 diffpairibias.n15 gnd 0.050681f
C208 diffpairibias.t14 gnd 0.084123f
C209 diffpairibias.n16 gnd 0.059977f
C210 diffpairibias.n17 gnd 0.226448f
C211 diffpairibias.t21 gnd 0.087239f
C212 diffpairibias.n18 gnd 0.050181f
C213 diffpairibias.t17 gnd 0.087239f
C214 diffpairibias.n19 gnd 0.050171f
C215 diffpairibias.t16 gnd 0.087239f
C216 diffpairibias.n20 gnd 0.050171f
C217 diffpairibias.t19 gnd 0.087239f
C218 diffpairibias.n21 gnd 0.045859f
C219 diffpairibias.n22 gnd 0.046268f
C220 minus.n0 gnd 0.030055f
C221 minus.t13 gnd 0.505366f
C222 minus.n1 gnd 0.204393f
C223 minus.n2 gnd 0.030055f
C224 minus.t20 gnd 0.505366f
C225 minus.n3 gnd 0.024893f
C226 minus.n4 gnd 0.030055f
C227 minus.t17 gnd 0.505366f
C228 minus.t23 gnd 0.505366f
C229 minus.n5 gnd 0.204393f
C230 minus.n6 gnd 0.030055f
C231 minus.t22 gnd 0.505366f
C232 minus.n7 gnd 0.204393f
C233 minus.n8 gnd 0.030055f
C234 minus.t5 gnd 0.505366f
C235 minus.n9 gnd 0.024893f
C236 minus.n10 gnd 0.030055f
C237 minus.t8 gnd 0.505366f
C238 minus.t10 gnd 0.505366f
C239 minus.n11 gnd 0.235043f
C240 minus.t16 gnd 0.566382f
C241 minus.n12 gnd 0.238051f
C242 minus.n13 gnd 0.128281f
C243 minus.n14 gnd 0.037948f
C244 minus.n15 gnd 0.034573f
C245 minus.n16 gnd 0.204393f
C246 minus.n17 gnd 0.036886f
C247 minus.n18 gnd 0.030055f
C248 minus.n19 gnd 0.030055f
C249 minus.n20 gnd 0.030055f
C250 minus.n21 gnd 0.038962f
C251 minus.n22 gnd 0.204393f
C252 minus.n23 gnd 0.036823f
C253 minus.n24 gnd 0.035698f
C254 minus.n25 gnd 0.030055f
C255 minus.n26 gnd 0.030055f
C256 minus.n27 gnd 0.038233f
C257 minus.n28 gnd 0.024274f
C258 minus.n29 gnd 0.038233f
C259 minus.n30 gnd 0.030055f
C260 minus.n31 gnd 0.030055f
C261 minus.n32 gnd 0.035698f
C262 minus.n33 gnd 0.036823f
C263 minus.n34 gnd 0.204393f
C264 minus.n35 gnd 0.038962f
C265 minus.n36 gnd 0.030055f
C266 minus.n37 gnd 0.030055f
C267 minus.n38 gnd 0.030055f
C268 minus.n39 gnd 0.036886f
C269 minus.n40 gnd 0.204393f
C270 minus.n41 gnd 0.034573f
C271 minus.n42 gnd 0.037948f
C272 minus.n43 gnd 0.030055f
C273 minus.n44 gnd 0.030055f
C274 minus.n45 gnd 0.03922f
C275 minus.n46 gnd 0.01164f
C276 minus.t9 gnd 0.546554f
C277 minus.n47 gnd 0.237023f
C278 minus.n48 gnd 0.352615f
C279 minus.n49 gnd 0.030055f
C280 minus.t14 gnd 0.546554f
C281 minus.t21 gnd 0.505366f
C282 minus.n50 gnd 0.204393f
C283 minus.n51 gnd 0.030055f
C284 minus.t18 gnd 0.505366f
C285 minus.n52 gnd 0.024893f
C286 minus.n53 gnd 0.030055f
C287 minus.t15 gnd 0.505366f
C288 minus.t7 gnd 0.505366f
C289 minus.n54 gnd 0.204393f
C290 minus.n55 gnd 0.030055f
C291 minus.t6 gnd 0.505366f
C292 minus.n56 gnd 0.204393f
C293 minus.n57 gnd 0.030055f
C294 minus.t12 gnd 0.505366f
C295 minus.n58 gnd 0.024893f
C296 minus.n59 gnd 0.030055f
C297 minus.t11 gnd 0.505366f
C298 minus.t19 gnd 0.505366f
C299 minus.n60 gnd 0.235043f
C300 minus.t24 gnd 0.566382f
C301 minus.n61 gnd 0.238051f
C302 minus.n62 gnd 0.128281f
C303 minus.n63 gnd 0.037948f
C304 minus.n64 gnd 0.034573f
C305 minus.n65 gnd 0.204393f
C306 minus.n66 gnd 0.036886f
C307 minus.n67 gnd 0.030055f
C308 minus.n68 gnd 0.030055f
C309 minus.n69 gnd 0.030055f
C310 minus.n70 gnd 0.038962f
C311 minus.n71 gnd 0.204393f
C312 minus.n72 gnd 0.036823f
C313 minus.n73 gnd 0.035698f
C314 minus.n74 gnd 0.030055f
C315 minus.n75 gnd 0.030055f
C316 minus.n76 gnd 0.038233f
C317 minus.n77 gnd 0.024274f
C318 minus.n78 gnd 0.038233f
C319 minus.n79 gnd 0.030055f
C320 minus.n80 gnd 0.030055f
C321 minus.n81 gnd 0.035698f
C322 minus.n82 gnd 0.036823f
C323 minus.n83 gnd 0.204393f
C324 minus.n84 gnd 0.038962f
C325 minus.n85 gnd 0.030055f
C326 minus.n86 gnd 0.030055f
C327 minus.n87 gnd 0.030055f
C328 minus.n88 gnd 0.036886f
C329 minus.n89 gnd 0.204393f
C330 minus.n90 gnd 0.034573f
C331 minus.n91 gnd 0.037948f
C332 minus.n92 gnd 0.030055f
C333 minus.n93 gnd 0.030055f
C334 minus.n94 gnd 0.03922f
C335 minus.n95 gnd 0.01164f
C336 minus.n96 gnd 0.237023f
C337 minus.n97 gnd 1.01584f
C338 minus.n98 gnd 1.50967f
C339 minus.t2 gnd 0.009265f
C340 minus.t1 gnd 0.009265f
C341 minus.n99 gnd 0.030465f
C342 minus.t3 gnd 0.009265f
C343 minus.t0 gnd 0.009265f
C344 minus.n100 gnd 0.030048f
C345 minus.n101 gnd 0.256447f
C346 minus.t4 gnd 0.051568f
C347 minus.n102 gnd 0.139941f
C348 minus.n103 gnd 2.01704f
C349 output.t0 gnd 0.464308f
C350 output.t10 gnd 0.044422f
C351 output.t8 gnd 0.044422f
C352 output.n0 gnd 0.364624f
C353 output.n1 gnd 0.614102f
C354 output.t15 gnd 0.044422f
C355 output.t2 gnd 0.044422f
C356 output.n2 gnd 0.364624f
C357 output.n3 gnd 0.350265f
C358 output.t4 gnd 0.044422f
C359 output.t12 gnd 0.044422f
C360 output.n4 gnd 0.364624f
C361 output.n5 gnd 0.350265f
C362 output.t14 gnd 0.044422f
C363 output.t5 gnd 0.044422f
C364 output.n6 gnd 0.364624f
C365 output.n7 gnd 0.350265f
C366 output.t6 gnd 0.044422f
C367 output.t11 gnd 0.044422f
C368 output.n8 gnd 0.364624f
C369 output.n9 gnd 0.350265f
C370 output.t13 gnd 0.044422f
C371 output.t3 gnd 0.044422f
C372 output.n10 gnd 0.364624f
C373 output.n11 gnd 0.350265f
C374 output.t9 gnd 0.044422f
C375 output.t7 gnd 0.044422f
C376 output.n12 gnd 0.364624f
C377 output.n13 gnd 0.350265f
C378 output.t1 gnd 0.462979f
C379 output.n14 gnd 0.28994f
C380 output.n15 gnd 0.015803f
C381 output.n16 gnd 0.011243f
C382 output.n17 gnd 0.006041f
C383 output.n18 gnd 0.01428f
C384 output.n19 gnd 0.006397f
C385 output.n20 gnd 0.011243f
C386 output.n21 gnd 0.006041f
C387 output.n22 gnd 0.01428f
C388 output.n23 gnd 0.006397f
C389 output.n24 gnd 0.048111f
C390 output.t18 gnd 0.023274f
C391 output.n25 gnd 0.01071f
C392 output.n26 gnd 0.008435f
C393 output.n27 gnd 0.006041f
C394 output.n28 gnd 0.267512f
C395 output.n29 gnd 0.011243f
C396 output.n30 gnd 0.006041f
C397 output.n31 gnd 0.006397f
C398 output.n32 gnd 0.01428f
C399 output.n33 gnd 0.01428f
C400 output.n34 gnd 0.006397f
C401 output.n35 gnd 0.006041f
C402 output.n36 gnd 0.011243f
C403 output.n37 gnd 0.011243f
C404 output.n38 gnd 0.006041f
C405 output.n39 gnd 0.006397f
C406 output.n40 gnd 0.01428f
C407 output.n41 gnd 0.030913f
C408 output.n42 gnd 0.006397f
C409 output.n43 gnd 0.006041f
C410 output.n44 gnd 0.025987f
C411 output.n45 gnd 0.097665f
C412 output.n46 gnd 0.015803f
C413 output.n47 gnd 0.011243f
C414 output.n48 gnd 0.006041f
C415 output.n49 gnd 0.01428f
C416 output.n50 gnd 0.006397f
C417 output.n51 gnd 0.011243f
C418 output.n52 gnd 0.006041f
C419 output.n53 gnd 0.01428f
C420 output.n54 gnd 0.006397f
C421 output.n55 gnd 0.048111f
C422 output.t17 gnd 0.023274f
C423 output.n56 gnd 0.01071f
C424 output.n57 gnd 0.008435f
C425 output.n58 gnd 0.006041f
C426 output.n59 gnd 0.267512f
C427 output.n60 gnd 0.011243f
C428 output.n61 gnd 0.006041f
C429 output.n62 gnd 0.006397f
C430 output.n63 gnd 0.01428f
C431 output.n64 gnd 0.01428f
C432 output.n65 gnd 0.006397f
C433 output.n66 gnd 0.006041f
C434 output.n67 gnd 0.011243f
C435 output.n68 gnd 0.011243f
C436 output.n69 gnd 0.006041f
C437 output.n70 gnd 0.006397f
C438 output.n71 gnd 0.01428f
C439 output.n72 gnd 0.030913f
C440 output.n73 gnd 0.006397f
C441 output.n74 gnd 0.006041f
C442 output.n75 gnd 0.025987f
C443 output.n76 gnd 0.09306f
C444 output.n77 gnd 1.65264f
C445 output.n78 gnd 0.015803f
C446 output.n79 gnd 0.011243f
C447 output.n80 gnd 0.006041f
C448 output.n81 gnd 0.01428f
C449 output.n82 gnd 0.006397f
C450 output.n83 gnd 0.011243f
C451 output.n84 gnd 0.006041f
C452 output.n85 gnd 0.01428f
C453 output.n86 gnd 0.006397f
C454 output.n87 gnd 0.048111f
C455 output.t16 gnd 0.023274f
C456 output.n88 gnd 0.01071f
C457 output.n89 gnd 0.008435f
C458 output.n90 gnd 0.006041f
C459 output.n91 gnd 0.267512f
C460 output.n92 gnd 0.011243f
C461 output.n93 gnd 0.006041f
C462 output.n94 gnd 0.006397f
C463 output.n95 gnd 0.01428f
C464 output.n96 gnd 0.01428f
C465 output.n97 gnd 0.006397f
C466 output.n98 gnd 0.006041f
C467 output.n99 gnd 0.011243f
C468 output.n100 gnd 0.011243f
C469 output.n101 gnd 0.006041f
C470 output.n102 gnd 0.006397f
C471 output.n103 gnd 0.01428f
C472 output.n104 gnd 0.030913f
C473 output.n105 gnd 0.006397f
C474 output.n106 gnd 0.006041f
C475 output.n107 gnd 0.025987f
C476 output.n108 gnd 0.09306f
C477 output.n109 gnd 0.713089f
C478 output.n110 gnd 0.015803f
C479 output.n111 gnd 0.011243f
C480 output.n112 gnd 0.006041f
C481 output.n113 gnd 0.01428f
C482 output.n114 gnd 0.006397f
C483 output.n115 gnd 0.011243f
C484 output.n116 gnd 0.006041f
C485 output.n117 gnd 0.01428f
C486 output.n118 gnd 0.006397f
C487 output.n119 gnd 0.048111f
C488 output.t19 gnd 0.023274f
C489 output.n120 gnd 0.01071f
C490 output.n121 gnd 0.008435f
C491 output.n122 gnd 0.006041f
C492 output.n123 gnd 0.267512f
C493 output.n124 gnd 0.011243f
C494 output.n125 gnd 0.006041f
C495 output.n126 gnd 0.006397f
C496 output.n127 gnd 0.01428f
C497 output.n128 gnd 0.01428f
C498 output.n129 gnd 0.006397f
C499 output.n130 gnd 0.006041f
C500 output.n131 gnd 0.011243f
C501 output.n132 gnd 0.011243f
C502 output.n133 gnd 0.006041f
C503 output.n134 gnd 0.006397f
C504 output.n135 gnd 0.01428f
C505 output.n136 gnd 0.030913f
C506 output.n137 gnd 0.006397f
C507 output.n138 gnd 0.006041f
C508 output.n139 gnd 0.025987f
C509 output.n140 gnd 0.09306f
C510 output.n141 gnd 1.67353f
C511 a_n2982_8322.t13 gnd 0.100149f
C512 a_n2982_8322.t1 gnd 20.7769f
C513 a_n2982_8322.t2 gnd 20.631199f
C514 a_n2982_8322.t4 gnd 20.631199f
C515 a_n2982_8322.t0 gnd 20.7769f
C516 a_n2982_8322.t3 gnd 20.631199f
C517 a_n2982_8322.t5 gnd 29.5576f
C518 a_n2982_8322.t12 gnd 0.937748f
C519 a_n2982_8322.t25 gnd 0.100149f
C520 a_n2982_8322.t21 gnd 0.100149f
C521 a_n2982_8322.n0 gnd 0.705452f
C522 a_n2982_8322.n1 gnd 0.788239f
C523 a_n2982_8322.t28 gnd 0.100149f
C524 a_n2982_8322.t18 gnd 0.100149f
C525 a_n2982_8322.n2 gnd 0.705452f
C526 a_n2982_8322.n3 gnd 0.400494f
C527 a_n2982_8322.t9 gnd 0.100149f
C528 a_n2982_8322.t8 gnd 0.100149f
C529 a_n2982_8322.n4 gnd 0.705452f
C530 a_n2982_8322.n5 gnd 0.400494f
C531 a_n2982_8322.t22 gnd 0.100149f
C532 a_n2982_8322.t15 gnd 0.100149f
C533 a_n2982_8322.n6 gnd 0.705452f
C534 a_n2982_8322.n7 gnd 0.400494f
C535 a_n2982_8322.t19 gnd 0.100149f
C536 a_n2982_8322.t17 gnd 0.100149f
C537 a_n2982_8322.n8 gnd 0.705452f
C538 a_n2982_8322.n9 gnd 0.400494f
C539 a_n2982_8322.t6 gnd 0.935881f
C540 a_n2982_8322.n10 gnd 1.8712f
C541 a_n2982_8322.t33 gnd 0.937748f
C542 a_n2982_8322.t37 gnd 0.100149f
C543 a_n2982_8322.t36 gnd 0.100149f
C544 a_n2982_8322.n11 gnd 0.705452f
C545 a_n2982_8322.n12 gnd 0.788239f
C546 a_n2982_8322.t31 gnd 0.935881f
C547 a_n2982_8322.n13 gnd 0.396653f
C548 a_n2982_8322.t34 gnd 0.935881f
C549 a_n2982_8322.n14 gnd 0.396653f
C550 a_n2982_8322.t32 gnd 0.100149f
C551 a_n2982_8322.t30 gnd 0.100149f
C552 a_n2982_8322.n15 gnd 0.705452f
C553 a_n2982_8322.n16 gnd 0.400494f
C554 a_n2982_8322.t35 gnd 0.935881f
C555 a_n2982_8322.n17 gnd 1.47125f
C556 a_n2982_8322.n18 gnd 2.3511f
C557 a_n2982_8322.n19 gnd 3.56583f
C558 a_n2982_8322.t7 gnd 0.935881f
C559 a_n2982_8322.n20 gnd 1.11135f
C560 a_n2982_8322.t24 gnd 0.100149f
C561 a_n2982_8322.t23 gnd 0.100149f
C562 a_n2982_8322.n21 gnd 0.705452f
C563 a_n2982_8322.n22 gnd 0.400494f
C564 a_n2982_8322.t11 gnd 0.100149f
C565 a_n2982_8322.t10 gnd 0.100149f
C566 a_n2982_8322.n23 gnd 0.705452f
C567 a_n2982_8322.n24 gnd 0.400494f
C568 a_n2982_8322.t26 gnd 0.100149f
C569 a_n2982_8322.t14 gnd 0.100149f
C570 a_n2982_8322.n25 gnd 0.705452f
C571 a_n2982_8322.n26 gnd 0.400494f
C572 a_n2982_8322.t27 gnd 0.937745f
C573 a_n2982_8322.t20 gnd 0.100149f
C574 a_n2982_8322.t16 gnd 0.100149f
C575 a_n2982_8322.n27 gnd 0.705452f
C576 a_n2982_8322.n28 gnd 0.788241f
C577 a_n2982_8322.n29 gnd 0.400492f
C578 a_n2982_8322.n30 gnd 0.705454f
C579 a_n2982_8322.t29 gnd 0.100149f
C580 a_n2903_n3924.t4 gnd 0.094851f
C581 a_n2903_n3924.t14 gnd 0.985803f
C582 a_n2903_n3924.n0 gnd 0.372677f
C583 a_n2903_n3924.t23 gnd 1.22484f
C584 a_n2903_n3924.n1 gnd 1.15477f
C585 a_n2903_n3924.t39 gnd 0.985803f
C586 a_n2903_n3924.n2 gnd 0.372677f
C587 a_n2903_n3924.t30 gnd 0.094851f
C588 a_n2903_n3924.t44 gnd 0.094851f
C589 a_n2903_n3924.n3 gnd 0.774663f
C590 a_n2903_n3924.n4 gnd 0.390386f
C591 a_n2903_n3924.t25 gnd 0.094851f
C592 a_n2903_n3924.t31 gnd 0.094851f
C593 a_n2903_n3924.n5 gnd 0.774663f
C594 a_n2903_n3924.n6 gnd 0.390386f
C595 a_n2903_n3924.t40 gnd 0.094851f
C596 a_n2903_n3924.t28 gnd 0.094851f
C597 a_n2903_n3924.n7 gnd 0.774663f
C598 a_n2903_n3924.n8 gnd 0.390386f
C599 a_n2903_n3924.t47 gnd 0.094851f
C600 a_n2903_n3924.t32 gnd 0.094851f
C601 a_n2903_n3924.n9 gnd 0.774663f
C602 a_n2903_n3924.n10 gnd 0.390386f
C603 a_n2903_n3924.t21 gnd 0.985803f
C604 a_n2903_n3924.n11 gnd 0.922787f
C605 a_n2903_n3924.t34 gnd 1.22537f
C606 a_n2903_n3924.t43 gnd 1.22484f
C607 a_n2903_n3924.n12 gnd 0.862674f
C608 a_n2903_n3924.t46 gnd 1.22484f
C609 a_n2903_n3924.n13 gnd 0.862674f
C610 a_n2903_n3924.t29 gnd 1.22484f
C611 a_n2903_n3924.n14 gnd 0.862674f
C612 a_n2903_n3924.t37 gnd 1.22484f
C613 a_n2903_n3924.n15 gnd 0.862674f
C614 a_n2903_n3924.t35 gnd 1.22484f
C615 a_n2903_n3924.n16 gnd 0.862674f
C616 a_n2903_n3924.t26 gnd 1.22484f
C617 a_n2903_n3924.n17 gnd 0.716127f
C618 a_n2903_n3924.n18 gnd 0.845678f
C619 a_n2903_n3924.n19 gnd 0.894202f
C620 a_n2903_n3924.t19 gnd 0.985799f
C621 a_n2903_n3924.n20 gnd 0.612329f
C622 a_n2903_n3924.t13 gnd 0.094851f
C623 a_n2903_n3924.t17 gnd 0.094851f
C624 a_n2903_n3924.n21 gnd 0.774662f
C625 a_n2903_n3924.n22 gnd 0.390388f
C626 a_n2903_n3924.t18 gnd 0.094851f
C627 a_n2903_n3924.t6 gnd 0.094851f
C628 a_n2903_n3924.n23 gnd 0.774662f
C629 a_n2903_n3924.n24 gnd 0.390388f
C630 a_n2903_n3924.t7 gnd 0.094851f
C631 a_n2903_n3924.t1 gnd 0.094851f
C632 a_n2903_n3924.n25 gnd 0.774662f
C633 a_n2903_n3924.n26 gnd 0.390388f
C634 a_n2903_n3924.t3 gnd 0.094851f
C635 a_n2903_n3924.t16 gnd 0.094851f
C636 a_n2903_n3924.n27 gnd 0.774662f
C637 a_n2903_n3924.n28 gnd 0.390388f
C638 a_n2903_n3924.t11 gnd 0.985799f
C639 a_n2903_n3924.n29 gnd 0.372681f
C640 a_n2903_n3924.t24 gnd 0.985799f
C641 a_n2903_n3924.n30 gnd 0.372681f
C642 a_n2903_n3924.t45 gnd 0.094851f
C643 a_n2903_n3924.t0 gnd 0.094851f
C644 a_n2903_n3924.n31 gnd 0.774662f
C645 a_n2903_n3924.n32 gnd 0.390388f
C646 a_n2903_n3924.t42 gnd 0.094851f
C647 a_n2903_n3924.t22 gnd 0.094851f
C648 a_n2903_n3924.n33 gnd 0.774662f
C649 a_n2903_n3924.n34 gnd 0.390388f
C650 a_n2903_n3924.t27 gnd 0.094851f
C651 a_n2903_n3924.t41 gnd 0.094851f
C652 a_n2903_n3924.n35 gnd 0.774662f
C653 a_n2903_n3924.n36 gnd 0.390388f
C654 a_n2903_n3924.t38 gnd 0.094851f
C655 a_n2903_n3924.t33 gnd 0.094851f
C656 a_n2903_n3924.n37 gnd 0.774662f
C657 a_n2903_n3924.n38 gnd 0.390388f
C658 a_n2903_n3924.t36 gnd 0.985799f
C659 a_n2903_n3924.n39 gnd 0.612329f
C660 a_n2903_n3924.n40 gnd 0.953249f
C661 a_n2903_n3924.t2 gnd 0.985799f
C662 a_n2903_n3924.n41 gnd 0.922791f
C663 a_n2903_n3924.t10 gnd 0.094851f
C664 a_n2903_n3924.t15 gnd 0.094851f
C665 a_n2903_n3924.n42 gnd 0.774663f
C666 a_n2903_n3924.n43 gnd 0.390386f
C667 a_n2903_n3924.t8 gnd 0.094851f
C668 a_n2903_n3924.t12 gnd 0.094851f
C669 a_n2903_n3924.n44 gnd 0.774663f
C670 a_n2903_n3924.n45 gnd 0.390386f
C671 a_n2903_n3924.t5 gnd 0.094851f
C672 a_n2903_n3924.t9 gnd 0.094851f
C673 a_n2903_n3924.n46 gnd 0.774663f
C674 a_n2903_n3924.n47 gnd 0.390386f
C675 a_n2903_n3924.n48 gnd 0.390385f
C676 a_n2903_n3924.n49 gnd 0.774665f
C677 a_n2903_n3924.t20 gnd 0.094851f
C678 plus.n0 gnd 0.022304f
C679 plus.t6 gnd 0.405612f
C680 plus.t12 gnd 0.375046f
C681 plus.n1 gnd 0.151685f
C682 plus.n2 gnd 0.022304f
C683 plus.t8 gnd 0.375046f
C684 plus.n3 gnd 0.018474f
C685 plus.n4 gnd 0.022304f
C686 plus.t7 gnd 0.375046f
C687 plus.t19 gnd 0.375046f
C688 plus.n5 gnd 0.151685f
C689 plus.n6 gnd 0.022304f
C690 plus.t18 gnd 0.375046f
C691 plus.n7 gnd 0.151685f
C692 plus.n8 gnd 0.022304f
C693 plus.t24 gnd 0.375046f
C694 plus.n9 gnd 0.018474f
C695 plus.n10 gnd 0.022304f
C696 plus.t22 gnd 0.375046f
C697 plus.t9 gnd 0.375046f
C698 plus.n11 gnd 0.174432f
C699 plus.t14 gnd 0.420328f
C700 plus.n12 gnd 0.176664f
C701 plus.n13 gnd 0.095201f
C702 plus.n14 gnd 0.028162f
C703 plus.n15 gnd 0.025657f
C704 plus.n16 gnd 0.151685f
C705 plus.n17 gnd 0.027374f
C706 plus.n18 gnd 0.022304f
C707 plus.n19 gnd 0.022304f
C708 plus.n20 gnd 0.022304f
C709 plus.n21 gnd 0.028914f
C710 plus.n22 gnd 0.151685f
C711 plus.n23 gnd 0.027327f
C712 plus.n24 gnd 0.026492f
C713 plus.n25 gnd 0.022304f
C714 plus.n26 gnd 0.022304f
C715 plus.n27 gnd 0.028374f
C716 plus.n28 gnd 0.018015f
C717 plus.n29 gnd 0.028374f
C718 plus.n30 gnd 0.022304f
C719 plus.n31 gnd 0.022304f
C720 plus.n32 gnd 0.026492f
C721 plus.n33 gnd 0.027327f
C722 plus.n34 gnd 0.151685f
C723 plus.n35 gnd 0.028914f
C724 plus.n36 gnd 0.022304f
C725 plus.n37 gnd 0.022304f
C726 plus.n38 gnd 0.022304f
C727 plus.n39 gnd 0.027374f
C728 plus.n40 gnd 0.151685f
C729 plus.n41 gnd 0.025657f
C730 plus.n42 gnd 0.028162f
C731 plus.n43 gnd 0.022304f
C732 plus.n44 gnd 0.022304f
C733 plus.n45 gnd 0.029106f
C734 plus.n46 gnd 0.008638f
C735 plus.n47 gnd 0.175901f
C736 plus.n48 gnd 0.255948f
C737 plus.n49 gnd 0.022304f
C738 plus.t10 gnd 0.375046f
C739 plus.n50 gnd 0.151685f
C740 plus.n51 gnd 0.022304f
C741 plus.t15 gnd 0.375046f
C742 plus.n52 gnd 0.018474f
C743 plus.n53 gnd 0.022304f
C744 plus.t13 gnd 0.375046f
C745 plus.t17 gnd 0.375046f
C746 plus.n54 gnd 0.151685f
C747 plus.n55 gnd 0.022304f
C748 plus.t16 gnd 0.375046f
C749 plus.n56 gnd 0.151685f
C750 plus.n57 gnd 0.022304f
C751 plus.t20 gnd 0.375046f
C752 plus.n58 gnd 0.018474f
C753 plus.n59 gnd 0.022304f
C754 plus.t21 gnd 0.375046f
C755 plus.t5 gnd 0.375046f
C756 plus.n60 gnd 0.174432f
C757 plus.t11 gnd 0.420328f
C758 plus.n61 gnd 0.176664f
C759 plus.n62 gnd 0.095201f
C760 plus.n63 gnd 0.028162f
C761 plus.n64 gnd 0.025657f
C762 plus.n65 gnd 0.151685f
C763 plus.n66 gnd 0.027374f
C764 plus.n67 gnd 0.022304f
C765 plus.n68 gnd 0.022304f
C766 plus.n69 gnd 0.022304f
C767 plus.n70 gnd 0.028914f
C768 plus.n71 gnd 0.151685f
C769 plus.n72 gnd 0.027327f
C770 plus.n73 gnd 0.026492f
C771 plus.n74 gnd 0.022304f
C772 plus.n75 gnd 0.022304f
C773 plus.n76 gnd 0.028374f
C774 plus.n77 gnd 0.018015f
C775 plus.n78 gnd 0.028374f
C776 plus.n79 gnd 0.022304f
C777 plus.n80 gnd 0.022304f
C778 plus.n81 gnd 0.026492f
C779 plus.n82 gnd 0.027327f
C780 plus.n83 gnd 0.151685f
C781 plus.n84 gnd 0.028914f
C782 plus.n85 gnd 0.022304f
C783 plus.n86 gnd 0.022304f
C784 plus.n87 gnd 0.022304f
C785 plus.n88 gnd 0.027374f
C786 plus.n89 gnd 0.151685f
C787 plus.n90 gnd 0.025657f
C788 plus.n91 gnd 0.028162f
C789 plus.n92 gnd 0.022304f
C790 plus.n93 gnd 0.022304f
C791 plus.n94 gnd 0.029106f
C792 plus.n95 gnd 0.008638f
C793 plus.t23 gnd 0.405612f
C794 plus.n96 gnd 0.175901f
C795 plus.n97 gnd 0.744951f
C796 plus.n98 gnd 1.11152f
C797 plus.t1 gnd 0.038504f
C798 plus.t2 gnd 0.006876f
C799 plus.t4 gnd 0.006876f
C800 plus.n99 gnd 0.022299f
C801 plus.n100 gnd 0.173113f
C802 plus.t0 gnd 0.006876f
C803 plus.t3 gnd 0.006876f
C804 plus.n101 gnd 0.022299f
C805 plus.n102 gnd 0.129942f
C806 plus.n103 gnd 2.84863f
C807 a_n8964_8799.n0 gnd 0.88507f
C808 a_n8964_8799.n1 gnd 3.63716f
C809 a_n8964_8799.n2 gnd 3.37643f
C810 a_n8964_8799.n3 gnd 1.67796f
C811 a_n8964_8799.n4 gnd 0.209378f
C812 a_n8964_8799.n5 gnd 0.292646f
C813 a_n8964_8799.n6 gnd 0.209378f
C814 a_n8964_8799.n7 gnd 0.209378f
C815 a_n8964_8799.n8 gnd 0.209378f
C816 a_n8964_8799.n9 gnd 0.275847f
C817 a_n8964_8799.n10 gnd 0.209378f
C818 a_n8964_8799.n11 gnd 0.292646f
C819 a_n8964_8799.n12 gnd 0.209378f
C820 a_n8964_8799.n13 gnd 0.209378f
C821 a_n8964_8799.n14 gnd 0.209378f
C822 a_n8964_8799.n15 gnd 0.275847f
C823 a_n8964_8799.n16 gnd 0.209378f
C824 a_n8964_8799.n17 gnd 0.458634f
C825 a_n8964_8799.n18 gnd 0.209378f
C826 a_n8964_8799.n19 gnd 0.209378f
C827 a_n8964_8799.n20 gnd 0.209378f
C828 a_n8964_8799.n21 gnd 0.275847f
C829 a_n8964_8799.n22 gnd 0.328191f
C830 a_n8964_8799.n23 gnd 0.209378f
C831 a_n8964_8799.n24 gnd 0.209378f
C832 a_n8964_8799.n25 gnd 0.209378f
C833 a_n8964_8799.n26 gnd 0.209378f
C834 a_n8964_8799.n27 gnd 0.240302f
C835 a_n8964_8799.n28 gnd 0.328191f
C836 a_n8964_8799.n29 gnd 0.209378f
C837 a_n8964_8799.n30 gnd 0.209378f
C838 a_n8964_8799.n31 gnd 0.209378f
C839 a_n8964_8799.n32 gnd 0.209378f
C840 a_n8964_8799.n33 gnd 0.240302f
C841 a_n8964_8799.n34 gnd 0.328191f
C842 a_n8964_8799.n35 gnd 0.209378f
C843 a_n8964_8799.n36 gnd 0.209378f
C844 a_n8964_8799.n37 gnd 0.209378f
C845 a_n8964_8799.n38 gnd 0.209378f
C846 a_n8964_8799.n39 gnd 0.406289f
C847 a_n8964_8799.n40 gnd 1.0279f
C848 a_n8964_8799.n41 gnd 1.01334f
C849 a_n8964_8799.n42 gnd 3.00818f
C850 a_n8964_8799.n43 gnd 1.53458f
C851 a_n8964_8799.n44 gnd 3.73985f
C852 a_n8964_8799.n45 gnd 1.01334f
C853 a_n8964_8799.n46 gnd 0.008684f
C854 a_n8964_8799.n47 gnd 0.001166f
C855 a_n8964_8799.n49 gnd 0.007799f
C856 a_n8964_8799.n50 gnd 0.011788f
C857 a_n8964_8799.n51 gnd 0.008106f
C858 a_n8964_8799.n53 gnd 4.05e-19
C859 a_n8964_8799.n54 gnd 0.008401f
C860 a_n8964_8799.n55 gnd 0.011603f
C861 a_n8964_8799.n56 gnd 0.007477f
C862 a_n8964_8799.n57 gnd 0.008684f
C863 a_n8964_8799.n58 gnd 0.001166f
C864 a_n8964_8799.n60 gnd 0.007799f
C865 a_n8964_8799.n61 gnd 0.011788f
C866 a_n8964_8799.n62 gnd 0.008106f
C867 a_n8964_8799.n64 gnd 4.05e-19
C868 a_n8964_8799.n65 gnd 0.008401f
C869 a_n8964_8799.n66 gnd 0.011603f
C870 a_n8964_8799.n67 gnd 0.007477f
C871 a_n8964_8799.n68 gnd 0.008684f
C872 a_n8964_8799.n69 gnd 0.001166f
C873 a_n8964_8799.n71 gnd 0.007799f
C874 a_n8964_8799.n72 gnd 0.011788f
C875 a_n8964_8799.n73 gnd 0.008106f
C876 a_n8964_8799.n75 gnd 4.05e-19
C877 a_n8964_8799.n76 gnd 0.008401f
C878 a_n8964_8799.n77 gnd 0.011603f
C879 a_n8964_8799.n78 gnd 0.007477f
C880 a_n8964_8799.n79 gnd 0.001166f
C881 a_n8964_8799.n81 gnd 0.007799f
C882 a_n8964_8799.n82 gnd 0.011788f
C883 a_n8964_8799.n83 gnd 0.008106f
C884 a_n8964_8799.n85 gnd 4.05e-19
C885 a_n8964_8799.n86 gnd 0.008401f
C886 a_n8964_8799.n87 gnd 0.011603f
C887 a_n8964_8799.n88 gnd 0.007477f
C888 a_n8964_8799.n89 gnd 0.252072f
C889 a_n8964_8799.n90 gnd 0.001166f
C890 a_n8964_8799.n92 gnd 0.007799f
C891 a_n8964_8799.n93 gnd 0.011788f
C892 a_n8964_8799.n94 gnd 0.008106f
C893 a_n8964_8799.n96 gnd 4.05e-19
C894 a_n8964_8799.n97 gnd 0.008401f
C895 a_n8964_8799.n98 gnd 0.011603f
C896 a_n8964_8799.n99 gnd 0.007477f
C897 a_n8964_8799.n100 gnd 0.252072f
C898 a_n8964_8799.n101 gnd 0.001166f
C899 a_n8964_8799.n103 gnd 0.007799f
C900 a_n8964_8799.n104 gnd 0.011788f
C901 a_n8964_8799.n105 gnd 0.008106f
C902 a_n8964_8799.n107 gnd 4.05e-19
C903 a_n8964_8799.n108 gnd 0.008401f
C904 a_n8964_8799.n109 gnd 0.011603f
C905 a_n8964_8799.n110 gnd 0.007477f
C906 a_n8964_8799.n111 gnd 0.252072f
C907 a_n8964_8799.t33 gnd 0.145227f
C908 a_n8964_8799.t21 gnd 0.145227f
C909 a_n8964_8799.t16 gnd 0.145227f
C910 a_n8964_8799.n112 gnd 1.14543f
C911 a_n8964_8799.t18 gnd 0.145227f
C912 a_n8964_8799.t29 gnd 0.145227f
C913 a_n8964_8799.n113 gnd 1.14354f
C914 a_n8964_8799.t20 gnd 0.145227f
C915 a_n8964_8799.t24 gnd 0.145227f
C916 a_n8964_8799.n114 gnd 1.14354f
C917 a_n8964_8799.t23 gnd 0.145227f
C918 a_n8964_8799.t35 gnd 0.145227f
C919 a_n8964_8799.n115 gnd 1.14354f
C920 a_n8964_8799.t15 gnd 0.145227f
C921 a_n8964_8799.t28 gnd 0.145227f
C922 a_n8964_8799.n116 gnd 1.14354f
C923 a_n8964_8799.t32 gnd 0.145227f
C924 a_n8964_8799.t25 gnd 0.145227f
C925 a_n8964_8799.n117 gnd 1.14354f
C926 a_n8964_8799.t6 gnd 0.112954f
C927 a_n8964_8799.t11 gnd 0.112954f
C928 a_n8964_8799.n118 gnd 1.00105f
C929 a_n8964_8799.t8 gnd 0.112954f
C930 a_n8964_8799.t10 gnd 0.112954f
C931 a_n8964_8799.n119 gnd 0.998105f
C932 a_n8964_8799.t40 gnd 0.112954f
C933 a_n8964_8799.t37 gnd 0.112954f
C934 a_n8964_8799.n120 gnd 0.998105f
C935 a_n8964_8799.t0 gnd 0.112954f
C936 a_n8964_8799.t3 gnd 0.112954f
C937 a_n8964_8799.n121 gnd 1.00105f
C938 a_n8964_8799.t39 gnd 0.112954f
C939 a_n8964_8799.t42 gnd 0.112954f
C940 a_n8964_8799.n122 gnd 0.998104f
C941 a_n8964_8799.t38 gnd 0.112954f
C942 a_n8964_8799.t41 gnd 0.112954f
C943 a_n8964_8799.n123 gnd 0.998104f
C944 a_n8964_8799.t4 gnd 0.112954f
C945 a_n8964_8799.t9 gnd 0.112954f
C946 a_n8964_8799.n124 gnd 1.00105f
C947 a_n8964_8799.t7 gnd 0.112954f
C948 a_n8964_8799.t1 gnd 0.112954f
C949 a_n8964_8799.n125 gnd 0.998104f
C950 a_n8964_8799.t43 gnd 0.112954f
C951 a_n8964_8799.t12 gnd 0.112954f
C952 a_n8964_8799.n126 gnd 0.998105f
C953 a_n8964_8799.t2 gnd 0.112954f
C954 a_n8964_8799.t5 gnd 0.112954f
C955 a_n8964_8799.n127 gnd 0.998105f
C956 a_n8964_8799.t81 gnd 0.602179f
C957 a_n8964_8799.n128 gnd 0.269219f
C958 a_n8964_8799.t110 gnd 0.602179f
C959 a_n8964_8799.t126 gnd 0.602179f
C960 a_n8964_8799.n129 gnd 0.272555f
C961 a_n8964_8799.t127 gnd 0.602179f
C962 a_n8964_8799.t69 gnd 0.602179f
C963 a_n8964_8799.t70 gnd 0.602179f
C964 a_n8964_8799.n130 gnd 0.274655f
C965 a_n8964_8799.t103 gnd 0.602179f
C966 a_n8964_8799.t108 gnd 0.602179f
C967 a_n8964_8799.n131 gnd 0.268138f
C968 a_n8964_8799.t83 gnd 0.613577f
C969 a_n8964_8799.n132 gnd 0.25246f
C970 a_n8964_8799.n133 gnd 0.011878f
C971 a_n8964_8799.t46 gnd 0.602179f
C972 a_n8964_8799.n134 gnd 0.268945f
C973 a_n8964_8799.n135 gnd 0.27254f
C974 a_n8964_8799.t130 gnd 0.602179f
C975 a_n8964_8799.n136 gnd 0.269035f
C976 a_n8964_8799.n137 gnd 0.26362f
C977 a_n8964_8799.t99 gnd 0.602179f
C978 a_n8964_8799.n138 gnd 0.268783f
C979 a_n8964_8799.n139 gnd 0.275093f
C980 a_n8964_8799.t84 gnd 0.602179f
C981 a_n8964_8799.n140 gnd 0.272422f
C982 a_n8964_8799.n141 gnd 0.268461f
C983 a_n8964_8799.t125 gnd 0.602179f
C984 a_n8964_8799.n142 gnd 0.263943f
C985 a_n8964_8799.t82 gnd 0.602179f
C986 a_n8964_8799.n143 gnd 0.272539f
C987 a_n8964_8799.t107 gnd 0.613566f
C988 a_n8964_8799.t90 gnd 0.602179f
C989 a_n8964_8799.n144 gnd 0.269219f
C990 a_n8964_8799.t122 gnd 0.602179f
C991 a_n8964_8799.t136 gnd 0.602179f
C992 a_n8964_8799.n145 gnd 0.272555f
C993 a_n8964_8799.t138 gnd 0.602179f
C994 a_n8964_8799.t76 gnd 0.602179f
C995 a_n8964_8799.t79 gnd 0.602179f
C996 a_n8964_8799.n146 gnd 0.274655f
C997 a_n8964_8799.t112 gnd 0.602179f
C998 a_n8964_8799.t118 gnd 0.602179f
C999 a_n8964_8799.n147 gnd 0.268138f
C1000 a_n8964_8799.t91 gnd 0.613577f
C1001 a_n8964_8799.n148 gnd 0.25246f
C1002 a_n8964_8799.n149 gnd 0.011878f
C1003 a_n8964_8799.t56 gnd 0.602179f
C1004 a_n8964_8799.n150 gnd 0.268945f
C1005 a_n8964_8799.n151 gnd 0.27254f
C1006 a_n8964_8799.t139 gnd 0.602179f
C1007 a_n8964_8799.n152 gnd 0.269035f
C1008 a_n8964_8799.n153 gnd 0.26362f
C1009 a_n8964_8799.t109 gnd 0.602179f
C1010 a_n8964_8799.n154 gnd 0.268783f
C1011 a_n8964_8799.n155 gnd 0.275093f
C1012 a_n8964_8799.t95 gnd 0.602179f
C1013 a_n8964_8799.n156 gnd 0.272422f
C1014 a_n8964_8799.n157 gnd 0.268461f
C1015 a_n8964_8799.t135 gnd 0.602179f
C1016 a_n8964_8799.n158 gnd 0.263943f
C1017 a_n8964_8799.t92 gnd 0.602179f
C1018 a_n8964_8799.n159 gnd 0.272539f
C1019 a_n8964_8799.t119 gnd 0.613566f
C1020 a_n8964_8799.n160 gnd 0.906949f
C1021 a_n8964_8799.t62 gnd 0.602179f
C1022 a_n8964_8799.n161 gnd 0.269219f
C1023 a_n8964_8799.t77 gnd 0.602179f
C1024 a_n8964_8799.t105 gnd 0.602179f
C1025 a_n8964_8799.n162 gnd 0.272555f
C1026 a_n8964_8799.t89 gnd 0.602179f
C1027 a_n8964_8799.t93 gnd 0.602179f
C1028 a_n8964_8799.t60 gnd 0.602179f
C1029 a_n8964_8799.n163 gnd 0.274655f
C1030 a_n8964_8799.t114 gnd 0.602179f
C1031 a_n8964_8799.t47 gnd 0.602179f
C1032 a_n8964_8799.n164 gnd 0.268138f
C1033 a_n8964_8799.t85 gnd 0.613577f
C1034 a_n8964_8799.n165 gnd 0.25246f
C1035 a_n8964_8799.n166 gnd 0.011878f
C1036 a_n8964_8799.t100 gnd 0.602179f
C1037 a_n8964_8799.n167 gnd 0.268945f
C1038 a_n8964_8799.n168 gnd 0.27254f
C1039 a_n8964_8799.t72 gnd 0.602179f
C1040 a_n8964_8799.n169 gnd 0.269035f
C1041 a_n8964_8799.n170 gnd 0.26362f
C1042 a_n8964_8799.t54 gnd 0.602179f
C1043 a_n8964_8799.n171 gnd 0.268783f
C1044 a_n8964_8799.n172 gnd 0.275093f
C1045 a_n8964_8799.t121 gnd 0.602179f
C1046 a_n8964_8799.n173 gnd 0.272422f
C1047 a_n8964_8799.n174 gnd 0.268461f
C1048 a_n8964_8799.t128 gnd 0.602179f
C1049 a_n8964_8799.n175 gnd 0.263943f
C1050 a_n8964_8799.t44 gnd 0.602179f
C1051 a_n8964_8799.n176 gnd 0.272539f
C1052 a_n8964_8799.t96 gnd 0.613566f
C1053 a_n8964_8799.n177 gnd 1.91248f
C1054 a_n8964_8799.t51 gnd 0.602179f
C1055 a_n8964_8799.t49 gnd 0.602179f
C1056 a_n8964_8799.t117 gnd 0.602179f
C1057 a_n8964_8799.n178 gnd 0.272139f
C1058 a_n8964_8799.t65 gnd 0.602179f
C1059 a_n8964_8799.t53 gnd 0.602179f
C1060 a_n8964_8799.t123 gnd 0.602179f
C1061 a_n8964_8799.n179 gnd 0.269035f
C1062 a_n8964_8799.t86 gnd 0.602179f
C1063 a_n8964_8799.t66 gnd 0.602179f
C1064 a_n8964_8799.t137 gnd 0.602179f
C1065 a_n8964_8799.n180 gnd 0.272555f
C1066 a_n8964_8799.t102 gnd 0.602179f
C1067 a_n8964_8799.t68 gnd 0.602179f
C1068 a_n8964_8799.t133 gnd 0.602179f
C1069 a_n8964_8799.n181 gnd 0.268461f
C1070 a_n8964_8799.t104 gnd 0.602179f
C1071 a_n8964_8799.t80 gnd 0.602179f
C1072 a_n8964_8799.t50 gnd 0.602179f
C1073 a_n8964_8799.n182 gnd 0.272539f
C1074 a_n8964_8799.t120 gnd 0.613577f
C1075 a_n8964_8799.n183 gnd 0.25246f
C1076 a_n8964_8799.n184 gnd 0.269219f
C1077 a_n8964_8799.n185 gnd 0.263943f
C1078 a_n8964_8799.n186 gnd 0.272422f
C1079 a_n8964_8799.n187 gnd 0.275093f
C1080 a_n8964_8799.n188 gnd 0.268783f
C1081 a_n8964_8799.n189 gnd 0.26362f
C1082 a_n8964_8799.n190 gnd 0.27254f
C1083 a_n8964_8799.n191 gnd 0.274655f
C1084 a_n8964_8799.n192 gnd 0.268138f
C1085 a_n8964_8799.n193 gnd 0.263458f
C1086 a_n8964_8799.t59 gnd 0.602179f
C1087 a_n8964_8799.t57 gnd 0.602179f
C1088 a_n8964_8799.t131 gnd 0.602179f
C1089 a_n8964_8799.n194 gnd 0.272139f
C1090 a_n8964_8799.t71 gnd 0.602179f
C1091 a_n8964_8799.t63 gnd 0.602179f
C1092 a_n8964_8799.t134 gnd 0.602179f
C1093 a_n8964_8799.n195 gnd 0.269035f
C1094 a_n8964_8799.t98 gnd 0.602179f
C1095 a_n8964_8799.t74 gnd 0.602179f
C1096 a_n8964_8799.t52 gnd 0.602179f
C1097 a_n8964_8799.n196 gnd 0.272555f
C1098 a_n8964_8799.t111 gnd 0.602179f
C1099 a_n8964_8799.t75 gnd 0.602179f
C1100 a_n8964_8799.t45 gnd 0.602179f
C1101 a_n8964_8799.n197 gnd 0.268461f
C1102 a_n8964_8799.t116 gnd 0.602179f
C1103 a_n8964_8799.t88 gnd 0.602179f
C1104 a_n8964_8799.t58 gnd 0.602179f
C1105 a_n8964_8799.n198 gnd 0.272539f
C1106 a_n8964_8799.t132 gnd 0.613577f
C1107 a_n8964_8799.n199 gnd 0.25246f
C1108 a_n8964_8799.n200 gnd 0.269219f
C1109 a_n8964_8799.n201 gnd 0.263943f
C1110 a_n8964_8799.n202 gnd 0.272422f
C1111 a_n8964_8799.n203 gnd 0.275093f
C1112 a_n8964_8799.n204 gnd 0.268783f
C1113 a_n8964_8799.n205 gnd 0.26362f
C1114 a_n8964_8799.n206 gnd 0.27254f
C1115 a_n8964_8799.n207 gnd 0.274655f
C1116 a_n8964_8799.n208 gnd 0.268138f
C1117 a_n8964_8799.n209 gnd 0.263458f
C1118 a_n8964_8799.n210 gnd 0.906949f
C1119 a_n8964_8799.t97 gnd 0.602179f
C1120 a_n8964_8799.t115 gnd 0.602179f
C1121 a_n8964_8799.t64 gnd 0.602179f
C1122 a_n8964_8799.n211 gnd 0.272139f
C1123 a_n8964_8799.t129 gnd 0.602179f
C1124 a_n8964_8799.t78 gnd 0.602179f
C1125 a_n8964_8799.t124 gnd 0.602179f
C1126 a_n8964_8799.n212 gnd 0.269035f
C1127 a_n8964_8799.t67 gnd 0.602179f
C1128 a_n8964_8799.t106 gnd 0.602179f
C1129 a_n8964_8799.t55 gnd 0.602179f
C1130 a_n8964_8799.n213 gnd 0.272555f
C1131 a_n8964_8799.t94 gnd 0.602179f
C1132 a_n8964_8799.t73 gnd 0.602179f
C1133 a_n8964_8799.t113 gnd 0.602179f
C1134 a_n8964_8799.n214 gnd 0.268461f
C1135 a_n8964_8799.t61 gnd 0.602179f
C1136 a_n8964_8799.t101 gnd 0.602179f
C1137 a_n8964_8799.t48 gnd 0.602179f
C1138 a_n8964_8799.n215 gnd 0.272539f
C1139 a_n8964_8799.t87 gnd 0.613577f
C1140 a_n8964_8799.n216 gnd 0.25246f
C1141 a_n8964_8799.n217 gnd 0.269219f
C1142 a_n8964_8799.n218 gnd 0.263943f
C1143 a_n8964_8799.n219 gnd 0.272422f
C1144 a_n8964_8799.n220 gnd 0.275093f
C1145 a_n8964_8799.n221 gnd 0.268783f
C1146 a_n8964_8799.n222 gnd 0.26362f
C1147 a_n8964_8799.n223 gnd 0.27254f
C1148 a_n8964_8799.n224 gnd 0.274655f
C1149 a_n8964_8799.n225 gnd 0.268138f
C1150 a_n8964_8799.n226 gnd 0.263458f
C1151 a_n8964_8799.n227 gnd 1.38861f
C1152 a_n8964_8799.n228 gnd 17.488302f
C1153 a_n8964_8799.n229 gnd 4.40708f
C1154 a_n8964_8799.n230 gnd 7.68272f
C1155 a_n8964_8799.t22 gnd 0.145227f
C1156 a_n8964_8799.t27 gnd 0.145227f
C1157 a_n8964_8799.n231 gnd 1.14354f
C1158 a_n8964_8799.t30 gnd 0.145227f
C1159 a_n8964_8799.t14 gnd 0.145227f
C1160 a_n8964_8799.n232 gnd 1.14354f
C1161 a_n8964_8799.t17 gnd 0.145227f
C1162 a_n8964_8799.t34 gnd 0.145227f
C1163 a_n8964_8799.n233 gnd 1.14543f
C1164 a_n8964_8799.t36 gnd 0.145227f
C1165 a_n8964_8799.t31 gnd 0.145227f
C1166 a_n8964_8799.n234 gnd 1.14354f
C1167 a_n8964_8799.t19 gnd 0.145227f
C1168 a_n8964_8799.t26 gnd 0.145227f
C1169 a_n8964_8799.n235 gnd 1.14354f
C1170 a_n8964_8799.n236 gnd 1.14354f
C1171 a_n8964_8799.t13 gnd 0.145227f
C1172 CSoutput.n0 gnd 0.045852f
C1173 CSoutput.t226 gnd 0.303299f
C1174 CSoutput.n1 gnd 0.136954f
C1175 CSoutput.n2 gnd 0.045852f
C1176 CSoutput.t224 gnd 0.303299f
C1177 CSoutput.n3 gnd 0.036341f
C1178 CSoutput.n4 gnd 0.045852f
C1179 CSoutput.t217 gnd 0.303299f
C1180 CSoutput.n5 gnd 0.031337f
C1181 CSoutput.n6 gnd 0.045852f
C1182 CSoutput.t221 gnd 0.303299f
C1183 CSoutput.t231 gnd 0.303299f
C1184 CSoutput.n7 gnd 0.135462f
C1185 CSoutput.n8 gnd 0.045852f
C1186 CSoutput.t229 gnd 0.303299f
C1187 CSoutput.n9 gnd 0.029878f
C1188 CSoutput.n10 gnd 0.045852f
C1189 CSoutput.t218 gnd 0.303299f
C1190 CSoutput.t223 gnd 0.303299f
C1191 CSoutput.n11 gnd 0.135462f
C1192 CSoutput.n12 gnd 0.045852f
C1193 CSoutput.t228 gnd 0.303299f
C1194 CSoutput.n13 gnd 0.031337f
C1195 CSoutput.n14 gnd 0.045852f
C1196 CSoutput.t233 gnd 0.303299f
C1197 CSoutput.t220 gnd 0.303299f
C1198 CSoutput.n15 gnd 0.135462f
C1199 CSoutput.n16 gnd 0.045852f
C1200 CSoutput.t227 gnd 0.303299f
C1201 CSoutput.n17 gnd 0.03347f
C1202 CSoutput.t235 gnd 0.36245f
C1203 CSoutput.t225 gnd 0.303299f
C1204 CSoutput.n18 gnd 0.172932f
C1205 CSoutput.n19 gnd 0.167804f
C1206 CSoutput.n20 gnd 0.194673f
C1207 CSoutput.n21 gnd 0.045852f
C1208 CSoutput.n22 gnd 0.038268f
C1209 CSoutput.n23 gnd 0.135462f
C1210 CSoutput.n24 gnd 0.03689f
C1211 CSoutput.n25 gnd 0.036341f
C1212 CSoutput.n26 gnd 0.045852f
C1213 CSoutput.n27 gnd 0.045852f
C1214 CSoutput.n28 gnd 0.037974f
C1215 CSoutput.n29 gnd 0.032241f
C1216 CSoutput.n30 gnd 0.138477f
C1217 CSoutput.n31 gnd 0.032685f
C1218 CSoutput.n32 gnd 0.045852f
C1219 CSoutput.n33 gnd 0.045852f
C1220 CSoutput.n34 gnd 0.045852f
C1221 CSoutput.n35 gnd 0.03757f
C1222 CSoutput.n36 gnd 0.135462f
C1223 CSoutput.n37 gnd 0.03593f
C1224 CSoutput.n38 gnd 0.037301f
C1225 CSoutput.n39 gnd 0.045852f
C1226 CSoutput.n40 gnd 0.045852f
C1227 CSoutput.n41 gnd 0.03826f
C1228 CSoutput.n42 gnd 0.03497f
C1229 CSoutput.n43 gnd 0.135462f
C1230 CSoutput.n44 gnd 0.035857f
C1231 CSoutput.n45 gnd 0.045852f
C1232 CSoutput.n46 gnd 0.045852f
C1233 CSoutput.n47 gnd 0.045852f
C1234 CSoutput.n48 gnd 0.035857f
C1235 CSoutput.n49 gnd 0.135462f
C1236 CSoutput.n50 gnd 0.03497f
C1237 CSoutput.n51 gnd 0.03826f
C1238 CSoutput.n52 gnd 0.045852f
C1239 CSoutput.n53 gnd 0.045852f
C1240 CSoutput.n54 gnd 0.037301f
C1241 CSoutput.n55 gnd 0.03593f
C1242 CSoutput.n56 gnd 0.135462f
C1243 CSoutput.n57 gnd 0.03757f
C1244 CSoutput.n58 gnd 0.045852f
C1245 CSoutput.n59 gnd 0.045852f
C1246 CSoutput.n60 gnd 0.045852f
C1247 CSoutput.n61 gnd 0.032685f
C1248 CSoutput.n62 gnd 0.138477f
C1249 CSoutput.n63 gnd 0.032241f
C1250 CSoutput.t234 gnd 0.303299f
C1251 CSoutput.n64 gnd 0.135462f
C1252 CSoutput.n65 gnd 0.037974f
C1253 CSoutput.n66 gnd 0.045852f
C1254 CSoutput.n67 gnd 0.045852f
C1255 CSoutput.n68 gnd 0.045852f
C1256 CSoutput.n69 gnd 0.03689f
C1257 CSoutput.n70 gnd 0.135462f
C1258 CSoutput.n71 gnd 0.038268f
C1259 CSoutput.n72 gnd 0.03347f
C1260 CSoutput.n73 gnd 0.045852f
C1261 CSoutput.n74 gnd 0.045852f
C1262 CSoutput.n75 gnd 0.034711f
C1263 CSoutput.n76 gnd 0.020615f
C1264 CSoutput.t236 gnd 0.340778f
C1265 CSoutput.n77 gnd 0.169285f
C1266 CSoutput.n78 gnd 0.692536f
C1267 CSoutput.t2 gnd 0.057193f
C1268 CSoutput.t174 gnd 0.057193f
C1269 CSoutput.n79 gnd 0.442811f
C1270 CSoutput.t126 gnd 0.057193f
C1271 CSoutput.t178 gnd 0.057193f
C1272 CSoutput.n80 gnd 0.442021f
C1273 CSoutput.n81 gnd 0.448651f
C1274 CSoutput.t149 gnd 0.057193f
C1275 CSoutput.t197 gnd 0.057193f
C1276 CSoutput.n82 gnd 0.442021f
C1277 CSoutput.n83 gnd 0.221076f
C1278 CSoutput.t141 gnd 0.057193f
C1279 CSoutput.t187 gnd 0.057193f
C1280 CSoutput.n84 gnd 0.442021f
C1281 CSoutput.n85 gnd 0.221076f
C1282 CSoutput.t131 gnd 0.057193f
C1283 CSoutput.t188 gnd 0.057193f
C1284 CSoutput.n86 gnd 0.442021f
C1285 CSoutput.n87 gnd 0.221076f
C1286 CSoutput.t150 gnd 0.057193f
C1287 CSoutput.t154 gnd 0.057193f
C1288 CSoutput.n88 gnd 0.442021f
C1289 CSoutput.n89 gnd 0.221076f
C1290 CSoutput.t194 gnd 0.057193f
C1291 CSoutput.t166 gnd 0.057193f
C1292 CSoutput.n90 gnd 0.442021f
C1293 CSoutput.n91 gnd 0.221076f
C1294 CSoutput.t171 gnd 0.057193f
C1295 CSoutput.t181 gnd 0.057193f
C1296 CSoutput.n92 gnd 0.442021f
C1297 CSoutput.n93 gnd 0.405403f
C1298 CSoutput.t130 gnd 0.057193f
C1299 CSoutput.t183 gnd 0.057193f
C1300 CSoutput.n94 gnd 0.442811f
C1301 CSoutput.t159 gnd 0.057193f
C1302 CSoutput.t176 gnd 0.057193f
C1303 CSoutput.n95 gnd 0.442021f
C1304 CSoutput.n96 gnd 0.448651f
C1305 CSoutput.t1 gnd 0.057193f
C1306 CSoutput.t214 gnd 0.057193f
C1307 CSoutput.n97 gnd 0.442021f
C1308 CSoutput.n98 gnd 0.221076f
C1309 CSoutput.t200 gnd 0.057193f
C1310 CSoutput.t124 gnd 0.057193f
C1311 CSoutput.n99 gnd 0.442021f
C1312 CSoutput.n100 gnd 0.221076f
C1313 CSoutput.t196 gnd 0.057193f
C1314 CSoutput.t185 gnd 0.057193f
C1315 CSoutput.n101 gnd 0.442021f
C1316 CSoutput.n102 gnd 0.221076f
C1317 CSoutput.t208 gnd 0.057193f
C1318 CSoutput.t125 gnd 0.057193f
C1319 CSoutput.n103 gnd 0.442021f
C1320 CSoutput.n104 gnd 0.221076f
C1321 CSoutput.t206 gnd 0.057193f
C1322 CSoutput.t193 gnd 0.057193f
C1323 CSoutput.n105 gnd 0.442021f
C1324 CSoutput.n106 gnd 0.221076f
C1325 CSoutput.t177 gnd 0.057193f
C1326 CSoutput.t182 gnd 0.057193f
C1327 CSoutput.n107 gnd 0.442021f
C1328 CSoutput.n108 gnd 0.32968f
C1329 CSoutput.n109 gnd 0.415725f
C1330 CSoutput.t142 gnd 0.057193f
C1331 CSoutput.t169 gnd 0.057193f
C1332 CSoutput.n110 gnd 0.442811f
C1333 CSoutput.t147 gnd 0.057193f
C1334 CSoutput.t133 gnd 0.057193f
C1335 CSoutput.n111 gnd 0.442021f
C1336 CSoutput.n112 gnd 0.448651f
C1337 CSoutput.t170 gnd 0.057193f
C1338 CSoutput.t136 gnd 0.057193f
C1339 CSoutput.n113 gnd 0.442021f
C1340 CSoutput.n114 gnd 0.221076f
C1341 CSoutput.t128 gnd 0.057193f
C1342 CSoutput.t129 gnd 0.057193f
C1343 CSoutput.n115 gnd 0.442021f
C1344 CSoutput.n116 gnd 0.221076f
C1345 CSoutput.t205 gnd 0.057193f
C1346 CSoutput.t153 gnd 0.057193f
C1347 CSoutput.n117 gnd 0.442021f
C1348 CSoutput.n118 gnd 0.221076f
C1349 CSoutput.t191 gnd 0.057193f
C1350 CSoutput.t138 gnd 0.057193f
C1351 CSoutput.n119 gnd 0.442021f
C1352 CSoutput.n120 gnd 0.221076f
C1353 CSoutput.t180 gnd 0.057193f
C1354 CSoutput.t210 gnd 0.057193f
C1355 CSoutput.n121 gnd 0.442021f
C1356 CSoutput.n122 gnd 0.221076f
C1357 CSoutput.t143 gnd 0.057193f
C1358 CSoutput.t184 gnd 0.057193f
C1359 CSoutput.n123 gnd 0.442021f
C1360 CSoutput.n124 gnd 0.32968f
C1361 CSoutput.n125 gnd 0.464674f
C1362 CSoutput.n126 gnd 9.31196f
C1363 CSoutput.n128 gnd 0.811108f
C1364 CSoutput.n129 gnd 0.608331f
C1365 CSoutput.n130 gnd 0.811108f
C1366 CSoutput.n131 gnd 0.811108f
C1367 CSoutput.n132 gnd 2.18375f
C1368 CSoutput.n133 gnd 0.811108f
C1369 CSoutput.n134 gnd 0.811108f
C1370 CSoutput.t230 gnd 1.01388f
C1371 CSoutput.n135 gnd 0.811108f
C1372 CSoutput.n136 gnd 0.811108f
C1373 CSoutput.n140 gnd 0.811108f
C1374 CSoutput.n144 gnd 0.811108f
C1375 CSoutput.n145 gnd 0.811108f
C1376 CSoutput.n147 gnd 0.811108f
C1377 CSoutput.n152 gnd 0.811108f
C1378 CSoutput.n154 gnd 0.811108f
C1379 CSoutput.n155 gnd 0.811108f
C1380 CSoutput.n157 gnd 0.811108f
C1381 CSoutput.n158 gnd 0.811108f
C1382 CSoutput.n160 gnd 0.811108f
C1383 CSoutput.t219 gnd 13.5535f
C1384 CSoutput.n162 gnd 0.811108f
C1385 CSoutput.n163 gnd 0.608331f
C1386 CSoutput.n164 gnd 0.811108f
C1387 CSoutput.n165 gnd 0.811108f
C1388 CSoutput.n166 gnd 2.18375f
C1389 CSoutput.n167 gnd 0.811108f
C1390 CSoutput.n168 gnd 0.811108f
C1391 CSoutput.t237 gnd 1.01388f
C1392 CSoutput.n169 gnd 0.811108f
C1393 CSoutput.n170 gnd 0.811108f
C1394 CSoutput.n174 gnd 0.811108f
C1395 CSoutput.n178 gnd 0.811108f
C1396 CSoutput.n179 gnd 0.811108f
C1397 CSoutput.n181 gnd 0.811108f
C1398 CSoutput.n186 gnd 0.811108f
C1399 CSoutput.n188 gnd 0.811108f
C1400 CSoutput.n189 gnd 0.811108f
C1401 CSoutput.n191 gnd 0.811108f
C1402 CSoutput.n192 gnd 0.811108f
C1403 CSoutput.n194 gnd 0.811108f
C1404 CSoutput.n195 gnd 0.608331f
C1405 CSoutput.n197 gnd 0.811108f
C1406 CSoutput.n198 gnd 0.608331f
C1407 CSoutput.n199 gnd 0.811108f
C1408 CSoutput.n200 gnd 0.811108f
C1409 CSoutput.n201 gnd 2.18375f
C1410 CSoutput.n202 gnd 0.811108f
C1411 CSoutput.n203 gnd 0.811108f
C1412 CSoutput.t232 gnd 1.01388f
C1413 CSoutput.n204 gnd 0.811108f
C1414 CSoutput.n205 gnd 2.18375f
C1415 CSoutput.n207 gnd 0.811108f
C1416 CSoutput.n208 gnd 0.811108f
C1417 CSoutput.n210 gnd 0.811108f
C1418 CSoutput.n211 gnd 0.811108f
C1419 CSoutput.t216 gnd 13.3326f
C1420 CSoutput.t222 gnd 13.5535f
C1421 CSoutput.n217 gnd 2.54456f
C1422 CSoutput.n218 gnd 10.3656f
C1423 CSoutput.n219 gnd 10.7994f
C1424 CSoutput.n224 gnd 2.75645f
C1425 CSoutput.n230 gnd 0.811108f
C1426 CSoutput.n232 gnd 0.811108f
C1427 CSoutput.n234 gnd 0.811108f
C1428 CSoutput.n236 gnd 0.811108f
C1429 CSoutput.n238 gnd 0.811108f
C1430 CSoutput.n244 gnd 0.811108f
C1431 CSoutput.n251 gnd 1.48807f
C1432 CSoutput.n252 gnd 1.48807f
C1433 CSoutput.n253 gnd 0.811108f
C1434 CSoutput.n254 gnd 0.811108f
C1435 CSoutput.n256 gnd 0.608331f
C1436 CSoutput.n257 gnd 0.520981f
C1437 CSoutput.n259 gnd 0.608331f
C1438 CSoutput.n260 gnd 0.520981f
C1439 CSoutput.n261 gnd 0.608331f
C1440 CSoutput.n263 gnd 0.811108f
C1441 CSoutput.n265 gnd 2.18375f
C1442 CSoutput.n266 gnd 2.54456f
C1443 CSoutput.n267 gnd 9.53371f
C1444 CSoutput.n269 gnd 0.608331f
C1445 CSoutput.n270 gnd 1.56527f
C1446 CSoutput.n271 gnd 0.608331f
C1447 CSoutput.n273 gnd 0.811108f
C1448 CSoutput.n275 gnd 2.18375f
C1449 CSoutput.n276 gnd 4.75656f
C1450 CSoutput.t175 gnd 0.057193f
C1451 CSoutput.t151 gnd 0.057193f
C1452 CSoutput.n277 gnd 0.442811f
C1453 CSoutput.t134 gnd 0.057193f
C1454 CSoutput.t127 gnd 0.057193f
C1455 CSoutput.n278 gnd 0.442021f
C1456 CSoutput.n279 gnd 0.448651f
C1457 CSoutput.t192 gnd 0.057193f
C1458 CSoutput.t146 gnd 0.057193f
C1459 CSoutput.n280 gnd 0.442021f
C1460 CSoutput.n281 gnd 0.221076f
C1461 CSoutput.t163 gnd 0.057193f
C1462 CSoutput.t168 gnd 0.057193f
C1463 CSoutput.n282 gnd 0.442021f
C1464 CSoutput.n283 gnd 0.221076f
C1465 CSoutput.t189 gnd 0.057193f
C1466 CSoutput.t0 gnd 0.057193f
C1467 CSoutput.n284 gnd 0.442021f
C1468 CSoutput.n285 gnd 0.221076f
C1469 CSoutput.t155 gnd 0.057193f
C1470 CSoutput.t209 gnd 0.057193f
C1471 CSoutput.n286 gnd 0.442021f
C1472 CSoutput.n287 gnd 0.221076f
C1473 CSoutput.t167 gnd 0.057193f
C1474 CSoutput.t195 gnd 0.057193f
C1475 CSoutput.n288 gnd 0.442021f
C1476 CSoutput.n289 gnd 0.221076f
C1477 CSoutput.t198 gnd 0.057193f
C1478 CSoutput.t165 gnd 0.057193f
C1479 CSoutput.n290 gnd 0.442021f
C1480 CSoutput.n291 gnd 0.405403f
C1481 CSoutput.t213 gnd 0.057193f
C1482 CSoutput.t207 gnd 0.057193f
C1483 CSoutput.n292 gnd 0.442811f
C1484 CSoutput.t139 gnd 0.057193f
C1485 CSoutput.t211 gnd 0.057193f
C1486 CSoutput.n293 gnd 0.442021f
C1487 CSoutput.n294 gnd 0.448651f
C1488 CSoutput.t179 gnd 0.057193f
C1489 CSoutput.t158 gnd 0.057193f
C1490 CSoutput.n295 gnd 0.442021f
C1491 CSoutput.n296 gnd 0.221076f
C1492 CSoutput.t152 gnd 0.057193f
C1493 CSoutput.t160 gnd 0.057193f
C1494 CSoutput.n297 gnd 0.442021f
C1495 CSoutput.n298 gnd 0.221076f
C1496 CSoutput.t172 gnd 0.057193f
C1497 CSoutput.t137 gnd 0.057193f
C1498 CSoutput.n299 gnd 0.442021f
C1499 CSoutput.n300 gnd 0.221076f
C1500 CSoutput.t161 gnd 0.057193f
C1501 CSoutput.t3 gnd 0.057193f
C1502 CSoutput.n301 gnd 0.442021f
C1503 CSoutput.n302 gnd 0.221076f
C1504 CSoutput.t202 gnd 0.057193f
C1505 CSoutput.t186 gnd 0.057193f
C1506 CSoutput.n303 gnd 0.442021f
C1507 CSoutput.n304 gnd 0.221076f
C1508 CSoutput.t212 gnd 0.057193f
C1509 CSoutput.t156 gnd 0.057193f
C1510 CSoutput.n305 gnd 0.442021f
C1511 CSoutput.n306 gnd 0.32968f
C1512 CSoutput.n307 gnd 0.415725f
C1513 CSoutput.t145 gnd 0.057193f
C1514 CSoutput.t199 gnd 0.057193f
C1515 CSoutput.n308 gnd 0.442811f
C1516 CSoutput.t203 gnd 0.057193f
C1517 CSoutput.t135 gnd 0.057193f
C1518 CSoutput.n309 gnd 0.442021f
C1519 CSoutput.n310 gnd 0.448651f
C1520 CSoutput.t173 gnd 0.057193f
C1521 CSoutput.t215 gnd 0.057193f
C1522 CSoutput.n311 gnd 0.442021f
C1523 CSoutput.n312 gnd 0.221076f
C1524 CSoutput.t164 gnd 0.057193f
C1525 CSoutput.t162 gnd 0.057193f
C1526 CSoutput.n313 gnd 0.442021f
C1527 CSoutput.n314 gnd 0.221076f
C1528 CSoutput.t201 gnd 0.057193f
C1529 CSoutput.t190 gnd 0.057193f
C1530 CSoutput.n315 gnd 0.442021f
C1531 CSoutput.n316 gnd 0.221076f
C1532 CSoutput.t204 gnd 0.057193f
C1533 CSoutput.t157 gnd 0.057193f
C1534 CSoutput.n317 gnd 0.442021f
C1535 CSoutput.n318 gnd 0.221076f
C1536 CSoutput.t140 gnd 0.057193f
C1537 CSoutput.t132 gnd 0.057193f
C1538 CSoutput.n319 gnd 0.442021f
C1539 CSoutput.n320 gnd 0.221076f
C1540 CSoutput.t144 gnd 0.057193f
C1541 CSoutput.t148 gnd 0.057193f
C1542 CSoutput.n321 gnd 0.44202f
C1543 CSoutput.n322 gnd 0.329682f
C1544 CSoutput.n323 gnd 0.464674f
C1545 CSoutput.n324 gnd 13.004299f
C1546 CSoutput.t52 gnd 0.050044f
C1547 CSoutput.t120 gnd 0.050044f
C1548 CSoutput.n325 gnd 0.443689f
C1549 CSoutput.t42 gnd 0.050044f
C1550 CSoutput.t51 gnd 0.050044f
C1551 CSoutput.n326 gnd 0.442209f
C1552 CSoutput.n327 gnd 0.412056f
C1553 CSoutput.t32 gnd 0.050044f
C1554 CSoutput.t58 gnd 0.050044f
C1555 CSoutput.n328 gnd 0.442209f
C1556 CSoutput.n329 gnd 0.203124f
C1557 CSoutput.t79 gnd 0.050044f
C1558 CSoutput.t45 gnd 0.050044f
C1559 CSoutput.n330 gnd 0.442209f
C1560 CSoutput.n331 gnd 0.203124f
C1561 CSoutput.t55 gnd 0.050044f
C1562 CSoutput.t110 gnd 0.050044f
C1563 CSoutput.n332 gnd 0.442209f
C1564 CSoutput.n333 gnd 0.203124f
C1565 CSoutput.t72 gnd 0.050044f
C1566 CSoutput.t86 gnd 0.050044f
C1567 CSoutput.n334 gnd 0.442209f
C1568 CSoutput.n335 gnd 0.203124f
C1569 CSoutput.t27 gnd 0.050044f
C1570 CSoutput.t59 gnd 0.050044f
C1571 CSoutput.n336 gnd 0.442209f
C1572 CSoutput.n337 gnd 0.203124f
C1573 CSoutput.t13 gnd 0.050044f
C1574 CSoutput.t39 gnd 0.050044f
C1575 CSoutput.n338 gnd 0.442209f
C1576 CSoutput.n339 gnd 0.203124f
C1577 CSoutput.t92 gnd 0.050044f
C1578 CSoutput.t103 gnd 0.050044f
C1579 CSoutput.n340 gnd 0.442209f
C1580 CSoutput.n341 gnd 0.203124f
C1581 CSoutput.t119 gnd 0.050044f
C1582 CSoutput.t63 gnd 0.050044f
C1583 CSoutput.n342 gnd 0.442209f
C1584 CSoutput.n343 gnd 0.374652f
C1585 CSoutput.t115 gnd 0.050044f
C1586 CSoutput.t5 gnd 0.050044f
C1587 CSoutput.n344 gnd 0.443689f
C1588 CSoutput.t17 gnd 0.050044f
C1589 CSoutput.t108 gnd 0.050044f
C1590 CSoutput.n345 gnd 0.442209f
C1591 CSoutput.n346 gnd 0.412056f
C1592 CSoutput.t7 gnd 0.050044f
C1593 CSoutput.t98 gnd 0.050044f
C1594 CSoutput.n347 gnd 0.442209f
C1595 CSoutput.n348 gnd 0.203124f
C1596 CSoutput.t109 gnd 0.050044f
C1597 CSoutput.t6 gnd 0.050044f
C1598 CSoutput.n349 gnd 0.442209f
C1599 CSoutput.n350 gnd 0.203124f
C1600 CSoutput.t88 gnd 0.050044f
C1601 CSoutput.t62 gnd 0.050044f
C1602 CSoutput.n351 gnd 0.442209f
C1603 CSoutput.n352 gnd 0.203124f
C1604 CSoutput.t8 gnd 0.050044f
C1605 CSoutput.t90 gnd 0.050044f
C1606 CSoutput.n353 gnd 0.442209f
C1607 CSoutput.n354 gnd 0.203124f
C1608 CSoutput.t65 gnd 0.050044f
C1609 CSoutput.t73 gnd 0.050044f
C1610 CSoutput.n355 gnd 0.442209f
C1611 CSoutput.n356 gnd 0.203124f
C1612 CSoutput.t89 gnd 0.050044f
C1613 CSoutput.t64 gnd 0.050044f
C1614 CSoutput.n357 gnd 0.442209f
C1615 CSoutput.n358 gnd 0.203124f
C1616 CSoutput.t74 gnd 0.050044f
C1617 CSoutput.t78 gnd 0.050044f
C1618 CSoutput.n359 gnd 0.442209f
C1619 CSoutput.n360 gnd 0.203124f
C1620 CSoutput.t56 gnd 0.050044f
C1621 CSoutput.t69 gnd 0.050044f
C1622 CSoutput.n361 gnd 0.442209f
C1623 CSoutput.n362 gnd 0.308386f
C1624 CSoutput.n363 gnd 0.388971f
C1625 CSoutput.t20 gnd 0.050044f
C1626 CSoutput.t111 gnd 0.050044f
C1627 CSoutput.n364 gnd 0.443689f
C1628 CSoutput.t40 gnd 0.050044f
C1629 CSoutput.t46 gnd 0.050044f
C1630 CSoutput.n365 gnd 0.442209f
C1631 CSoutput.n366 gnd 0.412056f
C1632 CSoutput.t9 gnd 0.050044f
C1633 CSoutput.t93 gnd 0.050044f
C1634 CSoutput.n367 gnd 0.442209f
C1635 CSoutput.n368 gnd 0.203124f
C1636 CSoutput.t54 gnd 0.050044f
C1637 CSoutput.t21 gnd 0.050044f
C1638 CSoutput.n369 gnd 0.442209f
C1639 CSoutput.n370 gnd 0.203124f
C1640 CSoutput.t30 gnd 0.050044f
C1641 CSoutput.t123 gnd 0.050044f
C1642 CSoutput.n371 gnd 0.442209f
C1643 CSoutput.n372 gnd 0.203124f
C1644 CSoutput.t31 gnd 0.050044f
C1645 CSoutput.t35 gnd 0.050044f
C1646 CSoutput.n373 gnd 0.442209f
C1647 CSoutput.n374 gnd 0.203124f
C1648 CSoutput.t16 gnd 0.050044f
C1649 CSoutput.t107 gnd 0.050044f
C1650 CSoutput.n375 gnd 0.442209f
C1651 CSoutput.n376 gnd 0.203124f
C1652 CSoutput.t38 gnd 0.050044f
C1653 CSoutput.t28 gnd 0.050044f
C1654 CSoutput.n377 gnd 0.442209f
C1655 CSoutput.n378 gnd 0.203124f
C1656 CSoutput.t4 gnd 0.050044f
C1657 CSoutput.t48 gnd 0.050044f
C1658 CSoutput.n379 gnd 0.442209f
C1659 CSoutput.n380 gnd 0.203124f
C1660 CSoutput.t53 gnd 0.050044f
C1661 CSoutput.t19 gnd 0.050044f
C1662 CSoutput.n381 gnd 0.442209f
C1663 CSoutput.n382 gnd 0.308386f
C1664 CSoutput.n383 gnd 0.417694f
C1665 CSoutput.n384 gnd 13.2702f
C1666 CSoutput.t34 gnd 0.050044f
C1667 CSoutput.t91 gnd 0.050044f
C1668 CSoutput.n385 gnd 0.443689f
C1669 CSoutput.t87 gnd 0.050044f
C1670 CSoutput.t61 gnd 0.050044f
C1671 CSoutput.n386 gnd 0.442209f
C1672 CSoutput.n387 gnd 0.412056f
C1673 CSoutput.t95 gnd 0.050044f
C1674 CSoutput.t49 gnd 0.050044f
C1675 CSoutput.n388 gnd 0.442209f
C1676 CSoutput.n389 gnd 0.203124f
C1677 CSoutput.t75 gnd 0.050044f
C1678 CSoutput.t113 gnd 0.050044f
C1679 CSoutput.n390 gnd 0.442209f
C1680 CSoutput.n391 gnd 0.203124f
C1681 CSoutput.t29 gnd 0.050044f
C1682 CSoutput.t94 gnd 0.050044f
C1683 CSoutput.n392 gnd 0.442209f
C1684 CSoutput.n393 gnd 0.203124f
C1685 CSoutput.t15 gnd 0.050044f
C1686 CSoutput.t101 gnd 0.050044f
C1687 CSoutput.n394 gnd 0.442209f
C1688 CSoutput.n395 gnd 0.203124f
C1689 CSoutput.t100 gnd 0.050044f
C1690 CSoutput.t41 gnd 0.050044f
C1691 CSoutput.n396 gnd 0.442209f
C1692 CSoutput.n397 gnd 0.203124f
C1693 CSoutput.t68 gnd 0.050044f
C1694 CSoutput.t37 gnd 0.050044f
C1695 CSoutput.n398 gnd 0.442209f
C1696 CSoutput.n399 gnd 0.203124f
C1697 CSoutput.t43 gnd 0.050044f
C1698 CSoutput.t18 gnd 0.050044f
C1699 CSoutput.n400 gnd 0.442209f
C1700 CSoutput.n401 gnd 0.203124f
C1701 CSoutput.t26 gnd 0.050044f
C1702 CSoutput.t44 gnd 0.050044f
C1703 CSoutput.n402 gnd 0.442209f
C1704 CSoutput.n403 gnd 0.374652f
C1705 CSoutput.t23 gnd 0.050044f
C1706 CSoutput.t14 gnd 0.050044f
C1707 CSoutput.n404 gnd 0.443689f
C1708 CSoutput.t10 gnd 0.050044f
C1709 CSoutput.t121 gnd 0.050044f
C1710 CSoutput.n405 gnd 0.442209f
C1711 CSoutput.n406 gnd 0.412056f
C1712 CSoutput.t122 gnd 0.050044f
C1713 CSoutput.t24 gnd 0.050044f
C1714 CSoutput.n407 gnd 0.442209f
C1715 CSoutput.n408 gnd 0.203124f
C1716 CSoutput.t25 gnd 0.050044f
C1717 CSoutput.t82 gnd 0.050044f
C1718 CSoutput.n409 gnd 0.442209f
C1719 CSoutput.n410 gnd 0.203124f
C1720 CSoutput.t83 gnd 0.050044f
C1721 CSoutput.t114 gnd 0.050044f
C1722 CSoutput.n411 gnd 0.442209f
C1723 CSoutput.n412 gnd 0.203124f
C1724 CSoutput.t117 gnd 0.050044f
C1725 CSoutput.t106 gnd 0.050044f
C1726 CSoutput.n413 gnd 0.442209f
C1727 CSoutput.n414 gnd 0.203124f
C1728 CSoutput.t97 gnd 0.050044f
C1729 CSoutput.t84 gnd 0.050044f
C1730 CSoutput.n415 gnd 0.442209f
C1731 CSoutput.n416 gnd 0.203124f
C1732 CSoutput.t85 gnd 0.050044f
C1733 CSoutput.t118 gnd 0.050044f
C1734 CSoutput.n417 gnd 0.442209f
C1735 CSoutput.n418 gnd 0.203124f
C1736 CSoutput.t71 gnd 0.050044f
C1737 CSoutput.t99 gnd 0.050044f
C1738 CSoutput.n419 gnd 0.442209f
C1739 CSoutput.n420 gnd 0.203124f
C1740 CSoutput.t105 gnd 0.050044f
C1741 CSoutput.t80 gnd 0.050044f
C1742 CSoutput.n421 gnd 0.442209f
C1743 CSoutput.n422 gnd 0.308386f
C1744 CSoutput.n423 gnd 0.388971f
C1745 CSoutput.t70 gnd 0.050044f
C1746 CSoutput.t102 gnd 0.050044f
C1747 CSoutput.n424 gnd 0.443689f
C1748 CSoutput.t33 gnd 0.050044f
C1749 CSoutput.t50 gnd 0.050044f
C1750 CSoutput.n425 gnd 0.442209f
C1751 CSoutput.n426 gnd 0.412056f
C1752 CSoutput.t60 gnd 0.050044f
C1753 CSoutput.t81 gnd 0.050044f
C1754 CSoutput.n427 gnd 0.442209f
C1755 CSoutput.n428 gnd 0.203124f
C1756 CSoutput.t104 gnd 0.050044f
C1757 CSoutput.t66 gnd 0.050044f
C1758 CSoutput.n429 gnd 0.442209f
C1759 CSoutput.n430 gnd 0.203124f
C1760 CSoutput.t76 gnd 0.050044f
C1761 CSoutput.t116 gnd 0.050044f
C1762 CSoutput.n431 gnd 0.442209f
C1763 CSoutput.n432 gnd 0.203124f
C1764 CSoutput.t11 gnd 0.050044f
C1765 CSoutput.t36 gnd 0.050044f
C1766 CSoutput.n433 gnd 0.442209f
C1767 CSoutput.n434 gnd 0.203124f
C1768 CSoutput.t67 gnd 0.050044f
C1769 CSoutput.t96 gnd 0.050044f
C1770 CSoutput.n435 gnd 0.442209f
C1771 CSoutput.n436 gnd 0.203124f
C1772 CSoutput.t112 gnd 0.050044f
C1773 CSoutput.t22 gnd 0.050044f
C1774 CSoutput.n437 gnd 0.442209f
C1775 CSoutput.n438 gnd 0.203124f
C1776 CSoutput.t57 gnd 0.050044f
C1777 CSoutput.t77 gnd 0.050044f
C1778 CSoutput.n439 gnd 0.442209f
C1779 CSoutput.n440 gnd 0.203124f
C1780 CSoutput.t12 gnd 0.050044f
C1781 CSoutput.t47 gnd 0.050044f
C1782 CSoutput.n441 gnd 0.442209f
C1783 CSoutput.n442 gnd 0.308386f
C1784 CSoutput.n443 gnd 0.417694f
C1785 CSoutput.n444 gnd 7.97774f
C1786 CSoutput.n445 gnd 13.8895f
C1787 commonsourceibias.n0 gnd 0.012817f
C1788 commonsourceibias.t151 gnd 0.194086f
C1789 commonsourceibias.t83 gnd 0.17946f
C1790 commonsourceibias.n1 gnd 0.009349f
C1791 commonsourceibias.n2 gnd 0.009605f
C1792 commonsourceibias.t161 gnd 0.17946f
C1793 commonsourceibias.n3 gnd 0.012358f
C1794 commonsourceibias.n4 gnd 0.009605f
C1795 commonsourceibias.t152 gnd 0.17946f
C1796 commonsourceibias.n5 gnd 0.071604f
C1797 commonsourceibias.t171 gnd 0.17946f
C1798 commonsourceibias.n6 gnd 0.009057f
C1799 commonsourceibias.n7 gnd 0.009605f
C1800 commonsourceibias.t145 gnd 0.17946f
C1801 commonsourceibias.n8 gnd 0.012174f
C1802 commonsourceibias.n9 gnd 0.009605f
C1803 commonsourceibias.t124 gnd 0.17946f
C1804 commonsourceibias.n10 gnd 0.071604f
C1805 commonsourceibias.t158 gnd 0.17946f
C1806 commonsourceibias.n11 gnd 0.008798f
C1807 commonsourceibias.n12 gnd 0.009605f
C1808 commonsourceibias.t148 gnd 0.17946f
C1809 commonsourceibias.n13 gnd 0.01197f
C1810 commonsourceibias.n14 gnd 0.012817f
C1811 commonsourceibias.t66 gnd 0.194086f
C1812 commonsourceibias.t10 gnd 0.17946f
C1813 commonsourceibias.n15 gnd 0.009349f
C1814 commonsourceibias.n16 gnd 0.009605f
C1815 commonsourceibias.t58 gnd 0.17946f
C1816 commonsourceibias.n17 gnd 0.012358f
C1817 commonsourceibias.n18 gnd 0.009605f
C1818 commonsourceibias.t64 gnd 0.17946f
C1819 commonsourceibias.n19 gnd 0.071604f
C1820 commonsourceibias.t2 gnd 0.17946f
C1821 commonsourceibias.n20 gnd 0.009057f
C1822 commonsourceibias.n21 gnd 0.009605f
C1823 commonsourceibias.t70 gnd 0.17946f
C1824 commonsourceibias.n22 gnd 0.012174f
C1825 commonsourceibias.n23 gnd 0.009605f
C1826 commonsourceibias.t54 gnd 0.17946f
C1827 commonsourceibias.n24 gnd 0.071604f
C1828 commonsourceibias.t60 gnd 0.17946f
C1829 commonsourceibias.n25 gnd 0.008798f
C1830 commonsourceibias.n26 gnd 0.009605f
C1831 commonsourceibias.t68 gnd 0.17946f
C1832 commonsourceibias.n27 gnd 0.01197f
C1833 commonsourceibias.n28 gnd 0.009605f
C1834 commonsourceibias.t30 gnd 0.17946f
C1835 commonsourceibias.n29 gnd 0.071604f
C1836 commonsourceibias.t50 gnd 0.17946f
C1837 commonsourceibias.n30 gnd 0.008571f
C1838 commonsourceibias.n31 gnd 0.009605f
C1839 commonsourceibias.t24 gnd 0.17946f
C1840 commonsourceibias.n32 gnd 0.011742f
C1841 commonsourceibias.n33 gnd 0.009605f
C1842 commonsourceibias.t78 gnd 0.17946f
C1843 commonsourceibias.n34 gnd 0.071604f
C1844 commonsourceibias.t18 gnd 0.17946f
C1845 commonsourceibias.n35 gnd 0.008375f
C1846 commonsourceibias.n36 gnd 0.009605f
C1847 commonsourceibias.t6 gnd 0.17946f
C1848 commonsourceibias.n37 gnd 0.011489f
C1849 commonsourceibias.n38 gnd 0.009605f
C1850 commonsourceibias.t14 gnd 0.17946f
C1851 commonsourceibias.n39 gnd 0.071604f
C1852 commonsourceibias.t42 gnd 0.17946f
C1853 commonsourceibias.n40 gnd 0.008208f
C1854 commonsourceibias.n41 gnd 0.009605f
C1855 commonsourceibias.t28 gnd 0.17946f
C1856 commonsourceibias.n42 gnd 0.011208f
C1857 commonsourceibias.t22 gnd 0.199526f
C1858 commonsourceibias.t4 gnd 0.17946f
C1859 commonsourceibias.n43 gnd 0.078221f
C1860 commonsourceibias.n44 gnd 0.085838f
C1861 commonsourceibias.n45 gnd 0.03983f
C1862 commonsourceibias.n46 gnd 0.009605f
C1863 commonsourceibias.n47 gnd 0.009349f
C1864 commonsourceibias.n48 gnd 0.013398f
C1865 commonsourceibias.n49 gnd 0.071604f
C1866 commonsourceibias.n50 gnd 0.013389f
C1867 commonsourceibias.n51 gnd 0.009605f
C1868 commonsourceibias.n52 gnd 0.009605f
C1869 commonsourceibias.n53 gnd 0.009605f
C1870 commonsourceibias.n54 gnd 0.012358f
C1871 commonsourceibias.n55 gnd 0.071604f
C1872 commonsourceibias.n56 gnd 0.012648f
C1873 commonsourceibias.n57 gnd 0.012288f
C1874 commonsourceibias.n58 gnd 0.009605f
C1875 commonsourceibias.n59 gnd 0.009605f
C1876 commonsourceibias.n60 gnd 0.009605f
C1877 commonsourceibias.n61 gnd 0.009057f
C1878 commonsourceibias.n62 gnd 0.01341f
C1879 commonsourceibias.n63 gnd 0.071604f
C1880 commonsourceibias.n64 gnd 0.013406f
C1881 commonsourceibias.n65 gnd 0.009605f
C1882 commonsourceibias.n66 gnd 0.009605f
C1883 commonsourceibias.n67 gnd 0.009605f
C1884 commonsourceibias.n68 gnd 0.012174f
C1885 commonsourceibias.n69 gnd 0.071604f
C1886 commonsourceibias.n70 gnd 0.012558f
C1887 commonsourceibias.n71 gnd 0.012378f
C1888 commonsourceibias.n72 gnd 0.009605f
C1889 commonsourceibias.n73 gnd 0.009605f
C1890 commonsourceibias.n74 gnd 0.009605f
C1891 commonsourceibias.n75 gnd 0.008798f
C1892 commonsourceibias.n76 gnd 0.013415f
C1893 commonsourceibias.n77 gnd 0.071604f
C1894 commonsourceibias.n78 gnd 0.013414f
C1895 commonsourceibias.n79 gnd 0.009605f
C1896 commonsourceibias.n80 gnd 0.009605f
C1897 commonsourceibias.n81 gnd 0.009605f
C1898 commonsourceibias.n82 gnd 0.01197f
C1899 commonsourceibias.n83 gnd 0.071604f
C1900 commonsourceibias.n84 gnd 0.012468f
C1901 commonsourceibias.n85 gnd 0.012468f
C1902 commonsourceibias.n86 gnd 0.009605f
C1903 commonsourceibias.n87 gnd 0.009605f
C1904 commonsourceibias.n88 gnd 0.009605f
C1905 commonsourceibias.n89 gnd 0.008571f
C1906 commonsourceibias.n90 gnd 0.013414f
C1907 commonsourceibias.n91 gnd 0.071604f
C1908 commonsourceibias.n92 gnd 0.013415f
C1909 commonsourceibias.n93 gnd 0.009605f
C1910 commonsourceibias.n94 gnd 0.009605f
C1911 commonsourceibias.n95 gnd 0.009605f
C1912 commonsourceibias.n96 gnd 0.011742f
C1913 commonsourceibias.n97 gnd 0.071604f
C1914 commonsourceibias.n98 gnd 0.012378f
C1915 commonsourceibias.n99 gnd 0.012558f
C1916 commonsourceibias.n100 gnd 0.009605f
C1917 commonsourceibias.n101 gnd 0.009605f
C1918 commonsourceibias.n102 gnd 0.009605f
C1919 commonsourceibias.n103 gnd 0.008375f
C1920 commonsourceibias.n104 gnd 0.013406f
C1921 commonsourceibias.n105 gnd 0.071604f
C1922 commonsourceibias.n106 gnd 0.01341f
C1923 commonsourceibias.n107 gnd 0.009605f
C1924 commonsourceibias.n108 gnd 0.009605f
C1925 commonsourceibias.n109 gnd 0.009605f
C1926 commonsourceibias.n110 gnd 0.011489f
C1927 commonsourceibias.n111 gnd 0.071604f
C1928 commonsourceibias.n112 gnd 0.012288f
C1929 commonsourceibias.n113 gnd 0.012648f
C1930 commonsourceibias.n114 gnd 0.009605f
C1931 commonsourceibias.n115 gnd 0.009605f
C1932 commonsourceibias.n116 gnd 0.009605f
C1933 commonsourceibias.n117 gnd 0.008208f
C1934 commonsourceibias.n118 gnd 0.013389f
C1935 commonsourceibias.n119 gnd 0.071604f
C1936 commonsourceibias.n120 gnd 0.013398f
C1937 commonsourceibias.n121 gnd 0.009605f
C1938 commonsourceibias.n122 gnd 0.009605f
C1939 commonsourceibias.n123 gnd 0.009605f
C1940 commonsourceibias.n124 gnd 0.011208f
C1941 commonsourceibias.n125 gnd 0.071604f
C1942 commonsourceibias.n126 gnd 0.011785f
C1943 commonsourceibias.n127 gnd 0.085919f
C1944 commonsourceibias.n128 gnd 0.095702f
C1945 commonsourceibias.t67 gnd 0.020728f
C1946 commonsourceibias.t11 gnd 0.020728f
C1947 commonsourceibias.n129 gnd 0.183157f
C1948 commonsourceibias.n130 gnd 0.158432f
C1949 commonsourceibias.t59 gnd 0.020728f
C1950 commonsourceibias.t65 gnd 0.020728f
C1951 commonsourceibias.n131 gnd 0.183157f
C1952 commonsourceibias.n132 gnd 0.084131f
C1953 commonsourceibias.t3 gnd 0.020728f
C1954 commonsourceibias.t71 gnd 0.020728f
C1955 commonsourceibias.n133 gnd 0.183157f
C1956 commonsourceibias.n134 gnd 0.084131f
C1957 commonsourceibias.t55 gnd 0.020728f
C1958 commonsourceibias.t61 gnd 0.020728f
C1959 commonsourceibias.n135 gnd 0.183157f
C1960 commonsourceibias.n136 gnd 0.084131f
C1961 commonsourceibias.t69 gnd 0.020728f
C1962 commonsourceibias.t31 gnd 0.020728f
C1963 commonsourceibias.n137 gnd 0.183157f
C1964 commonsourceibias.n138 gnd 0.070287f
C1965 commonsourceibias.t5 gnd 0.020728f
C1966 commonsourceibias.t23 gnd 0.020728f
C1967 commonsourceibias.n139 gnd 0.18377f
C1968 commonsourceibias.t43 gnd 0.020728f
C1969 commonsourceibias.t29 gnd 0.020728f
C1970 commonsourceibias.n140 gnd 0.183157f
C1971 commonsourceibias.n141 gnd 0.170668f
C1972 commonsourceibias.t7 gnd 0.020728f
C1973 commonsourceibias.t15 gnd 0.020728f
C1974 commonsourceibias.n142 gnd 0.183157f
C1975 commonsourceibias.n143 gnd 0.084131f
C1976 commonsourceibias.t79 gnd 0.020728f
C1977 commonsourceibias.t19 gnd 0.020728f
C1978 commonsourceibias.n144 gnd 0.183157f
C1979 commonsourceibias.n145 gnd 0.084131f
C1980 commonsourceibias.t51 gnd 0.020728f
C1981 commonsourceibias.t25 gnd 0.020728f
C1982 commonsourceibias.n146 gnd 0.183157f
C1983 commonsourceibias.n147 gnd 0.070287f
C1984 commonsourceibias.n148 gnd 0.085111f
C1985 commonsourceibias.n149 gnd 0.062167f
C1986 commonsourceibias.t93 gnd 0.17946f
C1987 commonsourceibias.n150 gnd 0.071604f
C1988 commonsourceibias.t131 gnd 0.17946f
C1989 commonsourceibias.n151 gnd 0.071604f
C1990 commonsourceibias.n152 gnd 0.009605f
C1991 commonsourceibias.t117 gnd 0.17946f
C1992 commonsourceibias.n153 gnd 0.071604f
C1993 commonsourceibias.n154 gnd 0.009605f
C1994 commonsourceibias.t176 gnd 0.17946f
C1995 commonsourceibias.n155 gnd 0.071604f
C1996 commonsourceibias.n156 gnd 0.009605f
C1997 commonsourceibias.t144 gnd 0.17946f
C1998 commonsourceibias.n157 gnd 0.008375f
C1999 commonsourceibias.n158 gnd 0.009605f
C2000 commonsourceibias.t190 gnd 0.17946f
C2001 commonsourceibias.n159 gnd 0.011489f
C2002 commonsourceibias.n160 gnd 0.009605f
C2003 commonsourceibias.t164 gnd 0.17946f
C2004 commonsourceibias.n161 gnd 0.071604f
C2005 commonsourceibias.t111 gnd 0.17946f
C2006 commonsourceibias.n162 gnd 0.008208f
C2007 commonsourceibias.n163 gnd 0.009605f
C2008 commonsourceibias.t100 gnd 0.17946f
C2009 commonsourceibias.n164 gnd 0.011208f
C2010 commonsourceibias.t140 gnd 0.199526f
C2011 commonsourceibias.t84 gnd 0.17946f
C2012 commonsourceibias.n165 gnd 0.078221f
C2013 commonsourceibias.n166 gnd 0.085838f
C2014 commonsourceibias.n167 gnd 0.03983f
C2015 commonsourceibias.n168 gnd 0.009605f
C2016 commonsourceibias.n169 gnd 0.009349f
C2017 commonsourceibias.n170 gnd 0.013398f
C2018 commonsourceibias.n171 gnd 0.071604f
C2019 commonsourceibias.n172 gnd 0.013389f
C2020 commonsourceibias.n173 gnd 0.009605f
C2021 commonsourceibias.n174 gnd 0.009605f
C2022 commonsourceibias.n175 gnd 0.009605f
C2023 commonsourceibias.n176 gnd 0.012358f
C2024 commonsourceibias.n177 gnd 0.071604f
C2025 commonsourceibias.n178 gnd 0.012648f
C2026 commonsourceibias.n179 gnd 0.012288f
C2027 commonsourceibias.n180 gnd 0.009605f
C2028 commonsourceibias.n181 gnd 0.009605f
C2029 commonsourceibias.n182 gnd 0.009605f
C2030 commonsourceibias.n183 gnd 0.009057f
C2031 commonsourceibias.n184 gnd 0.01341f
C2032 commonsourceibias.n185 gnd 0.071604f
C2033 commonsourceibias.n186 gnd 0.013406f
C2034 commonsourceibias.n187 gnd 0.009605f
C2035 commonsourceibias.n188 gnd 0.009605f
C2036 commonsourceibias.n189 gnd 0.009605f
C2037 commonsourceibias.n190 gnd 0.012174f
C2038 commonsourceibias.n191 gnd 0.071604f
C2039 commonsourceibias.n192 gnd 0.012558f
C2040 commonsourceibias.n193 gnd 0.012378f
C2041 commonsourceibias.n194 gnd 0.009605f
C2042 commonsourceibias.n195 gnd 0.009605f
C2043 commonsourceibias.n196 gnd 0.011742f
C2044 commonsourceibias.n197 gnd 0.008798f
C2045 commonsourceibias.n198 gnd 0.013415f
C2046 commonsourceibias.n199 gnd 0.009605f
C2047 commonsourceibias.n200 gnd 0.009605f
C2048 commonsourceibias.n201 gnd 0.013414f
C2049 commonsourceibias.n202 gnd 0.008571f
C2050 commonsourceibias.n203 gnd 0.01197f
C2051 commonsourceibias.n204 gnd 0.009605f
C2052 commonsourceibias.n205 gnd 0.008391f
C2053 commonsourceibias.n206 gnd 0.012468f
C2054 commonsourceibias.n207 gnd 0.012468f
C2055 commonsourceibias.n208 gnd 0.008391f
C2056 commonsourceibias.n209 gnd 0.009605f
C2057 commonsourceibias.n210 gnd 0.009605f
C2058 commonsourceibias.n211 gnd 0.008571f
C2059 commonsourceibias.n212 gnd 0.013414f
C2060 commonsourceibias.n213 gnd 0.071604f
C2061 commonsourceibias.n214 gnd 0.013415f
C2062 commonsourceibias.n215 gnd 0.009605f
C2063 commonsourceibias.n216 gnd 0.009605f
C2064 commonsourceibias.n217 gnd 0.009605f
C2065 commonsourceibias.n218 gnd 0.011742f
C2066 commonsourceibias.n219 gnd 0.071604f
C2067 commonsourceibias.n220 gnd 0.012378f
C2068 commonsourceibias.n221 gnd 0.012558f
C2069 commonsourceibias.n222 gnd 0.009605f
C2070 commonsourceibias.n223 gnd 0.009605f
C2071 commonsourceibias.n224 gnd 0.009605f
C2072 commonsourceibias.n225 gnd 0.008375f
C2073 commonsourceibias.n226 gnd 0.013406f
C2074 commonsourceibias.n227 gnd 0.071604f
C2075 commonsourceibias.n228 gnd 0.01341f
C2076 commonsourceibias.n229 gnd 0.009605f
C2077 commonsourceibias.n230 gnd 0.009605f
C2078 commonsourceibias.n231 gnd 0.009605f
C2079 commonsourceibias.n232 gnd 0.011489f
C2080 commonsourceibias.n233 gnd 0.071604f
C2081 commonsourceibias.n234 gnd 0.012288f
C2082 commonsourceibias.n235 gnd 0.012648f
C2083 commonsourceibias.n236 gnd 0.009605f
C2084 commonsourceibias.n237 gnd 0.009605f
C2085 commonsourceibias.n238 gnd 0.009605f
C2086 commonsourceibias.n239 gnd 0.008208f
C2087 commonsourceibias.n240 gnd 0.013389f
C2088 commonsourceibias.n241 gnd 0.071604f
C2089 commonsourceibias.n242 gnd 0.013398f
C2090 commonsourceibias.n243 gnd 0.009605f
C2091 commonsourceibias.n244 gnd 0.009605f
C2092 commonsourceibias.n245 gnd 0.009605f
C2093 commonsourceibias.n246 gnd 0.011208f
C2094 commonsourceibias.n247 gnd 0.071604f
C2095 commonsourceibias.n248 gnd 0.011785f
C2096 commonsourceibias.n249 gnd 0.085919f
C2097 commonsourceibias.n250 gnd 0.056156f
C2098 commonsourceibias.n251 gnd 0.012817f
C2099 commonsourceibias.t88 gnd 0.194086f
C2100 commonsourceibias.t198 gnd 0.17946f
C2101 commonsourceibias.n252 gnd 0.009349f
C2102 commonsourceibias.n253 gnd 0.009605f
C2103 commonsourceibias.t186 gnd 0.17946f
C2104 commonsourceibias.n254 gnd 0.012358f
C2105 commonsourceibias.n255 gnd 0.009605f
C2106 commonsourceibias.t95 gnd 0.17946f
C2107 commonsourceibias.n256 gnd 0.071604f
C2108 commonsourceibias.t196 gnd 0.17946f
C2109 commonsourceibias.n257 gnd 0.009057f
C2110 commonsourceibias.n258 gnd 0.009605f
C2111 commonsourceibias.t105 gnd 0.17946f
C2112 commonsourceibias.n259 gnd 0.012174f
C2113 commonsourceibias.n260 gnd 0.009605f
C2114 commonsourceibias.t94 gnd 0.17946f
C2115 commonsourceibias.n261 gnd 0.071604f
C2116 commonsourceibias.t197 gnd 0.17946f
C2117 commonsourceibias.n262 gnd 0.008798f
C2118 commonsourceibias.n263 gnd 0.009605f
C2119 commonsourceibias.t115 gnd 0.17946f
C2120 commonsourceibias.n264 gnd 0.01197f
C2121 commonsourceibias.n265 gnd 0.009605f
C2122 commonsourceibias.t141 gnd 0.17946f
C2123 commonsourceibias.n266 gnd 0.071604f
C2124 commonsourceibias.t195 gnd 0.17946f
C2125 commonsourceibias.n267 gnd 0.008571f
C2126 commonsourceibias.n268 gnd 0.009605f
C2127 commonsourceibias.t113 gnd 0.17946f
C2128 commonsourceibias.n269 gnd 0.011742f
C2129 commonsourceibias.n270 gnd 0.009605f
C2130 commonsourceibias.t138 gnd 0.17946f
C2131 commonsourceibias.n271 gnd 0.071604f
C2132 commonsourceibias.t130 gnd 0.17946f
C2133 commonsourceibias.n272 gnd 0.008375f
C2134 commonsourceibias.n273 gnd 0.009605f
C2135 commonsourceibias.t114 gnd 0.17946f
C2136 commonsourceibias.n274 gnd 0.011489f
C2137 commonsourceibias.n275 gnd 0.009605f
C2138 commonsourceibias.t139 gnd 0.17946f
C2139 commonsourceibias.n276 gnd 0.071604f
C2140 commonsourceibias.t129 gnd 0.17946f
C2141 commonsourceibias.n277 gnd 0.008208f
C2142 commonsourceibias.n278 gnd 0.009605f
C2143 commonsourceibias.t125 gnd 0.17946f
C2144 commonsourceibias.n279 gnd 0.011208f
C2145 commonsourceibias.t134 gnd 0.199526f
C2146 commonsourceibias.t147 gnd 0.17946f
C2147 commonsourceibias.n280 gnd 0.078221f
C2148 commonsourceibias.n281 gnd 0.085838f
C2149 commonsourceibias.n282 gnd 0.03983f
C2150 commonsourceibias.n283 gnd 0.009605f
C2151 commonsourceibias.n284 gnd 0.009349f
C2152 commonsourceibias.n285 gnd 0.013398f
C2153 commonsourceibias.n286 gnd 0.071604f
C2154 commonsourceibias.n287 gnd 0.013389f
C2155 commonsourceibias.n288 gnd 0.009605f
C2156 commonsourceibias.n289 gnd 0.009605f
C2157 commonsourceibias.n290 gnd 0.009605f
C2158 commonsourceibias.n291 gnd 0.012358f
C2159 commonsourceibias.n292 gnd 0.071604f
C2160 commonsourceibias.n293 gnd 0.012648f
C2161 commonsourceibias.n294 gnd 0.012288f
C2162 commonsourceibias.n295 gnd 0.009605f
C2163 commonsourceibias.n296 gnd 0.009605f
C2164 commonsourceibias.n297 gnd 0.009605f
C2165 commonsourceibias.n298 gnd 0.009057f
C2166 commonsourceibias.n299 gnd 0.01341f
C2167 commonsourceibias.n300 gnd 0.071604f
C2168 commonsourceibias.n301 gnd 0.013406f
C2169 commonsourceibias.n302 gnd 0.009605f
C2170 commonsourceibias.n303 gnd 0.009605f
C2171 commonsourceibias.n304 gnd 0.009605f
C2172 commonsourceibias.n305 gnd 0.012174f
C2173 commonsourceibias.n306 gnd 0.071604f
C2174 commonsourceibias.n307 gnd 0.012558f
C2175 commonsourceibias.n308 gnd 0.012378f
C2176 commonsourceibias.n309 gnd 0.009605f
C2177 commonsourceibias.n310 gnd 0.009605f
C2178 commonsourceibias.n311 gnd 0.009605f
C2179 commonsourceibias.n312 gnd 0.008798f
C2180 commonsourceibias.n313 gnd 0.013415f
C2181 commonsourceibias.n314 gnd 0.071604f
C2182 commonsourceibias.n315 gnd 0.013414f
C2183 commonsourceibias.n316 gnd 0.009605f
C2184 commonsourceibias.n317 gnd 0.009605f
C2185 commonsourceibias.n318 gnd 0.009605f
C2186 commonsourceibias.n319 gnd 0.01197f
C2187 commonsourceibias.n320 gnd 0.071604f
C2188 commonsourceibias.n321 gnd 0.012468f
C2189 commonsourceibias.n322 gnd 0.012468f
C2190 commonsourceibias.n323 gnd 0.009605f
C2191 commonsourceibias.n324 gnd 0.009605f
C2192 commonsourceibias.n325 gnd 0.009605f
C2193 commonsourceibias.n326 gnd 0.008571f
C2194 commonsourceibias.n327 gnd 0.013414f
C2195 commonsourceibias.n328 gnd 0.071604f
C2196 commonsourceibias.n329 gnd 0.013415f
C2197 commonsourceibias.n330 gnd 0.009605f
C2198 commonsourceibias.n331 gnd 0.009605f
C2199 commonsourceibias.n332 gnd 0.009605f
C2200 commonsourceibias.n333 gnd 0.011742f
C2201 commonsourceibias.n334 gnd 0.071604f
C2202 commonsourceibias.n335 gnd 0.012378f
C2203 commonsourceibias.n336 gnd 0.012558f
C2204 commonsourceibias.n337 gnd 0.009605f
C2205 commonsourceibias.n338 gnd 0.009605f
C2206 commonsourceibias.n339 gnd 0.009605f
C2207 commonsourceibias.n340 gnd 0.008375f
C2208 commonsourceibias.n341 gnd 0.013406f
C2209 commonsourceibias.n342 gnd 0.071604f
C2210 commonsourceibias.n343 gnd 0.01341f
C2211 commonsourceibias.n344 gnd 0.009605f
C2212 commonsourceibias.n345 gnd 0.009605f
C2213 commonsourceibias.n346 gnd 0.009605f
C2214 commonsourceibias.n347 gnd 0.011489f
C2215 commonsourceibias.n348 gnd 0.071604f
C2216 commonsourceibias.n349 gnd 0.012288f
C2217 commonsourceibias.n350 gnd 0.012648f
C2218 commonsourceibias.n351 gnd 0.009605f
C2219 commonsourceibias.n352 gnd 0.009605f
C2220 commonsourceibias.n353 gnd 0.009605f
C2221 commonsourceibias.n354 gnd 0.008208f
C2222 commonsourceibias.n355 gnd 0.013389f
C2223 commonsourceibias.n356 gnd 0.071604f
C2224 commonsourceibias.n357 gnd 0.013398f
C2225 commonsourceibias.n358 gnd 0.009605f
C2226 commonsourceibias.n359 gnd 0.009605f
C2227 commonsourceibias.n360 gnd 0.009605f
C2228 commonsourceibias.n361 gnd 0.011208f
C2229 commonsourceibias.n362 gnd 0.071604f
C2230 commonsourceibias.n363 gnd 0.011785f
C2231 commonsourceibias.n364 gnd 0.085919f
C2232 commonsourceibias.n365 gnd 0.029883f
C2233 commonsourceibias.n366 gnd 0.153509f
C2234 commonsourceibias.n367 gnd 0.012817f
C2235 commonsourceibias.t92 gnd 0.17946f
C2236 commonsourceibias.n368 gnd 0.009349f
C2237 commonsourceibias.n369 gnd 0.009605f
C2238 commonsourceibias.t163 gnd 0.17946f
C2239 commonsourceibias.n370 gnd 0.012358f
C2240 commonsourceibias.n371 gnd 0.009605f
C2241 commonsourceibias.t157 gnd 0.17946f
C2242 commonsourceibias.n372 gnd 0.071604f
C2243 commonsourceibias.t194 gnd 0.17946f
C2244 commonsourceibias.n373 gnd 0.009057f
C2245 commonsourceibias.n374 gnd 0.009605f
C2246 commonsourceibias.t110 gnd 0.17946f
C2247 commonsourceibias.n375 gnd 0.012174f
C2248 commonsourceibias.n376 gnd 0.009605f
C2249 commonsourceibias.t149 gnd 0.17946f
C2250 commonsourceibias.n377 gnd 0.071604f
C2251 commonsourceibias.t182 gnd 0.17946f
C2252 commonsourceibias.n378 gnd 0.008798f
C2253 commonsourceibias.n379 gnd 0.009605f
C2254 commonsourceibias.t173 gnd 0.17946f
C2255 commonsourceibias.n380 gnd 0.01197f
C2256 commonsourceibias.n381 gnd 0.009605f
C2257 commonsourceibias.t80 gnd 0.17946f
C2258 commonsourceibias.n382 gnd 0.071604f
C2259 commonsourceibias.t172 gnd 0.17946f
C2260 commonsourceibias.n383 gnd 0.008571f
C2261 commonsourceibias.n384 gnd 0.009605f
C2262 commonsourceibias.t168 gnd 0.17946f
C2263 commonsourceibias.n385 gnd 0.011742f
C2264 commonsourceibias.n386 gnd 0.009605f
C2265 commonsourceibias.t187 gnd 0.17946f
C2266 commonsourceibias.n387 gnd 0.071604f
C2267 commonsourceibias.t96 gnd 0.17946f
C2268 commonsourceibias.n388 gnd 0.008375f
C2269 commonsourceibias.n389 gnd 0.009605f
C2270 commonsourceibias.t165 gnd 0.17946f
C2271 commonsourceibias.n390 gnd 0.011489f
C2272 commonsourceibias.n391 gnd 0.009605f
C2273 commonsourceibias.t175 gnd 0.17946f
C2274 commonsourceibias.n392 gnd 0.071604f
C2275 commonsourceibias.t199 gnd 0.17946f
C2276 commonsourceibias.n393 gnd 0.008208f
C2277 commonsourceibias.n394 gnd 0.009605f
C2278 commonsourceibias.t155 gnd 0.17946f
C2279 commonsourceibias.n395 gnd 0.011208f
C2280 commonsourceibias.t184 gnd 0.199526f
C2281 commonsourceibias.t150 gnd 0.17946f
C2282 commonsourceibias.n396 gnd 0.078221f
C2283 commonsourceibias.n397 gnd 0.085838f
C2284 commonsourceibias.n398 gnd 0.03983f
C2285 commonsourceibias.n399 gnd 0.009605f
C2286 commonsourceibias.n400 gnd 0.009349f
C2287 commonsourceibias.n401 gnd 0.013398f
C2288 commonsourceibias.n402 gnd 0.071604f
C2289 commonsourceibias.n403 gnd 0.013389f
C2290 commonsourceibias.n404 gnd 0.009605f
C2291 commonsourceibias.n405 gnd 0.009605f
C2292 commonsourceibias.n406 gnd 0.009605f
C2293 commonsourceibias.n407 gnd 0.012358f
C2294 commonsourceibias.n408 gnd 0.071604f
C2295 commonsourceibias.n409 gnd 0.012648f
C2296 commonsourceibias.n410 gnd 0.012288f
C2297 commonsourceibias.n411 gnd 0.009605f
C2298 commonsourceibias.n412 gnd 0.009605f
C2299 commonsourceibias.n413 gnd 0.009605f
C2300 commonsourceibias.n414 gnd 0.009057f
C2301 commonsourceibias.n415 gnd 0.01341f
C2302 commonsourceibias.n416 gnd 0.071604f
C2303 commonsourceibias.n417 gnd 0.013406f
C2304 commonsourceibias.n418 gnd 0.009605f
C2305 commonsourceibias.n419 gnd 0.009605f
C2306 commonsourceibias.n420 gnd 0.009605f
C2307 commonsourceibias.n421 gnd 0.012174f
C2308 commonsourceibias.n422 gnd 0.071604f
C2309 commonsourceibias.n423 gnd 0.012558f
C2310 commonsourceibias.n424 gnd 0.012378f
C2311 commonsourceibias.n425 gnd 0.009605f
C2312 commonsourceibias.n426 gnd 0.009605f
C2313 commonsourceibias.n427 gnd 0.009605f
C2314 commonsourceibias.n428 gnd 0.008798f
C2315 commonsourceibias.n429 gnd 0.013415f
C2316 commonsourceibias.n430 gnd 0.071604f
C2317 commonsourceibias.n431 gnd 0.013414f
C2318 commonsourceibias.n432 gnd 0.009605f
C2319 commonsourceibias.n433 gnd 0.009605f
C2320 commonsourceibias.n434 gnd 0.009605f
C2321 commonsourceibias.n435 gnd 0.01197f
C2322 commonsourceibias.n436 gnd 0.071604f
C2323 commonsourceibias.n437 gnd 0.012468f
C2324 commonsourceibias.n438 gnd 0.012468f
C2325 commonsourceibias.n439 gnd 0.009605f
C2326 commonsourceibias.n440 gnd 0.009605f
C2327 commonsourceibias.n441 gnd 0.009605f
C2328 commonsourceibias.n442 gnd 0.008571f
C2329 commonsourceibias.n443 gnd 0.013414f
C2330 commonsourceibias.n444 gnd 0.071604f
C2331 commonsourceibias.n445 gnd 0.013415f
C2332 commonsourceibias.n446 gnd 0.009605f
C2333 commonsourceibias.n447 gnd 0.009605f
C2334 commonsourceibias.n448 gnd 0.009605f
C2335 commonsourceibias.n449 gnd 0.011742f
C2336 commonsourceibias.n450 gnd 0.071604f
C2337 commonsourceibias.n451 gnd 0.012378f
C2338 commonsourceibias.n452 gnd 0.012558f
C2339 commonsourceibias.n453 gnd 0.009605f
C2340 commonsourceibias.n454 gnd 0.009605f
C2341 commonsourceibias.n455 gnd 0.009605f
C2342 commonsourceibias.n456 gnd 0.008375f
C2343 commonsourceibias.n457 gnd 0.013406f
C2344 commonsourceibias.n458 gnd 0.071604f
C2345 commonsourceibias.n459 gnd 0.01341f
C2346 commonsourceibias.n460 gnd 0.009605f
C2347 commonsourceibias.n461 gnd 0.009605f
C2348 commonsourceibias.n462 gnd 0.009605f
C2349 commonsourceibias.n463 gnd 0.011489f
C2350 commonsourceibias.n464 gnd 0.071604f
C2351 commonsourceibias.n465 gnd 0.012288f
C2352 commonsourceibias.n466 gnd 0.012648f
C2353 commonsourceibias.n467 gnd 0.009605f
C2354 commonsourceibias.n468 gnd 0.009605f
C2355 commonsourceibias.n469 gnd 0.009605f
C2356 commonsourceibias.n470 gnd 0.008208f
C2357 commonsourceibias.n471 gnd 0.013389f
C2358 commonsourceibias.n472 gnd 0.071604f
C2359 commonsourceibias.n473 gnd 0.013398f
C2360 commonsourceibias.n474 gnd 0.009605f
C2361 commonsourceibias.n475 gnd 0.009605f
C2362 commonsourceibias.n476 gnd 0.009605f
C2363 commonsourceibias.n477 gnd 0.011208f
C2364 commonsourceibias.n478 gnd 0.071604f
C2365 commonsourceibias.n479 gnd 0.011785f
C2366 commonsourceibias.t183 gnd 0.194086f
C2367 commonsourceibias.n480 gnd 0.085919f
C2368 commonsourceibias.n481 gnd 0.029883f
C2369 commonsourceibias.n482 gnd 0.456424f
C2370 commonsourceibias.n483 gnd 0.012817f
C2371 commonsourceibias.t112 gnd 0.194086f
C2372 commonsourceibias.t169 gnd 0.17946f
C2373 commonsourceibias.n484 gnd 0.009349f
C2374 commonsourceibias.n485 gnd 0.009605f
C2375 commonsourceibias.t142 gnd 0.17946f
C2376 commonsourceibias.n486 gnd 0.012358f
C2377 commonsourceibias.n487 gnd 0.009605f
C2378 commonsourceibias.t154 gnd 0.17946f
C2379 commonsourceibias.n488 gnd 0.009057f
C2380 commonsourceibias.n489 gnd 0.009605f
C2381 commonsourceibias.t108 gnd 0.17946f
C2382 commonsourceibias.n490 gnd 0.012174f
C2383 commonsourceibias.n491 gnd 0.009605f
C2384 commonsourceibias.t128 gnd 0.17946f
C2385 commonsourceibias.n492 gnd 0.008798f
C2386 commonsourceibias.n493 gnd 0.009605f
C2387 commonsourceibias.t109 gnd 0.17946f
C2388 commonsourceibias.n494 gnd 0.01197f
C2389 commonsourceibias.t77 gnd 0.020728f
C2390 commonsourceibias.t17 gnd 0.020728f
C2391 commonsourceibias.n495 gnd 0.18377f
C2392 commonsourceibias.t63 gnd 0.020728f
C2393 commonsourceibias.t75 gnd 0.020728f
C2394 commonsourceibias.n496 gnd 0.183157f
C2395 commonsourceibias.n497 gnd 0.170668f
C2396 commonsourceibias.t49 gnd 0.020728f
C2397 commonsourceibias.t13 gnd 0.020728f
C2398 commonsourceibias.n498 gnd 0.183157f
C2399 commonsourceibias.n499 gnd 0.084131f
C2400 commonsourceibias.t47 gnd 0.020728f
C2401 commonsourceibias.t57 gnd 0.020728f
C2402 commonsourceibias.n500 gnd 0.183157f
C2403 commonsourceibias.n501 gnd 0.084131f
C2404 commonsourceibias.t73 gnd 0.020728f
C2405 commonsourceibias.t27 gnd 0.020728f
C2406 commonsourceibias.n502 gnd 0.183157f
C2407 commonsourceibias.n503 gnd 0.070287f
C2408 commonsourceibias.n504 gnd 0.012817f
C2409 commonsourceibias.t0 gnd 0.17946f
C2410 commonsourceibias.n505 gnd 0.009349f
C2411 commonsourceibias.n506 gnd 0.009605f
C2412 commonsourceibias.t20 gnd 0.17946f
C2413 commonsourceibias.n507 gnd 0.012358f
C2414 commonsourceibias.n508 gnd 0.009605f
C2415 commonsourceibias.t32 gnd 0.17946f
C2416 commonsourceibias.n509 gnd 0.009057f
C2417 commonsourceibias.n510 gnd 0.009605f
C2418 commonsourceibias.t44 gnd 0.17946f
C2419 commonsourceibias.n511 gnd 0.012174f
C2420 commonsourceibias.n512 gnd 0.009605f
C2421 commonsourceibias.t52 gnd 0.17946f
C2422 commonsourceibias.n513 gnd 0.008798f
C2423 commonsourceibias.n514 gnd 0.009605f
C2424 commonsourceibias.t36 gnd 0.17946f
C2425 commonsourceibias.n515 gnd 0.01197f
C2426 commonsourceibias.n516 gnd 0.009605f
C2427 commonsourceibias.t26 gnd 0.17946f
C2428 commonsourceibias.n517 gnd 0.008571f
C2429 commonsourceibias.n518 gnd 0.009605f
C2430 commonsourceibias.t72 gnd 0.17946f
C2431 commonsourceibias.n519 gnd 0.011742f
C2432 commonsourceibias.n520 gnd 0.009605f
C2433 commonsourceibias.t46 gnd 0.17946f
C2434 commonsourceibias.n521 gnd 0.008375f
C2435 commonsourceibias.n522 gnd 0.009605f
C2436 commonsourceibias.t12 gnd 0.17946f
C2437 commonsourceibias.n523 gnd 0.011489f
C2438 commonsourceibias.n524 gnd 0.009605f
C2439 commonsourceibias.t74 gnd 0.17946f
C2440 commonsourceibias.n525 gnd 0.008208f
C2441 commonsourceibias.n526 gnd 0.009605f
C2442 commonsourceibias.t62 gnd 0.17946f
C2443 commonsourceibias.n527 gnd 0.011208f
C2444 commonsourceibias.t76 gnd 0.199526f
C2445 commonsourceibias.t16 gnd 0.17946f
C2446 commonsourceibias.n528 gnd 0.078221f
C2447 commonsourceibias.n529 gnd 0.085838f
C2448 commonsourceibias.n530 gnd 0.03983f
C2449 commonsourceibias.n531 gnd 0.009605f
C2450 commonsourceibias.n532 gnd 0.009349f
C2451 commonsourceibias.n533 gnd 0.013398f
C2452 commonsourceibias.n534 gnd 0.071604f
C2453 commonsourceibias.n535 gnd 0.013389f
C2454 commonsourceibias.n536 gnd 0.009605f
C2455 commonsourceibias.n537 gnd 0.009605f
C2456 commonsourceibias.n538 gnd 0.009605f
C2457 commonsourceibias.n539 gnd 0.012358f
C2458 commonsourceibias.n540 gnd 0.071604f
C2459 commonsourceibias.n541 gnd 0.012648f
C2460 commonsourceibias.t48 gnd 0.17946f
C2461 commonsourceibias.n542 gnd 0.071604f
C2462 commonsourceibias.n543 gnd 0.012288f
C2463 commonsourceibias.n544 gnd 0.009605f
C2464 commonsourceibias.n545 gnd 0.009605f
C2465 commonsourceibias.n546 gnd 0.009605f
C2466 commonsourceibias.n547 gnd 0.009057f
C2467 commonsourceibias.n548 gnd 0.01341f
C2468 commonsourceibias.n549 gnd 0.071604f
C2469 commonsourceibias.n550 gnd 0.013406f
C2470 commonsourceibias.n551 gnd 0.009605f
C2471 commonsourceibias.n552 gnd 0.009605f
C2472 commonsourceibias.n553 gnd 0.009605f
C2473 commonsourceibias.n554 gnd 0.012174f
C2474 commonsourceibias.n555 gnd 0.071604f
C2475 commonsourceibias.n556 gnd 0.012558f
C2476 commonsourceibias.t56 gnd 0.17946f
C2477 commonsourceibias.n557 gnd 0.071604f
C2478 commonsourceibias.n558 gnd 0.012378f
C2479 commonsourceibias.n559 gnd 0.009605f
C2480 commonsourceibias.n560 gnd 0.009605f
C2481 commonsourceibias.n561 gnd 0.009605f
C2482 commonsourceibias.n562 gnd 0.008798f
C2483 commonsourceibias.n563 gnd 0.013415f
C2484 commonsourceibias.n564 gnd 0.071604f
C2485 commonsourceibias.n565 gnd 0.013414f
C2486 commonsourceibias.n566 gnd 0.009605f
C2487 commonsourceibias.n567 gnd 0.009605f
C2488 commonsourceibias.n568 gnd 0.009605f
C2489 commonsourceibias.n569 gnd 0.01197f
C2490 commonsourceibias.n570 gnd 0.071604f
C2491 commonsourceibias.n571 gnd 0.012468f
C2492 commonsourceibias.t34 gnd 0.17946f
C2493 commonsourceibias.n572 gnd 0.071604f
C2494 commonsourceibias.n573 gnd 0.012468f
C2495 commonsourceibias.n574 gnd 0.009605f
C2496 commonsourceibias.n575 gnd 0.009605f
C2497 commonsourceibias.n576 gnd 0.009605f
C2498 commonsourceibias.n577 gnd 0.008571f
C2499 commonsourceibias.n578 gnd 0.013414f
C2500 commonsourceibias.n579 gnd 0.071604f
C2501 commonsourceibias.n580 gnd 0.013415f
C2502 commonsourceibias.n581 gnd 0.009605f
C2503 commonsourceibias.n582 gnd 0.009605f
C2504 commonsourceibias.n583 gnd 0.009605f
C2505 commonsourceibias.n584 gnd 0.011742f
C2506 commonsourceibias.n585 gnd 0.071604f
C2507 commonsourceibias.n586 gnd 0.012378f
C2508 commonsourceibias.t8 gnd 0.17946f
C2509 commonsourceibias.n587 gnd 0.071604f
C2510 commonsourceibias.n588 gnd 0.012558f
C2511 commonsourceibias.n589 gnd 0.009605f
C2512 commonsourceibias.n590 gnd 0.009605f
C2513 commonsourceibias.n591 gnd 0.009605f
C2514 commonsourceibias.n592 gnd 0.008375f
C2515 commonsourceibias.n593 gnd 0.013406f
C2516 commonsourceibias.n594 gnd 0.071604f
C2517 commonsourceibias.n595 gnd 0.01341f
C2518 commonsourceibias.n596 gnd 0.009605f
C2519 commonsourceibias.n597 gnd 0.009605f
C2520 commonsourceibias.n598 gnd 0.009605f
C2521 commonsourceibias.n599 gnd 0.011489f
C2522 commonsourceibias.n600 gnd 0.071604f
C2523 commonsourceibias.n601 gnd 0.012288f
C2524 commonsourceibias.t38 gnd 0.17946f
C2525 commonsourceibias.n602 gnd 0.071604f
C2526 commonsourceibias.n603 gnd 0.012648f
C2527 commonsourceibias.n604 gnd 0.009605f
C2528 commonsourceibias.n605 gnd 0.009605f
C2529 commonsourceibias.n606 gnd 0.009605f
C2530 commonsourceibias.n607 gnd 0.008208f
C2531 commonsourceibias.n608 gnd 0.013389f
C2532 commonsourceibias.n609 gnd 0.071604f
C2533 commonsourceibias.n610 gnd 0.013398f
C2534 commonsourceibias.n611 gnd 0.009605f
C2535 commonsourceibias.n612 gnd 0.009605f
C2536 commonsourceibias.n613 gnd 0.009605f
C2537 commonsourceibias.n614 gnd 0.011208f
C2538 commonsourceibias.n615 gnd 0.071604f
C2539 commonsourceibias.n616 gnd 0.011785f
C2540 commonsourceibias.t40 gnd 0.194086f
C2541 commonsourceibias.n617 gnd 0.085919f
C2542 commonsourceibias.n618 gnd 0.095702f
C2543 commonsourceibias.t1 gnd 0.020728f
C2544 commonsourceibias.t41 gnd 0.020728f
C2545 commonsourceibias.n619 gnd 0.183157f
C2546 commonsourceibias.n620 gnd 0.158432f
C2547 commonsourceibias.t39 gnd 0.020728f
C2548 commonsourceibias.t21 gnd 0.020728f
C2549 commonsourceibias.n621 gnd 0.183157f
C2550 commonsourceibias.n622 gnd 0.084131f
C2551 commonsourceibias.t45 gnd 0.020728f
C2552 commonsourceibias.t33 gnd 0.020728f
C2553 commonsourceibias.n623 gnd 0.183157f
C2554 commonsourceibias.n624 gnd 0.084131f
C2555 commonsourceibias.t53 gnd 0.020728f
C2556 commonsourceibias.t9 gnd 0.020728f
C2557 commonsourceibias.n625 gnd 0.183157f
C2558 commonsourceibias.n626 gnd 0.084131f
C2559 commonsourceibias.t35 gnd 0.020728f
C2560 commonsourceibias.t37 gnd 0.020728f
C2561 commonsourceibias.n627 gnd 0.183157f
C2562 commonsourceibias.n628 gnd 0.070287f
C2563 commonsourceibias.n629 gnd 0.085111f
C2564 commonsourceibias.n630 gnd 0.062167f
C2565 commonsourceibias.t102 gnd 0.17946f
C2566 commonsourceibias.n631 gnd 0.071604f
C2567 commonsourceibias.n632 gnd 0.009605f
C2568 commonsourceibias.t188 gnd 0.17946f
C2569 commonsourceibias.n633 gnd 0.071604f
C2570 commonsourceibias.n634 gnd 0.009605f
C2571 commonsourceibias.t162 gnd 0.17946f
C2572 commonsourceibias.n635 gnd 0.071604f
C2573 commonsourceibias.n636 gnd 0.009605f
C2574 commonsourceibias.t103 gnd 0.17946f
C2575 commonsourceibias.n637 gnd 0.008375f
C2576 commonsourceibias.n638 gnd 0.009605f
C2577 commonsourceibias.t166 gnd 0.17946f
C2578 commonsourceibias.n639 gnd 0.011489f
C2579 commonsourceibias.n640 gnd 0.009605f
C2580 commonsourceibias.t185 gnd 0.17946f
C2581 commonsourceibias.n641 gnd 0.008208f
C2582 commonsourceibias.n642 gnd 0.009605f
C2583 commonsourceibias.t160 gnd 0.17946f
C2584 commonsourceibias.n643 gnd 0.011208f
C2585 commonsourceibias.t177 gnd 0.199526f
C2586 commonsourceibias.t159 gnd 0.17946f
C2587 commonsourceibias.n644 gnd 0.078221f
C2588 commonsourceibias.n645 gnd 0.085838f
C2589 commonsourceibias.n646 gnd 0.03983f
C2590 commonsourceibias.n647 gnd 0.009605f
C2591 commonsourceibias.n648 gnd 0.009349f
C2592 commonsourceibias.n649 gnd 0.013398f
C2593 commonsourceibias.n650 gnd 0.071604f
C2594 commonsourceibias.n651 gnd 0.013389f
C2595 commonsourceibias.n652 gnd 0.009605f
C2596 commonsourceibias.n653 gnd 0.009605f
C2597 commonsourceibias.n654 gnd 0.009605f
C2598 commonsourceibias.n655 gnd 0.012358f
C2599 commonsourceibias.n656 gnd 0.071604f
C2600 commonsourceibias.n657 gnd 0.012648f
C2601 commonsourceibias.t135 gnd 0.17946f
C2602 commonsourceibias.n658 gnd 0.071604f
C2603 commonsourceibias.n659 gnd 0.012288f
C2604 commonsourceibias.n660 gnd 0.009605f
C2605 commonsourceibias.n661 gnd 0.009605f
C2606 commonsourceibias.n662 gnd 0.009605f
C2607 commonsourceibias.n663 gnd 0.009057f
C2608 commonsourceibias.n664 gnd 0.01341f
C2609 commonsourceibias.n665 gnd 0.071604f
C2610 commonsourceibias.n666 gnd 0.013406f
C2611 commonsourceibias.n667 gnd 0.009605f
C2612 commonsourceibias.n668 gnd 0.009605f
C2613 commonsourceibias.n669 gnd 0.009605f
C2614 commonsourceibias.n670 gnd 0.012174f
C2615 commonsourceibias.n671 gnd 0.071604f
C2616 commonsourceibias.n672 gnd 0.012558f
C2617 commonsourceibias.n673 gnd 0.012378f
C2618 commonsourceibias.n674 gnd 0.009605f
C2619 commonsourceibias.n675 gnd 0.009605f
C2620 commonsourceibias.n676 gnd 0.011742f
C2621 commonsourceibias.n677 gnd 0.008798f
C2622 commonsourceibias.n678 gnd 0.013415f
C2623 commonsourceibias.n679 gnd 0.009605f
C2624 commonsourceibias.n680 gnd 0.009605f
C2625 commonsourceibias.n681 gnd 0.013414f
C2626 commonsourceibias.n682 gnd 0.008571f
C2627 commonsourceibias.n683 gnd 0.01197f
C2628 commonsourceibias.n684 gnd 0.009605f
C2629 commonsourceibias.n685 gnd 0.008391f
C2630 commonsourceibias.n686 gnd 0.012468f
C2631 commonsourceibias.t174 gnd 0.17946f
C2632 commonsourceibias.n687 gnd 0.071604f
C2633 commonsourceibias.n688 gnd 0.012468f
C2634 commonsourceibias.n689 gnd 0.008391f
C2635 commonsourceibias.n690 gnd 0.009605f
C2636 commonsourceibias.n691 gnd 0.009605f
C2637 commonsourceibias.n692 gnd 0.008571f
C2638 commonsourceibias.n693 gnd 0.013414f
C2639 commonsourceibias.n694 gnd 0.071604f
C2640 commonsourceibias.n695 gnd 0.013415f
C2641 commonsourceibias.n696 gnd 0.009605f
C2642 commonsourceibias.n697 gnd 0.009605f
C2643 commonsourceibias.n698 gnd 0.009605f
C2644 commonsourceibias.n699 gnd 0.011742f
C2645 commonsourceibias.n700 gnd 0.071604f
C2646 commonsourceibias.n701 gnd 0.012378f
C2647 commonsourceibias.t90 gnd 0.17946f
C2648 commonsourceibias.n702 gnd 0.071604f
C2649 commonsourceibias.n703 gnd 0.012558f
C2650 commonsourceibias.n704 gnd 0.009605f
C2651 commonsourceibias.n705 gnd 0.009605f
C2652 commonsourceibias.n706 gnd 0.009605f
C2653 commonsourceibias.n707 gnd 0.008375f
C2654 commonsourceibias.n708 gnd 0.013406f
C2655 commonsourceibias.n709 gnd 0.071604f
C2656 commonsourceibias.n710 gnd 0.01341f
C2657 commonsourceibias.n711 gnd 0.009605f
C2658 commonsourceibias.n712 gnd 0.009605f
C2659 commonsourceibias.n713 gnd 0.009605f
C2660 commonsourceibias.n714 gnd 0.011489f
C2661 commonsourceibias.n715 gnd 0.071604f
C2662 commonsourceibias.n716 gnd 0.012288f
C2663 commonsourceibias.t116 gnd 0.17946f
C2664 commonsourceibias.n717 gnd 0.071604f
C2665 commonsourceibias.n718 gnd 0.012648f
C2666 commonsourceibias.n719 gnd 0.009605f
C2667 commonsourceibias.n720 gnd 0.009605f
C2668 commonsourceibias.n721 gnd 0.009605f
C2669 commonsourceibias.n722 gnd 0.008208f
C2670 commonsourceibias.n723 gnd 0.013389f
C2671 commonsourceibias.n724 gnd 0.071604f
C2672 commonsourceibias.n725 gnd 0.013398f
C2673 commonsourceibias.n726 gnd 0.009605f
C2674 commonsourceibias.n727 gnd 0.009605f
C2675 commonsourceibias.n728 gnd 0.009605f
C2676 commonsourceibias.n729 gnd 0.011208f
C2677 commonsourceibias.n730 gnd 0.071604f
C2678 commonsourceibias.n731 gnd 0.011785f
C2679 commonsourceibias.n732 gnd 0.085919f
C2680 commonsourceibias.n733 gnd 0.056156f
C2681 commonsourceibias.n734 gnd 0.012817f
C2682 commonsourceibias.t180 gnd 0.17946f
C2683 commonsourceibias.n735 gnd 0.009349f
C2684 commonsourceibias.n736 gnd 0.009605f
C2685 commonsourceibias.t82 gnd 0.17946f
C2686 commonsourceibias.n737 gnd 0.012358f
C2687 commonsourceibias.n738 gnd 0.009605f
C2688 commonsourceibias.t179 gnd 0.17946f
C2689 commonsourceibias.n739 gnd 0.009057f
C2690 commonsourceibias.n740 gnd 0.009605f
C2691 commonsourceibias.t81 gnd 0.17946f
C2692 commonsourceibias.n741 gnd 0.012174f
C2693 commonsourceibias.n742 gnd 0.009605f
C2694 commonsourceibias.t178 gnd 0.17946f
C2695 commonsourceibias.n743 gnd 0.008798f
C2696 commonsourceibias.n744 gnd 0.009605f
C2697 commonsourceibias.t89 gnd 0.17946f
C2698 commonsourceibias.n745 gnd 0.01197f
C2699 commonsourceibias.n746 gnd 0.009605f
C2700 commonsourceibias.t97 gnd 0.17946f
C2701 commonsourceibias.n747 gnd 0.008571f
C2702 commonsourceibias.n748 gnd 0.009605f
C2703 commonsourceibias.t86 gnd 0.17946f
C2704 commonsourceibias.n749 gnd 0.011742f
C2705 commonsourceibias.n750 gnd 0.009605f
C2706 commonsourceibias.t106 gnd 0.17946f
C2707 commonsourceibias.n751 gnd 0.008375f
C2708 commonsourceibias.n752 gnd 0.009605f
C2709 commonsourceibias.t85 gnd 0.17946f
C2710 commonsourceibias.n753 gnd 0.011489f
C2711 commonsourceibias.n754 gnd 0.009605f
C2712 commonsourceibias.t104 gnd 0.17946f
C2713 commonsourceibias.n755 gnd 0.008208f
C2714 commonsourceibias.n756 gnd 0.009605f
C2715 commonsourceibias.t132 gnd 0.17946f
C2716 commonsourceibias.n757 gnd 0.011208f
C2717 commonsourceibias.t98 gnd 0.199526f
C2718 commonsourceibias.t123 gnd 0.17946f
C2719 commonsourceibias.n758 gnd 0.078221f
C2720 commonsourceibias.n759 gnd 0.085838f
C2721 commonsourceibias.n760 gnd 0.03983f
C2722 commonsourceibias.n761 gnd 0.009605f
C2723 commonsourceibias.n762 gnd 0.009349f
C2724 commonsourceibias.n763 gnd 0.013398f
C2725 commonsourceibias.n764 gnd 0.071604f
C2726 commonsourceibias.n765 gnd 0.013389f
C2727 commonsourceibias.n766 gnd 0.009605f
C2728 commonsourceibias.n767 gnd 0.009605f
C2729 commonsourceibias.n768 gnd 0.009605f
C2730 commonsourceibias.n769 gnd 0.012358f
C2731 commonsourceibias.n770 gnd 0.071604f
C2732 commonsourceibias.n771 gnd 0.012648f
C2733 commonsourceibias.t118 gnd 0.17946f
C2734 commonsourceibias.n772 gnd 0.071604f
C2735 commonsourceibias.n773 gnd 0.012288f
C2736 commonsourceibias.n774 gnd 0.009605f
C2737 commonsourceibias.n775 gnd 0.009605f
C2738 commonsourceibias.n776 gnd 0.009605f
C2739 commonsourceibias.n777 gnd 0.009057f
C2740 commonsourceibias.n778 gnd 0.01341f
C2741 commonsourceibias.n779 gnd 0.071604f
C2742 commonsourceibias.n780 gnd 0.013406f
C2743 commonsourceibias.n781 gnd 0.009605f
C2744 commonsourceibias.n782 gnd 0.009605f
C2745 commonsourceibias.n783 gnd 0.009605f
C2746 commonsourceibias.n784 gnd 0.012174f
C2747 commonsourceibias.n785 gnd 0.071604f
C2748 commonsourceibias.n786 gnd 0.012558f
C2749 commonsourceibias.t119 gnd 0.17946f
C2750 commonsourceibias.n787 gnd 0.071604f
C2751 commonsourceibias.n788 gnd 0.012378f
C2752 commonsourceibias.n789 gnd 0.009605f
C2753 commonsourceibias.n790 gnd 0.009605f
C2754 commonsourceibias.n791 gnd 0.009605f
C2755 commonsourceibias.n792 gnd 0.008798f
C2756 commonsourceibias.n793 gnd 0.013415f
C2757 commonsourceibias.n794 gnd 0.071604f
C2758 commonsourceibias.n795 gnd 0.013414f
C2759 commonsourceibias.n796 gnd 0.009605f
C2760 commonsourceibias.n797 gnd 0.009605f
C2761 commonsourceibias.n798 gnd 0.009605f
C2762 commonsourceibias.n799 gnd 0.01197f
C2763 commonsourceibias.n800 gnd 0.071604f
C2764 commonsourceibias.n801 gnd 0.012468f
C2765 commonsourceibias.t120 gnd 0.17946f
C2766 commonsourceibias.n802 gnd 0.071604f
C2767 commonsourceibias.n803 gnd 0.012468f
C2768 commonsourceibias.n804 gnd 0.009605f
C2769 commonsourceibias.n805 gnd 0.009605f
C2770 commonsourceibias.n806 gnd 0.009605f
C2771 commonsourceibias.n807 gnd 0.008571f
C2772 commonsourceibias.n808 gnd 0.013414f
C2773 commonsourceibias.n809 gnd 0.071604f
C2774 commonsourceibias.n810 gnd 0.013415f
C2775 commonsourceibias.n811 gnd 0.009605f
C2776 commonsourceibias.n812 gnd 0.009605f
C2777 commonsourceibias.n813 gnd 0.009605f
C2778 commonsourceibias.n814 gnd 0.011742f
C2779 commonsourceibias.n815 gnd 0.071604f
C2780 commonsourceibias.n816 gnd 0.012378f
C2781 commonsourceibias.t121 gnd 0.17946f
C2782 commonsourceibias.n817 gnd 0.071604f
C2783 commonsourceibias.n818 gnd 0.012558f
C2784 commonsourceibias.n819 gnd 0.009605f
C2785 commonsourceibias.n820 gnd 0.009605f
C2786 commonsourceibias.n821 gnd 0.009605f
C2787 commonsourceibias.n822 gnd 0.008375f
C2788 commonsourceibias.n823 gnd 0.013406f
C2789 commonsourceibias.n824 gnd 0.071604f
C2790 commonsourceibias.n825 gnd 0.01341f
C2791 commonsourceibias.n826 gnd 0.009605f
C2792 commonsourceibias.n827 gnd 0.009605f
C2793 commonsourceibias.n828 gnd 0.009605f
C2794 commonsourceibias.n829 gnd 0.011489f
C2795 commonsourceibias.n830 gnd 0.071604f
C2796 commonsourceibias.n831 gnd 0.012288f
C2797 commonsourceibias.t193 gnd 0.17946f
C2798 commonsourceibias.n832 gnd 0.071604f
C2799 commonsourceibias.n833 gnd 0.012648f
C2800 commonsourceibias.n834 gnd 0.009605f
C2801 commonsourceibias.n835 gnd 0.009605f
C2802 commonsourceibias.n836 gnd 0.009605f
C2803 commonsourceibias.n837 gnd 0.008208f
C2804 commonsourceibias.n838 gnd 0.013389f
C2805 commonsourceibias.n839 gnd 0.071604f
C2806 commonsourceibias.n840 gnd 0.013398f
C2807 commonsourceibias.n841 gnd 0.009605f
C2808 commonsourceibias.n842 gnd 0.009605f
C2809 commonsourceibias.n843 gnd 0.009605f
C2810 commonsourceibias.n844 gnd 0.011208f
C2811 commonsourceibias.n845 gnd 0.071604f
C2812 commonsourceibias.n846 gnd 0.011785f
C2813 commonsourceibias.t189 gnd 0.194086f
C2814 commonsourceibias.n847 gnd 0.085919f
C2815 commonsourceibias.n848 gnd 0.029883f
C2816 commonsourceibias.n849 gnd 0.153509f
C2817 commonsourceibias.n850 gnd 0.012817f
C2818 commonsourceibias.t133 gnd 0.17946f
C2819 commonsourceibias.n851 gnd 0.009349f
C2820 commonsourceibias.n852 gnd 0.009605f
C2821 commonsourceibias.t153 gnd 0.17946f
C2822 commonsourceibias.n853 gnd 0.012358f
C2823 commonsourceibias.n854 gnd 0.009605f
C2824 commonsourceibias.t122 gnd 0.17946f
C2825 commonsourceibias.n855 gnd 0.009057f
C2826 commonsourceibias.n856 gnd 0.009605f
C2827 commonsourceibias.t143 gnd 0.17946f
C2828 commonsourceibias.n857 gnd 0.012174f
C2829 commonsourceibias.n858 gnd 0.009605f
C2830 commonsourceibias.t99 gnd 0.17946f
C2831 commonsourceibias.n859 gnd 0.008798f
C2832 commonsourceibias.n860 gnd 0.009605f
C2833 commonsourceibias.t87 gnd 0.17946f
C2834 commonsourceibias.n861 gnd 0.01197f
C2835 commonsourceibias.n862 gnd 0.009605f
C2836 commonsourceibias.t167 gnd 0.17946f
C2837 commonsourceibias.n863 gnd 0.008571f
C2838 commonsourceibias.n864 gnd 0.009605f
C2839 commonsourceibias.t192 gnd 0.17946f
C2840 commonsourceibias.n865 gnd 0.011742f
C2841 commonsourceibias.n866 gnd 0.009605f
C2842 commonsourceibias.t136 gnd 0.17946f
C2843 commonsourceibias.n867 gnd 0.008375f
C2844 commonsourceibias.n868 gnd 0.009605f
C2845 commonsourceibias.t181 gnd 0.17946f
C2846 commonsourceibias.n869 gnd 0.011489f
C2847 commonsourceibias.n870 gnd 0.009605f
C2848 commonsourceibias.t126 gnd 0.17946f
C2849 commonsourceibias.n871 gnd 0.008208f
C2850 commonsourceibias.n872 gnd 0.009605f
C2851 commonsourceibias.t146 gnd 0.17946f
C2852 commonsourceibias.n873 gnd 0.011208f
C2853 commonsourceibias.t191 gnd 0.199526f
C2854 commonsourceibias.t156 gnd 0.17946f
C2855 commonsourceibias.n874 gnd 0.078221f
C2856 commonsourceibias.n875 gnd 0.085838f
C2857 commonsourceibias.n876 gnd 0.03983f
C2858 commonsourceibias.n877 gnd 0.009605f
C2859 commonsourceibias.n878 gnd 0.009349f
C2860 commonsourceibias.n879 gnd 0.013398f
C2861 commonsourceibias.n880 gnd 0.071604f
C2862 commonsourceibias.n881 gnd 0.013389f
C2863 commonsourceibias.n882 gnd 0.009605f
C2864 commonsourceibias.n883 gnd 0.009605f
C2865 commonsourceibias.n884 gnd 0.009605f
C2866 commonsourceibias.n885 gnd 0.012358f
C2867 commonsourceibias.n886 gnd 0.071604f
C2868 commonsourceibias.n887 gnd 0.012648f
C2869 commonsourceibias.t91 gnd 0.17946f
C2870 commonsourceibias.n888 gnd 0.071604f
C2871 commonsourceibias.n889 gnd 0.012288f
C2872 commonsourceibias.n890 gnd 0.009605f
C2873 commonsourceibias.n891 gnd 0.009605f
C2874 commonsourceibias.n892 gnd 0.009605f
C2875 commonsourceibias.n893 gnd 0.009057f
C2876 commonsourceibias.n894 gnd 0.01341f
C2877 commonsourceibias.n895 gnd 0.071604f
C2878 commonsourceibias.n896 gnd 0.013406f
C2879 commonsourceibias.n897 gnd 0.009605f
C2880 commonsourceibias.n898 gnd 0.009605f
C2881 commonsourceibias.n899 gnd 0.009605f
C2882 commonsourceibias.n900 gnd 0.012174f
C2883 commonsourceibias.n901 gnd 0.071604f
C2884 commonsourceibias.n902 gnd 0.012558f
C2885 commonsourceibias.t107 gnd 0.17946f
C2886 commonsourceibias.n903 gnd 0.071604f
C2887 commonsourceibias.n904 gnd 0.012378f
C2888 commonsourceibias.n905 gnd 0.009605f
C2889 commonsourceibias.n906 gnd 0.009605f
C2890 commonsourceibias.n907 gnd 0.009605f
C2891 commonsourceibias.n908 gnd 0.008798f
C2892 commonsourceibias.n909 gnd 0.013415f
C2893 commonsourceibias.n910 gnd 0.071604f
C2894 commonsourceibias.n911 gnd 0.013414f
C2895 commonsourceibias.n912 gnd 0.009605f
C2896 commonsourceibias.n913 gnd 0.009605f
C2897 commonsourceibias.n914 gnd 0.009605f
C2898 commonsourceibias.n915 gnd 0.01197f
C2899 commonsourceibias.n916 gnd 0.071604f
C2900 commonsourceibias.n917 gnd 0.012468f
C2901 commonsourceibias.t127 gnd 0.17946f
C2902 commonsourceibias.n918 gnd 0.071604f
C2903 commonsourceibias.n919 gnd 0.012468f
C2904 commonsourceibias.n920 gnd 0.009605f
C2905 commonsourceibias.n921 gnd 0.009605f
C2906 commonsourceibias.n922 gnd 0.009605f
C2907 commonsourceibias.n923 gnd 0.008571f
C2908 commonsourceibias.n924 gnd 0.013414f
C2909 commonsourceibias.n925 gnd 0.071604f
C2910 commonsourceibias.n926 gnd 0.013415f
C2911 commonsourceibias.n927 gnd 0.009605f
C2912 commonsourceibias.n928 gnd 0.009605f
C2913 commonsourceibias.n929 gnd 0.009605f
C2914 commonsourceibias.n930 gnd 0.011742f
C2915 commonsourceibias.n931 gnd 0.071604f
C2916 commonsourceibias.n932 gnd 0.012378f
C2917 commonsourceibias.t137 gnd 0.17946f
C2918 commonsourceibias.n933 gnd 0.071604f
C2919 commonsourceibias.n934 gnd 0.012558f
C2920 commonsourceibias.n935 gnd 0.009605f
C2921 commonsourceibias.n936 gnd 0.009605f
C2922 commonsourceibias.n937 gnd 0.009605f
C2923 commonsourceibias.n938 gnd 0.008375f
C2924 commonsourceibias.n939 gnd 0.013406f
C2925 commonsourceibias.n940 gnd 0.071604f
C2926 commonsourceibias.n941 gnd 0.01341f
C2927 commonsourceibias.n942 gnd 0.009605f
C2928 commonsourceibias.n943 gnd 0.009605f
C2929 commonsourceibias.n944 gnd 0.009605f
C2930 commonsourceibias.n945 gnd 0.011489f
C2931 commonsourceibias.n946 gnd 0.071604f
C2932 commonsourceibias.n947 gnd 0.012288f
C2933 commonsourceibias.t170 gnd 0.17946f
C2934 commonsourceibias.n948 gnd 0.071604f
C2935 commonsourceibias.n949 gnd 0.012648f
C2936 commonsourceibias.n950 gnd 0.009605f
C2937 commonsourceibias.n951 gnd 0.009605f
C2938 commonsourceibias.n952 gnd 0.009605f
C2939 commonsourceibias.n953 gnd 0.008208f
C2940 commonsourceibias.n954 gnd 0.013389f
C2941 commonsourceibias.n955 gnd 0.071604f
C2942 commonsourceibias.n956 gnd 0.013398f
C2943 commonsourceibias.n957 gnd 0.009605f
C2944 commonsourceibias.n958 gnd 0.009605f
C2945 commonsourceibias.n959 gnd 0.009605f
C2946 commonsourceibias.n960 gnd 0.011208f
C2947 commonsourceibias.n961 gnd 0.071604f
C2948 commonsourceibias.n962 gnd 0.011785f
C2949 commonsourceibias.t101 gnd 0.194086f
C2950 commonsourceibias.n963 gnd 0.085919f
C2951 commonsourceibias.n964 gnd 0.029883f
C2952 commonsourceibias.n965 gnd 0.202572f
C2953 commonsourceibias.n966 gnd 5.28148f
C2954 vdd.t238 gnd 0.034846f
C2955 vdd.t218 gnd 0.034846f
C2956 vdd.n0 gnd 0.274839f
C2957 vdd.t197 gnd 0.034846f
C2958 vdd.t234 gnd 0.034846f
C2959 vdd.n1 gnd 0.274385f
C2960 vdd.n2 gnd 0.253035f
C2961 vdd.t215 gnd 0.034846f
C2962 vdd.t245 gnd 0.034846f
C2963 vdd.n3 gnd 0.274385f
C2964 vdd.n4 gnd 0.127969f
C2965 vdd.t243 gnd 0.034846f
C2966 vdd.t223 gnd 0.034846f
C2967 vdd.n5 gnd 0.274385f
C2968 vdd.n6 gnd 0.120076f
C2969 vdd.t249 gnd 0.034846f
C2970 vdd.t213 gnd 0.034846f
C2971 vdd.n7 gnd 0.274839f
C2972 vdd.t221 gnd 0.034846f
C2973 vdd.t241 gnd 0.034846f
C2974 vdd.n8 gnd 0.274385f
C2975 vdd.n9 gnd 0.253035f
C2976 vdd.t230 gnd 0.034846f
C2977 vdd.t201 gnd 0.034846f
C2978 vdd.n10 gnd 0.274385f
C2979 vdd.n11 gnd 0.127969f
C2980 vdd.t210 gnd 0.034846f
C2981 vdd.t228 gnd 0.034846f
C2982 vdd.n12 gnd 0.274385f
C2983 vdd.n13 gnd 0.120076f
C2984 vdd.n14 gnd 0.084891f
C2985 vdd.t14 gnd 0.019359f
C2986 vdd.t193 gnd 0.019359f
C2987 vdd.n15 gnd 0.178192f
C2988 vdd.t60 gnd 0.019359f
C2989 vdd.t10 gnd 0.019359f
C2990 vdd.n16 gnd 0.177671f
C2991 vdd.n17 gnd 0.309202f
C2992 vdd.t8 gnd 0.019359f
C2993 vdd.t157 gnd 0.019359f
C2994 vdd.n18 gnd 0.177671f
C2995 vdd.n19 gnd 0.127921f
C2996 vdd.t192 gnd 0.019359f
C2997 vdd.t13 gnd 0.019359f
C2998 vdd.n20 gnd 0.178192f
C2999 vdd.t11 gnd 0.019359f
C3000 vdd.t173 gnd 0.019359f
C3001 vdd.n21 gnd 0.177671f
C3002 vdd.n22 gnd 0.309202f
C3003 vdd.t59 gnd 0.019359f
C3004 vdd.t12 gnd 0.019359f
C3005 vdd.n23 gnd 0.177671f
C3006 vdd.n24 gnd 0.127921f
C3007 vdd.t9 gnd 0.019359f
C3008 vdd.t158 gnd 0.019359f
C3009 vdd.n25 gnd 0.177671f
C3010 vdd.t40 gnd 0.019359f
C3011 vdd.t36 gnd 0.019359f
C3012 vdd.n26 gnd 0.177671f
C3013 vdd.n27 gnd 19.6921f
C3014 vdd.n28 gnd 7.906759f
C3015 vdd.n29 gnd 0.00528f
C3016 vdd.n30 gnd 0.0049f
C3017 vdd.n31 gnd 0.00271f
C3018 vdd.n32 gnd 0.006223f
C3019 vdd.n33 gnd 0.002633f
C3020 vdd.n34 gnd 0.002788f
C3021 vdd.n35 gnd 0.0049f
C3022 vdd.n36 gnd 0.002633f
C3023 vdd.n37 gnd 0.006223f
C3024 vdd.n38 gnd 0.002788f
C3025 vdd.n39 gnd 0.0049f
C3026 vdd.n40 gnd 0.002633f
C3027 vdd.n41 gnd 0.004667f
C3028 vdd.n42 gnd 0.004681f
C3029 vdd.t175 gnd 0.01337f
C3030 vdd.n43 gnd 0.029747f
C3031 vdd.n44 gnd 0.154813f
C3032 vdd.n45 gnd 0.002633f
C3033 vdd.n46 gnd 0.002788f
C3034 vdd.n47 gnd 0.006223f
C3035 vdd.n48 gnd 0.006223f
C3036 vdd.n49 gnd 0.002788f
C3037 vdd.n50 gnd 0.002633f
C3038 vdd.n51 gnd 0.0049f
C3039 vdd.n52 gnd 0.0049f
C3040 vdd.n53 gnd 0.002633f
C3041 vdd.n54 gnd 0.002788f
C3042 vdd.n55 gnd 0.006223f
C3043 vdd.n56 gnd 0.006223f
C3044 vdd.n57 gnd 0.002788f
C3045 vdd.n58 gnd 0.002633f
C3046 vdd.n59 gnd 0.0049f
C3047 vdd.n60 gnd 0.0049f
C3048 vdd.n61 gnd 0.002633f
C3049 vdd.n62 gnd 0.002788f
C3050 vdd.n63 gnd 0.006223f
C3051 vdd.n64 gnd 0.006223f
C3052 vdd.n65 gnd 0.014713f
C3053 vdd.n66 gnd 0.00271f
C3054 vdd.n67 gnd 0.002633f
C3055 vdd.n68 gnd 0.012664f
C3056 vdd.n69 gnd 0.008841f
C3057 vdd.t64 gnd 0.030974f
C3058 vdd.t34 gnd 0.030974f
C3059 vdd.n70 gnd 0.212878f
C3060 vdd.n71 gnd 0.167396f
C3061 vdd.t22 gnd 0.030974f
C3062 vdd.t252 gnd 0.030974f
C3063 vdd.n72 gnd 0.212878f
C3064 vdd.n73 gnd 0.135088f
C3065 vdd.t54 gnd 0.030974f
C3066 vdd.t156 gnd 0.030974f
C3067 vdd.n74 gnd 0.212878f
C3068 vdd.n75 gnd 0.135088f
C3069 vdd.t164 gnd 0.030974f
C3070 vdd.t191 gnd 0.030974f
C3071 vdd.n76 gnd 0.212878f
C3072 vdd.n77 gnd 0.135088f
C3073 vdd.t1 gnd 0.030974f
C3074 vdd.t147 gnd 0.030974f
C3075 vdd.n78 gnd 0.212878f
C3076 vdd.n79 gnd 0.135088f
C3077 vdd.t269 gnd 0.030974f
C3078 vdd.t163 gnd 0.030974f
C3079 vdd.n80 gnd 0.212878f
C3080 vdd.n81 gnd 0.135088f
C3081 vdd.t255 gnd 0.030974f
C3082 vdd.t258 gnd 0.030974f
C3083 vdd.n82 gnd 0.212878f
C3084 vdd.n83 gnd 0.135088f
C3085 vdd.n84 gnd 0.00528f
C3086 vdd.n85 gnd 0.0049f
C3087 vdd.n86 gnd 0.00271f
C3088 vdd.n87 gnd 0.006223f
C3089 vdd.n88 gnd 0.002633f
C3090 vdd.n89 gnd 0.002788f
C3091 vdd.n90 gnd 0.0049f
C3092 vdd.n91 gnd 0.002633f
C3093 vdd.n92 gnd 0.006223f
C3094 vdd.n93 gnd 0.002788f
C3095 vdd.n94 gnd 0.0049f
C3096 vdd.n95 gnd 0.002633f
C3097 vdd.n96 gnd 0.004667f
C3098 vdd.n97 gnd 0.004681f
C3099 vdd.t160 gnd 0.01337f
C3100 vdd.n98 gnd 0.029747f
C3101 vdd.n99 gnd 0.154813f
C3102 vdd.n100 gnd 0.002633f
C3103 vdd.n101 gnd 0.002788f
C3104 vdd.n102 gnd 0.006223f
C3105 vdd.n103 gnd 0.006223f
C3106 vdd.n104 gnd 0.002788f
C3107 vdd.n105 gnd 0.002633f
C3108 vdd.n106 gnd 0.0049f
C3109 vdd.n107 gnd 0.0049f
C3110 vdd.n108 gnd 0.002633f
C3111 vdd.n109 gnd 0.002788f
C3112 vdd.n110 gnd 0.006223f
C3113 vdd.n111 gnd 0.006223f
C3114 vdd.n112 gnd 0.002788f
C3115 vdd.n113 gnd 0.002633f
C3116 vdd.n114 gnd 0.0049f
C3117 vdd.n115 gnd 0.0049f
C3118 vdd.n116 gnd 0.002633f
C3119 vdd.n117 gnd 0.002788f
C3120 vdd.n118 gnd 0.006223f
C3121 vdd.n119 gnd 0.006223f
C3122 vdd.n120 gnd 0.014713f
C3123 vdd.n121 gnd 0.00271f
C3124 vdd.n122 gnd 0.002633f
C3125 vdd.n123 gnd 0.012664f
C3126 vdd.n124 gnd 0.008564f
C3127 vdd.n125 gnd 0.100506f
C3128 vdd.n126 gnd 0.00528f
C3129 vdd.n127 gnd 0.0049f
C3130 vdd.n128 gnd 0.00271f
C3131 vdd.n129 gnd 0.006223f
C3132 vdd.n130 gnd 0.002633f
C3133 vdd.n131 gnd 0.002788f
C3134 vdd.n132 gnd 0.0049f
C3135 vdd.n133 gnd 0.002633f
C3136 vdd.n134 gnd 0.006223f
C3137 vdd.n135 gnd 0.002788f
C3138 vdd.n136 gnd 0.0049f
C3139 vdd.n137 gnd 0.002633f
C3140 vdd.n138 gnd 0.004667f
C3141 vdd.n139 gnd 0.004681f
C3142 vdd.t273 gnd 0.01337f
C3143 vdd.n140 gnd 0.029747f
C3144 vdd.n141 gnd 0.154813f
C3145 vdd.n142 gnd 0.002633f
C3146 vdd.n143 gnd 0.002788f
C3147 vdd.n144 gnd 0.006223f
C3148 vdd.n145 gnd 0.006223f
C3149 vdd.n146 gnd 0.002788f
C3150 vdd.n147 gnd 0.002633f
C3151 vdd.n148 gnd 0.0049f
C3152 vdd.n149 gnd 0.0049f
C3153 vdd.n150 gnd 0.002633f
C3154 vdd.n151 gnd 0.002788f
C3155 vdd.n152 gnd 0.006223f
C3156 vdd.n153 gnd 0.006223f
C3157 vdd.n154 gnd 0.002788f
C3158 vdd.n155 gnd 0.002633f
C3159 vdd.n156 gnd 0.0049f
C3160 vdd.n157 gnd 0.0049f
C3161 vdd.n158 gnd 0.002633f
C3162 vdd.n159 gnd 0.002788f
C3163 vdd.n160 gnd 0.006223f
C3164 vdd.n161 gnd 0.006223f
C3165 vdd.n162 gnd 0.014713f
C3166 vdd.n163 gnd 0.00271f
C3167 vdd.n164 gnd 0.002633f
C3168 vdd.n165 gnd 0.012664f
C3169 vdd.n166 gnd 0.008841f
C3170 vdd.t267 gnd 0.030974f
C3171 vdd.t42 gnd 0.030974f
C3172 vdd.n167 gnd 0.212878f
C3173 vdd.n168 gnd 0.167396f
C3174 vdd.t271 gnd 0.030974f
C3175 vdd.t179 gnd 0.030974f
C3176 vdd.n169 gnd 0.212878f
C3177 vdd.n170 gnd 0.135088f
C3178 vdd.t150 gnd 0.030974f
C3179 vdd.t142 gnd 0.030974f
C3180 vdd.n171 gnd 0.212878f
C3181 vdd.n172 gnd 0.135088f
C3182 vdd.t153 gnd 0.030974f
C3183 vdd.t170 gnd 0.030974f
C3184 vdd.n173 gnd 0.212878f
C3185 vdd.n174 gnd 0.135088f
C3186 vdd.t39 gnd 0.030974f
C3187 vdd.t154 gnd 0.030974f
C3188 vdd.n175 gnd 0.212878f
C3189 vdd.n176 gnd 0.135088f
C3190 vdd.t7 gnd 0.030974f
C3191 vdd.t262 gnd 0.030974f
C3192 vdd.n177 gnd 0.212878f
C3193 vdd.n178 gnd 0.135088f
C3194 vdd.t188 gnd 0.030974f
C3195 vdd.t272 gnd 0.030974f
C3196 vdd.n179 gnd 0.212878f
C3197 vdd.n180 gnd 0.135088f
C3198 vdd.n181 gnd 0.00528f
C3199 vdd.n182 gnd 0.0049f
C3200 vdd.n183 gnd 0.00271f
C3201 vdd.n184 gnd 0.006223f
C3202 vdd.n185 gnd 0.002633f
C3203 vdd.n186 gnd 0.002788f
C3204 vdd.n187 gnd 0.0049f
C3205 vdd.n188 gnd 0.002633f
C3206 vdd.n189 gnd 0.006223f
C3207 vdd.n190 gnd 0.002788f
C3208 vdd.n191 gnd 0.0049f
C3209 vdd.n192 gnd 0.002633f
C3210 vdd.n193 gnd 0.004667f
C3211 vdd.n194 gnd 0.004681f
C3212 vdd.t148 gnd 0.01337f
C3213 vdd.n195 gnd 0.029747f
C3214 vdd.n196 gnd 0.154813f
C3215 vdd.n197 gnd 0.002633f
C3216 vdd.n198 gnd 0.002788f
C3217 vdd.n199 gnd 0.006223f
C3218 vdd.n200 gnd 0.006223f
C3219 vdd.n201 gnd 0.002788f
C3220 vdd.n202 gnd 0.002633f
C3221 vdd.n203 gnd 0.0049f
C3222 vdd.n204 gnd 0.0049f
C3223 vdd.n205 gnd 0.002633f
C3224 vdd.n206 gnd 0.002788f
C3225 vdd.n207 gnd 0.006223f
C3226 vdd.n208 gnd 0.006223f
C3227 vdd.n209 gnd 0.002788f
C3228 vdd.n210 gnd 0.002633f
C3229 vdd.n211 gnd 0.0049f
C3230 vdd.n212 gnd 0.0049f
C3231 vdd.n213 gnd 0.002633f
C3232 vdd.n214 gnd 0.002788f
C3233 vdd.n215 gnd 0.006223f
C3234 vdd.n216 gnd 0.006223f
C3235 vdd.n217 gnd 0.014713f
C3236 vdd.n218 gnd 0.00271f
C3237 vdd.n219 gnd 0.002633f
C3238 vdd.n220 gnd 0.012664f
C3239 vdd.n221 gnd 0.008564f
C3240 vdd.n222 gnd 0.059791f
C3241 vdd.n223 gnd 0.215442f
C3242 vdd.n224 gnd 0.00528f
C3243 vdd.n225 gnd 0.0049f
C3244 vdd.n226 gnd 0.00271f
C3245 vdd.n227 gnd 0.006223f
C3246 vdd.n228 gnd 0.002633f
C3247 vdd.n229 gnd 0.002788f
C3248 vdd.n230 gnd 0.0049f
C3249 vdd.n231 gnd 0.002633f
C3250 vdd.n232 gnd 0.006223f
C3251 vdd.n233 gnd 0.002788f
C3252 vdd.n234 gnd 0.0049f
C3253 vdd.n235 gnd 0.002633f
C3254 vdd.n236 gnd 0.004667f
C3255 vdd.n237 gnd 0.004681f
C3256 vdd.t52 gnd 0.01337f
C3257 vdd.n238 gnd 0.029747f
C3258 vdd.n239 gnd 0.154813f
C3259 vdd.n240 gnd 0.002633f
C3260 vdd.n241 gnd 0.002788f
C3261 vdd.n242 gnd 0.006223f
C3262 vdd.n243 gnd 0.006223f
C3263 vdd.n244 gnd 0.002788f
C3264 vdd.n245 gnd 0.002633f
C3265 vdd.n246 gnd 0.0049f
C3266 vdd.n247 gnd 0.0049f
C3267 vdd.n248 gnd 0.002633f
C3268 vdd.n249 gnd 0.002788f
C3269 vdd.n250 gnd 0.006223f
C3270 vdd.n251 gnd 0.006223f
C3271 vdd.n252 gnd 0.002788f
C3272 vdd.n253 gnd 0.002633f
C3273 vdd.n254 gnd 0.0049f
C3274 vdd.n255 gnd 0.0049f
C3275 vdd.n256 gnd 0.002633f
C3276 vdd.n257 gnd 0.002788f
C3277 vdd.n258 gnd 0.006223f
C3278 vdd.n259 gnd 0.006223f
C3279 vdd.n260 gnd 0.014713f
C3280 vdd.n261 gnd 0.00271f
C3281 vdd.n262 gnd 0.002633f
C3282 vdd.n263 gnd 0.012664f
C3283 vdd.n264 gnd 0.008841f
C3284 vdd.t259 gnd 0.030974f
C3285 vdd.t263 gnd 0.030974f
C3286 vdd.n265 gnd 0.212878f
C3287 vdd.n266 gnd 0.167396f
C3288 vdd.t35 gnd 0.030974f
C3289 vdd.t172 gnd 0.030974f
C3290 vdd.n267 gnd 0.212878f
C3291 vdd.n268 gnd 0.135088f
C3292 vdd.t275 gnd 0.030974f
C3293 vdd.t159 gnd 0.030974f
C3294 vdd.n269 gnd 0.212878f
C3295 vdd.n270 gnd 0.135088f
C3296 vdd.t155 gnd 0.030974f
C3297 vdd.t261 gnd 0.030974f
C3298 vdd.n271 gnd 0.212878f
C3299 vdd.n272 gnd 0.135088f
C3300 vdd.t250 gnd 0.030974f
C3301 vdd.t264 gnd 0.030974f
C3302 vdd.n273 gnd 0.212878f
C3303 vdd.n274 gnd 0.135088f
C3304 vdd.t149 gnd 0.030974f
C3305 vdd.t44 gnd 0.030974f
C3306 vdd.n275 gnd 0.212878f
C3307 vdd.n276 gnd 0.135088f
C3308 vdd.t30 gnd 0.030974f
C3309 vdd.t50 gnd 0.030974f
C3310 vdd.n277 gnd 0.212878f
C3311 vdd.n278 gnd 0.135088f
C3312 vdd.n279 gnd 0.00528f
C3313 vdd.n280 gnd 0.0049f
C3314 vdd.n281 gnd 0.00271f
C3315 vdd.n282 gnd 0.006223f
C3316 vdd.n283 gnd 0.002633f
C3317 vdd.n284 gnd 0.002788f
C3318 vdd.n285 gnd 0.0049f
C3319 vdd.n286 gnd 0.002633f
C3320 vdd.n287 gnd 0.006223f
C3321 vdd.n288 gnd 0.002788f
C3322 vdd.n289 gnd 0.0049f
C3323 vdd.n290 gnd 0.002633f
C3324 vdd.n291 gnd 0.004667f
C3325 vdd.n292 gnd 0.004681f
C3326 vdd.t57 gnd 0.01337f
C3327 vdd.n293 gnd 0.029747f
C3328 vdd.n294 gnd 0.154813f
C3329 vdd.n295 gnd 0.002633f
C3330 vdd.n296 gnd 0.002788f
C3331 vdd.n297 gnd 0.006223f
C3332 vdd.n298 gnd 0.006223f
C3333 vdd.n299 gnd 0.002788f
C3334 vdd.n300 gnd 0.002633f
C3335 vdd.n301 gnd 0.0049f
C3336 vdd.n302 gnd 0.0049f
C3337 vdd.n303 gnd 0.002633f
C3338 vdd.n304 gnd 0.002788f
C3339 vdd.n305 gnd 0.006223f
C3340 vdd.n306 gnd 0.006223f
C3341 vdd.n307 gnd 0.002788f
C3342 vdd.n308 gnd 0.002633f
C3343 vdd.n309 gnd 0.0049f
C3344 vdd.n310 gnd 0.0049f
C3345 vdd.n311 gnd 0.002633f
C3346 vdd.n312 gnd 0.002788f
C3347 vdd.n313 gnd 0.006223f
C3348 vdd.n314 gnd 0.006223f
C3349 vdd.n315 gnd 0.014713f
C3350 vdd.n316 gnd 0.00271f
C3351 vdd.n317 gnd 0.002633f
C3352 vdd.n318 gnd 0.012664f
C3353 vdd.n319 gnd 0.008564f
C3354 vdd.n320 gnd 0.059791f
C3355 vdd.n321 gnd 0.241267f
C3356 vdd.n322 gnd 0.007394f
C3357 vdd.n323 gnd 0.009621f
C3358 vdd.n324 gnd 0.007744f
C3359 vdd.n325 gnd 0.007744f
C3360 vdd.n326 gnd 0.009621f
C3361 vdd.n327 gnd 0.009621f
C3362 vdd.n328 gnd 0.702993f
C3363 vdd.n329 gnd 0.009621f
C3364 vdd.n330 gnd 0.009621f
C3365 vdd.n331 gnd 0.009621f
C3366 vdd.n332 gnd 0.761985f
C3367 vdd.n333 gnd 0.009621f
C3368 vdd.n334 gnd 0.009621f
C3369 vdd.n335 gnd 0.009621f
C3370 vdd.n336 gnd 0.009621f
C3371 vdd.n337 gnd 0.007744f
C3372 vdd.n338 gnd 0.009621f
C3373 vdd.t146 gnd 0.491603f
C3374 vdd.n339 gnd 0.009621f
C3375 vdd.n340 gnd 0.009621f
C3376 vdd.n341 gnd 0.009621f
C3377 vdd.t43 gnd 0.491603f
C3378 vdd.n342 gnd 0.009621f
C3379 vdd.n343 gnd 0.009621f
C3380 vdd.n344 gnd 0.009621f
C3381 vdd.n345 gnd 0.009621f
C3382 vdd.n346 gnd 0.009621f
C3383 vdd.n347 gnd 0.007744f
C3384 vdd.n348 gnd 0.009621f
C3385 vdd.n349 gnd 0.555512f
C3386 vdd.n350 gnd 0.009621f
C3387 vdd.n351 gnd 0.009621f
C3388 vdd.n352 gnd 0.009621f
C3389 vdd.t49 gnd 0.491603f
C3390 vdd.n353 gnd 0.009621f
C3391 vdd.n354 gnd 0.009621f
C3392 vdd.n355 gnd 0.009621f
C3393 vdd.n356 gnd 0.009621f
C3394 vdd.n357 gnd 0.009621f
C3395 vdd.n358 gnd 0.007744f
C3396 vdd.n359 gnd 0.009621f
C3397 vdd.t56 gnd 0.491603f
C3398 vdd.n360 gnd 0.009621f
C3399 vdd.n361 gnd 0.009621f
C3400 vdd.n362 gnd 0.009621f
C3401 vdd.n363 gnd 0.830809f
C3402 vdd.n364 gnd 0.009621f
C3403 vdd.n365 gnd 0.009621f
C3404 vdd.n366 gnd 0.009621f
C3405 vdd.n367 gnd 0.009621f
C3406 vdd.n368 gnd 0.009621f
C3407 vdd.n369 gnd 0.006427f
C3408 vdd.n370 gnd 0.021909f
C3409 vdd.t84 gnd 0.491603f
C3410 vdd.n371 gnd 0.009621f
C3411 vdd.n372 gnd 0.021909f
C3412 vdd.n404 gnd 0.009621f
C3413 vdd.t109 gnd 0.118362f
C3414 vdd.t108 gnd 0.126496f
C3415 vdd.t107 gnd 0.154579f
C3416 vdd.n405 gnd 0.198149f
C3417 vdd.n406 gnd 0.167255f
C3418 vdd.n407 gnd 0.0127f
C3419 vdd.n408 gnd 0.009621f
C3420 vdd.n409 gnd 0.007744f
C3421 vdd.n410 gnd 0.009621f
C3422 vdd.n411 gnd 0.007744f
C3423 vdd.n412 gnd 0.009621f
C3424 vdd.n413 gnd 0.007744f
C3425 vdd.n414 gnd 0.009621f
C3426 vdd.n415 gnd 0.007744f
C3427 vdd.n416 gnd 0.009621f
C3428 vdd.n417 gnd 0.007744f
C3429 vdd.n418 gnd 0.009621f
C3430 vdd.t86 gnd 0.118362f
C3431 vdd.t85 gnd 0.126496f
C3432 vdd.t83 gnd 0.154579f
C3433 vdd.n419 gnd 0.198149f
C3434 vdd.n420 gnd 0.167255f
C3435 vdd.n421 gnd 0.007744f
C3436 vdd.n422 gnd 0.009621f
C3437 vdd.n423 gnd 0.007744f
C3438 vdd.n424 gnd 0.009621f
C3439 vdd.n425 gnd 0.007744f
C3440 vdd.n426 gnd 0.009621f
C3441 vdd.n427 gnd 0.007744f
C3442 vdd.n428 gnd 0.009621f
C3443 vdd.n429 gnd 0.007744f
C3444 vdd.n430 gnd 0.009621f
C3445 vdd.t100 gnd 0.118362f
C3446 vdd.t99 gnd 0.126496f
C3447 vdd.t98 gnd 0.154579f
C3448 vdd.n431 gnd 0.198149f
C3449 vdd.n432 gnd 0.167255f
C3450 vdd.n433 gnd 0.016571f
C3451 vdd.n434 gnd 0.009621f
C3452 vdd.n435 gnd 0.007744f
C3453 vdd.n436 gnd 0.009621f
C3454 vdd.n437 gnd 0.007744f
C3455 vdd.n438 gnd 0.009621f
C3456 vdd.n439 gnd 0.007744f
C3457 vdd.n440 gnd 0.009621f
C3458 vdd.n441 gnd 0.007744f
C3459 vdd.n442 gnd 0.009621f
C3460 vdd.n443 gnd 0.021909f
C3461 vdd.n444 gnd 0.022059f
C3462 vdd.n445 gnd 0.022059f
C3463 vdd.n446 gnd 0.006427f
C3464 vdd.n447 gnd 0.007744f
C3465 vdd.n448 gnd 0.009621f
C3466 vdd.n449 gnd 0.009621f
C3467 vdd.n450 gnd 0.007744f
C3468 vdd.n451 gnd 0.009621f
C3469 vdd.n452 gnd 0.009621f
C3470 vdd.n453 gnd 0.009621f
C3471 vdd.n454 gnd 0.009621f
C3472 vdd.n455 gnd 0.009621f
C3473 vdd.n456 gnd 0.007744f
C3474 vdd.n457 gnd 0.007744f
C3475 vdd.n458 gnd 0.009621f
C3476 vdd.n459 gnd 0.009621f
C3477 vdd.n460 gnd 0.007744f
C3478 vdd.n461 gnd 0.009621f
C3479 vdd.n462 gnd 0.009621f
C3480 vdd.n463 gnd 0.009621f
C3481 vdd.n464 gnd 0.009621f
C3482 vdd.n465 gnd 0.009621f
C3483 vdd.n466 gnd 0.007744f
C3484 vdd.n467 gnd 0.007744f
C3485 vdd.n468 gnd 0.009621f
C3486 vdd.n469 gnd 0.009621f
C3487 vdd.n470 gnd 0.007744f
C3488 vdd.n471 gnd 0.009621f
C3489 vdd.n472 gnd 0.009621f
C3490 vdd.n473 gnd 0.009621f
C3491 vdd.n474 gnd 0.009621f
C3492 vdd.n475 gnd 0.009621f
C3493 vdd.n476 gnd 0.007744f
C3494 vdd.n477 gnd 0.007744f
C3495 vdd.n478 gnd 0.009621f
C3496 vdd.n479 gnd 0.009621f
C3497 vdd.n480 gnd 0.007744f
C3498 vdd.n481 gnd 0.009621f
C3499 vdd.n482 gnd 0.009621f
C3500 vdd.n483 gnd 0.009621f
C3501 vdd.n484 gnd 0.009621f
C3502 vdd.n485 gnd 0.009621f
C3503 vdd.n486 gnd 0.007744f
C3504 vdd.n487 gnd 0.007744f
C3505 vdd.n488 gnd 0.009621f
C3506 vdd.n489 gnd 0.009621f
C3507 vdd.n490 gnd 0.006466f
C3508 vdd.n491 gnd 0.009621f
C3509 vdd.n492 gnd 0.009621f
C3510 vdd.n493 gnd 0.009621f
C3511 vdd.n494 gnd 0.009621f
C3512 vdd.n495 gnd 0.009621f
C3513 vdd.n496 gnd 0.006466f
C3514 vdd.n497 gnd 0.007744f
C3515 vdd.n498 gnd 0.009621f
C3516 vdd.n499 gnd 0.009621f
C3517 vdd.n500 gnd 0.007744f
C3518 vdd.n501 gnd 0.009621f
C3519 vdd.n502 gnd 0.009621f
C3520 vdd.n503 gnd 0.009621f
C3521 vdd.n504 gnd 0.009621f
C3522 vdd.n505 gnd 0.009621f
C3523 vdd.n506 gnd 0.007744f
C3524 vdd.n507 gnd 0.007744f
C3525 vdd.n508 gnd 0.009621f
C3526 vdd.n509 gnd 0.009621f
C3527 vdd.n510 gnd 0.007744f
C3528 vdd.n511 gnd 0.009621f
C3529 vdd.n512 gnd 0.009621f
C3530 vdd.n513 gnd 0.009621f
C3531 vdd.n514 gnd 0.009621f
C3532 vdd.n515 gnd 0.009621f
C3533 vdd.n516 gnd 0.007744f
C3534 vdd.n517 gnd 0.007744f
C3535 vdd.n518 gnd 0.009621f
C3536 vdd.n519 gnd 0.009621f
C3537 vdd.n520 gnd 0.007744f
C3538 vdd.n521 gnd 0.009621f
C3539 vdd.n522 gnd 0.009621f
C3540 vdd.n523 gnd 0.009621f
C3541 vdd.n524 gnd 0.009621f
C3542 vdd.n525 gnd 0.009621f
C3543 vdd.n526 gnd 0.007744f
C3544 vdd.n527 gnd 0.007744f
C3545 vdd.n528 gnd 0.009621f
C3546 vdd.n529 gnd 0.009621f
C3547 vdd.n530 gnd 0.007744f
C3548 vdd.n531 gnd 0.009621f
C3549 vdd.n532 gnd 0.009621f
C3550 vdd.n533 gnd 0.009621f
C3551 vdd.n534 gnd 0.009621f
C3552 vdd.n535 gnd 0.009621f
C3553 vdd.n536 gnd 0.007744f
C3554 vdd.n537 gnd 0.007744f
C3555 vdd.n538 gnd 0.009621f
C3556 vdd.n539 gnd 0.009621f
C3557 vdd.n540 gnd 0.007744f
C3558 vdd.n541 gnd 0.009621f
C3559 vdd.n542 gnd 0.009621f
C3560 vdd.n543 gnd 0.009621f
C3561 vdd.n544 gnd 0.009621f
C3562 vdd.n545 gnd 0.009621f
C3563 vdd.n546 gnd 0.005266f
C3564 vdd.n547 gnd 0.016571f
C3565 vdd.n548 gnd 0.009621f
C3566 vdd.n549 gnd 0.009621f
C3567 vdd.n550 gnd 0.007666f
C3568 vdd.n551 gnd 0.009621f
C3569 vdd.n552 gnd 0.009621f
C3570 vdd.n553 gnd 0.009621f
C3571 vdd.n554 gnd 0.009621f
C3572 vdd.n555 gnd 0.009621f
C3573 vdd.n556 gnd 0.007744f
C3574 vdd.n557 gnd 0.007744f
C3575 vdd.n558 gnd 0.009621f
C3576 vdd.n559 gnd 0.009621f
C3577 vdd.n560 gnd 0.007744f
C3578 vdd.n561 gnd 0.009621f
C3579 vdd.n562 gnd 0.009621f
C3580 vdd.n563 gnd 0.009621f
C3581 vdd.n564 gnd 0.009621f
C3582 vdd.n565 gnd 0.009621f
C3583 vdd.n566 gnd 0.007744f
C3584 vdd.n567 gnd 0.007744f
C3585 vdd.n568 gnd 0.009621f
C3586 vdd.n569 gnd 0.009621f
C3587 vdd.n570 gnd 0.007744f
C3588 vdd.n571 gnd 0.009621f
C3589 vdd.n572 gnd 0.009621f
C3590 vdd.n573 gnd 0.009621f
C3591 vdd.n574 gnd 0.009621f
C3592 vdd.n575 gnd 0.009621f
C3593 vdd.n576 gnd 0.007744f
C3594 vdd.n577 gnd 0.007744f
C3595 vdd.n578 gnd 0.009621f
C3596 vdd.n579 gnd 0.009621f
C3597 vdd.n580 gnd 0.007744f
C3598 vdd.n581 gnd 0.009621f
C3599 vdd.n582 gnd 0.009621f
C3600 vdd.n583 gnd 0.009621f
C3601 vdd.n584 gnd 0.009621f
C3602 vdd.n585 gnd 0.009621f
C3603 vdd.n586 gnd 0.007744f
C3604 vdd.n587 gnd 0.007744f
C3605 vdd.n588 gnd 0.009621f
C3606 vdd.n589 gnd 0.009621f
C3607 vdd.n590 gnd 0.007744f
C3608 vdd.n591 gnd 0.009621f
C3609 vdd.n592 gnd 0.009621f
C3610 vdd.n593 gnd 0.009621f
C3611 vdd.n594 gnd 0.009621f
C3612 vdd.n595 gnd 0.009621f
C3613 vdd.n596 gnd 0.007744f
C3614 vdd.n597 gnd 0.009621f
C3615 vdd.n598 gnd 0.007744f
C3616 vdd.n599 gnd 0.004065f
C3617 vdd.n600 gnd 0.009621f
C3618 vdd.n601 gnd 0.009621f
C3619 vdd.n602 gnd 0.007744f
C3620 vdd.n603 gnd 0.009621f
C3621 vdd.n604 gnd 0.007744f
C3622 vdd.n605 gnd 0.009621f
C3623 vdd.n606 gnd 0.007744f
C3624 vdd.n607 gnd 0.009621f
C3625 vdd.n608 gnd 0.007744f
C3626 vdd.n609 gnd 0.009621f
C3627 vdd.n610 gnd 0.007744f
C3628 vdd.n611 gnd 0.009621f
C3629 vdd.n612 gnd 0.009621f
C3630 vdd.n613 gnd 0.535848f
C3631 vdd.t152 gnd 0.491603f
C3632 vdd.n614 gnd 0.009621f
C3633 vdd.n615 gnd 0.007744f
C3634 vdd.n616 gnd 0.009621f
C3635 vdd.n617 gnd 0.007744f
C3636 vdd.n618 gnd 0.009621f
C3637 vdd.t53 gnd 0.491603f
C3638 vdd.n619 gnd 0.009621f
C3639 vdd.n620 gnd 0.007744f
C3640 vdd.n621 gnd 0.009621f
C3641 vdd.n622 gnd 0.007744f
C3642 vdd.n623 gnd 0.009621f
C3643 vdd.t171 gnd 0.491603f
C3644 vdd.n624 gnd 0.614504f
C3645 vdd.n625 gnd 0.009621f
C3646 vdd.n626 gnd 0.007744f
C3647 vdd.n627 gnd 0.009621f
C3648 vdd.n628 gnd 0.007744f
C3649 vdd.n629 gnd 0.009621f
C3650 vdd.t21 gnd 0.491603f
C3651 vdd.n630 gnd 0.009621f
C3652 vdd.n631 gnd 0.007744f
C3653 vdd.n632 gnd 0.009621f
C3654 vdd.n633 gnd 0.007744f
C3655 vdd.n634 gnd 0.009621f
C3656 vdd.n635 gnd 0.683328f
C3657 vdd.n636 gnd 0.816061f
C3658 vdd.t33 gnd 0.491603f
C3659 vdd.n637 gnd 0.009621f
C3660 vdd.n638 gnd 0.007744f
C3661 vdd.n639 gnd 0.009621f
C3662 vdd.n640 gnd 0.007744f
C3663 vdd.n641 gnd 0.009621f
C3664 vdd.n642 gnd 0.516183f
C3665 vdd.n643 gnd 0.009621f
C3666 vdd.n644 gnd 0.007744f
C3667 vdd.n645 gnd 0.009621f
C3668 vdd.n646 gnd 0.007744f
C3669 vdd.n647 gnd 0.009621f
C3670 vdd.n648 gnd 0.983206f
C3671 vdd.t51 gnd 0.491603f
C3672 vdd.n649 gnd 0.009621f
C3673 vdd.n650 gnd 0.007744f
C3674 vdd.n651 gnd 0.009621f
C3675 vdd.n652 gnd 0.007744f
C3676 vdd.n653 gnd 0.009621f
C3677 vdd.t88 gnd 0.491603f
C3678 vdd.n654 gnd 0.009621f
C3679 vdd.n655 gnd 0.007744f
C3680 vdd.n656 gnd 0.022059f
C3681 vdd.n657 gnd 0.022059f
C3682 vdd.n658 gnd 11.8476f
C3683 vdd.n659 gnd 0.54568f
C3684 vdd.n660 gnd 0.022059f
C3685 vdd.n661 gnd 0.008274f
C3686 vdd.n662 gnd 0.007744f
C3687 vdd.n667 gnd 0.006157f
C3688 vdd.n668 gnd 0.007744f
C3689 vdd.n669 gnd 0.009621f
C3690 vdd.n670 gnd 0.009621f
C3691 vdd.n671 gnd 0.009621f
C3692 vdd.n672 gnd 0.009621f
C3693 vdd.n673 gnd 0.009621f
C3694 vdd.n674 gnd 0.007744f
C3695 vdd.n675 gnd 0.009621f
C3696 vdd.n676 gnd 0.009621f
C3697 vdd.n677 gnd 0.009621f
C3698 vdd.n678 gnd 0.009621f
C3699 vdd.n679 gnd 0.009621f
C3700 vdd.n680 gnd 0.007744f
C3701 vdd.n681 gnd 0.009621f
C3702 vdd.n682 gnd 0.009621f
C3703 vdd.n683 gnd 0.009621f
C3704 vdd.n684 gnd 0.009621f
C3705 vdd.n685 gnd 0.009621f
C3706 vdd.t119 gnd 0.118362f
C3707 vdd.t120 gnd 0.126496f
C3708 vdd.t118 gnd 0.154579f
C3709 vdd.n686 gnd 0.198149f
C3710 vdd.n687 gnd 0.166481f
C3711 vdd.n688 gnd 0.015797f
C3712 vdd.n689 gnd 0.009621f
C3713 vdd.n690 gnd 0.009621f
C3714 vdd.n691 gnd 0.009621f
C3715 vdd.n692 gnd 0.009621f
C3716 vdd.n693 gnd 0.009621f
C3717 vdd.n694 gnd 0.007744f
C3718 vdd.n695 gnd 0.009621f
C3719 vdd.n696 gnd 0.009621f
C3720 vdd.n697 gnd 0.009621f
C3721 vdd.n698 gnd 0.009621f
C3722 vdd.n699 gnd 0.009621f
C3723 vdd.n700 gnd 0.007744f
C3724 vdd.n701 gnd 0.009621f
C3725 vdd.n702 gnd 0.009621f
C3726 vdd.n703 gnd 0.009621f
C3727 vdd.n704 gnd 0.009621f
C3728 vdd.n705 gnd 0.009621f
C3729 vdd.n706 gnd 0.007744f
C3730 vdd.n707 gnd 0.009621f
C3731 vdd.n708 gnd 0.009621f
C3732 vdd.n709 gnd 0.009621f
C3733 vdd.n710 gnd 0.009621f
C3734 vdd.n711 gnd 0.009621f
C3735 vdd.n712 gnd 0.007744f
C3736 vdd.n713 gnd 0.009621f
C3737 vdd.n714 gnd 0.009621f
C3738 vdd.n715 gnd 0.009621f
C3739 vdd.n716 gnd 0.009621f
C3740 vdd.n717 gnd 0.009621f
C3741 vdd.n718 gnd 0.007744f
C3742 vdd.n719 gnd 0.009621f
C3743 vdd.n720 gnd 0.009621f
C3744 vdd.n721 gnd 0.009621f
C3745 vdd.n722 gnd 0.007666f
C3746 vdd.t102 gnd 0.118362f
C3747 vdd.t103 gnd 0.126496f
C3748 vdd.t101 gnd 0.154579f
C3749 vdd.n723 gnd 0.198149f
C3750 vdd.n724 gnd 0.166481f
C3751 vdd.n725 gnd 0.009621f
C3752 vdd.n726 gnd 0.007744f
C3753 vdd.n728 gnd 0.009621f
C3754 vdd.n730 gnd 0.009621f
C3755 vdd.n731 gnd 0.009621f
C3756 vdd.n732 gnd 0.007744f
C3757 vdd.n733 gnd 0.009621f
C3758 vdd.n734 gnd 0.009621f
C3759 vdd.n735 gnd 0.009621f
C3760 vdd.n736 gnd 0.009621f
C3761 vdd.n737 gnd 0.009621f
C3762 vdd.n738 gnd 0.007744f
C3763 vdd.n739 gnd 0.009621f
C3764 vdd.n740 gnd 0.009621f
C3765 vdd.n741 gnd 0.009621f
C3766 vdd.n742 gnd 0.009621f
C3767 vdd.n743 gnd 0.009621f
C3768 vdd.n744 gnd 0.007744f
C3769 vdd.n745 gnd 0.009621f
C3770 vdd.n746 gnd 0.009621f
C3771 vdd.n747 gnd 0.009621f
C3772 vdd.n748 gnd 0.006157f
C3773 vdd.n753 gnd 0.006542f
C3774 vdd.n754 gnd 0.006542f
C3775 vdd.n755 gnd 0.006542f
C3776 vdd.n756 gnd 11.6117f
C3777 vdd.n757 gnd 0.006542f
C3778 vdd.n758 gnd 0.006542f
C3779 vdd.n759 gnd 0.006542f
C3780 vdd.n761 gnd 0.006542f
C3781 vdd.n762 gnd 0.006542f
C3782 vdd.n764 gnd 0.006542f
C3783 vdd.n765 gnd 0.004762f
C3784 vdd.n767 gnd 0.006542f
C3785 vdd.t68 gnd 0.264369f
C3786 vdd.t67 gnd 0.270614f
C3787 vdd.t65 gnd 0.17259f
C3788 vdd.n768 gnd 0.093276f
C3789 vdd.n769 gnd 0.052909f
C3790 vdd.n770 gnd 0.00935f
C3791 vdd.n771 gnd 0.014855f
C3792 vdd.n773 gnd 0.006542f
C3793 vdd.n774 gnd 0.66858f
C3794 vdd.n775 gnd 0.014008f
C3795 vdd.n776 gnd 0.014008f
C3796 vdd.n777 gnd 0.006542f
C3797 vdd.n778 gnd 0.014855f
C3798 vdd.n779 gnd 0.006542f
C3799 vdd.n780 gnd 0.006542f
C3800 vdd.n781 gnd 0.006542f
C3801 vdd.n782 gnd 0.006542f
C3802 vdd.n783 gnd 0.006542f
C3803 vdd.n785 gnd 0.006542f
C3804 vdd.n786 gnd 0.006542f
C3805 vdd.n788 gnd 0.006542f
C3806 vdd.n789 gnd 0.006542f
C3807 vdd.n791 gnd 0.006542f
C3808 vdd.n792 gnd 0.006542f
C3809 vdd.n794 gnd 0.006542f
C3810 vdd.n795 gnd 0.006542f
C3811 vdd.n797 gnd 0.006542f
C3812 vdd.n798 gnd 0.006542f
C3813 vdd.n800 gnd 0.006542f
C3814 vdd.n801 gnd 0.004762f
C3815 vdd.n803 gnd 0.006542f
C3816 vdd.t82 gnd 0.264369f
C3817 vdd.t81 gnd 0.270614f
C3818 vdd.t80 gnd 0.17259f
C3819 vdd.n804 gnd 0.093276f
C3820 vdd.n805 gnd 0.052909f
C3821 vdd.n806 gnd 0.00935f
C3822 vdd.n807 gnd 0.006542f
C3823 vdd.n808 gnd 0.006542f
C3824 vdd.t66 gnd 0.33429f
C3825 vdd.n809 gnd 0.006542f
C3826 vdd.n810 gnd 0.006542f
C3827 vdd.n811 gnd 0.006542f
C3828 vdd.n812 gnd 0.006542f
C3829 vdd.n813 gnd 0.006542f
C3830 vdd.n814 gnd 0.66858f
C3831 vdd.n815 gnd 0.006542f
C3832 vdd.n816 gnd 0.006542f
C3833 vdd.n817 gnd 0.526015f
C3834 vdd.n818 gnd 0.006542f
C3835 vdd.n819 gnd 0.006542f
C3836 vdd.n820 gnd 0.006542f
C3837 vdd.n821 gnd 0.006542f
C3838 vdd.n822 gnd 0.66858f
C3839 vdd.n823 gnd 0.006542f
C3840 vdd.n824 gnd 0.006542f
C3841 vdd.n825 gnd 0.006542f
C3842 vdd.n826 gnd 0.006542f
C3843 vdd.n827 gnd 0.006542f
C3844 vdd.t208 gnd 0.33429f
C3845 vdd.n828 gnd 0.006542f
C3846 vdd.n829 gnd 0.006542f
C3847 vdd.n830 gnd 0.006542f
C3848 vdd.n831 gnd 0.006542f
C3849 vdd.n832 gnd 0.006542f
C3850 vdd.t225 gnd 0.33429f
C3851 vdd.n833 gnd 0.006542f
C3852 vdd.n834 gnd 0.006542f
C3853 vdd.n835 gnd 0.644f
C3854 vdd.n836 gnd 0.006542f
C3855 vdd.n837 gnd 0.006542f
C3856 vdd.n838 gnd 0.006542f
C3857 vdd.t224 gnd 0.33429f
C3858 vdd.n839 gnd 0.006542f
C3859 vdd.n840 gnd 0.006542f
C3860 vdd.n841 gnd 0.496519f
C3861 vdd.n842 gnd 0.006542f
C3862 vdd.n843 gnd 0.006542f
C3863 vdd.n844 gnd 0.006542f
C3864 vdd.n845 gnd 0.467023f
C3865 vdd.n846 gnd 0.006542f
C3866 vdd.n847 gnd 0.006542f
C3867 vdd.n848 gnd 0.349038f
C3868 vdd.n849 gnd 0.006542f
C3869 vdd.n850 gnd 0.006542f
C3870 vdd.n851 gnd 0.006542f
C3871 vdd.n852 gnd 0.614504f
C3872 vdd.n853 gnd 0.006542f
C3873 vdd.n854 gnd 0.006542f
C3874 vdd.t231 gnd 0.33429f
C3875 vdd.n855 gnd 0.006542f
C3876 vdd.n856 gnd 0.006542f
C3877 vdd.n857 gnd 0.006542f
C3878 vdd.n858 gnd 0.66858f
C3879 vdd.n859 gnd 0.006542f
C3880 vdd.n860 gnd 0.006542f
C3881 vdd.t232 gnd 0.33429f
C3882 vdd.n861 gnd 0.006542f
C3883 vdd.n862 gnd 0.006542f
C3884 vdd.n863 gnd 0.006542f
C3885 vdd.t202 gnd 0.33429f
C3886 vdd.n864 gnd 0.006542f
C3887 vdd.n865 gnd 0.006542f
C3888 vdd.n866 gnd 0.006542f
C3889 vdd.t93 gnd 0.270614f
C3890 vdd.t91 gnd 0.17259f
C3891 vdd.t94 gnd 0.270614f
C3892 vdd.n867 gnd 0.152096f
C3893 vdd.n868 gnd 0.018952f
C3894 vdd.n869 gnd 0.006542f
C3895 vdd.t92 gnd 0.240886f
C3896 vdd.n870 gnd 0.006542f
C3897 vdd.n871 gnd 0.006542f
C3898 vdd.n872 gnd 0.575176f
C3899 vdd.n873 gnd 0.006542f
C3900 vdd.n874 gnd 0.006542f
C3901 vdd.n875 gnd 0.006542f
C3902 vdd.n876 gnd 0.388367f
C3903 vdd.n877 gnd 0.006542f
C3904 vdd.n878 gnd 0.006542f
C3905 vdd.t203 gnd 0.137649f
C3906 vdd.n879 gnd 0.427695f
C3907 vdd.n880 gnd 0.006542f
C3908 vdd.n881 gnd 0.006542f
C3909 vdd.n882 gnd 0.006542f
C3910 vdd.n883 gnd 0.535848f
C3911 vdd.n884 gnd 0.006542f
C3912 vdd.n885 gnd 0.006542f
C3913 vdd.t216 gnd 0.33429f
C3914 vdd.n886 gnd 0.006542f
C3915 vdd.n887 gnd 0.006542f
C3916 vdd.n888 gnd 0.006542f
C3917 vdd.t212 gnd 0.33429f
C3918 vdd.n889 gnd 0.006542f
C3919 vdd.n890 gnd 0.006542f
C3920 vdd.t235 gnd 0.33429f
C3921 vdd.n891 gnd 0.006542f
C3922 vdd.n892 gnd 0.006542f
C3923 vdd.n893 gnd 0.006542f
C3924 vdd.t194 gnd 0.226137f
C3925 vdd.n894 gnd 0.006542f
C3926 vdd.n895 gnd 0.006542f
C3927 vdd.n896 gnd 0.589924f
C3928 vdd.n897 gnd 0.006542f
C3929 vdd.n898 gnd 0.006542f
C3930 vdd.n899 gnd 0.006542f
C3931 vdd.t236 gnd 0.33429f
C3932 vdd.n900 gnd 0.006542f
C3933 vdd.n901 gnd 0.006542f
C3934 vdd.t248 gnd 0.319542f
C3935 vdd.n902 gnd 0.442443f
C3936 vdd.n903 gnd 0.006542f
C3937 vdd.n904 gnd 0.006542f
C3938 vdd.n905 gnd 0.006542f
C3939 vdd.t198 gnd 0.33429f
C3940 vdd.n906 gnd 0.006542f
C3941 vdd.n907 gnd 0.006542f
C3942 vdd.t240 gnd 0.33429f
C3943 vdd.n908 gnd 0.006542f
C3944 vdd.n909 gnd 0.006542f
C3945 vdd.n910 gnd 0.006542f
C3946 vdd.n911 gnd 0.66858f
C3947 vdd.n912 gnd 0.006542f
C3948 vdd.n913 gnd 0.006542f
C3949 vdd.t220 gnd 0.33429f
C3950 vdd.n914 gnd 0.006542f
C3951 vdd.n915 gnd 0.006542f
C3952 vdd.n916 gnd 0.006542f
C3953 vdd.n917 gnd 0.462107f
C3954 vdd.n918 gnd 0.006542f
C3955 vdd.n919 gnd 0.006542f
C3956 vdd.n920 gnd 0.006542f
C3957 vdd.n921 gnd 0.006542f
C3958 vdd.n922 gnd 0.006542f
C3959 vdd.t122 gnd 0.33429f
C3960 vdd.n923 gnd 0.006542f
C3961 vdd.n924 gnd 0.006542f
C3962 vdd.t200 gnd 0.33429f
C3963 vdd.n925 gnd 0.006542f
C3964 vdd.n926 gnd 0.014008f
C3965 vdd.n927 gnd 0.014008f
C3966 vdd.n928 gnd 0.757069f
C3967 vdd.n929 gnd 0.006542f
C3968 vdd.n930 gnd 0.006542f
C3969 vdd.t229 gnd 0.33429f
C3970 vdd.n931 gnd 0.014008f
C3971 vdd.n932 gnd 0.006542f
C3972 vdd.n933 gnd 0.006542f
C3973 vdd.t242 gnd 0.57026f
C3974 vdd.n951 gnd 0.014855f
C3975 vdd.n969 gnd 0.014008f
C3976 vdd.n970 gnd 0.006542f
C3977 vdd.n971 gnd 0.014008f
C3978 vdd.t140 gnd 0.264369f
C3979 vdd.t139 gnd 0.270614f
C3980 vdd.t138 gnd 0.17259f
C3981 vdd.n972 gnd 0.093276f
C3982 vdd.n973 gnd 0.052909f
C3983 vdd.n974 gnd 0.014855f
C3984 vdd.n975 gnd 0.006542f
C3985 vdd.n976 gnd 0.393283f
C3986 vdd.n977 gnd 0.014008f
C3987 vdd.n978 gnd 0.006542f
C3988 vdd.n979 gnd 0.014855f
C3989 vdd.n980 gnd 0.006542f
C3990 vdd.t117 gnd 0.264369f
C3991 vdd.t116 gnd 0.270614f
C3992 vdd.t114 gnd 0.17259f
C3993 vdd.n981 gnd 0.093276f
C3994 vdd.n982 gnd 0.052909f
C3995 vdd.n983 gnd 0.00935f
C3996 vdd.n984 gnd 0.006542f
C3997 vdd.n985 gnd 0.006542f
C3998 vdd.t115 gnd 0.33429f
C3999 vdd.n986 gnd 0.006542f
C4000 vdd.t244 gnd 0.33429f
C4001 vdd.n987 gnd 0.006542f
C4002 vdd.n988 gnd 0.006542f
C4003 vdd.n989 gnd 0.006542f
C4004 vdd.n990 gnd 0.006542f
C4005 vdd.n991 gnd 0.006542f
C4006 vdd.n992 gnd 0.66858f
C4007 vdd.n993 gnd 0.006542f
C4008 vdd.n994 gnd 0.006542f
C4009 vdd.t214 gnd 0.33429f
C4010 vdd.n995 gnd 0.006542f
C4011 vdd.n996 gnd 0.006542f
C4012 vdd.n997 gnd 0.006542f
C4013 vdd.n998 gnd 0.006542f
C4014 vdd.n999 gnd 0.481771f
C4015 vdd.n1000 gnd 0.006542f
C4016 vdd.n1001 gnd 0.006542f
C4017 vdd.n1002 gnd 0.006542f
C4018 vdd.n1003 gnd 0.006542f
C4019 vdd.n1004 gnd 0.006542f
C4020 vdd.t195 gnd 0.33429f
C4021 vdd.n1005 gnd 0.006542f
C4022 vdd.n1006 gnd 0.006542f
C4023 vdd.t233 gnd 0.33429f
C4024 vdd.n1007 gnd 0.006542f
C4025 vdd.n1008 gnd 0.006542f
C4026 vdd.n1009 gnd 0.006542f
C4027 vdd.t219 gnd 0.33429f
C4028 vdd.n1010 gnd 0.006542f
C4029 vdd.n1011 gnd 0.006542f
C4030 vdd.t196 gnd 0.33429f
C4031 vdd.n1012 gnd 0.006542f
C4032 vdd.n1013 gnd 0.006542f
C4033 vdd.n1014 gnd 0.006542f
C4034 vdd.t217 gnd 0.319542f
C4035 vdd.n1015 gnd 0.006542f
C4036 vdd.n1016 gnd 0.006542f
C4037 vdd.n1017 gnd 0.496519f
C4038 vdd.n1018 gnd 0.006542f
C4039 vdd.n1019 gnd 0.006542f
C4040 vdd.n1020 gnd 0.006542f
C4041 vdd.t237 gnd 0.33429f
C4042 vdd.n1021 gnd 0.006542f
C4043 vdd.n1022 gnd 0.006542f
C4044 vdd.t205 gnd 0.226137f
C4045 vdd.n1023 gnd 0.349038f
C4046 vdd.n1024 gnd 0.006542f
C4047 vdd.n1025 gnd 0.006542f
C4048 vdd.n1026 gnd 0.006542f
C4049 vdd.n1027 gnd 0.614504f
C4050 vdd.n1028 gnd 0.006542f
C4051 vdd.n1029 gnd 0.006542f
C4052 vdd.t246 gnd 0.33429f
C4053 vdd.n1030 gnd 0.006542f
C4054 vdd.n1031 gnd 0.006542f
C4055 vdd.n1032 gnd 0.006542f
C4056 vdd.n1033 gnd 0.66858f
C4057 vdd.n1034 gnd 0.006542f
C4058 vdd.n1035 gnd 0.006542f
C4059 vdd.t211 gnd 0.33429f
C4060 vdd.n1036 gnd 0.006542f
C4061 vdd.n1037 gnd 0.006542f
C4062 vdd.n1038 gnd 0.006542f
C4063 vdd.t204 gnd 0.137649f
C4064 vdd.n1039 gnd 0.006542f
C4065 vdd.n1040 gnd 0.006542f
C4066 vdd.n1041 gnd 0.006542f
C4067 vdd.t130 gnd 0.270614f
C4068 vdd.t128 gnd 0.17259f
C4069 vdd.t131 gnd 0.270614f
C4070 vdd.n1042 gnd 0.152096f
C4071 vdd.n1043 gnd 0.006542f
C4072 vdd.n1044 gnd 0.006542f
C4073 vdd.t226 gnd 0.33429f
C4074 vdd.n1045 gnd 0.006542f
C4075 vdd.n1046 gnd 0.006542f
C4076 vdd.t129 gnd 0.240886f
C4077 vdd.n1047 gnd 0.530931f
C4078 vdd.n1048 gnd 0.006542f
C4079 vdd.n1049 gnd 0.006542f
C4080 vdd.n1050 gnd 0.006542f
C4081 vdd.n1051 gnd 0.388367f
C4082 vdd.n1052 gnd 0.006542f
C4083 vdd.n1053 gnd 0.006542f
C4084 vdd.n1054 gnd 0.427695f
C4085 vdd.n1055 gnd 0.006542f
C4086 vdd.n1056 gnd 0.006542f
C4087 vdd.n1057 gnd 0.006542f
C4088 vdd.n1058 gnd 0.535848f
C4089 vdd.n1059 gnd 0.006542f
C4090 vdd.n1060 gnd 0.006542f
C4091 vdd.t206 gnd 0.33429f
C4092 vdd.n1061 gnd 0.006542f
C4093 vdd.n1062 gnd 0.006542f
C4094 vdd.n1063 gnd 0.006542f
C4095 vdd.n1064 gnd 0.66858f
C4096 vdd.n1065 gnd 0.006542f
C4097 vdd.n1066 gnd 0.006542f
C4098 vdd.t207 gnd 0.33429f
C4099 vdd.n1067 gnd 0.006542f
C4100 vdd.n1068 gnd 0.006542f
C4101 vdd.n1069 gnd 0.006542f
C4102 vdd.t247 gnd 0.33429f
C4103 vdd.n1070 gnd 0.006542f
C4104 vdd.n1071 gnd 0.006542f
C4105 vdd.n1072 gnd 0.006542f
C4106 vdd.n1073 gnd 0.006542f
C4107 vdd.n1074 gnd 0.006542f
C4108 vdd.t239 gnd 0.33429f
C4109 vdd.n1075 gnd 0.006542f
C4110 vdd.n1076 gnd 0.006542f
C4111 vdd.n1077 gnd 0.653832f
C4112 vdd.n1078 gnd 0.006542f
C4113 vdd.n1079 gnd 0.006542f
C4114 vdd.n1080 gnd 0.006542f
C4115 vdd.t199 gnd 0.33429f
C4116 vdd.n1081 gnd 0.006542f
C4117 vdd.n1082 gnd 0.006542f
C4118 vdd.n1083 gnd 0.506351f
C4119 vdd.n1084 gnd 0.006542f
C4120 vdd.n1085 gnd 0.006542f
C4121 vdd.n1086 gnd 0.006542f
C4122 vdd.n1087 gnd 0.66858f
C4123 vdd.n1088 gnd 0.006542f
C4124 vdd.n1089 gnd 0.006542f
C4125 vdd.n1090 gnd 0.35887f
C4126 vdd.n1091 gnd 0.006542f
C4127 vdd.n1092 gnd 0.006542f
C4128 vdd.n1093 gnd 0.006542f
C4129 vdd.n1094 gnd 0.66858f
C4130 vdd.n1095 gnd 0.006542f
C4131 vdd.n1096 gnd 0.006542f
C4132 vdd.n1097 gnd 0.006542f
C4133 vdd.n1098 gnd 0.006542f
C4134 vdd.n1099 gnd 0.006542f
C4135 vdd.t70 gnd 0.33429f
C4136 vdd.n1100 gnd 0.006542f
C4137 vdd.n1101 gnd 0.006542f
C4138 vdd.n1102 gnd 0.006542f
C4139 vdd.n1103 gnd 0.014008f
C4140 vdd.n1104 gnd 0.014008f
C4141 vdd.n1105 gnd 0.90455f
C4142 vdd.n1106 gnd 0.006542f
C4143 vdd.n1107 gnd 0.006542f
C4144 vdd.n1108 gnd 0.476855f
C4145 vdd.n1109 gnd 0.014008f
C4146 vdd.n1110 gnd 0.006542f
C4147 vdd.n1111 gnd 0.006542f
C4148 vdd.n1112 gnd 11.8476f
C4149 vdd.n1146 gnd 0.014855f
C4150 vdd.n1147 gnd 0.006542f
C4151 vdd.n1148 gnd 0.006542f
C4152 vdd.n1149 gnd 0.006157f
C4153 vdd.n1152 gnd 0.022059f
C4154 vdd.n1153 gnd 0.006427f
C4155 vdd.n1154 gnd 0.007744f
C4156 vdd.n1156 gnd 0.009621f
C4157 vdd.n1157 gnd 0.009621f
C4158 vdd.n1158 gnd 0.007744f
C4159 vdd.n1160 gnd 0.009621f
C4160 vdd.n1161 gnd 0.009621f
C4161 vdd.n1162 gnd 0.009621f
C4162 vdd.n1163 gnd 0.009621f
C4163 vdd.n1164 gnd 0.009621f
C4164 vdd.n1165 gnd 0.007744f
C4165 vdd.n1167 gnd 0.009621f
C4166 vdd.n1168 gnd 0.009621f
C4167 vdd.n1169 gnd 0.009621f
C4168 vdd.n1170 gnd 0.009621f
C4169 vdd.n1171 gnd 0.009621f
C4170 vdd.n1172 gnd 0.007744f
C4171 vdd.n1174 gnd 0.009621f
C4172 vdd.n1175 gnd 0.009621f
C4173 vdd.n1176 gnd 0.009621f
C4174 vdd.n1177 gnd 0.009621f
C4175 vdd.n1178 gnd 0.006466f
C4176 vdd.t79 gnd 0.118362f
C4177 vdd.t78 gnd 0.126496f
C4178 vdd.t77 gnd 0.154579f
C4179 vdd.n1179 gnd 0.198149f
C4180 vdd.n1180 gnd 0.166481f
C4181 vdd.n1182 gnd 0.009621f
C4182 vdd.n1183 gnd 0.009621f
C4183 vdd.n1184 gnd 0.007744f
C4184 vdd.n1185 gnd 0.009621f
C4185 vdd.n1187 gnd 0.009621f
C4186 vdd.n1188 gnd 0.009621f
C4187 vdd.n1189 gnd 0.009621f
C4188 vdd.n1190 gnd 0.009621f
C4189 vdd.n1191 gnd 0.007744f
C4190 vdd.n1193 gnd 0.009621f
C4191 vdd.n1194 gnd 0.009621f
C4192 vdd.n1195 gnd 0.009621f
C4193 vdd.n1196 gnd 0.009621f
C4194 vdd.n1197 gnd 0.009621f
C4195 vdd.n1198 gnd 0.007744f
C4196 vdd.n1200 gnd 0.009621f
C4197 vdd.n1201 gnd 0.009621f
C4198 vdd.n1202 gnd 0.009621f
C4199 vdd.n1203 gnd 0.009621f
C4200 vdd.n1204 gnd 0.009621f
C4201 vdd.n1205 gnd 0.007744f
C4202 vdd.n1207 gnd 0.009621f
C4203 vdd.n1208 gnd 0.009621f
C4204 vdd.n1209 gnd 0.009621f
C4205 vdd.n1210 gnd 0.009621f
C4206 vdd.n1211 gnd 0.009621f
C4207 vdd.n1212 gnd 0.007744f
C4208 vdd.n1214 gnd 0.009621f
C4209 vdd.n1215 gnd 0.009621f
C4210 vdd.n1216 gnd 0.009621f
C4211 vdd.n1217 gnd 0.009621f
C4212 vdd.n1218 gnd 0.007666f
C4213 vdd.t76 gnd 0.118362f
C4214 vdd.t75 gnd 0.126496f
C4215 vdd.t73 gnd 0.154579f
C4216 vdd.n1219 gnd 0.198149f
C4217 vdd.n1220 gnd 0.166481f
C4218 vdd.n1222 gnd 0.009621f
C4219 vdd.n1223 gnd 0.009621f
C4220 vdd.n1224 gnd 0.007744f
C4221 vdd.n1225 gnd 0.009621f
C4222 vdd.n1227 gnd 0.009621f
C4223 vdd.n1228 gnd 0.009621f
C4224 vdd.n1229 gnd 0.009621f
C4225 vdd.n1230 gnd 0.009621f
C4226 vdd.n1231 gnd 0.007744f
C4227 vdd.n1233 gnd 0.009621f
C4228 vdd.n1234 gnd 0.009621f
C4229 vdd.n1235 gnd 0.009621f
C4230 vdd.n1236 gnd 0.009621f
C4231 vdd.n1237 gnd 0.009621f
C4232 vdd.n1238 gnd 0.007744f
C4233 vdd.n1240 gnd 0.009621f
C4234 vdd.n1241 gnd 0.009621f
C4235 vdd.n1242 gnd 0.009621f
C4236 vdd.n1243 gnd 0.009621f
C4237 vdd.n1244 gnd 0.009621f
C4238 vdd.n1245 gnd 0.007744f
C4239 vdd.n1247 gnd 0.009621f
C4240 vdd.n1248 gnd 0.009621f
C4241 vdd.n1249 gnd 0.006157f
C4242 vdd.n1250 gnd 0.007744f
C4243 vdd.n1251 gnd 0.014855f
C4244 vdd.n1252 gnd 0.014855f
C4245 vdd.n1253 gnd 0.006542f
C4246 vdd.n1254 gnd 0.006542f
C4247 vdd.n1255 gnd 0.006542f
C4248 vdd.n1256 gnd 0.006542f
C4249 vdd.n1257 gnd 0.006542f
C4250 vdd.n1258 gnd 0.006542f
C4251 vdd.n1259 gnd 0.006542f
C4252 vdd.n1260 gnd 0.006542f
C4253 vdd.n1261 gnd 0.006542f
C4254 vdd.n1262 gnd 0.006542f
C4255 vdd.n1263 gnd 0.006542f
C4256 vdd.n1264 gnd 0.006542f
C4257 vdd.n1265 gnd 0.006542f
C4258 vdd.n1266 gnd 0.006542f
C4259 vdd.n1267 gnd 0.006542f
C4260 vdd.n1268 gnd 0.006542f
C4261 vdd.n1269 gnd 0.006542f
C4262 vdd.n1270 gnd 0.006542f
C4263 vdd.n1271 gnd 0.006542f
C4264 vdd.n1272 gnd 0.006542f
C4265 vdd.n1273 gnd 0.006542f
C4266 vdd.n1274 gnd 0.006542f
C4267 vdd.n1275 gnd 0.006542f
C4268 vdd.n1276 gnd 0.006542f
C4269 vdd.n1277 gnd 0.006542f
C4270 vdd.n1278 gnd 0.006542f
C4271 vdd.n1279 gnd 0.006542f
C4272 vdd.n1280 gnd 0.006542f
C4273 vdd.n1281 gnd 0.006542f
C4274 vdd.n1282 gnd 0.006542f
C4275 vdd.n1283 gnd 0.006542f
C4276 vdd.n1284 gnd 0.006542f
C4277 vdd.n1285 gnd 0.006542f
C4278 vdd.t71 gnd 0.264369f
C4279 vdd.t72 gnd 0.270614f
C4280 vdd.t69 gnd 0.17259f
C4281 vdd.n1286 gnd 0.093276f
C4282 vdd.n1287 gnd 0.052909f
C4283 vdd.n1288 gnd 0.00935f
C4284 vdd.n1289 gnd 0.006542f
C4285 vdd.t105 gnd 0.264369f
C4286 vdd.t106 gnd 0.270614f
C4287 vdd.t104 gnd 0.17259f
C4288 vdd.n1290 gnd 0.093276f
C4289 vdd.n1291 gnd 0.052909f
C4290 vdd.n1292 gnd 0.006542f
C4291 vdd.n1293 gnd 0.006542f
C4292 vdd.n1294 gnd 0.006542f
C4293 vdd.n1295 gnd 0.006542f
C4294 vdd.n1296 gnd 0.006542f
C4295 vdd.n1297 gnd 0.006542f
C4296 vdd.n1298 gnd 0.006542f
C4297 vdd.n1299 gnd 0.006542f
C4298 vdd.n1300 gnd 0.006542f
C4299 vdd.n1301 gnd 0.006542f
C4300 vdd.n1302 gnd 0.006542f
C4301 vdd.n1303 gnd 0.006542f
C4302 vdd.n1304 gnd 0.006542f
C4303 vdd.n1305 gnd 0.006542f
C4304 vdd.n1306 gnd 0.006542f
C4305 vdd.n1307 gnd 0.006542f
C4306 vdd.n1308 gnd 0.006542f
C4307 vdd.n1309 gnd 0.006542f
C4308 vdd.n1310 gnd 0.006542f
C4309 vdd.n1311 gnd 0.006542f
C4310 vdd.n1312 gnd 0.006542f
C4311 vdd.n1313 gnd 0.006542f
C4312 vdd.n1314 gnd 0.006542f
C4313 vdd.n1315 gnd 0.006542f
C4314 vdd.n1316 gnd 0.006542f
C4315 vdd.n1317 gnd 0.006542f
C4316 vdd.n1318 gnd 0.004762f
C4317 vdd.n1319 gnd 0.00935f
C4318 vdd.n1320 gnd 0.005051f
C4319 vdd.n1321 gnd 0.006542f
C4320 vdd.n1322 gnd 0.006542f
C4321 vdd.n1323 gnd 0.006542f
C4322 vdd.n1324 gnd 0.014855f
C4323 vdd.n1325 gnd 0.014855f
C4324 vdd.n1326 gnd 0.014008f
C4325 vdd.n1327 gnd 0.014008f
C4326 vdd.n1328 gnd 0.006542f
C4327 vdd.n1329 gnd 0.006542f
C4328 vdd.n1330 gnd 0.006542f
C4329 vdd.n1331 gnd 0.006542f
C4330 vdd.n1332 gnd 0.006542f
C4331 vdd.n1333 gnd 0.006542f
C4332 vdd.n1334 gnd 0.006542f
C4333 vdd.n1335 gnd 0.006542f
C4334 vdd.n1336 gnd 0.006542f
C4335 vdd.n1337 gnd 0.006542f
C4336 vdd.n1338 gnd 0.006542f
C4337 vdd.n1339 gnd 0.006542f
C4338 vdd.n1340 gnd 0.006542f
C4339 vdd.n1341 gnd 0.006542f
C4340 vdd.n1342 gnd 0.006542f
C4341 vdd.n1343 gnd 0.006542f
C4342 vdd.n1344 gnd 0.006542f
C4343 vdd.n1345 gnd 0.006542f
C4344 vdd.n1346 gnd 0.006542f
C4345 vdd.n1347 gnd 0.006542f
C4346 vdd.n1348 gnd 0.006542f
C4347 vdd.n1349 gnd 0.006542f
C4348 vdd.n1350 gnd 0.006542f
C4349 vdd.n1351 gnd 0.006542f
C4350 vdd.n1352 gnd 0.006542f
C4351 vdd.n1353 gnd 0.006542f
C4352 vdd.n1354 gnd 0.006542f
C4353 vdd.n1355 gnd 0.006542f
C4354 vdd.n1356 gnd 0.006542f
C4355 vdd.n1357 gnd 0.006542f
C4356 vdd.n1358 gnd 0.006542f
C4357 vdd.n1359 gnd 0.006542f
C4358 vdd.n1360 gnd 0.006542f
C4359 vdd.n1361 gnd 0.006542f
C4360 vdd.n1362 gnd 0.006542f
C4361 vdd.n1363 gnd 0.006542f
C4362 vdd.n1364 gnd 0.006542f
C4363 vdd.n1365 gnd 0.006542f
C4364 vdd.n1366 gnd 0.006542f
C4365 vdd.n1367 gnd 0.006542f
C4366 vdd.n1368 gnd 0.006542f
C4367 vdd.n1369 gnd 0.006542f
C4368 vdd.n1370 gnd 0.398199f
C4369 vdd.n1371 gnd 0.006542f
C4370 vdd.n1372 gnd 0.006542f
C4371 vdd.n1373 gnd 0.006542f
C4372 vdd.n1374 gnd 0.006542f
C4373 vdd.n1375 gnd 0.006542f
C4374 vdd.n1376 gnd 0.006542f
C4375 vdd.n1377 gnd 0.006542f
C4376 vdd.n1378 gnd 0.006542f
C4377 vdd.n1379 gnd 0.006542f
C4378 vdd.n1380 gnd 0.006542f
C4379 vdd.n1381 gnd 0.006542f
C4380 vdd.n1382 gnd 0.006542f
C4381 vdd.n1383 gnd 0.006542f
C4382 vdd.n1384 gnd 0.006542f
C4383 vdd.n1385 gnd 0.006542f
C4384 vdd.n1386 gnd 0.006542f
C4385 vdd.n1387 gnd 0.006542f
C4386 vdd.n1388 gnd 0.006542f
C4387 vdd.n1389 gnd 0.006542f
C4388 vdd.n1390 gnd 0.006542f
C4389 vdd.n1391 gnd 0.006542f
C4390 vdd.n1392 gnd 0.006542f
C4391 vdd.n1393 gnd 0.006542f
C4392 vdd.n1394 gnd 0.006542f
C4393 vdd.n1395 gnd 0.006542f
C4394 vdd.n1396 gnd 0.604672f
C4395 vdd.n1397 gnd 0.006542f
C4396 vdd.n1398 gnd 0.006542f
C4397 vdd.n1399 gnd 0.006542f
C4398 vdd.n1400 gnd 0.006542f
C4399 vdd.n1401 gnd 0.006542f
C4400 vdd.n1402 gnd 0.006542f
C4401 vdd.n1403 gnd 0.006542f
C4402 vdd.n1404 gnd 0.006542f
C4403 vdd.n1405 gnd 0.006542f
C4404 vdd.n1406 gnd 0.006542f
C4405 vdd.n1407 gnd 0.006542f
C4406 vdd.n1408 gnd 0.211389f
C4407 vdd.n1409 gnd 0.006542f
C4408 vdd.n1410 gnd 0.006542f
C4409 vdd.n1411 gnd 0.006542f
C4410 vdd.n1412 gnd 0.006542f
C4411 vdd.n1413 gnd 0.006542f
C4412 vdd.n1414 gnd 0.006542f
C4413 vdd.n1415 gnd 0.006542f
C4414 vdd.n1416 gnd 0.006542f
C4415 vdd.n1417 gnd 0.006542f
C4416 vdd.n1418 gnd 0.006542f
C4417 vdd.n1419 gnd 0.006542f
C4418 vdd.n1420 gnd 0.006542f
C4419 vdd.n1421 gnd 0.006542f
C4420 vdd.n1422 gnd 0.006542f
C4421 vdd.n1423 gnd 0.006542f
C4422 vdd.n1424 gnd 0.006542f
C4423 vdd.n1425 gnd 0.006542f
C4424 vdd.n1426 gnd 0.006542f
C4425 vdd.n1427 gnd 0.006542f
C4426 vdd.n1428 gnd 0.006542f
C4427 vdd.n1429 gnd 0.006542f
C4428 vdd.n1430 gnd 0.006542f
C4429 vdd.n1431 gnd 0.006542f
C4430 vdd.n1432 gnd 0.006542f
C4431 vdd.n1433 gnd 0.006542f
C4432 vdd.n1434 gnd 0.006542f
C4433 vdd.n1435 gnd 0.006542f
C4434 vdd.n1436 gnd 0.006542f
C4435 vdd.n1437 gnd 0.006542f
C4436 vdd.n1438 gnd 0.006542f
C4437 vdd.n1439 gnd 0.006542f
C4438 vdd.n1440 gnd 0.006542f
C4439 vdd.n1441 gnd 0.006542f
C4440 vdd.n1442 gnd 0.006542f
C4441 vdd.n1443 gnd 0.006542f
C4442 vdd.n1444 gnd 0.006542f
C4443 vdd.n1445 gnd 0.006542f
C4444 vdd.n1446 gnd 0.006542f
C4445 vdd.n1447 gnd 0.006542f
C4446 vdd.n1448 gnd 0.006542f
C4447 vdd.n1449 gnd 0.006542f
C4448 vdd.n1450 gnd 0.006542f
C4449 vdd.n1451 gnd 0.014008f
C4450 vdd.n1452 gnd 0.014008f
C4451 vdd.n1453 gnd 0.014855f
C4452 vdd.n1454 gnd 0.006542f
C4453 vdd.n1455 gnd 0.006542f
C4454 vdd.n1456 gnd 0.005051f
C4455 vdd.n1457 gnd 0.006542f
C4456 vdd.n1458 gnd 0.006542f
C4457 vdd.n1459 gnd 0.004762f
C4458 vdd.n1460 gnd 0.006542f
C4459 vdd.n1461 gnd 0.006542f
C4460 vdd.n1462 gnd 0.006542f
C4461 vdd.n1463 gnd 0.006542f
C4462 vdd.n1464 gnd 0.006542f
C4463 vdd.n1465 gnd 0.006542f
C4464 vdd.n1466 gnd 0.006542f
C4465 vdd.n1467 gnd 0.006542f
C4466 vdd.n1468 gnd 0.006542f
C4467 vdd.n1469 gnd 0.006542f
C4468 vdd.n1470 gnd 0.006542f
C4469 vdd.n1471 gnd 0.006542f
C4470 vdd.n1472 gnd 0.006542f
C4471 vdd.n1473 gnd 0.006542f
C4472 vdd.n1474 gnd 0.006542f
C4473 vdd.n1475 gnd 0.006542f
C4474 vdd.n1476 gnd 0.006542f
C4475 vdd.n1477 gnd 0.006542f
C4476 vdd.n1478 gnd 0.006542f
C4477 vdd.n1479 gnd 0.006542f
C4478 vdd.n1480 gnd 0.006542f
C4479 vdd.n1481 gnd 0.006542f
C4480 vdd.n1482 gnd 0.006542f
C4481 vdd.n1483 gnd 0.006542f
C4482 vdd.n1484 gnd 0.006542f
C4483 vdd.n1485 gnd 0.006542f
C4484 vdd.n1486 gnd 0.044072f
C4485 vdd.n1488 gnd 0.022059f
C4486 vdd.n1489 gnd 0.007744f
C4487 vdd.n1491 gnd 0.009621f
C4488 vdd.n1492 gnd 0.007744f
C4489 vdd.n1493 gnd 0.009621f
C4490 vdd.n1495 gnd 0.009621f
C4491 vdd.n1496 gnd 0.009621f
C4492 vdd.n1498 gnd 0.009621f
C4493 vdd.n1499 gnd 0.006427f
C4494 vdd.n1500 gnd 0.54568f
C4495 vdd.n1501 gnd 0.009621f
C4496 vdd.n1502 gnd 0.022059f
C4497 vdd.n1503 gnd 0.007744f
C4498 vdd.n1504 gnd 0.009621f
C4499 vdd.n1505 gnd 0.007744f
C4500 vdd.n1506 gnd 0.009621f
C4501 vdd.n1507 gnd 0.983206f
C4502 vdd.n1508 gnd 0.009621f
C4503 vdd.n1509 gnd 0.007744f
C4504 vdd.n1510 gnd 0.007744f
C4505 vdd.n1511 gnd 0.009621f
C4506 vdd.n1512 gnd 0.007744f
C4507 vdd.n1513 gnd 0.009621f
C4508 vdd.t165 gnd 0.491603f
C4509 vdd.n1514 gnd 0.009621f
C4510 vdd.n1515 gnd 0.007744f
C4511 vdd.n1516 gnd 0.009621f
C4512 vdd.n1517 gnd 0.007744f
C4513 vdd.n1518 gnd 0.009621f
C4514 vdd.t4 gnd 0.491603f
C4515 vdd.n1519 gnd 0.009621f
C4516 vdd.n1520 gnd 0.007744f
C4517 vdd.n1521 gnd 0.009621f
C4518 vdd.n1522 gnd 0.007744f
C4519 vdd.n1523 gnd 0.009621f
C4520 vdd.t31 gnd 0.491603f
C4521 vdd.n1524 gnd 0.683328f
C4522 vdd.n1525 gnd 0.009621f
C4523 vdd.n1526 gnd 0.007744f
C4524 vdd.n1527 gnd 0.009621f
C4525 vdd.n1528 gnd 0.007744f
C4526 vdd.n1529 gnd 0.009621f
C4527 vdd.n1530 gnd 0.781649f
C4528 vdd.n1531 gnd 0.009621f
C4529 vdd.n1532 gnd 0.007744f
C4530 vdd.n1533 gnd 0.009621f
C4531 vdd.n1534 gnd 0.007744f
C4532 vdd.n1535 gnd 0.009621f
C4533 vdd.n1536 gnd 0.614504f
C4534 vdd.t37 gnd 0.491603f
C4535 vdd.n1537 gnd 0.009621f
C4536 vdd.n1538 gnd 0.007744f
C4537 vdd.n1539 gnd 0.009621f
C4538 vdd.n1540 gnd 0.007744f
C4539 vdd.n1541 gnd 0.009621f
C4540 vdd.t15 gnd 0.491603f
C4541 vdd.n1542 gnd 0.009621f
C4542 vdd.n1543 gnd 0.007744f
C4543 vdd.n1544 gnd 0.009621f
C4544 vdd.n1545 gnd 0.007744f
C4545 vdd.n1546 gnd 0.009621f
C4546 vdd.t23 gnd 0.491603f
C4547 vdd.n1547 gnd 0.535848f
C4548 vdd.n1548 gnd 0.009621f
C4549 vdd.n1549 gnd 0.007744f
C4550 vdd.n1550 gnd 0.009621f
C4551 vdd.n1551 gnd 0.007744f
C4552 vdd.n1552 gnd 0.009621f
C4553 vdd.t143 gnd 0.491603f
C4554 vdd.n1553 gnd 0.009621f
C4555 vdd.n1554 gnd 0.007744f
C4556 vdd.n1555 gnd 0.009621f
C4557 vdd.n1556 gnd 0.007744f
C4558 vdd.n1557 gnd 0.009621f
C4559 vdd.n1558 gnd 0.761985f
C4560 vdd.n1559 gnd 0.816061f
C4561 vdd.t27 gnd 0.491603f
C4562 vdd.n1560 gnd 0.009621f
C4563 vdd.n1561 gnd 0.007744f
C4564 vdd.n1562 gnd 0.009621f
C4565 vdd.n1563 gnd 0.007744f
C4566 vdd.n1564 gnd 0.009621f
C4567 vdd.n1565 gnd 0.59484f
C4568 vdd.n1566 gnd 0.009621f
C4569 vdd.n1567 gnd 0.007744f
C4570 vdd.n1568 gnd 0.009621f
C4571 vdd.n1569 gnd 0.007744f
C4572 vdd.n1570 gnd 0.009621f
C4573 vdd.t161 gnd 0.491603f
C4574 vdd.t61 gnd 0.491603f
C4575 vdd.n1571 gnd 0.009621f
C4576 vdd.n1572 gnd 0.007744f
C4577 vdd.n1573 gnd 0.009621f
C4578 vdd.n1574 gnd 0.007744f
C4579 vdd.n1575 gnd 0.009621f
C4580 vdd.t180 gnd 0.491603f
C4581 vdd.n1576 gnd 0.009621f
C4582 vdd.n1577 gnd 0.007744f
C4583 vdd.n1578 gnd 0.009621f
C4584 vdd.n1579 gnd 0.007744f
C4585 vdd.n1580 gnd 0.009621f
C4586 vdd.t182 gnd 0.491603f
C4587 vdd.n1581 gnd 0.722657f
C4588 vdd.n1582 gnd 0.009621f
C4589 vdd.n1583 gnd 0.007744f
C4590 vdd.n1584 gnd 0.009621f
C4591 vdd.n1585 gnd 0.007744f
C4592 vdd.n1586 gnd 0.009621f
C4593 vdd.n1587 gnd 0.983206f
C4594 vdd.n1588 gnd 0.009621f
C4595 vdd.n1589 gnd 0.007744f
C4596 vdd.n1590 gnd 0.009621f
C4597 vdd.n1591 gnd 0.007744f
C4598 vdd.n1592 gnd 0.009621f
C4599 vdd.n1593 gnd 0.830809f
C4600 vdd.n1594 gnd 0.009621f
C4601 vdd.n1595 gnd 0.007744f
C4602 vdd.n1596 gnd 0.021909f
C4603 vdd.n1597 gnd 0.006427f
C4604 vdd.n1598 gnd 0.021909f
C4605 vdd.n1599 gnd 1.29783f
C4606 vdd.n1600 gnd 0.021909f
C4607 vdd.n1601 gnd 0.006427f
C4608 vdd.n1602 gnd 0.009621f
C4609 vdd.t112 gnd 0.118362f
C4610 vdd.t113 gnd 0.126496f
C4611 vdd.t110 gnd 0.154579f
C4612 vdd.n1603 gnd 0.198149f
C4613 vdd.n1604 gnd 0.167255f
C4614 vdd.n1605 gnd 0.0127f
C4615 vdd.n1606 gnd 0.009621f
C4616 vdd.n1637 gnd 0.009621f
C4617 vdd.n1638 gnd 0.009621f
C4618 vdd.n1639 gnd 0.022059f
C4619 vdd.n1640 gnd 0.007744f
C4620 vdd.n1641 gnd 0.009621f
C4621 vdd.n1642 gnd 0.009621f
C4622 vdd.n1643 gnd 0.009621f
C4623 vdd.n1644 gnd 0.009621f
C4624 vdd.n1645 gnd 0.007744f
C4625 vdd.n1646 gnd 0.009621f
C4626 vdd.n1647 gnd 0.009621f
C4627 vdd.n1648 gnd 0.009621f
C4628 vdd.n1649 gnd 0.009621f
C4629 vdd.n1650 gnd 0.009621f
C4630 vdd.n1651 gnd 0.007744f
C4631 vdd.n1652 gnd 0.009621f
C4632 vdd.n1653 gnd 0.009621f
C4633 vdd.n1654 gnd 0.009621f
C4634 vdd.n1655 gnd 0.009621f
C4635 vdd.n1656 gnd 0.009621f
C4636 vdd.n1657 gnd 0.007744f
C4637 vdd.n1658 gnd 0.009621f
C4638 vdd.n1659 gnd 0.009621f
C4639 vdd.n1660 gnd 0.009621f
C4640 vdd.n1661 gnd 0.009621f
C4641 vdd.n1662 gnd 0.009621f
C4642 vdd.n1663 gnd 0.006466f
C4643 vdd.n1664 gnd 0.009621f
C4644 vdd.n1665 gnd 0.009621f
C4645 vdd.n1666 gnd 0.009621f
C4646 vdd.n1667 gnd 0.007744f
C4647 vdd.n1668 gnd 0.009621f
C4648 vdd.n1669 gnd 0.009621f
C4649 vdd.n1670 gnd 0.009621f
C4650 vdd.n1671 gnd 0.009621f
C4651 vdd.n1672 gnd 0.009621f
C4652 vdd.n1673 gnd 0.007744f
C4653 vdd.n1674 gnd 0.009621f
C4654 vdd.n1675 gnd 0.009621f
C4655 vdd.n1676 gnd 0.009621f
C4656 vdd.n1677 gnd 0.009621f
C4657 vdd.n1678 gnd 0.009621f
C4658 vdd.n1679 gnd 0.007744f
C4659 vdd.n1680 gnd 0.009621f
C4660 vdd.n1681 gnd 0.009621f
C4661 vdd.n1682 gnd 0.009621f
C4662 vdd.n1683 gnd 0.009621f
C4663 vdd.n1684 gnd 0.009621f
C4664 vdd.n1685 gnd 0.007744f
C4665 vdd.n1686 gnd 0.009621f
C4666 vdd.n1687 gnd 0.009621f
C4667 vdd.n1688 gnd 0.009621f
C4668 vdd.n1689 gnd 0.009621f
C4669 vdd.n1690 gnd 0.009621f
C4670 vdd.n1691 gnd 0.007744f
C4671 vdd.n1692 gnd 0.009621f
C4672 vdd.n1693 gnd 0.009621f
C4673 vdd.n1694 gnd 0.009621f
C4674 vdd.n1695 gnd 0.009621f
C4675 vdd.n1696 gnd 0.007666f
C4676 vdd.n1697 gnd 0.009621f
C4677 vdd.n1698 gnd 0.009621f
C4678 vdd.n1699 gnd 0.009621f
C4679 vdd.n1700 gnd 0.009621f
C4680 vdd.n1701 gnd 0.009621f
C4681 vdd.n1702 gnd 0.007744f
C4682 vdd.n1703 gnd 0.009621f
C4683 vdd.n1704 gnd 0.009621f
C4684 vdd.n1705 gnd 0.009621f
C4685 vdd.n1706 gnd 0.009621f
C4686 vdd.n1707 gnd 0.009621f
C4687 vdd.n1708 gnd 0.007744f
C4688 vdd.n1709 gnd 0.009621f
C4689 vdd.n1710 gnd 0.009621f
C4690 vdd.n1711 gnd 0.009621f
C4691 vdd.n1712 gnd 0.009621f
C4692 vdd.n1713 gnd 0.009621f
C4693 vdd.n1714 gnd 0.007744f
C4694 vdd.n1715 gnd 0.009621f
C4695 vdd.n1716 gnd 0.009621f
C4696 vdd.n1717 gnd 0.009621f
C4697 vdd.n1718 gnd 0.009621f
C4698 vdd.n1719 gnd 0.009621f
C4699 vdd.n1720 gnd 0.007744f
C4700 vdd.n1721 gnd 0.009621f
C4701 vdd.n1722 gnd 0.009621f
C4702 vdd.n1723 gnd 0.009621f
C4703 vdd.n1724 gnd 0.009621f
C4704 vdd.n1725 gnd 0.009621f
C4705 vdd.n1726 gnd 0.004065f
C4706 vdd.n1727 gnd 0.009621f
C4707 vdd.n1728 gnd 0.007744f
C4708 vdd.n1729 gnd 0.007744f
C4709 vdd.n1730 gnd 0.007744f
C4710 vdd.n1731 gnd 0.009621f
C4711 vdd.n1732 gnd 0.009621f
C4712 vdd.n1733 gnd 0.009621f
C4713 vdd.n1734 gnd 0.007744f
C4714 vdd.n1735 gnd 0.007744f
C4715 vdd.n1736 gnd 0.007744f
C4716 vdd.n1737 gnd 0.009621f
C4717 vdd.n1738 gnd 0.009621f
C4718 vdd.n1739 gnd 0.009621f
C4719 vdd.n1740 gnd 0.007744f
C4720 vdd.n1741 gnd 0.007744f
C4721 vdd.n1742 gnd 0.007744f
C4722 vdd.n1743 gnd 0.009621f
C4723 vdd.n1744 gnd 0.009621f
C4724 vdd.n1745 gnd 0.009621f
C4725 vdd.n1746 gnd 0.007744f
C4726 vdd.n1747 gnd 0.007744f
C4727 vdd.n1748 gnd 0.007744f
C4728 vdd.n1749 gnd 0.009621f
C4729 vdd.n1750 gnd 0.009621f
C4730 vdd.n1751 gnd 0.009621f
C4731 vdd.n1752 gnd 0.007744f
C4732 vdd.n1753 gnd 0.007744f
C4733 vdd.n1754 gnd 0.007744f
C4734 vdd.n1755 gnd 0.009621f
C4735 vdd.n1756 gnd 0.009621f
C4736 vdd.n1757 gnd 0.009621f
C4737 vdd.n1758 gnd 0.009621f
C4738 vdd.t126 gnd 0.118362f
C4739 vdd.t127 gnd 0.126496f
C4740 vdd.t125 gnd 0.154579f
C4741 vdd.n1759 gnd 0.198149f
C4742 vdd.n1760 gnd 0.167255f
C4743 vdd.n1761 gnd 0.016571f
C4744 vdd.n1762 gnd 0.005266f
C4745 vdd.n1763 gnd 0.007744f
C4746 vdd.n1764 gnd 0.009621f
C4747 vdd.n1765 gnd 0.009621f
C4748 vdd.n1766 gnd 0.009621f
C4749 vdd.n1767 gnd 0.007744f
C4750 vdd.n1768 gnd 0.007744f
C4751 vdd.n1769 gnd 0.007744f
C4752 vdd.n1770 gnd 0.009621f
C4753 vdd.n1771 gnd 0.009621f
C4754 vdd.n1772 gnd 0.009621f
C4755 vdd.n1773 gnd 0.007744f
C4756 vdd.n1774 gnd 0.007744f
C4757 vdd.n1775 gnd 0.007744f
C4758 vdd.n1776 gnd 0.009621f
C4759 vdd.n1777 gnd 0.009621f
C4760 vdd.n1778 gnd 0.009621f
C4761 vdd.n1779 gnd 0.007744f
C4762 vdd.n1780 gnd 0.007744f
C4763 vdd.n1781 gnd 0.007744f
C4764 vdd.n1782 gnd 0.009621f
C4765 vdd.n1783 gnd 0.009621f
C4766 vdd.n1784 gnd 0.009621f
C4767 vdd.n1785 gnd 0.007744f
C4768 vdd.n1786 gnd 0.007744f
C4769 vdd.n1787 gnd 0.007744f
C4770 vdd.n1788 gnd 0.009621f
C4771 vdd.n1789 gnd 0.009621f
C4772 vdd.n1790 gnd 0.009621f
C4773 vdd.n1791 gnd 0.007744f
C4774 vdd.n1792 gnd 0.006466f
C4775 vdd.n1793 gnd 0.009621f
C4776 vdd.n1794 gnd 0.009621f
C4777 vdd.t136 gnd 0.118362f
C4778 vdd.t137 gnd 0.126496f
C4779 vdd.t135 gnd 0.154579f
C4780 vdd.n1795 gnd 0.198149f
C4781 vdd.n1796 gnd 0.167255f
C4782 vdd.n1797 gnd 0.016571f
C4783 vdd.n1798 gnd 0.009621f
C4784 vdd.n1799 gnd 0.009621f
C4785 vdd.n1800 gnd 0.009621f
C4786 vdd.n1801 gnd 0.007744f
C4787 vdd.n1802 gnd 0.007744f
C4788 vdd.n1803 gnd 0.007744f
C4789 vdd.n1804 gnd 0.009621f
C4790 vdd.n1805 gnd 0.009621f
C4791 vdd.n1806 gnd 0.009621f
C4792 vdd.n1807 gnd 0.007744f
C4793 vdd.n1808 gnd 0.007744f
C4794 vdd.n1809 gnd 0.007744f
C4795 vdd.n1810 gnd 0.009621f
C4796 vdd.n1811 gnd 0.009621f
C4797 vdd.n1812 gnd 0.009621f
C4798 vdd.n1813 gnd 0.007744f
C4799 vdd.n1814 gnd 0.007744f
C4800 vdd.n1815 gnd 0.007744f
C4801 vdd.n1816 gnd 0.009621f
C4802 vdd.n1817 gnd 0.009621f
C4803 vdd.n1818 gnd 0.009621f
C4804 vdd.n1819 gnd 0.007744f
C4805 vdd.n1820 gnd 0.007744f
C4806 vdd.n1821 gnd 0.007744f
C4807 vdd.n1822 gnd 0.009621f
C4808 vdd.n1823 gnd 0.009621f
C4809 vdd.n1824 gnd 0.009621f
C4810 vdd.n1825 gnd 0.007744f
C4811 vdd.n1826 gnd 0.006427f
C4812 vdd.n1827 gnd 0.022059f
C4813 vdd.n1829 gnd 2.17289f
C4814 vdd.n1830 gnd 0.022059f
C4815 vdd.n1831 gnd 0.003678f
C4816 vdd.n1832 gnd 0.022059f
C4817 vdd.n1833 gnd 0.021909f
C4818 vdd.n1834 gnd 0.009621f
C4819 vdd.n1835 gnd 0.007744f
C4820 vdd.n1836 gnd 0.009621f
C4821 vdd.t111 gnd 0.491603f
C4822 vdd.n1837 gnd 0.644f
C4823 vdd.n1838 gnd 0.009621f
C4824 vdd.n1839 gnd 0.007744f
C4825 vdd.n1840 gnd 0.009621f
C4826 vdd.n1841 gnd 0.009621f
C4827 vdd.n1842 gnd 0.009621f
C4828 vdd.n1843 gnd 0.007744f
C4829 vdd.n1844 gnd 0.009621f
C4830 vdd.n1845 gnd 0.983206f
C4831 vdd.n1846 gnd 0.009621f
C4832 vdd.n1847 gnd 0.007744f
C4833 vdd.n1848 gnd 0.009621f
C4834 vdd.n1849 gnd 0.009621f
C4835 vdd.n1850 gnd 0.009621f
C4836 vdd.n1851 gnd 0.007744f
C4837 vdd.n1852 gnd 0.009621f
C4838 vdd.n1853 gnd 0.816061f
C4839 vdd.t47 gnd 0.491603f
C4840 vdd.n1854 gnd 0.565344f
C4841 vdd.n1855 gnd 0.009621f
C4842 vdd.n1856 gnd 0.007744f
C4843 vdd.n1857 gnd 0.009621f
C4844 vdd.n1858 gnd 0.009621f
C4845 vdd.n1859 gnd 0.009621f
C4846 vdd.n1860 gnd 0.007744f
C4847 vdd.n1861 gnd 0.009621f
C4848 vdd.n1862 gnd 0.585008f
C4849 vdd.n1863 gnd 0.009621f
C4850 vdd.n1864 gnd 0.007744f
C4851 vdd.n1865 gnd 0.009621f
C4852 vdd.n1866 gnd 0.009621f
C4853 vdd.n1867 gnd 0.009621f
C4854 vdd.n1868 gnd 0.007744f
C4855 vdd.n1869 gnd 0.009621f
C4856 vdd.n1870 gnd 0.555512f
C4857 vdd.n1871 gnd 0.752153f
C4858 vdd.n1872 gnd 0.009621f
C4859 vdd.n1873 gnd 0.007744f
C4860 vdd.n1874 gnd 0.009621f
C4861 vdd.n1875 gnd 0.009621f
C4862 vdd.n1876 gnd 0.009621f
C4863 vdd.n1877 gnd 0.007744f
C4864 vdd.n1878 gnd 0.009621f
C4865 vdd.n1879 gnd 0.816061f
C4866 vdd.n1880 gnd 0.009621f
C4867 vdd.n1881 gnd 0.007744f
C4868 vdd.n1882 gnd 0.009621f
C4869 vdd.n1883 gnd 0.009621f
C4870 vdd.n1884 gnd 0.009621f
C4871 vdd.n1885 gnd 0.007744f
C4872 vdd.n1886 gnd 0.009621f
C4873 vdd.t17 gnd 0.491603f
C4874 vdd.n1887 gnd 0.712825f
C4875 vdd.n1888 gnd 0.009621f
C4876 vdd.n1889 gnd 0.007744f
C4877 vdd.n1890 gnd 0.009621f
C4878 vdd.n1891 gnd 0.009621f
C4879 vdd.n1892 gnd 0.009621f
C4880 vdd.n1893 gnd 0.007744f
C4881 vdd.n1894 gnd 0.009621f
C4882 vdd.n1895 gnd 0.54568f
C4883 vdd.n1896 gnd 0.009621f
C4884 vdd.n1897 gnd 0.007744f
C4885 vdd.n1898 gnd 0.009621f
C4886 vdd.n1899 gnd 0.009621f
C4887 vdd.n1900 gnd 0.009621f
C4888 vdd.n1901 gnd 0.007744f
C4889 vdd.n1902 gnd 0.009621f
C4890 vdd.n1903 gnd 0.702993f
C4891 vdd.n1904 gnd 0.604672f
C4892 vdd.n1905 gnd 0.009621f
C4893 vdd.n1906 gnd 0.007744f
C4894 vdd.n1907 gnd 0.007394f
C4895 vdd.n1908 gnd 0.00528f
C4896 vdd.n1909 gnd 0.0049f
C4897 vdd.n1910 gnd 0.00271f
C4898 vdd.n1911 gnd 0.006223f
C4899 vdd.n1912 gnd 0.002633f
C4900 vdd.n1913 gnd 0.002788f
C4901 vdd.n1914 gnd 0.0049f
C4902 vdd.n1915 gnd 0.002633f
C4903 vdd.n1916 gnd 0.006223f
C4904 vdd.n1917 gnd 0.002788f
C4905 vdd.n1918 gnd 0.0049f
C4906 vdd.n1919 gnd 0.002633f
C4907 vdd.n1920 gnd 0.004667f
C4908 vdd.n1921 gnd 0.004681f
C4909 vdd.t174 gnd 0.01337f
C4910 vdd.n1922 gnd 0.029747f
C4911 vdd.n1923 gnd 0.154813f
C4912 vdd.n1924 gnd 0.002633f
C4913 vdd.n1925 gnd 0.002788f
C4914 vdd.n1926 gnd 0.006223f
C4915 vdd.n1927 gnd 0.006223f
C4916 vdd.n1928 gnd 0.002788f
C4917 vdd.n1929 gnd 0.002633f
C4918 vdd.n1930 gnd 0.0049f
C4919 vdd.n1931 gnd 0.0049f
C4920 vdd.n1932 gnd 0.002633f
C4921 vdd.n1933 gnd 0.002788f
C4922 vdd.n1934 gnd 0.006223f
C4923 vdd.n1935 gnd 0.006223f
C4924 vdd.n1936 gnd 0.002788f
C4925 vdd.n1937 gnd 0.002633f
C4926 vdd.n1938 gnd 0.0049f
C4927 vdd.n1939 gnd 0.0049f
C4928 vdd.n1940 gnd 0.002633f
C4929 vdd.n1941 gnd 0.002788f
C4930 vdd.n1942 gnd 0.006223f
C4931 vdd.n1943 gnd 0.006223f
C4932 vdd.n1944 gnd 0.014713f
C4933 vdd.n1945 gnd 0.00271f
C4934 vdd.n1946 gnd 0.002633f
C4935 vdd.n1947 gnd 0.012664f
C4936 vdd.n1948 gnd 0.008841f
C4937 vdd.t178 gnd 0.030974f
C4938 vdd.t5 gnd 0.030974f
C4939 vdd.n1949 gnd 0.212878f
C4940 vdd.n1950 gnd 0.167396f
C4941 vdd.t257 gnd 0.030974f
C4942 vdd.t20 gnd 0.030974f
C4943 vdd.n1951 gnd 0.212878f
C4944 vdd.n1952 gnd 0.135088f
C4945 vdd.t189 gnd 0.030974f
C4946 vdd.t58 gnd 0.030974f
C4947 vdd.n1953 gnd 0.212878f
C4948 vdd.n1954 gnd 0.135088f
C4949 vdd.t190 gnd 0.030974f
C4950 vdd.t45 gnd 0.030974f
C4951 vdd.n1955 gnd 0.212878f
C4952 vdd.n1956 gnd 0.135088f
C4953 vdd.t145 gnd 0.030974f
C4954 vdd.t28 gnd 0.030974f
C4955 vdd.n1957 gnd 0.212878f
C4956 vdd.n1958 gnd 0.135088f
C4957 vdd.t162 gnd 0.030974f
C4958 vdd.t62 gnd 0.030974f
C4959 vdd.n1959 gnd 0.212878f
C4960 vdd.n1960 gnd 0.135088f
C4961 vdd.t183 gnd 0.030974f
C4962 vdd.t254 gnd 0.030974f
C4963 vdd.n1961 gnd 0.212878f
C4964 vdd.n1962 gnd 0.135088f
C4965 vdd.n1963 gnd 0.00528f
C4966 vdd.n1964 gnd 0.0049f
C4967 vdd.n1965 gnd 0.00271f
C4968 vdd.n1966 gnd 0.006223f
C4969 vdd.n1967 gnd 0.002633f
C4970 vdd.n1968 gnd 0.002788f
C4971 vdd.n1969 gnd 0.0049f
C4972 vdd.n1970 gnd 0.002633f
C4973 vdd.n1971 gnd 0.006223f
C4974 vdd.n1972 gnd 0.002788f
C4975 vdd.n1973 gnd 0.0049f
C4976 vdd.n1974 gnd 0.002633f
C4977 vdd.n1975 gnd 0.004667f
C4978 vdd.n1976 gnd 0.004681f
C4979 vdd.t168 gnd 0.01337f
C4980 vdd.n1977 gnd 0.029747f
C4981 vdd.n1978 gnd 0.154813f
C4982 vdd.n1979 gnd 0.002633f
C4983 vdd.n1980 gnd 0.002788f
C4984 vdd.n1981 gnd 0.006223f
C4985 vdd.n1982 gnd 0.006223f
C4986 vdd.n1983 gnd 0.002788f
C4987 vdd.n1984 gnd 0.002633f
C4988 vdd.n1985 gnd 0.0049f
C4989 vdd.n1986 gnd 0.0049f
C4990 vdd.n1987 gnd 0.002633f
C4991 vdd.n1988 gnd 0.002788f
C4992 vdd.n1989 gnd 0.006223f
C4993 vdd.n1990 gnd 0.006223f
C4994 vdd.n1991 gnd 0.002788f
C4995 vdd.n1992 gnd 0.002633f
C4996 vdd.n1993 gnd 0.0049f
C4997 vdd.n1994 gnd 0.0049f
C4998 vdd.n1995 gnd 0.002633f
C4999 vdd.n1996 gnd 0.002788f
C5000 vdd.n1997 gnd 0.006223f
C5001 vdd.n1998 gnd 0.006223f
C5002 vdd.n1999 gnd 0.014713f
C5003 vdd.n2000 gnd 0.00271f
C5004 vdd.n2001 gnd 0.002633f
C5005 vdd.n2002 gnd 0.012664f
C5006 vdd.n2003 gnd 0.008564f
C5007 vdd.n2004 gnd 0.100506f
C5008 vdd.n2005 gnd 0.00528f
C5009 vdd.n2006 gnd 0.0049f
C5010 vdd.n2007 gnd 0.00271f
C5011 vdd.n2008 gnd 0.006223f
C5012 vdd.n2009 gnd 0.002633f
C5013 vdd.n2010 gnd 0.002788f
C5014 vdd.n2011 gnd 0.0049f
C5015 vdd.n2012 gnd 0.002633f
C5016 vdd.n2013 gnd 0.006223f
C5017 vdd.n2014 gnd 0.002788f
C5018 vdd.n2015 gnd 0.0049f
C5019 vdd.n2016 gnd 0.002633f
C5020 vdd.n2017 gnd 0.004667f
C5021 vdd.n2018 gnd 0.004681f
C5022 vdd.t185 gnd 0.01337f
C5023 vdd.n2019 gnd 0.029747f
C5024 vdd.n2020 gnd 0.154813f
C5025 vdd.n2021 gnd 0.002633f
C5026 vdd.n2022 gnd 0.002788f
C5027 vdd.n2023 gnd 0.006223f
C5028 vdd.n2024 gnd 0.006223f
C5029 vdd.n2025 gnd 0.002788f
C5030 vdd.n2026 gnd 0.002633f
C5031 vdd.n2027 gnd 0.0049f
C5032 vdd.n2028 gnd 0.0049f
C5033 vdd.n2029 gnd 0.002633f
C5034 vdd.n2030 gnd 0.002788f
C5035 vdd.n2031 gnd 0.006223f
C5036 vdd.n2032 gnd 0.006223f
C5037 vdd.n2033 gnd 0.002788f
C5038 vdd.n2034 gnd 0.002633f
C5039 vdd.n2035 gnd 0.0049f
C5040 vdd.n2036 gnd 0.0049f
C5041 vdd.n2037 gnd 0.002633f
C5042 vdd.n2038 gnd 0.002788f
C5043 vdd.n2039 gnd 0.006223f
C5044 vdd.n2040 gnd 0.006223f
C5045 vdd.n2041 gnd 0.014713f
C5046 vdd.n2042 gnd 0.00271f
C5047 vdd.n2043 gnd 0.002633f
C5048 vdd.n2044 gnd 0.012664f
C5049 vdd.n2045 gnd 0.008841f
C5050 vdd.t176 gnd 0.030974f
C5051 vdd.t26 gnd 0.030974f
C5052 vdd.n2046 gnd 0.212878f
C5053 vdd.n2047 gnd 0.167396f
C5054 vdd.t274 gnd 0.030974f
C5055 vdd.t151 gnd 0.030974f
C5056 vdd.n2048 gnd 0.212878f
C5057 vdd.n2049 gnd 0.135088f
C5058 vdd.t16 gnd 0.030974f
C5059 vdd.t3 gnd 0.030974f
C5060 vdd.n2050 gnd 0.212878f
C5061 vdd.n2051 gnd 0.135088f
C5062 vdd.t187 gnd 0.030974f
C5063 vdd.t260 gnd 0.030974f
C5064 vdd.n2052 gnd 0.212878f
C5065 vdd.n2053 gnd 0.135088f
C5066 vdd.t18 gnd 0.030974f
C5067 vdd.t256 gnd 0.030974f
C5068 vdd.n2054 gnd 0.212878f
C5069 vdd.n2055 gnd 0.135088f
C5070 vdd.t253 gnd 0.030974f
C5071 vdd.t268 gnd 0.030974f
C5072 vdd.n2056 gnd 0.212878f
C5073 vdd.n2057 gnd 0.135088f
C5074 vdd.t184 gnd 0.030974f
C5075 vdd.t266 gnd 0.030974f
C5076 vdd.n2058 gnd 0.212878f
C5077 vdd.n2059 gnd 0.135088f
C5078 vdd.n2060 gnd 0.00528f
C5079 vdd.n2061 gnd 0.0049f
C5080 vdd.n2062 gnd 0.00271f
C5081 vdd.n2063 gnd 0.006223f
C5082 vdd.n2064 gnd 0.002633f
C5083 vdd.n2065 gnd 0.002788f
C5084 vdd.n2066 gnd 0.0049f
C5085 vdd.n2067 gnd 0.002633f
C5086 vdd.n2068 gnd 0.006223f
C5087 vdd.n2069 gnd 0.002788f
C5088 vdd.n2070 gnd 0.0049f
C5089 vdd.n2071 gnd 0.002633f
C5090 vdd.n2072 gnd 0.004667f
C5091 vdd.n2073 gnd 0.004681f
C5092 vdd.t177 gnd 0.01337f
C5093 vdd.n2074 gnd 0.029747f
C5094 vdd.n2075 gnd 0.154813f
C5095 vdd.n2076 gnd 0.002633f
C5096 vdd.n2077 gnd 0.002788f
C5097 vdd.n2078 gnd 0.006223f
C5098 vdd.n2079 gnd 0.006223f
C5099 vdd.n2080 gnd 0.002788f
C5100 vdd.n2081 gnd 0.002633f
C5101 vdd.n2082 gnd 0.0049f
C5102 vdd.n2083 gnd 0.0049f
C5103 vdd.n2084 gnd 0.002633f
C5104 vdd.n2085 gnd 0.002788f
C5105 vdd.n2086 gnd 0.006223f
C5106 vdd.n2087 gnd 0.006223f
C5107 vdd.n2088 gnd 0.002788f
C5108 vdd.n2089 gnd 0.002633f
C5109 vdd.n2090 gnd 0.0049f
C5110 vdd.n2091 gnd 0.0049f
C5111 vdd.n2092 gnd 0.002633f
C5112 vdd.n2093 gnd 0.002788f
C5113 vdd.n2094 gnd 0.006223f
C5114 vdd.n2095 gnd 0.006223f
C5115 vdd.n2096 gnd 0.014713f
C5116 vdd.n2097 gnd 0.00271f
C5117 vdd.n2098 gnd 0.002633f
C5118 vdd.n2099 gnd 0.012664f
C5119 vdd.n2100 gnd 0.008564f
C5120 vdd.n2101 gnd 0.059791f
C5121 vdd.n2102 gnd 0.215442f
C5122 vdd.n2103 gnd 0.00528f
C5123 vdd.n2104 gnd 0.0049f
C5124 vdd.n2105 gnd 0.00271f
C5125 vdd.n2106 gnd 0.006223f
C5126 vdd.n2107 gnd 0.002633f
C5127 vdd.n2108 gnd 0.002788f
C5128 vdd.n2109 gnd 0.0049f
C5129 vdd.n2110 gnd 0.002633f
C5130 vdd.n2111 gnd 0.006223f
C5131 vdd.n2112 gnd 0.002788f
C5132 vdd.n2113 gnd 0.0049f
C5133 vdd.n2114 gnd 0.002633f
C5134 vdd.n2115 gnd 0.004667f
C5135 vdd.n2116 gnd 0.004681f
C5136 vdd.t166 gnd 0.01337f
C5137 vdd.n2117 gnd 0.029747f
C5138 vdd.n2118 gnd 0.154813f
C5139 vdd.n2119 gnd 0.002633f
C5140 vdd.n2120 gnd 0.002788f
C5141 vdd.n2121 gnd 0.006223f
C5142 vdd.n2122 gnd 0.006223f
C5143 vdd.n2123 gnd 0.002788f
C5144 vdd.n2124 gnd 0.002633f
C5145 vdd.n2125 gnd 0.0049f
C5146 vdd.n2126 gnd 0.0049f
C5147 vdd.n2127 gnd 0.002633f
C5148 vdd.n2128 gnd 0.002788f
C5149 vdd.n2129 gnd 0.006223f
C5150 vdd.n2130 gnd 0.006223f
C5151 vdd.n2131 gnd 0.002788f
C5152 vdd.n2132 gnd 0.002633f
C5153 vdd.n2133 gnd 0.0049f
C5154 vdd.n2134 gnd 0.0049f
C5155 vdd.n2135 gnd 0.002633f
C5156 vdd.n2136 gnd 0.002788f
C5157 vdd.n2137 gnd 0.006223f
C5158 vdd.n2138 gnd 0.006223f
C5159 vdd.n2139 gnd 0.014713f
C5160 vdd.n2140 gnd 0.00271f
C5161 vdd.n2141 gnd 0.002633f
C5162 vdd.n2142 gnd 0.012664f
C5163 vdd.n2143 gnd 0.008841f
C5164 vdd.t32 gnd 0.030974f
C5165 vdd.t46 gnd 0.030974f
C5166 vdd.n2144 gnd 0.212878f
C5167 vdd.n2145 gnd 0.167396f
C5168 vdd.t38 gnd 0.030974f
C5169 vdd.t55 gnd 0.030974f
C5170 vdd.n2146 gnd 0.212878f
C5171 vdd.n2147 gnd 0.135088f
C5172 vdd.t25 gnd 0.030974f
C5173 vdd.t167 gnd 0.030974f
C5174 vdd.n2148 gnd 0.212878f
C5175 vdd.n2149 gnd 0.135088f
C5176 vdd.t144 gnd 0.030974f
C5177 vdd.t24 gnd 0.030974f
C5178 vdd.n2150 gnd 0.212878f
C5179 vdd.n2151 gnd 0.135088f
C5180 vdd.t41 gnd 0.030974f
C5181 vdd.t265 gnd 0.030974f
C5182 vdd.n2152 gnd 0.212878f
C5183 vdd.n2153 gnd 0.135088f
C5184 vdd.t270 gnd 0.030974f
C5185 vdd.t251 gnd 0.030974f
C5186 vdd.n2154 gnd 0.212878f
C5187 vdd.n2155 gnd 0.135088f
C5188 vdd.t186 gnd 0.030974f
C5189 vdd.t181 gnd 0.030974f
C5190 vdd.n2156 gnd 0.212878f
C5191 vdd.n2157 gnd 0.135088f
C5192 vdd.n2158 gnd 0.00528f
C5193 vdd.n2159 gnd 0.0049f
C5194 vdd.n2160 gnd 0.00271f
C5195 vdd.n2161 gnd 0.006223f
C5196 vdd.n2162 gnd 0.002633f
C5197 vdd.n2163 gnd 0.002788f
C5198 vdd.n2164 gnd 0.0049f
C5199 vdd.n2165 gnd 0.002633f
C5200 vdd.n2166 gnd 0.006223f
C5201 vdd.n2167 gnd 0.002788f
C5202 vdd.n2168 gnd 0.0049f
C5203 vdd.n2169 gnd 0.002633f
C5204 vdd.n2170 gnd 0.004667f
C5205 vdd.n2171 gnd 0.004681f
C5206 vdd.t48 gnd 0.01337f
C5207 vdd.n2172 gnd 0.029747f
C5208 vdd.n2173 gnd 0.154813f
C5209 vdd.n2174 gnd 0.002633f
C5210 vdd.n2175 gnd 0.002788f
C5211 vdd.n2176 gnd 0.006223f
C5212 vdd.n2177 gnd 0.006223f
C5213 vdd.n2178 gnd 0.002788f
C5214 vdd.n2179 gnd 0.002633f
C5215 vdd.n2180 gnd 0.0049f
C5216 vdd.n2181 gnd 0.0049f
C5217 vdd.n2182 gnd 0.002633f
C5218 vdd.n2183 gnd 0.002788f
C5219 vdd.n2184 gnd 0.006223f
C5220 vdd.n2185 gnd 0.006223f
C5221 vdd.n2186 gnd 0.002788f
C5222 vdd.n2187 gnd 0.002633f
C5223 vdd.n2188 gnd 0.0049f
C5224 vdd.n2189 gnd 0.0049f
C5225 vdd.n2190 gnd 0.002633f
C5226 vdd.n2191 gnd 0.002788f
C5227 vdd.n2192 gnd 0.006223f
C5228 vdd.n2193 gnd 0.006223f
C5229 vdd.n2194 gnd 0.014713f
C5230 vdd.n2195 gnd 0.00271f
C5231 vdd.n2196 gnd 0.002633f
C5232 vdd.n2197 gnd 0.012664f
C5233 vdd.n2198 gnd 0.008564f
C5234 vdd.n2199 gnd 0.059791f
C5235 vdd.n2200 gnd 0.241267f
C5236 vdd.n2201 gnd 2.6504f
C5237 vdd.n2202 gnd 0.567475f
C5238 vdd.n2203 gnd 0.007394f
C5239 vdd.n2204 gnd 0.009621f
C5240 vdd.n2205 gnd 0.007744f
C5241 vdd.n2206 gnd 0.009621f
C5242 vdd.n2207 gnd 0.771817f
C5243 vdd.n2208 gnd 0.009621f
C5244 vdd.n2209 gnd 0.007744f
C5245 vdd.n2210 gnd 0.009621f
C5246 vdd.n2211 gnd 0.009621f
C5247 vdd.n2212 gnd 0.009621f
C5248 vdd.n2213 gnd 0.007744f
C5249 vdd.n2214 gnd 0.009621f
C5250 vdd.t2 gnd 0.491603f
C5251 vdd.n2215 gnd 0.816061f
C5252 vdd.n2216 gnd 0.009621f
C5253 vdd.n2217 gnd 0.007744f
C5254 vdd.n2218 gnd 0.009621f
C5255 vdd.n2219 gnd 0.009621f
C5256 vdd.n2220 gnd 0.009621f
C5257 vdd.n2221 gnd 0.007744f
C5258 vdd.n2222 gnd 0.009621f
C5259 vdd.n2223 gnd 0.693161f
C5260 vdd.n2224 gnd 0.009621f
C5261 vdd.n2225 gnd 0.007744f
C5262 vdd.n2226 gnd 0.009621f
C5263 vdd.n2227 gnd 0.009621f
C5264 vdd.n2228 gnd 0.009621f
C5265 vdd.n2229 gnd 0.007744f
C5266 vdd.n2230 gnd 0.009621f
C5267 vdd.n2231 gnd 0.816061f
C5268 vdd.t19 gnd 0.491603f
C5269 vdd.n2232 gnd 0.526015f
C5270 vdd.n2233 gnd 0.009621f
C5271 vdd.n2234 gnd 0.007744f
C5272 vdd.n2235 gnd 0.009621f
C5273 vdd.n2236 gnd 0.009621f
C5274 vdd.n2237 gnd 0.009621f
C5275 vdd.n2238 gnd 0.007744f
C5276 vdd.n2239 gnd 0.009621f
C5277 vdd.n2240 gnd 0.624336f
C5278 vdd.n2241 gnd 0.009621f
C5279 vdd.n2242 gnd 0.007744f
C5280 vdd.n2243 gnd 0.009621f
C5281 vdd.n2244 gnd 0.009621f
C5282 vdd.n2245 gnd 0.009621f
C5283 vdd.n2246 gnd 0.007744f
C5284 vdd.n2247 gnd 0.009621f
C5285 vdd.n2248 gnd 0.516183f
C5286 vdd.n2249 gnd 0.791481f
C5287 vdd.n2250 gnd 0.009621f
C5288 vdd.n2251 gnd 0.007744f
C5289 vdd.n2252 gnd 0.009621f
C5290 vdd.n2253 gnd 0.009621f
C5291 vdd.n2254 gnd 0.009621f
C5292 vdd.n2255 gnd 0.007744f
C5293 vdd.n2256 gnd 0.009621f
C5294 vdd.n2257 gnd 0.958626f
C5295 vdd.n2258 gnd 0.009621f
C5296 vdd.n2259 gnd 0.007744f
C5297 vdd.n2260 gnd 0.009621f
C5298 vdd.n2261 gnd 0.009621f
C5299 vdd.n2262 gnd 0.021909f
C5300 vdd.n2263 gnd 0.009621f
C5301 vdd.n2264 gnd 0.009621f
C5302 vdd.n2265 gnd 0.007744f
C5303 vdd.n2266 gnd 0.009621f
C5304 vdd.t74 gnd 0.491603f
C5305 vdd.n2267 gnd 0.92913f
C5306 vdd.n2268 gnd 0.009621f
C5307 vdd.n2269 gnd 0.007744f
C5308 vdd.n2270 gnd 0.009621f
C5309 vdd.n2271 gnd 0.009621f
C5310 vdd.n2272 gnd 0.021909f
C5311 vdd.n2273 gnd 0.006427f
C5312 vdd.n2274 gnd 0.021909f
C5313 vdd.n2275 gnd 1.29783f
C5314 vdd.n2276 gnd 0.021909f
C5315 vdd.n2277 gnd 0.022059f
C5316 vdd.n2278 gnd 0.003678f
C5317 vdd.t97 gnd 0.118362f
C5318 vdd.t96 gnd 0.126496f
C5319 vdd.t95 gnd 0.154579f
C5320 vdd.n2279 gnd 0.198149f
C5321 vdd.n2280 gnd 0.166481f
C5322 vdd.n2281 gnd 0.011925f
C5323 vdd.n2282 gnd 0.004065f
C5324 vdd.n2283 gnd 0.008274f
C5325 vdd.n2284 gnd 1.02135f
C5326 vdd.n2286 gnd 0.007744f
C5327 vdd.n2287 gnd 0.007744f
C5328 vdd.n2288 gnd 0.009621f
C5329 vdd.n2290 gnd 0.009621f
C5330 vdd.n2291 gnd 0.009621f
C5331 vdd.n2292 gnd 0.007744f
C5332 vdd.n2293 gnd 0.007744f
C5333 vdd.n2294 gnd 0.007744f
C5334 vdd.n2295 gnd 0.009621f
C5335 vdd.n2297 gnd 0.009621f
C5336 vdd.n2298 gnd 0.009621f
C5337 vdd.n2299 gnd 0.007744f
C5338 vdd.n2300 gnd 0.007744f
C5339 vdd.n2301 gnd 0.007744f
C5340 vdd.n2302 gnd 0.009621f
C5341 vdd.n2304 gnd 0.009621f
C5342 vdd.n2305 gnd 0.009621f
C5343 vdd.n2306 gnd 0.007744f
C5344 vdd.n2307 gnd 0.007744f
C5345 vdd.n2308 gnd 0.007744f
C5346 vdd.n2309 gnd 0.009621f
C5347 vdd.n2311 gnd 0.009621f
C5348 vdd.n2312 gnd 0.009621f
C5349 vdd.n2313 gnd 0.007744f
C5350 vdd.n2314 gnd 0.009621f
C5351 vdd.n2315 gnd 0.009621f
C5352 vdd.n2316 gnd 0.009621f
C5353 vdd.n2317 gnd 0.015797f
C5354 vdd.n2318 gnd 0.005266f
C5355 vdd.n2319 gnd 0.007744f
C5356 vdd.n2320 gnd 0.009621f
C5357 vdd.n2322 gnd 0.009621f
C5358 vdd.n2323 gnd 0.009621f
C5359 vdd.n2324 gnd 0.007744f
C5360 vdd.n2325 gnd 0.007744f
C5361 vdd.n2326 gnd 0.007744f
C5362 vdd.n2327 gnd 0.009621f
C5363 vdd.n2329 gnd 0.009621f
C5364 vdd.n2330 gnd 0.009621f
C5365 vdd.n2331 gnd 0.007744f
C5366 vdd.n2332 gnd 0.007744f
C5367 vdd.n2333 gnd 0.007744f
C5368 vdd.n2334 gnd 0.009621f
C5369 vdd.n2336 gnd 0.009621f
C5370 vdd.n2337 gnd 0.009621f
C5371 vdd.n2338 gnd 0.007744f
C5372 vdd.n2339 gnd 0.007744f
C5373 vdd.n2340 gnd 0.007744f
C5374 vdd.n2341 gnd 0.009621f
C5375 vdd.n2343 gnd 0.009621f
C5376 vdd.n2344 gnd 0.009621f
C5377 vdd.n2345 gnd 0.007744f
C5378 vdd.n2346 gnd 0.007744f
C5379 vdd.n2347 gnd 0.007744f
C5380 vdd.n2348 gnd 0.009621f
C5381 vdd.n2350 gnd 0.009621f
C5382 vdd.n2351 gnd 0.009621f
C5383 vdd.n2352 gnd 0.007744f
C5384 vdd.n2353 gnd 0.009621f
C5385 vdd.n2354 gnd 0.009621f
C5386 vdd.n2355 gnd 0.009621f
C5387 vdd.n2356 gnd 0.015797f
C5388 vdd.n2357 gnd 0.006466f
C5389 vdd.n2358 gnd 0.007744f
C5390 vdd.n2359 gnd 0.009621f
C5391 vdd.n2361 gnd 0.009621f
C5392 vdd.n2362 gnd 0.009621f
C5393 vdd.n2363 gnd 0.007744f
C5394 vdd.n2364 gnd 0.007744f
C5395 vdd.n2365 gnd 0.007744f
C5396 vdd.n2366 gnd 0.009621f
C5397 vdd.n2368 gnd 0.009621f
C5398 vdd.n2369 gnd 0.009621f
C5399 vdd.n2370 gnd 0.007744f
C5400 vdd.n2371 gnd 0.007744f
C5401 vdd.n2372 gnd 0.007744f
C5402 vdd.n2373 gnd 0.009621f
C5403 vdd.n2375 gnd 0.009621f
C5404 vdd.n2376 gnd 0.009621f
C5405 vdd.n2377 gnd 0.007744f
C5406 vdd.n2378 gnd 0.007744f
C5407 vdd.n2379 gnd 0.007744f
C5408 vdd.n2380 gnd 0.009621f
C5409 vdd.n2382 gnd 0.009621f
C5410 vdd.n2383 gnd 0.007744f
C5411 vdd.n2384 gnd 0.007744f
C5412 vdd.n2385 gnd 0.009621f
C5413 vdd.n2387 gnd 0.009621f
C5414 vdd.n2388 gnd 0.009621f
C5415 vdd.n2389 gnd 0.007744f
C5416 vdd.n2390 gnd 0.008274f
C5417 vdd.n2391 gnd 1.02135f
C5418 vdd.n2392 gnd 0.044072f
C5419 vdd.n2393 gnd 0.006542f
C5420 vdd.n2394 gnd 0.006542f
C5421 vdd.n2395 gnd 0.006542f
C5422 vdd.n2396 gnd 0.006542f
C5423 vdd.n2397 gnd 0.006542f
C5424 vdd.n2398 gnd 0.006542f
C5425 vdd.n2399 gnd 0.006542f
C5426 vdd.n2400 gnd 0.006542f
C5427 vdd.n2401 gnd 0.006542f
C5428 vdd.n2402 gnd 0.006542f
C5429 vdd.n2403 gnd 0.006542f
C5430 vdd.n2404 gnd 0.006542f
C5431 vdd.n2405 gnd 0.006542f
C5432 vdd.n2406 gnd 0.006542f
C5433 vdd.n2407 gnd 0.006542f
C5434 vdd.n2408 gnd 0.006542f
C5435 vdd.n2409 gnd 0.006542f
C5436 vdd.n2410 gnd 0.006542f
C5437 vdd.n2411 gnd 0.006542f
C5438 vdd.n2412 gnd 0.006542f
C5439 vdd.n2413 gnd 0.006542f
C5440 vdd.n2414 gnd 0.006542f
C5441 vdd.n2415 gnd 0.006542f
C5442 vdd.n2416 gnd 0.006542f
C5443 vdd.n2417 gnd 0.006542f
C5444 vdd.n2418 gnd 0.006542f
C5445 vdd.n2419 gnd 0.006542f
C5446 vdd.n2420 gnd 0.006542f
C5447 vdd.n2421 gnd 0.006542f
C5448 vdd.n2422 gnd 0.006542f
C5449 vdd.n2423 gnd 11.6117f
C5450 vdd.n2425 gnd 0.014855f
C5451 vdd.n2426 gnd 0.014855f
C5452 vdd.n2427 gnd 0.014008f
C5453 vdd.n2428 gnd 0.006542f
C5454 vdd.n2429 gnd 0.006542f
C5455 vdd.n2430 gnd 0.66858f
C5456 vdd.n2431 gnd 0.006542f
C5457 vdd.n2432 gnd 0.006542f
C5458 vdd.n2433 gnd 0.006542f
C5459 vdd.n2434 gnd 0.006542f
C5460 vdd.n2435 gnd 0.006542f
C5461 vdd.n2436 gnd 0.526015f
C5462 vdd.n2437 gnd 0.006542f
C5463 vdd.n2438 gnd 0.006542f
C5464 vdd.n2439 gnd 0.006542f
C5465 vdd.n2440 gnd 0.006542f
C5466 vdd.n2441 gnd 0.006542f
C5467 vdd.n2442 gnd 0.66858f
C5468 vdd.n2443 gnd 0.006542f
C5469 vdd.n2444 gnd 0.006542f
C5470 vdd.n2445 gnd 0.006542f
C5471 vdd.n2446 gnd 0.006542f
C5472 vdd.n2447 gnd 0.006542f
C5473 vdd.n2448 gnd 0.66858f
C5474 vdd.n2449 gnd 0.006542f
C5475 vdd.n2450 gnd 0.006542f
C5476 vdd.n2451 gnd 0.006542f
C5477 vdd.n2452 gnd 0.006542f
C5478 vdd.n2453 gnd 0.006542f
C5479 vdd.n2454 gnd 0.644f
C5480 vdd.n2455 gnd 0.006542f
C5481 vdd.n2456 gnd 0.006542f
C5482 vdd.n2457 gnd 0.006542f
C5483 vdd.n2458 gnd 0.006542f
C5484 vdd.n2459 gnd 0.006542f
C5485 vdd.n2460 gnd 0.496519f
C5486 vdd.n2461 gnd 0.006542f
C5487 vdd.n2462 gnd 0.006542f
C5488 vdd.n2463 gnd 0.006542f
C5489 vdd.n2464 gnd 0.006542f
C5490 vdd.n2465 gnd 0.006542f
C5491 vdd.n2466 gnd 0.349038f
C5492 vdd.n2467 gnd 0.006542f
C5493 vdd.n2468 gnd 0.006542f
C5494 vdd.n2469 gnd 0.006542f
C5495 vdd.n2470 gnd 0.006542f
C5496 vdd.n2471 gnd 0.006542f
C5497 vdd.n2472 gnd 0.467023f
C5498 vdd.n2473 gnd 0.006542f
C5499 vdd.n2474 gnd 0.006542f
C5500 vdd.n2475 gnd 0.006542f
C5501 vdd.n2476 gnd 0.006542f
C5502 vdd.n2477 gnd 0.006542f
C5503 vdd.n2478 gnd 0.614504f
C5504 vdd.n2479 gnd 0.006542f
C5505 vdd.n2480 gnd 0.006542f
C5506 vdd.n2481 gnd 0.006542f
C5507 vdd.n2482 gnd 0.006542f
C5508 vdd.n2483 gnd 0.006542f
C5509 vdd.n2484 gnd 0.66858f
C5510 vdd.n2485 gnd 0.006542f
C5511 vdd.n2486 gnd 0.006542f
C5512 vdd.n2487 gnd 0.006542f
C5513 vdd.n2488 gnd 0.006542f
C5514 vdd.n2489 gnd 0.006542f
C5515 vdd.n2490 gnd 0.575176f
C5516 vdd.n2491 gnd 0.006542f
C5517 vdd.n2492 gnd 0.006542f
C5518 vdd.n2493 gnd 0.005195f
C5519 vdd.n2494 gnd 0.018952f
C5520 vdd.n2495 gnd 0.004618f
C5521 vdd.n2496 gnd 0.006542f
C5522 vdd.n2497 gnd 0.427695f
C5523 vdd.n2498 gnd 0.006542f
C5524 vdd.n2499 gnd 0.006542f
C5525 vdd.n2500 gnd 0.006542f
C5526 vdd.n2501 gnd 0.006542f
C5527 vdd.n2502 gnd 0.006542f
C5528 vdd.n2503 gnd 0.388367f
C5529 vdd.n2504 gnd 0.006542f
C5530 vdd.n2505 gnd 0.006542f
C5531 vdd.n2506 gnd 0.006542f
C5532 vdd.n2507 gnd 0.006542f
C5533 vdd.n2508 gnd 0.006542f
C5534 vdd.n2509 gnd 0.535848f
C5535 vdd.n2510 gnd 0.006542f
C5536 vdd.n2511 gnd 0.006542f
C5537 vdd.n2512 gnd 0.006542f
C5538 vdd.n2513 gnd 0.006542f
C5539 vdd.n2514 gnd 0.006542f
C5540 vdd.n2515 gnd 0.589924f
C5541 vdd.n2516 gnd 0.006542f
C5542 vdd.n2517 gnd 0.006542f
C5543 vdd.n2518 gnd 0.006542f
C5544 vdd.n2519 gnd 0.006542f
C5545 vdd.n2520 gnd 0.006542f
C5546 vdd.n2521 gnd 0.442443f
C5547 vdd.n2522 gnd 0.006542f
C5548 vdd.n2523 gnd 0.006542f
C5549 vdd.n2524 gnd 0.006542f
C5550 vdd.n2525 gnd 0.006542f
C5551 vdd.n2526 gnd 0.006542f
C5552 vdd.n2527 gnd 0.211389f
C5553 vdd.n2528 gnd 0.006542f
C5554 vdd.n2529 gnd 0.006542f
C5555 vdd.n2530 gnd 0.006542f
C5556 vdd.n2531 gnd 0.006542f
C5557 vdd.n2532 gnd 0.006542f
C5558 vdd.n2533 gnd 0.211389f
C5559 vdd.n2534 gnd 0.006542f
C5560 vdd.n2535 gnd 0.006542f
C5561 vdd.n2536 gnd 0.006542f
C5562 vdd.n2537 gnd 0.006542f
C5563 vdd.n2538 gnd 0.006542f
C5564 vdd.n2539 gnd 0.66858f
C5565 vdd.n2540 gnd 0.006542f
C5566 vdd.n2541 gnd 0.006542f
C5567 vdd.n2542 gnd 0.006542f
C5568 vdd.n2543 gnd 0.006542f
C5569 vdd.n2544 gnd 0.006542f
C5570 vdd.n2545 gnd 0.006542f
C5571 vdd.n2546 gnd 0.006542f
C5572 vdd.n2547 gnd 0.462107f
C5573 vdd.n2548 gnd 0.006542f
C5574 vdd.n2549 gnd 0.006542f
C5575 vdd.n2550 gnd 0.006542f
C5576 vdd.n2551 gnd 0.006542f
C5577 vdd.n2552 gnd 0.006542f
C5578 vdd.n2553 gnd 0.006542f
C5579 vdd.n2554 gnd 0.417863f
C5580 vdd.n2555 gnd 0.006542f
C5581 vdd.n2556 gnd 0.006542f
C5582 vdd.n2557 gnd 0.006542f
C5583 vdd.n2558 gnd 0.014855f
C5584 vdd.n2559 gnd 0.014008f
C5585 vdd.n2560 gnd 0.006542f
C5586 vdd.n2561 gnd 0.006542f
C5587 vdd.n2562 gnd 0.005051f
C5588 vdd.n2563 gnd 0.006542f
C5589 vdd.n2564 gnd 0.006542f
C5590 vdd.n2565 gnd 0.004762f
C5591 vdd.n2566 gnd 0.006542f
C5592 vdd.n2567 gnd 0.006542f
C5593 vdd.n2568 gnd 0.006542f
C5594 vdd.n2569 gnd 0.006542f
C5595 vdd.n2570 gnd 0.006542f
C5596 vdd.n2571 gnd 0.006542f
C5597 vdd.n2572 gnd 0.006542f
C5598 vdd.n2573 gnd 0.006542f
C5599 vdd.n2574 gnd 0.006542f
C5600 vdd.n2575 gnd 0.006542f
C5601 vdd.n2576 gnd 0.006542f
C5602 vdd.n2577 gnd 0.006542f
C5603 vdd.n2578 gnd 0.006542f
C5604 vdd.n2579 gnd 0.006542f
C5605 vdd.n2580 gnd 0.006542f
C5606 vdd.n2581 gnd 0.006542f
C5607 vdd.n2582 gnd 0.006542f
C5608 vdd.n2583 gnd 0.006542f
C5609 vdd.n2584 gnd 0.006542f
C5610 vdd.n2585 gnd 0.006542f
C5611 vdd.n2586 gnd 0.006542f
C5612 vdd.n2587 gnd 0.006542f
C5613 vdd.n2588 gnd 0.006542f
C5614 vdd.n2589 gnd 0.006542f
C5615 vdd.n2590 gnd 0.006542f
C5616 vdd.n2591 gnd 0.006542f
C5617 vdd.n2592 gnd 0.006542f
C5618 vdd.n2593 gnd 0.006542f
C5619 vdd.n2594 gnd 0.006542f
C5620 vdd.n2595 gnd 0.006542f
C5621 vdd.n2596 gnd 0.006542f
C5622 vdd.n2597 gnd 0.006542f
C5623 vdd.n2598 gnd 0.006542f
C5624 vdd.n2599 gnd 0.006542f
C5625 vdd.n2600 gnd 0.006542f
C5626 vdd.n2601 gnd 0.006542f
C5627 vdd.n2602 gnd 0.006542f
C5628 vdd.n2603 gnd 0.006542f
C5629 vdd.n2604 gnd 0.006542f
C5630 vdd.n2605 gnd 0.006542f
C5631 vdd.n2606 gnd 0.006542f
C5632 vdd.n2607 gnd 0.006542f
C5633 vdd.n2608 gnd 0.006542f
C5634 vdd.n2609 gnd 0.006542f
C5635 vdd.n2610 gnd 0.006542f
C5636 vdd.n2611 gnd 0.006542f
C5637 vdd.n2612 gnd 0.006542f
C5638 vdd.n2613 gnd 0.006542f
C5639 vdd.n2614 gnd 0.006542f
C5640 vdd.n2615 gnd 0.006542f
C5641 vdd.n2616 gnd 0.006542f
C5642 vdd.n2617 gnd 0.006542f
C5643 vdd.n2618 gnd 0.006542f
C5644 vdd.n2619 gnd 0.006542f
C5645 vdd.n2620 gnd 0.006542f
C5646 vdd.n2621 gnd 0.006542f
C5647 vdd.n2622 gnd 0.006542f
C5648 vdd.n2623 gnd 0.006542f
C5649 vdd.n2624 gnd 0.006542f
C5650 vdd.n2625 gnd 0.006542f
C5651 vdd.n2626 gnd 0.014855f
C5652 vdd.n2627 gnd 0.014008f
C5653 vdd.n2628 gnd 0.014008f
C5654 vdd.n2629 gnd 0.757069f
C5655 vdd.n2630 gnd 0.014008f
C5656 vdd.n2631 gnd 0.014855f
C5657 vdd.n2632 gnd 0.014008f
C5658 vdd.n2633 gnd 0.006542f
C5659 vdd.n2634 gnd 0.006542f
C5660 vdd.n2635 gnd 0.006542f
C5661 vdd.n2636 gnd 0.005051f
C5662 vdd.n2637 gnd 0.00935f
C5663 vdd.n2638 gnd 0.004762f
C5664 vdd.n2639 gnd 0.006542f
C5665 vdd.n2640 gnd 0.006542f
C5666 vdd.n2641 gnd 0.006542f
C5667 vdd.n2642 gnd 0.006542f
C5668 vdd.n2643 gnd 0.006542f
C5669 vdd.n2644 gnd 0.006542f
C5670 vdd.n2645 gnd 0.006542f
C5671 vdd.n2646 gnd 0.006542f
C5672 vdd.n2647 gnd 0.006542f
C5673 vdd.n2648 gnd 0.006542f
C5674 vdd.n2649 gnd 0.006542f
C5675 vdd.n2650 gnd 0.006542f
C5676 vdd.n2651 gnd 0.006542f
C5677 vdd.n2652 gnd 0.006542f
C5678 vdd.n2653 gnd 0.006542f
C5679 vdd.n2654 gnd 0.006542f
C5680 vdd.n2655 gnd 0.006542f
C5681 vdd.n2656 gnd 0.006542f
C5682 vdd.n2657 gnd 0.006542f
C5683 vdd.n2658 gnd 0.006542f
C5684 vdd.n2659 gnd 0.006542f
C5685 vdd.n2660 gnd 0.006542f
C5686 vdd.n2661 gnd 0.006542f
C5687 vdd.n2662 gnd 0.006542f
C5688 vdd.n2663 gnd 0.006542f
C5689 vdd.n2664 gnd 0.006542f
C5690 vdd.n2665 gnd 0.006542f
C5691 vdd.n2666 gnd 0.006542f
C5692 vdd.n2667 gnd 0.006542f
C5693 vdd.n2668 gnd 0.006542f
C5694 vdd.n2669 gnd 0.006542f
C5695 vdd.n2670 gnd 0.006542f
C5696 vdd.n2671 gnd 0.006542f
C5697 vdd.n2672 gnd 0.006542f
C5698 vdd.n2673 gnd 0.006542f
C5699 vdd.n2674 gnd 0.006542f
C5700 vdd.n2675 gnd 0.006542f
C5701 vdd.n2676 gnd 0.006542f
C5702 vdd.n2677 gnd 0.006542f
C5703 vdd.n2678 gnd 0.006542f
C5704 vdd.n2679 gnd 0.006542f
C5705 vdd.n2680 gnd 0.006542f
C5706 vdd.n2681 gnd 0.006542f
C5707 vdd.n2682 gnd 0.006542f
C5708 vdd.n2683 gnd 0.006542f
C5709 vdd.n2684 gnd 0.006542f
C5710 vdd.n2685 gnd 0.006542f
C5711 vdd.n2686 gnd 0.006542f
C5712 vdd.n2687 gnd 0.006542f
C5713 vdd.n2688 gnd 0.006542f
C5714 vdd.n2689 gnd 0.006542f
C5715 vdd.n2690 gnd 0.006542f
C5716 vdd.n2691 gnd 0.006542f
C5717 vdd.n2692 gnd 0.006542f
C5718 vdd.n2693 gnd 0.006542f
C5719 vdd.n2694 gnd 0.006542f
C5720 vdd.n2695 gnd 0.006542f
C5721 vdd.n2696 gnd 0.006542f
C5722 vdd.n2697 gnd 0.006542f
C5723 vdd.n2698 gnd 0.006542f
C5724 vdd.n2699 gnd 0.014855f
C5725 vdd.n2700 gnd 0.014855f
C5726 vdd.n2701 gnd 0.816061f
C5727 vdd.t222 gnd 2.90046f
C5728 vdd.t209 gnd 2.90046f
C5729 vdd.n2735 gnd 0.014855f
C5730 vdd.t227 gnd 0.57026f
C5731 vdd.n2736 gnd 0.006542f
C5732 vdd.t123 gnd 0.264369f
C5733 vdd.t124 gnd 0.270614f
C5734 vdd.t121 gnd 0.17259f
C5735 vdd.n2737 gnd 0.093276f
C5736 vdd.n2738 gnd 0.052909f
C5737 vdd.n2739 gnd 0.006542f
C5738 vdd.t133 gnd 0.264369f
C5739 vdd.t134 gnd 0.270614f
C5740 vdd.t132 gnd 0.17259f
C5741 vdd.n2740 gnd 0.093276f
C5742 vdd.n2741 gnd 0.052909f
C5743 vdd.n2742 gnd 0.00935f
C5744 vdd.n2743 gnd 0.014855f
C5745 vdd.n2744 gnd 0.014855f
C5746 vdd.n2745 gnd 0.006542f
C5747 vdd.n2746 gnd 0.006542f
C5748 vdd.n2747 gnd 0.006542f
C5749 vdd.n2748 gnd 0.006542f
C5750 vdd.n2749 gnd 0.006542f
C5751 vdd.n2750 gnd 0.006542f
C5752 vdd.n2751 gnd 0.006542f
C5753 vdd.n2752 gnd 0.006542f
C5754 vdd.n2753 gnd 0.006542f
C5755 vdd.n2754 gnd 0.006542f
C5756 vdd.n2755 gnd 0.006542f
C5757 vdd.n2756 gnd 0.006542f
C5758 vdd.n2757 gnd 0.006542f
C5759 vdd.n2758 gnd 0.006542f
C5760 vdd.n2759 gnd 0.006542f
C5761 vdd.n2760 gnd 0.006542f
C5762 vdd.n2761 gnd 0.006542f
C5763 vdd.n2762 gnd 0.006542f
C5764 vdd.n2763 gnd 0.006542f
C5765 vdd.n2764 gnd 0.006542f
C5766 vdd.n2765 gnd 0.006542f
C5767 vdd.n2766 gnd 0.006542f
C5768 vdd.n2767 gnd 0.006542f
C5769 vdd.n2768 gnd 0.006542f
C5770 vdd.n2769 gnd 0.006542f
C5771 vdd.n2770 gnd 0.006542f
C5772 vdd.n2771 gnd 0.006542f
C5773 vdd.n2772 gnd 0.006542f
C5774 vdd.n2773 gnd 0.006542f
C5775 vdd.n2774 gnd 0.006542f
C5776 vdd.n2775 gnd 0.006542f
C5777 vdd.n2776 gnd 0.006542f
C5778 vdd.n2777 gnd 0.006542f
C5779 vdd.n2778 gnd 0.006542f
C5780 vdd.n2779 gnd 0.006542f
C5781 vdd.n2780 gnd 0.006542f
C5782 vdd.n2781 gnd 0.006542f
C5783 vdd.n2782 gnd 0.006542f
C5784 vdd.n2783 gnd 0.006542f
C5785 vdd.n2784 gnd 0.006542f
C5786 vdd.n2785 gnd 0.006542f
C5787 vdd.n2786 gnd 0.006542f
C5788 vdd.n2787 gnd 0.006542f
C5789 vdd.n2788 gnd 0.006542f
C5790 vdd.n2789 gnd 0.006542f
C5791 vdd.n2790 gnd 0.006542f
C5792 vdd.n2791 gnd 0.006542f
C5793 vdd.n2792 gnd 0.006542f
C5794 vdd.n2793 gnd 0.006542f
C5795 vdd.n2794 gnd 0.006542f
C5796 vdd.n2795 gnd 0.006542f
C5797 vdd.n2796 gnd 0.006542f
C5798 vdd.n2797 gnd 0.006542f
C5799 vdd.n2798 gnd 0.006542f
C5800 vdd.n2799 gnd 0.006542f
C5801 vdd.n2800 gnd 0.006542f
C5802 vdd.n2801 gnd 0.006542f
C5803 vdd.n2802 gnd 0.006542f
C5804 vdd.n2803 gnd 0.006542f
C5805 vdd.n2804 gnd 0.006542f
C5806 vdd.n2805 gnd 0.004762f
C5807 vdd.n2806 gnd 0.006542f
C5808 vdd.n2807 gnd 0.006542f
C5809 vdd.n2808 gnd 0.005051f
C5810 vdd.n2809 gnd 0.006542f
C5811 vdd.n2810 gnd 0.006542f
C5812 vdd.n2811 gnd 0.014855f
C5813 vdd.n2812 gnd 0.014008f
C5814 vdd.n2813 gnd 0.014008f
C5815 vdd.n2814 gnd 0.006542f
C5816 vdd.n2815 gnd 0.006542f
C5817 vdd.n2816 gnd 0.006542f
C5818 vdd.n2817 gnd 0.006542f
C5819 vdd.n2818 gnd 0.006542f
C5820 vdd.n2819 gnd 0.006542f
C5821 vdd.n2820 gnd 0.006542f
C5822 vdd.n2821 gnd 0.006542f
C5823 vdd.n2822 gnd 0.006542f
C5824 vdd.n2823 gnd 0.006542f
C5825 vdd.n2824 gnd 0.006542f
C5826 vdd.n2825 gnd 0.006542f
C5827 vdd.n2826 gnd 0.006542f
C5828 vdd.n2827 gnd 0.006542f
C5829 vdd.n2828 gnd 0.006542f
C5830 vdd.n2829 gnd 0.006542f
C5831 vdd.n2830 gnd 0.006542f
C5832 vdd.n2831 gnd 0.006542f
C5833 vdd.n2832 gnd 0.006542f
C5834 vdd.n2833 gnd 0.006542f
C5835 vdd.n2834 gnd 0.006542f
C5836 vdd.n2835 gnd 0.006542f
C5837 vdd.n2836 gnd 0.006542f
C5838 vdd.n2837 gnd 0.006542f
C5839 vdd.n2838 gnd 0.006542f
C5840 vdd.n2839 gnd 0.006542f
C5841 vdd.n2840 gnd 0.006542f
C5842 vdd.n2841 gnd 0.006542f
C5843 vdd.n2842 gnd 0.006542f
C5844 vdd.n2843 gnd 0.006542f
C5845 vdd.n2844 gnd 0.006542f
C5846 vdd.n2845 gnd 0.006542f
C5847 vdd.n2846 gnd 0.006542f
C5848 vdd.n2847 gnd 0.006542f
C5849 vdd.n2848 gnd 0.006542f
C5850 vdd.n2849 gnd 0.006542f
C5851 vdd.n2850 gnd 0.006542f
C5852 vdd.n2851 gnd 0.006542f
C5853 vdd.n2852 gnd 0.006542f
C5854 vdd.n2853 gnd 0.006542f
C5855 vdd.n2854 gnd 0.006542f
C5856 vdd.n2855 gnd 0.006542f
C5857 vdd.n2856 gnd 0.006542f
C5858 vdd.n2857 gnd 0.006542f
C5859 vdd.n2858 gnd 0.006542f
C5860 vdd.n2859 gnd 0.006542f
C5861 vdd.n2860 gnd 0.006542f
C5862 vdd.n2861 gnd 0.006542f
C5863 vdd.n2862 gnd 0.006542f
C5864 vdd.n2863 gnd 0.006542f
C5865 vdd.n2864 gnd 0.006542f
C5866 vdd.n2865 gnd 0.006542f
C5867 vdd.n2866 gnd 0.006542f
C5868 vdd.n2867 gnd 0.006542f
C5869 vdd.n2868 gnd 0.006542f
C5870 vdd.n2869 gnd 0.006542f
C5871 vdd.n2870 gnd 0.006542f
C5872 vdd.n2871 gnd 0.006542f
C5873 vdd.n2872 gnd 0.006542f
C5874 vdd.n2873 gnd 0.006542f
C5875 vdd.n2874 gnd 0.006542f
C5876 vdd.n2875 gnd 0.006542f
C5877 vdd.n2876 gnd 0.006542f
C5878 vdd.n2877 gnd 0.006542f
C5879 vdd.n2878 gnd 0.006542f
C5880 vdd.n2879 gnd 0.006542f
C5881 vdd.n2880 gnd 0.006542f
C5882 vdd.n2881 gnd 0.006542f
C5883 vdd.n2882 gnd 0.006542f
C5884 vdd.n2883 gnd 0.006542f
C5885 vdd.n2884 gnd 0.006542f
C5886 vdd.n2885 gnd 0.006542f
C5887 vdd.n2886 gnd 0.006542f
C5888 vdd.n2887 gnd 0.006542f
C5889 vdd.n2888 gnd 0.006542f
C5890 vdd.n2889 gnd 0.006542f
C5891 vdd.n2890 gnd 0.006542f
C5892 vdd.n2891 gnd 0.006542f
C5893 vdd.n2892 gnd 0.006542f
C5894 vdd.n2893 gnd 0.006542f
C5895 vdd.n2894 gnd 0.006542f
C5896 vdd.n2895 gnd 0.006542f
C5897 vdd.n2896 gnd 0.006542f
C5898 vdd.n2897 gnd 0.006542f
C5899 vdd.n2898 gnd 0.006542f
C5900 vdd.n2899 gnd 0.006542f
C5901 vdd.n2900 gnd 0.006542f
C5902 vdd.n2901 gnd 0.006542f
C5903 vdd.n2902 gnd 0.006542f
C5904 vdd.n2903 gnd 0.006542f
C5905 vdd.n2904 gnd 0.006542f
C5906 vdd.n2905 gnd 0.006542f
C5907 vdd.n2906 gnd 0.006542f
C5908 vdd.n2907 gnd 0.006542f
C5909 vdd.n2908 gnd 0.006542f
C5910 vdd.n2909 gnd 0.006542f
C5911 vdd.n2910 gnd 0.006542f
C5912 vdd.n2911 gnd 0.006542f
C5913 vdd.n2912 gnd 0.006542f
C5914 vdd.n2913 gnd 0.006542f
C5915 vdd.n2914 gnd 0.006542f
C5916 vdd.n2915 gnd 0.211389f
C5917 vdd.n2916 gnd 0.006542f
C5918 vdd.n2917 gnd 0.006542f
C5919 vdd.n2918 gnd 0.006542f
C5920 vdd.n2919 gnd 0.006542f
C5921 vdd.n2920 gnd 0.006542f
C5922 vdd.n2921 gnd 0.211389f
C5923 vdd.n2922 gnd 0.006542f
C5924 vdd.n2923 gnd 0.006542f
C5925 vdd.n2924 gnd 0.006542f
C5926 vdd.n2925 gnd 0.006542f
C5927 vdd.n2926 gnd 0.006542f
C5928 vdd.n2927 gnd 0.006542f
C5929 vdd.n2928 gnd 0.006542f
C5930 vdd.n2929 gnd 0.006542f
C5931 vdd.n2930 gnd 0.006542f
C5932 vdd.n2931 gnd 0.006542f
C5933 vdd.n2932 gnd 0.006542f
C5934 vdd.n2933 gnd 0.417863f
C5935 vdd.n2934 gnd 0.006542f
C5936 vdd.n2935 gnd 0.006542f
C5937 vdd.n2936 gnd 0.006542f
C5938 vdd.n2937 gnd 0.014008f
C5939 vdd.n2938 gnd 0.014008f
C5940 vdd.n2939 gnd 0.014855f
C5941 vdd.n2940 gnd 0.014855f
C5942 vdd.n2941 gnd 0.006542f
C5943 vdd.n2942 gnd 0.006542f
C5944 vdd.n2943 gnd 0.006542f
C5945 vdd.n2944 gnd 0.005051f
C5946 vdd.n2945 gnd 0.00935f
C5947 vdd.n2946 gnd 0.004762f
C5948 vdd.n2947 gnd 0.006542f
C5949 vdd.n2948 gnd 0.006542f
C5950 vdd.n2949 gnd 0.006542f
C5951 vdd.n2950 gnd 0.006542f
C5952 vdd.n2951 gnd 0.006542f
C5953 vdd.n2952 gnd 0.006542f
C5954 vdd.n2953 gnd 0.006542f
C5955 vdd.n2954 gnd 0.006542f
C5956 vdd.n2955 gnd 0.006542f
C5957 vdd.n2956 gnd 0.006542f
C5958 vdd.n2957 gnd 0.006542f
C5959 vdd.n2958 gnd 0.006542f
C5960 vdd.n2959 gnd 0.006542f
C5961 vdd.n2960 gnd 0.006542f
C5962 vdd.n2961 gnd 0.006542f
C5963 vdd.n2962 gnd 0.006542f
C5964 vdd.n2963 gnd 0.006542f
C5965 vdd.n2964 gnd 0.006542f
C5966 vdd.n2965 gnd 0.006542f
C5967 vdd.n2966 gnd 0.006542f
C5968 vdd.n2967 gnd 0.006542f
C5969 vdd.n2968 gnd 0.006542f
C5970 vdd.n2969 gnd 0.006542f
C5971 vdd.n2970 gnd 0.006542f
C5972 vdd.n2971 gnd 0.006542f
C5973 vdd.n2972 gnd 0.006542f
C5974 vdd.n2973 gnd 0.006542f
C5975 vdd.n2974 gnd 0.006542f
C5976 vdd.n2975 gnd 0.006542f
C5977 vdd.n2976 gnd 0.006542f
C5978 vdd.n2977 gnd 0.006542f
C5979 vdd.n2978 gnd 0.006542f
C5980 vdd.n2979 gnd 0.006542f
C5981 vdd.n2980 gnd 0.006542f
C5982 vdd.n2981 gnd 0.006542f
C5983 vdd.n2982 gnd 0.006542f
C5984 vdd.n2983 gnd 0.006542f
C5985 vdd.n2984 gnd 0.006542f
C5986 vdd.n2985 gnd 0.006542f
C5987 vdd.n2986 gnd 0.006542f
C5988 vdd.n2987 gnd 0.006542f
C5989 vdd.n2988 gnd 0.006542f
C5990 vdd.n2989 gnd 0.006542f
C5991 vdd.n2990 gnd 0.006542f
C5992 vdd.n2991 gnd 0.006542f
C5993 vdd.n2992 gnd 0.006542f
C5994 vdd.n2993 gnd 0.006542f
C5995 vdd.n2994 gnd 0.006542f
C5996 vdd.n2995 gnd 0.006542f
C5997 vdd.n2996 gnd 0.006542f
C5998 vdd.n2997 gnd 0.006542f
C5999 vdd.n2998 gnd 0.006542f
C6000 vdd.n2999 gnd 0.006542f
C6001 vdd.n3000 gnd 0.006542f
C6002 vdd.n3001 gnd 0.006542f
C6003 vdd.n3002 gnd 0.006542f
C6004 vdd.n3003 gnd 0.006542f
C6005 vdd.n3004 gnd 0.006542f
C6006 vdd.n3005 gnd 0.816061f
C6007 vdd.n3007 gnd 0.014855f
C6008 vdd.n3008 gnd 0.014855f
C6009 vdd.n3009 gnd 0.014008f
C6010 vdd.n3010 gnd 0.006542f
C6011 vdd.n3011 gnd 0.006542f
C6012 vdd.n3012 gnd 0.393283f
C6013 vdd.n3013 gnd 0.006542f
C6014 vdd.n3014 gnd 0.006542f
C6015 vdd.n3015 gnd 0.006542f
C6016 vdd.n3016 gnd 0.006542f
C6017 vdd.n3017 gnd 0.006542f
C6018 vdd.n3018 gnd 0.398199f
C6019 vdd.n3019 gnd 0.006542f
C6020 vdd.n3020 gnd 0.006542f
C6021 vdd.n3021 gnd 0.006542f
C6022 vdd.n3022 gnd 0.006542f
C6023 vdd.n3023 gnd 0.006542f
C6024 vdd.n3024 gnd 0.66858f
C6025 vdd.n3025 gnd 0.006542f
C6026 vdd.n3026 gnd 0.006542f
C6027 vdd.n3027 gnd 0.006542f
C6028 vdd.n3028 gnd 0.006542f
C6029 vdd.n3029 gnd 0.006542f
C6030 vdd.n3030 gnd 0.481771f
C6031 vdd.n3031 gnd 0.006542f
C6032 vdd.n3032 gnd 0.006542f
C6033 vdd.n3033 gnd 0.006542f
C6034 vdd.n3034 gnd 0.006542f
C6035 vdd.n3035 gnd 0.006542f
C6036 vdd.n3036 gnd 0.604672f
C6037 vdd.n3037 gnd 0.006542f
C6038 vdd.n3038 gnd 0.006542f
C6039 vdd.n3039 gnd 0.006542f
C6040 vdd.n3040 gnd 0.006542f
C6041 vdd.n3041 gnd 0.006542f
C6042 vdd.n3042 gnd 0.496519f
C6043 vdd.n3043 gnd 0.006542f
C6044 vdd.n3044 gnd 0.006542f
C6045 vdd.n3045 gnd 0.006542f
C6046 vdd.n3046 gnd 0.006542f
C6047 vdd.n3047 gnd 0.006542f
C6048 vdd.n3048 gnd 0.349038f
C6049 vdd.n3049 gnd 0.006542f
C6050 vdd.n3050 gnd 0.006542f
C6051 vdd.n3051 gnd 0.006542f
C6052 vdd.n3052 gnd 0.006542f
C6053 vdd.n3053 gnd 0.006542f
C6054 vdd.n3054 gnd 0.211389f
C6055 vdd.n3055 gnd 0.006542f
C6056 vdd.n3056 gnd 0.006542f
C6057 vdd.n3057 gnd 0.006542f
C6058 vdd.n3058 gnd 0.006542f
C6059 vdd.n3059 gnd 0.006542f
C6060 vdd.n3060 gnd 0.614504f
C6061 vdd.n3061 gnd 0.006542f
C6062 vdd.n3062 gnd 0.006542f
C6063 vdd.n3063 gnd 0.006542f
C6064 vdd.n3064 gnd 0.004618f
C6065 vdd.n3065 gnd 0.006542f
C6066 vdd.n3066 gnd 0.006542f
C6067 vdd.n3067 gnd 0.66858f
C6068 vdd.n3068 gnd 0.006542f
C6069 vdd.n3069 gnd 0.006542f
C6070 vdd.n3070 gnd 0.006542f
C6071 vdd.n3071 gnd 0.006542f
C6072 vdd.n3072 gnd 0.006542f
C6073 vdd.n3073 gnd 0.530931f
C6074 vdd.n3074 gnd 0.006542f
C6075 vdd.n3075 gnd 0.005195f
C6076 vdd.n3076 gnd 0.006542f
C6077 vdd.n3077 gnd 0.006542f
C6078 vdd.n3078 gnd 0.006542f
C6079 vdd.n3079 gnd 0.427695f
C6080 vdd.n3080 gnd 0.006542f
C6081 vdd.n3081 gnd 0.006542f
C6082 vdd.n3082 gnd 0.006542f
C6083 vdd.n3083 gnd 0.006542f
C6084 vdd.n3084 gnd 0.006542f
C6085 vdd.n3085 gnd 0.388367f
C6086 vdd.n3086 gnd 0.006542f
C6087 vdd.n3087 gnd 0.006542f
C6088 vdd.n3088 gnd 0.006542f
C6089 vdd.n3089 gnd 0.006542f
C6090 vdd.n3090 gnd 0.006542f
C6091 vdd.n3091 gnd 0.535848f
C6092 vdd.n3092 gnd 0.006542f
C6093 vdd.n3093 gnd 0.006542f
C6094 vdd.n3094 gnd 0.006542f
C6095 vdd.n3095 gnd 0.006542f
C6096 vdd.n3096 gnd 0.006542f
C6097 vdd.n3097 gnd 0.66858f
C6098 vdd.n3098 gnd 0.006542f
C6099 vdd.n3099 gnd 0.006542f
C6100 vdd.n3100 gnd 0.006542f
C6101 vdd.n3101 gnd 0.006542f
C6102 vdd.n3102 gnd 0.006542f
C6103 vdd.n3103 gnd 0.653832f
C6104 vdd.n3104 gnd 0.006542f
C6105 vdd.n3105 gnd 0.006542f
C6106 vdd.n3106 gnd 0.006542f
C6107 vdd.n3107 gnd 0.006542f
C6108 vdd.n3108 gnd 0.006542f
C6109 vdd.n3109 gnd 0.506351f
C6110 vdd.n3110 gnd 0.006542f
C6111 vdd.n3111 gnd 0.006542f
C6112 vdd.n3112 gnd 0.006542f
C6113 vdd.n3113 gnd 0.006542f
C6114 vdd.n3114 gnd 0.006542f
C6115 vdd.n3115 gnd 0.35887f
C6116 vdd.n3116 gnd 0.006542f
C6117 vdd.n3117 gnd 0.006542f
C6118 vdd.n3118 gnd 0.006542f
C6119 vdd.n3119 gnd 0.006542f
C6120 vdd.n3120 gnd 0.006542f
C6121 vdd.n3121 gnd 0.66858f
C6122 vdd.n3122 gnd 0.006542f
C6123 vdd.n3123 gnd 0.006542f
C6124 vdd.n3124 gnd 0.006542f
C6125 vdd.n3125 gnd 0.006542f
C6126 vdd.n3126 gnd 0.006542f
C6127 vdd.n3127 gnd 0.006542f
C6128 vdd.n3129 gnd 0.006542f
C6129 vdd.n3130 gnd 0.006542f
C6130 vdd.n3132 gnd 0.006542f
C6131 vdd.n3133 gnd 0.006542f
C6132 vdd.n3136 gnd 0.006542f
C6133 vdd.n3137 gnd 0.006542f
C6134 vdd.n3138 gnd 0.006542f
C6135 vdd.n3139 gnd 0.006542f
C6136 vdd.n3141 gnd 0.006542f
C6137 vdd.n3142 gnd 0.006542f
C6138 vdd.n3143 gnd 0.006542f
C6139 vdd.n3144 gnd 0.006542f
C6140 vdd.n3145 gnd 0.006542f
C6141 vdd.n3146 gnd 0.006542f
C6142 vdd.n3148 gnd 0.006542f
C6143 vdd.n3149 gnd 0.006542f
C6144 vdd.n3150 gnd 0.006542f
C6145 vdd.n3151 gnd 0.006542f
C6146 vdd.n3152 gnd 0.006542f
C6147 vdd.n3153 gnd 0.006542f
C6148 vdd.n3155 gnd 0.006542f
C6149 vdd.n3156 gnd 0.006542f
C6150 vdd.n3157 gnd 0.006542f
C6151 vdd.n3158 gnd 0.006542f
C6152 vdd.n3159 gnd 0.006542f
C6153 vdd.n3160 gnd 0.006542f
C6154 vdd.n3162 gnd 0.006542f
C6155 vdd.n3163 gnd 0.014855f
C6156 vdd.n3164 gnd 0.014855f
C6157 vdd.n3165 gnd 0.014008f
C6158 vdd.n3166 gnd 0.006542f
C6159 vdd.n3167 gnd 0.006542f
C6160 vdd.n3168 gnd 0.006542f
C6161 vdd.n3169 gnd 0.006542f
C6162 vdd.n3170 gnd 0.006542f
C6163 vdd.n3171 gnd 0.006542f
C6164 vdd.n3172 gnd 0.66858f
C6165 vdd.n3173 gnd 0.006542f
C6166 vdd.n3174 gnd 0.006542f
C6167 vdd.n3175 gnd 0.006542f
C6168 vdd.n3176 gnd 0.006542f
C6169 vdd.n3177 gnd 0.006542f
C6170 vdd.n3178 gnd 0.476855f
C6171 vdd.n3179 gnd 0.006542f
C6172 vdd.n3180 gnd 0.006542f
C6173 vdd.n3181 gnd 0.006542f
C6174 vdd.n3182 gnd 0.014855f
C6175 vdd.n3184 gnd 0.014855f
C6176 vdd.n3185 gnd 0.014008f
C6177 vdd.n3186 gnd 0.006542f
C6178 vdd.n3187 gnd 0.005051f
C6179 vdd.n3188 gnd 0.006542f
C6180 vdd.n3190 gnd 0.006542f
C6181 vdd.n3191 gnd 0.006542f
C6182 vdd.n3192 gnd 0.006542f
C6183 vdd.n3193 gnd 0.006542f
C6184 vdd.n3194 gnd 0.006542f
C6185 vdd.n3195 gnd 0.006542f
C6186 vdd.n3197 gnd 0.006542f
C6187 vdd.n3198 gnd 0.006542f
C6188 vdd.n3199 gnd 0.006542f
C6189 vdd.n3200 gnd 0.006542f
C6190 vdd.n3201 gnd 0.006542f
C6191 vdd.n3202 gnd 0.006542f
C6192 vdd.n3204 gnd 0.006542f
C6193 vdd.n3205 gnd 0.006542f
C6194 vdd.n3206 gnd 0.006542f
C6195 vdd.n3207 gnd 0.006542f
C6196 vdd.n3208 gnd 0.006542f
C6197 vdd.n3209 gnd 0.006542f
C6198 vdd.n3211 gnd 0.006542f
C6199 vdd.n3212 gnd 0.006542f
C6200 vdd.n3213 gnd 0.006542f
C6201 vdd.n3214 gnd 1.02503f
C6202 vdd.n3215 gnd 0.040397f
C6203 vdd.n3216 gnd 0.006542f
C6204 vdd.n3217 gnd 0.006542f
C6205 vdd.n3219 gnd 0.006542f
C6206 vdd.n3220 gnd 0.006542f
C6207 vdd.n3221 gnd 0.006542f
C6208 vdd.n3222 gnd 0.006542f
C6209 vdd.n3223 gnd 0.006542f
C6210 vdd.n3224 gnd 0.006542f
C6211 vdd.n3226 gnd 0.006542f
C6212 vdd.n3227 gnd 0.006542f
C6213 vdd.n3228 gnd 0.006542f
C6214 vdd.n3229 gnd 0.006542f
C6215 vdd.n3230 gnd 0.006542f
C6216 vdd.n3231 gnd 0.006542f
C6217 vdd.n3233 gnd 0.006542f
C6218 vdd.n3234 gnd 0.006542f
C6219 vdd.n3235 gnd 0.006542f
C6220 vdd.n3236 gnd 0.006542f
C6221 vdd.n3237 gnd 0.006542f
C6222 vdd.n3238 gnd 0.006542f
C6223 vdd.n3240 gnd 0.006542f
C6224 vdd.n3241 gnd 0.006542f
C6225 vdd.n3243 gnd 0.006542f
C6226 vdd.n3244 gnd 0.006542f
C6227 vdd.n3245 gnd 0.014855f
C6228 vdd.n3246 gnd 0.014008f
C6229 vdd.n3247 gnd 0.014008f
C6230 vdd.n3248 gnd 0.90455f
C6231 vdd.n3249 gnd 0.014008f
C6232 vdd.n3250 gnd 0.014855f
C6233 vdd.n3251 gnd 0.014008f
C6234 vdd.n3252 gnd 0.006542f
C6235 vdd.n3253 gnd 0.005051f
C6236 vdd.n3254 gnd 0.006542f
C6237 vdd.n3256 gnd 0.006542f
C6238 vdd.n3257 gnd 0.006542f
C6239 vdd.n3258 gnd 0.006542f
C6240 vdd.n3259 gnd 0.006542f
C6241 vdd.n3260 gnd 0.006542f
C6242 vdd.n3261 gnd 0.006542f
C6243 vdd.n3263 gnd 0.006542f
C6244 vdd.n3264 gnd 0.006542f
C6245 vdd.n3265 gnd 0.006542f
C6246 vdd.n3266 gnd 0.006542f
C6247 vdd.n3267 gnd 0.006542f
C6248 vdd.n3268 gnd 0.006542f
C6249 vdd.n3270 gnd 0.006542f
C6250 vdd.n3271 gnd 0.006542f
C6251 vdd.n3272 gnd 0.006542f
C6252 vdd.n3273 gnd 0.006542f
C6253 vdd.n3274 gnd 0.006542f
C6254 vdd.n3275 gnd 0.006542f
C6255 vdd.n3277 gnd 0.006542f
C6256 vdd.n3278 gnd 0.006542f
C6257 vdd.n3280 gnd 0.006542f
C6258 vdd.n3281 gnd 0.040397f
C6259 vdd.n3282 gnd 1.02503f
C6260 vdd.n3283 gnd 0.008274f
C6261 vdd.n3284 gnd 0.003678f
C6262 vdd.t89 gnd 0.118362f
C6263 vdd.t90 gnd 0.126496f
C6264 vdd.t87 gnd 0.154579f
C6265 vdd.n3285 gnd 0.198149f
C6266 vdd.n3286 gnd 0.166481f
C6267 vdd.n3287 gnd 0.011925f
C6268 vdd.n3288 gnd 0.009621f
C6269 vdd.n3289 gnd 0.004065f
C6270 vdd.n3290 gnd 0.007744f
C6271 vdd.n3291 gnd 0.009621f
C6272 vdd.n3292 gnd 0.009621f
C6273 vdd.n3293 gnd 0.007744f
C6274 vdd.n3294 gnd 0.007744f
C6275 vdd.n3295 gnd 0.009621f
C6276 vdd.n3297 gnd 0.009621f
C6277 vdd.n3298 gnd 0.007744f
C6278 vdd.n3299 gnd 0.007744f
C6279 vdd.n3300 gnd 0.007744f
C6280 vdd.n3301 gnd 0.009621f
C6281 vdd.n3303 gnd 0.009621f
C6282 vdd.n3305 gnd 0.009621f
C6283 vdd.n3306 gnd 0.007744f
C6284 vdd.n3307 gnd 0.007744f
C6285 vdd.n3308 gnd 0.007744f
C6286 vdd.n3309 gnd 0.009621f
C6287 vdd.n3311 gnd 0.009621f
C6288 vdd.n3313 gnd 0.009621f
C6289 vdd.n3314 gnd 0.007744f
C6290 vdd.n3315 gnd 0.007744f
C6291 vdd.n3316 gnd 0.007744f
C6292 vdd.n3317 gnd 0.009621f
C6293 vdd.n3319 gnd 0.009621f
C6294 vdd.n3320 gnd 0.009621f
C6295 vdd.n3321 gnd 0.007744f
C6296 vdd.n3322 gnd 0.007744f
C6297 vdd.n3323 gnd 0.009621f
C6298 vdd.n3324 gnd 0.009621f
C6299 vdd.n3326 gnd 0.009621f
C6300 vdd.n3327 gnd 0.007744f
C6301 vdd.n3328 gnd 0.009621f
C6302 vdd.n3329 gnd 0.009621f
C6303 vdd.n3330 gnd 0.009621f
C6304 vdd.n3331 gnd 0.015797f
C6305 vdd.n3332 gnd 0.005266f
C6306 vdd.n3333 gnd 0.009621f
C6307 vdd.n3335 gnd 0.009621f
C6308 vdd.n3337 gnd 0.009621f
C6309 vdd.n3338 gnd 0.007744f
C6310 vdd.n3339 gnd 0.007744f
C6311 vdd.n3340 gnd 0.007744f
C6312 vdd.n3341 gnd 0.009621f
C6313 vdd.n3343 gnd 0.009621f
C6314 vdd.n3345 gnd 0.009621f
C6315 vdd.n3346 gnd 0.007744f
C6316 vdd.n3347 gnd 0.007744f
C6317 vdd.n3348 gnd 0.007744f
C6318 vdd.n3349 gnd 0.009621f
C6319 vdd.n3351 gnd 0.009621f
C6320 vdd.n3353 gnd 0.009621f
C6321 vdd.n3354 gnd 0.007744f
C6322 vdd.n3355 gnd 0.007744f
C6323 vdd.n3356 gnd 0.007744f
C6324 vdd.n3357 gnd 0.009621f
C6325 vdd.n3359 gnd 0.009621f
C6326 vdd.n3361 gnd 0.009621f
C6327 vdd.n3362 gnd 0.007744f
C6328 vdd.n3363 gnd 0.007744f
C6329 vdd.n3364 gnd 0.007744f
C6330 vdd.n3365 gnd 0.009621f
C6331 vdd.n3367 gnd 0.009621f
C6332 vdd.n3369 gnd 0.009621f
C6333 vdd.n3370 gnd 0.007744f
C6334 vdd.n3371 gnd 0.007744f
C6335 vdd.n3372 gnd 0.006466f
C6336 vdd.n3373 gnd 0.009621f
C6337 vdd.n3375 gnd 0.009621f
C6338 vdd.n3377 gnd 0.009621f
C6339 vdd.n3378 gnd 0.006466f
C6340 vdd.n3379 gnd 0.007744f
C6341 vdd.n3380 gnd 0.007744f
C6342 vdd.n3381 gnd 0.009621f
C6343 vdd.n3383 gnd 0.009621f
C6344 vdd.n3385 gnd 0.009621f
C6345 vdd.n3386 gnd 0.007744f
C6346 vdd.n3387 gnd 0.007744f
C6347 vdd.n3388 gnd 0.007744f
C6348 vdd.n3389 gnd 0.009621f
C6349 vdd.n3391 gnd 0.009621f
C6350 vdd.n3393 gnd 0.009621f
C6351 vdd.n3394 gnd 0.007744f
C6352 vdd.n3395 gnd 0.007744f
C6353 vdd.n3396 gnd 0.007744f
C6354 vdd.n3397 gnd 0.009621f
C6355 vdd.n3399 gnd 0.009621f
C6356 vdd.n3400 gnd 0.009621f
C6357 vdd.n3401 gnd 0.007744f
C6358 vdd.n3402 gnd 0.007744f
C6359 vdd.n3403 gnd 0.009621f
C6360 vdd.n3404 gnd 0.009621f
C6361 vdd.n3405 gnd 0.007744f
C6362 vdd.n3406 gnd 0.007744f
C6363 vdd.n3407 gnd 0.009621f
C6364 vdd.n3408 gnd 0.009621f
C6365 vdd.n3410 gnd 0.009621f
C6366 vdd.n3411 gnd 0.007744f
C6367 vdd.n3412 gnd 0.006427f
C6368 vdd.n3413 gnd 0.022059f
C6369 vdd.n3414 gnd 0.021909f
C6370 vdd.n3415 gnd 0.006427f
C6371 vdd.n3416 gnd 0.021909f
C6372 vdd.n3417 gnd 1.29783f
C6373 vdd.n3418 gnd 0.021909f
C6374 vdd.n3419 gnd 0.006427f
C6375 vdd.n3420 gnd 0.021909f
C6376 vdd.n3421 gnd 0.009621f
C6377 vdd.n3422 gnd 0.009621f
C6378 vdd.n3423 gnd 0.007744f
C6379 vdd.n3424 gnd 0.009621f
C6380 vdd.n3425 gnd 0.92913f
C6381 vdd.n3426 gnd 0.009621f
C6382 vdd.n3427 gnd 0.007744f
C6383 vdd.n3428 gnd 0.009621f
C6384 vdd.n3429 gnd 0.009621f
C6385 vdd.n3430 gnd 0.009621f
C6386 vdd.n3431 gnd 0.007744f
C6387 vdd.n3432 gnd 0.009621f
C6388 vdd.n3433 gnd 0.958626f
C6389 vdd.n3434 gnd 0.009621f
C6390 vdd.n3435 gnd 0.007744f
C6391 vdd.n3436 gnd 0.009621f
C6392 vdd.n3437 gnd 0.009621f
C6393 vdd.n3438 gnd 0.009621f
C6394 vdd.n3439 gnd 0.007744f
C6395 vdd.n3440 gnd 0.009621f
C6396 vdd.t63 gnd 0.491603f
C6397 vdd.n3441 gnd 0.791481f
C6398 vdd.n3442 gnd 0.009621f
C6399 vdd.n3443 gnd 0.007744f
C6400 vdd.n3444 gnd 0.009621f
C6401 vdd.n3445 gnd 0.009621f
C6402 vdd.n3446 gnd 0.009621f
C6403 vdd.n3447 gnd 0.007744f
C6404 vdd.n3448 gnd 0.009621f
C6405 vdd.n3449 gnd 0.624336f
C6406 vdd.n3450 gnd 0.009621f
C6407 vdd.n3451 gnd 0.007744f
C6408 vdd.n3452 gnd 0.009621f
C6409 vdd.n3453 gnd 0.009621f
C6410 vdd.n3454 gnd 0.009621f
C6411 vdd.n3455 gnd 0.007744f
C6412 vdd.n3456 gnd 0.009621f
C6413 vdd.n3457 gnd 0.781649f
C6414 vdd.n3458 gnd 0.526015f
C6415 vdd.n3459 gnd 0.009621f
C6416 vdd.n3460 gnd 0.007744f
C6417 vdd.n3461 gnd 0.009621f
C6418 vdd.n3462 gnd 0.009621f
C6419 vdd.n3463 gnd 0.009621f
C6420 vdd.n3464 gnd 0.007744f
C6421 vdd.n3465 gnd 0.009621f
C6422 vdd.n3466 gnd 0.693161f
C6423 vdd.n3467 gnd 0.009621f
C6424 vdd.n3468 gnd 0.007744f
C6425 vdd.n3469 gnd 0.009621f
C6426 vdd.n3470 gnd 0.009621f
C6427 vdd.n3471 gnd 0.009621f
C6428 vdd.n3472 gnd 0.009621f
C6429 vdd.n3473 gnd 0.009621f
C6430 vdd.n3474 gnd 0.007744f
C6431 vdd.n3475 gnd 0.007744f
C6432 vdd.n3476 gnd 0.009621f
C6433 vdd.t141 gnd 0.491603f
C6434 vdd.n3477 gnd 0.816061f
C6435 vdd.n3478 gnd 0.009621f
C6436 vdd.n3479 gnd 0.007744f
C6437 vdd.n3480 gnd 0.009621f
C6438 vdd.n3481 gnd 0.009621f
C6439 vdd.n3482 gnd 0.009621f
C6440 vdd.n3483 gnd 0.007744f
C6441 vdd.n3484 gnd 0.009621f
C6442 vdd.n3485 gnd 0.771817f
C6443 vdd.n3486 gnd 0.009621f
C6444 vdd.n3487 gnd 0.009621f
C6445 vdd.n3488 gnd 0.007744f
C6446 vdd.n3489 gnd 0.007744f
C6447 vdd.n3490 gnd 0.007744f
C6448 vdd.n3491 gnd 0.009621f
C6449 vdd.n3492 gnd 0.009621f
C6450 vdd.n3493 gnd 0.009621f
C6451 vdd.n3494 gnd 0.009621f
C6452 vdd.n3495 gnd 0.007744f
C6453 vdd.n3496 gnd 0.007744f
C6454 vdd.n3497 gnd 0.007744f
C6455 vdd.n3498 gnd 0.009621f
C6456 vdd.n3499 gnd 0.009621f
C6457 vdd.n3500 gnd 0.009621f
C6458 vdd.n3501 gnd 0.009621f
C6459 vdd.n3502 gnd 0.007744f
C6460 vdd.n3503 gnd 0.007744f
C6461 vdd.n3504 gnd 0.007744f
C6462 vdd.n3505 gnd 0.009621f
C6463 vdd.n3506 gnd 0.009621f
C6464 vdd.n3507 gnd 0.009621f
C6465 vdd.n3508 gnd 0.816061f
C6466 vdd.n3509 gnd 0.009621f
C6467 vdd.n3510 gnd 0.007744f
C6468 vdd.n3511 gnd 0.007744f
C6469 vdd.n3512 gnd 0.007744f
C6470 vdd.n3513 gnd 0.009621f
C6471 vdd.n3514 gnd 0.009621f
C6472 vdd.n3515 gnd 0.009621f
C6473 vdd.n3516 gnd 0.009621f
C6474 vdd.n3517 gnd 0.007744f
C6475 vdd.n3518 gnd 0.007744f
C6476 vdd.n3519 gnd 0.006427f
C6477 vdd.n3520 gnd 0.021909f
C6478 vdd.n3521 gnd 0.022059f
C6479 vdd.n3522 gnd 0.003678f
C6480 vdd.n3523 gnd 0.022059f
C6481 vdd.n3525 gnd 2.17289f
C6482 vdd.n3526 gnd 1.29783f
C6483 vdd.n3527 gnd 0.644f
C6484 vdd.n3528 gnd 0.009621f
C6485 vdd.n3529 gnd 0.007744f
C6486 vdd.n3530 gnd 0.007744f
C6487 vdd.n3531 gnd 0.007744f
C6488 vdd.n3532 gnd 0.009621f
C6489 vdd.n3533 gnd 0.983206f
C6490 vdd.n3534 gnd 0.983206f
C6491 vdd.n3535 gnd 0.565344f
C6492 vdd.n3536 gnd 0.009621f
C6493 vdd.n3537 gnd 0.007744f
C6494 vdd.n3538 gnd 0.007744f
C6495 vdd.n3539 gnd 0.007744f
C6496 vdd.n3540 gnd 0.009621f
C6497 vdd.n3541 gnd 0.585008f
C6498 vdd.n3542 gnd 0.722657f
C6499 vdd.t29 gnd 0.491603f
C6500 vdd.n3543 gnd 0.752153f
C6501 vdd.n3544 gnd 0.009621f
C6502 vdd.n3545 gnd 0.007744f
C6503 vdd.n3546 gnd 0.007744f
C6504 vdd.n3547 gnd 0.007744f
C6505 vdd.n3548 gnd 0.009621f
C6506 vdd.n3549 gnd 0.816061f
C6507 vdd.t6 gnd 0.491603f
C6508 vdd.n3550 gnd 0.59484f
C6509 vdd.n3551 gnd 0.712825f
C6510 vdd.n3552 gnd 0.009621f
C6511 vdd.n3553 gnd 0.007744f
C6512 vdd.n3554 gnd 0.007744f
C6513 vdd.n3555 gnd 0.007744f
C6514 vdd.n3556 gnd 0.009621f
C6515 vdd.n3557 gnd 0.54568f
C6516 vdd.t0 gnd 0.491603f
C6517 vdd.n3558 gnd 0.816061f
C6518 vdd.t169 gnd 0.491603f
C6519 vdd.n3559 gnd 0.604672f
C6520 vdd.n3560 gnd 0.009621f
C6521 vdd.n3561 gnd 0.007744f
C6522 vdd.n3562 gnd 0.007394f
C6523 vdd.n3563 gnd 0.567475f
C6524 vdd.n3564 gnd 2.64002f
C6525 a_n2804_13878.t23 gnd 0.194556f
C6526 a_n2804_13878.t10 gnd 0.194556f
C6527 a_n2804_13878.t20 gnd 0.194556f
C6528 a_n2804_13878.n0 gnd 1.53358f
C6529 a_n2804_13878.t25 gnd 0.194556f
C6530 a_n2804_13878.t15 gnd 0.194556f
C6531 a_n2804_13878.n1 gnd 1.53196f
C6532 a_n2804_13878.n2 gnd 2.14061f
C6533 a_n2804_13878.t21 gnd 0.194556f
C6534 a_n2804_13878.t14 gnd 0.194556f
C6535 a_n2804_13878.n3 gnd 1.53196f
C6536 a_n2804_13878.n4 gnd 1.04414f
C6537 a_n2804_13878.t8 gnd 0.194556f
C6538 a_n2804_13878.t11 gnd 0.194556f
C6539 a_n2804_13878.n5 gnd 1.53196f
C6540 a_n2804_13878.n6 gnd 1.04414f
C6541 a_n2804_13878.t24 gnd 0.194556f
C6542 a_n2804_13878.t9 gnd 0.194556f
C6543 a_n2804_13878.n7 gnd 1.53196f
C6544 a_n2804_13878.n8 gnd 1.04414f
C6545 a_n2804_13878.t19 gnd 0.194556f
C6546 a_n2804_13878.t7 gnd 0.194556f
C6547 a_n2804_13878.n9 gnd 1.53196f
C6548 a_n2804_13878.n10 gnd 4.90178f
C6549 a_n2804_13878.t1 gnd 1.82172f
C6550 a_n2804_13878.t4 gnd 0.194556f
C6551 a_n2804_13878.t31 gnd 0.194556f
C6552 a_n2804_13878.n11 gnd 1.37045f
C6553 a_n2804_13878.n12 gnd 1.53128f
C6554 a_n2804_13878.t0 gnd 1.81809f
C6555 a_n2804_13878.n13 gnd 0.770559f
C6556 a_n2804_13878.t5 gnd 1.81809f
C6557 a_n2804_13878.n14 gnd 0.770559f
C6558 a_n2804_13878.t30 gnd 0.194556f
C6559 a_n2804_13878.t3 gnd 0.194556f
C6560 a_n2804_13878.n15 gnd 1.37045f
C6561 a_n2804_13878.n16 gnd 0.778022f
C6562 a_n2804_13878.t2 gnd 1.81809f
C6563 a_n2804_13878.n17 gnd 2.85814f
C6564 a_n2804_13878.n18 gnd 3.74876f
C6565 a_n2804_13878.t13 gnd 0.194556f
C6566 a_n2804_13878.t22 gnd 0.194556f
C6567 a_n2804_13878.n19 gnd 1.53195f
C6568 a_n2804_13878.n20 gnd 2.50239f
C6569 a_n2804_13878.t26 gnd 0.194556f
C6570 a_n2804_13878.t12 gnd 0.194556f
C6571 a_n2804_13878.n21 gnd 1.53196f
C6572 a_n2804_13878.n22 gnd 0.678771f
C6573 a_n2804_13878.t16 gnd 0.194556f
C6574 a_n2804_13878.t17 gnd 0.194556f
C6575 a_n2804_13878.n23 gnd 1.53196f
C6576 a_n2804_13878.n24 gnd 0.678771f
C6577 a_n2804_13878.t27 gnd 0.194556f
C6578 a_n2804_13878.t28 gnd 0.194556f
C6579 a_n2804_13878.n25 gnd 1.53196f
C6580 a_n2804_13878.n26 gnd 0.678771f
C6581 a_n2804_13878.t6 gnd 0.194556f
C6582 a_n2804_13878.t18 gnd 0.194556f
C6583 a_n2804_13878.n27 gnd 1.53196f
C6584 a_n2804_13878.n28 gnd 1.37704f
C6585 a_n2804_13878.n29 gnd 1.5345f
C6586 a_n2804_13878.t29 gnd 0.194556f
C6587 a_n2982_13878.n0 gnd 0.883913f
C6588 a_n2982_13878.n1 gnd 3.58469f
C6589 a_n2982_13878.n2 gnd 3.31432f
C6590 a_n2982_13878.n3 gnd 3.91444f
C6591 a_n2982_13878.n4 gnd 0.902552f
C6592 a_n2982_13878.n5 gnd 0.198406f
C6593 a_n2982_13878.n6 gnd 0.14613f
C6594 a_n2982_13878.n7 gnd 0.22967f
C6595 a_n2982_13878.n8 gnd 0.177393f
C6596 a_n2982_13878.n9 gnd 0.198406f
C6597 a_n2982_13878.n10 gnd 1.32168f
C6598 a_n2982_13878.n11 gnd 0.14613f
C6599 a_n2982_13878.n12 gnd 0.954828f
C6600 a_n2982_13878.n13 gnd 0.209105f
C6601 a_n2982_13878.n14 gnd 0.735977f
C6602 a_n2982_13878.n15 gnd 0.209105f
C6603 a_n2982_13878.n16 gnd 0.209105f
C6604 a_n2982_13878.n17 gnd 0.476233f
C6605 a_n2982_13878.n18 gnd 0.274168f
C6606 a_n2982_13878.n19 gnd 0.209105f
C6607 a_n2982_13878.n20 gnd 0.528509f
C6608 a_n2982_13878.n21 gnd 0.209105f
C6609 a_n2982_13878.n22 gnd 0.209105f
C6610 a_n2982_13878.n23 gnd 0.930364f
C6611 a_n2982_13878.n24 gnd 0.274168f
C6612 a_n2982_13878.n25 gnd 0.970217f
C6613 a_n2982_13878.n26 gnd 0.209105f
C6614 a_n2982_13878.n27 gnd 0.209105f
C6615 a_n2982_13878.n28 gnd 0.476233f
C6616 a_n2982_13878.n29 gnd 0.209105f
C6617 a_n2982_13878.n30 gnd 0.274168f
C6618 a_n2982_13878.n31 gnd 3.21642f
C6619 a_n2982_13878.n32 gnd 0.104552f
C6620 a_n2982_13878.n33 gnd 0.209105f
C6621 a_n2982_13878.n34 gnd 0.842549f
C6622 a_n2982_13878.n35 gnd 0.209105f
C6623 a_n2982_13878.n36 gnd 0.274168f
C6624 a_n2982_13878.n37 gnd 1.72153f
C6625 a_n2982_13878.n38 gnd 1.16f
C6626 a_n2982_13878.n39 gnd 2.31679f
C6627 a_n2982_13878.n40 gnd 1.16f
C6628 a_n2982_13878.n41 gnd 2.11818f
C6629 a_n2982_13878.n42 gnd 1.72153f
C6630 a_n2982_13878.n43 gnd 0.00839f
C6631 a_n2982_13878.n44 gnd 4.04e-19
C6632 a_n2982_13878.n46 gnd 0.008096f
C6633 a_n2982_13878.n47 gnd 0.011772f
C6634 a_n2982_13878.n48 gnd 0.007788f
C6635 a_n2982_13878.n49 gnd 0.277359f
C6636 a_n2982_13878.n50 gnd 0.00839f
C6637 a_n2982_13878.n51 gnd 4.04e-19
C6638 a_n2982_13878.n53 gnd 0.008096f
C6639 a_n2982_13878.n54 gnd 0.011772f
C6640 a_n2982_13878.n55 gnd 0.007788f
C6641 a_n2982_13878.n57 gnd 0.277359f
C6642 a_n2982_13878.n58 gnd 0.00839f
C6643 a_n2982_13878.n59 gnd 4.04e-19
C6644 a_n2982_13878.n61 gnd 0.008096f
C6645 a_n2982_13878.n62 gnd 0.011772f
C6646 a_n2982_13878.n63 gnd 0.007788f
C6647 a_n2982_13878.n65 gnd 0.277359f
C6648 a_n2982_13878.n66 gnd 0.00839f
C6649 a_n2982_13878.n67 gnd 4.04e-19
C6650 a_n2982_13878.n69 gnd 0.008096f
C6651 a_n2982_13878.n70 gnd 0.011772f
C6652 a_n2982_13878.n71 gnd 0.007788f
C6653 a_n2982_13878.n73 gnd 0.277359f
C6654 a_n2982_13878.n74 gnd 0.008096f
C6655 a_n2982_13878.n75 gnd 0.276227f
C6656 a_n2982_13878.n76 gnd 0.008096f
C6657 a_n2982_13878.n77 gnd 0.276227f
C6658 a_n2982_13878.n78 gnd 0.008096f
C6659 a_n2982_13878.n79 gnd 0.276227f
C6660 a_n2982_13878.n80 gnd 0.008096f
C6661 a_n2982_13878.n81 gnd 0.276227f
C6662 a_n2982_13878.n83 gnd 0.296601f
C6663 a_n2982_13878.t17 gnd 0.688688f
C6664 a_n2982_13878.t23 gnd 0.674643f
C6665 a_n2982_13878.t21 gnd 0.674643f
C6666 a_n2982_13878.t63 gnd 0.674643f
C6667 a_n2982_13878.n84 gnd 0.296483f
C6668 a_n2982_13878.t25 gnd 0.674643f
C6669 a_n2982_13878.t57 gnd 0.674643f
C6670 a_n2982_13878.t61 gnd 0.674643f
C6671 a_n2982_13878.n85 gnd 0.292849f
C6672 a_n2982_13878.t59 gnd 0.674643f
C6673 a_n2982_13878.t45 gnd 0.674643f
C6674 a_n2982_13878.t51 gnd 0.674643f
C6675 a_n2982_13878.t31 gnd 0.685497f
C6676 a_n2982_13878.t106 gnd 0.688688f
C6677 a_n2982_13878.t83 gnd 0.674643f
C6678 a_n2982_13878.t88 gnd 0.674643f
C6679 a_n2982_13878.t76 gnd 0.674643f
C6680 a_n2982_13878.n86 gnd 0.296483f
C6681 a_n2982_13878.t93 gnd 0.674643f
C6682 a_n2982_13878.t102 gnd 0.674643f
C6683 a_n2982_13878.t103 gnd 0.674643f
C6684 a_n2982_13878.n87 gnd 0.292849f
C6685 a_n2982_13878.t70 gnd 0.674643f
C6686 a_n2982_13878.t85 gnd 0.674643f
C6687 a_n2982_13878.t73 gnd 0.674643f
C6688 a_n2982_13878.n88 gnd 0.296601f
C6689 a_n2982_13878.t80 gnd 0.674643f
C6690 a_n2982_13878.t99 gnd 0.685497f
C6691 a_n2982_13878.t50 gnd 1.35806f
C6692 a_n2982_13878.t34 gnd 0.145037f
C6693 a_n2982_13878.t40 gnd 0.145037f
C6694 a_n2982_13878.n89 gnd 1.02164f
C6695 a_n2982_13878.t38 gnd 0.145037f
C6696 a_n2982_13878.t44 gnd 0.145037f
C6697 a_n2982_13878.n90 gnd 1.02164f
C6698 a_n2982_13878.t48 gnd 0.145037f
C6699 a_n2982_13878.t28 gnd 0.145037f
C6700 a_n2982_13878.n91 gnd 1.02164f
C6701 a_n2982_13878.t42 gnd 0.145037f
C6702 a_n2982_13878.t36 gnd 0.145037f
C6703 a_n2982_13878.n92 gnd 1.02164f
C6704 a_n2982_13878.t56 gnd 0.145037f
C6705 a_n2982_13878.t20 gnd 0.145037f
C6706 a_n2982_13878.n93 gnd 1.02164f
C6707 a_n2982_13878.t30 gnd 1.35535f
C6708 a_n2982_13878.t55 gnd 0.674643f
C6709 a_n2982_13878.n94 gnd 0.296601f
C6710 a_n2982_13878.t19 gnd 0.674643f
C6711 a_n2982_13878.t41 gnd 0.674643f
C6712 a_n2982_13878.n95 gnd 0.287692f
C6713 a_n2982_13878.t43 gnd 0.674643f
C6714 a_n2982_13878.n96 gnd 0.29915f
C6715 a_n2982_13878.t47 gnd 0.674643f
C6716 a_n2982_13878.t39 gnd 0.674643f
C6717 a_n2982_13878.n97 gnd 0.292527f
C6718 a_n2982_13878.t49 gnd 0.688688f
C6719 a_n2982_13878.t82 gnd 0.674643f
C6720 a_n2982_13878.n98 gnd 0.296601f
C6721 a_n2982_13878.t91 gnd 0.674643f
C6722 a_n2982_13878.t97 gnd 0.674643f
C6723 a_n2982_13878.n99 gnd 0.287692f
C6724 a_n2982_13878.t101 gnd 0.674643f
C6725 a_n2982_13878.n100 gnd 0.29915f
C6726 a_n2982_13878.t72 gnd 0.674643f
C6727 a_n2982_13878.t75 gnd 0.674643f
C6728 a_n2982_13878.n101 gnd 0.292527f
C6729 a_n2982_13878.t105 gnd 0.688688f
C6730 a_n2982_13878.t74 gnd 0.674643f
C6731 a_n2982_13878.n102 gnd 0.298713f
C6732 a_n2982_13878.t100 gnd 0.674643f
C6733 a_n2982_13878.n103 gnd 0.296483f
C6734 a_n2982_13878.n104 gnd 0.296616f
C6735 a_n2982_13878.t96 gnd 0.674643f
C6736 a_n2982_13878.n105 gnd 0.292849f
C6737 a_n2982_13878.t69 gnd 0.674643f
C6738 a_n2982_13878.n106 gnd 0.293101f
C6739 a_n2982_13878.n107 gnd 0.298713f
C6740 a_n2982_13878.t71 gnd 0.685497f
C6741 a_n2982_13878.t33 gnd 0.674643f
C6742 a_n2982_13878.n108 gnd 0.298713f
C6743 a_n2982_13878.t37 gnd 0.674643f
C6744 a_n2982_13878.n109 gnd 0.296483f
C6745 a_n2982_13878.n110 gnd 0.296616f
C6746 a_n2982_13878.t27 gnd 0.674643f
C6747 a_n2982_13878.n111 gnd 0.292849f
C6748 a_n2982_13878.t35 gnd 0.674643f
C6749 a_n2982_13878.n112 gnd 0.293101f
C6750 a_n2982_13878.n113 gnd 0.298713f
C6751 a_n2982_13878.t29 gnd 0.685497f
C6752 a_n2982_13878.n114 gnd 1.30619f
C6753 a_n2982_13878.t79 gnd 0.674643f
C6754 a_n2982_13878.n115 gnd 0.292849f
C6755 a_n2982_13878.t87 gnd 0.674643f
C6756 a_n2982_13878.n116 gnd 0.292849f
C6757 a_n2982_13878.t77 gnd 0.674643f
C6758 a_n2982_13878.n117 gnd 0.292849f
C6759 a_n2982_13878.t92 gnd 0.674643f
C6760 a_n2982_13878.n118 gnd 0.292849f
C6761 a_n2982_13878.t81 gnd 0.674643f
C6762 a_n2982_13878.n119 gnd 0.287531f
C6763 a_n2982_13878.t107 gnd 0.674643f
C6764 a_n2982_13878.n120 gnd 0.296616f
C6765 a_n2982_13878.t84 gnd 0.685948f
C6766 a_n2982_13878.t94 gnd 0.674643f
C6767 a_n2982_13878.n121 gnd 0.287531f
C6768 a_n2982_13878.t78 gnd 0.674643f
C6769 a_n2982_13878.n122 gnd 0.296616f
C6770 a_n2982_13878.t89 gnd 0.685948f
C6771 a_n2982_13878.t98 gnd 0.674643f
C6772 a_n2982_13878.n123 gnd 0.287531f
C6773 a_n2982_13878.t86 gnd 0.674643f
C6774 a_n2982_13878.n124 gnd 0.296616f
C6775 a_n2982_13878.t104 gnd 0.685948f
C6776 a_n2982_13878.t90 gnd 0.674643f
C6777 a_n2982_13878.n125 gnd 0.287531f
C6778 a_n2982_13878.t68 gnd 0.674643f
C6779 a_n2982_13878.n126 gnd 0.296616f
C6780 a_n2982_13878.t95 gnd 0.685948f
C6781 a_n2982_13878.n127 gnd 1.64303f
C6782 a_n2982_13878.n128 gnd 0.298713f
C6783 a_n2982_13878.n129 gnd 0.293101f
C6784 a_n2982_13878.n130 gnd 0.287692f
C6785 a_n2982_13878.n131 gnd 0.296616f
C6786 a_n2982_13878.n132 gnd 0.29915f
C6787 a_n2982_13878.n133 gnd 0.292527f
C6788 a_n2982_13878.n134 gnd 0.298713f
C6789 a_n2982_13878.t53 gnd 0.674643f
C6790 a_n2982_13878.n135 gnd 0.298713f
C6791 a_n2982_13878.t3 gnd 0.112807f
C6792 a_n2982_13878.t66 gnd 0.112807f
C6793 a_n2982_13878.n136 gnd 0.999739f
C6794 a_n2982_13878.t0 gnd 0.112807f
C6795 a_n2982_13878.t16 gnd 0.112807f
C6796 a_n2982_13878.n137 gnd 0.9968f
C6797 a_n2982_13878.t2 gnd 0.112807f
C6798 a_n2982_13878.t5 gnd 0.112807f
C6799 a_n2982_13878.n138 gnd 0.9968f
C6800 a_n2982_13878.t10 gnd 0.112807f
C6801 a_n2982_13878.t11 gnd 0.112807f
C6802 a_n2982_13878.n139 gnd 0.999739f
C6803 a_n2982_13878.t15 gnd 0.112807f
C6804 a_n2982_13878.t12 gnd 0.112807f
C6805 a_n2982_13878.n140 gnd 0.9968f
C6806 a_n2982_13878.t1 gnd 0.112807f
C6807 a_n2982_13878.t67 gnd 0.112807f
C6808 a_n2982_13878.n141 gnd 0.996801f
C6809 a_n2982_13878.t9 gnd 0.112807f
C6810 a_n2982_13878.t14 gnd 0.112807f
C6811 a_n2982_13878.n142 gnd 0.996801f
C6812 a_n2982_13878.t6 gnd 0.112807f
C6813 a_n2982_13878.t4 gnd 0.112807f
C6814 a_n2982_13878.n143 gnd 0.996801f
C6815 a_n2982_13878.t65 gnd 0.112807f
C6816 a_n2982_13878.t13 gnd 0.112807f
C6817 a_n2982_13878.n144 gnd 0.99974f
C6818 a_n2982_13878.t8 gnd 0.112807f
C6819 a_n2982_13878.t7 gnd 0.112807f
C6820 a_n2982_13878.n145 gnd 0.996801f
C6821 a_n2982_13878.n146 gnd 0.293101f
C6822 a_n2982_13878.n147 gnd 0.287692f
C6823 a_n2982_13878.n148 gnd 0.296616f
C6824 a_n2982_13878.n149 gnd 0.29915f
C6825 a_n2982_13878.n150 gnd 0.292527f
C6826 a_n2982_13878.n151 gnd 0.298713f
C6827 a_n2982_13878.n152 gnd 0.993167f
C6828 a_n2982_13878.t32 gnd 1.35806f
C6829 a_n2982_13878.t52 gnd 0.145037f
C6830 a_n2982_13878.t54 gnd 0.145037f
C6831 a_n2982_13878.n153 gnd 1.02164f
C6832 a_n2982_13878.t60 gnd 0.145037f
C6833 a_n2982_13878.t46 gnd 0.145037f
C6834 a_n2982_13878.n154 gnd 1.02164f
C6835 a_n2982_13878.t58 gnd 0.145037f
C6836 a_n2982_13878.t62 gnd 0.145037f
C6837 a_n2982_13878.n155 gnd 1.02164f
C6838 a_n2982_13878.t64 gnd 0.145037f
C6839 a_n2982_13878.t26 gnd 0.145037f
C6840 a_n2982_13878.n156 gnd 1.02164f
C6841 a_n2982_13878.t24 gnd 0.145037f
C6842 a_n2982_13878.t22 gnd 0.145037f
C6843 a_n2982_13878.n157 gnd 1.02164f
C6844 a_n2982_13878.t18 gnd 1.35535f
.ends

