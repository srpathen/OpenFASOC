* NGSPICE file created from opamp517.ext - technology: sky130A

.subckt opamp517 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n6972_8799.t30 plus.t5 a_n3827_n3924.t33 gnd.t118 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X1 CSoutput.t141 a_n6972_8799.t32 vdd.t255 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X2 a_n1808_13878.t7 a_n1996_n452.t44 vdd.t118 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 a_n1808_13878.t19 a_n1996_n452.t37 a_n1996_n452.t38 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 vdd.t254 a_n6972_8799.t33 CSoutput.t140 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X5 CSoutput.t139 a_n6972_8799.t34 vdd.t253 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 vdd.t98 vdd.t96 vdd.t97 vdd.t32 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X7 outputibias.t7 outputibias.t6 gnd.t181 gnd.t180 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X8 gnd.t334 gnd.t332 plus.t1 gnd.t333 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X9 a_n3827_n3924.t20 diffpairibias.t20 gnd.t134 gnd.t133 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X10 gnd.t86 commonsourceibias.t80 CSoutput.t27 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 gnd.t331 gnd.t329 gnd.t330 gnd.t310 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X12 CSoutput.t138 a_n6972_8799.t35 vdd.t252 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X13 commonsourceibias.t79 commonsourceibias.t78 gnd.t219 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X14 a_n3827_n3924.t26 plus.t6 a_n6972_8799.t29 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X15 commonsourceibias.t77 commonsourceibias.t76 gnd.t89 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 gnd.t328 gnd.t326 gnd.t327 gnd.t310 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X17 a_n3827_n3924.t46 minus.t5 a_n1996_n452.t43 gnd.t337 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X18 vdd.t123 CSoutput.t176 output.t15 gnd.t162 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X19 a_n1986_8322.t21 a_n1996_n452.t45 a_n6972_8799.t4 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X20 gnd.t325 gnd.t323 gnd.t324 gnd.t242 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X21 CSoutput.t28 commonsourceibias.t81 gnd.t87 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 CSoutput.t137 a_n6972_8799.t36 vdd.t251 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X23 gnd.t62 commonsourceibias.t74 commonsourceibias.t75 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X24 CSoutput.t151 commonsourceibias.t82 gnd.t194 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 vdd.t250 a_n6972_8799.t37 CSoutput.t136 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X26 gnd.t322 gnd.t320 gnd.t321 gnd.t242 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X27 a_n1996_n452.t7 minus.t6 a_n3827_n3924.t8 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X28 commonsourceibias.t73 commonsourceibias.t72 gnd.t202 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X29 vdd.t124 CSoutput.t177 output.t14 gnd.t163 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X30 CSoutput.t152 commonsourceibias.t83 gnd.t195 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X31 vdd.t249 a_n6972_8799.t38 CSoutput.t135 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X32 a_n1996_n452.t6 minus.t7 a_n3827_n3924.t6 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X33 CSoutput.t134 a_n6972_8799.t39 vdd.t248 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X34 vdd.t247 a_n6972_8799.t40 CSoutput.t133 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X35 a_n6972_8799.t3 a_n1996_n452.t46 a_n1986_8322.t20 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X36 CSoutput.t132 a_n6972_8799.t41 vdd.t246 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X37 gnd.t319 gnd.t316 gnd.t318 gnd.t317 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X38 commonsourceibias.t71 commonsourceibias.t70 gnd.t101 gnd.t100 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X39 a_n3827_n3924.t22 minus.t8 a_n1996_n452.t16 gnd.t137 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X40 CSoutput.t131 a_n6972_8799.t42 vdd.t245 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X41 vdd.t95 vdd.t93 vdd.t94 vdd.t28 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X42 a_n3827_n3924.t25 diffpairibias.t21 gnd.t225 gnd.t224 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X43 CSoutput.t158 commonsourceibias.t84 gnd.t217 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X44 CSoutput.t130 a_n6972_8799.t43 vdd.t244 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X45 vdd.t92 vdd.t90 vdd.t91 vdd.t32 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X46 gnd.t218 commonsourceibias.t85 CSoutput.t159 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X47 gnd.t315 gnd.t313 gnd.t314 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X48 gnd.t148 commonsourceibias.t68 commonsourceibias.t69 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 CSoutput.t129 a_n6972_8799.t44 vdd.t227 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X50 commonsourceibias.t67 commonsourceibias.t66 gnd.t103 gnd.t102 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 a_n3827_n3924.t41 plus.t7 a_n6972_8799.t28 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X52 gnd.t84 commonsourceibias.t86 CSoutput.t25 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X53 vdd.t243 a_n6972_8799.t45 CSoutput.t128 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X54 a_n1808_13878.t18 a_n1996_n452.t27 a_n1996_n452.t28 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X55 gnd.t85 commonsourceibias.t87 CSoutput.t26 gnd.t74 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 CSoutput.t127 a_n6972_8799.t46 vdd.t242 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X57 a_n1996_n452.t40 a_n1996_n452.t39 a_n1808_13878.t17 vdd.t99 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X58 gnd.t192 commonsourceibias.t88 CSoutput.t149 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X59 a_n6972_8799.t27 plus.t8 a_n3827_n3924.t42 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X60 CSoutput.t126 a_n6972_8799.t47 vdd.t241 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 output.t13 CSoutput.t178 vdd.t19 gnd.t80 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X62 vdd.t89 vdd.t87 vdd.t88 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X63 vdd.t240 a_n6972_8799.t48 CSoutput.t125 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X64 gnd.t149 commonsourceibias.t64 commonsourceibias.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X65 diffpairibias.t19 diffpairibias.t18 gnd.t48 gnd.t47 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X66 commonsourceibias.t63 commonsourceibias.t62 gnd.t203 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 a_n1996_n452.t2 minus.t9 a_n3827_n3924.t2 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X68 CSoutput.t124 a_n6972_8799.t49 vdd.t239 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X69 commonsourceibias.t61 commonsourceibias.t60 gnd.t204 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 vdd.t238 a_n6972_8799.t50 CSoutput.t123 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 vdd.t237 a_n6972_8799.t51 CSoutput.t122 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 vdd.t235 a_n6972_8799.t52 CSoutput.t121 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X73 gnd.t312 gnd.t309 gnd.t311 gnd.t310 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X74 plus.t0 gnd.t306 gnd.t308 gnd.t307 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X75 diffpairibias.t17 diffpairibias.t16 gnd.t197 gnd.t196 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X76 gnd.t104 commonsourceibias.t58 commonsourceibias.t59 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X77 CSoutput.t120 a_n6972_8799.t53 vdd.t234 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X78 CSoutput.t119 a_n6972_8799.t54 vdd.t233 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X79 CSoutput.t150 commonsourceibias.t89 gnd.t193 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 gnd.t305 gnd.t303 gnd.t304 gnd.t250 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X81 vdd.t232 a_n6972_8799.t55 CSoutput.t118 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 CSoutput.t117 a_n6972_8799.t56 vdd.t231 vdd.t218 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 CSoutput.t156 commonsourceibias.t90 gnd.t215 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 CSoutput.t116 a_n6972_8799.t57 vdd.t228 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X85 CSoutput.t115 a_n6972_8799.t58 vdd.t230 vdd.t218 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 gnd.t63 commonsourceibias.t56 commonsourceibias.t57 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 vdd.t20 CSoutput.t179 output.t12 gnd.t81 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X88 CSoutput.t157 commonsourceibias.t91 gnd.t216 gnd.t102 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 CSoutput.t169 commonsourceibias.t92 gnd.t345 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 vdd.t229 a_n6972_8799.t59 CSoutput.t114 vdd.t216 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X91 a_n3827_n3924.t43 plus.t9 a_n6972_8799.t26 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X92 CSoutput.t170 commonsourceibias.t93 gnd.t346 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X93 CSoutput.t11 commonsourceibias.t94 gnd.t42 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 a_n3827_n3924.t10 diffpairibias.t22 gnd.t93 gnd.t92 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X95 a_n1996_n452.t34 a_n1996_n452.t33 a_n1808_13878.t16 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X96 vdd.t226 a_n6972_8799.t60 CSoutput.t113 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X97 output.t11 CSoutput.t180 vdd.t21 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X98 a_n6972_8799.t5 a_n1996_n452.t47 a_n1986_8322.t19 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X99 vdd.t225 a_n6972_8799.t61 CSoutput.t112 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X100 a_n1996_n452.t24 a_n1996_n452.t23 a_n1808_13878.t15 vdd.t105 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X101 vdd.t224 a_n6972_8799.t62 CSoutput.t111 vdd.t216 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 gnd.t205 commonsourceibias.t54 commonsourceibias.t55 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X103 gnd.t106 commonsourceibias.t52 commonsourceibias.t53 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 gnd.t150 commonsourceibias.t50 commonsourceibias.t51 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X105 output.t19 outputibias.t8 gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X106 CSoutput.t181 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X107 vdd.t223 a_n6972_8799.t63 CSoutput.t110 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X108 CSoutput.t109 a_n6972_8799.t64 vdd.t222 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X109 gnd.t302 gnd.t299 gnd.t301 gnd.t300 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X110 diffpairibias.t15 diffpairibias.t14 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X111 a_n1996_n452.t5 minus.t10 a_n3827_n3924.t5 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X112 output.t18 outputibias.t9 gnd.t336 gnd.t335 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X113 vdd.t86 vdd.t84 vdd.t85 vdd.t71 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X114 vdd.t221 a_n6972_8799.t65 CSoutput.t108 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X115 CSoutput.t107 a_n6972_8799.t66 vdd.t220 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X116 gnd.t44 commonsourceibias.t95 CSoutput.t12 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 vdd.t83 vdd.t80 vdd.t82 vdd.t81 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X118 gnd.t5 commonsourceibias.t96 CSoutput.t1 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X119 gnd.t7 commonsourceibias.t97 CSoutput.t2 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 gnd.t73 commonsourceibias.t98 CSoutput.t23 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X121 a_n3827_n3924.t9 minus.t11 a_n1996_n452.t8 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X122 vdd.t79 vdd.t77 vdd.t78 vdd.t24 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X123 gnd.t75 commonsourceibias.t99 CSoutput.t24 gnd.t74 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X124 output.t10 CSoutput.t182 vdd.t125 gnd.t166 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X125 vdd.t76 vdd.t74 vdd.t75 vdd.t67 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X126 vdd.t126 CSoutput.t183 output.t9 gnd.t167 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X127 vdd.t257 a_n1996_n452.t48 a_n1986_8322.t9 vdd.t256 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X128 gnd.t351 commonsourceibias.t100 CSoutput.t173 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X129 gnd.t298 gnd.t296 gnd.t297 gnd.t246 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X130 a_n1986_8322.t8 a_n1996_n452.t49 vdd.t110 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X131 a_n3827_n3924.t48 diffpairibias.t23 gnd.t354 gnd.t353 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X132 CSoutput.t106 a_n6972_8799.t67 vdd.t219 vdd.t218 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X133 gnd.t295 gnd.t293 gnd.t294 gnd.t257 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X134 CSoutput.t174 commonsourceibias.t101 gnd.t352 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X135 vdd.t217 a_n6972_8799.t68 CSoutput.t105 vdd.t216 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X136 a_n3827_n3924.t24 minus.t12 a_n1996_n452.t18 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X137 gnd.t206 commonsourceibias.t48 commonsourceibias.t49 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 vdd.t104 a_n1996_n452.t50 a_n1808_13878.t6 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X139 a_n1996_n452.t4 minus.t13 a_n3827_n3924.t4 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X140 a_n3827_n3924.t28 plus.t10 a_n6972_8799.t25 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X141 a_n3827_n3924.t32 plus.t11 a_n6972_8799.t24 gnd.t128 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X142 gnd.t30 commonsourceibias.t102 CSoutput.t8 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X143 vdd.t73 vdd.t70 vdd.t72 vdd.t71 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X144 vdd.t215 a_n6972_8799.t69 CSoutput.t104 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X145 vdd.t69 vdd.t66 vdd.t68 vdd.t67 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X146 gnd.t151 commonsourceibias.t46 commonsourceibias.t47 gnd.t74 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X147 a_n6972_8799.t23 plus.t12 a_n3827_n3924.t39 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X148 a_n6972_8799.t22 plus.t13 a_n3827_n3924.t30 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X149 vdd.t65 vdd.t62 vdd.t64 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X150 a_n1986_8322.t7 a_n1996_n452.t51 vdd.t259 vdd.t258 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X151 a_n6972_8799.t6 a_n1996_n452.t52 a_n1986_8322.t18 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X152 diffpairibias.t13 diffpairibias.t12 gnd.t132 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X153 CSoutput.t184 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X154 CSoutput.t9 commonsourceibias.t103 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X155 a_n1996_n452.t17 minus.t14 a_n3827_n3924.t23 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X156 a_n1996_n452.t26 a_n1996_n452.t25 a_n1808_13878.t14 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X157 vdd.t213 a_n6972_8799.t70 CSoutput.t103 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X158 a_n6972_8799.t2 a_n1996_n452.t53 a_n1986_8322.t17 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X159 CSoutput.t102 a_n6972_8799.t71 vdd.t212 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X160 CSoutput.t144 commonsourceibias.t104 gnd.t186 gnd.t102 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 commonsourceibias.t45 commonsourceibias.t44 gnd.t34 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X162 CSoutput.t32 commonsourceibias.t105 gnd.t122 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X163 a_n1808_13878.t13 a_n1996_n452.t35 a_n1996_n452.t36 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X164 gnd.t292 gnd.t290 minus.t4 gnd.t291 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X165 gnd.t226 commonsourceibias.t106 CSoutput.t161 gnd.t142 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X166 a_n3827_n3924.t12 minus.t15 a_n1996_n452.t10 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X167 CSoutput.t148 commonsourceibias.t107 gnd.t191 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 vdd.t127 CSoutput.t185 output.t8 gnd.t168 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X169 CSoutput.t5 commonsourceibias.t108 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X170 gnd.t190 commonsourceibias.t109 CSoutput.t147 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X171 CSoutput.t101 a_n6972_8799.t72 vdd.t211 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X172 gnd.t107 commonsourceibias.t42 commonsourceibias.t43 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X173 vdd.t5 a_n1996_n452.t54 a_n1986_8322.t6 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X174 gnd.t40 commonsourceibias.t110 CSoutput.t10 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X175 vdd.t210 a_n6972_8799.t73 CSoutput.t100 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X176 commonsourceibias.t41 commonsourceibias.t40 gnd.t108 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X177 gnd.t152 commonsourceibias.t38 commonsourceibias.t39 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X178 CSoutput.t99 a_n6972_8799.t74 vdd.t209 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X179 vdd.t205 a_n6972_8799.t75 CSoutput.t98 vdd.t134 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X180 a_n3827_n3924.t31 plus.t14 a_n6972_8799.t21 gnd.t337 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X181 gnd.t289 gnd.t287 minus.t3 gnd.t288 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X182 gnd.t207 commonsourceibias.t36 commonsourceibias.t37 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 a_n3827_n3924.t47 diffpairibias.t24 gnd.t348 gnd.t347 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X184 commonsourceibias.t35 commonsourceibias.t34 gnd.t208 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X185 a_n3827_n3924.t7 diffpairibias.t25 gnd.t50 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X186 gnd.t3 commonsourceibias.t111 CSoutput.t0 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 vdd.t208 a_n6972_8799.t76 CSoutput.t97 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X188 a_n6972_8799.t20 plus.t15 a_n3827_n3924.t34 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X189 gnd.t222 commonsourceibias.t112 CSoutput.t160 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X190 gnd.t147 commonsourceibias.t113 CSoutput.t40 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X191 gnd.t350 commonsourceibias.t114 CSoutput.t172 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X192 gnd.t28 commonsourceibias.t115 CSoutput.t7 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X193 CSoutput.t186 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X194 CSoutput.t143 commonsourceibias.t116 gnd.t185 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 commonsourceibias.t33 commonsourceibias.t32 gnd.t109 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 CSoutput.t31 commonsourceibias.t117 gnd.t120 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X197 CSoutput.t96 a_n6972_8799.t77 vdd.t207 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X198 CSoutput.t95 a_n6972_8799.t78 vdd.t204 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X199 CSoutput.t187 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X200 gnd.t146 commonsourceibias.t118 CSoutput.t39 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 CSoutput.t146 commonsourceibias.t119 gnd.t188 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X202 gnd.t286 gnd.t284 gnd.t285 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X203 diffpairibias.t11 diffpairibias.t10 gnd.t356 gnd.t355 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X204 a_n1808_13878.t5 a_n1996_n452.t55 vdd.t261 vdd.t260 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X205 gnd.t187 commonsourceibias.t120 CSoutput.t145 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X206 vdd.t107 a_n1996_n452.t56 a_n1808_13878.t4 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X207 vdd.t61 vdd.t59 vdd.t60 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X208 output.t17 outputibias.t10 gnd.t165 gnd.t164 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X209 gnd.t153 commonsourceibias.t30 commonsourceibias.t31 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 CSoutput.t94 a_n6972_8799.t79 vdd.t203 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X211 gnd.t209 commonsourceibias.t28 commonsourceibias.t29 gnd.t142 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X212 vdd.t201 a_n6972_8799.t80 CSoutput.t93 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X213 commonsourceibias.t27 commonsourceibias.t26 gnd.t154 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X214 CSoutput.t38 commonsourceibias.t121 gnd.t145 gnd.t100 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 diffpairibias.t9 diffpairibias.t8 gnd.t126 gnd.t125 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X216 a_n3827_n3924.t11 minus.t16 a_n1996_n452.t9 gnd.t94 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X217 CSoutput.t92 a_n6972_8799.t81 vdd.t199 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X218 vdd.t197 a_n6972_8799.t82 CSoutput.t91 vdd.t134 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X219 gnd.t223 commonsourceibias.t24 commonsourceibias.t25 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 CSoutput.t37 commonsourceibias.t122 gnd.t144 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X221 a_n1986_8322.t16 a_n1996_n452.t57 a_n6972_8799.t9 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X222 CSoutput.t90 a_n6972_8799.t83 vdd.t196 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X223 diffpairibias.t7 diffpairibias.t6 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X224 vdd.t195 a_n6972_8799.t84 CSoutput.t89 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X225 a_n1996_n452.t15 minus.t17 a_n3827_n3924.t19 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X226 CSoutput.t88 a_n6972_8799.t85 vdd.t193 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X227 a_n1996_n452.t11 minus.t18 a_n3827_n3924.t14 gnd.t118 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X228 gnd.t143 commonsourceibias.t123 CSoutput.t36 gnd.t142 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X229 vdd.t192 a_n6972_8799.t86 CSoutput.t87 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X230 plus.t2 gnd.t281 gnd.t283 gnd.t282 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X231 vdd.t14 a_n1996_n452.t58 a_n1986_8322.t5 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X232 vdd.t185 a_n6972_8799.t87 CSoutput.t86 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X233 vdd.t111 CSoutput.t188 output.t7 gnd.t156 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X234 CSoutput.t35 commonsourceibias.t124 gnd.t141 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 a_n6972_8799.t19 plus.t16 a_n3827_n3924.t36 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X236 CSoutput.t168 commonsourceibias.t125 gnd.t344 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X237 gnd.t280 gnd.t277 gnd.t279 gnd.t278 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X238 gnd.t276 gnd.t274 minus.t2 gnd.t275 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X239 gnd.t343 commonsourceibias.t126 CSoutput.t167 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 a_n3827_n3924.t1 minus.t19 a_n1996_n452.t1 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X241 gnd.t273 gnd.t270 gnd.t272 gnd.t271 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X242 gnd.t342 commonsourceibias.t127 CSoutput.t166 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 a_n1808_13878.t3 a_n1996_n452.t59 vdd.t11 vdd.t10 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X244 CSoutput.t162 commonsourceibias.t128 gnd.t338 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X245 commonsourceibias.t23 commonsourceibias.t22 gnd.t46 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 CSoutput.t165 commonsourceibias.t129 gnd.t341 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X247 vdd.t190 a_n6972_8799.t88 CSoutput.t85 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X248 CSoutput.t84 a_n6972_8799.t89 vdd.t189 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X249 CSoutput.t83 a_n6972_8799.t90 vdd.t188 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X250 gnd.t269 gnd.t267 gnd.t268 gnd.t246 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X251 minus.t1 gnd.t264 gnd.t266 gnd.t265 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X252 vdd.t58 vdd.t56 vdd.t57 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X253 a_n3827_n3924.t49 diffpairibias.t26 gnd.t358 gnd.t357 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X254 vdd.t102 a_n1996_n452.t60 a_n1986_8322.t4 vdd.t101 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X255 a_n1986_8322.t15 a_n1996_n452.t61 a_n6972_8799.t1 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X256 CSoutput.t82 a_n6972_8799.t91 vdd.t187 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X257 gnd.t340 commonsourceibias.t130 CSoutput.t164 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X258 vdd.t184 a_n6972_8799.t92 CSoutput.t81 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X259 vdd.t55 vdd.t53 vdd.t54 vdd.t36 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X260 CSoutput.t80 a_n6972_8799.t93 vdd.t183 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X261 vdd.t182 a_n6972_8799.t94 CSoutput.t79 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X262 vdd.t181 a_n6972_8799.t95 CSoutput.t78 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X263 a_n6972_8799.t18 plus.t17 a_n3827_n3924.t38 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X264 gnd.t174 commonsourceibias.t131 CSoutput.t43 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X265 CSoutput.t163 commonsourceibias.t132 gnd.t339 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X266 vdd.t52 vdd.t49 vdd.t51 vdd.t50 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X267 CSoutput.t22 commonsourceibias.t133 gnd.t71 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X268 a_n3827_n3924.t40 plus.t18 a_n6972_8799.t17 gnd.t137 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X269 gnd.t61 commonsourceibias.t134 CSoutput.t18 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X270 gnd.t69 commonsourceibias.t135 CSoutput.t21 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X271 a_n1808_13878.t12 a_n1996_n452.t19 a_n1996_n452.t20 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X272 CSoutput.t77 a_n6972_8799.t96 vdd.t180 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 vdd.t112 CSoutput.t189 output.t6 gnd.t157 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X274 CSoutput.t17 commonsourceibias.t136 gnd.t60 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 a_n1986_8322.t14 a_n1996_n452.t62 a_n6972_8799.t7 vdd.t99 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X276 diffpairibias.t5 diffpairibias.t4 gnd.t21 gnd.t20 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X277 commonsourceibias.t21 commonsourceibias.t20 gnd.t173 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 gnd.t263 gnd.t260 gnd.t262 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X279 gnd.t67 commonsourceibias.t137 CSoutput.t20 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X280 CSoutput.t16 commonsourceibias.t138 gnd.t58 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X281 gnd.t172 commonsourceibias.t18 commonsourceibias.t19 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X282 CSoutput.t76 a_n6972_8799.t97 vdd.t179 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X283 a_n3827_n3924.t13 diffpairibias.t27 gnd.t117 gnd.t116 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X284 vdd.t177 a_n6972_8799.t98 CSoutput.t75 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 CSoutput.t44 commonsourceibias.t139 gnd.t175 gnd.t100 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 CSoutput.t190 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X287 vdd.t176 a_n6972_8799.t99 CSoutput.t74 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 a_n1986_8322.t3 a_n1996_n452.t63 vdd.t116 vdd.t115 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X289 CSoutput.t73 a_n6972_8799.t100 vdd.t174 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X290 CSoutput.t45 commonsourceibias.t140 gnd.t176 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X291 vdd.t122 a_n1996_n452.t64 a_n1808_13878.t2 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X292 gnd.t36 commonsourceibias.t16 commonsourceibias.t17 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X293 output.t16 outputibias.t11 gnd.t9 gnd.t8 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X294 CSoutput.t72 a_n6972_8799.t101 vdd.t172 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X295 vdd.t48 vdd.t46 vdd.t47 vdd.t36 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X296 CSoutput.t41 commonsourceibias.t141 gnd.t169 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X297 CSoutput.t71 a_n6972_8799.t102 vdd.t170 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X298 gnd.t214 commonsourceibias.t142 CSoutput.t155 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X299 gnd.t259 gnd.t256 gnd.t258 gnd.t257 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X300 vdd.t169 a_n6972_8799.t103 CSoutput.t70 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 vdd.t167 a_n6972_8799.t104 CSoutput.t69 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X302 CSoutput.t154 commonsourceibias.t143 gnd.t213 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X303 vdd.t45 vdd.t42 vdd.t44 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X304 minus.t0 gnd.t253 gnd.t255 gnd.t254 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X305 commonsourceibias.t15 commonsourceibias.t14 gnd.t111 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X306 a_n3827_n3924.t3 minus.t20 a_n1996_n452.t3 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X307 commonsourceibias.t13 commonsourceibias.t12 gnd.t112 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X308 a_n1986_8322.t13 a_n1996_n452.t65 a_n6972_8799.t0 vdd.t1 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X309 CSoutput.t68 a_n6972_8799.t105 vdd.t166 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X310 vdd.t41 vdd.t39 vdd.t40 vdd.t28 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X311 CSoutput.t153 commonsourceibias.t144 gnd.t212 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X312 a_n6972_8799.t8 a_n1996_n452.t66 a_n1986_8322.t12 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X313 gnd.t155 commonsourceibias.t10 commonsourceibias.t11 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 output.t5 CSoutput.t191 vdd.t113 gnd.t158 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X315 vdd.t164 a_n6972_8799.t106 CSoutput.t67 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X316 a_n1808_13878.t1 a_n1996_n452.t67 vdd.t263 vdd.t262 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X317 gnd.t349 commonsourceibias.t145 CSoutput.t171 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X318 CSoutput.t175 commonsourceibias.t146 gnd.t359 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X319 gnd.t252 gnd.t249 gnd.t251 gnd.t250 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X320 vdd.t162 a_n6972_8799.t107 CSoutput.t66 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X321 a_n1996_n452.t0 minus.t21 a_n3827_n3924.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X322 CSoutput.t65 a_n6972_8799.t108 vdd.t161 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X323 gnd.t248 gnd.t245 gnd.t247 gnd.t246 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X324 commonsourceibias.t9 commonsourceibias.t8 gnd.t210 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X325 vdd.t38 vdd.t35 vdd.t37 vdd.t36 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X326 a_n6972_8799.t16 plus.t19 a_n3827_n3924.t35 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X327 vdd.t34 vdd.t31 vdd.t33 vdd.t32 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X328 a_n3827_n3924.t18 minus.t22 a_n1996_n452.t14 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X329 gnd.t211 commonsourceibias.t6 commonsourceibias.t7 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 a_n1808_13878.t11 a_n1996_n452.t29 a_n1996_n452.t30 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X331 CSoutput.t64 a_n6972_8799.t109 vdd.t159 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X332 commonsourceibias.t5 commonsourceibias.t4 gnd.t179 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X333 a_n3827_n3924.t44 plus.t20 a_n6972_8799.t15 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X334 vdd.t158 a_n6972_8799.t110 CSoutput.t63 vdd.t140 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X335 gnd.t184 commonsourceibias.t147 CSoutput.t142 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 CSoutput.t42 commonsourceibias.t148 gnd.t171 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X337 CSoutput.t192 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X338 output.t4 CSoutput.t193 vdd.t114 gnd.t159 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X339 CSoutput.t62 a_n6972_8799.t111 vdd.t157 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 gnd.t139 commonsourceibias.t149 CSoutput.t34 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X341 a_n3827_n3924.t15 diffpairibias.t28 gnd.t124 gnd.t123 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X342 vdd.t156 a_n6972_8799.t112 CSoutput.t61 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X343 gnd.t56 commonsourceibias.t150 CSoutput.t15 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X344 a_n1996_n452.t22 a_n1996_n452.t21 a_n1808_13878.t10 vdd.t1 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X345 gnd.t244 gnd.t241 gnd.t243 gnd.t242 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X346 a_n6972_8799.t10 a_n1996_n452.t68 a_n1986_8322.t11 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X347 vdd.t155 a_n6972_8799.t113 CSoutput.t60 vdd.t140 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X348 output.t3 CSoutput.t194 vdd.t15 gnd.t76 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X349 gnd.t138 commonsourceibias.t151 CSoutput.t33 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X350 CSoutput.t59 a_n6972_8799.t114 vdd.t154 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X351 a_n6972_8799.t14 plus.t21 a_n3827_n3924.t27 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X352 vdd.t16 CSoutput.t195 output.t2 gnd.t77 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X353 vdd.t152 a_n6972_8799.t115 CSoutput.t58 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X354 gnd.t240 gnd.t237 gnd.t239 gnd.t238 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X355 CSoutput.t30 commonsourceibias.t152 gnd.t99 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X356 CSoutput.t4 commonsourceibias.t153 gnd.t13 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X357 commonsourceibias.t3 commonsourceibias.t2 gnd.t177 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X358 gnd.t236 gnd.t234 plus.t4 gnd.t235 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X359 outputibias.t5 outputibias.t4 gnd.t91 gnd.t90 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X360 diffpairibias.t3 diffpairibias.t2 gnd.t183 gnd.t182 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X361 vdd.t151 a_n6972_8799.t116 CSoutput.t57 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X362 vdd.t30 vdd.t27 vdd.t29 vdd.t28 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X363 CSoutput.t56 a_n6972_8799.t117 vdd.t149 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X364 a_n3827_n3924.t45 plus.t22 a_n6972_8799.t13 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X365 gnd.t233 gnd.t231 plus.t3 gnd.t232 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X366 vdd.t147 a_n6972_8799.t118 CSoutput.t55 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X367 outputibias.t3 outputibias.t2 gnd.t115 gnd.t114 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X368 diffpairibias.t1 diffpairibias.t0 gnd.t221 gnd.t220 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X369 a_n3827_n3924.t37 plus.t23 a_n6972_8799.t12 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X370 CSoutput.t14 commonsourceibias.t154 gnd.t54 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X371 outputibias.t1 outputibias.t0 gnd.t161 gnd.t160 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X372 vdd.t120 a_n1996_n452.t69 a_n1808_13878.t0 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X373 gnd.t97 commonsourceibias.t155 CSoutput.t29 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X374 a_n6972_8799.t11 plus.t24 a_n3827_n3924.t29 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X375 a_n3827_n3924.t17 minus.t23 a_n1996_n452.t13 gnd.t128 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X376 CSoutput.t54 a_n6972_8799.t119 vdd.t145 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X377 vdd.t143 a_n6972_8799.t120 CSoutput.t53 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X378 vdd.t141 a_n6972_8799.t121 CSoutput.t52 vdd.t140 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X379 CSoutput.t6 commonsourceibias.t156 gnd.t26 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X380 CSoutput.t51 a_n6972_8799.t122 vdd.t133 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X381 output.t1 CSoutput.t196 vdd.t17 gnd.t78 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X382 gnd.t65 commonsourceibias.t157 CSoutput.t19 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X383 gnd.t230 gnd.t227 gnd.t229 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X384 a_n1996_n452.t12 minus.t24 a_n3827_n3924.t16 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X385 CSoutput.t50 a_n6972_8799.t123 vdd.t131 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X386 gnd.t52 commonsourceibias.t158 CSoutput.t13 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X387 a_n1986_8322.t10 a_n1996_n452.t70 a_n6972_8799.t31 vdd.t105 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X388 vdd.t139 a_n6972_8799.t124 CSoutput.t49 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X389 CSoutput.t48 a_n6972_8799.t125 vdd.t137 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X390 output.t0 CSoutput.t197 vdd.t18 gnd.t79 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X391 vdd.t135 a_n6972_8799.t126 CSoutput.t47 vdd.t134 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X392 gnd.t11 commonsourceibias.t159 CSoutput.t3 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X393 a_n1986_8322.t2 a_n1996_n452.t71 vdd.t3 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X394 a_n1808_13878.t9 a_n1996_n452.t31 a_n1996_n452.t32 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X395 vdd.t129 a_n6972_8799.t127 CSoutput.t46 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X396 commonsourceibias.t1 commonsourceibias.t0 gnd.t113 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X397 a_n3827_n3924.t21 diffpairibias.t29 gnd.t136 gnd.t135 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X398 a_n1996_n452.t42 a_n1996_n452.t41 a_n1808_13878.t8 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X399 vdd.t26 vdd.t23 vdd.t25 vdd.t24 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
R0 plus.n43 plus.t18 322.512
R1 plus.n9 plus.t13 322.512
R2 plus.n42 plus.t17 297.12
R3 plus.n46 plus.t22 297.12
R4 plus.n48 plus.t21 297.12
R5 plus.n52 plus.t23 297.12
R6 plus.n54 plus.t8 297.12
R7 plus.n58 plus.t7 297.12
R8 plus.n60 plus.t12 297.12
R9 plus.n64 plus.t10 297.12
R10 plus.n66 plus.t24 297.12
R11 plus.n32 plus.t14 297.12
R12 plus.n30 plus.t15 297.12
R13 plus.n2 plus.t9 297.12
R14 plus.n24 plus.t5 297.12
R15 plus.n4 plus.t6 297.12
R16 plus.n18 plus.t19 297.12
R17 plus.n6 plus.t20 297.12
R18 plus.n12 plus.t16 297.12
R19 plus.n8 plus.t11 297.12
R20 plus.n70 plus.t3 243.97
R21 plus.n70 plus.n69 223.454
R22 plus.n72 plus.n71 223.454
R23 plus.n67 plus.n66 161.3
R24 plus.n65 plus.n34 161.3
R25 plus.n64 plus.n63 161.3
R26 plus.n62 plus.n35 161.3
R27 plus.n61 plus.n60 161.3
R28 plus.n59 plus.n36 161.3
R29 plus.n58 plus.n57 161.3
R30 plus.n56 plus.n37 161.3
R31 plus.n55 plus.n54 161.3
R32 plus.n53 plus.n38 161.3
R33 plus.n52 plus.n51 161.3
R34 plus.n50 plus.n39 161.3
R35 plus.n49 plus.n48 161.3
R36 plus.n47 plus.n40 161.3
R37 plus.n46 plus.n45 161.3
R38 plus.n44 plus.n41 161.3
R39 plus.n11 plus.n10 161.3
R40 plus.n12 plus.n7 161.3
R41 plus.n14 plus.n13 161.3
R42 plus.n15 plus.n6 161.3
R43 plus.n17 plus.n16 161.3
R44 plus.n18 plus.n5 161.3
R45 plus.n20 plus.n19 161.3
R46 plus.n21 plus.n4 161.3
R47 plus.n23 plus.n22 161.3
R48 plus.n24 plus.n3 161.3
R49 plus.n26 plus.n25 161.3
R50 plus.n27 plus.n2 161.3
R51 plus.n29 plus.n28 161.3
R52 plus.n30 plus.n1 161.3
R53 plus.n31 plus.n0 161.3
R54 plus.n33 plus.n32 161.3
R55 plus.n44 plus.n43 45.0031
R56 plus.n10 plus.n9 45.0031
R57 plus.n66 plus.n65 41.6278
R58 plus.n32 plus.n31 41.6278
R59 plus.n42 plus.n41 37.246
R60 plus.n64 plus.n35 37.246
R61 plus.n30 plus.n29 37.246
R62 plus.n11 plus.n8 37.246
R63 plus.n47 plus.n46 32.8641
R64 plus.n60 plus.n59 32.8641
R65 plus.n25 plus.n2 32.8641
R66 plus.n13 plus.n12 32.8641
R67 plus.n68 plus.n67 31.6047
R68 plus.n48 plus.n39 28.4823
R69 plus.n58 plus.n37 28.4823
R70 plus.n24 plus.n23 28.4823
R71 plus.n17 plus.n6 28.4823
R72 plus.n53 plus.n52 24.1005
R73 plus.n54 plus.n53 24.1005
R74 plus.n19 plus.n4 24.1005
R75 plus.n19 plus.n18 24.1005
R76 plus.n69 plus.t1 19.8005
R77 plus.n69 plus.t2 19.8005
R78 plus.n71 plus.t4 19.8005
R79 plus.n71 plus.t0 19.8005
R80 plus.n52 plus.n39 19.7187
R81 plus.n54 plus.n37 19.7187
R82 plus.n23 plus.n4 19.7187
R83 plus.n18 plus.n17 19.7187
R84 plus.n43 plus.n42 15.6319
R85 plus.n9 plus.n8 15.6319
R86 plus.n48 plus.n47 15.3369
R87 plus.n59 plus.n58 15.3369
R88 plus.n25 plus.n24 15.3369
R89 plus.n13 plus.n6 15.3369
R90 plus plus.n73 15.0665
R91 plus.n68 plus.n33 11.866
R92 plus.n46 plus.n41 10.955
R93 plus.n60 plus.n35 10.955
R94 plus.n29 plus.n2 10.955
R95 plus.n12 plus.n11 10.955
R96 plus.n65 plus.n64 6.57323
R97 plus.n31 plus.n30 6.57323
R98 plus.n73 plus.n72 5.40567
R99 plus.n73 plus.n68 1.188
R100 plus.n72 plus.n70 0.716017
R101 plus.n45 plus.n44 0.189894
R102 plus.n45 plus.n40 0.189894
R103 plus.n49 plus.n40 0.189894
R104 plus.n50 plus.n49 0.189894
R105 plus.n51 plus.n50 0.189894
R106 plus.n51 plus.n38 0.189894
R107 plus.n55 plus.n38 0.189894
R108 plus.n56 plus.n55 0.189894
R109 plus.n57 plus.n56 0.189894
R110 plus.n57 plus.n36 0.189894
R111 plus.n61 plus.n36 0.189894
R112 plus.n62 plus.n61 0.189894
R113 plus.n63 plus.n62 0.189894
R114 plus.n63 plus.n34 0.189894
R115 plus.n67 plus.n34 0.189894
R116 plus.n33 plus.n0 0.189894
R117 plus.n1 plus.n0 0.189894
R118 plus.n28 plus.n1 0.189894
R119 plus.n28 plus.n27 0.189894
R120 plus.n27 plus.n26 0.189894
R121 plus.n26 plus.n3 0.189894
R122 plus.n22 plus.n3 0.189894
R123 plus.n22 plus.n21 0.189894
R124 plus.n21 plus.n20 0.189894
R125 plus.n20 plus.n5 0.189894
R126 plus.n16 plus.n5 0.189894
R127 plus.n16 plus.n15 0.189894
R128 plus.n15 plus.n14 0.189894
R129 plus.n14 plus.n7 0.189894
R130 plus.n10 plus.n7 0.189894
R131 a_n3827_n3924.n10 a_n3827_n3924.t13 214.994
R132 a_n3827_n3924.n7 a_n3827_n3924.t20 214.994
R133 a_n3827_n3924.n10 a_n3827_n3924.t48 214.321
R134 a_n3827_n3924.n10 a_n3827_n3924.t15 214.321
R135 a_n3827_n3924.n9 a_n3827_n3924.t7 214.321
R136 a_n3827_n3924.n9 a_n3827_n3924.t21 214.321
R137 a_n3827_n3924.n8 a_n3827_n3924.t47 214.321
R138 a_n3827_n3924.n8 a_n3827_n3924.t25 214.321
R139 a_n3827_n3924.n7 a_n3827_n3924.t10 214.321
R140 a_n3827_n3924.n7 a_n3827_n3924.t49 214.321
R141 a_n3827_n3924.n4 a_n3827_n3924.t40 55.8337
R142 a_n3827_n3924.n4 a_n3827_n3924.t16 55.8337
R143 a_n3827_n3924.n6 a_n3827_n3924.t46 55.8337
R144 a_n3827_n3924.n3 a_n3827_n3924.t29 55.8335
R145 a_n3827_n3924.n11 a_n3827_n3924.t4 55.8335
R146 a_n3827_n3924.n0 a_n3827_n3924.t22 55.8335
R147 a_n3827_n3924.n0 a_n3827_n3924.t30 55.8335
R148 a_n3827_n3924.n2 a_n3827_n3924.t31 55.8335
R149 a_n3827_n3924.n29 a_n3827_n3924.n11 53.0054
R150 a_n3827_n3924.n3 a_n3827_n3924.n13 53.0052
R151 a_n3827_n3924.n4 a_n3827_n3924.n14 53.0052
R152 a_n3827_n3924.n4 a_n3827_n3924.n15 53.0052
R153 a_n3827_n3924.n4 a_n3827_n3924.n16 53.0052
R154 a_n3827_n3924.n5 a_n3827_n3924.n17 53.0052
R155 a_n3827_n3924.n5 a_n3827_n3924.n18 53.0052
R156 a_n3827_n3924.n6 a_n3827_n3924.n19 53.0052
R157 a_n3827_n3924.n6 a_n3827_n3924.n20 53.0052
R158 a_n3827_n3924.n0 a_n3827_n3924.n12 53.0051
R159 a_n3827_n3924.n0 a_n3827_n3924.n21 53.0051
R160 a_n3827_n3924.n0 a_n3827_n3924.n22 53.0051
R161 a_n3827_n3924.n1 a_n3827_n3924.n23 53.0051
R162 a_n3827_n3924.n1 a_n3827_n3924.n24 53.0051
R163 a_n3827_n3924.n2 a_n3827_n3924.n25 53.0051
R164 a_n3827_n3924.n2 a_n3827_n3924.n26 53.0051
R165 a_n3827_n3924.n27 a_n3827_n3924.n6 12.1986
R166 a_n3827_n3924.n28 a_n3827_n3924.n3 12.1986
R167 a_n3827_n3924.n27 a_n3827_n3924.n2 5.11903
R168 a_n3827_n3924.n11 a_n3827_n3924.n28 5.11903
R169 a_n3827_n3924.n12 a_n3827_n3924.t19 2.82907
R170 a_n3827_n3924.n12 a_n3827_n3924.t11 2.82907
R171 a_n3827_n3924.n21 a_n3827_n3924.t5 2.82907
R172 a_n3827_n3924.n21 a_n3827_n3924.t24 2.82907
R173 a_n3827_n3924.n22 a_n3827_n3924.t6 2.82907
R174 a_n3827_n3924.n22 a_n3827_n3924.t9 2.82907
R175 a_n3827_n3924.n23 a_n3827_n3924.t36 2.82907
R176 a_n3827_n3924.n23 a_n3827_n3924.t32 2.82907
R177 a_n3827_n3924.n24 a_n3827_n3924.t35 2.82907
R178 a_n3827_n3924.n24 a_n3827_n3924.t44 2.82907
R179 a_n3827_n3924.n25 a_n3827_n3924.t33 2.82907
R180 a_n3827_n3924.n25 a_n3827_n3924.t26 2.82907
R181 a_n3827_n3924.n26 a_n3827_n3924.t34 2.82907
R182 a_n3827_n3924.n26 a_n3827_n3924.t43 2.82907
R183 a_n3827_n3924.n13 a_n3827_n3924.t39 2.82907
R184 a_n3827_n3924.n13 a_n3827_n3924.t28 2.82907
R185 a_n3827_n3924.n14 a_n3827_n3924.t42 2.82907
R186 a_n3827_n3924.n14 a_n3827_n3924.t41 2.82907
R187 a_n3827_n3924.n15 a_n3827_n3924.t27 2.82907
R188 a_n3827_n3924.n15 a_n3827_n3924.t37 2.82907
R189 a_n3827_n3924.n16 a_n3827_n3924.t38 2.82907
R190 a_n3827_n3924.n16 a_n3827_n3924.t45 2.82907
R191 a_n3827_n3924.n17 a_n3827_n3924.t2 2.82907
R192 a_n3827_n3924.n17 a_n3827_n3924.t17 2.82907
R193 a_n3827_n3924.n18 a_n3827_n3924.t23 2.82907
R194 a_n3827_n3924.n18 a_n3827_n3924.t12 2.82907
R195 a_n3827_n3924.n19 a_n3827_n3924.t14 2.82907
R196 a_n3827_n3924.n19 a_n3827_n3924.t1 2.82907
R197 a_n3827_n3924.n20 a_n3827_n3924.t8 2.82907
R198 a_n3827_n3924.n20 a_n3827_n3924.t18 2.82907
R199 a_n3827_n3924.t0 a_n3827_n3924.n29 2.82907
R200 a_n3827_n3924.n29 a_n3827_n3924.t3 2.82907
R201 a_n3827_n3924.n8 a_n3827_n3924.n7 2.01503
R202 a_n3827_n3924.n7 a_n3827_n3924.n27 1.95694
R203 a_n3827_n3924.n28 a_n3827_n3924.n10 1.95694
R204 a_n3827_n3924.n6 a_n3827_n3924.n5 1.77636
R205 a_n3827_n3924.n4 a_n3827_n3924.n3 1.77636
R206 a_n3827_n3924.n2 a_n3827_n3924.n1 1.77636
R207 a_n3827_n3924.n11 a_n3827_n3924.n0 1.77636
R208 a_n3827_n3924.n9 a_n3827_n3924.n8 1.34352
R209 a_n3827_n3924.n10 a_n3827_n3924.n9 1.34352
R210 a_n3827_n3924.n1 a_n3827_n3924.n0 1.12334
R211 a_n3827_n3924.n5 a_n3827_n3924.n4 1.12334
R212 a_n6972_8799.n172 a_n6972_8799.t54 485.149
R213 a_n6972_8799.n220 a_n6972_8799.t66 485.149
R214 a_n6972_8799.n269 a_n6972_8799.t114 485.149
R215 a_n6972_8799.n24 a_n6972_8799.t110 485.149
R216 a_n6972_8799.n72 a_n6972_8799.t121 485.149
R217 a_n6972_8799.n121 a_n6972_8799.t113 485.149
R218 a_n6972_8799.n204 a_n6972_8799.t75 464.166
R219 a_n6972_8799.n203 a_n6972_8799.t74 464.166
R220 a_n6972_8799.n159 a_n6972_8799.t52 464.166
R221 a_n6972_8799.n197 a_n6972_8799.t111 464.166
R222 a_n6972_8799.n196 a_n6972_8799.t76 464.166
R223 a_n6972_8799.n162 a_n6972_8799.t58 464.166
R224 a_n6972_8799.n190 a_n6972_8799.t115 464.166
R225 a_n6972_8799.n189 a_n6972_8799.t90 464.166
R226 a_n6972_8799.n165 a_n6972_8799.t88 464.166
R227 a_n6972_8799.n184 a_n6972_8799.t35 464.166
R228 a_n6972_8799.n182 a_n6972_8799.t94 464.166
R229 a_n6972_8799.n168 a_n6972_8799.t93 464.166
R230 a_n6972_8799.n177 a_n6972_8799.t37 464.166
R231 a_n6972_8799.n175 a_n6972_8799.t36 464.166
R232 a_n6972_8799.n171 a_n6972_8799.t107 464.166
R233 a_n6972_8799.n252 a_n6972_8799.t82 464.166
R234 a_n6972_8799.n251 a_n6972_8799.t81 464.166
R235 a_n6972_8799.n207 a_n6972_8799.t65 464.166
R236 a_n6972_8799.n245 a_n6972_8799.t123 464.166
R237 a_n6972_8799.n244 a_n6972_8799.t87 464.166
R238 a_n6972_8799.n210 a_n6972_8799.t67 464.166
R239 a_n6972_8799.n238 a_n6972_8799.t127 464.166
R240 a_n6972_8799.n237 a_n6972_8799.t100 464.166
R241 a_n6972_8799.n213 a_n6972_8799.t99 464.166
R242 a_n6972_8799.n232 a_n6972_8799.t44 464.166
R243 a_n6972_8799.n230 a_n6972_8799.t103 464.166
R244 a_n6972_8799.n216 a_n6972_8799.t102 464.166
R245 a_n6972_8799.n225 a_n6972_8799.t48 464.166
R246 a_n6972_8799.n223 a_n6972_8799.t47 464.166
R247 a_n6972_8799.n219 a_n6972_8799.t118 464.166
R248 a_n6972_8799.n301 a_n6972_8799.t126 464.166
R249 a_n6972_8799.n300 a_n6972_8799.t46 464.166
R250 a_n6972_8799.n256 a_n6972_8799.t86 464.166
R251 a_n6972_8799.n294 a_n6972_8799.t34 464.166
R252 a_n6972_8799.n293 a_n6972_8799.t106 464.166
R253 a_n6972_8799.n259 a_n6972_8799.t56 464.166
R254 a_n6972_8799.n287 a_n6972_8799.t92 464.166
R255 a_n6972_8799.n286 a_n6972_8799.t39 464.166
R256 a_n6972_8799.n262 a_n6972_8799.t60 464.166
R257 a_n6972_8799.n281 a_n6972_8799.t122 464.166
R258 a_n6972_8799.n279 a_n6972_8799.t98 464.166
R259 a_n6972_8799.n265 a_n6972_8799.t117 464.166
R260 a_n6972_8799.n274 a_n6972_8799.t84 464.166
R261 a_n6972_8799.n272 a_n6972_8799.t101 464.166
R262 a_n6972_8799.n268 a_n6972_8799.t50 464.166
R263 a_n6972_8799.n23 a_n6972_8799.t72 464.166
R264 a_n6972_8799.n27 a_n6972_8799.t73 464.166
R265 a_n6972_8799.n21 a_n6972_8799.t96 464.166
R266 a_n6972_8799.n32 a_n6972_8799.t63 464.166
R267 a_n6972_8799.n34 a_n6972_8799.t64 464.166
R268 a_n6972_8799.n38 a_n6972_8799.t95 464.166
R269 a_n6972_8799.n39 a_n6972_8799.t32 464.166
R270 a_n6972_8799.n17 a_n6972_8799.t61 464.166
R271 a_n6972_8799.n44 a_n6972_8799.t78 464.166
R272 a_n6972_8799.n46 a_n6972_8799.t112 464.166
R273 a_n6972_8799.n50 a_n6972_8799.t43 464.166
R274 a_n6972_8799.n51 a_n6972_8799.t59 464.166
R275 a_n6972_8799.n13 a_n6972_8799.t109 464.166
R276 a_n6972_8799.n57 a_n6972_8799.t40 464.166
R277 a_n6972_8799.n58 a_n6972_8799.t41 464.166
R278 a_n6972_8799.n71 a_n6972_8799.t79 464.166
R279 a_n6972_8799.n75 a_n6972_8799.t80 464.166
R280 a_n6972_8799.n69 a_n6972_8799.t108 464.166
R281 a_n6972_8799.n80 a_n6972_8799.t70 464.166
R282 a_n6972_8799.n82 a_n6972_8799.t71 464.166
R283 a_n6972_8799.n86 a_n6972_8799.t104 464.166
R284 a_n6972_8799.n87 a_n6972_8799.t42 464.166
R285 a_n6972_8799.n65 a_n6972_8799.t69 464.166
R286 a_n6972_8799.n92 a_n6972_8799.t89 464.166
R287 a_n6972_8799.n94 a_n6972_8799.t124 464.166
R288 a_n6972_8799.n98 a_n6972_8799.t57 464.166
R289 a_n6972_8799.n99 a_n6972_8799.t68 464.166
R290 a_n6972_8799.n61 a_n6972_8799.t119 464.166
R291 a_n6972_8799.n105 a_n6972_8799.t51 464.166
R292 a_n6972_8799.n106 a_n6972_8799.t53 464.166
R293 a_n6972_8799.n120 a_n6972_8799.t49 464.166
R294 a_n6972_8799.n124 a_n6972_8799.t33 464.166
R295 a_n6972_8799.n118 a_n6972_8799.t83 464.166
R296 a_n6972_8799.n129 a_n6972_8799.t116 464.166
R297 a_n6972_8799.n131 a_n6972_8799.t97 464.166
R298 a_n6972_8799.n135 a_n6972_8799.t120 464.166
R299 a_n6972_8799.n136 a_n6972_8799.t77 464.166
R300 a_n6972_8799.n114 a_n6972_8799.t38 464.166
R301 a_n6972_8799.n141 a_n6972_8799.t91 464.166
R302 a_n6972_8799.n143 a_n6972_8799.t55 464.166
R303 a_n6972_8799.n147 a_n6972_8799.t105 464.166
R304 a_n6972_8799.n148 a_n6972_8799.t62 464.166
R305 a_n6972_8799.n110 a_n6972_8799.t85 464.166
R306 a_n6972_8799.n154 a_n6972_8799.t45 464.166
R307 a_n6972_8799.n155 a_n6972_8799.t125 464.166
R308 a_n6972_8799.n174 a_n6972_8799.n173 161.3
R309 a_n6972_8799.n175 a_n6972_8799.n170 161.3
R310 a_n6972_8799.n176 a_n6972_8799.n169 161.3
R311 a_n6972_8799.n178 a_n6972_8799.n177 161.3
R312 a_n6972_8799.n179 a_n6972_8799.n168 161.3
R313 a_n6972_8799.n181 a_n6972_8799.n180 161.3
R314 a_n6972_8799.n182 a_n6972_8799.n167 161.3
R315 a_n6972_8799.n183 a_n6972_8799.n166 161.3
R316 a_n6972_8799.n185 a_n6972_8799.n184 161.3
R317 a_n6972_8799.n186 a_n6972_8799.n165 161.3
R318 a_n6972_8799.n188 a_n6972_8799.n187 161.3
R319 a_n6972_8799.n189 a_n6972_8799.n164 161.3
R320 a_n6972_8799.n190 a_n6972_8799.n163 161.3
R321 a_n6972_8799.n192 a_n6972_8799.n191 161.3
R322 a_n6972_8799.n193 a_n6972_8799.n162 161.3
R323 a_n6972_8799.n195 a_n6972_8799.n194 161.3
R324 a_n6972_8799.n196 a_n6972_8799.n161 161.3
R325 a_n6972_8799.n197 a_n6972_8799.n160 161.3
R326 a_n6972_8799.n199 a_n6972_8799.n198 161.3
R327 a_n6972_8799.n200 a_n6972_8799.n159 161.3
R328 a_n6972_8799.n202 a_n6972_8799.n201 161.3
R329 a_n6972_8799.n203 a_n6972_8799.n158 161.3
R330 a_n6972_8799.n205 a_n6972_8799.n204 161.3
R331 a_n6972_8799.n222 a_n6972_8799.n221 161.3
R332 a_n6972_8799.n223 a_n6972_8799.n218 161.3
R333 a_n6972_8799.n224 a_n6972_8799.n217 161.3
R334 a_n6972_8799.n226 a_n6972_8799.n225 161.3
R335 a_n6972_8799.n227 a_n6972_8799.n216 161.3
R336 a_n6972_8799.n229 a_n6972_8799.n228 161.3
R337 a_n6972_8799.n230 a_n6972_8799.n215 161.3
R338 a_n6972_8799.n231 a_n6972_8799.n214 161.3
R339 a_n6972_8799.n233 a_n6972_8799.n232 161.3
R340 a_n6972_8799.n234 a_n6972_8799.n213 161.3
R341 a_n6972_8799.n236 a_n6972_8799.n235 161.3
R342 a_n6972_8799.n237 a_n6972_8799.n212 161.3
R343 a_n6972_8799.n238 a_n6972_8799.n211 161.3
R344 a_n6972_8799.n240 a_n6972_8799.n239 161.3
R345 a_n6972_8799.n241 a_n6972_8799.n210 161.3
R346 a_n6972_8799.n243 a_n6972_8799.n242 161.3
R347 a_n6972_8799.n244 a_n6972_8799.n209 161.3
R348 a_n6972_8799.n245 a_n6972_8799.n208 161.3
R349 a_n6972_8799.n247 a_n6972_8799.n246 161.3
R350 a_n6972_8799.n248 a_n6972_8799.n207 161.3
R351 a_n6972_8799.n250 a_n6972_8799.n249 161.3
R352 a_n6972_8799.n251 a_n6972_8799.n206 161.3
R353 a_n6972_8799.n253 a_n6972_8799.n252 161.3
R354 a_n6972_8799.n271 a_n6972_8799.n270 161.3
R355 a_n6972_8799.n272 a_n6972_8799.n267 161.3
R356 a_n6972_8799.n273 a_n6972_8799.n266 161.3
R357 a_n6972_8799.n275 a_n6972_8799.n274 161.3
R358 a_n6972_8799.n276 a_n6972_8799.n265 161.3
R359 a_n6972_8799.n278 a_n6972_8799.n277 161.3
R360 a_n6972_8799.n279 a_n6972_8799.n264 161.3
R361 a_n6972_8799.n280 a_n6972_8799.n263 161.3
R362 a_n6972_8799.n282 a_n6972_8799.n281 161.3
R363 a_n6972_8799.n283 a_n6972_8799.n262 161.3
R364 a_n6972_8799.n285 a_n6972_8799.n284 161.3
R365 a_n6972_8799.n286 a_n6972_8799.n261 161.3
R366 a_n6972_8799.n287 a_n6972_8799.n260 161.3
R367 a_n6972_8799.n289 a_n6972_8799.n288 161.3
R368 a_n6972_8799.n290 a_n6972_8799.n259 161.3
R369 a_n6972_8799.n292 a_n6972_8799.n291 161.3
R370 a_n6972_8799.n293 a_n6972_8799.n258 161.3
R371 a_n6972_8799.n294 a_n6972_8799.n257 161.3
R372 a_n6972_8799.n296 a_n6972_8799.n295 161.3
R373 a_n6972_8799.n297 a_n6972_8799.n256 161.3
R374 a_n6972_8799.n299 a_n6972_8799.n298 161.3
R375 a_n6972_8799.n300 a_n6972_8799.n255 161.3
R376 a_n6972_8799.n302 a_n6972_8799.n301 161.3
R377 a_n6972_8799.n59 a_n6972_8799.n58 161.3
R378 a_n6972_8799.n57 a_n6972_8799.n12 161.3
R379 a_n6972_8799.n56 a_n6972_8799.n55 161.3
R380 a_n6972_8799.n54 a_n6972_8799.n13 161.3
R381 a_n6972_8799.n53 a_n6972_8799.n52 161.3
R382 a_n6972_8799.n51 a_n6972_8799.n14 161.3
R383 a_n6972_8799.n50 a_n6972_8799.n49 161.3
R384 a_n6972_8799.n48 a_n6972_8799.n15 161.3
R385 a_n6972_8799.n47 a_n6972_8799.n46 161.3
R386 a_n6972_8799.n45 a_n6972_8799.n16 161.3
R387 a_n6972_8799.n44 a_n6972_8799.n43 161.3
R388 a_n6972_8799.n42 a_n6972_8799.n17 161.3
R389 a_n6972_8799.n41 a_n6972_8799.n40 161.3
R390 a_n6972_8799.n39 a_n6972_8799.n18 161.3
R391 a_n6972_8799.n38 a_n6972_8799.n37 161.3
R392 a_n6972_8799.n36 a_n6972_8799.n19 161.3
R393 a_n6972_8799.n35 a_n6972_8799.n34 161.3
R394 a_n6972_8799.n33 a_n6972_8799.n20 161.3
R395 a_n6972_8799.n32 a_n6972_8799.n31 161.3
R396 a_n6972_8799.n30 a_n6972_8799.n21 161.3
R397 a_n6972_8799.n29 a_n6972_8799.n28 161.3
R398 a_n6972_8799.n27 a_n6972_8799.n22 161.3
R399 a_n6972_8799.n26 a_n6972_8799.n25 161.3
R400 a_n6972_8799.n107 a_n6972_8799.n106 161.3
R401 a_n6972_8799.n105 a_n6972_8799.n60 161.3
R402 a_n6972_8799.n104 a_n6972_8799.n103 161.3
R403 a_n6972_8799.n102 a_n6972_8799.n61 161.3
R404 a_n6972_8799.n101 a_n6972_8799.n100 161.3
R405 a_n6972_8799.n99 a_n6972_8799.n62 161.3
R406 a_n6972_8799.n98 a_n6972_8799.n97 161.3
R407 a_n6972_8799.n96 a_n6972_8799.n63 161.3
R408 a_n6972_8799.n95 a_n6972_8799.n94 161.3
R409 a_n6972_8799.n93 a_n6972_8799.n64 161.3
R410 a_n6972_8799.n92 a_n6972_8799.n91 161.3
R411 a_n6972_8799.n90 a_n6972_8799.n65 161.3
R412 a_n6972_8799.n89 a_n6972_8799.n88 161.3
R413 a_n6972_8799.n87 a_n6972_8799.n66 161.3
R414 a_n6972_8799.n86 a_n6972_8799.n85 161.3
R415 a_n6972_8799.n84 a_n6972_8799.n67 161.3
R416 a_n6972_8799.n83 a_n6972_8799.n82 161.3
R417 a_n6972_8799.n81 a_n6972_8799.n68 161.3
R418 a_n6972_8799.n80 a_n6972_8799.n79 161.3
R419 a_n6972_8799.n78 a_n6972_8799.n69 161.3
R420 a_n6972_8799.n77 a_n6972_8799.n76 161.3
R421 a_n6972_8799.n75 a_n6972_8799.n70 161.3
R422 a_n6972_8799.n74 a_n6972_8799.n73 161.3
R423 a_n6972_8799.n156 a_n6972_8799.n155 161.3
R424 a_n6972_8799.n154 a_n6972_8799.n109 161.3
R425 a_n6972_8799.n153 a_n6972_8799.n152 161.3
R426 a_n6972_8799.n151 a_n6972_8799.n110 161.3
R427 a_n6972_8799.n150 a_n6972_8799.n149 161.3
R428 a_n6972_8799.n148 a_n6972_8799.n111 161.3
R429 a_n6972_8799.n147 a_n6972_8799.n146 161.3
R430 a_n6972_8799.n145 a_n6972_8799.n112 161.3
R431 a_n6972_8799.n144 a_n6972_8799.n143 161.3
R432 a_n6972_8799.n142 a_n6972_8799.n113 161.3
R433 a_n6972_8799.n141 a_n6972_8799.n140 161.3
R434 a_n6972_8799.n139 a_n6972_8799.n114 161.3
R435 a_n6972_8799.n138 a_n6972_8799.n137 161.3
R436 a_n6972_8799.n136 a_n6972_8799.n115 161.3
R437 a_n6972_8799.n135 a_n6972_8799.n134 161.3
R438 a_n6972_8799.n133 a_n6972_8799.n116 161.3
R439 a_n6972_8799.n132 a_n6972_8799.n131 161.3
R440 a_n6972_8799.n130 a_n6972_8799.n117 161.3
R441 a_n6972_8799.n129 a_n6972_8799.n128 161.3
R442 a_n6972_8799.n127 a_n6972_8799.n118 161.3
R443 a_n6972_8799.n126 a_n6972_8799.n125 161.3
R444 a_n6972_8799.n124 a_n6972_8799.n119 161.3
R445 a_n6972_8799.n123 a_n6972_8799.n122 161.3
R446 a_n6972_8799.n8 a_n6972_8799.n6 98.9633
R447 a_n6972_8799.n3 a_n6972_8799.n1 98.9631
R448 a_n6972_8799.n10 a_n6972_8799.n9 98.6055
R449 a_n6972_8799.n8 a_n6972_8799.n7 98.6055
R450 a_n6972_8799.n3 a_n6972_8799.n2 98.6055
R451 a_n6972_8799.n5 a_n6972_8799.n4 98.6055
R452 a_n6972_8799.n308 a_n6972_8799.n306 81.3764
R453 a_n6972_8799.n317 a_n6972_8799.n315 81.3764
R454 a_n6972_8799.n320 a_n6972_8799.n0 81.3764
R455 a_n6972_8799.n321 a_n6972_8799.n320 80.9326
R456 a_n6972_8799.n314 a_n6972_8799.n313 80.9324
R457 a_n6972_8799.n312 a_n6972_8799.n311 80.9324
R458 a_n6972_8799.n310 a_n6972_8799.n309 80.9324
R459 a_n6972_8799.n308 a_n6972_8799.n307 80.9324
R460 a_n6972_8799.n317 a_n6972_8799.n316 80.9324
R461 a_n6972_8799.n319 a_n6972_8799.n318 80.9324
R462 a_n6972_8799.n173 a_n6972_8799.n172 70.4033
R463 a_n6972_8799.n221 a_n6972_8799.n220 70.4033
R464 a_n6972_8799.n270 a_n6972_8799.n269 70.4033
R465 a_n6972_8799.n25 a_n6972_8799.n24 70.4033
R466 a_n6972_8799.n73 a_n6972_8799.n72 70.4033
R467 a_n6972_8799.n122 a_n6972_8799.n121 70.4033
R468 a_n6972_8799.n204 a_n6972_8799.n203 48.2005
R469 a_n6972_8799.n197 a_n6972_8799.n196 48.2005
R470 a_n6972_8799.n190 a_n6972_8799.n189 48.2005
R471 a_n6972_8799.n184 a_n6972_8799.n165 48.2005
R472 a_n6972_8799.n177 a_n6972_8799.n168 48.2005
R473 a_n6972_8799.n252 a_n6972_8799.n251 48.2005
R474 a_n6972_8799.n245 a_n6972_8799.n244 48.2005
R475 a_n6972_8799.n238 a_n6972_8799.n237 48.2005
R476 a_n6972_8799.n232 a_n6972_8799.n213 48.2005
R477 a_n6972_8799.n225 a_n6972_8799.n216 48.2005
R478 a_n6972_8799.n301 a_n6972_8799.n300 48.2005
R479 a_n6972_8799.n294 a_n6972_8799.n293 48.2005
R480 a_n6972_8799.n287 a_n6972_8799.n286 48.2005
R481 a_n6972_8799.n281 a_n6972_8799.n262 48.2005
R482 a_n6972_8799.n274 a_n6972_8799.n265 48.2005
R483 a_n6972_8799.n32 a_n6972_8799.n21 48.2005
R484 a_n6972_8799.n39 a_n6972_8799.n38 48.2005
R485 a_n6972_8799.n44 a_n6972_8799.n17 48.2005
R486 a_n6972_8799.n51 a_n6972_8799.n50 48.2005
R487 a_n6972_8799.n58 a_n6972_8799.n57 48.2005
R488 a_n6972_8799.n80 a_n6972_8799.n69 48.2005
R489 a_n6972_8799.n87 a_n6972_8799.n86 48.2005
R490 a_n6972_8799.n92 a_n6972_8799.n65 48.2005
R491 a_n6972_8799.n99 a_n6972_8799.n98 48.2005
R492 a_n6972_8799.n106 a_n6972_8799.n105 48.2005
R493 a_n6972_8799.n129 a_n6972_8799.n118 48.2005
R494 a_n6972_8799.n136 a_n6972_8799.n135 48.2005
R495 a_n6972_8799.n141 a_n6972_8799.n114 48.2005
R496 a_n6972_8799.n148 a_n6972_8799.n147 48.2005
R497 a_n6972_8799.n155 a_n6972_8799.n154 48.2005
R498 a_n6972_8799.n191 a_n6972_8799.n162 47.4702
R499 a_n6972_8799.n183 a_n6972_8799.n182 47.4702
R500 a_n6972_8799.n239 a_n6972_8799.n210 47.4702
R501 a_n6972_8799.n231 a_n6972_8799.n230 47.4702
R502 a_n6972_8799.n288 a_n6972_8799.n259 47.4702
R503 a_n6972_8799.n280 a_n6972_8799.n279 47.4702
R504 a_n6972_8799.n34 a_n6972_8799.n19 47.4702
R505 a_n6972_8799.n46 a_n6972_8799.n45 47.4702
R506 a_n6972_8799.n82 a_n6972_8799.n67 47.4702
R507 a_n6972_8799.n94 a_n6972_8799.n93 47.4702
R508 a_n6972_8799.n131 a_n6972_8799.n116 47.4702
R509 a_n6972_8799.n143 a_n6972_8799.n142 47.4702
R510 a_n6972_8799.n198 a_n6972_8799.n159 46.0096
R511 a_n6972_8799.n176 a_n6972_8799.n175 46.0096
R512 a_n6972_8799.n246 a_n6972_8799.n207 46.0096
R513 a_n6972_8799.n224 a_n6972_8799.n223 46.0096
R514 a_n6972_8799.n295 a_n6972_8799.n256 46.0096
R515 a_n6972_8799.n273 a_n6972_8799.n272 46.0096
R516 a_n6972_8799.n28 a_n6972_8799.n27 46.0096
R517 a_n6972_8799.n52 a_n6972_8799.n13 46.0096
R518 a_n6972_8799.n76 a_n6972_8799.n75 46.0096
R519 a_n6972_8799.n100 a_n6972_8799.n61 46.0096
R520 a_n6972_8799.n125 a_n6972_8799.n124 46.0096
R521 a_n6972_8799.n149 a_n6972_8799.n110 46.0096
R522 a_n6972_8799.n319 a_n6972_8799.n314 32.7526
R523 a_n6972_8799.n11 a_n6972_8799.n5 30.7135
R524 a_n6972_8799.n202 a_n6972_8799.n159 27.0217
R525 a_n6972_8799.n175 a_n6972_8799.n174 27.0217
R526 a_n6972_8799.n250 a_n6972_8799.n207 27.0217
R527 a_n6972_8799.n223 a_n6972_8799.n222 27.0217
R528 a_n6972_8799.n299 a_n6972_8799.n256 27.0217
R529 a_n6972_8799.n272 a_n6972_8799.n271 27.0217
R530 a_n6972_8799.n27 a_n6972_8799.n26 27.0217
R531 a_n6972_8799.n56 a_n6972_8799.n13 27.0217
R532 a_n6972_8799.n75 a_n6972_8799.n74 27.0217
R533 a_n6972_8799.n104 a_n6972_8799.n61 27.0217
R534 a_n6972_8799.n124 a_n6972_8799.n123 27.0217
R535 a_n6972_8799.n153 a_n6972_8799.n110 27.0217
R536 a_n6972_8799.n195 a_n6972_8799.n162 25.5611
R537 a_n6972_8799.n182 a_n6972_8799.n181 25.5611
R538 a_n6972_8799.n243 a_n6972_8799.n210 25.5611
R539 a_n6972_8799.n230 a_n6972_8799.n229 25.5611
R540 a_n6972_8799.n292 a_n6972_8799.n259 25.5611
R541 a_n6972_8799.n279 a_n6972_8799.n278 25.5611
R542 a_n6972_8799.n34 a_n6972_8799.n33 25.5611
R543 a_n6972_8799.n46 a_n6972_8799.n15 25.5611
R544 a_n6972_8799.n82 a_n6972_8799.n81 25.5611
R545 a_n6972_8799.n94 a_n6972_8799.n63 25.5611
R546 a_n6972_8799.n131 a_n6972_8799.n130 25.5611
R547 a_n6972_8799.n143 a_n6972_8799.n112 25.5611
R548 a_n6972_8799.n189 a_n6972_8799.n188 24.1005
R549 a_n6972_8799.n188 a_n6972_8799.n165 24.1005
R550 a_n6972_8799.n237 a_n6972_8799.n236 24.1005
R551 a_n6972_8799.n236 a_n6972_8799.n213 24.1005
R552 a_n6972_8799.n286 a_n6972_8799.n285 24.1005
R553 a_n6972_8799.n285 a_n6972_8799.n262 24.1005
R554 a_n6972_8799.n40 a_n6972_8799.n39 24.1005
R555 a_n6972_8799.n40 a_n6972_8799.n17 24.1005
R556 a_n6972_8799.n88 a_n6972_8799.n87 24.1005
R557 a_n6972_8799.n88 a_n6972_8799.n65 24.1005
R558 a_n6972_8799.n137 a_n6972_8799.n136 24.1005
R559 a_n6972_8799.n137 a_n6972_8799.n114 24.1005
R560 a_n6972_8799.n196 a_n6972_8799.n195 22.6399
R561 a_n6972_8799.n181 a_n6972_8799.n168 22.6399
R562 a_n6972_8799.n244 a_n6972_8799.n243 22.6399
R563 a_n6972_8799.n229 a_n6972_8799.n216 22.6399
R564 a_n6972_8799.n293 a_n6972_8799.n292 22.6399
R565 a_n6972_8799.n278 a_n6972_8799.n265 22.6399
R566 a_n6972_8799.n33 a_n6972_8799.n32 22.6399
R567 a_n6972_8799.n50 a_n6972_8799.n15 22.6399
R568 a_n6972_8799.n81 a_n6972_8799.n80 22.6399
R569 a_n6972_8799.n98 a_n6972_8799.n63 22.6399
R570 a_n6972_8799.n130 a_n6972_8799.n129 22.6399
R571 a_n6972_8799.n147 a_n6972_8799.n112 22.6399
R572 a_n6972_8799.n203 a_n6972_8799.n202 21.1793
R573 a_n6972_8799.n174 a_n6972_8799.n171 21.1793
R574 a_n6972_8799.n251 a_n6972_8799.n250 21.1793
R575 a_n6972_8799.n222 a_n6972_8799.n219 21.1793
R576 a_n6972_8799.n300 a_n6972_8799.n299 21.1793
R577 a_n6972_8799.n271 a_n6972_8799.n268 21.1793
R578 a_n6972_8799.n26 a_n6972_8799.n23 21.1793
R579 a_n6972_8799.n57 a_n6972_8799.n56 21.1793
R580 a_n6972_8799.n74 a_n6972_8799.n71 21.1793
R581 a_n6972_8799.n105 a_n6972_8799.n104 21.1793
R582 a_n6972_8799.n123 a_n6972_8799.n120 21.1793
R583 a_n6972_8799.n154 a_n6972_8799.n153 21.1793
R584 a_n6972_8799.n172 a_n6972_8799.n171 20.9576
R585 a_n6972_8799.n220 a_n6972_8799.n219 20.9576
R586 a_n6972_8799.n269 a_n6972_8799.n268 20.9576
R587 a_n6972_8799.n24 a_n6972_8799.n23 20.9576
R588 a_n6972_8799.n72 a_n6972_8799.n71 20.9576
R589 a_n6972_8799.n121 a_n6972_8799.n120 20.9576
R590 a_n6972_8799.n11 a_n6972_8799.n10 17.7361
R591 a_n6972_8799.n310 a_n6972_8799.n305 12.3339
R592 a_n6972_8799.n305 a_n6972_8799.n11 11.4887
R593 a_n6972_8799.n254 a_n6972_8799.n205 9.07815
R594 a_n6972_8799.n108 a_n6972_8799.n59 9.07815
R595 a_n6972_8799.n304 a_n6972_8799.n157 6.86985
R596 a_n6972_8799.n304 a_n6972_8799.n303 6.51296
R597 a_n6972_8799.n254 a_n6972_8799.n253 4.9702
R598 a_n6972_8799.n303 a_n6972_8799.n302 4.9702
R599 a_n6972_8799.n108 a_n6972_8799.n107 4.9702
R600 a_n6972_8799.n157 a_n6972_8799.n156 4.9702
R601 a_n6972_8799.n303 a_n6972_8799.n254 4.10845
R602 a_n6972_8799.n157 a_n6972_8799.n108 4.10845
R603 a_n6972_8799.n9 a_n6972_8799.t7 3.61217
R604 a_n6972_8799.n9 a_n6972_8799.t10 3.61217
R605 a_n6972_8799.n7 a_n6972_8799.t9 3.61217
R606 a_n6972_8799.n7 a_n6972_8799.t5 3.61217
R607 a_n6972_8799.n6 a_n6972_8799.t31 3.61217
R608 a_n6972_8799.n6 a_n6972_8799.t2 3.61217
R609 a_n6972_8799.n1 a_n6972_8799.t1 3.61217
R610 a_n6972_8799.n1 a_n6972_8799.t3 3.61217
R611 a_n6972_8799.n2 a_n6972_8799.t4 3.61217
R612 a_n6972_8799.n2 a_n6972_8799.t6 3.61217
R613 a_n6972_8799.n4 a_n6972_8799.t0 3.61217
R614 a_n6972_8799.n4 a_n6972_8799.t8 3.61217
R615 a_n6972_8799.n305 a_n6972_8799.n304 3.4105
R616 a_n6972_8799.n315 a_n6972_8799.t24 2.82907
R617 a_n6972_8799.n315 a_n6972_8799.t22 2.82907
R618 a_n6972_8799.n316 a_n6972_8799.t15 2.82907
R619 a_n6972_8799.n316 a_n6972_8799.t19 2.82907
R620 a_n6972_8799.n318 a_n6972_8799.t29 2.82907
R621 a_n6972_8799.n318 a_n6972_8799.t16 2.82907
R622 a_n6972_8799.n313 a_n6972_8799.t25 2.82907
R623 a_n6972_8799.n313 a_n6972_8799.t11 2.82907
R624 a_n6972_8799.n311 a_n6972_8799.t28 2.82907
R625 a_n6972_8799.n311 a_n6972_8799.t23 2.82907
R626 a_n6972_8799.n309 a_n6972_8799.t12 2.82907
R627 a_n6972_8799.n309 a_n6972_8799.t27 2.82907
R628 a_n6972_8799.n307 a_n6972_8799.t13 2.82907
R629 a_n6972_8799.n307 a_n6972_8799.t14 2.82907
R630 a_n6972_8799.n306 a_n6972_8799.t17 2.82907
R631 a_n6972_8799.n306 a_n6972_8799.t18 2.82907
R632 a_n6972_8799.n0 a_n6972_8799.t21 2.82907
R633 a_n6972_8799.n0 a_n6972_8799.t20 2.82907
R634 a_n6972_8799.n321 a_n6972_8799.t26 2.82907
R635 a_n6972_8799.t30 a_n6972_8799.n321 2.82907
R636 a_n6972_8799.n198 a_n6972_8799.n197 2.19141
R637 a_n6972_8799.n177 a_n6972_8799.n176 2.19141
R638 a_n6972_8799.n246 a_n6972_8799.n245 2.19141
R639 a_n6972_8799.n225 a_n6972_8799.n224 2.19141
R640 a_n6972_8799.n295 a_n6972_8799.n294 2.19141
R641 a_n6972_8799.n274 a_n6972_8799.n273 2.19141
R642 a_n6972_8799.n28 a_n6972_8799.n21 2.19141
R643 a_n6972_8799.n52 a_n6972_8799.n51 2.19141
R644 a_n6972_8799.n76 a_n6972_8799.n69 2.19141
R645 a_n6972_8799.n100 a_n6972_8799.n99 2.19141
R646 a_n6972_8799.n125 a_n6972_8799.n118 2.19141
R647 a_n6972_8799.n149 a_n6972_8799.n148 2.19141
R648 a_n6972_8799.n191 a_n6972_8799.n190 0.730803
R649 a_n6972_8799.n184 a_n6972_8799.n183 0.730803
R650 a_n6972_8799.n239 a_n6972_8799.n238 0.730803
R651 a_n6972_8799.n232 a_n6972_8799.n231 0.730803
R652 a_n6972_8799.n288 a_n6972_8799.n287 0.730803
R653 a_n6972_8799.n281 a_n6972_8799.n280 0.730803
R654 a_n6972_8799.n38 a_n6972_8799.n19 0.730803
R655 a_n6972_8799.n45 a_n6972_8799.n44 0.730803
R656 a_n6972_8799.n86 a_n6972_8799.n67 0.730803
R657 a_n6972_8799.n93 a_n6972_8799.n92 0.730803
R658 a_n6972_8799.n135 a_n6972_8799.n116 0.730803
R659 a_n6972_8799.n142 a_n6972_8799.n141 0.730803
R660 a_n6972_8799.n310 a_n6972_8799.n308 0.444466
R661 a_n6972_8799.n312 a_n6972_8799.n310 0.444466
R662 a_n6972_8799.n314 a_n6972_8799.n312 0.444466
R663 a_n6972_8799.n320 a_n6972_8799.n319 0.444466
R664 a_n6972_8799.n319 a_n6972_8799.n317 0.444466
R665 a_n6972_8799.n10 a_n6972_8799.n8 0.358259
R666 a_n6972_8799.n5 a_n6972_8799.n3 0.358259
R667 a_n6972_8799.n205 a_n6972_8799.n158 0.189894
R668 a_n6972_8799.n201 a_n6972_8799.n158 0.189894
R669 a_n6972_8799.n201 a_n6972_8799.n200 0.189894
R670 a_n6972_8799.n200 a_n6972_8799.n199 0.189894
R671 a_n6972_8799.n199 a_n6972_8799.n160 0.189894
R672 a_n6972_8799.n161 a_n6972_8799.n160 0.189894
R673 a_n6972_8799.n194 a_n6972_8799.n161 0.189894
R674 a_n6972_8799.n194 a_n6972_8799.n193 0.189894
R675 a_n6972_8799.n193 a_n6972_8799.n192 0.189894
R676 a_n6972_8799.n192 a_n6972_8799.n163 0.189894
R677 a_n6972_8799.n164 a_n6972_8799.n163 0.189894
R678 a_n6972_8799.n187 a_n6972_8799.n164 0.189894
R679 a_n6972_8799.n187 a_n6972_8799.n186 0.189894
R680 a_n6972_8799.n186 a_n6972_8799.n185 0.189894
R681 a_n6972_8799.n185 a_n6972_8799.n166 0.189894
R682 a_n6972_8799.n167 a_n6972_8799.n166 0.189894
R683 a_n6972_8799.n180 a_n6972_8799.n167 0.189894
R684 a_n6972_8799.n180 a_n6972_8799.n179 0.189894
R685 a_n6972_8799.n179 a_n6972_8799.n178 0.189894
R686 a_n6972_8799.n178 a_n6972_8799.n169 0.189894
R687 a_n6972_8799.n170 a_n6972_8799.n169 0.189894
R688 a_n6972_8799.n173 a_n6972_8799.n170 0.189894
R689 a_n6972_8799.n253 a_n6972_8799.n206 0.189894
R690 a_n6972_8799.n249 a_n6972_8799.n206 0.189894
R691 a_n6972_8799.n249 a_n6972_8799.n248 0.189894
R692 a_n6972_8799.n248 a_n6972_8799.n247 0.189894
R693 a_n6972_8799.n247 a_n6972_8799.n208 0.189894
R694 a_n6972_8799.n209 a_n6972_8799.n208 0.189894
R695 a_n6972_8799.n242 a_n6972_8799.n209 0.189894
R696 a_n6972_8799.n242 a_n6972_8799.n241 0.189894
R697 a_n6972_8799.n241 a_n6972_8799.n240 0.189894
R698 a_n6972_8799.n240 a_n6972_8799.n211 0.189894
R699 a_n6972_8799.n212 a_n6972_8799.n211 0.189894
R700 a_n6972_8799.n235 a_n6972_8799.n212 0.189894
R701 a_n6972_8799.n235 a_n6972_8799.n234 0.189894
R702 a_n6972_8799.n234 a_n6972_8799.n233 0.189894
R703 a_n6972_8799.n233 a_n6972_8799.n214 0.189894
R704 a_n6972_8799.n215 a_n6972_8799.n214 0.189894
R705 a_n6972_8799.n228 a_n6972_8799.n215 0.189894
R706 a_n6972_8799.n228 a_n6972_8799.n227 0.189894
R707 a_n6972_8799.n227 a_n6972_8799.n226 0.189894
R708 a_n6972_8799.n226 a_n6972_8799.n217 0.189894
R709 a_n6972_8799.n218 a_n6972_8799.n217 0.189894
R710 a_n6972_8799.n221 a_n6972_8799.n218 0.189894
R711 a_n6972_8799.n302 a_n6972_8799.n255 0.189894
R712 a_n6972_8799.n298 a_n6972_8799.n255 0.189894
R713 a_n6972_8799.n298 a_n6972_8799.n297 0.189894
R714 a_n6972_8799.n297 a_n6972_8799.n296 0.189894
R715 a_n6972_8799.n296 a_n6972_8799.n257 0.189894
R716 a_n6972_8799.n258 a_n6972_8799.n257 0.189894
R717 a_n6972_8799.n291 a_n6972_8799.n258 0.189894
R718 a_n6972_8799.n291 a_n6972_8799.n290 0.189894
R719 a_n6972_8799.n290 a_n6972_8799.n289 0.189894
R720 a_n6972_8799.n289 a_n6972_8799.n260 0.189894
R721 a_n6972_8799.n261 a_n6972_8799.n260 0.189894
R722 a_n6972_8799.n284 a_n6972_8799.n261 0.189894
R723 a_n6972_8799.n284 a_n6972_8799.n283 0.189894
R724 a_n6972_8799.n283 a_n6972_8799.n282 0.189894
R725 a_n6972_8799.n282 a_n6972_8799.n263 0.189894
R726 a_n6972_8799.n264 a_n6972_8799.n263 0.189894
R727 a_n6972_8799.n277 a_n6972_8799.n264 0.189894
R728 a_n6972_8799.n277 a_n6972_8799.n276 0.189894
R729 a_n6972_8799.n276 a_n6972_8799.n275 0.189894
R730 a_n6972_8799.n275 a_n6972_8799.n266 0.189894
R731 a_n6972_8799.n267 a_n6972_8799.n266 0.189894
R732 a_n6972_8799.n270 a_n6972_8799.n267 0.189894
R733 a_n6972_8799.n25 a_n6972_8799.n22 0.189894
R734 a_n6972_8799.n29 a_n6972_8799.n22 0.189894
R735 a_n6972_8799.n30 a_n6972_8799.n29 0.189894
R736 a_n6972_8799.n31 a_n6972_8799.n30 0.189894
R737 a_n6972_8799.n31 a_n6972_8799.n20 0.189894
R738 a_n6972_8799.n35 a_n6972_8799.n20 0.189894
R739 a_n6972_8799.n36 a_n6972_8799.n35 0.189894
R740 a_n6972_8799.n37 a_n6972_8799.n36 0.189894
R741 a_n6972_8799.n37 a_n6972_8799.n18 0.189894
R742 a_n6972_8799.n41 a_n6972_8799.n18 0.189894
R743 a_n6972_8799.n42 a_n6972_8799.n41 0.189894
R744 a_n6972_8799.n43 a_n6972_8799.n42 0.189894
R745 a_n6972_8799.n43 a_n6972_8799.n16 0.189894
R746 a_n6972_8799.n47 a_n6972_8799.n16 0.189894
R747 a_n6972_8799.n48 a_n6972_8799.n47 0.189894
R748 a_n6972_8799.n49 a_n6972_8799.n48 0.189894
R749 a_n6972_8799.n49 a_n6972_8799.n14 0.189894
R750 a_n6972_8799.n53 a_n6972_8799.n14 0.189894
R751 a_n6972_8799.n54 a_n6972_8799.n53 0.189894
R752 a_n6972_8799.n55 a_n6972_8799.n54 0.189894
R753 a_n6972_8799.n55 a_n6972_8799.n12 0.189894
R754 a_n6972_8799.n59 a_n6972_8799.n12 0.189894
R755 a_n6972_8799.n73 a_n6972_8799.n70 0.189894
R756 a_n6972_8799.n77 a_n6972_8799.n70 0.189894
R757 a_n6972_8799.n78 a_n6972_8799.n77 0.189894
R758 a_n6972_8799.n79 a_n6972_8799.n78 0.189894
R759 a_n6972_8799.n79 a_n6972_8799.n68 0.189894
R760 a_n6972_8799.n83 a_n6972_8799.n68 0.189894
R761 a_n6972_8799.n84 a_n6972_8799.n83 0.189894
R762 a_n6972_8799.n85 a_n6972_8799.n84 0.189894
R763 a_n6972_8799.n85 a_n6972_8799.n66 0.189894
R764 a_n6972_8799.n89 a_n6972_8799.n66 0.189894
R765 a_n6972_8799.n90 a_n6972_8799.n89 0.189894
R766 a_n6972_8799.n91 a_n6972_8799.n90 0.189894
R767 a_n6972_8799.n91 a_n6972_8799.n64 0.189894
R768 a_n6972_8799.n95 a_n6972_8799.n64 0.189894
R769 a_n6972_8799.n96 a_n6972_8799.n95 0.189894
R770 a_n6972_8799.n97 a_n6972_8799.n96 0.189894
R771 a_n6972_8799.n97 a_n6972_8799.n62 0.189894
R772 a_n6972_8799.n101 a_n6972_8799.n62 0.189894
R773 a_n6972_8799.n102 a_n6972_8799.n101 0.189894
R774 a_n6972_8799.n103 a_n6972_8799.n102 0.189894
R775 a_n6972_8799.n103 a_n6972_8799.n60 0.189894
R776 a_n6972_8799.n107 a_n6972_8799.n60 0.189894
R777 a_n6972_8799.n122 a_n6972_8799.n119 0.189894
R778 a_n6972_8799.n126 a_n6972_8799.n119 0.189894
R779 a_n6972_8799.n127 a_n6972_8799.n126 0.189894
R780 a_n6972_8799.n128 a_n6972_8799.n127 0.189894
R781 a_n6972_8799.n128 a_n6972_8799.n117 0.189894
R782 a_n6972_8799.n132 a_n6972_8799.n117 0.189894
R783 a_n6972_8799.n133 a_n6972_8799.n132 0.189894
R784 a_n6972_8799.n134 a_n6972_8799.n133 0.189894
R785 a_n6972_8799.n134 a_n6972_8799.n115 0.189894
R786 a_n6972_8799.n138 a_n6972_8799.n115 0.189894
R787 a_n6972_8799.n139 a_n6972_8799.n138 0.189894
R788 a_n6972_8799.n140 a_n6972_8799.n139 0.189894
R789 a_n6972_8799.n140 a_n6972_8799.n113 0.189894
R790 a_n6972_8799.n144 a_n6972_8799.n113 0.189894
R791 a_n6972_8799.n145 a_n6972_8799.n144 0.189894
R792 a_n6972_8799.n146 a_n6972_8799.n145 0.189894
R793 a_n6972_8799.n146 a_n6972_8799.n111 0.189894
R794 a_n6972_8799.n150 a_n6972_8799.n111 0.189894
R795 a_n6972_8799.n151 a_n6972_8799.n150 0.189894
R796 a_n6972_8799.n152 a_n6972_8799.n151 0.189894
R797 a_n6972_8799.n152 a_n6972_8799.n109 0.189894
R798 a_n6972_8799.n156 a_n6972_8799.n109 0.189894
R799 gnd.n6708 gnd.n746 838.101
R800 gnd.n3538 gnd.n2158 766.379
R801 gnd.n3541 gnd.n3540 766.379
R802 gnd.n2780 gnd.n2683 766.379
R803 gnd.n2776 gnd.n2681 766.379
R804 gnd.n3629 gnd.n2180 756.769
R805 gnd.n3532 gnd.n3531 756.769
R806 gnd.n2873 gnd.n2590 756.769
R807 gnd.n2871 gnd.n2593 756.769
R808 gnd.n7473 gnd.n129 751.963
R809 gnd.n7631 gnd.n7630 751.963
R810 gnd.n7179 gnd.n457 751.963
R811 gnd.n7232 gnd.n459 751.963
R812 gnd.n6256 gnd.n1087 751.963
R813 gnd.n4723 gnd.n1090 751.963
R814 gnd.n4061 gnd.n3633 751.963
R815 gnd.n4102 gnd.n3635 751.963
R816 gnd.n7628 gnd.n131 732.745
R817 gnd.n199 gnd.n127 732.745
R818 gnd.n7105 gnd.n456 732.745
R819 gnd.n7234 gnd.n454 732.745
R820 gnd.n6254 gnd.n1092 732.745
R821 gnd.n6185 gnd.n1089 732.745
R822 gnd.n3867 gnd.n3632 732.745
R823 gnd.n4104 gnd.n2156 732.745
R824 gnd.n4531 gnd.n978 723.135
R825 gnd.n6707 gnd.n747 723.135
R826 gnd.n6921 gnd.n6919 723.135
R827 gnd.n4535 gnd.n980 723.135
R828 gnd.n4769 gnd.n1897 711.122
R829 gnd.n6000 gnd.n464 711.122
R830 gnd.n4648 gnd.n1188 711.122
R831 gnd.n6002 gnd.n1314 711.122
R832 gnd.n6316 gnd.n980 587.962
R833 gnd.n4268 gnd.n4267 585
R834 gnd.n4267 gnd.n979 585
R835 gnd.n4269 gnd.n1990 585
R836 gnd.n4282 gnd.n1990 585
R837 gnd.n4270 gnd.n2001 585
R838 gnd.n2001 gnd.n1999 585
R839 gnd.n4272 gnd.n4271 585
R840 gnd.n4273 gnd.n4272 585
R841 gnd.n2002 gnd.n2000 585
R842 gnd.n2000 gnd.n1996 585
R843 gnd.n4257 gnd.n4256 585
R844 gnd.n4256 gnd.n4255 585
R845 gnd.n2005 gnd.n2004 585
R846 gnd.n2006 gnd.n2005 585
R847 gnd.n4246 gnd.n4245 585
R848 gnd.n4247 gnd.n4246 585
R849 gnd.n2017 gnd.n2016 585
R850 gnd.n2023 gnd.n2016 585
R851 gnd.n4241 gnd.n4240 585
R852 gnd.n4240 gnd.n4239 585
R853 gnd.n2020 gnd.n2019 585
R854 gnd.n2032 gnd.n2020 585
R855 gnd.n4230 gnd.n4229 585
R856 gnd.n4231 gnd.n4230 585
R857 gnd.n2034 gnd.n2033 585
R858 gnd.n2033 gnd.n2029 585
R859 gnd.n4225 gnd.n4224 585
R860 gnd.n4224 gnd.n4223 585
R861 gnd.n2038 gnd.n2037 585
R862 gnd.n2039 gnd.n2038 585
R863 gnd.n4214 gnd.n4213 585
R864 gnd.n4215 gnd.n4214 585
R865 gnd.n2051 gnd.n2050 585
R866 gnd.n2050 gnd.n2047 585
R867 gnd.n4209 gnd.n4208 585
R868 gnd.n4208 gnd.n4207 585
R869 gnd.n2054 gnd.n2053 585
R870 gnd.n2065 gnd.n2054 585
R871 gnd.n4198 gnd.n4197 585
R872 gnd.n4199 gnd.n4198 585
R873 gnd.n2067 gnd.n2066 585
R874 gnd.n2066 gnd.n2062 585
R875 gnd.n4193 gnd.n4192 585
R876 gnd.n4192 gnd.n4191 585
R877 gnd.n2070 gnd.n2069 585
R878 gnd.n2071 gnd.n2070 585
R879 gnd.n4182 gnd.n4181 585
R880 gnd.n4183 gnd.n4182 585
R881 gnd.n2083 gnd.n2082 585
R882 gnd.n2082 gnd.n2079 585
R883 gnd.n4177 gnd.n4176 585
R884 gnd.n4176 gnd.n4175 585
R885 gnd.n2086 gnd.n2085 585
R886 gnd.n2097 gnd.n2086 585
R887 gnd.n4166 gnd.n4165 585
R888 gnd.n4167 gnd.n4166 585
R889 gnd.n2099 gnd.n2098 585
R890 gnd.n2098 gnd.n2094 585
R891 gnd.n4161 gnd.n4160 585
R892 gnd.n4160 gnd.n4159 585
R893 gnd.n2102 gnd.n2101 585
R894 gnd.n2103 gnd.n2102 585
R895 gnd.n4150 gnd.n4149 585
R896 gnd.n4151 gnd.n4150 585
R897 gnd.n2115 gnd.n2114 585
R898 gnd.n2114 gnd.n2111 585
R899 gnd.n4145 gnd.n4144 585
R900 gnd.n4144 gnd.n4143 585
R901 gnd.n2118 gnd.n2117 585
R902 gnd.n2129 gnd.n2118 585
R903 gnd.n4134 gnd.n4133 585
R904 gnd.n4135 gnd.n4134 585
R905 gnd.n2131 gnd.n2130 585
R906 gnd.n2130 gnd.n2126 585
R907 gnd.n4129 gnd.n4128 585
R908 gnd.n4128 gnd.n4127 585
R909 gnd.n2134 gnd.n2133 585
R910 gnd.n2135 gnd.n2134 585
R911 gnd.n4118 gnd.n4117 585
R912 gnd.n4119 gnd.n4118 585
R913 gnd.n2147 gnd.n2146 585
R914 gnd.n2146 gnd.n2143 585
R915 gnd.n4113 gnd.n4112 585
R916 gnd.n4112 gnd.n4111 585
R917 gnd.n2150 gnd.n2149 585
R918 gnd.n3634 gnd.n2150 585
R919 gnd.n4102 gnd.n4101 585
R920 gnd.n4103 gnd.n4102 585
R921 gnd.n4098 gnd.n3635 585
R922 gnd.n4097 gnd.n4096 585
R923 gnd.n4094 gnd.n3637 585
R924 gnd.n4092 gnd.n4091 585
R925 gnd.n4090 gnd.n3638 585
R926 gnd.n4089 gnd.n4088 585
R927 gnd.n4086 gnd.n3643 585
R928 gnd.n4084 gnd.n4083 585
R929 gnd.n4082 gnd.n3644 585
R930 gnd.n4081 gnd.n4080 585
R931 gnd.n4078 gnd.n3649 585
R932 gnd.n4076 gnd.n4075 585
R933 gnd.n4074 gnd.n3650 585
R934 gnd.n4073 gnd.n4072 585
R935 gnd.n4070 gnd.n3655 585
R936 gnd.n4068 gnd.n4067 585
R937 gnd.n4066 gnd.n3656 585
R938 gnd.n4060 gnd.n3661 585
R939 gnd.n4062 gnd.n4061 585
R940 gnd.n4061 gnd.n3631 585
R941 gnd.n3992 gnd.n3704 585
R942 gnd.n3704 gnd.n979 585
R943 gnd.n3993 gnd.n1989 585
R944 gnd.n4282 gnd.n1989 585
R945 gnd.n3702 gnd.n3701 585
R946 gnd.n3701 gnd.n1999 585
R947 gnd.n3997 gnd.n1998 585
R948 gnd.n4273 gnd.n1998 585
R949 gnd.n3998 gnd.n3700 585
R950 gnd.n3700 gnd.n1996 585
R951 gnd.n3999 gnd.n2008 585
R952 gnd.n4255 gnd.n2008 585
R953 gnd.n3698 gnd.n3697 585
R954 gnd.n3697 gnd.n2006 585
R955 gnd.n4003 gnd.n2015 585
R956 gnd.n4247 gnd.n2015 585
R957 gnd.n4004 gnd.n3696 585
R958 gnd.n3696 gnd.n2023 585
R959 gnd.n4005 gnd.n2022 585
R960 gnd.n4239 gnd.n2022 585
R961 gnd.n3694 gnd.n3693 585
R962 gnd.n3693 gnd.n2032 585
R963 gnd.n4009 gnd.n2031 585
R964 gnd.n4231 gnd.n2031 585
R965 gnd.n4011 gnd.n4010 585
R966 gnd.n4010 gnd.n2029 585
R967 gnd.n4012 gnd.n2041 585
R968 gnd.n4223 gnd.n2041 585
R969 gnd.n4014 gnd.n4013 585
R970 gnd.n4013 gnd.n2039 585
R971 gnd.n4015 gnd.n2049 585
R972 gnd.n4215 gnd.n2049 585
R973 gnd.n4017 gnd.n4016 585
R974 gnd.n4016 gnd.n2047 585
R975 gnd.n4018 gnd.n2056 585
R976 gnd.n4207 gnd.n2056 585
R977 gnd.n4020 gnd.n4019 585
R978 gnd.n4019 gnd.n2065 585
R979 gnd.n4021 gnd.n2064 585
R980 gnd.n4199 gnd.n2064 585
R981 gnd.n4023 gnd.n4022 585
R982 gnd.n4022 gnd.n2062 585
R983 gnd.n4024 gnd.n2073 585
R984 gnd.n4191 gnd.n2073 585
R985 gnd.n4026 gnd.n4025 585
R986 gnd.n4025 gnd.n2071 585
R987 gnd.n4027 gnd.n2081 585
R988 gnd.n4183 gnd.n2081 585
R989 gnd.n4029 gnd.n4028 585
R990 gnd.n4028 gnd.n2079 585
R991 gnd.n4030 gnd.n2088 585
R992 gnd.n4175 gnd.n2088 585
R993 gnd.n4032 gnd.n4031 585
R994 gnd.n4031 gnd.n2097 585
R995 gnd.n4033 gnd.n2096 585
R996 gnd.n4167 gnd.n2096 585
R997 gnd.n4035 gnd.n4034 585
R998 gnd.n4034 gnd.n2094 585
R999 gnd.n4036 gnd.n2105 585
R1000 gnd.n4159 gnd.n2105 585
R1001 gnd.n4038 gnd.n4037 585
R1002 gnd.n4037 gnd.n2103 585
R1003 gnd.n4039 gnd.n2113 585
R1004 gnd.n4151 gnd.n2113 585
R1005 gnd.n4041 gnd.n4040 585
R1006 gnd.n4040 gnd.n2111 585
R1007 gnd.n4042 gnd.n2120 585
R1008 gnd.n4143 gnd.n2120 585
R1009 gnd.n4044 gnd.n4043 585
R1010 gnd.n4043 gnd.n2129 585
R1011 gnd.n4045 gnd.n2128 585
R1012 gnd.n4135 gnd.n2128 585
R1013 gnd.n4047 gnd.n4046 585
R1014 gnd.n4046 gnd.n2126 585
R1015 gnd.n4048 gnd.n2137 585
R1016 gnd.n4127 gnd.n2137 585
R1017 gnd.n4050 gnd.n4049 585
R1018 gnd.n4049 gnd.n2135 585
R1019 gnd.n4051 gnd.n2145 585
R1020 gnd.n4119 gnd.n2145 585
R1021 gnd.n4053 gnd.n4052 585
R1022 gnd.n4052 gnd.n2143 585
R1023 gnd.n4054 gnd.n2152 585
R1024 gnd.n4111 gnd.n2152 585
R1025 gnd.n4056 gnd.n4055 585
R1026 gnd.n4055 gnd.n3634 585
R1027 gnd.n4057 gnd.n3633 585
R1028 gnd.n4103 gnd.n3633 585
R1029 gnd.n3538 gnd.n3537 585
R1030 gnd.n3539 gnd.n3538 585
R1031 gnd.n2233 gnd.n2232 585
R1032 gnd.n2239 gnd.n2232 585
R1033 gnd.n3513 gnd.n2251 585
R1034 gnd.n2251 gnd.n2238 585
R1035 gnd.n3515 gnd.n3514 585
R1036 gnd.n3516 gnd.n3515 585
R1037 gnd.n2252 gnd.n2250 585
R1038 gnd.n2250 gnd.n2246 585
R1039 gnd.n3247 gnd.n3246 585
R1040 gnd.n3246 gnd.n3245 585
R1041 gnd.n2257 gnd.n2256 585
R1042 gnd.n3216 gnd.n2257 585
R1043 gnd.n3236 gnd.n3235 585
R1044 gnd.n3235 gnd.n3234 585
R1045 gnd.n2264 gnd.n2263 585
R1046 gnd.n3222 gnd.n2264 585
R1047 gnd.n3192 gnd.n2284 585
R1048 gnd.n2284 gnd.n2283 585
R1049 gnd.n3194 gnd.n3193 585
R1050 gnd.n3195 gnd.n3194 585
R1051 gnd.n2285 gnd.n2282 585
R1052 gnd.n2293 gnd.n2282 585
R1053 gnd.n3170 gnd.n2305 585
R1054 gnd.n2305 gnd.n2292 585
R1055 gnd.n3172 gnd.n3171 585
R1056 gnd.n3173 gnd.n3172 585
R1057 gnd.n2306 gnd.n2304 585
R1058 gnd.n2304 gnd.n2300 585
R1059 gnd.n3158 gnd.n3157 585
R1060 gnd.n3157 gnd.n3156 585
R1061 gnd.n2311 gnd.n2310 585
R1062 gnd.n2321 gnd.n2311 585
R1063 gnd.n3147 gnd.n3146 585
R1064 gnd.n3146 gnd.n3145 585
R1065 gnd.n2318 gnd.n2317 585
R1066 gnd.n3133 gnd.n2318 585
R1067 gnd.n3107 gnd.n2339 585
R1068 gnd.n2339 gnd.n2328 585
R1069 gnd.n3109 gnd.n3108 585
R1070 gnd.n3110 gnd.n3109 585
R1071 gnd.n2340 gnd.n2338 585
R1072 gnd.n2348 gnd.n2338 585
R1073 gnd.n3085 gnd.n2360 585
R1074 gnd.n2360 gnd.n2347 585
R1075 gnd.n3087 gnd.n3086 585
R1076 gnd.n3088 gnd.n3087 585
R1077 gnd.n2361 gnd.n2359 585
R1078 gnd.n2359 gnd.n2355 585
R1079 gnd.n3073 gnd.n3072 585
R1080 gnd.n3072 gnd.n3071 585
R1081 gnd.n2366 gnd.n2365 585
R1082 gnd.n2375 gnd.n2366 585
R1083 gnd.n3062 gnd.n3061 585
R1084 gnd.n3061 gnd.n3060 585
R1085 gnd.n2373 gnd.n2372 585
R1086 gnd.n3048 gnd.n2373 585
R1087 gnd.n2486 gnd.n2485 585
R1088 gnd.n2486 gnd.n2382 585
R1089 gnd.n3005 gnd.n3004 585
R1090 gnd.n3004 gnd.n3003 585
R1091 gnd.n3006 gnd.n2480 585
R1092 gnd.n2491 gnd.n2480 585
R1093 gnd.n3008 gnd.n3007 585
R1094 gnd.n3009 gnd.n3008 585
R1095 gnd.n2481 gnd.n2479 585
R1096 gnd.n2504 gnd.n2479 585
R1097 gnd.n2464 gnd.n2463 585
R1098 gnd.n2467 gnd.n2464 585
R1099 gnd.n3019 gnd.n3018 585
R1100 gnd.n3018 gnd.n3017 585
R1101 gnd.n3020 gnd.n2458 585
R1102 gnd.n2979 gnd.n2458 585
R1103 gnd.n3022 gnd.n3021 585
R1104 gnd.n3023 gnd.n3022 585
R1105 gnd.n2459 gnd.n2457 585
R1106 gnd.n2518 gnd.n2457 585
R1107 gnd.n2971 gnd.n2970 585
R1108 gnd.n2970 gnd.n2969 585
R1109 gnd.n2515 gnd.n2514 585
R1110 gnd.n2953 gnd.n2515 585
R1111 gnd.n2940 gnd.n2534 585
R1112 gnd.n2534 gnd.n2533 585
R1113 gnd.n2942 gnd.n2941 585
R1114 gnd.n2943 gnd.n2942 585
R1115 gnd.n2535 gnd.n2532 585
R1116 gnd.n2541 gnd.n2532 585
R1117 gnd.n2921 gnd.n2920 585
R1118 gnd.n2922 gnd.n2921 585
R1119 gnd.n2552 gnd.n2551 585
R1120 gnd.n2551 gnd.n2547 585
R1121 gnd.n2911 gnd.n2910 585
R1122 gnd.n2912 gnd.n2911 585
R1123 gnd.n2562 gnd.n2561 585
R1124 gnd.n2567 gnd.n2561 585
R1125 gnd.n2889 gnd.n2580 585
R1126 gnd.n2580 gnd.n2566 585
R1127 gnd.n2891 gnd.n2890 585
R1128 gnd.n2892 gnd.n2891 585
R1129 gnd.n2581 gnd.n2579 585
R1130 gnd.n2579 gnd.n2575 585
R1131 gnd.n2880 gnd.n2879 585
R1132 gnd.n2881 gnd.n2880 585
R1133 gnd.n2588 gnd.n2587 585
R1134 gnd.n2592 gnd.n2587 585
R1135 gnd.n2857 gnd.n2609 585
R1136 gnd.n2609 gnd.n2591 585
R1137 gnd.n2859 gnd.n2858 585
R1138 gnd.n2860 gnd.n2859 585
R1139 gnd.n2610 gnd.n2608 585
R1140 gnd.n2608 gnd.n2599 585
R1141 gnd.n2852 gnd.n2851 585
R1142 gnd.n2851 gnd.n2850 585
R1143 gnd.n2657 gnd.n2656 585
R1144 gnd.n2658 gnd.n2657 585
R1145 gnd.n2811 gnd.n2810 585
R1146 gnd.n2812 gnd.n2811 585
R1147 gnd.n2667 gnd.n2666 585
R1148 gnd.n2666 gnd.n2665 585
R1149 gnd.n2806 gnd.n2805 585
R1150 gnd.n2805 gnd.n2804 585
R1151 gnd.n2670 gnd.n2669 585
R1152 gnd.n2671 gnd.n2670 585
R1153 gnd.n2795 gnd.n2794 585
R1154 gnd.n2796 gnd.n2795 585
R1155 gnd.n2678 gnd.n2677 585
R1156 gnd.n2787 gnd.n2677 585
R1157 gnd.n2790 gnd.n2789 585
R1158 gnd.n2789 gnd.n2788 585
R1159 gnd.n2681 gnd.n2680 585
R1160 gnd.n2682 gnd.n2681 585
R1161 gnd.n2776 gnd.n2775 585
R1162 gnd.n2774 gnd.n2700 585
R1163 gnd.n2773 gnd.n2699 585
R1164 gnd.n2778 gnd.n2699 585
R1165 gnd.n2772 gnd.n2771 585
R1166 gnd.n2770 gnd.n2769 585
R1167 gnd.n2768 gnd.n2767 585
R1168 gnd.n2766 gnd.n2765 585
R1169 gnd.n2764 gnd.n2763 585
R1170 gnd.n2762 gnd.n2761 585
R1171 gnd.n2760 gnd.n2759 585
R1172 gnd.n2758 gnd.n2757 585
R1173 gnd.n2756 gnd.n2755 585
R1174 gnd.n2754 gnd.n2753 585
R1175 gnd.n2752 gnd.n2751 585
R1176 gnd.n2750 gnd.n2749 585
R1177 gnd.n2748 gnd.n2747 585
R1178 gnd.n2746 gnd.n2745 585
R1179 gnd.n2744 gnd.n2743 585
R1180 gnd.n2742 gnd.n2741 585
R1181 gnd.n2740 gnd.n2739 585
R1182 gnd.n2738 gnd.n2737 585
R1183 gnd.n2736 gnd.n2735 585
R1184 gnd.n2734 gnd.n2733 585
R1185 gnd.n2732 gnd.n2731 585
R1186 gnd.n2730 gnd.n2729 585
R1187 gnd.n2687 gnd.n2686 585
R1188 gnd.n2781 gnd.n2780 585
R1189 gnd.n3542 gnd.n3541 585
R1190 gnd.n3544 gnd.n3543 585
R1191 gnd.n3546 gnd.n3545 585
R1192 gnd.n3548 gnd.n3547 585
R1193 gnd.n3550 gnd.n3549 585
R1194 gnd.n3552 gnd.n3551 585
R1195 gnd.n3554 gnd.n3553 585
R1196 gnd.n3556 gnd.n3555 585
R1197 gnd.n3558 gnd.n3557 585
R1198 gnd.n3560 gnd.n3559 585
R1199 gnd.n3562 gnd.n3561 585
R1200 gnd.n3564 gnd.n3563 585
R1201 gnd.n3566 gnd.n3565 585
R1202 gnd.n3568 gnd.n3567 585
R1203 gnd.n3570 gnd.n3569 585
R1204 gnd.n3572 gnd.n3571 585
R1205 gnd.n3574 gnd.n3573 585
R1206 gnd.n3576 gnd.n3575 585
R1207 gnd.n3578 gnd.n3577 585
R1208 gnd.n3580 gnd.n3579 585
R1209 gnd.n3582 gnd.n3581 585
R1210 gnd.n3584 gnd.n3583 585
R1211 gnd.n3586 gnd.n3585 585
R1212 gnd.n3588 gnd.n3587 585
R1213 gnd.n3590 gnd.n3589 585
R1214 gnd.n3591 gnd.n2200 585
R1215 gnd.n3592 gnd.n2158 585
R1216 gnd.n3630 gnd.n2158 585
R1217 gnd.n3540 gnd.n2230 585
R1218 gnd.n3540 gnd.n3539 585
R1219 gnd.n3209 gnd.n2229 585
R1220 gnd.n2239 gnd.n2229 585
R1221 gnd.n3211 gnd.n3210 585
R1222 gnd.n3210 gnd.n2238 585
R1223 gnd.n3212 gnd.n2248 585
R1224 gnd.n3516 gnd.n2248 585
R1225 gnd.n3214 gnd.n3213 585
R1226 gnd.n3213 gnd.n2246 585
R1227 gnd.n3215 gnd.n2259 585
R1228 gnd.n3245 gnd.n2259 585
R1229 gnd.n3218 gnd.n3217 585
R1230 gnd.n3217 gnd.n3216 585
R1231 gnd.n3219 gnd.n2266 585
R1232 gnd.n3234 gnd.n2266 585
R1233 gnd.n3221 gnd.n3220 585
R1234 gnd.n3222 gnd.n3221 585
R1235 gnd.n2276 gnd.n2275 585
R1236 gnd.n2283 gnd.n2275 585
R1237 gnd.n3197 gnd.n3196 585
R1238 gnd.n3196 gnd.n3195 585
R1239 gnd.n2279 gnd.n2278 585
R1240 gnd.n2293 gnd.n2279 585
R1241 gnd.n3123 gnd.n3122 585
R1242 gnd.n3122 gnd.n2292 585
R1243 gnd.n3124 gnd.n2302 585
R1244 gnd.n3173 gnd.n2302 585
R1245 gnd.n3126 gnd.n3125 585
R1246 gnd.n3125 gnd.n2300 585
R1247 gnd.n3127 gnd.n2313 585
R1248 gnd.n3156 gnd.n2313 585
R1249 gnd.n3129 gnd.n3128 585
R1250 gnd.n3128 gnd.n2321 585
R1251 gnd.n3130 gnd.n2320 585
R1252 gnd.n3145 gnd.n2320 585
R1253 gnd.n3132 gnd.n3131 585
R1254 gnd.n3133 gnd.n3132 585
R1255 gnd.n2332 gnd.n2331 585
R1256 gnd.n2331 gnd.n2328 585
R1257 gnd.n3112 gnd.n3111 585
R1258 gnd.n3111 gnd.n3110 585
R1259 gnd.n2335 gnd.n2334 585
R1260 gnd.n2348 gnd.n2335 585
R1261 gnd.n3036 gnd.n3035 585
R1262 gnd.n3035 gnd.n2347 585
R1263 gnd.n3037 gnd.n2357 585
R1264 gnd.n3088 gnd.n2357 585
R1265 gnd.n3039 gnd.n3038 585
R1266 gnd.n3038 gnd.n2355 585
R1267 gnd.n3040 gnd.n2368 585
R1268 gnd.n3071 gnd.n2368 585
R1269 gnd.n3042 gnd.n3041 585
R1270 gnd.n3041 gnd.n2375 585
R1271 gnd.n3043 gnd.n2374 585
R1272 gnd.n3060 gnd.n2374 585
R1273 gnd.n3045 gnd.n3044 585
R1274 gnd.n3048 gnd.n3045 585
R1275 gnd.n2385 gnd.n2384 585
R1276 gnd.n2384 gnd.n2382 585
R1277 gnd.n2488 gnd.n2487 585
R1278 gnd.n3003 gnd.n2487 585
R1279 gnd.n2490 gnd.n2489 585
R1280 gnd.n2491 gnd.n2490 585
R1281 gnd.n2501 gnd.n2477 585
R1282 gnd.n3009 gnd.n2477 585
R1283 gnd.n2503 gnd.n2502 585
R1284 gnd.n2504 gnd.n2503 585
R1285 gnd.n2500 gnd.n2499 585
R1286 gnd.n2500 gnd.n2467 585
R1287 gnd.n2498 gnd.n2465 585
R1288 gnd.n3017 gnd.n2465 585
R1289 gnd.n2454 gnd.n2452 585
R1290 gnd.n2979 gnd.n2454 585
R1291 gnd.n3025 gnd.n3024 585
R1292 gnd.n3024 gnd.n3023 585
R1293 gnd.n2453 gnd.n2451 585
R1294 gnd.n2518 gnd.n2453 585
R1295 gnd.n2950 gnd.n2517 585
R1296 gnd.n2969 gnd.n2517 585
R1297 gnd.n2952 gnd.n2951 585
R1298 gnd.n2953 gnd.n2952 585
R1299 gnd.n2527 gnd.n2526 585
R1300 gnd.n2533 gnd.n2526 585
R1301 gnd.n2945 gnd.n2944 585
R1302 gnd.n2944 gnd.n2943 585
R1303 gnd.n2530 gnd.n2529 585
R1304 gnd.n2541 gnd.n2530 585
R1305 gnd.n2830 gnd.n2549 585
R1306 gnd.n2922 gnd.n2549 585
R1307 gnd.n2832 gnd.n2831 585
R1308 gnd.n2831 gnd.n2547 585
R1309 gnd.n2833 gnd.n2560 585
R1310 gnd.n2912 gnd.n2560 585
R1311 gnd.n2835 gnd.n2834 585
R1312 gnd.n2835 gnd.n2567 585
R1313 gnd.n2837 gnd.n2836 585
R1314 gnd.n2836 gnd.n2566 585
R1315 gnd.n2838 gnd.n2577 585
R1316 gnd.n2892 gnd.n2577 585
R1317 gnd.n2840 gnd.n2839 585
R1318 gnd.n2839 gnd.n2575 585
R1319 gnd.n2841 gnd.n2586 585
R1320 gnd.n2881 gnd.n2586 585
R1321 gnd.n2843 gnd.n2842 585
R1322 gnd.n2843 gnd.n2592 585
R1323 gnd.n2845 gnd.n2844 585
R1324 gnd.n2844 gnd.n2591 585
R1325 gnd.n2846 gnd.n2607 585
R1326 gnd.n2860 gnd.n2607 585
R1327 gnd.n2847 gnd.n2660 585
R1328 gnd.n2660 gnd.n2599 585
R1329 gnd.n2849 gnd.n2848 585
R1330 gnd.n2850 gnd.n2849 585
R1331 gnd.n2661 gnd.n2659 585
R1332 gnd.n2659 gnd.n2658 585
R1333 gnd.n2814 gnd.n2813 585
R1334 gnd.n2813 gnd.n2812 585
R1335 gnd.n2664 gnd.n2663 585
R1336 gnd.n2665 gnd.n2664 585
R1337 gnd.n2803 gnd.n2802 585
R1338 gnd.n2804 gnd.n2803 585
R1339 gnd.n2673 gnd.n2672 585
R1340 gnd.n2672 gnd.n2671 585
R1341 gnd.n2798 gnd.n2797 585
R1342 gnd.n2797 gnd.n2796 585
R1343 gnd.n2676 gnd.n2675 585
R1344 gnd.n2787 gnd.n2676 585
R1345 gnd.n2786 gnd.n2785 585
R1346 gnd.n2788 gnd.n2786 585
R1347 gnd.n2684 gnd.n2683 585
R1348 gnd.n2683 gnd.n2682 585
R1349 gnd.n3525 gnd.n2180 585
R1350 gnd.n2180 gnd.n2157 585
R1351 gnd.n3526 gnd.n2241 585
R1352 gnd.n2241 gnd.n2231 585
R1353 gnd.n3528 gnd.n3527 585
R1354 gnd.n3529 gnd.n3528 585
R1355 gnd.n2242 gnd.n2240 585
R1356 gnd.n2249 gnd.n2240 585
R1357 gnd.n3519 gnd.n3518 585
R1358 gnd.n3518 gnd.n3517 585
R1359 gnd.n2245 gnd.n2244 585
R1360 gnd.n3244 gnd.n2245 585
R1361 gnd.n3230 gnd.n2268 585
R1362 gnd.n2268 gnd.n2258 585
R1363 gnd.n3232 gnd.n3231 585
R1364 gnd.n3233 gnd.n3232 585
R1365 gnd.n2269 gnd.n2267 585
R1366 gnd.n2267 gnd.n2265 585
R1367 gnd.n3225 gnd.n3224 585
R1368 gnd.n3224 gnd.n3223 585
R1369 gnd.n2272 gnd.n2271 585
R1370 gnd.n2281 gnd.n2272 585
R1371 gnd.n3181 gnd.n2295 585
R1372 gnd.n2295 gnd.n2280 585
R1373 gnd.n3183 gnd.n3182 585
R1374 gnd.n3184 gnd.n3183 585
R1375 gnd.n2296 gnd.n2294 585
R1376 gnd.n2303 gnd.n2294 585
R1377 gnd.n3176 gnd.n3175 585
R1378 gnd.n3175 gnd.n3174 585
R1379 gnd.n2299 gnd.n2298 585
R1380 gnd.n3155 gnd.n2299 585
R1381 gnd.n3141 gnd.n2323 585
R1382 gnd.n2323 gnd.n2312 585
R1383 gnd.n3143 gnd.n3142 585
R1384 gnd.n3144 gnd.n3143 585
R1385 gnd.n2324 gnd.n2322 585
R1386 gnd.n2322 gnd.n2319 585
R1387 gnd.n3136 gnd.n3135 585
R1388 gnd.n3135 gnd.n3134 585
R1389 gnd.n2327 gnd.n2326 585
R1390 gnd.n2337 gnd.n2327 585
R1391 gnd.n3096 gnd.n2350 585
R1392 gnd.n2350 gnd.n2336 585
R1393 gnd.n3098 gnd.n3097 585
R1394 gnd.n3099 gnd.n3098 585
R1395 gnd.n2351 gnd.n2349 585
R1396 gnd.n2358 gnd.n2349 585
R1397 gnd.n3091 gnd.n3090 585
R1398 gnd.n3090 gnd.n3089 585
R1399 gnd.n2354 gnd.n2353 585
R1400 gnd.n3070 gnd.n2354 585
R1401 gnd.n3056 gnd.n2377 585
R1402 gnd.n2377 gnd.n2367 585
R1403 gnd.n3058 gnd.n3057 585
R1404 gnd.n3059 gnd.n3058 585
R1405 gnd.n2378 gnd.n2376 585
R1406 gnd.n3047 gnd.n2376 585
R1407 gnd.n3051 gnd.n3050 585
R1408 gnd.n3050 gnd.n3049 585
R1409 gnd.n2381 gnd.n2380 585
R1410 gnd.n3002 gnd.n2381 585
R1411 gnd.n2495 gnd.n2494 585
R1412 gnd.n2496 gnd.n2495 585
R1413 gnd.n2475 gnd.n2474 585
R1414 gnd.n2478 gnd.n2475 585
R1415 gnd.n3012 gnd.n3011 585
R1416 gnd.n3011 gnd.n3010 585
R1417 gnd.n3013 gnd.n2469 585
R1418 gnd.n2505 gnd.n2469 585
R1419 gnd.n3015 gnd.n3014 585
R1420 gnd.n3016 gnd.n3015 585
R1421 gnd.n2470 gnd.n2468 585
R1422 gnd.n2980 gnd.n2468 585
R1423 gnd.n2964 gnd.n2963 585
R1424 gnd.n2963 gnd.n2456 585
R1425 gnd.n2965 gnd.n2520 585
R1426 gnd.n2520 gnd.n2455 585
R1427 gnd.n2967 gnd.n2966 585
R1428 gnd.n2968 gnd.n2967 585
R1429 gnd.n2521 gnd.n2519 585
R1430 gnd.n2519 gnd.n2516 585
R1431 gnd.n2956 gnd.n2955 585
R1432 gnd.n2955 gnd.n2954 585
R1433 gnd.n2524 gnd.n2523 585
R1434 gnd.n2531 gnd.n2524 585
R1435 gnd.n2930 gnd.n2929 585
R1436 gnd.n2931 gnd.n2930 585
R1437 gnd.n2543 gnd.n2542 585
R1438 gnd.n2550 gnd.n2542 585
R1439 gnd.n2925 gnd.n2924 585
R1440 gnd.n2924 gnd.n2923 585
R1441 gnd.n2546 gnd.n2545 585
R1442 gnd.n2913 gnd.n2546 585
R1443 gnd.n2900 gnd.n2570 585
R1444 gnd.n2570 gnd.n2569 585
R1445 gnd.n2902 gnd.n2901 585
R1446 gnd.n2903 gnd.n2902 585
R1447 gnd.n2571 gnd.n2568 585
R1448 gnd.n2578 gnd.n2568 585
R1449 gnd.n2895 gnd.n2894 585
R1450 gnd.n2894 gnd.n2893 585
R1451 gnd.n2574 gnd.n2573 585
R1452 gnd.n2882 gnd.n2574 585
R1453 gnd.n2869 gnd.n2595 585
R1454 gnd.n2595 gnd.n2594 585
R1455 gnd.n2871 gnd.n2870 585
R1456 gnd.n2872 gnd.n2871 585
R1457 gnd.n2865 gnd.n2593 585
R1458 gnd.n2864 gnd.n2863 585
R1459 gnd.n2598 gnd.n2597 585
R1460 gnd.n2861 gnd.n2598 585
R1461 gnd.n2620 gnd.n2619 585
R1462 gnd.n2623 gnd.n2622 585
R1463 gnd.n2621 gnd.n2616 585
R1464 gnd.n2628 gnd.n2627 585
R1465 gnd.n2630 gnd.n2629 585
R1466 gnd.n2633 gnd.n2632 585
R1467 gnd.n2631 gnd.n2614 585
R1468 gnd.n2638 gnd.n2637 585
R1469 gnd.n2640 gnd.n2639 585
R1470 gnd.n2643 gnd.n2642 585
R1471 gnd.n2641 gnd.n2612 585
R1472 gnd.n2648 gnd.n2647 585
R1473 gnd.n2652 gnd.n2649 585
R1474 gnd.n2653 gnd.n2590 585
R1475 gnd.n3531 gnd.n2195 585
R1476 gnd.n3598 gnd.n3597 585
R1477 gnd.n3600 gnd.n3599 585
R1478 gnd.n3602 gnd.n3601 585
R1479 gnd.n3604 gnd.n3603 585
R1480 gnd.n3606 gnd.n3605 585
R1481 gnd.n3608 gnd.n3607 585
R1482 gnd.n3610 gnd.n3609 585
R1483 gnd.n3612 gnd.n3611 585
R1484 gnd.n3614 gnd.n3613 585
R1485 gnd.n3616 gnd.n3615 585
R1486 gnd.n3618 gnd.n3617 585
R1487 gnd.n3620 gnd.n3619 585
R1488 gnd.n3623 gnd.n3622 585
R1489 gnd.n3621 gnd.n2183 585
R1490 gnd.n3627 gnd.n2181 585
R1491 gnd.n3629 gnd.n3628 585
R1492 gnd.n3630 gnd.n3629 585
R1493 gnd.n3532 gnd.n2236 585
R1494 gnd.n3532 gnd.n2157 585
R1495 gnd.n3534 gnd.n3533 585
R1496 gnd.n3533 gnd.n2231 585
R1497 gnd.n3530 gnd.n2235 585
R1498 gnd.n3530 gnd.n3529 585
R1499 gnd.n3509 gnd.n2237 585
R1500 gnd.n2249 gnd.n2237 585
R1501 gnd.n3508 gnd.n2247 585
R1502 gnd.n3517 gnd.n2247 585
R1503 gnd.n3243 gnd.n2254 585
R1504 gnd.n3244 gnd.n3243 585
R1505 gnd.n3242 gnd.n3241 585
R1506 gnd.n3242 gnd.n2258 585
R1507 gnd.n3240 gnd.n2260 585
R1508 gnd.n3233 gnd.n2260 585
R1509 gnd.n2273 gnd.n2261 585
R1510 gnd.n2273 gnd.n2265 585
R1511 gnd.n3189 gnd.n2274 585
R1512 gnd.n3223 gnd.n2274 585
R1513 gnd.n3188 gnd.n3187 585
R1514 gnd.n3187 gnd.n2281 585
R1515 gnd.n3186 gnd.n2289 585
R1516 gnd.n3186 gnd.n2280 585
R1517 gnd.n3185 gnd.n2291 585
R1518 gnd.n3185 gnd.n3184 585
R1519 gnd.n3164 gnd.n2290 585
R1520 gnd.n2303 gnd.n2290 585
R1521 gnd.n3163 gnd.n2301 585
R1522 gnd.n3174 gnd.n2301 585
R1523 gnd.n3154 gnd.n2308 585
R1524 gnd.n3155 gnd.n3154 585
R1525 gnd.n3153 gnd.n3152 585
R1526 gnd.n3153 gnd.n2312 585
R1527 gnd.n3151 gnd.n2314 585
R1528 gnd.n3144 gnd.n2314 585
R1529 gnd.n2329 gnd.n2315 585
R1530 gnd.n2329 gnd.n2319 585
R1531 gnd.n3104 gnd.n2330 585
R1532 gnd.n3134 gnd.n2330 585
R1533 gnd.n3103 gnd.n3102 585
R1534 gnd.n3102 gnd.n2337 585
R1535 gnd.n3101 gnd.n2344 585
R1536 gnd.n3101 gnd.n2336 585
R1537 gnd.n3100 gnd.n2346 585
R1538 gnd.n3100 gnd.n3099 585
R1539 gnd.n3079 gnd.n2345 585
R1540 gnd.n2358 gnd.n2345 585
R1541 gnd.n3078 gnd.n2356 585
R1542 gnd.n3089 gnd.n2356 585
R1543 gnd.n3069 gnd.n2363 585
R1544 gnd.n3070 gnd.n3069 585
R1545 gnd.n3068 gnd.n3067 585
R1546 gnd.n3068 gnd.n2367 585
R1547 gnd.n3066 gnd.n2369 585
R1548 gnd.n3059 gnd.n2369 585
R1549 gnd.n3046 gnd.n2370 585
R1550 gnd.n3047 gnd.n3046 585
R1551 gnd.n2999 gnd.n2383 585
R1552 gnd.n3049 gnd.n2383 585
R1553 gnd.n3001 gnd.n3000 585
R1554 gnd.n3002 gnd.n3001 585
R1555 gnd.n2994 gnd.n2497 585
R1556 gnd.n2497 gnd.n2496 585
R1557 gnd.n2992 gnd.n2991 585
R1558 gnd.n2991 gnd.n2478 585
R1559 gnd.n2989 gnd.n2476 585
R1560 gnd.n3010 gnd.n2476 585
R1561 gnd.n2507 gnd.n2506 585
R1562 gnd.n2506 gnd.n2505 585
R1563 gnd.n2983 gnd.n2466 585
R1564 gnd.n3016 gnd.n2466 585
R1565 gnd.n2982 gnd.n2981 585
R1566 gnd.n2981 gnd.n2980 585
R1567 gnd.n2978 gnd.n2509 585
R1568 gnd.n2978 gnd.n2456 585
R1569 gnd.n2977 gnd.n2976 585
R1570 gnd.n2977 gnd.n2455 585
R1571 gnd.n2512 gnd.n2511 585
R1572 gnd.n2968 gnd.n2511 585
R1573 gnd.n2936 gnd.n2935 585
R1574 gnd.n2935 gnd.n2516 585
R1575 gnd.n2937 gnd.n2525 585
R1576 gnd.n2954 gnd.n2525 585
R1577 gnd.n2934 gnd.n2933 585
R1578 gnd.n2933 gnd.n2531 585
R1579 gnd.n2932 gnd.n2539 585
R1580 gnd.n2932 gnd.n2931 585
R1581 gnd.n2917 gnd.n2540 585
R1582 gnd.n2550 gnd.n2540 585
R1583 gnd.n2916 gnd.n2548 585
R1584 gnd.n2923 gnd.n2548 585
R1585 gnd.n2915 gnd.n2914 585
R1586 gnd.n2914 gnd.n2913 585
R1587 gnd.n2559 gnd.n2556 585
R1588 gnd.n2569 gnd.n2559 585
R1589 gnd.n2905 gnd.n2904 585
R1590 gnd.n2904 gnd.n2903 585
R1591 gnd.n2565 gnd.n2564 585
R1592 gnd.n2578 gnd.n2565 585
R1593 gnd.n2885 gnd.n2576 585
R1594 gnd.n2893 gnd.n2576 585
R1595 gnd.n2884 gnd.n2883 585
R1596 gnd.n2883 gnd.n2882 585
R1597 gnd.n2585 gnd.n2583 585
R1598 gnd.n2594 gnd.n2585 585
R1599 gnd.n2874 gnd.n2873 585
R1600 gnd.n2873 gnd.n2872 585
R1601 gnd.n987 gnd.n985 585
R1602 gnd.n985 gnd.n979 585
R1603 gnd.n4281 gnd.n4280 585
R1604 gnd.n4282 gnd.n4281 585
R1605 gnd.n1992 gnd.n1991 585
R1606 gnd.n1999 gnd.n1991 585
R1607 gnd.n4275 gnd.n4274 585
R1608 gnd.n4274 gnd.n4273 585
R1609 gnd.n1995 gnd.n1994 585
R1610 gnd.n1996 gnd.n1995 585
R1611 gnd.n4254 gnd.n4253 585
R1612 gnd.n4255 gnd.n4254 585
R1613 gnd.n2010 gnd.n2009 585
R1614 gnd.n2009 gnd.n2006 585
R1615 gnd.n4249 gnd.n4248 585
R1616 gnd.n4248 gnd.n4247 585
R1617 gnd.n2013 gnd.n2012 585
R1618 gnd.n2023 gnd.n2013 585
R1619 gnd.n4238 gnd.n4237 585
R1620 gnd.n4239 gnd.n4238 585
R1621 gnd.n2025 gnd.n2024 585
R1622 gnd.n2032 gnd.n2024 585
R1623 gnd.n4233 gnd.n4232 585
R1624 gnd.n4232 gnd.n4231 585
R1625 gnd.n2028 gnd.n2027 585
R1626 gnd.n2029 gnd.n2028 585
R1627 gnd.n4222 gnd.n4221 585
R1628 gnd.n4223 gnd.n4222 585
R1629 gnd.n2043 gnd.n2042 585
R1630 gnd.n2042 gnd.n2039 585
R1631 gnd.n4217 gnd.n4216 585
R1632 gnd.n4216 gnd.n4215 585
R1633 gnd.n2046 gnd.n2045 585
R1634 gnd.n2047 gnd.n2046 585
R1635 gnd.n4206 gnd.n4205 585
R1636 gnd.n4207 gnd.n4206 585
R1637 gnd.n2058 gnd.n2057 585
R1638 gnd.n2065 gnd.n2057 585
R1639 gnd.n4201 gnd.n4200 585
R1640 gnd.n4200 gnd.n4199 585
R1641 gnd.n2061 gnd.n2060 585
R1642 gnd.n2062 gnd.n2061 585
R1643 gnd.n4190 gnd.n4189 585
R1644 gnd.n4191 gnd.n4190 585
R1645 gnd.n2075 gnd.n2074 585
R1646 gnd.n2074 gnd.n2071 585
R1647 gnd.n4185 gnd.n4184 585
R1648 gnd.n4184 gnd.n4183 585
R1649 gnd.n2078 gnd.n2077 585
R1650 gnd.n2079 gnd.n2078 585
R1651 gnd.n4174 gnd.n4173 585
R1652 gnd.n4175 gnd.n4174 585
R1653 gnd.n2090 gnd.n2089 585
R1654 gnd.n2097 gnd.n2089 585
R1655 gnd.n4169 gnd.n4168 585
R1656 gnd.n4168 gnd.n4167 585
R1657 gnd.n2093 gnd.n2092 585
R1658 gnd.n2094 gnd.n2093 585
R1659 gnd.n4158 gnd.n4157 585
R1660 gnd.n4159 gnd.n4158 585
R1661 gnd.n2107 gnd.n2106 585
R1662 gnd.n2106 gnd.n2103 585
R1663 gnd.n4153 gnd.n4152 585
R1664 gnd.n4152 gnd.n4151 585
R1665 gnd.n2110 gnd.n2109 585
R1666 gnd.n2111 gnd.n2110 585
R1667 gnd.n4142 gnd.n4141 585
R1668 gnd.n4143 gnd.n4142 585
R1669 gnd.n2122 gnd.n2121 585
R1670 gnd.n2129 gnd.n2121 585
R1671 gnd.n4137 gnd.n4136 585
R1672 gnd.n4136 gnd.n4135 585
R1673 gnd.n2125 gnd.n2124 585
R1674 gnd.n2126 gnd.n2125 585
R1675 gnd.n4126 gnd.n4125 585
R1676 gnd.n4127 gnd.n4126 585
R1677 gnd.n2139 gnd.n2138 585
R1678 gnd.n2138 gnd.n2135 585
R1679 gnd.n4121 gnd.n4120 585
R1680 gnd.n4120 gnd.n4119 585
R1681 gnd.n2142 gnd.n2141 585
R1682 gnd.n2143 gnd.n2142 585
R1683 gnd.n4110 gnd.n4109 585
R1684 gnd.n4111 gnd.n4110 585
R1685 gnd.n2154 gnd.n2153 585
R1686 gnd.n3634 gnd.n2153 585
R1687 gnd.n4105 gnd.n4104 585
R1688 gnd.n4104 gnd.n4103 585
R1689 gnd.n3773 gnd.n2156 585
R1690 gnd.n3776 gnd.n3775 585
R1691 gnd.n3772 gnd.n3771 585
R1692 gnd.n3771 gnd.n3631 585
R1693 gnd.n3781 gnd.n3780 585
R1694 gnd.n3783 gnd.n3770 585
R1695 gnd.n3786 gnd.n3785 585
R1696 gnd.n3768 gnd.n3767 585
R1697 gnd.n3791 gnd.n3790 585
R1698 gnd.n3793 gnd.n3766 585
R1699 gnd.n3796 gnd.n3795 585
R1700 gnd.n3764 gnd.n3763 585
R1701 gnd.n3801 gnd.n3800 585
R1702 gnd.n3803 gnd.n3762 585
R1703 gnd.n3806 gnd.n3805 585
R1704 gnd.n3760 gnd.n3759 585
R1705 gnd.n3811 gnd.n3810 585
R1706 gnd.n3813 gnd.n3755 585
R1707 gnd.n3816 gnd.n3815 585
R1708 gnd.n3753 gnd.n3752 585
R1709 gnd.n3821 gnd.n3820 585
R1710 gnd.n3823 gnd.n3751 585
R1711 gnd.n3826 gnd.n3825 585
R1712 gnd.n3749 gnd.n3748 585
R1713 gnd.n3831 gnd.n3830 585
R1714 gnd.n3833 gnd.n3747 585
R1715 gnd.n3836 gnd.n3835 585
R1716 gnd.n3745 gnd.n3744 585
R1717 gnd.n3841 gnd.n3840 585
R1718 gnd.n3843 gnd.n3743 585
R1719 gnd.n3846 gnd.n3845 585
R1720 gnd.n3741 gnd.n3740 585
R1721 gnd.n3851 gnd.n3850 585
R1722 gnd.n3853 gnd.n3739 585
R1723 gnd.n3856 gnd.n3855 585
R1724 gnd.n3737 gnd.n3736 585
R1725 gnd.n3862 gnd.n3861 585
R1726 gnd.n3864 gnd.n3735 585
R1727 gnd.n3865 gnd.n3734 585
R1728 gnd.n3868 gnd.n3867 585
R1729 gnd.n3957 gnd.n3956 585
R1730 gnd.n3956 gnd.n979 585
R1731 gnd.n3955 gnd.n1988 585
R1732 gnd.n4282 gnd.n1988 585
R1733 gnd.n3954 gnd.n3953 585
R1734 gnd.n3953 gnd.n1999 585
R1735 gnd.n3712 gnd.n1997 585
R1736 gnd.n4273 gnd.n1997 585
R1737 gnd.n3949 gnd.n3948 585
R1738 gnd.n3948 gnd.n1996 585
R1739 gnd.n3947 gnd.n2007 585
R1740 gnd.n4255 gnd.n2007 585
R1741 gnd.n3946 gnd.n3945 585
R1742 gnd.n3945 gnd.n2006 585
R1743 gnd.n3714 gnd.n2014 585
R1744 gnd.n4247 gnd.n2014 585
R1745 gnd.n3941 gnd.n3940 585
R1746 gnd.n3940 gnd.n2023 585
R1747 gnd.n3939 gnd.n2021 585
R1748 gnd.n4239 gnd.n2021 585
R1749 gnd.n3938 gnd.n3937 585
R1750 gnd.n3937 gnd.n2032 585
R1751 gnd.n3935 gnd.n2030 585
R1752 gnd.n4231 gnd.n2030 585
R1753 gnd.n3934 gnd.n3933 585
R1754 gnd.n3933 gnd.n2029 585
R1755 gnd.n3716 gnd.n2040 585
R1756 gnd.n4223 gnd.n2040 585
R1757 gnd.n3929 gnd.n3928 585
R1758 gnd.n3928 gnd.n2039 585
R1759 gnd.n3927 gnd.n2048 585
R1760 gnd.n4215 gnd.n2048 585
R1761 gnd.n3926 gnd.n3925 585
R1762 gnd.n3925 gnd.n2047 585
R1763 gnd.n3718 gnd.n2055 585
R1764 gnd.n4207 gnd.n2055 585
R1765 gnd.n3921 gnd.n3920 585
R1766 gnd.n3920 gnd.n2065 585
R1767 gnd.n3919 gnd.n2063 585
R1768 gnd.n4199 gnd.n2063 585
R1769 gnd.n3918 gnd.n3917 585
R1770 gnd.n3917 gnd.n2062 585
R1771 gnd.n3720 gnd.n2072 585
R1772 gnd.n4191 gnd.n2072 585
R1773 gnd.n3913 gnd.n3912 585
R1774 gnd.n3912 gnd.n2071 585
R1775 gnd.n3911 gnd.n2080 585
R1776 gnd.n4183 gnd.n2080 585
R1777 gnd.n3910 gnd.n3909 585
R1778 gnd.n3909 gnd.n2079 585
R1779 gnd.n3722 gnd.n2087 585
R1780 gnd.n4175 gnd.n2087 585
R1781 gnd.n3905 gnd.n3904 585
R1782 gnd.n3904 gnd.n2097 585
R1783 gnd.n3903 gnd.n2095 585
R1784 gnd.n4167 gnd.n2095 585
R1785 gnd.n3902 gnd.n3901 585
R1786 gnd.n3901 gnd.n2094 585
R1787 gnd.n3724 gnd.n2104 585
R1788 gnd.n4159 gnd.n2104 585
R1789 gnd.n3897 gnd.n3896 585
R1790 gnd.n3896 gnd.n2103 585
R1791 gnd.n3895 gnd.n2112 585
R1792 gnd.n4151 gnd.n2112 585
R1793 gnd.n3894 gnd.n3893 585
R1794 gnd.n3893 gnd.n2111 585
R1795 gnd.n3726 gnd.n2119 585
R1796 gnd.n4143 gnd.n2119 585
R1797 gnd.n3889 gnd.n3888 585
R1798 gnd.n3888 gnd.n2129 585
R1799 gnd.n3887 gnd.n2127 585
R1800 gnd.n4135 gnd.n2127 585
R1801 gnd.n3886 gnd.n3885 585
R1802 gnd.n3885 gnd.n2126 585
R1803 gnd.n3728 gnd.n2136 585
R1804 gnd.n4127 gnd.n2136 585
R1805 gnd.n3881 gnd.n3880 585
R1806 gnd.n3880 gnd.n2135 585
R1807 gnd.n3879 gnd.n2144 585
R1808 gnd.n4119 gnd.n2144 585
R1809 gnd.n3878 gnd.n3877 585
R1810 gnd.n3877 gnd.n2143 585
R1811 gnd.n3730 gnd.n2151 585
R1812 gnd.n4111 gnd.n2151 585
R1813 gnd.n3873 gnd.n3872 585
R1814 gnd.n3872 gnd.n3634 585
R1815 gnd.n3871 gnd.n3632 585
R1816 gnd.n4103 gnd.n3632 585
R1817 gnd.n4531 gnd.n4530 585
R1818 gnd.n4529 gnd.n4284 585
R1819 gnd.n4528 gnd.n4283 585
R1820 gnd.n4533 gnd.n4283 585
R1821 gnd.n4527 gnd.n4526 585
R1822 gnd.n4525 gnd.n4524 585
R1823 gnd.n4523 gnd.n4522 585
R1824 gnd.n4521 gnd.n4520 585
R1825 gnd.n4519 gnd.n4518 585
R1826 gnd.n4517 gnd.n4516 585
R1827 gnd.n4515 gnd.n4514 585
R1828 gnd.n4513 gnd.n4512 585
R1829 gnd.n4511 gnd.n4510 585
R1830 gnd.n4509 gnd.n4508 585
R1831 gnd.n4507 gnd.n4506 585
R1832 gnd.n4505 gnd.n4504 585
R1833 gnd.n4503 gnd.n4502 585
R1834 gnd.n4501 gnd.n4500 585
R1835 gnd.n4499 gnd.n4498 585
R1836 gnd.n4497 gnd.n4496 585
R1837 gnd.n4495 gnd.n4494 585
R1838 gnd.n4493 gnd.n4492 585
R1839 gnd.n4491 gnd.n4490 585
R1840 gnd.n4489 gnd.n4488 585
R1841 gnd.n4487 gnd.n4486 585
R1842 gnd.n4485 gnd.n4484 585
R1843 gnd.n4483 gnd.n4482 585
R1844 gnd.n4481 gnd.n4480 585
R1845 gnd.n4479 gnd.n4478 585
R1846 gnd.n4477 gnd.n4476 585
R1847 gnd.n4475 gnd.n4474 585
R1848 gnd.n4473 gnd.n4472 585
R1849 gnd.n4471 gnd.n4470 585
R1850 gnd.n4469 gnd.n4468 585
R1851 gnd.n4467 gnd.n4466 585
R1852 gnd.n4465 gnd.n4464 585
R1853 gnd.n4463 gnd.n4462 585
R1854 gnd.n4461 gnd.n4460 585
R1855 gnd.n4459 gnd.n4458 585
R1856 gnd.n4457 gnd.n4456 585
R1857 gnd.n4455 gnd.n4454 585
R1858 gnd.n4453 gnd.n4452 585
R1859 gnd.n4451 gnd.n4450 585
R1860 gnd.n4449 gnd.n4448 585
R1861 gnd.n4447 gnd.n4446 585
R1862 gnd.n4445 gnd.n4444 585
R1863 gnd.n4443 gnd.n4442 585
R1864 gnd.n4441 gnd.n4440 585
R1865 gnd.n4439 gnd.n4438 585
R1866 gnd.n4437 gnd.n4436 585
R1867 gnd.n4435 gnd.n4434 585
R1868 gnd.n4433 gnd.n4432 585
R1869 gnd.n4431 gnd.n4430 585
R1870 gnd.n4429 gnd.n4428 585
R1871 gnd.n4427 gnd.n4426 585
R1872 gnd.n4425 gnd.n4424 585
R1873 gnd.n4423 gnd.n4422 585
R1874 gnd.n4421 gnd.n4420 585
R1875 gnd.n4419 gnd.n4418 585
R1876 gnd.n4417 gnd.n4416 585
R1877 gnd.n4415 gnd.n4414 585
R1878 gnd.n4413 gnd.n4412 585
R1879 gnd.n4411 gnd.n4410 585
R1880 gnd.n4409 gnd.n4408 585
R1881 gnd.n4407 gnd.n4406 585
R1882 gnd.n4405 gnd.n4404 585
R1883 gnd.n4403 gnd.n4402 585
R1884 gnd.n4401 gnd.n4400 585
R1885 gnd.n4399 gnd.n4398 585
R1886 gnd.n4397 gnd.n4396 585
R1887 gnd.n4395 gnd.n4394 585
R1888 gnd.n4393 gnd.n4392 585
R1889 gnd.n4391 gnd.n4390 585
R1890 gnd.n4389 gnd.n4388 585
R1891 gnd.n4387 gnd.n4386 585
R1892 gnd.n4385 gnd.n4384 585
R1893 gnd.n4383 gnd.n4382 585
R1894 gnd.n4381 gnd.n4380 585
R1895 gnd.n4379 gnd.n4378 585
R1896 gnd.n4377 gnd.n4376 585
R1897 gnd.n4375 gnd.n4374 585
R1898 gnd.n4373 gnd.n4372 585
R1899 gnd.n4371 gnd.n4370 585
R1900 gnd.n4369 gnd.n4368 585
R1901 gnd.n1947 gnd.n1946 585
R1902 gnd.n4536 gnd.n4535 585
R1903 gnd.n978 gnd.n977 585
R1904 gnd.n6318 gnd.n978 585
R1905 gnd.n6321 gnd.n6320 585
R1906 gnd.n6320 gnd.n6319 585
R1907 gnd.n975 gnd.n974 585
R1908 gnd.n974 gnd.n973 585
R1909 gnd.n6326 gnd.n6325 585
R1910 gnd.n6327 gnd.n6326 585
R1911 gnd.n972 gnd.n971 585
R1912 gnd.n6328 gnd.n972 585
R1913 gnd.n6331 gnd.n6330 585
R1914 gnd.n6330 gnd.n6329 585
R1915 gnd.n969 gnd.n968 585
R1916 gnd.n968 gnd.n967 585
R1917 gnd.n6336 gnd.n6335 585
R1918 gnd.n6337 gnd.n6336 585
R1919 gnd.n966 gnd.n965 585
R1920 gnd.n6338 gnd.n966 585
R1921 gnd.n6341 gnd.n6340 585
R1922 gnd.n6340 gnd.n6339 585
R1923 gnd.n963 gnd.n962 585
R1924 gnd.n962 gnd.n961 585
R1925 gnd.n6346 gnd.n6345 585
R1926 gnd.n6347 gnd.n6346 585
R1927 gnd.n960 gnd.n959 585
R1928 gnd.n6348 gnd.n960 585
R1929 gnd.n6351 gnd.n6350 585
R1930 gnd.n6350 gnd.n6349 585
R1931 gnd.n957 gnd.n956 585
R1932 gnd.n956 gnd.n955 585
R1933 gnd.n6356 gnd.n6355 585
R1934 gnd.n6357 gnd.n6356 585
R1935 gnd.n954 gnd.n953 585
R1936 gnd.n6358 gnd.n954 585
R1937 gnd.n6361 gnd.n6360 585
R1938 gnd.n6360 gnd.n6359 585
R1939 gnd.n951 gnd.n950 585
R1940 gnd.n950 gnd.n949 585
R1941 gnd.n6366 gnd.n6365 585
R1942 gnd.n6367 gnd.n6366 585
R1943 gnd.n948 gnd.n947 585
R1944 gnd.n6368 gnd.n948 585
R1945 gnd.n6371 gnd.n6370 585
R1946 gnd.n6370 gnd.n6369 585
R1947 gnd.n945 gnd.n944 585
R1948 gnd.n944 gnd.n943 585
R1949 gnd.n6376 gnd.n6375 585
R1950 gnd.n6377 gnd.n6376 585
R1951 gnd.n942 gnd.n941 585
R1952 gnd.n6378 gnd.n942 585
R1953 gnd.n6381 gnd.n6380 585
R1954 gnd.n6380 gnd.n6379 585
R1955 gnd.n939 gnd.n938 585
R1956 gnd.n938 gnd.n937 585
R1957 gnd.n6386 gnd.n6385 585
R1958 gnd.n6387 gnd.n6386 585
R1959 gnd.n936 gnd.n935 585
R1960 gnd.n6388 gnd.n936 585
R1961 gnd.n6391 gnd.n6390 585
R1962 gnd.n6390 gnd.n6389 585
R1963 gnd.n933 gnd.n932 585
R1964 gnd.n932 gnd.n931 585
R1965 gnd.n6396 gnd.n6395 585
R1966 gnd.n6397 gnd.n6396 585
R1967 gnd.n930 gnd.n929 585
R1968 gnd.n6398 gnd.n930 585
R1969 gnd.n6401 gnd.n6400 585
R1970 gnd.n6400 gnd.n6399 585
R1971 gnd.n927 gnd.n926 585
R1972 gnd.n926 gnd.n925 585
R1973 gnd.n6406 gnd.n6405 585
R1974 gnd.n6407 gnd.n6406 585
R1975 gnd.n924 gnd.n923 585
R1976 gnd.n6408 gnd.n924 585
R1977 gnd.n6411 gnd.n6410 585
R1978 gnd.n6410 gnd.n6409 585
R1979 gnd.n921 gnd.n920 585
R1980 gnd.n920 gnd.n919 585
R1981 gnd.n6416 gnd.n6415 585
R1982 gnd.n6417 gnd.n6416 585
R1983 gnd.n918 gnd.n917 585
R1984 gnd.n6418 gnd.n918 585
R1985 gnd.n6421 gnd.n6420 585
R1986 gnd.n6420 gnd.n6419 585
R1987 gnd.n915 gnd.n914 585
R1988 gnd.n914 gnd.n913 585
R1989 gnd.n6426 gnd.n6425 585
R1990 gnd.n6427 gnd.n6426 585
R1991 gnd.n912 gnd.n911 585
R1992 gnd.n6428 gnd.n912 585
R1993 gnd.n6431 gnd.n6430 585
R1994 gnd.n6430 gnd.n6429 585
R1995 gnd.n909 gnd.n908 585
R1996 gnd.n908 gnd.n907 585
R1997 gnd.n6436 gnd.n6435 585
R1998 gnd.n6437 gnd.n6436 585
R1999 gnd.n906 gnd.n905 585
R2000 gnd.n6438 gnd.n906 585
R2001 gnd.n6441 gnd.n6440 585
R2002 gnd.n6440 gnd.n6439 585
R2003 gnd.n903 gnd.n902 585
R2004 gnd.n902 gnd.n901 585
R2005 gnd.n6446 gnd.n6445 585
R2006 gnd.n6447 gnd.n6446 585
R2007 gnd.n900 gnd.n899 585
R2008 gnd.n6448 gnd.n900 585
R2009 gnd.n6451 gnd.n6450 585
R2010 gnd.n6450 gnd.n6449 585
R2011 gnd.n897 gnd.n896 585
R2012 gnd.n896 gnd.n895 585
R2013 gnd.n6456 gnd.n6455 585
R2014 gnd.n6457 gnd.n6456 585
R2015 gnd.n894 gnd.n893 585
R2016 gnd.n6458 gnd.n894 585
R2017 gnd.n6461 gnd.n6460 585
R2018 gnd.n6460 gnd.n6459 585
R2019 gnd.n891 gnd.n890 585
R2020 gnd.n890 gnd.n889 585
R2021 gnd.n6466 gnd.n6465 585
R2022 gnd.n6467 gnd.n6466 585
R2023 gnd.n888 gnd.n887 585
R2024 gnd.n6468 gnd.n888 585
R2025 gnd.n6471 gnd.n6470 585
R2026 gnd.n6470 gnd.n6469 585
R2027 gnd.n885 gnd.n884 585
R2028 gnd.n884 gnd.n883 585
R2029 gnd.n6476 gnd.n6475 585
R2030 gnd.n6477 gnd.n6476 585
R2031 gnd.n882 gnd.n881 585
R2032 gnd.n6478 gnd.n882 585
R2033 gnd.n6481 gnd.n6480 585
R2034 gnd.n6480 gnd.n6479 585
R2035 gnd.n879 gnd.n878 585
R2036 gnd.n878 gnd.n877 585
R2037 gnd.n6486 gnd.n6485 585
R2038 gnd.n6487 gnd.n6486 585
R2039 gnd.n876 gnd.n875 585
R2040 gnd.n6488 gnd.n876 585
R2041 gnd.n6491 gnd.n6490 585
R2042 gnd.n6490 gnd.n6489 585
R2043 gnd.n873 gnd.n872 585
R2044 gnd.n872 gnd.n871 585
R2045 gnd.n6496 gnd.n6495 585
R2046 gnd.n6497 gnd.n6496 585
R2047 gnd.n870 gnd.n869 585
R2048 gnd.n6498 gnd.n870 585
R2049 gnd.n6501 gnd.n6500 585
R2050 gnd.n6500 gnd.n6499 585
R2051 gnd.n867 gnd.n866 585
R2052 gnd.n866 gnd.n865 585
R2053 gnd.n6506 gnd.n6505 585
R2054 gnd.n6507 gnd.n6506 585
R2055 gnd.n864 gnd.n863 585
R2056 gnd.n6508 gnd.n864 585
R2057 gnd.n6511 gnd.n6510 585
R2058 gnd.n6510 gnd.n6509 585
R2059 gnd.n861 gnd.n860 585
R2060 gnd.n860 gnd.n859 585
R2061 gnd.n6516 gnd.n6515 585
R2062 gnd.n6517 gnd.n6516 585
R2063 gnd.n858 gnd.n857 585
R2064 gnd.n6518 gnd.n858 585
R2065 gnd.n6521 gnd.n6520 585
R2066 gnd.n6520 gnd.n6519 585
R2067 gnd.n855 gnd.n854 585
R2068 gnd.n854 gnd.n853 585
R2069 gnd.n6526 gnd.n6525 585
R2070 gnd.n6527 gnd.n6526 585
R2071 gnd.n852 gnd.n851 585
R2072 gnd.n6528 gnd.n852 585
R2073 gnd.n6531 gnd.n6530 585
R2074 gnd.n6530 gnd.n6529 585
R2075 gnd.n849 gnd.n848 585
R2076 gnd.n848 gnd.n847 585
R2077 gnd.n6536 gnd.n6535 585
R2078 gnd.n6537 gnd.n6536 585
R2079 gnd.n846 gnd.n845 585
R2080 gnd.n6538 gnd.n846 585
R2081 gnd.n6541 gnd.n6540 585
R2082 gnd.n6540 gnd.n6539 585
R2083 gnd.n843 gnd.n842 585
R2084 gnd.n842 gnd.n841 585
R2085 gnd.n6546 gnd.n6545 585
R2086 gnd.n6547 gnd.n6546 585
R2087 gnd.n840 gnd.n839 585
R2088 gnd.n6548 gnd.n840 585
R2089 gnd.n6551 gnd.n6550 585
R2090 gnd.n6550 gnd.n6549 585
R2091 gnd.n837 gnd.n836 585
R2092 gnd.n836 gnd.n835 585
R2093 gnd.n6556 gnd.n6555 585
R2094 gnd.n6557 gnd.n6556 585
R2095 gnd.n834 gnd.n833 585
R2096 gnd.n6558 gnd.n834 585
R2097 gnd.n6561 gnd.n6560 585
R2098 gnd.n6560 gnd.n6559 585
R2099 gnd.n831 gnd.n830 585
R2100 gnd.n830 gnd.n829 585
R2101 gnd.n6566 gnd.n6565 585
R2102 gnd.n6567 gnd.n6566 585
R2103 gnd.n828 gnd.n827 585
R2104 gnd.n6568 gnd.n828 585
R2105 gnd.n6571 gnd.n6570 585
R2106 gnd.n6570 gnd.n6569 585
R2107 gnd.n825 gnd.n824 585
R2108 gnd.n824 gnd.n823 585
R2109 gnd.n6576 gnd.n6575 585
R2110 gnd.n6577 gnd.n6576 585
R2111 gnd.n822 gnd.n821 585
R2112 gnd.n6578 gnd.n822 585
R2113 gnd.n6581 gnd.n6580 585
R2114 gnd.n6580 gnd.n6579 585
R2115 gnd.n819 gnd.n818 585
R2116 gnd.n818 gnd.n817 585
R2117 gnd.n6586 gnd.n6585 585
R2118 gnd.n6587 gnd.n6586 585
R2119 gnd.n816 gnd.n815 585
R2120 gnd.n6588 gnd.n816 585
R2121 gnd.n6591 gnd.n6590 585
R2122 gnd.n6590 gnd.n6589 585
R2123 gnd.n813 gnd.n812 585
R2124 gnd.n812 gnd.n811 585
R2125 gnd.n6596 gnd.n6595 585
R2126 gnd.n6597 gnd.n6596 585
R2127 gnd.n810 gnd.n809 585
R2128 gnd.n6598 gnd.n810 585
R2129 gnd.n6601 gnd.n6600 585
R2130 gnd.n6600 gnd.n6599 585
R2131 gnd.n807 gnd.n806 585
R2132 gnd.n806 gnd.n805 585
R2133 gnd.n6606 gnd.n6605 585
R2134 gnd.n6607 gnd.n6606 585
R2135 gnd.n804 gnd.n803 585
R2136 gnd.n6608 gnd.n804 585
R2137 gnd.n6611 gnd.n6610 585
R2138 gnd.n6610 gnd.n6609 585
R2139 gnd.n801 gnd.n800 585
R2140 gnd.n800 gnd.n799 585
R2141 gnd.n6616 gnd.n6615 585
R2142 gnd.n6617 gnd.n6616 585
R2143 gnd.n798 gnd.n797 585
R2144 gnd.n6618 gnd.n798 585
R2145 gnd.n6621 gnd.n6620 585
R2146 gnd.n6620 gnd.n6619 585
R2147 gnd.n795 gnd.n794 585
R2148 gnd.n794 gnd.n793 585
R2149 gnd.n6626 gnd.n6625 585
R2150 gnd.n6627 gnd.n6626 585
R2151 gnd.n792 gnd.n791 585
R2152 gnd.n6628 gnd.n792 585
R2153 gnd.n6631 gnd.n6630 585
R2154 gnd.n6630 gnd.n6629 585
R2155 gnd.n789 gnd.n788 585
R2156 gnd.n788 gnd.n787 585
R2157 gnd.n6636 gnd.n6635 585
R2158 gnd.n6637 gnd.n6636 585
R2159 gnd.n786 gnd.n785 585
R2160 gnd.n6638 gnd.n786 585
R2161 gnd.n6641 gnd.n6640 585
R2162 gnd.n6640 gnd.n6639 585
R2163 gnd.n783 gnd.n782 585
R2164 gnd.n782 gnd.n781 585
R2165 gnd.n6646 gnd.n6645 585
R2166 gnd.n6647 gnd.n6646 585
R2167 gnd.n780 gnd.n779 585
R2168 gnd.n6648 gnd.n780 585
R2169 gnd.n6651 gnd.n6650 585
R2170 gnd.n6650 gnd.n6649 585
R2171 gnd.n777 gnd.n776 585
R2172 gnd.n776 gnd.n775 585
R2173 gnd.n6656 gnd.n6655 585
R2174 gnd.n6657 gnd.n6656 585
R2175 gnd.n774 gnd.n773 585
R2176 gnd.n6658 gnd.n774 585
R2177 gnd.n6661 gnd.n6660 585
R2178 gnd.n6660 gnd.n6659 585
R2179 gnd.n771 gnd.n770 585
R2180 gnd.n770 gnd.n769 585
R2181 gnd.n6666 gnd.n6665 585
R2182 gnd.n6667 gnd.n6666 585
R2183 gnd.n768 gnd.n767 585
R2184 gnd.n6668 gnd.n768 585
R2185 gnd.n6671 gnd.n6670 585
R2186 gnd.n6670 gnd.n6669 585
R2187 gnd.n765 gnd.n764 585
R2188 gnd.n764 gnd.n763 585
R2189 gnd.n6676 gnd.n6675 585
R2190 gnd.n6677 gnd.n6676 585
R2191 gnd.n762 gnd.n761 585
R2192 gnd.n6678 gnd.n762 585
R2193 gnd.n6681 gnd.n6680 585
R2194 gnd.n6680 gnd.n6679 585
R2195 gnd.n759 gnd.n758 585
R2196 gnd.n758 gnd.n757 585
R2197 gnd.n6686 gnd.n6685 585
R2198 gnd.n6687 gnd.n6686 585
R2199 gnd.n756 gnd.n755 585
R2200 gnd.n6688 gnd.n756 585
R2201 gnd.n6691 gnd.n6690 585
R2202 gnd.n6690 gnd.n6689 585
R2203 gnd.n753 gnd.n752 585
R2204 gnd.n752 gnd.n751 585
R2205 gnd.n6697 gnd.n6696 585
R2206 gnd.n6698 gnd.n6697 585
R2207 gnd.n750 gnd.n749 585
R2208 gnd.n6699 gnd.n750 585
R2209 gnd.n6702 gnd.n6701 585
R2210 gnd.n6701 gnd.n6700 585
R2211 gnd.n6703 gnd.n747 585
R2212 gnd.n747 gnd.n746 585
R2213 gnd.n622 gnd.n621 585
R2214 gnd.n6910 gnd.n621 585
R2215 gnd.n6913 gnd.n6912 585
R2216 gnd.n6912 gnd.n6911 585
R2217 gnd.n625 gnd.n624 585
R2218 gnd.n6909 gnd.n625 585
R2219 gnd.n6907 gnd.n6906 585
R2220 gnd.n6908 gnd.n6907 585
R2221 gnd.n628 gnd.n627 585
R2222 gnd.n627 gnd.n626 585
R2223 gnd.n6902 gnd.n6901 585
R2224 gnd.n6901 gnd.n6900 585
R2225 gnd.n631 gnd.n630 585
R2226 gnd.n6899 gnd.n631 585
R2227 gnd.n6897 gnd.n6896 585
R2228 gnd.n6898 gnd.n6897 585
R2229 gnd.n634 gnd.n633 585
R2230 gnd.n633 gnd.n632 585
R2231 gnd.n6892 gnd.n6891 585
R2232 gnd.n6891 gnd.n6890 585
R2233 gnd.n637 gnd.n636 585
R2234 gnd.n6889 gnd.n637 585
R2235 gnd.n6887 gnd.n6886 585
R2236 gnd.n6888 gnd.n6887 585
R2237 gnd.n640 gnd.n639 585
R2238 gnd.n639 gnd.n638 585
R2239 gnd.n6882 gnd.n6881 585
R2240 gnd.n6881 gnd.n6880 585
R2241 gnd.n643 gnd.n642 585
R2242 gnd.n6879 gnd.n643 585
R2243 gnd.n6877 gnd.n6876 585
R2244 gnd.n6878 gnd.n6877 585
R2245 gnd.n646 gnd.n645 585
R2246 gnd.n645 gnd.n644 585
R2247 gnd.n6872 gnd.n6871 585
R2248 gnd.n6871 gnd.n6870 585
R2249 gnd.n649 gnd.n648 585
R2250 gnd.n6869 gnd.n649 585
R2251 gnd.n6867 gnd.n6866 585
R2252 gnd.n6868 gnd.n6867 585
R2253 gnd.n652 gnd.n651 585
R2254 gnd.n651 gnd.n650 585
R2255 gnd.n6862 gnd.n6861 585
R2256 gnd.n6861 gnd.n6860 585
R2257 gnd.n655 gnd.n654 585
R2258 gnd.n6859 gnd.n655 585
R2259 gnd.n6857 gnd.n6856 585
R2260 gnd.n6858 gnd.n6857 585
R2261 gnd.n658 gnd.n657 585
R2262 gnd.n657 gnd.n656 585
R2263 gnd.n6852 gnd.n6851 585
R2264 gnd.n6851 gnd.n6850 585
R2265 gnd.n661 gnd.n660 585
R2266 gnd.n6849 gnd.n661 585
R2267 gnd.n6847 gnd.n6846 585
R2268 gnd.n6848 gnd.n6847 585
R2269 gnd.n664 gnd.n663 585
R2270 gnd.n663 gnd.n662 585
R2271 gnd.n6842 gnd.n6841 585
R2272 gnd.n6841 gnd.n6840 585
R2273 gnd.n667 gnd.n666 585
R2274 gnd.n6839 gnd.n667 585
R2275 gnd.n6837 gnd.n6836 585
R2276 gnd.n6838 gnd.n6837 585
R2277 gnd.n670 gnd.n669 585
R2278 gnd.n669 gnd.n668 585
R2279 gnd.n6832 gnd.n6831 585
R2280 gnd.n6831 gnd.n6830 585
R2281 gnd.n673 gnd.n672 585
R2282 gnd.n6829 gnd.n673 585
R2283 gnd.n6827 gnd.n6826 585
R2284 gnd.n6828 gnd.n6827 585
R2285 gnd.n676 gnd.n675 585
R2286 gnd.n675 gnd.n674 585
R2287 gnd.n6822 gnd.n6821 585
R2288 gnd.n6821 gnd.n6820 585
R2289 gnd.n679 gnd.n678 585
R2290 gnd.n6819 gnd.n679 585
R2291 gnd.n6817 gnd.n6816 585
R2292 gnd.n6818 gnd.n6817 585
R2293 gnd.n682 gnd.n681 585
R2294 gnd.n681 gnd.n680 585
R2295 gnd.n6812 gnd.n6811 585
R2296 gnd.n6811 gnd.n6810 585
R2297 gnd.n685 gnd.n684 585
R2298 gnd.n6809 gnd.n685 585
R2299 gnd.n6807 gnd.n6806 585
R2300 gnd.n6808 gnd.n6807 585
R2301 gnd.n688 gnd.n687 585
R2302 gnd.n687 gnd.n686 585
R2303 gnd.n6802 gnd.n6801 585
R2304 gnd.n6801 gnd.n6800 585
R2305 gnd.n691 gnd.n690 585
R2306 gnd.n6799 gnd.n691 585
R2307 gnd.n6797 gnd.n6796 585
R2308 gnd.n6798 gnd.n6797 585
R2309 gnd.n694 gnd.n693 585
R2310 gnd.n693 gnd.n692 585
R2311 gnd.n6792 gnd.n6791 585
R2312 gnd.n6791 gnd.n6790 585
R2313 gnd.n697 gnd.n696 585
R2314 gnd.n6789 gnd.n697 585
R2315 gnd.n6787 gnd.n6786 585
R2316 gnd.n6788 gnd.n6787 585
R2317 gnd.n700 gnd.n699 585
R2318 gnd.n699 gnd.n698 585
R2319 gnd.n6782 gnd.n6781 585
R2320 gnd.n6781 gnd.n6780 585
R2321 gnd.n703 gnd.n702 585
R2322 gnd.n6779 gnd.n703 585
R2323 gnd.n6777 gnd.n6776 585
R2324 gnd.n6778 gnd.n6777 585
R2325 gnd.n706 gnd.n705 585
R2326 gnd.n705 gnd.n704 585
R2327 gnd.n6772 gnd.n6771 585
R2328 gnd.n6771 gnd.n6770 585
R2329 gnd.n709 gnd.n708 585
R2330 gnd.n6769 gnd.n709 585
R2331 gnd.n6767 gnd.n6766 585
R2332 gnd.n6768 gnd.n6767 585
R2333 gnd.n712 gnd.n711 585
R2334 gnd.n711 gnd.n710 585
R2335 gnd.n6762 gnd.n6761 585
R2336 gnd.n6761 gnd.n6760 585
R2337 gnd.n715 gnd.n714 585
R2338 gnd.n6759 gnd.n715 585
R2339 gnd.n6757 gnd.n6756 585
R2340 gnd.n6758 gnd.n6757 585
R2341 gnd.n718 gnd.n717 585
R2342 gnd.n717 gnd.n716 585
R2343 gnd.n6752 gnd.n6751 585
R2344 gnd.n6751 gnd.n6750 585
R2345 gnd.n721 gnd.n720 585
R2346 gnd.n6749 gnd.n721 585
R2347 gnd.n6747 gnd.n6746 585
R2348 gnd.n6748 gnd.n6747 585
R2349 gnd.n724 gnd.n723 585
R2350 gnd.n723 gnd.n722 585
R2351 gnd.n6742 gnd.n6741 585
R2352 gnd.n6741 gnd.n6740 585
R2353 gnd.n727 gnd.n726 585
R2354 gnd.n6739 gnd.n727 585
R2355 gnd.n6737 gnd.n6736 585
R2356 gnd.n6738 gnd.n6737 585
R2357 gnd.n730 gnd.n729 585
R2358 gnd.n729 gnd.n728 585
R2359 gnd.n6732 gnd.n6731 585
R2360 gnd.n6731 gnd.n6730 585
R2361 gnd.n733 gnd.n732 585
R2362 gnd.n6729 gnd.n733 585
R2363 gnd.n6727 gnd.n6726 585
R2364 gnd.n6728 gnd.n6727 585
R2365 gnd.n736 gnd.n735 585
R2366 gnd.n735 gnd.n734 585
R2367 gnd.n6722 gnd.n6721 585
R2368 gnd.n6721 gnd.n6720 585
R2369 gnd.n739 gnd.n738 585
R2370 gnd.n6719 gnd.n739 585
R2371 gnd.n6717 gnd.n6716 585
R2372 gnd.n6718 gnd.n6717 585
R2373 gnd.n742 gnd.n741 585
R2374 gnd.n741 gnd.n740 585
R2375 gnd.n6712 gnd.n6711 585
R2376 gnd.n6711 gnd.n6710 585
R2377 gnd.n745 gnd.n744 585
R2378 gnd.n6709 gnd.n745 585
R2379 gnd.n6707 gnd.n6706 585
R2380 gnd.n6708 gnd.n6707 585
R2381 gnd.n6257 gnd.n6256 585
R2382 gnd.n6256 gnd.n6255 585
R2383 gnd.n6258 gnd.n1082 585
R2384 gnd.n6178 gnd.n1082 585
R2385 gnd.n6260 gnd.n6259 585
R2386 gnd.n6261 gnd.n6260 585
R2387 gnd.n1067 gnd.n1066 585
R2388 gnd.n4592 gnd.n1067 585
R2389 gnd.n6269 gnd.n6268 585
R2390 gnd.n6268 gnd.n6267 585
R2391 gnd.n6270 gnd.n1061 585
R2392 gnd.n4583 gnd.n1061 585
R2393 gnd.n6272 gnd.n6271 585
R2394 gnd.n6273 gnd.n6272 585
R2395 gnd.n1045 gnd.n1044 585
R2396 gnd.n4579 gnd.n1045 585
R2397 gnd.n6281 gnd.n6280 585
R2398 gnd.n6280 gnd.n6279 585
R2399 gnd.n6282 gnd.n1039 585
R2400 gnd.n4606 gnd.n1039 585
R2401 gnd.n6284 gnd.n6283 585
R2402 gnd.n6285 gnd.n6284 585
R2403 gnd.n1025 gnd.n1024 585
R2404 gnd.n4571 gnd.n1025 585
R2405 gnd.n6293 gnd.n6292 585
R2406 gnd.n6292 gnd.n6291 585
R2407 gnd.n6294 gnd.n1019 585
R2408 gnd.n4563 gnd.n1019 585
R2409 gnd.n6296 gnd.n6295 585
R2410 gnd.n6297 gnd.n6296 585
R2411 gnd.n1003 gnd.n1002 585
R2412 gnd.n3980 gnd.n1003 585
R2413 gnd.n6305 gnd.n6304 585
R2414 gnd.n6304 gnd.n6303 585
R2415 gnd.n6306 gnd.n997 585
R2416 gnd.n3967 gnd.n997 585
R2417 gnd.n6308 gnd.n6307 585
R2418 gnd.n6309 gnd.n6308 585
R2419 gnd.n998 gnd.n996 585
R2420 gnd.n3962 gnd.n996 585
R2421 gnd.n4266 gnd.n984 585
R2422 gnd.n6315 gnd.n984 585
R2423 gnd.n4724 gnd.n4723 585
R2424 gnd.n4721 gnd.n4715 585
R2425 gnd.n4731 gnd.n4712 585
R2426 gnd.n4732 gnd.n4710 585
R2427 gnd.n4709 gnd.n4702 585
R2428 gnd.n4739 gnd.n4701 585
R2429 gnd.n4740 gnd.n4700 585
R2430 gnd.n4698 gnd.n4690 585
R2431 gnd.n4747 gnd.n4689 585
R2432 gnd.n4748 gnd.n4687 585
R2433 gnd.n4686 gnd.n4679 585
R2434 gnd.n4755 gnd.n4678 585
R2435 gnd.n4756 gnd.n4677 585
R2436 gnd.n4675 gnd.n4668 585
R2437 gnd.n4763 gnd.n4667 585
R2438 gnd.n4764 gnd.n4665 585
R2439 gnd.n4664 gnd.n4656 585
R2440 gnd.n4662 gnd.n4661 585
R2441 gnd.n4657 gnd.n1087 585
R2442 gnd.n1096 gnd.n1087 585
R2443 gnd.n1166 gnd.n1090 585
R2444 gnd.n6255 gnd.n1090 585
R2445 gnd.n6177 gnd.n6176 585
R2446 gnd.n6178 gnd.n6177 585
R2447 gnd.n1165 gnd.n1081 585
R2448 gnd.n6261 gnd.n1081 585
R2449 gnd.n4594 gnd.n4593 585
R2450 gnd.n4593 gnd.n4592 585
R2451 gnd.n1926 gnd.n1070 585
R2452 gnd.n6267 gnd.n1070 585
R2453 gnd.n4598 gnd.n1925 585
R2454 gnd.n4583 gnd.n1925 585
R2455 gnd.n4599 gnd.n1059 585
R2456 gnd.n6273 gnd.n1059 585
R2457 gnd.n4600 gnd.n1924 585
R2458 gnd.n4579 gnd.n1924 585
R2459 gnd.n1921 gnd.n1048 585
R2460 gnd.n6279 gnd.n1048 585
R2461 gnd.n4605 gnd.n4604 585
R2462 gnd.n4606 gnd.n4605 585
R2463 gnd.n1920 gnd.n1038 585
R2464 gnd.n6285 gnd.n1038 585
R2465 gnd.n4570 gnd.n4569 585
R2466 gnd.n4571 gnd.n4570 585
R2467 gnd.n1933 gnd.n1027 585
R2468 gnd.n6291 gnd.n1027 585
R2469 gnd.n4565 gnd.n4564 585
R2470 gnd.n4564 gnd.n4563 585
R2471 gnd.n1935 gnd.n1017 585
R2472 gnd.n6297 gnd.n1017 585
R2473 gnd.n3982 gnd.n3981 585
R2474 gnd.n3981 gnd.n3980 585
R2475 gnd.n3985 gnd.n1006 585
R2476 gnd.n6303 gnd.n1006 585
R2477 gnd.n3986 gnd.n3707 585
R2478 gnd.n3967 gnd.n3707 585
R2479 gnd.n3987 gnd.n995 585
R2480 gnd.n6309 gnd.n995 585
R2481 gnd.n3961 gnd.n3705 585
R2482 gnd.n3962 gnd.n3961 585
R2483 gnd.n3991 gnd.n982 585
R2484 gnd.n6315 gnd.n982 585
R2485 gnd.n7533 gnd.n129 585
R2486 gnd.n7629 gnd.n129 585
R2487 gnd.n7534 gnd.n7471 585
R2488 gnd.n7471 gnd.n126 585
R2489 gnd.n7535 gnd.n207 585
R2490 gnd.n7549 gnd.n207 585
R2491 gnd.n219 gnd.n217 585
R2492 gnd.n217 gnd.n206 585
R2493 gnd.n7540 gnd.n7539 585
R2494 gnd.n7541 gnd.n7540 585
R2495 gnd.n218 gnd.n216 585
R2496 gnd.n216 gnd.n213 585
R2497 gnd.n7467 gnd.n7466 585
R2498 gnd.n7466 gnd.n7465 585
R2499 gnd.n222 gnd.n221 585
R2500 gnd.n232 gnd.n222 585
R2501 gnd.n7456 gnd.n7455 585
R2502 gnd.n7457 gnd.n7456 585
R2503 gnd.n234 gnd.n233 585
R2504 gnd.n233 gnd.n229 585
R2505 gnd.n7451 gnd.n7450 585
R2506 gnd.n7450 gnd.n7449 585
R2507 gnd.n237 gnd.n236 585
R2508 gnd.n238 gnd.n237 585
R2509 gnd.n7440 gnd.n7439 585
R2510 gnd.n7441 gnd.n7440 585
R2511 gnd.n248 gnd.n247 585
R2512 gnd.n254 gnd.n247 585
R2513 gnd.n7435 gnd.n7434 585
R2514 gnd.n7434 gnd.n7433 585
R2515 gnd.n251 gnd.n250 585
R2516 gnd.n263 gnd.n251 585
R2517 gnd.n7424 gnd.n7423 585
R2518 gnd.n7425 gnd.n7424 585
R2519 gnd.n265 gnd.n264 585
R2520 gnd.n264 gnd.n260 585
R2521 gnd.n7419 gnd.n7418 585
R2522 gnd.n7418 gnd.n7417 585
R2523 gnd.n268 gnd.n267 585
R2524 gnd.n269 gnd.n268 585
R2525 gnd.n7408 gnd.n7407 585
R2526 gnd.n7409 gnd.n7408 585
R2527 gnd.n279 gnd.n278 585
R2528 gnd.n284 gnd.n278 585
R2529 gnd.n7403 gnd.n7402 585
R2530 gnd.n7402 gnd.n7401 585
R2531 gnd.n282 gnd.n281 585
R2532 gnd.n293 gnd.n282 585
R2533 gnd.n7392 gnd.n7391 585
R2534 gnd.n7393 gnd.n7392 585
R2535 gnd.n295 gnd.n294 585
R2536 gnd.n294 gnd.n290 585
R2537 gnd.n7387 gnd.n7386 585
R2538 gnd.n7386 gnd.n7385 585
R2539 gnd.n298 gnd.n297 585
R2540 gnd.n299 gnd.n298 585
R2541 gnd.n7376 gnd.n7375 585
R2542 gnd.n7377 gnd.n7376 585
R2543 gnd.n309 gnd.n308 585
R2544 gnd.n314 gnd.n308 585
R2545 gnd.n7371 gnd.n7370 585
R2546 gnd.n7370 gnd.n7369 585
R2547 gnd.n312 gnd.n311 585
R2548 gnd.n323 gnd.n312 585
R2549 gnd.n7360 gnd.n7359 585
R2550 gnd.n7361 gnd.n7360 585
R2551 gnd.n325 gnd.n324 585
R2552 gnd.n324 gnd.n320 585
R2553 gnd.n7355 gnd.n7354 585
R2554 gnd.n7354 gnd.n7353 585
R2555 gnd.n329 gnd.n328 585
R2556 gnd.n330 gnd.n329 585
R2557 gnd.n7344 gnd.n7343 585
R2558 gnd.n7345 gnd.n7344 585
R2559 gnd.n342 gnd.n341 585
R2560 gnd.n341 gnd.n338 585
R2561 gnd.n7339 gnd.n7338 585
R2562 gnd.n7338 gnd.n7337 585
R2563 gnd.n345 gnd.n344 585
R2564 gnd.n356 gnd.n345 585
R2565 gnd.n7328 gnd.n7327 585
R2566 gnd.n7329 gnd.n7328 585
R2567 gnd.n358 gnd.n357 585
R2568 gnd.n357 gnd.n353 585
R2569 gnd.n7323 gnd.n7322 585
R2570 gnd.n7322 gnd.n7321 585
R2571 gnd.n361 gnd.n360 585
R2572 gnd.n362 gnd.n361 585
R2573 gnd.n7312 gnd.n7311 585
R2574 gnd.n7313 gnd.n7312 585
R2575 gnd.n375 gnd.n374 585
R2576 gnd.n7040 gnd.n374 585
R2577 gnd.n7307 gnd.n7306 585
R2578 gnd.n7306 gnd.n7305 585
R2579 gnd.n378 gnd.n377 585
R2580 gnd.n6928 gnd.n378 585
R2581 gnd.n7296 gnd.n7295 585
R2582 gnd.n7297 gnd.n7296 585
R2583 gnd.n392 gnd.n391 585
R2584 gnd.n5882 gnd.n391 585
R2585 gnd.n7291 gnd.n7290 585
R2586 gnd.n7290 gnd.n7289 585
R2587 gnd.n395 gnd.n394 585
R2588 gnd.n5907 gnd.n395 585
R2589 gnd.n7280 gnd.n7279 585
R2590 gnd.n7281 gnd.n7280 585
R2591 gnd.n409 gnd.n408 585
R2592 gnd.n5911 gnd.n408 585
R2593 gnd.n7275 gnd.n7274 585
R2594 gnd.n7274 gnd.n7273 585
R2595 gnd.n412 gnd.n411 585
R2596 gnd.n5917 gnd.n412 585
R2597 gnd.n7264 gnd.n7263 585
R2598 gnd.n7265 gnd.n7264 585
R2599 gnd.n426 gnd.n425 585
R2600 gnd.n5870 gnd.n425 585
R2601 gnd.n7259 gnd.n7258 585
R2602 gnd.n7258 gnd.n7257 585
R2603 gnd.n429 gnd.n428 585
R2604 gnd.n5866 gnd.n429 585
R2605 gnd.n7248 gnd.n7247 585
R2606 gnd.n7249 gnd.n7248 585
R2607 gnd.n444 gnd.n443 585
R2608 gnd.n7098 gnd.n443 585
R2609 gnd.n7243 gnd.n7242 585
R2610 gnd.n7242 gnd.n7241 585
R2611 gnd.n447 gnd.n446 585
R2612 gnd.n5973 gnd.n447 585
R2613 gnd.n7232 gnd.n7231 585
R2614 gnd.n7233 gnd.n7232 585
R2615 gnd.n7228 gnd.n459 585
R2616 gnd.n7227 gnd.n461 585
R2617 gnd.n531 gnd.n462 585
R2618 gnd.n7220 gnd.n468 585
R2619 gnd.n7219 gnd.n469 585
R2620 gnd.n533 gnd.n470 585
R2621 gnd.n7212 gnd.n476 585
R2622 gnd.n7211 gnd.n477 585
R2623 gnd.n536 gnd.n478 585
R2624 gnd.n7204 gnd.n484 585
R2625 gnd.n7203 gnd.n485 585
R2626 gnd.n538 gnd.n486 585
R2627 gnd.n7196 gnd.n492 585
R2628 gnd.n7195 gnd.n493 585
R2629 gnd.n541 gnd.n494 585
R2630 gnd.n7188 gnd.n500 585
R2631 gnd.n7187 gnd.n501 585
R2632 gnd.n510 gnd.n504 585
R2633 gnd.n7180 gnd.n7179 585
R2634 gnd.n7179 gnd.n7178 585
R2635 gnd.n7632 gnd.n7631 585
R2636 gnd.n7504 gnd.n124 585
R2637 gnd.n7506 gnd.n7505 585
R2638 gnd.n7502 gnd.n7501 585
R2639 gnd.n7510 gnd.n7500 585
R2640 gnd.n7511 gnd.n7498 585
R2641 gnd.n7512 gnd.n7497 585
R2642 gnd.n7495 gnd.n7493 585
R2643 gnd.n7516 gnd.n7492 585
R2644 gnd.n7517 gnd.n7490 585
R2645 gnd.n7518 gnd.n7489 585
R2646 gnd.n7487 gnd.n7485 585
R2647 gnd.n7522 gnd.n7484 585
R2648 gnd.n7523 gnd.n7482 585
R2649 gnd.n7524 gnd.n7481 585
R2650 gnd.n7479 gnd.n7477 585
R2651 gnd.n7528 gnd.n7476 585
R2652 gnd.n7529 gnd.n7474 585
R2653 gnd.n7530 gnd.n7473 585
R2654 gnd.n7473 gnd.n128 585
R2655 gnd.n7630 gnd.n120 585
R2656 gnd.n7630 gnd.n7629 585
R2657 gnd.n7636 gnd.n119 585
R2658 gnd.n126 gnd.n119 585
R2659 gnd.n7637 gnd.n118 585
R2660 gnd.n7549 gnd.n118 585
R2661 gnd.n7638 gnd.n117 585
R2662 gnd.n206 gnd.n117 585
R2663 gnd.n215 gnd.n115 585
R2664 gnd.n7541 gnd.n215 585
R2665 gnd.n7642 gnd.n114 585
R2666 gnd.n213 gnd.n114 585
R2667 gnd.n7643 gnd.n113 585
R2668 gnd.n7465 gnd.n113 585
R2669 gnd.n7644 gnd.n112 585
R2670 gnd.n232 gnd.n112 585
R2671 gnd.n231 gnd.n110 585
R2672 gnd.n7457 gnd.n231 585
R2673 gnd.n7648 gnd.n109 585
R2674 gnd.n229 gnd.n109 585
R2675 gnd.n7649 gnd.n108 585
R2676 gnd.n7449 gnd.n108 585
R2677 gnd.n7650 gnd.n107 585
R2678 gnd.n238 gnd.n107 585
R2679 gnd.n246 gnd.n105 585
R2680 gnd.n7441 gnd.n246 585
R2681 gnd.n7654 gnd.n104 585
R2682 gnd.n254 gnd.n104 585
R2683 gnd.n7655 gnd.n103 585
R2684 gnd.n7433 gnd.n103 585
R2685 gnd.n7656 gnd.n102 585
R2686 gnd.n263 gnd.n102 585
R2687 gnd.n262 gnd.n100 585
R2688 gnd.n7425 gnd.n262 585
R2689 gnd.n7660 gnd.n99 585
R2690 gnd.n260 gnd.n99 585
R2691 gnd.n7661 gnd.n98 585
R2692 gnd.n7417 gnd.n98 585
R2693 gnd.n7662 gnd.n97 585
R2694 gnd.n269 gnd.n97 585
R2695 gnd.n277 gnd.n95 585
R2696 gnd.n7409 gnd.n277 585
R2697 gnd.n7666 gnd.n94 585
R2698 gnd.n284 gnd.n94 585
R2699 gnd.n7667 gnd.n93 585
R2700 gnd.n7401 gnd.n93 585
R2701 gnd.n7668 gnd.n92 585
R2702 gnd.n293 gnd.n92 585
R2703 gnd.n292 gnd.n90 585
R2704 gnd.n7393 gnd.n292 585
R2705 gnd.n7672 gnd.n89 585
R2706 gnd.n290 gnd.n89 585
R2707 gnd.n7673 gnd.n88 585
R2708 gnd.n7385 gnd.n88 585
R2709 gnd.n7674 gnd.n87 585
R2710 gnd.n299 gnd.n87 585
R2711 gnd.n307 gnd.n85 585
R2712 gnd.n7377 gnd.n307 585
R2713 gnd.n7678 gnd.n84 585
R2714 gnd.n314 gnd.n84 585
R2715 gnd.n7679 gnd.n83 585
R2716 gnd.n7369 gnd.n83 585
R2717 gnd.n7680 gnd.n82 585
R2718 gnd.n323 gnd.n82 585
R2719 gnd.n322 gnd.n80 585
R2720 gnd.n7361 gnd.n322 585
R2721 gnd.n7054 gnd.n7053 585
R2722 gnd.n7053 gnd.n320 585
R2723 gnd.n7055 gnd.n332 585
R2724 gnd.n7353 gnd.n332 585
R2725 gnd.n7056 gnd.n7052 585
R2726 gnd.n7052 gnd.n330 585
R2727 gnd.n7050 gnd.n340 585
R2728 gnd.n7345 gnd.n340 585
R2729 gnd.n7060 gnd.n7049 585
R2730 gnd.n7049 gnd.n338 585
R2731 gnd.n7061 gnd.n347 585
R2732 gnd.n7337 gnd.n347 585
R2733 gnd.n7062 gnd.n7048 585
R2734 gnd.n7048 gnd.n356 585
R2735 gnd.n7046 gnd.n355 585
R2736 gnd.n7329 gnd.n355 585
R2737 gnd.n7066 gnd.n7045 585
R2738 gnd.n7045 gnd.n353 585
R2739 gnd.n7067 gnd.n364 585
R2740 gnd.n7321 gnd.n364 585
R2741 gnd.n7068 gnd.n7044 585
R2742 gnd.n7044 gnd.n362 585
R2743 gnd.n7042 gnd.n373 585
R2744 gnd.n7313 gnd.n373 585
R2745 gnd.n7072 gnd.n7041 585
R2746 gnd.n7041 gnd.n7040 585
R2747 gnd.n7073 gnd.n380 585
R2748 gnd.n7305 gnd.n380 585
R2749 gnd.n7074 gnd.n610 585
R2750 gnd.n6928 gnd.n610 585
R2751 gnd.n608 gnd.n389 585
R2752 gnd.n7297 gnd.n389 585
R2753 gnd.n7078 gnd.n607 585
R2754 gnd.n5882 gnd.n607 585
R2755 gnd.n7079 gnd.n398 585
R2756 gnd.n7289 gnd.n398 585
R2757 gnd.n7080 gnd.n606 585
R2758 gnd.n5907 gnd.n606 585
R2759 gnd.n604 gnd.n407 585
R2760 gnd.n7281 gnd.n407 585
R2761 gnd.n7084 gnd.n603 585
R2762 gnd.n5911 gnd.n603 585
R2763 gnd.n7085 gnd.n414 585
R2764 gnd.n7273 gnd.n414 585
R2765 gnd.n7086 gnd.n602 585
R2766 gnd.n5917 gnd.n602 585
R2767 gnd.n600 gnd.n423 585
R2768 gnd.n7265 gnd.n423 585
R2769 gnd.n7090 gnd.n599 585
R2770 gnd.n5870 gnd.n599 585
R2771 gnd.n7091 gnd.n432 585
R2772 gnd.n7257 gnd.n432 585
R2773 gnd.n7092 gnd.n598 585
R2774 gnd.n5866 gnd.n598 585
R2775 gnd.n595 gnd.n441 585
R2776 gnd.n7249 gnd.n441 585
R2777 gnd.n7097 gnd.n7096 585
R2778 gnd.n7098 gnd.n7097 585
R2779 gnd.n594 gnd.n449 585
R2780 gnd.n7241 gnd.n449 585
R2781 gnd.n5972 gnd.n5971 585
R2782 gnd.n5973 gnd.n5972 585
R2783 gnd.n5931 gnd.n457 585
R2784 gnd.n7233 gnd.n457 585
R2785 gnd.n6254 gnd.n6253 585
R2786 gnd.n6255 gnd.n6254 585
R2787 gnd.n1078 gnd.n1077 585
R2788 gnd.n6178 gnd.n1078 585
R2789 gnd.n6263 gnd.n6262 585
R2790 gnd.n6262 gnd.n6261 585
R2791 gnd.n6264 gnd.n1072 585
R2792 gnd.n4592 gnd.n1072 585
R2793 gnd.n6266 gnd.n6265 585
R2794 gnd.n6267 gnd.n6266 585
R2795 gnd.n1056 gnd.n1055 585
R2796 gnd.n4583 gnd.n1056 585
R2797 gnd.n6275 gnd.n6274 585
R2798 gnd.n6274 gnd.n6273 585
R2799 gnd.n6276 gnd.n1050 585
R2800 gnd.n4579 gnd.n1050 585
R2801 gnd.n6278 gnd.n6277 585
R2802 gnd.n6279 gnd.n6278 585
R2803 gnd.n1035 gnd.n1034 585
R2804 gnd.n4606 gnd.n1035 585
R2805 gnd.n6287 gnd.n6286 585
R2806 gnd.n6286 gnd.n6285 585
R2807 gnd.n6288 gnd.n1029 585
R2808 gnd.n4571 gnd.n1029 585
R2809 gnd.n6290 gnd.n6289 585
R2810 gnd.n6291 gnd.n6290 585
R2811 gnd.n1014 gnd.n1013 585
R2812 gnd.n4563 gnd.n1014 585
R2813 gnd.n6299 gnd.n6298 585
R2814 gnd.n6298 gnd.n6297 585
R2815 gnd.n6300 gnd.n1008 585
R2816 gnd.n3980 gnd.n1008 585
R2817 gnd.n6302 gnd.n6301 585
R2818 gnd.n6303 gnd.n6302 585
R2819 gnd.n992 gnd.n991 585
R2820 gnd.n3967 gnd.n992 585
R2821 gnd.n6311 gnd.n6310 585
R2822 gnd.n6310 gnd.n6309 585
R2823 gnd.n6312 gnd.n986 585
R2824 gnd.n3962 gnd.n986 585
R2825 gnd.n6314 gnd.n6313 585
R2826 gnd.n6315 gnd.n6314 585
R2827 gnd.n6185 gnd.n6184 585
R2828 gnd.n6187 gnd.n1159 585
R2829 gnd.n6189 gnd.n6188 585
R2830 gnd.n6190 gnd.n1152 585
R2831 gnd.n6192 gnd.n6191 585
R2832 gnd.n6194 gnd.n1150 585
R2833 gnd.n6196 gnd.n6195 585
R2834 gnd.n6197 gnd.n1145 585
R2835 gnd.n6199 gnd.n6198 585
R2836 gnd.n6201 gnd.n1143 585
R2837 gnd.n6203 gnd.n6202 585
R2838 gnd.n6204 gnd.n1138 585
R2839 gnd.n6206 gnd.n6205 585
R2840 gnd.n6208 gnd.n1136 585
R2841 gnd.n6210 gnd.n6209 585
R2842 gnd.n6211 gnd.n1131 585
R2843 gnd.n6213 gnd.n6212 585
R2844 gnd.n6215 gnd.n1129 585
R2845 gnd.n6217 gnd.n6216 585
R2846 gnd.n6218 gnd.n1123 585
R2847 gnd.n6220 gnd.n6219 585
R2848 gnd.n6224 gnd.n1118 585
R2849 gnd.n6226 gnd.n6225 585
R2850 gnd.n6227 gnd.n1113 585
R2851 gnd.n6229 gnd.n6228 585
R2852 gnd.n6231 gnd.n1111 585
R2853 gnd.n6233 gnd.n6232 585
R2854 gnd.n6234 gnd.n1106 585
R2855 gnd.n6236 gnd.n6235 585
R2856 gnd.n6238 gnd.n1104 585
R2857 gnd.n6240 gnd.n6239 585
R2858 gnd.n6241 gnd.n1098 585
R2859 gnd.n6243 gnd.n6242 585
R2860 gnd.n6245 gnd.n1097 585
R2861 gnd.n6246 gnd.n1095 585
R2862 gnd.n6249 gnd.n6248 585
R2863 gnd.n6250 gnd.n1092 585
R2864 gnd.n1096 gnd.n1092 585
R2865 gnd.n6181 gnd.n1089 585
R2866 gnd.n6255 gnd.n1089 585
R2867 gnd.n6180 gnd.n6179 585
R2868 gnd.n6179 gnd.n6178 585
R2869 gnd.n1163 gnd.n1080 585
R2870 gnd.n6261 gnd.n1080 585
R2871 gnd.n4591 gnd.n4590 585
R2872 gnd.n4592 gnd.n4591 585
R2873 gnd.n1927 gnd.n1069 585
R2874 gnd.n6267 gnd.n1069 585
R2875 gnd.n4585 gnd.n4584 585
R2876 gnd.n4584 gnd.n4583 585
R2877 gnd.n4582 gnd.n1058 585
R2878 gnd.n6273 gnd.n1058 585
R2879 gnd.n4581 gnd.n4580 585
R2880 gnd.n4580 gnd.n4579 585
R2881 gnd.n1929 gnd.n1047 585
R2882 gnd.n6279 gnd.n1047 585
R2883 gnd.n4575 gnd.n1919 585
R2884 gnd.n4606 gnd.n1919 585
R2885 gnd.n4574 gnd.n1037 585
R2886 gnd.n6285 gnd.n1037 585
R2887 gnd.n4573 gnd.n4572 585
R2888 gnd.n4572 gnd.n4571 585
R2889 gnd.n1931 gnd.n1026 585
R2890 gnd.n6291 gnd.n1026 585
R2891 gnd.n3976 gnd.n1936 585
R2892 gnd.n4563 gnd.n1936 585
R2893 gnd.n3977 gnd.n1016 585
R2894 gnd.n6297 gnd.n1016 585
R2895 gnd.n3979 gnd.n3978 585
R2896 gnd.n3980 gnd.n3979 585
R2897 gnd.n3708 gnd.n1005 585
R2898 gnd.n6303 gnd.n1005 585
R2899 gnd.n3969 gnd.n3968 585
R2900 gnd.n3968 gnd.n3967 585
R2901 gnd.n3965 gnd.n994 585
R2902 gnd.n6309 gnd.n994 585
R2903 gnd.n3964 gnd.n3963 585
R2904 gnd.n3963 gnd.n3962 585
R2905 gnd.n3710 gnd.n981 585
R2906 gnd.n6315 gnd.n981 585
R2907 gnd.n7628 gnd.n7627 585
R2908 gnd.n7629 gnd.n7628 585
R2909 gnd.n132 gnd.n130 585
R2910 gnd.n130 gnd.n126 585
R2911 gnd.n7548 gnd.n7547 585
R2912 gnd.n7549 gnd.n7548 585
R2913 gnd.n209 gnd.n208 585
R2914 gnd.n208 gnd.n206 585
R2915 gnd.n7543 gnd.n7542 585
R2916 gnd.n7542 gnd.n7541 585
R2917 gnd.n212 gnd.n211 585
R2918 gnd.n213 gnd.n212 585
R2919 gnd.n7464 gnd.n7463 585
R2920 gnd.n7465 gnd.n7464 585
R2921 gnd.n225 gnd.n224 585
R2922 gnd.n232 gnd.n224 585
R2923 gnd.n7459 gnd.n7458 585
R2924 gnd.n7458 gnd.n7457 585
R2925 gnd.n228 gnd.n227 585
R2926 gnd.n229 gnd.n228 585
R2927 gnd.n7448 gnd.n7447 585
R2928 gnd.n7449 gnd.n7448 585
R2929 gnd.n241 gnd.n240 585
R2930 gnd.n240 gnd.n238 585
R2931 gnd.n7443 gnd.n7442 585
R2932 gnd.n7442 gnd.n7441 585
R2933 gnd.n244 gnd.n243 585
R2934 gnd.n254 gnd.n244 585
R2935 gnd.n7432 gnd.n7431 585
R2936 gnd.n7433 gnd.n7432 585
R2937 gnd.n256 gnd.n255 585
R2938 gnd.n263 gnd.n255 585
R2939 gnd.n7427 gnd.n7426 585
R2940 gnd.n7426 gnd.n7425 585
R2941 gnd.n259 gnd.n258 585
R2942 gnd.n260 gnd.n259 585
R2943 gnd.n7416 gnd.n7415 585
R2944 gnd.n7417 gnd.n7416 585
R2945 gnd.n272 gnd.n271 585
R2946 gnd.n271 gnd.n269 585
R2947 gnd.n7411 gnd.n7410 585
R2948 gnd.n7410 gnd.n7409 585
R2949 gnd.n275 gnd.n274 585
R2950 gnd.n284 gnd.n275 585
R2951 gnd.n7400 gnd.n7399 585
R2952 gnd.n7401 gnd.n7400 585
R2953 gnd.n286 gnd.n285 585
R2954 gnd.n293 gnd.n285 585
R2955 gnd.n7395 gnd.n7394 585
R2956 gnd.n7394 gnd.n7393 585
R2957 gnd.n289 gnd.n288 585
R2958 gnd.n290 gnd.n289 585
R2959 gnd.n7384 gnd.n7383 585
R2960 gnd.n7385 gnd.n7384 585
R2961 gnd.n302 gnd.n301 585
R2962 gnd.n301 gnd.n299 585
R2963 gnd.n7379 gnd.n7378 585
R2964 gnd.n7378 gnd.n7377 585
R2965 gnd.n305 gnd.n304 585
R2966 gnd.n314 gnd.n305 585
R2967 gnd.n7368 gnd.n7367 585
R2968 gnd.n7369 gnd.n7368 585
R2969 gnd.n316 gnd.n315 585
R2970 gnd.n323 gnd.n315 585
R2971 gnd.n7363 gnd.n7362 585
R2972 gnd.n7362 gnd.n7361 585
R2973 gnd.n319 gnd.n318 585
R2974 gnd.n320 gnd.n319 585
R2975 gnd.n7352 gnd.n7351 585
R2976 gnd.n7353 gnd.n7352 585
R2977 gnd.n334 gnd.n333 585
R2978 gnd.n333 gnd.n330 585
R2979 gnd.n7347 gnd.n7346 585
R2980 gnd.n7346 gnd.n7345 585
R2981 gnd.n337 gnd.n336 585
R2982 gnd.n338 gnd.n337 585
R2983 gnd.n7336 gnd.n7335 585
R2984 gnd.n7337 gnd.n7336 585
R2985 gnd.n349 gnd.n348 585
R2986 gnd.n356 gnd.n348 585
R2987 gnd.n7331 gnd.n7330 585
R2988 gnd.n7330 gnd.n7329 585
R2989 gnd.n352 gnd.n351 585
R2990 gnd.n353 gnd.n352 585
R2991 gnd.n7320 gnd.n7319 585
R2992 gnd.n7321 gnd.n7320 585
R2993 gnd.n367 gnd.n366 585
R2994 gnd.n366 gnd.n362 585
R2995 gnd.n7315 gnd.n7314 585
R2996 gnd.n7314 gnd.n7313 585
R2997 gnd.n370 gnd.n369 585
R2998 gnd.n7040 gnd.n370 585
R2999 gnd.n7304 gnd.n7303 585
R3000 gnd.n7305 gnd.n7304 585
R3001 gnd.n383 gnd.n382 585
R3002 gnd.n6928 gnd.n382 585
R3003 gnd.n7299 gnd.n7298 585
R3004 gnd.n7298 gnd.n7297 585
R3005 gnd.n386 gnd.n385 585
R3006 gnd.n5882 gnd.n386 585
R3007 gnd.n7288 gnd.n7287 585
R3008 gnd.n7289 gnd.n7288 585
R3009 gnd.n401 gnd.n400 585
R3010 gnd.n5907 gnd.n400 585
R3011 gnd.n7283 gnd.n7282 585
R3012 gnd.n7282 gnd.n7281 585
R3013 gnd.n404 gnd.n403 585
R3014 gnd.n5911 gnd.n404 585
R3015 gnd.n7272 gnd.n7271 585
R3016 gnd.n7273 gnd.n7272 585
R3017 gnd.n417 gnd.n416 585
R3018 gnd.n5917 gnd.n416 585
R3019 gnd.n7267 gnd.n7266 585
R3020 gnd.n7266 gnd.n7265 585
R3021 gnd.n420 gnd.n419 585
R3022 gnd.n5870 gnd.n420 585
R3023 gnd.n7256 gnd.n7255 585
R3024 gnd.n7257 gnd.n7256 585
R3025 gnd.n435 gnd.n434 585
R3026 gnd.n5866 gnd.n434 585
R3027 gnd.n7251 gnd.n7250 585
R3028 gnd.n7250 gnd.n7249 585
R3029 gnd.n438 gnd.n437 585
R3030 gnd.n7098 gnd.n438 585
R3031 gnd.n7240 gnd.n7239 585
R3032 gnd.n7241 gnd.n7240 585
R3033 gnd.n452 gnd.n451 585
R3034 gnd.n5973 gnd.n451 585
R3035 gnd.n7235 gnd.n7234 585
R3036 gnd.n7234 gnd.n7233 585
R3037 gnd.n545 gnd.n454 585
R3038 gnd.n7176 gnd.n7175 585
R3039 gnd.n7174 gnd.n544 585
R3040 gnd.n7178 gnd.n544 585
R3041 gnd.n7173 gnd.n7172 585
R3042 gnd.n7171 gnd.n7170 585
R3043 gnd.n7169 gnd.n7168 585
R3044 gnd.n7167 gnd.n7166 585
R3045 gnd.n7165 gnd.n7164 585
R3046 gnd.n7163 gnd.n7162 585
R3047 gnd.n7161 gnd.n7160 585
R3048 gnd.n7159 gnd.n7158 585
R3049 gnd.n7157 gnd.n7156 585
R3050 gnd.n7155 gnd.n7154 585
R3051 gnd.n7153 gnd.n7152 585
R3052 gnd.n7151 gnd.n7150 585
R3053 gnd.n7149 gnd.n7148 585
R3054 gnd.n7146 gnd.n7145 585
R3055 gnd.n7144 gnd.n7143 585
R3056 gnd.n7142 gnd.n7141 585
R3057 gnd.n7140 gnd.n7139 585
R3058 gnd.n7138 gnd.n7137 585
R3059 gnd.n7136 gnd.n7135 585
R3060 gnd.n7134 gnd.n7133 585
R3061 gnd.n7132 gnd.n7131 585
R3062 gnd.n7130 gnd.n7129 585
R3063 gnd.n7128 gnd.n7127 585
R3064 gnd.n7126 gnd.n7125 585
R3065 gnd.n7124 gnd.n7123 585
R3066 gnd.n7122 gnd.n7121 585
R3067 gnd.n7120 gnd.n7119 585
R3068 gnd.n7118 gnd.n7117 585
R3069 gnd.n7116 gnd.n7115 585
R3070 gnd.n7114 gnd.n7113 585
R3071 gnd.n7112 gnd.n7111 585
R3072 gnd.n7110 gnd.n584 585
R3073 gnd.n588 gnd.n585 585
R3074 gnd.n7106 gnd.n7105 585
R3075 gnd.n200 gnd.n199 585
R3076 gnd.n7557 gnd.n195 585
R3077 gnd.n7559 gnd.n7558 585
R3078 gnd.n7561 gnd.n193 585
R3079 gnd.n7563 gnd.n7562 585
R3080 gnd.n7564 gnd.n188 585
R3081 gnd.n7566 gnd.n7565 585
R3082 gnd.n7568 gnd.n186 585
R3083 gnd.n7570 gnd.n7569 585
R3084 gnd.n7571 gnd.n181 585
R3085 gnd.n7573 gnd.n7572 585
R3086 gnd.n7575 gnd.n179 585
R3087 gnd.n7577 gnd.n7576 585
R3088 gnd.n7578 gnd.n174 585
R3089 gnd.n7580 gnd.n7579 585
R3090 gnd.n7582 gnd.n172 585
R3091 gnd.n7584 gnd.n7583 585
R3092 gnd.n7585 gnd.n167 585
R3093 gnd.n7587 gnd.n7586 585
R3094 gnd.n7589 gnd.n165 585
R3095 gnd.n7591 gnd.n7590 585
R3096 gnd.n7595 gnd.n160 585
R3097 gnd.n7597 gnd.n7596 585
R3098 gnd.n7599 gnd.n158 585
R3099 gnd.n7601 gnd.n7600 585
R3100 gnd.n7602 gnd.n153 585
R3101 gnd.n7604 gnd.n7603 585
R3102 gnd.n7606 gnd.n151 585
R3103 gnd.n7608 gnd.n7607 585
R3104 gnd.n7609 gnd.n146 585
R3105 gnd.n7611 gnd.n7610 585
R3106 gnd.n7613 gnd.n144 585
R3107 gnd.n7615 gnd.n7614 585
R3108 gnd.n7616 gnd.n139 585
R3109 gnd.n7618 gnd.n7617 585
R3110 gnd.n7620 gnd.n137 585
R3111 gnd.n7622 gnd.n7621 585
R3112 gnd.n7623 gnd.n135 585
R3113 gnd.n7624 gnd.n131 585
R3114 gnd.n131 gnd.n128 585
R3115 gnd.n7553 gnd.n127 585
R3116 gnd.n7629 gnd.n127 585
R3117 gnd.n7552 gnd.n7551 585
R3118 gnd.n7551 gnd.n126 585
R3119 gnd.n7550 gnd.n204 585
R3120 gnd.n7550 gnd.n7549 585
R3121 gnd.n6976 gnd.n205 585
R3122 gnd.n206 gnd.n205 585
R3123 gnd.n6977 gnd.n214 585
R3124 gnd.n7541 gnd.n214 585
R3125 gnd.n6979 gnd.n6978 585
R3126 gnd.n6978 gnd.n213 585
R3127 gnd.n6980 gnd.n223 585
R3128 gnd.n7465 gnd.n223 585
R3129 gnd.n6982 gnd.n6981 585
R3130 gnd.n6981 gnd.n232 585
R3131 gnd.n6983 gnd.n230 585
R3132 gnd.n7457 gnd.n230 585
R3133 gnd.n6985 gnd.n6984 585
R3134 gnd.n6984 gnd.n229 585
R3135 gnd.n6986 gnd.n239 585
R3136 gnd.n7449 gnd.n239 585
R3137 gnd.n6988 gnd.n6987 585
R3138 gnd.n6987 gnd.n238 585
R3139 gnd.n6989 gnd.n245 585
R3140 gnd.n7441 gnd.n245 585
R3141 gnd.n6991 gnd.n6990 585
R3142 gnd.n6990 gnd.n254 585
R3143 gnd.n6992 gnd.n253 585
R3144 gnd.n7433 gnd.n253 585
R3145 gnd.n6994 gnd.n6993 585
R3146 gnd.n6993 gnd.n263 585
R3147 gnd.n6995 gnd.n261 585
R3148 gnd.n7425 gnd.n261 585
R3149 gnd.n6997 gnd.n6996 585
R3150 gnd.n6996 gnd.n260 585
R3151 gnd.n6998 gnd.n270 585
R3152 gnd.n7417 gnd.n270 585
R3153 gnd.n7000 gnd.n6999 585
R3154 gnd.n6999 gnd.n269 585
R3155 gnd.n7001 gnd.n276 585
R3156 gnd.n7409 gnd.n276 585
R3157 gnd.n7003 gnd.n7002 585
R3158 gnd.n7002 gnd.n284 585
R3159 gnd.n7004 gnd.n283 585
R3160 gnd.n7401 gnd.n283 585
R3161 gnd.n7006 gnd.n7005 585
R3162 gnd.n7005 gnd.n293 585
R3163 gnd.n7007 gnd.n291 585
R3164 gnd.n7393 gnd.n291 585
R3165 gnd.n7009 gnd.n7008 585
R3166 gnd.n7008 gnd.n290 585
R3167 gnd.n7010 gnd.n300 585
R3168 gnd.n7385 gnd.n300 585
R3169 gnd.n7012 gnd.n7011 585
R3170 gnd.n7011 gnd.n299 585
R3171 gnd.n7013 gnd.n306 585
R3172 gnd.n7377 gnd.n306 585
R3173 gnd.n7015 gnd.n7014 585
R3174 gnd.n7014 gnd.n314 585
R3175 gnd.n7016 gnd.n313 585
R3176 gnd.n7369 gnd.n313 585
R3177 gnd.n7018 gnd.n7017 585
R3178 gnd.n7017 gnd.n323 585
R3179 gnd.n7019 gnd.n321 585
R3180 gnd.n7361 gnd.n321 585
R3181 gnd.n7021 gnd.n7020 585
R3182 gnd.n7020 gnd.n320 585
R3183 gnd.n7022 gnd.n331 585
R3184 gnd.n7353 gnd.n331 585
R3185 gnd.n7024 gnd.n7023 585
R3186 gnd.n7023 gnd.n330 585
R3187 gnd.n7025 gnd.n339 585
R3188 gnd.n7345 gnd.n339 585
R3189 gnd.n7027 gnd.n7026 585
R3190 gnd.n7026 gnd.n338 585
R3191 gnd.n7028 gnd.n346 585
R3192 gnd.n7337 gnd.n346 585
R3193 gnd.n7030 gnd.n7029 585
R3194 gnd.n7029 gnd.n356 585
R3195 gnd.n7031 gnd.n354 585
R3196 gnd.n7329 gnd.n354 585
R3197 gnd.n7033 gnd.n7032 585
R3198 gnd.n7032 gnd.n353 585
R3199 gnd.n7034 gnd.n363 585
R3200 gnd.n7321 gnd.n363 585
R3201 gnd.n7036 gnd.n7035 585
R3202 gnd.n7035 gnd.n362 585
R3203 gnd.n7037 gnd.n372 585
R3204 gnd.n7313 gnd.n372 585
R3205 gnd.n7039 gnd.n7038 585
R3206 gnd.n7040 gnd.n7039 585
R3207 gnd.n611 gnd.n379 585
R3208 gnd.n7305 gnd.n379 585
R3209 gnd.n6930 gnd.n6929 585
R3210 gnd.n6929 gnd.n6928 585
R3211 gnd.n613 gnd.n388 585
R3212 gnd.n7297 gnd.n388 585
R3213 gnd.n5884 gnd.n5883 585
R3214 gnd.n5883 gnd.n5882 585
R3215 gnd.n5885 gnd.n397 585
R3216 gnd.n7289 gnd.n397 585
R3217 gnd.n5909 gnd.n5908 585
R3218 gnd.n5908 gnd.n5907 585
R3219 gnd.n5910 gnd.n406 585
R3220 gnd.n7281 gnd.n406 585
R3221 gnd.n5913 gnd.n5912 585
R3222 gnd.n5912 gnd.n5911 585
R3223 gnd.n5914 gnd.n413 585
R3224 gnd.n7273 gnd.n413 585
R3225 gnd.n5916 gnd.n5915 585
R3226 gnd.n5917 gnd.n5916 585
R3227 gnd.n5862 gnd.n422 585
R3228 gnd.n7265 gnd.n422 585
R3229 gnd.n5872 gnd.n5871 585
R3230 gnd.n5871 gnd.n5870 585
R3231 gnd.n5869 gnd.n431 585
R3232 gnd.n7257 gnd.n431 585
R3233 gnd.n5868 gnd.n5867 585
R3234 gnd.n5867 gnd.n5866 585
R3235 gnd.n593 gnd.n440 585
R3236 gnd.n7249 gnd.n440 585
R3237 gnd.n7100 gnd.n7099 585
R3238 gnd.n7099 gnd.n7098 585
R3239 gnd.n7101 gnd.n448 585
R3240 gnd.n7241 gnd.n448 585
R3241 gnd.n7102 gnd.n590 585
R3242 gnd.n5973 gnd.n590 585
R3243 gnd.n7103 gnd.n456 585
R3244 gnd.n7233 gnd.n456 585
R3245 gnd.n5711 gnd.n1406 585
R3246 gnd.n1406 gnd.n1392 585
R3247 gnd.n5713 gnd.n5712 585
R3248 gnd.n5714 gnd.n5713 585
R3249 gnd.n1407 gnd.n1405 585
R3250 gnd.n1405 gnd.n1402 585
R3251 gnd.n5582 gnd.n5581 585
R3252 gnd.n5583 gnd.n5582 585
R3253 gnd.n5580 gnd.n1480 585
R3254 gnd.n5547 gnd.n1480 585
R3255 gnd.n5579 gnd.n5578 585
R3256 gnd.n5578 gnd.n5577 585
R3257 gnd.n1482 gnd.n1481 585
R3258 gnd.n5543 gnd.n1482 585
R3259 gnd.n5566 gnd.n5565 585
R3260 gnd.n5567 gnd.n5566 585
R3261 gnd.n5564 gnd.n1491 585
R3262 gnd.n1496 gnd.n1491 585
R3263 gnd.n5563 gnd.n5562 585
R3264 gnd.n5562 gnd.n5561 585
R3265 gnd.n1493 gnd.n1492 585
R3266 gnd.n5532 gnd.n1493 585
R3267 gnd.n5517 gnd.n5516 585
R3268 gnd.n5516 gnd.n5515 585
R3269 gnd.n5518 gnd.n1515 585
R3270 gnd.n1518 gnd.n1515 585
R3271 gnd.n5520 gnd.n5519 585
R3272 gnd.n5521 gnd.n5520 585
R3273 gnd.n1516 gnd.n1514 585
R3274 gnd.n1514 gnd.n1511 585
R3275 gnd.n5504 gnd.n5503 585
R3276 gnd.n5505 gnd.n5504 585
R3277 gnd.n5502 gnd.n1527 585
R3278 gnd.n1532 gnd.n1527 585
R3279 gnd.n5501 gnd.n5500 585
R3280 gnd.n5500 gnd.n5499 585
R3281 gnd.n1529 gnd.n1528 585
R3282 gnd.n5470 gnd.n1529 585
R3283 gnd.n5488 gnd.n5487 585
R3284 gnd.n5489 gnd.n5488 585
R3285 gnd.n5486 gnd.n1541 585
R3286 gnd.n1541 gnd.n1538 585
R3287 gnd.n5485 gnd.n5484 585
R3288 gnd.n5484 gnd.n5483 585
R3289 gnd.n1543 gnd.n1542 585
R3290 gnd.n5452 gnd.n1543 585
R3291 gnd.n5438 gnd.n5437 585
R3292 gnd.n5437 gnd.n1553 585
R3293 gnd.n5439 gnd.n1563 585
R3294 gnd.n5420 gnd.n1563 585
R3295 gnd.n5441 gnd.n5440 585
R3296 gnd.n5442 gnd.n5441 585
R3297 gnd.n5436 gnd.n1562 585
R3298 gnd.n1562 gnd.n1559 585
R3299 gnd.n5435 gnd.n5434 585
R3300 gnd.n5434 gnd.n5433 585
R3301 gnd.n1565 gnd.n1564 585
R3302 gnd.n5411 gnd.n1565 585
R3303 gnd.n5397 gnd.n5396 585
R3304 gnd.n5396 gnd.n1576 585
R3305 gnd.n5398 gnd.n1585 585
R3306 gnd.n5340 gnd.n1585 585
R3307 gnd.n5400 gnd.n5399 585
R3308 gnd.n5401 gnd.n5400 585
R3309 gnd.n5395 gnd.n1584 585
R3310 gnd.n5390 gnd.n1584 585
R3311 gnd.n5394 gnd.n5393 585
R3312 gnd.n5393 gnd.n5392 585
R3313 gnd.n1587 gnd.n1586 585
R3314 gnd.n1600 gnd.n1587 585
R3315 gnd.n5363 gnd.n5362 585
R3316 gnd.n5362 gnd.n1598 585
R3317 gnd.n5364 gnd.n1610 585
R3318 gnd.n5350 gnd.n1610 585
R3319 gnd.n5366 gnd.n5365 585
R3320 gnd.n5367 gnd.n5366 585
R3321 gnd.n5361 gnd.n1609 585
R3322 gnd.n5356 gnd.n1609 585
R3323 gnd.n5360 gnd.n5359 585
R3324 gnd.n5359 gnd.n5358 585
R3325 gnd.n1612 gnd.n1611 585
R3326 gnd.n5334 gnd.n1612 585
R3327 gnd.n5301 gnd.n5298 585
R3328 gnd.n5301 gnd.n5300 585
R3329 gnd.n5302 gnd.n5297 585
R3330 gnd.n5302 gnd.n1625 585
R3331 gnd.n5304 gnd.n5303 585
R3332 gnd.n5303 gnd.n1624 585
R3333 gnd.n5305 gnd.n1636 585
R3334 gnd.n5285 gnd.n1636 585
R3335 gnd.n5307 gnd.n5306 585
R3336 gnd.n5308 gnd.n5307 585
R3337 gnd.n5296 gnd.n1635 585
R3338 gnd.n5291 gnd.n1635 585
R3339 gnd.n5295 gnd.n5294 585
R3340 gnd.n5294 gnd.n5293 585
R3341 gnd.n1638 gnd.n1637 585
R3342 gnd.n5275 gnd.n1638 585
R3343 gnd.n5261 gnd.n5260 585
R3344 gnd.n5260 gnd.n5259 585
R3345 gnd.n5262 gnd.n1652 585
R3346 gnd.n5257 gnd.n1652 585
R3347 gnd.n5264 gnd.n5263 585
R3348 gnd.n5265 gnd.n5264 585
R3349 gnd.n1653 gnd.n1651 585
R3350 gnd.n5251 gnd.n1651 585
R3351 gnd.n5227 gnd.n1671 585
R3352 gnd.n1671 gnd.n1670 585
R3353 gnd.n5229 gnd.n5228 585
R3354 gnd.n5230 gnd.n5229 585
R3355 gnd.n5226 gnd.n1668 585
R3356 gnd.n1668 gnd.n1665 585
R3357 gnd.n5225 gnd.n5224 585
R3358 gnd.n5224 gnd.n5223 585
R3359 gnd.n1673 gnd.n1672 585
R3360 gnd.n1775 gnd.n1673 585
R3361 gnd.n5211 gnd.n5210 585
R3362 gnd.n5212 gnd.n5211 585
R3363 gnd.n5209 gnd.n1685 585
R3364 gnd.n1690 gnd.n1685 585
R3365 gnd.n5208 gnd.n5207 585
R3366 gnd.n5207 gnd.n5206 585
R3367 gnd.n1687 gnd.n1686 585
R3368 gnd.n1782 gnd.n1687 585
R3369 gnd.n5192 gnd.n5191 585
R3370 gnd.n5193 gnd.n5192 585
R3371 gnd.n5190 gnd.n1699 585
R3372 gnd.n5185 gnd.n1699 585
R3373 gnd.n5189 gnd.n5188 585
R3374 gnd.n5188 gnd.n5187 585
R3375 gnd.n1701 gnd.n1700 585
R3376 gnd.n1713 gnd.n1701 585
R3377 gnd.n5161 gnd.n1723 585
R3378 gnd.n1790 gnd.n1723 585
R3379 gnd.n5163 gnd.n5162 585
R3380 gnd.n5164 gnd.n5163 585
R3381 gnd.n5160 gnd.n1722 585
R3382 gnd.n1722 gnd.n1719 585
R3383 gnd.n5159 gnd.n5158 585
R3384 gnd.n5158 gnd.n5157 585
R3385 gnd.n1725 gnd.n1724 585
R3386 gnd.n1799 gnd.n1725 585
R3387 gnd.n5146 gnd.n5145 585
R3388 gnd.n5147 gnd.n5146 585
R3389 gnd.n5144 gnd.n1735 585
R3390 gnd.n1803 gnd.n1735 585
R3391 gnd.n5143 gnd.n5142 585
R3392 gnd.n5142 gnd.n5141 585
R3393 gnd.n1737 gnd.n1736 585
R3394 gnd.n1808 gnd.n1737 585
R3395 gnd.n5128 gnd.n5127 585
R3396 gnd.n5129 gnd.n5128 585
R3397 gnd.n5126 gnd.n1748 585
R3398 gnd.n1754 gnd.n1748 585
R3399 gnd.n5125 gnd.n5124 585
R3400 gnd.n5124 gnd.n5123 585
R3401 gnd.n1750 gnd.n1749 585
R3402 gnd.n5098 gnd.n1750 585
R3403 gnd.n5111 gnd.n5110 585
R3404 gnd.n5112 gnd.n5111 585
R3405 gnd.n5109 gnd.n1764 585
R3406 gnd.n5104 gnd.n1764 585
R3407 gnd.n5108 gnd.n5107 585
R3408 gnd.n5107 gnd.n5106 585
R3409 gnd.n1766 gnd.n1765 585
R3410 gnd.n5087 gnd.n1766 585
R3411 gnd.n4936 gnd.n4915 585
R3412 gnd.n4915 gnd.n1820 585
R3413 gnd.n5075 gnd.n5074 585
R3414 gnd.n5073 gnd.n4914 585
R3415 gnd.n5072 gnd.n4913 585
R3416 gnd.n5077 gnd.n4913 585
R3417 gnd.n5071 gnd.n5070 585
R3418 gnd.n5069 gnd.n5068 585
R3419 gnd.n5067 gnd.n5066 585
R3420 gnd.n5065 gnd.n5064 585
R3421 gnd.n5063 gnd.n5062 585
R3422 gnd.n5061 gnd.n5060 585
R3423 gnd.n5059 gnd.n5058 585
R3424 gnd.n5057 gnd.n5056 585
R3425 gnd.n5055 gnd.n5054 585
R3426 gnd.n5053 gnd.n5052 585
R3427 gnd.n5051 gnd.n5050 585
R3428 gnd.n5049 gnd.n5048 585
R3429 gnd.n5047 gnd.n5046 585
R3430 gnd.n5045 gnd.n5044 585
R3431 gnd.n5043 gnd.n5042 585
R3432 gnd.n5041 gnd.n5040 585
R3433 gnd.n5039 gnd.n5038 585
R3434 gnd.n5037 gnd.n5036 585
R3435 gnd.n5035 gnd.n5034 585
R3436 gnd.n5033 gnd.n5032 585
R3437 gnd.n5031 gnd.n5030 585
R3438 gnd.n5029 gnd.n5028 585
R3439 gnd.n5027 gnd.n5026 585
R3440 gnd.n5025 gnd.n5024 585
R3441 gnd.n5023 gnd.n5022 585
R3442 gnd.n5021 gnd.n5020 585
R3443 gnd.n5019 gnd.n5018 585
R3444 gnd.n5017 gnd.n5016 585
R3445 gnd.n5015 gnd.n5014 585
R3446 gnd.n5013 gnd.n5012 585
R3447 gnd.n5011 gnd.n5009 585
R3448 gnd.n5008 gnd.n5007 585
R3449 gnd.n5006 gnd.n5005 585
R3450 gnd.n5003 gnd.n5002 585
R3451 gnd.n5001 gnd.n5000 585
R3452 gnd.n4999 gnd.n4998 585
R3453 gnd.n4997 gnd.n4996 585
R3454 gnd.n4995 gnd.n4994 585
R3455 gnd.n4993 gnd.n4992 585
R3456 gnd.n4991 gnd.n4990 585
R3457 gnd.n4989 gnd.n4988 585
R3458 gnd.n4987 gnd.n4986 585
R3459 gnd.n4985 gnd.n4984 585
R3460 gnd.n4983 gnd.n4982 585
R3461 gnd.n4981 gnd.n4980 585
R3462 gnd.n4979 gnd.n4978 585
R3463 gnd.n4977 gnd.n4976 585
R3464 gnd.n4975 gnd.n4974 585
R3465 gnd.n4973 gnd.n4972 585
R3466 gnd.n4971 gnd.n4970 585
R3467 gnd.n4969 gnd.n4968 585
R3468 gnd.n4967 gnd.n4966 585
R3469 gnd.n4965 gnd.n4964 585
R3470 gnd.n4963 gnd.n4962 585
R3471 gnd.n4961 gnd.n4960 585
R3472 gnd.n4959 gnd.n4958 585
R3473 gnd.n4957 gnd.n4956 585
R3474 gnd.n4955 gnd.n4954 585
R3475 gnd.n4953 gnd.n4952 585
R3476 gnd.n4951 gnd.n4950 585
R3477 gnd.n4949 gnd.n4948 585
R3478 gnd.n4947 gnd.n4946 585
R3479 gnd.n5592 gnd.n5591 585
R3480 gnd.n5593 gnd.n1476 585
R3481 gnd.n5595 gnd.n5594 585
R3482 gnd.n5597 gnd.n1474 585
R3483 gnd.n5599 gnd.n5598 585
R3484 gnd.n5600 gnd.n1473 585
R3485 gnd.n5602 gnd.n5601 585
R3486 gnd.n5604 gnd.n1471 585
R3487 gnd.n5606 gnd.n5605 585
R3488 gnd.n5607 gnd.n1470 585
R3489 gnd.n5609 gnd.n5608 585
R3490 gnd.n5611 gnd.n1468 585
R3491 gnd.n5613 gnd.n5612 585
R3492 gnd.n5614 gnd.n1467 585
R3493 gnd.n5616 gnd.n5615 585
R3494 gnd.n5618 gnd.n1465 585
R3495 gnd.n5620 gnd.n5619 585
R3496 gnd.n5621 gnd.n1464 585
R3497 gnd.n5623 gnd.n5622 585
R3498 gnd.n5625 gnd.n1462 585
R3499 gnd.n5627 gnd.n5626 585
R3500 gnd.n5628 gnd.n1461 585
R3501 gnd.n5630 gnd.n5629 585
R3502 gnd.n5632 gnd.n1459 585
R3503 gnd.n5634 gnd.n5633 585
R3504 gnd.n5635 gnd.n1458 585
R3505 gnd.n5637 gnd.n5636 585
R3506 gnd.n5639 gnd.n1456 585
R3507 gnd.n5641 gnd.n5640 585
R3508 gnd.n5643 gnd.n1453 585
R3509 gnd.n5645 gnd.n5644 585
R3510 gnd.n5647 gnd.n1452 585
R3511 gnd.n5648 gnd.n1396 585
R3512 gnd.n5651 gnd.n561 585
R3513 gnd.n5653 gnd.n5652 585
R3514 gnd.n5655 gnd.n1450 585
R3515 gnd.n5657 gnd.n5656 585
R3516 gnd.n5659 gnd.n1447 585
R3517 gnd.n5661 gnd.n5660 585
R3518 gnd.n5663 gnd.n1445 585
R3519 gnd.n5665 gnd.n5664 585
R3520 gnd.n5666 gnd.n1444 585
R3521 gnd.n5668 gnd.n5667 585
R3522 gnd.n5670 gnd.n1442 585
R3523 gnd.n5672 gnd.n5671 585
R3524 gnd.n5673 gnd.n1441 585
R3525 gnd.n5675 gnd.n5674 585
R3526 gnd.n5677 gnd.n1439 585
R3527 gnd.n5679 gnd.n5678 585
R3528 gnd.n5680 gnd.n1438 585
R3529 gnd.n5682 gnd.n5681 585
R3530 gnd.n5684 gnd.n1436 585
R3531 gnd.n5686 gnd.n5685 585
R3532 gnd.n5687 gnd.n1435 585
R3533 gnd.n5689 gnd.n5688 585
R3534 gnd.n5691 gnd.n1433 585
R3535 gnd.n5693 gnd.n5692 585
R3536 gnd.n5694 gnd.n1432 585
R3537 gnd.n5696 gnd.n5695 585
R3538 gnd.n5698 gnd.n1430 585
R3539 gnd.n5700 gnd.n5699 585
R3540 gnd.n5701 gnd.n1429 585
R3541 gnd.n5703 gnd.n5702 585
R3542 gnd.n5705 gnd.n1428 585
R3543 gnd.n5706 gnd.n1427 585
R3544 gnd.n5709 gnd.n5708 585
R3545 gnd.n5590 gnd.n5588 585
R3546 gnd.n5590 gnd.n1392 585
R3547 gnd.n5587 gnd.n1403 585
R3548 gnd.n5714 gnd.n1403 585
R3549 gnd.n5586 gnd.n5585 585
R3550 gnd.n5585 gnd.n1402 585
R3551 gnd.n5584 gnd.n1477 585
R3552 gnd.n5584 gnd.n5583 585
R3553 gnd.n5539 gnd.n1478 585
R3554 gnd.n5547 gnd.n1478 585
R3555 gnd.n5540 gnd.n1483 585
R3556 gnd.n5577 gnd.n1483 585
R3557 gnd.n5542 gnd.n5541 585
R3558 gnd.n5543 gnd.n5542 585
R3559 gnd.n5538 gnd.n1489 585
R3560 gnd.n5567 gnd.n1489 585
R3561 gnd.n5537 gnd.n5536 585
R3562 gnd.n5536 gnd.n1496 585
R3563 gnd.n5535 gnd.n1495 585
R3564 gnd.n5561 gnd.n1495 585
R3565 gnd.n5534 gnd.n5533 585
R3566 gnd.n5533 gnd.n5532 585
R3567 gnd.n1505 gnd.n1504 585
R3568 gnd.n5515 gnd.n1505 585
R3569 gnd.n5460 gnd.n5459 585
R3570 gnd.n5459 gnd.n1518 585
R3571 gnd.n5461 gnd.n1512 585
R3572 gnd.n5521 gnd.n1512 585
R3573 gnd.n5463 gnd.n5462 585
R3574 gnd.n5462 gnd.n1511 585
R3575 gnd.n5464 gnd.n1526 585
R3576 gnd.n5505 gnd.n1526 585
R3577 gnd.n5466 gnd.n5465 585
R3578 gnd.n5465 gnd.n1532 585
R3579 gnd.n5467 gnd.n1530 585
R3580 gnd.n5499 gnd.n1530 585
R3581 gnd.n5469 gnd.n5468 585
R3582 gnd.n5470 gnd.n5469 585
R3583 gnd.n5458 gnd.n1539 585
R3584 gnd.n5489 gnd.n1539 585
R3585 gnd.n5457 gnd.n5456 585
R3586 gnd.n5456 gnd.n1538 585
R3587 gnd.n5455 gnd.n1545 585
R3588 gnd.n5483 gnd.n1545 585
R3589 gnd.n5454 gnd.n5453 585
R3590 gnd.n5453 gnd.n5452 585
R3591 gnd.n1552 gnd.n1551 585
R3592 gnd.n1553 gnd.n1552 585
R3593 gnd.n5419 gnd.n5418 585
R3594 gnd.n5420 gnd.n5419 585
R3595 gnd.n5417 gnd.n1560 585
R3596 gnd.n5442 gnd.n1560 585
R3597 gnd.n5416 gnd.n5415 585
R3598 gnd.n5415 gnd.n1559 585
R3599 gnd.n5414 gnd.n1567 585
R3600 gnd.n5433 gnd.n1567 585
R3601 gnd.n5413 gnd.n5412 585
R3602 gnd.n5412 gnd.n5411 585
R3603 gnd.n1574 gnd.n1573 585
R3604 gnd.n1576 gnd.n1574 585
R3605 gnd.n5342 gnd.n5341 585
R3606 gnd.n5341 gnd.n5340 585
R3607 gnd.n5343 gnd.n1582 585
R3608 gnd.n5401 gnd.n1582 585
R3609 gnd.n5344 gnd.n1590 585
R3610 gnd.n5390 gnd.n1590 585
R3611 gnd.n5345 gnd.n1589 585
R3612 gnd.n5392 gnd.n1589 585
R3613 gnd.n5347 gnd.n5346 585
R3614 gnd.n5347 gnd.n1600 585
R3615 gnd.n5348 gnd.n5338 585
R3616 gnd.n5348 gnd.n1598 585
R3617 gnd.n5352 gnd.n5351 585
R3618 gnd.n5351 gnd.n5350 585
R3619 gnd.n5353 gnd.n1607 585
R3620 gnd.n5367 gnd.n1607 585
R3621 gnd.n5355 gnd.n5354 585
R3622 gnd.n5356 gnd.n5355 585
R3623 gnd.n5337 gnd.n1614 585
R3624 gnd.n5358 gnd.n1614 585
R3625 gnd.n5336 gnd.n5335 585
R3626 gnd.n5335 gnd.n5334 585
R3627 gnd.n1616 gnd.n1615 585
R3628 gnd.n5300 gnd.n1616 585
R3629 gnd.n5281 gnd.n5280 585
R3630 gnd.n5281 gnd.n1625 585
R3631 gnd.n5282 gnd.n5279 585
R3632 gnd.n5282 gnd.n1624 585
R3633 gnd.n5287 gnd.n5286 585
R3634 gnd.n5286 gnd.n5285 585
R3635 gnd.n5288 gnd.n1634 585
R3636 gnd.n5308 gnd.n1634 585
R3637 gnd.n5290 gnd.n5289 585
R3638 gnd.n5291 gnd.n5290 585
R3639 gnd.n5278 gnd.n1640 585
R3640 gnd.n5293 gnd.n1640 585
R3641 gnd.n5277 gnd.n5276 585
R3642 gnd.n5276 gnd.n5275 585
R3643 gnd.n1643 gnd.n1642 585
R3644 gnd.n5259 gnd.n1643 585
R3645 gnd.n5256 gnd.n5255 585
R3646 gnd.n5257 gnd.n5256 585
R3647 gnd.n5254 gnd.n1650 585
R3648 gnd.n5265 gnd.n1650 585
R3649 gnd.n5253 gnd.n5252 585
R3650 gnd.n5252 gnd.n5251 585
R3651 gnd.n1656 gnd.n1655 585
R3652 gnd.n1670 gnd.n1656 585
R3653 gnd.n1770 gnd.n1666 585
R3654 gnd.n5230 gnd.n1666 585
R3655 gnd.n1772 gnd.n1771 585
R3656 gnd.n1771 gnd.n1665 585
R3657 gnd.n1773 gnd.n1675 585
R3658 gnd.n5223 gnd.n1675 585
R3659 gnd.n1777 gnd.n1776 585
R3660 gnd.n1776 gnd.n1775 585
R3661 gnd.n1778 gnd.n1683 585
R3662 gnd.n5212 gnd.n1683 585
R3663 gnd.n1780 gnd.n1779 585
R3664 gnd.n1779 gnd.n1690 585
R3665 gnd.n1781 gnd.n1689 585
R3666 gnd.n5206 gnd.n1689 585
R3667 gnd.n1784 gnd.n1783 585
R3668 gnd.n1783 gnd.n1782 585
R3669 gnd.n1785 gnd.n1697 585
R3670 gnd.n5193 gnd.n1697 585
R3671 gnd.n1786 gnd.n1705 585
R3672 gnd.n5185 gnd.n1705 585
R3673 gnd.n1787 gnd.n1704 585
R3674 gnd.n5187 gnd.n1704 585
R3675 gnd.n1789 gnd.n1788 585
R3676 gnd.n1789 gnd.n1713 585
R3677 gnd.n1792 gnd.n1791 585
R3678 gnd.n1791 gnd.n1790 585
R3679 gnd.n1793 gnd.n1720 585
R3680 gnd.n5164 gnd.n1720 585
R3681 gnd.n1795 gnd.n1794 585
R3682 gnd.n1794 gnd.n1719 585
R3683 gnd.n1796 gnd.n1727 585
R3684 gnd.n5157 gnd.n1727 585
R3685 gnd.n1801 gnd.n1800 585
R3686 gnd.n1800 gnd.n1799 585
R3687 gnd.n1802 gnd.n1733 585
R3688 gnd.n5147 gnd.n1733 585
R3689 gnd.n1805 gnd.n1804 585
R3690 gnd.n1804 gnd.n1803 585
R3691 gnd.n1806 gnd.n1739 585
R3692 gnd.n5141 gnd.n1739 585
R3693 gnd.n1810 gnd.n1809 585
R3694 gnd.n1809 gnd.n1808 585
R3695 gnd.n1811 gnd.n1746 585
R3696 gnd.n5129 gnd.n1746 585
R3697 gnd.n1813 gnd.n1812 585
R3698 gnd.n1812 gnd.n1754 585
R3699 gnd.n1814 gnd.n1752 585
R3700 gnd.n5123 gnd.n1752 585
R3701 gnd.n5100 gnd.n5099 585
R3702 gnd.n5099 gnd.n5098 585
R3703 gnd.n5101 gnd.n1763 585
R3704 gnd.n5112 gnd.n1763 585
R3705 gnd.n5103 gnd.n5102 585
R3706 gnd.n5104 gnd.n5103 585
R3707 gnd.n1769 gnd.n1768 585
R3708 gnd.n5106 gnd.n1768 585
R3709 gnd.n4943 gnd.n1821 585
R3710 gnd.n5087 gnd.n1821 585
R3711 gnd.n4945 gnd.n4944 585
R3712 gnd.n4945 gnd.n1820 585
R3713 gnd.n6919 gnd.n6918 585
R3714 gnd.n6919 gnd.n365 585
R3715 gnd.n6921 gnd.n620 585
R3716 gnd.n6921 gnd.n6920 585
R3717 gnd.n6923 gnd.n6922 585
R3718 gnd.n6922 gnd.n371 585
R3719 gnd.n6924 gnd.n615 585
R3720 gnd.n615 gnd.n381 585
R3721 gnd.n6926 gnd.n6925 585
R3722 gnd.n6927 gnd.n6926 585
R3723 gnd.n616 gnd.n614 585
R3724 gnd.n614 gnd.n390 585
R3725 gnd.n5900 gnd.n5899 585
R3726 gnd.n5900 gnd.n387 585
R3727 gnd.n5902 gnd.n5901 585
R3728 gnd.n5901 gnd.n399 585
R3729 gnd.n5903 gnd.n5887 585
R3730 gnd.n5887 gnd.n396 585
R3731 gnd.n5905 gnd.n5904 585
R3732 gnd.n5906 gnd.n5905 585
R3733 gnd.n5888 gnd.n5886 585
R3734 gnd.n5886 gnd.n405 585
R3735 gnd.n5891 gnd.n5860 585
R3736 gnd.n5860 gnd.n415 585
R3737 gnd.n5919 gnd.n5861 585
R3738 gnd.n5919 gnd.n5918 585
R3739 gnd.n5920 gnd.n5859 585
R3740 gnd.n5920 gnd.n424 585
R3741 gnd.n5922 gnd.n5921 585
R3742 gnd.n5921 gnd.n421 585
R3743 gnd.n5923 gnd.n5854 585
R3744 gnd.n5854 gnd.n433 585
R3745 gnd.n5925 gnd.n5924 585
R3746 gnd.n5925 gnd.n430 585
R3747 gnd.n5926 gnd.n5853 585
R3748 gnd.n5926 gnd.n442 585
R3749 gnd.n5928 gnd.n5927 585
R3750 gnd.n5927 gnd.n439 585
R3751 gnd.n5929 gnd.n5848 585
R3752 gnd.n5848 gnd.n450 585
R3753 gnd.n5975 gnd.n5930 585
R3754 gnd.n5975 gnd.n5974 585
R3755 gnd.n5976 gnd.n5847 585
R3756 gnd.n5976 gnd.n458 585
R3757 gnd.n5978 gnd.n5977 585
R3758 gnd.n5977 gnd.n455 585
R3759 gnd.n5979 gnd.n5840 585
R3760 gnd.n5840 gnd.n511 585
R3761 gnd.n5981 gnd.n5980 585
R3762 gnd.n5982 gnd.n5981 585
R3763 gnd.n5841 gnd.n5820 585
R3764 gnd.n5983 gnd.n5820 585
R3765 gnd.n5986 gnd.n5819 585
R3766 gnd.n5986 gnd.n5985 585
R3767 gnd.n5988 gnd.n5987 585
R3768 gnd.n5987 gnd.n1316 585
R3769 gnd.n5989 gnd.n1326 585
R3770 gnd.n1326 gnd.n1315 585
R3771 gnd.n5991 gnd.n5990 585
R3772 gnd.n5992 gnd.n5991 585
R3773 gnd.n1327 gnd.n1325 585
R3774 gnd.n1325 gnd.n1322 585
R3775 gnd.n5813 gnd.n5812 585
R3776 gnd.n5812 gnd.n5811 585
R3777 gnd.n1330 gnd.n1329 585
R3778 gnd.n1331 gnd.n1330 585
R3779 gnd.n5799 gnd.n5798 585
R3780 gnd.n5800 gnd.n5799 585
R3781 gnd.n1341 gnd.n1340 585
R3782 gnd.n1340 gnd.n1337 585
R3783 gnd.n5794 gnd.n5793 585
R3784 gnd.n5793 gnd.n5792 585
R3785 gnd.n1344 gnd.n1343 585
R3786 gnd.n1345 gnd.n1344 585
R3787 gnd.n5780 gnd.n5779 585
R3788 gnd.n5781 gnd.n5780 585
R3789 gnd.n1355 gnd.n1354 585
R3790 gnd.n1354 gnd.n1351 585
R3791 gnd.n5775 gnd.n5774 585
R3792 gnd.n5774 gnd.n5773 585
R3793 gnd.n1358 gnd.n1357 585
R3794 gnd.n1359 gnd.n1358 585
R3795 gnd.n5761 gnd.n5760 585
R3796 gnd.n5762 gnd.n5761 585
R3797 gnd.n1369 gnd.n1368 585
R3798 gnd.n1368 gnd.n1365 585
R3799 gnd.n5756 gnd.n5755 585
R3800 gnd.n5755 gnd.n5754 585
R3801 gnd.n1372 gnd.n1371 585
R3802 gnd.n1373 gnd.n1372 585
R3803 gnd.n5742 gnd.n5741 585
R3804 gnd.n5743 gnd.n5742 585
R3805 gnd.n1383 gnd.n1382 585
R3806 gnd.n1382 gnd.n1379 585
R3807 gnd.n5737 gnd.n5736 585
R3808 gnd.n5736 gnd.n5735 585
R3809 gnd.n1386 gnd.n1385 585
R3810 gnd.n1394 gnd.n1386 585
R3811 gnd.n5723 gnd.n5722 585
R3812 gnd.n5724 gnd.n5723 585
R3813 gnd.n1398 gnd.n1397 585
R3814 gnd.n1404 gnd.n1397 585
R3815 gnd.n5718 gnd.n5717 585
R3816 gnd.n5717 gnd.n5716 585
R3817 gnd.n1401 gnd.n1400 585
R3818 gnd.n1479 gnd.n1401 585
R3819 gnd.n5575 gnd.n5574 585
R3820 gnd.n5576 gnd.n5575 585
R3821 gnd.n1485 gnd.n1484 585
R3822 gnd.n1503 gnd.n1484 585
R3823 gnd.n5570 gnd.n5569 585
R3824 gnd.n5569 gnd.n5568 585
R3825 gnd.n1488 gnd.n1487 585
R3826 gnd.n1494 gnd.n1488 585
R3827 gnd.n5529 gnd.n5528 585
R3828 gnd.n5530 gnd.n5529 585
R3829 gnd.n1507 gnd.n1506 585
R3830 gnd.n1517 gnd.n1506 585
R3831 gnd.n5524 gnd.n5523 585
R3832 gnd.n5523 gnd.n5522 585
R3833 gnd.n1510 gnd.n1509 585
R3834 gnd.n1525 gnd.n1510 585
R3835 gnd.n5497 gnd.n5496 585
R3836 gnd.n5498 gnd.n5497 585
R3837 gnd.n1534 gnd.n1533 585
R3838 gnd.n5471 gnd.n1533 585
R3839 gnd.n5492 gnd.n5491 585
R3840 gnd.n5491 gnd.n5490 585
R3841 gnd.n1537 gnd.n1536 585
R3842 gnd.n5482 gnd.n1537 585
R3843 gnd.n5450 gnd.n5449 585
R3844 gnd.n5451 gnd.n5450 585
R3845 gnd.n1555 gnd.n1554 585
R3846 gnd.n5421 gnd.n1554 585
R3847 gnd.n5445 gnd.n5444 585
R3848 gnd.n5444 gnd.n5443 585
R3849 gnd.n1558 gnd.n1557 585
R3850 gnd.n5432 gnd.n1558 585
R3851 gnd.n5409 gnd.n5408 585
R3852 gnd.n5410 gnd.n5409 585
R3853 gnd.n1578 gnd.n1577 585
R3854 gnd.n5339 gnd.n1577 585
R3855 gnd.n5404 gnd.n5403 585
R3856 gnd.n5403 gnd.n5402 585
R3857 gnd.n1581 gnd.n1580 585
R3858 gnd.n5391 gnd.n1581 585
R3859 gnd.n5375 gnd.n5374 585
R3860 gnd.n5376 gnd.n5375 585
R3861 gnd.n1602 gnd.n1601 585
R3862 gnd.n5349 gnd.n1601 585
R3863 gnd.n5370 gnd.n5369 585
R3864 gnd.n5369 gnd.n5368 585
R3865 gnd.n1605 gnd.n1604 585
R3866 gnd.n5357 gnd.n1605 585
R3867 gnd.n5332 gnd.n5331 585
R3868 gnd.n5333 gnd.n5332 585
R3869 gnd.n1620 gnd.n1619 585
R3870 gnd.n5299 gnd.n1619 585
R3871 gnd.n5327 gnd.n5326 585
R3872 gnd.n5326 gnd.n5325 585
R3873 gnd.n1623 gnd.n1622 585
R3874 gnd.n5283 gnd.n1623 585
R3875 gnd.n5243 gnd.n5242 585
R3876 gnd.n5243 gnd.n1633 585
R3877 gnd.n5244 gnd.n5239 585
R3878 gnd.n5244 gnd.n1639 585
R3879 gnd.n5246 gnd.n5245 585
R3880 gnd.n5245 gnd.n1644 585
R3881 gnd.n5247 gnd.n1660 585
R3882 gnd.n1660 gnd.n1654 585
R3883 gnd.n5249 gnd.n5248 585
R3884 gnd.n5250 gnd.n5249 585
R3885 gnd.n1661 gnd.n1659 585
R3886 gnd.n1669 gnd.n1659 585
R3887 gnd.n5233 gnd.n5232 585
R3888 gnd.n5232 gnd.n5231 585
R3889 gnd.n1664 gnd.n1663 585
R3890 gnd.n1674 gnd.n1664 585
R3891 gnd.n5201 gnd.n1692 585
R3892 gnd.n1692 gnd.n1684 585
R3893 gnd.n5203 gnd.n5202 585
R3894 gnd.n5204 gnd.n5203 585
R3895 gnd.n1693 gnd.n1691 585
R3896 gnd.n1691 gnd.n1688 585
R3897 gnd.n5196 gnd.n5195 585
R3898 gnd.n5195 gnd.n5194 585
R3899 gnd.n1696 gnd.n1695 585
R3900 gnd.n5186 gnd.n1696 585
R3901 gnd.n5173 gnd.n5172 585
R3902 gnd.n5174 gnd.n5173 585
R3903 gnd.n1715 gnd.n1714 585
R3904 gnd.n1721 gnd.n1714 585
R3905 gnd.n5168 gnd.n5167 585
R3906 gnd.n5167 gnd.n5166 585
R3907 gnd.n1718 gnd.n1717 585
R3908 gnd.n1726 gnd.n1718 585
R3909 gnd.n5137 gnd.n1741 585
R3910 gnd.n1741 gnd.n1734 585
R3911 gnd.n5139 gnd.n5138 585
R3912 gnd.n5140 gnd.n5139 585
R3913 gnd.n1742 gnd.n1740 585
R3914 gnd.n1807 gnd.n1740 585
R3915 gnd.n5132 gnd.n5131 585
R3916 gnd.n5131 gnd.n5130 585
R3917 gnd.n1745 gnd.n1744 585
R3918 gnd.n5122 gnd.n1745 585
R3919 gnd.n5096 gnd.n5095 585
R3920 gnd.n5097 gnd.n5096 585
R3921 gnd.n1816 gnd.n1815 585
R3922 gnd.n1815 gnd.n1762 585
R3923 gnd.n5091 gnd.n5090 585
R3924 gnd.n5090 gnd.n1767 585
R3925 gnd.n5089 gnd.n1818 585
R3926 gnd.n5089 gnd.n5088 585
R3927 gnd.n4875 gnd.n1819 585
R3928 gnd.n4912 gnd.n1819 585
R3929 gnd.n4877 gnd.n4876 585
R3930 gnd.n4878 gnd.n4877 585
R3931 gnd.n1829 gnd.n1828 585
R3932 gnd.n1836 gnd.n1828 585
R3933 gnd.n4870 gnd.n4869 585
R3934 gnd.n4869 gnd.n4868 585
R3935 gnd.n1832 gnd.n1831 585
R3936 gnd.n4858 gnd.n1832 585
R3937 gnd.n4856 gnd.n4855 585
R3938 gnd.n4857 gnd.n4856 585
R3939 gnd.n1844 gnd.n1843 585
R3940 gnd.n1850 gnd.n1843 585
R3941 gnd.n4851 gnd.n4850 585
R3942 gnd.n4850 gnd.n4849 585
R3943 gnd.n1847 gnd.n1846 585
R3944 gnd.n4839 gnd.n1847 585
R3945 gnd.n4837 gnd.n4836 585
R3946 gnd.n4838 gnd.n4837 585
R3947 gnd.n1858 gnd.n1857 585
R3948 gnd.n1864 gnd.n1857 585
R3949 gnd.n4832 gnd.n4831 585
R3950 gnd.n4831 gnd.n4830 585
R3951 gnd.n1861 gnd.n1860 585
R3952 gnd.n4820 gnd.n1861 585
R3953 gnd.n4818 gnd.n4817 585
R3954 gnd.n4819 gnd.n4818 585
R3955 gnd.n1872 gnd.n1871 585
R3956 gnd.n1878 gnd.n1871 585
R3957 gnd.n4813 gnd.n4812 585
R3958 gnd.n4812 gnd.n4811 585
R3959 gnd.n1875 gnd.n1874 585
R3960 gnd.n4801 gnd.n1875 585
R3961 gnd.n4799 gnd.n4798 585
R3962 gnd.n4800 gnd.n4799 585
R3963 gnd.n1886 gnd.n1885 585
R3964 gnd.n1892 gnd.n1885 585
R3965 gnd.n4794 gnd.n4793 585
R3966 gnd.n4793 gnd.n4792 585
R3967 gnd.n1889 gnd.n1888 585
R3968 gnd.n4782 gnd.n1889 585
R3969 gnd.n4780 gnd.n4779 585
R3970 gnd.n4781 gnd.n4780 585
R3971 gnd.n1900 gnd.n1899 585
R3972 gnd.n4772 gnd.n1899 585
R3973 gnd.n4775 gnd.n4774 585
R3974 gnd.n4774 gnd.n4773 585
R3975 gnd.n1903 gnd.n1902 585
R3976 gnd.n4634 gnd.n1903 585
R3977 gnd.n4632 gnd.n4631 585
R3978 gnd.n4633 gnd.n4632 585
R3979 gnd.n1906 gnd.n1905 585
R3980 gnd.n1905 gnd.n1904 585
R3981 gnd.n4627 gnd.n4626 585
R3982 gnd.n4626 gnd.n1091 585
R3983 gnd.n4625 gnd.n1908 585
R3984 gnd.n4625 gnd.n1088 585
R3985 gnd.n4624 gnd.n4623 585
R3986 gnd.n4624 gnd.n1164 585
R3987 gnd.n1910 gnd.n1909 585
R3988 gnd.n1909 gnd.n1079 585
R3989 gnd.n4619 gnd.n4618 585
R3990 gnd.n4618 gnd.n1071 585
R3991 gnd.n4617 gnd.n1912 585
R3992 gnd.n4617 gnd.n1068 585
R3993 gnd.n4616 gnd.n4615 585
R3994 gnd.n4616 gnd.n1060 585
R3995 gnd.n1914 gnd.n1913 585
R3996 gnd.n1913 gnd.n1057 585
R3997 gnd.n4611 gnd.n4610 585
R3998 gnd.n4610 gnd.n1049 585
R3999 gnd.n4609 gnd.n1916 585
R4000 gnd.n4609 gnd.n1046 585
R4001 gnd.n4608 gnd.n1918 585
R4002 gnd.n4608 gnd.n4607 585
R4003 gnd.n4558 gnd.n1917 585
R4004 gnd.n1917 gnd.n1036 585
R4005 gnd.n4559 gnd.n1938 585
R4006 gnd.n1938 gnd.n1028 585
R4007 gnd.n4561 gnd.n4560 585
R4008 gnd.n4562 gnd.n4561 585
R4009 gnd.n1939 gnd.n1937 585
R4010 gnd.n1937 gnd.n1018 585
R4011 gnd.n4551 gnd.n4550 585
R4012 gnd.n4550 gnd.n1015 585
R4013 gnd.n4549 gnd.n1941 585
R4014 gnd.n4549 gnd.n1007 585
R4015 gnd.n4548 gnd.n4547 585
R4016 gnd.n4548 gnd.n1004 585
R4017 gnd.n1943 gnd.n1942 585
R4018 gnd.n3966 gnd.n1942 585
R4019 gnd.n4543 gnd.n4542 585
R4020 gnd.n4542 gnd.n993 585
R4021 gnd.n4541 gnd.n4540 585
R4022 gnd.n4541 gnd.n983 585
R4023 gnd.n4539 gnd.n980 585
R4024 gnd.n6000 gnd.n5999 585
R4025 gnd.n6001 gnd.n6000 585
R4026 gnd.n1318 gnd.n1317 585
R4027 gnd.n1324 gnd.n1317 585
R4028 gnd.n5995 gnd.n5994 585
R4029 gnd.n5994 gnd.n5993 585
R4030 gnd.n1321 gnd.n1320 585
R4031 gnd.n5810 gnd.n1321 585
R4032 gnd.n5808 gnd.n5807 585
R4033 gnd.n5809 gnd.n5808 585
R4034 gnd.n1333 gnd.n1332 585
R4035 gnd.n1339 gnd.n1332 585
R4036 gnd.n5803 gnd.n5802 585
R4037 gnd.n5802 gnd.n5801 585
R4038 gnd.n1336 gnd.n1335 585
R4039 gnd.n5791 gnd.n1336 585
R4040 gnd.n5789 gnd.n5788 585
R4041 gnd.n5790 gnd.n5789 585
R4042 gnd.n1347 gnd.n1346 585
R4043 gnd.n1353 gnd.n1346 585
R4044 gnd.n5784 gnd.n5783 585
R4045 gnd.n5783 gnd.n5782 585
R4046 gnd.n1350 gnd.n1349 585
R4047 gnd.n5772 gnd.n1350 585
R4048 gnd.n5770 gnd.n5769 585
R4049 gnd.n5771 gnd.n5770 585
R4050 gnd.n1361 gnd.n1360 585
R4051 gnd.n1367 gnd.n1360 585
R4052 gnd.n5765 gnd.n5764 585
R4053 gnd.n5764 gnd.n5763 585
R4054 gnd.n1364 gnd.n1363 585
R4055 gnd.n5753 gnd.n1364 585
R4056 gnd.n5751 gnd.n5750 585
R4057 gnd.n5752 gnd.n5751 585
R4058 gnd.n1375 gnd.n1374 585
R4059 gnd.n1381 gnd.n1374 585
R4060 gnd.n5746 gnd.n5745 585
R4061 gnd.n5745 gnd.n5744 585
R4062 gnd.n1378 gnd.n1377 585
R4063 gnd.n5734 gnd.n1378 585
R4064 gnd.n5732 gnd.n5731 585
R4065 gnd.n5733 gnd.n5732 585
R4066 gnd.n1388 gnd.n1387 585
R4067 gnd.n1395 gnd.n1387 585
R4068 gnd.n5727 gnd.n5726 585
R4069 gnd.n5726 gnd.n5725 585
R4070 gnd.n1391 gnd.n1390 585
R4071 gnd.n5715 gnd.n1391 585
R4072 gnd.n5552 gnd.n5550 585
R4073 gnd.n5550 gnd.n5549 585
R4074 gnd.n5553 gnd.n5548 585
R4075 gnd.n5548 gnd.n5547 585
R4076 gnd.n5554 gnd.n5546 585
R4077 gnd.n5546 gnd.n5545 585
R4078 gnd.n1500 gnd.n1498 585
R4079 gnd.n1498 gnd.n1490 585
R4080 gnd.n5559 gnd.n5558 585
R4081 gnd.n5560 gnd.n5559 585
R4082 gnd.n1499 gnd.n1497 585
R4083 gnd.n5531 gnd.n1497 585
R4084 gnd.n5513 gnd.n5512 585
R4085 gnd.n5514 gnd.n5513 585
R4086 gnd.n1521 gnd.n1520 585
R4087 gnd.n1520 gnd.n1513 585
R4088 gnd.n5508 gnd.n5507 585
R4089 gnd.n5507 gnd.n5506 585
R4090 gnd.n1524 gnd.n1523 585
R4091 gnd.n1531 gnd.n1524 585
R4092 gnd.n5475 gnd.n5474 585
R4093 gnd.n5474 gnd.n5473 585
R4094 gnd.n1549 gnd.n1547 585
R4095 gnd.n1547 gnd.n1540 585
R4096 gnd.n5480 gnd.n5479 585
R4097 gnd.n5481 gnd.n5480 585
R4098 gnd.n1548 gnd.n1546 585
R4099 gnd.n1546 gnd.n1544 585
R4100 gnd.n5425 gnd.n5424 585
R4101 gnd.n5424 gnd.n5423 585
R4102 gnd.n1571 gnd.n1569 585
R4103 gnd.n1569 gnd.n1561 585
R4104 gnd.n5430 gnd.n5429 585
R4105 gnd.n5431 gnd.n5430 585
R4106 gnd.n1570 gnd.n1568 585
R4107 gnd.n1568 gnd.n1566 585
R4108 gnd.n5383 gnd.n5382 585
R4109 gnd.n5382 gnd.n1576 585
R4110 gnd.n1594 gnd.n1592 585
R4111 gnd.n1592 gnd.n1583 585
R4112 gnd.n5388 gnd.n5387 585
R4113 gnd.n5389 gnd.n5388 585
R4114 gnd.n1593 gnd.n1591 585
R4115 gnd.n1591 gnd.n1588 585
R4116 gnd.n5379 gnd.n5378 585
R4117 gnd.n5378 gnd.n5377 585
R4118 gnd.n1597 gnd.n1596 585
R4119 gnd.n1608 gnd.n1597 585
R4120 gnd.n5317 gnd.n5316 585
R4121 gnd.n5316 gnd.n1606 585
R4122 gnd.n5318 gnd.n5315 585
R4123 gnd.n5315 gnd.n1613 585
R4124 gnd.n1629 gnd.n1627 585
R4125 gnd.n1627 gnd.n1618 585
R4126 gnd.n5323 gnd.n5322 585
R4127 gnd.n5324 gnd.n5323 585
R4128 gnd.n1628 gnd.n1626 585
R4129 gnd.n5284 gnd.n1626 585
R4130 gnd.n5311 gnd.n5310 585
R4131 gnd.n5310 gnd.n5309 585
R4132 gnd.n1632 gnd.n1631 585
R4133 gnd.n5292 gnd.n1632 585
R4134 gnd.n5273 gnd.n5272 585
R4135 gnd.n5274 gnd.n5273 585
R4136 gnd.n1646 gnd.n1645 585
R4137 gnd.n5258 gnd.n1645 585
R4138 gnd.n5268 gnd.n5267 585
R4139 gnd.n5267 gnd.n5266 585
R4140 gnd.n1649 gnd.n1648 585
R4141 gnd.n1658 gnd.n1649 585
R4142 gnd.n1678 gnd.n1667 585
R4143 gnd.n5230 gnd.n1667 585
R4144 gnd.n5221 gnd.n5220 585
R4145 gnd.n5222 gnd.n5221 585
R4146 gnd.n1677 gnd.n1676 585
R4147 gnd.n1774 gnd.n1676 585
R4148 gnd.n5215 gnd.n5214 585
R4149 gnd.n5214 gnd.n5213 585
R4150 gnd.n1681 gnd.n1680 585
R4151 gnd.n5205 gnd.n1681 585
R4152 gnd.n1709 gnd.n1707 585
R4153 gnd.n1707 gnd.n1698 585
R4154 gnd.n5183 gnd.n5182 585
R4155 gnd.n5184 gnd.n5183 585
R4156 gnd.n1708 gnd.n1706 585
R4157 gnd.n1706 gnd.n1703 585
R4158 gnd.n5177 gnd.n5176 585
R4159 gnd.n5176 gnd.n5175 585
R4160 gnd.n1712 gnd.n1711 585
R4161 gnd.n5165 gnd.n1712 585
R4162 gnd.n5155 gnd.n5154 585
R4163 gnd.n5156 gnd.n5155 585
R4164 gnd.n1729 gnd.n1728 585
R4165 gnd.n1798 gnd.n1728 585
R4166 gnd.n5150 gnd.n5149 585
R4167 gnd.n5149 gnd.n5148 585
R4168 gnd.n1732 gnd.n1731 585
R4169 gnd.n1738 gnd.n1732 585
R4170 gnd.n1758 gnd.n1756 585
R4171 gnd.n1756 gnd.n1747 585
R4172 gnd.n5120 gnd.n5119 585
R4173 gnd.n5121 gnd.n5120 585
R4174 gnd.n1757 gnd.n1755 585
R4175 gnd.n1755 gnd.n1751 585
R4176 gnd.n5114 gnd.n5113 585
R4177 gnd.n5113 gnd.n5112 585
R4178 gnd.n1761 gnd.n1760 585
R4179 gnd.n5105 gnd.n1761 585
R4180 gnd.n5085 gnd.n5084 585
R4181 gnd.n5086 gnd.n5085 585
R4182 gnd.n1824 gnd.n1823 585
R4183 gnd.n4911 gnd.n1823 585
R4184 gnd.n5080 gnd.n5079 585
R4185 gnd.n5079 gnd.n5078 585
R4186 gnd.n1827 gnd.n1826 585
R4187 gnd.n1835 gnd.n1827 585
R4188 gnd.n4866 gnd.n4865 585
R4189 gnd.n4867 gnd.n4866 585
R4190 gnd.n1838 gnd.n1837 585
R4191 gnd.n1837 gnd.n1833 585
R4192 gnd.n4861 gnd.n4860 585
R4193 gnd.n4860 gnd.n4859 585
R4194 gnd.n1841 gnd.n1840 585
R4195 gnd.n1842 gnd.n1841 585
R4196 gnd.n4847 gnd.n4846 585
R4197 gnd.n4848 gnd.n4847 585
R4198 gnd.n1852 gnd.n1851 585
R4199 gnd.n1851 gnd.n1848 585
R4200 gnd.n4842 gnd.n4841 585
R4201 gnd.n4841 gnd.n4840 585
R4202 gnd.n1855 gnd.n1854 585
R4203 gnd.n1856 gnd.n1855 585
R4204 gnd.n4828 gnd.n4827 585
R4205 gnd.n4829 gnd.n4828 585
R4206 gnd.n1866 gnd.n1865 585
R4207 gnd.n1865 gnd.n1862 585
R4208 gnd.n4823 gnd.n4822 585
R4209 gnd.n4822 gnd.n4821 585
R4210 gnd.n1869 gnd.n1868 585
R4211 gnd.n1870 gnd.n1869 585
R4212 gnd.n4809 gnd.n4808 585
R4213 gnd.n4810 gnd.n4809 585
R4214 gnd.n1880 gnd.n1879 585
R4215 gnd.n1879 gnd.n1876 585
R4216 gnd.n4804 gnd.n4803 585
R4217 gnd.n4803 gnd.n4802 585
R4218 gnd.n1883 gnd.n1882 585
R4219 gnd.n1884 gnd.n1883 585
R4220 gnd.n4790 gnd.n4789 585
R4221 gnd.n4791 gnd.n4790 585
R4222 gnd.n1894 gnd.n1893 585
R4223 gnd.n1893 gnd.n1890 585
R4224 gnd.n4785 gnd.n4784 585
R4225 gnd.n4784 gnd.n4783 585
R4226 gnd.n1897 gnd.n1896 585
R4227 gnd.n1898 gnd.n1897 585
R4228 gnd.n4769 gnd.n4768 585
R4229 gnd.n4767 gnd.n4651 585
R4230 gnd.n4653 gnd.n4650 585
R4231 gnd.n4771 gnd.n4650 585
R4232 gnd.n4760 gnd.n4670 585
R4233 gnd.n4759 gnd.n4671 585
R4234 gnd.n4673 gnd.n4672 585
R4235 gnd.n4752 gnd.n4681 585
R4236 gnd.n4751 gnd.n4682 585
R4237 gnd.n4692 gnd.n4683 585
R4238 gnd.n4744 gnd.n4693 585
R4239 gnd.n4743 gnd.n4694 585
R4240 gnd.n4696 gnd.n4695 585
R4241 gnd.n4736 gnd.n4704 585
R4242 gnd.n4735 gnd.n4705 585
R4243 gnd.n4717 gnd.n4706 585
R4244 gnd.n4728 gnd.n4718 585
R4245 gnd.n4727 gnd.n4720 585
R4246 gnd.n4719 gnd.n1170 585
R4247 gnd.n6171 gnd.n1171 585
R4248 gnd.n6170 gnd.n1172 585
R4249 gnd.n6169 gnd.n1173 585
R4250 gnd.n4644 gnd.n1174 585
R4251 gnd.n6165 gnd.n1176 585
R4252 gnd.n6164 gnd.n1177 585
R4253 gnd.n6163 gnd.n1178 585
R4254 gnd.n6160 gnd.n1183 585
R4255 gnd.n6159 gnd.n1184 585
R4256 gnd.n6158 gnd.n1185 585
R4257 gnd.n4648 gnd.n1186 585
R4258 gnd.n6003 gnd.n6002 585
R4259 gnd.n6002 gnd.n6001 585
R4260 gnd.n6004 gnd.n1313 585
R4261 gnd.n1324 gnd.n1313 585
R4262 gnd.n1323 gnd.n1311 585
R4263 gnd.n5993 gnd.n1323 585
R4264 gnd.n6008 gnd.n1310 585
R4265 gnd.n5810 gnd.n1310 585
R4266 gnd.n6009 gnd.n1309 585
R4267 gnd.n5809 gnd.n1309 585
R4268 gnd.n6010 gnd.n1308 585
R4269 gnd.n1339 gnd.n1308 585
R4270 gnd.n1338 gnd.n1306 585
R4271 gnd.n5801 gnd.n1338 585
R4272 gnd.n6014 gnd.n1305 585
R4273 gnd.n5791 gnd.n1305 585
R4274 gnd.n6015 gnd.n1304 585
R4275 gnd.n5790 gnd.n1304 585
R4276 gnd.n6016 gnd.n1303 585
R4277 gnd.n1353 gnd.n1303 585
R4278 gnd.n1352 gnd.n1301 585
R4279 gnd.n5782 gnd.n1352 585
R4280 gnd.n6020 gnd.n1300 585
R4281 gnd.n5772 gnd.n1300 585
R4282 gnd.n6021 gnd.n1299 585
R4283 gnd.n5771 gnd.n1299 585
R4284 gnd.n6022 gnd.n1298 585
R4285 gnd.n1367 gnd.n1298 585
R4286 gnd.n1366 gnd.n1296 585
R4287 gnd.n5763 gnd.n1366 585
R4288 gnd.n6026 gnd.n1295 585
R4289 gnd.n5753 gnd.n1295 585
R4290 gnd.n6027 gnd.n1294 585
R4291 gnd.n5752 gnd.n1294 585
R4292 gnd.n6028 gnd.n1293 585
R4293 gnd.n1381 gnd.n1293 585
R4294 gnd.n1380 gnd.n1291 585
R4295 gnd.n5744 gnd.n1380 585
R4296 gnd.n6032 gnd.n1290 585
R4297 gnd.n5734 gnd.n1290 585
R4298 gnd.n6033 gnd.n1289 585
R4299 gnd.n5733 gnd.n1289 585
R4300 gnd.n6034 gnd.n1288 585
R4301 gnd.n1395 gnd.n1288 585
R4302 gnd.n1393 gnd.n1286 585
R4303 gnd.n5725 gnd.n1393 585
R4304 gnd.n6038 gnd.n1285 585
R4305 gnd.n5715 gnd.n1285 585
R4306 gnd.n6039 gnd.n1284 585
R4307 gnd.n5549 gnd.n1284 585
R4308 gnd.n6040 gnd.n1283 585
R4309 gnd.n5547 gnd.n1283 585
R4310 gnd.n5544 gnd.n1281 585
R4311 gnd.n5545 gnd.n5544 585
R4312 gnd.n6044 gnd.n1280 585
R4313 gnd.n1490 gnd.n1280 585
R4314 gnd.n6045 gnd.n1279 585
R4315 gnd.n5560 gnd.n1279 585
R4316 gnd.n6046 gnd.n1278 585
R4317 gnd.n5531 gnd.n1278 585
R4318 gnd.n1519 gnd.n1276 585
R4319 gnd.n5514 gnd.n1519 585
R4320 gnd.n6050 gnd.n1275 585
R4321 gnd.n1513 gnd.n1275 585
R4322 gnd.n6051 gnd.n1274 585
R4323 gnd.n5506 gnd.n1274 585
R4324 gnd.n6052 gnd.n1273 585
R4325 gnd.n1531 gnd.n1273 585
R4326 gnd.n5472 gnd.n1271 585
R4327 gnd.n5473 gnd.n5472 585
R4328 gnd.n6056 gnd.n1270 585
R4329 gnd.n1540 gnd.n1270 585
R4330 gnd.n6057 gnd.n1269 585
R4331 gnd.n5481 gnd.n1269 585
R4332 gnd.n6058 gnd.n1268 585
R4333 gnd.n1544 gnd.n1268 585
R4334 gnd.n5422 gnd.n1266 585
R4335 gnd.n5423 gnd.n5422 585
R4336 gnd.n6062 gnd.n1265 585
R4337 gnd.n1561 gnd.n1265 585
R4338 gnd.n6063 gnd.n1264 585
R4339 gnd.n5431 gnd.n1264 585
R4340 gnd.n6064 gnd.n1263 585
R4341 gnd.n1566 gnd.n1263 585
R4342 gnd.n1575 gnd.n1261 585
R4343 gnd.n1576 gnd.n1575 585
R4344 gnd.n6068 gnd.n1260 585
R4345 gnd.n1583 gnd.n1260 585
R4346 gnd.n6069 gnd.n1259 585
R4347 gnd.n5389 gnd.n1259 585
R4348 gnd.n6070 gnd.n1258 585
R4349 gnd.n1588 gnd.n1258 585
R4350 gnd.n1599 gnd.n1256 585
R4351 gnd.n5377 gnd.n1599 585
R4352 gnd.n6074 gnd.n1255 585
R4353 gnd.n1608 gnd.n1255 585
R4354 gnd.n6075 gnd.n1254 585
R4355 gnd.n1606 gnd.n1254 585
R4356 gnd.n6076 gnd.n1253 585
R4357 gnd.n1613 gnd.n1253 585
R4358 gnd.n1617 gnd.n1251 585
R4359 gnd.n1618 gnd.n1617 585
R4360 gnd.n6080 gnd.n1250 585
R4361 gnd.n5324 gnd.n1250 585
R4362 gnd.n6081 gnd.n1249 585
R4363 gnd.n5284 gnd.n1249 585
R4364 gnd.n6082 gnd.n1248 585
R4365 gnd.n5309 gnd.n1248 585
R4366 gnd.n1641 gnd.n1246 585
R4367 gnd.n5292 gnd.n1641 585
R4368 gnd.n6086 gnd.n1245 585
R4369 gnd.n5274 gnd.n1245 585
R4370 gnd.n6087 gnd.n1244 585
R4371 gnd.n5258 gnd.n1244 585
R4372 gnd.n6088 gnd.n1243 585
R4373 gnd.n5266 gnd.n1243 585
R4374 gnd.n1657 gnd.n1241 585
R4375 gnd.n1658 gnd.n1657 585
R4376 gnd.n6092 gnd.n1240 585
R4377 gnd.n5230 gnd.n1240 585
R4378 gnd.n6093 gnd.n1239 585
R4379 gnd.n5222 gnd.n1239 585
R4380 gnd.n6094 gnd.n1238 585
R4381 gnd.n1774 gnd.n1238 585
R4382 gnd.n1682 gnd.n1236 585
R4383 gnd.n5213 gnd.n1682 585
R4384 gnd.n6098 gnd.n1235 585
R4385 gnd.n5205 gnd.n1235 585
R4386 gnd.n6099 gnd.n1234 585
R4387 gnd.n1698 gnd.n1234 585
R4388 gnd.n6100 gnd.n1233 585
R4389 gnd.n5184 gnd.n1233 585
R4390 gnd.n1702 gnd.n1231 585
R4391 gnd.n1703 gnd.n1702 585
R4392 gnd.n6104 gnd.n1230 585
R4393 gnd.n5175 gnd.n1230 585
R4394 gnd.n6105 gnd.n1229 585
R4395 gnd.n5165 gnd.n1229 585
R4396 gnd.n6106 gnd.n1228 585
R4397 gnd.n5156 gnd.n1228 585
R4398 gnd.n1797 gnd.n1226 585
R4399 gnd.n1798 gnd.n1797 585
R4400 gnd.n6110 gnd.n1225 585
R4401 gnd.n5148 gnd.n1225 585
R4402 gnd.n6111 gnd.n1224 585
R4403 gnd.n1738 gnd.n1224 585
R4404 gnd.n6112 gnd.n1223 585
R4405 gnd.n1747 gnd.n1223 585
R4406 gnd.n1753 gnd.n1221 585
R4407 gnd.n5121 gnd.n1753 585
R4408 gnd.n6116 gnd.n1220 585
R4409 gnd.n1751 gnd.n1220 585
R4410 gnd.n6117 gnd.n1219 585
R4411 gnd.n5112 gnd.n1219 585
R4412 gnd.n6118 gnd.n1218 585
R4413 gnd.n5105 gnd.n1218 585
R4414 gnd.n1822 gnd.n1216 585
R4415 gnd.n5086 gnd.n1822 585
R4416 gnd.n6122 gnd.n1215 585
R4417 gnd.n4911 gnd.n1215 585
R4418 gnd.n6123 gnd.n1214 585
R4419 gnd.n5078 gnd.n1214 585
R4420 gnd.n6124 gnd.n1213 585
R4421 gnd.n1835 gnd.n1213 585
R4422 gnd.n1834 gnd.n1211 585
R4423 gnd.n4867 gnd.n1834 585
R4424 gnd.n6128 gnd.n1210 585
R4425 gnd.n1833 gnd.n1210 585
R4426 gnd.n6129 gnd.n1209 585
R4427 gnd.n4859 gnd.n1209 585
R4428 gnd.n6130 gnd.n1208 585
R4429 gnd.n1842 gnd.n1208 585
R4430 gnd.n1849 gnd.n1206 585
R4431 gnd.n4848 gnd.n1849 585
R4432 gnd.n6134 gnd.n1205 585
R4433 gnd.n1848 gnd.n1205 585
R4434 gnd.n6135 gnd.n1204 585
R4435 gnd.n4840 gnd.n1204 585
R4436 gnd.n6136 gnd.n1203 585
R4437 gnd.n1856 gnd.n1203 585
R4438 gnd.n1863 gnd.n1201 585
R4439 gnd.n4829 gnd.n1863 585
R4440 gnd.n6140 gnd.n1200 585
R4441 gnd.n1862 gnd.n1200 585
R4442 gnd.n6141 gnd.n1199 585
R4443 gnd.n4821 gnd.n1199 585
R4444 gnd.n6142 gnd.n1198 585
R4445 gnd.n1870 gnd.n1198 585
R4446 gnd.n1877 gnd.n1196 585
R4447 gnd.n4810 gnd.n1877 585
R4448 gnd.n6146 gnd.n1195 585
R4449 gnd.n1876 gnd.n1195 585
R4450 gnd.n6147 gnd.n1194 585
R4451 gnd.n4802 gnd.n1194 585
R4452 gnd.n6148 gnd.n1193 585
R4453 gnd.n1884 gnd.n1193 585
R4454 gnd.n1891 gnd.n1191 585
R4455 gnd.n4791 gnd.n1891 585
R4456 gnd.n6152 gnd.n1190 585
R4457 gnd.n1890 gnd.n1190 585
R4458 gnd.n6153 gnd.n1189 585
R4459 gnd.n4783 gnd.n1189 585
R4460 gnd.n6154 gnd.n1188 585
R4461 gnd.n1898 gnd.n1188 585
R4462 gnd.n5950 gnd.n1314 585
R4463 gnd.n5984 gnd.n1314 585
R4464 gnd.n5951 gnd.n5949 585
R4465 gnd.n5947 gnd.n5946 585
R4466 gnd.n5955 gnd.n5945 585
R4467 gnd.n5959 gnd.n5944 585
R4468 gnd.n5960 gnd.n5943 585
R4469 gnd.n5941 gnd.n5940 585
R4470 gnd.n5964 gnd.n5939 585
R4471 gnd.n5965 gnd.n5938 585
R4472 gnd.n5966 gnd.n5937 585
R4473 gnd.n5936 gnd.n5935 585
R4474 gnd.n5934 gnd.n508 585
R4475 gnd.n7183 gnd.n507 585
R4476 gnd.n7184 gnd.n506 585
R4477 gnd.n5832 gnd.n498 585
R4478 gnd.n7191 gnd.n497 585
R4479 gnd.n7192 gnd.n496 585
R4480 gnd.n5829 gnd.n490 585
R4481 gnd.n7199 gnd.n489 585
R4482 gnd.n7200 gnd.n488 585
R4483 gnd.n5827 gnd.n482 585
R4484 gnd.n7207 gnd.n481 585
R4485 gnd.n7208 gnd.n480 585
R4486 gnd.n5824 gnd.n474 585
R4487 gnd.n7215 gnd.n473 585
R4488 gnd.n7216 gnd.n472 585
R4489 gnd.n5822 gnd.n466 585
R4490 gnd.n7223 gnd.n465 585
R4491 gnd.n7224 gnd.n464 585
R4492 gnd.n3631 gnd.n3630 537.605
R4493 gnd.n5708 gnd.n1406 473.281
R4494 gnd.n5591 gnd.n5590 473.281
R4495 gnd.n4946 gnd.n4945 473.281
R4496 gnd.n5075 gnd.n4915 473.281
R4497 gnd.n4941 gnd.t303 443.966
R4498 gnd.n1454 gnd.t256 443.966
R4499 gnd.n4938 gnd.t249 443.966
R4500 gnd.n1448 gnd.t293 443.966
R4501 gnd.n1179 gnd.t270 371.625
R4502 gnd.n564 gnd.t267 371.625
R4503 gnd.n586 gnd.t245 371.625
R4504 gnd.n201 gnd.t313 371.625
R4505 gnd.n7592 gnd.t227 371.625
R4506 gnd.n122 gnd.t284 371.625
R4507 gnd.n502 gnd.t296 371.625
R4508 gnd.n4713 gnd.t320 371.625
R4509 gnd.n1157 gnd.t323 371.625
R4510 gnd.n1120 gnd.t241 371.625
R4511 gnd.n3756 gnd.t329 371.625
R4512 gnd.n3732 gnd.t309 371.625
R4513 gnd.n3659 gnd.t326 371.625
R4514 gnd.n5956 gnd.t237 371.625
R4515 gnd.n2650 gnd.t316 323.425
R4516 gnd.n2196 gnd.t260 323.425
R4517 gnd.n3498 gnd.n3472 289.615
R4518 gnd.n3466 gnd.n3440 289.615
R4519 gnd.n3434 gnd.n3408 289.615
R4520 gnd.n3403 gnd.n3377 289.615
R4521 gnd.n3371 gnd.n3345 289.615
R4522 gnd.n3339 gnd.n3313 289.615
R4523 gnd.n3307 gnd.n3281 289.615
R4524 gnd.n3276 gnd.n3250 289.615
R4525 gnd.n2724 gnd.t299 279.217
R4526 gnd.n2222 gnd.t277 279.217
R4527 gnd.n4922 gnd.t236 260.649
R4528 gnd.n1419 gnd.t276 260.649
R4529 gnd.n5077 gnd.n5076 256.663
R4530 gnd.n5077 gnd.n4879 256.663
R4531 gnd.n5077 gnd.n4880 256.663
R4532 gnd.n5077 gnd.n4881 256.663
R4533 gnd.n5077 gnd.n4882 256.663
R4534 gnd.n5077 gnd.n4883 256.663
R4535 gnd.n5077 gnd.n4884 256.663
R4536 gnd.n5077 gnd.n4885 256.663
R4537 gnd.n5077 gnd.n4886 256.663
R4538 gnd.n5077 gnd.n4887 256.663
R4539 gnd.n5077 gnd.n4888 256.663
R4540 gnd.n5077 gnd.n4889 256.663
R4541 gnd.n5077 gnd.n4890 256.663
R4542 gnd.n5077 gnd.n4891 256.663
R4543 gnd.n5077 gnd.n4892 256.663
R4544 gnd.n5077 gnd.n4893 256.663
R4545 gnd.n5013 gnd.n5010 256.663
R4546 gnd.n5077 gnd.n4894 256.663
R4547 gnd.n5077 gnd.n4895 256.663
R4548 gnd.n5077 gnd.n4896 256.663
R4549 gnd.n5077 gnd.n4897 256.663
R4550 gnd.n5077 gnd.n4898 256.663
R4551 gnd.n5077 gnd.n4899 256.663
R4552 gnd.n5077 gnd.n4900 256.663
R4553 gnd.n5077 gnd.n4901 256.663
R4554 gnd.n5077 gnd.n4902 256.663
R4555 gnd.n5077 gnd.n4903 256.663
R4556 gnd.n5077 gnd.n4904 256.663
R4557 gnd.n5077 gnd.n4905 256.663
R4558 gnd.n5077 gnd.n4906 256.663
R4559 gnd.n5077 gnd.n4907 256.663
R4560 gnd.n5077 gnd.n4908 256.663
R4561 gnd.n5077 gnd.n4909 256.663
R4562 gnd.n5077 gnd.n4910 256.663
R4563 gnd.n5589 gnd.n1396 256.663
R4564 gnd.n5596 gnd.n1396 256.663
R4565 gnd.n1475 gnd.n1396 256.663
R4566 gnd.n5603 gnd.n1396 256.663
R4567 gnd.n1472 gnd.n1396 256.663
R4568 gnd.n5610 gnd.n1396 256.663
R4569 gnd.n1469 gnd.n1396 256.663
R4570 gnd.n5617 gnd.n1396 256.663
R4571 gnd.n1466 gnd.n1396 256.663
R4572 gnd.n5624 gnd.n1396 256.663
R4573 gnd.n1463 gnd.n1396 256.663
R4574 gnd.n5631 gnd.n1396 256.663
R4575 gnd.n1460 gnd.n1396 256.663
R4576 gnd.n5638 gnd.n1396 256.663
R4577 gnd.n1457 gnd.n1396 256.663
R4578 gnd.n5646 gnd.n1396 256.663
R4579 gnd.n5649 gnd.n561 256.663
R4580 gnd.n5650 gnd.n1396 256.663
R4581 gnd.n5654 gnd.n1396 256.663
R4582 gnd.n1451 gnd.n1396 256.663
R4583 gnd.n5662 gnd.n1396 256.663
R4584 gnd.n1446 gnd.n1396 256.663
R4585 gnd.n5669 gnd.n1396 256.663
R4586 gnd.n1443 gnd.n1396 256.663
R4587 gnd.n5676 gnd.n1396 256.663
R4588 gnd.n1440 gnd.n1396 256.663
R4589 gnd.n5683 gnd.n1396 256.663
R4590 gnd.n1437 gnd.n1396 256.663
R4591 gnd.n5690 gnd.n1396 256.663
R4592 gnd.n1434 gnd.n1396 256.663
R4593 gnd.n5697 gnd.n1396 256.663
R4594 gnd.n1431 gnd.n1396 256.663
R4595 gnd.n5704 gnd.n1396 256.663
R4596 gnd.n5707 gnd.n1396 256.663
R4597 gnd.n4095 gnd.n3631 242.672
R4598 gnd.n4093 gnd.n3631 242.672
R4599 gnd.n4087 gnd.n3631 242.672
R4600 gnd.n4085 gnd.n3631 242.672
R4601 gnd.n4079 gnd.n3631 242.672
R4602 gnd.n4077 gnd.n3631 242.672
R4603 gnd.n4071 gnd.n3631 242.672
R4604 gnd.n4069 gnd.n3631 242.672
R4605 gnd.n4059 gnd.n3631 242.672
R4606 gnd.n2778 gnd.n2777 242.672
R4607 gnd.n2778 gnd.n2688 242.672
R4608 gnd.n2778 gnd.n2689 242.672
R4609 gnd.n2778 gnd.n2690 242.672
R4610 gnd.n2778 gnd.n2691 242.672
R4611 gnd.n2778 gnd.n2692 242.672
R4612 gnd.n2778 gnd.n2693 242.672
R4613 gnd.n2778 gnd.n2694 242.672
R4614 gnd.n2778 gnd.n2695 242.672
R4615 gnd.n2778 gnd.n2696 242.672
R4616 gnd.n2778 gnd.n2697 242.672
R4617 gnd.n2778 gnd.n2698 242.672
R4618 gnd.n2779 gnd.n2778 242.672
R4619 gnd.n3630 gnd.n2171 242.672
R4620 gnd.n3630 gnd.n2170 242.672
R4621 gnd.n3630 gnd.n2169 242.672
R4622 gnd.n3630 gnd.n2168 242.672
R4623 gnd.n3630 gnd.n2167 242.672
R4624 gnd.n3630 gnd.n2166 242.672
R4625 gnd.n3630 gnd.n2165 242.672
R4626 gnd.n3630 gnd.n2164 242.672
R4627 gnd.n3630 gnd.n2163 242.672
R4628 gnd.n3630 gnd.n2162 242.672
R4629 gnd.n3630 gnd.n2161 242.672
R4630 gnd.n3630 gnd.n2160 242.672
R4631 gnd.n3630 gnd.n2159 242.672
R4632 gnd.n2862 gnd.n2861 242.672
R4633 gnd.n2861 gnd.n2600 242.672
R4634 gnd.n2861 gnd.n2601 242.672
R4635 gnd.n2861 gnd.n2602 242.672
R4636 gnd.n2861 gnd.n2603 242.672
R4637 gnd.n2861 gnd.n2604 242.672
R4638 gnd.n2861 gnd.n2605 242.672
R4639 gnd.n2861 gnd.n2606 242.672
R4640 gnd.n3630 gnd.n2172 242.672
R4641 gnd.n3630 gnd.n2173 242.672
R4642 gnd.n3630 gnd.n2174 242.672
R4643 gnd.n3630 gnd.n2175 242.672
R4644 gnd.n3630 gnd.n2176 242.672
R4645 gnd.n3630 gnd.n2177 242.672
R4646 gnd.n3630 gnd.n2178 242.672
R4647 gnd.n3630 gnd.n2179 242.672
R4648 gnd.n3774 gnd.n3631 242.672
R4649 gnd.n3782 gnd.n3631 242.672
R4650 gnd.n3784 gnd.n3631 242.672
R4651 gnd.n3792 gnd.n3631 242.672
R4652 gnd.n3794 gnd.n3631 242.672
R4653 gnd.n3802 gnd.n3631 242.672
R4654 gnd.n3804 gnd.n3631 242.672
R4655 gnd.n3812 gnd.n3631 242.672
R4656 gnd.n3814 gnd.n3631 242.672
R4657 gnd.n3822 gnd.n3631 242.672
R4658 gnd.n3824 gnd.n3631 242.672
R4659 gnd.n3832 gnd.n3631 242.672
R4660 gnd.n3834 gnd.n3631 242.672
R4661 gnd.n3842 gnd.n3631 242.672
R4662 gnd.n3844 gnd.n3631 242.672
R4663 gnd.n3852 gnd.n3631 242.672
R4664 gnd.n3854 gnd.n3631 242.672
R4665 gnd.n3863 gnd.n3631 242.672
R4666 gnd.n3866 gnd.n3631 242.672
R4667 gnd.n4533 gnd.n4532 242.672
R4668 gnd.n4533 gnd.n1948 242.672
R4669 gnd.n4533 gnd.n1949 242.672
R4670 gnd.n4533 gnd.n1950 242.672
R4671 gnd.n4533 gnd.n1951 242.672
R4672 gnd.n4533 gnd.n1952 242.672
R4673 gnd.n4533 gnd.n1953 242.672
R4674 gnd.n4533 gnd.n1954 242.672
R4675 gnd.n4533 gnd.n1955 242.672
R4676 gnd.n4533 gnd.n1956 242.672
R4677 gnd.n4533 gnd.n1957 242.672
R4678 gnd.n4533 gnd.n1958 242.672
R4679 gnd.n4533 gnd.n1959 242.672
R4680 gnd.n4533 gnd.n1960 242.672
R4681 gnd.n4533 gnd.n1961 242.672
R4682 gnd.n4533 gnd.n1962 242.672
R4683 gnd.n4533 gnd.n1963 242.672
R4684 gnd.n4533 gnd.n1964 242.672
R4685 gnd.n4533 gnd.n1965 242.672
R4686 gnd.n4533 gnd.n1966 242.672
R4687 gnd.n4533 gnd.n1967 242.672
R4688 gnd.n4533 gnd.n1968 242.672
R4689 gnd.n4533 gnd.n1969 242.672
R4690 gnd.n4533 gnd.n1970 242.672
R4691 gnd.n4533 gnd.n1971 242.672
R4692 gnd.n4533 gnd.n1972 242.672
R4693 gnd.n4533 gnd.n1973 242.672
R4694 gnd.n4533 gnd.n1974 242.672
R4695 gnd.n4533 gnd.n1975 242.672
R4696 gnd.n4533 gnd.n1976 242.672
R4697 gnd.n4533 gnd.n1977 242.672
R4698 gnd.n4533 gnd.n1978 242.672
R4699 gnd.n4533 gnd.n1979 242.672
R4700 gnd.n4533 gnd.n1980 242.672
R4701 gnd.n4533 gnd.n1981 242.672
R4702 gnd.n4533 gnd.n1982 242.672
R4703 gnd.n4533 gnd.n1983 242.672
R4704 gnd.n4533 gnd.n1984 242.672
R4705 gnd.n4533 gnd.n1985 242.672
R4706 gnd.n4533 gnd.n1986 242.672
R4707 gnd.n4533 gnd.n1987 242.672
R4708 gnd.n4534 gnd.n4533 242.672
R4709 gnd.n4722 gnd.n1096 242.672
R4710 gnd.n4711 gnd.n1096 242.672
R4711 gnd.n4708 gnd.n1096 242.672
R4712 gnd.n4699 gnd.n1096 242.672
R4713 gnd.n4688 gnd.n1096 242.672
R4714 gnd.n4685 gnd.n1096 242.672
R4715 gnd.n4676 gnd.n1096 242.672
R4716 gnd.n4666 gnd.n1096 242.672
R4717 gnd.n4663 gnd.n1096 242.672
R4718 gnd.n7178 gnd.n530 242.672
R4719 gnd.n7178 gnd.n532 242.672
R4720 gnd.n7178 gnd.n534 242.672
R4721 gnd.n7178 gnd.n535 242.672
R4722 gnd.n7178 gnd.n537 242.672
R4723 gnd.n7178 gnd.n539 242.672
R4724 gnd.n7178 gnd.n540 242.672
R4725 gnd.n7178 gnd.n542 242.672
R4726 gnd.n7178 gnd.n543 242.672
R4727 gnd.n128 gnd.n125 242.672
R4728 gnd.n7503 gnd.n128 242.672
R4729 gnd.n7499 gnd.n128 242.672
R4730 gnd.n7496 gnd.n128 242.672
R4731 gnd.n7491 gnd.n128 242.672
R4732 gnd.n7488 gnd.n128 242.672
R4733 gnd.n7483 gnd.n128 242.672
R4734 gnd.n7480 gnd.n128 242.672
R4735 gnd.n7475 gnd.n128 242.672
R4736 gnd.n6186 gnd.n1096 242.672
R4737 gnd.n1160 gnd.n1096 242.672
R4738 gnd.n6193 gnd.n1096 242.672
R4739 gnd.n1151 gnd.n1096 242.672
R4740 gnd.n6200 gnd.n1096 242.672
R4741 gnd.n1144 gnd.n1096 242.672
R4742 gnd.n6207 gnd.n1096 242.672
R4743 gnd.n1137 gnd.n1096 242.672
R4744 gnd.n6214 gnd.n1096 242.672
R4745 gnd.n1130 gnd.n1096 242.672
R4746 gnd.n6221 gnd.n1096 242.672
R4747 gnd.n6222 gnd.n1122 242.672
R4748 gnd.n6223 gnd.n1096 242.672
R4749 gnd.n1119 gnd.n1096 242.672
R4750 gnd.n6230 gnd.n1096 242.672
R4751 gnd.n1112 gnd.n1096 242.672
R4752 gnd.n6237 gnd.n1096 242.672
R4753 gnd.n1105 gnd.n1096 242.672
R4754 gnd.n6244 gnd.n1096 242.672
R4755 gnd.n6247 gnd.n1096 242.672
R4756 gnd.n7178 gnd.n7177 242.672
R4757 gnd.n7178 gnd.n512 242.672
R4758 gnd.n7178 gnd.n513 242.672
R4759 gnd.n7178 gnd.n514 242.672
R4760 gnd.n7178 gnd.n515 242.672
R4761 gnd.n7178 gnd.n516 242.672
R4762 gnd.n7178 gnd.n517 242.672
R4763 gnd.n7178 gnd.n518 242.672
R4764 gnd.n7147 gnd.n562 242.672
R4765 gnd.n7178 gnd.n519 242.672
R4766 gnd.n7178 gnd.n520 242.672
R4767 gnd.n7178 gnd.n521 242.672
R4768 gnd.n7178 gnd.n522 242.672
R4769 gnd.n7178 gnd.n523 242.672
R4770 gnd.n7178 gnd.n524 242.672
R4771 gnd.n7178 gnd.n525 242.672
R4772 gnd.n7178 gnd.n526 242.672
R4773 gnd.n7178 gnd.n527 242.672
R4774 gnd.n7178 gnd.n528 242.672
R4775 gnd.n7178 gnd.n529 242.672
R4776 gnd.n198 gnd.n128 242.672
R4777 gnd.n7560 gnd.n128 242.672
R4778 gnd.n194 gnd.n128 242.672
R4779 gnd.n7567 gnd.n128 242.672
R4780 gnd.n187 gnd.n128 242.672
R4781 gnd.n7574 gnd.n128 242.672
R4782 gnd.n180 gnd.n128 242.672
R4783 gnd.n7581 gnd.n128 242.672
R4784 gnd.n173 gnd.n128 242.672
R4785 gnd.n7588 gnd.n128 242.672
R4786 gnd.n166 gnd.n128 242.672
R4787 gnd.n7598 gnd.n128 242.672
R4788 gnd.n159 gnd.n128 242.672
R4789 gnd.n7605 gnd.n128 242.672
R4790 gnd.n152 gnd.n128 242.672
R4791 gnd.n7612 gnd.n128 242.672
R4792 gnd.n145 gnd.n128 242.672
R4793 gnd.n7619 gnd.n128 242.672
R4794 gnd.n138 gnd.n128 242.672
R4795 gnd.n4771 gnd.n4770 242.672
R4796 gnd.n4771 gnd.n4635 242.672
R4797 gnd.n4771 gnd.n4636 242.672
R4798 gnd.n4771 gnd.n4637 242.672
R4799 gnd.n4771 gnd.n4638 242.672
R4800 gnd.n4771 gnd.n4639 242.672
R4801 gnd.n4771 gnd.n4640 242.672
R4802 gnd.n4771 gnd.n4641 242.672
R4803 gnd.n4771 gnd.n4642 242.672
R4804 gnd.n4771 gnd.n4643 242.672
R4805 gnd.n4771 gnd.n4645 242.672
R4806 gnd.n4771 gnd.n4646 242.672
R4807 gnd.n4771 gnd.n4647 242.672
R4808 gnd.n4771 gnd.n4649 242.672
R4809 gnd.n5984 gnd.n5839 242.672
R4810 gnd.n5984 gnd.n5838 242.672
R4811 gnd.n5984 gnd.n5837 242.672
R4812 gnd.n5984 gnd.n5836 242.672
R4813 gnd.n5984 gnd.n5835 242.672
R4814 gnd.n5984 gnd.n5834 242.672
R4815 gnd.n5984 gnd.n5833 242.672
R4816 gnd.n5984 gnd.n5831 242.672
R4817 gnd.n5984 gnd.n5830 242.672
R4818 gnd.n5984 gnd.n5828 242.672
R4819 gnd.n5984 gnd.n5826 242.672
R4820 gnd.n5984 gnd.n5825 242.672
R4821 gnd.n5984 gnd.n5823 242.672
R4822 gnd.n5984 gnd.n5821 242.672
R4823 gnd.n135 gnd.n131 240.244
R4824 gnd.n7621 gnd.n7620 240.244
R4825 gnd.n7618 gnd.n139 240.244
R4826 gnd.n7614 gnd.n7613 240.244
R4827 gnd.n7611 gnd.n146 240.244
R4828 gnd.n7607 gnd.n7606 240.244
R4829 gnd.n7604 gnd.n153 240.244
R4830 gnd.n7600 gnd.n7599 240.244
R4831 gnd.n7597 gnd.n160 240.244
R4832 gnd.n7590 gnd.n7589 240.244
R4833 gnd.n7587 gnd.n167 240.244
R4834 gnd.n7583 gnd.n7582 240.244
R4835 gnd.n7580 gnd.n174 240.244
R4836 gnd.n7576 gnd.n7575 240.244
R4837 gnd.n7573 gnd.n181 240.244
R4838 gnd.n7569 gnd.n7568 240.244
R4839 gnd.n7566 gnd.n188 240.244
R4840 gnd.n7562 gnd.n7561 240.244
R4841 gnd.n7559 gnd.n195 240.244
R4842 gnd.n590 gnd.n456 240.244
R4843 gnd.n590 gnd.n448 240.244
R4844 gnd.n7099 gnd.n448 240.244
R4845 gnd.n7099 gnd.n440 240.244
R4846 gnd.n5867 gnd.n440 240.244
R4847 gnd.n5867 gnd.n431 240.244
R4848 gnd.n5871 gnd.n431 240.244
R4849 gnd.n5871 gnd.n422 240.244
R4850 gnd.n5916 gnd.n422 240.244
R4851 gnd.n5916 gnd.n413 240.244
R4852 gnd.n5912 gnd.n413 240.244
R4853 gnd.n5912 gnd.n406 240.244
R4854 gnd.n5908 gnd.n406 240.244
R4855 gnd.n5908 gnd.n397 240.244
R4856 gnd.n5883 gnd.n397 240.244
R4857 gnd.n5883 gnd.n388 240.244
R4858 gnd.n6929 gnd.n388 240.244
R4859 gnd.n6929 gnd.n379 240.244
R4860 gnd.n7039 gnd.n379 240.244
R4861 gnd.n7039 gnd.n372 240.244
R4862 gnd.n7035 gnd.n372 240.244
R4863 gnd.n7035 gnd.n363 240.244
R4864 gnd.n7032 gnd.n363 240.244
R4865 gnd.n7032 gnd.n354 240.244
R4866 gnd.n7029 gnd.n354 240.244
R4867 gnd.n7029 gnd.n346 240.244
R4868 gnd.n7026 gnd.n346 240.244
R4869 gnd.n7026 gnd.n339 240.244
R4870 gnd.n7023 gnd.n339 240.244
R4871 gnd.n7023 gnd.n331 240.244
R4872 gnd.n7020 gnd.n331 240.244
R4873 gnd.n7020 gnd.n321 240.244
R4874 gnd.n7017 gnd.n321 240.244
R4875 gnd.n7017 gnd.n313 240.244
R4876 gnd.n7014 gnd.n313 240.244
R4877 gnd.n7014 gnd.n306 240.244
R4878 gnd.n7011 gnd.n306 240.244
R4879 gnd.n7011 gnd.n300 240.244
R4880 gnd.n7008 gnd.n300 240.244
R4881 gnd.n7008 gnd.n291 240.244
R4882 gnd.n7005 gnd.n291 240.244
R4883 gnd.n7005 gnd.n283 240.244
R4884 gnd.n7002 gnd.n283 240.244
R4885 gnd.n7002 gnd.n276 240.244
R4886 gnd.n6999 gnd.n276 240.244
R4887 gnd.n6999 gnd.n270 240.244
R4888 gnd.n6996 gnd.n270 240.244
R4889 gnd.n6996 gnd.n261 240.244
R4890 gnd.n6993 gnd.n261 240.244
R4891 gnd.n6993 gnd.n253 240.244
R4892 gnd.n6990 gnd.n253 240.244
R4893 gnd.n6990 gnd.n245 240.244
R4894 gnd.n6987 gnd.n245 240.244
R4895 gnd.n6987 gnd.n239 240.244
R4896 gnd.n6984 gnd.n239 240.244
R4897 gnd.n6984 gnd.n230 240.244
R4898 gnd.n6981 gnd.n230 240.244
R4899 gnd.n6981 gnd.n223 240.244
R4900 gnd.n6978 gnd.n223 240.244
R4901 gnd.n6978 gnd.n214 240.244
R4902 gnd.n214 gnd.n205 240.244
R4903 gnd.n7550 gnd.n205 240.244
R4904 gnd.n7551 gnd.n7550 240.244
R4905 gnd.n7551 gnd.n127 240.244
R4906 gnd.n7176 gnd.n544 240.244
R4907 gnd.n7172 gnd.n544 240.244
R4908 gnd.n7170 gnd.n7169 240.244
R4909 gnd.n7166 gnd.n7165 240.244
R4910 gnd.n7162 gnd.n7161 240.244
R4911 gnd.n7158 gnd.n7157 240.244
R4912 gnd.n7154 gnd.n7153 240.244
R4913 gnd.n7150 gnd.n7149 240.244
R4914 gnd.n7145 gnd.n7144 240.244
R4915 gnd.n7141 gnd.n7140 240.244
R4916 gnd.n7137 gnd.n7136 240.244
R4917 gnd.n7133 gnd.n7132 240.244
R4918 gnd.n7129 gnd.n7128 240.244
R4919 gnd.n7125 gnd.n7124 240.244
R4920 gnd.n7121 gnd.n7120 240.244
R4921 gnd.n7117 gnd.n7116 240.244
R4922 gnd.n7113 gnd.n7112 240.244
R4923 gnd.n585 gnd.n584 240.244
R4924 gnd.n7234 gnd.n451 240.244
R4925 gnd.n7240 gnd.n451 240.244
R4926 gnd.n7240 gnd.n438 240.244
R4927 gnd.n7250 gnd.n438 240.244
R4928 gnd.n7250 gnd.n434 240.244
R4929 gnd.n7256 gnd.n434 240.244
R4930 gnd.n7256 gnd.n420 240.244
R4931 gnd.n7266 gnd.n420 240.244
R4932 gnd.n7266 gnd.n416 240.244
R4933 gnd.n7272 gnd.n416 240.244
R4934 gnd.n7272 gnd.n404 240.244
R4935 gnd.n7282 gnd.n404 240.244
R4936 gnd.n7282 gnd.n400 240.244
R4937 gnd.n7288 gnd.n400 240.244
R4938 gnd.n7288 gnd.n386 240.244
R4939 gnd.n7298 gnd.n386 240.244
R4940 gnd.n7298 gnd.n382 240.244
R4941 gnd.n7304 gnd.n382 240.244
R4942 gnd.n7304 gnd.n370 240.244
R4943 gnd.n7314 gnd.n370 240.244
R4944 gnd.n7314 gnd.n366 240.244
R4945 gnd.n7320 gnd.n366 240.244
R4946 gnd.n7320 gnd.n352 240.244
R4947 gnd.n7330 gnd.n352 240.244
R4948 gnd.n7330 gnd.n348 240.244
R4949 gnd.n7336 gnd.n348 240.244
R4950 gnd.n7336 gnd.n337 240.244
R4951 gnd.n7346 gnd.n337 240.244
R4952 gnd.n7346 gnd.n333 240.244
R4953 gnd.n7352 gnd.n333 240.244
R4954 gnd.n7352 gnd.n319 240.244
R4955 gnd.n7362 gnd.n319 240.244
R4956 gnd.n7362 gnd.n315 240.244
R4957 gnd.n7368 gnd.n315 240.244
R4958 gnd.n7368 gnd.n305 240.244
R4959 gnd.n7378 gnd.n305 240.244
R4960 gnd.n7378 gnd.n301 240.244
R4961 gnd.n7384 gnd.n301 240.244
R4962 gnd.n7384 gnd.n289 240.244
R4963 gnd.n7394 gnd.n289 240.244
R4964 gnd.n7394 gnd.n285 240.244
R4965 gnd.n7400 gnd.n285 240.244
R4966 gnd.n7400 gnd.n275 240.244
R4967 gnd.n7410 gnd.n275 240.244
R4968 gnd.n7410 gnd.n271 240.244
R4969 gnd.n7416 gnd.n271 240.244
R4970 gnd.n7416 gnd.n259 240.244
R4971 gnd.n7426 gnd.n259 240.244
R4972 gnd.n7426 gnd.n255 240.244
R4973 gnd.n7432 gnd.n255 240.244
R4974 gnd.n7432 gnd.n244 240.244
R4975 gnd.n7442 gnd.n244 240.244
R4976 gnd.n7442 gnd.n240 240.244
R4977 gnd.n7448 gnd.n240 240.244
R4978 gnd.n7448 gnd.n228 240.244
R4979 gnd.n7458 gnd.n228 240.244
R4980 gnd.n7458 gnd.n224 240.244
R4981 gnd.n7464 gnd.n224 240.244
R4982 gnd.n7464 gnd.n212 240.244
R4983 gnd.n7542 gnd.n212 240.244
R4984 gnd.n7542 gnd.n208 240.244
R4985 gnd.n7548 gnd.n208 240.244
R4986 gnd.n7548 gnd.n130 240.244
R4987 gnd.n7628 gnd.n130 240.244
R4988 gnd.n7474 gnd.n7473 240.244
R4989 gnd.n7479 gnd.n7476 240.244
R4990 gnd.n7482 gnd.n7481 240.244
R4991 gnd.n7487 gnd.n7484 240.244
R4992 gnd.n7490 gnd.n7489 240.244
R4993 gnd.n7495 gnd.n7492 240.244
R4994 gnd.n7498 gnd.n7497 240.244
R4995 gnd.n7502 gnd.n7500 240.244
R4996 gnd.n7505 gnd.n7504 240.244
R4997 gnd.n5972 gnd.n457 240.244
R4998 gnd.n5972 gnd.n449 240.244
R4999 gnd.n7097 gnd.n449 240.244
R5000 gnd.n7097 gnd.n441 240.244
R5001 gnd.n598 gnd.n441 240.244
R5002 gnd.n598 gnd.n432 240.244
R5003 gnd.n599 gnd.n432 240.244
R5004 gnd.n599 gnd.n423 240.244
R5005 gnd.n602 gnd.n423 240.244
R5006 gnd.n602 gnd.n414 240.244
R5007 gnd.n603 gnd.n414 240.244
R5008 gnd.n603 gnd.n407 240.244
R5009 gnd.n606 gnd.n407 240.244
R5010 gnd.n606 gnd.n398 240.244
R5011 gnd.n607 gnd.n398 240.244
R5012 gnd.n607 gnd.n389 240.244
R5013 gnd.n610 gnd.n389 240.244
R5014 gnd.n610 gnd.n380 240.244
R5015 gnd.n7041 gnd.n380 240.244
R5016 gnd.n7041 gnd.n373 240.244
R5017 gnd.n7044 gnd.n373 240.244
R5018 gnd.n7044 gnd.n364 240.244
R5019 gnd.n7045 gnd.n364 240.244
R5020 gnd.n7045 gnd.n355 240.244
R5021 gnd.n7048 gnd.n355 240.244
R5022 gnd.n7048 gnd.n347 240.244
R5023 gnd.n7049 gnd.n347 240.244
R5024 gnd.n7049 gnd.n340 240.244
R5025 gnd.n7052 gnd.n340 240.244
R5026 gnd.n7052 gnd.n332 240.244
R5027 gnd.n7053 gnd.n332 240.244
R5028 gnd.n7053 gnd.n322 240.244
R5029 gnd.n322 gnd.n82 240.244
R5030 gnd.n83 gnd.n82 240.244
R5031 gnd.n84 gnd.n83 240.244
R5032 gnd.n307 gnd.n84 240.244
R5033 gnd.n307 gnd.n87 240.244
R5034 gnd.n88 gnd.n87 240.244
R5035 gnd.n89 gnd.n88 240.244
R5036 gnd.n292 gnd.n89 240.244
R5037 gnd.n292 gnd.n92 240.244
R5038 gnd.n93 gnd.n92 240.244
R5039 gnd.n94 gnd.n93 240.244
R5040 gnd.n277 gnd.n94 240.244
R5041 gnd.n277 gnd.n97 240.244
R5042 gnd.n98 gnd.n97 240.244
R5043 gnd.n99 gnd.n98 240.244
R5044 gnd.n262 gnd.n99 240.244
R5045 gnd.n262 gnd.n102 240.244
R5046 gnd.n103 gnd.n102 240.244
R5047 gnd.n104 gnd.n103 240.244
R5048 gnd.n246 gnd.n104 240.244
R5049 gnd.n246 gnd.n107 240.244
R5050 gnd.n108 gnd.n107 240.244
R5051 gnd.n109 gnd.n108 240.244
R5052 gnd.n231 gnd.n109 240.244
R5053 gnd.n231 gnd.n112 240.244
R5054 gnd.n113 gnd.n112 240.244
R5055 gnd.n114 gnd.n113 240.244
R5056 gnd.n215 gnd.n114 240.244
R5057 gnd.n215 gnd.n117 240.244
R5058 gnd.n118 gnd.n117 240.244
R5059 gnd.n119 gnd.n118 240.244
R5060 gnd.n7630 gnd.n119 240.244
R5061 gnd.n531 gnd.n461 240.244
R5062 gnd.n469 gnd.n468 240.244
R5063 gnd.n533 gnd.n476 240.244
R5064 gnd.n536 gnd.n477 240.244
R5065 gnd.n485 gnd.n484 240.244
R5066 gnd.n538 gnd.n492 240.244
R5067 gnd.n541 gnd.n493 240.244
R5068 gnd.n501 gnd.n500 240.244
R5069 gnd.n7179 gnd.n510 240.244
R5070 gnd.n7232 gnd.n447 240.244
R5071 gnd.n7242 gnd.n447 240.244
R5072 gnd.n7242 gnd.n443 240.244
R5073 gnd.n7248 gnd.n443 240.244
R5074 gnd.n7248 gnd.n429 240.244
R5075 gnd.n7258 gnd.n429 240.244
R5076 gnd.n7258 gnd.n425 240.244
R5077 gnd.n7264 gnd.n425 240.244
R5078 gnd.n7264 gnd.n412 240.244
R5079 gnd.n7274 gnd.n412 240.244
R5080 gnd.n7274 gnd.n408 240.244
R5081 gnd.n7280 gnd.n408 240.244
R5082 gnd.n7280 gnd.n395 240.244
R5083 gnd.n7290 gnd.n395 240.244
R5084 gnd.n7290 gnd.n391 240.244
R5085 gnd.n7296 gnd.n391 240.244
R5086 gnd.n7296 gnd.n378 240.244
R5087 gnd.n7306 gnd.n378 240.244
R5088 gnd.n7306 gnd.n374 240.244
R5089 gnd.n7312 gnd.n374 240.244
R5090 gnd.n7312 gnd.n361 240.244
R5091 gnd.n7322 gnd.n361 240.244
R5092 gnd.n7322 gnd.n357 240.244
R5093 gnd.n7328 gnd.n357 240.244
R5094 gnd.n7328 gnd.n345 240.244
R5095 gnd.n7338 gnd.n345 240.244
R5096 gnd.n7338 gnd.n341 240.244
R5097 gnd.n7344 gnd.n341 240.244
R5098 gnd.n7344 gnd.n329 240.244
R5099 gnd.n7354 gnd.n329 240.244
R5100 gnd.n7354 gnd.n324 240.244
R5101 gnd.n7360 gnd.n324 240.244
R5102 gnd.n7360 gnd.n312 240.244
R5103 gnd.n7370 gnd.n312 240.244
R5104 gnd.n7370 gnd.n308 240.244
R5105 gnd.n7376 gnd.n308 240.244
R5106 gnd.n7376 gnd.n298 240.244
R5107 gnd.n7386 gnd.n298 240.244
R5108 gnd.n7386 gnd.n294 240.244
R5109 gnd.n7392 gnd.n294 240.244
R5110 gnd.n7392 gnd.n282 240.244
R5111 gnd.n7402 gnd.n282 240.244
R5112 gnd.n7402 gnd.n278 240.244
R5113 gnd.n7408 gnd.n278 240.244
R5114 gnd.n7408 gnd.n268 240.244
R5115 gnd.n7418 gnd.n268 240.244
R5116 gnd.n7418 gnd.n264 240.244
R5117 gnd.n7424 gnd.n264 240.244
R5118 gnd.n7424 gnd.n251 240.244
R5119 gnd.n7434 gnd.n251 240.244
R5120 gnd.n7434 gnd.n247 240.244
R5121 gnd.n7440 gnd.n247 240.244
R5122 gnd.n7440 gnd.n237 240.244
R5123 gnd.n7450 gnd.n237 240.244
R5124 gnd.n7450 gnd.n233 240.244
R5125 gnd.n7456 gnd.n233 240.244
R5126 gnd.n7456 gnd.n222 240.244
R5127 gnd.n7466 gnd.n222 240.244
R5128 gnd.n7466 gnd.n216 240.244
R5129 gnd.n7540 gnd.n216 240.244
R5130 gnd.n7540 gnd.n217 240.244
R5131 gnd.n217 gnd.n207 240.244
R5132 gnd.n7471 gnd.n207 240.244
R5133 gnd.n7471 gnd.n129 240.244
R5134 gnd.n6320 gnd.n978 240.244
R5135 gnd.n6320 gnd.n974 240.244
R5136 gnd.n6326 gnd.n974 240.244
R5137 gnd.n6326 gnd.n972 240.244
R5138 gnd.n6330 gnd.n972 240.244
R5139 gnd.n6330 gnd.n968 240.244
R5140 gnd.n6336 gnd.n968 240.244
R5141 gnd.n6336 gnd.n966 240.244
R5142 gnd.n6340 gnd.n966 240.244
R5143 gnd.n6340 gnd.n962 240.244
R5144 gnd.n6346 gnd.n962 240.244
R5145 gnd.n6346 gnd.n960 240.244
R5146 gnd.n6350 gnd.n960 240.244
R5147 gnd.n6350 gnd.n956 240.244
R5148 gnd.n6356 gnd.n956 240.244
R5149 gnd.n6356 gnd.n954 240.244
R5150 gnd.n6360 gnd.n954 240.244
R5151 gnd.n6360 gnd.n950 240.244
R5152 gnd.n6366 gnd.n950 240.244
R5153 gnd.n6366 gnd.n948 240.244
R5154 gnd.n6370 gnd.n948 240.244
R5155 gnd.n6370 gnd.n944 240.244
R5156 gnd.n6376 gnd.n944 240.244
R5157 gnd.n6376 gnd.n942 240.244
R5158 gnd.n6380 gnd.n942 240.244
R5159 gnd.n6380 gnd.n938 240.244
R5160 gnd.n6386 gnd.n938 240.244
R5161 gnd.n6386 gnd.n936 240.244
R5162 gnd.n6390 gnd.n936 240.244
R5163 gnd.n6390 gnd.n932 240.244
R5164 gnd.n6396 gnd.n932 240.244
R5165 gnd.n6396 gnd.n930 240.244
R5166 gnd.n6400 gnd.n930 240.244
R5167 gnd.n6400 gnd.n926 240.244
R5168 gnd.n6406 gnd.n926 240.244
R5169 gnd.n6406 gnd.n924 240.244
R5170 gnd.n6410 gnd.n924 240.244
R5171 gnd.n6410 gnd.n920 240.244
R5172 gnd.n6416 gnd.n920 240.244
R5173 gnd.n6416 gnd.n918 240.244
R5174 gnd.n6420 gnd.n918 240.244
R5175 gnd.n6420 gnd.n914 240.244
R5176 gnd.n6426 gnd.n914 240.244
R5177 gnd.n6426 gnd.n912 240.244
R5178 gnd.n6430 gnd.n912 240.244
R5179 gnd.n6430 gnd.n908 240.244
R5180 gnd.n6436 gnd.n908 240.244
R5181 gnd.n6436 gnd.n906 240.244
R5182 gnd.n6440 gnd.n906 240.244
R5183 gnd.n6440 gnd.n902 240.244
R5184 gnd.n6446 gnd.n902 240.244
R5185 gnd.n6446 gnd.n900 240.244
R5186 gnd.n6450 gnd.n900 240.244
R5187 gnd.n6450 gnd.n896 240.244
R5188 gnd.n6456 gnd.n896 240.244
R5189 gnd.n6456 gnd.n894 240.244
R5190 gnd.n6460 gnd.n894 240.244
R5191 gnd.n6460 gnd.n890 240.244
R5192 gnd.n6466 gnd.n890 240.244
R5193 gnd.n6466 gnd.n888 240.244
R5194 gnd.n6470 gnd.n888 240.244
R5195 gnd.n6470 gnd.n884 240.244
R5196 gnd.n6476 gnd.n884 240.244
R5197 gnd.n6476 gnd.n882 240.244
R5198 gnd.n6480 gnd.n882 240.244
R5199 gnd.n6480 gnd.n878 240.244
R5200 gnd.n6486 gnd.n878 240.244
R5201 gnd.n6486 gnd.n876 240.244
R5202 gnd.n6490 gnd.n876 240.244
R5203 gnd.n6490 gnd.n872 240.244
R5204 gnd.n6496 gnd.n872 240.244
R5205 gnd.n6496 gnd.n870 240.244
R5206 gnd.n6500 gnd.n870 240.244
R5207 gnd.n6500 gnd.n866 240.244
R5208 gnd.n6506 gnd.n866 240.244
R5209 gnd.n6506 gnd.n864 240.244
R5210 gnd.n6510 gnd.n864 240.244
R5211 gnd.n6510 gnd.n860 240.244
R5212 gnd.n6516 gnd.n860 240.244
R5213 gnd.n6516 gnd.n858 240.244
R5214 gnd.n6520 gnd.n858 240.244
R5215 gnd.n6520 gnd.n854 240.244
R5216 gnd.n6526 gnd.n854 240.244
R5217 gnd.n6526 gnd.n852 240.244
R5218 gnd.n6530 gnd.n852 240.244
R5219 gnd.n6530 gnd.n848 240.244
R5220 gnd.n6536 gnd.n848 240.244
R5221 gnd.n6536 gnd.n846 240.244
R5222 gnd.n6540 gnd.n846 240.244
R5223 gnd.n6540 gnd.n842 240.244
R5224 gnd.n6546 gnd.n842 240.244
R5225 gnd.n6546 gnd.n840 240.244
R5226 gnd.n6550 gnd.n840 240.244
R5227 gnd.n6550 gnd.n836 240.244
R5228 gnd.n6556 gnd.n836 240.244
R5229 gnd.n6556 gnd.n834 240.244
R5230 gnd.n6560 gnd.n834 240.244
R5231 gnd.n6560 gnd.n830 240.244
R5232 gnd.n6566 gnd.n830 240.244
R5233 gnd.n6566 gnd.n828 240.244
R5234 gnd.n6570 gnd.n828 240.244
R5235 gnd.n6570 gnd.n824 240.244
R5236 gnd.n6576 gnd.n824 240.244
R5237 gnd.n6576 gnd.n822 240.244
R5238 gnd.n6580 gnd.n822 240.244
R5239 gnd.n6580 gnd.n818 240.244
R5240 gnd.n6586 gnd.n818 240.244
R5241 gnd.n6586 gnd.n816 240.244
R5242 gnd.n6590 gnd.n816 240.244
R5243 gnd.n6590 gnd.n812 240.244
R5244 gnd.n6596 gnd.n812 240.244
R5245 gnd.n6596 gnd.n810 240.244
R5246 gnd.n6600 gnd.n810 240.244
R5247 gnd.n6600 gnd.n806 240.244
R5248 gnd.n6606 gnd.n806 240.244
R5249 gnd.n6606 gnd.n804 240.244
R5250 gnd.n6610 gnd.n804 240.244
R5251 gnd.n6610 gnd.n800 240.244
R5252 gnd.n6616 gnd.n800 240.244
R5253 gnd.n6616 gnd.n798 240.244
R5254 gnd.n6620 gnd.n798 240.244
R5255 gnd.n6620 gnd.n794 240.244
R5256 gnd.n6626 gnd.n794 240.244
R5257 gnd.n6626 gnd.n792 240.244
R5258 gnd.n6630 gnd.n792 240.244
R5259 gnd.n6630 gnd.n788 240.244
R5260 gnd.n6636 gnd.n788 240.244
R5261 gnd.n6636 gnd.n786 240.244
R5262 gnd.n6640 gnd.n786 240.244
R5263 gnd.n6640 gnd.n782 240.244
R5264 gnd.n6646 gnd.n782 240.244
R5265 gnd.n6646 gnd.n780 240.244
R5266 gnd.n6650 gnd.n780 240.244
R5267 gnd.n6650 gnd.n776 240.244
R5268 gnd.n6656 gnd.n776 240.244
R5269 gnd.n6656 gnd.n774 240.244
R5270 gnd.n6660 gnd.n774 240.244
R5271 gnd.n6660 gnd.n770 240.244
R5272 gnd.n6666 gnd.n770 240.244
R5273 gnd.n6666 gnd.n768 240.244
R5274 gnd.n6670 gnd.n768 240.244
R5275 gnd.n6670 gnd.n764 240.244
R5276 gnd.n6676 gnd.n764 240.244
R5277 gnd.n6676 gnd.n762 240.244
R5278 gnd.n6680 gnd.n762 240.244
R5279 gnd.n6680 gnd.n758 240.244
R5280 gnd.n6686 gnd.n758 240.244
R5281 gnd.n6686 gnd.n756 240.244
R5282 gnd.n6690 gnd.n756 240.244
R5283 gnd.n6690 gnd.n752 240.244
R5284 gnd.n6697 gnd.n752 240.244
R5285 gnd.n6697 gnd.n750 240.244
R5286 gnd.n6701 gnd.n750 240.244
R5287 gnd.n6701 gnd.n747 240.244
R5288 gnd.n6707 gnd.n745 240.244
R5289 gnd.n6711 gnd.n745 240.244
R5290 gnd.n6711 gnd.n741 240.244
R5291 gnd.n6717 gnd.n741 240.244
R5292 gnd.n6717 gnd.n739 240.244
R5293 gnd.n6721 gnd.n739 240.244
R5294 gnd.n6721 gnd.n735 240.244
R5295 gnd.n6727 gnd.n735 240.244
R5296 gnd.n6727 gnd.n733 240.244
R5297 gnd.n6731 gnd.n733 240.244
R5298 gnd.n6731 gnd.n729 240.244
R5299 gnd.n6737 gnd.n729 240.244
R5300 gnd.n6737 gnd.n727 240.244
R5301 gnd.n6741 gnd.n727 240.244
R5302 gnd.n6741 gnd.n723 240.244
R5303 gnd.n6747 gnd.n723 240.244
R5304 gnd.n6747 gnd.n721 240.244
R5305 gnd.n6751 gnd.n721 240.244
R5306 gnd.n6751 gnd.n717 240.244
R5307 gnd.n6757 gnd.n717 240.244
R5308 gnd.n6757 gnd.n715 240.244
R5309 gnd.n6761 gnd.n715 240.244
R5310 gnd.n6761 gnd.n711 240.244
R5311 gnd.n6767 gnd.n711 240.244
R5312 gnd.n6767 gnd.n709 240.244
R5313 gnd.n6771 gnd.n709 240.244
R5314 gnd.n6771 gnd.n705 240.244
R5315 gnd.n6777 gnd.n705 240.244
R5316 gnd.n6777 gnd.n703 240.244
R5317 gnd.n6781 gnd.n703 240.244
R5318 gnd.n6781 gnd.n699 240.244
R5319 gnd.n6787 gnd.n699 240.244
R5320 gnd.n6787 gnd.n697 240.244
R5321 gnd.n6791 gnd.n697 240.244
R5322 gnd.n6791 gnd.n693 240.244
R5323 gnd.n6797 gnd.n693 240.244
R5324 gnd.n6797 gnd.n691 240.244
R5325 gnd.n6801 gnd.n691 240.244
R5326 gnd.n6801 gnd.n687 240.244
R5327 gnd.n6807 gnd.n687 240.244
R5328 gnd.n6807 gnd.n685 240.244
R5329 gnd.n6811 gnd.n685 240.244
R5330 gnd.n6811 gnd.n681 240.244
R5331 gnd.n6817 gnd.n681 240.244
R5332 gnd.n6817 gnd.n679 240.244
R5333 gnd.n6821 gnd.n679 240.244
R5334 gnd.n6821 gnd.n675 240.244
R5335 gnd.n6827 gnd.n675 240.244
R5336 gnd.n6827 gnd.n673 240.244
R5337 gnd.n6831 gnd.n673 240.244
R5338 gnd.n6831 gnd.n669 240.244
R5339 gnd.n6837 gnd.n669 240.244
R5340 gnd.n6837 gnd.n667 240.244
R5341 gnd.n6841 gnd.n667 240.244
R5342 gnd.n6841 gnd.n663 240.244
R5343 gnd.n6847 gnd.n663 240.244
R5344 gnd.n6847 gnd.n661 240.244
R5345 gnd.n6851 gnd.n661 240.244
R5346 gnd.n6851 gnd.n657 240.244
R5347 gnd.n6857 gnd.n657 240.244
R5348 gnd.n6857 gnd.n655 240.244
R5349 gnd.n6861 gnd.n655 240.244
R5350 gnd.n6861 gnd.n651 240.244
R5351 gnd.n6867 gnd.n651 240.244
R5352 gnd.n6867 gnd.n649 240.244
R5353 gnd.n6871 gnd.n649 240.244
R5354 gnd.n6871 gnd.n645 240.244
R5355 gnd.n6877 gnd.n645 240.244
R5356 gnd.n6877 gnd.n643 240.244
R5357 gnd.n6881 gnd.n643 240.244
R5358 gnd.n6881 gnd.n639 240.244
R5359 gnd.n6887 gnd.n639 240.244
R5360 gnd.n6887 gnd.n637 240.244
R5361 gnd.n6891 gnd.n637 240.244
R5362 gnd.n6891 gnd.n633 240.244
R5363 gnd.n6897 gnd.n633 240.244
R5364 gnd.n6897 gnd.n631 240.244
R5365 gnd.n6901 gnd.n631 240.244
R5366 gnd.n6901 gnd.n627 240.244
R5367 gnd.n6907 gnd.n627 240.244
R5368 gnd.n6907 gnd.n625 240.244
R5369 gnd.n6912 gnd.n625 240.244
R5370 gnd.n6912 gnd.n621 240.244
R5371 gnd.n6919 gnd.n621 240.244
R5372 gnd.n4541 gnd.n980 240.244
R5373 gnd.n4542 gnd.n4541 240.244
R5374 gnd.n4542 gnd.n1942 240.244
R5375 gnd.n4548 gnd.n1942 240.244
R5376 gnd.n4549 gnd.n4548 240.244
R5377 gnd.n4550 gnd.n4549 240.244
R5378 gnd.n4550 gnd.n1937 240.244
R5379 gnd.n4561 gnd.n1937 240.244
R5380 gnd.n4561 gnd.n1938 240.244
R5381 gnd.n1938 gnd.n1917 240.244
R5382 gnd.n4608 gnd.n1917 240.244
R5383 gnd.n4609 gnd.n4608 240.244
R5384 gnd.n4610 gnd.n4609 240.244
R5385 gnd.n4610 gnd.n1913 240.244
R5386 gnd.n4616 gnd.n1913 240.244
R5387 gnd.n4617 gnd.n4616 240.244
R5388 gnd.n4618 gnd.n4617 240.244
R5389 gnd.n4618 gnd.n1909 240.244
R5390 gnd.n4624 gnd.n1909 240.244
R5391 gnd.n4625 gnd.n4624 240.244
R5392 gnd.n4626 gnd.n4625 240.244
R5393 gnd.n4626 gnd.n1905 240.244
R5394 gnd.n4632 gnd.n1905 240.244
R5395 gnd.n4632 gnd.n1903 240.244
R5396 gnd.n4774 gnd.n1903 240.244
R5397 gnd.n4774 gnd.n1899 240.244
R5398 gnd.n4780 gnd.n1899 240.244
R5399 gnd.n4780 gnd.n1889 240.244
R5400 gnd.n4793 gnd.n1889 240.244
R5401 gnd.n4793 gnd.n1885 240.244
R5402 gnd.n4799 gnd.n1885 240.244
R5403 gnd.n4799 gnd.n1875 240.244
R5404 gnd.n4812 gnd.n1875 240.244
R5405 gnd.n4812 gnd.n1871 240.244
R5406 gnd.n4818 gnd.n1871 240.244
R5407 gnd.n4818 gnd.n1861 240.244
R5408 gnd.n4831 gnd.n1861 240.244
R5409 gnd.n4831 gnd.n1857 240.244
R5410 gnd.n4837 gnd.n1857 240.244
R5411 gnd.n4837 gnd.n1847 240.244
R5412 gnd.n4850 gnd.n1847 240.244
R5413 gnd.n4850 gnd.n1843 240.244
R5414 gnd.n4856 gnd.n1843 240.244
R5415 gnd.n4856 gnd.n1832 240.244
R5416 gnd.n4869 gnd.n1832 240.244
R5417 gnd.n4869 gnd.n1828 240.244
R5418 gnd.n4877 gnd.n1828 240.244
R5419 gnd.n4877 gnd.n1819 240.244
R5420 gnd.n5089 gnd.n1819 240.244
R5421 gnd.n5090 gnd.n5089 240.244
R5422 gnd.n5090 gnd.n1815 240.244
R5423 gnd.n5096 gnd.n1815 240.244
R5424 gnd.n5096 gnd.n1745 240.244
R5425 gnd.n5131 gnd.n1745 240.244
R5426 gnd.n5131 gnd.n1740 240.244
R5427 gnd.n5139 gnd.n1740 240.244
R5428 gnd.n5139 gnd.n1741 240.244
R5429 gnd.n1741 gnd.n1718 240.244
R5430 gnd.n5167 gnd.n1718 240.244
R5431 gnd.n5167 gnd.n1714 240.244
R5432 gnd.n5173 gnd.n1714 240.244
R5433 gnd.n5173 gnd.n1696 240.244
R5434 gnd.n5195 gnd.n1696 240.244
R5435 gnd.n5195 gnd.n1691 240.244
R5436 gnd.n5203 gnd.n1691 240.244
R5437 gnd.n5203 gnd.n1692 240.244
R5438 gnd.n1692 gnd.n1664 240.244
R5439 gnd.n5232 gnd.n1664 240.244
R5440 gnd.n5232 gnd.n1659 240.244
R5441 gnd.n5249 gnd.n1659 240.244
R5442 gnd.n5249 gnd.n1660 240.244
R5443 gnd.n5245 gnd.n1660 240.244
R5444 gnd.n5245 gnd.n5244 240.244
R5445 gnd.n5244 gnd.n5243 240.244
R5446 gnd.n5243 gnd.n1623 240.244
R5447 gnd.n5326 gnd.n1623 240.244
R5448 gnd.n5326 gnd.n1619 240.244
R5449 gnd.n5332 gnd.n1619 240.244
R5450 gnd.n5332 gnd.n1605 240.244
R5451 gnd.n5369 gnd.n1605 240.244
R5452 gnd.n5369 gnd.n1601 240.244
R5453 gnd.n5375 gnd.n1601 240.244
R5454 gnd.n5375 gnd.n1581 240.244
R5455 gnd.n5403 gnd.n1581 240.244
R5456 gnd.n5403 gnd.n1577 240.244
R5457 gnd.n5409 gnd.n1577 240.244
R5458 gnd.n5409 gnd.n1558 240.244
R5459 gnd.n5444 gnd.n1558 240.244
R5460 gnd.n5444 gnd.n1554 240.244
R5461 gnd.n5450 gnd.n1554 240.244
R5462 gnd.n5450 gnd.n1537 240.244
R5463 gnd.n5491 gnd.n1537 240.244
R5464 gnd.n5491 gnd.n1533 240.244
R5465 gnd.n5497 gnd.n1533 240.244
R5466 gnd.n5497 gnd.n1510 240.244
R5467 gnd.n5523 gnd.n1510 240.244
R5468 gnd.n5523 gnd.n1506 240.244
R5469 gnd.n5529 gnd.n1506 240.244
R5470 gnd.n5529 gnd.n1488 240.244
R5471 gnd.n5569 gnd.n1488 240.244
R5472 gnd.n5569 gnd.n1484 240.244
R5473 gnd.n5575 gnd.n1484 240.244
R5474 gnd.n5575 gnd.n1401 240.244
R5475 gnd.n5717 gnd.n1401 240.244
R5476 gnd.n5717 gnd.n1397 240.244
R5477 gnd.n5723 gnd.n1397 240.244
R5478 gnd.n5723 gnd.n1386 240.244
R5479 gnd.n5736 gnd.n1386 240.244
R5480 gnd.n5736 gnd.n1382 240.244
R5481 gnd.n5742 gnd.n1382 240.244
R5482 gnd.n5742 gnd.n1372 240.244
R5483 gnd.n5755 gnd.n1372 240.244
R5484 gnd.n5755 gnd.n1368 240.244
R5485 gnd.n5761 gnd.n1368 240.244
R5486 gnd.n5761 gnd.n1358 240.244
R5487 gnd.n5774 gnd.n1358 240.244
R5488 gnd.n5774 gnd.n1354 240.244
R5489 gnd.n5780 gnd.n1354 240.244
R5490 gnd.n5780 gnd.n1344 240.244
R5491 gnd.n5793 gnd.n1344 240.244
R5492 gnd.n5793 gnd.n1340 240.244
R5493 gnd.n5799 gnd.n1340 240.244
R5494 gnd.n5799 gnd.n1330 240.244
R5495 gnd.n5812 gnd.n1330 240.244
R5496 gnd.n5812 gnd.n1325 240.244
R5497 gnd.n5991 gnd.n1325 240.244
R5498 gnd.n5991 gnd.n1326 240.244
R5499 gnd.n5987 gnd.n1326 240.244
R5500 gnd.n5987 gnd.n5986 240.244
R5501 gnd.n5986 gnd.n5820 240.244
R5502 gnd.n5981 gnd.n5820 240.244
R5503 gnd.n5981 gnd.n5840 240.244
R5504 gnd.n5977 gnd.n5840 240.244
R5505 gnd.n5977 gnd.n5976 240.244
R5506 gnd.n5976 gnd.n5975 240.244
R5507 gnd.n5975 gnd.n5848 240.244
R5508 gnd.n5927 gnd.n5848 240.244
R5509 gnd.n5927 gnd.n5926 240.244
R5510 gnd.n5926 gnd.n5925 240.244
R5511 gnd.n5925 gnd.n5854 240.244
R5512 gnd.n5921 gnd.n5854 240.244
R5513 gnd.n5921 gnd.n5920 240.244
R5514 gnd.n5920 gnd.n5919 240.244
R5515 gnd.n5919 gnd.n5860 240.244
R5516 gnd.n5886 gnd.n5860 240.244
R5517 gnd.n5905 gnd.n5886 240.244
R5518 gnd.n5905 gnd.n5887 240.244
R5519 gnd.n5901 gnd.n5887 240.244
R5520 gnd.n5901 gnd.n5900 240.244
R5521 gnd.n5900 gnd.n614 240.244
R5522 gnd.n6926 gnd.n614 240.244
R5523 gnd.n6926 gnd.n615 240.244
R5524 gnd.n6922 gnd.n615 240.244
R5525 gnd.n6922 gnd.n6921 240.244
R5526 gnd.n4284 gnd.n4283 240.244
R5527 gnd.n4526 gnd.n4283 240.244
R5528 gnd.n4524 gnd.n4523 240.244
R5529 gnd.n4520 gnd.n4519 240.244
R5530 gnd.n4516 gnd.n4515 240.244
R5531 gnd.n4512 gnd.n4511 240.244
R5532 gnd.n4508 gnd.n4507 240.244
R5533 gnd.n4504 gnd.n4503 240.244
R5534 gnd.n4500 gnd.n4499 240.244
R5535 gnd.n4496 gnd.n4495 240.244
R5536 gnd.n4492 gnd.n4491 240.244
R5537 gnd.n4488 gnd.n4487 240.244
R5538 gnd.n4484 gnd.n4483 240.244
R5539 gnd.n4480 gnd.n4479 240.244
R5540 gnd.n4476 gnd.n4475 240.244
R5541 gnd.n4472 gnd.n4471 240.244
R5542 gnd.n4468 gnd.n4467 240.244
R5543 gnd.n4464 gnd.n4463 240.244
R5544 gnd.n4460 gnd.n4459 240.244
R5545 gnd.n4456 gnd.n4455 240.244
R5546 gnd.n4452 gnd.n4451 240.244
R5547 gnd.n4448 gnd.n4447 240.244
R5548 gnd.n4444 gnd.n4443 240.244
R5549 gnd.n4440 gnd.n4439 240.244
R5550 gnd.n4436 gnd.n4435 240.244
R5551 gnd.n4432 gnd.n4431 240.244
R5552 gnd.n4428 gnd.n4427 240.244
R5553 gnd.n4424 gnd.n4423 240.244
R5554 gnd.n4420 gnd.n4419 240.244
R5555 gnd.n4416 gnd.n4415 240.244
R5556 gnd.n4412 gnd.n4411 240.244
R5557 gnd.n4408 gnd.n4407 240.244
R5558 gnd.n4404 gnd.n4403 240.244
R5559 gnd.n4400 gnd.n4399 240.244
R5560 gnd.n4396 gnd.n4395 240.244
R5561 gnd.n4392 gnd.n4391 240.244
R5562 gnd.n4388 gnd.n4387 240.244
R5563 gnd.n4384 gnd.n4383 240.244
R5564 gnd.n4380 gnd.n4379 240.244
R5565 gnd.n4376 gnd.n4375 240.244
R5566 gnd.n4372 gnd.n4371 240.244
R5567 gnd.n4368 gnd.n1947 240.244
R5568 gnd.n6248 gnd.n1092 240.244
R5569 gnd.n6246 gnd.n6245 240.244
R5570 gnd.n6243 gnd.n1098 240.244
R5571 gnd.n6239 gnd.n6238 240.244
R5572 gnd.n6236 gnd.n1106 240.244
R5573 gnd.n6232 gnd.n6231 240.244
R5574 gnd.n6229 gnd.n1113 240.244
R5575 gnd.n6225 gnd.n6224 240.244
R5576 gnd.n6220 gnd.n1123 240.244
R5577 gnd.n6216 gnd.n6215 240.244
R5578 gnd.n6213 gnd.n1131 240.244
R5579 gnd.n6209 gnd.n6208 240.244
R5580 gnd.n6206 gnd.n1138 240.244
R5581 gnd.n6202 gnd.n6201 240.244
R5582 gnd.n6199 gnd.n1145 240.244
R5583 gnd.n6195 gnd.n6194 240.244
R5584 gnd.n6192 gnd.n1152 240.244
R5585 gnd.n6188 gnd.n6187 240.244
R5586 gnd.n3872 gnd.n3632 240.244
R5587 gnd.n3872 gnd.n2151 240.244
R5588 gnd.n3877 gnd.n2151 240.244
R5589 gnd.n3877 gnd.n2144 240.244
R5590 gnd.n3880 gnd.n2144 240.244
R5591 gnd.n3880 gnd.n2136 240.244
R5592 gnd.n3885 gnd.n2136 240.244
R5593 gnd.n3885 gnd.n2127 240.244
R5594 gnd.n3888 gnd.n2127 240.244
R5595 gnd.n3888 gnd.n2119 240.244
R5596 gnd.n3893 gnd.n2119 240.244
R5597 gnd.n3893 gnd.n2112 240.244
R5598 gnd.n3896 gnd.n2112 240.244
R5599 gnd.n3896 gnd.n2104 240.244
R5600 gnd.n3901 gnd.n2104 240.244
R5601 gnd.n3901 gnd.n2095 240.244
R5602 gnd.n3904 gnd.n2095 240.244
R5603 gnd.n3904 gnd.n2087 240.244
R5604 gnd.n3909 gnd.n2087 240.244
R5605 gnd.n3909 gnd.n2080 240.244
R5606 gnd.n3912 gnd.n2080 240.244
R5607 gnd.n3912 gnd.n2072 240.244
R5608 gnd.n3917 gnd.n2072 240.244
R5609 gnd.n3917 gnd.n2063 240.244
R5610 gnd.n3920 gnd.n2063 240.244
R5611 gnd.n3920 gnd.n2055 240.244
R5612 gnd.n3925 gnd.n2055 240.244
R5613 gnd.n3925 gnd.n2048 240.244
R5614 gnd.n3928 gnd.n2048 240.244
R5615 gnd.n3928 gnd.n2040 240.244
R5616 gnd.n3933 gnd.n2040 240.244
R5617 gnd.n3933 gnd.n2030 240.244
R5618 gnd.n3937 gnd.n2030 240.244
R5619 gnd.n3937 gnd.n2021 240.244
R5620 gnd.n3940 gnd.n2021 240.244
R5621 gnd.n3940 gnd.n2014 240.244
R5622 gnd.n3945 gnd.n2014 240.244
R5623 gnd.n3945 gnd.n2007 240.244
R5624 gnd.n3948 gnd.n2007 240.244
R5625 gnd.n3948 gnd.n1997 240.244
R5626 gnd.n3953 gnd.n1997 240.244
R5627 gnd.n3953 gnd.n1988 240.244
R5628 gnd.n3956 gnd.n1988 240.244
R5629 gnd.n3956 gnd.n981 240.244
R5630 gnd.n3963 gnd.n981 240.244
R5631 gnd.n3963 gnd.n994 240.244
R5632 gnd.n3968 gnd.n994 240.244
R5633 gnd.n3968 gnd.n1005 240.244
R5634 gnd.n3979 gnd.n1005 240.244
R5635 gnd.n3979 gnd.n1016 240.244
R5636 gnd.n1936 gnd.n1016 240.244
R5637 gnd.n1936 gnd.n1026 240.244
R5638 gnd.n4572 gnd.n1026 240.244
R5639 gnd.n4572 gnd.n1037 240.244
R5640 gnd.n1919 gnd.n1037 240.244
R5641 gnd.n1919 gnd.n1047 240.244
R5642 gnd.n4580 gnd.n1047 240.244
R5643 gnd.n4580 gnd.n1058 240.244
R5644 gnd.n4584 gnd.n1058 240.244
R5645 gnd.n4584 gnd.n1069 240.244
R5646 gnd.n4591 gnd.n1069 240.244
R5647 gnd.n4591 gnd.n1080 240.244
R5648 gnd.n6179 gnd.n1080 240.244
R5649 gnd.n6179 gnd.n1089 240.244
R5650 gnd.n3775 gnd.n3771 240.244
R5651 gnd.n3781 gnd.n3771 240.244
R5652 gnd.n3785 gnd.n3783 240.244
R5653 gnd.n3791 gnd.n3767 240.244
R5654 gnd.n3795 gnd.n3793 240.244
R5655 gnd.n3801 gnd.n3763 240.244
R5656 gnd.n3805 gnd.n3803 240.244
R5657 gnd.n3811 gnd.n3759 240.244
R5658 gnd.n3815 gnd.n3813 240.244
R5659 gnd.n3821 gnd.n3752 240.244
R5660 gnd.n3825 gnd.n3823 240.244
R5661 gnd.n3831 gnd.n3748 240.244
R5662 gnd.n3835 gnd.n3833 240.244
R5663 gnd.n3841 gnd.n3744 240.244
R5664 gnd.n3845 gnd.n3843 240.244
R5665 gnd.n3851 gnd.n3740 240.244
R5666 gnd.n3855 gnd.n3853 240.244
R5667 gnd.n3862 gnd.n3736 240.244
R5668 gnd.n3865 gnd.n3864 240.244
R5669 gnd.n4104 gnd.n2153 240.244
R5670 gnd.n4110 gnd.n2153 240.244
R5671 gnd.n4110 gnd.n2142 240.244
R5672 gnd.n4120 gnd.n2142 240.244
R5673 gnd.n4120 gnd.n2138 240.244
R5674 gnd.n4126 gnd.n2138 240.244
R5675 gnd.n4126 gnd.n2125 240.244
R5676 gnd.n4136 gnd.n2125 240.244
R5677 gnd.n4136 gnd.n2121 240.244
R5678 gnd.n4142 gnd.n2121 240.244
R5679 gnd.n4142 gnd.n2110 240.244
R5680 gnd.n4152 gnd.n2110 240.244
R5681 gnd.n4152 gnd.n2106 240.244
R5682 gnd.n4158 gnd.n2106 240.244
R5683 gnd.n4158 gnd.n2093 240.244
R5684 gnd.n4168 gnd.n2093 240.244
R5685 gnd.n4168 gnd.n2089 240.244
R5686 gnd.n4174 gnd.n2089 240.244
R5687 gnd.n4174 gnd.n2078 240.244
R5688 gnd.n4184 gnd.n2078 240.244
R5689 gnd.n4184 gnd.n2074 240.244
R5690 gnd.n4190 gnd.n2074 240.244
R5691 gnd.n4190 gnd.n2061 240.244
R5692 gnd.n4200 gnd.n2061 240.244
R5693 gnd.n4200 gnd.n2057 240.244
R5694 gnd.n4206 gnd.n2057 240.244
R5695 gnd.n4206 gnd.n2046 240.244
R5696 gnd.n4216 gnd.n2046 240.244
R5697 gnd.n4216 gnd.n2042 240.244
R5698 gnd.n4222 gnd.n2042 240.244
R5699 gnd.n4222 gnd.n2028 240.244
R5700 gnd.n4232 gnd.n2028 240.244
R5701 gnd.n4232 gnd.n2024 240.244
R5702 gnd.n4238 gnd.n2024 240.244
R5703 gnd.n4238 gnd.n2013 240.244
R5704 gnd.n4248 gnd.n2013 240.244
R5705 gnd.n4248 gnd.n2009 240.244
R5706 gnd.n4254 gnd.n2009 240.244
R5707 gnd.n4254 gnd.n1995 240.244
R5708 gnd.n4274 gnd.n1995 240.244
R5709 gnd.n4274 gnd.n1991 240.244
R5710 gnd.n4281 gnd.n1991 240.244
R5711 gnd.n4281 gnd.n985 240.244
R5712 gnd.n6314 gnd.n985 240.244
R5713 gnd.n6314 gnd.n986 240.244
R5714 gnd.n6310 gnd.n986 240.244
R5715 gnd.n6310 gnd.n992 240.244
R5716 gnd.n6302 gnd.n992 240.244
R5717 gnd.n6302 gnd.n1008 240.244
R5718 gnd.n6298 gnd.n1008 240.244
R5719 gnd.n6298 gnd.n1014 240.244
R5720 gnd.n6290 gnd.n1014 240.244
R5721 gnd.n6290 gnd.n1029 240.244
R5722 gnd.n6286 gnd.n1029 240.244
R5723 gnd.n6286 gnd.n1035 240.244
R5724 gnd.n6278 gnd.n1035 240.244
R5725 gnd.n6278 gnd.n1050 240.244
R5726 gnd.n6274 gnd.n1050 240.244
R5727 gnd.n6274 gnd.n1056 240.244
R5728 gnd.n6266 gnd.n1056 240.244
R5729 gnd.n6266 gnd.n1072 240.244
R5730 gnd.n6262 gnd.n1072 240.244
R5731 gnd.n6262 gnd.n1078 240.244
R5732 gnd.n6254 gnd.n1078 240.244
R5733 gnd.n3629 gnd.n2181 240.244
R5734 gnd.n3622 gnd.n3621 240.244
R5735 gnd.n3619 gnd.n3618 240.244
R5736 gnd.n3615 gnd.n3614 240.244
R5737 gnd.n3611 gnd.n3610 240.244
R5738 gnd.n3607 gnd.n3606 240.244
R5739 gnd.n3603 gnd.n3602 240.244
R5740 gnd.n3599 gnd.n3598 240.244
R5741 gnd.n2873 gnd.n2585 240.244
R5742 gnd.n2883 gnd.n2585 240.244
R5743 gnd.n2883 gnd.n2576 240.244
R5744 gnd.n2576 gnd.n2565 240.244
R5745 gnd.n2904 gnd.n2565 240.244
R5746 gnd.n2904 gnd.n2559 240.244
R5747 gnd.n2914 gnd.n2559 240.244
R5748 gnd.n2914 gnd.n2548 240.244
R5749 gnd.n2548 gnd.n2540 240.244
R5750 gnd.n2932 gnd.n2540 240.244
R5751 gnd.n2933 gnd.n2932 240.244
R5752 gnd.n2933 gnd.n2525 240.244
R5753 gnd.n2935 gnd.n2525 240.244
R5754 gnd.n2935 gnd.n2511 240.244
R5755 gnd.n2977 gnd.n2511 240.244
R5756 gnd.n2978 gnd.n2977 240.244
R5757 gnd.n2981 gnd.n2978 240.244
R5758 gnd.n2981 gnd.n2466 240.244
R5759 gnd.n2506 gnd.n2466 240.244
R5760 gnd.n2506 gnd.n2476 240.244
R5761 gnd.n2991 gnd.n2476 240.244
R5762 gnd.n2991 gnd.n2497 240.244
R5763 gnd.n3001 gnd.n2497 240.244
R5764 gnd.n3001 gnd.n2383 240.244
R5765 gnd.n3046 gnd.n2383 240.244
R5766 gnd.n3046 gnd.n2369 240.244
R5767 gnd.n3068 gnd.n2369 240.244
R5768 gnd.n3069 gnd.n3068 240.244
R5769 gnd.n3069 gnd.n2356 240.244
R5770 gnd.n2356 gnd.n2345 240.244
R5771 gnd.n3100 gnd.n2345 240.244
R5772 gnd.n3101 gnd.n3100 240.244
R5773 gnd.n3102 gnd.n3101 240.244
R5774 gnd.n3102 gnd.n2330 240.244
R5775 gnd.n2330 gnd.n2329 240.244
R5776 gnd.n2329 gnd.n2314 240.244
R5777 gnd.n3153 gnd.n2314 240.244
R5778 gnd.n3154 gnd.n3153 240.244
R5779 gnd.n3154 gnd.n2301 240.244
R5780 gnd.n2301 gnd.n2290 240.244
R5781 gnd.n3185 gnd.n2290 240.244
R5782 gnd.n3186 gnd.n3185 240.244
R5783 gnd.n3187 gnd.n3186 240.244
R5784 gnd.n3187 gnd.n2274 240.244
R5785 gnd.n2274 gnd.n2273 240.244
R5786 gnd.n2273 gnd.n2260 240.244
R5787 gnd.n3242 gnd.n2260 240.244
R5788 gnd.n3243 gnd.n3242 240.244
R5789 gnd.n3243 gnd.n2247 240.244
R5790 gnd.n2247 gnd.n2237 240.244
R5791 gnd.n3530 gnd.n2237 240.244
R5792 gnd.n3533 gnd.n3530 240.244
R5793 gnd.n3533 gnd.n3532 240.244
R5794 gnd.n2863 gnd.n2598 240.244
R5795 gnd.n2619 gnd.n2598 240.244
R5796 gnd.n2622 gnd.n2621 240.244
R5797 gnd.n2629 gnd.n2628 240.244
R5798 gnd.n2632 gnd.n2631 240.244
R5799 gnd.n2639 gnd.n2638 240.244
R5800 gnd.n2642 gnd.n2641 240.244
R5801 gnd.n2649 gnd.n2648 240.244
R5802 gnd.n2871 gnd.n2595 240.244
R5803 gnd.n2595 gnd.n2574 240.244
R5804 gnd.n2894 gnd.n2574 240.244
R5805 gnd.n2894 gnd.n2568 240.244
R5806 gnd.n2902 gnd.n2568 240.244
R5807 gnd.n2902 gnd.n2570 240.244
R5808 gnd.n2570 gnd.n2546 240.244
R5809 gnd.n2924 gnd.n2546 240.244
R5810 gnd.n2924 gnd.n2542 240.244
R5811 gnd.n2930 gnd.n2542 240.244
R5812 gnd.n2930 gnd.n2524 240.244
R5813 gnd.n2955 gnd.n2524 240.244
R5814 gnd.n2955 gnd.n2519 240.244
R5815 gnd.n2967 gnd.n2519 240.244
R5816 gnd.n2967 gnd.n2520 240.244
R5817 gnd.n2963 gnd.n2520 240.244
R5818 gnd.n2963 gnd.n2468 240.244
R5819 gnd.n3015 gnd.n2468 240.244
R5820 gnd.n3015 gnd.n2469 240.244
R5821 gnd.n3011 gnd.n2469 240.244
R5822 gnd.n3011 gnd.n2475 240.244
R5823 gnd.n2495 gnd.n2475 240.244
R5824 gnd.n2495 gnd.n2381 240.244
R5825 gnd.n3050 gnd.n2381 240.244
R5826 gnd.n3050 gnd.n2376 240.244
R5827 gnd.n3058 gnd.n2376 240.244
R5828 gnd.n3058 gnd.n2377 240.244
R5829 gnd.n2377 gnd.n2354 240.244
R5830 gnd.n3090 gnd.n2354 240.244
R5831 gnd.n3090 gnd.n2349 240.244
R5832 gnd.n3098 gnd.n2349 240.244
R5833 gnd.n3098 gnd.n2350 240.244
R5834 gnd.n2350 gnd.n2327 240.244
R5835 gnd.n3135 gnd.n2327 240.244
R5836 gnd.n3135 gnd.n2322 240.244
R5837 gnd.n3143 gnd.n2322 240.244
R5838 gnd.n3143 gnd.n2323 240.244
R5839 gnd.n2323 gnd.n2299 240.244
R5840 gnd.n3175 gnd.n2299 240.244
R5841 gnd.n3175 gnd.n2294 240.244
R5842 gnd.n3183 gnd.n2294 240.244
R5843 gnd.n3183 gnd.n2295 240.244
R5844 gnd.n2295 gnd.n2272 240.244
R5845 gnd.n3224 gnd.n2272 240.244
R5846 gnd.n3224 gnd.n2267 240.244
R5847 gnd.n3232 gnd.n2267 240.244
R5848 gnd.n3232 gnd.n2268 240.244
R5849 gnd.n2268 gnd.n2245 240.244
R5850 gnd.n3518 gnd.n2245 240.244
R5851 gnd.n3518 gnd.n2240 240.244
R5852 gnd.n3528 gnd.n2240 240.244
R5853 gnd.n3528 gnd.n2241 240.244
R5854 gnd.n2241 gnd.n2180 240.244
R5855 gnd.n2200 gnd.n2158 240.244
R5856 gnd.n3589 gnd.n3588 240.244
R5857 gnd.n3585 gnd.n3584 240.244
R5858 gnd.n3581 gnd.n3580 240.244
R5859 gnd.n3577 gnd.n3576 240.244
R5860 gnd.n3573 gnd.n3572 240.244
R5861 gnd.n3569 gnd.n3568 240.244
R5862 gnd.n3565 gnd.n3564 240.244
R5863 gnd.n3561 gnd.n3560 240.244
R5864 gnd.n3557 gnd.n3556 240.244
R5865 gnd.n3553 gnd.n3552 240.244
R5866 gnd.n3549 gnd.n3548 240.244
R5867 gnd.n3545 gnd.n3544 240.244
R5868 gnd.n2786 gnd.n2683 240.244
R5869 gnd.n2786 gnd.n2676 240.244
R5870 gnd.n2797 gnd.n2676 240.244
R5871 gnd.n2797 gnd.n2672 240.244
R5872 gnd.n2803 gnd.n2672 240.244
R5873 gnd.n2803 gnd.n2664 240.244
R5874 gnd.n2813 gnd.n2664 240.244
R5875 gnd.n2813 gnd.n2659 240.244
R5876 gnd.n2849 gnd.n2659 240.244
R5877 gnd.n2849 gnd.n2660 240.244
R5878 gnd.n2660 gnd.n2607 240.244
R5879 gnd.n2844 gnd.n2607 240.244
R5880 gnd.n2844 gnd.n2843 240.244
R5881 gnd.n2843 gnd.n2586 240.244
R5882 gnd.n2839 gnd.n2586 240.244
R5883 gnd.n2839 gnd.n2577 240.244
R5884 gnd.n2836 gnd.n2577 240.244
R5885 gnd.n2836 gnd.n2835 240.244
R5886 gnd.n2835 gnd.n2560 240.244
R5887 gnd.n2831 gnd.n2560 240.244
R5888 gnd.n2831 gnd.n2549 240.244
R5889 gnd.n2549 gnd.n2530 240.244
R5890 gnd.n2944 gnd.n2530 240.244
R5891 gnd.n2944 gnd.n2526 240.244
R5892 gnd.n2952 gnd.n2526 240.244
R5893 gnd.n2952 gnd.n2517 240.244
R5894 gnd.n2517 gnd.n2453 240.244
R5895 gnd.n3024 gnd.n2453 240.244
R5896 gnd.n3024 gnd.n2454 240.244
R5897 gnd.n2465 gnd.n2454 240.244
R5898 gnd.n2500 gnd.n2465 240.244
R5899 gnd.n2503 gnd.n2500 240.244
R5900 gnd.n2503 gnd.n2477 240.244
R5901 gnd.n2490 gnd.n2477 240.244
R5902 gnd.n2490 gnd.n2487 240.244
R5903 gnd.n2487 gnd.n2384 240.244
R5904 gnd.n3045 gnd.n2384 240.244
R5905 gnd.n3045 gnd.n2374 240.244
R5906 gnd.n3041 gnd.n2374 240.244
R5907 gnd.n3041 gnd.n2368 240.244
R5908 gnd.n3038 gnd.n2368 240.244
R5909 gnd.n3038 gnd.n2357 240.244
R5910 gnd.n3035 gnd.n2357 240.244
R5911 gnd.n3035 gnd.n2335 240.244
R5912 gnd.n3111 gnd.n2335 240.244
R5913 gnd.n3111 gnd.n2331 240.244
R5914 gnd.n3132 gnd.n2331 240.244
R5915 gnd.n3132 gnd.n2320 240.244
R5916 gnd.n3128 gnd.n2320 240.244
R5917 gnd.n3128 gnd.n2313 240.244
R5918 gnd.n3125 gnd.n2313 240.244
R5919 gnd.n3125 gnd.n2302 240.244
R5920 gnd.n3122 gnd.n2302 240.244
R5921 gnd.n3122 gnd.n2279 240.244
R5922 gnd.n3196 gnd.n2279 240.244
R5923 gnd.n3196 gnd.n2275 240.244
R5924 gnd.n3221 gnd.n2275 240.244
R5925 gnd.n3221 gnd.n2266 240.244
R5926 gnd.n3217 gnd.n2266 240.244
R5927 gnd.n3217 gnd.n2259 240.244
R5928 gnd.n3213 gnd.n2259 240.244
R5929 gnd.n3213 gnd.n2248 240.244
R5930 gnd.n3210 gnd.n2248 240.244
R5931 gnd.n3210 gnd.n2229 240.244
R5932 gnd.n3540 gnd.n2229 240.244
R5933 gnd.n2700 gnd.n2699 240.244
R5934 gnd.n2771 gnd.n2699 240.244
R5935 gnd.n2769 gnd.n2768 240.244
R5936 gnd.n2765 gnd.n2764 240.244
R5937 gnd.n2761 gnd.n2760 240.244
R5938 gnd.n2757 gnd.n2756 240.244
R5939 gnd.n2753 gnd.n2752 240.244
R5940 gnd.n2749 gnd.n2748 240.244
R5941 gnd.n2745 gnd.n2744 240.244
R5942 gnd.n2741 gnd.n2740 240.244
R5943 gnd.n2737 gnd.n2736 240.244
R5944 gnd.n2733 gnd.n2732 240.244
R5945 gnd.n2729 gnd.n2687 240.244
R5946 gnd.n2789 gnd.n2681 240.244
R5947 gnd.n2789 gnd.n2677 240.244
R5948 gnd.n2795 gnd.n2677 240.244
R5949 gnd.n2795 gnd.n2670 240.244
R5950 gnd.n2805 gnd.n2670 240.244
R5951 gnd.n2805 gnd.n2666 240.244
R5952 gnd.n2811 gnd.n2666 240.244
R5953 gnd.n2811 gnd.n2657 240.244
R5954 gnd.n2851 gnd.n2657 240.244
R5955 gnd.n2851 gnd.n2608 240.244
R5956 gnd.n2859 gnd.n2608 240.244
R5957 gnd.n2859 gnd.n2609 240.244
R5958 gnd.n2609 gnd.n2587 240.244
R5959 gnd.n2880 gnd.n2587 240.244
R5960 gnd.n2880 gnd.n2579 240.244
R5961 gnd.n2891 gnd.n2579 240.244
R5962 gnd.n2891 gnd.n2580 240.244
R5963 gnd.n2580 gnd.n2561 240.244
R5964 gnd.n2911 gnd.n2561 240.244
R5965 gnd.n2911 gnd.n2551 240.244
R5966 gnd.n2921 gnd.n2551 240.244
R5967 gnd.n2921 gnd.n2532 240.244
R5968 gnd.n2942 gnd.n2532 240.244
R5969 gnd.n2942 gnd.n2534 240.244
R5970 gnd.n2534 gnd.n2515 240.244
R5971 gnd.n2970 gnd.n2515 240.244
R5972 gnd.n2970 gnd.n2457 240.244
R5973 gnd.n3022 gnd.n2457 240.244
R5974 gnd.n3022 gnd.n2458 240.244
R5975 gnd.n3018 gnd.n2458 240.244
R5976 gnd.n3018 gnd.n2464 240.244
R5977 gnd.n2479 gnd.n2464 240.244
R5978 gnd.n3008 gnd.n2479 240.244
R5979 gnd.n3008 gnd.n2480 240.244
R5980 gnd.n3004 gnd.n2480 240.244
R5981 gnd.n3004 gnd.n2486 240.244
R5982 gnd.n2486 gnd.n2373 240.244
R5983 gnd.n3061 gnd.n2373 240.244
R5984 gnd.n3061 gnd.n2366 240.244
R5985 gnd.n3072 gnd.n2366 240.244
R5986 gnd.n3072 gnd.n2359 240.244
R5987 gnd.n3087 gnd.n2359 240.244
R5988 gnd.n3087 gnd.n2360 240.244
R5989 gnd.n2360 gnd.n2338 240.244
R5990 gnd.n3109 gnd.n2338 240.244
R5991 gnd.n3109 gnd.n2339 240.244
R5992 gnd.n2339 gnd.n2318 240.244
R5993 gnd.n3146 gnd.n2318 240.244
R5994 gnd.n3146 gnd.n2311 240.244
R5995 gnd.n3157 gnd.n2311 240.244
R5996 gnd.n3157 gnd.n2304 240.244
R5997 gnd.n3172 gnd.n2304 240.244
R5998 gnd.n3172 gnd.n2305 240.244
R5999 gnd.n2305 gnd.n2282 240.244
R6000 gnd.n3194 gnd.n2282 240.244
R6001 gnd.n3194 gnd.n2284 240.244
R6002 gnd.n2284 gnd.n2264 240.244
R6003 gnd.n3235 gnd.n2264 240.244
R6004 gnd.n3235 gnd.n2257 240.244
R6005 gnd.n3246 gnd.n2257 240.244
R6006 gnd.n3246 gnd.n2250 240.244
R6007 gnd.n3515 gnd.n2250 240.244
R6008 gnd.n3515 gnd.n2251 240.244
R6009 gnd.n2251 gnd.n2232 240.244
R6010 gnd.n3538 gnd.n2232 240.244
R6011 gnd.n4662 gnd.n1087 240.244
R6012 gnd.n4665 gnd.n4664 240.244
R6013 gnd.n4675 gnd.n4667 240.244
R6014 gnd.n4678 gnd.n4677 240.244
R6015 gnd.n4687 gnd.n4686 240.244
R6016 gnd.n4698 gnd.n4689 240.244
R6017 gnd.n4701 gnd.n4700 240.244
R6018 gnd.n4710 gnd.n4709 240.244
R6019 gnd.n4721 gnd.n4712 240.244
R6020 gnd.n4055 gnd.n3633 240.244
R6021 gnd.n4055 gnd.n2152 240.244
R6022 gnd.n4052 gnd.n2152 240.244
R6023 gnd.n4052 gnd.n2145 240.244
R6024 gnd.n4049 gnd.n2145 240.244
R6025 gnd.n4049 gnd.n2137 240.244
R6026 gnd.n4046 gnd.n2137 240.244
R6027 gnd.n4046 gnd.n2128 240.244
R6028 gnd.n4043 gnd.n2128 240.244
R6029 gnd.n4043 gnd.n2120 240.244
R6030 gnd.n4040 gnd.n2120 240.244
R6031 gnd.n4040 gnd.n2113 240.244
R6032 gnd.n4037 gnd.n2113 240.244
R6033 gnd.n4037 gnd.n2105 240.244
R6034 gnd.n4034 gnd.n2105 240.244
R6035 gnd.n4034 gnd.n2096 240.244
R6036 gnd.n4031 gnd.n2096 240.244
R6037 gnd.n4031 gnd.n2088 240.244
R6038 gnd.n4028 gnd.n2088 240.244
R6039 gnd.n4028 gnd.n2081 240.244
R6040 gnd.n4025 gnd.n2081 240.244
R6041 gnd.n4025 gnd.n2073 240.244
R6042 gnd.n4022 gnd.n2073 240.244
R6043 gnd.n4022 gnd.n2064 240.244
R6044 gnd.n4019 gnd.n2064 240.244
R6045 gnd.n4019 gnd.n2056 240.244
R6046 gnd.n4016 gnd.n2056 240.244
R6047 gnd.n4016 gnd.n2049 240.244
R6048 gnd.n4013 gnd.n2049 240.244
R6049 gnd.n4013 gnd.n2041 240.244
R6050 gnd.n4010 gnd.n2041 240.244
R6051 gnd.n4010 gnd.n2031 240.244
R6052 gnd.n3693 gnd.n2031 240.244
R6053 gnd.n3693 gnd.n2022 240.244
R6054 gnd.n3696 gnd.n2022 240.244
R6055 gnd.n3696 gnd.n2015 240.244
R6056 gnd.n3697 gnd.n2015 240.244
R6057 gnd.n3697 gnd.n2008 240.244
R6058 gnd.n3700 gnd.n2008 240.244
R6059 gnd.n3700 gnd.n1998 240.244
R6060 gnd.n3701 gnd.n1998 240.244
R6061 gnd.n3701 gnd.n1989 240.244
R6062 gnd.n3704 gnd.n1989 240.244
R6063 gnd.n3704 gnd.n982 240.244
R6064 gnd.n3961 gnd.n982 240.244
R6065 gnd.n3961 gnd.n995 240.244
R6066 gnd.n3707 gnd.n995 240.244
R6067 gnd.n3707 gnd.n1006 240.244
R6068 gnd.n3981 gnd.n1006 240.244
R6069 gnd.n3981 gnd.n1017 240.244
R6070 gnd.n4564 gnd.n1017 240.244
R6071 gnd.n4564 gnd.n1027 240.244
R6072 gnd.n4570 gnd.n1027 240.244
R6073 gnd.n4570 gnd.n1038 240.244
R6074 gnd.n4605 gnd.n1038 240.244
R6075 gnd.n4605 gnd.n1048 240.244
R6076 gnd.n1924 gnd.n1048 240.244
R6077 gnd.n1924 gnd.n1059 240.244
R6078 gnd.n1925 gnd.n1059 240.244
R6079 gnd.n1925 gnd.n1070 240.244
R6080 gnd.n4593 gnd.n1070 240.244
R6081 gnd.n4593 gnd.n1081 240.244
R6082 gnd.n6177 gnd.n1081 240.244
R6083 gnd.n6177 gnd.n1090 240.244
R6084 gnd.n4096 gnd.n4094 240.244
R6085 gnd.n4092 gnd.n3638 240.244
R6086 gnd.n4088 gnd.n4086 240.244
R6087 gnd.n4084 gnd.n3644 240.244
R6088 gnd.n4080 gnd.n4078 240.244
R6089 gnd.n4076 gnd.n3650 240.244
R6090 gnd.n4072 gnd.n4070 240.244
R6091 gnd.n4068 gnd.n3656 240.244
R6092 gnd.n4061 gnd.n4060 240.244
R6093 gnd.n4102 gnd.n2150 240.244
R6094 gnd.n4112 gnd.n2150 240.244
R6095 gnd.n4112 gnd.n2146 240.244
R6096 gnd.n4118 gnd.n2146 240.244
R6097 gnd.n4118 gnd.n2134 240.244
R6098 gnd.n4128 gnd.n2134 240.244
R6099 gnd.n4128 gnd.n2130 240.244
R6100 gnd.n4134 gnd.n2130 240.244
R6101 gnd.n4134 gnd.n2118 240.244
R6102 gnd.n4144 gnd.n2118 240.244
R6103 gnd.n4144 gnd.n2114 240.244
R6104 gnd.n4150 gnd.n2114 240.244
R6105 gnd.n4150 gnd.n2102 240.244
R6106 gnd.n4160 gnd.n2102 240.244
R6107 gnd.n4160 gnd.n2098 240.244
R6108 gnd.n4166 gnd.n2098 240.244
R6109 gnd.n4166 gnd.n2086 240.244
R6110 gnd.n4176 gnd.n2086 240.244
R6111 gnd.n4176 gnd.n2082 240.244
R6112 gnd.n4182 gnd.n2082 240.244
R6113 gnd.n4182 gnd.n2070 240.244
R6114 gnd.n4192 gnd.n2070 240.244
R6115 gnd.n4192 gnd.n2066 240.244
R6116 gnd.n4198 gnd.n2066 240.244
R6117 gnd.n4198 gnd.n2054 240.244
R6118 gnd.n4208 gnd.n2054 240.244
R6119 gnd.n4208 gnd.n2050 240.244
R6120 gnd.n4214 gnd.n2050 240.244
R6121 gnd.n4214 gnd.n2038 240.244
R6122 gnd.n4224 gnd.n2038 240.244
R6123 gnd.n4224 gnd.n2033 240.244
R6124 gnd.n4230 gnd.n2033 240.244
R6125 gnd.n4230 gnd.n2020 240.244
R6126 gnd.n4240 gnd.n2020 240.244
R6127 gnd.n4240 gnd.n2016 240.244
R6128 gnd.n4246 gnd.n2016 240.244
R6129 gnd.n4246 gnd.n2005 240.244
R6130 gnd.n4256 gnd.n2005 240.244
R6131 gnd.n4256 gnd.n2000 240.244
R6132 gnd.n4272 gnd.n2000 240.244
R6133 gnd.n4272 gnd.n2001 240.244
R6134 gnd.n2001 gnd.n1990 240.244
R6135 gnd.n4267 gnd.n1990 240.244
R6136 gnd.n4267 gnd.n984 240.244
R6137 gnd.n996 gnd.n984 240.244
R6138 gnd.n6308 gnd.n996 240.244
R6139 gnd.n6308 gnd.n997 240.244
R6140 gnd.n6304 gnd.n997 240.244
R6141 gnd.n6304 gnd.n1003 240.244
R6142 gnd.n6296 gnd.n1003 240.244
R6143 gnd.n6296 gnd.n1019 240.244
R6144 gnd.n6292 gnd.n1019 240.244
R6145 gnd.n6292 gnd.n1025 240.244
R6146 gnd.n6284 gnd.n1025 240.244
R6147 gnd.n6284 gnd.n1039 240.244
R6148 gnd.n6280 gnd.n1039 240.244
R6149 gnd.n6280 gnd.n1045 240.244
R6150 gnd.n6272 gnd.n1045 240.244
R6151 gnd.n6272 gnd.n1061 240.244
R6152 gnd.n6268 gnd.n1061 240.244
R6153 gnd.n6268 gnd.n1067 240.244
R6154 gnd.n6260 gnd.n1067 240.244
R6155 gnd.n6260 gnd.n1082 240.244
R6156 gnd.n6256 gnd.n1082 240.244
R6157 gnd.n4784 gnd.n1897 240.244
R6158 gnd.n4784 gnd.n1893 240.244
R6159 gnd.n4790 gnd.n1893 240.244
R6160 gnd.n4790 gnd.n1883 240.244
R6161 gnd.n4803 gnd.n1883 240.244
R6162 gnd.n4803 gnd.n1879 240.244
R6163 gnd.n4809 gnd.n1879 240.244
R6164 gnd.n4809 gnd.n1869 240.244
R6165 gnd.n4822 gnd.n1869 240.244
R6166 gnd.n4822 gnd.n1865 240.244
R6167 gnd.n4828 gnd.n1865 240.244
R6168 gnd.n4828 gnd.n1855 240.244
R6169 gnd.n4841 gnd.n1855 240.244
R6170 gnd.n4841 gnd.n1851 240.244
R6171 gnd.n4847 gnd.n1851 240.244
R6172 gnd.n4847 gnd.n1841 240.244
R6173 gnd.n4860 gnd.n1841 240.244
R6174 gnd.n4860 gnd.n1837 240.244
R6175 gnd.n4866 gnd.n1837 240.244
R6176 gnd.n4866 gnd.n1827 240.244
R6177 gnd.n5079 gnd.n1827 240.244
R6178 gnd.n5079 gnd.n1823 240.244
R6179 gnd.n5085 gnd.n1823 240.244
R6180 gnd.n5085 gnd.n1761 240.244
R6181 gnd.n5113 gnd.n1761 240.244
R6182 gnd.n5113 gnd.n1755 240.244
R6183 gnd.n5120 gnd.n1755 240.244
R6184 gnd.n5120 gnd.n1756 240.244
R6185 gnd.n1756 gnd.n1732 240.244
R6186 gnd.n5149 gnd.n1732 240.244
R6187 gnd.n5149 gnd.n1728 240.244
R6188 gnd.n5155 gnd.n1728 240.244
R6189 gnd.n5155 gnd.n1712 240.244
R6190 gnd.n5176 gnd.n1712 240.244
R6191 gnd.n5176 gnd.n1706 240.244
R6192 gnd.n5183 gnd.n1706 240.244
R6193 gnd.n5183 gnd.n1707 240.244
R6194 gnd.n1707 gnd.n1681 240.244
R6195 gnd.n5214 gnd.n1681 240.244
R6196 gnd.n5214 gnd.n1676 240.244
R6197 gnd.n5221 gnd.n1676 240.244
R6198 gnd.n5221 gnd.n1667 240.244
R6199 gnd.n1667 gnd.n1649 240.244
R6200 gnd.n5267 gnd.n1649 240.244
R6201 gnd.n5267 gnd.n1645 240.244
R6202 gnd.n5273 gnd.n1645 240.244
R6203 gnd.n5273 gnd.n1632 240.244
R6204 gnd.n5310 gnd.n1632 240.244
R6205 gnd.n5310 gnd.n1626 240.244
R6206 gnd.n5323 gnd.n1626 240.244
R6207 gnd.n5323 gnd.n1627 240.244
R6208 gnd.n5315 gnd.n1627 240.244
R6209 gnd.n5316 gnd.n5315 240.244
R6210 gnd.n5316 gnd.n1597 240.244
R6211 gnd.n5378 gnd.n1597 240.244
R6212 gnd.n5378 gnd.n1591 240.244
R6213 gnd.n5388 gnd.n1591 240.244
R6214 gnd.n5388 gnd.n1592 240.244
R6215 gnd.n5382 gnd.n1592 240.244
R6216 gnd.n5382 gnd.n1568 240.244
R6217 gnd.n5430 gnd.n1568 240.244
R6218 gnd.n5430 gnd.n1569 240.244
R6219 gnd.n5424 gnd.n1569 240.244
R6220 gnd.n5424 gnd.n1546 240.244
R6221 gnd.n5480 gnd.n1546 240.244
R6222 gnd.n5480 gnd.n1547 240.244
R6223 gnd.n5474 gnd.n1547 240.244
R6224 gnd.n5474 gnd.n1524 240.244
R6225 gnd.n5507 gnd.n1524 240.244
R6226 gnd.n5507 gnd.n1520 240.244
R6227 gnd.n5513 gnd.n1520 240.244
R6228 gnd.n5513 gnd.n1497 240.244
R6229 gnd.n5559 gnd.n1497 240.244
R6230 gnd.n5559 gnd.n1498 240.244
R6231 gnd.n5546 gnd.n1498 240.244
R6232 gnd.n5548 gnd.n5546 240.244
R6233 gnd.n5550 gnd.n5548 240.244
R6234 gnd.n5550 gnd.n1391 240.244
R6235 gnd.n5726 gnd.n1391 240.244
R6236 gnd.n5726 gnd.n1387 240.244
R6237 gnd.n5732 gnd.n1387 240.244
R6238 gnd.n5732 gnd.n1378 240.244
R6239 gnd.n5745 gnd.n1378 240.244
R6240 gnd.n5745 gnd.n1374 240.244
R6241 gnd.n5751 gnd.n1374 240.244
R6242 gnd.n5751 gnd.n1364 240.244
R6243 gnd.n5764 gnd.n1364 240.244
R6244 gnd.n5764 gnd.n1360 240.244
R6245 gnd.n5770 gnd.n1360 240.244
R6246 gnd.n5770 gnd.n1350 240.244
R6247 gnd.n5783 gnd.n1350 240.244
R6248 gnd.n5783 gnd.n1346 240.244
R6249 gnd.n5789 gnd.n1346 240.244
R6250 gnd.n5789 gnd.n1336 240.244
R6251 gnd.n5802 gnd.n1336 240.244
R6252 gnd.n5802 gnd.n1332 240.244
R6253 gnd.n5808 gnd.n1332 240.244
R6254 gnd.n5808 gnd.n1321 240.244
R6255 gnd.n5994 gnd.n1321 240.244
R6256 gnd.n5994 gnd.n1317 240.244
R6257 gnd.n6000 gnd.n1317 240.244
R6258 gnd.n4651 gnd.n4650 240.244
R6259 gnd.n4670 gnd.n4650 240.244
R6260 gnd.n4672 gnd.n4671 240.244
R6261 gnd.n4682 gnd.n4681 240.244
R6262 gnd.n4693 gnd.n4692 240.244
R6263 gnd.n4695 gnd.n4694 240.244
R6264 gnd.n4705 gnd.n4704 240.244
R6265 gnd.n4718 gnd.n4717 240.244
R6266 gnd.n4720 gnd.n4719 240.244
R6267 gnd.n1172 gnd.n1171 240.244
R6268 gnd.n4644 gnd.n1173 240.244
R6269 gnd.n1177 gnd.n1176 240.244
R6270 gnd.n1183 gnd.n1178 240.244
R6271 gnd.n1185 gnd.n1184 240.244
R6272 gnd.n1189 gnd.n1188 240.244
R6273 gnd.n1190 gnd.n1189 240.244
R6274 gnd.n1891 gnd.n1190 240.244
R6275 gnd.n1891 gnd.n1193 240.244
R6276 gnd.n1194 gnd.n1193 240.244
R6277 gnd.n1195 gnd.n1194 240.244
R6278 gnd.n1877 gnd.n1195 240.244
R6279 gnd.n1877 gnd.n1198 240.244
R6280 gnd.n1199 gnd.n1198 240.244
R6281 gnd.n1200 gnd.n1199 240.244
R6282 gnd.n1863 gnd.n1200 240.244
R6283 gnd.n1863 gnd.n1203 240.244
R6284 gnd.n1204 gnd.n1203 240.244
R6285 gnd.n1205 gnd.n1204 240.244
R6286 gnd.n1849 gnd.n1205 240.244
R6287 gnd.n1849 gnd.n1208 240.244
R6288 gnd.n1209 gnd.n1208 240.244
R6289 gnd.n1210 gnd.n1209 240.244
R6290 gnd.n1834 gnd.n1210 240.244
R6291 gnd.n1834 gnd.n1213 240.244
R6292 gnd.n1214 gnd.n1213 240.244
R6293 gnd.n1215 gnd.n1214 240.244
R6294 gnd.n1822 gnd.n1215 240.244
R6295 gnd.n1822 gnd.n1218 240.244
R6296 gnd.n1219 gnd.n1218 240.244
R6297 gnd.n1220 gnd.n1219 240.244
R6298 gnd.n1753 gnd.n1220 240.244
R6299 gnd.n1753 gnd.n1223 240.244
R6300 gnd.n1224 gnd.n1223 240.244
R6301 gnd.n1225 gnd.n1224 240.244
R6302 gnd.n1797 gnd.n1225 240.244
R6303 gnd.n1797 gnd.n1228 240.244
R6304 gnd.n1229 gnd.n1228 240.244
R6305 gnd.n1230 gnd.n1229 240.244
R6306 gnd.n1702 gnd.n1230 240.244
R6307 gnd.n1702 gnd.n1233 240.244
R6308 gnd.n1234 gnd.n1233 240.244
R6309 gnd.n1235 gnd.n1234 240.244
R6310 gnd.n1682 gnd.n1235 240.244
R6311 gnd.n1682 gnd.n1238 240.244
R6312 gnd.n1239 gnd.n1238 240.244
R6313 gnd.n1240 gnd.n1239 240.244
R6314 gnd.n1657 gnd.n1240 240.244
R6315 gnd.n1657 gnd.n1243 240.244
R6316 gnd.n1244 gnd.n1243 240.244
R6317 gnd.n1245 gnd.n1244 240.244
R6318 gnd.n1641 gnd.n1245 240.244
R6319 gnd.n1641 gnd.n1248 240.244
R6320 gnd.n1249 gnd.n1248 240.244
R6321 gnd.n1250 gnd.n1249 240.244
R6322 gnd.n1617 gnd.n1250 240.244
R6323 gnd.n1617 gnd.n1253 240.244
R6324 gnd.n1254 gnd.n1253 240.244
R6325 gnd.n1255 gnd.n1254 240.244
R6326 gnd.n1599 gnd.n1255 240.244
R6327 gnd.n1599 gnd.n1258 240.244
R6328 gnd.n1259 gnd.n1258 240.244
R6329 gnd.n1260 gnd.n1259 240.244
R6330 gnd.n1575 gnd.n1260 240.244
R6331 gnd.n1575 gnd.n1263 240.244
R6332 gnd.n1264 gnd.n1263 240.244
R6333 gnd.n1265 gnd.n1264 240.244
R6334 gnd.n5422 gnd.n1265 240.244
R6335 gnd.n5422 gnd.n1268 240.244
R6336 gnd.n1269 gnd.n1268 240.244
R6337 gnd.n1270 gnd.n1269 240.244
R6338 gnd.n5472 gnd.n1270 240.244
R6339 gnd.n5472 gnd.n1273 240.244
R6340 gnd.n1274 gnd.n1273 240.244
R6341 gnd.n1275 gnd.n1274 240.244
R6342 gnd.n1519 gnd.n1275 240.244
R6343 gnd.n1519 gnd.n1278 240.244
R6344 gnd.n1279 gnd.n1278 240.244
R6345 gnd.n1280 gnd.n1279 240.244
R6346 gnd.n5544 gnd.n1280 240.244
R6347 gnd.n5544 gnd.n1283 240.244
R6348 gnd.n1284 gnd.n1283 240.244
R6349 gnd.n1285 gnd.n1284 240.244
R6350 gnd.n1393 gnd.n1285 240.244
R6351 gnd.n1393 gnd.n1288 240.244
R6352 gnd.n1289 gnd.n1288 240.244
R6353 gnd.n1290 gnd.n1289 240.244
R6354 gnd.n1380 gnd.n1290 240.244
R6355 gnd.n1380 gnd.n1293 240.244
R6356 gnd.n1294 gnd.n1293 240.244
R6357 gnd.n1295 gnd.n1294 240.244
R6358 gnd.n1366 gnd.n1295 240.244
R6359 gnd.n1366 gnd.n1298 240.244
R6360 gnd.n1299 gnd.n1298 240.244
R6361 gnd.n1300 gnd.n1299 240.244
R6362 gnd.n1352 gnd.n1300 240.244
R6363 gnd.n1352 gnd.n1303 240.244
R6364 gnd.n1304 gnd.n1303 240.244
R6365 gnd.n1305 gnd.n1304 240.244
R6366 gnd.n1338 gnd.n1305 240.244
R6367 gnd.n1338 gnd.n1308 240.244
R6368 gnd.n1309 gnd.n1308 240.244
R6369 gnd.n1310 gnd.n1309 240.244
R6370 gnd.n1323 gnd.n1310 240.244
R6371 gnd.n1323 gnd.n1313 240.244
R6372 gnd.n6002 gnd.n1313 240.244
R6373 gnd.n5822 gnd.n465 240.244
R6374 gnd.n473 gnd.n472 240.244
R6375 gnd.n5824 gnd.n480 240.244
R6376 gnd.n5827 gnd.n481 240.244
R6377 gnd.n489 gnd.n488 240.244
R6378 gnd.n5829 gnd.n496 240.244
R6379 gnd.n5832 gnd.n497 240.244
R6380 gnd.n507 gnd.n506 240.244
R6381 gnd.n5935 gnd.n5934 240.244
R6382 gnd.n5938 gnd.n5937 240.244
R6383 gnd.n5940 gnd.n5939 240.244
R6384 gnd.n5944 gnd.n5943 240.244
R6385 gnd.n5946 gnd.n5945 240.244
R6386 gnd.n5949 gnd.n1314 240.244
R6387 gnd.n4922 gnd.n4921 240.132
R6388 gnd.n1419 gnd.n1418 240.132
R6389 gnd.n6319 gnd.n6318 225.874
R6390 gnd.n6319 gnd.n973 225.874
R6391 gnd.n6327 gnd.n973 225.874
R6392 gnd.n6328 gnd.n6327 225.874
R6393 gnd.n6329 gnd.n6328 225.874
R6394 gnd.n6329 gnd.n967 225.874
R6395 gnd.n6337 gnd.n967 225.874
R6396 gnd.n6338 gnd.n6337 225.874
R6397 gnd.n6339 gnd.n6338 225.874
R6398 gnd.n6339 gnd.n961 225.874
R6399 gnd.n6347 gnd.n961 225.874
R6400 gnd.n6348 gnd.n6347 225.874
R6401 gnd.n6349 gnd.n6348 225.874
R6402 gnd.n6349 gnd.n955 225.874
R6403 gnd.n6357 gnd.n955 225.874
R6404 gnd.n6358 gnd.n6357 225.874
R6405 gnd.n6359 gnd.n6358 225.874
R6406 gnd.n6359 gnd.n949 225.874
R6407 gnd.n6367 gnd.n949 225.874
R6408 gnd.n6368 gnd.n6367 225.874
R6409 gnd.n6369 gnd.n6368 225.874
R6410 gnd.n6369 gnd.n943 225.874
R6411 gnd.n6377 gnd.n943 225.874
R6412 gnd.n6378 gnd.n6377 225.874
R6413 gnd.n6379 gnd.n6378 225.874
R6414 gnd.n6379 gnd.n937 225.874
R6415 gnd.n6387 gnd.n937 225.874
R6416 gnd.n6388 gnd.n6387 225.874
R6417 gnd.n6389 gnd.n6388 225.874
R6418 gnd.n6389 gnd.n931 225.874
R6419 gnd.n6397 gnd.n931 225.874
R6420 gnd.n6398 gnd.n6397 225.874
R6421 gnd.n6399 gnd.n6398 225.874
R6422 gnd.n6399 gnd.n925 225.874
R6423 gnd.n6407 gnd.n925 225.874
R6424 gnd.n6408 gnd.n6407 225.874
R6425 gnd.n6409 gnd.n6408 225.874
R6426 gnd.n6409 gnd.n919 225.874
R6427 gnd.n6417 gnd.n919 225.874
R6428 gnd.n6418 gnd.n6417 225.874
R6429 gnd.n6419 gnd.n6418 225.874
R6430 gnd.n6419 gnd.n913 225.874
R6431 gnd.n6427 gnd.n913 225.874
R6432 gnd.n6428 gnd.n6427 225.874
R6433 gnd.n6429 gnd.n6428 225.874
R6434 gnd.n6429 gnd.n907 225.874
R6435 gnd.n6437 gnd.n907 225.874
R6436 gnd.n6438 gnd.n6437 225.874
R6437 gnd.n6439 gnd.n6438 225.874
R6438 gnd.n6439 gnd.n901 225.874
R6439 gnd.n6447 gnd.n901 225.874
R6440 gnd.n6448 gnd.n6447 225.874
R6441 gnd.n6449 gnd.n6448 225.874
R6442 gnd.n6449 gnd.n895 225.874
R6443 gnd.n6457 gnd.n895 225.874
R6444 gnd.n6458 gnd.n6457 225.874
R6445 gnd.n6459 gnd.n6458 225.874
R6446 gnd.n6459 gnd.n889 225.874
R6447 gnd.n6467 gnd.n889 225.874
R6448 gnd.n6468 gnd.n6467 225.874
R6449 gnd.n6469 gnd.n6468 225.874
R6450 gnd.n6469 gnd.n883 225.874
R6451 gnd.n6477 gnd.n883 225.874
R6452 gnd.n6478 gnd.n6477 225.874
R6453 gnd.n6479 gnd.n6478 225.874
R6454 gnd.n6479 gnd.n877 225.874
R6455 gnd.n6487 gnd.n877 225.874
R6456 gnd.n6488 gnd.n6487 225.874
R6457 gnd.n6489 gnd.n6488 225.874
R6458 gnd.n6489 gnd.n871 225.874
R6459 gnd.n6497 gnd.n871 225.874
R6460 gnd.n6498 gnd.n6497 225.874
R6461 gnd.n6499 gnd.n6498 225.874
R6462 gnd.n6499 gnd.n865 225.874
R6463 gnd.n6507 gnd.n865 225.874
R6464 gnd.n6508 gnd.n6507 225.874
R6465 gnd.n6509 gnd.n6508 225.874
R6466 gnd.n6509 gnd.n859 225.874
R6467 gnd.n6517 gnd.n859 225.874
R6468 gnd.n6518 gnd.n6517 225.874
R6469 gnd.n6519 gnd.n6518 225.874
R6470 gnd.n6519 gnd.n853 225.874
R6471 gnd.n6527 gnd.n853 225.874
R6472 gnd.n6528 gnd.n6527 225.874
R6473 gnd.n6529 gnd.n6528 225.874
R6474 gnd.n6529 gnd.n847 225.874
R6475 gnd.n6537 gnd.n847 225.874
R6476 gnd.n6538 gnd.n6537 225.874
R6477 gnd.n6539 gnd.n6538 225.874
R6478 gnd.n6539 gnd.n841 225.874
R6479 gnd.n6547 gnd.n841 225.874
R6480 gnd.n6548 gnd.n6547 225.874
R6481 gnd.n6549 gnd.n6548 225.874
R6482 gnd.n6549 gnd.n835 225.874
R6483 gnd.n6557 gnd.n835 225.874
R6484 gnd.n6558 gnd.n6557 225.874
R6485 gnd.n6559 gnd.n6558 225.874
R6486 gnd.n6559 gnd.n829 225.874
R6487 gnd.n6567 gnd.n829 225.874
R6488 gnd.n6568 gnd.n6567 225.874
R6489 gnd.n6569 gnd.n6568 225.874
R6490 gnd.n6569 gnd.n823 225.874
R6491 gnd.n6577 gnd.n823 225.874
R6492 gnd.n6578 gnd.n6577 225.874
R6493 gnd.n6579 gnd.n6578 225.874
R6494 gnd.n6579 gnd.n817 225.874
R6495 gnd.n6587 gnd.n817 225.874
R6496 gnd.n6588 gnd.n6587 225.874
R6497 gnd.n6589 gnd.n6588 225.874
R6498 gnd.n6589 gnd.n811 225.874
R6499 gnd.n6597 gnd.n811 225.874
R6500 gnd.n6598 gnd.n6597 225.874
R6501 gnd.n6599 gnd.n6598 225.874
R6502 gnd.n6599 gnd.n805 225.874
R6503 gnd.n6607 gnd.n805 225.874
R6504 gnd.n6608 gnd.n6607 225.874
R6505 gnd.n6609 gnd.n6608 225.874
R6506 gnd.n6609 gnd.n799 225.874
R6507 gnd.n6617 gnd.n799 225.874
R6508 gnd.n6618 gnd.n6617 225.874
R6509 gnd.n6619 gnd.n6618 225.874
R6510 gnd.n6619 gnd.n793 225.874
R6511 gnd.n6627 gnd.n793 225.874
R6512 gnd.n6628 gnd.n6627 225.874
R6513 gnd.n6629 gnd.n6628 225.874
R6514 gnd.n6629 gnd.n787 225.874
R6515 gnd.n6637 gnd.n787 225.874
R6516 gnd.n6638 gnd.n6637 225.874
R6517 gnd.n6639 gnd.n6638 225.874
R6518 gnd.n6639 gnd.n781 225.874
R6519 gnd.n6647 gnd.n781 225.874
R6520 gnd.n6648 gnd.n6647 225.874
R6521 gnd.n6649 gnd.n6648 225.874
R6522 gnd.n6649 gnd.n775 225.874
R6523 gnd.n6657 gnd.n775 225.874
R6524 gnd.n6658 gnd.n6657 225.874
R6525 gnd.n6659 gnd.n6658 225.874
R6526 gnd.n6659 gnd.n769 225.874
R6527 gnd.n6667 gnd.n769 225.874
R6528 gnd.n6668 gnd.n6667 225.874
R6529 gnd.n6669 gnd.n6668 225.874
R6530 gnd.n6669 gnd.n763 225.874
R6531 gnd.n6677 gnd.n763 225.874
R6532 gnd.n6678 gnd.n6677 225.874
R6533 gnd.n6679 gnd.n6678 225.874
R6534 gnd.n6679 gnd.n757 225.874
R6535 gnd.n6687 gnd.n757 225.874
R6536 gnd.n6688 gnd.n6687 225.874
R6537 gnd.n6689 gnd.n6688 225.874
R6538 gnd.n6689 gnd.n751 225.874
R6539 gnd.n6698 gnd.n751 225.874
R6540 gnd.n6699 gnd.n6698 225.874
R6541 gnd.n6700 gnd.n6699 225.874
R6542 gnd.n6700 gnd.n746 225.874
R6543 gnd.n2724 gnd.t302 224.174
R6544 gnd.n2222 gnd.t279 224.174
R6545 gnd.n562 gnd.n518 199.319
R6546 gnd.n562 gnd.n519 199.319
R6547 gnd.n6223 gnd.n6222 199.319
R6548 gnd.n6222 gnd.n6221 199.319
R6549 gnd.n4923 gnd.n4920 186.49
R6550 gnd.n1420 gnd.n1417 186.49
R6551 gnd.n3499 gnd.n3498 185
R6552 gnd.n3497 gnd.n3496 185
R6553 gnd.n3476 gnd.n3475 185
R6554 gnd.n3491 gnd.n3490 185
R6555 gnd.n3489 gnd.n3488 185
R6556 gnd.n3480 gnd.n3479 185
R6557 gnd.n3483 gnd.n3482 185
R6558 gnd.n3467 gnd.n3466 185
R6559 gnd.n3465 gnd.n3464 185
R6560 gnd.n3444 gnd.n3443 185
R6561 gnd.n3459 gnd.n3458 185
R6562 gnd.n3457 gnd.n3456 185
R6563 gnd.n3448 gnd.n3447 185
R6564 gnd.n3451 gnd.n3450 185
R6565 gnd.n3435 gnd.n3434 185
R6566 gnd.n3433 gnd.n3432 185
R6567 gnd.n3412 gnd.n3411 185
R6568 gnd.n3427 gnd.n3426 185
R6569 gnd.n3425 gnd.n3424 185
R6570 gnd.n3416 gnd.n3415 185
R6571 gnd.n3419 gnd.n3418 185
R6572 gnd.n3404 gnd.n3403 185
R6573 gnd.n3402 gnd.n3401 185
R6574 gnd.n3381 gnd.n3380 185
R6575 gnd.n3396 gnd.n3395 185
R6576 gnd.n3394 gnd.n3393 185
R6577 gnd.n3385 gnd.n3384 185
R6578 gnd.n3388 gnd.n3387 185
R6579 gnd.n3372 gnd.n3371 185
R6580 gnd.n3370 gnd.n3369 185
R6581 gnd.n3349 gnd.n3348 185
R6582 gnd.n3364 gnd.n3363 185
R6583 gnd.n3362 gnd.n3361 185
R6584 gnd.n3353 gnd.n3352 185
R6585 gnd.n3356 gnd.n3355 185
R6586 gnd.n3340 gnd.n3339 185
R6587 gnd.n3338 gnd.n3337 185
R6588 gnd.n3317 gnd.n3316 185
R6589 gnd.n3332 gnd.n3331 185
R6590 gnd.n3330 gnd.n3329 185
R6591 gnd.n3321 gnd.n3320 185
R6592 gnd.n3324 gnd.n3323 185
R6593 gnd.n3308 gnd.n3307 185
R6594 gnd.n3306 gnd.n3305 185
R6595 gnd.n3285 gnd.n3284 185
R6596 gnd.n3300 gnd.n3299 185
R6597 gnd.n3298 gnd.n3297 185
R6598 gnd.n3289 gnd.n3288 185
R6599 gnd.n3292 gnd.n3291 185
R6600 gnd.n3277 gnd.n3276 185
R6601 gnd.n3275 gnd.n3274 185
R6602 gnd.n3254 gnd.n3253 185
R6603 gnd.n3269 gnd.n3268 185
R6604 gnd.n3267 gnd.n3266 185
R6605 gnd.n3258 gnd.n3257 185
R6606 gnd.n3261 gnd.n3260 185
R6607 gnd.n2725 gnd.t301 178.987
R6608 gnd.n2223 gnd.t280 178.987
R6609 gnd.n1 gnd.t134 170.774
R6610 gnd.n9 gnd.t117 170.103
R6611 gnd.n8 gnd.t354 170.103
R6612 gnd.n7 gnd.t124 170.103
R6613 gnd.n6 gnd.t50 170.103
R6614 gnd.n5 gnd.t136 170.103
R6615 gnd.n4 gnd.t348 170.103
R6616 gnd.n3 gnd.t225 170.103
R6617 gnd.n2 gnd.t93 170.103
R6618 gnd.n1 gnd.t358 170.103
R6619 gnd.n7147 gnd.n561 164.544
R6620 gnd.n5013 gnd.n1122 164.544
R6621 gnd.n5706 gnd.n5705 163.367
R6622 gnd.n5703 gnd.n1429 163.367
R6623 gnd.n5699 gnd.n5698 163.367
R6624 gnd.n5696 gnd.n1432 163.367
R6625 gnd.n5692 gnd.n5691 163.367
R6626 gnd.n5689 gnd.n1435 163.367
R6627 gnd.n5685 gnd.n5684 163.367
R6628 gnd.n5682 gnd.n1438 163.367
R6629 gnd.n5678 gnd.n5677 163.367
R6630 gnd.n5675 gnd.n1441 163.367
R6631 gnd.n5671 gnd.n5670 163.367
R6632 gnd.n5668 gnd.n1444 163.367
R6633 gnd.n5664 gnd.n5663 163.367
R6634 gnd.n5661 gnd.n1447 163.367
R6635 gnd.n5656 gnd.n5655 163.367
R6636 gnd.n5653 gnd.n5651 163.367
R6637 gnd.n5648 gnd.n5647 163.367
R6638 gnd.n5645 gnd.n1453 163.367
R6639 gnd.n5640 gnd.n5639 163.367
R6640 gnd.n5637 gnd.n1458 163.367
R6641 gnd.n5633 gnd.n5632 163.367
R6642 gnd.n5630 gnd.n1461 163.367
R6643 gnd.n5626 gnd.n5625 163.367
R6644 gnd.n5623 gnd.n1464 163.367
R6645 gnd.n5619 gnd.n5618 163.367
R6646 gnd.n5616 gnd.n1467 163.367
R6647 gnd.n5612 gnd.n5611 163.367
R6648 gnd.n5609 gnd.n1470 163.367
R6649 gnd.n5605 gnd.n5604 163.367
R6650 gnd.n5602 gnd.n1473 163.367
R6651 gnd.n5598 gnd.n5597 163.367
R6652 gnd.n5595 gnd.n1476 163.367
R6653 gnd.n4945 gnd.n1821 163.367
R6654 gnd.n1821 gnd.n1768 163.367
R6655 gnd.n5103 gnd.n1768 163.367
R6656 gnd.n5103 gnd.n1763 163.367
R6657 gnd.n5099 gnd.n1763 163.367
R6658 gnd.n5099 gnd.n1752 163.367
R6659 gnd.n1812 gnd.n1752 163.367
R6660 gnd.n1812 gnd.n1746 163.367
R6661 gnd.n1809 gnd.n1746 163.367
R6662 gnd.n1809 gnd.n1739 163.367
R6663 gnd.n1804 gnd.n1739 163.367
R6664 gnd.n1804 gnd.n1733 163.367
R6665 gnd.n1800 gnd.n1733 163.367
R6666 gnd.n1800 gnd.n1727 163.367
R6667 gnd.n1794 gnd.n1727 163.367
R6668 gnd.n1794 gnd.n1720 163.367
R6669 gnd.n1791 gnd.n1720 163.367
R6670 gnd.n1791 gnd.n1789 163.367
R6671 gnd.n1789 gnd.n1704 163.367
R6672 gnd.n1705 gnd.n1704 163.367
R6673 gnd.n1705 gnd.n1697 163.367
R6674 gnd.n1783 gnd.n1697 163.367
R6675 gnd.n1783 gnd.n1689 163.367
R6676 gnd.n1779 gnd.n1689 163.367
R6677 gnd.n1779 gnd.n1683 163.367
R6678 gnd.n1776 gnd.n1683 163.367
R6679 gnd.n1776 gnd.n1675 163.367
R6680 gnd.n1771 gnd.n1675 163.367
R6681 gnd.n1771 gnd.n1666 163.367
R6682 gnd.n1666 gnd.n1656 163.367
R6683 gnd.n5252 gnd.n1656 163.367
R6684 gnd.n5252 gnd.n1650 163.367
R6685 gnd.n5256 gnd.n1650 163.367
R6686 gnd.n5256 gnd.n1643 163.367
R6687 gnd.n5276 gnd.n1643 163.367
R6688 gnd.n5276 gnd.n1640 163.367
R6689 gnd.n5290 gnd.n1640 163.367
R6690 gnd.n5290 gnd.n1634 163.367
R6691 gnd.n5286 gnd.n1634 163.367
R6692 gnd.n5286 gnd.n5282 163.367
R6693 gnd.n5282 gnd.n5281 163.367
R6694 gnd.n5281 gnd.n1616 163.367
R6695 gnd.n5335 gnd.n1616 163.367
R6696 gnd.n5335 gnd.n1614 163.367
R6697 gnd.n5355 gnd.n1614 163.367
R6698 gnd.n5355 gnd.n1607 163.367
R6699 gnd.n5351 gnd.n1607 163.367
R6700 gnd.n5351 gnd.n5348 163.367
R6701 gnd.n5348 gnd.n5347 163.367
R6702 gnd.n5347 gnd.n1589 163.367
R6703 gnd.n1590 gnd.n1589 163.367
R6704 gnd.n1590 gnd.n1582 163.367
R6705 gnd.n5341 gnd.n1582 163.367
R6706 gnd.n5341 gnd.n1574 163.367
R6707 gnd.n5412 gnd.n1574 163.367
R6708 gnd.n5412 gnd.n1567 163.367
R6709 gnd.n5415 gnd.n1567 163.367
R6710 gnd.n5415 gnd.n1560 163.367
R6711 gnd.n5419 gnd.n1560 163.367
R6712 gnd.n5419 gnd.n1552 163.367
R6713 gnd.n5453 gnd.n1552 163.367
R6714 gnd.n5453 gnd.n1545 163.367
R6715 gnd.n5456 gnd.n1545 163.367
R6716 gnd.n5456 gnd.n1539 163.367
R6717 gnd.n5469 gnd.n1539 163.367
R6718 gnd.n5469 gnd.n1530 163.367
R6719 gnd.n5465 gnd.n1530 163.367
R6720 gnd.n5465 gnd.n1526 163.367
R6721 gnd.n5462 gnd.n1526 163.367
R6722 gnd.n5462 gnd.n1512 163.367
R6723 gnd.n5459 gnd.n1512 163.367
R6724 gnd.n5459 gnd.n1505 163.367
R6725 gnd.n5533 gnd.n1505 163.367
R6726 gnd.n5533 gnd.n1495 163.367
R6727 gnd.n5536 gnd.n1495 163.367
R6728 gnd.n5536 gnd.n1489 163.367
R6729 gnd.n5542 gnd.n1489 163.367
R6730 gnd.n5542 gnd.n1483 163.367
R6731 gnd.n1483 gnd.n1478 163.367
R6732 gnd.n5584 gnd.n1478 163.367
R6733 gnd.n5585 gnd.n5584 163.367
R6734 gnd.n5585 gnd.n1403 163.367
R6735 gnd.n5590 gnd.n1403 163.367
R6736 gnd.n4914 gnd.n4913 163.367
R6737 gnd.n5070 gnd.n4913 163.367
R6738 gnd.n5068 gnd.n5067 163.367
R6739 gnd.n5064 gnd.n5063 163.367
R6740 gnd.n5060 gnd.n5059 163.367
R6741 gnd.n5056 gnd.n5055 163.367
R6742 gnd.n5052 gnd.n5051 163.367
R6743 gnd.n5048 gnd.n5047 163.367
R6744 gnd.n5044 gnd.n5043 163.367
R6745 gnd.n5040 gnd.n5039 163.367
R6746 gnd.n5036 gnd.n5035 163.367
R6747 gnd.n5032 gnd.n5031 163.367
R6748 gnd.n5028 gnd.n5027 163.367
R6749 gnd.n5024 gnd.n5023 163.367
R6750 gnd.n5020 gnd.n5019 163.367
R6751 gnd.n5016 gnd.n5015 163.367
R6752 gnd.n5012 gnd.n5011 163.367
R6753 gnd.n5007 gnd.n5006 163.367
R6754 gnd.n5002 gnd.n5001 163.367
R6755 gnd.n4998 gnd.n4997 163.367
R6756 gnd.n4994 gnd.n4993 163.367
R6757 gnd.n4990 gnd.n4989 163.367
R6758 gnd.n4986 gnd.n4985 163.367
R6759 gnd.n4982 gnd.n4981 163.367
R6760 gnd.n4978 gnd.n4977 163.367
R6761 gnd.n4974 gnd.n4973 163.367
R6762 gnd.n4970 gnd.n4969 163.367
R6763 gnd.n4966 gnd.n4965 163.367
R6764 gnd.n4962 gnd.n4961 163.367
R6765 gnd.n4958 gnd.n4957 163.367
R6766 gnd.n4954 gnd.n4953 163.367
R6767 gnd.n4950 gnd.n4949 163.367
R6768 gnd.n4915 gnd.n1766 163.367
R6769 gnd.n5107 gnd.n1766 163.367
R6770 gnd.n5107 gnd.n1764 163.367
R6771 gnd.n5111 gnd.n1764 163.367
R6772 gnd.n5111 gnd.n1750 163.367
R6773 gnd.n5124 gnd.n1750 163.367
R6774 gnd.n5124 gnd.n1748 163.367
R6775 gnd.n5128 gnd.n1748 163.367
R6776 gnd.n5128 gnd.n1737 163.367
R6777 gnd.n5142 gnd.n1737 163.367
R6778 gnd.n5142 gnd.n1735 163.367
R6779 gnd.n5146 gnd.n1735 163.367
R6780 gnd.n5146 gnd.n1725 163.367
R6781 gnd.n5158 gnd.n1725 163.367
R6782 gnd.n5158 gnd.n1722 163.367
R6783 gnd.n5163 gnd.n1722 163.367
R6784 gnd.n5163 gnd.n1723 163.367
R6785 gnd.n1723 gnd.n1701 163.367
R6786 gnd.n5188 gnd.n1701 163.367
R6787 gnd.n5188 gnd.n1699 163.367
R6788 gnd.n5192 gnd.n1699 163.367
R6789 gnd.n5192 gnd.n1687 163.367
R6790 gnd.n5207 gnd.n1687 163.367
R6791 gnd.n5207 gnd.n1685 163.367
R6792 gnd.n5211 gnd.n1685 163.367
R6793 gnd.n5211 gnd.n1673 163.367
R6794 gnd.n5224 gnd.n1673 163.367
R6795 gnd.n5224 gnd.n1668 163.367
R6796 gnd.n5229 gnd.n1668 163.367
R6797 gnd.n5229 gnd.n1671 163.367
R6798 gnd.n1671 gnd.n1651 163.367
R6799 gnd.n5264 gnd.n1651 163.367
R6800 gnd.n5264 gnd.n1652 163.367
R6801 gnd.n5260 gnd.n1652 163.367
R6802 gnd.n5260 gnd.n1638 163.367
R6803 gnd.n5294 gnd.n1638 163.367
R6804 gnd.n5294 gnd.n1635 163.367
R6805 gnd.n5307 gnd.n1635 163.367
R6806 gnd.n5307 gnd.n1636 163.367
R6807 gnd.n5303 gnd.n1636 163.367
R6808 gnd.n5303 gnd.n5302 163.367
R6809 gnd.n5302 gnd.n5301 163.367
R6810 gnd.n5301 gnd.n1612 163.367
R6811 gnd.n5359 gnd.n1612 163.367
R6812 gnd.n5359 gnd.n1609 163.367
R6813 gnd.n5366 gnd.n1609 163.367
R6814 gnd.n5366 gnd.n1610 163.367
R6815 gnd.n5362 gnd.n1610 163.367
R6816 gnd.n5362 gnd.n1587 163.367
R6817 gnd.n5393 gnd.n1587 163.367
R6818 gnd.n5393 gnd.n1584 163.367
R6819 gnd.n5400 gnd.n1584 163.367
R6820 gnd.n5400 gnd.n1585 163.367
R6821 gnd.n5396 gnd.n1585 163.367
R6822 gnd.n5396 gnd.n1565 163.367
R6823 gnd.n5434 gnd.n1565 163.367
R6824 gnd.n5434 gnd.n1562 163.367
R6825 gnd.n5441 gnd.n1562 163.367
R6826 gnd.n5441 gnd.n1563 163.367
R6827 gnd.n5437 gnd.n1563 163.367
R6828 gnd.n5437 gnd.n1543 163.367
R6829 gnd.n5484 gnd.n1543 163.367
R6830 gnd.n5484 gnd.n1541 163.367
R6831 gnd.n5488 gnd.n1541 163.367
R6832 gnd.n5488 gnd.n1529 163.367
R6833 gnd.n5500 gnd.n1529 163.367
R6834 gnd.n5500 gnd.n1527 163.367
R6835 gnd.n5504 gnd.n1527 163.367
R6836 gnd.n5504 gnd.n1514 163.367
R6837 gnd.n5520 gnd.n1514 163.367
R6838 gnd.n5520 gnd.n1515 163.367
R6839 gnd.n5516 gnd.n1515 163.367
R6840 gnd.n5516 gnd.n1493 163.367
R6841 gnd.n5562 gnd.n1493 163.367
R6842 gnd.n5562 gnd.n1491 163.367
R6843 gnd.n5566 gnd.n1491 163.367
R6844 gnd.n5566 gnd.n1482 163.367
R6845 gnd.n5578 gnd.n1482 163.367
R6846 gnd.n5578 gnd.n1480 163.367
R6847 gnd.n5582 gnd.n1480 163.367
R6848 gnd.n5582 gnd.n1405 163.367
R6849 gnd.n5713 gnd.n1405 163.367
R6850 gnd.n5713 gnd.n1406 163.367
R6851 gnd.n1426 gnd.n1425 156.462
R6852 gnd.n3439 gnd.n3407 153.042
R6853 gnd.n3503 gnd.n3502 152.079
R6854 gnd.n3471 gnd.n3470 152.079
R6855 gnd.n3439 gnd.n3438 152.079
R6856 gnd.n4928 gnd.n4927 152
R6857 gnd.n4929 gnd.n4918 152
R6858 gnd.n4931 gnd.n4930 152
R6859 gnd.n4933 gnd.n4916 152
R6860 gnd.n4935 gnd.n4934 152
R6861 gnd.n1424 gnd.n1408 152
R6862 gnd.n1416 gnd.n1409 152
R6863 gnd.n1415 gnd.n1414 152
R6864 gnd.n1413 gnd.n1410 152
R6865 gnd.n1411 gnd.t274 150.546
R6866 gnd.t38 gnd.n3481 147.661
R6867 gnd.t165 gnd.n3449 147.661
R6868 gnd.t336 gnd.n3417 147.661
R6869 gnd.t9 gnd.n3386 147.661
R6870 gnd.t91 gnd.n3354 147.661
R6871 gnd.t115 gnd.n3322 147.661
R6872 gnd.t161 gnd.n3290 147.661
R6873 gnd.t181 gnd.n3259 147.661
R6874 gnd.n5650 gnd.n5649 143.351
R6875 gnd.n5010 gnd.n4893 143.351
R6876 gnd.n5010 gnd.n4894 143.351
R6877 gnd.n4925 gnd.t231 130.484
R6878 gnd.n4934 gnd.t234 126.766
R6879 gnd.n4932 gnd.t306 126.766
R6880 gnd.n4918 gnd.t332 126.766
R6881 gnd.n4926 gnd.t281 126.766
R6882 gnd.n1412 gnd.t253 126.766
R6883 gnd.n1414 gnd.t287 126.766
R6884 gnd.n1423 gnd.t264 126.766
R6885 gnd.n1425 gnd.t290 126.766
R6886 gnd.n3498 gnd.n3497 104.615
R6887 gnd.n3497 gnd.n3475 104.615
R6888 gnd.n3490 gnd.n3475 104.615
R6889 gnd.n3490 gnd.n3489 104.615
R6890 gnd.n3489 gnd.n3479 104.615
R6891 gnd.n3482 gnd.n3479 104.615
R6892 gnd.n3466 gnd.n3465 104.615
R6893 gnd.n3465 gnd.n3443 104.615
R6894 gnd.n3458 gnd.n3443 104.615
R6895 gnd.n3458 gnd.n3457 104.615
R6896 gnd.n3457 gnd.n3447 104.615
R6897 gnd.n3450 gnd.n3447 104.615
R6898 gnd.n3434 gnd.n3433 104.615
R6899 gnd.n3433 gnd.n3411 104.615
R6900 gnd.n3426 gnd.n3411 104.615
R6901 gnd.n3426 gnd.n3425 104.615
R6902 gnd.n3425 gnd.n3415 104.615
R6903 gnd.n3418 gnd.n3415 104.615
R6904 gnd.n3403 gnd.n3402 104.615
R6905 gnd.n3402 gnd.n3380 104.615
R6906 gnd.n3395 gnd.n3380 104.615
R6907 gnd.n3395 gnd.n3394 104.615
R6908 gnd.n3394 gnd.n3384 104.615
R6909 gnd.n3387 gnd.n3384 104.615
R6910 gnd.n3371 gnd.n3370 104.615
R6911 gnd.n3370 gnd.n3348 104.615
R6912 gnd.n3363 gnd.n3348 104.615
R6913 gnd.n3363 gnd.n3362 104.615
R6914 gnd.n3362 gnd.n3352 104.615
R6915 gnd.n3355 gnd.n3352 104.615
R6916 gnd.n3339 gnd.n3338 104.615
R6917 gnd.n3338 gnd.n3316 104.615
R6918 gnd.n3331 gnd.n3316 104.615
R6919 gnd.n3331 gnd.n3330 104.615
R6920 gnd.n3330 gnd.n3320 104.615
R6921 gnd.n3323 gnd.n3320 104.615
R6922 gnd.n3307 gnd.n3306 104.615
R6923 gnd.n3306 gnd.n3284 104.615
R6924 gnd.n3299 gnd.n3284 104.615
R6925 gnd.n3299 gnd.n3298 104.615
R6926 gnd.n3298 gnd.n3288 104.615
R6927 gnd.n3291 gnd.n3288 104.615
R6928 gnd.n3276 gnd.n3275 104.615
R6929 gnd.n3275 gnd.n3253 104.615
R6930 gnd.n3268 gnd.n3253 104.615
R6931 gnd.n3268 gnd.n3267 104.615
R6932 gnd.n3267 gnd.n3257 104.615
R6933 gnd.n3260 gnd.n3257 104.615
R6934 gnd.n2650 gnd.t319 100.632
R6935 gnd.n2196 gnd.t262 100.632
R6936 gnd.n7621 gnd.n138 99.6594
R6937 gnd.n7619 gnd.n7618 99.6594
R6938 gnd.n7614 gnd.n145 99.6594
R6939 gnd.n7612 gnd.n7611 99.6594
R6940 gnd.n7607 gnd.n152 99.6594
R6941 gnd.n7605 gnd.n7604 99.6594
R6942 gnd.n7600 gnd.n159 99.6594
R6943 gnd.n7598 gnd.n7597 99.6594
R6944 gnd.n7590 gnd.n166 99.6594
R6945 gnd.n7588 gnd.n7587 99.6594
R6946 gnd.n7583 gnd.n173 99.6594
R6947 gnd.n7581 gnd.n7580 99.6594
R6948 gnd.n7576 gnd.n180 99.6594
R6949 gnd.n7574 gnd.n7573 99.6594
R6950 gnd.n7569 gnd.n187 99.6594
R6951 gnd.n7567 gnd.n7566 99.6594
R6952 gnd.n7562 gnd.n194 99.6594
R6953 gnd.n7560 gnd.n7559 99.6594
R6954 gnd.n199 gnd.n198 99.6594
R6955 gnd.n7177 gnd.n454 99.6594
R6956 gnd.n7172 gnd.n512 99.6594
R6957 gnd.n7169 gnd.n513 99.6594
R6958 gnd.n7165 gnd.n514 99.6594
R6959 gnd.n7161 gnd.n515 99.6594
R6960 gnd.n7157 gnd.n516 99.6594
R6961 gnd.n7153 gnd.n517 99.6594
R6962 gnd.n7149 gnd.n518 99.6594
R6963 gnd.n7144 gnd.n520 99.6594
R6964 gnd.n7140 gnd.n521 99.6594
R6965 gnd.n7136 gnd.n522 99.6594
R6966 gnd.n7132 gnd.n523 99.6594
R6967 gnd.n7128 gnd.n524 99.6594
R6968 gnd.n7124 gnd.n525 99.6594
R6969 gnd.n7120 gnd.n526 99.6594
R6970 gnd.n7116 gnd.n527 99.6594
R6971 gnd.n7112 gnd.n528 99.6594
R6972 gnd.n585 gnd.n529 99.6594
R6973 gnd.n7476 gnd.n7475 99.6594
R6974 gnd.n7481 gnd.n7480 99.6594
R6975 gnd.n7484 gnd.n7483 99.6594
R6976 gnd.n7489 gnd.n7488 99.6594
R6977 gnd.n7492 gnd.n7491 99.6594
R6978 gnd.n7497 gnd.n7496 99.6594
R6979 gnd.n7500 gnd.n7499 99.6594
R6980 gnd.n7505 gnd.n7503 99.6594
R6981 gnd.n7631 gnd.n125 99.6594
R6982 gnd.n530 gnd.n459 99.6594
R6983 gnd.n532 gnd.n531 99.6594
R6984 gnd.n534 gnd.n469 99.6594
R6985 gnd.n535 gnd.n476 99.6594
R6986 gnd.n537 gnd.n536 99.6594
R6987 gnd.n539 gnd.n485 99.6594
R6988 gnd.n540 gnd.n492 99.6594
R6989 gnd.n542 gnd.n541 99.6594
R6990 gnd.n543 gnd.n501 99.6594
R6991 gnd.n4532 gnd.n4531 99.6594
R6992 gnd.n4526 gnd.n1948 99.6594
R6993 gnd.n4523 gnd.n1949 99.6594
R6994 gnd.n4519 gnd.n1950 99.6594
R6995 gnd.n4515 gnd.n1951 99.6594
R6996 gnd.n4511 gnd.n1952 99.6594
R6997 gnd.n4507 gnd.n1953 99.6594
R6998 gnd.n4503 gnd.n1954 99.6594
R6999 gnd.n4499 gnd.n1955 99.6594
R7000 gnd.n4495 gnd.n1956 99.6594
R7001 gnd.n4491 gnd.n1957 99.6594
R7002 gnd.n4487 gnd.n1958 99.6594
R7003 gnd.n4483 gnd.n1959 99.6594
R7004 gnd.n4479 gnd.n1960 99.6594
R7005 gnd.n4475 gnd.n1961 99.6594
R7006 gnd.n4471 gnd.n1962 99.6594
R7007 gnd.n4467 gnd.n1963 99.6594
R7008 gnd.n4463 gnd.n1964 99.6594
R7009 gnd.n4459 gnd.n1965 99.6594
R7010 gnd.n4455 gnd.n1966 99.6594
R7011 gnd.n4451 gnd.n1967 99.6594
R7012 gnd.n4447 gnd.n1968 99.6594
R7013 gnd.n4443 gnd.n1969 99.6594
R7014 gnd.n4439 gnd.n1970 99.6594
R7015 gnd.n4435 gnd.n1971 99.6594
R7016 gnd.n4431 gnd.n1972 99.6594
R7017 gnd.n4427 gnd.n1973 99.6594
R7018 gnd.n4423 gnd.n1974 99.6594
R7019 gnd.n4419 gnd.n1975 99.6594
R7020 gnd.n4415 gnd.n1976 99.6594
R7021 gnd.n4411 gnd.n1977 99.6594
R7022 gnd.n4407 gnd.n1978 99.6594
R7023 gnd.n4403 gnd.n1979 99.6594
R7024 gnd.n4399 gnd.n1980 99.6594
R7025 gnd.n4395 gnd.n1981 99.6594
R7026 gnd.n4391 gnd.n1982 99.6594
R7027 gnd.n4387 gnd.n1983 99.6594
R7028 gnd.n4383 gnd.n1984 99.6594
R7029 gnd.n4379 gnd.n1985 99.6594
R7030 gnd.n4375 gnd.n1986 99.6594
R7031 gnd.n4371 gnd.n1987 99.6594
R7032 gnd.n4534 gnd.n1947 99.6594
R7033 gnd.n6247 gnd.n6246 99.6594
R7034 gnd.n6244 gnd.n6243 99.6594
R7035 gnd.n6239 gnd.n1105 99.6594
R7036 gnd.n6237 gnd.n6236 99.6594
R7037 gnd.n6232 gnd.n1112 99.6594
R7038 gnd.n6230 gnd.n6229 99.6594
R7039 gnd.n6225 gnd.n1119 99.6594
R7040 gnd.n6221 gnd.n6220 99.6594
R7041 gnd.n6216 gnd.n1130 99.6594
R7042 gnd.n6214 gnd.n6213 99.6594
R7043 gnd.n6209 gnd.n1137 99.6594
R7044 gnd.n6207 gnd.n6206 99.6594
R7045 gnd.n6202 gnd.n1144 99.6594
R7046 gnd.n6200 gnd.n6199 99.6594
R7047 gnd.n6195 gnd.n1151 99.6594
R7048 gnd.n6193 gnd.n6192 99.6594
R7049 gnd.n6188 gnd.n1160 99.6594
R7050 gnd.n6186 gnd.n6185 99.6594
R7051 gnd.n3774 gnd.n2156 99.6594
R7052 gnd.n3782 gnd.n3781 99.6594
R7053 gnd.n3785 gnd.n3784 99.6594
R7054 gnd.n3792 gnd.n3791 99.6594
R7055 gnd.n3795 gnd.n3794 99.6594
R7056 gnd.n3802 gnd.n3801 99.6594
R7057 gnd.n3805 gnd.n3804 99.6594
R7058 gnd.n3812 gnd.n3811 99.6594
R7059 gnd.n3815 gnd.n3814 99.6594
R7060 gnd.n3822 gnd.n3821 99.6594
R7061 gnd.n3825 gnd.n3824 99.6594
R7062 gnd.n3832 gnd.n3831 99.6594
R7063 gnd.n3835 gnd.n3834 99.6594
R7064 gnd.n3842 gnd.n3841 99.6594
R7065 gnd.n3845 gnd.n3844 99.6594
R7066 gnd.n3852 gnd.n3851 99.6594
R7067 gnd.n3855 gnd.n3854 99.6594
R7068 gnd.n3863 gnd.n3862 99.6594
R7069 gnd.n3866 gnd.n3865 99.6594
R7070 gnd.n3621 gnd.n2179 99.6594
R7071 gnd.n3619 gnd.n2178 99.6594
R7072 gnd.n3615 gnd.n2177 99.6594
R7073 gnd.n3611 gnd.n2176 99.6594
R7074 gnd.n3607 gnd.n2175 99.6594
R7075 gnd.n3603 gnd.n2174 99.6594
R7076 gnd.n3599 gnd.n2173 99.6594
R7077 gnd.n3531 gnd.n2172 99.6594
R7078 gnd.n2862 gnd.n2593 99.6594
R7079 gnd.n2619 gnd.n2600 99.6594
R7080 gnd.n2621 gnd.n2601 99.6594
R7081 gnd.n2629 gnd.n2602 99.6594
R7082 gnd.n2631 gnd.n2603 99.6594
R7083 gnd.n2639 gnd.n2604 99.6594
R7084 gnd.n2641 gnd.n2605 99.6594
R7085 gnd.n2649 gnd.n2606 99.6594
R7086 gnd.n3589 gnd.n2159 99.6594
R7087 gnd.n3585 gnd.n2160 99.6594
R7088 gnd.n3581 gnd.n2161 99.6594
R7089 gnd.n3577 gnd.n2162 99.6594
R7090 gnd.n3573 gnd.n2163 99.6594
R7091 gnd.n3569 gnd.n2164 99.6594
R7092 gnd.n3565 gnd.n2165 99.6594
R7093 gnd.n3561 gnd.n2166 99.6594
R7094 gnd.n3557 gnd.n2167 99.6594
R7095 gnd.n3553 gnd.n2168 99.6594
R7096 gnd.n3549 gnd.n2169 99.6594
R7097 gnd.n3545 gnd.n2170 99.6594
R7098 gnd.n3541 gnd.n2171 99.6594
R7099 gnd.n2777 gnd.n2776 99.6594
R7100 gnd.n2771 gnd.n2688 99.6594
R7101 gnd.n2768 gnd.n2689 99.6594
R7102 gnd.n2764 gnd.n2690 99.6594
R7103 gnd.n2760 gnd.n2691 99.6594
R7104 gnd.n2756 gnd.n2692 99.6594
R7105 gnd.n2752 gnd.n2693 99.6594
R7106 gnd.n2748 gnd.n2694 99.6594
R7107 gnd.n2744 gnd.n2695 99.6594
R7108 gnd.n2740 gnd.n2696 99.6594
R7109 gnd.n2736 gnd.n2697 99.6594
R7110 gnd.n2732 gnd.n2698 99.6594
R7111 gnd.n2779 gnd.n2687 99.6594
R7112 gnd.n4664 gnd.n4663 99.6594
R7113 gnd.n4667 gnd.n4666 99.6594
R7114 gnd.n4677 gnd.n4676 99.6594
R7115 gnd.n4686 gnd.n4685 99.6594
R7116 gnd.n4689 gnd.n4688 99.6594
R7117 gnd.n4700 gnd.n4699 99.6594
R7118 gnd.n4709 gnd.n4708 99.6594
R7119 gnd.n4712 gnd.n4711 99.6594
R7120 gnd.n4723 gnd.n4722 99.6594
R7121 gnd.n4095 gnd.n3635 99.6594
R7122 gnd.n4094 gnd.n4093 99.6594
R7123 gnd.n4087 gnd.n3638 99.6594
R7124 gnd.n4086 gnd.n4085 99.6594
R7125 gnd.n4079 gnd.n3644 99.6594
R7126 gnd.n4078 gnd.n4077 99.6594
R7127 gnd.n4071 gnd.n3650 99.6594
R7128 gnd.n4070 gnd.n4069 99.6594
R7129 gnd.n4059 gnd.n3656 99.6594
R7130 gnd.n4096 gnd.n4095 99.6594
R7131 gnd.n4093 gnd.n4092 99.6594
R7132 gnd.n4088 gnd.n4087 99.6594
R7133 gnd.n4085 gnd.n4084 99.6594
R7134 gnd.n4080 gnd.n4079 99.6594
R7135 gnd.n4077 gnd.n4076 99.6594
R7136 gnd.n4072 gnd.n4071 99.6594
R7137 gnd.n4069 gnd.n4068 99.6594
R7138 gnd.n4060 gnd.n4059 99.6594
R7139 gnd.n2777 gnd.n2700 99.6594
R7140 gnd.n2769 gnd.n2688 99.6594
R7141 gnd.n2765 gnd.n2689 99.6594
R7142 gnd.n2761 gnd.n2690 99.6594
R7143 gnd.n2757 gnd.n2691 99.6594
R7144 gnd.n2753 gnd.n2692 99.6594
R7145 gnd.n2749 gnd.n2693 99.6594
R7146 gnd.n2745 gnd.n2694 99.6594
R7147 gnd.n2741 gnd.n2695 99.6594
R7148 gnd.n2737 gnd.n2696 99.6594
R7149 gnd.n2733 gnd.n2697 99.6594
R7150 gnd.n2729 gnd.n2698 99.6594
R7151 gnd.n2780 gnd.n2779 99.6594
R7152 gnd.n3544 gnd.n2171 99.6594
R7153 gnd.n3548 gnd.n2170 99.6594
R7154 gnd.n3552 gnd.n2169 99.6594
R7155 gnd.n3556 gnd.n2168 99.6594
R7156 gnd.n3560 gnd.n2167 99.6594
R7157 gnd.n3564 gnd.n2166 99.6594
R7158 gnd.n3568 gnd.n2165 99.6594
R7159 gnd.n3572 gnd.n2164 99.6594
R7160 gnd.n3576 gnd.n2163 99.6594
R7161 gnd.n3580 gnd.n2162 99.6594
R7162 gnd.n3584 gnd.n2161 99.6594
R7163 gnd.n3588 gnd.n2160 99.6594
R7164 gnd.n2200 gnd.n2159 99.6594
R7165 gnd.n2863 gnd.n2862 99.6594
R7166 gnd.n2622 gnd.n2600 99.6594
R7167 gnd.n2628 gnd.n2601 99.6594
R7168 gnd.n2632 gnd.n2602 99.6594
R7169 gnd.n2638 gnd.n2603 99.6594
R7170 gnd.n2642 gnd.n2604 99.6594
R7171 gnd.n2648 gnd.n2605 99.6594
R7172 gnd.n2606 gnd.n2590 99.6594
R7173 gnd.n3598 gnd.n2172 99.6594
R7174 gnd.n3602 gnd.n2173 99.6594
R7175 gnd.n3606 gnd.n2174 99.6594
R7176 gnd.n3610 gnd.n2175 99.6594
R7177 gnd.n3614 gnd.n2176 99.6594
R7178 gnd.n3618 gnd.n2177 99.6594
R7179 gnd.n3622 gnd.n2178 99.6594
R7180 gnd.n2181 gnd.n2179 99.6594
R7181 gnd.n3775 gnd.n3774 99.6594
R7182 gnd.n3783 gnd.n3782 99.6594
R7183 gnd.n3784 gnd.n3767 99.6594
R7184 gnd.n3793 gnd.n3792 99.6594
R7185 gnd.n3794 gnd.n3763 99.6594
R7186 gnd.n3803 gnd.n3802 99.6594
R7187 gnd.n3804 gnd.n3759 99.6594
R7188 gnd.n3813 gnd.n3812 99.6594
R7189 gnd.n3814 gnd.n3752 99.6594
R7190 gnd.n3823 gnd.n3822 99.6594
R7191 gnd.n3824 gnd.n3748 99.6594
R7192 gnd.n3833 gnd.n3832 99.6594
R7193 gnd.n3834 gnd.n3744 99.6594
R7194 gnd.n3843 gnd.n3842 99.6594
R7195 gnd.n3844 gnd.n3740 99.6594
R7196 gnd.n3853 gnd.n3852 99.6594
R7197 gnd.n3854 gnd.n3736 99.6594
R7198 gnd.n3864 gnd.n3863 99.6594
R7199 gnd.n3867 gnd.n3866 99.6594
R7200 gnd.n4532 gnd.n4284 99.6594
R7201 gnd.n4524 gnd.n1948 99.6594
R7202 gnd.n4520 gnd.n1949 99.6594
R7203 gnd.n4516 gnd.n1950 99.6594
R7204 gnd.n4512 gnd.n1951 99.6594
R7205 gnd.n4508 gnd.n1952 99.6594
R7206 gnd.n4504 gnd.n1953 99.6594
R7207 gnd.n4500 gnd.n1954 99.6594
R7208 gnd.n4496 gnd.n1955 99.6594
R7209 gnd.n4492 gnd.n1956 99.6594
R7210 gnd.n4488 gnd.n1957 99.6594
R7211 gnd.n4484 gnd.n1958 99.6594
R7212 gnd.n4480 gnd.n1959 99.6594
R7213 gnd.n4476 gnd.n1960 99.6594
R7214 gnd.n4472 gnd.n1961 99.6594
R7215 gnd.n4468 gnd.n1962 99.6594
R7216 gnd.n4464 gnd.n1963 99.6594
R7217 gnd.n4460 gnd.n1964 99.6594
R7218 gnd.n4456 gnd.n1965 99.6594
R7219 gnd.n4452 gnd.n1966 99.6594
R7220 gnd.n4448 gnd.n1967 99.6594
R7221 gnd.n4444 gnd.n1968 99.6594
R7222 gnd.n4440 gnd.n1969 99.6594
R7223 gnd.n4436 gnd.n1970 99.6594
R7224 gnd.n4432 gnd.n1971 99.6594
R7225 gnd.n4428 gnd.n1972 99.6594
R7226 gnd.n4424 gnd.n1973 99.6594
R7227 gnd.n4420 gnd.n1974 99.6594
R7228 gnd.n4416 gnd.n1975 99.6594
R7229 gnd.n4412 gnd.n1976 99.6594
R7230 gnd.n4408 gnd.n1977 99.6594
R7231 gnd.n4404 gnd.n1978 99.6594
R7232 gnd.n4400 gnd.n1979 99.6594
R7233 gnd.n4396 gnd.n1980 99.6594
R7234 gnd.n4392 gnd.n1981 99.6594
R7235 gnd.n4388 gnd.n1982 99.6594
R7236 gnd.n4384 gnd.n1983 99.6594
R7237 gnd.n4380 gnd.n1984 99.6594
R7238 gnd.n4376 gnd.n1985 99.6594
R7239 gnd.n4372 gnd.n1986 99.6594
R7240 gnd.n4368 gnd.n1987 99.6594
R7241 gnd.n4535 gnd.n4534 99.6594
R7242 gnd.n4722 gnd.n4721 99.6594
R7243 gnd.n4711 gnd.n4710 99.6594
R7244 gnd.n4708 gnd.n4701 99.6594
R7245 gnd.n4699 gnd.n4698 99.6594
R7246 gnd.n4688 gnd.n4687 99.6594
R7247 gnd.n4685 gnd.n4678 99.6594
R7248 gnd.n4676 gnd.n4675 99.6594
R7249 gnd.n4666 gnd.n4665 99.6594
R7250 gnd.n4663 gnd.n4662 99.6594
R7251 gnd.n530 gnd.n461 99.6594
R7252 gnd.n532 gnd.n468 99.6594
R7253 gnd.n534 gnd.n533 99.6594
R7254 gnd.n535 gnd.n477 99.6594
R7255 gnd.n537 gnd.n484 99.6594
R7256 gnd.n539 gnd.n538 99.6594
R7257 gnd.n540 gnd.n493 99.6594
R7258 gnd.n542 gnd.n500 99.6594
R7259 gnd.n543 gnd.n510 99.6594
R7260 gnd.n7504 gnd.n125 99.6594
R7261 gnd.n7503 gnd.n7502 99.6594
R7262 gnd.n7499 gnd.n7498 99.6594
R7263 gnd.n7496 gnd.n7495 99.6594
R7264 gnd.n7491 gnd.n7490 99.6594
R7265 gnd.n7488 gnd.n7487 99.6594
R7266 gnd.n7483 gnd.n7482 99.6594
R7267 gnd.n7480 gnd.n7479 99.6594
R7268 gnd.n7475 gnd.n7474 99.6594
R7269 gnd.n6187 gnd.n6186 99.6594
R7270 gnd.n1160 gnd.n1152 99.6594
R7271 gnd.n6194 gnd.n6193 99.6594
R7272 gnd.n1151 gnd.n1145 99.6594
R7273 gnd.n6201 gnd.n6200 99.6594
R7274 gnd.n1144 gnd.n1138 99.6594
R7275 gnd.n6208 gnd.n6207 99.6594
R7276 gnd.n1137 gnd.n1131 99.6594
R7277 gnd.n6215 gnd.n6214 99.6594
R7278 gnd.n1130 gnd.n1123 99.6594
R7279 gnd.n6224 gnd.n6223 99.6594
R7280 gnd.n1119 gnd.n1113 99.6594
R7281 gnd.n6231 gnd.n6230 99.6594
R7282 gnd.n1112 gnd.n1106 99.6594
R7283 gnd.n6238 gnd.n6237 99.6594
R7284 gnd.n1105 gnd.n1098 99.6594
R7285 gnd.n6245 gnd.n6244 99.6594
R7286 gnd.n6248 gnd.n6247 99.6594
R7287 gnd.n7177 gnd.n7176 99.6594
R7288 gnd.n7170 gnd.n512 99.6594
R7289 gnd.n7166 gnd.n513 99.6594
R7290 gnd.n7162 gnd.n514 99.6594
R7291 gnd.n7158 gnd.n515 99.6594
R7292 gnd.n7154 gnd.n516 99.6594
R7293 gnd.n7150 gnd.n517 99.6594
R7294 gnd.n7145 gnd.n519 99.6594
R7295 gnd.n7141 gnd.n520 99.6594
R7296 gnd.n7137 gnd.n521 99.6594
R7297 gnd.n7133 gnd.n522 99.6594
R7298 gnd.n7129 gnd.n523 99.6594
R7299 gnd.n7125 gnd.n524 99.6594
R7300 gnd.n7121 gnd.n525 99.6594
R7301 gnd.n7117 gnd.n526 99.6594
R7302 gnd.n7113 gnd.n527 99.6594
R7303 gnd.n584 gnd.n528 99.6594
R7304 gnd.n7105 gnd.n529 99.6594
R7305 gnd.n198 gnd.n195 99.6594
R7306 gnd.n7561 gnd.n7560 99.6594
R7307 gnd.n194 gnd.n188 99.6594
R7308 gnd.n7568 gnd.n7567 99.6594
R7309 gnd.n187 gnd.n181 99.6594
R7310 gnd.n7575 gnd.n7574 99.6594
R7311 gnd.n180 gnd.n174 99.6594
R7312 gnd.n7582 gnd.n7581 99.6594
R7313 gnd.n173 gnd.n167 99.6594
R7314 gnd.n7589 gnd.n7588 99.6594
R7315 gnd.n166 gnd.n160 99.6594
R7316 gnd.n7599 gnd.n7598 99.6594
R7317 gnd.n159 gnd.n153 99.6594
R7318 gnd.n7606 gnd.n7605 99.6594
R7319 gnd.n152 gnd.n146 99.6594
R7320 gnd.n7613 gnd.n7612 99.6594
R7321 gnd.n145 gnd.n139 99.6594
R7322 gnd.n7620 gnd.n7619 99.6594
R7323 gnd.n138 gnd.n135 99.6594
R7324 gnd.n4770 gnd.n4769 99.6594
R7325 gnd.n4670 gnd.n4635 99.6594
R7326 gnd.n4672 gnd.n4636 99.6594
R7327 gnd.n4682 gnd.n4637 99.6594
R7328 gnd.n4693 gnd.n4638 99.6594
R7329 gnd.n4695 gnd.n4639 99.6594
R7330 gnd.n4705 gnd.n4640 99.6594
R7331 gnd.n4718 gnd.n4641 99.6594
R7332 gnd.n4719 gnd.n4642 99.6594
R7333 gnd.n4643 gnd.n1172 99.6594
R7334 gnd.n4645 gnd.n4644 99.6594
R7335 gnd.n4646 gnd.n1177 99.6594
R7336 gnd.n4647 gnd.n1183 99.6594
R7337 gnd.n4649 gnd.n1185 99.6594
R7338 gnd.n4770 gnd.n4651 99.6594
R7339 gnd.n4671 gnd.n4635 99.6594
R7340 gnd.n4681 gnd.n4636 99.6594
R7341 gnd.n4692 gnd.n4637 99.6594
R7342 gnd.n4694 gnd.n4638 99.6594
R7343 gnd.n4704 gnd.n4639 99.6594
R7344 gnd.n4717 gnd.n4640 99.6594
R7345 gnd.n4720 gnd.n4641 99.6594
R7346 gnd.n4642 gnd.n1171 99.6594
R7347 gnd.n4643 gnd.n1173 99.6594
R7348 gnd.n4645 gnd.n1176 99.6594
R7349 gnd.n4646 gnd.n1178 99.6594
R7350 gnd.n4647 gnd.n1184 99.6594
R7351 gnd.n4649 gnd.n4648 99.6594
R7352 gnd.n5821 gnd.n465 99.6594
R7353 gnd.n5823 gnd.n472 99.6594
R7354 gnd.n5825 gnd.n5824 99.6594
R7355 gnd.n5826 gnd.n481 99.6594
R7356 gnd.n5828 gnd.n488 99.6594
R7357 gnd.n5830 gnd.n5829 99.6594
R7358 gnd.n5831 gnd.n497 99.6594
R7359 gnd.n5833 gnd.n506 99.6594
R7360 gnd.n5934 gnd.n5834 99.6594
R7361 gnd.n5937 gnd.n5835 99.6594
R7362 gnd.n5939 gnd.n5836 99.6594
R7363 gnd.n5943 gnd.n5837 99.6594
R7364 gnd.n5945 gnd.n5838 99.6594
R7365 gnd.n5949 gnd.n5839 99.6594
R7366 gnd.n5946 gnd.n5839 99.6594
R7367 gnd.n5944 gnd.n5838 99.6594
R7368 gnd.n5940 gnd.n5837 99.6594
R7369 gnd.n5938 gnd.n5836 99.6594
R7370 gnd.n5935 gnd.n5835 99.6594
R7371 gnd.n5834 gnd.n507 99.6594
R7372 gnd.n5833 gnd.n5832 99.6594
R7373 gnd.n5831 gnd.n496 99.6594
R7374 gnd.n5830 gnd.n489 99.6594
R7375 gnd.n5828 gnd.n5827 99.6594
R7376 gnd.n5826 gnd.n480 99.6594
R7377 gnd.n5825 gnd.n473 99.6594
R7378 gnd.n5823 gnd.n5822 99.6594
R7379 gnd.n5821 gnd.n464 99.6594
R7380 gnd.n1179 gnd.t273 98.63
R7381 gnd.n564 gnd.t269 98.63
R7382 gnd.n586 gnd.t248 98.63
R7383 gnd.n201 gnd.t314 98.63
R7384 gnd.n7592 gnd.t229 98.63
R7385 gnd.n122 gnd.t285 98.63
R7386 gnd.n502 gnd.t298 98.63
R7387 gnd.n4713 gnd.t321 98.63
R7388 gnd.n1157 gnd.t324 98.63
R7389 gnd.n1120 gnd.t243 98.63
R7390 gnd.n3756 gnd.t331 98.63
R7391 gnd.n3732 gnd.t312 98.63
R7392 gnd.n3659 gnd.t328 98.63
R7393 gnd.n5956 gnd.t239 98.63
R7394 gnd.n4941 gnd.t305 92.8196
R7395 gnd.n1454 gnd.t258 92.8196
R7396 gnd.n4938 gnd.t252 92.8118
R7397 gnd.n1448 gnd.t294 92.8118
R7398 gnd.n6318 gnd.n6317 90.3496
R7399 gnd.n4925 gnd.n4924 81.8399
R7400 gnd.n6709 gnd.n6708 75.227
R7401 gnd.n6710 gnd.n6709 75.227
R7402 gnd.n6710 gnd.n740 75.227
R7403 gnd.n6718 gnd.n740 75.227
R7404 gnd.n6719 gnd.n6718 75.227
R7405 gnd.n6720 gnd.n6719 75.227
R7406 gnd.n6720 gnd.n734 75.227
R7407 gnd.n6728 gnd.n734 75.227
R7408 gnd.n6729 gnd.n6728 75.227
R7409 gnd.n6730 gnd.n6729 75.227
R7410 gnd.n6730 gnd.n728 75.227
R7411 gnd.n6738 gnd.n728 75.227
R7412 gnd.n6739 gnd.n6738 75.227
R7413 gnd.n6740 gnd.n6739 75.227
R7414 gnd.n6740 gnd.n722 75.227
R7415 gnd.n6748 gnd.n722 75.227
R7416 gnd.n6749 gnd.n6748 75.227
R7417 gnd.n6750 gnd.n6749 75.227
R7418 gnd.n6750 gnd.n716 75.227
R7419 gnd.n6758 gnd.n716 75.227
R7420 gnd.n6759 gnd.n6758 75.227
R7421 gnd.n6760 gnd.n6759 75.227
R7422 gnd.n6760 gnd.n710 75.227
R7423 gnd.n6768 gnd.n710 75.227
R7424 gnd.n6769 gnd.n6768 75.227
R7425 gnd.n6770 gnd.n6769 75.227
R7426 gnd.n6770 gnd.n704 75.227
R7427 gnd.n6778 gnd.n704 75.227
R7428 gnd.n6779 gnd.n6778 75.227
R7429 gnd.n6780 gnd.n6779 75.227
R7430 gnd.n6780 gnd.n698 75.227
R7431 gnd.n6788 gnd.n698 75.227
R7432 gnd.n6789 gnd.n6788 75.227
R7433 gnd.n6790 gnd.n6789 75.227
R7434 gnd.n6790 gnd.n692 75.227
R7435 gnd.n6798 gnd.n692 75.227
R7436 gnd.n6799 gnd.n6798 75.227
R7437 gnd.n6800 gnd.n6799 75.227
R7438 gnd.n6800 gnd.n686 75.227
R7439 gnd.n6808 gnd.n686 75.227
R7440 gnd.n6809 gnd.n6808 75.227
R7441 gnd.n6810 gnd.n6809 75.227
R7442 gnd.n6810 gnd.n680 75.227
R7443 gnd.n6818 gnd.n680 75.227
R7444 gnd.n6819 gnd.n6818 75.227
R7445 gnd.n6820 gnd.n6819 75.227
R7446 gnd.n6820 gnd.n674 75.227
R7447 gnd.n6828 gnd.n674 75.227
R7448 gnd.n6829 gnd.n6828 75.227
R7449 gnd.n6830 gnd.n6829 75.227
R7450 gnd.n6830 gnd.n668 75.227
R7451 gnd.n6838 gnd.n668 75.227
R7452 gnd.n6839 gnd.n6838 75.227
R7453 gnd.n6840 gnd.n6839 75.227
R7454 gnd.n6840 gnd.n662 75.227
R7455 gnd.n6848 gnd.n662 75.227
R7456 gnd.n6849 gnd.n6848 75.227
R7457 gnd.n6850 gnd.n6849 75.227
R7458 gnd.n6850 gnd.n656 75.227
R7459 gnd.n6858 gnd.n656 75.227
R7460 gnd.n6859 gnd.n6858 75.227
R7461 gnd.n6860 gnd.n6859 75.227
R7462 gnd.n6860 gnd.n650 75.227
R7463 gnd.n6868 gnd.n650 75.227
R7464 gnd.n6869 gnd.n6868 75.227
R7465 gnd.n6870 gnd.n6869 75.227
R7466 gnd.n6870 gnd.n644 75.227
R7467 gnd.n6878 gnd.n644 75.227
R7468 gnd.n6879 gnd.n6878 75.227
R7469 gnd.n6880 gnd.n6879 75.227
R7470 gnd.n6880 gnd.n638 75.227
R7471 gnd.n6888 gnd.n638 75.227
R7472 gnd.n6889 gnd.n6888 75.227
R7473 gnd.n6890 gnd.n6889 75.227
R7474 gnd.n6890 gnd.n632 75.227
R7475 gnd.n6898 gnd.n632 75.227
R7476 gnd.n6899 gnd.n6898 75.227
R7477 gnd.n6900 gnd.n6899 75.227
R7478 gnd.n6900 gnd.n626 75.227
R7479 gnd.n6908 gnd.n626 75.227
R7480 gnd.n6909 gnd.n6908 75.227
R7481 gnd.n6911 gnd.n6909 75.227
R7482 gnd.n6911 gnd.n6910 75.227
R7483 gnd.n2651 gnd.t318 74.8376
R7484 gnd.n2197 gnd.t263 74.8376
R7485 gnd.n4942 gnd.t304 72.8438
R7486 gnd.n1455 gnd.t259 72.8438
R7487 gnd.n4926 gnd.n4919 72.8411
R7488 gnd.n4932 gnd.n4917 72.8411
R7489 gnd.n1423 gnd.n1422 72.8411
R7490 gnd.n1180 gnd.t272 72.836
R7491 gnd.n4939 gnd.t251 72.836
R7492 gnd.n1449 gnd.t295 72.836
R7493 gnd.n565 gnd.t268 72.836
R7494 gnd.n587 gnd.t247 72.836
R7495 gnd.n202 gnd.t315 72.836
R7496 gnd.n7593 gnd.t230 72.836
R7497 gnd.n123 gnd.t286 72.836
R7498 gnd.n503 gnd.t297 72.836
R7499 gnd.n4714 gnd.t322 72.836
R7500 gnd.n1158 gnd.t325 72.836
R7501 gnd.n1121 gnd.t244 72.836
R7502 gnd.n3757 gnd.t330 72.836
R7503 gnd.n3733 gnd.t311 72.836
R7504 gnd.n3660 gnd.t327 72.836
R7505 gnd.n5957 gnd.t240 72.836
R7506 gnd.n5707 gnd.n5706 71.676
R7507 gnd.n5704 gnd.n5703 71.676
R7508 gnd.n5699 gnd.n1431 71.676
R7509 gnd.n5697 gnd.n5696 71.676
R7510 gnd.n5692 gnd.n1434 71.676
R7511 gnd.n5690 gnd.n5689 71.676
R7512 gnd.n5685 gnd.n1437 71.676
R7513 gnd.n5683 gnd.n5682 71.676
R7514 gnd.n5678 gnd.n1440 71.676
R7515 gnd.n5676 gnd.n5675 71.676
R7516 gnd.n5671 gnd.n1443 71.676
R7517 gnd.n5669 gnd.n5668 71.676
R7518 gnd.n5664 gnd.n1446 71.676
R7519 gnd.n5662 gnd.n5661 71.676
R7520 gnd.n5656 gnd.n1451 71.676
R7521 gnd.n5654 gnd.n5653 71.676
R7522 gnd.n5649 gnd.n5648 71.676
R7523 gnd.n5646 gnd.n5645 71.676
R7524 gnd.n5640 gnd.n1457 71.676
R7525 gnd.n5638 gnd.n5637 71.676
R7526 gnd.n5633 gnd.n1460 71.676
R7527 gnd.n5631 gnd.n5630 71.676
R7528 gnd.n5626 gnd.n1463 71.676
R7529 gnd.n5624 gnd.n5623 71.676
R7530 gnd.n5619 gnd.n1466 71.676
R7531 gnd.n5617 gnd.n5616 71.676
R7532 gnd.n5612 gnd.n1469 71.676
R7533 gnd.n5610 gnd.n5609 71.676
R7534 gnd.n5605 gnd.n1472 71.676
R7535 gnd.n5603 gnd.n5602 71.676
R7536 gnd.n5598 gnd.n1475 71.676
R7537 gnd.n5596 gnd.n5595 71.676
R7538 gnd.n5591 gnd.n5589 71.676
R7539 gnd.n5076 gnd.n5075 71.676
R7540 gnd.n5070 gnd.n4879 71.676
R7541 gnd.n5067 gnd.n4880 71.676
R7542 gnd.n5063 gnd.n4881 71.676
R7543 gnd.n5059 gnd.n4882 71.676
R7544 gnd.n5055 gnd.n4883 71.676
R7545 gnd.n5051 gnd.n4884 71.676
R7546 gnd.n5047 gnd.n4885 71.676
R7547 gnd.n5043 gnd.n4886 71.676
R7548 gnd.n5039 gnd.n4887 71.676
R7549 gnd.n5035 gnd.n4888 71.676
R7550 gnd.n5031 gnd.n4889 71.676
R7551 gnd.n5027 gnd.n4890 71.676
R7552 gnd.n5023 gnd.n4891 71.676
R7553 gnd.n5019 gnd.n4892 71.676
R7554 gnd.n5015 gnd.n4893 71.676
R7555 gnd.n5011 gnd.n4895 71.676
R7556 gnd.n5006 gnd.n4896 71.676
R7557 gnd.n5001 gnd.n4897 71.676
R7558 gnd.n4997 gnd.n4898 71.676
R7559 gnd.n4993 gnd.n4899 71.676
R7560 gnd.n4989 gnd.n4900 71.676
R7561 gnd.n4985 gnd.n4901 71.676
R7562 gnd.n4981 gnd.n4902 71.676
R7563 gnd.n4977 gnd.n4903 71.676
R7564 gnd.n4973 gnd.n4904 71.676
R7565 gnd.n4969 gnd.n4905 71.676
R7566 gnd.n4965 gnd.n4906 71.676
R7567 gnd.n4961 gnd.n4907 71.676
R7568 gnd.n4957 gnd.n4908 71.676
R7569 gnd.n4953 gnd.n4909 71.676
R7570 gnd.n4949 gnd.n4910 71.676
R7571 gnd.n5076 gnd.n4914 71.676
R7572 gnd.n5068 gnd.n4879 71.676
R7573 gnd.n5064 gnd.n4880 71.676
R7574 gnd.n5060 gnd.n4881 71.676
R7575 gnd.n5056 gnd.n4882 71.676
R7576 gnd.n5052 gnd.n4883 71.676
R7577 gnd.n5048 gnd.n4884 71.676
R7578 gnd.n5044 gnd.n4885 71.676
R7579 gnd.n5040 gnd.n4886 71.676
R7580 gnd.n5036 gnd.n4887 71.676
R7581 gnd.n5032 gnd.n4888 71.676
R7582 gnd.n5028 gnd.n4889 71.676
R7583 gnd.n5024 gnd.n4890 71.676
R7584 gnd.n5020 gnd.n4891 71.676
R7585 gnd.n5016 gnd.n4892 71.676
R7586 gnd.n5012 gnd.n4894 71.676
R7587 gnd.n5007 gnd.n4895 71.676
R7588 gnd.n5002 gnd.n4896 71.676
R7589 gnd.n4998 gnd.n4897 71.676
R7590 gnd.n4994 gnd.n4898 71.676
R7591 gnd.n4990 gnd.n4899 71.676
R7592 gnd.n4986 gnd.n4900 71.676
R7593 gnd.n4982 gnd.n4901 71.676
R7594 gnd.n4978 gnd.n4902 71.676
R7595 gnd.n4974 gnd.n4903 71.676
R7596 gnd.n4970 gnd.n4904 71.676
R7597 gnd.n4966 gnd.n4905 71.676
R7598 gnd.n4962 gnd.n4906 71.676
R7599 gnd.n4958 gnd.n4907 71.676
R7600 gnd.n4954 gnd.n4908 71.676
R7601 gnd.n4950 gnd.n4909 71.676
R7602 gnd.n4946 gnd.n4910 71.676
R7603 gnd.n5589 gnd.n1476 71.676
R7604 gnd.n5597 gnd.n5596 71.676
R7605 gnd.n1475 gnd.n1473 71.676
R7606 gnd.n5604 gnd.n5603 71.676
R7607 gnd.n1472 gnd.n1470 71.676
R7608 gnd.n5611 gnd.n5610 71.676
R7609 gnd.n1469 gnd.n1467 71.676
R7610 gnd.n5618 gnd.n5617 71.676
R7611 gnd.n1466 gnd.n1464 71.676
R7612 gnd.n5625 gnd.n5624 71.676
R7613 gnd.n1463 gnd.n1461 71.676
R7614 gnd.n5632 gnd.n5631 71.676
R7615 gnd.n1460 gnd.n1458 71.676
R7616 gnd.n5639 gnd.n5638 71.676
R7617 gnd.n1457 gnd.n1453 71.676
R7618 gnd.n5647 gnd.n5646 71.676
R7619 gnd.n5651 gnd.n5650 71.676
R7620 gnd.n5655 gnd.n5654 71.676
R7621 gnd.n1451 gnd.n1447 71.676
R7622 gnd.n5663 gnd.n5662 71.676
R7623 gnd.n1446 gnd.n1444 71.676
R7624 gnd.n5670 gnd.n5669 71.676
R7625 gnd.n1443 gnd.n1441 71.676
R7626 gnd.n5677 gnd.n5676 71.676
R7627 gnd.n1440 gnd.n1438 71.676
R7628 gnd.n5684 gnd.n5683 71.676
R7629 gnd.n1437 gnd.n1435 71.676
R7630 gnd.n5691 gnd.n5690 71.676
R7631 gnd.n1434 gnd.n1432 71.676
R7632 gnd.n5698 gnd.n5697 71.676
R7633 gnd.n1431 gnd.n1429 71.676
R7634 gnd.n5705 gnd.n5704 71.676
R7635 gnd.n5708 gnd.n5707 71.676
R7636 gnd.n10 gnd.t126 69.1507
R7637 gnd.n18 gnd.t199 68.4792
R7638 gnd.n17 gnd.t221 68.4792
R7639 gnd.n16 gnd.t356 68.4792
R7640 gnd.n15 gnd.t132 68.4792
R7641 gnd.n14 gnd.t19 68.4792
R7642 gnd.n13 gnd.t183 68.4792
R7643 gnd.n12 gnd.t197 68.4792
R7644 gnd.n11 gnd.t21 68.4792
R7645 gnd.n10 gnd.t48 68.4792
R7646 gnd.n5004 gnd.n4942 59.5399
R7647 gnd.n5642 gnd.n1455 59.5399
R7648 gnd.n4940 gnd.n4939 59.5399
R7649 gnd.n5658 gnd.n1449 59.5399
R7650 gnd.n4937 gnd.n4935 59.1804
R7651 gnd.n2429 gnd.t111 56.607
R7652 gnd.n60 gnd.t62 56.607
R7653 gnd.n2390 gnd.t144 56.407
R7654 gnd.n2409 gnd.t176 56.407
R7655 gnd.n21 gnd.t351 56.407
R7656 gnd.n40 gnd.t28 56.407
R7657 gnd.n2446 gnd.t209 55.8337
R7658 gnd.n2407 gnd.t226 55.8337
R7659 gnd.n2426 gnd.t143 55.8337
R7660 gnd.n77 gnd.t219 55.8337
R7661 gnd.n38 gnd.t352 55.8337
R7662 gnd.n57 gnd.t120 55.8337
R7663 gnd.n4923 gnd.n4922 54.358
R7664 gnd.n1420 gnd.n1419 54.358
R7665 gnd.n2429 gnd.n2428 53.0052
R7666 gnd.n2431 gnd.n2430 53.0052
R7667 gnd.n2433 gnd.n2432 53.0052
R7668 gnd.n2435 gnd.n2434 53.0052
R7669 gnd.n2437 gnd.n2436 53.0052
R7670 gnd.n2439 gnd.n2438 53.0052
R7671 gnd.n2441 gnd.n2440 53.0052
R7672 gnd.n2443 gnd.n2442 53.0052
R7673 gnd.n2445 gnd.n2444 53.0052
R7674 gnd.n2390 gnd.n2389 53.0052
R7675 gnd.n2392 gnd.n2391 53.0052
R7676 gnd.n2394 gnd.n2393 53.0052
R7677 gnd.n2396 gnd.n2395 53.0052
R7678 gnd.n2398 gnd.n2397 53.0052
R7679 gnd.n2400 gnd.n2399 53.0052
R7680 gnd.n2402 gnd.n2401 53.0052
R7681 gnd.n2404 gnd.n2403 53.0052
R7682 gnd.n2406 gnd.n2405 53.0052
R7683 gnd.n2409 gnd.n2408 53.0052
R7684 gnd.n2411 gnd.n2410 53.0052
R7685 gnd.n2413 gnd.n2412 53.0052
R7686 gnd.n2415 gnd.n2414 53.0052
R7687 gnd.n2417 gnd.n2416 53.0052
R7688 gnd.n2419 gnd.n2418 53.0052
R7689 gnd.n2421 gnd.n2420 53.0052
R7690 gnd.n2423 gnd.n2422 53.0052
R7691 gnd.n2425 gnd.n2424 53.0052
R7692 gnd.n76 gnd.n75 53.0052
R7693 gnd.n74 gnd.n73 53.0052
R7694 gnd.n72 gnd.n71 53.0052
R7695 gnd.n70 gnd.n69 53.0052
R7696 gnd.n68 gnd.n67 53.0052
R7697 gnd.n66 gnd.n65 53.0052
R7698 gnd.n64 gnd.n63 53.0052
R7699 gnd.n62 gnd.n61 53.0052
R7700 gnd.n60 gnd.n59 53.0052
R7701 gnd.n37 gnd.n36 53.0052
R7702 gnd.n35 gnd.n34 53.0052
R7703 gnd.n33 gnd.n32 53.0052
R7704 gnd.n31 gnd.n30 53.0052
R7705 gnd.n29 gnd.n28 53.0052
R7706 gnd.n27 gnd.n26 53.0052
R7707 gnd.n25 gnd.n24 53.0052
R7708 gnd.n23 gnd.n22 53.0052
R7709 gnd.n21 gnd.n20 53.0052
R7710 gnd.n56 gnd.n55 53.0052
R7711 gnd.n54 gnd.n53 53.0052
R7712 gnd.n52 gnd.n51 53.0052
R7713 gnd.n50 gnd.n49 53.0052
R7714 gnd.n48 gnd.n47 53.0052
R7715 gnd.n46 gnd.n45 53.0052
R7716 gnd.n44 gnd.n43 53.0052
R7717 gnd.n42 gnd.n41 53.0052
R7718 gnd.n40 gnd.n39 53.0052
R7719 gnd.n1411 gnd.n1410 52.4801
R7720 gnd.n3482 gnd.t38 52.3082
R7721 gnd.n3450 gnd.t165 52.3082
R7722 gnd.n3418 gnd.t336 52.3082
R7723 gnd.n3387 gnd.t9 52.3082
R7724 gnd.n3355 gnd.t91 52.3082
R7725 gnd.n3323 gnd.t115 52.3082
R7726 gnd.n3291 gnd.t161 52.3082
R7727 gnd.n3260 gnd.t181 52.3082
R7728 gnd.n7629 gnd.n128 51.6227
R7729 gnd.n3312 gnd.n3280 51.4173
R7730 gnd.n3376 gnd.n3375 50.455
R7731 gnd.n3344 gnd.n3343 50.455
R7732 gnd.n3312 gnd.n3311 50.455
R7733 gnd.n2725 gnd.n2724 45.1884
R7734 gnd.n2223 gnd.n2222 45.1884
R7735 gnd.n6910 gnd.n252 45.1364
R7736 gnd.n5710 gnd.n1426 44.3322
R7737 gnd.n4926 gnd.n4925 44.3189
R7738 gnd.n1181 gnd.n1180 42.4732
R7739 gnd.n5958 gnd.n5957 42.4732
R7740 gnd.n588 gnd.n587 42.2793
R7741 gnd.n7557 gnd.n202 42.2793
R7742 gnd.n7594 gnd.n7593 42.2793
R7743 gnd.n124 gnd.n123 42.2793
R7744 gnd.n504 gnd.n503 42.2793
R7745 gnd.n4715 gnd.n4714 42.2793
R7746 gnd.n2726 gnd.n2725 42.2793
R7747 gnd.n2224 gnd.n2223 42.2793
R7748 gnd.n2652 gnd.n2651 42.2793
R7749 gnd.n3597 gnd.n2197 42.2793
R7750 gnd.n1159 gnd.n1158 42.2793
R7751 gnd.n3758 gnd.n3757 42.2793
R7752 gnd.n3734 gnd.n3733 42.2793
R7753 gnd.n3661 gnd.n3660 42.2793
R7754 gnd.n4924 gnd.n4923 41.6274
R7755 gnd.n1421 gnd.n1420 41.6274
R7756 gnd.n4933 gnd.n4932 40.8975
R7757 gnd.n1424 gnd.n1423 40.8975
R7758 gnd.n7147 gnd.n565 36.9518
R7759 gnd.n1122 gnd.n1121 36.9518
R7760 gnd.n2778 gnd.n2682 36.8252
R7761 gnd.n4932 gnd.n4931 35.055
R7762 gnd.n4927 gnd.n4926 35.055
R7763 gnd.n1413 gnd.n1412 35.055
R7764 gnd.n1423 gnd.n1409 35.055
R7765 gnd.n3630 gnd.n2157 32.8146
R7766 gnd.n4633 gnd.n1904 31.8661
R7767 gnd.n4634 gnd.n4633 31.8661
R7768 gnd.n4773 gnd.n4772 31.8661
R7769 gnd.n5985 gnd.n1316 31.8661
R7770 gnd.n5983 gnd.n5982 31.8661
R7771 gnd.n5982 gnd.n511 31.8661
R7772 gnd.n7321 gnd.n362 31.8661
R7773 gnd.n7329 gnd.n353 31.8661
R7774 gnd.n7329 gnd.n356 31.8661
R7775 gnd.n7337 gnd.n338 31.8661
R7776 gnd.n7345 gnd.n338 31.8661
R7777 gnd.n7353 gnd.n330 31.8661
R7778 gnd.n7361 gnd.n320 31.8661
R7779 gnd.n7361 gnd.n323 31.8661
R7780 gnd.n7369 gnd.n314 31.8661
R7781 gnd.n7377 gnd.n299 31.8661
R7782 gnd.n7385 gnd.n299 31.8661
R7783 gnd.n7393 gnd.n290 31.8661
R7784 gnd.n7393 gnd.n293 31.8661
R7785 gnd.n7401 gnd.n284 31.8661
R7786 gnd.n7409 gnd.n269 31.8661
R7787 gnd.n7417 gnd.n269 31.8661
R7788 gnd.n7425 gnd.n260 31.8661
R7789 gnd.n7425 gnd.n263 31.8661
R7790 gnd.n7433 gnd.n254 31.8661
R7791 gnd.n7441 gnd.n238 31.8661
R7792 gnd.n7449 gnd.n238 31.8661
R7793 gnd.n7457 gnd.n229 31.8661
R7794 gnd.n7457 gnd.n232 31.8661
R7795 gnd.n7465 gnd.n213 31.8661
R7796 gnd.n7541 gnd.n213 31.8661
R7797 gnd.n7541 gnd.n206 31.8661
R7798 gnd.n7549 gnd.n206 31.8661
R7799 gnd.n7629 gnd.n126 31.8661
R7800 gnd.t68 gnd.n330 31.5474
R7801 gnd.n314 gnd.t15 31.5474
R7802 gnd.n284 gnd.t43 30.9101
R7803 gnd.n5592 gnd.n5588 30.7517
R7804 gnd.n4947 gnd.n4944 30.7517
R7805 gnd.n254 gnd.t178 30.2728
R7806 gnd.n4103 gnd.n3631 29.5331
R7807 gnd.t228 gnd.n126 28.3609
R7808 gnd.n1096 gnd.n1091 28.0422
R7809 gnd.n7178 gnd.n455 28.0422
R7810 gnd.n1180 gnd.n1179 25.7944
R7811 gnd.n565 gnd.n564 25.7944
R7812 gnd.n587 gnd.n586 25.7944
R7813 gnd.n202 gnd.n201 25.7944
R7814 gnd.n7593 gnd.n7592 25.7944
R7815 gnd.n123 gnd.n122 25.7944
R7816 gnd.n503 gnd.n502 25.7944
R7817 gnd.n4714 gnd.n4713 25.7944
R7818 gnd.n2651 gnd.n2650 25.7944
R7819 gnd.n2197 gnd.n2196 25.7944
R7820 gnd.n1158 gnd.n1157 25.7944
R7821 gnd.n1121 gnd.n1120 25.7944
R7822 gnd.n3757 gnd.n3756 25.7944
R7823 gnd.n3733 gnd.n3732 25.7944
R7824 gnd.n3660 gnd.n3659 25.7944
R7825 gnd.n5957 gnd.n5956 25.7944
R7826 gnd.n4771 gnd.n4634 23.8997
R7827 gnd.n5984 gnd.n5983 23.8997
R7828 gnd.n6315 gnd.n983 23.581
R7829 gnd.n3962 gnd.n993 23.581
R7830 gnd.n3967 gnd.n1004 23.581
R7831 gnd.n6303 gnd.n1007 23.581
R7832 gnd.n6297 gnd.n1018 23.581
R7833 gnd.n4563 gnd.n4562 23.581
R7834 gnd.n6291 gnd.n1028 23.581
R7835 gnd.n4571 gnd.n1036 23.581
R7836 gnd.n4606 gnd.n1046 23.581
R7837 gnd.n6279 gnd.n1049 23.581
R7838 gnd.n6273 gnd.n1060 23.581
R7839 gnd.n4583 gnd.n1068 23.581
R7840 gnd.n6267 gnd.n1071 23.581
R7841 gnd.n4592 gnd.n1079 23.581
R7842 gnd.n6178 gnd.n1088 23.581
R7843 gnd.n6255 gnd.n1091 23.581
R7844 gnd.n7233 gnd.n455 23.581
R7845 gnd.n5973 gnd.n458 23.581
R7846 gnd.n7098 gnd.n450 23.581
R7847 gnd.n7249 gnd.n439 23.581
R7848 gnd.n5866 gnd.n442 23.581
R7849 gnd.n7257 gnd.n430 23.581
R7850 gnd.n7265 gnd.n421 23.581
R7851 gnd.n5917 gnd.n424 23.581
R7852 gnd.n5911 gnd.n415 23.581
R7853 gnd.n7281 gnd.n405 23.581
R7854 gnd.n5907 gnd.n5906 23.581
R7855 gnd.n7289 gnd.n396 23.581
R7856 gnd.n7297 gnd.n387 23.581
R7857 gnd.n6928 gnd.n390 23.581
R7858 gnd.n7040 gnd.n381 23.581
R7859 gnd.n7313 gnd.n371 23.581
R7860 gnd.n6920 gnd.n362 23.581
R7861 gnd.n7465 gnd.t119 23.2624
R7862 gnd.n7401 gnd.t100 21.9878
R7863 gnd.n7353 gnd.t12 21.3504
R7864 gnd.n7369 gnd.t10 21.3504
R7865 gnd.n7337 gnd.t41 20.7131
R7866 gnd.n7385 gnd.t29 20.7131
R7867 gnd.n6309 gnd.t170 20.0758
R7868 gnd.n1164 gnd.t242 20.0758
R7869 gnd.n5974 gnd.t246 20.0758
R7870 gnd.n7305 gnd.t189 20.0758
R7871 gnd.n7417 gnd.t45 20.0758
R7872 gnd.n4942 gnd.n4941 19.9763
R7873 gnd.n1455 gnd.n1454 19.9763
R7874 gnd.n4939 gnd.n4938 19.9763
R7875 gnd.n1449 gnd.n1448 19.9763
R7876 gnd.n4920 gnd.t283 19.8005
R7877 gnd.n4920 gnd.t233 19.8005
R7878 gnd.n4921 gnd.t308 19.8005
R7879 gnd.n4921 gnd.t334 19.8005
R7880 gnd.n1417 gnd.t266 19.8005
R7881 gnd.n1417 gnd.t292 19.8005
R7882 gnd.n1418 gnd.t255 19.8005
R7883 gnd.n1418 gnd.t289 19.8005
R7884 gnd.n365 gnd.t72 19.7572
R7885 gnd.t39 gnd.n252 19.7572
R7886 gnd.n4917 gnd.n4916 19.5087
R7887 gnd.n4930 gnd.n4917 19.5087
R7888 gnd.n4928 gnd.n4919 19.5087
R7889 gnd.n1422 gnd.n1416 19.5087
R7890 gnd.n6285 gnd.t96 19.4385
R7891 gnd.n7273 gnd.t59 19.4385
R7892 gnd.n7449 gnd.t74 19.4385
R7893 gnd.n6154 gnd.n6153 19.3944
R7894 gnd.n6153 gnd.n6152 19.3944
R7895 gnd.n6152 gnd.n1191 19.3944
R7896 gnd.n6148 gnd.n1191 19.3944
R7897 gnd.n6148 gnd.n6147 19.3944
R7898 gnd.n6147 gnd.n6146 19.3944
R7899 gnd.n6146 gnd.n1196 19.3944
R7900 gnd.n6142 gnd.n1196 19.3944
R7901 gnd.n6142 gnd.n6141 19.3944
R7902 gnd.n6141 gnd.n6140 19.3944
R7903 gnd.n6140 gnd.n1201 19.3944
R7904 gnd.n6136 gnd.n1201 19.3944
R7905 gnd.n6136 gnd.n6135 19.3944
R7906 gnd.n6135 gnd.n6134 19.3944
R7907 gnd.n6134 gnd.n1206 19.3944
R7908 gnd.n6130 gnd.n1206 19.3944
R7909 gnd.n6130 gnd.n6129 19.3944
R7910 gnd.n6129 gnd.n6128 19.3944
R7911 gnd.n6128 gnd.n1211 19.3944
R7912 gnd.n6124 gnd.n1211 19.3944
R7913 gnd.n6124 gnd.n6123 19.3944
R7914 gnd.n6123 gnd.n6122 19.3944
R7915 gnd.n6122 gnd.n1216 19.3944
R7916 gnd.n6118 gnd.n1216 19.3944
R7917 gnd.n6118 gnd.n6117 19.3944
R7918 gnd.n6117 gnd.n6116 19.3944
R7919 gnd.n6116 gnd.n1221 19.3944
R7920 gnd.n6112 gnd.n1221 19.3944
R7921 gnd.n6112 gnd.n6111 19.3944
R7922 gnd.n6111 gnd.n6110 19.3944
R7923 gnd.n6110 gnd.n1226 19.3944
R7924 gnd.n6106 gnd.n1226 19.3944
R7925 gnd.n6106 gnd.n6105 19.3944
R7926 gnd.n6105 gnd.n6104 19.3944
R7927 gnd.n6104 gnd.n1231 19.3944
R7928 gnd.n6100 gnd.n1231 19.3944
R7929 gnd.n6100 gnd.n6099 19.3944
R7930 gnd.n6099 gnd.n6098 19.3944
R7931 gnd.n6098 gnd.n1236 19.3944
R7932 gnd.n6094 gnd.n1236 19.3944
R7933 gnd.n6094 gnd.n6093 19.3944
R7934 gnd.n6093 gnd.n6092 19.3944
R7935 gnd.n6092 gnd.n1241 19.3944
R7936 gnd.n6088 gnd.n1241 19.3944
R7937 gnd.n6088 gnd.n6087 19.3944
R7938 gnd.n6087 gnd.n6086 19.3944
R7939 gnd.n6086 gnd.n1246 19.3944
R7940 gnd.n6082 gnd.n1246 19.3944
R7941 gnd.n6082 gnd.n6081 19.3944
R7942 gnd.n6081 gnd.n6080 19.3944
R7943 gnd.n6080 gnd.n1251 19.3944
R7944 gnd.n6076 gnd.n1251 19.3944
R7945 gnd.n6076 gnd.n6075 19.3944
R7946 gnd.n6075 gnd.n6074 19.3944
R7947 gnd.n6074 gnd.n1256 19.3944
R7948 gnd.n6070 gnd.n1256 19.3944
R7949 gnd.n6070 gnd.n6069 19.3944
R7950 gnd.n6069 gnd.n6068 19.3944
R7951 gnd.n6068 gnd.n1261 19.3944
R7952 gnd.n6064 gnd.n1261 19.3944
R7953 gnd.n6064 gnd.n6063 19.3944
R7954 gnd.n6063 gnd.n6062 19.3944
R7955 gnd.n6062 gnd.n1266 19.3944
R7956 gnd.n6058 gnd.n1266 19.3944
R7957 gnd.n6058 gnd.n6057 19.3944
R7958 gnd.n6057 gnd.n6056 19.3944
R7959 gnd.n6056 gnd.n1271 19.3944
R7960 gnd.n6052 gnd.n1271 19.3944
R7961 gnd.n6052 gnd.n6051 19.3944
R7962 gnd.n6051 gnd.n6050 19.3944
R7963 gnd.n6050 gnd.n1276 19.3944
R7964 gnd.n6046 gnd.n1276 19.3944
R7965 gnd.n6046 gnd.n6045 19.3944
R7966 gnd.n6045 gnd.n6044 19.3944
R7967 gnd.n6044 gnd.n1281 19.3944
R7968 gnd.n6040 gnd.n1281 19.3944
R7969 gnd.n6040 gnd.n6039 19.3944
R7970 gnd.n6039 gnd.n6038 19.3944
R7971 gnd.n6038 gnd.n1286 19.3944
R7972 gnd.n6034 gnd.n1286 19.3944
R7973 gnd.n6034 gnd.n6033 19.3944
R7974 gnd.n6033 gnd.n6032 19.3944
R7975 gnd.n6032 gnd.n1291 19.3944
R7976 gnd.n6028 gnd.n1291 19.3944
R7977 gnd.n6028 gnd.n6027 19.3944
R7978 gnd.n6027 gnd.n6026 19.3944
R7979 gnd.n6026 gnd.n1296 19.3944
R7980 gnd.n6022 gnd.n1296 19.3944
R7981 gnd.n6022 gnd.n6021 19.3944
R7982 gnd.n6021 gnd.n6020 19.3944
R7983 gnd.n6020 gnd.n1301 19.3944
R7984 gnd.n6016 gnd.n1301 19.3944
R7985 gnd.n6016 gnd.n6015 19.3944
R7986 gnd.n6015 gnd.n6014 19.3944
R7987 gnd.n6014 gnd.n1306 19.3944
R7988 gnd.n6010 gnd.n1306 19.3944
R7989 gnd.n6010 gnd.n6009 19.3944
R7990 gnd.n6009 gnd.n6008 19.3944
R7991 gnd.n6008 gnd.n1311 19.3944
R7992 gnd.n6004 gnd.n1311 19.3944
R7993 gnd.n6004 gnd.n6003 19.3944
R7994 gnd.n6160 gnd.n6159 19.3944
R7995 gnd.n6159 gnd.n6158 19.3944
R7996 gnd.n6158 gnd.n1186 19.3944
R7997 gnd.n4768 gnd.n4767 19.3944
R7998 gnd.n4767 gnd.n4653 19.3944
R7999 gnd.n4760 gnd.n4653 19.3944
R8000 gnd.n4760 gnd.n4759 19.3944
R8001 gnd.n4759 gnd.n4673 19.3944
R8002 gnd.n4752 gnd.n4673 19.3944
R8003 gnd.n4752 gnd.n4751 19.3944
R8004 gnd.n4751 gnd.n4683 19.3944
R8005 gnd.n4744 gnd.n4683 19.3944
R8006 gnd.n4744 gnd.n4743 19.3944
R8007 gnd.n4743 gnd.n4696 19.3944
R8008 gnd.n4736 gnd.n4696 19.3944
R8009 gnd.n4736 gnd.n4735 19.3944
R8010 gnd.n4735 gnd.n4706 19.3944
R8011 gnd.n4728 gnd.n4706 19.3944
R8012 gnd.n4728 gnd.n4727 19.3944
R8013 gnd.n4727 gnd.n1170 19.3944
R8014 gnd.n6171 gnd.n1170 19.3944
R8015 gnd.n6171 gnd.n6170 19.3944
R8016 gnd.n6170 gnd.n6169 19.3944
R8017 gnd.n6169 gnd.n1174 19.3944
R8018 gnd.n6165 gnd.n1174 19.3944
R8019 gnd.n6165 gnd.n6164 19.3944
R8020 gnd.n6164 gnd.n6163 19.3944
R8021 gnd.n7175 gnd.n545 19.3944
R8022 gnd.n7175 gnd.n7174 19.3944
R8023 gnd.n7174 gnd.n7173 19.3944
R8024 gnd.n7173 gnd.n7171 19.3944
R8025 gnd.n7171 gnd.n7168 19.3944
R8026 gnd.n7168 gnd.n7167 19.3944
R8027 gnd.n7167 gnd.n7164 19.3944
R8028 gnd.n7164 gnd.n7163 19.3944
R8029 gnd.n7163 gnd.n7160 19.3944
R8030 gnd.n7160 gnd.n7159 19.3944
R8031 gnd.n7159 gnd.n7156 19.3944
R8032 gnd.n7156 gnd.n7155 19.3944
R8033 gnd.n7155 gnd.n7152 19.3944
R8034 gnd.n7152 gnd.n7151 19.3944
R8035 gnd.n7151 gnd.n7148 19.3944
R8036 gnd.n7146 gnd.n7143 19.3944
R8037 gnd.n7143 gnd.n7142 19.3944
R8038 gnd.n7142 gnd.n7139 19.3944
R8039 gnd.n7139 gnd.n7138 19.3944
R8040 gnd.n7138 gnd.n7135 19.3944
R8041 gnd.n7135 gnd.n7134 19.3944
R8042 gnd.n7134 gnd.n7131 19.3944
R8043 gnd.n7131 gnd.n7130 19.3944
R8044 gnd.n7130 gnd.n7127 19.3944
R8045 gnd.n7127 gnd.n7126 19.3944
R8046 gnd.n7126 gnd.n7123 19.3944
R8047 gnd.n7123 gnd.n7122 19.3944
R8048 gnd.n7122 gnd.n7119 19.3944
R8049 gnd.n7119 gnd.n7118 19.3944
R8050 gnd.n7118 gnd.n7115 19.3944
R8051 gnd.n7115 gnd.n7114 19.3944
R8052 gnd.n7114 gnd.n7111 19.3944
R8053 gnd.n7111 gnd.n7110 19.3944
R8054 gnd.n7103 gnd.n7102 19.3944
R8055 gnd.n7102 gnd.n7101 19.3944
R8056 gnd.n7101 gnd.n7100 19.3944
R8057 gnd.n7100 gnd.n593 19.3944
R8058 gnd.n5868 gnd.n593 19.3944
R8059 gnd.n5869 gnd.n5868 19.3944
R8060 gnd.n5872 gnd.n5869 19.3944
R8061 gnd.n5872 gnd.n5862 19.3944
R8062 gnd.n5915 gnd.n5862 19.3944
R8063 gnd.n5915 gnd.n5914 19.3944
R8064 gnd.n5914 gnd.n5913 19.3944
R8065 gnd.n5913 gnd.n5910 19.3944
R8066 gnd.n5910 gnd.n5909 19.3944
R8067 gnd.n5909 gnd.n5885 19.3944
R8068 gnd.n5885 gnd.n5884 19.3944
R8069 gnd.n5884 gnd.n613 19.3944
R8070 gnd.n6930 gnd.n613 19.3944
R8071 gnd.n6930 gnd.n611 19.3944
R8072 gnd.n7038 gnd.n611 19.3944
R8073 gnd.n7038 gnd.n7037 19.3944
R8074 gnd.n7037 gnd.n7036 19.3944
R8075 gnd.n7036 gnd.n7034 19.3944
R8076 gnd.n7034 gnd.n7033 19.3944
R8077 gnd.n7033 gnd.n7031 19.3944
R8078 gnd.n7031 gnd.n7030 19.3944
R8079 gnd.n7030 gnd.n7028 19.3944
R8080 gnd.n7028 gnd.n7027 19.3944
R8081 gnd.n7027 gnd.n7025 19.3944
R8082 gnd.n7025 gnd.n7024 19.3944
R8083 gnd.n7024 gnd.n7022 19.3944
R8084 gnd.n7022 gnd.n7021 19.3944
R8085 gnd.n7021 gnd.n7019 19.3944
R8086 gnd.n7019 gnd.n7018 19.3944
R8087 gnd.n7018 gnd.n7016 19.3944
R8088 gnd.n7016 gnd.n7015 19.3944
R8089 gnd.n7015 gnd.n7013 19.3944
R8090 gnd.n7013 gnd.n7012 19.3944
R8091 gnd.n7012 gnd.n7010 19.3944
R8092 gnd.n7010 gnd.n7009 19.3944
R8093 gnd.n7009 gnd.n7007 19.3944
R8094 gnd.n7007 gnd.n7006 19.3944
R8095 gnd.n7006 gnd.n7004 19.3944
R8096 gnd.n7004 gnd.n7003 19.3944
R8097 gnd.n7003 gnd.n7001 19.3944
R8098 gnd.n7001 gnd.n7000 19.3944
R8099 gnd.n7000 gnd.n6998 19.3944
R8100 gnd.n6998 gnd.n6997 19.3944
R8101 gnd.n6997 gnd.n6995 19.3944
R8102 gnd.n6995 gnd.n6994 19.3944
R8103 gnd.n6994 gnd.n6992 19.3944
R8104 gnd.n6992 gnd.n6991 19.3944
R8105 gnd.n6991 gnd.n6989 19.3944
R8106 gnd.n6989 gnd.n6988 19.3944
R8107 gnd.n6988 gnd.n6986 19.3944
R8108 gnd.n6986 gnd.n6985 19.3944
R8109 gnd.n6985 gnd.n6983 19.3944
R8110 gnd.n6983 gnd.n6982 19.3944
R8111 gnd.n6982 gnd.n6980 19.3944
R8112 gnd.n6980 gnd.n6979 19.3944
R8113 gnd.n6979 gnd.n6977 19.3944
R8114 gnd.n6977 gnd.n6976 19.3944
R8115 gnd.n6976 gnd.n204 19.3944
R8116 gnd.n7552 gnd.n204 19.3944
R8117 gnd.n7553 gnd.n7552 19.3944
R8118 gnd.n7591 gnd.n165 19.3944
R8119 gnd.n7586 gnd.n165 19.3944
R8120 gnd.n7586 gnd.n7585 19.3944
R8121 gnd.n7585 gnd.n7584 19.3944
R8122 gnd.n7584 gnd.n172 19.3944
R8123 gnd.n7579 gnd.n172 19.3944
R8124 gnd.n7579 gnd.n7578 19.3944
R8125 gnd.n7578 gnd.n7577 19.3944
R8126 gnd.n7577 gnd.n179 19.3944
R8127 gnd.n7572 gnd.n179 19.3944
R8128 gnd.n7572 gnd.n7571 19.3944
R8129 gnd.n7571 gnd.n7570 19.3944
R8130 gnd.n7570 gnd.n186 19.3944
R8131 gnd.n7565 gnd.n186 19.3944
R8132 gnd.n7565 gnd.n7564 19.3944
R8133 gnd.n7564 gnd.n7563 19.3944
R8134 gnd.n7563 gnd.n193 19.3944
R8135 gnd.n7558 gnd.n193 19.3944
R8136 gnd.n7624 gnd.n7623 19.3944
R8137 gnd.n7623 gnd.n7622 19.3944
R8138 gnd.n7622 gnd.n137 19.3944
R8139 gnd.n7617 gnd.n137 19.3944
R8140 gnd.n7617 gnd.n7616 19.3944
R8141 gnd.n7616 gnd.n7615 19.3944
R8142 gnd.n7615 gnd.n144 19.3944
R8143 gnd.n7610 gnd.n144 19.3944
R8144 gnd.n7610 gnd.n7609 19.3944
R8145 gnd.n7609 gnd.n7608 19.3944
R8146 gnd.n7608 gnd.n151 19.3944
R8147 gnd.n7603 gnd.n151 19.3944
R8148 gnd.n7603 gnd.n7602 19.3944
R8149 gnd.n7602 gnd.n7601 19.3944
R8150 gnd.n7601 gnd.n158 19.3944
R8151 gnd.n7596 gnd.n158 19.3944
R8152 gnd.n7596 gnd.n7595 19.3944
R8153 gnd.n7235 gnd.n452 19.3944
R8154 gnd.n7239 gnd.n452 19.3944
R8155 gnd.n7239 gnd.n437 19.3944
R8156 gnd.n7251 gnd.n437 19.3944
R8157 gnd.n7251 gnd.n435 19.3944
R8158 gnd.n7255 gnd.n435 19.3944
R8159 gnd.n7255 gnd.n419 19.3944
R8160 gnd.n7267 gnd.n419 19.3944
R8161 gnd.n7267 gnd.n417 19.3944
R8162 gnd.n7271 gnd.n417 19.3944
R8163 gnd.n7271 gnd.n403 19.3944
R8164 gnd.n7283 gnd.n403 19.3944
R8165 gnd.n7283 gnd.n401 19.3944
R8166 gnd.n7287 gnd.n401 19.3944
R8167 gnd.n7287 gnd.n385 19.3944
R8168 gnd.n7299 gnd.n385 19.3944
R8169 gnd.n7299 gnd.n383 19.3944
R8170 gnd.n7303 gnd.n383 19.3944
R8171 gnd.n7303 gnd.n369 19.3944
R8172 gnd.n7315 gnd.n369 19.3944
R8173 gnd.n7315 gnd.n367 19.3944
R8174 gnd.n7319 gnd.n367 19.3944
R8175 gnd.n7319 gnd.n351 19.3944
R8176 gnd.n7331 gnd.n351 19.3944
R8177 gnd.n7331 gnd.n349 19.3944
R8178 gnd.n7335 gnd.n349 19.3944
R8179 gnd.n7335 gnd.n336 19.3944
R8180 gnd.n7347 gnd.n336 19.3944
R8181 gnd.n7347 gnd.n334 19.3944
R8182 gnd.n7351 gnd.n334 19.3944
R8183 gnd.n7351 gnd.n318 19.3944
R8184 gnd.n7363 gnd.n318 19.3944
R8185 gnd.n7363 gnd.n316 19.3944
R8186 gnd.n7367 gnd.n316 19.3944
R8187 gnd.n7367 gnd.n304 19.3944
R8188 gnd.n7379 gnd.n304 19.3944
R8189 gnd.n7379 gnd.n302 19.3944
R8190 gnd.n7383 gnd.n302 19.3944
R8191 gnd.n7383 gnd.n288 19.3944
R8192 gnd.n7395 gnd.n288 19.3944
R8193 gnd.n7395 gnd.n286 19.3944
R8194 gnd.n7399 gnd.n286 19.3944
R8195 gnd.n7399 gnd.n274 19.3944
R8196 gnd.n7411 gnd.n274 19.3944
R8197 gnd.n7411 gnd.n272 19.3944
R8198 gnd.n7415 gnd.n272 19.3944
R8199 gnd.n7415 gnd.n258 19.3944
R8200 gnd.n7427 gnd.n258 19.3944
R8201 gnd.n7427 gnd.n256 19.3944
R8202 gnd.n7431 gnd.n256 19.3944
R8203 gnd.n7431 gnd.n243 19.3944
R8204 gnd.n7443 gnd.n243 19.3944
R8205 gnd.n7443 gnd.n241 19.3944
R8206 gnd.n7447 gnd.n241 19.3944
R8207 gnd.n7447 gnd.n227 19.3944
R8208 gnd.n7459 gnd.n227 19.3944
R8209 gnd.n7459 gnd.n225 19.3944
R8210 gnd.n7463 gnd.n225 19.3944
R8211 gnd.n7463 gnd.n211 19.3944
R8212 gnd.n7543 gnd.n211 19.3944
R8213 gnd.n7543 gnd.n209 19.3944
R8214 gnd.n7547 gnd.n209 19.3944
R8215 gnd.n7547 gnd.n132 19.3944
R8216 gnd.n7627 gnd.n132 19.3944
R8217 gnd.n5971 gnd.n5931 19.3944
R8218 gnd.n5971 gnd.n594 19.3944
R8219 gnd.n7096 gnd.n594 19.3944
R8220 gnd.n7096 gnd.n595 19.3944
R8221 gnd.n7092 gnd.n595 19.3944
R8222 gnd.n7092 gnd.n7091 19.3944
R8223 gnd.n7091 gnd.n7090 19.3944
R8224 gnd.n7090 gnd.n600 19.3944
R8225 gnd.n7086 gnd.n600 19.3944
R8226 gnd.n7086 gnd.n7085 19.3944
R8227 gnd.n7085 gnd.n7084 19.3944
R8228 gnd.n7084 gnd.n604 19.3944
R8229 gnd.n7080 gnd.n604 19.3944
R8230 gnd.n7080 gnd.n7079 19.3944
R8231 gnd.n7079 gnd.n7078 19.3944
R8232 gnd.n7078 gnd.n608 19.3944
R8233 gnd.n7074 gnd.n608 19.3944
R8234 gnd.n7074 gnd.n7073 19.3944
R8235 gnd.n7073 gnd.n7072 19.3944
R8236 gnd.n7072 gnd.n7042 19.3944
R8237 gnd.n7068 gnd.n7042 19.3944
R8238 gnd.n7068 gnd.n7067 19.3944
R8239 gnd.n7067 gnd.n7066 19.3944
R8240 gnd.n7066 gnd.n7046 19.3944
R8241 gnd.n7062 gnd.n7046 19.3944
R8242 gnd.n7062 gnd.n7061 19.3944
R8243 gnd.n7061 gnd.n7060 19.3944
R8244 gnd.n7060 gnd.n7050 19.3944
R8245 gnd.n7056 gnd.n7050 19.3944
R8246 gnd.n7056 gnd.n7055 19.3944
R8247 gnd.n7055 gnd.n7054 19.3944
R8248 gnd.n7054 gnd.n80 19.3944
R8249 gnd.n7680 gnd.n80 19.3944
R8250 gnd.n7680 gnd.n7679 19.3944
R8251 gnd.n7679 gnd.n7678 19.3944
R8252 gnd.n7678 gnd.n85 19.3944
R8253 gnd.n7674 gnd.n85 19.3944
R8254 gnd.n7674 gnd.n7673 19.3944
R8255 gnd.n7673 gnd.n7672 19.3944
R8256 gnd.n7672 gnd.n90 19.3944
R8257 gnd.n7668 gnd.n90 19.3944
R8258 gnd.n7668 gnd.n7667 19.3944
R8259 gnd.n7667 gnd.n7666 19.3944
R8260 gnd.n7666 gnd.n95 19.3944
R8261 gnd.n7662 gnd.n95 19.3944
R8262 gnd.n7662 gnd.n7661 19.3944
R8263 gnd.n7661 gnd.n7660 19.3944
R8264 gnd.n7660 gnd.n100 19.3944
R8265 gnd.n7656 gnd.n100 19.3944
R8266 gnd.n7656 gnd.n7655 19.3944
R8267 gnd.n7655 gnd.n7654 19.3944
R8268 gnd.n7654 gnd.n105 19.3944
R8269 gnd.n7650 gnd.n105 19.3944
R8270 gnd.n7650 gnd.n7649 19.3944
R8271 gnd.n7649 gnd.n7648 19.3944
R8272 gnd.n7648 gnd.n110 19.3944
R8273 gnd.n7644 gnd.n110 19.3944
R8274 gnd.n7644 gnd.n7643 19.3944
R8275 gnd.n7643 gnd.n7642 19.3944
R8276 gnd.n7642 gnd.n115 19.3944
R8277 gnd.n7638 gnd.n115 19.3944
R8278 gnd.n7638 gnd.n7637 19.3944
R8279 gnd.n7637 gnd.n7636 19.3944
R8280 gnd.n7636 gnd.n120 19.3944
R8281 gnd.n7530 gnd.n7529 19.3944
R8282 gnd.n7529 gnd.n7528 19.3944
R8283 gnd.n7528 gnd.n7477 19.3944
R8284 gnd.n7524 gnd.n7477 19.3944
R8285 gnd.n7524 gnd.n7523 19.3944
R8286 gnd.n7523 gnd.n7522 19.3944
R8287 gnd.n7522 gnd.n7485 19.3944
R8288 gnd.n7518 gnd.n7485 19.3944
R8289 gnd.n7518 gnd.n7517 19.3944
R8290 gnd.n7517 gnd.n7516 19.3944
R8291 gnd.n7516 gnd.n7493 19.3944
R8292 gnd.n7512 gnd.n7493 19.3944
R8293 gnd.n7512 gnd.n7511 19.3944
R8294 gnd.n7511 gnd.n7510 19.3944
R8295 gnd.n7510 gnd.n7501 19.3944
R8296 gnd.n7506 gnd.n7501 19.3944
R8297 gnd.n7228 gnd.n7227 19.3944
R8298 gnd.n7227 gnd.n462 19.3944
R8299 gnd.n7220 gnd.n462 19.3944
R8300 gnd.n7220 gnd.n7219 19.3944
R8301 gnd.n7219 gnd.n470 19.3944
R8302 gnd.n7212 gnd.n470 19.3944
R8303 gnd.n7212 gnd.n7211 19.3944
R8304 gnd.n7211 gnd.n478 19.3944
R8305 gnd.n7204 gnd.n478 19.3944
R8306 gnd.n7204 gnd.n7203 19.3944
R8307 gnd.n7203 gnd.n486 19.3944
R8308 gnd.n7196 gnd.n486 19.3944
R8309 gnd.n7196 gnd.n7195 19.3944
R8310 gnd.n7195 gnd.n494 19.3944
R8311 gnd.n7188 gnd.n494 19.3944
R8312 gnd.n7188 gnd.n7187 19.3944
R8313 gnd.n7231 gnd.n446 19.3944
R8314 gnd.n7243 gnd.n446 19.3944
R8315 gnd.n7243 gnd.n444 19.3944
R8316 gnd.n7247 gnd.n444 19.3944
R8317 gnd.n7247 gnd.n428 19.3944
R8318 gnd.n7259 gnd.n428 19.3944
R8319 gnd.n7259 gnd.n426 19.3944
R8320 gnd.n7263 gnd.n426 19.3944
R8321 gnd.n7263 gnd.n411 19.3944
R8322 gnd.n7275 gnd.n411 19.3944
R8323 gnd.n7275 gnd.n409 19.3944
R8324 gnd.n7279 gnd.n409 19.3944
R8325 gnd.n7279 gnd.n394 19.3944
R8326 gnd.n7291 gnd.n394 19.3944
R8327 gnd.n7291 gnd.n392 19.3944
R8328 gnd.n7295 gnd.n392 19.3944
R8329 gnd.n7295 gnd.n377 19.3944
R8330 gnd.n7307 gnd.n377 19.3944
R8331 gnd.n7307 gnd.n375 19.3944
R8332 gnd.n7311 gnd.n375 19.3944
R8333 gnd.n7311 gnd.n360 19.3944
R8334 gnd.n7323 gnd.n360 19.3944
R8335 gnd.n7323 gnd.n358 19.3944
R8336 gnd.n7327 gnd.n358 19.3944
R8337 gnd.n7327 gnd.n344 19.3944
R8338 gnd.n7339 gnd.n344 19.3944
R8339 gnd.n7339 gnd.n342 19.3944
R8340 gnd.n7343 gnd.n342 19.3944
R8341 gnd.n7343 gnd.n328 19.3944
R8342 gnd.n7355 gnd.n328 19.3944
R8343 gnd.n7355 gnd.n325 19.3944
R8344 gnd.n7359 gnd.n325 19.3944
R8345 gnd.n7359 gnd.n311 19.3944
R8346 gnd.n7371 gnd.n311 19.3944
R8347 gnd.n7371 gnd.n309 19.3944
R8348 gnd.n7375 gnd.n309 19.3944
R8349 gnd.n7375 gnd.n297 19.3944
R8350 gnd.n7387 gnd.n297 19.3944
R8351 gnd.n7387 gnd.n295 19.3944
R8352 gnd.n7391 gnd.n295 19.3944
R8353 gnd.n7391 gnd.n281 19.3944
R8354 gnd.n7403 gnd.n281 19.3944
R8355 gnd.n7403 gnd.n279 19.3944
R8356 gnd.n7407 gnd.n279 19.3944
R8357 gnd.n7407 gnd.n267 19.3944
R8358 gnd.n7419 gnd.n267 19.3944
R8359 gnd.n7419 gnd.n265 19.3944
R8360 gnd.n7423 gnd.n265 19.3944
R8361 gnd.n7423 gnd.n250 19.3944
R8362 gnd.n7435 gnd.n250 19.3944
R8363 gnd.n7435 gnd.n248 19.3944
R8364 gnd.n7439 gnd.n248 19.3944
R8365 gnd.n7439 gnd.n236 19.3944
R8366 gnd.n7451 gnd.n236 19.3944
R8367 gnd.n7451 gnd.n234 19.3944
R8368 gnd.n7455 gnd.n234 19.3944
R8369 gnd.n7455 gnd.n221 19.3944
R8370 gnd.n7467 gnd.n221 19.3944
R8371 gnd.n7467 gnd.n218 19.3944
R8372 gnd.n7539 gnd.n218 19.3944
R8373 gnd.n7539 gnd.n219 19.3944
R8374 gnd.n7535 gnd.n219 19.3944
R8375 gnd.n7535 gnd.n7534 19.3944
R8376 gnd.n7534 gnd.n7533 19.3944
R8377 gnd.n4661 gnd.n4657 19.3944
R8378 gnd.n4661 gnd.n4656 19.3944
R8379 gnd.n4764 gnd.n4656 19.3944
R8380 gnd.n4764 gnd.n4763 19.3944
R8381 gnd.n4763 gnd.n4668 19.3944
R8382 gnd.n4756 gnd.n4668 19.3944
R8383 gnd.n4756 gnd.n4755 19.3944
R8384 gnd.n4755 gnd.n4679 19.3944
R8385 gnd.n4748 gnd.n4679 19.3944
R8386 gnd.n4748 gnd.n4747 19.3944
R8387 gnd.n4747 gnd.n4690 19.3944
R8388 gnd.n4740 gnd.n4690 19.3944
R8389 gnd.n4740 gnd.n4739 19.3944
R8390 gnd.n4739 gnd.n4702 19.3944
R8391 gnd.n4732 gnd.n4702 19.3944
R8392 gnd.n4732 gnd.n4731 19.3944
R8393 gnd.n4540 gnd.n4539 19.3944
R8394 gnd.n4543 gnd.n4540 19.3944
R8395 gnd.n4543 gnd.n1943 19.3944
R8396 gnd.n4547 gnd.n1943 19.3944
R8397 gnd.n4547 gnd.n1941 19.3944
R8398 gnd.n4551 gnd.n1941 19.3944
R8399 gnd.n4551 gnd.n1939 19.3944
R8400 gnd.n4560 gnd.n1939 19.3944
R8401 gnd.n4560 gnd.n4559 19.3944
R8402 gnd.n4559 gnd.n4558 19.3944
R8403 gnd.n4558 gnd.n1918 19.3944
R8404 gnd.n1918 gnd.n1916 19.3944
R8405 gnd.n4611 gnd.n1916 19.3944
R8406 gnd.n4611 gnd.n1914 19.3944
R8407 gnd.n4615 gnd.n1914 19.3944
R8408 gnd.n4615 gnd.n1912 19.3944
R8409 gnd.n4619 gnd.n1912 19.3944
R8410 gnd.n4619 gnd.n1910 19.3944
R8411 gnd.n4623 gnd.n1910 19.3944
R8412 gnd.n4623 gnd.n1908 19.3944
R8413 gnd.n4627 gnd.n1908 19.3944
R8414 gnd.n4627 gnd.n1906 19.3944
R8415 gnd.n4631 gnd.n1906 19.3944
R8416 gnd.n4631 gnd.n1902 19.3944
R8417 gnd.n4775 gnd.n1902 19.3944
R8418 gnd.n4775 gnd.n1900 19.3944
R8419 gnd.n4779 gnd.n1900 19.3944
R8420 gnd.n4779 gnd.n1888 19.3944
R8421 gnd.n4794 gnd.n1888 19.3944
R8422 gnd.n4794 gnd.n1886 19.3944
R8423 gnd.n4798 gnd.n1886 19.3944
R8424 gnd.n4798 gnd.n1874 19.3944
R8425 gnd.n4813 gnd.n1874 19.3944
R8426 gnd.n4813 gnd.n1872 19.3944
R8427 gnd.n4817 gnd.n1872 19.3944
R8428 gnd.n4817 gnd.n1860 19.3944
R8429 gnd.n4832 gnd.n1860 19.3944
R8430 gnd.n4832 gnd.n1858 19.3944
R8431 gnd.n4836 gnd.n1858 19.3944
R8432 gnd.n4836 gnd.n1846 19.3944
R8433 gnd.n4851 gnd.n1846 19.3944
R8434 gnd.n4851 gnd.n1844 19.3944
R8435 gnd.n4855 gnd.n1844 19.3944
R8436 gnd.n4855 gnd.n1831 19.3944
R8437 gnd.n4870 gnd.n1831 19.3944
R8438 gnd.n4870 gnd.n1829 19.3944
R8439 gnd.n4876 gnd.n1829 19.3944
R8440 gnd.n4876 gnd.n4875 19.3944
R8441 gnd.n4875 gnd.n1818 19.3944
R8442 gnd.n5091 gnd.n1818 19.3944
R8443 gnd.n5091 gnd.n1816 19.3944
R8444 gnd.n5095 gnd.n1816 19.3944
R8445 gnd.n5095 gnd.n1744 19.3944
R8446 gnd.n5132 gnd.n1744 19.3944
R8447 gnd.n5132 gnd.n1742 19.3944
R8448 gnd.n5138 gnd.n1742 19.3944
R8449 gnd.n5138 gnd.n5137 19.3944
R8450 gnd.n5137 gnd.n1717 19.3944
R8451 gnd.n5168 gnd.n1717 19.3944
R8452 gnd.n5168 gnd.n1715 19.3944
R8453 gnd.n5172 gnd.n1715 19.3944
R8454 gnd.n5172 gnd.n1695 19.3944
R8455 gnd.n5196 gnd.n1695 19.3944
R8456 gnd.n5196 gnd.n1693 19.3944
R8457 gnd.n5202 gnd.n1693 19.3944
R8458 gnd.n5202 gnd.n5201 19.3944
R8459 gnd.n5201 gnd.n1663 19.3944
R8460 gnd.n5233 gnd.n1663 19.3944
R8461 gnd.n5233 gnd.n1661 19.3944
R8462 gnd.n5248 gnd.n1661 19.3944
R8463 gnd.n5248 gnd.n5247 19.3944
R8464 gnd.n5247 gnd.n5246 19.3944
R8465 gnd.n5246 gnd.n5239 19.3944
R8466 gnd.n5242 gnd.n5239 19.3944
R8467 gnd.n5242 gnd.n1622 19.3944
R8468 gnd.n5327 gnd.n1622 19.3944
R8469 gnd.n5327 gnd.n1620 19.3944
R8470 gnd.n5331 gnd.n1620 19.3944
R8471 gnd.n5331 gnd.n1604 19.3944
R8472 gnd.n5370 gnd.n1604 19.3944
R8473 gnd.n5370 gnd.n1602 19.3944
R8474 gnd.n5374 gnd.n1602 19.3944
R8475 gnd.n5374 gnd.n1580 19.3944
R8476 gnd.n5404 gnd.n1580 19.3944
R8477 gnd.n5404 gnd.n1578 19.3944
R8478 gnd.n5408 gnd.n1578 19.3944
R8479 gnd.n5408 gnd.n1557 19.3944
R8480 gnd.n5445 gnd.n1557 19.3944
R8481 gnd.n5445 gnd.n1555 19.3944
R8482 gnd.n5449 gnd.n1555 19.3944
R8483 gnd.n5449 gnd.n1536 19.3944
R8484 gnd.n5492 gnd.n1536 19.3944
R8485 gnd.n5492 gnd.n1534 19.3944
R8486 gnd.n5496 gnd.n1534 19.3944
R8487 gnd.n5496 gnd.n1509 19.3944
R8488 gnd.n5524 gnd.n1509 19.3944
R8489 gnd.n5524 gnd.n1507 19.3944
R8490 gnd.n5528 gnd.n1507 19.3944
R8491 gnd.n5528 gnd.n1487 19.3944
R8492 gnd.n5570 gnd.n1487 19.3944
R8493 gnd.n5570 gnd.n1485 19.3944
R8494 gnd.n5574 gnd.n1485 19.3944
R8495 gnd.n5574 gnd.n1400 19.3944
R8496 gnd.n5718 gnd.n1400 19.3944
R8497 gnd.n5718 gnd.n1398 19.3944
R8498 gnd.n5722 gnd.n1398 19.3944
R8499 gnd.n5722 gnd.n1385 19.3944
R8500 gnd.n5737 gnd.n1385 19.3944
R8501 gnd.n5737 gnd.n1383 19.3944
R8502 gnd.n5741 gnd.n1383 19.3944
R8503 gnd.n5741 gnd.n1371 19.3944
R8504 gnd.n5756 gnd.n1371 19.3944
R8505 gnd.n5756 gnd.n1369 19.3944
R8506 gnd.n5760 gnd.n1369 19.3944
R8507 gnd.n5760 gnd.n1357 19.3944
R8508 gnd.n5775 gnd.n1357 19.3944
R8509 gnd.n5775 gnd.n1355 19.3944
R8510 gnd.n5779 gnd.n1355 19.3944
R8511 gnd.n5779 gnd.n1343 19.3944
R8512 gnd.n5794 gnd.n1343 19.3944
R8513 gnd.n5794 gnd.n1341 19.3944
R8514 gnd.n5798 gnd.n1341 19.3944
R8515 gnd.n5798 gnd.n1329 19.3944
R8516 gnd.n5813 gnd.n1329 19.3944
R8517 gnd.n5813 gnd.n1327 19.3944
R8518 gnd.n5990 gnd.n1327 19.3944
R8519 gnd.n5990 gnd.n5989 19.3944
R8520 gnd.n5989 gnd.n5988 19.3944
R8521 gnd.n5988 gnd.n5819 19.3944
R8522 gnd.n5841 gnd.n5819 19.3944
R8523 gnd.n5980 gnd.n5841 19.3944
R8524 gnd.n5980 gnd.n5979 19.3944
R8525 gnd.n5979 gnd.n5978 19.3944
R8526 gnd.n5978 gnd.n5847 19.3944
R8527 gnd.n5930 gnd.n5847 19.3944
R8528 gnd.n5930 gnd.n5929 19.3944
R8529 gnd.n5929 gnd.n5928 19.3944
R8530 gnd.n5928 gnd.n5853 19.3944
R8531 gnd.n5924 gnd.n5853 19.3944
R8532 gnd.n5924 gnd.n5923 19.3944
R8533 gnd.n5923 gnd.n5922 19.3944
R8534 gnd.n5922 gnd.n5859 19.3944
R8535 gnd.n5861 gnd.n5859 19.3944
R8536 gnd.n5891 gnd.n5861 19.3944
R8537 gnd.n5891 gnd.n5888 19.3944
R8538 gnd.n5904 gnd.n5888 19.3944
R8539 gnd.n5904 gnd.n5903 19.3944
R8540 gnd.n5903 gnd.n5902 19.3944
R8541 gnd.n5902 gnd.n5899 19.3944
R8542 gnd.n5899 gnd.n616 19.3944
R8543 gnd.n6925 gnd.n616 19.3944
R8544 gnd.n6925 gnd.n6924 19.3944
R8545 gnd.n6924 gnd.n6923 19.3944
R8546 gnd.n6923 gnd.n620 19.3944
R8547 gnd.n6706 gnd.n744 19.3944
R8548 gnd.n6712 gnd.n744 19.3944
R8549 gnd.n6712 gnd.n742 19.3944
R8550 gnd.n6716 gnd.n742 19.3944
R8551 gnd.n6716 gnd.n738 19.3944
R8552 gnd.n6722 gnd.n738 19.3944
R8553 gnd.n6722 gnd.n736 19.3944
R8554 gnd.n6726 gnd.n736 19.3944
R8555 gnd.n6726 gnd.n732 19.3944
R8556 gnd.n6732 gnd.n732 19.3944
R8557 gnd.n6732 gnd.n730 19.3944
R8558 gnd.n6736 gnd.n730 19.3944
R8559 gnd.n6736 gnd.n726 19.3944
R8560 gnd.n6742 gnd.n726 19.3944
R8561 gnd.n6742 gnd.n724 19.3944
R8562 gnd.n6746 gnd.n724 19.3944
R8563 gnd.n6746 gnd.n720 19.3944
R8564 gnd.n6752 gnd.n720 19.3944
R8565 gnd.n6752 gnd.n718 19.3944
R8566 gnd.n6756 gnd.n718 19.3944
R8567 gnd.n6756 gnd.n714 19.3944
R8568 gnd.n6762 gnd.n714 19.3944
R8569 gnd.n6762 gnd.n712 19.3944
R8570 gnd.n6766 gnd.n712 19.3944
R8571 gnd.n6766 gnd.n708 19.3944
R8572 gnd.n6772 gnd.n708 19.3944
R8573 gnd.n6772 gnd.n706 19.3944
R8574 gnd.n6776 gnd.n706 19.3944
R8575 gnd.n6776 gnd.n702 19.3944
R8576 gnd.n6782 gnd.n702 19.3944
R8577 gnd.n6782 gnd.n700 19.3944
R8578 gnd.n6786 gnd.n700 19.3944
R8579 gnd.n6786 gnd.n696 19.3944
R8580 gnd.n6792 gnd.n696 19.3944
R8581 gnd.n6792 gnd.n694 19.3944
R8582 gnd.n6796 gnd.n694 19.3944
R8583 gnd.n6796 gnd.n690 19.3944
R8584 gnd.n6802 gnd.n690 19.3944
R8585 gnd.n6802 gnd.n688 19.3944
R8586 gnd.n6806 gnd.n688 19.3944
R8587 gnd.n6806 gnd.n684 19.3944
R8588 gnd.n6812 gnd.n684 19.3944
R8589 gnd.n6812 gnd.n682 19.3944
R8590 gnd.n6816 gnd.n682 19.3944
R8591 gnd.n6816 gnd.n678 19.3944
R8592 gnd.n6822 gnd.n678 19.3944
R8593 gnd.n6822 gnd.n676 19.3944
R8594 gnd.n6826 gnd.n676 19.3944
R8595 gnd.n6826 gnd.n672 19.3944
R8596 gnd.n6832 gnd.n672 19.3944
R8597 gnd.n6832 gnd.n670 19.3944
R8598 gnd.n6836 gnd.n670 19.3944
R8599 gnd.n6836 gnd.n666 19.3944
R8600 gnd.n6842 gnd.n666 19.3944
R8601 gnd.n6842 gnd.n664 19.3944
R8602 gnd.n6846 gnd.n664 19.3944
R8603 gnd.n6846 gnd.n660 19.3944
R8604 gnd.n6852 gnd.n660 19.3944
R8605 gnd.n6852 gnd.n658 19.3944
R8606 gnd.n6856 gnd.n658 19.3944
R8607 gnd.n6856 gnd.n654 19.3944
R8608 gnd.n6862 gnd.n654 19.3944
R8609 gnd.n6862 gnd.n652 19.3944
R8610 gnd.n6866 gnd.n652 19.3944
R8611 gnd.n6866 gnd.n648 19.3944
R8612 gnd.n6872 gnd.n648 19.3944
R8613 gnd.n6872 gnd.n646 19.3944
R8614 gnd.n6876 gnd.n646 19.3944
R8615 gnd.n6876 gnd.n642 19.3944
R8616 gnd.n6882 gnd.n642 19.3944
R8617 gnd.n6882 gnd.n640 19.3944
R8618 gnd.n6886 gnd.n640 19.3944
R8619 gnd.n6886 gnd.n636 19.3944
R8620 gnd.n6892 gnd.n636 19.3944
R8621 gnd.n6892 gnd.n634 19.3944
R8622 gnd.n6896 gnd.n634 19.3944
R8623 gnd.n6896 gnd.n630 19.3944
R8624 gnd.n6902 gnd.n630 19.3944
R8625 gnd.n6902 gnd.n628 19.3944
R8626 gnd.n6906 gnd.n628 19.3944
R8627 gnd.n6906 gnd.n624 19.3944
R8628 gnd.n6913 gnd.n624 19.3944
R8629 gnd.n6913 gnd.n622 19.3944
R8630 gnd.n6918 gnd.n622 19.3944
R8631 gnd.n6321 gnd.n977 19.3944
R8632 gnd.n6321 gnd.n975 19.3944
R8633 gnd.n6325 gnd.n975 19.3944
R8634 gnd.n6325 gnd.n971 19.3944
R8635 gnd.n6331 gnd.n971 19.3944
R8636 gnd.n6331 gnd.n969 19.3944
R8637 gnd.n6335 gnd.n969 19.3944
R8638 gnd.n6335 gnd.n965 19.3944
R8639 gnd.n6341 gnd.n965 19.3944
R8640 gnd.n6341 gnd.n963 19.3944
R8641 gnd.n6345 gnd.n963 19.3944
R8642 gnd.n6345 gnd.n959 19.3944
R8643 gnd.n6351 gnd.n959 19.3944
R8644 gnd.n6351 gnd.n957 19.3944
R8645 gnd.n6355 gnd.n957 19.3944
R8646 gnd.n6355 gnd.n953 19.3944
R8647 gnd.n6361 gnd.n953 19.3944
R8648 gnd.n6361 gnd.n951 19.3944
R8649 gnd.n6365 gnd.n951 19.3944
R8650 gnd.n6365 gnd.n947 19.3944
R8651 gnd.n6371 gnd.n947 19.3944
R8652 gnd.n6371 gnd.n945 19.3944
R8653 gnd.n6375 gnd.n945 19.3944
R8654 gnd.n6375 gnd.n941 19.3944
R8655 gnd.n6381 gnd.n941 19.3944
R8656 gnd.n6381 gnd.n939 19.3944
R8657 gnd.n6385 gnd.n939 19.3944
R8658 gnd.n6385 gnd.n935 19.3944
R8659 gnd.n6391 gnd.n935 19.3944
R8660 gnd.n6391 gnd.n933 19.3944
R8661 gnd.n6395 gnd.n933 19.3944
R8662 gnd.n6395 gnd.n929 19.3944
R8663 gnd.n6401 gnd.n929 19.3944
R8664 gnd.n6401 gnd.n927 19.3944
R8665 gnd.n6405 gnd.n927 19.3944
R8666 gnd.n6405 gnd.n923 19.3944
R8667 gnd.n6411 gnd.n923 19.3944
R8668 gnd.n6411 gnd.n921 19.3944
R8669 gnd.n6415 gnd.n921 19.3944
R8670 gnd.n6415 gnd.n917 19.3944
R8671 gnd.n6421 gnd.n917 19.3944
R8672 gnd.n6421 gnd.n915 19.3944
R8673 gnd.n6425 gnd.n915 19.3944
R8674 gnd.n6425 gnd.n911 19.3944
R8675 gnd.n6431 gnd.n911 19.3944
R8676 gnd.n6431 gnd.n909 19.3944
R8677 gnd.n6435 gnd.n909 19.3944
R8678 gnd.n6435 gnd.n905 19.3944
R8679 gnd.n6441 gnd.n905 19.3944
R8680 gnd.n6441 gnd.n903 19.3944
R8681 gnd.n6445 gnd.n903 19.3944
R8682 gnd.n6445 gnd.n899 19.3944
R8683 gnd.n6451 gnd.n899 19.3944
R8684 gnd.n6451 gnd.n897 19.3944
R8685 gnd.n6455 gnd.n897 19.3944
R8686 gnd.n6455 gnd.n893 19.3944
R8687 gnd.n6461 gnd.n893 19.3944
R8688 gnd.n6461 gnd.n891 19.3944
R8689 gnd.n6465 gnd.n891 19.3944
R8690 gnd.n6465 gnd.n887 19.3944
R8691 gnd.n6471 gnd.n887 19.3944
R8692 gnd.n6471 gnd.n885 19.3944
R8693 gnd.n6475 gnd.n885 19.3944
R8694 gnd.n6475 gnd.n881 19.3944
R8695 gnd.n6481 gnd.n881 19.3944
R8696 gnd.n6481 gnd.n879 19.3944
R8697 gnd.n6485 gnd.n879 19.3944
R8698 gnd.n6485 gnd.n875 19.3944
R8699 gnd.n6491 gnd.n875 19.3944
R8700 gnd.n6491 gnd.n873 19.3944
R8701 gnd.n6495 gnd.n873 19.3944
R8702 gnd.n6495 gnd.n869 19.3944
R8703 gnd.n6501 gnd.n869 19.3944
R8704 gnd.n6501 gnd.n867 19.3944
R8705 gnd.n6505 gnd.n867 19.3944
R8706 gnd.n6505 gnd.n863 19.3944
R8707 gnd.n6511 gnd.n863 19.3944
R8708 gnd.n6511 gnd.n861 19.3944
R8709 gnd.n6515 gnd.n861 19.3944
R8710 gnd.n6515 gnd.n857 19.3944
R8711 gnd.n6521 gnd.n857 19.3944
R8712 gnd.n6521 gnd.n855 19.3944
R8713 gnd.n6525 gnd.n855 19.3944
R8714 gnd.n6525 gnd.n851 19.3944
R8715 gnd.n6531 gnd.n851 19.3944
R8716 gnd.n6531 gnd.n849 19.3944
R8717 gnd.n6535 gnd.n849 19.3944
R8718 gnd.n6535 gnd.n845 19.3944
R8719 gnd.n6541 gnd.n845 19.3944
R8720 gnd.n6541 gnd.n843 19.3944
R8721 gnd.n6545 gnd.n843 19.3944
R8722 gnd.n6545 gnd.n839 19.3944
R8723 gnd.n6551 gnd.n839 19.3944
R8724 gnd.n6551 gnd.n837 19.3944
R8725 gnd.n6555 gnd.n837 19.3944
R8726 gnd.n6555 gnd.n833 19.3944
R8727 gnd.n6561 gnd.n833 19.3944
R8728 gnd.n6561 gnd.n831 19.3944
R8729 gnd.n6565 gnd.n831 19.3944
R8730 gnd.n6565 gnd.n827 19.3944
R8731 gnd.n6571 gnd.n827 19.3944
R8732 gnd.n6571 gnd.n825 19.3944
R8733 gnd.n6575 gnd.n825 19.3944
R8734 gnd.n6575 gnd.n821 19.3944
R8735 gnd.n6581 gnd.n821 19.3944
R8736 gnd.n6581 gnd.n819 19.3944
R8737 gnd.n6585 gnd.n819 19.3944
R8738 gnd.n6585 gnd.n815 19.3944
R8739 gnd.n6591 gnd.n815 19.3944
R8740 gnd.n6591 gnd.n813 19.3944
R8741 gnd.n6595 gnd.n813 19.3944
R8742 gnd.n6595 gnd.n809 19.3944
R8743 gnd.n6601 gnd.n809 19.3944
R8744 gnd.n6601 gnd.n807 19.3944
R8745 gnd.n6605 gnd.n807 19.3944
R8746 gnd.n6605 gnd.n803 19.3944
R8747 gnd.n6611 gnd.n803 19.3944
R8748 gnd.n6611 gnd.n801 19.3944
R8749 gnd.n6615 gnd.n801 19.3944
R8750 gnd.n6615 gnd.n797 19.3944
R8751 gnd.n6621 gnd.n797 19.3944
R8752 gnd.n6621 gnd.n795 19.3944
R8753 gnd.n6625 gnd.n795 19.3944
R8754 gnd.n6625 gnd.n791 19.3944
R8755 gnd.n6631 gnd.n791 19.3944
R8756 gnd.n6631 gnd.n789 19.3944
R8757 gnd.n6635 gnd.n789 19.3944
R8758 gnd.n6635 gnd.n785 19.3944
R8759 gnd.n6641 gnd.n785 19.3944
R8760 gnd.n6641 gnd.n783 19.3944
R8761 gnd.n6645 gnd.n783 19.3944
R8762 gnd.n6645 gnd.n779 19.3944
R8763 gnd.n6651 gnd.n779 19.3944
R8764 gnd.n6651 gnd.n777 19.3944
R8765 gnd.n6655 gnd.n777 19.3944
R8766 gnd.n6655 gnd.n773 19.3944
R8767 gnd.n6661 gnd.n773 19.3944
R8768 gnd.n6661 gnd.n771 19.3944
R8769 gnd.n6665 gnd.n771 19.3944
R8770 gnd.n6665 gnd.n767 19.3944
R8771 gnd.n6671 gnd.n767 19.3944
R8772 gnd.n6671 gnd.n765 19.3944
R8773 gnd.n6675 gnd.n765 19.3944
R8774 gnd.n6675 gnd.n761 19.3944
R8775 gnd.n6681 gnd.n761 19.3944
R8776 gnd.n6681 gnd.n759 19.3944
R8777 gnd.n6685 gnd.n759 19.3944
R8778 gnd.n6685 gnd.n755 19.3944
R8779 gnd.n6691 gnd.n755 19.3944
R8780 gnd.n6691 gnd.n753 19.3944
R8781 gnd.n6696 gnd.n753 19.3944
R8782 gnd.n6696 gnd.n749 19.3944
R8783 gnd.n6702 gnd.n749 19.3944
R8784 gnd.n6703 gnd.n6702 19.3944
R8785 gnd.n4530 gnd.n4529 19.3944
R8786 gnd.n4529 gnd.n4528 19.3944
R8787 gnd.n4528 gnd.n4527 19.3944
R8788 gnd.n4527 gnd.n4525 19.3944
R8789 gnd.n4525 gnd.n4522 19.3944
R8790 gnd.n4522 gnd.n4521 19.3944
R8791 gnd.n4521 gnd.n4518 19.3944
R8792 gnd.n4518 gnd.n4517 19.3944
R8793 gnd.n4517 gnd.n4514 19.3944
R8794 gnd.n4514 gnd.n4513 19.3944
R8795 gnd.n4513 gnd.n4510 19.3944
R8796 gnd.n4510 gnd.n4509 19.3944
R8797 gnd.n4509 gnd.n4506 19.3944
R8798 gnd.n4506 gnd.n4505 19.3944
R8799 gnd.n4505 gnd.n4502 19.3944
R8800 gnd.n4502 gnd.n4501 19.3944
R8801 gnd.n4501 gnd.n4498 19.3944
R8802 gnd.n4498 gnd.n4497 19.3944
R8803 gnd.n4497 gnd.n4494 19.3944
R8804 gnd.n4494 gnd.n4493 19.3944
R8805 gnd.n4493 gnd.n4490 19.3944
R8806 gnd.n4490 gnd.n4489 19.3944
R8807 gnd.n4489 gnd.n4486 19.3944
R8808 gnd.n4486 gnd.n4485 19.3944
R8809 gnd.n4485 gnd.n4482 19.3944
R8810 gnd.n4482 gnd.n4481 19.3944
R8811 gnd.n4481 gnd.n4478 19.3944
R8812 gnd.n4478 gnd.n4477 19.3944
R8813 gnd.n4477 gnd.n4474 19.3944
R8814 gnd.n4474 gnd.n4473 19.3944
R8815 gnd.n4473 gnd.n4470 19.3944
R8816 gnd.n4470 gnd.n4469 19.3944
R8817 gnd.n4469 gnd.n4466 19.3944
R8818 gnd.n4466 gnd.n4465 19.3944
R8819 gnd.n4465 gnd.n4462 19.3944
R8820 gnd.n4462 gnd.n4461 19.3944
R8821 gnd.n4461 gnd.n4458 19.3944
R8822 gnd.n4458 gnd.n4457 19.3944
R8823 gnd.n4457 gnd.n4454 19.3944
R8824 gnd.n4454 gnd.n4453 19.3944
R8825 gnd.n4453 gnd.n4450 19.3944
R8826 gnd.n4450 gnd.n4449 19.3944
R8827 gnd.n4449 gnd.n4446 19.3944
R8828 gnd.n4446 gnd.n4445 19.3944
R8829 gnd.n4445 gnd.n4442 19.3944
R8830 gnd.n4442 gnd.n4441 19.3944
R8831 gnd.n4441 gnd.n4438 19.3944
R8832 gnd.n4438 gnd.n4437 19.3944
R8833 gnd.n4437 gnd.n4434 19.3944
R8834 gnd.n4434 gnd.n4433 19.3944
R8835 gnd.n4433 gnd.n4430 19.3944
R8836 gnd.n4430 gnd.n4429 19.3944
R8837 gnd.n4429 gnd.n4426 19.3944
R8838 gnd.n4426 gnd.n4425 19.3944
R8839 gnd.n4425 gnd.n4422 19.3944
R8840 gnd.n4422 gnd.n4421 19.3944
R8841 gnd.n4421 gnd.n4418 19.3944
R8842 gnd.n4418 gnd.n4417 19.3944
R8843 gnd.n4417 gnd.n4414 19.3944
R8844 gnd.n4414 gnd.n4413 19.3944
R8845 gnd.n4413 gnd.n4410 19.3944
R8846 gnd.n4410 gnd.n4409 19.3944
R8847 gnd.n4409 gnd.n4406 19.3944
R8848 gnd.n4406 gnd.n4405 19.3944
R8849 gnd.n4405 gnd.n4402 19.3944
R8850 gnd.n4402 gnd.n4401 19.3944
R8851 gnd.n4401 gnd.n4398 19.3944
R8852 gnd.n4398 gnd.n4397 19.3944
R8853 gnd.n4397 gnd.n4394 19.3944
R8854 gnd.n4394 gnd.n4393 19.3944
R8855 gnd.n4393 gnd.n4390 19.3944
R8856 gnd.n4390 gnd.n4389 19.3944
R8857 gnd.n4389 gnd.n4386 19.3944
R8858 gnd.n4386 gnd.n4385 19.3944
R8859 gnd.n4385 gnd.n4382 19.3944
R8860 gnd.n4382 gnd.n4381 19.3944
R8861 gnd.n4381 gnd.n4378 19.3944
R8862 gnd.n4378 gnd.n4377 19.3944
R8863 gnd.n4377 gnd.n4374 19.3944
R8864 gnd.n4374 gnd.n4373 19.3944
R8865 gnd.n4373 gnd.n4370 19.3944
R8866 gnd.n4370 gnd.n4369 19.3944
R8867 gnd.n4369 gnd.n1946 19.3944
R8868 gnd.n4536 gnd.n1946 19.3944
R8869 gnd.n2775 gnd.n2774 19.3944
R8870 gnd.n2774 gnd.n2773 19.3944
R8871 gnd.n2773 gnd.n2772 19.3944
R8872 gnd.n2772 gnd.n2770 19.3944
R8873 gnd.n2770 gnd.n2767 19.3944
R8874 gnd.n2767 gnd.n2766 19.3944
R8875 gnd.n2766 gnd.n2763 19.3944
R8876 gnd.n2763 gnd.n2762 19.3944
R8877 gnd.n2762 gnd.n2759 19.3944
R8878 gnd.n2759 gnd.n2758 19.3944
R8879 gnd.n2758 gnd.n2755 19.3944
R8880 gnd.n2755 gnd.n2754 19.3944
R8881 gnd.n2754 gnd.n2751 19.3944
R8882 gnd.n2751 gnd.n2750 19.3944
R8883 gnd.n2750 gnd.n2747 19.3944
R8884 gnd.n2747 gnd.n2746 19.3944
R8885 gnd.n2746 gnd.n2743 19.3944
R8886 gnd.n2743 gnd.n2742 19.3944
R8887 gnd.n2742 gnd.n2739 19.3944
R8888 gnd.n2739 gnd.n2738 19.3944
R8889 gnd.n2738 gnd.n2735 19.3944
R8890 gnd.n2735 gnd.n2734 19.3944
R8891 gnd.n2731 gnd.n2730 19.3944
R8892 gnd.n2730 gnd.n2686 19.3944
R8893 gnd.n2781 gnd.n2686 19.3944
R8894 gnd.n3547 gnd.n3546 19.3944
R8895 gnd.n3546 gnd.n3543 19.3944
R8896 gnd.n3543 gnd.n3542 19.3944
R8897 gnd.n3592 gnd.n3591 19.3944
R8898 gnd.n3591 gnd.n3590 19.3944
R8899 gnd.n3590 gnd.n3587 19.3944
R8900 gnd.n3587 gnd.n3586 19.3944
R8901 gnd.n3586 gnd.n3583 19.3944
R8902 gnd.n3583 gnd.n3582 19.3944
R8903 gnd.n3582 gnd.n3579 19.3944
R8904 gnd.n3579 gnd.n3578 19.3944
R8905 gnd.n3578 gnd.n3575 19.3944
R8906 gnd.n3575 gnd.n3574 19.3944
R8907 gnd.n3574 gnd.n3571 19.3944
R8908 gnd.n3571 gnd.n3570 19.3944
R8909 gnd.n3570 gnd.n3567 19.3944
R8910 gnd.n3567 gnd.n3566 19.3944
R8911 gnd.n3566 gnd.n3563 19.3944
R8912 gnd.n3563 gnd.n3562 19.3944
R8913 gnd.n3562 gnd.n3559 19.3944
R8914 gnd.n3559 gnd.n3558 19.3944
R8915 gnd.n3558 gnd.n3555 19.3944
R8916 gnd.n3555 gnd.n3554 19.3944
R8917 gnd.n3554 gnd.n3551 19.3944
R8918 gnd.n3551 gnd.n3550 19.3944
R8919 gnd.n2874 gnd.n2583 19.3944
R8920 gnd.n2884 gnd.n2583 19.3944
R8921 gnd.n2885 gnd.n2884 19.3944
R8922 gnd.n2885 gnd.n2564 19.3944
R8923 gnd.n2905 gnd.n2564 19.3944
R8924 gnd.n2905 gnd.n2556 19.3944
R8925 gnd.n2915 gnd.n2556 19.3944
R8926 gnd.n2916 gnd.n2915 19.3944
R8927 gnd.n2917 gnd.n2916 19.3944
R8928 gnd.n2917 gnd.n2539 19.3944
R8929 gnd.n2934 gnd.n2539 19.3944
R8930 gnd.n2937 gnd.n2934 19.3944
R8931 gnd.n2937 gnd.n2936 19.3944
R8932 gnd.n2936 gnd.n2512 19.3944
R8933 gnd.n2976 gnd.n2512 19.3944
R8934 gnd.n2976 gnd.n2509 19.3944
R8935 gnd.n2982 gnd.n2509 19.3944
R8936 gnd.n2983 gnd.n2982 19.3944
R8937 gnd.n2983 gnd.n2507 19.3944
R8938 gnd.n2989 gnd.n2507 19.3944
R8939 gnd.n2992 gnd.n2989 19.3944
R8940 gnd.n2994 gnd.n2992 19.3944
R8941 gnd.n3000 gnd.n2994 19.3944
R8942 gnd.n3000 gnd.n2999 19.3944
R8943 gnd.n2999 gnd.n2370 19.3944
R8944 gnd.n3066 gnd.n2370 19.3944
R8945 gnd.n3067 gnd.n3066 19.3944
R8946 gnd.n3067 gnd.n2363 19.3944
R8947 gnd.n3078 gnd.n2363 19.3944
R8948 gnd.n3079 gnd.n3078 19.3944
R8949 gnd.n3079 gnd.n2346 19.3944
R8950 gnd.n2346 gnd.n2344 19.3944
R8951 gnd.n3103 gnd.n2344 19.3944
R8952 gnd.n3104 gnd.n3103 19.3944
R8953 gnd.n3104 gnd.n2315 19.3944
R8954 gnd.n3151 gnd.n2315 19.3944
R8955 gnd.n3152 gnd.n3151 19.3944
R8956 gnd.n3152 gnd.n2308 19.3944
R8957 gnd.n3163 gnd.n2308 19.3944
R8958 gnd.n3164 gnd.n3163 19.3944
R8959 gnd.n3164 gnd.n2291 19.3944
R8960 gnd.n2291 gnd.n2289 19.3944
R8961 gnd.n3188 gnd.n2289 19.3944
R8962 gnd.n3189 gnd.n3188 19.3944
R8963 gnd.n3189 gnd.n2261 19.3944
R8964 gnd.n3240 gnd.n2261 19.3944
R8965 gnd.n3241 gnd.n3240 19.3944
R8966 gnd.n3241 gnd.n2254 19.3944
R8967 gnd.n3508 gnd.n2254 19.3944
R8968 gnd.n3509 gnd.n3508 19.3944
R8969 gnd.n3509 gnd.n2235 19.3944
R8970 gnd.n3534 gnd.n2235 19.3944
R8971 gnd.n3534 gnd.n2236 19.3944
R8972 gnd.n2865 gnd.n2864 19.3944
R8973 gnd.n2864 gnd.n2597 19.3944
R8974 gnd.n2620 gnd.n2597 19.3944
R8975 gnd.n2623 gnd.n2620 19.3944
R8976 gnd.n2623 gnd.n2616 19.3944
R8977 gnd.n2627 gnd.n2616 19.3944
R8978 gnd.n2630 gnd.n2627 19.3944
R8979 gnd.n2633 gnd.n2630 19.3944
R8980 gnd.n2633 gnd.n2614 19.3944
R8981 gnd.n2637 gnd.n2614 19.3944
R8982 gnd.n2640 gnd.n2637 19.3944
R8983 gnd.n2643 gnd.n2640 19.3944
R8984 gnd.n2643 gnd.n2612 19.3944
R8985 gnd.n2647 gnd.n2612 19.3944
R8986 gnd.n2870 gnd.n2869 19.3944
R8987 gnd.n2869 gnd.n2573 19.3944
R8988 gnd.n2895 gnd.n2573 19.3944
R8989 gnd.n2895 gnd.n2571 19.3944
R8990 gnd.n2901 gnd.n2571 19.3944
R8991 gnd.n2901 gnd.n2900 19.3944
R8992 gnd.n2900 gnd.n2545 19.3944
R8993 gnd.n2925 gnd.n2545 19.3944
R8994 gnd.n2925 gnd.n2543 19.3944
R8995 gnd.n2929 gnd.n2543 19.3944
R8996 gnd.n2929 gnd.n2523 19.3944
R8997 gnd.n2956 gnd.n2523 19.3944
R8998 gnd.n2956 gnd.n2521 19.3944
R8999 gnd.n2966 gnd.n2521 19.3944
R9000 gnd.n2966 gnd.n2965 19.3944
R9001 gnd.n2965 gnd.n2964 19.3944
R9002 gnd.n2964 gnd.n2470 19.3944
R9003 gnd.n3014 gnd.n2470 19.3944
R9004 gnd.n3014 gnd.n3013 19.3944
R9005 gnd.n3013 gnd.n3012 19.3944
R9006 gnd.n3012 gnd.n2474 19.3944
R9007 gnd.n2494 gnd.n2474 19.3944
R9008 gnd.n2494 gnd.n2380 19.3944
R9009 gnd.n3051 gnd.n2380 19.3944
R9010 gnd.n3051 gnd.n2378 19.3944
R9011 gnd.n3057 gnd.n2378 19.3944
R9012 gnd.n3057 gnd.n3056 19.3944
R9013 gnd.n3056 gnd.n2353 19.3944
R9014 gnd.n3091 gnd.n2353 19.3944
R9015 gnd.n3091 gnd.n2351 19.3944
R9016 gnd.n3097 gnd.n2351 19.3944
R9017 gnd.n3097 gnd.n3096 19.3944
R9018 gnd.n3096 gnd.n2326 19.3944
R9019 gnd.n3136 gnd.n2326 19.3944
R9020 gnd.n3136 gnd.n2324 19.3944
R9021 gnd.n3142 gnd.n2324 19.3944
R9022 gnd.n3142 gnd.n3141 19.3944
R9023 gnd.n3141 gnd.n2298 19.3944
R9024 gnd.n3176 gnd.n2298 19.3944
R9025 gnd.n3176 gnd.n2296 19.3944
R9026 gnd.n3182 gnd.n2296 19.3944
R9027 gnd.n3182 gnd.n3181 19.3944
R9028 gnd.n3181 gnd.n2271 19.3944
R9029 gnd.n3225 gnd.n2271 19.3944
R9030 gnd.n3225 gnd.n2269 19.3944
R9031 gnd.n3231 gnd.n2269 19.3944
R9032 gnd.n3231 gnd.n3230 19.3944
R9033 gnd.n3230 gnd.n2244 19.3944
R9034 gnd.n3519 gnd.n2244 19.3944
R9035 gnd.n3519 gnd.n2242 19.3944
R9036 gnd.n3527 gnd.n2242 19.3944
R9037 gnd.n3527 gnd.n3526 19.3944
R9038 gnd.n3526 gnd.n3525 19.3944
R9039 gnd.n3628 gnd.n3627 19.3944
R9040 gnd.n3627 gnd.n2183 19.3944
R9041 gnd.n3623 gnd.n2183 19.3944
R9042 gnd.n3623 gnd.n3620 19.3944
R9043 gnd.n3620 gnd.n3617 19.3944
R9044 gnd.n3617 gnd.n3616 19.3944
R9045 gnd.n3616 gnd.n3613 19.3944
R9046 gnd.n3613 gnd.n3612 19.3944
R9047 gnd.n3612 gnd.n3609 19.3944
R9048 gnd.n3609 gnd.n3608 19.3944
R9049 gnd.n3608 gnd.n3605 19.3944
R9050 gnd.n3605 gnd.n3604 19.3944
R9051 gnd.n3604 gnd.n3601 19.3944
R9052 gnd.n3601 gnd.n3600 19.3944
R9053 gnd.n2785 gnd.n2684 19.3944
R9054 gnd.n2785 gnd.n2675 19.3944
R9055 gnd.n2798 gnd.n2675 19.3944
R9056 gnd.n2798 gnd.n2673 19.3944
R9057 gnd.n2802 gnd.n2673 19.3944
R9058 gnd.n2802 gnd.n2663 19.3944
R9059 gnd.n2814 gnd.n2663 19.3944
R9060 gnd.n2814 gnd.n2661 19.3944
R9061 gnd.n2848 gnd.n2661 19.3944
R9062 gnd.n2848 gnd.n2847 19.3944
R9063 gnd.n2847 gnd.n2846 19.3944
R9064 gnd.n2846 gnd.n2845 19.3944
R9065 gnd.n2845 gnd.n2842 19.3944
R9066 gnd.n2842 gnd.n2841 19.3944
R9067 gnd.n2841 gnd.n2840 19.3944
R9068 gnd.n2840 gnd.n2838 19.3944
R9069 gnd.n2838 gnd.n2837 19.3944
R9070 gnd.n2837 gnd.n2834 19.3944
R9071 gnd.n2834 gnd.n2833 19.3944
R9072 gnd.n2833 gnd.n2832 19.3944
R9073 gnd.n2832 gnd.n2830 19.3944
R9074 gnd.n2830 gnd.n2529 19.3944
R9075 gnd.n2945 gnd.n2529 19.3944
R9076 gnd.n2945 gnd.n2527 19.3944
R9077 gnd.n2951 gnd.n2527 19.3944
R9078 gnd.n2951 gnd.n2950 19.3944
R9079 gnd.n2950 gnd.n2451 19.3944
R9080 gnd.n3025 gnd.n2451 19.3944
R9081 gnd.n3025 gnd.n2452 19.3944
R9082 gnd.n2499 gnd.n2498 19.3944
R9083 gnd.n2502 gnd.n2501 19.3944
R9084 gnd.n2489 gnd.n2488 19.3944
R9085 gnd.n3044 gnd.n2385 19.3944
R9086 gnd.n3044 gnd.n3043 19.3944
R9087 gnd.n3043 gnd.n3042 19.3944
R9088 gnd.n3042 gnd.n3040 19.3944
R9089 gnd.n3040 gnd.n3039 19.3944
R9090 gnd.n3039 gnd.n3037 19.3944
R9091 gnd.n3037 gnd.n3036 19.3944
R9092 gnd.n3036 gnd.n2334 19.3944
R9093 gnd.n3112 gnd.n2334 19.3944
R9094 gnd.n3112 gnd.n2332 19.3944
R9095 gnd.n3131 gnd.n2332 19.3944
R9096 gnd.n3131 gnd.n3130 19.3944
R9097 gnd.n3130 gnd.n3129 19.3944
R9098 gnd.n3129 gnd.n3127 19.3944
R9099 gnd.n3127 gnd.n3126 19.3944
R9100 gnd.n3126 gnd.n3124 19.3944
R9101 gnd.n3124 gnd.n3123 19.3944
R9102 gnd.n3123 gnd.n2278 19.3944
R9103 gnd.n3197 gnd.n2278 19.3944
R9104 gnd.n3197 gnd.n2276 19.3944
R9105 gnd.n3220 gnd.n2276 19.3944
R9106 gnd.n3220 gnd.n3219 19.3944
R9107 gnd.n3219 gnd.n3218 19.3944
R9108 gnd.n3218 gnd.n3215 19.3944
R9109 gnd.n3215 gnd.n3214 19.3944
R9110 gnd.n3214 gnd.n3212 19.3944
R9111 gnd.n3212 gnd.n3211 19.3944
R9112 gnd.n3211 gnd.n3209 19.3944
R9113 gnd.n3209 gnd.n2230 19.3944
R9114 gnd.n2790 gnd.n2680 19.3944
R9115 gnd.n2790 gnd.n2678 19.3944
R9116 gnd.n2794 gnd.n2678 19.3944
R9117 gnd.n2794 gnd.n2669 19.3944
R9118 gnd.n2806 gnd.n2669 19.3944
R9119 gnd.n2806 gnd.n2667 19.3944
R9120 gnd.n2810 gnd.n2667 19.3944
R9121 gnd.n2810 gnd.n2656 19.3944
R9122 gnd.n2852 gnd.n2656 19.3944
R9123 gnd.n2852 gnd.n2610 19.3944
R9124 gnd.n2858 gnd.n2610 19.3944
R9125 gnd.n2858 gnd.n2857 19.3944
R9126 gnd.n2857 gnd.n2588 19.3944
R9127 gnd.n2879 gnd.n2588 19.3944
R9128 gnd.n2879 gnd.n2581 19.3944
R9129 gnd.n2890 gnd.n2581 19.3944
R9130 gnd.n2890 gnd.n2889 19.3944
R9131 gnd.n2889 gnd.n2562 19.3944
R9132 gnd.n2910 gnd.n2562 19.3944
R9133 gnd.n2910 gnd.n2552 19.3944
R9134 gnd.n2920 gnd.n2552 19.3944
R9135 gnd.n2920 gnd.n2535 19.3944
R9136 gnd.n2941 gnd.n2535 19.3944
R9137 gnd.n2941 gnd.n2940 19.3944
R9138 gnd.n2940 gnd.n2514 19.3944
R9139 gnd.n2971 gnd.n2514 19.3944
R9140 gnd.n2971 gnd.n2459 19.3944
R9141 gnd.n3021 gnd.n2459 19.3944
R9142 gnd.n3021 gnd.n3020 19.3944
R9143 gnd.n3020 gnd.n3019 19.3944
R9144 gnd.n3019 gnd.n2463 19.3944
R9145 gnd.n2481 gnd.n2463 19.3944
R9146 gnd.n3007 gnd.n2481 19.3944
R9147 gnd.n3007 gnd.n3006 19.3944
R9148 gnd.n3006 gnd.n3005 19.3944
R9149 gnd.n3005 gnd.n2485 19.3944
R9150 gnd.n2485 gnd.n2372 19.3944
R9151 gnd.n3062 gnd.n2372 19.3944
R9152 gnd.n3062 gnd.n2365 19.3944
R9153 gnd.n3073 gnd.n2365 19.3944
R9154 gnd.n3073 gnd.n2361 19.3944
R9155 gnd.n3086 gnd.n2361 19.3944
R9156 gnd.n3086 gnd.n3085 19.3944
R9157 gnd.n3085 gnd.n2340 19.3944
R9158 gnd.n3108 gnd.n2340 19.3944
R9159 gnd.n3108 gnd.n3107 19.3944
R9160 gnd.n3107 gnd.n2317 19.3944
R9161 gnd.n3147 gnd.n2317 19.3944
R9162 gnd.n3147 gnd.n2310 19.3944
R9163 gnd.n3158 gnd.n2310 19.3944
R9164 gnd.n3158 gnd.n2306 19.3944
R9165 gnd.n3171 gnd.n2306 19.3944
R9166 gnd.n3171 gnd.n3170 19.3944
R9167 gnd.n3170 gnd.n2285 19.3944
R9168 gnd.n3193 gnd.n2285 19.3944
R9169 gnd.n3193 gnd.n3192 19.3944
R9170 gnd.n3192 gnd.n2263 19.3944
R9171 gnd.n3236 gnd.n2263 19.3944
R9172 gnd.n3236 gnd.n2256 19.3944
R9173 gnd.n3247 gnd.n2256 19.3944
R9174 gnd.n3247 gnd.n2252 19.3944
R9175 gnd.n3514 gnd.n2252 19.3944
R9176 gnd.n3514 gnd.n3513 19.3944
R9177 gnd.n3513 gnd.n2233 19.3944
R9178 gnd.n3537 gnd.n2233 19.3944
R9179 gnd.n3873 gnd.n3871 19.3944
R9180 gnd.n3873 gnd.n3730 19.3944
R9181 gnd.n3878 gnd.n3730 19.3944
R9182 gnd.n3879 gnd.n3878 19.3944
R9183 gnd.n3881 gnd.n3879 19.3944
R9184 gnd.n3881 gnd.n3728 19.3944
R9185 gnd.n3886 gnd.n3728 19.3944
R9186 gnd.n3887 gnd.n3886 19.3944
R9187 gnd.n3889 gnd.n3887 19.3944
R9188 gnd.n3889 gnd.n3726 19.3944
R9189 gnd.n3894 gnd.n3726 19.3944
R9190 gnd.n3895 gnd.n3894 19.3944
R9191 gnd.n3897 gnd.n3895 19.3944
R9192 gnd.n3897 gnd.n3724 19.3944
R9193 gnd.n3902 gnd.n3724 19.3944
R9194 gnd.n3903 gnd.n3902 19.3944
R9195 gnd.n3905 gnd.n3903 19.3944
R9196 gnd.n3905 gnd.n3722 19.3944
R9197 gnd.n3910 gnd.n3722 19.3944
R9198 gnd.n3911 gnd.n3910 19.3944
R9199 gnd.n3913 gnd.n3911 19.3944
R9200 gnd.n3913 gnd.n3720 19.3944
R9201 gnd.n3918 gnd.n3720 19.3944
R9202 gnd.n3919 gnd.n3918 19.3944
R9203 gnd.n3921 gnd.n3919 19.3944
R9204 gnd.n3921 gnd.n3718 19.3944
R9205 gnd.n3926 gnd.n3718 19.3944
R9206 gnd.n3927 gnd.n3926 19.3944
R9207 gnd.n3929 gnd.n3927 19.3944
R9208 gnd.n3929 gnd.n3716 19.3944
R9209 gnd.n3934 gnd.n3716 19.3944
R9210 gnd.n3935 gnd.n3934 19.3944
R9211 gnd.n3938 gnd.n3935 19.3944
R9212 gnd.n3939 gnd.n3938 19.3944
R9213 gnd.n3941 gnd.n3939 19.3944
R9214 gnd.n3941 gnd.n3714 19.3944
R9215 gnd.n3946 gnd.n3714 19.3944
R9216 gnd.n3947 gnd.n3946 19.3944
R9217 gnd.n3949 gnd.n3947 19.3944
R9218 gnd.n3949 gnd.n3712 19.3944
R9219 gnd.n3954 gnd.n3712 19.3944
R9220 gnd.n3955 gnd.n3954 19.3944
R9221 gnd.n3957 gnd.n3955 19.3944
R9222 gnd.n3957 gnd.n3710 19.3944
R9223 gnd.n3964 gnd.n3710 19.3944
R9224 gnd.n3965 gnd.n3964 19.3944
R9225 gnd.n3969 gnd.n3965 19.3944
R9226 gnd.n3969 gnd.n3708 19.3944
R9227 gnd.n3978 gnd.n3708 19.3944
R9228 gnd.n3978 gnd.n3977 19.3944
R9229 gnd.n3977 gnd.n3976 19.3944
R9230 gnd.n3976 gnd.n1931 19.3944
R9231 gnd.n4573 gnd.n1931 19.3944
R9232 gnd.n4574 gnd.n4573 19.3944
R9233 gnd.n4575 gnd.n4574 19.3944
R9234 gnd.n4575 gnd.n1929 19.3944
R9235 gnd.n4581 gnd.n1929 19.3944
R9236 gnd.n4582 gnd.n4581 19.3944
R9237 gnd.n4585 gnd.n4582 19.3944
R9238 gnd.n4585 gnd.n1927 19.3944
R9239 gnd.n4590 gnd.n1927 19.3944
R9240 gnd.n4590 gnd.n1163 19.3944
R9241 gnd.n6180 gnd.n1163 19.3944
R9242 gnd.n6181 gnd.n6180 19.3944
R9243 gnd.n6219 gnd.n6218 19.3944
R9244 gnd.n6218 gnd.n6217 19.3944
R9245 gnd.n6217 gnd.n1129 19.3944
R9246 gnd.n6212 gnd.n1129 19.3944
R9247 gnd.n6212 gnd.n6211 19.3944
R9248 gnd.n6211 gnd.n6210 19.3944
R9249 gnd.n6210 gnd.n1136 19.3944
R9250 gnd.n6205 gnd.n1136 19.3944
R9251 gnd.n6205 gnd.n6204 19.3944
R9252 gnd.n6204 gnd.n6203 19.3944
R9253 gnd.n6203 gnd.n1143 19.3944
R9254 gnd.n6198 gnd.n1143 19.3944
R9255 gnd.n6198 gnd.n6197 19.3944
R9256 gnd.n6197 gnd.n6196 19.3944
R9257 gnd.n6196 gnd.n1150 19.3944
R9258 gnd.n6191 gnd.n1150 19.3944
R9259 gnd.n6191 gnd.n6190 19.3944
R9260 gnd.n6190 gnd.n6189 19.3944
R9261 gnd.n6250 gnd.n6249 19.3944
R9262 gnd.n6249 gnd.n1095 19.3944
R9263 gnd.n1097 gnd.n1095 19.3944
R9264 gnd.n6242 gnd.n1097 19.3944
R9265 gnd.n6242 gnd.n6241 19.3944
R9266 gnd.n6241 gnd.n6240 19.3944
R9267 gnd.n6240 gnd.n1104 19.3944
R9268 gnd.n6235 gnd.n1104 19.3944
R9269 gnd.n6235 gnd.n6234 19.3944
R9270 gnd.n6234 gnd.n6233 19.3944
R9271 gnd.n6233 gnd.n1111 19.3944
R9272 gnd.n6228 gnd.n1111 19.3944
R9273 gnd.n6228 gnd.n6227 19.3944
R9274 gnd.n6227 gnd.n6226 19.3944
R9275 gnd.n6226 gnd.n1118 19.3944
R9276 gnd.n4105 gnd.n2154 19.3944
R9277 gnd.n4109 gnd.n2154 19.3944
R9278 gnd.n4109 gnd.n2141 19.3944
R9279 gnd.n4121 gnd.n2141 19.3944
R9280 gnd.n4121 gnd.n2139 19.3944
R9281 gnd.n4125 gnd.n2139 19.3944
R9282 gnd.n4125 gnd.n2124 19.3944
R9283 gnd.n4137 gnd.n2124 19.3944
R9284 gnd.n4137 gnd.n2122 19.3944
R9285 gnd.n4141 gnd.n2122 19.3944
R9286 gnd.n4141 gnd.n2109 19.3944
R9287 gnd.n4153 gnd.n2109 19.3944
R9288 gnd.n4153 gnd.n2107 19.3944
R9289 gnd.n4157 gnd.n2107 19.3944
R9290 gnd.n4157 gnd.n2092 19.3944
R9291 gnd.n4169 gnd.n2092 19.3944
R9292 gnd.n4169 gnd.n2090 19.3944
R9293 gnd.n4173 gnd.n2090 19.3944
R9294 gnd.n4173 gnd.n2077 19.3944
R9295 gnd.n4185 gnd.n2077 19.3944
R9296 gnd.n4185 gnd.n2075 19.3944
R9297 gnd.n4189 gnd.n2075 19.3944
R9298 gnd.n4189 gnd.n2060 19.3944
R9299 gnd.n4201 gnd.n2060 19.3944
R9300 gnd.n4201 gnd.n2058 19.3944
R9301 gnd.n4205 gnd.n2058 19.3944
R9302 gnd.n4205 gnd.n2045 19.3944
R9303 gnd.n4217 gnd.n2045 19.3944
R9304 gnd.n4217 gnd.n2043 19.3944
R9305 gnd.n4221 gnd.n2043 19.3944
R9306 gnd.n4221 gnd.n2027 19.3944
R9307 gnd.n4233 gnd.n2027 19.3944
R9308 gnd.n4233 gnd.n2025 19.3944
R9309 gnd.n4237 gnd.n2025 19.3944
R9310 gnd.n4237 gnd.n2012 19.3944
R9311 gnd.n4249 gnd.n2012 19.3944
R9312 gnd.n4249 gnd.n2010 19.3944
R9313 gnd.n4253 gnd.n2010 19.3944
R9314 gnd.n4253 gnd.n1994 19.3944
R9315 gnd.n4275 gnd.n1994 19.3944
R9316 gnd.n4275 gnd.n1992 19.3944
R9317 gnd.n4280 gnd.n1992 19.3944
R9318 gnd.n4280 gnd.n987 19.3944
R9319 gnd.n6313 gnd.n987 19.3944
R9320 gnd.n6313 gnd.n6312 19.3944
R9321 gnd.n6312 gnd.n6311 19.3944
R9322 gnd.n6311 gnd.n991 19.3944
R9323 gnd.n6301 gnd.n991 19.3944
R9324 gnd.n6301 gnd.n6300 19.3944
R9325 gnd.n6300 gnd.n6299 19.3944
R9326 gnd.n6299 gnd.n1013 19.3944
R9327 gnd.n6289 gnd.n1013 19.3944
R9328 gnd.n6289 gnd.n6288 19.3944
R9329 gnd.n6288 gnd.n6287 19.3944
R9330 gnd.n6287 gnd.n1034 19.3944
R9331 gnd.n6277 gnd.n1034 19.3944
R9332 gnd.n6277 gnd.n6276 19.3944
R9333 gnd.n6276 gnd.n6275 19.3944
R9334 gnd.n6275 gnd.n1055 19.3944
R9335 gnd.n6265 gnd.n1055 19.3944
R9336 gnd.n6265 gnd.n6264 19.3944
R9337 gnd.n6264 gnd.n6263 19.3944
R9338 gnd.n6263 gnd.n1077 19.3944
R9339 gnd.n6253 gnd.n1077 19.3944
R9340 gnd.n3776 gnd.n3773 19.3944
R9341 gnd.n3776 gnd.n3772 19.3944
R9342 gnd.n3780 gnd.n3772 19.3944
R9343 gnd.n3780 gnd.n3770 19.3944
R9344 gnd.n3786 gnd.n3770 19.3944
R9345 gnd.n3786 gnd.n3768 19.3944
R9346 gnd.n3790 gnd.n3768 19.3944
R9347 gnd.n3790 gnd.n3766 19.3944
R9348 gnd.n3796 gnd.n3766 19.3944
R9349 gnd.n3796 gnd.n3764 19.3944
R9350 gnd.n3800 gnd.n3764 19.3944
R9351 gnd.n3800 gnd.n3762 19.3944
R9352 gnd.n3806 gnd.n3762 19.3944
R9353 gnd.n3806 gnd.n3760 19.3944
R9354 gnd.n3810 gnd.n3760 19.3944
R9355 gnd.n3810 gnd.n3755 19.3944
R9356 gnd.n3816 gnd.n3755 19.3944
R9357 gnd.n3820 gnd.n3753 19.3944
R9358 gnd.n3820 gnd.n3751 19.3944
R9359 gnd.n3826 gnd.n3751 19.3944
R9360 gnd.n3826 gnd.n3749 19.3944
R9361 gnd.n3830 gnd.n3749 19.3944
R9362 gnd.n3830 gnd.n3747 19.3944
R9363 gnd.n3836 gnd.n3747 19.3944
R9364 gnd.n3836 gnd.n3745 19.3944
R9365 gnd.n3840 gnd.n3745 19.3944
R9366 gnd.n3840 gnd.n3743 19.3944
R9367 gnd.n3846 gnd.n3743 19.3944
R9368 gnd.n3846 gnd.n3741 19.3944
R9369 gnd.n3850 gnd.n3741 19.3944
R9370 gnd.n3850 gnd.n3739 19.3944
R9371 gnd.n3856 gnd.n3739 19.3944
R9372 gnd.n3856 gnd.n3737 19.3944
R9373 gnd.n3861 gnd.n3737 19.3944
R9374 gnd.n3861 gnd.n3735 19.3944
R9375 gnd.n4098 gnd.n4097 19.3944
R9376 gnd.n4097 gnd.n3637 19.3944
R9377 gnd.n4091 gnd.n3637 19.3944
R9378 gnd.n4091 gnd.n4090 19.3944
R9379 gnd.n4090 gnd.n4089 19.3944
R9380 gnd.n4089 gnd.n3643 19.3944
R9381 gnd.n4083 gnd.n3643 19.3944
R9382 gnd.n4083 gnd.n4082 19.3944
R9383 gnd.n4082 gnd.n4081 19.3944
R9384 gnd.n4081 gnd.n3649 19.3944
R9385 gnd.n4075 gnd.n3649 19.3944
R9386 gnd.n4075 gnd.n4074 19.3944
R9387 gnd.n4074 gnd.n4073 19.3944
R9388 gnd.n4073 gnd.n3655 19.3944
R9389 gnd.n4067 gnd.n3655 19.3944
R9390 gnd.n4067 gnd.n4066 19.3944
R9391 gnd.n4057 gnd.n4056 19.3944
R9392 gnd.n4056 gnd.n4054 19.3944
R9393 gnd.n4054 gnd.n4053 19.3944
R9394 gnd.n4053 gnd.n4051 19.3944
R9395 gnd.n4051 gnd.n4050 19.3944
R9396 gnd.n4050 gnd.n4048 19.3944
R9397 gnd.n4048 gnd.n4047 19.3944
R9398 gnd.n4047 gnd.n4045 19.3944
R9399 gnd.n4045 gnd.n4044 19.3944
R9400 gnd.n4044 gnd.n4042 19.3944
R9401 gnd.n4042 gnd.n4041 19.3944
R9402 gnd.n4041 gnd.n4039 19.3944
R9403 gnd.n4039 gnd.n4038 19.3944
R9404 gnd.n4038 gnd.n4036 19.3944
R9405 gnd.n4036 gnd.n4035 19.3944
R9406 gnd.n4035 gnd.n4033 19.3944
R9407 gnd.n4033 gnd.n4032 19.3944
R9408 gnd.n4032 gnd.n4030 19.3944
R9409 gnd.n4030 gnd.n4029 19.3944
R9410 gnd.n4029 gnd.n4027 19.3944
R9411 gnd.n4027 gnd.n4026 19.3944
R9412 gnd.n4026 gnd.n4024 19.3944
R9413 gnd.n4024 gnd.n4023 19.3944
R9414 gnd.n4023 gnd.n4021 19.3944
R9415 gnd.n4021 gnd.n4020 19.3944
R9416 gnd.n4020 gnd.n4018 19.3944
R9417 gnd.n4018 gnd.n4017 19.3944
R9418 gnd.n4017 gnd.n4015 19.3944
R9419 gnd.n4015 gnd.n4014 19.3944
R9420 gnd.n4014 gnd.n4012 19.3944
R9421 gnd.n4012 gnd.n4011 19.3944
R9422 gnd.n4011 gnd.n4009 19.3944
R9423 gnd.n4009 gnd.n3694 19.3944
R9424 gnd.n4005 gnd.n3694 19.3944
R9425 gnd.n4005 gnd.n4004 19.3944
R9426 gnd.n4004 gnd.n4003 19.3944
R9427 gnd.n4003 gnd.n3698 19.3944
R9428 gnd.n3999 gnd.n3698 19.3944
R9429 gnd.n3999 gnd.n3998 19.3944
R9430 gnd.n3998 gnd.n3997 19.3944
R9431 gnd.n3997 gnd.n3702 19.3944
R9432 gnd.n3993 gnd.n3702 19.3944
R9433 gnd.n3993 gnd.n3992 19.3944
R9434 gnd.n3992 gnd.n3991 19.3944
R9435 gnd.n3991 gnd.n3705 19.3944
R9436 gnd.n3987 gnd.n3705 19.3944
R9437 gnd.n3987 gnd.n3986 19.3944
R9438 gnd.n3986 gnd.n3985 19.3944
R9439 gnd.n3985 gnd.n3982 19.3944
R9440 gnd.n3982 gnd.n1935 19.3944
R9441 gnd.n4565 gnd.n1935 19.3944
R9442 gnd.n4565 gnd.n1933 19.3944
R9443 gnd.n4569 gnd.n1933 19.3944
R9444 gnd.n4569 gnd.n1920 19.3944
R9445 gnd.n4604 gnd.n1920 19.3944
R9446 gnd.n4604 gnd.n1921 19.3944
R9447 gnd.n4600 gnd.n1921 19.3944
R9448 gnd.n4600 gnd.n4599 19.3944
R9449 gnd.n4599 gnd.n4598 19.3944
R9450 gnd.n4598 gnd.n1926 19.3944
R9451 gnd.n4594 gnd.n1926 19.3944
R9452 gnd.n4594 gnd.n1165 19.3944
R9453 gnd.n6176 gnd.n1165 19.3944
R9454 gnd.n6176 gnd.n1166 19.3944
R9455 gnd.n4101 gnd.n2149 19.3944
R9456 gnd.n4113 gnd.n2149 19.3944
R9457 gnd.n4113 gnd.n2147 19.3944
R9458 gnd.n4117 gnd.n2147 19.3944
R9459 gnd.n4117 gnd.n2133 19.3944
R9460 gnd.n4129 gnd.n2133 19.3944
R9461 gnd.n4129 gnd.n2131 19.3944
R9462 gnd.n4133 gnd.n2131 19.3944
R9463 gnd.n4133 gnd.n2117 19.3944
R9464 gnd.n4145 gnd.n2117 19.3944
R9465 gnd.n4145 gnd.n2115 19.3944
R9466 gnd.n4149 gnd.n2115 19.3944
R9467 gnd.n4149 gnd.n2101 19.3944
R9468 gnd.n4161 gnd.n2101 19.3944
R9469 gnd.n4161 gnd.n2099 19.3944
R9470 gnd.n4165 gnd.n2099 19.3944
R9471 gnd.n4165 gnd.n2085 19.3944
R9472 gnd.n4177 gnd.n2085 19.3944
R9473 gnd.n4177 gnd.n2083 19.3944
R9474 gnd.n4181 gnd.n2083 19.3944
R9475 gnd.n4181 gnd.n2069 19.3944
R9476 gnd.n4193 gnd.n2069 19.3944
R9477 gnd.n4193 gnd.n2067 19.3944
R9478 gnd.n4197 gnd.n2067 19.3944
R9479 gnd.n4197 gnd.n2053 19.3944
R9480 gnd.n4209 gnd.n2053 19.3944
R9481 gnd.n4209 gnd.n2051 19.3944
R9482 gnd.n4213 gnd.n2051 19.3944
R9483 gnd.n4213 gnd.n2037 19.3944
R9484 gnd.n4225 gnd.n2037 19.3944
R9485 gnd.n4225 gnd.n2034 19.3944
R9486 gnd.n4229 gnd.n2034 19.3944
R9487 gnd.n4229 gnd.n2019 19.3944
R9488 gnd.n4241 gnd.n2019 19.3944
R9489 gnd.n4241 gnd.n2017 19.3944
R9490 gnd.n4245 gnd.n2017 19.3944
R9491 gnd.n4245 gnd.n2004 19.3944
R9492 gnd.n4257 gnd.n2004 19.3944
R9493 gnd.n4257 gnd.n2002 19.3944
R9494 gnd.n4271 gnd.n2002 19.3944
R9495 gnd.n4271 gnd.n4270 19.3944
R9496 gnd.n4270 gnd.n4269 19.3944
R9497 gnd.n4269 gnd.n4268 19.3944
R9498 gnd.n4268 gnd.n4266 19.3944
R9499 gnd.n4266 gnd.n998 19.3944
R9500 gnd.n6307 gnd.n998 19.3944
R9501 gnd.n6307 gnd.n6306 19.3944
R9502 gnd.n6306 gnd.n6305 19.3944
R9503 gnd.n6305 gnd.n1002 19.3944
R9504 gnd.n6295 gnd.n1002 19.3944
R9505 gnd.n6295 gnd.n6294 19.3944
R9506 gnd.n6294 gnd.n6293 19.3944
R9507 gnd.n6293 gnd.n1024 19.3944
R9508 gnd.n6283 gnd.n1024 19.3944
R9509 gnd.n6283 gnd.n6282 19.3944
R9510 gnd.n6282 gnd.n6281 19.3944
R9511 gnd.n6281 gnd.n1044 19.3944
R9512 gnd.n6271 gnd.n1044 19.3944
R9513 gnd.n6271 gnd.n6270 19.3944
R9514 gnd.n6270 gnd.n6269 19.3944
R9515 gnd.n6269 gnd.n1066 19.3944
R9516 gnd.n6259 gnd.n1066 19.3944
R9517 gnd.n6259 gnd.n6258 19.3944
R9518 gnd.n6258 gnd.n6257 19.3944
R9519 gnd.n4785 gnd.n1896 19.3944
R9520 gnd.n4785 gnd.n1894 19.3944
R9521 gnd.n4789 gnd.n1894 19.3944
R9522 gnd.n4789 gnd.n1882 19.3944
R9523 gnd.n4804 gnd.n1882 19.3944
R9524 gnd.n4804 gnd.n1880 19.3944
R9525 gnd.n4808 gnd.n1880 19.3944
R9526 gnd.n4808 gnd.n1868 19.3944
R9527 gnd.n4823 gnd.n1868 19.3944
R9528 gnd.n4823 gnd.n1866 19.3944
R9529 gnd.n4827 gnd.n1866 19.3944
R9530 gnd.n4827 gnd.n1854 19.3944
R9531 gnd.n4842 gnd.n1854 19.3944
R9532 gnd.n4842 gnd.n1852 19.3944
R9533 gnd.n4846 gnd.n1852 19.3944
R9534 gnd.n4846 gnd.n1840 19.3944
R9535 gnd.n4861 gnd.n1840 19.3944
R9536 gnd.n4861 gnd.n1838 19.3944
R9537 gnd.n4865 gnd.n1838 19.3944
R9538 gnd.n4865 gnd.n1826 19.3944
R9539 gnd.n5080 gnd.n1826 19.3944
R9540 gnd.n5080 gnd.n1824 19.3944
R9541 gnd.n5084 gnd.n1824 19.3944
R9542 gnd.n5084 gnd.n1760 19.3944
R9543 gnd.n5114 gnd.n1760 19.3944
R9544 gnd.n5114 gnd.n1757 19.3944
R9545 gnd.n5119 gnd.n1757 19.3944
R9546 gnd.n5119 gnd.n1758 19.3944
R9547 gnd.n1758 gnd.n1731 19.3944
R9548 gnd.n5150 gnd.n1731 19.3944
R9549 gnd.n5150 gnd.n1729 19.3944
R9550 gnd.n5154 gnd.n1729 19.3944
R9551 gnd.n5154 gnd.n1711 19.3944
R9552 gnd.n5177 gnd.n1711 19.3944
R9553 gnd.n5177 gnd.n1708 19.3944
R9554 gnd.n5182 gnd.n1708 19.3944
R9555 gnd.n5182 gnd.n1709 19.3944
R9556 gnd.n1709 gnd.n1680 19.3944
R9557 gnd.n5215 gnd.n1680 19.3944
R9558 gnd.n5215 gnd.n1677 19.3944
R9559 gnd.n5220 gnd.n1677 19.3944
R9560 gnd.n5220 gnd.n1678 19.3944
R9561 gnd.n1678 gnd.n1648 19.3944
R9562 gnd.n5268 gnd.n1648 19.3944
R9563 gnd.n5268 gnd.n1646 19.3944
R9564 gnd.n5272 gnd.n1646 19.3944
R9565 gnd.n5272 gnd.n1631 19.3944
R9566 gnd.n5311 gnd.n1631 19.3944
R9567 gnd.n5311 gnd.n1628 19.3944
R9568 gnd.n5322 gnd.n1628 19.3944
R9569 gnd.n5322 gnd.n1629 19.3944
R9570 gnd.n5318 gnd.n1629 19.3944
R9571 gnd.n5318 gnd.n5317 19.3944
R9572 gnd.n5317 gnd.n1596 19.3944
R9573 gnd.n5379 gnd.n1596 19.3944
R9574 gnd.n5379 gnd.n1593 19.3944
R9575 gnd.n5387 gnd.n1593 19.3944
R9576 gnd.n5387 gnd.n1594 19.3944
R9577 gnd.n5383 gnd.n1594 19.3944
R9578 gnd.n5383 gnd.n1570 19.3944
R9579 gnd.n5429 gnd.n1570 19.3944
R9580 gnd.n5429 gnd.n1571 19.3944
R9581 gnd.n5425 gnd.n1571 19.3944
R9582 gnd.n5425 gnd.n1548 19.3944
R9583 gnd.n5479 gnd.n1548 19.3944
R9584 gnd.n5479 gnd.n1549 19.3944
R9585 gnd.n5475 gnd.n1549 19.3944
R9586 gnd.n5475 gnd.n1523 19.3944
R9587 gnd.n5508 gnd.n1523 19.3944
R9588 gnd.n5508 gnd.n1521 19.3944
R9589 gnd.n5512 gnd.n1521 19.3944
R9590 gnd.n5512 gnd.n1499 19.3944
R9591 gnd.n5558 gnd.n1499 19.3944
R9592 gnd.n5558 gnd.n1500 19.3944
R9593 gnd.n5554 gnd.n1500 19.3944
R9594 gnd.n5554 gnd.n5553 19.3944
R9595 gnd.n5553 gnd.n5552 19.3944
R9596 gnd.n5552 gnd.n1390 19.3944
R9597 gnd.n5727 gnd.n1390 19.3944
R9598 gnd.n5727 gnd.n1388 19.3944
R9599 gnd.n5731 gnd.n1388 19.3944
R9600 gnd.n5731 gnd.n1377 19.3944
R9601 gnd.n5746 gnd.n1377 19.3944
R9602 gnd.n5746 gnd.n1375 19.3944
R9603 gnd.n5750 gnd.n1375 19.3944
R9604 gnd.n5750 gnd.n1363 19.3944
R9605 gnd.n5765 gnd.n1363 19.3944
R9606 gnd.n5765 gnd.n1361 19.3944
R9607 gnd.n5769 gnd.n1361 19.3944
R9608 gnd.n5769 gnd.n1349 19.3944
R9609 gnd.n5784 gnd.n1349 19.3944
R9610 gnd.n5784 gnd.n1347 19.3944
R9611 gnd.n5788 gnd.n1347 19.3944
R9612 gnd.n5788 gnd.n1335 19.3944
R9613 gnd.n5803 gnd.n1335 19.3944
R9614 gnd.n5803 gnd.n1333 19.3944
R9615 gnd.n5807 gnd.n1333 19.3944
R9616 gnd.n5807 gnd.n1320 19.3944
R9617 gnd.n5995 gnd.n1320 19.3944
R9618 gnd.n5995 gnd.n1318 19.3944
R9619 gnd.n5999 gnd.n1318 19.3944
R9620 gnd.n5955 gnd.n5947 19.3944
R9621 gnd.n5951 gnd.n5947 19.3944
R9622 gnd.n5951 gnd.n5950 19.3944
R9623 gnd.n7224 gnd.n7223 19.3944
R9624 gnd.n7223 gnd.n466 19.3944
R9625 gnd.n7216 gnd.n466 19.3944
R9626 gnd.n7216 gnd.n7215 19.3944
R9627 gnd.n7215 gnd.n474 19.3944
R9628 gnd.n7208 gnd.n474 19.3944
R9629 gnd.n7208 gnd.n7207 19.3944
R9630 gnd.n7207 gnd.n482 19.3944
R9631 gnd.n7200 gnd.n482 19.3944
R9632 gnd.n7200 gnd.n7199 19.3944
R9633 gnd.n7199 gnd.n490 19.3944
R9634 gnd.n7192 gnd.n490 19.3944
R9635 gnd.n7192 gnd.n7191 19.3944
R9636 gnd.n7191 gnd.n498 19.3944
R9637 gnd.n7184 gnd.n498 19.3944
R9638 gnd.n7184 gnd.n7183 19.3944
R9639 gnd.n7183 gnd.n508 19.3944
R9640 gnd.n5936 gnd.n508 19.3944
R9641 gnd.n5966 gnd.n5936 19.3944
R9642 gnd.n5966 gnd.n5965 19.3944
R9643 gnd.n5965 gnd.n5964 19.3944
R9644 gnd.n5964 gnd.n5941 19.3944
R9645 gnd.n5960 gnd.n5941 19.3944
R9646 gnd.n5960 gnd.n5959 19.3944
R9647 gnd.n4937 gnd.n4936 18.5761
R9648 gnd.n5711 gnd.n5710 18.5761
R9649 gnd.n7148 gnd.n7147 18.4247
R9650 gnd.n1122 gnd.n1118 18.4247
R9651 gnd.n7506 gnd.n124 18.2308
R9652 gnd.n7187 gnd.n504 18.2308
R9653 gnd.n4731 gnd.n4715 18.2308
R9654 gnd.n4066 gnd.n3661 18.2308
R9655 gnd.n2788 gnd.n2682 18.2305
R9656 gnd.n2788 gnd.n2787 18.2305
R9657 gnd.n2796 gnd.n2671 18.2305
R9658 gnd.n2804 gnd.n2671 18.2305
R9659 gnd.n2804 gnd.n2665 18.2305
R9660 gnd.n2812 gnd.n2665 18.2305
R9661 gnd.n2812 gnd.n2658 18.2305
R9662 gnd.n2850 gnd.n2658 18.2305
R9663 gnd.n2860 gnd.n2591 18.2305
R9664 gnd.n4103 gnd.n3634 18.2305
R9665 gnd.n4111 gnd.n2143 18.2305
R9666 gnd.n4119 gnd.n2143 18.2305
R9667 gnd.n4119 gnd.n2135 18.2305
R9668 gnd.n4127 gnd.n2135 18.2305
R9669 gnd.n4135 gnd.n2126 18.2305
R9670 gnd.n4135 gnd.n2129 18.2305
R9671 gnd.n4143 gnd.n2111 18.2305
R9672 gnd.n4151 gnd.n2111 18.2305
R9673 gnd.n4159 gnd.n2103 18.2305
R9674 gnd.n4167 gnd.n2094 18.2305
R9675 gnd.n4167 gnd.n2097 18.2305
R9676 gnd.n4175 gnd.n2079 18.2305
R9677 gnd.n4183 gnd.n2079 18.2305
R9678 gnd.n4191 gnd.n2071 18.2305
R9679 gnd.n4199 gnd.n2062 18.2305
R9680 gnd.n4199 gnd.n2065 18.2305
R9681 gnd.n4207 gnd.n2047 18.2305
R9682 gnd.n4215 gnd.n2047 18.2305
R9683 gnd.n4223 gnd.n2039 18.2305
R9684 gnd.n4231 gnd.n2029 18.2305
R9685 gnd.n4231 gnd.n2032 18.2305
R9686 gnd.n4239 gnd.n2023 18.2305
R9687 gnd.n4247 gnd.n2006 18.2305
R9688 gnd.n4255 gnd.n2006 18.2305
R9689 gnd.n4273 gnd.n1996 18.2305
R9690 gnd.n4273 gnd.n1999 18.2305
R9691 gnd.n4282 gnd.n979 18.2305
R9692 gnd.t105 gnd.n2039 18.0482
R9693 gnd.n2023 gnd.t53 18.0482
R9694 gnd.t102 gnd.n2071 17.6836
R9695 gnd.t55 gnd.n2103 17.319
R9696 gnd.n3634 gnd.t310 16.2252
R9697 gnd.n4772 gnd.n1898 15.9333
R9698 gnd.n4781 gnd.n1898 15.9333
R9699 gnd.n4783 gnd.n4781 15.9333
R9700 gnd.n4783 gnd.n4782 15.9333
R9701 gnd.n4792 gnd.n1890 15.9333
R9702 gnd.n4792 gnd.n4791 15.9333
R9703 gnd.n4791 gnd.n1892 15.9333
R9704 gnd.n1892 gnd.n1884 15.9333
R9705 gnd.n4800 gnd.n1884 15.9333
R9706 gnd.n4802 gnd.n4800 15.9333
R9707 gnd.n4802 gnd.n4801 15.9333
R9708 gnd.n4801 gnd.n1876 15.9333
R9709 gnd.n4811 gnd.n1876 15.9333
R9710 gnd.n4810 gnd.n1878 15.9333
R9711 gnd.n1878 gnd.n1870 15.9333
R9712 gnd.n4819 gnd.n1870 15.9333
R9713 gnd.n4821 gnd.n4819 15.9333
R9714 gnd.n4821 gnd.n4820 15.9333
R9715 gnd.n4820 gnd.n1862 15.9333
R9716 gnd.n4830 gnd.n1862 15.9333
R9717 gnd.n4830 gnd.n4829 15.9333
R9718 gnd.n1864 gnd.n1856 15.9333
R9719 gnd.n4838 gnd.n1856 15.9333
R9720 gnd.n4840 gnd.n4838 15.9333
R9721 gnd.n4840 gnd.n4839 15.9333
R9722 gnd.n4839 gnd.n1848 15.9333
R9723 gnd.n4849 gnd.n1848 15.9333
R9724 gnd.n4849 gnd.n4848 15.9333
R9725 gnd.n4848 gnd.n1850 15.9333
R9726 gnd.n4857 gnd.n1842 15.9333
R9727 gnd.n4859 gnd.n4857 15.9333
R9728 gnd.n4859 gnd.n4858 15.9333
R9729 gnd.n4858 gnd.n1833 15.9333
R9730 gnd.n4868 gnd.n1833 15.9333
R9731 gnd.n4868 gnd.n4867 15.9333
R9732 gnd.n4867 gnd.n1836 15.9333
R9733 gnd.n1836 gnd.n1835 15.9333
R9734 gnd.n5078 gnd.n4878 15.9333
R9735 gnd.n4912 gnd.n4911 15.9333
R9736 gnd.n5086 gnd.n1767 15.9333
R9737 gnd.n5112 gnd.n1762 15.9333
R9738 gnd.n5122 gnd.n5121 15.9333
R9739 gnd.n1798 gnd.n1734 15.9333
R9740 gnd.n5166 gnd.n5165 15.9333
R9741 gnd.n5231 gnd.n5230 15.9333
R9742 gnd.n5274 gnd.n1644 15.9333
R9743 gnd.n5309 gnd.n1633 15.9333
R9744 gnd.n5325 gnd.n5324 15.9333
R9745 gnd.n5333 gnd.n1618 15.9333
R9746 gnd.n5368 gnd.n1606 15.9333
R9747 gnd.n5377 gnd.n5376 15.9333
R9748 gnd.n5410 gnd.n1576 15.9333
R9749 gnd.n1531 gnd.n1525 15.9333
R9750 gnd.n1517 gnd.n1513 15.9333
R9751 gnd.n5531 gnd.n1494 15.9333
R9752 gnd.n1503 gnd.n1490 15.9333
R9753 gnd.n5547 gnd.n1479 15.9333
R9754 gnd.n5716 gnd.n5715 15.9333
R9755 gnd.n5725 gnd.n5724 15.9333
R9756 gnd.n5735 gnd.n5733 15.9333
R9757 gnd.n5735 gnd.n5734 15.9333
R9758 gnd.n5734 gnd.n1379 15.9333
R9759 gnd.n5744 gnd.n1379 15.9333
R9760 gnd.n5744 gnd.n5743 15.9333
R9761 gnd.n5743 gnd.n1381 15.9333
R9762 gnd.n1381 gnd.n1373 15.9333
R9763 gnd.n5752 gnd.n1373 15.9333
R9764 gnd.n5754 gnd.n5753 15.9333
R9765 gnd.n5753 gnd.n1365 15.9333
R9766 gnd.n5763 gnd.n1365 15.9333
R9767 gnd.n5763 gnd.n5762 15.9333
R9768 gnd.n5762 gnd.n1367 15.9333
R9769 gnd.n1367 gnd.n1359 15.9333
R9770 gnd.n5771 gnd.n1359 15.9333
R9771 gnd.n5773 gnd.n5771 15.9333
R9772 gnd.n5772 gnd.n1351 15.9333
R9773 gnd.n5782 gnd.n1351 15.9333
R9774 gnd.n5782 gnd.n5781 15.9333
R9775 gnd.n5781 gnd.n1353 15.9333
R9776 gnd.n1353 gnd.n1345 15.9333
R9777 gnd.n5790 gnd.n1345 15.9333
R9778 gnd.n5792 gnd.n5790 15.9333
R9779 gnd.n5792 gnd.n5791 15.9333
R9780 gnd.n5801 gnd.n1337 15.9333
R9781 gnd.n5801 gnd.n5800 15.9333
R9782 gnd.n5800 gnd.n1339 15.9333
R9783 gnd.n1339 gnd.n1331 15.9333
R9784 gnd.n5809 gnd.n1331 15.9333
R9785 gnd.n5811 gnd.n5809 15.9333
R9786 gnd.n5811 gnd.n5810 15.9333
R9787 gnd.n5810 gnd.n1322 15.9333
R9788 gnd.n5993 gnd.n1322 15.9333
R9789 gnd.n5992 gnd.n1324 15.9333
R9790 gnd.n1324 gnd.n1315 15.9333
R9791 gnd.n6001 gnd.n1315 15.9333
R9792 gnd.n6001 gnd.n1316 15.9333
R9793 gnd.n3483 gnd.n3481 15.6674
R9794 gnd.n3451 gnd.n3449 15.6674
R9795 gnd.n3419 gnd.n3417 15.6674
R9796 gnd.n3388 gnd.n3386 15.6674
R9797 gnd.n3356 gnd.n3354 15.6674
R9798 gnd.n3324 gnd.n3322 15.6674
R9799 gnd.n3292 gnd.n3290 15.6674
R9800 gnd.n3261 gnd.n3259 15.6674
R9801 gnd.n5156 gnd.n1719 15.296
R9802 gnd.n1713 gnd.n1703 15.296
R9803 gnd.n5194 gnd.t118 15.296
R9804 gnd.n5284 gnd.n1624 15.296
R9805 gnd.n5334 gnd.n1613 15.296
R9806 gnd.n5482 gnd.t94 15.296
R9807 gnd.n5470 gnd.n1540 15.296
R9808 gnd.n5506 gnd.n5505 15.296
R9809 gnd.n1412 gnd.n1411 15.0827
R9810 gnd.n4924 gnd.n4919 15.0481
R9811 gnd.n1422 gnd.n1421 15.0481
R9812 gnd.t110 gnd.n1057 14.9773
R9813 gnd.n1835 gnd.t47 14.9773
R9814 gnd.n5733 gnd.t353 14.9773
R9815 gnd.t27 gnd.n433 14.9773
R9816 gnd.n5088 gnd.n5087 14.6587
R9817 gnd.n1775 gnd.n1684 14.6587
R9818 gnd.n5443 gnd.n1559 14.6587
R9819 gnd.n5568 gnd.n5567 14.6587
R9820 gnd.t2 gnd.n1015 14.34
R9821 gnd.t121 gnd.n399 14.34
R9822 gnd.n2872 gnd.n2592 14.2199
R9823 gnd.n2882 gnd.n2575 14.2199
R9824 gnd.n2578 gnd.n2566 14.2199
R9825 gnd.n2903 gnd.n2567 14.2199
R9826 gnd.n2913 gnd.n2547 14.2199
R9827 gnd.n2923 gnd.n2922 14.2199
R9828 gnd.n2533 gnd.n2531 14.2199
R9829 gnd.n2954 gnd.n2953 14.2199
R9830 gnd.n2969 gnd.n2516 14.2199
R9831 gnd.n3023 gnd.n2455 14.2199
R9832 gnd.n2979 gnd.n2456 14.2199
R9833 gnd.n3016 gnd.n2467 14.2199
R9834 gnd.n2505 gnd.n2504 14.2199
R9835 gnd.n3010 gnd.n3009 14.2199
R9836 gnd.n2491 gnd.n2478 14.2199
R9837 gnd.n3049 gnd.n3048 14.2199
R9838 gnd.n3059 gnd.n2375 14.2199
R9839 gnd.n3071 gnd.n2367 14.2199
R9840 gnd.n3070 gnd.n2355 14.2199
R9841 gnd.n3089 gnd.n3088 14.2199
R9842 gnd.n3099 gnd.n2348 14.2199
R9843 gnd.n3110 gnd.n2336 14.2199
R9844 gnd.n3134 gnd.n3133 14.2199
R9845 gnd.n3145 gnd.n2319 14.2199
R9846 gnd.n3144 gnd.n2321 14.2199
R9847 gnd.n3156 gnd.n2312 14.2199
R9848 gnd.n3174 gnd.n3173 14.2199
R9849 gnd.n2303 gnd.n2292 14.2199
R9850 gnd.n3195 gnd.n2280 14.2199
R9851 gnd.n3223 gnd.n3222 14.2199
R9852 gnd.n3234 gnd.n2265 14.2199
R9853 gnd.n3245 gnd.n2258 14.2199
R9854 gnd.n3244 gnd.n2246 14.2199
R9855 gnd.n3517 gnd.n3516 14.2199
R9856 gnd.n3539 gnd.n2231 14.2199
R9857 gnd.n5130 gnd.t282 14.0214
R9858 gnd.n5148 gnd.n5147 14.0214
R9859 gnd.n5193 gnd.n1698 14.0214
R9860 gnd.n5292 gnd.n5291 14.0214
R9861 gnd.n5367 gnd.n1608 14.0214
R9862 gnd.n5483 gnd.n1544 14.0214
R9863 gnd.n5514 gnd.n1518 14.0214
R9864 gnd.t291 gnd.n1394 14.0214
R9865 gnd.n5266 gnd.t347 13.7027
R9866 gnd.n5389 gnd.t18 13.7027
R9867 gnd.n7110 gnd.n588 13.5763
R9868 gnd.n7558 gnd.n7557 13.5763
R9869 gnd.n2653 gnd.n2652 13.5763
R9870 gnd.n3597 gnd.n2195 13.5763
R9871 gnd.n6189 gnd.n1159 13.5763
R9872 gnd.n3735 gnd.n3734 13.5763
R9873 gnd.n5141 gnd.n5140 13.384
R9874 gnd.n5206 gnd.n1688 13.384
R9875 gnd.t1 gnd.n5204 13.384
R9876 gnd.t130 gnd.n5421 13.384
R9877 gnd.n5451 gnd.n1553 13.384
R9878 gnd.n5532 gnd.n5530 13.384
R9879 gnd.n2893 gnd.t180 13.3084
R9880 gnd.n4127 gnd.t142 13.3084
R9881 gnd.n4935 gnd.n4916 13.1884
R9882 gnd.n4930 gnd.n4929 13.1884
R9883 gnd.n4929 gnd.n4928 13.1884
R9884 gnd.n1415 gnd.n1410 13.1884
R9885 gnd.n1416 gnd.n1415 13.1884
R9886 gnd.n4931 gnd.n4918 13.146
R9887 gnd.n4927 gnd.n4918 13.146
R9888 gnd.n1414 gnd.n1413 13.146
R9889 gnd.n1414 gnd.n1409 13.146
R9890 gnd.n5077 gnd.n4912 13.0654
R9891 gnd.n5576 gnd.t355 13.0654
R9892 gnd.n5724 gnd.n1396 13.0654
R9893 gnd.n2594 gnd.t317 12.9438
R9894 gnd.n4159 gnd.t70 12.9438
R9895 gnd.n3484 gnd.n3480 12.8005
R9896 gnd.n3452 gnd.n3448 12.8005
R9897 gnd.n3420 gnd.n3416 12.8005
R9898 gnd.n3389 gnd.n3385 12.8005
R9899 gnd.n3357 gnd.n3353 12.8005
R9900 gnd.n3325 gnd.n3321 12.8005
R9901 gnd.n3293 gnd.n3289 12.8005
R9902 gnd.n3262 gnd.n3258 12.8005
R9903 gnd.n1808 gnd.n1747 12.7467
R9904 gnd.n5259 gnd.n5258 12.7467
R9905 gnd.n1600 gnd.n1588 12.7467
R9906 gnd.n5561 gnd.n5560 12.7467
R9907 gnd.n4191 gnd.t51 12.5792
R9908 gnd.t133 gnd.n4810 12.4281
R9909 gnd.n5791 gnd.t198 12.4281
R9910 gnd.t74 gnd.n229 12.4281
R9911 gnd.n7106 gnd.n588 12.4126
R9912 gnd.n7557 gnd.n200 12.4126
R9913 gnd.n2652 gnd.n2647 12.4126
R9914 gnd.n3600 gnd.n3597 12.4126
R9915 gnd.n6184 gnd.n1159 12.4126
R9916 gnd.n3868 gnd.n3734 12.4126
R9917 gnd.t8 gnd.n2599 12.2146
R9918 gnd.n4223 gnd.t98 12.2146
R9919 gnd.n4239 gnd.t64 12.2146
R9920 gnd.n5074 gnd.n4937 12.1761
R9921 gnd.n5710 gnd.n5709 12.1761
R9922 gnd.n1799 gnd.n1726 12.1094
R9923 gnd.n5186 gnd.n5185 12.1094
R9924 gnd.n5490 gnd.n1538 12.1094
R9925 gnd.n5522 gnd.n5521 12.1094
R9926 gnd.n3488 gnd.n3487 12.0247
R9927 gnd.n3456 gnd.n3455 12.0247
R9928 gnd.n3424 gnd.n3423 12.0247
R9929 gnd.n3393 gnd.n3392 12.0247
R9930 gnd.n3361 gnd.n3360 12.0247
R9931 gnd.n3329 gnd.n3328 12.0247
R9932 gnd.n3297 gnd.n3296 12.0247
R9933 gnd.n3266 gnd.n3265 12.0247
R9934 gnd.t162 gnd.n2293 11.85
R9935 gnd.n4207 gnd.t140 11.85
R9936 gnd.n4255 gnd.t6 11.85
R9937 gnd.t45 gnd.n260 11.7908
R9938 gnd.t78 gnd.n2328 11.4854
R9939 gnd.n4175 gnd.t4 11.4854
R9940 gnd.n5123 gnd.n1751 11.4721
R9941 gnd.t200 gnd.n1674 11.4721
R9942 gnd.n5223 gnd.n5222 11.4721
R9943 gnd.n5251 gnd.n1658 11.4721
R9944 gnd.n5401 gnd.n1583 11.4721
R9945 gnd.n5433 gnd.n1566 11.4721
R9946 gnd.n5432 gnd.t201 11.4721
R9947 gnd.n5545 gnd.n5543 11.4721
R9948 gnd.n5549 gnd.n1402 11.4721
R9949 gnd.n5714 gnd.t265 11.4721
R9950 gnd.n4533 gnd.t33 11.3031
R9951 gnd.n3491 gnd.n3478 11.249
R9952 gnd.n3459 gnd.n3446 11.249
R9953 gnd.n3427 gnd.n3414 11.249
R9954 gnd.n3396 gnd.n3383 11.249
R9955 gnd.n3364 gnd.n3351 11.249
R9956 gnd.n3332 gnd.n3319 11.249
R9957 gnd.n3300 gnd.n3287 11.249
R9958 gnd.n3269 gnd.n3256 11.249
R9959 gnd.n1850 gnd.t357 11.1535
R9960 gnd.n1690 gnd.t196 11.1535
R9961 gnd.n5420 gnd.t49 11.1535
R9962 gnd.n5754 gnd.t220 11.1535
R9963 gnd.n356 gnd.t41 11.1535
R9964 gnd.t29 gnd.n290 11.1535
R9965 gnd.n3060 gnd.t156 11.1208
R9966 gnd.n4143 gnd.t31 11.1208
R9967 gnd.n5164 gnd.n1721 10.8348
R9968 gnd.n1790 gnd.n1721 10.8348
R9969 gnd.n5299 gnd.n1625 10.8348
R9970 gnd.n5300 gnd.n5299 10.8348
R9971 gnd.n5499 gnd.n5498 10.8348
R9972 gnd.n5498 gnd.n1532 10.8348
R9973 gnd.n3017 gnd.t80 10.7562
R9974 gnd.n3002 gnd.t164 10.7562
R9975 gnd.n5644 gnd.n1452 10.6151
R9976 gnd.n5644 gnd.n5643 10.6151
R9977 gnd.n5641 gnd.n1456 10.6151
R9978 gnd.n5636 gnd.n1456 10.6151
R9979 gnd.n5636 gnd.n5635 10.6151
R9980 gnd.n5635 gnd.n5634 10.6151
R9981 gnd.n5634 gnd.n1459 10.6151
R9982 gnd.n5629 gnd.n1459 10.6151
R9983 gnd.n5629 gnd.n5628 10.6151
R9984 gnd.n5628 gnd.n5627 10.6151
R9985 gnd.n5627 gnd.n1462 10.6151
R9986 gnd.n5622 gnd.n1462 10.6151
R9987 gnd.n5622 gnd.n5621 10.6151
R9988 gnd.n5621 gnd.n5620 10.6151
R9989 gnd.n5620 gnd.n1465 10.6151
R9990 gnd.n5615 gnd.n1465 10.6151
R9991 gnd.n5615 gnd.n5614 10.6151
R9992 gnd.n5614 gnd.n5613 10.6151
R9993 gnd.n5613 gnd.n1468 10.6151
R9994 gnd.n5608 gnd.n1468 10.6151
R9995 gnd.n5608 gnd.n5607 10.6151
R9996 gnd.n5607 gnd.n5606 10.6151
R9997 gnd.n5606 gnd.n1471 10.6151
R9998 gnd.n5601 gnd.n1471 10.6151
R9999 gnd.n5601 gnd.n5600 10.6151
R10000 gnd.n5600 gnd.n5599 10.6151
R10001 gnd.n5599 gnd.n1474 10.6151
R10002 gnd.n5594 gnd.n1474 10.6151
R10003 gnd.n5594 gnd.n5593 10.6151
R10004 gnd.n5593 gnd.n5592 10.6151
R10005 gnd.n4944 gnd.n4943 10.6151
R10006 gnd.n4943 gnd.n1769 10.6151
R10007 gnd.n5102 gnd.n1769 10.6151
R10008 gnd.n5102 gnd.n5101 10.6151
R10009 gnd.n5101 gnd.n5100 10.6151
R10010 gnd.n5100 gnd.n1814 10.6151
R10011 gnd.n1814 gnd.n1813 10.6151
R10012 gnd.n1813 gnd.n1811 10.6151
R10013 gnd.n1811 gnd.n1810 10.6151
R10014 gnd.n1810 gnd.n1806 10.6151
R10015 gnd.n1806 gnd.n1805 10.6151
R10016 gnd.n1805 gnd.n1802 10.6151
R10017 gnd.n1802 gnd.n1801 10.6151
R10018 gnd.n1801 gnd.n1796 10.6151
R10019 gnd.n1796 gnd.n1795 10.6151
R10020 gnd.n1795 gnd.n1793 10.6151
R10021 gnd.n1793 gnd.n1792 10.6151
R10022 gnd.n1792 gnd.n1788 10.6151
R10023 gnd.n1788 gnd.n1787 10.6151
R10024 gnd.n1787 gnd.n1786 10.6151
R10025 gnd.n1786 gnd.n1785 10.6151
R10026 gnd.n1785 gnd.n1784 10.6151
R10027 gnd.n1784 gnd.n1781 10.6151
R10028 gnd.n1781 gnd.n1780 10.6151
R10029 gnd.n1780 gnd.n1778 10.6151
R10030 gnd.n1778 gnd.n1777 10.6151
R10031 gnd.n1777 gnd.n1773 10.6151
R10032 gnd.n1773 gnd.n1772 10.6151
R10033 gnd.n1772 gnd.n1770 10.6151
R10034 gnd.n1770 gnd.n1655 10.6151
R10035 gnd.n5253 gnd.n1655 10.6151
R10036 gnd.n5254 gnd.n5253 10.6151
R10037 gnd.n5255 gnd.n5254 10.6151
R10038 gnd.n5255 gnd.n1642 10.6151
R10039 gnd.n5277 gnd.n1642 10.6151
R10040 gnd.n5278 gnd.n5277 10.6151
R10041 gnd.n5289 gnd.n5278 10.6151
R10042 gnd.n5289 gnd.n5288 10.6151
R10043 gnd.n5288 gnd.n5287 10.6151
R10044 gnd.n5287 gnd.n5279 10.6151
R10045 gnd.n5280 gnd.n5279 10.6151
R10046 gnd.n5280 gnd.n1615 10.6151
R10047 gnd.n5336 gnd.n1615 10.6151
R10048 gnd.n5337 gnd.n5336 10.6151
R10049 gnd.n5354 gnd.n5337 10.6151
R10050 gnd.n5354 gnd.n5353 10.6151
R10051 gnd.n5353 gnd.n5352 10.6151
R10052 gnd.n5352 gnd.n5338 10.6151
R10053 gnd.n5346 gnd.n5338 10.6151
R10054 gnd.n5346 gnd.n5345 10.6151
R10055 gnd.n5345 gnd.n5344 10.6151
R10056 gnd.n5344 gnd.n5343 10.6151
R10057 gnd.n5343 gnd.n5342 10.6151
R10058 gnd.n5342 gnd.n1573 10.6151
R10059 gnd.n5413 gnd.n1573 10.6151
R10060 gnd.n5414 gnd.n5413 10.6151
R10061 gnd.n5416 gnd.n5414 10.6151
R10062 gnd.n5417 gnd.n5416 10.6151
R10063 gnd.n5418 gnd.n5417 10.6151
R10064 gnd.n5418 gnd.n1551 10.6151
R10065 gnd.n5454 gnd.n1551 10.6151
R10066 gnd.n5455 gnd.n5454 10.6151
R10067 gnd.n5457 gnd.n5455 10.6151
R10068 gnd.n5458 gnd.n5457 10.6151
R10069 gnd.n5468 gnd.n5458 10.6151
R10070 gnd.n5468 gnd.n5467 10.6151
R10071 gnd.n5467 gnd.n5466 10.6151
R10072 gnd.n5466 gnd.n5464 10.6151
R10073 gnd.n5464 gnd.n5463 10.6151
R10074 gnd.n5463 gnd.n5461 10.6151
R10075 gnd.n5461 gnd.n5460 10.6151
R10076 gnd.n5460 gnd.n1504 10.6151
R10077 gnd.n5534 gnd.n1504 10.6151
R10078 gnd.n5535 gnd.n5534 10.6151
R10079 gnd.n5537 gnd.n5535 10.6151
R10080 gnd.n5538 gnd.n5537 10.6151
R10081 gnd.n5541 gnd.n5538 10.6151
R10082 gnd.n5541 gnd.n5540 10.6151
R10083 gnd.n5540 gnd.n5539 10.6151
R10084 gnd.n5539 gnd.n1477 10.6151
R10085 gnd.n5586 gnd.n1477 10.6151
R10086 gnd.n5587 gnd.n5586 10.6151
R10087 gnd.n5588 gnd.n5587 10.6151
R10088 gnd.n5009 gnd.n5008 10.6151
R10089 gnd.n5008 gnd.n5005 10.6151
R10090 gnd.n5003 gnd.n5000 10.6151
R10091 gnd.n5000 gnd.n4999 10.6151
R10092 gnd.n4999 gnd.n4996 10.6151
R10093 gnd.n4996 gnd.n4995 10.6151
R10094 gnd.n4995 gnd.n4992 10.6151
R10095 gnd.n4992 gnd.n4991 10.6151
R10096 gnd.n4991 gnd.n4988 10.6151
R10097 gnd.n4988 gnd.n4987 10.6151
R10098 gnd.n4987 gnd.n4984 10.6151
R10099 gnd.n4984 gnd.n4983 10.6151
R10100 gnd.n4983 gnd.n4980 10.6151
R10101 gnd.n4980 gnd.n4979 10.6151
R10102 gnd.n4979 gnd.n4976 10.6151
R10103 gnd.n4976 gnd.n4975 10.6151
R10104 gnd.n4975 gnd.n4972 10.6151
R10105 gnd.n4972 gnd.n4971 10.6151
R10106 gnd.n4971 gnd.n4968 10.6151
R10107 gnd.n4968 gnd.n4967 10.6151
R10108 gnd.n4967 gnd.n4964 10.6151
R10109 gnd.n4964 gnd.n4963 10.6151
R10110 gnd.n4963 gnd.n4960 10.6151
R10111 gnd.n4960 gnd.n4959 10.6151
R10112 gnd.n4959 gnd.n4956 10.6151
R10113 gnd.n4956 gnd.n4955 10.6151
R10114 gnd.n4955 gnd.n4952 10.6151
R10115 gnd.n4952 gnd.n4951 10.6151
R10116 gnd.n4951 gnd.n4948 10.6151
R10117 gnd.n4948 gnd.n4947 10.6151
R10118 gnd.n5074 gnd.n5073 10.6151
R10119 gnd.n5073 gnd.n5072 10.6151
R10120 gnd.n5072 gnd.n5071 10.6151
R10121 gnd.n5071 gnd.n5069 10.6151
R10122 gnd.n5069 gnd.n5066 10.6151
R10123 gnd.n5066 gnd.n5065 10.6151
R10124 gnd.n5065 gnd.n5062 10.6151
R10125 gnd.n5062 gnd.n5061 10.6151
R10126 gnd.n5061 gnd.n5058 10.6151
R10127 gnd.n5058 gnd.n5057 10.6151
R10128 gnd.n5057 gnd.n5054 10.6151
R10129 gnd.n5054 gnd.n5053 10.6151
R10130 gnd.n5053 gnd.n5050 10.6151
R10131 gnd.n5050 gnd.n5049 10.6151
R10132 gnd.n5049 gnd.n5046 10.6151
R10133 gnd.n5046 gnd.n5045 10.6151
R10134 gnd.n5045 gnd.n5042 10.6151
R10135 gnd.n5042 gnd.n5041 10.6151
R10136 gnd.n5041 gnd.n5038 10.6151
R10137 gnd.n5038 gnd.n5037 10.6151
R10138 gnd.n5037 gnd.n5034 10.6151
R10139 gnd.n5034 gnd.n5033 10.6151
R10140 gnd.n5033 gnd.n5030 10.6151
R10141 gnd.n5030 gnd.n5029 10.6151
R10142 gnd.n5029 gnd.n5026 10.6151
R10143 gnd.n5026 gnd.n5025 10.6151
R10144 gnd.n5025 gnd.n5022 10.6151
R10145 gnd.n5022 gnd.n5021 10.6151
R10146 gnd.n5018 gnd.n5017 10.6151
R10147 gnd.n5017 gnd.n5014 10.6151
R10148 gnd.n5709 gnd.n1427 10.6151
R10149 gnd.n1428 gnd.n1427 10.6151
R10150 gnd.n5702 gnd.n1428 10.6151
R10151 gnd.n5702 gnd.n5701 10.6151
R10152 gnd.n5701 gnd.n5700 10.6151
R10153 gnd.n5700 gnd.n1430 10.6151
R10154 gnd.n5695 gnd.n1430 10.6151
R10155 gnd.n5695 gnd.n5694 10.6151
R10156 gnd.n5694 gnd.n5693 10.6151
R10157 gnd.n5693 gnd.n1433 10.6151
R10158 gnd.n5688 gnd.n1433 10.6151
R10159 gnd.n5688 gnd.n5687 10.6151
R10160 gnd.n5687 gnd.n5686 10.6151
R10161 gnd.n5686 gnd.n1436 10.6151
R10162 gnd.n5681 gnd.n1436 10.6151
R10163 gnd.n5681 gnd.n5680 10.6151
R10164 gnd.n5680 gnd.n5679 10.6151
R10165 gnd.n5679 gnd.n1439 10.6151
R10166 gnd.n5674 gnd.n1439 10.6151
R10167 gnd.n5674 gnd.n5673 10.6151
R10168 gnd.n5673 gnd.n5672 10.6151
R10169 gnd.n5672 gnd.n1442 10.6151
R10170 gnd.n5667 gnd.n1442 10.6151
R10171 gnd.n5667 gnd.n5666 10.6151
R10172 gnd.n5666 gnd.n5665 10.6151
R10173 gnd.n5665 gnd.n1445 10.6151
R10174 gnd.n5660 gnd.n1445 10.6151
R10175 gnd.n5660 gnd.n5659 10.6151
R10176 gnd.n5657 gnd.n1450 10.6151
R10177 gnd.n5652 gnd.n1450 10.6151
R10178 gnd.n4936 gnd.n1765 10.6151
R10179 gnd.n5108 gnd.n1765 10.6151
R10180 gnd.n5109 gnd.n5108 10.6151
R10181 gnd.n5110 gnd.n5109 10.6151
R10182 gnd.n5110 gnd.n1749 10.6151
R10183 gnd.n5125 gnd.n1749 10.6151
R10184 gnd.n5126 gnd.n5125 10.6151
R10185 gnd.n5127 gnd.n5126 10.6151
R10186 gnd.n5127 gnd.n1736 10.6151
R10187 gnd.n5143 gnd.n1736 10.6151
R10188 gnd.n5144 gnd.n5143 10.6151
R10189 gnd.n5145 gnd.n5144 10.6151
R10190 gnd.n5145 gnd.n1724 10.6151
R10191 gnd.n5159 gnd.n1724 10.6151
R10192 gnd.n5160 gnd.n5159 10.6151
R10193 gnd.n5162 gnd.n5160 10.6151
R10194 gnd.n5162 gnd.n5161 10.6151
R10195 gnd.n5161 gnd.n1700 10.6151
R10196 gnd.n5189 gnd.n1700 10.6151
R10197 gnd.n5190 gnd.n5189 10.6151
R10198 gnd.n5191 gnd.n5190 10.6151
R10199 gnd.n5191 gnd.n1686 10.6151
R10200 gnd.n5208 gnd.n1686 10.6151
R10201 gnd.n5209 gnd.n5208 10.6151
R10202 gnd.n5210 gnd.n5209 10.6151
R10203 gnd.n5210 gnd.n1672 10.6151
R10204 gnd.n5225 gnd.n1672 10.6151
R10205 gnd.n5226 gnd.n5225 10.6151
R10206 gnd.n5228 gnd.n5226 10.6151
R10207 gnd.n5228 gnd.n5227 10.6151
R10208 gnd.n5227 gnd.n1653 10.6151
R10209 gnd.n5263 gnd.n1653 10.6151
R10210 gnd.n5263 gnd.n5262 10.6151
R10211 gnd.n5262 gnd.n5261 10.6151
R10212 gnd.n5261 gnd.n1637 10.6151
R10213 gnd.n5295 gnd.n1637 10.6151
R10214 gnd.n5296 gnd.n5295 10.6151
R10215 gnd.n5306 gnd.n5296 10.6151
R10216 gnd.n5306 gnd.n5305 10.6151
R10217 gnd.n5305 gnd.n5304 10.6151
R10218 gnd.n5304 gnd.n5297 10.6151
R10219 gnd.n5298 gnd.n5297 10.6151
R10220 gnd.n5298 gnd.n1611 10.6151
R10221 gnd.n5360 gnd.n1611 10.6151
R10222 gnd.n5361 gnd.n5360 10.6151
R10223 gnd.n5365 gnd.n5361 10.6151
R10224 gnd.n5365 gnd.n5364 10.6151
R10225 gnd.n5364 gnd.n5363 10.6151
R10226 gnd.n5363 gnd.n1586 10.6151
R10227 gnd.n5394 gnd.n1586 10.6151
R10228 gnd.n5395 gnd.n5394 10.6151
R10229 gnd.n5399 gnd.n5395 10.6151
R10230 gnd.n5399 gnd.n5398 10.6151
R10231 gnd.n5398 gnd.n5397 10.6151
R10232 gnd.n5397 gnd.n1564 10.6151
R10233 gnd.n5435 gnd.n1564 10.6151
R10234 gnd.n5436 gnd.n5435 10.6151
R10235 gnd.n5440 gnd.n5436 10.6151
R10236 gnd.n5440 gnd.n5439 10.6151
R10237 gnd.n5439 gnd.n5438 10.6151
R10238 gnd.n5438 gnd.n1542 10.6151
R10239 gnd.n5485 gnd.n1542 10.6151
R10240 gnd.n5486 gnd.n5485 10.6151
R10241 gnd.n5487 gnd.n5486 10.6151
R10242 gnd.n5487 gnd.n1528 10.6151
R10243 gnd.n5501 gnd.n1528 10.6151
R10244 gnd.n5502 gnd.n5501 10.6151
R10245 gnd.n5503 gnd.n5502 10.6151
R10246 gnd.n5503 gnd.n1516 10.6151
R10247 gnd.n5519 gnd.n1516 10.6151
R10248 gnd.n5519 gnd.n5518 10.6151
R10249 gnd.n5518 gnd.n5517 10.6151
R10250 gnd.n5517 gnd.n1492 10.6151
R10251 gnd.n5563 gnd.n1492 10.6151
R10252 gnd.n5564 gnd.n5563 10.6151
R10253 gnd.n5565 gnd.n5564 10.6151
R10254 gnd.n5565 gnd.n1481 10.6151
R10255 gnd.n5579 gnd.n1481 10.6151
R10256 gnd.n5580 gnd.n5579 10.6151
R10257 gnd.n5581 gnd.n5580 10.6151
R10258 gnd.n5581 gnd.n1407 10.6151
R10259 gnd.n5712 gnd.n1407 10.6151
R10260 gnd.n5712 gnd.n5711 10.6151
R10261 gnd.n2861 gnd.n2860 10.5739
R10262 gnd.n5175 gnd.t224 10.5161
R10263 gnd.n5473 gnd.t131 10.5161
R10264 gnd.t12 gnd.n320 10.5161
R10265 gnd.n323 gnd.t10 10.5161
R10266 gnd.n3492 gnd.n3476 10.4732
R10267 gnd.n3460 gnd.n3444 10.4732
R10268 gnd.n3428 gnd.n3412 10.4732
R10269 gnd.n3397 gnd.n3381 10.4732
R10270 gnd.n3365 gnd.n3349 10.4732
R10271 gnd.n3333 gnd.n3317 10.4732
R10272 gnd.n3301 gnd.n3285 10.4732
R10273 gnd.n3270 gnd.n3254 10.4732
R10274 gnd.t163 gnd.n2541 10.3916
R10275 gnd.n5105 gnd.n5104 10.1975
R10276 gnd.n5098 gnd.n1751 10.1975
R10277 gnd.n5222 gnd.n1665 10.1975
R10278 gnd.n1670 gnd.n1658 10.1975
R10279 gnd.n5340 gnd.n1583 10.1975
R10280 gnd.n5411 gnd.n1566 10.1975
R10281 gnd.n2569 gnd.t82 10.027
R10282 gnd.t333 gnd.t92 9.87883
R10283 gnd.t72 gnd.n353 9.87883
R10284 gnd.n293 gnd.t100 9.87883
R10285 gnd.n7683 gnd.n78 9.81789
R10286 gnd.n3496 gnd.n3495 9.69747
R10287 gnd.n3464 gnd.n3463 9.69747
R10288 gnd.n3432 gnd.n3431 9.69747
R10289 gnd.n3401 gnd.n3400 9.69747
R10290 gnd.n3369 gnd.n3368 9.69747
R10291 gnd.n3337 gnd.n3336 9.69747
R10292 gnd.n3305 gnd.n3304 9.69747
R10293 gnd.n3274 gnd.n3273 9.69747
R10294 gnd.n2968 gnd.t157 9.66242
R10295 gnd.n5157 gnd.n1726 9.56018
R10296 gnd.n5187 gnd.n5186 9.56018
R10297 gnd.n1669 gnd.t95 9.56018
R10298 gnd.n5285 gnd.n5283 9.56018
R10299 gnd.n5358 gnd.n5357 9.56018
R10300 gnd.n5339 gnd.t23 9.56018
R10301 gnd.n5490 gnd.n5489 9.56018
R10302 gnd.n5522 gnd.n1511 9.56018
R10303 gnd.n4658 gnd.n4657 9.45751
R10304 gnd.n7229 gnd.n7228 9.45599
R10305 gnd.n3502 gnd.n3501 9.45567
R10306 gnd.n3470 gnd.n3469 9.45567
R10307 gnd.n3438 gnd.n3437 9.45567
R10308 gnd.n3407 gnd.n3406 9.45567
R10309 gnd.n3375 gnd.n3374 9.45567
R10310 gnd.n3343 gnd.n3342 9.45567
R10311 gnd.n3311 gnd.n3310 9.45567
R10312 gnd.n3280 gnd.n3279 9.45567
R10313 gnd.n2448 gnd.n2447 9.39724
R10314 gnd.n7623 gnd.n134 9.3005
R10315 gnd.n7622 gnd.n136 9.3005
R10316 gnd.n140 gnd.n137 9.3005
R10317 gnd.n7617 gnd.n141 9.3005
R10318 gnd.n7616 gnd.n142 9.3005
R10319 gnd.n7615 gnd.n143 9.3005
R10320 gnd.n147 gnd.n144 9.3005
R10321 gnd.n7610 gnd.n148 9.3005
R10322 gnd.n7609 gnd.n149 9.3005
R10323 gnd.n7608 gnd.n150 9.3005
R10324 gnd.n154 gnd.n151 9.3005
R10325 gnd.n7603 gnd.n155 9.3005
R10326 gnd.n7602 gnd.n156 9.3005
R10327 gnd.n7601 gnd.n157 9.3005
R10328 gnd.n161 gnd.n158 9.3005
R10329 gnd.n7596 gnd.n162 9.3005
R10330 gnd.n7595 gnd.n163 9.3005
R10331 gnd.n7591 gnd.n164 9.3005
R10332 gnd.n168 gnd.n165 9.3005
R10333 gnd.n7586 gnd.n169 9.3005
R10334 gnd.n7585 gnd.n170 9.3005
R10335 gnd.n7584 gnd.n171 9.3005
R10336 gnd.n175 gnd.n172 9.3005
R10337 gnd.n7579 gnd.n176 9.3005
R10338 gnd.n7578 gnd.n177 9.3005
R10339 gnd.n7577 gnd.n178 9.3005
R10340 gnd.n182 gnd.n179 9.3005
R10341 gnd.n7572 gnd.n183 9.3005
R10342 gnd.n7571 gnd.n184 9.3005
R10343 gnd.n7570 gnd.n185 9.3005
R10344 gnd.n189 gnd.n186 9.3005
R10345 gnd.n7565 gnd.n190 9.3005
R10346 gnd.n7564 gnd.n191 9.3005
R10347 gnd.n7563 gnd.n192 9.3005
R10348 gnd.n196 gnd.n193 9.3005
R10349 gnd.n7558 gnd.n197 9.3005
R10350 gnd.n7557 gnd.n7556 9.3005
R10351 gnd.n7555 gnd.n200 9.3005
R10352 gnd.n7625 gnd.n7624 9.3005
R10353 gnd.n7102 gnd.n589 9.3005
R10354 gnd.n7101 gnd.n591 9.3005
R10355 gnd.n7100 gnd.n592 9.3005
R10356 gnd.n5864 gnd.n593 9.3005
R10357 gnd.n5868 gnd.n5865 9.3005
R10358 gnd.n5869 gnd.n5863 9.3005
R10359 gnd.n5873 gnd.n5872 9.3005
R10360 gnd.n5874 gnd.n5862 9.3005
R10361 gnd.n5915 gnd.n5875 9.3005
R10362 gnd.n5914 gnd.n5876 9.3005
R10363 gnd.n5913 gnd.n5877 9.3005
R10364 gnd.n5910 gnd.n5878 9.3005
R10365 gnd.n5909 gnd.n5879 9.3005
R10366 gnd.n5885 gnd.n5880 9.3005
R10367 gnd.n5884 gnd.n5881 9.3005
R10368 gnd.n613 gnd.n612 9.3005
R10369 gnd.n6931 gnd.n6930 9.3005
R10370 gnd.n6932 gnd.n611 9.3005
R10371 gnd.n7038 gnd.n6933 9.3005
R10372 gnd.n7037 gnd.n6934 9.3005
R10373 gnd.n7036 gnd.n6935 9.3005
R10374 gnd.n7034 gnd.n6936 9.3005
R10375 gnd.n7033 gnd.n6937 9.3005
R10376 gnd.n7031 gnd.n6938 9.3005
R10377 gnd.n7030 gnd.n6939 9.3005
R10378 gnd.n7028 gnd.n6940 9.3005
R10379 gnd.n7027 gnd.n6941 9.3005
R10380 gnd.n7025 gnd.n6942 9.3005
R10381 gnd.n7024 gnd.n6943 9.3005
R10382 gnd.n7022 gnd.n6944 9.3005
R10383 gnd.n7021 gnd.n6945 9.3005
R10384 gnd.n7019 gnd.n326 9.3005
R10385 gnd.n7018 gnd.n6946 9.3005
R10386 gnd.n7016 gnd.n6947 9.3005
R10387 gnd.n7015 gnd.n6948 9.3005
R10388 gnd.n7013 gnd.n6949 9.3005
R10389 gnd.n7012 gnd.n6950 9.3005
R10390 gnd.n7010 gnd.n6951 9.3005
R10391 gnd.n7009 gnd.n6952 9.3005
R10392 gnd.n7007 gnd.n6953 9.3005
R10393 gnd.n7006 gnd.n6954 9.3005
R10394 gnd.n7004 gnd.n6955 9.3005
R10395 gnd.n7003 gnd.n6956 9.3005
R10396 gnd.n7001 gnd.n6957 9.3005
R10397 gnd.n7000 gnd.n6958 9.3005
R10398 gnd.n6998 gnd.n6959 9.3005
R10399 gnd.n6997 gnd.n6960 9.3005
R10400 gnd.n6995 gnd.n6961 9.3005
R10401 gnd.n6994 gnd.n6962 9.3005
R10402 gnd.n6992 gnd.n6963 9.3005
R10403 gnd.n6991 gnd.n6964 9.3005
R10404 gnd.n6989 gnd.n6965 9.3005
R10405 gnd.n6988 gnd.n6966 9.3005
R10406 gnd.n6986 gnd.n6967 9.3005
R10407 gnd.n6985 gnd.n6968 9.3005
R10408 gnd.n6983 gnd.n6969 9.3005
R10409 gnd.n6982 gnd.n6970 9.3005
R10410 gnd.n6980 gnd.n6971 9.3005
R10411 gnd.n6979 gnd.n6972 9.3005
R10412 gnd.n6977 gnd.n6973 9.3005
R10413 gnd.n6976 gnd.n6975 9.3005
R10414 gnd.n6974 gnd.n204 9.3005
R10415 gnd.n7552 gnd.n203 9.3005
R10416 gnd.n7554 gnd.n7553 9.3005
R10417 gnd.n7104 gnd.n7103 9.3005
R10418 gnd.n7110 gnd.n7109 9.3005
R10419 gnd.n7111 gnd.n583 9.3005
R10420 gnd.n7114 gnd.n582 9.3005
R10421 gnd.n7115 gnd.n581 9.3005
R10422 gnd.n7118 gnd.n580 9.3005
R10423 gnd.n7119 gnd.n579 9.3005
R10424 gnd.n7122 gnd.n578 9.3005
R10425 gnd.n7123 gnd.n577 9.3005
R10426 gnd.n7126 gnd.n576 9.3005
R10427 gnd.n7127 gnd.n575 9.3005
R10428 gnd.n7130 gnd.n574 9.3005
R10429 gnd.n7131 gnd.n573 9.3005
R10430 gnd.n7134 gnd.n572 9.3005
R10431 gnd.n7135 gnd.n571 9.3005
R10432 gnd.n7138 gnd.n570 9.3005
R10433 gnd.n7139 gnd.n569 9.3005
R10434 gnd.n7142 gnd.n568 9.3005
R10435 gnd.n7143 gnd.n567 9.3005
R10436 gnd.n7146 gnd.n566 9.3005
R10437 gnd.n7148 gnd.n560 9.3005
R10438 gnd.n7151 gnd.n559 9.3005
R10439 gnd.n7152 gnd.n558 9.3005
R10440 gnd.n7155 gnd.n557 9.3005
R10441 gnd.n7156 gnd.n556 9.3005
R10442 gnd.n7159 gnd.n555 9.3005
R10443 gnd.n7160 gnd.n554 9.3005
R10444 gnd.n7163 gnd.n553 9.3005
R10445 gnd.n7164 gnd.n552 9.3005
R10446 gnd.n7167 gnd.n551 9.3005
R10447 gnd.n7168 gnd.n550 9.3005
R10448 gnd.n7171 gnd.n549 9.3005
R10449 gnd.n7173 gnd.n548 9.3005
R10450 gnd.n7174 gnd.n547 9.3005
R10451 gnd.n7175 gnd.n546 9.3005
R10452 gnd.n545 gnd.n453 9.3005
R10453 gnd.n7108 gnd.n588 9.3005
R10454 gnd.n7107 gnd.n7106 9.3005
R10455 gnd.n7237 gnd.n452 9.3005
R10456 gnd.n7239 gnd.n7238 9.3005
R10457 gnd.n437 gnd.n436 9.3005
R10458 gnd.n7252 gnd.n7251 9.3005
R10459 gnd.n7253 gnd.n435 9.3005
R10460 gnd.n7255 gnd.n7254 9.3005
R10461 gnd.n419 gnd.n418 9.3005
R10462 gnd.n7268 gnd.n7267 9.3005
R10463 gnd.n7269 gnd.n417 9.3005
R10464 gnd.n7271 gnd.n7270 9.3005
R10465 gnd.n403 gnd.n402 9.3005
R10466 gnd.n7284 gnd.n7283 9.3005
R10467 gnd.n7285 gnd.n401 9.3005
R10468 gnd.n7287 gnd.n7286 9.3005
R10469 gnd.n385 gnd.n384 9.3005
R10470 gnd.n7300 gnd.n7299 9.3005
R10471 gnd.n7301 gnd.n383 9.3005
R10472 gnd.n7303 gnd.n7302 9.3005
R10473 gnd.n369 gnd.n368 9.3005
R10474 gnd.n7316 gnd.n7315 9.3005
R10475 gnd.n7317 gnd.n367 9.3005
R10476 gnd.n7319 gnd.n7318 9.3005
R10477 gnd.n351 gnd.n350 9.3005
R10478 gnd.n7332 gnd.n7331 9.3005
R10479 gnd.n7333 gnd.n349 9.3005
R10480 gnd.n7335 gnd.n7334 9.3005
R10481 gnd.n336 gnd.n335 9.3005
R10482 gnd.n7348 gnd.n7347 9.3005
R10483 gnd.n7349 gnd.n334 9.3005
R10484 gnd.n7351 gnd.n7350 9.3005
R10485 gnd.n318 gnd.n317 9.3005
R10486 gnd.n7364 gnd.n7363 9.3005
R10487 gnd.n7365 gnd.n316 9.3005
R10488 gnd.n7367 gnd.n7366 9.3005
R10489 gnd.n304 gnd.n303 9.3005
R10490 gnd.n7380 gnd.n7379 9.3005
R10491 gnd.n7381 gnd.n302 9.3005
R10492 gnd.n7383 gnd.n7382 9.3005
R10493 gnd.n288 gnd.n287 9.3005
R10494 gnd.n7396 gnd.n7395 9.3005
R10495 gnd.n7397 gnd.n286 9.3005
R10496 gnd.n7399 gnd.n7398 9.3005
R10497 gnd.n274 gnd.n273 9.3005
R10498 gnd.n7412 gnd.n7411 9.3005
R10499 gnd.n7413 gnd.n272 9.3005
R10500 gnd.n7415 gnd.n7414 9.3005
R10501 gnd.n258 gnd.n257 9.3005
R10502 gnd.n7428 gnd.n7427 9.3005
R10503 gnd.n7429 gnd.n256 9.3005
R10504 gnd.n7431 gnd.n7430 9.3005
R10505 gnd.n243 gnd.n242 9.3005
R10506 gnd.n7444 gnd.n7443 9.3005
R10507 gnd.n7445 gnd.n241 9.3005
R10508 gnd.n7447 gnd.n7446 9.3005
R10509 gnd.n227 gnd.n226 9.3005
R10510 gnd.n7460 gnd.n7459 9.3005
R10511 gnd.n7461 gnd.n225 9.3005
R10512 gnd.n7463 gnd.n7462 9.3005
R10513 gnd.n211 gnd.n210 9.3005
R10514 gnd.n7544 gnd.n7543 9.3005
R10515 gnd.n7545 gnd.n209 9.3005
R10516 gnd.n7547 gnd.n7546 9.3005
R10517 gnd.n133 gnd.n132 9.3005
R10518 gnd.n7627 gnd.n7626 9.3005
R10519 gnd.n7236 gnd.n7235 9.3005
R10520 gnd.n977 gnd.n976 9.3005
R10521 gnd.n6322 gnd.n6321 9.3005
R10522 gnd.n6323 gnd.n975 9.3005
R10523 gnd.n6325 gnd.n6324 9.3005
R10524 gnd.n971 gnd.n970 9.3005
R10525 gnd.n6332 gnd.n6331 9.3005
R10526 gnd.n6333 gnd.n969 9.3005
R10527 gnd.n6335 gnd.n6334 9.3005
R10528 gnd.n965 gnd.n964 9.3005
R10529 gnd.n6342 gnd.n6341 9.3005
R10530 gnd.n6343 gnd.n963 9.3005
R10531 gnd.n6345 gnd.n6344 9.3005
R10532 gnd.n959 gnd.n958 9.3005
R10533 gnd.n6352 gnd.n6351 9.3005
R10534 gnd.n6353 gnd.n957 9.3005
R10535 gnd.n6355 gnd.n6354 9.3005
R10536 gnd.n953 gnd.n952 9.3005
R10537 gnd.n6362 gnd.n6361 9.3005
R10538 gnd.n6363 gnd.n951 9.3005
R10539 gnd.n6365 gnd.n6364 9.3005
R10540 gnd.n947 gnd.n946 9.3005
R10541 gnd.n6372 gnd.n6371 9.3005
R10542 gnd.n6373 gnd.n945 9.3005
R10543 gnd.n6375 gnd.n6374 9.3005
R10544 gnd.n941 gnd.n940 9.3005
R10545 gnd.n6382 gnd.n6381 9.3005
R10546 gnd.n6383 gnd.n939 9.3005
R10547 gnd.n6385 gnd.n6384 9.3005
R10548 gnd.n935 gnd.n934 9.3005
R10549 gnd.n6392 gnd.n6391 9.3005
R10550 gnd.n6393 gnd.n933 9.3005
R10551 gnd.n6395 gnd.n6394 9.3005
R10552 gnd.n929 gnd.n928 9.3005
R10553 gnd.n6402 gnd.n6401 9.3005
R10554 gnd.n6403 gnd.n927 9.3005
R10555 gnd.n6405 gnd.n6404 9.3005
R10556 gnd.n923 gnd.n922 9.3005
R10557 gnd.n6412 gnd.n6411 9.3005
R10558 gnd.n6413 gnd.n921 9.3005
R10559 gnd.n6415 gnd.n6414 9.3005
R10560 gnd.n917 gnd.n916 9.3005
R10561 gnd.n6422 gnd.n6421 9.3005
R10562 gnd.n6423 gnd.n915 9.3005
R10563 gnd.n6425 gnd.n6424 9.3005
R10564 gnd.n911 gnd.n910 9.3005
R10565 gnd.n6432 gnd.n6431 9.3005
R10566 gnd.n6433 gnd.n909 9.3005
R10567 gnd.n6435 gnd.n6434 9.3005
R10568 gnd.n905 gnd.n904 9.3005
R10569 gnd.n6442 gnd.n6441 9.3005
R10570 gnd.n6443 gnd.n903 9.3005
R10571 gnd.n6445 gnd.n6444 9.3005
R10572 gnd.n899 gnd.n898 9.3005
R10573 gnd.n6452 gnd.n6451 9.3005
R10574 gnd.n6453 gnd.n897 9.3005
R10575 gnd.n6455 gnd.n6454 9.3005
R10576 gnd.n893 gnd.n892 9.3005
R10577 gnd.n6462 gnd.n6461 9.3005
R10578 gnd.n6463 gnd.n891 9.3005
R10579 gnd.n6465 gnd.n6464 9.3005
R10580 gnd.n887 gnd.n886 9.3005
R10581 gnd.n6472 gnd.n6471 9.3005
R10582 gnd.n6473 gnd.n885 9.3005
R10583 gnd.n6475 gnd.n6474 9.3005
R10584 gnd.n881 gnd.n880 9.3005
R10585 gnd.n6482 gnd.n6481 9.3005
R10586 gnd.n6483 gnd.n879 9.3005
R10587 gnd.n6485 gnd.n6484 9.3005
R10588 gnd.n875 gnd.n874 9.3005
R10589 gnd.n6492 gnd.n6491 9.3005
R10590 gnd.n6493 gnd.n873 9.3005
R10591 gnd.n6495 gnd.n6494 9.3005
R10592 gnd.n869 gnd.n868 9.3005
R10593 gnd.n6502 gnd.n6501 9.3005
R10594 gnd.n6503 gnd.n867 9.3005
R10595 gnd.n6505 gnd.n6504 9.3005
R10596 gnd.n863 gnd.n862 9.3005
R10597 gnd.n6512 gnd.n6511 9.3005
R10598 gnd.n6513 gnd.n861 9.3005
R10599 gnd.n6515 gnd.n6514 9.3005
R10600 gnd.n857 gnd.n856 9.3005
R10601 gnd.n6522 gnd.n6521 9.3005
R10602 gnd.n6523 gnd.n855 9.3005
R10603 gnd.n6525 gnd.n6524 9.3005
R10604 gnd.n851 gnd.n850 9.3005
R10605 gnd.n6532 gnd.n6531 9.3005
R10606 gnd.n6533 gnd.n849 9.3005
R10607 gnd.n6535 gnd.n6534 9.3005
R10608 gnd.n845 gnd.n844 9.3005
R10609 gnd.n6542 gnd.n6541 9.3005
R10610 gnd.n6543 gnd.n843 9.3005
R10611 gnd.n6545 gnd.n6544 9.3005
R10612 gnd.n839 gnd.n838 9.3005
R10613 gnd.n6552 gnd.n6551 9.3005
R10614 gnd.n6553 gnd.n837 9.3005
R10615 gnd.n6555 gnd.n6554 9.3005
R10616 gnd.n833 gnd.n832 9.3005
R10617 gnd.n6562 gnd.n6561 9.3005
R10618 gnd.n6563 gnd.n831 9.3005
R10619 gnd.n6565 gnd.n6564 9.3005
R10620 gnd.n827 gnd.n826 9.3005
R10621 gnd.n6572 gnd.n6571 9.3005
R10622 gnd.n6573 gnd.n825 9.3005
R10623 gnd.n6575 gnd.n6574 9.3005
R10624 gnd.n821 gnd.n820 9.3005
R10625 gnd.n6582 gnd.n6581 9.3005
R10626 gnd.n6583 gnd.n819 9.3005
R10627 gnd.n6585 gnd.n6584 9.3005
R10628 gnd.n815 gnd.n814 9.3005
R10629 gnd.n6592 gnd.n6591 9.3005
R10630 gnd.n6593 gnd.n813 9.3005
R10631 gnd.n6595 gnd.n6594 9.3005
R10632 gnd.n809 gnd.n808 9.3005
R10633 gnd.n6602 gnd.n6601 9.3005
R10634 gnd.n6603 gnd.n807 9.3005
R10635 gnd.n6605 gnd.n6604 9.3005
R10636 gnd.n803 gnd.n802 9.3005
R10637 gnd.n6612 gnd.n6611 9.3005
R10638 gnd.n6613 gnd.n801 9.3005
R10639 gnd.n6615 gnd.n6614 9.3005
R10640 gnd.n797 gnd.n796 9.3005
R10641 gnd.n6622 gnd.n6621 9.3005
R10642 gnd.n6623 gnd.n795 9.3005
R10643 gnd.n6625 gnd.n6624 9.3005
R10644 gnd.n791 gnd.n790 9.3005
R10645 gnd.n6632 gnd.n6631 9.3005
R10646 gnd.n6633 gnd.n789 9.3005
R10647 gnd.n6635 gnd.n6634 9.3005
R10648 gnd.n785 gnd.n784 9.3005
R10649 gnd.n6642 gnd.n6641 9.3005
R10650 gnd.n6643 gnd.n783 9.3005
R10651 gnd.n6645 gnd.n6644 9.3005
R10652 gnd.n779 gnd.n778 9.3005
R10653 gnd.n6652 gnd.n6651 9.3005
R10654 gnd.n6653 gnd.n777 9.3005
R10655 gnd.n6655 gnd.n6654 9.3005
R10656 gnd.n773 gnd.n772 9.3005
R10657 gnd.n6662 gnd.n6661 9.3005
R10658 gnd.n6663 gnd.n771 9.3005
R10659 gnd.n6665 gnd.n6664 9.3005
R10660 gnd.n767 gnd.n766 9.3005
R10661 gnd.n6672 gnd.n6671 9.3005
R10662 gnd.n6673 gnd.n765 9.3005
R10663 gnd.n6675 gnd.n6674 9.3005
R10664 gnd.n761 gnd.n760 9.3005
R10665 gnd.n6682 gnd.n6681 9.3005
R10666 gnd.n6683 gnd.n759 9.3005
R10667 gnd.n6685 gnd.n6684 9.3005
R10668 gnd.n755 gnd.n754 9.3005
R10669 gnd.n6692 gnd.n6691 9.3005
R10670 gnd.n6693 gnd.n753 9.3005
R10671 gnd.n6696 gnd.n6695 9.3005
R10672 gnd.n6694 gnd.n749 9.3005
R10673 gnd.n6702 gnd.n748 9.3005
R10674 gnd.n6704 gnd.n6703 9.3005
R10675 gnd.n744 gnd.n743 9.3005
R10676 gnd.n6713 gnd.n6712 9.3005
R10677 gnd.n6714 gnd.n742 9.3005
R10678 gnd.n6716 gnd.n6715 9.3005
R10679 gnd.n738 gnd.n737 9.3005
R10680 gnd.n6723 gnd.n6722 9.3005
R10681 gnd.n6724 gnd.n736 9.3005
R10682 gnd.n6726 gnd.n6725 9.3005
R10683 gnd.n732 gnd.n731 9.3005
R10684 gnd.n6733 gnd.n6732 9.3005
R10685 gnd.n6734 gnd.n730 9.3005
R10686 gnd.n6736 gnd.n6735 9.3005
R10687 gnd.n726 gnd.n725 9.3005
R10688 gnd.n6743 gnd.n6742 9.3005
R10689 gnd.n6744 gnd.n724 9.3005
R10690 gnd.n6746 gnd.n6745 9.3005
R10691 gnd.n720 gnd.n719 9.3005
R10692 gnd.n6753 gnd.n6752 9.3005
R10693 gnd.n6754 gnd.n718 9.3005
R10694 gnd.n6756 gnd.n6755 9.3005
R10695 gnd.n714 gnd.n713 9.3005
R10696 gnd.n6763 gnd.n6762 9.3005
R10697 gnd.n6764 gnd.n712 9.3005
R10698 gnd.n6766 gnd.n6765 9.3005
R10699 gnd.n708 gnd.n707 9.3005
R10700 gnd.n6773 gnd.n6772 9.3005
R10701 gnd.n6774 gnd.n706 9.3005
R10702 gnd.n6776 gnd.n6775 9.3005
R10703 gnd.n702 gnd.n701 9.3005
R10704 gnd.n6783 gnd.n6782 9.3005
R10705 gnd.n6784 gnd.n700 9.3005
R10706 gnd.n6786 gnd.n6785 9.3005
R10707 gnd.n696 gnd.n695 9.3005
R10708 gnd.n6793 gnd.n6792 9.3005
R10709 gnd.n6794 gnd.n694 9.3005
R10710 gnd.n6796 gnd.n6795 9.3005
R10711 gnd.n690 gnd.n689 9.3005
R10712 gnd.n6803 gnd.n6802 9.3005
R10713 gnd.n6804 gnd.n688 9.3005
R10714 gnd.n6806 gnd.n6805 9.3005
R10715 gnd.n684 gnd.n683 9.3005
R10716 gnd.n6813 gnd.n6812 9.3005
R10717 gnd.n6814 gnd.n682 9.3005
R10718 gnd.n6816 gnd.n6815 9.3005
R10719 gnd.n678 gnd.n677 9.3005
R10720 gnd.n6823 gnd.n6822 9.3005
R10721 gnd.n6824 gnd.n676 9.3005
R10722 gnd.n6826 gnd.n6825 9.3005
R10723 gnd.n672 gnd.n671 9.3005
R10724 gnd.n6833 gnd.n6832 9.3005
R10725 gnd.n6834 gnd.n670 9.3005
R10726 gnd.n6836 gnd.n6835 9.3005
R10727 gnd.n666 gnd.n665 9.3005
R10728 gnd.n6843 gnd.n6842 9.3005
R10729 gnd.n6844 gnd.n664 9.3005
R10730 gnd.n6846 gnd.n6845 9.3005
R10731 gnd.n660 gnd.n659 9.3005
R10732 gnd.n6853 gnd.n6852 9.3005
R10733 gnd.n6854 gnd.n658 9.3005
R10734 gnd.n6856 gnd.n6855 9.3005
R10735 gnd.n654 gnd.n653 9.3005
R10736 gnd.n6863 gnd.n6862 9.3005
R10737 gnd.n6864 gnd.n652 9.3005
R10738 gnd.n6866 gnd.n6865 9.3005
R10739 gnd.n648 gnd.n647 9.3005
R10740 gnd.n6873 gnd.n6872 9.3005
R10741 gnd.n6874 gnd.n646 9.3005
R10742 gnd.n6876 gnd.n6875 9.3005
R10743 gnd.n642 gnd.n641 9.3005
R10744 gnd.n6883 gnd.n6882 9.3005
R10745 gnd.n6884 gnd.n640 9.3005
R10746 gnd.n6886 gnd.n6885 9.3005
R10747 gnd.n636 gnd.n635 9.3005
R10748 gnd.n6893 gnd.n6892 9.3005
R10749 gnd.n6894 gnd.n634 9.3005
R10750 gnd.n6896 gnd.n6895 9.3005
R10751 gnd.n630 gnd.n629 9.3005
R10752 gnd.n6903 gnd.n6902 9.3005
R10753 gnd.n6904 gnd.n628 9.3005
R10754 gnd.n6906 gnd.n6905 9.3005
R10755 gnd.n624 gnd.n623 9.3005
R10756 gnd.n6914 gnd.n6913 9.3005
R10757 gnd.n6915 gnd.n622 9.3005
R10758 gnd.n6918 gnd.n6917 9.3005
R10759 gnd.n6706 gnd.n6705 9.3005
R10760 gnd.n4540 gnd.n1944 9.3005
R10761 gnd.n4544 gnd.n4543 9.3005
R10762 gnd.n4545 gnd.n1943 9.3005
R10763 gnd.n4547 gnd.n4546 9.3005
R10764 gnd.n1941 gnd.n1940 9.3005
R10765 gnd.n4552 gnd.n4551 9.3005
R10766 gnd.n4553 gnd.n1939 9.3005
R10767 gnd.n4560 gnd.n4554 9.3005
R10768 gnd.n4559 gnd.n4555 9.3005
R10769 gnd.n4558 gnd.n4557 9.3005
R10770 gnd.n4556 gnd.n1918 9.3005
R10771 gnd.n1916 gnd.n1915 9.3005
R10772 gnd.n4612 gnd.n4611 9.3005
R10773 gnd.n4613 gnd.n1914 9.3005
R10774 gnd.n4615 gnd.n4614 9.3005
R10775 gnd.n1912 gnd.n1911 9.3005
R10776 gnd.n4620 gnd.n4619 9.3005
R10777 gnd.n4621 gnd.n1910 9.3005
R10778 gnd.n4623 gnd.n4622 9.3005
R10779 gnd.n1908 gnd.n1907 9.3005
R10780 gnd.n4628 gnd.n4627 9.3005
R10781 gnd.n4629 gnd.n1906 9.3005
R10782 gnd.n4631 gnd.n4630 9.3005
R10783 gnd.n1902 gnd.n1901 9.3005
R10784 gnd.n4776 gnd.n4775 9.3005
R10785 gnd.n4777 gnd.n1900 9.3005
R10786 gnd.n4779 gnd.n4778 9.3005
R10787 gnd.n1888 gnd.n1887 9.3005
R10788 gnd.n4795 gnd.n4794 9.3005
R10789 gnd.n4796 gnd.n1886 9.3005
R10790 gnd.n4798 gnd.n4797 9.3005
R10791 gnd.n1874 gnd.n1873 9.3005
R10792 gnd.n4814 gnd.n4813 9.3005
R10793 gnd.n4815 gnd.n1872 9.3005
R10794 gnd.n4817 gnd.n4816 9.3005
R10795 gnd.n1860 gnd.n1859 9.3005
R10796 gnd.n4833 gnd.n4832 9.3005
R10797 gnd.n4834 gnd.n1858 9.3005
R10798 gnd.n4836 gnd.n4835 9.3005
R10799 gnd.n1846 gnd.n1845 9.3005
R10800 gnd.n4852 gnd.n4851 9.3005
R10801 gnd.n4853 gnd.n1844 9.3005
R10802 gnd.n4855 gnd.n4854 9.3005
R10803 gnd.n1831 gnd.n1830 9.3005
R10804 gnd.n4871 gnd.n4870 9.3005
R10805 gnd.n4872 gnd.n1829 9.3005
R10806 gnd.n4876 gnd.n4873 9.3005
R10807 gnd.n4875 gnd.n4874 9.3005
R10808 gnd.n1818 gnd.n1817 9.3005
R10809 gnd.n5092 gnd.n5091 9.3005
R10810 gnd.n5093 gnd.n1816 9.3005
R10811 gnd.n5095 gnd.n5094 9.3005
R10812 gnd.n1744 gnd.n1743 9.3005
R10813 gnd.n5133 gnd.n5132 9.3005
R10814 gnd.n5134 gnd.n1742 9.3005
R10815 gnd.n5138 gnd.n5135 9.3005
R10816 gnd.n5137 gnd.n5136 9.3005
R10817 gnd.n1717 gnd.n1716 9.3005
R10818 gnd.n5169 gnd.n5168 9.3005
R10819 gnd.n5170 gnd.n1715 9.3005
R10820 gnd.n5172 gnd.n5171 9.3005
R10821 gnd.n1695 gnd.n1694 9.3005
R10822 gnd.n5197 gnd.n5196 9.3005
R10823 gnd.n5198 gnd.n1693 9.3005
R10824 gnd.n5202 gnd.n5199 9.3005
R10825 gnd.n5201 gnd.n5200 9.3005
R10826 gnd.n1663 gnd.n1662 9.3005
R10827 gnd.n5234 gnd.n5233 9.3005
R10828 gnd.n5235 gnd.n1661 9.3005
R10829 gnd.n5248 gnd.n5236 9.3005
R10830 gnd.n5247 gnd.n5237 9.3005
R10831 gnd.n5246 gnd.n5238 9.3005
R10832 gnd.n5240 gnd.n5239 9.3005
R10833 gnd.n5242 gnd.n5241 9.3005
R10834 gnd.n1622 gnd.n1621 9.3005
R10835 gnd.n5328 gnd.n5327 9.3005
R10836 gnd.n5329 gnd.n1620 9.3005
R10837 gnd.n5331 gnd.n5330 9.3005
R10838 gnd.n1604 gnd.n1603 9.3005
R10839 gnd.n5371 gnd.n5370 9.3005
R10840 gnd.n5372 gnd.n1602 9.3005
R10841 gnd.n5374 gnd.n5373 9.3005
R10842 gnd.n1580 gnd.n1579 9.3005
R10843 gnd.n5405 gnd.n5404 9.3005
R10844 gnd.n5406 gnd.n1578 9.3005
R10845 gnd.n5408 gnd.n5407 9.3005
R10846 gnd.n1557 gnd.n1556 9.3005
R10847 gnd.n5446 gnd.n5445 9.3005
R10848 gnd.n5447 gnd.n1555 9.3005
R10849 gnd.n5449 gnd.n5448 9.3005
R10850 gnd.n1536 gnd.n1535 9.3005
R10851 gnd.n5493 gnd.n5492 9.3005
R10852 gnd.n5494 gnd.n1534 9.3005
R10853 gnd.n5496 gnd.n5495 9.3005
R10854 gnd.n1509 gnd.n1508 9.3005
R10855 gnd.n5525 gnd.n5524 9.3005
R10856 gnd.n5526 gnd.n1507 9.3005
R10857 gnd.n5528 gnd.n5527 9.3005
R10858 gnd.n1487 gnd.n1486 9.3005
R10859 gnd.n5571 gnd.n5570 9.3005
R10860 gnd.n5572 gnd.n1485 9.3005
R10861 gnd.n5574 gnd.n5573 9.3005
R10862 gnd.n1400 gnd.n1399 9.3005
R10863 gnd.n5719 gnd.n5718 9.3005
R10864 gnd.n5720 gnd.n1398 9.3005
R10865 gnd.n5722 gnd.n5721 9.3005
R10866 gnd.n1385 gnd.n1384 9.3005
R10867 gnd.n5738 gnd.n5737 9.3005
R10868 gnd.n5739 gnd.n1383 9.3005
R10869 gnd.n5741 gnd.n5740 9.3005
R10870 gnd.n1371 gnd.n1370 9.3005
R10871 gnd.n5757 gnd.n5756 9.3005
R10872 gnd.n5758 gnd.n1369 9.3005
R10873 gnd.n5760 gnd.n5759 9.3005
R10874 gnd.n1357 gnd.n1356 9.3005
R10875 gnd.n5776 gnd.n5775 9.3005
R10876 gnd.n5777 gnd.n1355 9.3005
R10877 gnd.n5779 gnd.n5778 9.3005
R10878 gnd.n1343 gnd.n1342 9.3005
R10879 gnd.n5795 gnd.n5794 9.3005
R10880 gnd.n5796 gnd.n1341 9.3005
R10881 gnd.n5798 gnd.n5797 9.3005
R10882 gnd.n1329 gnd.n1328 9.3005
R10883 gnd.n5814 gnd.n5813 9.3005
R10884 gnd.n5815 gnd.n1327 9.3005
R10885 gnd.n5990 gnd.n5816 9.3005
R10886 gnd.n5989 gnd.n5817 9.3005
R10887 gnd.n5988 gnd.n5818 9.3005
R10888 gnd.n5842 gnd.n5819 9.3005
R10889 gnd.n5843 gnd.n5841 9.3005
R10890 gnd.n5980 gnd.n5844 9.3005
R10891 gnd.n5979 gnd.n5845 9.3005
R10892 gnd.n5978 gnd.n5846 9.3005
R10893 gnd.n5849 gnd.n5847 9.3005
R10894 gnd.n5930 gnd.n5850 9.3005
R10895 gnd.n5929 gnd.n5851 9.3005
R10896 gnd.n5928 gnd.n5852 9.3005
R10897 gnd.n5855 gnd.n5853 9.3005
R10898 gnd.n5924 gnd.n5856 9.3005
R10899 gnd.n5923 gnd.n5857 9.3005
R10900 gnd.n5922 gnd.n5858 9.3005
R10901 gnd.n5889 gnd.n5859 9.3005
R10902 gnd.n5890 gnd.n5861 9.3005
R10903 gnd.n5892 gnd.n5891 9.3005
R10904 gnd.n5893 gnd.n5888 9.3005
R10905 gnd.n5904 gnd.n5894 9.3005
R10906 gnd.n5903 gnd.n5895 9.3005
R10907 gnd.n5902 gnd.n5896 9.3005
R10908 gnd.n5899 gnd.n5898 9.3005
R10909 gnd.n5897 gnd.n616 9.3005
R10910 gnd.n6925 gnd.n617 9.3005
R10911 gnd.n6924 gnd.n618 9.3005
R10912 gnd.n6923 gnd.n619 9.3005
R10913 gnd.n6916 gnd.n620 9.3005
R10914 gnd.n4539 gnd.n4538 9.3005
R10915 gnd.n1946 gnd.n1945 9.3005
R10916 gnd.n4369 gnd.n4367 9.3005
R10917 gnd.n4370 gnd.n4366 9.3005
R10918 gnd.n4373 gnd.n4365 9.3005
R10919 gnd.n4374 gnd.n4364 9.3005
R10920 gnd.n4377 gnd.n4363 9.3005
R10921 gnd.n4378 gnd.n4362 9.3005
R10922 gnd.n4381 gnd.n4361 9.3005
R10923 gnd.n4382 gnd.n4360 9.3005
R10924 gnd.n4385 gnd.n4359 9.3005
R10925 gnd.n4386 gnd.n4358 9.3005
R10926 gnd.n4389 gnd.n4357 9.3005
R10927 gnd.n4390 gnd.n4356 9.3005
R10928 gnd.n4393 gnd.n4355 9.3005
R10929 gnd.n4394 gnd.n4354 9.3005
R10930 gnd.n4397 gnd.n4353 9.3005
R10931 gnd.n4398 gnd.n4352 9.3005
R10932 gnd.n4401 gnd.n4351 9.3005
R10933 gnd.n4402 gnd.n4350 9.3005
R10934 gnd.n4405 gnd.n4349 9.3005
R10935 gnd.n4406 gnd.n4348 9.3005
R10936 gnd.n4409 gnd.n4347 9.3005
R10937 gnd.n4410 gnd.n4346 9.3005
R10938 gnd.n4413 gnd.n4345 9.3005
R10939 gnd.n4414 gnd.n4344 9.3005
R10940 gnd.n4417 gnd.n4343 9.3005
R10941 gnd.n4418 gnd.n4342 9.3005
R10942 gnd.n4421 gnd.n4341 9.3005
R10943 gnd.n4422 gnd.n4340 9.3005
R10944 gnd.n4425 gnd.n4339 9.3005
R10945 gnd.n4426 gnd.n4338 9.3005
R10946 gnd.n4429 gnd.n4337 9.3005
R10947 gnd.n4430 gnd.n4336 9.3005
R10948 gnd.n4433 gnd.n4335 9.3005
R10949 gnd.n4434 gnd.n4334 9.3005
R10950 gnd.n4437 gnd.n4333 9.3005
R10951 gnd.n4438 gnd.n4332 9.3005
R10952 gnd.n4441 gnd.n4331 9.3005
R10953 gnd.n4442 gnd.n4330 9.3005
R10954 gnd.n4445 gnd.n4329 9.3005
R10955 gnd.n4446 gnd.n4328 9.3005
R10956 gnd.n4449 gnd.n4327 9.3005
R10957 gnd.n4450 gnd.n4326 9.3005
R10958 gnd.n4453 gnd.n4325 9.3005
R10959 gnd.n4454 gnd.n4324 9.3005
R10960 gnd.n4457 gnd.n4323 9.3005
R10961 gnd.n4458 gnd.n4322 9.3005
R10962 gnd.n4461 gnd.n4321 9.3005
R10963 gnd.n4462 gnd.n4320 9.3005
R10964 gnd.n4465 gnd.n4319 9.3005
R10965 gnd.n4466 gnd.n4318 9.3005
R10966 gnd.n4469 gnd.n4317 9.3005
R10967 gnd.n4470 gnd.n4316 9.3005
R10968 gnd.n4473 gnd.n4315 9.3005
R10969 gnd.n4474 gnd.n4314 9.3005
R10970 gnd.n4477 gnd.n4313 9.3005
R10971 gnd.n4478 gnd.n4312 9.3005
R10972 gnd.n4481 gnd.n4311 9.3005
R10973 gnd.n4482 gnd.n4310 9.3005
R10974 gnd.n4485 gnd.n4309 9.3005
R10975 gnd.n4486 gnd.n4308 9.3005
R10976 gnd.n4489 gnd.n4307 9.3005
R10977 gnd.n4490 gnd.n4306 9.3005
R10978 gnd.n4493 gnd.n4305 9.3005
R10979 gnd.n4494 gnd.n4304 9.3005
R10980 gnd.n4497 gnd.n4303 9.3005
R10981 gnd.n4498 gnd.n4302 9.3005
R10982 gnd.n4501 gnd.n4301 9.3005
R10983 gnd.n4502 gnd.n4300 9.3005
R10984 gnd.n4505 gnd.n4299 9.3005
R10985 gnd.n4506 gnd.n4298 9.3005
R10986 gnd.n4509 gnd.n4297 9.3005
R10987 gnd.n4510 gnd.n4296 9.3005
R10988 gnd.n4513 gnd.n4295 9.3005
R10989 gnd.n4514 gnd.n4294 9.3005
R10990 gnd.n4517 gnd.n4293 9.3005
R10991 gnd.n4518 gnd.n4292 9.3005
R10992 gnd.n4521 gnd.n4291 9.3005
R10993 gnd.n4522 gnd.n4290 9.3005
R10994 gnd.n4525 gnd.n4289 9.3005
R10995 gnd.n4527 gnd.n4288 9.3005
R10996 gnd.n4528 gnd.n4287 9.3005
R10997 gnd.n4529 gnd.n4286 9.3005
R10998 gnd.n4530 gnd.n4285 9.3005
R10999 gnd.n4537 gnd.n4536 9.3005
R11000 gnd.n3501 gnd.n3500 9.3005
R11001 gnd.n3474 gnd.n3473 9.3005
R11002 gnd.n3495 gnd.n3494 9.3005
R11003 gnd.n3493 gnd.n3492 9.3005
R11004 gnd.n3478 gnd.n3477 9.3005
R11005 gnd.n3487 gnd.n3486 9.3005
R11006 gnd.n3485 gnd.n3484 9.3005
R11007 gnd.n3469 gnd.n3468 9.3005
R11008 gnd.n3442 gnd.n3441 9.3005
R11009 gnd.n3463 gnd.n3462 9.3005
R11010 gnd.n3461 gnd.n3460 9.3005
R11011 gnd.n3446 gnd.n3445 9.3005
R11012 gnd.n3455 gnd.n3454 9.3005
R11013 gnd.n3453 gnd.n3452 9.3005
R11014 gnd.n3437 gnd.n3436 9.3005
R11015 gnd.n3410 gnd.n3409 9.3005
R11016 gnd.n3431 gnd.n3430 9.3005
R11017 gnd.n3429 gnd.n3428 9.3005
R11018 gnd.n3414 gnd.n3413 9.3005
R11019 gnd.n3423 gnd.n3422 9.3005
R11020 gnd.n3421 gnd.n3420 9.3005
R11021 gnd.n3406 gnd.n3405 9.3005
R11022 gnd.n3379 gnd.n3378 9.3005
R11023 gnd.n3400 gnd.n3399 9.3005
R11024 gnd.n3398 gnd.n3397 9.3005
R11025 gnd.n3383 gnd.n3382 9.3005
R11026 gnd.n3392 gnd.n3391 9.3005
R11027 gnd.n3390 gnd.n3389 9.3005
R11028 gnd.n3374 gnd.n3373 9.3005
R11029 gnd.n3347 gnd.n3346 9.3005
R11030 gnd.n3368 gnd.n3367 9.3005
R11031 gnd.n3366 gnd.n3365 9.3005
R11032 gnd.n3351 gnd.n3350 9.3005
R11033 gnd.n3360 gnd.n3359 9.3005
R11034 gnd.n3358 gnd.n3357 9.3005
R11035 gnd.n3342 gnd.n3341 9.3005
R11036 gnd.n3315 gnd.n3314 9.3005
R11037 gnd.n3336 gnd.n3335 9.3005
R11038 gnd.n3334 gnd.n3333 9.3005
R11039 gnd.n3319 gnd.n3318 9.3005
R11040 gnd.n3328 gnd.n3327 9.3005
R11041 gnd.n3326 gnd.n3325 9.3005
R11042 gnd.n3310 gnd.n3309 9.3005
R11043 gnd.n3283 gnd.n3282 9.3005
R11044 gnd.n3304 gnd.n3303 9.3005
R11045 gnd.n3302 gnd.n3301 9.3005
R11046 gnd.n3287 gnd.n3286 9.3005
R11047 gnd.n3296 gnd.n3295 9.3005
R11048 gnd.n3294 gnd.n3293 9.3005
R11049 gnd.n3279 gnd.n3278 9.3005
R11050 gnd.n3252 gnd.n3251 9.3005
R11051 gnd.n3273 gnd.n3272 9.3005
R11052 gnd.n3271 gnd.n3270 9.3005
R11053 gnd.n3256 gnd.n3255 9.3005
R11054 gnd.n3265 gnd.n3264 9.3005
R11055 gnd.n3263 gnd.n3262 9.3005
R11056 gnd.n3627 gnd.n3626 9.3005
R11057 gnd.n3625 gnd.n2183 9.3005
R11058 gnd.n3624 gnd.n3623 9.3005
R11059 gnd.n3620 gnd.n2184 9.3005
R11060 gnd.n3617 gnd.n2185 9.3005
R11061 gnd.n3616 gnd.n2186 9.3005
R11062 gnd.n3613 gnd.n2187 9.3005
R11063 gnd.n3612 gnd.n2188 9.3005
R11064 gnd.n3609 gnd.n2189 9.3005
R11065 gnd.n3608 gnd.n2190 9.3005
R11066 gnd.n3605 gnd.n2191 9.3005
R11067 gnd.n3604 gnd.n2192 9.3005
R11068 gnd.n3601 gnd.n2193 9.3005
R11069 gnd.n3600 gnd.n2194 9.3005
R11070 gnd.n3597 gnd.n3596 9.3005
R11071 gnd.n3595 gnd.n2195 9.3005
R11072 gnd.n3628 gnd.n2182 9.3005
R11073 gnd.n2869 gnd.n2868 9.3005
R11074 gnd.n2573 gnd.n2572 9.3005
R11075 gnd.n2896 gnd.n2895 9.3005
R11076 gnd.n2897 gnd.n2571 9.3005
R11077 gnd.n2901 gnd.n2898 9.3005
R11078 gnd.n2900 gnd.n2899 9.3005
R11079 gnd.n2545 gnd.n2544 9.3005
R11080 gnd.n2926 gnd.n2925 9.3005
R11081 gnd.n2927 gnd.n2543 9.3005
R11082 gnd.n2929 gnd.n2928 9.3005
R11083 gnd.n2523 gnd.n2522 9.3005
R11084 gnd.n2957 gnd.n2956 9.3005
R11085 gnd.n2958 gnd.n2521 9.3005
R11086 gnd.n2966 gnd.n2959 9.3005
R11087 gnd.n2965 gnd.n2960 9.3005
R11088 gnd.n2964 gnd.n2962 9.3005
R11089 gnd.n2961 gnd.n2470 9.3005
R11090 gnd.n3014 gnd.n2471 9.3005
R11091 gnd.n3013 gnd.n2472 9.3005
R11092 gnd.n3012 gnd.n2473 9.3005
R11093 gnd.n2492 gnd.n2474 9.3005
R11094 gnd.n2494 gnd.n2493 9.3005
R11095 gnd.n2380 gnd.n2379 9.3005
R11096 gnd.n3052 gnd.n3051 9.3005
R11097 gnd.n3053 gnd.n2378 9.3005
R11098 gnd.n3057 gnd.n3054 9.3005
R11099 gnd.n3056 gnd.n3055 9.3005
R11100 gnd.n2353 gnd.n2352 9.3005
R11101 gnd.n3092 gnd.n3091 9.3005
R11102 gnd.n3093 gnd.n2351 9.3005
R11103 gnd.n3097 gnd.n3094 9.3005
R11104 gnd.n3096 gnd.n3095 9.3005
R11105 gnd.n2326 gnd.n2325 9.3005
R11106 gnd.n3137 gnd.n3136 9.3005
R11107 gnd.n3138 gnd.n2324 9.3005
R11108 gnd.n3142 gnd.n3139 9.3005
R11109 gnd.n3141 gnd.n3140 9.3005
R11110 gnd.n2298 gnd.n2297 9.3005
R11111 gnd.n3177 gnd.n3176 9.3005
R11112 gnd.n3178 gnd.n2296 9.3005
R11113 gnd.n3182 gnd.n3179 9.3005
R11114 gnd.n3181 gnd.n3180 9.3005
R11115 gnd.n2271 gnd.n2270 9.3005
R11116 gnd.n3226 gnd.n3225 9.3005
R11117 gnd.n3227 gnd.n2269 9.3005
R11118 gnd.n3231 gnd.n3228 9.3005
R11119 gnd.n3230 gnd.n3229 9.3005
R11120 gnd.n2244 gnd.n2243 9.3005
R11121 gnd.n3520 gnd.n3519 9.3005
R11122 gnd.n3521 gnd.n2242 9.3005
R11123 gnd.n3527 gnd.n3522 9.3005
R11124 gnd.n3526 gnd.n3523 9.3005
R11125 gnd.n3525 gnd.n3524 9.3005
R11126 gnd.n2870 gnd.n2867 9.3005
R11127 gnd.n2652 gnd.n2611 9.3005
R11128 gnd.n2647 gnd.n2646 9.3005
R11129 gnd.n2645 gnd.n2612 9.3005
R11130 gnd.n2644 gnd.n2643 9.3005
R11131 gnd.n2640 gnd.n2613 9.3005
R11132 gnd.n2637 gnd.n2636 9.3005
R11133 gnd.n2635 gnd.n2614 9.3005
R11134 gnd.n2634 gnd.n2633 9.3005
R11135 gnd.n2630 gnd.n2615 9.3005
R11136 gnd.n2627 gnd.n2626 9.3005
R11137 gnd.n2625 gnd.n2616 9.3005
R11138 gnd.n2624 gnd.n2623 9.3005
R11139 gnd.n2620 gnd.n2618 9.3005
R11140 gnd.n2617 gnd.n2597 9.3005
R11141 gnd.n2864 gnd.n2596 9.3005
R11142 gnd.n2866 gnd.n2865 9.3005
R11143 gnd.n2654 gnd.n2653 9.3005
R11144 gnd.n2877 gnd.n2583 9.3005
R11145 gnd.n2884 gnd.n2584 9.3005
R11146 gnd.n2886 gnd.n2885 9.3005
R11147 gnd.n2887 gnd.n2564 9.3005
R11148 gnd.n2906 gnd.n2905 9.3005
R11149 gnd.n2908 gnd.n2556 9.3005
R11150 gnd.n2915 gnd.n2558 9.3005
R11151 gnd.n2916 gnd.n2553 9.3005
R11152 gnd.n2918 gnd.n2917 9.3005
R11153 gnd.n2554 gnd.n2539 9.3005
R11154 gnd.n2934 gnd.n2537 9.3005
R11155 gnd.n2938 gnd.n2937 9.3005
R11156 gnd.n2936 gnd.n2513 9.3005
R11157 gnd.n2973 gnd.n2512 9.3005
R11158 gnd.n2976 gnd.n2975 9.3005
R11159 gnd.n2509 gnd.n2508 9.3005
R11160 gnd.n2982 gnd.n2510 9.3005
R11161 gnd.n2984 gnd.n2983 9.3005
R11162 gnd.n2986 gnd.n2507 9.3005
R11163 gnd.n2989 gnd.n2988 9.3005
R11164 gnd.n2992 gnd.n2990 9.3005
R11165 gnd.n2994 gnd.n2993 9.3005
R11166 gnd.n3000 gnd.n2995 9.3005
R11167 gnd.n2999 gnd.n2998 9.3005
R11168 gnd.n2371 gnd.n2370 9.3005
R11169 gnd.n3066 gnd.n3065 9.3005
R11170 gnd.n3067 gnd.n2364 9.3005
R11171 gnd.n3075 gnd.n2363 9.3005
R11172 gnd.n3078 gnd.n3077 9.3005
R11173 gnd.n3080 gnd.n3079 9.3005
R11174 gnd.n3083 gnd.n2346 9.3005
R11175 gnd.n3081 gnd.n2344 9.3005
R11176 gnd.n3103 gnd.n2342 9.3005
R11177 gnd.n3105 gnd.n3104 9.3005
R11178 gnd.n2316 gnd.n2315 9.3005
R11179 gnd.n3151 gnd.n3150 9.3005
R11180 gnd.n3152 gnd.n2309 9.3005
R11181 gnd.n3160 gnd.n2308 9.3005
R11182 gnd.n3163 gnd.n3162 9.3005
R11183 gnd.n3165 gnd.n3164 9.3005
R11184 gnd.n3168 gnd.n2291 9.3005
R11185 gnd.n3166 gnd.n2289 9.3005
R11186 gnd.n3188 gnd.n2287 9.3005
R11187 gnd.n3190 gnd.n3189 9.3005
R11188 gnd.n2262 gnd.n2261 9.3005
R11189 gnd.n3240 gnd.n3239 9.3005
R11190 gnd.n3241 gnd.n2255 9.3005
R11191 gnd.n3249 gnd.n2254 9.3005
R11192 gnd.n3508 gnd.n3507 9.3005
R11193 gnd.n3510 gnd.n3509 9.3005
R11194 gnd.n3511 gnd.n2235 9.3005
R11195 gnd.n3535 gnd.n3534 9.3005
R11196 gnd.n2236 gnd.n2198 9.3005
R11197 gnd.n2875 gnd.n2874 9.3005
R11198 gnd.n3591 gnd.n2199 9.3005
R11199 gnd.n3590 gnd.n2201 9.3005
R11200 gnd.n3587 gnd.n2202 9.3005
R11201 gnd.n3586 gnd.n2203 9.3005
R11202 gnd.n3583 gnd.n2204 9.3005
R11203 gnd.n3582 gnd.n2205 9.3005
R11204 gnd.n3579 gnd.n2206 9.3005
R11205 gnd.n3578 gnd.n2207 9.3005
R11206 gnd.n3575 gnd.n2208 9.3005
R11207 gnd.n3574 gnd.n2209 9.3005
R11208 gnd.n3571 gnd.n2210 9.3005
R11209 gnd.n3570 gnd.n2211 9.3005
R11210 gnd.n3567 gnd.n2212 9.3005
R11211 gnd.n3566 gnd.n2213 9.3005
R11212 gnd.n3563 gnd.n2214 9.3005
R11213 gnd.n3562 gnd.n2215 9.3005
R11214 gnd.n3559 gnd.n2216 9.3005
R11215 gnd.n3558 gnd.n2217 9.3005
R11216 gnd.n3555 gnd.n2218 9.3005
R11217 gnd.n3554 gnd.n2219 9.3005
R11218 gnd.n3551 gnd.n2220 9.3005
R11219 gnd.n3550 gnd.n2221 9.3005
R11220 gnd.n3547 gnd.n2225 9.3005
R11221 gnd.n3546 gnd.n2226 9.3005
R11222 gnd.n3543 gnd.n2227 9.3005
R11223 gnd.n3542 gnd.n2228 9.3005
R11224 gnd.n3593 gnd.n3592 9.3005
R11225 gnd.n3044 gnd.n3028 9.3005
R11226 gnd.n3043 gnd.n3029 9.3005
R11227 gnd.n3042 gnd.n3030 9.3005
R11228 gnd.n3040 gnd.n3031 9.3005
R11229 gnd.n3039 gnd.n3032 9.3005
R11230 gnd.n3037 gnd.n3033 9.3005
R11231 gnd.n3036 gnd.n3034 9.3005
R11232 gnd.n2334 gnd.n2333 9.3005
R11233 gnd.n3113 gnd.n3112 9.3005
R11234 gnd.n3114 gnd.n2332 9.3005
R11235 gnd.n3131 gnd.n3115 9.3005
R11236 gnd.n3130 gnd.n3116 9.3005
R11237 gnd.n3129 gnd.n3117 9.3005
R11238 gnd.n3127 gnd.n3118 9.3005
R11239 gnd.n3126 gnd.n3119 9.3005
R11240 gnd.n3124 gnd.n3120 9.3005
R11241 gnd.n3123 gnd.n3121 9.3005
R11242 gnd.n2278 gnd.n2277 9.3005
R11243 gnd.n3198 gnd.n3197 9.3005
R11244 gnd.n3199 gnd.n2276 9.3005
R11245 gnd.n3220 gnd.n3200 9.3005
R11246 gnd.n3219 gnd.n3201 9.3005
R11247 gnd.n3218 gnd.n3202 9.3005
R11248 gnd.n3215 gnd.n3203 9.3005
R11249 gnd.n3214 gnd.n3204 9.3005
R11250 gnd.n3212 gnd.n3205 9.3005
R11251 gnd.n3211 gnd.n3206 9.3005
R11252 gnd.n3209 gnd.n3208 9.3005
R11253 gnd.n3207 gnd.n2230 9.3005
R11254 gnd.n2785 gnd.n2784 9.3005
R11255 gnd.n2675 gnd.n2674 9.3005
R11256 gnd.n2799 gnd.n2798 9.3005
R11257 gnd.n2800 gnd.n2673 9.3005
R11258 gnd.n2802 gnd.n2801 9.3005
R11259 gnd.n2663 gnd.n2662 9.3005
R11260 gnd.n2815 gnd.n2814 9.3005
R11261 gnd.n2816 gnd.n2661 9.3005
R11262 gnd.n2848 gnd.n2817 9.3005
R11263 gnd.n2847 gnd.n2818 9.3005
R11264 gnd.n2846 gnd.n2819 9.3005
R11265 gnd.n2845 gnd.n2820 9.3005
R11266 gnd.n2842 gnd.n2821 9.3005
R11267 gnd.n2841 gnd.n2822 9.3005
R11268 gnd.n2840 gnd.n2823 9.3005
R11269 gnd.n2838 gnd.n2824 9.3005
R11270 gnd.n2837 gnd.n2825 9.3005
R11271 gnd.n2834 gnd.n2826 9.3005
R11272 gnd.n2833 gnd.n2827 9.3005
R11273 gnd.n2832 gnd.n2828 9.3005
R11274 gnd.n2830 gnd.n2829 9.3005
R11275 gnd.n2529 gnd.n2528 9.3005
R11276 gnd.n2946 gnd.n2945 9.3005
R11277 gnd.n2947 gnd.n2527 9.3005
R11278 gnd.n2951 gnd.n2948 9.3005
R11279 gnd.n2950 gnd.n2949 9.3005
R11280 gnd.n2451 gnd.n2450 9.3005
R11281 gnd.n3026 gnd.n3025 9.3005
R11282 gnd.n2783 gnd.n2684 9.3005
R11283 gnd.n2686 gnd.n2685 9.3005
R11284 gnd.n2730 gnd.n2728 9.3005
R11285 gnd.n2731 gnd.n2727 9.3005
R11286 gnd.n2734 gnd.n2723 9.3005
R11287 gnd.n2735 gnd.n2722 9.3005
R11288 gnd.n2738 gnd.n2721 9.3005
R11289 gnd.n2739 gnd.n2720 9.3005
R11290 gnd.n2742 gnd.n2719 9.3005
R11291 gnd.n2743 gnd.n2718 9.3005
R11292 gnd.n2746 gnd.n2717 9.3005
R11293 gnd.n2747 gnd.n2716 9.3005
R11294 gnd.n2750 gnd.n2715 9.3005
R11295 gnd.n2751 gnd.n2714 9.3005
R11296 gnd.n2754 gnd.n2713 9.3005
R11297 gnd.n2755 gnd.n2712 9.3005
R11298 gnd.n2758 gnd.n2711 9.3005
R11299 gnd.n2759 gnd.n2710 9.3005
R11300 gnd.n2762 gnd.n2709 9.3005
R11301 gnd.n2763 gnd.n2708 9.3005
R11302 gnd.n2766 gnd.n2707 9.3005
R11303 gnd.n2767 gnd.n2706 9.3005
R11304 gnd.n2770 gnd.n2705 9.3005
R11305 gnd.n2772 gnd.n2704 9.3005
R11306 gnd.n2773 gnd.n2703 9.3005
R11307 gnd.n2774 gnd.n2702 9.3005
R11308 gnd.n2775 gnd.n2701 9.3005
R11309 gnd.n2782 gnd.n2781 9.3005
R11310 gnd.n2791 gnd.n2790 9.3005
R11311 gnd.n2792 gnd.n2678 9.3005
R11312 gnd.n2794 gnd.n2793 9.3005
R11313 gnd.n2669 gnd.n2668 9.3005
R11314 gnd.n2807 gnd.n2806 9.3005
R11315 gnd.n2808 gnd.n2667 9.3005
R11316 gnd.n2810 gnd.n2809 9.3005
R11317 gnd.n2656 gnd.n2655 9.3005
R11318 gnd.n2853 gnd.n2852 9.3005
R11319 gnd.n2854 gnd.n2610 9.3005
R11320 gnd.n2858 gnd.n2856 9.3005
R11321 gnd.n2857 gnd.n2589 9.3005
R11322 gnd.n2876 gnd.n2588 9.3005
R11323 gnd.n2879 gnd.n2878 9.3005
R11324 gnd.n2582 gnd.n2581 9.3005
R11325 gnd.n2890 gnd.n2888 9.3005
R11326 gnd.n2889 gnd.n2563 9.3005
R11327 gnd.n2907 gnd.n2562 9.3005
R11328 gnd.n2910 gnd.n2909 9.3005
R11329 gnd.n2557 gnd.n2552 9.3005
R11330 gnd.n2920 gnd.n2919 9.3005
R11331 gnd.n2555 gnd.n2535 9.3005
R11332 gnd.n2941 gnd.n2536 9.3005
R11333 gnd.n2940 gnd.n2939 9.3005
R11334 gnd.n2538 gnd.n2514 9.3005
R11335 gnd.n2972 gnd.n2971 9.3005
R11336 gnd.n2974 gnd.n2459 9.3005
R11337 gnd.n3021 gnd.n2460 9.3005
R11338 gnd.n3020 gnd.n2461 9.3005
R11339 gnd.n3019 gnd.n2462 9.3005
R11340 gnd.n2985 gnd.n2463 9.3005
R11341 gnd.n2987 gnd.n2481 9.3005
R11342 gnd.n3007 gnd.n2482 9.3005
R11343 gnd.n3006 gnd.n2483 9.3005
R11344 gnd.n3005 gnd.n2484 9.3005
R11345 gnd.n2996 gnd.n2485 9.3005
R11346 gnd.n2997 gnd.n2372 9.3005
R11347 gnd.n3063 gnd.n3062 9.3005
R11348 gnd.n3064 gnd.n2365 9.3005
R11349 gnd.n3074 gnd.n3073 9.3005
R11350 gnd.n3076 gnd.n2361 9.3005
R11351 gnd.n3086 gnd.n2362 9.3005
R11352 gnd.n3085 gnd.n3084 9.3005
R11353 gnd.n3082 gnd.n2340 9.3005
R11354 gnd.n3108 gnd.n2341 9.3005
R11355 gnd.n3107 gnd.n3106 9.3005
R11356 gnd.n2343 gnd.n2317 9.3005
R11357 gnd.n3148 gnd.n3147 9.3005
R11358 gnd.n3149 gnd.n2310 9.3005
R11359 gnd.n3159 gnd.n3158 9.3005
R11360 gnd.n3161 gnd.n2306 9.3005
R11361 gnd.n3171 gnd.n2307 9.3005
R11362 gnd.n3170 gnd.n3169 9.3005
R11363 gnd.n3167 gnd.n2285 9.3005
R11364 gnd.n3193 gnd.n2286 9.3005
R11365 gnd.n3192 gnd.n3191 9.3005
R11366 gnd.n2288 gnd.n2263 9.3005
R11367 gnd.n3237 gnd.n3236 9.3005
R11368 gnd.n3238 gnd.n2256 9.3005
R11369 gnd.n3248 gnd.n3247 9.3005
R11370 gnd.n3506 gnd.n2252 9.3005
R11371 gnd.n3514 gnd.n2253 9.3005
R11372 gnd.n3513 gnd.n3512 9.3005
R11373 gnd.n2234 gnd.n2233 9.3005
R11374 gnd.n3537 gnd.n3536 9.3005
R11375 gnd.n2680 gnd.n2679 9.3005
R11376 gnd.n3859 gnd.n3735 9.3005
R11377 gnd.n3861 gnd.n3860 9.3005
R11378 gnd.n3858 gnd.n3737 9.3005
R11379 gnd.n3857 gnd.n3856 9.3005
R11380 gnd.n3739 gnd.n3738 9.3005
R11381 gnd.n3850 gnd.n3849 9.3005
R11382 gnd.n3848 gnd.n3741 9.3005
R11383 gnd.n3847 gnd.n3846 9.3005
R11384 gnd.n3743 gnd.n3742 9.3005
R11385 gnd.n3840 gnd.n3839 9.3005
R11386 gnd.n3838 gnd.n3745 9.3005
R11387 gnd.n3837 gnd.n3836 9.3005
R11388 gnd.n3747 gnd.n3746 9.3005
R11389 gnd.n3830 gnd.n3829 9.3005
R11390 gnd.n3828 gnd.n3749 9.3005
R11391 gnd.n3827 gnd.n3826 9.3005
R11392 gnd.n3751 gnd.n3750 9.3005
R11393 gnd.n3820 gnd.n3819 9.3005
R11394 gnd.n3818 gnd.n3753 9.3005
R11395 gnd.n3817 gnd.n3816 9.3005
R11396 gnd.n3755 gnd.n3754 9.3005
R11397 gnd.n3810 gnd.n3809 9.3005
R11398 gnd.n3808 gnd.n3760 9.3005
R11399 gnd.n3807 gnd.n3806 9.3005
R11400 gnd.n3762 gnd.n3761 9.3005
R11401 gnd.n3800 gnd.n3799 9.3005
R11402 gnd.n3798 gnd.n3764 9.3005
R11403 gnd.n3797 gnd.n3796 9.3005
R11404 gnd.n3766 gnd.n3765 9.3005
R11405 gnd.n3790 gnd.n3789 9.3005
R11406 gnd.n3788 gnd.n3768 9.3005
R11407 gnd.n3787 gnd.n3786 9.3005
R11408 gnd.n3770 gnd.n3769 9.3005
R11409 gnd.n3780 gnd.n3779 9.3005
R11410 gnd.n3778 gnd.n3772 9.3005
R11411 gnd.n3777 gnd.n3776 9.3005
R11412 gnd.n3773 gnd.n2155 9.3005
R11413 gnd.n3734 gnd.n3731 9.3005
R11414 gnd.n3869 gnd.n3868 9.3005
R11415 gnd.n4107 gnd.n2154 9.3005
R11416 gnd.n4109 gnd.n4108 9.3005
R11417 gnd.n2141 gnd.n2140 9.3005
R11418 gnd.n4122 gnd.n4121 9.3005
R11419 gnd.n4123 gnd.n2139 9.3005
R11420 gnd.n4125 gnd.n4124 9.3005
R11421 gnd.n2124 gnd.n2123 9.3005
R11422 gnd.n4138 gnd.n4137 9.3005
R11423 gnd.n4139 gnd.n2122 9.3005
R11424 gnd.n4141 gnd.n4140 9.3005
R11425 gnd.n2109 gnd.n2108 9.3005
R11426 gnd.n4154 gnd.n4153 9.3005
R11427 gnd.n4155 gnd.n2107 9.3005
R11428 gnd.n4157 gnd.n4156 9.3005
R11429 gnd.n2092 gnd.n2091 9.3005
R11430 gnd.n4170 gnd.n4169 9.3005
R11431 gnd.n4171 gnd.n2090 9.3005
R11432 gnd.n4173 gnd.n4172 9.3005
R11433 gnd.n2077 gnd.n2076 9.3005
R11434 gnd.n4186 gnd.n4185 9.3005
R11435 gnd.n4187 gnd.n2075 9.3005
R11436 gnd.n4189 gnd.n4188 9.3005
R11437 gnd.n2060 gnd.n2059 9.3005
R11438 gnd.n4202 gnd.n4201 9.3005
R11439 gnd.n4203 gnd.n2058 9.3005
R11440 gnd.n4205 gnd.n4204 9.3005
R11441 gnd.n2045 gnd.n2044 9.3005
R11442 gnd.n4106 gnd.n4105 9.3005
R11443 gnd.n4218 gnd.n4217 9.3005
R11444 gnd.n4219 gnd.n2043 9.3005
R11445 gnd.n4221 gnd.n4220 9.3005
R11446 gnd.n2027 gnd.n2026 9.3005
R11447 gnd.n4234 gnd.n4233 9.3005
R11448 gnd.n4235 gnd.n2025 9.3005
R11449 gnd.n4237 gnd.n4236 9.3005
R11450 gnd.n2012 gnd.n2011 9.3005
R11451 gnd.n4250 gnd.n4249 9.3005
R11452 gnd.n4251 gnd.n2010 9.3005
R11453 gnd.n4253 gnd.n4252 9.3005
R11454 gnd.n1994 gnd.n1993 9.3005
R11455 gnd.n4276 gnd.n4275 9.3005
R11456 gnd.n4277 gnd.n1992 9.3005
R11457 gnd.n4280 gnd.n4279 9.3005
R11458 gnd.n4278 gnd.n987 9.3005
R11459 gnd.n6313 gnd.n988 9.3005
R11460 gnd.n6312 gnd.n989 9.3005
R11461 gnd.n6311 gnd.n990 9.3005
R11462 gnd.n1009 gnd.n991 9.3005
R11463 gnd.n6301 gnd.n1010 9.3005
R11464 gnd.n6300 gnd.n1011 9.3005
R11465 gnd.n6299 gnd.n1012 9.3005
R11466 gnd.n1030 gnd.n1013 9.3005
R11467 gnd.n6289 gnd.n1031 9.3005
R11468 gnd.n6288 gnd.n1032 9.3005
R11469 gnd.n6287 gnd.n1033 9.3005
R11470 gnd.n1051 gnd.n1034 9.3005
R11471 gnd.n6277 gnd.n1052 9.3005
R11472 gnd.n6276 gnd.n1053 9.3005
R11473 gnd.n6275 gnd.n1054 9.3005
R11474 gnd.n1073 gnd.n1055 9.3005
R11475 gnd.n6265 gnd.n1074 9.3005
R11476 gnd.n6264 gnd.n1075 9.3005
R11477 gnd.n6263 gnd.n1076 9.3005
R11478 gnd.n1093 gnd.n1077 9.3005
R11479 gnd.n6253 gnd.n6252 9.3005
R11480 gnd.n1124 gnd.n1118 9.3005
R11481 gnd.n6226 gnd.n1117 9.3005
R11482 gnd.n6227 gnd.n1116 9.3005
R11483 gnd.n6228 gnd.n1115 9.3005
R11484 gnd.n1114 gnd.n1111 9.3005
R11485 gnd.n6233 gnd.n1110 9.3005
R11486 gnd.n6234 gnd.n1109 9.3005
R11487 gnd.n6235 gnd.n1108 9.3005
R11488 gnd.n1107 gnd.n1104 9.3005
R11489 gnd.n6240 gnd.n1103 9.3005
R11490 gnd.n6241 gnd.n1102 9.3005
R11491 gnd.n6242 gnd.n1101 9.3005
R11492 gnd.n1100 gnd.n1097 9.3005
R11493 gnd.n1099 gnd.n1095 9.3005
R11494 gnd.n6249 gnd.n1094 9.3005
R11495 gnd.n6251 gnd.n6250 9.3005
R11496 gnd.n6218 gnd.n1127 9.3005
R11497 gnd.n6217 gnd.n1128 9.3005
R11498 gnd.n1132 gnd.n1129 9.3005
R11499 gnd.n6212 gnd.n1133 9.3005
R11500 gnd.n6211 gnd.n1134 9.3005
R11501 gnd.n6210 gnd.n1135 9.3005
R11502 gnd.n1139 gnd.n1136 9.3005
R11503 gnd.n6205 gnd.n1140 9.3005
R11504 gnd.n6204 gnd.n1141 9.3005
R11505 gnd.n6203 gnd.n1142 9.3005
R11506 gnd.n1146 gnd.n1143 9.3005
R11507 gnd.n6198 gnd.n1147 9.3005
R11508 gnd.n6197 gnd.n1148 9.3005
R11509 gnd.n6196 gnd.n1149 9.3005
R11510 gnd.n1153 gnd.n1150 9.3005
R11511 gnd.n6191 gnd.n1154 9.3005
R11512 gnd.n6190 gnd.n1155 9.3005
R11513 gnd.n6189 gnd.n1156 9.3005
R11514 gnd.n1161 gnd.n1159 9.3005
R11515 gnd.n6184 gnd.n6183 9.3005
R11516 gnd.n6219 gnd.n1126 9.3005
R11517 gnd.n3874 gnd.n3873 9.3005
R11518 gnd.n3875 gnd.n3730 9.3005
R11519 gnd.n3878 gnd.n3876 9.3005
R11520 gnd.n3879 gnd.n3729 9.3005
R11521 gnd.n3882 gnd.n3881 9.3005
R11522 gnd.n3883 gnd.n3728 9.3005
R11523 gnd.n3886 gnd.n3884 9.3005
R11524 gnd.n3887 gnd.n3727 9.3005
R11525 gnd.n3890 gnd.n3889 9.3005
R11526 gnd.n3891 gnd.n3726 9.3005
R11527 gnd.n3894 gnd.n3892 9.3005
R11528 gnd.n3895 gnd.n3725 9.3005
R11529 gnd.n3898 gnd.n3897 9.3005
R11530 gnd.n3899 gnd.n3724 9.3005
R11531 gnd.n3902 gnd.n3900 9.3005
R11532 gnd.n3903 gnd.n3723 9.3005
R11533 gnd.n3906 gnd.n3905 9.3005
R11534 gnd.n3907 gnd.n3722 9.3005
R11535 gnd.n3910 gnd.n3908 9.3005
R11536 gnd.n3911 gnd.n3721 9.3005
R11537 gnd.n3914 gnd.n3913 9.3005
R11538 gnd.n3915 gnd.n3720 9.3005
R11539 gnd.n3918 gnd.n3916 9.3005
R11540 gnd.n3919 gnd.n3719 9.3005
R11541 gnd.n3922 gnd.n3921 9.3005
R11542 gnd.n3923 gnd.n3718 9.3005
R11543 gnd.n3926 gnd.n3924 9.3005
R11544 gnd.n3927 gnd.n3717 9.3005
R11545 gnd.n3930 gnd.n3929 9.3005
R11546 gnd.n3931 gnd.n3716 9.3005
R11547 gnd.n3934 gnd.n3932 9.3005
R11548 gnd.n3935 gnd.n2035 9.3005
R11549 gnd.n3938 gnd.n3936 9.3005
R11550 gnd.n3939 gnd.n3715 9.3005
R11551 gnd.n3942 gnd.n3941 9.3005
R11552 gnd.n3943 gnd.n3714 9.3005
R11553 gnd.n3946 gnd.n3944 9.3005
R11554 gnd.n3947 gnd.n3713 9.3005
R11555 gnd.n3950 gnd.n3949 9.3005
R11556 gnd.n3951 gnd.n3712 9.3005
R11557 gnd.n3954 gnd.n3952 9.3005
R11558 gnd.n3955 gnd.n3711 9.3005
R11559 gnd.n3958 gnd.n3957 9.3005
R11560 gnd.n3959 gnd.n3710 9.3005
R11561 gnd.n3964 gnd.n3960 9.3005
R11562 gnd.n3965 gnd.n3709 9.3005
R11563 gnd.n3970 gnd.n3969 9.3005
R11564 gnd.n3971 gnd.n3708 9.3005
R11565 gnd.n3978 gnd.n3972 9.3005
R11566 gnd.n3977 gnd.n3973 9.3005
R11567 gnd.n3976 gnd.n3975 9.3005
R11568 gnd.n3974 gnd.n1931 9.3005
R11569 gnd.n4573 gnd.n1932 9.3005
R11570 gnd.n4574 gnd.n1930 9.3005
R11571 gnd.n4576 gnd.n4575 9.3005
R11572 gnd.n4577 gnd.n1929 9.3005
R11573 gnd.n4581 gnd.n4578 9.3005
R11574 gnd.n4582 gnd.n1928 9.3005
R11575 gnd.n4586 gnd.n4585 9.3005
R11576 gnd.n4587 gnd.n1927 9.3005
R11577 gnd.n4590 gnd.n4589 9.3005
R11578 gnd.n4588 gnd.n1163 9.3005
R11579 gnd.n6180 gnd.n1162 9.3005
R11580 gnd.n6182 gnd.n6181 9.3005
R11581 gnd.n3871 gnd.n3870 9.3005
R11582 gnd.n4009 gnd.n4008 9.3005
R11583 gnd.n4056 gnd.n3662 9.3005
R11584 gnd.n4054 gnd.n3663 9.3005
R11585 gnd.n4053 gnd.n3664 9.3005
R11586 gnd.n4051 gnd.n3665 9.3005
R11587 gnd.n4050 gnd.n3666 9.3005
R11588 gnd.n4048 gnd.n3667 9.3005
R11589 gnd.n4047 gnd.n3668 9.3005
R11590 gnd.n4045 gnd.n3669 9.3005
R11591 gnd.n4044 gnd.n3670 9.3005
R11592 gnd.n4042 gnd.n3671 9.3005
R11593 gnd.n4041 gnd.n3672 9.3005
R11594 gnd.n4039 gnd.n3673 9.3005
R11595 gnd.n4038 gnd.n3674 9.3005
R11596 gnd.n4036 gnd.n3675 9.3005
R11597 gnd.n4035 gnd.n3676 9.3005
R11598 gnd.n4033 gnd.n3677 9.3005
R11599 gnd.n4032 gnd.n3678 9.3005
R11600 gnd.n4030 gnd.n3679 9.3005
R11601 gnd.n4029 gnd.n3680 9.3005
R11602 gnd.n4027 gnd.n3681 9.3005
R11603 gnd.n4026 gnd.n3682 9.3005
R11604 gnd.n4024 gnd.n3683 9.3005
R11605 gnd.n4023 gnd.n3684 9.3005
R11606 gnd.n4021 gnd.n3685 9.3005
R11607 gnd.n4020 gnd.n3686 9.3005
R11608 gnd.n4018 gnd.n3687 9.3005
R11609 gnd.n4017 gnd.n3688 9.3005
R11610 gnd.n4015 gnd.n3689 9.3005
R11611 gnd.n4014 gnd.n3690 9.3005
R11612 gnd.n4012 gnd.n3691 9.3005
R11613 gnd.n4011 gnd.n3692 9.3005
R11614 gnd.n4058 gnd.n4057 9.3005
R11615 gnd.n4066 gnd.n4065 9.3005
R11616 gnd.n4067 gnd.n3658 9.3005
R11617 gnd.n3657 gnd.n3655 9.3005
R11618 gnd.n4073 gnd.n3654 9.3005
R11619 gnd.n4074 gnd.n3653 9.3005
R11620 gnd.n4075 gnd.n3652 9.3005
R11621 gnd.n3651 gnd.n3649 9.3005
R11622 gnd.n4081 gnd.n3648 9.3005
R11623 gnd.n4082 gnd.n3647 9.3005
R11624 gnd.n4083 gnd.n3646 9.3005
R11625 gnd.n3645 gnd.n3643 9.3005
R11626 gnd.n4089 gnd.n3642 9.3005
R11627 gnd.n4090 gnd.n3641 9.3005
R11628 gnd.n4091 gnd.n3640 9.3005
R11629 gnd.n3639 gnd.n3637 9.3005
R11630 gnd.n4097 gnd.n3636 9.3005
R11631 gnd.n4099 gnd.n4098 9.3005
R11632 gnd.n4064 gnd.n3661 9.3005
R11633 gnd.n4063 gnd.n4062 9.3005
R11634 gnd.n2149 gnd.n2148 9.3005
R11635 gnd.n4114 gnd.n4113 9.3005
R11636 gnd.n4115 gnd.n2147 9.3005
R11637 gnd.n4117 gnd.n4116 9.3005
R11638 gnd.n2133 gnd.n2132 9.3005
R11639 gnd.n4130 gnd.n4129 9.3005
R11640 gnd.n4131 gnd.n2131 9.3005
R11641 gnd.n4133 gnd.n4132 9.3005
R11642 gnd.n2117 gnd.n2116 9.3005
R11643 gnd.n4146 gnd.n4145 9.3005
R11644 gnd.n4147 gnd.n2115 9.3005
R11645 gnd.n4149 gnd.n4148 9.3005
R11646 gnd.n2101 gnd.n2100 9.3005
R11647 gnd.n4162 gnd.n4161 9.3005
R11648 gnd.n4163 gnd.n2099 9.3005
R11649 gnd.n4165 gnd.n4164 9.3005
R11650 gnd.n2085 gnd.n2084 9.3005
R11651 gnd.n4178 gnd.n4177 9.3005
R11652 gnd.n4179 gnd.n2083 9.3005
R11653 gnd.n4181 gnd.n4180 9.3005
R11654 gnd.n2069 gnd.n2068 9.3005
R11655 gnd.n4194 gnd.n4193 9.3005
R11656 gnd.n4195 gnd.n2067 9.3005
R11657 gnd.n4197 gnd.n4196 9.3005
R11658 gnd.n2053 gnd.n2052 9.3005
R11659 gnd.n4210 gnd.n4209 9.3005
R11660 gnd.n4211 gnd.n2051 9.3005
R11661 gnd.n4213 gnd.n4212 9.3005
R11662 gnd.n2037 gnd.n2036 9.3005
R11663 gnd.n4226 gnd.n4225 9.3005
R11664 gnd.n4227 gnd.n2034 9.3005
R11665 gnd.n4229 gnd.n4228 9.3005
R11666 gnd.n2019 gnd.n2018 9.3005
R11667 gnd.n4242 gnd.n4241 9.3005
R11668 gnd.n4243 gnd.n2017 9.3005
R11669 gnd.n4245 gnd.n4244 9.3005
R11670 gnd.n2004 gnd.n2003 9.3005
R11671 gnd.n4258 gnd.n4257 9.3005
R11672 gnd.n4259 gnd.n2002 9.3005
R11673 gnd.n4271 gnd.n4260 9.3005
R11674 gnd.n4270 gnd.n4261 9.3005
R11675 gnd.n4269 gnd.n4262 9.3005
R11676 gnd.n4268 gnd.n4263 9.3005
R11677 gnd.n4266 gnd.n4265 9.3005
R11678 gnd.n4264 gnd.n998 9.3005
R11679 gnd.n6307 gnd.n999 9.3005
R11680 gnd.n6306 gnd.n1000 9.3005
R11681 gnd.n6305 gnd.n1001 9.3005
R11682 gnd.n1020 gnd.n1002 9.3005
R11683 gnd.n6295 gnd.n1021 9.3005
R11684 gnd.n6294 gnd.n1022 9.3005
R11685 gnd.n6293 gnd.n1023 9.3005
R11686 gnd.n1040 gnd.n1024 9.3005
R11687 gnd.n6283 gnd.n1041 9.3005
R11688 gnd.n6282 gnd.n1042 9.3005
R11689 gnd.n6281 gnd.n1043 9.3005
R11690 gnd.n1062 gnd.n1044 9.3005
R11691 gnd.n6271 gnd.n1063 9.3005
R11692 gnd.n6270 gnd.n1064 9.3005
R11693 gnd.n6269 gnd.n1065 9.3005
R11694 gnd.n1083 gnd.n1066 9.3005
R11695 gnd.n6259 gnd.n1084 9.3005
R11696 gnd.n6258 gnd.n1085 9.3005
R11697 gnd.n6257 gnd.n1086 9.3005
R11698 gnd.n4101 gnd.n4100 9.3005
R11699 gnd.n7223 gnd.n7222 9.3005
R11700 gnd.n467 gnd.n466 9.3005
R11701 gnd.n7217 gnd.n7216 9.3005
R11702 gnd.n7215 gnd.n7214 9.3005
R11703 gnd.n475 gnd.n474 9.3005
R11704 gnd.n7209 gnd.n7208 9.3005
R11705 gnd.n7207 gnd.n7206 9.3005
R11706 gnd.n483 gnd.n482 9.3005
R11707 gnd.n7201 gnd.n7200 9.3005
R11708 gnd.n7199 gnd.n7198 9.3005
R11709 gnd.n491 gnd.n490 9.3005
R11710 gnd.n7193 gnd.n7192 9.3005
R11711 gnd.n7191 gnd.n7190 9.3005
R11712 gnd.n499 gnd.n498 9.3005
R11713 gnd.n7185 gnd.n7184 9.3005
R11714 gnd.n7183 gnd.n7182 9.3005
R11715 gnd.n509 gnd.n508 9.3005
R11716 gnd.n5936 gnd.n5932 9.3005
R11717 gnd.n7225 gnd.n7224 9.3005
R11718 gnd.n7187 gnd.n7186 9.3005
R11719 gnd.n7189 gnd.n7188 9.3005
R11720 gnd.n495 gnd.n494 9.3005
R11721 gnd.n7195 gnd.n7194 9.3005
R11722 gnd.n7197 gnd.n7196 9.3005
R11723 gnd.n487 gnd.n486 9.3005
R11724 gnd.n7203 gnd.n7202 9.3005
R11725 gnd.n7205 gnd.n7204 9.3005
R11726 gnd.n479 gnd.n478 9.3005
R11727 gnd.n7211 gnd.n7210 9.3005
R11728 gnd.n7213 gnd.n7212 9.3005
R11729 gnd.n471 gnd.n470 9.3005
R11730 gnd.n7219 gnd.n7218 9.3005
R11731 gnd.n7221 gnd.n7220 9.3005
R11732 gnd.n463 gnd.n462 9.3005
R11733 gnd.n7227 gnd.n7226 9.3005
R11734 gnd.n505 gnd.n504 9.3005
R11735 gnd.n7181 gnd.n7180 9.3005
R11736 gnd.n5967 gnd.n5966 9.3005
R11737 gnd.n5965 gnd.n5933 9.3005
R11738 gnd.n5964 gnd.n5963 9.3005
R11739 gnd.n5962 gnd.n5941 9.3005
R11740 gnd.n5961 gnd.n5960 9.3005
R11741 gnd.n5959 gnd.n5942 9.3005
R11742 gnd.n5955 gnd.n5954 9.3005
R11743 gnd.n5953 gnd.n5947 9.3005
R11744 gnd.n5952 gnd.n5951 9.3005
R11745 gnd.n5950 gnd.n5948 9.3005
R11746 gnd.n6153 gnd.n1187 9.3005
R11747 gnd.n6152 gnd.n6151 9.3005
R11748 gnd.n6150 gnd.n1191 9.3005
R11749 gnd.n6149 gnd.n6148 9.3005
R11750 gnd.n6147 gnd.n1192 9.3005
R11751 gnd.n6146 gnd.n6145 9.3005
R11752 gnd.n6144 gnd.n1196 9.3005
R11753 gnd.n6143 gnd.n6142 9.3005
R11754 gnd.n6141 gnd.n1197 9.3005
R11755 gnd.n6140 gnd.n6139 9.3005
R11756 gnd.n6138 gnd.n1201 9.3005
R11757 gnd.n6137 gnd.n6136 9.3005
R11758 gnd.n6135 gnd.n1202 9.3005
R11759 gnd.n6134 gnd.n6133 9.3005
R11760 gnd.n6132 gnd.n1206 9.3005
R11761 gnd.n6131 gnd.n6130 9.3005
R11762 gnd.n6129 gnd.n1207 9.3005
R11763 gnd.n6128 gnd.n6127 9.3005
R11764 gnd.n6126 gnd.n1211 9.3005
R11765 gnd.n6125 gnd.n6124 9.3005
R11766 gnd.n6123 gnd.n1212 9.3005
R11767 gnd.n6122 gnd.n6121 9.3005
R11768 gnd.n6120 gnd.n1216 9.3005
R11769 gnd.n6119 gnd.n6118 9.3005
R11770 gnd.n6117 gnd.n1217 9.3005
R11771 gnd.n6116 gnd.n6115 9.3005
R11772 gnd.n6114 gnd.n1221 9.3005
R11773 gnd.n6113 gnd.n6112 9.3005
R11774 gnd.n6111 gnd.n1222 9.3005
R11775 gnd.n6110 gnd.n6109 9.3005
R11776 gnd.n6108 gnd.n1226 9.3005
R11777 gnd.n6107 gnd.n6106 9.3005
R11778 gnd.n6105 gnd.n1227 9.3005
R11779 gnd.n6104 gnd.n6103 9.3005
R11780 gnd.n6102 gnd.n1231 9.3005
R11781 gnd.n6101 gnd.n6100 9.3005
R11782 gnd.n6099 gnd.n1232 9.3005
R11783 gnd.n6098 gnd.n6097 9.3005
R11784 gnd.n6096 gnd.n1236 9.3005
R11785 gnd.n6095 gnd.n6094 9.3005
R11786 gnd.n6093 gnd.n1237 9.3005
R11787 gnd.n6092 gnd.n6091 9.3005
R11788 gnd.n6090 gnd.n1241 9.3005
R11789 gnd.n6089 gnd.n6088 9.3005
R11790 gnd.n6087 gnd.n1242 9.3005
R11791 gnd.n6086 gnd.n6085 9.3005
R11792 gnd.n6084 gnd.n1246 9.3005
R11793 gnd.n6083 gnd.n6082 9.3005
R11794 gnd.n6081 gnd.n1247 9.3005
R11795 gnd.n6080 gnd.n6079 9.3005
R11796 gnd.n6078 gnd.n1251 9.3005
R11797 gnd.n6077 gnd.n6076 9.3005
R11798 gnd.n6075 gnd.n1252 9.3005
R11799 gnd.n6074 gnd.n6073 9.3005
R11800 gnd.n6072 gnd.n1256 9.3005
R11801 gnd.n6071 gnd.n6070 9.3005
R11802 gnd.n6069 gnd.n1257 9.3005
R11803 gnd.n6068 gnd.n6067 9.3005
R11804 gnd.n6066 gnd.n1261 9.3005
R11805 gnd.n6065 gnd.n6064 9.3005
R11806 gnd.n6063 gnd.n1262 9.3005
R11807 gnd.n6062 gnd.n6061 9.3005
R11808 gnd.n6060 gnd.n1266 9.3005
R11809 gnd.n6059 gnd.n6058 9.3005
R11810 gnd.n6057 gnd.n1267 9.3005
R11811 gnd.n6056 gnd.n6055 9.3005
R11812 gnd.n6054 gnd.n1271 9.3005
R11813 gnd.n6053 gnd.n6052 9.3005
R11814 gnd.n6051 gnd.n1272 9.3005
R11815 gnd.n6050 gnd.n6049 9.3005
R11816 gnd.n6048 gnd.n1276 9.3005
R11817 gnd.n6047 gnd.n6046 9.3005
R11818 gnd.n6045 gnd.n1277 9.3005
R11819 gnd.n6044 gnd.n6043 9.3005
R11820 gnd.n6042 gnd.n1281 9.3005
R11821 gnd.n6041 gnd.n6040 9.3005
R11822 gnd.n6039 gnd.n1282 9.3005
R11823 gnd.n6038 gnd.n6037 9.3005
R11824 gnd.n6036 gnd.n1286 9.3005
R11825 gnd.n6035 gnd.n6034 9.3005
R11826 gnd.n6033 gnd.n1287 9.3005
R11827 gnd.n6032 gnd.n6031 9.3005
R11828 gnd.n6030 gnd.n1291 9.3005
R11829 gnd.n6029 gnd.n6028 9.3005
R11830 gnd.n6027 gnd.n1292 9.3005
R11831 gnd.n6026 gnd.n6025 9.3005
R11832 gnd.n6024 gnd.n1296 9.3005
R11833 gnd.n6023 gnd.n6022 9.3005
R11834 gnd.n6021 gnd.n1297 9.3005
R11835 gnd.n6020 gnd.n6019 9.3005
R11836 gnd.n6018 gnd.n1301 9.3005
R11837 gnd.n6017 gnd.n6016 9.3005
R11838 gnd.n6015 gnd.n1302 9.3005
R11839 gnd.n6014 gnd.n6013 9.3005
R11840 gnd.n6012 gnd.n1306 9.3005
R11841 gnd.n6011 gnd.n6010 9.3005
R11842 gnd.n6009 gnd.n1307 9.3005
R11843 gnd.n6008 gnd.n6007 9.3005
R11844 gnd.n6006 gnd.n1311 9.3005
R11845 gnd.n6005 gnd.n6004 9.3005
R11846 gnd.n6003 gnd.n1312 9.3005
R11847 gnd.n6155 gnd.n6154 9.3005
R11848 gnd.n6158 gnd.n6157 9.3005
R11849 gnd.n6159 gnd.n1182 9.3005
R11850 gnd.n6161 gnd.n6160 9.3005
R11851 gnd.n6163 gnd.n6162 9.3005
R11852 gnd.n6164 gnd.n1175 9.3005
R11853 gnd.n6166 gnd.n6165 9.3005
R11854 gnd.n6167 gnd.n1174 9.3005
R11855 gnd.n6169 gnd.n6168 9.3005
R11856 gnd.n6170 gnd.n1168 9.3005
R11857 gnd.n6156 gnd.n1186 9.3005
R11858 gnd.n4007 gnd.n3694 9.3005
R11859 gnd.n4006 gnd.n4005 9.3005
R11860 gnd.n4004 gnd.n3695 9.3005
R11861 gnd.n4003 gnd.n4002 9.3005
R11862 gnd.n4001 gnd.n3698 9.3005
R11863 gnd.n4000 gnd.n3999 9.3005
R11864 gnd.n3998 gnd.n3699 9.3005
R11865 gnd.n3997 gnd.n3996 9.3005
R11866 gnd.n3995 gnd.n3702 9.3005
R11867 gnd.n3994 gnd.n3993 9.3005
R11868 gnd.n3992 gnd.n3703 9.3005
R11869 gnd.n3991 gnd.n3990 9.3005
R11870 gnd.n3989 gnd.n3705 9.3005
R11871 gnd.n3988 gnd.n3987 9.3005
R11872 gnd.n3986 gnd.n3706 9.3005
R11873 gnd.n3985 gnd.n3984 9.3005
R11874 gnd.n3983 gnd.n3982 9.3005
R11875 gnd.n1935 gnd.n1934 9.3005
R11876 gnd.n4566 gnd.n4565 9.3005
R11877 gnd.n4567 gnd.n1933 9.3005
R11878 gnd.n4569 gnd.n4568 9.3005
R11879 gnd.n1922 gnd.n1920 9.3005
R11880 gnd.n4604 gnd.n4603 9.3005
R11881 gnd.n4602 gnd.n1921 9.3005
R11882 gnd.n4601 gnd.n4600 9.3005
R11883 gnd.n4599 gnd.n1923 9.3005
R11884 gnd.n4598 gnd.n4597 9.3005
R11885 gnd.n4596 gnd.n1926 9.3005
R11886 gnd.n4595 gnd.n4594 9.3005
R11887 gnd.n1167 gnd.n1165 9.3005
R11888 gnd.n6176 gnd.n6175 9.3005
R11889 gnd.n6174 gnd.n1166 9.3005
R11890 gnd.n6172 gnd.n6171 9.3005
R11891 gnd.n1170 gnd.n1169 9.3005
R11892 gnd.n4727 gnd.n4726 9.3005
R11893 gnd.n4729 gnd.n4728 9.3005
R11894 gnd.n4707 gnd.n4706 9.3005
R11895 gnd.n4735 gnd.n4734 9.3005
R11896 gnd.n4737 gnd.n4736 9.3005
R11897 gnd.n4697 gnd.n4696 9.3005
R11898 gnd.n4743 gnd.n4742 9.3005
R11899 gnd.n4745 gnd.n4744 9.3005
R11900 gnd.n4684 gnd.n4683 9.3005
R11901 gnd.n4751 gnd.n4750 9.3005
R11902 gnd.n4753 gnd.n4752 9.3005
R11903 gnd.n4674 gnd.n4673 9.3005
R11904 gnd.n4759 gnd.n4758 9.3005
R11905 gnd.n4761 gnd.n4760 9.3005
R11906 gnd.n4655 gnd.n4653 9.3005
R11907 gnd.n4767 gnd.n4766 9.3005
R11908 gnd.n4768 gnd.n4652 9.3005
R11909 gnd.n4661 gnd.n4660 9.3005
R11910 gnd.n4656 gnd.n4654 9.3005
R11911 gnd.n4765 gnd.n4764 9.3005
R11912 gnd.n4763 gnd.n4762 9.3005
R11913 gnd.n4669 gnd.n4668 9.3005
R11914 gnd.n4757 gnd.n4756 9.3005
R11915 gnd.n4755 gnd.n4754 9.3005
R11916 gnd.n4680 gnd.n4679 9.3005
R11917 gnd.n4749 gnd.n4748 9.3005
R11918 gnd.n4747 gnd.n4746 9.3005
R11919 gnd.n4691 gnd.n4690 9.3005
R11920 gnd.n4741 gnd.n4740 9.3005
R11921 gnd.n4739 gnd.n4738 9.3005
R11922 gnd.n4703 gnd.n4702 9.3005
R11923 gnd.n4733 gnd.n4732 9.3005
R11924 gnd.n4731 gnd.n4730 9.3005
R11925 gnd.n4716 gnd.n4715 9.3005
R11926 gnd.n4725 gnd.n4724 9.3005
R11927 gnd.n4786 gnd.n4785 9.3005
R11928 gnd.n4787 gnd.n1894 9.3005
R11929 gnd.n4789 gnd.n4788 9.3005
R11930 gnd.n1882 gnd.n1881 9.3005
R11931 gnd.n4805 gnd.n4804 9.3005
R11932 gnd.n4806 gnd.n1880 9.3005
R11933 gnd.n4808 gnd.n4807 9.3005
R11934 gnd.n1868 gnd.n1867 9.3005
R11935 gnd.n4824 gnd.n4823 9.3005
R11936 gnd.n4825 gnd.n1866 9.3005
R11937 gnd.n4827 gnd.n4826 9.3005
R11938 gnd.n1854 gnd.n1853 9.3005
R11939 gnd.n4843 gnd.n4842 9.3005
R11940 gnd.n4844 gnd.n1852 9.3005
R11941 gnd.n4846 gnd.n4845 9.3005
R11942 gnd.n1840 gnd.n1839 9.3005
R11943 gnd.n4862 gnd.n4861 9.3005
R11944 gnd.n4863 gnd.n1838 9.3005
R11945 gnd.n4865 gnd.n4864 9.3005
R11946 gnd.n1826 gnd.n1825 9.3005
R11947 gnd.n5081 gnd.n5080 9.3005
R11948 gnd.n5082 gnd.n1824 9.3005
R11949 gnd.n5084 gnd.n5083 9.3005
R11950 gnd.n1760 gnd.n1759 9.3005
R11951 gnd.n5115 gnd.n5114 9.3005
R11952 gnd.n5116 gnd.n1757 9.3005
R11953 gnd.n5119 gnd.n5118 9.3005
R11954 gnd.n5117 gnd.n1758 9.3005
R11955 gnd.n1731 gnd.n1730 9.3005
R11956 gnd.n5151 gnd.n5150 9.3005
R11957 gnd.n5152 gnd.n1729 9.3005
R11958 gnd.n5154 gnd.n5153 9.3005
R11959 gnd.n1711 gnd.n1710 9.3005
R11960 gnd.n5178 gnd.n5177 9.3005
R11961 gnd.n5179 gnd.n1708 9.3005
R11962 gnd.n5182 gnd.n5181 9.3005
R11963 gnd.n5180 gnd.n1709 9.3005
R11964 gnd.n1680 gnd.n1679 9.3005
R11965 gnd.n5216 gnd.n5215 9.3005
R11966 gnd.n5217 gnd.n1677 9.3005
R11967 gnd.n5220 gnd.n5219 9.3005
R11968 gnd.n5218 gnd.n1678 9.3005
R11969 gnd.n1648 gnd.n1647 9.3005
R11970 gnd.n5269 gnd.n5268 9.3005
R11971 gnd.n5270 gnd.n1646 9.3005
R11972 gnd.n5272 gnd.n5271 9.3005
R11973 gnd.n1631 gnd.n1630 9.3005
R11974 gnd.n5312 gnd.n5311 9.3005
R11975 gnd.n5313 gnd.n1628 9.3005
R11976 gnd.n5322 gnd.n5321 9.3005
R11977 gnd.n5320 gnd.n1629 9.3005
R11978 gnd.n5319 gnd.n5318 9.3005
R11979 gnd.n5317 gnd.n5314 9.3005
R11980 gnd.n1596 gnd.n1595 9.3005
R11981 gnd.n5380 gnd.n5379 9.3005
R11982 gnd.n5381 gnd.n1593 9.3005
R11983 gnd.n5387 gnd.n5386 9.3005
R11984 gnd.n5385 gnd.n1594 9.3005
R11985 gnd.n5384 gnd.n5383 9.3005
R11986 gnd.n1572 gnd.n1570 9.3005
R11987 gnd.n5429 gnd.n5428 9.3005
R11988 gnd.n5427 gnd.n1571 9.3005
R11989 gnd.n5426 gnd.n5425 9.3005
R11990 gnd.n1550 gnd.n1548 9.3005
R11991 gnd.n5479 gnd.n5478 9.3005
R11992 gnd.n5477 gnd.n1549 9.3005
R11993 gnd.n5476 gnd.n5475 9.3005
R11994 gnd.n1523 gnd.n1522 9.3005
R11995 gnd.n5509 gnd.n5508 9.3005
R11996 gnd.n5510 gnd.n1521 9.3005
R11997 gnd.n5512 gnd.n5511 9.3005
R11998 gnd.n1501 gnd.n1499 9.3005
R11999 gnd.n5558 gnd.n5557 9.3005
R12000 gnd.n5556 gnd.n1500 9.3005
R12001 gnd.n5555 gnd.n5554 9.3005
R12002 gnd.n5553 gnd.n1502 9.3005
R12003 gnd.n5552 gnd.n5551 9.3005
R12004 gnd.n1390 gnd.n1389 9.3005
R12005 gnd.n5728 gnd.n5727 9.3005
R12006 gnd.n5729 gnd.n1388 9.3005
R12007 gnd.n5731 gnd.n5730 9.3005
R12008 gnd.n1377 gnd.n1376 9.3005
R12009 gnd.n5747 gnd.n5746 9.3005
R12010 gnd.n5748 gnd.n1375 9.3005
R12011 gnd.n5750 gnd.n5749 9.3005
R12012 gnd.n1363 gnd.n1362 9.3005
R12013 gnd.n5766 gnd.n5765 9.3005
R12014 gnd.n5767 gnd.n1361 9.3005
R12015 gnd.n5769 gnd.n5768 9.3005
R12016 gnd.n1349 gnd.n1348 9.3005
R12017 gnd.n5785 gnd.n5784 9.3005
R12018 gnd.n5786 gnd.n1347 9.3005
R12019 gnd.n5788 gnd.n5787 9.3005
R12020 gnd.n1335 gnd.n1334 9.3005
R12021 gnd.n5804 gnd.n5803 9.3005
R12022 gnd.n5805 gnd.n1333 9.3005
R12023 gnd.n5807 gnd.n5806 9.3005
R12024 gnd.n1320 gnd.n1319 9.3005
R12025 gnd.n5996 gnd.n5995 9.3005
R12026 gnd.n5997 gnd.n1318 9.3005
R12027 gnd.n5999 gnd.n5998 9.3005
R12028 gnd.n1896 gnd.n1895 9.3005
R12029 gnd.n446 gnd.n445 9.3005
R12030 gnd.n7244 gnd.n7243 9.3005
R12031 gnd.n7245 gnd.n444 9.3005
R12032 gnd.n7247 gnd.n7246 9.3005
R12033 gnd.n428 gnd.n427 9.3005
R12034 gnd.n7260 gnd.n7259 9.3005
R12035 gnd.n7261 gnd.n426 9.3005
R12036 gnd.n7263 gnd.n7262 9.3005
R12037 gnd.n411 gnd.n410 9.3005
R12038 gnd.n7276 gnd.n7275 9.3005
R12039 gnd.n7277 gnd.n409 9.3005
R12040 gnd.n7279 gnd.n7278 9.3005
R12041 gnd.n394 gnd.n393 9.3005
R12042 gnd.n7292 gnd.n7291 9.3005
R12043 gnd.n7293 gnd.n392 9.3005
R12044 gnd.n7295 gnd.n7294 9.3005
R12045 gnd.n377 gnd.n376 9.3005
R12046 gnd.n7308 gnd.n7307 9.3005
R12047 gnd.n7309 gnd.n375 9.3005
R12048 gnd.n7311 gnd.n7310 9.3005
R12049 gnd.n360 gnd.n359 9.3005
R12050 gnd.n7324 gnd.n7323 9.3005
R12051 gnd.n7325 gnd.n358 9.3005
R12052 gnd.n7327 gnd.n7326 9.3005
R12053 gnd.n344 gnd.n343 9.3005
R12054 gnd.n7340 gnd.n7339 9.3005
R12055 gnd.n7341 gnd.n342 9.3005
R12056 gnd.n7343 gnd.n7342 9.3005
R12057 gnd.n328 gnd.n327 9.3005
R12058 gnd.n7356 gnd.n7355 9.3005
R12059 gnd.n7357 gnd.n325 9.3005
R12060 gnd.n7359 gnd.n7358 9.3005
R12061 gnd.n311 gnd.n310 9.3005
R12062 gnd.n7372 gnd.n7371 9.3005
R12063 gnd.n7373 gnd.n309 9.3005
R12064 gnd.n7375 gnd.n7374 9.3005
R12065 gnd.n297 gnd.n296 9.3005
R12066 gnd.n7388 gnd.n7387 9.3005
R12067 gnd.n7389 gnd.n295 9.3005
R12068 gnd.n7391 gnd.n7390 9.3005
R12069 gnd.n281 gnd.n280 9.3005
R12070 gnd.n7404 gnd.n7403 9.3005
R12071 gnd.n7405 gnd.n279 9.3005
R12072 gnd.n7407 gnd.n7406 9.3005
R12073 gnd.n267 gnd.n266 9.3005
R12074 gnd.n7420 gnd.n7419 9.3005
R12075 gnd.n7421 gnd.n265 9.3005
R12076 gnd.n7423 gnd.n7422 9.3005
R12077 gnd.n250 gnd.n249 9.3005
R12078 gnd.n7436 gnd.n7435 9.3005
R12079 gnd.n7437 gnd.n248 9.3005
R12080 gnd.n7439 gnd.n7438 9.3005
R12081 gnd.n236 gnd.n235 9.3005
R12082 gnd.n7452 gnd.n7451 9.3005
R12083 gnd.n7453 gnd.n234 9.3005
R12084 gnd.n7455 gnd.n7454 9.3005
R12085 gnd.n221 gnd.n220 9.3005
R12086 gnd.n7468 gnd.n7467 9.3005
R12087 gnd.n7469 gnd.n218 9.3005
R12088 gnd.n7539 gnd.n7538 9.3005
R12089 gnd.n7537 gnd.n219 9.3005
R12090 gnd.n7536 gnd.n7535 9.3005
R12091 gnd.n7534 gnd.n7470 9.3005
R12092 gnd.n7533 gnd.n7532 9.3005
R12093 gnd.n7231 gnd.n7230 9.3005
R12094 gnd.n7529 gnd.n7472 9.3005
R12095 gnd.n7528 gnd.n7527 9.3005
R12096 gnd.n7526 gnd.n7477 9.3005
R12097 gnd.n7525 gnd.n7524 9.3005
R12098 gnd.n7523 gnd.n7478 9.3005
R12099 gnd.n7522 gnd.n7521 9.3005
R12100 gnd.n7520 gnd.n7485 9.3005
R12101 gnd.n7519 gnd.n7518 9.3005
R12102 gnd.n7517 gnd.n7486 9.3005
R12103 gnd.n7516 gnd.n7515 9.3005
R12104 gnd.n7514 gnd.n7493 9.3005
R12105 gnd.n7513 gnd.n7512 9.3005
R12106 gnd.n7511 gnd.n7494 9.3005
R12107 gnd.n7510 gnd.n7509 9.3005
R12108 gnd.n7508 gnd.n7501 9.3005
R12109 gnd.n7507 gnd.n7506 9.3005
R12110 gnd.n124 gnd.n121 9.3005
R12111 gnd.n7633 gnd.n7632 9.3005
R12112 gnd.n7531 gnd.n7530 9.3005
R12113 gnd.n5971 gnd.n5970 9.3005
R12114 gnd.n596 gnd.n594 9.3005
R12115 gnd.n7096 gnd.n7095 9.3005
R12116 gnd.n7094 gnd.n595 9.3005
R12117 gnd.n7093 gnd.n7092 9.3005
R12118 gnd.n7091 gnd.n597 9.3005
R12119 gnd.n7090 gnd.n7089 9.3005
R12120 gnd.n7088 gnd.n600 9.3005
R12121 gnd.n7087 gnd.n7086 9.3005
R12122 gnd.n7085 gnd.n601 9.3005
R12123 gnd.n7084 gnd.n7083 9.3005
R12124 gnd.n7082 gnd.n604 9.3005
R12125 gnd.n7081 gnd.n7080 9.3005
R12126 gnd.n7079 gnd.n605 9.3005
R12127 gnd.n7078 gnd.n7077 9.3005
R12128 gnd.n7076 gnd.n608 9.3005
R12129 gnd.n7075 gnd.n7074 9.3005
R12130 gnd.n7073 gnd.n609 9.3005
R12131 gnd.n7072 gnd.n7071 9.3005
R12132 gnd.n7070 gnd.n7042 9.3005
R12133 gnd.n7069 gnd.n7068 9.3005
R12134 gnd.n7067 gnd.n7043 9.3005
R12135 gnd.n7066 gnd.n7065 9.3005
R12136 gnd.n7064 gnd.n7046 9.3005
R12137 gnd.n7063 gnd.n7062 9.3005
R12138 gnd.n7061 gnd.n7047 9.3005
R12139 gnd.n7060 gnd.n7059 9.3005
R12140 gnd.n7058 gnd.n7050 9.3005
R12141 gnd.n7057 gnd.n7056 9.3005
R12142 gnd.n7055 gnd.n7051 9.3005
R12143 gnd.n7054 gnd.n79 9.3005
R12144 gnd.n7682 gnd.n80 9.3005
R12145 gnd.n7681 gnd.n7680 9.3005
R12146 gnd.n7679 gnd.n81 9.3005
R12147 gnd.n7678 gnd.n7677 9.3005
R12148 gnd.n7676 gnd.n85 9.3005
R12149 gnd.n7675 gnd.n7674 9.3005
R12150 gnd.n7673 gnd.n86 9.3005
R12151 gnd.n7672 gnd.n7671 9.3005
R12152 gnd.n7670 gnd.n90 9.3005
R12153 gnd.n7669 gnd.n7668 9.3005
R12154 gnd.n7667 gnd.n91 9.3005
R12155 gnd.n7666 gnd.n7665 9.3005
R12156 gnd.n7664 gnd.n95 9.3005
R12157 gnd.n7663 gnd.n7662 9.3005
R12158 gnd.n7661 gnd.n96 9.3005
R12159 gnd.n7660 gnd.n7659 9.3005
R12160 gnd.n7658 gnd.n100 9.3005
R12161 gnd.n7657 gnd.n7656 9.3005
R12162 gnd.n7655 gnd.n101 9.3005
R12163 gnd.n7654 gnd.n7653 9.3005
R12164 gnd.n7652 gnd.n105 9.3005
R12165 gnd.n7651 gnd.n7650 9.3005
R12166 gnd.n7649 gnd.n106 9.3005
R12167 gnd.n7648 gnd.n7647 9.3005
R12168 gnd.n7646 gnd.n110 9.3005
R12169 gnd.n7645 gnd.n7644 9.3005
R12170 gnd.n7643 gnd.n111 9.3005
R12171 gnd.n7642 gnd.n7641 9.3005
R12172 gnd.n7640 gnd.n115 9.3005
R12173 gnd.n7639 gnd.n7638 9.3005
R12174 gnd.n7637 gnd.n116 9.3005
R12175 gnd.n7636 gnd.n7635 9.3005
R12176 gnd.n7634 gnd.n120 9.3005
R12177 gnd.n5969 gnd.n5931 9.3005
R12178 gnd.n2796 gnd.t300 9.29782
R12179 gnd.n2496 gnd.t158 9.29782
R12180 gnd.n3980 gnd.t2 9.24152
R12181 gnd.n5882 gnd.t121 9.24152
R12182 gnd.n263 gnd.t39 9.24152
R12183 gnd.n2787 gnd.t300 8.93321
R12184 gnd.t278 gnd.n2238 8.93321
R12185 gnd.t261 gnd.n2239 8.93321
R12186 gnd.n5129 gnd.n1747 8.92286
R12187 gnd.t232 gnd.n1738 8.92286
R12188 gnd.n5213 gnd.n5212 8.92286
R12189 gnd.n5258 gnd.n5257 8.92286
R12190 gnd.n5392 gnd.n1588 8.92286
R12191 gnd.n5442 gnd.n1561 8.92286
R12192 gnd.n5560 gnd.n1496 8.92286
R12193 gnd.n5725 gnd.n1392 8.92286
R12194 gnd.n3499 gnd.n3474 8.92171
R12195 gnd.n3467 gnd.n3442 8.92171
R12196 gnd.n3435 gnd.n3410 8.92171
R12197 gnd.n3404 gnd.n3379 8.92171
R12198 gnd.n3372 gnd.n3347 8.92171
R12199 gnd.n3340 gnd.n3315 8.92171
R12200 gnd.n3308 gnd.n3283 8.92171
R12201 gnd.n3277 gnd.n3252 8.92171
R12202 gnd.n1426 gnd.n1408 8.72777
R12203 gnd.n4579 gnd.t110 8.60421
R12204 gnd.n4782 gnd.t271 8.60421
R12205 gnd.t125 gnd.n1864 8.60421
R12206 gnd.n5773 gnd.t116 8.60421
R12207 gnd.t238 gnd.n5992 8.60421
R12208 gnd.n5870 gnd.t27 8.60421
R12209 gnd.n232 gnd.t119 8.60421
R12210 gnd.n3155 gnd.t79 8.56861
R12211 gnd.n2427 gnd.n2407 8.43467
R12212 gnd.n58 gnd.n38 8.43467
R12213 gnd.n4008 gnd.n0 8.41456
R12214 gnd.n7683 gnd.n7682 8.41456
R12215 gnd.n3962 gnd.n983 8.28555
R12216 gnd.n6309 gnd.n993 8.28555
R12217 gnd.n3967 gnd.n3966 8.28555
R12218 gnd.n6303 gnd.n1004 8.28555
R12219 gnd.n3980 gnd.n1007 8.28555
R12220 gnd.n6297 gnd.n1015 8.28555
R12221 gnd.n4563 gnd.n1018 8.28555
R12222 gnd.n4571 gnd.n1028 8.28555
R12223 gnd.n6285 gnd.n1036 8.28555
R12224 gnd.n4607 gnd.n4606 8.28555
R12225 gnd.n6279 gnd.n1046 8.28555
R12226 gnd.n4579 gnd.n1049 8.28555
R12227 gnd.n6273 gnd.n1057 8.28555
R12228 gnd.n4583 gnd.n1060 8.28555
R12229 gnd.n6267 gnd.n1068 8.28555
R12230 gnd.n4592 gnd.n1071 8.28555
R12231 gnd.n6261 gnd.n1079 8.28555
R12232 gnd.n6178 gnd.n1164 8.28555
R12233 gnd.n6255 gnd.n1088 8.28555
R12234 gnd.t307 gnd.n5105 8.28555
R12235 gnd.n1782 gnd.n1688 8.28555
R12236 gnd.n5293 gnd.n1639 8.28555
R12237 gnd.n5350 gnd.n5349 8.28555
R12238 gnd.n5452 gnd.n5451 8.28555
R12239 gnd.n5549 gnd.t288 8.28555
R12240 gnd.n7233 gnd.n458 8.28555
R12241 gnd.n5974 gnd.n5973 8.28555
R12242 gnd.n7241 gnd.n450 8.28555
R12243 gnd.n7098 gnd.n439 8.28555
R12244 gnd.n7249 gnd.n442 8.28555
R12245 gnd.n5866 gnd.n430 8.28555
R12246 gnd.n7257 gnd.n433 8.28555
R12247 gnd.n5870 gnd.n421 8.28555
R12248 gnd.n7265 gnd.n424 8.28555
R12249 gnd.n5918 gnd.n5917 8.28555
R12250 gnd.n7273 gnd.n415 8.28555
R12251 gnd.n5911 gnd.n405 8.28555
R12252 gnd.n5907 gnd.n396 8.28555
R12253 gnd.n7289 gnd.n399 8.28555
R12254 gnd.n5882 gnd.n387 8.28555
R12255 gnd.n7297 gnd.n390 8.28555
R12256 gnd.n6928 gnd.n6927 8.28555
R12257 gnd.n7305 gnd.n381 8.28555
R12258 gnd.n7040 gnd.n371 8.28555
R12259 gnd.t90 gnd.n2281 8.20401
R12260 gnd.n3233 gnd.t167 8.20401
R12261 gnd.n3500 gnd.n3472 8.14595
R12262 gnd.n3468 gnd.n3440 8.14595
R12263 gnd.n3436 gnd.n3408 8.14595
R12264 gnd.n3405 gnd.n3377 8.14595
R12265 gnd.n3373 gnd.n3345 8.14595
R12266 gnd.n3341 gnd.n3313 8.14595
R12267 gnd.n3309 gnd.n3281 8.14595
R12268 gnd.n3278 gnd.n3250 8.14595
R12269 gnd.n3505 gnd.n3504 7.97301
R12270 gnd.n4773 gnd.n4771 7.9669
R12271 gnd.n5985 gnd.n5984 7.9669
R12272 gnd.n2943 gnd.t335 7.83941
R12273 gnd.n7632 gnd.n124 7.75808
R12274 gnd.n7180 gnd.n504 7.75808
R12275 gnd.n4724 gnd.n4715 7.75808
R12276 gnd.n4062 gnd.n3661 7.75808
R12277 gnd.n2861 gnd.n2599 7.65711
R12278 gnd.n1782 gnd.n1698 7.64824
R12279 gnd.n1654 gnd.t14 7.64824
R12280 gnd.n5275 gnd.t128 7.64824
R12281 gnd.n5293 gnd.n5292 7.64824
R12282 gnd.n5350 gnd.n1608 7.64824
R12283 gnd.t24 gnd.n1598 7.64824
R12284 gnd.n5391 gnd.t83 7.64824
R12285 gnd.n5452 gnd.n1544 7.64824
R12286 gnd.n5577 gnd.t254 7.64824
R12287 gnd.t271 gnd.n1890 7.32958
R12288 gnd.n4829 gnd.t125 7.32958
R12289 gnd.t116 gnd.n5772 7.32958
R12290 gnd.n5993 gnd.t238 7.32958
R12291 gnd.n6920 gnd.t88 7.32958
R12292 gnd.n4934 gnd.n4933 7.30353
R12293 gnd.n1425 gnd.n1424 7.30353
R12294 gnd.n2129 gnd.t31 7.11021
R12295 gnd.n5088 gnd.n1820 7.01093
R12296 gnd.n5130 gnd.n5129 7.01093
R12297 gnd.n1807 gnd.t232 7.01093
R12298 gnd.n5212 gnd.n1684 7.01093
R12299 gnd.n5265 gnd.t14 7.01093
R12300 gnd.n5257 gnd.n1654 7.01093
R12301 gnd.n5392 gnd.n5391 7.01093
R12302 gnd.t83 gnd.n5390 7.01093
R12303 gnd.n5443 gnd.n5442 7.01093
R12304 gnd.n1404 gnd.n1392 7.01093
R12305 gnd.n2097 gnd.t4 6.74561
R12306 gnd.n4562 gnd.t25 6.69227
R12307 gnd.n5140 gnd.t20 6.69227
R12308 gnd.n5530 gnd.t123 6.69227
R12309 gnd.n5906 gnd.t66 6.69227
R12310 gnd.n5643 gnd.n5642 6.5566
R12311 gnd.n5005 gnd.n5004 6.5566
R12312 gnd.n5018 gnd.n4940 6.5566
R12313 gnd.n5658 gnd.n5657 6.5566
R12314 gnd.n2931 gnd.t335 6.38101
R12315 gnd.n2065 gnd.t140 6.38101
R12316 gnd.t6 gnd.n1996 6.38101
R12317 gnd.t235 gnd.n1820 6.37362
R12318 gnd.n5187 gnd.n1703 6.37362
R12319 gnd.n5230 gnd.t95 6.37362
R12320 gnd.n5285 gnd.n5284 6.37362
R12321 gnd.n5358 gnd.n1613 6.37362
R12322 gnd.t23 gnd.n1576 6.37362
R12323 gnd.n5489 gnd.n1540 6.37362
R12324 gnd.n6160 gnd.n1181 6.20656
R12325 gnd.n7594 gnd.n7591 6.20656
R12326 gnd.n3758 gnd.n3753 6.20656
R12327 gnd.n5958 gnd.n5955 6.20656
R12328 gnd.n6317 gnd.n979 6.19871
R12329 gnd.t127 gnd.t182 6.05496
R12330 gnd.t137 gnd.t135 6.05496
R12331 gnd.n2850 gnd.t8 6.01641
R12332 gnd.n2283 gnd.t90 6.01641
R12333 gnd.n3216 gnd.t167 6.01641
R12334 gnd.t98 gnd.n2029 6.01641
R12335 gnd.n2032 gnd.t64 6.01641
R12336 gnd.n3502 gnd.n3472 5.81868
R12337 gnd.n3470 gnd.n3440 5.81868
R12338 gnd.n3438 gnd.n3408 5.81868
R12339 gnd.n3407 gnd.n3377 5.81868
R12340 gnd.n3375 gnd.n3345 5.81868
R12341 gnd.n3343 gnd.n3313 5.81868
R12342 gnd.n3311 gnd.n3281 5.81868
R12343 gnd.n3280 gnd.n3250 5.81868
R12344 gnd.n5104 gnd.n1762 5.73631
R12345 gnd.n5231 gnd.n1665 5.73631
R12346 gnd.n1670 gnd.n1669 5.73631
R12347 gnd.t128 gnd.n1639 5.73631
R12348 gnd.n5349 gnd.t24 5.73631
R12349 gnd.n5340 gnd.n5339 5.73631
R12350 gnd.n5411 gnd.n5410 5.73631
R12351 gnd.n5583 gnd.n1479 5.73631
R12352 gnd.t79 gnd.n2300 5.65181
R12353 gnd.t51 gnd.n2062 5.65181
R12354 gnd.n1999 gnd.t33 5.65181
R12355 gnd.n1452 gnd.n561 5.62001
R12356 gnd.n5013 gnd.n5009 5.62001
R12357 gnd.n5014 gnd.n5013 5.62001
R12358 gnd.n5652 gnd.n561 5.62001
R12359 gnd.n2731 gnd.n2726 5.4308
R12360 gnd.n3547 gnd.n2224 5.4308
R12361 gnd.t224 gnd.n5174 5.41765
R12362 gnd.t131 gnd.n5471 5.41765
R12363 gnd.t77 gnd.n2347 5.28721
R12364 gnd.n2249 gnd.t278 5.28721
R12365 gnd.n3529 gnd.t261 5.28721
R12366 gnd.t70 gnd.n2094 5.28721
R12367 gnd.t114 gnd.t77 5.10491
R12368 gnd.n5148 gnd.t337 5.09899
R12369 gnd.n5165 gnd.n5164 5.09899
R12370 gnd.n5324 gnd.n1625 5.09899
R12371 gnd.n5300 gnd.n1618 5.09899
R12372 gnd.n1532 gnd.n1531 5.09899
R12373 gnd.t22 gnd.n5514 5.09899
R12374 gnd.n3500 gnd.n3499 5.04292
R12375 gnd.n3468 gnd.n3467 5.04292
R12376 gnd.n3436 gnd.n3435 5.04292
R12377 gnd.n3405 gnd.n3404 5.04292
R12378 gnd.n3373 gnd.n3372 5.04292
R12379 gnd.n3341 gnd.n3340 5.04292
R12380 gnd.n3309 gnd.n3308 5.04292
R12381 gnd.n3278 gnd.n3277 5.04292
R12382 gnd.n3003 gnd.t158 4.92261
R12383 gnd.t142 gnd.n2126 4.92261
R12384 gnd.n2447 gnd.n2446 4.82753
R12385 gnd.n78 gnd.n77 4.82753
R12386 gnd.t357 gnd.n1842 4.78034
R12387 gnd.t220 gnd.n5752 4.78034
R12388 gnd.n2452 gnd.n2449 4.74817
R12389 gnd.n2502 gnd.n2388 4.74817
R12390 gnd.n2489 gnd.n2387 4.74817
R12391 gnd.n2386 gnd.n2385 4.74817
R12392 gnd.n2498 gnd.n2449 4.74817
R12393 gnd.n2499 gnd.n2388 4.74817
R12394 gnd.n2501 gnd.n2387 4.74817
R12395 gnd.n2488 gnd.n2386 4.74817
R12396 gnd.n2427 gnd.n2426 4.7074
R12397 gnd.n58 gnd.n57 4.7074
R12398 gnd.n2447 gnd.n2427 4.65959
R12399 gnd.n78 gnd.n58 4.65959
R12400 gnd.n6317 gnd.n6316 4.63942
R12401 gnd.n7147 gnd.n563 4.6132
R12402 gnd.n1125 gnd.n1122 4.6132
R12403 gnd.t157 gnd.n2518 4.55801
R12404 gnd.n5106 gnd.n1767 4.46168
R12405 gnd.n5123 gnd.n5122 4.46168
R12406 gnd.n1774 gnd.t200 4.46168
R12407 gnd.n5223 gnd.n1674 4.46168
R12408 gnd.n5251 gnd.n5250 4.46168
R12409 gnd.n5402 gnd.n5401 4.46168
R12410 gnd.n5433 gnd.n5432 4.46168
R12411 gnd.t201 gnd.n5431 4.46168
R12412 gnd.n1496 gnd.t275 4.46168
R12413 gnd.n5543 gnd.n1503 4.46168
R12414 gnd.n5716 gnd.n1402 4.46168
R12415 gnd.n1421 gnd.n1408 4.46111
R12416 gnd.n3485 gnd.n3481 4.38594
R12417 gnd.n3453 gnd.n3449 4.38594
R12418 gnd.n3421 gnd.n3417 4.38594
R12419 gnd.n3390 gnd.n3386 4.38594
R12420 gnd.n3358 gnd.n3354 4.38594
R12421 gnd.n3326 gnd.n3322 4.38594
R12422 gnd.n3294 gnd.n3290 4.38594
R12423 gnd.n3263 gnd.n3259 4.38594
R12424 gnd.n3496 gnd.n3474 4.26717
R12425 gnd.n3464 gnd.n3442 4.26717
R12426 gnd.n3432 gnd.n3410 4.26717
R12427 gnd.n3401 gnd.n3379 4.26717
R12428 gnd.n3369 gnd.n3347 4.26717
R12429 gnd.n3337 gnd.n3315 4.26717
R12430 gnd.n3305 gnd.n3283 4.26717
R12431 gnd.n3274 gnd.n3252 4.26717
R12432 gnd.n2912 gnd.t82 4.19341
R12433 gnd.n4607 gnd.t96 4.14303
R12434 gnd.n5918 gnd.t59 4.14303
R12435 gnd.n3504 gnd.n3503 4.08274
R12436 gnd.n5642 gnd.n5641 4.05904
R12437 gnd.n5004 gnd.n5003 4.05904
R12438 gnd.n5021 gnd.n4940 4.05904
R12439 gnd.n5659 gnd.n5658 4.05904
R12440 gnd.n2872 gnd.n2591 4.01111
R12441 gnd.n2594 gnd.n2592 4.01111
R12442 gnd.n2882 gnd.n2881 4.01111
R12443 gnd.n2893 gnd.n2575 4.01111
R12444 gnd.n2892 gnd.n2578 4.01111
R12445 gnd.n2903 gnd.n2566 4.01111
R12446 gnd.n2569 gnd.n2567 4.01111
R12447 gnd.n2913 gnd.n2912 4.01111
R12448 gnd.n2923 gnd.n2547 4.01111
R12449 gnd.n2922 gnd.n2550 4.01111
R12450 gnd.n2931 gnd.n2541 4.01111
R12451 gnd.n2943 gnd.n2531 4.01111
R12452 gnd.n2953 gnd.n2516 4.01111
R12453 gnd.n2969 gnd.n2968 4.01111
R12454 gnd.n2518 gnd.n2455 4.01111
R12455 gnd.n3023 gnd.n2456 4.01111
R12456 gnd.n3017 gnd.n3016 4.01111
R12457 gnd.n2505 gnd.n2467 4.01111
R12458 gnd.n3009 gnd.n2478 4.01111
R12459 gnd.n2496 gnd.n2491 4.01111
R12460 gnd.n3003 gnd.n3002 4.01111
R12461 gnd.n3049 gnd.n2382 4.01111
R12462 gnd.n3048 gnd.n3047 4.01111
R12463 gnd.n3060 gnd.n3059 4.01111
R12464 gnd.n2375 gnd.n2367 4.01111
R12465 gnd.n3089 gnd.n2355 4.01111
R12466 gnd.n3088 gnd.n2358 4.01111
R12467 gnd.n3099 gnd.n2347 4.01111
R12468 gnd.n2348 gnd.n2336 4.01111
R12469 gnd.n3110 gnd.n2337 4.01111
R12470 gnd.n3134 gnd.n2328 4.01111
R12471 gnd.n3133 gnd.n2319 4.01111
R12472 gnd.n3156 gnd.n3155 4.01111
R12473 gnd.n3174 gnd.n2300 4.01111
R12474 gnd.n3173 gnd.n2303 4.01111
R12475 gnd.n3184 gnd.n2292 4.01111
R12476 gnd.n2293 gnd.n2280 4.01111
R12477 gnd.n3195 gnd.n2281 4.01111
R12478 gnd.n3222 gnd.n2265 4.01111
R12479 gnd.n3234 gnd.n3233 4.01111
R12480 gnd.n3216 gnd.n2258 4.01111
R12481 gnd.n3245 gnd.n3244 4.01111
R12482 gnd.n3517 gnd.n2246 4.01111
R12483 gnd.n3516 gnd.n2249 4.01111
R12484 gnd.n3529 gnd.n2238 4.01111
R12485 gnd.n2239 gnd.n2231 4.01111
R12486 gnd.n3539 gnd.n2157 4.01111
R12487 gnd.n19 gnd.n9 3.99943
R12488 gnd.n2550 gnd.t163 3.82881
R12489 gnd.n2358 gnd.t114 3.82881
R12490 gnd.n3223 gnd.t159 3.82881
R12491 gnd.n1904 gnd.n1096 3.82437
R12492 gnd.n1799 gnd.n1798 3.82437
R12493 gnd.n1790 gnd.t129 3.82437
R12494 gnd.n5185 gnd.n5184 3.82437
R12495 gnd.n5309 gnd.n5308 3.82437
R12496 gnd.n5283 gnd.t127 3.82437
R12497 gnd.n5357 gnd.t137 3.82437
R12498 gnd.n5356 gnd.n1606 3.82437
R12499 gnd.n5481 gnd.n1538 3.82437
R12500 gnd.n5499 gnd.t0 3.82437
R12501 gnd.n5521 gnd.n1513 3.82437
R12502 gnd.n7178 gnd.n511 3.82437
R12503 gnd.n3504 gnd.n3376 3.70378
R12504 gnd.n3027 gnd.n2448 3.65935
R12505 gnd.n19 gnd.n18 3.60163
R12506 gnd.n3966 gnd.t170 3.50571
R12507 gnd.n6261 gnd.t242 3.50571
R12508 gnd.n4811 gnd.t133 3.50571
R12509 gnd.t198 gnd.n1337 3.50571
R12510 gnd.n7241 gnd.t246 3.50571
R12511 gnd.n6927 gnd.t189 3.50571
R12512 gnd.n7549 gnd.t228 3.50571
R12513 gnd.n3495 gnd.n3476 3.49141
R12514 gnd.n3463 gnd.n3444 3.49141
R12515 gnd.n3431 gnd.n3412 3.49141
R12516 gnd.n3400 gnd.n3381 3.49141
R12517 gnd.n3368 gnd.n3349 3.49141
R12518 gnd.n3336 gnd.n3317 3.49141
R12519 gnd.n3304 gnd.n3285 3.49141
R12520 gnd.n3273 gnd.n3254 3.49141
R12521 gnd.t160 gnd.n2979 3.46421
R12522 gnd.n2980 gnd.t80 3.46421
R12523 gnd.t164 gnd.n2382 3.46421
R12524 gnd.t168 gnd.n3144 3.46421
R12525 gnd.n5106 gnd.t307 3.18706
R12526 gnd.n5097 gnd.t333 3.18706
R12527 gnd.t250 gnd.n5097 3.18706
R12528 gnd.n1808 gnd.n1807 3.18706
R12529 gnd.n5157 gnd.t57 3.18706
R12530 gnd.t57 gnd.n5156 3.18706
R12531 gnd.n5204 gnd.n1690 3.18706
R12532 gnd.n5259 gnd.n1644 3.18706
R12533 gnd.n5376 gnd.n1600 3.18706
R12534 gnd.n5421 gnd.n5420 3.18706
R12535 gnd.n5506 gnd.t17 3.18706
R12536 gnd.t17 gnd.n1511 3.18706
R12537 gnd.n5561 gnd.n1494 3.18706
R12538 gnd.t257 gnd.n5576 3.18706
R12539 gnd.t265 gnd.n1404 3.18706
R12540 gnd.n3047 gnd.t156 3.0996
R12541 gnd.t166 gnd.n3070 3.0996
R12542 gnd.t37 gnd.n2312 3.0996
R12543 gnd.n5078 gnd.n5077 2.8684
R12544 gnd.n5112 gnd.t92 2.8684
R12545 gnd.n5547 gnd.t355 2.8684
R12546 gnd.n1396 gnd.n1395 2.8684
R12547 gnd.n7433 gnd.n252 2.8684
R12548 gnd.n2428 gnd.t113 2.82907
R12549 gnd.n2428 gnd.t107 2.82907
R12550 gnd.n2430 gnd.t204 2.82907
R12551 gnd.n2430 gnd.t153 2.82907
R12552 gnd.n2432 gnd.t34 2.82907
R12553 gnd.n2432 gnd.t36 2.82907
R12554 gnd.n2434 gnd.t109 2.82907
R12555 gnd.n2434 gnd.t104 2.82907
R12556 gnd.n2436 gnd.t202 2.82907
R12557 gnd.n2436 gnd.t149 2.82907
R12558 gnd.n2438 gnd.t203 2.82907
R12559 gnd.n2438 gnd.t106 2.82907
R12560 gnd.n2440 gnd.t103 2.82907
R12561 gnd.n2440 gnd.t211 2.82907
R12562 gnd.n2442 gnd.t112 2.82907
R12563 gnd.n2442 gnd.t148 2.82907
R12564 gnd.n2444 gnd.t177 2.82907
R12565 gnd.n2444 gnd.t206 2.82907
R12566 gnd.n2389 gnd.t26 2.82907
R12567 gnd.n2389 gnd.t214 2.82907
R12568 gnd.n2391 gnd.t339 2.82907
R12569 gnd.n2391 gnd.t3 2.82907
R12570 gnd.n2393 gnd.t87 2.82907
R12571 gnd.n2393 gnd.t139 2.82907
R12572 gnd.n2395 gnd.t169 2.82907
R12573 gnd.n2395 gnd.t7 2.82907
R12574 gnd.n2397 gnd.t99 2.82907
R12575 gnd.n2397 gnd.t65 2.82907
R12576 gnd.n2399 gnd.t141 2.82907
R12577 gnd.n2399 gnd.t174 2.82907
R12578 gnd.n2401 gnd.t216 2.82907
R12579 gnd.n2401 gnd.t349 2.82907
R12580 gnd.n2403 gnd.t185 2.82907
R12581 gnd.n2403 gnd.t5 2.82907
R12582 gnd.n2405 gnd.t215 2.82907
R12583 gnd.n2405 gnd.t61 2.82907
R12584 gnd.n2408 gnd.t217 2.82907
R12585 gnd.n2408 gnd.t97 2.82907
R12586 gnd.n2410 gnd.t171 2.82907
R12587 gnd.n2410 gnd.t340 2.82907
R12588 gnd.n2412 gnd.t193 2.82907
R12589 gnd.n2412 gnd.t86 2.82907
R12590 gnd.n2414 gnd.t54 2.82907
R12591 gnd.n2414 gnd.t147 2.82907
R12592 gnd.n2416 gnd.t194 2.82907
R12593 gnd.n2416 gnd.t218 2.82907
R12594 gnd.n2418 gnd.t213 2.82907
R12595 gnd.n2418 gnd.t184 2.82907
R12596 gnd.n2420 gnd.t186 2.82907
R12597 gnd.n2420 gnd.t52 2.82907
R12598 gnd.n2422 gnd.t71 2.82907
R12599 gnd.n2422 gnd.t350 2.82907
R12600 gnd.n2424 gnd.t32 2.82907
R12601 gnd.n2424 gnd.t56 2.82907
R12602 gnd.n75 gnd.t179 2.82907
R12603 gnd.n75 gnd.t151 2.82907
R12604 gnd.n73 gnd.t46 2.82907
R12605 gnd.n73 gnd.t205 2.82907
R12606 gnd.n71 gnd.t101 2.82907
R12607 gnd.n71 gnd.t172 2.82907
R12608 gnd.n69 gnd.t154 2.82907
R12609 gnd.n69 gnd.t152 2.82907
R12610 gnd.n67 gnd.t108 2.82907
R12611 gnd.n67 gnd.t63 2.82907
R12612 gnd.n65 gnd.t208 2.82907
R12613 gnd.n65 gnd.t155 2.82907
R12614 gnd.n63 gnd.t89 2.82907
R12615 gnd.n63 gnd.t223 2.82907
R12616 gnd.n61 gnd.t210 2.82907
R12617 gnd.n61 gnd.t207 2.82907
R12618 gnd.n59 gnd.t173 2.82907
R12619 gnd.n59 gnd.t150 2.82907
R12620 gnd.n36 gnd.t341 2.82907
R12621 gnd.n36 gnd.t85 2.82907
R12622 gnd.n34 gnd.t346 2.82907
R12623 gnd.n34 gnd.t40 2.82907
R12624 gnd.n32 gnd.t145 2.82907
R12625 gnd.n32 gnd.t44 2.82907
R12626 gnd.n30 gnd.t16 2.82907
R12627 gnd.n30 gnd.t30 2.82907
R12628 gnd.n28 gnd.t58 2.82907
R12629 gnd.n28 gnd.t11 2.82907
R12630 gnd.n26 gnd.t195 2.82907
R12631 gnd.n26 gnd.t146 2.82907
R12632 gnd.n24 gnd.t338 2.82907
R12633 gnd.n24 gnd.t84 2.82907
R12634 gnd.n22 gnd.t345 2.82907
R12635 gnd.n22 gnd.t190 2.82907
R12636 gnd.n20 gnd.t188 2.82907
R12637 gnd.n20 gnd.t67 2.82907
R12638 gnd.n55 gnd.t359 2.82907
R12639 gnd.n55 gnd.t75 2.82907
R12640 gnd.n53 gnd.t191 2.82907
R12641 gnd.n53 gnd.t342 2.82907
R12642 gnd.n51 gnd.t175 2.82907
R12643 gnd.n51 gnd.t222 2.82907
R12644 gnd.n49 gnd.t344 2.82907
R12645 gnd.n49 gnd.t187 2.82907
R12646 gnd.n47 gnd.t13 2.82907
R12647 gnd.n47 gnd.t192 2.82907
R12648 gnd.n45 gnd.t42 2.82907
R12649 gnd.n45 gnd.t69 2.82907
R12650 gnd.n43 gnd.t212 2.82907
R12651 gnd.n43 gnd.t73 2.82907
R12652 gnd.n41 gnd.t122 2.82907
R12653 gnd.n41 gnd.t343 2.82907
R12654 gnd.n39 gnd.t60 2.82907
R12655 gnd.n39 gnd.t138 2.82907
R12656 gnd.n3010 gnd.t81 2.735
R12657 gnd.n2337 gnd.t78 2.735
R12658 gnd.n3492 gnd.n3491 2.71565
R12659 gnd.n3460 gnd.n3459 2.71565
R12660 gnd.n3428 gnd.n3427 2.71565
R12661 gnd.n3397 gnd.n3396 2.71565
R12662 gnd.n3365 gnd.n3364 2.71565
R12663 gnd.n3333 gnd.n3332 2.71565
R12664 gnd.n3301 gnd.n3300 2.71565
R12665 gnd.n3270 gnd.n3269 2.71565
R12666 gnd.n6316 gnd.t35 2.66809
R12667 gnd.n4911 gnd.t235 2.54975
R12668 gnd.n5098 gnd.t250 2.54975
R12669 gnd.n5141 gnd.n1738 2.54975
R12670 gnd.n1803 gnd.t337 2.54975
R12671 gnd.n5206 gnd.n5205 2.54975
R12672 gnd.n5205 gnd.t1 2.54975
R12673 gnd.n5275 gnd.n5274 2.54975
R12674 gnd.n5377 gnd.n1598 2.54975
R12675 gnd.n5423 gnd.t130 2.54975
R12676 gnd.n5423 gnd.n1553 2.54975
R12677 gnd.n5515 gnd.t22 2.54975
R12678 gnd.n5532 gnd.n5531 2.54975
R12679 gnd.n5568 gnd.t275 2.54975
R12680 gnd.n5545 gnd.t254 2.54975
R12681 gnd.n5577 gnd.t257 2.54975
R12682 gnd.n2954 gnd.t76 2.3704
R12683 gnd.n3184 gnd.t162 2.3704
R12684 gnd.n3027 gnd.n2449 2.27742
R12685 gnd.n3027 gnd.n2388 2.27742
R12686 gnd.n3027 gnd.n2387 2.27742
R12687 gnd.n3027 gnd.n2386 2.27742
R12688 gnd.n5250 gnd.t347 2.23109
R12689 gnd.n5308 gnd.t182 2.23109
R12690 gnd.t135 gnd.n5356 2.23109
R12691 gnd.n5402 gnd.t18 2.23109
R12692 gnd.n7321 gnd.n365 2.23109
R12693 gnd.n4111 gnd.t310 2.0058
R12694 gnd.n3488 gnd.n3478 1.93989
R12695 gnd.n3456 gnd.n3446 1.93989
R12696 gnd.n3424 gnd.n3414 1.93989
R12697 gnd.n3393 gnd.n3383 1.93989
R12698 gnd.n3361 gnd.n3351 1.93989
R12699 gnd.n3329 gnd.n3319 1.93989
R12700 gnd.n3297 gnd.n3287 1.93989
R12701 gnd.n3266 gnd.n3256 1.93989
R12702 gnd.n5147 gnd.n1734 1.91244
R12703 gnd.n5194 gnd.n5193 1.91244
R12704 gnd.n5291 gnd.n1633 1.91244
R12705 gnd.n5368 gnd.n5367 1.91244
R12706 gnd.n5483 gnd.n5482 1.91244
R12707 gnd.n1518 gnd.n1517 1.91244
R12708 gnd.n5583 gnd.t288 1.91244
R12709 gnd.n1395 gnd.t291 1.91244
R12710 gnd.n2533 gnd.t76 1.6412
R12711 gnd.n6291 gnd.t25 1.59378
R12712 gnd.n1803 gnd.t20 1.59378
R12713 gnd.n5213 gnd.t196 1.59378
R12714 gnd.t49 gnd.n1561 1.59378
R12715 gnd.n5515 gnd.t123 1.59378
R12716 gnd.n7281 gnd.t66 1.59378
R12717 gnd.n7441 gnd.t178 1.59378
R12718 gnd.n2881 gnd.t317 1.2766
R12719 gnd.n2504 gnd.t81 1.2766
R12720 gnd.n4533 gnd.n4282 1.2766
R12721 gnd.n5087 gnd.n5086 1.27512
R12722 gnd.n5121 gnd.n1754 1.27512
R12723 gnd.n5175 gnd.t129 1.27512
R12724 gnd.n1775 gnd.n1774 1.27512
R12725 gnd.n5266 gnd.n5265 1.27512
R12726 gnd.n5390 gnd.n5389 1.27512
R12727 gnd.n5431 gnd.n1559 1.27512
R12728 gnd.n5473 gnd.t0 1.27512
R12729 gnd.n5567 gnd.n1490 1.27512
R12730 gnd.n5715 gnd.n5714 1.27512
R12731 gnd.n2734 gnd.n2726 1.16414
R12732 gnd.n3550 gnd.n2224 1.16414
R12733 gnd.n3487 gnd.n3480 1.16414
R12734 gnd.n3455 gnd.n3448 1.16414
R12735 gnd.n3423 gnd.n3416 1.16414
R12736 gnd.n3392 gnd.n3385 1.16414
R12737 gnd.n3360 gnd.n3353 1.16414
R12738 gnd.n3328 gnd.n3321 1.16414
R12739 gnd.n3296 gnd.n3289 1.16414
R12740 gnd.n3265 gnd.n3258 1.16414
R12741 gnd.n7147 gnd.n7146 0.970197
R12742 gnd.n6219 gnd.n1122 0.970197
R12743 gnd.n3471 gnd.n3439 0.962709
R12744 gnd.n3503 gnd.n3471 0.962709
R12745 gnd.n3344 gnd.n3312 0.962709
R12746 gnd.n3376 gnd.n3344 0.962709
R12747 gnd.t35 gnd.n6315 0.956468
R12748 gnd.n4878 gnd.t47 0.956468
R12749 gnd.n1394 gnd.t353 0.956468
R12750 gnd.n7313 gnd.t88 0.956468
R12751 gnd.n7409 gnd.t43 0.956468
R12752 gnd.t180 gnd.n2892 0.912001
R12753 gnd.n3071 gnd.t166 0.912001
R12754 gnd.n2321 gnd.t37 0.912001
R12755 gnd.n4151 gnd.t55 0.912001
R12756 gnd.n2439 gnd.n2437 0.773756
R12757 gnd.n70 gnd.n68 0.773756
R12758 gnd.n2446 gnd.n2445 0.773756
R12759 gnd.n2445 gnd.n2443 0.773756
R12760 gnd.n2443 gnd.n2441 0.773756
R12761 gnd.n2441 gnd.n2439 0.773756
R12762 gnd.n2437 gnd.n2435 0.773756
R12763 gnd.n2435 gnd.n2433 0.773756
R12764 gnd.n2433 gnd.n2431 0.773756
R12765 gnd.n2431 gnd.n2429 0.773756
R12766 gnd.n62 gnd.n60 0.773756
R12767 gnd.n64 gnd.n62 0.773756
R12768 gnd.n66 gnd.n64 0.773756
R12769 gnd.n68 gnd.n66 0.773756
R12770 gnd.n72 gnd.n70 0.773756
R12771 gnd.n74 gnd.n72 0.773756
R12772 gnd.n76 gnd.n74 0.773756
R12773 gnd.n77 gnd.n76 0.773756
R12774 gnd gnd.n0 0.70738
R12775 gnd.n2 gnd.n1 0.672012
R12776 gnd.n3 gnd.n2 0.672012
R12777 gnd.n4 gnd.n3 0.672012
R12778 gnd.n5 gnd.n4 0.672012
R12779 gnd.n6 gnd.n5 0.672012
R12780 gnd.n7 gnd.n6 0.672012
R12781 gnd.n8 gnd.n7 0.672012
R12782 gnd.n9 gnd.n8 0.672012
R12783 gnd.n11 gnd.n10 0.672012
R12784 gnd.n12 gnd.n11 0.672012
R12785 gnd.n13 gnd.n12 0.672012
R12786 gnd.n14 gnd.n13 0.672012
R12787 gnd.n15 gnd.n14 0.672012
R12788 gnd.n16 gnd.n15 0.672012
R12789 gnd.n17 gnd.n16 0.672012
R12790 gnd.n18 gnd.n17 0.672012
R12791 gnd.n1754 gnd.t282 0.637812
R12792 gnd.n5166 gnd.n1719 0.637812
R12793 gnd.n5174 gnd.n1713 0.637812
R12794 gnd.n5184 gnd.t118 0.637812
R12795 gnd.n5325 gnd.n1624 0.637812
R12796 gnd.n5334 gnd.n5333 0.637812
R12797 gnd.t94 gnd.n5481 0.637812
R12798 gnd.n5471 gnd.n5470 0.637812
R12799 gnd.n5505 gnd.n1525 0.637812
R12800 gnd.n7684 gnd.n7683 0.637193
R12801 gnd.n2407 gnd.n2406 0.573776
R12802 gnd.n2406 gnd.n2404 0.573776
R12803 gnd.n2404 gnd.n2402 0.573776
R12804 gnd.n2402 gnd.n2400 0.573776
R12805 gnd.n2400 gnd.n2398 0.573776
R12806 gnd.n2398 gnd.n2396 0.573776
R12807 gnd.n2396 gnd.n2394 0.573776
R12808 gnd.n2394 gnd.n2392 0.573776
R12809 gnd.n2392 gnd.n2390 0.573776
R12810 gnd.n2426 gnd.n2425 0.573776
R12811 gnd.n2425 gnd.n2423 0.573776
R12812 gnd.n2423 gnd.n2421 0.573776
R12813 gnd.n2421 gnd.n2419 0.573776
R12814 gnd.n2419 gnd.n2417 0.573776
R12815 gnd.n2417 gnd.n2415 0.573776
R12816 gnd.n2415 gnd.n2413 0.573776
R12817 gnd.n2413 gnd.n2411 0.573776
R12818 gnd.n2411 gnd.n2409 0.573776
R12819 gnd.n23 gnd.n21 0.573776
R12820 gnd.n25 gnd.n23 0.573776
R12821 gnd.n27 gnd.n25 0.573776
R12822 gnd.n29 gnd.n27 0.573776
R12823 gnd.n31 gnd.n29 0.573776
R12824 gnd.n33 gnd.n31 0.573776
R12825 gnd.n35 gnd.n33 0.573776
R12826 gnd.n37 gnd.n35 0.573776
R12827 gnd.n38 gnd.n37 0.573776
R12828 gnd.n42 gnd.n40 0.573776
R12829 gnd.n44 gnd.n42 0.573776
R12830 gnd.n46 gnd.n44 0.573776
R12831 gnd.n48 gnd.n46 0.573776
R12832 gnd.n50 gnd.n48 0.573776
R12833 gnd.n52 gnd.n50 0.573776
R12834 gnd.n54 gnd.n52 0.573776
R12835 gnd.n56 gnd.n54 0.573776
R12836 gnd.n57 gnd.n56 0.573776
R12837 gnd.n2980 gnd.t160 0.547401
R12838 gnd.n3145 gnd.t168 0.547401
R12839 gnd.n4183 gnd.t102 0.547401
R12840 gnd.n3207 gnd.n2228 0.486781
R12841 gnd.n5998 gnd.n460 0.486781
R12842 gnd.n2783 gnd.n2782 0.48678
R12843 gnd.n4659 gnd.n1895 0.485256
R12844 gnd.n3524 gnd.n2182 0.480683
R12845 gnd.n2867 gnd.n2866 0.480683
R12846 gnd.n4063 gnd.n4058 0.477634
R12847 gnd.n4100 gnd.n4099 0.477634
R12848 gnd.n7532 gnd.n7531 0.477634
R12849 gnd.n7634 gnd.n7633 0.477634
R12850 gnd.n7626 gnd.n7625 0.465439
R12851 gnd.n7555 gnd.n7554 0.465439
R12852 gnd.n7107 gnd.n7104 0.465439
R12853 gnd.n7236 gnd.n453 0.465439
R12854 gnd.n4106 gnd.n2155 0.465439
R12855 gnd.n3870 gnd.n3869 0.465439
R12856 gnd.n6252 gnd.n6251 0.465439
R12857 gnd.n6183 gnd.n6182 0.465439
R12858 gnd.n4285 gnd.n976 0.459342
R12859 gnd.n6705 gnd.n6704 0.459342
R12860 gnd.n6917 gnd.n6916 0.459342
R12861 gnd.n4538 gnd.n4537 0.459342
R12862 gnd.n5948 gnd.n1312 0.451719
R12863 gnd.n6156 gnd.n6155 0.451719
R12864 gnd.n6163 gnd.n1181 0.388379
R12865 gnd.n7595 gnd.n7594 0.388379
R12866 gnd.n3484 gnd.n3483 0.388379
R12867 gnd.n3452 gnd.n3451 0.388379
R12868 gnd.n3420 gnd.n3419 0.388379
R12869 gnd.n3389 gnd.n3388 0.388379
R12870 gnd.n3357 gnd.n3356 0.388379
R12871 gnd.n3325 gnd.n3324 0.388379
R12872 gnd.n3293 gnd.n3292 0.388379
R12873 gnd.n3262 gnd.n3261 0.388379
R12874 gnd.n3816 gnd.n3758 0.388379
R12875 gnd.n5959 gnd.n5958 0.388379
R12876 gnd.n4658 gnd.n1086 0.378829
R12877 gnd.n7230 gnd.n7229 0.377553
R12878 gnd.n7684 gnd.n19 0.374463
R12879 gnd gnd.n7684 0.367492
R12880 gnd.n7345 gnd.t68 0.319156
R12881 gnd.n7377 gnd.t15 0.319156
R12882 gnd.n2701 gnd.n2679 0.311721
R12883 gnd.n3595 gnd.n3594 0.268793
R12884 gnd.n6174 gnd.n6173 0.247451
R12885 gnd.n5969 gnd.n5968 0.247451
R12886 gnd.n3594 gnd.n3593 0.241354
R12887 gnd.n563 gnd.n560 0.229039
R12888 gnd.n566 gnd.n563 0.229039
R12889 gnd.n1125 gnd.n1124 0.229039
R12890 gnd.n1126 gnd.n1125 0.229039
R12891 gnd.n2448 gnd.n0 0.210825
R12892 gnd.n2855 gnd.n2654 0.206293
R12893 gnd.n2283 gnd.t159 0.1828
R12894 gnd.n4215 gnd.t105 0.1828
R12895 gnd.n4247 gnd.t53 0.1828
R12896 gnd.n3501 gnd.n3473 0.155672
R12897 gnd.n3494 gnd.n3473 0.155672
R12898 gnd.n3494 gnd.n3493 0.155672
R12899 gnd.n3493 gnd.n3477 0.155672
R12900 gnd.n3486 gnd.n3477 0.155672
R12901 gnd.n3486 gnd.n3485 0.155672
R12902 gnd.n3469 gnd.n3441 0.155672
R12903 gnd.n3462 gnd.n3441 0.155672
R12904 gnd.n3462 gnd.n3461 0.155672
R12905 gnd.n3461 gnd.n3445 0.155672
R12906 gnd.n3454 gnd.n3445 0.155672
R12907 gnd.n3454 gnd.n3453 0.155672
R12908 gnd.n3437 gnd.n3409 0.155672
R12909 gnd.n3430 gnd.n3409 0.155672
R12910 gnd.n3430 gnd.n3429 0.155672
R12911 gnd.n3429 gnd.n3413 0.155672
R12912 gnd.n3422 gnd.n3413 0.155672
R12913 gnd.n3422 gnd.n3421 0.155672
R12914 gnd.n3406 gnd.n3378 0.155672
R12915 gnd.n3399 gnd.n3378 0.155672
R12916 gnd.n3399 gnd.n3398 0.155672
R12917 gnd.n3398 gnd.n3382 0.155672
R12918 gnd.n3391 gnd.n3382 0.155672
R12919 gnd.n3391 gnd.n3390 0.155672
R12920 gnd.n3374 gnd.n3346 0.155672
R12921 gnd.n3367 gnd.n3346 0.155672
R12922 gnd.n3367 gnd.n3366 0.155672
R12923 gnd.n3366 gnd.n3350 0.155672
R12924 gnd.n3359 gnd.n3350 0.155672
R12925 gnd.n3359 gnd.n3358 0.155672
R12926 gnd.n3342 gnd.n3314 0.155672
R12927 gnd.n3335 gnd.n3314 0.155672
R12928 gnd.n3335 gnd.n3334 0.155672
R12929 gnd.n3334 gnd.n3318 0.155672
R12930 gnd.n3327 gnd.n3318 0.155672
R12931 gnd.n3327 gnd.n3326 0.155672
R12932 gnd.n3310 gnd.n3282 0.155672
R12933 gnd.n3303 gnd.n3282 0.155672
R12934 gnd.n3303 gnd.n3302 0.155672
R12935 gnd.n3302 gnd.n3286 0.155672
R12936 gnd.n3295 gnd.n3286 0.155672
R12937 gnd.n3295 gnd.n3294 0.155672
R12938 gnd.n3279 gnd.n3251 0.155672
R12939 gnd.n3272 gnd.n3251 0.155672
R12940 gnd.n3272 gnd.n3271 0.155672
R12941 gnd.n3271 gnd.n3255 0.155672
R12942 gnd.n3264 gnd.n3255 0.155672
R12943 gnd.n3264 gnd.n3263 0.155672
R12944 gnd.n7382 gnd.n7381 0.152939
R12945 gnd.n7382 gnd.n287 0.152939
R12946 gnd.n7396 gnd.n287 0.152939
R12947 gnd.n7397 gnd.n7396 0.152939
R12948 gnd.n7398 gnd.n7397 0.152939
R12949 gnd.n7398 gnd.n273 0.152939
R12950 gnd.n7412 gnd.n273 0.152939
R12951 gnd.n7413 gnd.n7412 0.152939
R12952 gnd.n7414 gnd.n7413 0.152939
R12953 gnd.n7414 gnd.n257 0.152939
R12954 gnd.n7428 gnd.n257 0.152939
R12955 gnd.n7429 gnd.n7428 0.152939
R12956 gnd.n7430 gnd.n7429 0.152939
R12957 gnd.n7430 gnd.n242 0.152939
R12958 gnd.n7444 gnd.n242 0.152939
R12959 gnd.n7445 gnd.n7444 0.152939
R12960 gnd.n7446 gnd.n7445 0.152939
R12961 gnd.n7446 gnd.n226 0.152939
R12962 gnd.n7460 gnd.n226 0.152939
R12963 gnd.n7461 gnd.n7460 0.152939
R12964 gnd.n7462 gnd.n7461 0.152939
R12965 gnd.n7462 gnd.n210 0.152939
R12966 gnd.n7544 gnd.n210 0.152939
R12967 gnd.n7545 gnd.n7544 0.152939
R12968 gnd.n7546 gnd.n7545 0.152939
R12969 gnd.n7546 gnd.n133 0.152939
R12970 gnd.n7626 gnd.n133 0.152939
R12971 gnd.n7625 gnd.n134 0.152939
R12972 gnd.n136 gnd.n134 0.152939
R12973 gnd.n140 gnd.n136 0.152939
R12974 gnd.n141 gnd.n140 0.152939
R12975 gnd.n142 gnd.n141 0.152939
R12976 gnd.n143 gnd.n142 0.152939
R12977 gnd.n147 gnd.n143 0.152939
R12978 gnd.n148 gnd.n147 0.152939
R12979 gnd.n149 gnd.n148 0.152939
R12980 gnd.n150 gnd.n149 0.152939
R12981 gnd.n154 gnd.n150 0.152939
R12982 gnd.n155 gnd.n154 0.152939
R12983 gnd.n156 gnd.n155 0.152939
R12984 gnd.n157 gnd.n156 0.152939
R12985 gnd.n161 gnd.n157 0.152939
R12986 gnd.n162 gnd.n161 0.152939
R12987 gnd.n163 gnd.n162 0.152939
R12988 gnd.n164 gnd.n163 0.152939
R12989 gnd.n168 gnd.n164 0.152939
R12990 gnd.n169 gnd.n168 0.152939
R12991 gnd.n170 gnd.n169 0.152939
R12992 gnd.n171 gnd.n170 0.152939
R12993 gnd.n175 gnd.n171 0.152939
R12994 gnd.n176 gnd.n175 0.152939
R12995 gnd.n177 gnd.n176 0.152939
R12996 gnd.n178 gnd.n177 0.152939
R12997 gnd.n182 gnd.n178 0.152939
R12998 gnd.n183 gnd.n182 0.152939
R12999 gnd.n184 gnd.n183 0.152939
R13000 gnd.n185 gnd.n184 0.152939
R13001 gnd.n189 gnd.n185 0.152939
R13002 gnd.n190 gnd.n189 0.152939
R13003 gnd.n191 gnd.n190 0.152939
R13004 gnd.n192 gnd.n191 0.152939
R13005 gnd.n196 gnd.n192 0.152939
R13006 gnd.n197 gnd.n196 0.152939
R13007 gnd.n7556 gnd.n197 0.152939
R13008 gnd.n7556 gnd.n7555 0.152939
R13009 gnd.n7104 gnd.n589 0.152939
R13010 gnd.n591 gnd.n589 0.152939
R13011 gnd.n592 gnd.n591 0.152939
R13012 gnd.n5864 gnd.n592 0.152939
R13013 gnd.n5865 gnd.n5864 0.152939
R13014 gnd.n5865 gnd.n5863 0.152939
R13015 gnd.n5873 gnd.n5863 0.152939
R13016 gnd.n5874 gnd.n5873 0.152939
R13017 gnd.n5875 gnd.n5874 0.152939
R13018 gnd.n5876 gnd.n5875 0.152939
R13019 gnd.n5877 gnd.n5876 0.152939
R13020 gnd.n5878 gnd.n5877 0.152939
R13021 gnd.n5879 gnd.n5878 0.152939
R13022 gnd.n5880 gnd.n5879 0.152939
R13023 gnd.n5881 gnd.n5880 0.152939
R13024 gnd.n5881 gnd.n612 0.152939
R13025 gnd.n6931 gnd.n612 0.152939
R13026 gnd.n6932 gnd.n6931 0.152939
R13027 gnd.n6933 gnd.n6932 0.152939
R13028 gnd.n6934 gnd.n6933 0.152939
R13029 gnd.n6935 gnd.n6934 0.152939
R13030 gnd.n6936 gnd.n6935 0.152939
R13031 gnd.n6937 gnd.n6936 0.152939
R13032 gnd.n6938 gnd.n6937 0.152939
R13033 gnd.n6939 gnd.n6938 0.152939
R13034 gnd.n6940 gnd.n6939 0.152939
R13035 gnd.n6941 gnd.n6940 0.152939
R13036 gnd.n6942 gnd.n6941 0.152939
R13037 gnd.n6943 gnd.n6942 0.152939
R13038 gnd.n6944 gnd.n6943 0.152939
R13039 gnd.n6945 gnd.n6944 0.152939
R13040 gnd.n6945 gnd.n326 0.152939
R13041 gnd.n6946 gnd.n326 0.152939
R13042 gnd.n6947 gnd.n6946 0.152939
R13043 gnd.n6948 gnd.n6947 0.152939
R13044 gnd.n6949 gnd.n6948 0.152939
R13045 gnd.n6950 gnd.n6949 0.152939
R13046 gnd.n6951 gnd.n6950 0.152939
R13047 gnd.n6952 gnd.n6951 0.152939
R13048 gnd.n6953 gnd.n6952 0.152939
R13049 gnd.n6954 gnd.n6953 0.152939
R13050 gnd.n6955 gnd.n6954 0.152939
R13051 gnd.n6956 gnd.n6955 0.152939
R13052 gnd.n6957 gnd.n6956 0.152939
R13053 gnd.n6958 gnd.n6957 0.152939
R13054 gnd.n6959 gnd.n6958 0.152939
R13055 gnd.n6960 gnd.n6959 0.152939
R13056 gnd.n6961 gnd.n6960 0.152939
R13057 gnd.n6962 gnd.n6961 0.152939
R13058 gnd.n6963 gnd.n6962 0.152939
R13059 gnd.n6964 gnd.n6963 0.152939
R13060 gnd.n6965 gnd.n6964 0.152939
R13061 gnd.n6966 gnd.n6965 0.152939
R13062 gnd.n6967 gnd.n6966 0.152939
R13063 gnd.n6968 gnd.n6967 0.152939
R13064 gnd.n6969 gnd.n6968 0.152939
R13065 gnd.n6970 gnd.n6969 0.152939
R13066 gnd.n6971 gnd.n6970 0.152939
R13067 gnd.n6972 gnd.n6971 0.152939
R13068 gnd.n6973 gnd.n6972 0.152939
R13069 gnd.n6975 gnd.n6973 0.152939
R13070 gnd.n6975 gnd.n6974 0.152939
R13071 gnd.n6974 gnd.n203 0.152939
R13072 gnd.n7554 gnd.n203 0.152939
R13073 gnd.n546 gnd.n453 0.152939
R13074 gnd.n547 gnd.n546 0.152939
R13075 gnd.n548 gnd.n547 0.152939
R13076 gnd.n549 gnd.n548 0.152939
R13077 gnd.n550 gnd.n549 0.152939
R13078 gnd.n551 gnd.n550 0.152939
R13079 gnd.n552 gnd.n551 0.152939
R13080 gnd.n553 gnd.n552 0.152939
R13081 gnd.n554 gnd.n553 0.152939
R13082 gnd.n555 gnd.n554 0.152939
R13083 gnd.n556 gnd.n555 0.152939
R13084 gnd.n557 gnd.n556 0.152939
R13085 gnd.n558 gnd.n557 0.152939
R13086 gnd.n559 gnd.n558 0.152939
R13087 gnd.n560 gnd.n559 0.152939
R13088 gnd.n567 gnd.n566 0.152939
R13089 gnd.n568 gnd.n567 0.152939
R13090 gnd.n569 gnd.n568 0.152939
R13091 gnd.n570 gnd.n569 0.152939
R13092 gnd.n571 gnd.n570 0.152939
R13093 gnd.n572 gnd.n571 0.152939
R13094 gnd.n573 gnd.n572 0.152939
R13095 gnd.n574 gnd.n573 0.152939
R13096 gnd.n575 gnd.n574 0.152939
R13097 gnd.n576 gnd.n575 0.152939
R13098 gnd.n577 gnd.n576 0.152939
R13099 gnd.n578 gnd.n577 0.152939
R13100 gnd.n579 gnd.n578 0.152939
R13101 gnd.n580 gnd.n579 0.152939
R13102 gnd.n581 gnd.n580 0.152939
R13103 gnd.n582 gnd.n581 0.152939
R13104 gnd.n583 gnd.n582 0.152939
R13105 gnd.n7109 gnd.n583 0.152939
R13106 gnd.n7109 gnd.n7108 0.152939
R13107 gnd.n7108 gnd.n7107 0.152939
R13108 gnd.n7237 gnd.n7236 0.152939
R13109 gnd.n7238 gnd.n7237 0.152939
R13110 gnd.n7238 gnd.n436 0.152939
R13111 gnd.n7252 gnd.n436 0.152939
R13112 gnd.n7253 gnd.n7252 0.152939
R13113 gnd.n7254 gnd.n7253 0.152939
R13114 gnd.n7254 gnd.n418 0.152939
R13115 gnd.n7268 gnd.n418 0.152939
R13116 gnd.n7269 gnd.n7268 0.152939
R13117 gnd.n7270 gnd.n7269 0.152939
R13118 gnd.n7270 gnd.n402 0.152939
R13119 gnd.n7284 gnd.n402 0.152939
R13120 gnd.n7285 gnd.n7284 0.152939
R13121 gnd.n7286 gnd.n7285 0.152939
R13122 gnd.n7286 gnd.n384 0.152939
R13123 gnd.n7300 gnd.n384 0.152939
R13124 gnd.n7301 gnd.n7300 0.152939
R13125 gnd.n7302 gnd.n7301 0.152939
R13126 gnd.n7302 gnd.n368 0.152939
R13127 gnd.n7316 gnd.n368 0.152939
R13128 gnd.n7317 gnd.n7316 0.152939
R13129 gnd.n7318 gnd.n7317 0.152939
R13130 gnd.n7318 gnd.n350 0.152939
R13131 gnd.n7332 gnd.n350 0.152939
R13132 gnd.n7333 gnd.n7332 0.152939
R13133 gnd.n7334 gnd.n7333 0.152939
R13134 gnd.n7334 gnd.n335 0.152939
R13135 gnd.n6322 gnd.n976 0.152939
R13136 gnd.n6323 gnd.n6322 0.152939
R13137 gnd.n6324 gnd.n6323 0.152939
R13138 gnd.n6324 gnd.n970 0.152939
R13139 gnd.n6332 gnd.n970 0.152939
R13140 gnd.n6333 gnd.n6332 0.152939
R13141 gnd.n6334 gnd.n6333 0.152939
R13142 gnd.n6334 gnd.n964 0.152939
R13143 gnd.n6342 gnd.n964 0.152939
R13144 gnd.n6343 gnd.n6342 0.152939
R13145 gnd.n6344 gnd.n6343 0.152939
R13146 gnd.n6344 gnd.n958 0.152939
R13147 gnd.n6352 gnd.n958 0.152939
R13148 gnd.n6353 gnd.n6352 0.152939
R13149 gnd.n6354 gnd.n6353 0.152939
R13150 gnd.n6354 gnd.n952 0.152939
R13151 gnd.n6362 gnd.n952 0.152939
R13152 gnd.n6363 gnd.n6362 0.152939
R13153 gnd.n6364 gnd.n6363 0.152939
R13154 gnd.n6364 gnd.n946 0.152939
R13155 gnd.n6372 gnd.n946 0.152939
R13156 gnd.n6373 gnd.n6372 0.152939
R13157 gnd.n6374 gnd.n6373 0.152939
R13158 gnd.n6374 gnd.n940 0.152939
R13159 gnd.n6382 gnd.n940 0.152939
R13160 gnd.n6383 gnd.n6382 0.152939
R13161 gnd.n6384 gnd.n6383 0.152939
R13162 gnd.n6384 gnd.n934 0.152939
R13163 gnd.n6392 gnd.n934 0.152939
R13164 gnd.n6393 gnd.n6392 0.152939
R13165 gnd.n6394 gnd.n6393 0.152939
R13166 gnd.n6394 gnd.n928 0.152939
R13167 gnd.n6402 gnd.n928 0.152939
R13168 gnd.n6403 gnd.n6402 0.152939
R13169 gnd.n6404 gnd.n6403 0.152939
R13170 gnd.n6404 gnd.n922 0.152939
R13171 gnd.n6412 gnd.n922 0.152939
R13172 gnd.n6413 gnd.n6412 0.152939
R13173 gnd.n6414 gnd.n6413 0.152939
R13174 gnd.n6414 gnd.n916 0.152939
R13175 gnd.n6422 gnd.n916 0.152939
R13176 gnd.n6423 gnd.n6422 0.152939
R13177 gnd.n6424 gnd.n6423 0.152939
R13178 gnd.n6424 gnd.n910 0.152939
R13179 gnd.n6432 gnd.n910 0.152939
R13180 gnd.n6433 gnd.n6432 0.152939
R13181 gnd.n6434 gnd.n6433 0.152939
R13182 gnd.n6434 gnd.n904 0.152939
R13183 gnd.n6442 gnd.n904 0.152939
R13184 gnd.n6443 gnd.n6442 0.152939
R13185 gnd.n6444 gnd.n6443 0.152939
R13186 gnd.n6444 gnd.n898 0.152939
R13187 gnd.n6452 gnd.n898 0.152939
R13188 gnd.n6453 gnd.n6452 0.152939
R13189 gnd.n6454 gnd.n6453 0.152939
R13190 gnd.n6454 gnd.n892 0.152939
R13191 gnd.n6462 gnd.n892 0.152939
R13192 gnd.n6463 gnd.n6462 0.152939
R13193 gnd.n6464 gnd.n6463 0.152939
R13194 gnd.n6464 gnd.n886 0.152939
R13195 gnd.n6472 gnd.n886 0.152939
R13196 gnd.n6473 gnd.n6472 0.152939
R13197 gnd.n6474 gnd.n6473 0.152939
R13198 gnd.n6474 gnd.n880 0.152939
R13199 gnd.n6482 gnd.n880 0.152939
R13200 gnd.n6483 gnd.n6482 0.152939
R13201 gnd.n6484 gnd.n6483 0.152939
R13202 gnd.n6484 gnd.n874 0.152939
R13203 gnd.n6492 gnd.n874 0.152939
R13204 gnd.n6493 gnd.n6492 0.152939
R13205 gnd.n6494 gnd.n6493 0.152939
R13206 gnd.n6494 gnd.n868 0.152939
R13207 gnd.n6502 gnd.n868 0.152939
R13208 gnd.n6503 gnd.n6502 0.152939
R13209 gnd.n6504 gnd.n6503 0.152939
R13210 gnd.n6504 gnd.n862 0.152939
R13211 gnd.n6512 gnd.n862 0.152939
R13212 gnd.n6513 gnd.n6512 0.152939
R13213 gnd.n6514 gnd.n6513 0.152939
R13214 gnd.n6514 gnd.n856 0.152939
R13215 gnd.n6522 gnd.n856 0.152939
R13216 gnd.n6523 gnd.n6522 0.152939
R13217 gnd.n6524 gnd.n6523 0.152939
R13218 gnd.n6524 gnd.n850 0.152939
R13219 gnd.n6532 gnd.n850 0.152939
R13220 gnd.n6533 gnd.n6532 0.152939
R13221 gnd.n6534 gnd.n6533 0.152939
R13222 gnd.n6534 gnd.n844 0.152939
R13223 gnd.n6542 gnd.n844 0.152939
R13224 gnd.n6543 gnd.n6542 0.152939
R13225 gnd.n6544 gnd.n6543 0.152939
R13226 gnd.n6544 gnd.n838 0.152939
R13227 gnd.n6552 gnd.n838 0.152939
R13228 gnd.n6553 gnd.n6552 0.152939
R13229 gnd.n6554 gnd.n6553 0.152939
R13230 gnd.n6554 gnd.n832 0.152939
R13231 gnd.n6562 gnd.n832 0.152939
R13232 gnd.n6563 gnd.n6562 0.152939
R13233 gnd.n6564 gnd.n6563 0.152939
R13234 gnd.n6564 gnd.n826 0.152939
R13235 gnd.n6572 gnd.n826 0.152939
R13236 gnd.n6573 gnd.n6572 0.152939
R13237 gnd.n6574 gnd.n6573 0.152939
R13238 gnd.n6574 gnd.n820 0.152939
R13239 gnd.n6582 gnd.n820 0.152939
R13240 gnd.n6583 gnd.n6582 0.152939
R13241 gnd.n6584 gnd.n6583 0.152939
R13242 gnd.n6584 gnd.n814 0.152939
R13243 gnd.n6592 gnd.n814 0.152939
R13244 gnd.n6593 gnd.n6592 0.152939
R13245 gnd.n6594 gnd.n6593 0.152939
R13246 gnd.n6594 gnd.n808 0.152939
R13247 gnd.n6602 gnd.n808 0.152939
R13248 gnd.n6603 gnd.n6602 0.152939
R13249 gnd.n6604 gnd.n6603 0.152939
R13250 gnd.n6604 gnd.n802 0.152939
R13251 gnd.n6612 gnd.n802 0.152939
R13252 gnd.n6613 gnd.n6612 0.152939
R13253 gnd.n6614 gnd.n6613 0.152939
R13254 gnd.n6614 gnd.n796 0.152939
R13255 gnd.n6622 gnd.n796 0.152939
R13256 gnd.n6623 gnd.n6622 0.152939
R13257 gnd.n6624 gnd.n6623 0.152939
R13258 gnd.n6624 gnd.n790 0.152939
R13259 gnd.n6632 gnd.n790 0.152939
R13260 gnd.n6633 gnd.n6632 0.152939
R13261 gnd.n6634 gnd.n6633 0.152939
R13262 gnd.n6634 gnd.n784 0.152939
R13263 gnd.n6642 gnd.n784 0.152939
R13264 gnd.n6643 gnd.n6642 0.152939
R13265 gnd.n6644 gnd.n6643 0.152939
R13266 gnd.n6644 gnd.n778 0.152939
R13267 gnd.n6652 gnd.n778 0.152939
R13268 gnd.n6653 gnd.n6652 0.152939
R13269 gnd.n6654 gnd.n6653 0.152939
R13270 gnd.n6654 gnd.n772 0.152939
R13271 gnd.n6662 gnd.n772 0.152939
R13272 gnd.n6663 gnd.n6662 0.152939
R13273 gnd.n6664 gnd.n6663 0.152939
R13274 gnd.n6664 gnd.n766 0.152939
R13275 gnd.n6672 gnd.n766 0.152939
R13276 gnd.n6673 gnd.n6672 0.152939
R13277 gnd.n6674 gnd.n6673 0.152939
R13278 gnd.n6674 gnd.n760 0.152939
R13279 gnd.n6682 gnd.n760 0.152939
R13280 gnd.n6683 gnd.n6682 0.152939
R13281 gnd.n6684 gnd.n6683 0.152939
R13282 gnd.n6684 gnd.n754 0.152939
R13283 gnd.n6692 gnd.n754 0.152939
R13284 gnd.n6693 gnd.n6692 0.152939
R13285 gnd.n6695 gnd.n6693 0.152939
R13286 gnd.n6695 gnd.n6694 0.152939
R13287 gnd.n6694 gnd.n748 0.152939
R13288 gnd.n6704 gnd.n748 0.152939
R13289 gnd.n6705 gnd.n743 0.152939
R13290 gnd.n6713 gnd.n743 0.152939
R13291 gnd.n6714 gnd.n6713 0.152939
R13292 gnd.n6715 gnd.n6714 0.152939
R13293 gnd.n6715 gnd.n737 0.152939
R13294 gnd.n6723 gnd.n737 0.152939
R13295 gnd.n6724 gnd.n6723 0.152939
R13296 gnd.n6725 gnd.n6724 0.152939
R13297 gnd.n6725 gnd.n731 0.152939
R13298 gnd.n6733 gnd.n731 0.152939
R13299 gnd.n6734 gnd.n6733 0.152939
R13300 gnd.n6735 gnd.n6734 0.152939
R13301 gnd.n6735 gnd.n725 0.152939
R13302 gnd.n6743 gnd.n725 0.152939
R13303 gnd.n6744 gnd.n6743 0.152939
R13304 gnd.n6745 gnd.n6744 0.152939
R13305 gnd.n6745 gnd.n719 0.152939
R13306 gnd.n6753 gnd.n719 0.152939
R13307 gnd.n6754 gnd.n6753 0.152939
R13308 gnd.n6755 gnd.n6754 0.152939
R13309 gnd.n6755 gnd.n713 0.152939
R13310 gnd.n6763 gnd.n713 0.152939
R13311 gnd.n6764 gnd.n6763 0.152939
R13312 gnd.n6765 gnd.n6764 0.152939
R13313 gnd.n6765 gnd.n707 0.152939
R13314 gnd.n6773 gnd.n707 0.152939
R13315 gnd.n6774 gnd.n6773 0.152939
R13316 gnd.n6775 gnd.n6774 0.152939
R13317 gnd.n6775 gnd.n701 0.152939
R13318 gnd.n6783 gnd.n701 0.152939
R13319 gnd.n6784 gnd.n6783 0.152939
R13320 gnd.n6785 gnd.n6784 0.152939
R13321 gnd.n6785 gnd.n695 0.152939
R13322 gnd.n6793 gnd.n695 0.152939
R13323 gnd.n6794 gnd.n6793 0.152939
R13324 gnd.n6795 gnd.n6794 0.152939
R13325 gnd.n6795 gnd.n689 0.152939
R13326 gnd.n6803 gnd.n689 0.152939
R13327 gnd.n6804 gnd.n6803 0.152939
R13328 gnd.n6805 gnd.n6804 0.152939
R13329 gnd.n6805 gnd.n683 0.152939
R13330 gnd.n6813 gnd.n683 0.152939
R13331 gnd.n6814 gnd.n6813 0.152939
R13332 gnd.n6815 gnd.n6814 0.152939
R13333 gnd.n6815 gnd.n677 0.152939
R13334 gnd.n6823 gnd.n677 0.152939
R13335 gnd.n6824 gnd.n6823 0.152939
R13336 gnd.n6825 gnd.n6824 0.152939
R13337 gnd.n6825 gnd.n671 0.152939
R13338 gnd.n6833 gnd.n671 0.152939
R13339 gnd.n6834 gnd.n6833 0.152939
R13340 gnd.n6835 gnd.n6834 0.152939
R13341 gnd.n6835 gnd.n665 0.152939
R13342 gnd.n6843 gnd.n665 0.152939
R13343 gnd.n6844 gnd.n6843 0.152939
R13344 gnd.n6845 gnd.n6844 0.152939
R13345 gnd.n6845 gnd.n659 0.152939
R13346 gnd.n6853 gnd.n659 0.152939
R13347 gnd.n6854 gnd.n6853 0.152939
R13348 gnd.n6855 gnd.n6854 0.152939
R13349 gnd.n6855 gnd.n653 0.152939
R13350 gnd.n6863 gnd.n653 0.152939
R13351 gnd.n6864 gnd.n6863 0.152939
R13352 gnd.n6865 gnd.n6864 0.152939
R13353 gnd.n6865 gnd.n647 0.152939
R13354 gnd.n6873 gnd.n647 0.152939
R13355 gnd.n6874 gnd.n6873 0.152939
R13356 gnd.n6875 gnd.n6874 0.152939
R13357 gnd.n6875 gnd.n641 0.152939
R13358 gnd.n6883 gnd.n641 0.152939
R13359 gnd.n6884 gnd.n6883 0.152939
R13360 gnd.n6885 gnd.n6884 0.152939
R13361 gnd.n6885 gnd.n635 0.152939
R13362 gnd.n6893 gnd.n635 0.152939
R13363 gnd.n6894 gnd.n6893 0.152939
R13364 gnd.n6895 gnd.n6894 0.152939
R13365 gnd.n6895 gnd.n629 0.152939
R13366 gnd.n6903 gnd.n629 0.152939
R13367 gnd.n6904 gnd.n6903 0.152939
R13368 gnd.n6905 gnd.n6904 0.152939
R13369 gnd.n6905 gnd.n623 0.152939
R13370 gnd.n6914 gnd.n623 0.152939
R13371 gnd.n6915 gnd.n6914 0.152939
R13372 gnd.n6917 gnd.n6915 0.152939
R13373 gnd.n4538 gnd.n1944 0.152939
R13374 gnd.n4544 gnd.n1944 0.152939
R13375 gnd.n4545 gnd.n4544 0.152939
R13376 gnd.n4546 gnd.n4545 0.152939
R13377 gnd.n4546 gnd.n1940 0.152939
R13378 gnd.n4552 gnd.n1940 0.152939
R13379 gnd.n4553 gnd.n4552 0.152939
R13380 gnd.n4554 gnd.n4553 0.152939
R13381 gnd.n4555 gnd.n4554 0.152939
R13382 gnd.n4557 gnd.n4555 0.152939
R13383 gnd.n4557 gnd.n4556 0.152939
R13384 gnd.n4556 gnd.n1915 0.152939
R13385 gnd.n4612 gnd.n1915 0.152939
R13386 gnd.n4613 gnd.n4612 0.152939
R13387 gnd.n4614 gnd.n4613 0.152939
R13388 gnd.n4614 gnd.n1911 0.152939
R13389 gnd.n4620 gnd.n1911 0.152939
R13390 gnd.n4621 gnd.n4620 0.152939
R13391 gnd.n4622 gnd.n4621 0.152939
R13392 gnd.n4622 gnd.n1907 0.152939
R13393 gnd.n4628 gnd.n1907 0.152939
R13394 gnd.n4629 gnd.n4628 0.152939
R13395 gnd.n4630 gnd.n4629 0.152939
R13396 gnd.n4630 gnd.n1901 0.152939
R13397 gnd.n4776 gnd.n1901 0.152939
R13398 gnd.n4777 gnd.n4776 0.152939
R13399 gnd.n4778 gnd.n4777 0.152939
R13400 gnd.n4778 gnd.n1887 0.152939
R13401 gnd.n4795 gnd.n1887 0.152939
R13402 gnd.n4796 gnd.n4795 0.152939
R13403 gnd.n4797 gnd.n4796 0.152939
R13404 gnd.n4797 gnd.n1873 0.152939
R13405 gnd.n4814 gnd.n1873 0.152939
R13406 gnd.n4815 gnd.n4814 0.152939
R13407 gnd.n4816 gnd.n4815 0.152939
R13408 gnd.n4816 gnd.n1859 0.152939
R13409 gnd.n4833 gnd.n1859 0.152939
R13410 gnd.n4834 gnd.n4833 0.152939
R13411 gnd.n4835 gnd.n4834 0.152939
R13412 gnd.n4835 gnd.n1845 0.152939
R13413 gnd.n4852 gnd.n1845 0.152939
R13414 gnd.n4853 gnd.n4852 0.152939
R13415 gnd.n4854 gnd.n4853 0.152939
R13416 gnd.n4854 gnd.n1830 0.152939
R13417 gnd.n4871 gnd.n1830 0.152939
R13418 gnd.n4872 gnd.n4871 0.152939
R13419 gnd.n4873 gnd.n4872 0.152939
R13420 gnd.n4874 gnd.n4873 0.152939
R13421 gnd.n4874 gnd.n1817 0.152939
R13422 gnd.n5092 gnd.n1817 0.152939
R13423 gnd.n5093 gnd.n5092 0.152939
R13424 gnd.n5094 gnd.n5093 0.152939
R13425 gnd.n5094 gnd.n1743 0.152939
R13426 gnd.n5133 gnd.n1743 0.152939
R13427 gnd.n5134 gnd.n5133 0.152939
R13428 gnd.n5135 gnd.n5134 0.152939
R13429 gnd.n5136 gnd.n5135 0.152939
R13430 gnd.n5136 gnd.n1716 0.152939
R13431 gnd.n5169 gnd.n1716 0.152939
R13432 gnd.n5170 gnd.n5169 0.152939
R13433 gnd.n5171 gnd.n5170 0.152939
R13434 gnd.n5171 gnd.n1694 0.152939
R13435 gnd.n5197 gnd.n1694 0.152939
R13436 gnd.n5198 gnd.n5197 0.152939
R13437 gnd.n5199 gnd.n5198 0.152939
R13438 gnd.n5200 gnd.n5199 0.152939
R13439 gnd.n5200 gnd.n1662 0.152939
R13440 gnd.n5234 gnd.n1662 0.152939
R13441 gnd.n5235 gnd.n5234 0.152939
R13442 gnd.n5236 gnd.n5235 0.152939
R13443 gnd.n5237 gnd.n5236 0.152939
R13444 gnd.n5238 gnd.n5237 0.152939
R13445 gnd.n5240 gnd.n5238 0.152939
R13446 gnd.n5241 gnd.n5240 0.152939
R13447 gnd.n5241 gnd.n1621 0.152939
R13448 gnd.n5328 gnd.n1621 0.152939
R13449 gnd.n5329 gnd.n5328 0.152939
R13450 gnd.n5330 gnd.n5329 0.152939
R13451 gnd.n5330 gnd.n1603 0.152939
R13452 gnd.n5371 gnd.n1603 0.152939
R13453 gnd.n5372 gnd.n5371 0.152939
R13454 gnd.n5373 gnd.n5372 0.152939
R13455 gnd.n5373 gnd.n1579 0.152939
R13456 gnd.n5405 gnd.n1579 0.152939
R13457 gnd.n5406 gnd.n5405 0.152939
R13458 gnd.n5407 gnd.n5406 0.152939
R13459 gnd.n5407 gnd.n1556 0.152939
R13460 gnd.n5446 gnd.n1556 0.152939
R13461 gnd.n5447 gnd.n5446 0.152939
R13462 gnd.n5448 gnd.n5447 0.152939
R13463 gnd.n5448 gnd.n1535 0.152939
R13464 gnd.n5493 gnd.n1535 0.152939
R13465 gnd.n5494 gnd.n5493 0.152939
R13466 gnd.n5495 gnd.n5494 0.152939
R13467 gnd.n5495 gnd.n1508 0.152939
R13468 gnd.n5525 gnd.n1508 0.152939
R13469 gnd.n5526 gnd.n5525 0.152939
R13470 gnd.n5527 gnd.n5526 0.152939
R13471 gnd.n5527 gnd.n1486 0.152939
R13472 gnd.n5571 gnd.n1486 0.152939
R13473 gnd.n5572 gnd.n5571 0.152939
R13474 gnd.n5573 gnd.n5572 0.152939
R13475 gnd.n5573 gnd.n1399 0.152939
R13476 gnd.n5719 gnd.n1399 0.152939
R13477 gnd.n5720 gnd.n5719 0.152939
R13478 gnd.n5721 gnd.n5720 0.152939
R13479 gnd.n5721 gnd.n1384 0.152939
R13480 gnd.n5738 gnd.n1384 0.152939
R13481 gnd.n5739 gnd.n5738 0.152939
R13482 gnd.n5740 gnd.n5739 0.152939
R13483 gnd.n5740 gnd.n1370 0.152939
R13484 gnd.n5757 gnd.n1370 0.152939
R13485 gnd.n5758 gnd.n5757 0.152939
R13486 gnd.n5759 gnd.n5758 0.152939
R13487 gnd.n5759 gnd.n1356 0.152939
R13488 gnd.n5776 gnd.n1356 0.152939
R13489 gnd.n5777 gnd.n5776 0.152939
R13490 gnd.n5778 gnd.n5777 0.152939
R13491 gnd.n5778 gnd.n1342 0.152939
R13492 gnd.n5795 gnd.n1342 0.152939
R13493 gnd.n5796 gnd.n5795 0.152939
R13494 gnd.n5797 gnd.n5796 0.152939
R13495 gnd.n5797 gnd.n1328 0.152939
R13496 gnd.n5814 gnd.n1328 0.152939
R13497 gnd.n5815 gnd.n5814 0.152939
R13498 gnd.n5816 gnd.n5815 0.152939
R13499 gnd.n5817 gnd.n5816 0.152939
R13500 gnd.n5818 gnd.n5817 0.152939
R13501 gnd.n5842 gnd.n5818 0.152939
R13502 gnd.n5843 gnd.n5842 0.152939
R13503 gnd.n5844 gnd.n5843 0.152939
R13504 gnd.n5845 gnd.n5844 0.152939
R13505 gnd.n5846 gnd.n5845 0.152939
R13506 gnd.n5849 gnd.n5846 0.152939
R13507 gnd.n5850 gnd.n5849 0.152939
R13508 gnd.n5851 gnd.n5850 0.152939
R13509 gnd.n5852 gnd.n5851 0.152939
R13510 gnd.n5855 gnd.n5852 0.152939
R13511 gnd.n5856 gnd.n5855 0.152939
R13512 gnd.n5857 gnd.n5856 0.152939
R13513 gnd.n5858 gnd.n5857 0.152939
R13514 gnd.n5889 gnd.n5858 0.152939
R13515 gnd.n5890 gnd.n5889 0.152939
R13516 gnd.n5892 gnd.n5890 0.152939
R13517 gnd.n5893 gnd.n5892 0.152939
R13518 gnd.n5894 gnd.n5893 0.152939
R13519 gnd.n5895 gnd.n5894 0.152939
R13520 gnd.n5896 gnd.n5895 0.152939
R13521 gnd.n5898 gnd.n5896 0.152939
R13522 gnd.n5898 gnd.n5897 0.152939
R13523 gnd.n5897 gnd.n617 0.152939
R13524 gnd.n618 gnd.n617 0.152939
R13525 gnd.n619 gnd.n618 0.152939
R13526 gnd.n6916 gnd.n619 0.152939
R13527 gnd.n4286 gnd.n4285 0.152939
R13528 gnd.n4287 gnd.n4286 0.152939
R13529 gnd.n4288 gnd.n4287 0.152939
R13530 gnd.n4289 gnd.n4288 0.152939
R13531 gnd.n4290 gnd.n4289 0.152939
R13532 gnd.n4291 gnd.n4290 0.152939
R13533 gnd.n4292 gnd.n4291 0.152939
R13534 gnd.n4293 gnd.n4292 0.152939
R13535 gnd.n4294 gnd.n4293 0.152939
R13536 gnd.n4295 gnd.n4294 0.152939
R13537 gnd.n4296 gnd.n4295 0.152939
R13538 gnd.n4297 gnd.n4296 0.152939
R13539 gnd.n4298 gnd.n4297 0.152939
R13540 gnd.n4299 gnd.n4298 0.152939
R13541 gnd.n4300 gnd.n4299 0.152939
R13542 gnd.n4301 gnd.n4300 0.152939
R13543 gnd.n4302 gnd.n4301 0.152939
R13544 gnd.n4303 gnd.n4302 0.152939
R13545 gnd.n4304 gnd.n4303 0.152939
R13546 gnd.n4305 gnd.n4304 0.152939
R13547 gnd.n4306 gnd.n4305 0.152939
R13548 gnd.n4307 gnd.n4306 0.152939
R13549 gnd.n4308 gnd.n4307 0.152939
R13550 gnd.n4309 gnd.n4308 0.152939
R13551 gnd.n4310 gnd.n4309 0.152939
R13552 gnd.n4311 gnd.n4310 0.152939
R13553 gnd.n4312 gnd.n4311 0.152939
R13554 gnd.n4313 gnd.n4312 0.152939
R13555 gnd.n4314 gnd.n4313 0.152939
R13556 gnd.n4315 gnd.n4314 0.152939
R13557 gnd.n4316 gnd.n4315 0.152939
R13558 gnd.n4317 gnd.n4316 0.152939
R13559 gnd.n4318 gnd.n4317 0.152939
R13560 gnd.n4319 gnd.n4318 0.152939
R13561 gnd.n4320 gnd.n4319 0.152939
R13562 gnd.n4321 gnd.n4320 0.152939
R13563 gnd.n4322 gnd.n4321 0.152939
R13564 gnd.n4323 gnd.n4322 0.152939
R13565 gnd.n4324 gnd.n4323 0.152939
R13566 gnd.n4325 gnd.n4324 0.152939
R13567 gnd.n4326 gnd.n4325 0.152939
R13568 gnd.n4327 gnd.n4326 0.152939
R13569 gnd.n4328 gnd.n4327 0.152939
R13570 gnd.n4329 gnd.n4328 0.152939
R13571 gnd.n4330 gnd.n4329 0.152939
R13572 gnd.n4331 gnd.n4330 0.152939
R13573 gnd.n4332 gnd.n4331 0.152939
R13574 gnd.n4333 gnd.n4332 0.152939
R13575 gnd.n4334 gnd.n4333 0.152939
R13576 gnd.n4335 gnd.n4334 0.152939
R13577 gnd.n4336 gnd.n4335 0.152939
R13578 gnd.n4337 gnd.n4336 0.152939
R13579 gnd.n4338 gnd.n4337 0.152939
R13580 gnd.n4339 gnd.n4338 0.152939
R13581 gnd.n4340 gnd.n4339 0.152939
R13582 gnd.n4341 gnd.n4340 0.152939
R13583 gnd.n4342 gnd.n4341 0.152939
R13584 gnd.n4343 gnd.n4342 0.152939
R13585 gnd.n4344 gnd.n4343 0.152939
R13586 gnd.n4345 gnd.n4344 0.152939
R13587 gnd.n4346 gnd.n4345 0.152939
R13588 gnd.n4347 gnd.n4346 0.152939
R13589 gnd.n4348 gnd.n4347 0.152939
R13590 gnd.n4349 gnd.n4348 0.152939
R13591 gnd.n4350 gnd.n4349 0.152939
R13592 gnd.n4351 gnd.n4350 0.152939
R13593 gnd.n4352 gnd.n4351 0.152939
R13594 gnd.n4353 gnd.n4352 0.152939
R13595 gnd.n4354 gnd.n4353 0.152939
R13596 gnd.n4355 gnd.n4354 0.152939
R13597 gnd.n4356 gnd.n4355 0.152939
R13598 gnd.n4357 gnd.n4356 0.152939
R13599 gnd.n4358 gnd.n4357 0.152939
R13600 gnd.n4359 gnd.n4358 0.152939
R13601 gnd.n4360 gnd.n4359 0.152939
R13602 gnd.n4361 gnd.n4360 0.152939
R13603 gnd.n4362 gnd.n4361 0.152939
R13604 gnd.n4363 gnd.n4362 0.152939
R13605 gnd.n4364 gnd.n4363 0.152939
R13606 gnd.n4365 gnd.n4364 0.152939
R13607 gnd.n4366 gnd.n4365 0.152939
R13608 gnd.n4367 gnd.n4366 0.152939
R13609 gnd.n4367 gnd.n1945 0.152939
R13610 gnd.n4537 gnd.n1945 0.152939
R13611 gnd.n3626 gnd.n2182 0.152939
R13612 gnd.n3626 gnd.n3625 0.152939
R13613 gnd.n3625 gnd.n3624 0.152939
R13614 gnd.n3624 gnd.n2184 0.152939
R13615 gnd.n2185 gnd.n2184 0.152939
R13616 gnd.n2186 gnd.n2185 0.152939
R13617 gnd.n2187 gnd.n2186 0.152939
R13618 gnd.n2188 gnd.n2187 0.152939
R13619 gnd.n2189 gnd.n2188 0.152939
R13620 gnd.n2190 gnd.n2189 0.152939
R13621 gnd.n2191 gnd.n2190 0.152939
R13622 gnd.n2192 gnd.n2191 0.152939
R13623 gnd.n2193 gnd.n2192 0.152939
R13624 gnd.n2194 gnd.n2193 0.152939
R13625 gnd.n3596 gnd.n2194 0.152939
R13626 gnd.n3596 gnd.n3595 0.152939
R13627 gnd.n2868 gnd.n2867 0.152939
R13628 gnd.n2868 gnd.n2572 0.152939
R13629 gnd.n2896 gnd.n2572 0.152939
R13630 gnd.n2897 gnd.n2896 0.152939
R13631 gnd.n2898 gnd.n2897 0.152939
R13632 gnd.n2899 gnd.n2898 0.152939
R13633 gnd.n2899 gnd.n2544 0.152939
R13634 gnd.n2926 gnd.n2544 0.152939
R13635 gnd.n2927 gnd.n2926 0.152939
R13636 gnd.n2928 gnd.n2927 0.152939
R13637 gnd.n2928 gnd.n2522 0.152939
R13638 gnd.n2957 gnd.n2522 0.152939
R13639 gnd.n2958 gnd.n2957 0.152939
R13640 gnd.n2959 gnd.n2958 0.152939
R13641 gnd.n2960 gnd.n2959 0.152939
R13642 gnd.n2962 gnd.n2960 0.152939
R13643 gnd.n2962 gnd.n2961 0.152939
R13644 gnd.n2961 gnd.n2471 0.152939
R13645 gnd.n2472 gnd.n2471 0.152939
R13646 gnd.n2473 gnd.n2472 0.152939
R13647 gnd.n2492 gnd.n2473 0.152939
R13648 gnd.n2493 gnd.n2492 0.152939
R13649 gnd.n2493 gnd.n2379 0.152939
R13650 gnd.n3052 gnd.n2379 0.152939
R13651 gnd.n3053 gnd.n3052 0.152939
R13652 gnd.n3054 gnd.n3053 0.152939
R13653 gnd.n3055 gnd.n3054 0.152939
R13654 gnd.n3055 gnd.n2352 0.152939
R13655 gnd.n3092 gnd.n2352 0.152939
R13656 gnd.n3093 gnd.n3092 0.152939
R13657 gnd.n3094 gnd.n3093 0.152939
R13658 gnd.n3095 gnd.n3094 0.152939
R13659 gnd.n3095 gnd.n2325 0.152939
R13660 gnd.n3137 gnd.n2325 0.152939
R13661 gnd.n3138 gnd.n3137 0.152939
R13662 gnd.n3139 gnd.n3138 0.152939
R13663 gnd.n3140 gnd.n3139 0.152939
R13664 gnd.n3140 gnd.n2297 0.152939
R13665 gnd.n3177 gnd.n2297 0.152939
R13666 gnd.n3178 gnd.n3177 0.152939
R13667 gnd.n3179 gnd.n3178 0.152939
R13668 gnd.n3180 gnd.n3179 0.152939
R13669 gnd.n3180 gnd.n2270 0.152939
R13670 gnd.n3226 gnd.n2270 0.152939
R13671 gnd.n3227 gnd.n3226 0.152939
R13672 gnd.n3228 gnd.n3227 0.152939
R13673 gnd.n3229 gnd.n3228 0.152939
R13674 gnd.n3229 gnd.n2243 0.152939
R13675 gnd.n3520 gnd.n2243 0.152939
R13676 gnd.n3521 gnd.n3520 0.152939
R13677 gnd.n3522 gnd.n3521 0.152939
R13678 gnd.n3523 gnd.n3522 0.152939
R13679 gnd.n3524 gnd.n3523 0.152939
R13680 gnd.n2866 gnd.n2596 0.152939
R13681 gnd.n2617 gnd.n2596 0.152939
R13682 gnd.n2618 gnd.n2617 0.152939
R13683 gnd.n2624 gnd.n2618 0.152939
R13684 gnd.n2625 gnd.n2624 0.152939
R13685 gnd.n2626 gnd.n2625 0.152939
R13686 gnd.n2626 gnd.n2615 0.152939
R13687 gnd.n2634 gnd.n2615 0.152939
R13688 gnd.n2635 gnd.n2634 0.152939
R13689 gnd.n2636 gnd.n2635 0.152939
R13690 gnd.n2636 gnd.n2613 0.152939
R13691 gnd.n2644 gnd.n2613 0.152939
R13692 gnd.n2645 gnd.n2644 0.152939
R13693 gnd.n2646 gnd.n2645 0.152939
R13694 gnd.n2646 gnd.n2611 0.152939
R13695 gnd.n2654 gnd.n2611 0.152939
R13696 gnd.n3593 gnd.n2199 0.152939
R13697 gnd.n2201 gnd.n2199 0.152939
R13698 gnd.n2202 gnd.n2201 0.152939
R13699 gnd.n2203 gnd.n2202 0.152939
R13700 gnd.n2204 gnd.n2203 0.152939
R13701 gnd.n2205 gnd.n2204 0.152939
R13702 gnd.n2206 gnd.n2205 0.152939
R13703 gnd.n2207 gnd.n2206 0.152939
R13704 gnd.n2208 gnd.n2207 0.152939
R13705 gnd.n2209 gnd.n2208 0.152939
R13706 gnd.n2210 gnd.n2209 0.152939
R13707 gnd.n2211 gnd.n2210 0.152939
R13708 gnd.n2212 gnd.n2211 0.152939
R13709 gnd.n2213 gnd.n2212 0.152939
R13710 gnd.n2214 gnd.n2213 0.152939
R13711 gnd.n2215 gnd.n2214 0.152939
R13712 gnd.n2216 gnd.n2215 0.152939
R13713 gnd.n2217 gnd.n2216 0.152939
R13714 gnd.n2218 gnd.n2217 0.152939
R13715 gnd.n2219 gnd.n2218 0.152939
R13716 gnd.n2220 gnd.n2219 0.152939
R13717 gnd.n2221 gnd.n2220 0.152939
R13718 gnd.n2225 gnd.n2221 0.152939
R13719 gnd.n2226 gnd.n2225 0.152939
R13720 gnd.n2227 gnd.n2226 0.152939
R13721 gnd.n2228 gnd.n2227 0.152939
R13722 gnd.n3029 gnd.n3028 0.152939
R13723 gnd.n3030 gnd.n3029 0.152939
R13724 gnd.n3031 gnd.n3030 0.152939
R13725 gnd.n3032 gnd.n3031 0.152939
R13726 gnd.n3033 gnd.n3032 0.152939
R13727 gnd.n3034 gnd.n3033 0.152939
R13728 gnd.n3034 gnd.n2333 0.152939
R13729 gnd.n3113 gnd.n2333 0.152939
R13730 gnd.n3114 gnd.n3113 0.152939
R13731 gnd.n3115 gnd.n3114 0.152939
R13732 gnd.n3116 gnd.n3115 0.152939
R13733 gnd.n3117 gnd.n3116 0.152939
R13734 gnd.n3118 gnd.n3117 0.152939
R13735 gnd.n3119 gnd.n3118 0.152939
R13736 gnd.n3120 gnd.n3119 0.152939
R13737 gnd.n3121 gnd.n3120 0.152939
R13738 gnd.n3121 gnd.n2277 0.152939
R13739 gnd.n3198 gnd.n2277 0.152939
R13740 gnd.n3199 gnd.n3198 0.152939
R13741 gnd.n3200 gnd.n3199 0.152939
R13742 gnd.n3201 gnd.n3200 0.152939
R13743 gnd.n3202 gnd.n3201 0.152939
R13744 gnd.n3203 gnd.n3202 0.152939
R13745 gnd.n3204 gnd.n3203 0.152939
R13746 gnd.n3205 gnd.n3204 0.152939
R13747 gnd.n3206 gnd.n3205 0.152939
R13748 gnd.n3208 gnd.n3206 0.152939
R13749 gnd.n3208 gnd.n3207 0.152939
R13750 gnd.n2784 gnd.n2783 0.152939
R13751 gnd.n2784 gnd.n2674 0.152939
R13752 gnd.n2799 gnd.n2674 0.152939
R13753 gnd.n2800 gnd.n2799 0.152939
R13754 gnd.n2801 gnd.n2800 0.152939
R13755 gnd.n2801 gnd.n2662 0.152939
R13756 gnd.n2815 gnd.n2662 0.152939
R13757 gnd.n2816 gnd.n2815 0.152939
R13758 gnd.n2817 gnd.n2816 0.152939
R13759 gnd.n2818 gnd.n2817 0.152939
R13760 gnd.n2819 gnd.n2818 0.152939
R13761 gnd.n2820 gnd.n2819 0.152939
R13762 gnd.n2821 gnd.n2820 0.152939
R13763 gnd.n2822 gnd.n2821 0.152939
R13764 gnd.n2823 gnd.n2822 0.152939
R13765 gnd.n2824 gnd.n2823 0.152939
R13766 gnd.n2825 gnd.n2824 0.152939
R13767 gnd.n2826 gnd.n2825 0.152939
R13768 gnd.n2827 gnd.n2826 0.152939
R13769 gnd.n2828 gnd.n2827 0.152939
R13770 gnd.n2829 gnd.n2828 0.152939
R13771 gnd.n2829 gnd.n2528 0.152939
R13772 gnd.n2946 gnd.n2528 0.152939
R13773 gnd.n2947 gnd.n2946 0.152939
R13774 gnd.n2948 gnd.n2947 0.152939
R13775 gnd.n2949 gnd.n2948 0.152939
R13776 gnd.n2949 gnd.n2450 0.152939
R13777 gnd.n3026 gnd.n2450 0.152939
R13778 gnd.n2702 gnd.n2701 0.152939
R13779 gnd.n2703 gnd.n2702 0.152939
R13780 gnd.n2704 gnd.n2703 0.152939
R13781 gnd.n2705 gnd.n2704 0.152939
R13782 gnd.n2706 gnd.n2705 0.152939
R13783 gnd.n2707 gnd.n2706 0.152939
R13784 gnd.n2708 gnd.n2707 0.152939
R13785 gnd.n2709 gnd.n2708 0.152939
R13786 gnd.n2710 gnd.n2709 0.152939
R13787 gnd.n2711 gnd.n2710 0.152939
R13788 gnd.n2712 gnd.n2711 0.152939
R13789 gnd.n2713 gnd.n2712 0.152939
R13790 gnd.n2714 gnd.n2713 0.152939
R13791 gnd.n2715 gnd.n2714 0.152939
R13792 gnd.n2716 gnd.n2715 0.152939
R13793 gnd.n2717 gnd.n2716 0.152939
R13794 gnd.n2718 gnd.n2717 0.152939
R13795 gnd.n2719 gnd.n2718 0.152939
R13796 gnd.n2720 gnd.n2719 0.152939
R13797 gnd.n2721 gnd.n2720 0.152939
R13798 gnd.n2722 gnd.n2721 0.152939
R13799 gnd.n2723 gnd.n2722 0.152939
R13800 gnd.n2727 gnd.n2723 0.152939
R13801 gnd.n2728 gnd.n2727 0.152939
R13802 gnd.n2728 gnd.n2685 0.152939
R13803 gnd.n2782 gnd.n2685 0.152939
R13804 gnd.n3777 gnd.n2155 0.152939
R13805 gnd.n3778 gnd.n3777 0.152939
R13806 gnd.n3779 gnd.n3778 0.152939
R13807 gnd.n3779 gnd.n3769 0.152939
R13808 gnd.n3787 gnd.n3769 0.152939
R13809 gnd.n3788 gnd.n3787 0.152939
R13810 gnd.n3789 gnd.n3788 0.152939
R13811 gnd.n3789 gnd.n3765 0.152939
R13812 gnd.n3797 gnd.n3765 0.152939
R13813 gnd.n3798 gnd.n3797 0.152939
R13814 gnd.n3799 gnd.n3798 0.152939
R13815 gnd.n3799 gnd.n3761 0.152939
R13816 gnd.n3807 gnd.n3761 0.152939
R13817 gnd.n3808 gnd.n3807 0.152939
R13818 gnd.n3809 gnd.n3808 0.152939
R13819 gnd.n3809 gnd.n3754 0.152939
R13820 gnd.n3817 gnd.n3754 0.152939
R13821 gnd.n3818 gnd.n3817 0.152939
R13822 gnd.n3819 gnd.n3818 0.152939
R13823 gnd.n3819 gnd.n3750 0.152939
R13824 gnd.n3827 gnd.n3750 0.152939
R13825 gnd.n3828 gnd.n3827 0.152939
R13826 gnd.n3829 gnd.n3828 0.152939
R13827 gnd.n3829 gnd.n3746 0.152939
R13828 gnd.n3837 gnd.n3746 0.152939
R13829 gnd.n3838 gnd.n3837 0.152939
R13830 gnd.n3839 gnd.n3838 0.152939
R13831 gnd.n3839 gnd.n3742 0.152939
R13832 gnd.n3847 gnd.n3742 0.152939
R13833 gnd.n3848 gnd.n3847 0.152939
R13834 gnd.n3849 gnd.n3848 0.152939
R13835 gnd.n3849 gnd.n3738 0.152939
R13836 gnd.n3857 gnd.n3738 0.152939
R13837 gnd.n3858 gnd.n3857 0.152939
R13838 gnd.n3860 gnd.n3858 0.152939
R13839 gnd.n3860 gnd.n3859 0.152939
R13840 gnd.n3859 gnd.n3731 0.152939
R13841 gnd.n3869 gnd.n3731 0.152939
R13842 gnd.n4107 gnd.n4106 0.152939
R13843 gnd.n4108 gnd.n4107 0.152939
R13844 gnd.n4108 gnd.n2140 0.152939
R13845 gnd.n4122 gnd.n2140 0.152939
R13846 gnd.n4123 gnd.n4122 0.152939
R13847 gnd.n4124 gnd.n4123 0.152939
R13848 gnd.n4124 gnd.n2123 0.152939
R13849 gnd.n4138 gnd.n2123 0.152939
R13850 gnd.n4139 gnd.n4138 0.152939
R13851 gnd.n4140 gnd.n4139 0.152939
R13852 gnd.n4140 gnd.n2108 0.152939
R13853 gnd.n4154 gnd.n2108 0.152939
R13854 gnd.n4155 gnd.n4154 0.152939
R13855 gnd.n4156 gnd.n4155 0.152939
R13856 gnd.n4156 gnd.n2091 0.152939
R13857 gnd.n4170 gnd.n2091 0.152939
R13858 gnd.n4171 gnd.n4170 0.152939
R13859 gnd.n4172 gnd.n4171 0.152939
R13860 gnd.n4172 gnd.n2076 0.152939
R13861 gnd.n4186 gnd.n2076 0.152939
R13862 gnd.n4187 gnd.n4186 0.152939
R13863 gnd.n4188 gnd.n4187 0.152939
R13864 gnd.n4188 gnd.n2059 0.152939
R13865 gnd.n4202 gnd.n2059 0.152939
R13866 gnd.n4203 gnd.n4202 0.152939
R13867 gnd.n4204 gnd.n4203 0.152939
R13868 gnd.n4204 gnd.n2044 0.152939
R13869 gnd.n4252 gnd.n4251 0.152939
R13870 gnd.n4252 gnd.n1993 0.152939
R13871 gnd.n4276 gnd.n1993 0.152939
R13872 gnd.n4277 gnd.n4276 0.152939
R13873 gnd.n4279 gnd.n4277 0.152939
R13874 gnd.n4279 gnd.n4278 0.152939
R13875 gnd.n4278 gnd.n988 0.152939
R13876 gnd.n989 gnd.n988 0.152939
R13877 gnd.n990 gnd.n989 0.152939
R13878 gnd.n1009 gnd.n990 0.152939
R13879 gnd.n1010 gnd.n1009 0.152939
R13880 gnd.n1011 gnd.n1010 0.152939
R13881 gnd.n1012 gnd.n1011 0.152939
R13882 gnd.n1030 gnd.n1012 0.152939
R13883 gnd.n1031 gnd.n1030 0.152939
R13884 gnd.n1032 gnd.n1031 0.152939
R13885 gnd.n1033 gnd.n1032 0.152939
R13886 gnd.n1051 gnd.n1033 0.152939
R13887 gnd.n1052 gnd.n1051 0.152939
R13888 gnd.n1053 gnd.n1052 0.152939
R13889 gnd.n1054 gnd.n1053 0.152939
R13890 gnd.n1073 gnd.n1054 0.152939
R13891 gnd.n1074 gnd.n1073 0.152939
R13892 gnd.n1075 gnd.n1074 0.152939
R13893 gnd.n1076 gnd.n1075 0.152939
R13894 gnd.n1093 gnd.n1076 0.152939
R13895 gnd.n6252 gnd.n1093 0.152939
R13896 gnd.n6251 gnd.n1094 0.152939
R13897 gnd.n1099 gnd.n1094 0.152939
R13898 gnd.n1100 gnd.n1099 0.152939
R13899 gnd.n1101 gnd.n1100 0.152939
R13900 gnd.n1102 gnd.n1101 0.152939
R13901 gnd.n1103 gnd.n1102 0.152939
R13902 gnd.n1107 gnd.n1103 0.152939
R13903 gnd.n1108 gnd.n1107 0.152939
R13904 gnd.n1109 gnd.n1108 0.152939
R13905 gnd.n1110 gnd.n1109 0.152939
R13906 gnd.n1114 gnd.n1110 0.152939
R13907 gnd.n1115 gnd.n1114 0.152939
R13908 gnd.n1116 gnd.n1115 0.152939
R13909 gnd.n1117 gnd.n1116 0.152939
R13910 gnd.n1124 gnd.n1117 0.152939
R13911 gnd.n1127 gnd.n1126 0.152939
R13912 gnd.n1128 gnd.n1127 0.152939
R13913 gnd.n1132 gnd.n1128 0.152939
R13914 gnd.n1133 gnd.n1132 0.152939
R13915 gnd.n1134 gnd.n1133 0.152939
R13916 gnd.n1135 gnd.n1134 0.152939
R13917 gnd.n1139 gnd.n1135 0.152939
R13918 gnd.n1140 gnd.n1139 0.152939
R13919 gnd.n1141 gnd.n1140 0.152939
R13920 gnd.n1142 gnd.n1141 0.152939
R13921 gnd.n1146 gnd.n1142 0.152939
R13922 gnd.n1147 gnd.n1146 0.152939
R13923 gnd.n1148 gnd.n1147 0.152939
R13924 gnd.n1149 gnd.n1148 0.152939
R13925 gnd.n1153 gnd.n1149 0.152939
R13926 gnd.n1154 gnd.n1153 0.152939
R13927 gnd.n1155 gnd.n1154 0.152939
R13928 gnd.n1156 gnd.n1155 0.152939
R13929 gnd.n1161 gnd.n1156 0.152939
R13930 gnd.n6183 gnd.n1161 0.152939
R13931 gnd.n3874 gnd.n3870 0.152939
R13932 gnd.n3875 gnd.n3874 0.152939
R13933 gnd.n3876 gnd.n3875 0.152939
R13934 gnd.n3876 gnd.n3729 0.152939
R13935 gnd.n3882 gnd.n3729 0.152939
R13936 gnd.n3883 gnd.n3882 0.152939
R13937 gnd.n3884 gnd.n3883 0.152939
R13938 gnd.n3884 gnd.n3727 0.152939
R13939 gnd.n3890 gnd.n3727 0.152939
R13940 gnd.n3891 gnd.n3890 0.152939
R13941 gnd.n3892 gnd.n3891 0.152939
R13942 gnd.n3892 gnd.n3725 0.152939
R13943 gnd.n3898 gnd.n3725 0.152939
R13944 gnd.n3899 gnd.n3898 0.152939
R13945 gnd.n3900 gnd.n3899 0.152939
R13946 gnd.n3900 gnd.n3723 0.152939
R13947 gnd.n3906 gnd.n3723 0.152939
R13948 gnd.n3907 gnd.n3906 0.152939
R13949 gnd.n3908 gnd.n3907 0.152939
R13950 gnd.n3908 gnd.n3721 0.152939
R13951 gnd.n3914 gnd.n3721 0.152939
R13952 gnd.n3915 gnd.n3914 0.152939
R13953 gnd.n3916 gnd.n3915 0.152939
R13954 gnd.n3916 gnd.n3719 0.152939
R13955 gnd.n3922 gnd.n3719 0.152939
R13956 gnd.n3923 gnd.n3922 0.152939
R13957 gnd.n3924 gnd.n3923 0.152939
R13958 gnd.n3924 gnd.n3717 0.152939
R13959 gnd.n3930 gnd.n3717 0.152939
R13960 gnd.n3931 gnd.n3930 0.152939
R13961 gnd.n3932 gnd.n3931 0.152939
R13962 gnd.n3932 gnd.n2035 0.152939
R13963 gnd.n3936 gnd.n2035 0.152939
R13964 gnd.n3936 gnd.n3715 0.152939
R13965 gnd.n3942 gnd.n3715 0.152939
R13966 gnd.n3943 gnd.n3942 0.152939
R13967 gnd.n3944 gnd.n3943 0.152939
R13968 gnd.n3944 gnd.n3713 0.152939
R13969 gnd.n3950 gnd.n3713 0.152939
R13970 gnd.n3951 gnd.n3950 0.152939
R13971 gnd.n3952 gnd.n3951 0.152939
R13972 gnd.n3952 gnd.n3711 0.152939
R13973 gnd.n3958 gnd.n3711 0.152939
R13974 gnd.n3959 gnd.n3958 0.152939
R13975 gnd.n3960 gnd.n3959 0.152939
R13976 gnd.n3960 gnd.n3709 0.152939
R13977 gnd.n3970 gnd.n3709 0.152939
R13978 gnd.n3971 gnd.n3970 0.152939
R13979 gnd.n3972 gnd.n3971 0.152939
R13980 gnd.n3973 gnd.n3972 0.152939
R13981 gnd.n3975 gnd.n3973 0.152939
R13982 gnd.n3975 gnd.n3974 0.152939
R13983 gnd.n3974 gnd.n1932 0.152939
R13984 gnd.n1932 gnd.n1930 0.152939
R13985 gnd.n4576 gnd.n1930 0.152939
R13986 gnd.n4577 gnd.n4576 0.152939
R13987 gnd.n4578 gnd.n4577 0.152939
R13988 gnd.n4578 gnd.n1928 0.152939
R13989 gnd.n4586 gnd.n1928 0.152939
R13990 gnd.n4587 gnd.n4586 0.152939
R13991 gnd.n4589 gnd.n4587 0.152939
R13992 gnd.n4589 gnd.n4588 0.152939
R13993 gnd.n4588 gnd.n1162 0.152939
R13994 gnd.n6182 gnd.n1162 0.152939
R13995 gnd.n4058 gnd.n3662 0.152939
R13996 gnd.n3663 gnd.n3662 0.152939
R13997 gnd.n3664 gnd.n3663 0.152939
R13998 gnd.n3665 gnd.n3664 0.152939
R13999 gnd.n3666 gnd.n3665 0.152939
R14000 gnd.n3667 gnd.n3666 0.152939
R14001 gnd.n3668 gnd.n3667 0.152939
R14002 gnd.n3669 gnd.n3668 0.152939
R14003 gnd.n3670 gnd.n3669 0.152939
R14004 gnd.n3671 gnd.n3670 0.152939
R14005 gnd.n3672 gnd.n3671 0.152939
R14006 gnd.n3673 gnd.n3672 0.152939
R14007 gnd.n3674 gnd.n3673 0.152939
R14008 gnd.n3675 gnd.n3674 0.152939
R14009 gnd.n3676 gnd.n3675 0.152939
R14010 gnd.n3677 gnd.n3676 0.152939
R14011 gnd.n3678 gnd.n3677 0.152939
R14012 gnd.n3679 gnd.n3678 0.152939
R14013 gnd.n3680 gnd.n3679 0.152939
R14014 gnd.n3681 gnd.n3680 0.152939
R14015 gnd.n3682 gnd.n3681 0.152939
R14016 gnd.n3683 gnd.n3682 0.152939
R14017 gnd.n3684 gnd.n3683 0.152939
R14018 gnd.n3685 gnd.n3684 0.152939
R14019 gnd.n3686 gnd.n3685 0.152939
R14020 gnd.n3687 gnd.n3686 0.152939
R14021 gnd.n3688 gnd.n3687 0.152939
R14022 gnd.n3689 gnd.n3688 0.152939
R14023 gnd.n3690 gnd.n3689 0.152939
R14024 gnd.n3691 gnd.n3690 0.152939
R14025 gnd.n3692 gnd.n3691 0.152939
R14026 gnd.n4099 gnd.n3636 0.152939
R14027 gnd.n3639 gnd.n3636 0.152939
R14028 gnd.n3640 gnd.n3639 0.152939
R14029 gnd.n3641 gnd.n3640 0.152939
R14030 gnd.n3642 gnd.n3641 0.152939
R14031 gnd.n3645 gnd.n3642 0.152939
R14032 gnd.n3646 gnd.n3645 0.152939
R14033 gnd.n3647 gnd.n3646 0.152939
R14034 gnd.n3648 gnd.n3647 0.152939
R14035 gnd.n3651 gnd.n3648 0.152939
R14036 gnd.n3652 gnd.n3651 0.152939
R14037 gnd.n3653 gnd.n3652 0.152939
R14038 gnd.n3654 gnd.n3653 0.152939
R14039 gnd.n3657 gnd.n3654 0.152939
R14040 gnd.n3658 gnd.n3657 0.152939
R14041 gnd.n4065 gnd.n3658 0.152939
R14042 gnd.n4065 gnd.n4064 0.152939
R14043 gnd.n4064 gnd.n4063 0.152939
R14044 gnd.n4100 gnd.n2148 0.152939
R14045 gnd.n4114 gnd.n2148 0.152939
R14046 gnd.n4115 gnd.n4114 0.152939
R14047 gnd.n4116 gnd.n4115 0.152939
R14048 gnd.n4116 gnd.n2132 0.152939
R14049 gnd.n4130 gnd.n2132 0.152939
R14050 gnd.n4131 gnd.n4130 0.152939
R14051 gnd.n4132 gnd.n4131 0.152939
R14052 gnd.n4132 gnd.n2116 0.152939
R14053 gnd.n4146 gnd.n2116 0.152939
R14054 gnd.n4147 gnd.n4146 0.152939
R14055 gnd.n4148 gnd.n4147 0.152939
R14056 gnd.n4148 gnd.n2100 0.152939
R14057 gnd.n4162 gnd.n2100 0.152939
R14058 gnd.n4163 gnd.n4162 0.152939
R14059 gnd.n4164 gnd.n4163 0.152939
R14060 gnd.n4164 gnd.n2084 0.152939
R14061 gnd.n4178 gnd.n2084 0.152939
R14062 gnd.n4179 gnd.n4178 0.152939
R14063 gnd.n4180 gnd.n4179 0.152939
R14064 gnd.n4180 gnd.n2068 0.152939
R14065 gnd.n4194 gnd.n2068 0.152939
R14066 gnd.n4195 gnd.n4194 0.152939
R14067 gnd.n4196 gnd.n4195 0.152939
R14068 gnd.n4196 gnd.n2052 0.152939
R14069 gnd.n4210 gnd.n2052 0.152939
R14070 gnd.n4211 gnd.n4210 0.152939
R14071 gnd.n4212 gnd.n4211 0.152939
R14072 gnd.n4212 gnd.n2036 0.152939
R14073 gnd.n4226 gnd.n2036 0.152939
R14074 gnd.n4227 gnd.n4226 0.152939
R14075 gnd.n4228 gnd.n4227 0.152939
R14076 gnd.n4228 gnd.n2018 0.152939
R14077 gnd.n4242 gnd.n2018 0.152939
R14078 gnd.n4243 gnd.n4242 0.152939
R14079 gnd.n4244 gnd.n4243 0.152939
R14080 gnd.n4244 gnd.n2003 0.152939
R14081 gnd.n4258 gnd.n2003 0.152939
R14082 gnd.n4259 gnd.n4258 0.152939
R14083 gnd.n4260 gnd.n4259 0.152939
R14084 gnd.n4261 gnd.n4260 0.152939
R14085 gnd.n4262 gnd.n4261 0.152939
R14086 gnd.n4263 gnd.n4262 0.152939
R14087 gnd.n4265 gnd.n4263 0.152939
R14088 gnd.n4265 gnd.n4264 0.152939
R14089 gnd.n4264 gnd.n999 0.152939
R14090 gnd.n1000 gnd.n999 0.152939
R14091 gnd.n1001 gnd.n1000 0.152939
R14092 gnd.n1020 gnd.n1001 0.152939
R14093 gnd.n1021 gnd.n1020 0.152939
R14094 gnd.n1022 gnd.n1021 0.152939
R14095 gnd.n1023 gnd.n1022 0.152939
R14096 gnd.n1040 gnd.n1023 0.152939
R14097 gnd.n1041 gnd.n1040 0.152939
R14098 gnd.n1042 gnd.n1041 0.152939
R14099 gnd.n1043 gnd.n1042 0.152939
R14100 gnd.n1062 gnd.n1043 0.152939
R14101 gnd.n1063 gnd.n1062 0.152939
R14102 gnd.n1064 gnd.n1063 0.152939
R14103 gnd.n1065 gnd.n1064 0.152939
R14104 gnd.n1083 gnd.n1065 0.152939
R14105 gnd.n1084 gnd.n1083 0.152939
R14106 gnd.n1085 gnd.n1084 0.152939
R14107 gnd.n1086 gnd.n1085 0.152939
R14108 gnd.n5967 gnd.n5933 0.152939
R14109 gnd.n5963 gnd.n5933 0.152939
R14110 gnd.n5963 gnd.n5962 0.152939
R14111 gnd.n5962 gnd.n5961 0.152939
R14112 gnd.n5961 gnd.n5942 0.152939
R14113 gnd.n5954 gnd.n5942 0.152939
R14114 gnd.n5954 gnd.n5953 0.152939
R14115 gnd.n5953 gnd.n5952 0.152939
R14116 gnd.n5952 gnd.n5948 0.152939
R14117 gnd.n6155 gnd.n1187 0.152939
R14118 gnd.n6151 gnd.n1187 0.152939
R14119 gnd.n6151 gnd.n6150 0.152939
R14120 gnd.n6150 gnd.n6149 0.152939
R14121 gnd.n6149 gnd.n1192 0.152939
R14122 gnd.n6145 gnd.n1192 0.152939
R14123 gnd.n6145 gnd.n6144 0.152939
R14124 gnd.n6144 gnd.n6143 0.152939
R14125 gnd.n6143 gnd.n1197 0.152939
R14126 gnd.n6139 gnd.n1197 0.152939
R14127 gnd.n6139 gnd.n6138 0.152939
R14128 gnd.n6138 gnd.n6137 0.152939
R14129 gnd.n6137 gnd.n1202 0.152939
R14130 gnd.n6133 gnd.n1202 0.152939
R14131 gnd.n6133 gnd.n6132 0.152939
R14132 gnd.n6132 gnd.n6131 0.152939
R14133 gnd.n6131 gnd.n1207 0.152939
R14134 gnd.n6127 gnd.n1207 0.152939
R14135 gnd.n6127 gnd.n6126 0.152939
R14136 gnd.n6126 gnd.n6125 0.152939
R14137 gnd.n6125 gnd.n1212 0.152939
R14138 gnd.n6121 gnd.n1212 0.152939
R14139 gnd.n6121 gnd.n6120 0.152939
R14140 gnd.n6120 gnd.n6119 0.152939
R14141 gnd.n6119 gnd.n1217 0.152939
R14142 gnd.n6115 gnd.n1217 0.152939
R14143 gnd.n6115 gnd.n6114 0.152939
R14144 gnd.n6114 gnd.n6113 0.152939
R14145 gnd.n6113 gnd.n1222 0.152939
R14146 gnd.n6109 gnd.n1222 0.152939
R14147 gnd.n6109 gnd.n6108 0.152939
R14148 gnd.n6108 gnd.n6107 0.152939
R14149 gnd.n6107 gnd.n1227 0.152939
R14150 gnd.n6103 gnd.n1227 0.152939
R14151 gnd.n6103 gnd.n6102 0.152939
R14152 gnd.n6102 gnd.n6101 0.152939
R14153 gnd.n6101 gnd.n1232 0.152939
R14154 gnd.n6097 gnd.n1232 0.152939
R14155 gnd.n6097 gnd.n6096 0.152939
R14156 gnd.n6096 gnd.n6095 0.152939
R14157 gnd.n6095 gnd.n1237 0.152939
R14158 gnd.n6091 gnd.n1237 0.152939
R14159 gnd.n6091 gnd.n6090 0.152939
R14160 gnd.n6090 gnd.n6089 0.152939
R14161 gnd.n6089 gnd.n1242 0.152939
R14162 gnd.n6085 gnd.n1242 0.152939
R14163 gnd.n6085 gnd.n6084 0.152939
R14164 gnd.n6084 gnd.n6083 0.152939
R14165 gnd.n6083 gnd.n1247 0.152939
R14166 gnd.n6079 gnd.n1247 0.152939
R14167 gnd.n6079 gnd.n6078 0.152939
R14168 gnd.n6078 gnd.n6077 0.152939
R14169 gnd.n6077 gnd.n1252 0.152939
R14170 gnd.n6073 gnd.n1252 0.152939
R14171 gnd.n6073 gnd.n6072 0.152939
R14172 gnd.n6072 gnd.n6071 0.152939
R14173 gnd.n6071 gnd.n1257 0.152939
R14174 gnd.n6067 gnd.n1257 0.152939
R14175 gnd.n6067 gnd.n6066 0.152939
R14176 gnd.n6066 gnd.n6065 0.152939
R14177 gnd.n6065 gnd.n1262 0.152939
R14178 gnd.n6061 gnd.n1262 0.152939
R14179 gnd.n6061 gnd.n6060 0.152939
R14180 gnd.n6060 gnd.n6059 0.152939
R14181 gnd.n6059 gnd.n1267 0.152939
R14182 gnd.n6055 gnd.n1267 0.152939
R14183 gnd.n6055 gnd.n6054 0.152939
R14184 gnd.n6054 gnd.n6053 0.152939
R14185 gnd.n6053 gnd.n1272 0.152939
R14186 gnd.n6049 gnd.n1272 0.152939
R14187 gnd.n6049 gnd.n6048 0.152939
R14188 gnd.n6048 gnd.n6047 0.152939
R14189 gnd.n6047 gnd.n1277 0.152939
R14190 gnd.n6043 gnd.n1277 0.152939
R14191 gnd.n6043 gnd.n6042 0.152939
R14192 gnd.n6042 gnd.n6041 0.152939
R14193 gnd.n6041 gnd.n1282 0.152939
R14194 gnd.n6037 gnd.n1282 0.152939
R14195 gnd.n6037 gnd.n6036 0.152939
R14196 gnd.n6036 gnd.n6035 0.152939
R14197 gnd.n6035 gnd.n1287 0.152939
R14198 gnd.n6031 gnd.n1287 0.152939
R14199 gnd.n6031 gnd.n6030 0.152939
R14200 gnd.n6030 gnd.n6029 0.152939
R14201 gnd.n6029 gnd.n1292 0.152939
R14202 gnd.n6025 gnd.n1292 0.152939
R14203 gnd.n6025 gnd.n6024 0.152939
R14204 gnd.n6024 gnd.n6023 0.152939
R14205 gnd.n6023 gnd.n1297 0.152939
R14206 gnd.n6019 gnd.n1297 0.152939
R14207 gnd.n6019 gnd.n6018 0.152939
R14208 gnd.n6018 gnd.n6017 0.152939
R14209 gnd.n6017 gnd.n1302 0.152939
R14210 gnd.n6013 gnd.n1302 0.152939
R14211 gnd.n6013 gnd.n6012 0.152939
R14212 gnd.n6012 gnd.n6011 0.152939
R14213 gnd.n6011 gnd.n1307 0.152939
R14214 gnd.n6007 gnd.n1307 0.152939
R14215 gnd.n6007 gnd.n6006 0.152939
R14216 gnd.n6006 gnd.n6005 0.152939
R14217 gnd.n6005 gnd.n1312 0.152939
R14218 gnd.n6168 gnd.n1168 0.152939
R14219 gnd.n6168 gnd.n6167 0.152939
R14220 gnd.n6167 gnd.n6166 0.152939
R14221 gnd.n6166 gnd.n1175 0.152939
R14222 gnd.n6162 gnd.n1175 0.152939
R14223 gnd.n6162 gnd.n6161 0.152939
R14224 gnd.n6161 gnd.n1182 0.152939
R14225 gnd.n6157 gnd.n1182 0.152939
R14226 gnd.n6157 gnd.n6156 0.152939
R14227 gnd.n4007 gnd.n4006 0.152939
R14228 gnd.n4006 gnd.n3695 0.152939
R14229 gnd.n4002 gnd.n3695 0.152939
R14230 gnd.n4002 gnd.n4001 0.152939
R14231 gnd.n4001 gnd.n4000 0.152939
R14232 gnd.n4000 gnd.n3699 0.152939
R14233 gnd.n3996 gnd.n3699 0.152939
R14234 gnd.n3996 gnd.n3995 0.152939
R14235 gnd.n3995 gnd.n3994 0.152939
R14236 gnd.n3994 gnd.n3703 0.152939
R14237 gnd.n3990 gnd.n3703 0.152939
R14238 gnd.n3990 gnd.n3989 0.152939
R14239 gnd.n3989 gnd.n3988 0.152939
R14240 gnd.n3988 gnd.n3706 0.152939
R14241 gnd.n3984 gnd.n3706 0.152939
R14242 gnd.n3984 gnd.n3983 0.152939
R14243 gnd.n3983 gnd.n1934 0.152939
R14244 gnd.n4566 gnd.n1934 0.152939
R14245 gnd.n4567 gnd.n4566 0.152939
R14246 gnd.n4568 gnd.n4567 0.152939
R14247 gnd.n4568 gnd.n1922 0.152939
R14248 gnd.n4603 gnd.n1922 0.152939
R14249 gnd.n4603 gnd.n4602 0.152939
R14250 gnd.n4602 gnd.n4601 0.152939
R14251 gnd.n4601 gnd.n1923 0.152939
R14252 gnd.n4597 gnd.n1923 0.152939
R14253 gnd.n4597 gnd.n4596 0.152939
R14254 gnd.n4596 gnd.n4595 0.152939
R14255 gnd.n4595 gnd.n1167 0.152939
R14256 gnd.n6175 gnd.n1167 0.152939
R14257 gnd.n6175 gnd.n6174 0.152939
R14258 gnd.n4786 gnd.n1895 0.152939
R14259 gnd.n4787 gnd.n4786 0.152939
R14260 gnd.n4788 gnd.n4787 0.152939
R14261 gnd.n4788 gnd.n1881 0.152939
R14262 gnd.n4805 gnd.n1881 0.152939
R14263 gnd.n4806 gnd.n4805 0.152939
R14264 gnd.n4807 gnd.n4806 0.152939
R14265 gnd.n4807 gnd.n1867 0.152939
R14266 gnd.n4824 gnd.n1867 0.152939
R14267 gnd.n4825 gnd.n4824 0.152939
R14268 gnd.n4826 gnd.n4825 0.152939
R14269 gnd.n4826 gnd.n1853 0.152939
R14270 gnd.n4843 gnd.n1853 0.152939
R14271 gnd.n4844 gnd.n4843 0.152939
R14272 gnd.n4845 gnd.n4844 0.152939
R14273 gnd.n4845 gnd.n1839 0.152939
R14274 gnd.n4862 gnd.n1839 0.152939
R14275 gnd.n4863 gnd.n4862 0.152939
R14276 gnd.n4864 gnd.n4863 0.152939
R14277 gnd.n4864 gnd.n1825 0.152939
R14278 gnd.n5081 gnd.n1825 0.152939
R14279 gnd.n5082 gnd.n5081 0.152939
R14280 gnd.n5083 gnd.n5082 0.152939
R14281 gnd.n5083 gnd.n1759 0.152939
R14282 gnd.n5115 gnd.n1759 0.152939
R14283 gnd.n5116 gnd.n5115 0.152939
R14284 gnd.n5118 gnd.n5116 0.152939
R14285 gnd.n5118 gnd.n5117 0.152939
R14286 gnd.n5117 gnd.n1730 0.152939
R14287 gnd.n5151 gnd.n1730 0.152939
R14288 gnd.n5152 gnd.n5151 0.152939
R14289 gnd.n5153 gnd.n5152 0.152939
R14290 gnd.n5153 gnd.n1710 0.152939
R14291 gnd.n5178 gnd.n1710 0.152939
R14292 gnd.n5179 gnd.n5178 0.152939
R14293 gnd.n5181 gnd.n5179 0.152939
R14294 gnd.n5181 gnd.n5180 0.152939
R14295 gnd.n5180 gnd.n1679 0.152939
R14296 gnd.n5216 gnd.n1679 0.152939
R14297 gnd.n5217 gnd.n5216 0.152939
R14298 gnd.n5219 gnd.n5217 0.152939
R14299 gnd.n5219 gnd.n5218 0.152939
R14300 gnd.n5218 gnd.n1647 0.152939
R14301 gnd.n5269 gnd.n1647 0.152939
R14302 gnd.n5270 gnd.n5269 0.152939
R14303 gnd.n5271 gnd.n5270 0.152939
R14304 gnd.n5271 gnd.n1630 0.152939
R14305 gnd.n5312 gnd.n1630 0.152939
R14306 gnd.n5313 gnd.n5312 0.152939
R14307 gnd.n5321 gnd.n5313 0.152939
R14308 gnd.n5321 gnd.n5320 0.152939
R14309 gnd.n5320 gnd.n5319 0.152939
R14310 gnd.n5319 gnd.n5314 0.152939
R14311 gnd.n5314 gnd.n1595 0.152939
R14312 gnd.n5380 gnd.n1595 0.152939
R14313 gnd.n5381 gnd.n5380 0.152939
R14314 gnd.n5386 gnd.n5381 0.152939
R14315 gnd.n5386 gnd.n5385 0.152939
R14316 gnd.n5385 gnd.n5384 0.152939
R14317 gnd.n5384 gnd.n1572 0.152939
R14318 gnd.n5428 gnd.n1572 0.152939
R14319 gnd.n5428 gnd.n5427 0.152939
R14320 gnd.n5427 gnd.n5426 0.152939
R14321 gnd.n5426 gnd.n1550 0.152939
R14322 gnd.n5478 gnd.n1550 0.152939
R14323 gnd.n5478 gnd.n5477 0.152939
R14324 gnd.n5477 gnd.n5476 0.152939
R14325 gnd.n5476 gnd.n1522 0.152939
R14326 gnd.n5509 gnd.n1522 0.152939
R14327 gnd.n5510 gnd.n5509 0.152939
R14328 gnd.n5511 gnd.n5510 0.152939
R14329 gnd.n5511 gnd.n1501 0.152939
R14330 gnd.n5557 gnd.n1501 0.152939
R14331 gnd.n5557 gnd.n5556 0.152939
R14332 gnd.n5556 gnd.n5555 0.152939
R14333 gnd.n5555 gnd.n1502 0.152939
R14334 gnd.n5551 gnd.n1502 0.152939
R14335 gnd.n5551 gnd.n1389 0.152939
R14336 gnd.n5728 gnd.n1389 0.152939
R14337 gnd.n5729 gnd.n5728 0.152939
R14338 gnd.n5730 gnd.n5729 0.152939
R14339 gnd.n5730 gnd.n1376 0.152939
R14340 gnd.n5747 gnd.n1376 0.152939
R14341 gnd.n5748 gnd.n5747 0.152939
R14342 gnd.n5749 gnd.n5748 0.152939
R14343 gnd.n5749 gnd.n1362 0.152939
R14344 gnd.n5766 gnd.n1362 0.152939
R14345 gnd.n5767 gnd.n5766 0.152939
R14346 gnd.n5768 gnd.n5767 0.152939
R14347 gnd.n5768 gnd.n1348 0.152939
R14348 gnd.n5785 gnd.n1348 0.152939
R14349 gnd.n5786 gnd.n5785 0.152939
R14350 gnd.n5787 gnd.n5786 0.152939
R14351 gnd.n5787 gnd.n1334 0.152939
R14352 gnd.n5804 gnd.n1334 0.152939
R14353 gnd.n5805 gnd.n5804 0.152939
R14354 gnd.n5806 gnd.n5805 0.152939
R14355 gnd.n5806 gnd.n1319 0.152939
R14356 gnd.n5996 gnd.n1319 0.152939
R14357 gnd.n5997 gnd.n5996 0.152939
R14358 gnd.n5998 gnd.n5997 0.152939
R14359 gnd.n7230 gnd.n445 0.152939
R14360 gnd.n7244 gnd.n445 0.152939
R14361 gnd.n7245 gnd.n7244 0.152939
R14362 gnd.n7246 gnd.n7245 0.152939
R14363 gnd.n7246 gnd.n427 0.152939
R14364 gnd.n7260 gnd.n427 0.152939
R14365 gnd.n7261 gnd.n7260 0.152939
R14366 gnd.n7262 gnd.n7261 0.152939
R14367 gnd.n7262 gnd.n410 0.152939
R14368 gnd.n7276 gnd.n410 0.152939
R14369 gnd.n7277 gnd.n7276 0.152939
R14370 gnd.n7278 gnd.n7277 0.152939
R14371 gnd.n7278 gnd.n393 0.152939
R14372 gnd.n7292 gnd.n393 0.152939
R14373 gnd.n7293 gnd.n7292 0.152939
R14374 gnd.n7294 gnd.n7293 0.152939
R14375 gnd.n7294 gnd.n376 0.152939
R14376 gnd.n7308 gnd.n376 0.152939
R14377 gnd.n7309 gnd.n7308 0.152939
R14378 gnd.n7310 gnd.n7309 0.152939
R14379 gnd.n7310 gnd.n359 0.152939
R14380 gnd.n7324 gnd.n359 0.152939
R14381 gnd.n7325 gnd.n7324 0.152939
R14382 gnd.n7326 gnd.n7325 0.152939
R14383 gnd.n7326 gnd.n343 0.152939
R14384 gnd.n7340 gnd.n343 0.152939
R14385 gnd.n7341 gnd.n7340 0.152939
R14386 gnd.n7342 gnd.n7341 0.152939
R14387 gnd.n7342 gnd.n327 0.152939
R14388 gnd.n7356 gnd.n327 0.152939
R14389 gnd.n7357 gnd.n7356 0.152939
R14390 gnd.n7358 gnd.n7357 0.152939
R14391 gnd.n7358 gnd.n310 0.152939
R14392 gnd.n7372 gnd.n310 0.152939
R14393 gnd.n7373 gnd.n7372 0.152939
R14394 gnd.n7374 gnd.n7373 0.152939
R14395 gnd.n7374 gnd.n296 0.152939
R14396 gnd.n7388 gnd.n296 0.152939
R14397 gnd.n7389 gnd.n7388 0.152939
R14398 gnd.n7390 gnd.n7389 0.152939
R14399 gnd.n7390 gnd.n280 0.152939
R14400 gnd.n7404 gnd.n280 0.152939
R14401 gnd.n7405 gnd.n7404 0.152939
R14402 gnd.n7406 gnd.n7405 0.152939
R14403 gnd.n7406 gnd.n266 0.152939
R14404 gnd.n7420 gnd.n266 0.152939
R14405 gnd.n7421 gnd.n7420 0.152939
R14406 gnd.n7422 gnd.n7421 0.152939
R14407 gnd.n7422 gnd.n249 0.152939
R14408 gnd.n7436 gnd.n249 0.152939
R14409 gnd.n7437 gnd.n7436 0.152939
R14410 gnd.n7438 gnd.n7437 0.152939
R14411 gnd.n7438 gnd.n235 0.152939
R14412 gnd.n7452 gnd.n235 0.152939
R14413 gnd.n7453 gnd.n7452 0.152939
R14414 gnd.n7454 gnd.n7453 0.152939
R14415 gnd.n7454 gnd.n220 0.152939
R14416 gnd.n7468 gnd.n220 0.152939
R14417 gnd.n7469 gnd.n7468 0.152939
R14418 gnd.n7538 gnd.n7469 0.152939
R14419 gnd.n7538 gnd.n7537 0.152939
R14420 gnd.n7537 gnd.n7536 0.152939
R14421 gnd.n7536 gnd.n7470 0.152939
R14422 gnd.n7532 gnd.n7470 0.152939
R14423 gnd.n7531 gnd.n7472 0.152939
R14424 gnd.n7527 gnd.n7472 0.152939
R14425 gnd.n7527 gnd.n7526 0.152939
R14426 gnd.n7526 gnd.n7525 0.152939
R14427 gnd.n7525 gnd.n7478 0.152939
R14428 gnd.n7521 gnd.n7478 0.152939
R14429 gnd.n7521 gnd.n7520 0.152939
R14430 gnd.n7520 gnd.n7519 0.152939
R14431 gnd.n7519 gnd.n7486 0.152939
R14432 gnd.n7515 gnd.n7486 0.152939
R14433 gnd.n7515 gnd.n7514 0.152939
R14434 gnd.n7514 gnd.n7513 0.152939
R14435 gnd.n7513 gnd.n7494 0.152939
R14436 gnd.n7509 gnd.n7494 0.152939
R14437 gnd.n7509 gnd.n7508 0.152939
R14438 gnd.n7508 gnd.n7507 0.152939
R14439 gnd.n7507 gnd.n121 0.152939
R14440 gnd.n7633 gnd.n121 0.152939
R14441 gnd.n5970 gnd.n5969 0.152939
R14442 gnd.n5970 gnd.n596 0.152939
R14443 gnd.n7095 gnd.n596 0.152939
R14444 gnd.n7095 gnd.n7094 0.152939
R14445 gnd.n7094 gnd.n7093 0.152939
R14446 gnd.n7093 gnd.n597 0.152939
R14447 gnd.n7089 gnd.n597 0.152939
R14448 gnd.n7089 gnd.n7088 0.152939
R14449 gnd.n7088 gnd.n7087 0.152939
R14450 gnd.n7087 gnd.n601 0.152939
R14451 gnd.n7083 gnd.n601 0.152939
R14452 gnd.n7083 gnd.n7082 0.152939
R14453 gnd.n7082 gnd.n7081 0.152939
R14454 gnd.n7081 gnd.n605 0.152939
R14455 gnd.n7077 gnd.n605 0.152939
R14456 gnd.n7077 gnd.n7076 0.152939
R14457 gnd.n7076 gnd.n7075 0.152939
R14458 gnd.n7075 gnd.n609 0.152939
R14459 gnd.n7071 gnd.n609 0.152939
R14460 gnd.n7071 gnd.n7070 0.152939
R14461 gnd.n7070 gnd.n7069 0.152939
R14462 gnd.n7069 gnd.n7043 0.152939
R14463 gnd.n7065 gnd.n7043 0.152939
R14464 gnd.n7065 gnd.n7064 0.152939
R14465 gnd.n7064 gnd.n7063 0.152939
R14466 gnd.n7063 gnd.n7047 0.152939
R14467 gnd.n7059 gnd.n7047 0.152939
R14468 gnd.n7059 gnd.n7058 0.152939
R14469 gnd.n7058 gnd.n7057 0.152939
R14470 gnd.n7057 gnd.n7051 0.152939
R14471 gnd.n7051 gnd.n79 0.152939
R14472 gnd.n7682 gnd.n79 0.152939
R14473 gnd.n7682 gnd.n7681 0.152939
R14474 gnd.n7681 gnd.n81 0.152939
R14475 gnd.n7677 gnd.n81 0.152939
R14476 gnd.n7677 gnd.n7676 0.152939
R14477 gnd.n7676 gnd.n7675 0.152939
R14478 gnd.n7675 gnd.n86 0.152939
R14479 gnd.n7671 gnd.n86 0.152939
R14480 gnd.n7671 gnd.n7670 0.152939
R14481 gnd.n7670 gnd.n7669 0.152939
R14482 gnd.n7669 gnd.n91 0.152939
R14483 gnd.n7665 gnd.n91 0.152939
R14484 gnd.n7665 gnd.n7664 0.152939
R14485 gnd.n7664 gnd.n7663 0.152939
R14486 gnd.n7663 gnd.n96 0.152939
R14487 gnd.n7659 gnd.n96 0.152939
R14488 gnd.n7659 gnd.n7658 0.152939
R14489 gnd.n7658 gnd.n7657 0.152939
R14490 gnd.n7657 gnd.n101 0.152939
R14491 gnd.n7653 gnd.n101 0.152939
R14492 gnd.n7653 gnd.n7652 0.152939
R14493 gnd.n7652 gnd.n7651 0.152939
R14494 gnd.n7651 gnd.n106 0.152939
R14495 gnd.n7647 gnd.n106 0.152939
R14496 gnd.n7647 gnd.n7646 0.152939
R14497 gnd.n7646 gnd.n7645 0.152939
R14498 gnd.n7645 gnd.n111 0.152939
R14499 gnd.n7641 gnd.n111 0.152939
R14500 gnd.n7641 gnd.n7640 0.152939
R14501 gnd.n7640 gnd.n7639 0.152939
R14502 gnd.n7639 gnd.n116 0.152939
R14503 gnd.n7635 gnd.n116 0.152939
R14504 gnd.n7635 gnd.n7634 0.152939
R14505 gnd.n5968 gnd.n5967 0.151415
R14506 gnd.n6173 gnd.n1168 0.151415
R14507 gnd.n4008 gnd.n3692 0.145814
R14508 gnd.n4008 gnd.n4007 0.145814
R14509 gnd.n3028 gnd.n3027 0.0767195
R14510 gnd.n3027 gnd.n3026 0.0767195
R14511 gnd.n4659 gnd.n4658 0.063
R14512 gnd.n7229 gnd.n460 0.063
R14513 gnd.n3594 gnd.n2198 0.0477147
R14514 gnd.n2791 gnd.n2679 0.0442063
R14515 gnd.n2792 gnd.n2791 0.0442063
R14516 gnd.n2793 gnd.n2792 0.0442063
R14517 gnd.n2793 gnd.n2668 0.0442063
R14518 gnd.n2807 gnd.n2668 0.0442063
R14519 gnd.n2808 gnd.n2807 0.0442063
R14520 gnd.n2809 gnd.n2808 0.0442063
R14521 gnd.n2809 gnd.n2655 0.0442063
R14522 gnd.n2853 gnd.n2655 0.0442063
R14523 gnd.n2854 gnd.n2853 0.0442063
R14524 gnd.n2856 gnd.n2589 0.0344674
R14525 gnd.n5932 gnd.n509 0.0343753
R14526 gnd.n6172 gnd.n1169 0.0343753
R14527 gnd.n2876 gnd.n2875 0.0269946
R14528 gnd.n2878 gnd.n2877 0.0269946
R14529 gnd.n2584 gnd.n2582 0.0269946
R14530 gnd.n2888 gnd.n2886 0.0269946
R14531 gnd.n2887 gnd.n2563 0.0269946
R14532 gnd.n2907 gnd.n2906 0.0269946
R14533 gnd.n2909 gnd.n2908 0.0269946
R14534 gnd.n2558 gnd.n2557 0.0269946
R14535 gnd.n2919 gnd.n2553 0.0269946
R14536 gnd.n2918 gnd.n2555 0.0269946
R14537 gnd.n2554 gnd.n2536 0.0269946
R14538 gnd.n2939 gnd.n2537 0.0269946
R14539 gnd.n2938 gnd.n2538 0.0269946
R14540 gnd.n2972 gnd.n2513 0.0269946
R14541 gnd.n2974 gnd.n2973 0.0269946
R14542 gnd.n2975 gnd.n2460 0.0269946
R14543 gnd.n2508 gnd.n2461 0.0269946
R14544 gnd.n2510 gnd.n2462 0.0269946
R14545 gnd.n2985 gnd.n2984 0.0269946
R14546 gnd.n2987 gnd.n2986 0.0269946
R14547 gnd.n2988 gnd.n2482 0.0269946
R14548 gnd.n2990 gnd.n2483 0.0269946
R14549 gnd.n2993 gnd.n2484 0.0269946
R14550 gnd.n2996 gnd.n2995 0.0269946
R14551 gnd.n2998 gnd.n2997 0.0269946
R14552 gnd.n3063 gnd.n2371 0.0269946
R14553 gnd.n3065 gnd.n3064 0.0269946
R14554 gnd.n3074 gnd.n2364 0.0269946
R14555 gnd.n3076 gnd.n3075 0.0269946
R14556 gnd.n3077 gnd.n2362 0.0269946
R14557 gnd.n3084 gnd.n3080 0.0269946
R14558 gnd.n3083 gnd.n3082 0.0269946
R14559 gnd.n3081 gnd.n2341 0.0269946
R14560 gnd.n3106 gnd.n2342 0.0269946
R14561 gnd.n3105 gnd.n2343 0.0269946
R14562 gnd.n3148 gnd.n2316 0.0269946
R14563 gnd.n3150 gnd.n3149 0.0269946
R14564 gnd.n3159 gnd.n2309 0.0269946
R14565 gnd.n3161 gnd.n3160 0.0269946
R14566 gnd.n3162 gnd.n2307 0.0269946
R14567 gnd.n3169 gnd.n3165 0.0269946
R14568 gnd.n3168 gnd.n3167 0.0269946
R14569 gnd.n3166 gnd.n2286 0.0269946
R14570 gnd.n3191 gnd.n2287 0.0269946
R14571 gnd.n3190 gnd.n2288 0.0269946
R14572 gnd.n3237 gnd.n2262 0.0269946
R14573 gnd.n3239 gnd.n3238 0.0269946
R14574 gnd.n3248 gnd.n2255 0.0269946
R14575 gnd.n3507 gnd.n2253 0.0269946
R14576 gnd.n3512 gnd.n3510 0.0269946
R14577 gnd.n3511 gnd.n2234 0.0269946
R14578 gnd.n3536 gnd.n3535 0.0269946
R14579 gnd.n7226 gnd.n460 0.0245515
R14580 gnd.n4660 gnd.n4659 0.0245515
R14581 gnd.n2856 gnd.n2855 0.0202011
R14582 gnd.n7226 gnd.n7225 0.0174377
R14583 gnd.n7225 gnd.n463 0.0174377
R14584 gnd.n7222 gnd.n463 0.0174377
R14585 gnd.n7222 gnd.n7221 0.0174377
R14586 gnd.n7221 gnd.n467 0.0174377
R14587 gnd.n7218 gnd.n467 0.0174377
R14588 gnd.n7218 gnd.n7217 0.0174377
R14589 gnd.n7217 gnd.n471 0.0174377
R14590 gnd.n7214 gnd.n471 0.0174377
R14591 gnd.n7214 gnd.n7213 0.0174377
R14592 gnd.n7213 gnd.n475 0.0174377
R14593 gnd.n7210 gnd.n475 0.0174377
R14594 gnd.n7210 gnd.n7209 0.0174377
R14595 gnd.n7209 gnd.n479 0.0174377
R14596 gnd.n7206 gnd.n479 0.0174377
R14597 gnd.n7206 gnd.n7205 0.0174377
R14598 gnd.n7205 gnd.n483 0.0174377
R14599 gnd.n7202 gnd.n483 0.0174377
R14600 gnd.n7202 gnd.n7201 0.0174377
R14601 gnd.n7201 gnd.n487 0.0174377
R14602 gnd.n7198 gnd.n487 0.0174377
R14603 gnd.n7198 gnd.n7197 0.0174377
R14604 gnd.n7197 gnd.n491 0.0174377
R14605 gnd.n7194 gnd.n491 0.0174377
R14606 gnd.n7194 gnd.n7193 0.0174377
R14607 gnd.n7193 gnd.n495 0.0174377
R14608 gnd.n7190 gnd.n495 0.0174377
R14609 gnd.n7190 gnd.n7189 0.0174377
R14610 gnd.n7189 gnd.n499 0.0174377
R14611 gnd.n7186 gnd.n499 0.0174377
R14612 gnd.n7186 gnd.n7185 0.0174377
R14613 gnd.n7185 gnd.n505 0.0174377
R14614 gnd.n7182 gnd.n505 0.0174377
R14615 gnd.n7182 gnd.n7181 0.0174377
R14616 gnd.n7181 gnd.n509 0.0174377
R14617 gnd.n4660 gnd.n4652 0.0174377
R14618 gnd.n4654 gnd.n4652 0.0174377
R14619 gnd.n4766 gnd.n4654 0.0174377
R14620 gnd.n4766 gnd.n4765 0.0174377
R14621 gnd.n4765 gnd.n4655 0.0174377
R14622 gnd.n4762 gnd.n4655 0.0174377
R14623 gnd.n4762 gnd.n4761 0.0174377
R14624 gnd.n4761 gnd.n4669 0.0174377
R14625 gnd.n4758 gnd.n4669 0.0174377
R14626 gnd.n4758 gnd.n4757 0.0174377
R14627 gnd.n4757 gnd.n4674 0.0174377
R14628 gnd.n4754 gnd.n4674 0.0174377
R14629 gnd.n4754 gnd.n4753 0.0174377
R14630 gnd.n4753 gnd.n4680 0.0174377
R14631 gnd.n4750 gnd.n4680 0.0174377
R14632 gnd.n4750 gnd.n4749 0.0174377
R14633 gnd.n4749 gnd.n4684 0.0174377
R14634 gnd.n4746 gnd.n4684 0.0174377
R14635 gnd.n4746 gnd.n4745 0.0174377
R14636 gnd.n4745 gnd.n4691 0.0174377
R14637 gnd.n4742 gnd.n4691 0.0174377
R14638 gnd.n4742 gnd.n4741 0.0174377
R14639 gnd.n4741 gnd.n4697 0.0174377
R14640 gnd.n4738 gnd.n4697 0.0174377
R14641 gnd.n4738 gnd.n4737 0.0174377
R14642 gnd.n4737 gnd.n4703 0.0174377
R14643 gnd.n4734 gnd.n4703 0.0174377
R14644 gnd.n4734 gnd.n4733 0.0174377
R14645 gnd.n4733 gnd.n4707 0.0174377
R14646 gnd.n4730 gnd.n4707 0.0174377
R14647 gnd.n4730 gnd.n4729 0.0174377
R14648 gnd.n4729 gnd.n4716 0.0174377
R14649 gnd.n4726 gnd.n4716 0.0174377
R14650 gnd.n4726 gnd.n4725 0.0174377
R14651 gnd.n4725 gnd.n1169 0.0174377
R14652 gnd.n2855 gnd.n2854 0.0148637
R14653 gnd.n3505 gnd.n3249 0.0144266
R14654 gnd.n3506 gnd.n3505 0.0130679
R14655 gnd.n2875 gnd.n2589 0.00797283
R14656 gnd.n2877 gnd.n2876 0.00797283
R14657 gnd.n2878 gnd.n2584 0.00797283
R14658 gnd.n2886 gnd.n2582 0.00797283
R14659 gnd.n2888 gnd.n2887 0.00797283
R14660 gnd.n2906 gnd.n2563 0.00797283
R14661 gnd.n2908 gnd.n2907 0.00797283
R14662 gnd.n2909 gnd.n2558 0.00797283
R14663 gnd.n2557 gnd.n2553 0.00797283
R14664 gnd.n2919 gnd.n2918 0.00797283
R14665 gnd.n2555 gnd.n2554 0.00797283
R14666 gnd.n2537 gnd.n2536 0.00797283
R14667 gnd.n2939 gnd.n2938 0.00797283
R14668 gnd.n2538 gnd.n2513 0.00797283
R14669 gnd.n2973 gnd.n2972 0.00797283
R14670 gnd.n2975 gnd.n2974 0.00797283
R14671 gnd.n2508 gnd.n2460 0.00797283
R14672 gnd.n2510 gnd.n2461 0.00797283
R14673 gnd.n2984 gnd.n2462 0.00797283
R14674 gnd.n2986 gnd.n2985 0.00797283
R14675 gnd.n2988 gnd.n2987 0.00797283
R14676 gnd.n2990 gnd.n2482 0.00797283
R14677 gnd.n2993 gnd.n2483 0.00797283
R14678 gnd.n2995 gnd.n2484 0.00797283
R14679 gnd.n2998 gnd.n2996 0.00797283
R14680 gnd.n2997 gnd.n2371 0.00797283
R14681 gnd.n3065 gnd.n3063 0.00797283
R14682 gnd.n3064 gnd.n2364 0.00797283
R14683 gnd.n3075 gnd.n3074 0.00797283
R14684 gnd.n3077 gnd.n3076 0.00797283
R14685 gnd.n3080 gnd.n2362 0.00797283
R14686 gnd.n3084 gnd.n3083 0.00797283
R14687 gnd.n3082 gnd.n3081 0.00797283
R14688 gnd.n2342 gnd.n2341 0.00797283
R14689 gnd.n3106 gnd.n3105 0.00797283
R14690 gnd.n2343 gnd.n2316 0.00797283
R14691 gnd.n3150 gnd.n3148 0.00797283
R14692 gnd.n3149 gnd.n2309 0.00797283
R14693 gnd.n3160 gnd.n3159 0.00797283
R14694 gnd.n3162 gnd.n3161 0.00797283
R14695 gnd.n3165 gnd.n2307 0.00797283
R14696 gnd.n3169 gnd.n3168 0.00797283
R14697 gnd.n3167 gnd.n3166 0.00797283
R14698 gnd.n2287 gnd.n2286 0.00797283
R14699 gnd.n3191 gnd.n3190 0.00797283
R14700 gnd.n2288 gnd.n2262 0.00797283
R14701 gnd.n3239 gnd.n3237 0.00797283
R14702 gnd.n3238 gnd.n2255 0.00797283
R14703 gnd.n3249 gnd.n3248 0.00797283
R14704 gnd.n3507 gnd.n3506 0.00797283
R14705 gnd.n3510 gnd.n2253 0.00797283
R14706 gnd.n3512 gnd.n3511 0.00797283
R14707 gnd.n3535 gnd.n2234 0.00797283
R14708 gnd.n3536 gnd.n2198 0.00797283
R14709 gnd.n7358 gnd.n326 0.00433921
R14710 gnd.n4228 gnd.n2035 0.00433921
R14711 gnd.n7348 gnd.n335 0.00335063
R14712 gnd.n7349 gnd.n7348 0.00335063
R14713 gnd.n7350 gnd.n7349 0.00335063
R14714 gnd.n7350 gnd.n317 0.00335063
R14715 gnd.n7364 gnd.n317 0.00335063
R14716 gnd.n7365 gnd.n7364 0.00335063
R14717 gnd.n7366 gnd.n7365 0.00335063
R14718 gnd.n7366 gnd.n303 0.00335063
R14719 gnd.n7380 gnd.n303 0.00335063
R14720 gnd.n7381 gnd.n7380 0.00335063
R14721 gnd.n4218 gnd.n2044 0.00335063
R14722 gnd.n4219 gnd.n4218 0.00335063
R14723 gnd.n4220 gnd.n4219 0.00335063
R14724 gnd.n4220 gnd.n2026 0.00335063
R14725 gnd.n4234 gnd.n2026 0.00335063
R14726 gnd.n4235 gnd.n4234 0.00335063
R14727 gnd.n4236 gnd.n4235 0.00335063
R14728 gnd.n4236 gnd.n2011 0.00335063
R14729 gnd.n4250 gnd.n2011 0.00335063
R14730 gnd.n4251 gnd.n4250 0.00335063
R14731 gnd.n5968 gnd.n5932 0.000838753
R14732 gnd.n6173 gnd.n6172 0.000838753
R14733 vdd.n315 vdd.n279 756.745
R14734 vdd.n260 vdd.n224 756.745
R14735 vdd.n217 vdd.n181 756.745
R14736 vdd.n162 vdd.n126 756.745
R14737 vdd.n120 vdd.n84 756.745
R14738 vdd.n65 vdd.n29 756.745
R14739 vdd.n1684 vdd.n1648 756.745
R14740 vdd.n1739 vdd.n1703 756.745
R14741 vdd.n1586 vdd.n1550 756.745
R14742 vdd.n1641 vdd.n1605 756.745
R14743 vdd.n1489 vdd.n1453 756.745
R14744 vdd.n1544 vdd.n1508 756.745
R14745 vdd.n2094 vdd.t77 640.208
R14746 vdd.n936 vdd.t62 640.208
R14747 vdd.n2068 vdd.t23 640.208
R14748 vdd.n928 vdd.t87 640.208
R14749 vdd.n2839 vdd.t49 640.208
R14750 vdd.n2559 vdd.t84 640.208
R14751 vdd.n804 vdd.t66 640.208
R14752 vdd.n2556 vdd.t70 640.208
R14753 vdd.n768 vdd.t74 640.208
R14754 vdd.n998 vdd.t80 640.208
R14755 vdd.n1148 vdd.t35 592.009
R14756 vdd.n1304 vdd.t46 592.009
R14757 vdd.n1340 vdd.t53 592.009
R14758 vdd.n2250 vdd.t42 592.009
R14759 vdd.n1887 vdd.t56 592.009
R14760 vdd.n1847 vdd.t59 592.009
R14761 vdd.n405 vdd.t31 592.009
R14762 vdd.n419 vdd.t90 592.009
R14763 vdd.n431 vdd.t96 592.009
R14764 vdd.n723 vdd.t27 592.009
R14765 vdd.n686 vdd.t39 592.009
R14766 vdd.n3013 vdd.t93 592.009
R14767 vdd.n316 vdd.n315 585
R14768 vdd.n314 vdd.n281 585
R14769 vdd.n313 vdd.n312 585
R14770 vdd.n284 vdd.n282 585
R14771 vdd.n307 vdd.n306 585
R14772 vdd.n305 vdd.n304 585
R14773 vdd.n288 vdd.n287 585
R14774 vdd.n299 vdd.n298 585
R14775 vdd.n297 vdd.n296 585
R14776 vdd.n292 vdd.n291 585
R14777 vdd.n261 vdd.n260 585
R14778 vdd.n259 vdd.n226 585
R14779 vdd.n258 vdd.n257 585
R14780 vdd.n229 vdd.n227 585
R14781 vdd.n252 vdd.n251 585
R14782 vdd.n250 vdd.n249 585
R14783 vdd.n233 vdd.n232 585
R14784 vdd.n244 vdd.n243 585
R14785 vdd.n242 vdd.n241 585
R14786 vdd.n237 vdd.n236 585
R14787 vdd.n218 vdd.n217 585
R14788 vdd.n216 vdd.n183 585
R14789 vdd.n215 vdd.n214 585
R14790 vdd.n186 vdd.n184 585
R14791 vdd.n209 vdd.n208 585
R14792 vdd.n207 vdd.n206 585
R14793 vdd.n190 vdd.n189 585
R14794 vdd.n201 vdd.n200 585
R14795 vdd.n199 vdd.n198 585
R14796 vdd.n194 vdd.n193 585
R14797 vdd.n163 vdd.n162 585
R14798 vdd.n161 vdd.n128 585
R14799 vdd.n160 vdd.n159 585
R14800 vdd.n131 vdd.n129 585
R14801 vdd.n154 vdd.n153 585
R14802 vdd.n152 vdd.n151 585
R14803 vdd.n135 vdd.n134 585
R14804 vdd.n146 vdd.n145 585
R14805 vdd.n144 vdd.n143 585
R14806 vdd.n139 vdd.n138 585
R14807 vdd.n121 vdd.n120 585
R14808 vdd.n119 vdd.n86 585
R14809 vdd.n118 vdd.n117 585
R14810 vdd.n89 vdd.n87 585
R14811 vdd.n112 vdd.n111 585
R14812 vdd.n110 vdd.n109 585
R14813 vdd.n93 vdd.n92 585
R14814 vdd.n104 vdd.n103 585
R14815 vdd.n102 vdd.n101 585
R14816 vdd.n97 vdd.n96 585
R14817 vdd.n66 vdd.n65 585
R14818 vdd.n64 vdd.n31 585
R14819 vdd.n63 vdd.n62 585
R14820 vdd.n34 vdd.n32 585
R14821 vdd.n57 vdd.n56 585
R14822 vdd.n55 vdd.n54 585
R14823 vdd.n38 vdd.n37 585
R14824 vdd.n49 vdd.n48 585
R14825 vdd.n47 vdd.n46 585
R14826 vdd.n42 vdd.n41 585
R14827 vdd.n1685 vdd.n1684 585
R14828 vdd.n1683 vdd.n1650 585
R14829 vdd.n1682 vdd.n1681 585
R14830 vdd.n1653 vdd.n1651 585
R14831 vdd.n1676 vdd.n1675 585
R14832 vdd.n1674 vdd.n1673 585
R14833 vdd.n1657 vdd.n1656 585
R14834 vdd.n1668 vdd.n1667 585
R14835 vdd.n1666 vdd.n1665 585
R14836 vdd.n1661 vdd.n1660 585
R14837 vdd.n1740 vdd.n1739 585
R14838 vdd.n1738 vdd.n1705 585
R14839 vdd.n1737 vdd.n1736 585
R14840 vdd.n1708 vdd.n1706 585
R14841 vdd.n1731 vdd.n1730 585
R14842 vdd.n1729 vdd.n1728 585
R14843 vdd.n1712 vdd.n1711 585
R14844 vdd.n1723 vdd.n1722 585
R14845 vdd.n1721 vdd.n1720 585
R14846 vdd.n1716 vdd.n1715 585
R14847 vdd.n1587 vdd.n1586 585
R14848 vdd.n1585 vdd.n1552 585
R14849 vdd.n1584 vdd.n1583 585
R14850 vdd.n1555 vdd.n1553 585
R14851 vdd.n1578 vdd.n1577 585
R14852 vdd.n1576 vdd.n1575 585
R14853 vdd.n1559 vdd.n1558 585
R14854 vdd.n1570 vdd.n1569 585
R14855 vdd.n1568 vdd.n1567 585
R14856 vdd.n1563 vdd.n1562 585
R14857 vdd.n1642 vdd.n1641 585
R14858 vdd.n1640 vdd.n1607 585
R14859 vdd.n1639 vdd.n1638 585
R14860 vdd.n1610 vdd.n1608 585
R14861 vdd.n1633 vdd.n1632 585
R14862 vdd.n1631 vdd.n1630 585
R14863 vdd.n1614 vdd.n1613 585
R14864 vdd.n1625 vdd.n1624 585
R14865 vdd.n1623 vdd.n1622 585
R14866 vdd.n1618 vdd.n1617 585
R14867 vdd.n1490 vdd.n1489 585
R14868 vdd.n1488 vdd.n1455 585
R14869 vdd.n1487 vdd.n1486 585
R14870 vdd.n1458 vdd.n1456 585
R14871 vdd.n1481 vdd.n1480 585
R14872 vdd.n1479 vdd.n1478 585
R14873 vdd.n1462 vdd.n1461 585
R14874 vdd.n1473 vdd.n1472 585
R14875 vdd.n1471 vdd.n1470 585
R14876 vdd.n1466 vdd.n1465 585
R14877 vdd.n1545 vdd.n1544 585
R14878 vdd.n1543 vdd.n1510 585
R14879 vdd.n1542 vdd.n1541 585
R14880 vdd.n1513 vdd.n1511 585
R14881 vdd.n1536 vdd.n1535 585
R14882 vdd.n1534 vdd.n1533 585
R14883 vdd.n1517 vdd.n1516 585
R14884 vdd.n1528 vdd.n1527 585
R14885 vdd.n1526 vdd.n1525 585
R14886 vdd.n1521 vdd.n1520 585
R14887 vdd.n445 vdd.n370 462.44
R14888 vdd.n3251 vdd.n372 462.44
R14889 vdd.n3146 vdd.n657 462.44
R14890 vdd.n3144 vdd.n660 462.44
R14891 vdd.n2245 vdd.n1047 462.44
R14892 vdd.n2248 vdd.n2247 462.44
R14893 vdd.n1375 vdd.n1145 462.44
R14894 vdd.n1372 vdd.n1143 462.44
R14895 vdd.n293 vdd.t233 329.043
R14896 vdd.n238 vdd.t205 329.043
R14897 vdd.n195 vdd.t220 329.043
R14898 vdd.n140 vdd.t197 329.043
R14899 vdd.n98 vdd.t154 329.043
R14900 vdd.n43 vdd.t135 329.043
R14901 vdd.n1662 vdd.t246 329.043
R14902 vdd.n1717 vdd.t158 329.043
R14903 vdd.n1564 vdd.t234 329.043
R14904 vdd.n1619 vdd.t141 329.043
R14905 vdd.n1467 vdd.t137 329.043
R14906 vdd.n1522 vdd.t155 329.043
R14907 vdd.n1148 vdd.t38 319.788
R14908 vdd.n1304 vdd.t48 319.788
R14909 vdd.n1340 vdd.t55 319.788
R14910 vdd.n2250 vdd.t44 319.788
R14911 vdd.n1887 vdd.t57 319.788
R14912 vdd.n1847 vdd.t60 319.788
R14913 vdd.n405 vdd.t33 319.788
R14914 vdd.n419 vdd.t91 319.788
R14915 vdd.n431 vdd.t97 319.788
R14916 vdd.n723 vdd.t30 319.788
R14917 vdd.n686 vdd.t41 319.788
R14918 vdd.n3013 vdd.t95 319.788
R14919 vdd.n1149 vdd.t37 303.69
R14920 vdd.n1305 vdd.t47 303.69
R14921 vdd.n1341 vdd.t54 303.69
R14922 vdd.n2251 vdd.t45 303.69
R14923 vdd.n1888 vdd.t58 303.69
R14924 vdd.n1848 vdd.t61 303.69
R14925 vdd.n406 vdd.t34 303.69
R14926 vdd.n420 vdd.t92 303.69
R14927 vdd.n432 vdd.t98 303.69
R14928 vdd.n724 vdd.t29 303.69
R14929 vdd.n687 vdd.t40 303.69
R14930 vdd.n3014 vdd.t94 303.69
R14931 vdd.n2782 vdd.n884 297.074
R14932 vdd.n2975 vdd.n778 297.074
R14933 vdd.n2912 vdd.n775 297.074
R14934 vdd.n2705 vdd.n885 297.074
R14935 vdd.n2520 vdd.n925 297.074
R14936 vdd.n2451 vdd.n2450 297.074
R14937 vdd.n2197 vdd.n1021 297.074
R14938 vdd.n2293 vdd.n1019 297.074
R14939 vdd.n2891 vdd.n776 297.074
R14940 vdd.n2978 vdd.n2977 297.074
R14941 vdd.n2554 vdd.n886 297.074
R14942 vdd.n2780 vdd.n887 297.074
R14943 vdd.n2448 vdd.n934 297.074
R14944 vdd.n932 vdd.n907 297.074
R14945 vdd.n2134 vdd.n1022 297.074
R14946 vdd.n2291 vdd.n1023 297.074
R14947 vdd.n2893 vdd.n776 185
R14948 vdd.n2976 vdd.n776 185
R14949 vdd.n2895 vdd.n2894 185
R14950 vdd.n2894 vdd.n774 185
R14951 vdd.n2896 vdd.n810 185
R14952 vdd.n2906 vdd.n810 185
R14953 vdd.n2897 vdd.n819 185
R14954 vdd.n819 vdd.n817 185
R14955 vdd.n2899 vdd.n2898 185
R14956 vdd.n2900 vdd.n2899 185
R14957 vdd.n2852 vdd.n818 185
R14958 vdd.n818 vdd.n814 185
R14959 vdd.n2851 vdd.n2850 185
R14960 vdd.n2850 vdd.n2849 185
R14961 vdd.n821 vdd.n820 185
R14962 vdd.n822 vdd.n821 185
R14963 vdd.n2842 vdd.n2841 185
R14964 vdd.n2843 vdd.n2842 185
R14965 vdd.n2838 vdd.n831 185
R14966 vdd.n831 vdd.n828 185
R14967 vdd.n2837 vdd.n2836 185
R14968 vdd.n2836 vdd.n2835 185
R14969 vdd.n833 vdd.n832 185
R14970 vdd.n841 vdd.n833 185
R14971 vdd.n2828 vdd.n2827 185
R14972 vdd.n2829 vdd.n2828 185
R14973 vdd.n2826 vdd.n842 185
R14974 vdd.n2677 vdd.n842 185
R14975 vdd.n2825 vdd.n2824 185
R14976 vdd.n2824 vdd.n2823 185
R14977 vdd.n844 vdd.n843 185
R14978 vdd.n845 vdd.n844 185
R14979 vdd.n2816 vdd.n2815 185
R14980 vdd.n2817 vdd.n2816 185
R14981 vdd.n2814 vdd.n854 185
R14982 vdd.n854 vdd.n851 185
R14983 vdd.n2813 vdd.n2812 185
R14984 vdd.n2812 vdd.n2811 185
R14985 vdd.n856 vdd.n855 185
R14986 vdd.n864 vdd.n856 185
R14987 vdd.n2804 vdd.n2803 185
R14988 vdd.n2805 vdd.n2804 185
R14989 vdd.n2802 vdd.n865 185
R14990 vdd.n871 vdd.n865 185
R14991 vdd.n2801 vdd.n2800 185
R14992 vdd.n2800 vdd.n2799 185
R14993 vdd.n867 vdd.n866 185
R14994 vdd.n868 vdd.n867 185
R14995 vdd.n2792 vdd.n2791 185
R14996 vdd.n2793 vdd.n2792 185
R14997 vdd.n2790 vdd.n877 185
R14998 vdd.n2698 vdd.n877 185
R14999 vdd.n2789 vdd.n2788 185
R15000 vdd.n2788 vdd.n2787 185
R15001 vdd.n879 vdd.n878 185
R15002 vdd.t260 vdd.n879 185
R15003 vdd.n2780 vdd.n2779 185
R15004 vdd.n2781 vdd.n2780 185
R15005 vdd.n2778 vdd.n887 185
R15006 vdd.n2777 vdd.n2776 185
R15007 vdd.n889 vdd.n888 185
R15008 vdd.n2563 vdd.n2562 185
R15009 vdd.n2565 vdd.n2564 185
R15010 vdd.n2567 vdd.n2566 185
R15011 vdd.n2569 vdd.n2568 185
R15012 vdd.n2571 vdd.n2570 185
R15013 vdd.n2573 vdd.n2572 185
R15014 vdd.n2575 vdd.n2574 185
R15015 vdd.n2577 vdd.n2576 185
R15016 vdd.n2579 vdd.n2578 185
R15017 vdd.n2581 vdd.n2580 185
R15018 vdd.n2583 vdd.n2582 185
R15019 vdd.n2585 vdd.n2584 185
R15020 vdd.n2587 vdd.n2586 185
R15021 vdd.n2589 vdd.n2588 185
R15022 vdd.n2591 vdd.n2590 185
R15023 vdd.n2593 vdd.n2592 185
R15024 vdd.n2595 vdd.n2594 185
R15025 vdd.n2597 vdd.n2596 185
R15026 vdd.n2599 vdd.n2598 185
R15027 vdd.n2601 vdd.n2600 185
R15028 vdd.n2603 vdd.n2602 185
R15029 vdd.n2605 vdd.n2604 185
R15030 vdd.n2607 vdd.n2606 185
R15031 vdd.n2609 vdd.n2608 185
R15032 vdd.n2611 vdd.n2610 185
R15033 vdd.n2613 vdd.n2612 185
R15034 vdd.n2615 vdd.n2614 185
R15035 vdd.n2617 vdd.n2616 185
R15036 vdd.n2619 vdd.n2618 185
R15037 vdd.n2621 vdd.n2620 185
R15038 vdd.n2623 vdd.n2622 185
R15039 vdd.n2624 vdd.n2554 185
R15040 vdd.n2774 vdd.n2554 185
R15041 vdd.n2979 vdd.n2978 185
R15042 vdd.n2980 vdd.n767 185
R15043 vdd.n2982 vdd.n2981 185
R15044 vdd.n2984 vdd.n765 185
R15045 vdd.n2986 vdd.n2985 185
R15046 vdd.n2987 vdd.n764 185
R15047 vdd.n2989 vdd.n2988 185
R15048 vdd.n2991 vdd.n762 185
R15049 vdd.n2993 vdd.n2992 185
R15050 vdd.n2994 vdd.n761 185
R15051 vdd.n2996 vdd.n2995 185
R15052 vdd.n2998 vdd.n759 185
R15053 vdd.n3000 vdd.n2999 185
R15054 vdd.n3001 vdd.n758 185
R15055 vdd.n3003 vdd.n3002 185
R15056 vdd.n3005 vdd.n757 185
R15057 vdd.n3006 vdd.n754 185
R15058 vdd.n3009 vdd.n3008 185
R15059 vdd.n755 vdd.n753 185
R15060 vdd.n2865 vdd.n2864 185
R15061 vdd.n2867 vdd.n2866 185
R15062 vdd.n2869 vdd.n2861 185
R15063 vdd.n2871 vdd.n2870 185
R15064 vdd.n2872 vdd.n2860 185
R15065 vdd.n2874 vdd.n2873 185
R15066 vdd.n2876 vdd.n2858 185
R15067 vdd.n2878 vdd.n2877 185
R15068 vdd.n2879 vdd.n2857 185
R15069 vdd.n2881 vdd.n2880 185
R15070 vdd.n2883 vdd.n2855 185
R15071 vdd.n2885 vdd.n2884 185
R15072 vdd.n2886 vdd.n2854 185
R15073 vdd.n2888 vdd.n2887 185
R15074 vdd.n2890 vdd.n2853 185
R15075 vdd.n2892 vdd.n2891 185
R15076 vdd.n2891 vdd.n756 185
R15077 vdd.n2977 vdd.n771 185
R15078 vdd.n2977 vdd.n2976 185
R15079 vdd.n2629 vdd.n773 185
R15080 vdd.n774 vdd.n773 185
R15081 vdd.n2630 vdd.n809 185
R15082 vdd.n2906 vdd.n809 185
R15083 vdd.n2632 vdd.n2631 185
R15084 vdd.n2631 vdd.n817 185
R15085 vdd.n2633 vdd.n816 185
R15086 vdd.n2900 vdd.n816 185
R15087 vdd.n2635 vdd.n2634 185
R15088 vdd.n2634 vdd.n814 185
R15089 vdd.n2636 vdd.n824 185
R15090 vdd.n2849 vdd.n824 185
R15091 vdd.n2638 vdd.n2637 185
R15092 vdd.n2637 vdd.n822 185
R15093 vdd.n2639 vdd.n830 185
R15094 vdd.n2843 vdd.n830 185
R15095 vdd.n2641 vdd.n2640 185
R15096 vdd.n2640 vdd.n828 185
R15097 vdd.n2642 vdd.n835 185
R15098 vdd.n2835 vdd.n835 185
R15099 vdd.n2644 vdd.n2643 185
R15100 vdd.n2643 vdd.n841 185
R15101 vdd.n2645 vdd.n840 185
R15102 vdd.n2829 vdd.n840 185
R15103 vdd.n2679 vdd.n2678 185
R15104 vdd.n2678 vdd.n2677 185
R15105 vdd.n2680 vdd.n847 185
R15106 vdd.n2823 vdd.n847 185
R15107 vdd.n2682 vdd.n2681 185
R15108 vdd.n2681 vdd.n845 185
R15109 vdd.n2683 vdd.n853 185
R15110 vdd.n2817 vdd.n853 185
R15111 vdd.n2685 vdd.n2684 185
R15112 vdd.n2684 vdd.n851 185
R15113 vdd.n2686 vdd.n858 185
R15114 vdd.n2811 vdd.n858 185
R15115 vdd.n2688 vdd.n2687 185
R15116 vdd.n2687 vdd.n864 185
R15117 vdd.n2689 vdd.n863 185
R15118 vdd.n2805 vdd.n863 185
R15119 vdd.n2691 vdd.n2690 185
R15120 vdd.n2690 vdd.n871 185
R15121 vdd.n2692 vdd.n870 185
R15122 vdd.n2799 vdd.n870 185
R15123 vdd.n2694 vdd.n2693 185
R15124 vdd.n2693 vdd.n868 185
R15125 vdd.n2695 vdd.n876 185
R15126 vdd.n2793 vdd.n876 185
R15127 vdd.n2697 vdd.n2696 185
R15128 vdd.n2698 vdd.n2697 185
R15129 vdd.n2628 vdd.n881 185
R15130 vdd.n2787 vdd.n881 185
R15131 vdd.n2627 vdd.n2626 185
R15132 vdd.n2626 vdd.t260 185
R15133 vdd.n2625 vdd.n886 185
R15134 vdd.n2781 vdd.n886 185
R15135 vdd.n2245 vdd.n2244 185
R15136 vdd.n2246 vdd.n2245 185
R15137 vdd.n1048 vdd.n1046 185
R15138 vdd.n1046 vdd.n1044 185
R15139 vdd.n1814 vdd.n1813 185
R15140 vdd.n1813 vdd.n1812 185
R15141 vdd.n1051 vdd.n1050 185
R15142 vdd.n1052 vdd.n1051 185
R15143 vdd.n1801 vdd.n1800 185
R15144 vdd.n1802 vdd.n1801 185
R15145 vdd.n1060 vdd.n1059 185
R15146 vdd.n1793 vdd.n1059 185
R15147 vdd.n1796 vdd.n1795 185
R15148 vdd.n1795 vdd.n1794 185
R15149 vdd.n1063 vdd.n1062 185
R15150 vdd.n1069 vdd.n1063 185
R15151 vdd.n1784 vdd.n1783 185
R15152 vdd.n1785 vdd.n1784 185
R15153 vdd.n1071 vdd.n1070 185
R15154 vdd.n1776 vdd.n1070 185
R15155 vdd.n1779 vdd.n1778 185
R15156 vdd.n1778 vdd.n1777 185
R15157 vdd.n1074 vdd.n1073 185
R15158 vdd.n1075 vdd.n1074 185
R15159 vdd.n1767 vdd.n1766 185
R15160 vdd.n1768 vdd.n1767 185
R15161 vdd.n1083 vdd.n1082 185
R15162 vdd.n1082 vdd.n1081 185
R15163 vdd.n1762 vdd.n1761 185
R15164 vdd.n1761 vdd.n1760 185
R15165 vdd.n1086 vdd.n1085 185
R15166 vdd.n1092 vdd.n1086 185
R15167 vdd.n1751 vdd.n1750 185
R15168 vdd.n1752 vdd.n1751 185
R15169 vdd.n1094 vdd.n1093 185
R15170 vdd.n1448 vdd.n1093 185
R15171 vdd.n1451 vdd.n1450 185
R15172 vdd.n1450 vdd.n1449 185
R15173 vdd.n1097 vdd.n1096 185
R15174 vdd.n1104 vdd.n1097 185
R15175 vdd.n1439 vdd.n1438 185
R15176 vdd.n1440 vdd.n1439 185
R15177 vdd.n1106 vdd.n1105 185
R15178 vdd.n1105 vdd.n1103 185
R15179 vdd.n1434 vdd.n1433 185
R15180 vdd.n1433 vdd.n1432 185
R15181 vdd.n1109 vdd.n1108 185
R15182 vdd.n1110 vdd.n1109 185
R15183 vdd.n1423 vdd.n1422 185
R15184 vdd.n1424 vdd.n1423 185
R15185 vdd.n1117 vdd.n1116 185
R15186 vdd.n1415 vdd.n1116 185
R15187 vdd.n1418 vdd.n1417 185
R15188 vdd.n1417 vdd.n1416 185
R15189 vdd.n1120 vdd.n1119 185
R15190 vdd.n1126 vdd.n1120 185
R15191 vdd.n1406 vdd.n1405 185
R15192 vdd.n1407 vdd.n1406 185
R15193 vdd.n1128 vdd.n1127 185
R15194 vdd.n1398 vdd.n1127 185
R15195 vdd.n1401 vdd.n1400 185
R15196 vdd.n1400 vdd.n1399 185
R15197 vdd.n1131 vdd.n1130 185
R15198 vdd.n1132 vdd.n1131 185
R15199 vdd.n1389 vdd.n1388 185
R15200 vdd.n1390 vdd.n1389 185
R15201 vdd.n1140 vdd.n1139 185
R15202 vdd.n1139 vdd.n1138 185
R15203 vdd.n1384 vdd.n1383 185
R15204 vdd.n1383 vdd.n1382 185
R15205 vdd.n1143 vdd.n1142 185
R15206 vdd.n1144 vdd.n1143 185
R15207 vdd.n1372 vdd.n1371 185
R15208 vdd.n1370 vdd.n1183 185
R15209 vdd.n1185 vdd.n1182 185
R15210 vdd.n1374 vdd.n1182 185
R15211 vdd.n1366 vdd.n1187 185
R15212 vdd.n1365 vdd.n1188 185
R15213 vdd.n1364 vdd.n1189 185
R15214 vdd.n1192 vdd.n1190 185
R15215 vdd.n1360 vdd.n1193 185
R15216 vdd.n1359 vdd.n1194 185
R15217 vdd.n1358 vdd.n1195 185
R15218 vdd.n1198 vdd.n1196 185
R15219 vdd.n1354 vdd.n1199 185
R15220 vdd.n1353 vdd.n1200 185
R15221 vdd.n1352 vdd.n1201 185
R15222 vdd.n1204 vdd.n1202 185
R15223 vdd.n1348 vdd.n1205 185
R15224 vdd.n1347 vdd.n1206 185
R15225 vdd.n1346 vdd.n1207 185
R15226 vdd.n1338 vdd.n1208 185
R15227 vdd.n1342 vdd.n1339 185
R15228 vdd.n1337 vdd.n1210 185
R15229 vdd.n1336 vdd.n1211 185
R15230 vdd.n1214 vdd.n1212 185
R15231 vdd.n1332 vdd.n1215 185
R15232 vdd.n1331 vdd.n1216 185
R15233 vdd.n1330 vdd.n1217 185
R15234 vdd.n1220 vdd.n1218 185
R15235 vdd.n1326 vdd.n1221 185
R15236 vdd.n1325 vdd.n1222 185
R15237 vdd.n1324 vdd.n1223 185
R15238 vdd.n1226 vdd.n1224 185
R15239 vdd.n1320 vdd.n1227 185
R15240 vdd.n1319 vdd.n1228 185
R15241 vdd.n1318 vdd.n1229 185
R15242 vdd.n1232 vdd.n1230 185
R15243 vdd.n1314 vdd.n1233 185
R15244 vdd.n1313 vdd.n1234 185
R15245 vdd.n1312 vdd.n1235 185
R15246 vdd.n1238 vdd.n1236 185
R15247 vdd.n1308 vdd.n1239 185
R15248 vdd.n1307 vdd.n1240 185
R15249 vdd.n1306 vdd.n1303 185
R15250 vdd.n1243 vdd.n1241 185
R15251 vdd.n1299 vdd.n1244 185
R15252 vdd.n1298 vdd.n1245 185
R15253 vdd.n1297 vdd.n1246 185
R15254 vdd.n1249 vdd.n1247 185
R15255 vdd.n1293 vdd.n1250 185
R15256 vdd.n1292 vdd.n1251 185
R15257 vdd.n1291 vdd.n1252 185
R15258 vdd.n1255 vdd.n1253 185
R15259 vdd.n1287 vdd.n1256 185
R15260 vdd.n1286 vdd.n1257 185
R15261 vdd.n1285 vdd.n1258 185
R15262 vdd.n1261 vdd.n1259 185
R15263 vdd.n1281 vdd.n1262 185
R15264 vdd.n1280 vdd.n1263 185
R15265 vdd.n1279 vdd.n1264 185
R15266 vdd.n1267 vdd.n1265 185
R15267 vdd.n1275 vdd.n1268 185
R15268 vdd.n1274 vdd.n1269 185
R15269 vdd.n1273 vdd.n1270 185
R15270 vdd.n1271 vdd.n1151 185
R15271 vdd.n1376 vdd.n1375 185
R15272 vdd.n1375 vdd.n1374 185
R15273 vdd.n2249 vdd.n2248 185
R15274 vdd.n2253 vdd.n1040 185
R15275 vdd.n1916 vdd.n1039 185
R15276 vdd.n1919 vdd.n1918 185
R15277 vdd.n1921 vdd.n1920 185
R15278 vdd.n1924 vdd.n1923 185
R15279 vdd.n1926 vdd.n1925 185
R15280 vdd.n1928 vdd.n1914 185
R15281 vdd.n1930 vdd.n1929 185
R15282 vdd.n1931 vdd.n1908 185
R15283 vdd.n1933 vdd.n1932 185
R15284 vdd.n1935 vdd.n1906 185
R15285 vdd.n1937 vdd.n1936 185
R15286 vdd.n1938 vdd.n1901 185
R15287 vdd.n1940 vdd.n1939 185
R15288 vdd.n1942 vdd.n1899 185
R15289 vdd.n1944 vdd.n1943 185
R15290 vdd.n1945 vdd.n1895 185
R15291 vdd.n1947 vdd.n1946 185
R15292 vdd.n1949 vdd.n1892 185
R15293 vdd.n1951 vdd.n1950 185
R15294 vdd.n1893 vdd.n1886 185
R15295 vdd.n1955 vdd.n1890 185
R15296 vdd.n1956 vdd.n1882 185
R15297 vdd.n1958 vdd.n1957 185
R15298 vdd.n1960 vdd.n1880 185
R15299 vdd.n1962 vdd.n1961 185
R15300 vdd.n1963 vdd.n1875 185
R15301 vdd.n1965 vdd.n1964 185
R15302 vdd.n1967 vdd.n1873 185
R15303 vdd.n1969 vdd.n1968 185
R15304 vdd.n1970 vdd.n1868 185
R15305 vdd.n1972 vdd.n1971 185
R15306 vdd.n1974 vdd.n1866 185
R15307 vdd.n1976 vdd.n1975 185
R15308 vdd.n1977 vdd.n1861 185
R15309 vdd.n1979 vdd.n1978 185
R15310 vdd.n1981 vdd.n1859 185
R15311 vdd.n1983 vdd.n1982 185
R15312 vdd.n1984 vdd.n1855 185
R15313 vdd.n1986 vdd.n1985 185
R15314 vdd.n1988 vdd.n1852 185
R15315 vdd.n1990 vdd.n1989 185
R15316 vdd.n1853 vdd.n1846 185
R15317 vdd.n1994 vdd.n1850 185
R15318 vdd.n1995 vdd.n1842 185
R15319 vdd.n1997 vdd.n1996 185
R15320 vdd.n1999 vdd.n1840 185
R15321 vdd.n2001 vdd.n2000 185
R15322 vdd.n2002 vdd.n1835 185
R15323 vdd.n2004 vdd.n2003 185
R15324 vdd.n2006 vdd.n1833 185
R15325 vdd.n2008 vdd.n2007 185
R15326 vdd.n2009 vdd.n1828 185
R15327 vdd.n2011 vdd.n2010 185
R15328 vdd.n2013 vdd.n1827 185
R15329 vdd.n2014 vdd.n1824 185
R15330 vdd.n2017 vdd.n2016 185
R15331 vdd.n1826 vdd.n1822 185
R15332 vdd.n2234 vdd.n1820 185
R15333 vdd.n2236 vdd.n2235 185
R15334 vdd.n2238 vdd.n1818 185
R15335 vdd.n2240 vdd.n2239 185
R15336 vdd.n2241 vdd.n1047 185
R15337 vdd.n2247 vdd.n1043 185
R15338 vdd.n2247 vdd.n2246 185
R15339 vdd.n1055 vdd.n1042 185
R15340 vdd.n1044 vdd.n1042 185
R15341 vdd.n1811 vdd.n1810 185
R15342 vdd.n1812 vdd.n1811 185
R15343 vdd.n1054 vdd.n1053 185
R15344 vdd.n1053 vdd.n1052 185
R15345 vdd.n1804 vdd.n1803 185
R15346 vdd.n1803 vdd.n1802 185
R15347 vdd.n1058 vdd.n1057 185
R15348 vdd.n1793 vdd.n1058 185
R15349 vdd.n1792 vdd.n1791 185
R15350 vdd.n1794 vdd.n1792 185
R15351 vdd.n1065 vdd.n1064 185
R15352 vdd.n1069 vdd.n1064 185
R15353 vdd.n1787 vdd.n1786 185
R15354 vdd.n1786 vdd.n1785 185
R15355 vdd.n1068 vdd.n1067 185
R15356 vdd.n1776 vdd.n1068 185
R15357 vdd.n1775 vdd.n1774 185
R15358 vdd.n1777 vdd.n1775 185
R15359 vdd.n1077 vdd.n1076 185
R15360 vdd.n1076 vdd.n1075 185
R15361 vdd.n1770 vdd.n1769 185
R15362 vdd.n1769 vdd.n1768 185
R15363 vdd.n1080 vdd.n1079 185
R15364 vdd.n1081 vdd.n1080 185
R15365 vdd.n1759 vdd.n1758 185
R15366 vdd.n1760 vdd.n1759 185
R15367 vdd.n1088 vdd.n1087 185
R15368 vdd.n1092 vdd.n1087 185
R15369 vdd.n1754 vdd.n1753 185
R15370 vdd.n1753 vdd.n1752 185
R15371 vdd.n1091 vdd.n1090 185
R15372 vdd.n1448 vdd.n1091 185
R15373 vdd.n1447 vdd.n1446 185
R15374 vdd.n1449 vdd.n1447 185
R15375 vdd.n1099 vdd.n1098 185
R15376 vdd.n1104 vdd.n1098 185
R15377 vdd.n1442 vdd.n1441 185
R15378 vdd.n1441 vdd.n1440 185
R15379 vdd.n1102 vdd.n1101 185
R15380 vdd.n1103 vdd.n1102 185
R15381 vdd.n1431 vdd.n1430 185
R15382 vdd.n1432 vdd.n1431 185
R15383 vdd.n1112 vdd.n1111 185
R15384 vdd.n1111 vdd.n1110 185
R15385 vdd.n1426 vdd.n1425 185
R15386 vdd.n1425 vdd.n1424 185
R15387 vdd.n1115 vdd.n1114 185
R15388 vdd.n1415 vdd.n1115 185
R15389 vdd.n1414 vdd.n1413 185
R15390 vdd.n1416 vdd.n1414 185
R15391 vdd.n1122 vdd.n1121 185
R15392 vdd.n1126 vdd.n1121 185
R15393 vdd.n1409 vdd.n1408 185
R15394 vdd.n1408 vdd.n1407 185
R15395 vdd.n1125 vdd.n1124 185
R15396 vdd.n1398 vdd.n1125 185
R15397 vdd.n1397 vdd.n1396 185
R15398 vdd.n1399 vdd.n1397 185
R15399 vdd.n1134 vdd.n1133 185
R15400 vdd.n1133 vdd.n1132 185
R15401 vdd.n1392 vdd.n1391 185
R15402 vdd.n1391 vdd.n1390 185
R15403 vdd.n1137 vdd.n1136 185
R15404 vdd.n1138 vdd.n1137 185
R15405 vdd.n1381 vdd.n1380 185
R15406 vdd.n1382 vdd.n1381 185
R15407 vdd.n1146 vdd.n1145 185
R15408 vdd.n1145 vdd.n1144 185
R15409 vdd.n927 vdd.n925 185
R15410 vdd.n2449 vdd.n925 185
R15411 vdd.n2371 vdd.n944 185
R15412 vdd.n944 vdd.t256 185
R15413 vdd.n2373 vdd.n2372 185
R15414 vdd.n2374 vdd.n2373 185
R15415 vdd.n2370 vdd.n943 185
R15416 vdd.n2073 vdd.n943 185
R15417 vdd.n2369 vdd.n2368 185
R15418 vdd.n2368 vdd.n2367 185
R15419 vdd.n946 vdd.n945 185
R15420 vdd.n947 vdd.n946 185
R15421 vdd.n2358 vdd.n2357 185
R15422 vdd.n2359 vdd.n2358 185
R15423 vdd.n2356 vdd.n957 185
R15424 vdd.n957 vdd.n954 185
R15425 vdd.n2355 vdd.n2354 185
R15426 vdd.n2354 vdd.n2353 185
R15427 vdd.n959 vdd.n958 185
R15428 vdd.n960 vdd.n959 185
R15429 vdd.n2346 vdd.n2345 185
R15430 vdd.n2347 vdd.n2346 185
R15431 vdd.n2344 vdd.n968 185
R15432 vdd.n973 vdd.n968 185
R15433 vdd.n2343 vdd.n2342 185
R15434 vdd.n2342 vdd.n2341 185
R15435 vdd.n970 vdd.n969 185
R15436 vdd.n979 vdd.n970 185
R15437 vdd.n2334 vdd.n2333 185
R15438 vdd.n2335 vdd.n2334 185
R15439 vdd.n2332 vdd.n980 185
R15440 vdd.n2174 vdd.n980 185
R15441 vdd.n2331 vdd.n2330 185
R15442 vdd.n2330 vdd.n2329 185
R15443 vdd.n982 vdd.n981 185
R15444 vdd.n983 vdd.n982 185
R15445 vdd.n2322 vdd.n2321 185
R15446 vdd.n2323 vdd.n2322 185
R15447 vdd.n2320 vdd.n992 185
R15448 vdd.n992 vdd.n989 185
R15449 vdd.n2319 vdd.n2318 185
R15450 vdd.n2318 vdd.n2317 185
R15451 vdd.n994 vdd.n993 185
R15452 vdd.n1004 vdd.n994 185
R15453 vdd.n2309 vdd.n2308 185
R15454 vdd.n2310 vdd.n2309 185
R15455 vdd.n2307 vdd.n1005 185
R15456 vdd.n1005 vdd.n1001 185
R15457 vdd.n2306 vdd.n2305 185
R15458 vdd.n2305 vdd.n2304 185
R15459 vdd.n1007 vdd.n1006 185
R15460 vdd.n1008 vdd.n1007 185
R15461 vdd.n2297 vdd.n2296 185
R15462 vdd.n2298 vdd.n2297 185
R15463 vdd.n2295 vdd.n1017 185
R15464 vdd.n1017 vdd.n1014 185
R15465 vdd.n2294 vdd.n2293 185
R15466 vdd.n2293 vdd.n2292 185
R15467 vdd.n1019 vdd.n1018 185
R15468 vdd.n2029 vdd.n2028 185
R15469 vdd.n2030 vdd.n2026 185
R15470 vdd.n2026 vdd.n1020 185
R15471 vdd.n2032 vdd.n2031 185
R15472 vdd.n2034 vdd.n2025 185
R15473 vdd.n2037 vdd.n2036 185
R15474 vdd.n2038 vdd.n2024 185
R15475 vdd.n2040 vdd.n2039 185
R15476 vdd.n2042 vdd.n2023 185
R15477 vdd.n2045 vdd.n2044 185
R15478 vdd.n2046 vdd.n2022 185
R15479 vdd.n2048 vdd.n2047 185
R15480 vdd.n2050 vdd.n2021 185
R15481 vdd.n2053 vdd.n2052 185
R15482 vdd.n2054 vdd.n2020 185
R15483 vdd.n2056 vdd.n2055 185
R15484 vdd.n2058 vdd.n2019 185
R15485 vdd.n2231 vdd.n2059 185
R15486 vdd.n2230 vdd.n2229 185
R15487 vdd.n2227 vdd.n2060 185
R15488 vdd.n2225 vdd.n2224 185
R15489 vdd.n2223 vdd.n2061 185
R15490 vdd.n2222 vdd.n2221 185
R15491 vdd.n2219 vdd.n2062 185
R15492 vdd.n2217 vdd.n2216 185
R15493 vdd.n2215 vdd.n2063 185
R15494 vdd.n2214 vdd.n2213 185
R15495 vdd.n2211 vdd.n2064 185
R15496 vdd.n2209 vdd.n2208 185
R15497 vdd.n2207 vdd.n2065 185
R15498 vdd.n2206 vdd.n2205 185
R15499 vdd.n2203 vdd.n2066 185
R15500 vdd.n2201 vdd.n2200 185
R15501 vdd.n2199 vdd.n2067 185
R15502 vdd.n2198 vdd.n2197 185
R15503 vdd.n2452 vdd.n2451 185
R15504 vdd.n2454 vdd.n2453 185
R15505 vdd.n2456 vdd.n2455 185
R15506 vdd.n2459 vdd.n2458 185
R15507 vdd.n2461 vdd.n2460 185
R15508 vdd.n2463 vdd.n2462 185
R15509 vdd.n2465 vdd.n2464 185
R15510 vdd.n2467 vdd.n2466 185
R15511 vdd.n2469 vdd.n2468 185
R15512 vdd.n2471 vdd.n2470 185
R15513 vdd.n2473 vdd.n2472 185
R15514 vdd.n2475 vdd.n2474 185
R15515 vdd.n2477 vdd.n2476 185
R15516 vdd.n2479 vdd.n2478 185
R15517 vdd.n2481 vdd.n2480 185
R15518 vdd.n2483 vdd.n2482 185
R15519 vdd.n2485 vdd.n2484 185
R15520 vdd.n2487 vdd.n2486 185
R15521 vdd.n2489 vdd.n2488 185
R15522 vdd.n2491 vdd.n2490 185
R15523 vdd.n2493 vdd.n2492 185
R15524 vdd.n2495 vdd.n2494 185
R15525 vdd.n2497 vdd.n2496 185
R15526 vdd.n2499 vdd.n2498 185
R15527 vdd.n2501 vdd.n2500 185
R15528 vdd.n2503 vdd.n2502 185
R15529 vdd.n2505 vdd.n2504 185
R15530 vdd.n2507 vdd.n2506 185
R15531 vdd.n2509 vdd.n2508 185
R15532 vdd.n2511 vdd.n2510 185
R15533 vdd.n2513 vdd.n2512 185
R15534 vdd.n2515 vdd.n2514 185
R15535 vdd.n2517 vdd.n2516 185
R15536 vdd.n2518 vdd.n926 185
R15537 vdd.n2520 vdd.n2519 185
R15538 vdd.n2521 vdd.n2520 185
R15539 vdd.n2450 vdd.n930 185
R15540 vdd.n2450 vdd.n2449 185
R15541 vdd.n2071 vdd.n931 185
R15542 vdd.t256 vdd.n931 185
R15543 vdd.n2072 vdd.n941 185
R15544 vdd.n2374 vdd.n941 185
R15545 vdd.n2075 vdd.n2074 185
R15546 vdd.n2074 vdd.n2073 185
R15547 vdd.n2076 vdd.n948 185
R15548 vdd.n2367 vdd.n948 185
R15549 vdd.n2078 vdd.n2077 185
R15550 vdd.n2077 vdd.n947 185
R15551 vdd.n2079 vdd.n955 185
R15552 vdd.n2359 vdd.n955 185
R15553 vdd.n2081 vdd.n2080 185
R15554 vdd.n2080 vdd.n954 185
R15555 vdd.n2082 vdd.n961 185
R15556 vdd.n2353 vdd.n961 185
R15557 vdd.n2084 vdd.n2083 185
R15558 vdd.n2083 vdd.n960 185
R15559 vdd.n2085 vdd.n966 185
R15560 vdd.n2347 vdd.n966 185
R15561 vdd.n2087 vdd.n2086 185
R15562 vdd.n2086 vdd.n973 185
R15563 vdd.n2088 vdd.n971 185
R15564 vdd.n2341 vdd.n971 185
R15565 vdd.n2090 vdd.n2089 185
R15566 vdd.n2089 vdd.n979 185
R15567 vdd.n2091 vdd.n977 185
R15568 vdd.n2335 vdd.n977 185
R15569 vdd.n2176 vdd.n2175 185
R15570 vdd.n2175 vdd.n2174 185
R15571 vdd.n2177 vdd.n984 185
R15572 vdd.n2329 vdd.n984 185
R15573 vdd.n2179 vdd.n2178 185
R15574 vdd.n2178 vdd.n983 185
R15575 vdd.n2180 vdd.n990 185
R15576 vdd.n2323 vdd.n990 185
R15577 vdd.n2182 vdd.n2181 185
R15578 vdd.n2181 vdd.n989 185
R15579 vdd.n2183 vdd.n995 185
R15580 vdd.n2317 vdd.n995 185
R15581 vdd.n2185 vdd.n2184 185
R15582 vdd.n2184 vdd.n1004 185
R15583 vdd.n2186 vdd.n1002 185
R15584 vdd.n2310 vdd.n1002 185
R15585 vdd.n2188 vdd.n2187 185
R15586 vdd.n2187 vdd.n1001 185
R15587 vdd.n2189 vdd.n1009 185
R15588 vdd.n2304 vdd.n1009 185
R15589 vdd.n2191 vdd.n2190 185
R15590 vdd.n2190 vdd.n1008 185
R15591 vdd.n2192 vdd.n1015 185
R15592 vdd.n2298 vdd.n1015 185
R15593 vdd.n2194 vdd.n2193 185
R15594 vdd.n2193 vdd.n1014 185
R15595 vdd.n2195 vdd.n1021 185
R15596 vdd.n2292 vdd.n1021 185
R15597 vdd.n370 vdd.n369 185
R15598 vdd.n3254 vdd.n370 185
R15599 vdd.n3257 vdd.n3256 185
R15600 vdd.n3256 vdd.n3255 185
R15601 vdd.n3258 vdd.n364 185
R15602 vdd.n364 vdd.n363 185
R15603 vdd.n3260 vdd.n3259 185
R15604 vdd.n3261 vdd.n3260 185
R15605 vdd.n359 vdd.n358 185
R15606 vdd.n3262 vdd.n359 185
R15607 vdd.n3265 vdd.n3264 185
R15608 vdd.n3264 vdd.n3263 185
R15609 vdd.n3266 vdd.n353 185
R15610 vdd.n3236 vdd.n353 185
R15611 vdd.n3268 vdd.n3267 185
R15612 vdd.n3269 vdd.n3268 185
R15613 vdd.n348 vdd.n347 185
R15614 vdd.n3270 vdd.n348 185
R15615 vdd.n3273 vdd.n3272 185
R15616 vdd.n3272 vdd.n3271 185
R15617 vdd.n3274 vdd.n342 185
R15618 vdd.n349 vdd.n342 185
R15619 vdd.n3276 vdd.n3275 185
R15620 vdd.n3277 vdd.n3276 185
R15621 vdd.n338 vdd.n337 185
R15622 vdd.n3278 vdd.n338 185
R15623 vdd.n3281 vdd.n3280 185
R15624 vdd.n3280 vdd.n3279 185
R15625 vdd.n3282 vdd.n333 185
R15626 vdd.n333 vdd.n332 185
R15627 vdd.n3284 vdd.n3283 185
R15628 vdd.n3285 vdd.n3284 185
R15629 vdd.n327 vdd.n325 185
R15630 vdd.n3286 vdd.n327 185
R15631 vdd.n3289 vdd.n3288 185
R15632 vdd.n3288 vdd.n3287 185
R15633 vdd.n326 vdd.n324 185
R15634 vdd.n328 vdd.n326 185
R15635 vdd.n3212 vdd.n3211 185
R15636 vdd.n3213 vdd.n3212 185
R15637 vdd.n615 vdd.n614 185
R15638 vdd.n614 vdd.n613 185
R15639 vdd.n3207 vdd.n3206 185
R15640 vdd.n3206 vdd.n3205 185
R15641 vdd.n618 vdd.n617 185
R15642 vdd.n624 vdd.n618 185
R15643 vdd.n3193 vdd.n3192 185
R15644 vdd.n3194 vdd.n3193 185
R15645 vdd.n626 vdd.n625 185
R15646 vdd.n3185 vdd.n625 185
R15647 vdd.n3188 vdd.n3187 185
R15648 vdd.n3187 vdd.n3186 185
R15649 vdd.n629 vdd.n628 185
R15650 vdd.n636 vdd.n629 185
R15651 vdd.n3176 vdd.n3175 185
R15652 vdd.n3177 vdd.n3176 185
R15653 vdd.n638 vdd.n637 185
R15654 vdd.n637 vdd.n635 185
R15655 vdd.n3171 vdd.n3170 185
R15656 vdd.n3170 vdd.n3169 185
R15657 vdd.n641 vdd.n640 185
R15658 vdd.n642 vdd.n641 185
R15659 vdd.n3160 vdd.n3159 185
R15660 vdd.n3161 vdd.n3160 185
R15661 vdd.n650 vdd.n649 185
R15662 vdd.n649 vdd.n648 185
R15663 vdd.n3155 vdd.n3154 185
R15664 vdd.n3154 vdd.n3153 185
R15665 vdd.n653 vdd.n652 185
R15666 vdd.n659 vdd.n653 185
R15667 vdd.n3144 vdd.n3143 185
R15668 vdd.n3145 vdd.n3144 185
R15669 vdd.n3140 vdd.n660 185
R15670 vdd.n3139 vdd.n3138 185
R15671 vdd.n3136 vdd.n662 185
R15672 vdd.n3136 vdd.n658 185
R15673 vdd.n3135 vdd.n3134 185
R15674 vdd.n3133 vdd.n3132 185
R15675 vdd.n3131 vdd.n3130 185
R15676 vdd.n3129 vdd.n3128 185
R15677 vdd.n3127 vdd.n668 185
R15678 vdd.n3125 vdd.n3124 185
R15679 vdd.n3123 vdd.n669 185
R15680 vdd.n3122 vdd.n3121 185
R15681 vdd.n3119 vdd.n674 185
R15682 vdd.n3117 vdd.n3116 185
R15683 vdd.n3115 vdd.n675 185
R15684 vdd.n3114 vdd.n3113 185
R15685 vdd.n3111 vdd.n680 185
R15686 vdd.n3109 vdd.n3108 185
R15687 vdd.n3107 vdd.n681 185
R15688 vdd.n3106 vdd.n3105 185
R15689 vdd.n3103 vdd.n688 185
R15690 vdd.n3101 vdd.n3100 185
R15691 vdd.n3099 vdd.n689 185
R15692 vdd.n3098 vdd.n3097 185
R15693 vdd.n3095 vdd.n694 185
R15694 vdd.n3093 vdd.n3092 185
R15695 vdd.n3091 vdd.n695 185
R15696 vdd.n3090 vdd.n3089 185
R15697 vdd.n3087 vdd.n700 185
R15698 vdd.n3085 vdd.n3084 185
R15699 vdd.n3083 vdd.n701 185
R15700 vdd.n3082 vdd.n3081 185
R15701 vdd.n3079 vdd.n706 185
R15702 vdd.n3077 vdd.n3076 185
R15703 vdd.n3075 vdd.n707 185
R15704 vdd.n3074 vdd.n3073 185
R15705 vdd.n3071 vdd.n712 185
R15706 vdd.n3069 vdd.n3068 185
R15707 vdd.n3067 vdd.n713 185
R15708 vdd.n3066 vdd.n3065 185
R15709 vdd.n3063 vdd.n718 185
R15710 vdd.n3061 vdd.n3060 185
R15711 vdd.n3059 vdd.n719 185
R15712 vdd.n728 vdd.n722 185
R15713 vdd.n3055 vdd.n3054 185
R15714 vdd.n3052 vdd.n726 185
R15715 vdd.n3051 vdd.n3050 185
R15716 vdd.n3049 vdd.n3048 185
R15717 vdd.n3047 vdd.n732 185
R15718 vdd.n3045 vdd.n3044 185
R15719 vdd.n3043 vdd.n733 185
R15720 vdd.n3042 vdd.n3041 185
R15721 vdd.n3039 vdd.n738 185
R15722 vdd.n3037 vdd.n3036 185
R15723 vdd.n3035 vdd.n739 185
R15724 vdd.n3034 vdd.n3033 185
R15725 vdd.n3031 vdd.n744 185
R15726 vdd.n3029 vdd.n3028 185
R15727 vdd.n3027 vdd.n745 185
R15728 vdd.n3026 vdd.n3025 185
R15729 vdd.n3023 vdd.n3022 185
R15730 vdd.n3021 vdd.n3020 185
R15731 vdd.n3019 vdd.n3018 185
R15732 vdd.n3017 vdd.n3016 185
R15733 vdd.n3012 vdd.n657 185
R15734 vdd.n658 vdd.n657 185
R15735 vdd.n3251 vdd.n3250 185
R15736 vdd.n599 vdd.n404 185
R15737 vdd.n598 vdd.n597 185
R15738 vdd.n596 vdd.n595 185
R15739 vdd.n594 vdd.n409 185
R15740 vdd.n590 vdd.n589 185
R15741 vdd.n588 vdd.n587 185
R15742 vdd.n586 vdd.n585 185
R15743 vdd.n584 vdd.n411 185
R15744 vdd.n580 vdd.n579 185
R15745 vdd.n578 vdd.n577 185
R15746 vdd.n576 vdd.n575 185
R15747 vdd.n574 vdd.n413 185
R15748 vdd.n570 vdd.n569 185
R15749 vdd.n568 vdd.n567 185
R15750 vdd.n566 vdd.n565 185
R15751 vdd.n564 vdd.n415 185
R15752 vdd.n560 vdd.n559 185
R15753 vdd.n558 vdd.n557 185
R15754 vdd.n556 vdd.n555 185
R15755 vdd.n554 vdd.n417 185
R15756 vdd.n550 vdd.n549 185
R15757 vdd.n548 vdd.n547 185
R15758 vdd.n546 vdd.n545 185
R15759 vdd.n544 vdd.n421 185
R15760 vdd.n540 vdd.n539 185
R15761 vdd.n538 vdd.n537 185
R15762 vdd.n536 vdd.n535 185
R15763 vdd.n534 vdd.n423 185
R15764 vdd.n530 vdd.n529 185
R15765 vdd.n528 vdd.n527 185
R15766 vdd.n526 vdd.n525 185
R15767 vdd.n524 vdd.n425 185
R15768 vdd.n520 vdd.n519 185
R15769 vdd.n518 vdd.n517 185
R15770 vdd.n516 vdd.n515 185
R15771 vdd.n514 vdd.n427 185
R15772 vdd.n510 vdd.n509 185
R15773 vdd.n508 vdd.n507 185
R15774 vdd.n506 vdd.n505 185
R15775 vdd.n504 vdd.n429 185
R15776 vdd.n500 vdd.n499 185
R15777 vdd.n498 vdd.n497 185
R15778 vdd.n496 vdd.n495 185
R15779 vdd.n494 vdd.n433 185
R15780 vdd.n490 vdd.n489 185
R15781 vdd.n488 vdd.n487 185
R15782 vdd.n486 vdd.n485 185
R15783 vdd.n484 vdd.n435 185
R15784 vdd.n480 vdd.n479 185
R15785 vdd.n478 vdd.n477 185
R15786 vdd.n476 vdd.n475 185
R15787 vdd.n474 vdd.n437 185
R15788 vdd.n470 vdd.n469 185
R15789 vdd.n468 vdd.n467 185
R15790 vdd.n466 vdd.n465 185
R15791 vdd.n464 vdd.n439 185
R15792 vdd.n460 vdd.n459 185
R15793 vdd.n458 vdd.n457 185
R15794 vdd.n456 vdd.n455 185
R15795 vdd.n454 vdd.n441 185
R15796 vdd.n450 vdd.n449 185
R15797 vdd.n448 vdd.n447 185
R15798 vdd.n446 vdd.n445 185
R15799 vdd.n3247 vdd.n372 185
R15800 vdd.n3254 vdd.n372 185
R15801 vdd.n3246 vdd.n371 185
R15802 vdd.n3255 vdd.n371 185
R15803 vdd.n3245 vdd.n3244 185
R15804 vdd.n3244 vdd.n363 185
R15805 vdd.n602 vdd.n362 185
R15806 vdd.n3261 vdd.n362 185
R15807 vdd.n3240 vdd.n361 185
R15808 vdd.n3262 vdd.n361 185
R15809 vdd.n3239 vdd.n360 185
R15810 vdd.n3263 vdd.n360 185
R15811 vdd.n3238 vdd.n3237 185
R15812 vdd.n3237 vdd.n3236 185
R15813 vdd.n604 vdd.n352 185
R15814 vdd.n3269 vdd.n352 185
R15815 vdd.n3232 vdd.n351 185
R15816 vdd.n3270 vdd.n351 185
R15817 vdd.n3231 vdd.n350 185
R15818 vdd.n3271 vdd.n350 185
R15819 vdd.n3230 vdd.n3229 185
R15820 vdd.n3229 vdd.n349 185
R15821 vdd.n606 vdd.n341 185
R15822 vdd.n3277 vdd.n341 185
R15823 vdd.n3225 vdd.n340 185
R15824 vdd.n3278 vdd.n340 185
R15825 vdd.n3224 vdd.n339 185
R15826 vdd.n3279 vdd.n339 185
R15827 vdd.n3223 vdd.n3222 185
R15828 vdd.n3222 vdd.n332 185
R15829 vdd.n608 vdd.n331 185
R15830 vdd.n3285 vdd.n331 185
R15831 vdd.n3218 vdd.n330 185
R15832 vdd.n3286 vdd.n330 185
R15833 vdd.n3217 vdd.n329 185
R15834 vdd.n3287 vdd.n329 185
R15835 vdd.n3216 vdd.n3215 185
R15836 vdd.n3215 vdd.n328 185
R15837 vdd.n3214 vdd.n610 185
R15838 vdd.n3214 vdd.n3213 185
R15839 vdd.n3202 vdd.n612 185
R15840 vdd.n613 vdd.n612 185
R15841 vdd.n3204 vdd.n3203 185
R15842 vdd.n3205 vdd.n3204 185
R15843 vdd.n620 vdd.n619 185
R15844 vdd.n624 vdd.n619 185
R15845 vdd.n3196 vdd.n3195 185
R15846 vdd.n3195 vdd.n3194 185
R15847 vdd.n623 vdd.n622 185
R15848 vdd.n3185 vdd.n623 185
R15849 vdd.n3184 vdd.n3183 185
R15850 vdd.n3186 vdd.n3184 185
R15851 vdd.n631 vdd.n630 185
R15852 vdd.n636 vdd.n630 185
R15853 vdd.n3179 vdd.n3178 185
R15854 vdd.n3178 vdd.n3177 185
R15855 vdd.n634 vdd.n633 185
R15856 vdd.n635 vdd.n634 185
R15857 vdd.n3168 vdd.n3167 185
R15858 vdd.n3169 vdd.n3168 185
R15859 vdd.n644 vdd.n643 185
R15860 vdd.n643 vdd.n642 185
R15861 vdd.n3163 vdd.n3162 185
R15862 vdd.n3162 vdd.n3161 185
R15863 vdd.n647 vdd.n646 185
R15864 vdd.n648 vdd.n647 185
R15865 vdd.n3152 vdd.n3151 185
R15866 vdd.n3153 vdd.n3152 185
R15867 vdd.n655 vdd.n654 185
R15868 vdd.n659 vdd.n654 185
R15869 vdd.n3147 vdd.n3146 185
R15870 vdd.n3146 vdd.n3145 185
R15871 vdd.n884 vdd.n883 185
R15872 vdd.n2772 vdd.n2771 185
R15873 vdd.n2770 vdd.n2555 185
R15874 vdd.n2774 vdd.n2555 185
R15875 vdd.n2769 vdd.n2768 185
R15876 vdd.n2767 vdd.n2766 185
R15877 vdd.n2765 vdd.n2764 185
R15878 vdd.n2763 vdd.n2762 185
R15879 vdd.n2761 vdd.n2760 185
R15880 vdd.n2759 vdd.n2758 185
R15881 vdd.n2757 vdd.n2756 185
R15882 vdd.n2755 vdd.n2754 185
R15883 vdd.n2753 vdd.n2752 185
R15884 vdd.n2751 vdd.n2750 185
R15885 vdd.n2749 vdd.n2748 185
R15886 vdd.n2747 vdd.n2746 185
R15887 vdd.n2745 vdd.n2744 185
R15888 vdd.n2743 vdd.n2742 185
R15889 vdd.n2741 vdd.n2740 185
R15890 vdd.n2739 vdd.n2738 185
R15891 vdd.n2737 vdd.n2736 185
R15892 vdd.n2735 vdd.n2734 185
R15893 vdd.n2733 vdd.n2732 185
R15894 vdd.n2731 vdd.n2730 185
R15895 vdd.n2729 vdd.n2728 185
R15896 vdd.n2727 vdd.n2726 185
R15897 vdd.n2725 vdd.n2724 185
R15898 vdd.n2723 vdd.n2722 185
R15899 vdd.n2721 vdd.n2720 185
R15900 vdd.n2719 vdd.n2718 185
R15901 vdd.n2717 vdd.n2716 185
R15902 vdd.n2715 vdd.n2714 185
R15903 vdd.n2713 vdd.n2712 185
R15904 vdd.n2710 vdd.n2709 185
R15905 vdd.n2708 vdd.n2707 185
R15906 vdd.n2706 vdd.n2705 185
R15907 vdd.n2913 vdd.n2912 185
R15908 vdd.n2914 vdd.n803 185
R15909 vdd.n2916 vdd.n2915 185
R15910 vdd.n2918 vdd.n801 185
R15911 vdd.n2920 vdd.n2919 185
R15912 vdd.n2921 vdd.n800 185
R15913 vdd.n2923 vdd.n2922 185
R15914 vdd.n2925 vdd.n798 185
R15915 vdd.n2927 vdd.n2926 185
R15916 vdd.n2928 vdd.n797 185
R15917 vdd.n2930 vdd.n2929 185
R15918 vdd.n2932 vdd.n795 185
R15919 vdd.n2934 vdd.n2933 185
R15920 vdd.n2935 vdd.n794 185
R15921 vdd.n2937 vdd.n2936 185
R15922 vdd.n2939 vdd.n792 185
R15923 vdd.n2941 vdd.n2940 185
R15924 vdd.n2943 vdd.n791 185
R15925 vdd.n2945 vdd.n2944 185
R15926 vdd.n2947 vdd.n789 185
R15927 vdd.n2949 vdd.n2948 185
R15928 vdd.n2950 vdd.n788 185
R15929 vdd.n2952 vdd.n2951 185
R15930 vdd.n2954 vdd.n786 185
R15931 vdd.n2956 vdd.n2955 185
R15932 vdd.n2957 vdd.n785 185
R15933 vdd.n2959 vdd.n2958 185
R15934 vdd.n2961 vdd.n783 185
R15935 vdd.n2963 vdd.n2962 185
R15936 vdd.n2964 vdd.n782 185
R15937 vdd.n2966 vdd.n2965 185
R15938 vdd.n2968 vdd.n781 185
R15939 vdd.n2969 vdd.n780 185
R15940 vdd.n2972 vdd.n2971 185
R15941 vdd.n2973 vdd.n778 185
R15942 vdd.n778 vdd.n756 185
R15943 vdd.n2910 vdd.n775 185
R15944 vdd.n2976 vdd.n775 185
R15945 vdd.n2909 vdd.n2908 185
R15946 vdd.n2908 vdd.n774 185
R15947 vdd.n2907 vdd.n807 185
R15948 vdd.n2907 vdd.n2906 185
R15949 vdd.n2661 vdd.n808 185
R15950 vdd.n817 vdd.n808 185
R15951 vdd.n2662 vdd.n815 185
R15952 vdd.n2900 vdd.n815 185
R15953 vdd.n2664 vdd.n2663 185
R15954 vdd.n2663 vdd.n814 185
R15955 vdd.n2665 vdd.n823 185
R15956 vdd.n2849 vdd.n823 185
R15957 vdd.n2667 vdd.n2666 185
R15958 vdd.n2666 vdd.n822 185
R15959 vdd.n2668 vdd.n829 185
R15960 vdd.n2843 vdd.n829 185
R15961 vdd.n2670 vdd.n2669 185
R15962 vdd.n2669 vdd.n828 185
R15963 vdd.n2671 vdd.n834 185
R15964 vdd.n2835 vdd.n834 185
R15965 vdd.n2673 vdd.n2672 185
R15966 vdd.n2672 vdd.n841 185
R15967 vdd.n2674 vdd.n839 185
R15968 vdd.n2829 vdd.n839 185
R15969 vdd.n2676 vdd.n2675 185
R15970 vdd.n2677 vdd.n2676 185
R15971 vdd.n2660 vdd.n846 185
R15972 vdd.n2823 vdd.n846 185
R15973 vdd.n2659 vdd.n2658 185
R15974 vdd.n2658 vdd.n845 185
R15975 vdd.n2657 vdd.n852 185
R15976 vdd.n2817 vdd.n852 185
R15977 vdd.n2656 vdd.n2655 185
R15978 vdd.n2655 vdd.n851 185
R15979 vdd.n2654 vdd.n857 185
R15980 vdd.n2811 vdd.n857 185
R15981 vdd.n2653 vdd.n2652 185
R15982 vdd.n2652 vdd.n864 185
R15983 vdd.n2651 vdd.n862 185
R15984 vdd.n2805 vdd.n862 185
R15985 vdd.n2650 vdd.n2649 185
R15986 vdd.n2649 vdd.n871 185
R15987 vdd.n2648 vdd.n869 185
R15988 vdd.n2799 vdd.n869 185
R15989 vdd.n2647 vdd.n2646 185
R15990 vdd.n2646 vdd.n868 185
R15991 vdd.n2558 vdd.n875 185
R15992 vdd.n2793 vdd.n875 185
R15993 vdd.n2700 vdd.n2699 185
R15994 vdd.n2699 vdd.n2698 185
R15995 vdd.n2701 vdd.n880 185
R15996 vdd.n2787 vdd.n880 185
R15997 vdd.n2703 vdd.n2702 185
R15998 vdd.n2702 vdd.t260 185
R15999 vdd.n2704 vdd.n885 185
R16000 vdd.n2781 vdd.n885 185
R16001 vdd.n2783 vdd.n2782 185
R16002 vdd.n2782 vdd.n2781 185
R16003 vdd.n2784 vdd.n882 185
R16004 vdd.n882 vdd.t260 185
R16005 vdd.n2786 vdd.n2785 185
R16006 vdd.n2787 vdd.n2786 185
R16007 vdd.n874 vdd.n873 185
R16008 vdd.n2698 vdd.n874 185
R16009 vdd.n2795 vdd.n2794 185
R16010 vdd.n2794 vdd.n2793 185
R16011 vdd.n2796 vdd.n872 185
R16012 vdd.n872 vdd.n868 185
R16013 vdd.n2798 vdd.n2797 185
R16014 vdd.n2799 vdd.n2798 185
R16015 vdd.n861 vdd.n860 185
R16016 vdd.n871 vdd.n861 185
R16017 vdd.n2807 vdd.n2806 185
R16018 vdd.n2806 vdd.n2805 185
R16019 vdd.n2808 vdd.n859 185
R16020 vdd.n864 vdd.n859 185
R16021 vdd.n2810 vdd.n2809 185
R16022 vdd.n2811 vdd.n2810 185
R16023 vdd.n850 vdd.n849 185
R16024 vdd.n851 vdd.n850 185
R16025 vdd.n2819 vdd.n2818 185
R16026 vdd.n2818 vdd.n2817 185
R16027 vdd.n2820 vdd.n848 185
R16028 vdd.n848 vdd.n845 185
R16029 vdd.n2822 vdd.n2821 185
R16030 vdd.n2823 vdd.n2822 185
R16031 vdd.n838 vdd.n837 185
R16032 vdd.n2677 vdd.n838 185
R16033 vdd.n2831 vdd.n2830 185
R16034 vdd.n2830 vdd.n2829 185
R16035 vdd.n2832 vdd.n836 185
R16036 vdd.n841 vdd.n836 185
R16037 vdd.n2834 vdd.n2833 185
R16038 vdd.n2835 vdd.n2834 185
R16039 vdd.n827 vdd.n826 185
R16040 vdd.n828 vdd.n827 185
R16041 vdd.n2845 vdd.n2844 185
R16042 vdd.n2844 vdd.n2843 185
R16043 vdd.n2846 vdd.n825 185
R16044 vdd.n825 vdd.n822 185
R16045 vdd.n2848 vdd.n2847 185
R16046 vdd.n2849 vdd.n2848 185
R16047 vdd.n813 vdd.n812 185
R16048 vdd.n814 vdd.n813 185
R16049 vdd.n2902 vdd.n2901 185
R16050 vdd.n2901 vdd.n2900 185
R16051 vdd.n2903 vdd.n811 185
R16052 vdd.n817 vdd.n811 185
R16053 vdd.n2905 vdd.n2904 185
R16054 vdd.n2906 vdd.n2905 185
R16055 vdd.n779 vdd.n777 185
R16056 vdd.n777 vdd.n774 185
R16057 vdd.n2975 vdd.n2974 185
R16058 vdd.n2976 vdd.n2975 185
R16059 vdd.n2448 vdd.n2447 185
R16060 vdd.n2449 vdd.n2448 185
R16061 vdd.n935 vdd.n933 185
R16062 vdd.n933 vdd.t256 185
R16063 vdd.n2363 vdd.n942 185
R16064 vdd.n2374 vdd.n942 185
R16065 vdd.n2364 vdd.n951 185
R16066 vdd.n2073 vdd.n951 185
R16067 vdd.n2366 vdd.n2365 185
R16068 vdd.n2367 vdd.n2366 185
R16069 vdd.n2362 vdd.n950 185
R16070 vdd.n950 vdd.n947 185
R16071 vdd.n2361 vdd.n2360 185
R16072 vdd.n2360 vdd.n2359 185
R16073 vdd.n953 vdd.n952 185
R16074 vdd.n954 vdd.n953 185
R16075 vdd.n2352 vdd.n2351 185
R16076 vdd.n2353 vdd.n2352 185
R16077 vdd.n2350 vdd.n963 185
R16078 vdd.n963 vdd.n960 185
R16079 vdd.n2349 vdd.n2348 185
R16080 vdd.n2348 vdd.n2347 185
R16081 vdd.n965 vdd.n964 185
R16082 vdd.n973 vdd.n965 185
R16083 vdd.n2340 vdd.n2339 185
R16084 vdd.n2341 vdd.n2340 185
R16085 vdd.n2338 vdd.n974 185
R16086 vdd.n979 vdd.n974 185
R16087 vdd.n2337 vdd.n2336 185
R16088 vdd.n2336 vdd.n2335 185
R16089 vdd.n976 vdd.n975 185
R16090 vdd.n2174 vdd.n976 185
R16091 vdd.n2328 vdd.n2327 185
R16092 vdd.n2329 vdd.n2328 185
R16093 vdd.n2326 vdd.n986 185
R16094 vdd.n986 vdd.n983 185
R16095 vdd.n2325 vdd.n2324 185
R16096 vdd.n2324 vdd.n2323 185
R16097 vdd.n988 vdd.n987 185
R16098 vdd.n989 vdd.n988 185
R16099 vdd.n2316 vdd.n2315 185
R16100 vdd.n2317 vdd.n2316 185
R16101 vdd.n2313 vdd.n997 185
R16102 vdd.n1004 vdd.n997 185
R16103 vdd.n2312 vdd.n2311 185
R16104 vdd.n2311 vdd.n2310 185
R16105 vdd.n1000 vdd.n999 185
R16106 vdd.n1001 vdd.n1000 185
R16107 vdd.n2303 vdd.n2302 185
R16108 vdd.n2304 vdd.n2303 185
R16109 vdd.n2301 vdd.n1011 185
R16110 vdd.n1011 vdd.n1008 185
R16111 vdd.n2300 vdd.n2299 185
R16112 vdd.n2299 vdd.n2298 185
R16113 vdd.n1013 vdd.n1012 185
R16114 vdd.n1014 vdd.n1013 185
R16115 vdd.n2291 vdd.n2290 185
R16116 vdd.n2292 vdd.n2291 185
R16117 vdd.n2379 vdd.n907 185
R16118 vdd.n2521 vdd.n907 185
R16119 vdd.n2381 vdd.n2380 185
R16120 vdd.n2383 vdd.n2382 185
R16121 vdd.n2385 vdd.n2384 185
R16122 vdd.n2387 vdd.n2386 185
R16123 vdd.n2389 vdd.n2388 185
R16124 vdd.n2391 vdd.n2390 185
R16125 vdd.n2393 vdd.n2392 185
R16126 vdd.n2395 vdd.n2394 185
R16127 vdd.n2397 vdd.n2396 185
R16128 vdd.n2399 vdd.n2398 185
R16129 vdd.n2401 vdd.n2400 185
R16130 vdd.n2403 vdd.n2402 185
R16131 vdd.n2405 vdd.n2404 185
R16132 vdd.n2407 vdd.n2406 185
R16133 vdd.n2409 vdd.n2408 185
R16134 vdd.n2411 vdd.n2410 185
R16135 vdd.n2413 vdd.n2412 185
R16136 vdd.n2415 vdd.n2414 185
R16137 vdd.n2417 vdd.n2416 185
R16138 vdd.n2419 vdd.n2418 185
R16139 vdd.n2421 vdd.n2420 185
R16140 vdd.n2423 vdd.n2422 185
R16141 vdd.n2425 vdd.n2424 185
R16142 vdd.n2427 vdd.n2426 185
R16143 vdd.n2429 vdd.n2428 185
R16144 vdd.n2431 vdd.n2430 185
R16145 vdd.n2433 vdd.n2432 185
R16146 vdd.n2435 vdd.n2434 185
R16147 vdd.n2437 vdd.n2436 185
R16148 vdd.n2439 vdd.n2438 185
R16149 vdd.n2441 vdd.n2440 185
R16150 vdd.n2443 vdd.n2442 185
R16151 vdd.n2445 vdd.n2444 185
R16152 vdd.n2446 vdd.n934 185
R16153 vdd.n2378 vdd.n932 185
R16154 vdd.n2449 vdd.n932 185
R16155 vdd.n2377 vdd.n2376 185
R16156 vdd.n2376 vdd.t256 185
R16157 vdd.n2375 vdd.n939 185
R16158 vdd.n2375 vdd.n2374 185
R16159 vdd.n2155 vdd.n940 185
R16160 vdd.n2073 vdd.n940 185
R16161 vdd.n2156 vdd.n949 185
R16162 vdd.n2367 vdd.n949 185
R16163 vdd.n2158 vdd.n2157 185
R16164 vdd.n2157 vdd.n947 185
R16165 vdd.n2159 vdd.n956 185
R16166 vdd.n2359 vdd.n956 185
R16167 vdd.n2161 vdd.n2160 185
R16168 vdd.n2160 vdd.n954 185
R16169 vdd.n2162 vdd.n962 185
R16170 vdd.n2353 vdd.n962 185
R16171 vdd.n2164 vdd.n2163 185
R16172 vdd.n2163 vdd.n960 185
R16173 vdd.n2165 vdd.n967 185
R16174 vdd.n2347 vdd.n967 185
R16175 vdd.n2167 vdd.n2166 185
R16176 vdd.n2166 vdd.n973 185
R16177 vdd.n2168 vdd.n972 185
R16178 vdd.n2341 vdd.n972 185
R16179 vdd.n2170 vdd.n2169 185
R16180 vdd.n2169 vdd.n979 185
R16181 vdd.n2171 vdd.n978 185
R16182 vdd.n2335 vdd.n978 185
R16183 vdd.n2173 vdd.n2172 185
R16184 vdd.n2174 vdd.n2173 185
R16185 vdd.n2154 vdd.n985 185
R16186 vdd.n2329 vdd.n985 185
R16187 vdd.n2153 vdd.n2152 185
R16188 vdd.n2152 vdd.n983 185
R16189 vdd.n2151 vdd.n991 185
R16190 vdd.n2323 vdd.n991 185
R16191 vdd.n2150 vdd.n2149 185
R16192 vdd.n2149 vdd.n989 185
R16193 vdd.n2148 vdd.n996 185
R16194 vdd.n2317 vdd.n996 185
R16195 vdd.n2147 vdd.n2146 185
R16196 vdd.n2146 vdd.n1004 185
R16197 vdd.n2145 vdd.n1003 185
R16198 vdd.n2310 vdd.n1003 185
R16199 vdd.n2144 vdd.n2143 185
R16200 vdd.n2143 vdd.n1001 185
R16201 vdd.n2142 vdd.n1010 185
R16202 vdd.n2304 vdd.n1010 185
R16203 vdd.n2141 vdd.n2140 185
R16204 vdd.n2140 vdd.n1008 185
R16205 vdd.n2139 vdd.n1016 185
R16206 vdd.n2298 vdd.n1016 185
R16207 vdd.n2138 vdd.n2137 185
R16208 vdd.n2137 vdd.n1014 185
R16209 vdd.n2136 vdd.n1022 185
R16210 vdd.n2292 vdd.n1022 185
R16211 vdd.n2289 vdd.n1023 185
R16212 vdd.n2288 vdd.n2287 185
R16213 vdd.n2285 vdd.n1024 185
R16214 vdd.n2283 vdd.n2282 185
R16215 vdd.n2281 vdd.n1025 185
R16216 vdd.n2280 vdd.n2279 185
R16217 vdd.n2277 vdd.n1026 185
R16218 vdd.n2275 vdd.n2274 185
R16219 vdd.n2273 vdd.n1027 185
R16220 vdd.n2272 vdd.n2271 185
R16221 vdd.n2269 vdd.n1028 185
R16222 vdd.n2267 vdd.n2266 185
R16223 vdd.n2265 vdd.n1029 185
R16224 vdd.n2264 vdd.n2263 185
R16225 vdd.n2261 vdd.n1030 185
R16226 vdd.n2259 vdd.n2258 185
R16227 vdd.n2257 vdd.n1031 185
R16228 vdd.n2256 vdd.n1033 185
R16229 vdd.n2101 vdd.n1034 185
R16230 vdd.n2104 vdd.n2103 185
R16231 vdd.n2106 vdd.n2105 185
R16232 vdd.n2108 vdd.n2100 185
R16233 vdd.n2111 vdd.n2110 185
R16234 vdd.n2112 vdd.n2099 185
R16235 vdd.n2114 vdd.n2113 185
R16236 vdd.n2116 vdd.n2098 185
R16237 vdd.n2119 vdd.n2118 185
R16238 vdd.n2120 vdd.n2097 185
R16239 vdd.n2122 vdd.n2121 185
R16240 vdd.n2124 vdd.n2096 185
R16241 vdd.n2127 vdd.n2126 185
R16242 vdd.n2128 vdd.n2093 185
R16243 vdd.n2131 vdd.n2130 185
R16244 vdd.n2133 vdd.n2092 185
R16245 vdd.n2135 vdd.n2134 185
R16246 vdd.n2134 vdd.n1020 185
R16247 vdd.n315 vdd.n314 171.744
R16248 vdd.n314 vdd.n313 171.744
R16249 vdd.n313 vdd.n282 171.744
R16250 vdd.n306 vdd.n282 171.744
R16251 vdd.n306 vdd.n305 171.744
R16252 vdd.n305 vdd.n287 171.744
R16253 vdd.n298 vdd.n287 171.744
R16254 vdd.n298 vdd.n297 171.744
R16255 vdd.n297 vdd.n291 171.744
R16256 vdd.n260 vdd.n259 171.744
R16257 vdd.n259 vdd.n258 171.744
R16258 vdd.n258 vdd.n227 171.744
R16259 vdd.n251 vdd.n227 171.744
R16260 vdd.n251 vdd.n250 171.744
R16261 vdd.n250 vdd.n232 171.744
R16262 vdd.n243 vdd.n232 171.744
R16263 vdd.n243 vdd.n242 171.744
R16264 vdd.n242 vdd.n236 171.744
R16265 vdd.n217 vdd.n216 171.744
R16266 vdd.n216 vdd.n215 171.744
R16267 vdd.n215 vdd.n184 171.744
R16268 vdd.n208 vdd.n184 171.744
R16269 vdd.n208 vdd.n207 171.744
R16270 vdd.n207 vdd.n189 171.744
R16271 vdd.n200 vdd.n189 171.744
R16272 vdd.n200 vdd.n199 171.744
R16273 vdd.n199 vdd.n193 171.744
R16274 vdd.n162 vdd.n161 171.744
R16275 vdd.n161 vdd.n160 171.744
R16276 vdd.n160 vdd.n129 171.744
R16277 vdd.n153 vdd.n129 171.744
R16278 vdd.n153 vdd.n152 171.744
R16279 vdd.n152 vdd.n134 171.744
R16280 vdd.n145 vdd.n134 171.744
R16281 vdd.n145 vdd.n144 171.744
R16282 vdd.n144 vdd.n138 171.744
R16283 vdd.n120 vdd.n119 171.744
R16284 vdd.n119 vdd.n118 171.744
R16285 vdd.n118 vdd.n87 171.744
R16286 vdd.n111 vdd.n87 171.744
R16287 vdd.n111 vdd.n110 171.744
R16288 vdd.n110 vdd.n92 171.744
R16289 vdd.n103 vdd.n92 171.744
R16290 vdd.n103 vdd.n102 171.744
R16291 vdd.n102 vdd.n96 171.744
R16292 vdd.n65 vdd.n64 171.744
R16293 vdd.n64 vdd.n63 171.744
R16294 vdd.n63 vdd.n32 171.744
R16295 vdd.n56 vdd.n32 171.744
R16296 vdd.n56 vdd.n55 171.744
R16297 vdd.n55 vdd.n37 171.744
R16298 vdd.n48 vdd.n37 171.744
R16299 vdd.n48 vdd.n47 171.744
R16300 vdd.n47 vdd.n41 171.744
R16301 vdd.n1684 vdd.n1683 171.744
R16302 vdd.n1683 vdd.n1682 171.744
R16303 vdd.n1682 vdd.n1651 171.744
R16304 vdd.n1675 vdd.n1651 171.744
R16305 vdd.n1675 vdd.n1674 171.744
R16306 vdd.n1674 vdd.n1656 171.744
R16307 vdd.n1667 vdd.n1656 171.744
R16308 vdd.n1667 vdd.n1666 171.744
R16309 vdd.n1666 vdd.n1660 171.744
R16310 vdd.n1739 vdd.n1738 171.744
R16311 vdd.n1738 vdd.n1737 171.744
R16312 vdd.n1737 vdd.n1706 171.744
R16313 vdd.n1730 vdd.n1706 171.744
R16314 vdd.n1730 vdd.n1729 171.744
R16315 vdd.n1729 vdd.n1711 171.744
R16316 vdd.n1722 vdd.n1711 171.744
R16317 vdd.n1722 vdd.n1721 171.744
R16318 vdd.n1721 vdd.n1715 171.744
R16319 vdd.n1586 vdd.n1585 171.744
R16320 vdd.n1585 vdd.n1584 171.744
R16321 vdd.n1584 vdd.n1553 171.744
R16322 vdd.n1577 vdd.n1553 171.744
R16323 vdd.n1577 vdd.n1576 171.744
R16324 vdd.n1576 vdd.n1558 171.744
R16325 vdd.n1569 vdd.n1558 171.744
R16326 vdd.n1569 vdd.n1568 171.744
R16327 vdd.n1568 vdd.n1562 171.744
R16328 vdd.n1641 vdd.n1640 171.744
R16329 vdd.n1640 vdd.n1639 171.744
R16330 vdd.n1639 vdd.n1608 171.744
R16331 vdd.n1632 vdd.n1608 171.744
R16332 vdd.n1632 vdd.n1631 171.744
R16333 vdd.n1631 vdd.n1613 171.744
R16334 vdd.n1624 vdd.n1613 171.744
R16335 vdd.n1624 vdd.n1623 171.744
R16336 vdd.n1623 vdd.n1617 171.744
R16337 vdd.n1489 vdd.n1488 171.744
R16338 vdd.n1488 vdd.n1487 171.744
R16339 vdd.n1487 vdd.n1456 171.744
R16340 vdd.n1480 vdd.n1456 171.744
R16341 vdd.n1480 vdd.n1479 171.744
R16342 vdd.n1479 vdd.n1461 171.744
R16343 vdd.n1472 vdd.n1461 171.744
R16344 vdd.n1472 vdd.n1471 171.744
R16345 vdd.n1471 vdd.n1465 171.744
R16346 vdd.n1544 vdd.n1543 171.744
R16347 vdd.n1543 vdd.n1542 171.744
R16348 vdd.n1542 vdd.n1511 171.744
R16349 vdd.n1535 vdd.n1511 171.744
R16350 vdd.n1535 vdd.n1534 171.744
R16351 vdd.n1534 vdd.n1516 171.744
R16352 vdd.n1527 vdd.n1516 171.744
R16353 vdd.n1527 vdd.n1526 171.744
R16354 vdd.n1526 vdd.n1520 171.744
R16355 vdd.n449 vdd.n448 146.341
R16356 vdd.n455 vdd.n454 146.341
R16357 vdd.n459 vdd.n458 146.341
R16358 vdd.n465 vdd.n464 146.341
R16359 vdd.n469 vdd.n468 146.341
R16360 vdd.n475 vdd.n474 146.341
R16361 vdd.n479 vdd.n478 146.341
R16362 vdd.n485 vdd.n484 146.341
R16363 vdd.n489 vdd.n488 146.341
R16364 vdd.n495 vdd.n494 146.341
R16365 vdd.n499 vdd.n498 146.341
R16366 vdd.n505 vdd.n504 146.341
R16367 vdd.n509 vdd.n508 146.341
R16368 vdd.n515 vdd.n514 146.341
R16369 vdd.n519 vdd.n518 146.341
R16370 vdd.n525 vdd.n524 146.341
R16371 vdd.n529 vdd.n528 146.341
R16372 vdd.n535 vdd.n534 146.341
R16373 vdd.n539 vdd.n538 146.341
R16374 vdd.n545 vdd.n544 146.341
R16375 vdd.n549 vdd.n548 146.341
R16376 vdd.n555 vdd.n554 146.341
R16377 vdd.n559 vdd.n558 146.341
R16378 vdd.n565 vdd.n564 146.341
R16379 vdd.n569 vdd.n568 146.341
R16380 vdd.n575 vdd.n574 146.341
R16381 vdd.n579 vdd.n578 146.341
R16382 vdd.n585 vdd.n584 146.341
R16383 vdd.n589 vdd.n588 146.341
R16384 vdd.n595 vdd.n594 146.341
R16385 vdd.n597 vdd.n404 146.341
R16386 vdd.n3146 vdd.n654 146.341
R16387 vdd.n3152 vdd.n654 146.341
R16388 vdd.n3152 vdd.n647 146.341
R16389 vdd.n3162 vdd.n647 146.341
R16390 vdd.n3162 vdd.n643 146.341
R16391 vdd.n3168 vdd.n643 146.341
R16392 vdd.n3168 vdd.n634 146.341
R16393 vdd.n3178 vdd.n634 146.341
R16394 vdd.n3178 vdd.n630 146.341
R16395 vdd.n3184 vdd.n630 146.341
R16396 vdd.n3184 vdd.n623 146.341
R16397 vdd.n3195 vdd.n623 146.341
R16398 vdd.n3195 vdd.n619 146.341
R16399 vdd.n3204 vdd.n619 146.341
R16400 vdd.n3204 vdd.n612 146.341
R16401 vdd.n3214 vdd.n612 146.341
R16402 vdd.n3215 vdd.n3214 146.341
R16403 vdd.n3215 vdd.n329 146.341
R16404 vdd.n330 vdd.n329 146.341
R16405 vdd.n331 vdd.n330 146.341
R16406 vdd.n3222 vdd.n331 146.341
R16407 vdd.n3222 vdd.n339 146.341
R16408 vdd.n340 vdd.n339 146.341
R16409 vdd.n341 vdd.n340 146.341
R16410 vdd.n3229 vdd.n341 146.341
R16411 vdd.n3229 vdd.n350 146.341
R16412 vdd.n351 vdd.n350 146.341
R16413 vdd.n352 vdd.n351 146.341
R16414 vdd.n3237 vdd.n352 146.341
R16415 vdd.n3237 vdd.n360 146.341
R16416 vdd.n361 vdd.n360 146.341
R16417 vdd.n362 vdd.n361 146.341
R16418 vdd.n3244 vdd.n362 146.341
R16419 vdd.n3244 vdd.n371 146.341
R16420 vdd.n372 vdd.n371 146.341
R16421 vdd.n3138 vdd.n3136 146.341
R16422 vdd.n3136 vdd.n3135 146.341
R16423 vdd.n3132 vdd.n3131 146.341
R16424 vdd.n3128 vdd.n3127 146.341
R16425 vdd.n3125 vdd.n669 146.341
R16426 vdd.n3121 vdd.n3119 146.341
R16427 vdd.n3117 vdd.n675 146.341
R16428 vdd.n3113 vdd.n3111 146.341
R16429 vdd.n3109 vdd.n681 146.341
R16430 vdd.n3105 vdd.n3103 146.341
R16431 vdd.n3101 vdd.n689 146.341
R16432 vdd.n3097 vdd.n3095 146.341
R16433 vdd.n3093 vdd.n695 146.341
R16434 vdd.n3089 vdd.n3087 146.341
R16435 vdd.n3085 vdd.n701 146.341
R16436 vdd.n3081 vdd.n3079 146.341
R16437 vdd.n3077 vdd.n707 146.341
R16438 vdd.n3073 vdd.n3071 146.341
R16439 vdd.n3069 vdd.n713 146.341
R16440 vdd.n3065 vdd.n3063 146.341
R16441 vdd.n3061 vdd.n719 146.341
R16442 vdd.n3054 vdd.n728 146.341
R16443 vdd.n3052 vdd.n3051 146.341
R16444 vdd.n3048 vdd.n3047 146.341
R16445 vdd.n3045 vdd.n733 146.341
R16446 vdd.n3041 vdd.n3039 146.341
R16447 vdd.n3037 vdd.n739 146.341
R16448 vdd.n3033 vdd.n3031 146.341
R16449 vdd.n3029 vdd.n745 146.341
R16450 vdd.n3025 vdd.n3023 146.341
R16451 vdd.n3020 vdd.n3019 146.341
R16452 vdd.n3016 vdd.n657 146.341
R16453 vdd.n3144 vdd.n653 146.341
R16454 vdd.n3154 vdd.n653 146.341
R16455 vdd.n3154 vdd.n649 146.341
R16456 vdd.n3160 vdd.n649 146.341
R16457 vdd.n3160 vdd.n641 146.341
R16458 vdd.n3170 vdd.n641 146.341
R16459 vdd.n3170 vdd.n637 146.341
R16460 vdd.n3176 vdd.n637 146.341
R16461 vdd.n3176 vdd.n629 146.341
R16462 vdd.n3187 vdd.n629 146.341
R16463 vdd.n3187 vdd.n625 146.341
R16464 vdd.n3193 vdd.n625 146.341
R16465 vdd.n3193 vdd.n618 146.341
R16466 vdd.n3206 vdd.n618 146.341
R16467 vdd.n3206 vdd.n614 146.341
R16468 vdd.n3212 vdd.n614 146.341
R16469 vdd.n3212 vdd.n326 146.341
R16470 vdd.n3288 vdd.n326 146.341
R16471 vdd.n3288 vdd.n327 146.341
R16472 vdd.n3284 vdd.n327 146.341
R16473 vdd.n3284 vdd.n333 146.341
R16474 vdd.n3280 vdd.n333 146.341
R16475 vdd.n3280 vdd.n338 146.341
R16476 vdd.n3276 vdd.n338 146.341
R16477 vdd.n3276 vdd.n342 146.341
R16478 vdd.n3272 vdd.n342 146.341
R16479 vdd.n3272 vdd.n348 146.341
R16480 vdd.n3268 vdd.n348 146.341
R16481 vdd.n3268 vdd.n353 146.341
R16482 vdd.n3264 vdd.n353 146.341
R16483 vdd.n3264 vdd.n359 146.341
R16484 vdd.n3260 vdd.n359 146.341
R16485 vdd.n3260 vdd.n364 146.341
R16486 vdd.n3256 vdd.n364 146.341
R16487 vdd.n3256 vdd.n370 146.341
R16488 vdd.n2239 vdd.n2238 146.341
R16489 vdd.n2236 vdd.n1820 146.341
R16490 vdd.n2016 vdd.n1826 146.341
R16491 vdd.n2014 vdd.n2013 146.341
R16492 vdd.n2011 vdd.n1828 146.341
R16493 vdd.n2007 vdd.n2006 146.341
R16494 vdd.n2004 vdd.n1835 146.341
R16495 vdd.n2000 vdd.n1999 146.341
R16496 vdd.n1997 vdd.n1842 146.341
R16497 vdd.n1853 vdd.n1850 146.341
R16498 vdd.n1989 vdd.n1988 146.341
R16499 vdd.n1986 vdd.n1855 146.341
R16500 vdd.n1982 vdd.n1981 146.341
R16501 vdd.n1979 vdd.n1861 146.341
R16502 vdd.n1975 vdd.n1974 146.341
R16503 vdd.n1972 vdd.n1868 146.341
R16504 vdd.n1968 vdd.n1967 146.341
R16505 vdd.n1965 vdd.n1875 146.341
R16506 vdd.n1961 vdd.n1960 146.341
R16507 vdd.n1958 vdd.n1882 146.341
R16508 vdd.n1893 vdd.n1890 146.341
R16509 vdd.n1950 vdd.n1949 146.341
R16510 vdd.n1947 vdd.n1895 146.341
R16511 vdd.n1943 vdd.n1942 146.341
R16512 vdd.n1940 vdd.n1901 146.341
R16513 vdd.n1936 vdd.n1935 146.341
R16514 vdd.n1933 vdd.n1908 146.341
R16515 vdd.n1929 vdd.n1928 146.341
R16516 vdd.n1926 vdd.n1923 146.341
R16517 vdd.n1921 vdd.n1918 146.341
R16518 vdd.n1916 vdd.n1040 146.341
R16519 vdd.n1381 vdd.n1145 146.341
R16520 vdd.n1381 vdd.n1137 146.341
R16521 vdd.n1391 vdd.n1137 146.341
R16522 vdd.n1391 vdd.n1133 146.341
R16523 vdd.n1397 vdd.n1133 146.341
R16524 vdd.n1397 vdd.n1125 146.341
R16525 vdd.n1408 vdd.n1125 146.341
R16526 vdd.n1408 vdd.n1121 146.341
R16527 vdd.n1414 vdd.n1121 146.341
R16528 vdd.n1414 vdd.n1115 146.341
R16529 vdd.n1425 vdd.n1115 146.341
R16530 vdd.n1425 vdd.n1111 146.341
R16531 vdd.n1431 vdd.n1111 146.341
R16532 vdd.n1431 vdd.n1102 146.341
R16533 vdd.n1441 vdd.n1102 146.341
R16534 vdd.n1441 vdd.n1098 146.341
R16535 vdd.n1447 vdd.n1098 146.341
R16536 vdd.n1447 vdd.n1091 146.341
R16537 vdd.n1753 vdd.n1091 146.341
R16538 vdd.n1753 vdd.n1087 146.341
R16539 vdd.n1759 vdd.n1087 146.341
R16540 vdd.n1759 vdd.n1080 146.341
R16541 vdd.n1769 vdd.n1080 146.341
R16542 vdd.n1769 vdd.n1076 146.341
R16543 vdd.n1775 vdd.n1076 146.341
R16544 vdd.n1775 vdd.n1068 146.341
R16545 vdd.n1786 vdd.n1068 146.341
R16546 vdd.n1786 vdd.n1064 146.341
R16547 vdd.n1792 vdd.n1064 146.341
R16548 vdd.n1792 vdd.n1058 146.341
R16549 vdd.n1803 vdd.n1058 146.341
R16550 vdd.n1803 vdd.n1053 146.341
R16551 vdd.n1811 vdd.n1053 146.341
R16552 vdd.n1811 vdd.n1042 146.341
R16553 vdd.n2247 vdd.n1042 146.341
R16554 vdd.n1183 vdd.n1182 146.341
R16555 vdd.n1187 vdd.n1182 146.341
R16556 vdd.n1189 vdd.n1188 146.341
R16557 vdd.n1193 vdd.n1192 146.341
R16558 vdd.n1195 vdd.n1194 146.341
R16559 vdd.n1199 vdd.n1198 146.341
R16560 vdd.n1201 vdd.n1200 146.341
R16561 vdd.n1205 vdd.n1204 146.341
R16562 vdd.n1207 vdd.n1206 146.341
R16563 vdd.n1339 vdd.n1338 146.341
R16564 vdd.n1211 vdd.n1210 146.341
R16565 vdd.n1215 vdd.n1214 146.341
R16566 vdd.n1217 vdd.n1216 146.341
R16567 vdd.n1221 vdd.n1220 146.341
R16568 vdd.n1223 vdd.n1222 146.341
R16569 vdd.n1227 vdd.n1226 146.341
R16570 vdd.n1229 vdd.n1228 146.341
R16571 vdd.n1233 vdd.n1232 146.341
R16572 vdd.n1235 vdd.n1234 146.341
R16573 vdd.n1239 vdd.n1238 146.341
R16574 vdd.n1303 vdd.n1240 146.341
R16575 vdd.n1244 vdd.n1243 146.341
R16576 vdd.n1246 vdd.n1245 146.341
R16577 vdd.n1250 vdd.n1249 146.341
R16578 vdd.n1252 vdd.n1251 146.341
R16579 vdd.n1256 vdd.n1255 146.341
R16580 vdd.n1258 vdd.n1257 146.341
R16581 vdd.n1262 vdd.n1261 146.341
R16582 vdd.n1264 vdd.n1263 146.341
R16583 vdd.n1268 vdd.n1267 146.341
R16584 vdd.n1270 vdd.n1269 146.341
R16585 vdd.n1375 vdd.n1151 146.341
R16586 vdd.n1383 vdd.n1143 146.341
R16587 vdd.n1383 vdd.n1139 146.341
R16588 vdd.n1389 vdd.n1139 146.341
R16589 vdd.n1389 vdd.n1131 146.341
R16590 vdd.n1400 vdd.n1131 146.341
R16591 vdd.n1400 vdd.n1127 146.341
R16592 vdd.n1406 vdd.n1127 146.341
R16593 vdd.n1406 vdd.n1120 146.341
R16594 vdd.n1417 vdd.n1120 146.341
R16595 vdd.n1417 vdd.n1116 146.341
R16596 vdd.n1423 vdd.n1116 146.341
R16597 vdd.n1423 vdd.n1109 146.341
R16598 vdd.n1433 vdd.n1109 146.341
R16599 vdd.n1433 vdd.n1105 146.341
R16600 vdd.n1439 vdd.n1105 146.341
R16601 vdd.n1439 vdd.n1097 146.341
R16602 vdd.n1450 vdd.n1097 146.341
R16603 vdd.n1450 vdd.n1093 146.341
R16604 vdd.n1751 vdd.n1093 146.341
R16605 vdd.n1751 vdd.n1086 146.341
R16606 vdd.n1761 vdd.n1086 146.341
R16607 vdd.n1761 vdd.n1082 146.341
R16608 vdd.n1767 vdd.n1082 146.341
R16609 vdd.n1767 vdd.n1074 146.341
R16610 vdd.n1778 vdd.n1074 146.341
R16611 vdd.n1778 vdd.n1070 146.341
R16612 vdd.n1784 vdd.n1070 146.341
R16613 vdd.n1784 vdd.n1063 146.341
R16614 vdd.n1795 vdd.n1063 146.341
R16615 vdd.n1795 vdd.n1059 146.341
R16616 vdd.n1801 vdd.n1059 146.341
R16617 vdd.n1801 vdd.n1051 146.341
R16618 vdd.n1813 vdd.n1051 146.341
R16619 vdd.n1813 vdd.n1046 146.341
R16620 vdd.n2245 vdd.n1046 146.341
R16621 vdd.n1045 vdd.n1020 141.707
R16622 vdd.n756 vdd.n658 141.707
R16623 vdd.n2094 vdd.t79 127.284
R16624 vdd.n936 vdd.t64 127.284
R16625 vdd.n2068 vdd.t26 127.284
R16626 vdd.n928 vdd.t88 127.284
R16627 vdd.n2839 vdd.t51 127.284
R16628 vdd.n2839 vdd.t52 127.284
R16629 vdd.n2559 vdd.t86 127.284
R16630 vdd.n804 vdd.t68 127.284
R16631 vdd.n2556 vdd.t73 127.284
R16632 vdd.n768 vdd.t75 127.284
R16633 vdd.n998 vdd.t82 127.284
R16634 vdd.n998 vdd.t83 127.284
R16635 vdd.n22 vdd.n20 117.314
R16636 vdd.n17 vdd.n15 117.314
R16637 vdd.n27 vdd.n26 116.927
R16638 vdd.n24 vdd.n23 116.927
R16639 vdd.n22 vdd.n21 116.927
R16640 vdd.n17 vdd.n16 116.927
R16641 vdd.n19 vdd.n18 116.927
R16642 vdd.n27 vdd.n25 116.927
R16643 vdd.n2095 vdd.t78 111.188
R16644 vdd.n937 vdd.t65 111.188
R16645 vdd.n2069 vdd.t25 111.188
R16646 vdd.n929 vdd.t89 111.188
R16647 vdd.n2560 vdd.t85 111.188
R16648 vdd.n805 vdd.t69 111.188
R16649 vdd.n2557 vdd.t72 111.188
R16650 vdd.n769 vdd.t76 111.188
R16651 vdd.n2782 vdd.n882 99.5127
R16652 vdd.n2786 vdd.n882 99.5127
R16653 vdd.n2786 vdd.n874 99.5127
R16654 vdd.n2794 vdd.n874 99.5127
R16655 vdd.n2794 vdd.n872 99.5127
R16656 vdd.n2798 vdd.n872 99.5127
R16657 vdd.n2798 vdd.n861 99.5127
R16658 vdd.n2806 vdd.n861 99.5127
R16659 vdd.n2806 vdd.n859 99.5127
R16660 vdd.n2810 vdd.n859 99.5127
R16661 vdd.n2810 vdd.n850 99.5127
R16662 vdd.n2818 vdd.n850 99.5127
R16663 vdd.n2818 vdd.n848 99.5127
R16664 vdd.n2822 vdd.n848 99.5127
R16665 vdd.n2822 vdd.n838 99.5127
R16666 vdd.n2830 vdd.n838 99.5127
R16667 vdd.n2830 vdd.n836 99.5127
R16668 vdd.n2834 vdd.n836 99.5127
R16669 vdd.n2834 vdd.n827 99.5127
R16670 vdd.n2844 vdd.n827 99.5127
R16671 vdd.n2844 vdd.n825 99.5127
R16672 vdd.n2848 vdd.n825 99.5127
R16673 vdd.n2848 vdd.n813 99.5127
R16674 vdd.n2901 vdd.n813 99.5127
R16675 vdd.n2901 vdd.n811 99.5127
R16676 vdd.n2905 vdd.n811 99.5127
R16677 vdd.n2905 vdd.n777 99.5127
R16678 vdd.n2975 vdd.n777 99.5127
R16679 vdd.n2971 vdd.n778 99.5127
R16680 vdd.n2969 vdd.n2968 99.5127
R16681 vdd.n2966 vdd.n782 99.5127
R16682 vdd.n2962 vdd.n2961 99.5127
R16683 vdd.n2959 vdd.n785 99.5127
R16684 vdd.n2955 vdd.n2954 99.5127
R16685 vdd.n2952 vdd.n788 99.5127
R16686 vdd.n2948 vdd.n2947 99.5127
R16687 vdd.n2945 vdd.n791 99.5127
R16688 vdd.n2940 vdd.n2939 99.5127
R16689 vdd.n2937 vdd.n794 99.5127
R16690 vdd.n2933 vdd.n2932 99.5127
R16691 vdd.n2930 vdd.n797 99.5127
R16692 vdd.n2926 vdd.n2925 99.5127
R16693 vdd.n2923 vdd.n800 99.5127
R16694 vdd.n2919 vdd.n2918 99.5127
R16695 vdd.n2916 vdd.n803 99.5127
R16696 vdd.n2702 vdd.n885 99.5127
R16697 vdd.n2702 vdd.n880 99.5127
R16698 vdd.n2699 vdd.n880 99.5127
R16699 vdd.n2699 vdd.n875 99.5127
R16700 vdd.n2646 vdd.n875 99.5127
R16701 vdd.n2646 vdd.n869 99.5127
R16702 vdd.n2649 vdd.n869 99.5127
R16703 vdd.n2649 vdd.n862 99.5127
R16704 vdd.n2652 vdd.n862 99.5127
R16705 vdd.n2652 vdd.n857 99.5127
R16706 vdd.n2655 vdd.n857 99.5127
R16707 vdd.n2655 vdd.n852 99.5127
R16708 vdd.n2658 vdd.n852 99.5127
R16709 vdd.n2658 vdd.n846 99.5127
R16710 vdd.n2676 vdd.n846 99.5127
R16711 vdd.n2676 vdd.n839 99.5127
R16712 vdd.n2672 vdd.n839 99.5127
R16713 vdd.n2672 vdd.n834 99.5127
R16714 vdd.n2669 vdd.n834 99.5127
R16715 vdd.n2669 vdd.n829 99.5127
R16716 vdd.n2666 vdd.n829 99.5127
R16717 vdd.n2666 vdd.n823 99.5127
R16718 vdd.n2663 vdd.n823 99.5127
R16719 vdd.n2663 vdd.n815 99.5127
R16720 vdd.n815 vdd.n808 99.5127
R16721 vdd.n2907 vdd.n808 99.5127
R16722 vdd.n2908 vdd.n2907 99.5127
R16723 vdd.n2908 vdd.n775 99.5127
R16724 vdd.n2772 vdd.n2555 99.5127
R16725 vdd.n2768 vdd.n2555 99.5127
R16726 vdd.n2766 vdd.n2765 99.5127
R16727 vdd.n2762 vdd.n2761 99.5127
R16728 vdd.n2758 vdd.n2757 99.5127
R16729 vdd.n2754 vdd.n2753 99.5127
R16730 vdd.n2750 vdd.n2749 99.5127
R16731 vdd.n2746 vdd.n2745 99.5127
R16732 vdd.n2742 vdd.n2741 99.5127
R16733 vdd.n2738 vdd.n2737 99.5127
R16734 vdd.n2734 vdd.n2733 99.5127
R16735 vdd.n2730 vdd.n2729 99.5127
R16736 vdd.n2726 vdd.n2725 99.5127
R16737 vdd.n2722 vdd.n2721 99.5127
R16738 vdd.n2718 vdd.n2717 99.5127
R16739 vdd.n2714 vdd.n2713 99.5127
R16740 vdd.n2709 vdd.n2708 99.5127
R16741 vdd.n2520 vdd.n926 99.5127
R16742 vdd.n2516 vdd.n2515 99.5127
R16743 vdd.n2512 vdd.n2511 99.5127
R16744 vdd.n2508 vdd.n2507 99.5127
R16745 vdd.n2504 vdd.n2503 99.5127
R16746 vdd.n2500 vdd.n2499 99.5127
R16747 vdd.n2496 vdd.n2495 99.5127
R16748 vdd.n2492 vdd.n2491 99.5127
R16749 vdd.n2488 vdd.n2487 99.5127
R16750 vdd.n2484 vdd.n2483 99.5127
R16751 vdd.n2480 vdd.n2479 99.5127
R16752 vdd.n2476 vdd.n2475 99.5127
R16753 vdd.n2472 vdd.n2471 99.5127
R16754 vdd.n2468 vdd.n2467 99.5127
R16755 vdd.n2464 vdd.n2463 99.5127
R16756 vdd.n2460 vdd.n2459 99.5127
R16757 vdd.n2455 vdd.n2454 99.5127
R16758 vdd.n2193 vdd.n1021 99.5127
R16759 vdd.n2193 vdd.n1015 99.5127
R16760 vdd.n2190 vdd.n1015 99.5127
R16761 vdd.n2190 vdd.n1009 99.5127
R16762 vdd.n2187 vdd.n1009 99.5127
R16763 vdd.n2187 vdd.n1002 99.5127
R16764 vdd.n2184 vdd.n1002 99.5127
R16765 vdd.n2184 vdd.n995 99.5127
R16766 vdd.n2181 vdd.n995 99.5127
R16767 vdd.n2181 vdd.n990 99.5127
R16768 vdd.n2178 vdd.n990 99.5127
R16769 vdd.n2178 vdd.n984 99.5127
R16770 vdd.n2175 vdd.n984 99.5127
R16771 vdd.n2175 vdd.n977 99.5127
R16772 vdd.n2089 vdd.n977 99.5127
R16773 vdd.n2089 vdd.n971 99.5127
R16774 vdd.n2086 vdd.n971 99.5127
R16775 vdd.n2086 vdd.n966 99.5127
R16776 vdd.n2083 vdd.n966 99.5127
R16777 vdd.n2083 vdd.n961 99.5127
R16778 vdd.n2080 vdd.n961 99.5127
R16779 vdd.n2080 vdd.n955 99.5127
R16780 vdd.n2077 vdd.n955 99.5127
R16781 vdd.n2077 vdd.n948 99.5127
R16782 vdd.n2074 vdd.n948 99.5127
R16783 vdd.n2074 vdd.n941 99.5127
R16784 vdd.n941 vdd.n931 99.5127
R16785 vdd.n2450 vdd.n931 99.5127
R16786 vdd.n2028 vdd.n2026 99.5127
R16787 vdd.n2032 vdd.n2026 99.5127
R16788 vdd.n2036 vdd.n2034 99.5127
R16789 vdd.n2040 vdd.n2024 99.5127
R16790 vdd.n2044 vdd.n2042 99.5127
R16791 vdd.n2048 vdd.n2022 99.5127
R16792 vdd.n2052 vdd.n2050 99.5127
R16793 vdd.n2056 vdd.n2020 99.5127
R16794 vdd.n2059 vdd.n2058 99.5127
R16795 vdd.n2229 vdd.n2227 99.5127
R16796 vdd.n2225 vdd.n2061 99.5127
R16797 vdd.n2221 vdd.n2219 99.5127
R16798 vdd.n2217 vdd.n2063 99.5127
R16799 vdd.n2213 vdd.n2211 99.5127
R16800 vdd.n2209 vdd.n2065 99.5127
R16801 vdd.n2205 vdd.n2203 99.5127
R16802 vdd.n2201 vdd.n2067 99.5127
R16803 vdd.n2293 vdd.n1017 99.5127
R16804 vdd.n2297 vdd.n1017 99.5127
R16805 vdd.n2297 vdd.n1007 99.5127
R16806 vdd.n2305 vdd.n1007 99.5127
R16807 vdd.n2305 vdd.n1005 99.5127
R16808 vdd.n2309 vdd.n1005 99.5127
R16809 vdd.n2309 vdd.n994 99.5127
R16810 vdd.n2318 vdd.n994 99.5127
R16811 vdd.n2318 vdd.n992 99.5127
R16812 vdd.n2322 vdd.n992 99.5127
R16813 vdd.n2322 vdd.n982 99.5127
R16814 vdd.n2330 vdd.n982 99.5127
R16815 vdd.n2330 vdd.n980 99.5127
R16816 vdd.n2334 vdd.n980 99.5127
R16817 vdd.n2334 vdd.n970 99.5127
R16818 vdd.n2342 vdd.n970 99.5127
R16819 vdd.n2342 vdd.n968 99.5127
R16820 vdd.n2346 vdd.n968 99.5127
R16821 vdd.n2346 vdd.n959 99.5127
R16822 vdd.n2354 vdd.n959 99.5127
R16823 vdd.n2354 vdd.n957 99.5127
R16824 vdd.n2358 vdd.n957 99.5127
R16825 vdd.n2358 vdd.n946 99.5127
R16826 vdd.n2368 vdd.n946 99.5127
R16827 vdd.n2368 vdd.n943 99.5127
R16828 vdd.n2373 vdd.n943 99.5127
R16829 vdd.n2373 vdd.n944 99.5127
R16830 vdd.n944 vdd.n925 99.5127
R16831 vdd.n2891 vdd.n2890 99.5127
R16832 vdd.n2888 vdd.n2854 99.5127
R16833 vdd.n2884 vdd.n2883 99.5127
R16834 vdd.n2881 vdd.n2857 99.5127
R16835 vdd.n2877 vdd.n2876 99.5127
R16836 vdd.n2874 vdd.n2860 99.5127
R16837 vdd.n2870 vdd.n2869 99.5127
R16838 vdd.n2867 vdd.n2864 99.5127
R16839 vdd.n3008 vdd.n755 99.5127
R16840 vdd.n3006 vdd.n3005 99.5127
R16841 vdd.n3003 vdd.n758 99.5127
R16842 vdd.n2999 vdd.n2998 99.5127
R16843 vdd.n2996 vdd.n761 99.5127
R16844 vdd.n2992 vdd.n2991 99.5127
R16845 vdd.n2989 vdd.n764 99.5127
R16846 vdd.n2985 vdd.n2984 99.5127
R16847 vdd.n2982 vdd.n767 99.5127
R16848 vdd.n2626 vdd.n886 99.5127
R16849 vdd.n2626 vdd.n881 99.5127
R16850 vdd.n2697 vdd.n881 99.5127
R16851 vdd.n2697 vdd.n876 99.5127
R16852 vdd.n2693 vdd.n876 99.5127
R16853 vdd.n2693 vdd.n870 99.5127
R16854 vdd.n2690 vdd.n870 99.5127
R16855 vdd.n2690 vdd.n863 99.5127
R16856 vdd.n2687 vdd.n863 99.5127
R16857 vdd.n2687 vdd.n858 99.5127
R16858 vdd.n2684 vdd.n858 99.5127
R16859 vdd.n2684 vdd.n853 99.5127
R16860 vdd.n2681 vdd.n853 99.5127
R16861 vdd.n2681 vdd.n847 99.5127
R16862 vdd.n2678 vdd.n847 99.5127
R16863 vdd.n2678 vdd.n840 99.5127
R16864 vdd.n2643 vdd.n840 99.5127
R16865 vdd.n2643 vdd.n835 99.5127
R16866 vdd.n2640 vdd.n835 99.5127
R16867 vdd.n2640 vdd.n830 99.5127
R16868 vdd.n2637 vdd.n830 99.5127
R16869 vdd.n2637 vdd.n824 99.5127
R16870 vdd.n2634 vdd.n824 99.5127
R16871 vdd.n2634 vdd.n816 99.5127
R16872 vdd.n2631 vdd.n816 99.5127
R16873 vdd.n2631 vdd.n809 99.5127
R16874 vdd.n809 vdd.n773 99.5127
R16875 vdd.n2977 vdd.n773 99.5127
R16876 vdd.n2776 vdd.n889 99.5127
R16877 vdd.n2564 vdd.n2563 99.5127
R16878 vdd.n2568 vdd.n2567 99.5127
R16879 vdd.n2572 vdd.n2571 99.5127
R16880 vdd.n2576 vdd.n2575 99.5127
R16881 vdd.n2580 vdd.n2579 99.5127
R16882 vdd.n2584 vdd.n2583 99.5127
R16883 vdd.n2588 vdd.n2587 99.5127
R16884 vdd.n2592 vdd.n2591 99.5127
R16885 vdd.n2596 vdd.n2595 99.5127
R16886 vdd.n2600 vdd.n2599 99.5127
R16887 vdd.n2604 vdd.n2603 99.5127
R16888 vdd.n2608 vdd.n2607 99.5127
R16889 vdd.n2612 vdd.n2611 99.5127
R16890 vdd.n2616 vdd.n2615 99.5127
R16891 vdd.n2620 vdd.n2619 99.5127
R16892 vdd.n2622 vdd.n2554 99.5127
R16893 vdd.n2780 vdd.n879 99.5127
R16894 vdd.n2788 vdd.n879 99.5127
R16895 vdd.n2788 vdd.n877 99.5127
R16896 vdd.n2792 vdd.n877 99.5127
R16897 vdd.n2792 vdd.n867 99.5127
R16898 vdd.n2800 vdd.n867 99.5127
R16899 vdd.n2800 vdd.n865 99.5127
R16900 vdd.n2804 vdd.n865 99.5127
R16901 vdd.n2804 vdd.n856 99.5127
R16902 vdd.n2812 vdd.n856 99.5127
R16903 vdd.n2812 vdd.n854 99.5127
R16904 vdd.n2816 vdd.n854 99.5127
R16905 vdd.n2816 vdd.n844 99.5127
R16906 vdd.n2824 vdd.n844 99.5127
R16907 vdd.n2824 vdd.n842 99.5127
R16908 vdd.n2828 vdd.n842 99.5127
R16909 vdd.n2828 vdd.n833 99.5127
R16910 vdd.n2836 vdd.n833 99.5127
R16911 vdd.n2836 vdd.n831 99.5127
R16912 vdd.n2842 vdd.n831 99.5127
R16913 vdd.n2842 vdd.n821 99.5127
R16914 vdd.n2850 vdd.n821 99.5127
R16915 vdd.n2850 vdd.n818 99.5127
R16916 vdd.n2899 vdd.n818 99.5127
R16917 vdd.n2899 vdd.n819 99.5127
R16918 vdd.n819 vdd.n810 99.5127
R16919 vdd.n2894 vdd.n810 99.5127
R16920 vdd.n2894 vdd.n776 99.5127
R16921 vdd.n2444 vdd.n2443 99.5127
R16922 vdd.n2440 vdd.n2439 99.5127
R16923 vdd.n2436 vdd.n2435 99.5127
R16924 vdd.n2432 vdd.n2431 99.5127
R16925 vdd.n2428 vdd.n2427 99.5127
R16926 vdd.n2424 vdd.n2423 99.5127
R16927 vdd.n2420 vdd.n2419 99.5127
R16928 vdd.n2416 vdd.n2415 99.5127
R16929 vdd.n2412 vdd.n2411 99.5127
R16930 vdd.n2408 vdd.n2407 99.5127
R16931 vdd.n2404 vdd.n2403 99.5127
R16932 vdd.n2400 vdd.n2399 99.5127
R16933 vdd.n2396 vdd.n2395 99.5127
R16934 vdd.n2392 vdd.n2391 99.5127
R16935 vdd.n2388 vdd.n2387 99.5127
R16936 vdd.n2384 vdd.n2383 99.5127
R16937 vdd.n2380 vdd.n907 99.5127
R16938 vdd.n2137 vdd.n1022 99.5127
R16939 vdd.n2137 vdd.n1016 99.5127
R16940 vdd.n2140 vdd.n1016 99.5127
R16941 vdd.n2140 vdd.n1010 99.5127
R16942 vdd.n2143 vdd.n1010 99.5127
R16943 vdd.n2143 vdd.n1003 99.5127
R16944 vdd.n2146 vdd.n1003 99.5127
R16945 vdd.n2146 vdd.n996 99.5127
R16946 vdd.n2149 vdd.n996 99.5127
R16947 vdd.n2149 vdd.n991 99.5127
R16948 vdd.n2152 vdd.n991 99.5127
R16949 vdd.n2152 vdd.n985 99.5127
R16950 vdd.n2173 vdd.n985 99.5127
R16951 vdd.n2173 vdd.n978 99.5127
R16952 vdd.n2169 vdd.n978 99.5127
R16953 vdd.n2169 vdd.n972 99.5127
R16954 vdd.n2166 vdd.n972 99.5127
R16955 vdd.n2166 vdd.n967 99.5127
R16956 vdd.n2163 vdd.n967 99.5127
R16957 vdd.n2163 vdd.n962 99.5127
R16958 vdd.n2160 vdd.n962 99.5127
R16959 vdd.n2160 vdd.n956 99.5127
R16960 vdd.n2157 vdd.n956 99.5127
R16961 vdd.n2157 vdd.n949 99.5127
R16962 vdd.n949 vdd.n940 99.5127
R16963 vdd.n2375 vdd.n940 99.5127
R16964 vdd.n2376 vdd.n2375 99.5127
R16965 vdd.n2376 vdd.n932 99.5127
R16966 vdd.n2287 vdd.n2285 99.5127
R16967 vdd.n2283 vdd.n1025 99.5127
R16968 vdd.n2279 vdd.n2277 99.5127
R16969 vdd.n2275 vdd.n1027 99.5127
R16970 vdd.n2271 vdd.n2269 99.5127
R16971 vdd.n2267 vdd.n1029 99.5127
R16972 vdd.n2263 vdd.n2261 99.5127
R16973 vdd.n2259 vdd.n1031 99.5127
R16974 vdd.n2101 vdd.n1033 99.5127
R16975 vdd.n2106 vdd.n2103 99.5127
R16976 vdd.n2110 vdd.n2108 99.5127
R16977 vdd.n2114 vdd.n2099 99.5127
R16978 vdd.n2118 vdd.n2116 99.5127
R16979 vdd.n2122 vdd.n2097 99.5127
R16980 vdd.n2126 vdd.n2124 99.5127
R16981 vdd.n2131 vdd.n2093 99.5127
R16982 vdd.n2134 vdd.n2133 99.5127
R16983 vdd.n2291 vdd.n1013 99.5127
R16984 vdd.n2299 vdd.n1013 99.5127
R16985 vdd.n2299 vdd.n1011 99.5127
R16986 vdd.n2303 vdd.n1011 99.5127
R16987 vdd.n2303 vdd.n1000 99.5127
R16988 vdd.n2311 vdd.n1000 99.5127
R16989 vdd.n2311 vdd.n997 99.5127
R16990 vdd.n2316 vdd.n997 99.5127
R16991 vdd.n2316 vdd.n988 99.5127
R16992 vdd.n2324 vdd.n988 99.5127
R16993 vdd.n2324 vdd.n986 99.5127
R16994 vdd.n2328 vdd.n986 99.5127
R16995 vdd.n2328 vdd.n976 99.5127
R16996 vdd.n2336 vdd.n976 99.5127
R16997 vdd.n2336 vdd.n974 99.5127
R16998 vdd.n2340 vdd.n974 99.5127
R16999 vdd.n2340 vdd.n965 99.5127
R17000 vdd.n2348 vdd.n965 99.5127
R17001 vdd.n2348 vdd.n963 99.5127
R17002 vdd.n2352 vdd.n963 99.5127
R17003 vdd.n2352 vdd.n953 99.5127
R17004 vdd.n2360 vdd.n953 99.5127
R17005 vdd.n2360 vdd.n950 99.5127
R17006 vdd.n2366 vdd.n950 99.5127
R17007 vdd.n2366 vdd.n951 99.5127
R17008 vdd.n951 vdd.n942 99.5127
R17009 vdd.n942 vdd.n933 99.5127
R17010 vdd.n2448 vdd.n933 99.5127
R17011 vdd.n9 vdd.n7 98.9633
R17012 vdd.n2 vdd.n0 98.9633
R17013 vdd.n9 vdd.n8 98.6055
R17014 vdd.n11 vdd.n10 98.6055
R17015 vdd.n13 vdd.n12 98.6055
R17016 vdd.n6 vdd.n5 98.6055
R17017 vdd.n4 vdd.n3 98.6055
R17018 vdd.n2 vdd.n1 98.6055
R17019 vdd.t233 vdd.n291 85.8723
R17020 vdd.t205 vdd.n236 85.8723
R17021 vdd.t220 vdd.n193 85.8723
R17022 vdd.t197 vdd.n138 85.8723
R17023 vdd.t154 vdd.n96 85.8723
R17024 vdd.t135 vdd.n41 85.8723
R17025 vdd.t246 vdd.n1660 85.8723
R17026 vdd.t158 vdd.n1715 85.8723
R17027 vdd.t234 vdd.n1562 85.8723
R17028 vdd.t141 vdd.n1617 85.8723
R17029 vdd.t137 vdd.n1465 85.8723
R17030 vdd.t155 vdd.n1520 85.8723
R17031 vdd.n2840 vdd.n2839 78.546
R17032 vdd.n2314 vdd.n998 78.546
R17033 vdd.n278 vdd.n277 75.1835
R17034 vdd.n276 vdd.n275 75.1835
R17035 vdd.n274 vdd.n273 75.1835
R17036 vdd.n272 vdd.n271 75.1835
R17037 vdd.n270 vdd.n269 75.1835
R17038 vdd.n268 vdd.n267 75.1835
R17039 vdd.n266 vdd.n265 75.1835
R17040 vdd.n180 vdd.n179 75.1835
R17041 vdd.n178 vdd.n177 75.1835
R17042 vdd.n176 vdd.n175 75.1835
R17043 vdd.n174 vdd.n173 75.1835
R17044 vdd.n172 vdd.n171 75.1835
R17045 vdd.n170 vdd.n169 75.1835
R17046 vdd.n168 vdd.n167 75.1835
R17047 vdd.n83 vdd.n82 75.1835
R17048 vdd.n81 vdd.n80 75.1835
R17049 vdd.n79 vdd.n78 75.1835
R17050 vdd.n77 vdd.n76 75.1835
R17051 vdd.n75 vdd.n74 75.1835
R17052 vdd.n73 vdd.n72 75.1835
R17053 vdd.n71 vdd.n70 75.1835
R17054 vdd.n1690 vdd.n1689 75.1835
R17055 vdd.n1692 vdd.n1691 75.1835
R17056 vdd.n1694 vdd.n1693 75.1835
R17057 vdd.n1696 vdd.n1695 75.1835
R17058 vdd.n1698 vdd.n1697 75.1835
R17059 vdd.n1700 vdd.n1699 75.1835
R17060 vdd.n1702 vdd.n1701 75.1835
R17061 vdd.n1592 vdd.n1591 75.1835
R17062 vdd.n1594 vdd.n1593 75.1835
R17063 vdd.n1596 vdd.n1595 75.1835
R17064 vdd.n1598 vdd.n1597 75.1835
R17065 vdd.n1600 vdd.n1599 75.1835
R17066 vdd.n1602 vdd.n1601 75.1835
R17067 vdd.n1604 vdd.n1603 75.1835
R17068 vdd.n1495 vdd.n1494 75.1835
R17069 vdd.n1497 vdd.n1496 75.1835
R17070 vdd.n1499 vdd.n1498 75.1835
R17071 vdd.n1501 vdd.n1500 75.1835
R17072 vdd.n1503 vdd.n1502 75.1835
R17073 vdd.n1505 vdd.n1504 75.1835
R17074 vdd.n1507 vdd.n1506 75.1835
R17075 vdd.n2775 vdd.n2774 72.8958
R17076 vdd.n2774 vdd.n2538 72.8958
R17077 vdd.n2774 vdd.n2539 72.8958
R17078 vdd.n2774 vdd.n2540 72.8958
R17079 vdd.n2774 vdd.n2541 72.8958
R17080 vdd.n2774 vdd.n2542 72.8958
R17081 vdd.n2774 vdd.n2543 72.8958
R17082 vdd.n2774 vdd.n2544 72.8958
R17083 vdd.n2774 vdd.n2545 72.8958
R17084 vdd.n2774 vdd.n2546 72.8958
R17085 vdd.n2774 vdd.n2547 72.8958
R17086 vdd.n2774 vdd.n2548 72.8958
R17087 vdd.n2774 vdd.n2549 72.8958
R17088 vdd.n2774 vdd.n2550 72.8958
R17089 vdd.n2774 vdd.n2551 72.8958
R17090 vdd.n2774 vdd.n2552 72.8958
R17091 vdd.n2774 vdd.n2553 72.8958
R17092 vdd.n772 vdd.n756 72.8958
R17093 vdd.n2983 vdd.n756 72.8958
R17094 vdd.n766 vdd.n756 72.8958
R17095 vdd.n2990 vdd.n756 72.8958
R17096 vdd.n763 vdd.n756 72.8958
R17097 vdd.n2997 vdd.n756 72.8958
R17098 vdd.n760 vdd.n756 72.8958
R17099 vdd.n3004 vdd.n756 72.8958
R17100 vdd.n3007 vdd.n756 72.8958
R17101 vdd.n2863 vdd.n756 72.8958
R17102 vdd.n2868 vdd.n756 72.8958
R17103 vdd.n2862 vdd.n756 72.8958
R17104 vdd.n2875 vdd.n756 72.8958
R17105 vdd.n2859 vdd.n756 72.8958
R17106 vdd.n2882 vdd.n756 72.8958
R17107 vdd.n2856 vdd.n756 72.8958
R17108 vdd.n2889 vdd.n756 72.8958
R17109 vdd.n2027 vdd.n1020 72.8958
R17110 vdd.n2033 vdd.n1020 72.8958
R17111 vdd.n2035 vdd.n1020 72.8958
R17112 vdd.n2041 vdd.n1020 72.8958
R17113 vdd.n2043 vdd.n1020 72.8958
R17114 vdd.n2049 vdd.n1020 72.8958
R17115 vdd.n2051 vdd.n1020 72.8958
R17116 vdd.n2057 vdd.n1020 72.8958
R17117 vdd.n2228 vdd.n1020 72.8958
R17118 vdd.n2226 vdd.n1020 72.8958
R17119 vdd.n2220 vdd.n1020 72.8958
R17120 vdd.n2218 vdd.n1020 72.8958
R17121 vdd.n2212 vdd.n1020 72.8958
R17122 vdd.n2210 vdd.n1020 72.8958
R17123 vdd.n2204 vdd.n1020 72.8958
R17124 vdd.n2202 vdd.n1020 72.8958
R17125 vdd.n2196 vdd.n1020 72.8958
R17126 vdd.n2521 vdd.n908 72.8958
R17127 vdd.n2521 vdd.n909 72.8958
R17128 vdd.n2521 vdd.n910 72.8958
R17129 vdd.n2521 vdd.n911 72.8958
R17130 vdd.n2521 vdd.n912 72.8958
R17131 vdd.n2521 vdd.n913 72.8958
R17132 vdd.n2521 vdd.n914 72.8958
R17133 vdd.n2521 vdd.n915 72.8958
R17134 vdd.n2521 vdd.n916 72.8958
R17135 vdd.n2521 vdd.n917 72.8958
R17136 vdd.n2521 vdd.n918 72.8958
R17137 vdd.n2521 vdd.n919 72.8958
R17138 vdd.n2521 vdd.n920 72.8958
R17139 vdd.n2521 vdd.n921 72.8958
R17140 vdd.n2521 vdd.n922 72.8958
R17141 vdd.n2521 vdd.n923 72.8958
R17142 vdd.n2521 vdd.n924 72.8958
R17143 vdd.n2774 vdd.n2773 72.8958
R17144 vdd.n2774 vdd.n2522 72.8958
R17145 vdd.n2774 vdd.n2523 72.8958
R17146 vdd.n2774 vdd.n2524 72.8958
R17147 vdd.n2774 vdd.n2525 72.8958
R17148 vdd.n2774 vdd.n2526 72.8958
R17149 vdd.n2774 vdd.n2527 72.8958
R17150 vdd.n2774 vdd.n2528 72.8958
R17151 vdd.n2774 vdd.n2529 72.8958
R17152 vdd.n2774 vdd.n2530 72.8958
R17153 vdd.n2774 vdd.n2531 72.8958
R17154 vdd.n2774 vdd.n2532 72.8958
R17155 vdd.n2774 vdd.n2533 72.8958
R17156 vdd.n2774 vdd.n2534 72.8958
R17157 vdd.n2774 vdd.n2535 72.8958
R17158 vdd.n2774 vdd.n2536 72.8958
R17159 vdd.n2774 vdd.n2537 72.8958
R17160 vdd.n2911 vdd.n756 72.8958
R17161 vdd.n2917 vdd.n756 72.8958
R17162 vdd.n802 vdd.n756 72.8958
R17163 vdd.n2924 vdd.n756 72.8958
R17164 vdd.n799 vdd.n756 72.8958
R17165 vdd.n2931 vdd.n756 72.8958
R17166 vdd.n796 vdd.n756 72.8958
R17167 vdd.n2938 vdd.n756 72.8958
R17168 vdd.n793 vdd.n756 72.8958
R17169 vdd.n2946 vdd.n756 72.8958
R17170 vdd.n790 vdd.n756 72.8958
R17171 vdd.n2953 vdd.n756 72.8958
R17172 vdd.n787 vdd.n756 72.8958
R17173 vdd.n2960 vdd.n756 72.8958
R17174 vdd.n784 vdd.n756 72.8958
R17175 vdd.n2967 vdd.n756 72.8958
R17176 vdd.n2970 vdd.n756 72.8958
R17177 vdd.n2521 vdd.n906 72.8958
R17178 vdd.n2521 vdd.n905 72.8958
R17179 vdd.n2521 vdd.n904 72.8958
R17180 vdd.n2521 vdd.n903 72.8958
R17181 vdd.n2521 vdd.n902 72.8958
R17182 vdd.n2521 vdd.n901 72.8958
R17183 vdd.n2521 vdd.n900 72.8958
R17184 vdd.n2521 vdd.n899 72.8958
R17185 vdd.n2521 vdd.n898 72.8958
R17186 vdd.n2521 vdd.n897 72.8958
R17187 vdd.n2521 vdd.n896 72.8958
R17188 vdd.n2521 vdd.n895 72.8958
R17189 vdd.n2521 vdd.n894 72.8958
R17190 vdd.n2521 vdd.n893 72.8958
R17191 vdd.n2521 vdd.n892 72.8958
R17192 vdd.n2521 vdd.n891 72.8958
R17193 vdd.n2521 vdd.n890 72.8958
R17194 vdd.n2286 vdd.n1020 72.8958
R17195 vdd.n2284 vdd.n1020 72.8958
R17196 vdd.n2278 vdd.n1020 72.8958
R17197 vdd.n2276 vdd.n1020 72.8958
R17198 vdd.n2270 vdd.n1020 72.8958
R17199 vdd.n2268 vdd.n1020 72.8958
R17200 vdd.n2262 vdd.n1020 72.8958
R17201 vdd.n2260 vdd.n1020 72.8958
R17202 vdd.n1032 vdd.n1020 72.8958
R17203 vdd.n2102 vdd.n1020 72.8958
R17204 vdd.n2107 vdd.n1020 72.8958
R17205 vdd.n2109 vdd.n1020 72.8958
R17206 vdd.n2115 vdd.n1020 72.8958
R17207 vdd.n2117 vdd.n1020 72.8958
R17208 vdd.n2123 vdd.n1020 72.8958
R17209 vdd.n2125 vdd.n1020 72.8958
R17210 vdd.n2132 vdd.n1020 72.8958
R17211 vdd.n1374 vdd.n1373 66.2847
R17212 vdd.n1374 vdd.n1152 66.2847
R17213 vdd.n1374 vdd.n1153 66.2847
R17214 vdd.n1374 vdd.n1154 66.2847
R17215 vdd.n1374 vdd.n1155 66.2847
R17216 vdd.n1374 vdd.n1156 66.2847
R17217 vdd.n1374 vdd.n1157 66.2847
R17218 vdd.n1374 vdd.n1158 66.2847
R17219 vdd.n1374 vdd.n1159 66.2847
R17220 vdd.n1374 vdd.n1160 66.2847
R17221 vdd.n1374 vdd.n1161 66.2847
R17222 vdd.n1374 vdd.n1162 66.2847
R17223 vdd.n1374 vdd.n1163 66.2847
R17224 vdd.n1374 vdd.n1164 66.2847
R17225 vdd.n1374 vdd.n1165 66.2847
R17226 vdd.n1374 vdd.n1166 66.2847
R17227 vdd.n1374 vdd.n1167 66.2847
R17228 vdd.n1374 vdd.n1168 66.2847
R17229 vdd.n1374 vdd.n1169 66.2847
R17230 vdd.n1374 vdd.n1170 66.2847
R17231 vdd.n1374 vdd.n1171 66.2847
R17232 vdd.n1374 vdd.n1172 66.2847
R17233 vdd.n1374 vdd.n1173 66.2847
R17234 vdd.n1374 vdd.n1174 66.2847
R17235 vdd.n1374 vdd.n1175 66.2847
R17236 vdd.n1374 vdd.n1176 66.2847
R17237 vdd.n1374 vdd.n1177 66.2847
R17238 vdd.n1374 vdd.n1178 66.2847
R17239 vdd.n1374 vdd.n1179 66.2847
R17240 vdd.n1374 vdd.n1180 66.2847
R17241 vdd.n1374 vdd.n1181 66.2847
R17242 vdd.n1045 vdd.n1041 66.2847
R17243 vdd.n1917 vdd.n1045 66.2847
R17244 vdd.n1922 vdd.n1045 66.2847
R17245 vdd.n1927 vdd.n1045 66.2847
R17246 vdd.n1915 vdd.n1045 66.2847
R17247 vdd.n1934 vdd.n1045 66.2847
R17248 vdd.n1907 vdd.n1045 66.2847
R17249 vdd.n1941 vdd.n1045 66.2847
R17250 vdd.n1900 vdd.n1045 66.2847
R17251 vdd.n1948 vdd.n1045 66.2847
R17252 vdd.n1894 vdd.n1045 66.2847
R17253 vdd.n1889 vdd.n1045 66.2847
R17254 vdd.n1959 vdd.n1045 66.2847
R17255 vdd.n1881 vdd.n1045 66.2847
R17256 vdd.n1966 vdd.n1045 66.2847
R17257 vdd.n1874 vdd.n1045 66.2847
R17258 vdd.n1973 vdd.n1045 66.2847
R17259 vdd.n1867 vdd.n1045 66.2847
R17260 vdd.n1980 vdd.n1045 66.2847
R17261 vdd.n1860 vdd.n1045 66.2847
R17262 vdd.n1987 vdd.n1045 66.2847
R17263 vdd.n1854 vdd.n1045 66.2847
R17264 vdd.n1849 vdd.n1045 66.2847
R17265 vdd.n1998 vdd.n1045 66.2847
R17266 vdd.n1841 vdd.n1045 66.2847
R17267 vdd.n2005 vdd.n1045 66.2847
R17268 vdd.n1834 vdd.n1045 66.2847
R17269 vdd.n2012 vdd.n1045 66.2847
R17270 vdd.n2015 vdd.n1045 66.2847
R17271 vdd.n1825 vdd.n1045 66.2847
R17272 vdd.n2237 vdd.n1045 66.2847
R17273 vdd.n1819 vdd.n1045 66.2847
R17274 vdd.n3137 vdd.n658 66.2847
R17275 vdd.n663 vdd.n658 66.2847
R17276 vdd.n666 vdd.n658 66.2847
R17277 vdd.n3126 vdd.n658 66.2847
R17278 vdd.n3120 vdd.n658 66.2847
R17279 vdd.n3118 vdd.n658 66.2847
R17280 vdd.n3112 vdd.n658 66.2847
R17281 vdd.n3110 vdd.n658 66.2847
R17282 vdd.n3104 vdd.n658 66.2847
R17283 vdd.n3102 vdd.n658 66.2847
R17284 vdd.n3096 vdd.n658 66.2847
R17285 vdd.n3094 vdd.n658 66.2847
R17286 vdd.n3088 vdd.n658 66.2847
R17287 vdd.n3086 vdd.n658 66.2847
R17288 vdd.n3080 vdd.n658 66.2847
R17289 vdd.n3078 vdd.n658 66.2847
R17290 vdd.n3072 vdd.n658 66.2847
R17291 vdd.n3070 vdd.n658 66.2847
R17292 vdd.n3064 vdd.n658 66.2847
R17293 vdd.n3062 vdd.n658 66.2847
R17294 vdd.n727 vdd.n658 66.2847
R17295 vdd.n3053 vdd.n658 66.2847
R17296 vdd.n729 vdd.n658 66.2847
R17297 vdd.n3046 vdd.n658 66.2847
R17298 vdd.n3040 vdd.n658 66.2847
R17299 vdd.n3038 vdd.n658 66.2847
R17300 vdd.n3032 vdd.n658 66.2847
R17301 vdd.n3030 vdd.n658 66.2847
R17302 vdd.n3024 vdd.n658 66.2847
R17303 vdd.n750 vdd.n658 66.2847
R17304 vdd.n752 vdd.n658 66.2847
R17305 vdd.n3253 vdd.n3252 66.2847
R17306 vdd.n3253 vdd.n403 66.2847
R17307 vdd.n3253 vdd.n402 66.2847
R17308 vdd.n3253 vdd.n401 66.2847
R17309 vdd.n3253 vdd.n400 66.2847
R17310 vdd.n3253 vdd.n399 66.2847
R17311 vdd.n3253 vdd.n398 66.2847
R17312 vdd.n3253 vdd.n397 66.2847
R17313 vdd.n3253 vdd.n396 66.2847
R17314 vdd.n3253 vdd.n395 66.2847
R17315 vdd.n3253 vdd.n394 66.2847
R17316 vdd.n3253 vdd.n393 66.2847
R17317 vdd.n3253 vdd.n392 66.2847
R17318 vdd.n3253 vdd.n391 66.2847
R17319 vdd.n3253 vdd.n390 66.2847
R17320 vdd.n3253 vdd.n389 66.2847
R17321 vdd.n3253 vdd.n388 66.2847
R17322 vdd.n3253 vdd.n387 66.2847
R17323 vdd.n3253 vdd.n386 66.2847
R17324 vdd.n3253 vdd.n385 66.2847
R17325 vdd.n3253 vdd.n384 66.2847
R17326 vdd.n3253 vdd.n383 66.2847
R17327 vdd.n3253 vdd.n382 66.2847
R17328 vdd.n3253 vdd.n381 66.2847
R17329 vdd.n3253 vdd.n380 66.2847
R17330 vdd.n3253 vdd.n379 66.2847
R17331 vdd.n3253 vdd.n378 66.2847
R17332 vdd.n3253 vdd.n377 66.2847
R17333 vdd.n3253 vdd.n376 66.2847
R17334 vdd.n3253 vdd.n375 66.2847
R17335 vdd.n3253 vdd.n374 66.2847
R17336 vdd.n3253 vdd.n373 66.2847
R17337 vdd.n448 vdd.n373 52.4337
R17338 vdd.n454 vdd.n374 52.4337
R17339 vdd.n458 vdd.n375 52.4337
R17340 vdd.n464 vdd.n376 52.4337
R17341 vdd.n468 vdd.n377 52.4337
R17342 vdd.n474 vdd.n378 52.4337
R17343 vdd.n478 vdd.n379 52.4337
R17344 vdd.n484 vdd.n380 52.4337
R17345 vdd.n488 vdd.n381 52.4337
R17346 vdd.n494 vdd.n382 52.4337
R17347 vdd.n498 vdd.n383 52.4337
R17348 vdd.n504 vdd.n384 52.4337
R17349 vdd.n508 vdd.n385 52.4337
R17350 vdd.n514 vdd.n386 52.4337
R17351 vdd.n518 vdd.n387 52.4337
R17352 vdd.n524 vdd.n388 52.4337
R17353 vdd.n528 vdd.n389 52.4337
R17354 vdd.n534 vdd.n390 52.4337
R17355 vdd.n538 vdd.n391 52.4337
R17356 vdd.n544 vdd.n392 52.4337
R17357 vdd.n548 vdd.n393 52.4337
R17358 vdd.n554 vdd.n394 52.4337
R17359 vdd.n558 vdd.n395 52.4337
R17360 vdd.n564 vdd.n396 52.4337
R17361 vdd.n568 vdd.n397 52.4337
R17362 vdd.n574 vdd.n398 52.4337
R17363 vdd.n578 vdd.n399 52.4337
R17364 vdd.n584 vdd.n400 52.4337
R17365 vdd.n588 vdd.n401 52.4337
R17366 vdd.n594 vdd.n402 52.4337
R17367 vdd.n597 vdd.n403 52.4337
R17368 vdd.n3252 vdd.n3251 52.4337
R17369 vdd.n3137 vdd.n660 52.4337
R17370 vdd.n3135 vdd.n663 52.4337
R17371 vdd.n3131 vdd.n666 52.4337
R17372 vdd.n3127 vdd.n3126 52.4337
R17373 vdd.n3120 vdd.n669 52.4337
R17374 vdd.n3119 vdd.n3118 52.4337
R17375 vdd.n3112 vdd.n675 52.4337
R17376 vdd.n3111 vdd.n3110 52.4337
R17377 vdd.n3104 vdd.n681 52.4337
R17378 vdd.n3103 vdd.n3102 52.4337
R17379 vdd.n3096 vdd.n689 52.4337
R17380 vdd.n3095 vdd.n3094 52.4337
R17381 vdd.n3088 vdd.n695 52.4337
R17382 vdd.n3087 vdd.n3086 52.4337
R17383 vdd.n3080 vdd.n701 52.4337
R17384 vdd.n3079 vdd.n3078 52.4337
R17385 vdd.n3072 vdd.n707 52.4337
R17386 vdd.n3071 vdd.n3070 52.4337
R17387 vdd.n3064 vdd.n713 52.4337
R17388 vdd.n3063 vdd.n3062 52.4337
R17389 vdd.n727 vdd.n719 52.4337
R17390 vdd.n3054 vdd.n3053 52.4337
R17391 vdd.n3051 vdd.n729 52.4337
R17392 vdd.n3047 vdd.n3046 52.4337
R17393 vdd.n3040 vdd.n733 52.4337
R17394 vdd.n3039 vdd.n3038 52.4337
R17395 vdd.n3032 vdd.n739 52.4337
R17396 vdd.n3031 vdd.n3030 52.4337
R17397 vdd.n3024 vdd.n745 52.4337
R17398 vdd.n3023 vdd.n750 52.4337
R17399 vdd.n3019 vdd.n752 52.4337
R17400 vdd.n2239 vdd.n1819 52.4337
R17401 vdd.n2237 vdd.n2236 52.4337
R17402 vdd.n1826 vdd.n1825 52.4337
R17403 vdd.n2015 vdd.n2014 52.4337
R17404 vdd.n2012 vdd.n2011 52.4337
R17405 vdd.n2007 vdd.n1834 52.4337
R17406 vdd.n2005 vdd.n2004 52.4337
R17407 vdd.n2000 vdd.n1841 52.4337
R17408 vdd.n1998 vdd.n1997 52.4337
R17409 vdd.n1850 vdd.n1849 52.4337
R17410 vdd.n1989 vdd.n1854 52.4337
R17411 vdd.n1987 vdd.n1986 52.4337
R17412 vdd.n1982 vdd.n1860 52.4337
R17413 vdd.n1980 vdd.n1979 52.4337
R17414 vdd.n1975 vdd.n1867 52.4337
R17415 vdd.n1973 vdd.n1972 52.4337
R17416 vdd.n1968 vdd.n1874 52.4337
R17417 vdd.n1966 vdd.n1965 52.4337
R17418 vdd.n1961 vdd.n1881 52.4337
R17419 vdd.n1959 vdd.n1958 52.4337
R17420 vdd.n1890 vdd.n1889 52.4337
R17421 vdd.n1950 vdd.n1894 52.4337
R17422 vdd.n1948 vdd.n1947 52.4337
R17423 vdd.n1943 vdd.n1900 52.4337
R17424 vdd.n1941 vdd.n1940 52.4337
R17425 vdd.n1936 vdd.n1907 52.4337
R17426 vdd.n1934 vdd.n1933 52.4337
R17427 vdd.n1929 vdd.n1915 52.4337
R17428 vdd.n1927 vdd.n1926 52.4337
R17429 vdd.n1922 vdd.n1921 52.4337
R17430 vdd.n1917 vdd.n1916 52.4337
R17431 vdd.n2248 vdd.n1041 52.4337
R17432 vdd.n1373 vdd.n1372 52.4337
R17433 vdd.n1187 vdd.n1152 52.4337
R17434 vdd.n1189 vdd.n1153 52.4337
R17435 vdd.n1193 vdd.n1154 52.4337
R17436 vdd.n1195 vdd.n1155 52.4337
R17437 vdd.n1199 vdd.n1156 52.4337
R17438 vdd.n1201 vdd.n1157 52.4337
R17439 vdd.n1205 vdd.n1158 52.4337
R17440 vdd.n1207 vdd.n1159 52.4337
R17441 vdd.n1339 vdd.n1160 52.4337
R17442 vdd.n1211 vdd.n1161 52.4337
R17443 vdd.n1215 vdd.n1162 52.4337
R17444 vdd.n1217 vdd.n1163 52.4337
R17445 vdd.n1221 vdd.n1164 52.4337
R17446 vdd.n1223 vdd.n1165 52.4337
R17447 vdd.n1227 vdd.n1166 52.4337
R17448 vdd.n1229 vdd.n1167 52.4337
R17449 vdd.n1233 vdd.n1168 52.4337
R17450 vdd.n1235 vdd.n1169 52.4337
R17451 vdd.n1239 vdd.n1170 52.4337
R17452 vdd.n1303 vdd.n1171 52.4337
R17453 vdd.n1244 vdd.n1172 52.4337
R17454 vdd.n1246 vdd.n1173 52.4337
R17455 vdd.n1250 vdd.n1174 52.4337
R17456 vdd.n1252 vdd.n1175 52.4337
R17457 vdd.n1256 vdd.n1176 52.4337
R17458 vdd.n1258 vdd.n1177 52.4337
R17459 vdd.n1262 vdd.n1178 52.4337
R17460 vdd.n1264 vdd.n1179 52.4337
R17461 vdd.n1268 vdd.n1180 52.4337
R17462 vdd.n1270 vdd.n1181 52.4337
R17463 vdd.n1373 vdd.n1183 52.4337
R17464 vdd.n1188 vdd.n1152 52.4337
R17465 vdd.n1192 vdd.n1153 52.4337
R17466 vdd.n1194 vdd.n1154 52.4337
R17467 vdd.n1198 vdd.n1155 52.4337
R17468 vdd.n1200 vdd.n1156 52.4337
R17469 vdd.n1204 vdd.n1157 52.4337
R17470 vdd.n1206 vdd.n1158 52.4337
R17471 vdd.n1338 vdd.n1159 52.4337
R17472 vdd.n1210 vdd.n1160 52.4337
R17473 vdd.n1214 vdd.n1161 52.4337
R17474 vdd.n1216 vdd.n1162 52.4337
R17475 vdd.n1220 vdd.n1163 52.4337
R17476 vdd.n1222 vdd.n1164 52.4337
R17477 vdd.n1226 vdd.n1165 52.4337
R17478 vdd.n1228 vdd.n1166 52.4337
R17479 vdd.n1232 vdd.n1167 52.4337
R17480 vdd.n1234 vdd.n1168 52.4337
R17481 vdd.n1238 vdd.n1169 52.4337
R17482 vdd.n1240 vdd.n1170 52.4337
R17483 vdd.n1243 vdd.n1171 52.4337
R17484 vdd.n1245 vdd.n1172 52.4337
R17485 vdd.n1249 vdd.n1173 52.4337
R17486 vdd.n1251 vdd.n1174 52.4337
R17487 vdd.n1255 vdd.n1175 52.4337
R17488 vdd.n1257 vdd.n1176 52.4337
R17489 vdd.n1261 vdd.n1177 52.4337
R17490 vdd.n1263 vdd.n1178 52.4337
R17491 vdd.n1267 vdd.n1179 52.4337
R17492 vdd.n1269 vdd.n1180 52.4337
R17493 vdd.n1181 vdd.n1151 52.4337
R17494 vdd.n1041 vdd.n1040 52.4337
R17495 vdd.n1918 vdd.n1917 52.4337
R17496 vdd.n1923 vdd.n1922 52.4337
R17497 vdd.n1928 vdd.n1927 52.4337
R17498 vdd.n1915 vdd.n1908 52.4337
R17499 vdd.n1935 vdd.n1934 52.4337
R17500 vdd.n1907 vdd.n1901 52.4337
R17501 vdd.n1942 vdd.n1941 52.4337
R17502 vdd.n1900 vdd.n1895 52.4337
R17503 vdd.n1949 vdd.n1948 52.4337
R17504 vdd.n1894 vdd.n1893 52.4337
R17505 vdd.n1889 vdd.n1882 52.4337
R17506 vdd.n1960 vdd.n1959 52.4337
R17507 vdd.n1881 vdd.n1875 52.4337
R17508 vdd.n1967 vdd.n1966 52.4337
R17509 vdd.n1874 vdd.n1868 52.4337
R17510 vdd.n1974 vdd.n1973 52.4337
R17511 vdd.n1867 vdd.n1861 52.4337
R17512 vdd.n1981 vdd.n1980 52.4337
R17513 vdd.n1860 vdd.n1855 52.4337
R17514 vdd.n1988 vdd.n1987 52.4337
R17515 vdd.n1854 vdd.n1853 52.4337
R17516 vdd.n1849 vdd.n1842 52.4337
R17517 vdd.n1999 vdd.n1998 52.4337
R17518 vdd.n1841 vdd.n1835 52.4337
R17519 vdd.n2006 vdd.n2005 52.4337
R17520 vdd.n1834 vdd.n1828 52.4337
R17521 vdd.n2013 vdd.n2012 52.4337
R17522 vdd.n2016 vdd.n2015 52.4337
R17523 vdd.n1825 vdd.n1820 52.4337
R17524 vdd.n2238 vdd.n2237 52.4337
R17525 vdd.n1819 vdd.n1047 52.4337
R17526 vdd.n3138 vdd.n3137 52.4337
R17527 vdd.n3132 vdd.n663 52.4337
R17528 vdd.n3128 vdd.n666 52.4337
R17529 vdd.n3126 vdd.n3125 52.4337
R17530 vdd.n3121 vdd.n3120 52.4337
R17531 vdd.n3118 vdd.n3117 52.4337
R17532 vdd.n3113 vdd.n3112 52.4337
R17533 vdd.n3110 vdd.n3109 52.4337
R17534 vdd.n3105 vdd.n3104 52.4337
R17535 vdd.n3102 vdd.n3101 52.4337
R17536 vdd.n3097 vdd.n3096 52.4337
R17537 vdd.n3094 vdd.n3093 52.4337
R17538 vdd.n3089 vdd.n3088 52.4337
R17539 vdd.n3086 vdd.n3085 52.4337
R17540 vdd.n3081 vdd.n3080 52.4337
R17541 vdd.n3078 vdd.n3077 52.4337
R17542 vdd.n3073 vdd.n3072 52.4337
R17543 vdd.n3070 vdd.n3069 52.4337
R17544 vdd.n3065 vdd.n3064 52.4337
R17545 vdd.n3062 vdd.n3061 52.4337
R17546 vdd.n728 vdd.n727 52.4337
R17547 vdd.n3053 vdd.n3052 52.4337
R17548 vdd.n3048 vdd.n729 52.4337
R17549 vdd.n3046 vdd.n3045 52.4337
R17550 vdd.n3041 vdd.n3040 52.4337
R17551 vdd.n3038 vdd.n3037 52.4337
R17552 vdd.n3033 vdd.n3032 52.4337
R17553 vdd.n3030 vdd.n3029 52.4337
R17554 vdd.n3025 vdd.n3024 52.4337
R17555 vdd.n3020 vdd.n750 52.4337
R17556 vdd.n3016 vdd.n752 52.4337
R17557 vdd.n3252 vdd.n404 52.4337
R17558 vdd.n595 vdd.n403 52.4337
R17559 vdd.n589 vdd.n402 52.4337
R17560 vdd.n585 vdd.n401 52.4337
R17561 vdd.n579 vdd.n400 52.4337
R17562 vdd.n575 vdd.n399 52.4337
R17563 vdd.n569 vdd.n398 52.4337
R17564 vdd.n565 vdd.n397 52.4337
R17565 vdd.n559 vdd.n396 52.4337
R17566 vdd.n555 vdd.n395 52.4337
R17567 vdd.n549 vdd.n394 52.4337
R17568 vdd.n545 vdd.n393 52.4337
R17569 vdd.n539 vdd.n392 52.4337
R17570 vdd.n535 vdd.n391 52.4337
R17571 vdd.n529 vdd.n390 52.4337
R17572 vdd.n525 vdd.n389 52.4337
R17573 vdd.n519 vdd.n388 52.4337
R17574 vdd.n515 vdd.n387 52.4337
R17575 vdd.n509 vdd.n386 52.4337
R17576 vdd.n505 vdd.n385 52.4337
R17577 vdd.n499 vdd.n384 52.4337
R17578 vdd.n495 vdd.n383 52.4337
R17579 vdd.n489 vdd.n382 52.4337
R17580 vdd.n485 vdd.n381 52.4337
R17581 vdd.n479 vdd.n380 52.4337
R17582 vdd.n475 vdd.n379 52.4337
R17583 vdd.n469 vdd.n378 52.4337
R17584 vdd.n465 vdd.n377 52.4337
R17585 vdd.n459 vdd.n376 52.4337
R17586 vdd.n455 vdd.n375 52.4337
R17587 vdd.n449 vdd.n374 52.4337
R17588 vdd.n445 vdd.n373 52.4337
R17589 vdd.t262 vdd.t13 51.4683
R17590 vdd.n266 vdd.n264 42.0461
R17591 vdd.n168 vdd.n166 42.0461
R17592 vdd.n71 vdd.n69 42.0461
R17593 vdd.n1690 vdd.n1688 42.0461
R17594 vdd.n1592 vdd.n1590 42.0461
R17595 vdd.n1495 vdd.n1493 42.0461
R17596 vdd.n320 vdd.n319 41.6884
R17597 vdd.n222 vdd.n221 41.6884
R17598 vdd.n125 vdd.n124 41.6884
R17599 vdd.n1744 vdd.n1743 41.6884
R17600 vdd.n1646 vdd.n1645 41.6884
R17601 vdd.n1549 vdd.n1548 41.6884
R17602 vdd.n1150 vdd.n1149 41.1157
R17603 vdd.n1306 vdd.n1305 41.1157
R17604 vdd.n1342 vdd.n1341 41.1157
R17605 vdd.n407 vdd.n406 41.1157
R17606 vdd.n547 vdd.n420 41.1157
R17607 vdd.n433 vdd.n432 41.1157
R17608 vdd.n2970 vdd.n2969 39.2114
R17609 vdd.n2967 vdd.n2966 39.2114
R17610 vdd.n2962 vdd.n784 39.2114
R17611 vdd.n2960 vdd.n2959 39.2114
R17612 vdd.n2955 vdd.n787 39.2114
R17613 vdd.n2953 vdd.n2952 39.2114
R17614 vdd.n2948 vdd.n790 39.2114
R17615 vdd.n2946 vdd.n2945 39.2114
R17616 vdd.n2940 vdd.n793 39.2114
R17617 vdd.n2938 vdd.n2937 39.2114
R17618 vdd.n2933 vdd.n796 39.2114
R17619 vdd.n2931 vdd.n2930 39.2114
R17620 vdd.n2926 vdd.n799 39.2114
R17621 vdd.n2924 vdd.n2923 39.2114
R17622 vdd.n2919 vdd.n802 39.2114
R17623 vdd.n2917 vdd.n2916 39.2114
R17624 vdd.n2912 vdd.n2911 39.2114
R17625 vdd.n2773 vdd.n884 39.2114
R17626 vdd.n2768 vdd.n2522 39.2114
R17627 vdd.n2765 vdd.n2523 39.2114
R17628 vdd.n2761 vdd.n2524 39.2114
R17629 vdd.n2757 vdd.n2525 39.2114
R17630 vdd.n2753 vdd.n2526 39.2114
R17631 vdd.n2749 vdd.n2527 39.2114
R17632 vdd.n2745 vdd.n2528 39.2114
R17633 vdd.n2741 vdd.n2529 39.2114
R17634 vdd.n2737 vdd.n2530 39.2114
R17635 vdd.n2733 vdd.n2531 39.2114
R17636 vdd.n2729 vdd.n2532 39.2114
R17637 vdd.n2725 vdd.n2533 39.2114
R17638 vdd.n2721 vdd.n2534 39.2114
R17639 vdd.n2717 vdd.n2535 39.2114
R17640 vdd.n2713 vdd.n2536 39.2114
R17641 vdd.n2708 vdd.n2537 39.2114
R17642 vdd.n2516 vdd.n924 39.2114
R17643 vdd.n2512 vdd.n923 39.2114
R17644 vdd.n2508 vdd.n922 39.2114
R17645 vdd.n2504 vdd.n921 39.2114
R17646 vdd.n2500 vdd.n920 39.2114
R17647 vdd.n2496 vdd.n919 39.2114
R17648 vdd.n2492 vdd.n918 39.2114
R17649 vdd.n2488 vdd.n917 39.2114
R17650 vdd.n2484 vdd.n916 39.2114
R17651 vdd.n2480 vdd.n915 39.2114
R17652 vdd.n2476 vdd.n914 39.2114
R17653 vdd.n2472 vdd.n913 39.2114
R17654 vdd.n2468 vdd.n912 39.2114
R17655 vdd.n2464 vdd.n911 39.2114
R17656 vdd.n2460 vdd.n910 39.2114
R17657 vdd.n2455 vdd.n909 39.2114
R17658 vdd.n2451 vdd.n908 39.2114
R17659 vdd.n2027 vdd.n1019 39.2114
R17660 vdd.n2033 vdd.n2032 39.2114
R17661 vdd.n2036 vdd.n2035 39.2114
R17662 vdd.n2041 vdd.n2040 39.2114
R17663 vdd.n2044 vdd.n2043 39.2114
R17664 vdd.n2049 vdd.n2048 39.2114
R17665 vdd.n2052 vdd.n2051 39.2114
R17666 vdd.n2057 vdd.n2056 39.2114
R17667 vdd.n2228 vdd.n2059 39.2114
R17668 vdd.n2227 vdd.n2226 39.2114
R17669 vdd.n2220 vdd.n2061 39.2114
R17670 vdd.n2219 vdd.n2218 39.2114
R17671 vdd.n2212 vdd.n2063 39.2114
R17672 vdd.n2211 vdd.n2210 39.2114
R17673 vdd.n2204 vdd.n2065 39.2114
R17674 vdd.n2203 vdd.n2202 39.2114
R17675 vdd.n2196 vdd.n2067 39.2114
R17676 vdd.n2889 vdd.n2888 39.2114
R17677 vdd.n2884 vdd.n2856 39.2114
R17678 vdd.n2882 vdd.n2881 39.2114
R17679 vdd.n2877 vdd.n2859 39.2114
R17680 vdd.n2875 vdd.n2874 39.2114
R17681 vdd.n2870 vdd.n2862 39.2114
R17682 vdd.n2868 vdd.n2867 39.2114
R17683 vdd.n2863 vdd.n755 39.2114
R17684 vdd.n3007 vdd.n3006 39.2114
R17685 vdd.n3004 vdd.n3003 39.2114
R17686 vdd.n2999 vdd.n760 39.2114
R17687 vdd.n2997 vdd.n2996 39.2114
R17688 vdd.n2992 vdd.n763 39.2114
R17689 vdd.n2990 vdd.n2989 39.2114
R17690 vdd.n2985 vdd.n766 39.2114
R17691 vdd.n2983 vdd.n2982 39.2114
R17692 vdd.n2978 vdd.n772 39.2114
R17693 vdd.n2775 vdd.n887 39.2114
R17694 vdd.n2538 vdd.n889 39.2114
R17695 vdd.n2564 vdd.n2539 39.2114
R17696 vdd.n2568 vdd.n2540 39.2114
R17697 vdd.n2572 vdd.n2541 39.2114
R17698 vdd.n2576 vdd.n2542 39.2114
R17699 vdd.n2580 vdd.n2543 39.2114
R17700 vdd.n2584 vdd.n2544 39.2114
R17701 vdd.n2588 vdd.n2545 39.2114
R17702 vdd.n2592 vdd.n2546 39.2114
R17703 vdd.n2596 vdd.n2547 39.2114
R17704 vdd.n2600 vdd.n2548 39.2114
R17705 vdd.n2604 vdd.n2549 39.2114
R17706 vdd.n2608 vdd.n2550 39.2114
R17707 vdd.n2612 vdd.n2551 39.2114
R17708 vdd.n2616 vdd.n2552 39.2114
R17709 vdd.n2620 vdd.n2553 39.2114
R17710 vdd.n2776 vdd.n2775 39.2114
R17711 vdd.n2563 vdd.n2538 39.2114
R17712 vdd.n2567 vdd.n2539 39.2114
R17713 vdd.n2571 vdd.n2540 39.2114
R17714 vdd.n2575 vdd.n2541 39.2114
R17715 vdd.n2579 vdd.n2542 39.2114
R17716 vdd.n2583 vdd.n2543 39.2114
R17717 vdd.n2587 vdd.n2544 39.2114
R17718 vdd.n2591 vdd.n2545 39.2114
R17719 vdd.n2595 vdd.n2546 39.2114
R17720 vdd.n2599 vdd.n2547 39.2114
R17721 vdd.n2603 vdd.n2548 39.2114
R17722 vdd.n2607 vdd.n2549 39.2114
R17723 vdd.n2611 vdd.n2550 39.2114
R17724 vdd.n2615 vdd.n2551 39.2114
R17725 vdd.n2619 vdd.n2552 39.2114
R17726 vdd.n2622 vdd.n2553 39.2114
R17727 vdd.n772 vdd.n767 39.2114
R17728 vdd.n2984 vdd.n2983 39.2114
R17729 vdd.n766 vdd.n764 39.2114
R17730 vdd.n2991 vdd.n2990 39.2114
R17731 vdd.n763 vdd.n761 39.2114
R17732 vdd.n2998 vdd.n2997 39.2114
R17733 vdd.n760 vdd.n758 39.2114
R17734 vdd.n3005 vdd.n3004 39.2114
R17735 vdd.n3008 vdd.n3007 39.2114
R17736 vdd.n2864 vdd.n2863 39.2114
R17737 vdd.n2869 vdd.n2868 39.2114
R17738 vdd.n2862 vdd.n2860 39.2114
R17739 vdd.n2876 vdd.n2875 39.2114
R17740 vdd.n2859 vdd.n2857 39.2114
R17741 vdd.n2883 vdd.n2882 39.2114
R17742 vdd.n2856 vdd.n2854 39.2114
R17743 vdd.n2890 vdd.n2889 39.2114
R17744 vdd.n2028 vdd.n2027 39.2114
R17745 vdd.n2034 vdd.n2033 39.2114
R17746 vdd.n2035 vdd.n2024 39.2114
R17747 vdd.n2042 vdd.n2041 39.2114
R17748 vdd.n2043 vdd.n2022 39.2114
R17749 vdd.n2050 vdd.n2049 39.2114
R17750 vdd.n2051 vdd.n2020 39.2114
R17751 vdd.n2058 vdd.n2057 39.2114
R17752 vdd.n2229 vdd.n2228 39.2114
R17753 vdd.n2226 vdd.n2225 39.2114
R17754 vdd.n2221 vdd.n2220 39.2114
R17755 vdd.n2218 vdd.n2217 39.2114
R17756 vdd.n2213 vdd.n2212 39.2114
R17757 vdd.n2210 vdd.n2209 39.2114
R17758 vdd.n2205 vdd.n2204 39.2114
R17759 vdd.n2202 vdd.n2201 39.2114
R17760 vdd.n2197 vdd.n2196 39.2114
R17761 vdd.n2454 vdd.n908 39.2114
R17762 vdd.n2459 vdd.n909 39.2114
R17763 vdd.n2463 vdd.n910 39.2114
R17764 vdd.n2467 vdd.n911 39.2114
R17765 vdd.n2471 vdd.n912 39.2114
R17766 vdd.n2475 vdd.n913 39.2114
R17767 vdd.n2479 vdd.n914 39.2114
R17768 vdd.n2483 vdd.n915 39.2114
R17769 vdd.n2487 vdd.n916 39.2114
R17770 vdd.n2491 vdd.n917 39.2114
R17771 vdd.n2495 vdd.n918 39.2114
R17772 vdd.n2499 vdd.n919 39.2114
R17773 vdd.n2503 vdd.n920 39.2114
R17774 vdd.n2507 vdd.n921 39.2114
R17775 vdd.n2511 vdd.n922 39.2114
R17776 vdd.n2515 vdd.n923 39.2114
R17777 vdd.n926 vdd.n924 39.2114
R17778 vdd.n2773 vdd.n2772 39.2114
R17779 vdd.n2766 vdd.n2522 39.2114
R17780 vdd.n2762 vdd.n2523 39.2114
R17781 vdd.n2758 vdd.n2524 39.2114
R17782 vdd.n2754 vdd.n2525 39.2114
R17783 vdd.n2750 vdd.n2526 39.2114
R17784 vdd.n2746 vdd.n2527 39.2114
R17785 vdd.n2742 vdd.n2528 39.2114
R17786 vdd.n2738 vdd.n2529 39.2114
R17787 vdd.n2734 vdd.n2530 39.2114
R17788 vdd.n2730 vdd.n2531 39.2114
R17789 vdd.n2726 vdd.n2532 39.2114
R17790 vdd.n2722 vdd.n2533 39.2114
R17791 vdd.n2718 vdd.n2534 39.2114
R17792 vdd.n2714 vdd.n2535 39.2114
R17793 vdd.n2709 vdd.n2536 39.2114
R17794 vdd.n2705 vdd.n2537 39.2114
R17795 vdd.n2911 vdd.n803 39.2114
R17796 vdd.n2918 vdd.n2917 39.2114
R17797 vdd.n802 vdd.n800 39.2114
R17798 vdd.n2925 vdd.n2924 39.2114
R17799 vdd.n799 vdd.n797 39.2114
R17800 vdd.n2932 vdd.n2931 39.2114
R17801 vdd.n796 vdd.n794 39.2114
R17802 vdd.n2939 vdd.n2938 39.2114
R17803 vdd.n793 vdd.n791 39.2114
R17804 vdd.n2947 vdd.n2946 39.2114
R17805 vdd.n790 vdd.n788 39.2114
R17806 vdd.n2954 vdd.n2953 39.2114
R17807 vdd.n787 vdd.n785 39.2114
R17808 vdd.n2961 vdd.n2960 39.2114
R17809 vdd.n784 vdd.n782 39.2114
R17810 vdd.n2968 vdd.n2967 39.2114
R17811 vdd.n2971 vdd.n2970 39.2114
R17812 vdd.n934 vdd.n890 39.2114
R17813 vdd.n2443 vdd.n891 39.2114
R17814 vdd.n2439 vdd.n892 39.2114
R17815 vdd.n2435 vdd.n893 39.2114
R17816 vdd.n2431 vdd.n894 39.2114
R17817 vdd.n2427 vdd.n895 39.2114
R17818 vdd.n2423 vdd.n896 39.2114
R17819 vdd.n2419 vdd.n897 39.2114
R17820 vdd.n2415 vdd.n898 39.2114
R17821 vdd.n2411 vdd.n899 39.2114
R17822 vdd.n2407 vdd.n900 39.2114
R17823 vdd.n2403 vdd.n901 39.2114
R17824 vdd.n2399 vdd.n902 39.2114
R17825 vdd.n2395 vdd.n903 39.2114
R17826 vdd.n2391 vdd.n904 39.2114
R17827 vdd.n2387 vdd.n905 39.2114
R17828 vdd.n2383 vdd.n906 39.2114
R17829 vdd.n2286 vdd.n1023 39.2114
R17830 vdd.n2285 vdd.n2284 39.2114
R17831 vdd.n2278 vdd.n1025 39.2114
R17832 vdd.n2277 vdd.n2276 39.2114
R17833 vdd.n2270 vdd.n1027 39.2114
R17834 vdd.n2269 vdd.n2268 39.2114
R17835 vdd.n2262 vdd.n1029 39.2114
R17836 vdd.n2261 vdd.n2260 39.2114
R17837 vdd.n1032 vdd.n1031 39.2114
R17838 vdd.n2102 vdd.n2101 39.2114
R17839 vdd.n2107 vdd.n2106 39.2114
R17840 vdd.n2110 vdd.n2109 39.2114
R17841 vdd.n2115 vdd.n2114 39.2114
R17842 vdd.n2118 vdd.n2117 39.2114
R17843 vdd.n2123 vdd.n2122 39.2114
R17844 vdd.n2126 vdd.n2125 39.2114
R17845 vdd.n2132 vdd.n2131 39.2114
R17846 vdd.n2380 vdd.n906 39.2114
R17847 vdd.n2384 vdd.n905 39.2114
R17848 vdd.n2388 vdd.n904 39.2114
R17849 vdd.n2392 vdd.n903 39.2114
R17850 vdd.n2396 vdd.n902 39.2114
R17851 vdd.n2400 vdd.n901 39.2114
R17852 vdd.n2404 vdd.n900 39.2114
R17853 vdd.n2408 vdd.n899 39.2114
R17854 vdd.n2412 vdd.n898 39.2114
R17855 vdd.n2416 vdd.n897 39.2114
R17856 vdd.n2420 vdd.n896 39.2114
R17857 vdd.n2424 vdd.n895 39.2114
R17858 vdd.n2428 vdd.n894 39.2114
R17859 vdd.n2432 vdd.n893 39.2114
R17860 vdd.n2436 vdd.n892 39.2114
R17861 vdd.n2440 vdd.n891 39.2114
R17862 vdd.n2444 vdd.n890 39.2114
R17863 vdd.n2287 vdd.n2286 39.2114
R17864 vdd.n2284 vdd.n2283 39.2114
R17865 vdd.n2279 vdd.n2278 39.2114
R17866 vdd.n2276 vdd.n2275 39.2114
R17867 vdd.n2271 vdd.n2270 39.2114
R17868 vdd.n2268 vdd.n2267 39.2114
R17869 vdd.n2263 vdd.n2262 39.2114
R17870 vdd.n2260 vdd.n2259 39.2114
R17871 vdd.n1033 vdd.n1032 39.2114
R17872 vdd.n2103 vdd.n2102 39.2114
R17873 vdd.n2108 vdd.n2107 39.2114
R17874 vdd.n2109 vdd.n2099 39.2114
R17875 vdd.n2116 vdd.n2115 39.2114
R17876 vdd.n2117 vdd.n2097 39.2114
R17877 vdd.n2124 vdd.n2123 39.2114
R17878 vdd.n2125 vdd.n2093 39.2114
R17879 vdd.n2133 vdd.n2132 39.2114
R17880 vdd.n2252 vdd.n2251 37.2369
R17881 vdd.n1955 vdd.n1888 37.2369
R17882 vdd.n1994 vdd.n1848 37.2369
R17883 vdd.n3059 vdd.n724 37.2369
R17884 vdd.n688 vdd.n687 37.2369
R17885 vdd.n3015 vdd.n3014 37.2369
R17886 vdd.n2294 vdd.n1018 31.6883
R17887 vdd.n2519 vdd.n927 31.6883
R17888 vdd.n2452 vdd.n930 31.6883
R17889 vdd.n2198 vdd.n2195 31.6883
R17890 vdd.n2706 vdd.n2704 31.6883
R17891 vdd.n2913 vdd.n2910 31.6883
R17892 vdd.n2783 vdd.n883 31.6883
R17893 vdd.n2974 vdd.n2973 31.6883
R17894 vdd.n2893 vdd.n2892 31.6883
R17895 vdd.n2979 vdd.n771 31.6883
R17896 vdd.n2625 vdd.n2624 31.6883
R17897 vdd.n2779 vdd.n2778 31.6883
R17898 vdd.n2290 vdd.n2289 31.6883
R17899 vdd.n2447 vdd.n2446 31.6883
R17900 vdd.n2379 vdd.n2378 31.6883
R17901 vdd.n2136 vdd.n2135 31.6883
R17902 vdd.n2129 vdd.n2095 30.449
R17903 vdd.n938 vdd.n937 30.449
R17904 vdd.n2070 vdd.n2069 30.449
R17905 vdd.n2457 vdd.n929 30.449
R17906 vdd.n2561 vdd.n2560 30.449
R17907 vdd.n806 vdd.n805 30.449
R17908 vdd.n2711 vdd.n2557 30.449
R17909 vdd.n770 vdd.n769 30.449
R17910 vdd.n1380 vdd.n1146 19.3944
R17911 vdd.n1380 vdd.n1136 19.3944
R17912 vdd.n1392 vdd.n1136 19.3944
R17913 vdd.n1392 vdd.n1134 19.3944
R17914 vdd.n1396 vdd.n1134 19.3944
R17915 vdd.n1396 vdd.n1124 19.3944
R17916 vdd.n1409 vdd.n1124 19.3944
R17917 vdd.n1409 vdd.n1122 19.3944
R17918 vdd.n1413 vdd.n1122 19.3944
R17919 vdd.n1413 vdd.n1114 19.3944
R17920 vdd.n1426 vdd.n1114 19.3944
R17921 vdd.n1426 vdd.n1112 19.3944
R17922 vdd.n1430 vdd.n1112 19.3944
R17923 vdd.n1430 vdd.n1101 19.3944
R17924 vdd.n1442 vdd.n1101 19.3944
R17925 vdd.n1442 vdd.n1099 19.3944
R17926 vdd.n1446 vdd.n1099 19.3944
R17927 vdd.n1446 vdd.n1090 19.3944
R17928 vdd.n1754 vdd.n1090 19.3944
R17929 vdd.n1754 vdd.n1088 19.3944
R17930 vdd.n1758 vdd.n1088 19.3944
R17931 vdd.n1758 vdd.n1079 19.3944
R17932 vdd.n1770 vdd.n1079 19.3944
R17933 vdd.n1770 vdd.n1077 19.3944
R17934 vdd.n1774 vdd.n1077 19.3944
R17935 vdd.n1774 vdd.n1067 19.3944
R17936 vdd.n1787 vdd.n1067 19.3944
R17937 vdd.n1787 vdd.n1065 19.3944
R17938 vdd.n1791 vdd.n1065 19.3944
R17939 vdd.n1791 vdd.n1057 19.3944
R17940 vdd.n1804 vdd.n1057 19.3944
R17941 vdd.n1804 vdd.n1054 19.3944
R17942 vdd.n1810 vdd.n1054 19.3944
R17943 vdd.n1810 vdd.n1055 19.3944
R17944 vdd.n1055 vdd.n1043 19.3944
R17945 vdd.n1299 vdd.n1241 19.3944
R17946 vdd.n1299 vdd.n1298 19.3944
R17947 vdd.n1298 vdd.n1297 19.3944
R17948 vdd.n1297 vdd.n1247 19.3944
R17949 vdd.n1293 vdd.n1247 19.3944
R17950 vdd.n1293 vdd.n1292 19.3944
R17951 vdd.n1292 vdd.n1291 19.3944
R17952 vdd.n1291 vdd.n1253 19.3944
R17953 vdd.n1287 vdd.n1253 19.3944
R17954 vdd.n1287 vdd.n1286 19.3944
R17955 vdd.n1286 vdd.n1285 19.3944
R17956 vdd.n1285 vdd.n1259 19.3944
R17957 vdd.n1281 vdd.n1259 19.3944
R17958 vdd.n1281 vdd.n1280 19.3944
R17959 vdd.n1280 vdd.n1279 19.3944
R17960 vdd.n1279 vdd.n1265 19.3944
R17961 vdd.n1275 vdd.n1265 19.3944
R17962 vdd.n1275 vdd.n1274 19.3944
R17963 vdd.n1274 vdd.n1273 19.3944
R17964 vdd.n1273 vdd.n1271 19.3944
R17965 vdd.n1337 vdd.n1336 19.3944
R17966 vdd.n1336 vdd.n1212 19.3944
R17967 vdd.n1332 vdd.n1212 19.3944
R17968 vdd.n1332 vdd.n1331 19.3944
R17969 vdd.n1331 vdd.n1330 19.3944
R17970 vdd.n1330 vdd.n1218 19.3944
R17971 vdd.n1326 vdd.n1218 19.3944
R17972 vdd.n1326 vdd.n1325 19.3944
R17973 vdd.n1325 vdd.n1324 19.3944
R17974 vdd.n1324 vdd.n1224 19.3944
R17975 vdd.n1320 vdd.n1224 19.3944
R17976 vdd.n1320 vdd.n1319 19.3944
R17977 vdd.n1319 vdd.n1318 19.3944
R17978 vdd.n1318 vdd.n1230 19.3944
R17979 vdd.n1314 vdd.n1230 19.3944
R17980 vdd.n1314 vdd.n1313 19.3944
R17981 vdd.n1313 vdd.n1312 19.3944
R17982 vdd.n1312 vdd.n1236 19.3944
R17983 vdd.n1308 vdd.n1236 19.3944
R17984 vdd.n1308 vdd.n1307 19.3944
R17985 vdd.n1371 vdd.n1370 19.3944
R17986 vdd.n1370 vdd.n1185 19.3944
R17987 vdd.n1366 vdd.n1185 19.3944
R17988 vdd.n1366 vdd.n1365 19.3944
R17989 vdd.n1365 vdd.n1364 19.3944
R17990 vdd.n1364 vdd.n1190 19.3944
R17991 vdd.n1360 vdd.n1190 19.3944
R17992 vdd.n1360 vdd.n1359 19.3944
R17993 vdd.n1359 vdd.n1358 19.3944
R17994 vdd.n1358 vdd.n1196 19.3944
R17995 vdd.n1354 vdd.n1196 19.3944
R17996 vdd.n1354 vdd.n1353 19.3944
R17997 vdd.n1353 vdd.n1352 19.3944
R17998 vdd.n1352 vdd.n1202 19.3944
R17999 vdd.n1348 vdd.n1202 19.3944
R18000 vdd.n1348 vdd.n1347 19.3944
R18001 vdd.n1347 vdd.n1346 19.3944
R18002 vdd.n1346 vdd.n1208 19.3944
R18003 vdd.n1951 vdd.n1886 19.3944
R18004 vdd.n1951 vdd.n1892 19.3944
R18005 vdd.n1946 vdd.n1892 19.3944
R18006 vdd.n1946 vdd.n1945 19.3944
R18007 vdd.n1945 vdd.n1944 19.3944
R18008 vdd.n1944 vdd.n1899 19.3944
R18009 vdd.n1939 vdd.n1899 19.3944
R18010 vdd.n1939 vdd.n1938 19.3944
R18011 vdd.n1938 vdd.n1937 19.3944
R18012 vdd.n1937 vdd.n1906 19.3944
R18013 vdd.n1932 vdd.n1906 19.3944
R18014 vdd.n1932 vdd.n1931 19.3944
R18015 vdd.n1931 vdd.n1930 19.3944
R18016 vdd.n1930 vdd.n1914 19.3944
R18017 vdd.n1925 vdd.n1914 19.3944
R18018 vdd.n1925 vdd.n1924 19.3944
R18019 vdd.n1920 vdd.n1919 19.3944
R18020 vdd.n2253 vdd.n1039 19.3944
R18021 vdd.n1990 vdd.n1846 19.3944
R18022 vdd.n1990 vdd.n1852 19.3944
R18023 vdd.n1985 vdd.n1852 19.3944
R18024 vdd.n1985 vdd.n1984 19.3944
R18025 vdd.n1984 vdd.n1983 19.3944
R18026 vdd.n1983 vdd.n1859 19.3944
R18027 vdd.n1978 vdd.n1859 19.3944
R18028 vdd.n1978 vdd.n1977 19.3944
R18029 vdd.n1977 vdd.n1976 19.3944
R18030 vdd.n1976 vdd.n1866 19.3944
R18031 vdd.n1971 vdd.n1866 19.3944
R18032 vdd.n1971 vdd.n1970 19.3944
R18033 vdd.n1970 vdd.n1969 19.3944
R18034 vdd.n1969 vdd.n1873 19.3944
R18035 vdd.n1964 vdd.n1873 19.3944
R18036 vdd.n1964 vdd.n1963 19.3944
R18037 vdd.n1963 vdd.n1962 19.3944
R18038 vdd.n1962 vdd.n1880 19.3944
R18039 vdd.n1957 vdd.n1880 19.3944
R18040 vdd.n1957 vdd.n1956 19.3944
R18041 vdd.n2241 vdd.n2240 19.3944
R18042 vdd.n2240 vdd.n1818 19.3944
R18043 vdd.n2235 vdd.n2234 19.3944
R18044 vdd.n2017 vdd.n1822 19.3944
R18045 vdd.n2017 vdd.n1824 19.3944
R18046 vdd.n1827 vdd.n1824 19.3944
R18047 vdd.n2010 vdd.n1827 19.3944
R18048 vdd.n2010 vdd.n2009 19.3944
R18049 vdd.n2009 vdd.n2008 19.3944
R18050 vdd.n2008 vdd.n1833 19.3944
R18051 vdd.n2003 vdd.n1833 19.3944
R18052 vdd.n2003 vdd.n2002 19.3944
R18053 vdd.n2002 vdd.n2001 19.3944
R18054 vdd.n2001 vdd.n1840 19.3944
R18055 vdd.n1996 vdd.n1840 19.3944
R18056 vdd.n1996 vdd.n1995 19.3944
R18057 vdd.n1384 vdd.n1142 19.3944
R18058 vdd.n1384 vdd.n1140 19.3944
R18059 vdd.n1388 vdd.n1140 19.3944
R18060 vdd.n1388 vdd.n1130 19.3944
R18061 vdd.n1401 vdd.n1130 19.3944
R18062 vdd.n1401 vdd.n1128 19.3944
R18063 vdd.n1405 vdd.n1128 19.3944
R18064 vdd.n1405 vdd.n1119 19.3944
R18065 vdd.n1418 vdd.n1119 19.3944
R18066 vdd.n1418 vdd.n1117 19.3944
R18067 vdd.n1422 vdd.n1117 19.3944
R18068 vdd.n1422 vdd.n1108 19.3944
R18069 vdd.n1434 vdd.n1108 19.3944
R18070 vdd.n1434 vdd.n1106 19.3944
R18071 vdd.n1438 vdd.n1106 19.3944
R18072 vdd.n1438 vdd.n1096 19.3944
R18073 vdd.n1451 vdd.n1096 19.3944
R18074 vdd.n1451 vdd.n1094 19.3944
R18075 vdd.n1750 vdd.n1094 19.3944
R18076 vdd.n1750 vdd.n1085 19.3944
R18077 vdd.n1762 vdd.n1085 19.3944
R18078 vdd.n1762 vdd.n1083 19.3944
R18079 vdd.n1766 vdd.n1083 19.3944
R18080 vdd.n1766 vdd.n1073 19.3944
R18081 vdd.n1779 vdd.n1073 19.3944
R18082 vdd.n1779 vdd.n1071 19.3944
R18083 vdd.n1783 vdd.n1071 19.3944
R18084 vdd.n1783 vdd.n1062 19.3944
R18085 vdd.n1796 vdd.n1062 19.3944
R18086 vdd.n1796 vdd.n1060 19.3944
R18087 vdd.n1800 vdd.n1060 19.3944
R18088 vdd.n1800 vdd.n1050 19.3944
R18089 vdd.n1814 vdd.n1050 19.3944
R18090 vdd.n1814 vdd.n1048 19.3944
R18091 vdd.n2244 vdd.n1048 19.3944
R18092 vdd.n3147 vdd.n655 19.3944
R18093 vdd.n3151 vdd.n655 19.3944
R18094 vdd.n3151 vdd.n646 19.3944
R18095 vdd.n3163 vdd.n646 19.3944
R18096 vdd.n3163 vdd.n644 19.3944
R18097 vdd.n3167 vdd.n644 19.3944
R18098 vdd.n3167 vdd.n633 19.3944
R18099 vdd.n3179 vdd.n633 19.3944
R18100 vdd.n3179 vdd.n631 19.3944
R18101 vdd.n3183 vdd.n631 19.3944
R18102 vdd.n3183 vdd.n622 19.3944
R18103 vdd.n3196 vdd.n622 19.3944
R18104 vdd.n3196 vdd.n620 19.3944
R18105 vdd.n3203 vdd.n620 19.3944
R18106 vdd.n3203 vdd.n3202 19.3944
R18107 vdd.n3202 vdd.n610 19.3944
R18108 vdd.n3216 vdd.n610 19.3944
R18109 vdd.n3217 vdd.n3216 19.3944
R18110 vdd.n3218 vdd.n3217 19.3944
R18111 vdd.n3218 vdd.n608 19.3944
R18112 vdd.n3223 vdd.n608 19.3944
R18113 vdd.n3224 vdd.n3223 19.3944
R18114 vdd.n3225 vdd.n3224 19.3944
R18115 vdd.n3225 vdd.n606 19.3944
R18116 vdd.n3230 vdd.n606 19.3944
R18117 vdd.n3231 vdd.n3230 19.3944
R18118 vdd.n3232 vdd.n3231 19.3944
R18119 vdd.n3232 vdd.n604 19.3944
R18120 vdd.n3238 vdd.n604 19.3944
R18121 vdd.n3239 vdd.n3238 19.3944
R18122 vdd.n3240 vdd.n3239 19.3944
R18123 vdd.n3240 vdd.n602 19.3944
R18124 vdd.n3245 vdd.n602 19.3944
R18125 vdd.n3246 vdd.n3245 19.3944
R18126 vdd.n3247 vdd.n3246 19.3944
R18127 vdd.n550 vdd.n417 19.3944
R18128 vdd.n556 vdd.n417 19.3944
R18129 vdd.n557 vdd.n556 19.3944
R18130 vdd.n560 vdd.n557 19.3944
R18131 vdd.n560 vdd.n415 19.3944
R18132 vdd.n566 vdd.n415 19.3944
R18133 vdd.n567 vdd.n566 19.3944
R18134 vdd.n570 vdd.n567 19.3944
R18135 vdd.n570 vdd.n413 19.3944
R18136 vdd.n576 vdd.n413 19.3944
R18137 vdd.n577 vdd.n576 19.3944
R18138 vdd.n580 vdd.n577 19.3944
R18139 vdd.n580 vdd.n411 19.3944
R18140 vdd.n586 vdd.n411 19.3944
R18141 vdd.n587 vdd.n586 19.3944
R18142 vdd.n590 vdd.n587 19.3944
R18143 vdd.n590 vdd.n409 19.3944
R18144 vdd.n596 vdd.n409 19.3944
R18145 vdd.n598 vdd.n596 19.3944
R18146 vdd.n599 vdd.n598 19.3944
R18147 vdd.n497 vdd.n496 19.3944
R18148 vdd.n500 vdd.n497 19.3944
R18149 vdd.n500 vdd.n429 19.3944
R18150 vdd.n506 vdd.n429 19.3944
R18151 vdd.n507 vdd.n506 19.3944
R18152 vdd.n510 vdd.n507 19.3944
R18153 vdd.n510 vdd.n427 19.3944
R18154 vdd.n516 vdd.n427 19.3944
R18155 vdd.n517 vdd.n516 19.3944
R18156 vdd.n520 vdd.n517 19.3944
R18157 vdd.n520 vdd.n425 19.3944
R18158 vdd.n526 vdd.n425 19.3944
R18159 vdd.n527 vdd.n526 19.3944
R18160 vdd.n530 vdd.n527 19.3944
R18161 vdd.n530 vdd.n423 19.3944
R18162 vdd.n536 vdd.n423 19.3944
R18163 vdd.n537 vdd.n536 19.3944
R18164 vdd.n540 vdd.n537 19.3944
R18165 vdd.n540 vdd.n421 19.3944
R18166 vdd.n546 vdd.n421 19.3944
R18167 vdd.n447 vdd.n446 19.3944
R18168 vdd.n450 vdd.n447 19.3944
R18169 vdd.n450 vdd.n441 19.3944
R18170 vdd.n456 vdd.n441 19.3944
R18171 vdd.n457 vdd.n456 19.3944
R18172 vdd.n460 vdd.n457 19.3944
R18173 vdd.n460 vdd.n439 19.3944
R18174 vdd.n466 vdd.n439 19.3944
R18175 vdd.n467 vdd.n466 19.3944
R18176 vdd.n470 vdd.n467 19.3944
R18177 vdd.n470 vdd.n437 19.3944
R18178 vdd.n476 vdd.n437 19.3944
R18179 vdd.n477 vdd.n476 19.3944
R18180 vdd.n480 vdd.n477 19.3944
R18181 vdd.n480 vdd.n435 19.3944
R18182 vdd.n486 vdd.n435 19.3944
R18183 vdd.n487 vdd.n486 19.3944
R18184 vdd.n490 vdd.n487 19.3944
R18185 vdd.n3143 vdd.n652 19.3944
R18186 vdd.n3155 vdd.n652 19.3944
R18187 vdd.n3155 vdd.n650 19.3944
R18188 vdd.n3159 vdd.n650 19.3944
R18189 vdd.n3159 vdd.n640 19.3944
R18190 vdd.n3171 vdd.n640 19.3944
R18191 vdd.n3171 vdd.n638 19.3944
R18192 vdd.n3175 vdd.n638 19.3944
R18193 vdd.n3175 vdd.n628 19.3944
R18194 vdd.n3188 vdd.n628 19.3944
R18195 vdd.n3188 vdd.n626 19.3944
R18196 vdd.n3192 vdd.n626 19.3944
R18197 vdd.n3192 vdd.n617 19.3944
R18198 vdd.n3207 vdd.n617 19.3944
R18199 vdd.n3207 vdd.n615 19.3944
R18200 vdd.n3211 vdd.n615 19.3944
R18201 vdd.n3211 vdd.n324 19.3944
R18202 vdd.n3289 vdd.n324 19.3944
R18203 vdd.n3289 vdd.n325 19.3944
R18204 vdd.n3283 vdd.n325 19.3944
R18205 vdd.n3283 vdd.n3282 19.3944
R18206 vdd.n3282 vdd.n3281 19.3944
R18207 vdd.n3281 vdd.n337 19.3944
R18208 vdd.n3275 vdd.n337 19.3944
R18209 vdd.n3275 vdd.n3274 19.3944
R18210 vdd.n3274 vdd.n3273 19.3944
R18211 vdd.n3273 vdd.n347 19.3944
R18212 vdd.n3267 vdd.n347 19.3944
R18213 vdd.n3267 vdd.n3266 19.3944
R18214 vdd.n3266 vdd.n3265 19.3944
R18215 vdd.n3265 vdd.n358 19.3944
R18216 vdd.n3259 vdd.n358 19.3944
R18217 vdd.n3259 vdd.n3258 19.3944
R18218 vdd.n3258 vdd.n3257 19.3944
R18219 vdd.n3257 vdd.n369 19.3944
R18220 vdd.n3100 vdd.n3099 19.3944
R18221 vdd.n3099 vdd.n3098 19.3944
R18222 vdd.n3098 vdd.n694 19.3944
R18223 vdd.n3092 vdd.n694 19.3944
R18224 vdd.n3092 vdd.n3091 19.3944
R18225 vdd.n3091 vdd.n3090 19.3944
R18226 vdd.n3090 vdd.n700 19.3944
R18227 vdd.n3084 vdd.n700 19.3944
R18228 vdd.n3084 vdd.n3083 19.3944
R18229 vdd.n3083 vdd.n3082 19.3944
R18230 vdd.n3082 vdd.n706 19.3944
R18231 vdd.n3076 vdd.n706 19.3944
R18232 vdd.n3076 vdd.n3075 19.3944
R18233 vdd.n3075 vdd.n3074 19.3944
R18234 vdd.n3074 vdd.n712 19.3944
R18235 vdd.n3068 vdd.n712 19.3944
R18236 vdd.n3068 vdd.n3067 19.3944
R18237 vdd.n3067 vdd.n3066 19.3944
R18238 vdd.n3066 vdd.n718 19.3944
R18239 vdd.n3060 vdd.n718 19.3944
R18240 vdd.n3140 vdd.n3139 19.3944
R18241 vdd.n3139 vdd.n662 19.3944
R18242 vdd.n3134 vdd.n3133 19.3944
R18243 vdd.n3130 vdd.n3129 19.3944
R18244 vdd.n3129 vdd.n668 19.3944
R18245 vdd.n3124 vdd.n668 19.3944
R18246 vdd.n3124 vdd.n3123 19.3944
R18247 vdd.n3123 vdd.n3122 19.3944
R18248 vdd.n3122 vdd.n674 19.3944
R18249 vdd.n3116 vdd.n674 19.3944
R18250 vdd.n3116 vdd.n3115 19.3944
R18251 vdd.n3115 vdd.n3114 19.3944
R18252 vdd.n3114 vdd.n680 19.3944
R18253 vdd.n3108 vdd.n680 19.3944
R18254 vdd.n3108 vdd.n3107 19.3944
R18255 vdd.n3107 vdd.n3106 19.3944
R18256 vdd.n3055 vdd.n722 19.3944
R18257 vdd.n3055 vdd.n726 19.3944
R18258 vdd.n3050 vdd.n726 19.3944
R18259 vdd.n3050 vdd.n3049 19.3944
R18260 vdd.n3049 vdd.n732 19.3944
R18261 vdd.n3044 vdd.n732 19.3944
R18262 vdd.n3044 vdd.n3043 19.3944
R18263 vdd.n3043 vdd.n3042 19.3944
R18264 vdd.n3042 vdd.n738 19.3944
R18265 vdd.n3036 vdd.n738 19.3944
R18266 vdd.n3036 vdd.n3035 19.3944
R18267 vdd.n3035 vdd.n3034 19.3944
R18268 vdd.n3034 vdd.n744 19.3944
R18269 vdd.n3028 vdd.n744 19.3944
R18270 vdd.n3028 vdd.n3027 19.3944
R18271 vdd.n3027 vdd.n3026 19.3944
R18272 vdd.n3022 vdd.n3021 19.3944
R18273 vdd.n3018 vdd.n3017 19.3944
R18274 vdd.n1306 vdd.n1241 19.0066
R18275 vdd.n1955 vdd.n1886 19.0066
R18276 vdd.n550 vdd.n547 19.0066
R18277 vdd.n3059 vdd.n722 19.0066
R18278 vdd.n1374 vdd.n1144 18.5924
R18279 vdd.n2246 vdd.n1045 18.5924
R18280 vdd.n3145 vdd.n658 18.5924
R18281 vdd.n3254 vdd.n3253 18.5924
R18282 vdd.n2095 vdd.n2094 16.0975
R18283 vdd.n937 vdd.n936 16.0975
R18284 vdd.n1149 vdd.n1148 16.0975
R18285 vdd.n1305 vdd.n1304 16.0975
R18286 vdd.n1341 vdd.n1340 16.0975
R18287 vdd.n2251 vdd.n2250 16.0975
R18288 vdd.n1888 vdd.n1887 16.0975
R18289 vdd.n1848 vdd.n1847 16.0975
R18290 vdd.n2069 vdd.n2068 16.0975
R18291 vdd.n929 vdd.n928 16.0975
R18292 vdd.n2560 vdd.n2559 16.0975
R18293 vdd.n406 vdd.n405 16.0975
R18294 vdd.n420 vdd.n419 16.0975
R18295 vdd.n432 vdd.n431 16.0975
R18296 vdd.n724 vdd.n723 16.0975
R18297 vdd.n687 vdd.n686 16.0975
R18298 vdd.n805 vdd.n804 16.0975
R18299 vdd.n2557 vdd.n2556 16.0975
R18300 vdd.n3014 vdd.n3013 16.0975
R18301 vdd.n769 vdd.n768 16.0975
R18302 vdd.t13 vdd.n2521 15.4182
R18303 vdd.n2774 vdd.t262 15.4182
R18304 vdd.n28 vdd.n27 15.0023
R18305 vdd.n2292 vdd.n1020 14.5112
R18306 vdd.n2976 vdd.n756 14.5112
R18307 vdd.n316 vdd.n281 13.1884
R18308 vdd.n261 vdd.n226 13.1884
R18309 vdd.n218 vdd.n183 13.1884
R18310 vdd.n163 vdd.n128 13.1884
R18311 vdd.n121 vdd.n86 13.1884
R18312 vdd.n66 vdd.n31 13.1884
R18313 vdd.n1685 vdd.n1650 13.1884
R18314 vdd.n1740 vdd.n1705 13.1884
R18315 vdd.n1587 vdd.n1552 13.1884
R18316 vdd.n1642 vdd.n1607 13.1884
R18317 vdd.n1490 vdd.n1455 13.1884
R18318 vdd.n1545 vdd.n1510 13.1884
R18319 vdd.n1342 vdd.n1337 12.9944
R18320 vdd.n1342 vdd.n1208 12.9944
R18321 vdd.n1994 vdd.n1846 12.9944
R18322 vdd.n1995 vdd.n1994 12.9944
R18323 vdd.n496 vdd.n433 12.9944
R18324 vdd.n490 vdd.n433 12.9944
R18325 vdd.n3100 vdd.n688 12.9944
R18326 vdd.n3106 vdd.n688 12.9944
R18327 vdd.n317 vdd.n279 12.8005
R18328 vdd.n312 vdd.n283 12.8005
R18329 vdd.n262 vdd.n224 12.8005
R18330 vdd.n257 vdd.n228 12.8005
R18331 vdd.n219 vdd.n181 12.8005
R18332 vdd.n214 vdd.n185 12.8005
R18333 vdd.n164 vdd.n126 12.8005
R18334 vdd.n159 vdd.n130 12.8005
R18335 vdd.n122 vdd.n84 12.8005
R18336 vdd.n117 vdd.n88 12.8005
R18337 vdd.n67 vdd.n29 12.8005
R18338 vdd.n62 vdd.n33 12.8005
R18339 vdd.n1686 vdd.n1648 12.8005
R18340 vdd.n1681 vdd.n1652 12.8005
R18341 vdd.n1741 vdd.n1703 12.8005
R18342 vdd.n1736 vdd.n1707 12.8005
R18343 vdd.n1588 vdd.n1550 12.8005
R18344 vdd.n1583 vdd.n1554 12.8005
R18345 vdd.n1643 vdd.n1605 12.8005
R18346 vdd.n1638 vdd.n1609 12.8005
R18347 vdd.n1491 vdd.n1453 12.8005
R18348 vdd.n1486 vdd.n1457 12.8005
R18349 vdd.n1546 vdd.n1508 12.8005
R18350 vdd.n1541 vdd.n1512 12.8005
R18351 vdd.n311 vdd.n284 12.0247
R18352 vdd.n256 vdd.n229 12.0247
R18353 vdd.n213 vdd.n186 12.0247
R18354 vdd.n158 vdd.n131 12.0247
R18355 vdd.n116 vdd.n89 12.0247
R18356 vdd.n61 vdd.n34 12.0247
R18357 vdd.n1680 vdd.n1653 12.0247
R18358 vdd.n1735 vdd.n1708 12.0247
R18359 vdd.n1582 vdd.n1555 12.0247
R18360 vdd.n1637 vdd.n1610 12.0247
R18361 vdd.n1485 vdd.n1458 12.0247
R18362 vdd.n1540 vdd.n1513 12.0247
R18363 vdd.n1382 vdd.n1144 11.337
R18364 vdd.n1390 vdd.n1138 11.337
R18365 vdd.n1390 vdd.n1132 11.337
R18366 vdd.n1399 vdd.n1132 11.337
R18367 vdd.n1407 vdd.n1126 11.337
R18368 vdd.n1416 vdd.n1415 11.337
R18369 vdd.n1432 vdd.n1110 11.337
R18370 vdd.n1440 vdd.n1103 11.337
R18371 vdd.n1449 vdd.n1448 11.337
R18372 vdd.n1752 vdd.n1092 11.337
R18373 vdd.n1768 vdd.n1081 11.337
R18374 vdd.n1777 vdd.n1075 11.337
R18375 vdd.n1785 vdd.n1069 11.337
R18376 vdd.n1794 vdd.n1793 11.337
R18377 vdd.n1802 vdd.n1052 11.337
R18378 vdd.n1812 vdd.n1052 11.337
R18379 vdd.n2246 vdd.n1044 11.337
R18380 vdd.n3145 vdd.n659 11.337
R18381 vdd.n3153 vdd.n648 11.337
R18382 vdd.n3161 vdd.n648 11.337
R18383 vdd.n3169 vdd.n642 11.337
R18384 vdd.n3177 vdd.n635 11.337
R18385 vdd.n3186 vdd.n3185 11.337
R18386 vdd.n3194 vdd.n624 11.337
R18387 vdd.n3213 vdd.n613 11.337
R18388 vdd.n3287 vdd.n328 11.337
R18389 vdd.n3285 vdd.n332 11.337
R18390 vdd.n3279 vdd.n3278 11.337
R18391 vdd.n3271 vdd.n349 11.337
R18392 vdd.n3270 vdd.n3269 11.337
R18393 vdd.n3263 vdd.n3262 11.337
R18394 vdd.n3262 vdd.n3261 11.337
R18395 vdd.n3261 vdd.n363 11.337
R18396 vdd.n3255 vdd.n3254 11.337
R18397 vdd.n308 vdd.n307 11.249
R18398 vdd.n253 vdd.n252 11.249
R18399 vdd.n210 vdd.n209 11.249
R18400 vdd.n155 vdd.n154 11.249
R18401 vdd.n113 vdd.n112 11.249
R18402 vdd.n58 vdd.n57 11.249
R18403 vdd.n1677 vdd.n1676 11.249
R18404 vdd.n1732 vdd.n1731 11.249
R18405 vdd.n1579 vdd.n1578 11.249
R18406 vdd.n1634 vdd.n1633 11.249
R18407 vdd.n1482 vdd.n1481 11.249
R18408 vdd.n1537 vdd.n1536 11.249
R18409 vdd.n2449 vdd.t109 11.1103
R18410 vdd.n2781 vdd.t106 11.1103
R18411 vdd.n1802 vdd.t136 10.7702
R18412 vdd.n3161 vdd.t134 10.7702
R18413 vdd.n293 vdd.n292 10.7238
R18414 vdd.n238 vdd.n237 10.7238
R18415 vdd.n195 vdd.n194 10.7238
R18416 vdd.n140 vdd.n139 10.7238
R18417 vdd.n98 vdd.n97 10.7238
R18418 vdd.n43 vdd.n42 10.7238
R18419 vdd.n1662 vdd.n1661 10.7238
R18420 vdd.n1717 vdd.n1716 10.7238
R18421 vdd.n1564 vdd.n1563 10.7238
R18422 vdd.n1619 vdd.n1618 10.7238
R18423 vdd.n1467 vdd.n1466 10.7238
R18424 vdd.n1522 vdd.n1521 10.7238
R18425 vdd.n2295 vdd.n2294 10.6151
R18426 vdd.n2296 vdd.n2295 10.6151
R18427 vdd.n2296 vdd.n1006 10.6151
R18428 vdd.n2306 vdd.n1006 10.6151
R18429 vdd.n2307 vdd.n2306 10.6151
R18430 vdd.n2308 vdd.n2307 10.6151
R18431 vdd.n2308 vdd.n993 10.6151
R18432 vdd.n2319 vdd.n993 10.6151
R18433 vdd.n2320 vdd.n2319 10.6151
R18434 vdd.n2321 vdd.n2320 10.6151
R18435 vdd.n2321 vdd.n981 10.6151
R18436 vdd.n2331 vdd.n981 10.6151
R18437 vdd.n2332 vdd.n2331 10.6151
R18438 vdd.n2333 vdd.n2332 10.6151
R18439 vdd.n2333 vdd.n969 10.6151
R18440 vdd.n2343 vdd.n969 10.6151
R18441 vdd.n2344 vdd.n2343 10.6151
R18442 vdd.n2345 vdd.n2344 10.6151
R18443 vdd.n2345 vdd.n958 10.6151
R18444 vdd.n2355 vdd.n958 10.6151
R18445 vdd.n2356 vdd.n2355 10.6151
R18446 vdd.n2357 vdd.n2356 10.6151
R18447 vdd.n2357 vdd.n945 10.6151
R18448 vdd.n2369 vdd.n945 10.6151
R18449 vdd.n2370 vdd.n2369 10.6151
R18450 vdd.n2372 vdd.n2370 10.6151
R18451 vdd.n2372 vdd.n2371 10.6151
R18452 vdd.n2371 vdd.n927 10.6151
R18453 vdd.n2519 vdd.n2518 10.6151
R18454 vdd.n2518 vdd.n2517 10.6151
R18455 vdd.n2517 vdd.n2514 10.6151
R18456 vdd.n2514 vdd.n2513 10.6151
R18457 vdd.n2513 vdd.n2510 10.6151
R18458 vdd.n2510 vdd.n2509 10.6151
R18459 vdd.n2509 vdd.n2506 10.6151
R18460 vdd.n2506 vdd.n2505 10.6151
R18461 vdd.n2505 vdd.n2502 10.6151
R18462 vdd.n2502 vdd.n2501 10.6151
R18463 vdd.n2501 vdd.n2498 10.6151
R18464 vdd.n2498 vdd.n2497 10.6151
R18465 vdd.n2497 vdd.n2494 10.6151
R18466 vdd.n2494 vdd.n2493 10.6151
R18467 vdd.n2493 vdd.n2490 10.6151
R18468 vdd.n2490 vdd.n2489 10.6151
R18469 vdd.n2489 vdd.n2486 10.6151
R18470 vdd.n2486 vdd.n2485 10.6151
R18471 vdd.n2485 vdd.n2482 10.6151
R18472 vdd.n2482 vdd.n2481 10.6151
R18473 vdd.n2481 vdd.n2478 10.6151
R18474 vdd.n2478 vdd.n2477 10.6151
R18475 vdd.n2477 vdd.n2474 10.6151
R18476 vdd.n2474 vdd.n2473 10.6151
R18477 vdd.n2473 vdd.n2470 10.6151
R18478 vdd.n2470 vdd.n2469 10.6151
R18479 vdd.n2469 vdd.n2466 10.6151
R18480 vdd.n2466 vdd.n2465 10.6151
R18481 vdd.n2465 vdd.n2462 10.6151
R18482 vdd.n2462 vdd.n2461 10.6151
R18483 vdd.n2461 vdd.n2458 10.6151
R18484 vdd.n2456 vdd.n2453 10.6151
R18485 vdd.n2453 vdd.n2452 10.6151
R18486 vdd.n2195 vdd.n2194 10.6151
R18487 vdd.n2194 vdd.n2192 10.6151
R18488 vdd.n2192 vdd.n2191 10.6151
R18489 vdd.n2191 vdd.n2189 10.6151
R18490 vdd.n2189 vdd.n2188 10.6151
R18491 vdd.n2188 vdd.n2186 10.6151
R18492 vdd.n2186 vdd.n2185 10.6151
R18493 vdd.n2185 vdd.n2183 10.6151
R18494 vdd.n2183 vdd.n2182 10.6151
R18495 vdd.n2182 vdd.n2180 10.6151
R18496 vdd.n2180 vdd.n2179 10.6151
R18497 vdd.n2179 vdd.n2177 10.6151
R18498 vdd.n2177 vdd.n2176 10.6151
R18499 vdd.n2176 vdd.n2091 10.6151
R18500 vdd.n2091 vdd.n2090 10.6151
R18501 vdd.n2090 vdd.n2088 10.6151
R18502 vdd.n2088 vdd.n2087 10.6151
R18503 vdd.n2087 vdd.n2085 10.6151
R18504 vdd.n2085 vdd.n2084 10.6151
R18505 vdd.n2084 vdd.n2082 10.6151
R18506 vdd.n2082 vdd.n2081 10.6151
R18507 vdd.n2081 vdd.n2079 10.6151
R18508 vdd.n2079 vdd.n2078 10.6151
R18509 vdd.n2078 vdd.n2076 10.6151
R18510 vdd.n2076 vdd.n2075 10.6151
R18511 vdd.n2075 vdd.n2072 10.6151
R18512 vdd.n2072 vdd.n2071 10.6151
R18513 vdd.n2071 vdd.n930 10.6151
R18514 vdd.n2029 vdd.n1018 10.6151
R18515 vdd.n2030 vdd.n2029 10.6151
R18516 vdd.n2031 vdd.n2030 10.6151
R18517 vdd.n2031 vdd.n2025 10.6151
R18518 vdd.n2037 vdd.n2025 10.6151
R18519 vdd.n2038 vdd.n2037 10.6151
R18520 vdd.n2039 vdd.n2038 10.6151
R18521 vdd.n2039 vdd.n2023 10.6151
R18522 vdd.n2045 vdd.n2023 10.6151
R18523 vdd.n2046 vdd.n2045 10.6151
R18524 vdd.n2047 vdd.n2046 10.6151
R18525 vdd.n2047 vdd.n2021 10.6151
R18526 vdd.n2053 vdd.n2021 10.6151
R18527 vdd.n2054 vdd.n2053 10.6151
R18528 vdd.n2055 vdd.n2054 10.6151
R18529 vdd.n2055 vdd.n2019 10.6151
R18530 vdd.n2231 vdd.n2019 10.6151
R18531 vdd.n2231 vdd.n2230 10.6151
R18532 vdd.n2230 vdd.n2060 10.6151
R18533 vdd.n2224 vdd.n2060 10.6151
R18534 vdd.n2224 vdd.n2223 10.6151
R18535 vdd.n2223 vdd.n2222 10.6151
R18536 vdd.n2222 vdd.n2062 10.6151
R18537 vdd.n2216 vdd.n2062 10.6151
R18538 vdd.n2216 vdd.n2215 10.6151
R18539 vdd.n2215 vdd.n2214 10.6151
R18540 vdd.n2214 vdd.n2064 10.6151
R18541 vdd.n2208 vdd.n2064 10.6151
R18542 vdd.n2208 vdd.n2207 10.6151
R18543 vdd.n2207 vdd.n2206 10.6151
R18544 vdd.n2206 vdd.n2066 10.6151
R18545 vdd.n2200 vdd.n2199 10.6151
R18546 vdd.n2199 vdd.n2198 10.6151
R18547 vdd.n2704 vdd.n2703 10.6151
R18548 vdd.n2703 vdd.n2701 10.6151
R18549 vdd.n2701 vdd.n2700 10.6151
R18550 vdd.n2700 vdd.n2558 10.6151
R18551 vdd.n2647 vdd.n2558 10.6151
R18552 vdd.n2648 vdd.n2647 10.6151
R18553 vdd.n2650 vdd.n2648 10.6151
R18554 vdd.n2651 vdd.n2650 10.6151
R18555 vdd.n2653 vdd.n2651 10.6151
R18556 vdd.n2654 vdd.n2653 10.6151
R18557 vdd.n2656 vdd.n2654 10.6151
R18558 vdd.n2657 vdd.n2656 10.6151
R18559 vdd.n2659 vdd.n2657 10.6151
R18560 vdd.n2660 vdd.n2659 10.6151
R18561 vdd.n2675 vdd.n2660 10.6151
R18562 vdd.n2675 vdd.n2674 10.6151
R18563 vdd.n2674 vdd.n2673 10.6151
R18564 vdd.n2673 vdd.n2671 10.6151
R18565 vdd.n2671 vdd.n2670 10.6151
R18566 vdd.n2670 vdd.n2668 10.6151
R18567 vdd.n2668 vdd.n2667 10.6151
R18568 vdd.n2667 vdd.n2665 10.6151
R18569 vdd.n2665 vdd.n2664 10.6151
R18570 vdd.n2664 vdd.n2662 10.6151
R18571 vdd.n2662 vdd.n2661 10.6151
R18572 vdd.n2661 vdd.n807 10.6151
R18573 vdd.n2909 vdd.n807 10.6151
R18574 vdd.n2910 vdd.n2909 10.6151
R18575 vdd.n2771 vdd.n883 10.6151
R18576 vdd.n2771 vdd.n2770 10.6151
R18577 vdd.n2770 vdd.n2769 10.6151
R18578 vdd.n2769 vdd.n2767 10.6151
R18579 vdd.n2767 vdd.n2764 10.6151
R18580 vdd.n2764 vdd.n2763 10.6151
R18581 vdd.n2763 vdd.n2760 10.6151
R18582 vdd.n2760 vdd.n2759 10.6151
R18583 vdd.n2759 vdd.n2756 10.6151
R18584 vdd.n2756 vdd.n2755 10.6151
R18585 vdd.n2755 vdd.n2752 10.6151
R18586 vdd.n2752 vdd.n2751 10.6151
R18587 vdd.n2751 vdd.n2748 10.6151
R18588 vdd.n2748 vdd.n2747 10.6151
R18589 vdd.n2747 vdd.n2744 10.6151
R18590 vdd.n2744 vdd.n2743 10.6151
R18591 vdd.n2743 vdd.n2740 10.6151
R18592 vdd.n2740 vdd.n2739 10.6151
R18593 vdd.n2739 vdd.n2736 10.6151
R18594 vdd.n2736 vdd.n2735 10.6151
R18595 vdd.n2735 vdd.n2732 10.6151
R18596 vdd.n2732 vdd.n2731 10.6151
R18597 vdd.n2731 vdd.n2728 10.6151
R18598 vdd.n2728 vdd.n2727 10.6151
R18599 vdd.n2727 vdd.n2724 10.6151
R18600 vdd.n2724 vdd.n2723 10.6151
R18601 vdd.n2723 vdd.n2720 10.6151
R18602 vdd.n2720 vdd.n2719 10.6151
R18603 vdd.n2719 vdd.n2716 10.6151
R18604 vdd.n2716 vdd.n2715 10.6151
R18605 vdd.n2715 vdd.n2712 10.6151
R18606 vdd.n2710 vdd.n2707 10.6151
R18607 vdd.n2707 vdd.n2706 10.6151
R18608 vdd.n2784 vdd.n2783 10.6151
R18609 vdd.n2785 vdd.n2784 10.6151
R18610 vdd.n2785 vdd.n873 10.6151
R18611 vdd.n2795 vdd.n873 10.6151
R18612 vdd.n2796 vdd.n2795 10.6151
R18613 vdd.n2797 vdd.n2796 10.6151
R18614 vdd.n2797 vdd.n860 10.6151
R18615 vdd.n2807 vdd.n860 10.6151
R18616 vdd.n2808 vdd.n2807 10.6151
R18617 vdd.n2809 vdd.n2808 10.6151
R18618 vdd.n2809 vdd.n849 10.6151
R18619 vdd.n2819 vdd.n849 10.6151
R18620 vdd.n2820 vdd.n2819 10.6151
R18621 vdd.n2821 vdd.n2820 10.6151
R18622 vdd.n2821 vdd.n837 10.6151
R18623 vdd.n2831 vdd.n837 10.6151
R18624 vdd.n2832 vdd.n2831 10.6151
R18625 vdd.n2833 vdd.n2832 10.6151
R18626 vdd.n2833 vdd.n826 10.6151
R18627 vdd.n2845 vdd.n826 10.6151
R18628 vdd.n2846 vdd.n2845 10.6151
R18629 vdd.n2847 vdd.n2846 10.6151
R18630 vdd.n2847 vdd.n812 10.6151
R18631 vdd.n2902 vdd.n812 10.6151
R18632 vdd.n2903 vdd.n2902 10.6151
R18633 vdd.n2904 vdd.n2903 10.6151
R18634 vdd.n2904 vdd.n779 10.6151
R18635 vdd.n2974 vdd.n779 10.6151
R18636 vdd.n2973 vdd.n2972 10.6151
R18637 vdd.n2972 vdd.n780 10.6151
R18638 vdd.n781 vdd.n780 10.6151
R18639 vdd.n2965 vdd.n781 10.6151
R18640 vdd.n2965 vdd.n2964 10.6151
R18641 vdd.n2964 vdd.n2963 10.6151
R18642 vdd.n2963 vdd.n783 10.6151
R18643 vdd.n2958 vdd.n783 10.6151
R18644 vdd.n2958 vdd.n2957 10.6151
R18645 vdd.n2957 vdd.n2956 10.6151
R18646 vdd.n2956 vdd.n786 10.6151
R18647 vdd.n2951 vdd.n786 10.6151
R18648 vdd.n2951 vdd.n2950 10.6151
R18649 vdd.n2950 vdd.n2949 10.6151
R18650 vdd.n2949 vdd.n789 10.6151
R18651 vdd.n2944 vdd.n789 10.6151
R18652 vdd.n2944 vdd.n2943 10.6151
R18653 vdd.n2943 vdd.n2941 10.6151
R18654 vdd.n2941 vdd.n792 10.6151
R18655 vdd.n2936 vdd.n792 10.6151
R18656 vdd.n2936 vdd.n2935 10.6151
R18657 vdd.n2935 vdd.n2934 10.6151
R18658 vdd.n2934 vdd.n795 10.6151
R18659 vdd.n2929 vdd.n795 10.6151
R18660 vdd.n2929 vdd.n2928 10.6151
R18661 vdd.n2928 vdd.n2927 10.6151
R18662 vdd.n2927 vdd.n798 10.6151
R18663 vdd.n2922 vdd.n798 10.6151
R18664 vdd.n2922 vdd.n2921 10.6151
R18665 vdd.n2921 vdd.n2920 10.6151
R18666 vdd.n2920 vdd.n801 10.6151
R18667 vdd.n2915 vdd.n2914 10.6151
R18668 vdd.n2914 vdd.n2913 10.6151
R18669 vdd.n2892 vdd.n2853 10.6151
R18670 vdd.n2887 vdd.n2853 10.6151
R18671 vdd.n2887 vdd.n2886 10.6151
R18672 vdd.n2886 vdd.n2885 10.6151
R18673 vdd.n2885 vdd.n2855 10.6151
R18674 vdd.n2880 vdd.n2855 10.6151
R18675 vdd.n2880 vdd.n2879 10.6151
R18676 vdd.n2879 vdd.n2878 10.6151
R18677 vdd.n2878 vdd.n2858 10.6151
R18678 vdd.n2873 vdd.n2858 10.6151
R18679 vdd.n2873 vdd.n2872 10.6151
R18680 vdd.n2872 vdd.n2871 10.6151
R18681 vdd.n2871 vdd.n2861 10.6151
R18682 vdd.n2866 vdd.n2861 10.6151
R18683 vdd.n2866 vdd.n2865 10.6151
R18684 vdd.n2865 vdd.n753 10.6151
R18685 vdd.n3009 vdd.n753 10.6151
R18686 vdd.n3009 vdd.n754 10.6151
R18687 vdd.n757 vdd.n754 10.6151
R18688 vdd.n3002 vdd.n757 10.6151
R18689 vdd.n3002 vdd.n3001 10.6151
R18690 vdd.n3001 vdd.n3000 10.6151
R18691 vdd.n3000 vdd.n759 10.6151
R18692 vdd.n2995 vdd.n759 10.6151
R18693 vdd.n2995 vdd.n2994 10.6151
R18694 vdd.n2994 vdd.n2993 10.6151
R18695 vdd.n2993 vdd.n762 10.6151
R18696 vdd.n2988 vdd.n762 10.6151
R18697 vdd.n2988 vdd.n2987 10.6151
R18698 vdd.n2987 vdd.n2986 10.6151
R18699 vdd.n2986 vdd.n765 10.6151
R18700 vdd.n2981 vdd.n2980 10.6151
R18701 vdd.n2980 vdd.n2979 10.6151
R18702 vdd.n2627 vdd.n2625 10.6151
R18703 vdd.n2628 vdd.n2627 10.6151
R18704 vdd.n2696 vdd.n2628 10.6151
R18705 vdd.n2696 vdd.n2695 10.6151
R18706 vdd.n2695 vdd.n2694 10.6151
R18707 vdd.n2694 vdd.n2692 10.6151
R18708 vdd.n2692 vdd.n2691 10.6151
R18709 vdd.n2691 vdd.n2689 10.6151
R18710 vdd.n2689 vdd.n2688 10.6151
R18711 vdd.n2688 vdd.n2686 10.6151
R18712 vdd.n2686 vdd.n2685 10.6151
R18713 vdd.n2685 vdd.n2683 10.6151
R18714 vdd.n2683 vdd.n2682 10.6151
R18715 vdd.n2682 vdd.n2680 10.6151
R18716 vdd.n2680 vdd.n2679 10.6151
R18717 vdd.n2679 vdd.n2645 10.6151
R18718 vdd.n2645 vdd.n2644 10.6151
R18719 vdd.n2644 vdd.n2642 10.6151
R18720 vdd.n2642 vdd.n2641 10.6151
R18721 vdd.n2641 vdd.n2639 10.6151
R18722 vdd.n2639 vdd.n2638 10.6151
R18723 vdd.n2638 vdd.n2636 10.6151
R18724 vdd.n2636 vdd.n2635 10.6151
R18725 vdd.n2635 vdd.n2633 10.6151
R18726 vdd.n2633 vdd.n2632 10.6151
R18727 vdd.n2632 vdd.n2630 10.6151
R18728 vdd.n2630 vdd.n2629 10.6151
R18729 vdd.n2629 vdd.n771 10.6151
R18730 vdd.n2778 vdd.n2777 10.6151
R18731 vdd.n2777 vdd.n888 10.6151
R18732 vdd.n2562 vdd.n888 10.6151
R18733 vdd.n2565 vdd.n2562 10.6151
R18734 vdd.n2566 vdd.n2565 10.6151
R18735 vdd.n2569 vdd.n2566 10.6151
R18736 vdd.n2570 vdd.n2569 10.6151
R18737 vdd.n2573 vdd.n2570 10.6151
R18738 vdd.n2574 vdd.n2573 10.6151
R18739 vdd.n2577 vdd.n2574 10.6151
R18740 vdd.n2578 vdd.n2577 10.6151
R18741 vdd.n2581 vdd.n2578 10.6151
R18742 vdd.n2582 vdd.n2581 10.6151
R18743 vdd.n2585 vdd.n2582 10.6151
R18744 vdd.n2586 vdd.n2585 10.6151
R18745 vdd.n2589 vdd.n2586 10.6151
R18746 vdd.n2590 vdd.n2589 10.6151
R18747 vdd.n2593 vdd.n2590 10.6151
R18748 vdd.n2594 vdd.n2593 10.6151
R18749 vdd.n2597 vdd.n2594 10.6151
R18750 vdd.n2598 vdd.n2597 10.6151
R18751 vdd.n2601 vdd.n2598 10.6151
R18752 vdd.n2602 vdd.n2601 10.6151
R18753 vdd.n2605 vdd.n2602 10.6151
R18754 vdd.n2606 vdd.n2605 10.6151
R18755 vdd.n2609 vdd.n2606 10.6151
R18756 vdd.n2610 vdd.n2609 10.6151
R18757 vdd.n2613 vdd.n2610 10.6151
R18758 vdd.n2614 vdd.n2613 10.6151
R18759 vdd.n2617 vdd.n2614 10.6151
R18760 vdd.n2618 vdd.n2617 10.6151
R18761 vdd.n2623 vdd.n2621 10.6151
R18762 vdd.n2624 vdd.n2623 10.6151
R18763 vdd.n2779 vdd.n878 10.6151
R18764 vdd.n2789 vdd.n878 10.6151
R18765 vdd.n2790 vdd.n2789 10.6151
R18766 vdd.n2791 vdd.n2790 10.6151
R18767 vdd.n2791 vdd.n866 10.6151
R18768 vdd.n2801 vdd.n866 10.6151
R18769 vdd.n2802 vdd.n2801 10.6151
R18770 vdd.n2803 vdd.n2802 10.6151
R18771 vdd.n2803 vdd.n855 10.6151
R18772 vdd.n2813 vdd.n855 10.6151
R18773 vdd.n2814 vdd.n2813 10.6151
R18774 vdd.n2815 vdd.n2814 10.6151
R18775 vdd.n2815 vdd.n843 10.6151
R18776 vdd.n2825 vdd.n843 10.6151
R18777 vdd.n2826 vdd.n2825 10.6151
R18778 vdd.n2827 vdd.n2826 10.6151
R18779 vdd.n2827 vdd.n832 10.6151
R18780 vdd.n2837 vdd.n832 10.6151
R18781 vdd.n2838 vdd.n2837 10.6151
R18782 vdd.n2841 vdd.n2838 10.6151
R18783 vdd.n2851 vdd.n820 10.6151
R18784 vdd.n2852 vdd.n2851 10.6151
R18785 vdd.n2898 vdd.n2852 10.6151
R18786 vdd.n2898 vdd.n2897 10.6151
R18787 vdd.n2897 vdd.n2896 10.6151
R18788 vdd.n2896 vdd.n2895 10.6151
R18789 vdd.n2895 vdd.n2893 10.6151
R18790 vdd.n2290 vdd.n1012 10.6151
R18791 vdd.n2300 vdd.n1012 10.6151
R18792 vdd.n2301 vdd.n2300 10.6151
R18793 vdd.n2302 vdd.n2301 10.6151
R18794 vdd.n2302 vdd.n999 10.6151
R18795 vdd.n2312 vdd.n999 10.6151
R18796 vdd.n2313 vdd.n2312 10.6151
R18797 vdd.n2315 vdd.n987 10.6151
R18798 vdd.n2325 vdd.n987 10.6151
R18799 vdd.n2326 vdd.n2325 10.6151
R18800 vdd.n2327 vdd.n2326 10.6151
R18801 vdd.n2327 vdd.n975 10.6151
R18802 vdd.n2337 vdd.n975 10.6151
R18803 vdd.n2338 vdd.n2337 10.6151
R18804 vdd.n2339 vdd.n2338 10.6151
R18805 vdd.n2339 vdd.n964 10.6151
R18806 vdd.n2349 vdd.n964 10.6151
R18807 vdd.n2350 vdd.n2349 10.6151
R18808 vdd.n2351 vdd.n2350 10.6151
R18809 vdd.n2351 vdd.n952 10.6151
R18810 vdd.n2361 vdd.n952 10.6151
R18811 vdd.n2362 vdd.n2361 10.6151
R18812 vdd.n2365 vdd.n2362 10.6151
R18813 vdd.n2365 vdd.n2364 10.6151
R18814 vdd.n2364 vdd.n2363 10.6151
R18815 vdd.n2363 vdd.n935 10.6151
R18816 vdd.n2447 vdd.n935 10.6151
R18817 vdd.n2446 vdd.n2445 10.6151
R18818 vdd.n2445 vdd.n2442 10.6151
R18819 vdd.n2442 vdd.n2441 10.6151
R18820 vdd.n2441 vdd.n2438 10.6151
R18821 vdd.n2438 vdd.n2437 10.6151
R18822 vdd.n2437 vdd.n2434 10.6151
R18823 vdd.n2434 vdd.n2433 10.6151
R18824 vdd.n2433 vdd.n2430 10.6151
R18825 vdd.n2430 vdd.n2429 10.6151
R18826 vdd.n2429 vdd.n2426 10.6151
R18827 vdd.n2426 vdd.n2425 10.6151
R18828 vdd.n2425 vdd.n2422 10.6151
R18829 vdd.n2422 vdd.n2421 10.6151
R18830 vdd.n2421 vdd.n2418 10.6151
R18831 vdd.n2418 vdd.n2417 10.6151
R18832 vdd.n2417 vdd.n2414 10.6151
R18833 vdd.n2414 vdd.n2413 10.6151
R18834 vdd.n2413 vdd.n2410 10.6151
R18835 vdd.n2410 vdd.n2409 10.6151
R18836 vdd.n2409 vdd.n2406 10.6151
R18837 vdd.n2406 vdd.n2405 10.6151
R18838 vdd.n2405 vdd.n2402 10.6151
R18839 vdd.n2402 vdd.n2401 10.6151
R18840 vdd.n2401 vdd.n2398 10.6151
R18841 vdd.n2398 vdd.n2397 10.6151
R18842 vdd.n2397 vdd.n2394 10.6151
R18843 vdd.n2394 vdd.n2393 10.6151
R18844 vdd.n2393 vdd.n2390 10.6151
R18845 vdd.n2390 vdd.n2389 10.6151
R18846 vdd.n2389 vdd.n2386 10.6151
R18847 vdd.n2386 vdd.n2385 10.6151
R18848 vdd.n2382 vdd.n2381 10.6151
R18849 vdd.n2381 vdd.n2379 10.6151
R18850 vdd.n2138 vdd.n2136 10.6151
R18851 vdd.n2139 vdd.n2138 10.6151
R18852 vdd.n2141 vdd.n2139 10.6151
R18853 vdd.n2142 vdd.n2141 10.6151
R18854 vdd.n2144 vdd.n2142 10.6151
R18855 vdd.n2145 vdd.n2144 10.6151
R18856 vdd.n2147 vdd.n2145 10.6151
R18857 vdd.n2148 vdd.n2147 10.6151
R18858 vdd.n2150 vdd.n2148 10.6151
R18859 vdd.n2151 vdd.n2150 10.6151
R18860 vdd.n2153 vdd.n2151 10.6151
R18861 vdd.n2154 vdd.n2153 10.6151
R18862 vdd.n2172 vdd.n2154 10.6151
R18863 vdd.n2172 vdd.n2171 10.6151
R18864 vdd.n2171 vdd.n2170 10.6151
R18865 vdd.n2170 vdd.n2168 10.6151
R18866 vdd.n2168 vdd.n2167 10.6151
R18867 vdd.n2167 vdd.n2165 10.6151
R18868 vdd.n2165 vdd.n2164 10.6151
R18869 vdd.n2164 vdd.n2162 10.6151
R18870 vdd.n2162 vdd.n2161 10.6151
R18871 vdd.n2161 vdd.n2159 10.6151
R18872 vdd.n2159 vdd.n2158 10.6151
R18873 vdd.n2158 vdd.n2156 10.6151
R18874 vdd.n2156 vdd.n2155 10.6151
R18875 vdd.n2155 vdd.n939 10.6151
R18876 vdd.n2377 vdd.n939 10.6151
R18877 vdd.n2378 vdd.n2377 10.6151
R18878 vdd.n2289 vdd.n2288 10.6151
R18879 vdd.n2288 vdd.n1024 10.6151
R18880 vdd.n2282 vdd.n1024 10.6151
R18881 vdd.n2282 vdd.n2281 10.6151
R18882 vdd.n2281 vdd.n2280 10.6151
R18883 vdd.n2280 vdd.n1026 10.6151
R18884 vdd.n2274 vdd.n1026 10.6151
R18885 vdd.n2274 vdd.n2273 10.6151
R18886 vdd.n2273 vdd.n2272 10.6151
R18887 vdd.n2272 vdd.n1028 10.6151
R18888 vdd.n2266 vdd.n1028 10.6151
R18889 vdd.n2266 vdd.n2265 10.6151
R18890 vdd.n2265 vdd.n2264 10.6151
R18891 vdd.n2264 vdd.n1030 10.6151
R18892 vdd.n2258 vdd.n1030 10.6151
R18893 vdd.n2258 vdd.n2257 10.6151
R18894 vdd.n2257 vdd.n2256 10.6151
R18895 vdd.n2256 vdd.n1034 10.6151
R18896 vdd.n2104 vdd.n1034 10.6151
R18897 vdd.n2105 vdd.n2104 10.6151
R18898 vdd.n2105 vdd.n2100 10.6151
R18899 vdd.n2111 vdd.n2100 10.6151
R18900 vdd.n2112 vdd.n2111 10.6151
R18901 vdd.n2113 vdd.n2112 10.6151
R18902 vdd.n2113 vdd.n2098 10.6151
R18903 vdd.n2119 vdd.n2098 10.6151
R18904 vdd.n2120 vdd.n2119 10.6151
R18905 vdd.n2121 vdd.n2120 10.6151
R18906 vdd.n2121 vdd.n2096 10.6151
R18907 vdd.n2127 vdd.n2096 10.6151
R18908 vdd.n2128 vdd.n2127 10.6151
R18909 vdd.n2130 vdd.n2092 10.6151
R18910 vdd.n2135 vdd.n2092 10.6151
R18911 vdd.t216 vdd.n1776 10.5435
R18912 vdd.n636 vdd.t130 10.5435
R18913 vdd.n304 vdd.n286 10.4732
R18914 vdd.n249 vdd.n231 10.4732
R18915 vdd.n206 vdd.n188 10.4732
R18916 vdd.n151 vdd.n133 10.4732
R18917 vdd.n109 vdd.n91 10.4732
R18918 vdd.n54 vdd.n36 10.4732
R18919 vdd.n1673 vdd.n1655 10.4732
R18920 vdd.n1728 vdd.n1710 10.4732
R18921 vdd.n1575 vdd.n1557 10.4732
R18922 vdd.n1630 vdd.n1612 10.4732
R18923 vdd.n1478 vdd.n1460 10.4732
R18924 vdd.n1533 vdd.n1515 10.4732
R18925 vdd.n1760 vdd.t186 10.3167
R18926 vdd.n3205 vdd.t128 10.3167
R18927 vdd.t142 vdd.n1104 10.09
R18928 vdd.n1812 vdd.t43 10.09
R18929 vdd.n3153 vdd.t28 10.09
R18930 vdd.n3286 vdd.t132 10.09
R18931 vdd.n1424 vdd.t160 9.86327
R18932 vdd.n3277 vdd.t194 9.86327
R18933 vdd.n303 vdd.n288 9.69747
R18934 vdd.n248 vdd.n233 9.69747
R18935 vdd.n205 vdd.n190 9.69747
R18936 vdd.n150 vdd.n135 9.69747
R18937 vdd.n108 vdd.n93 9.69747
R18938 vdd.n53 vdd.n38 9.69747
R18939 vdd.n1672 vdd.n1657 9.69747
R18940 vdd.n1727 vdd.n1712 9.69747
R18941 vdd.n1574 vdd.n1559 9.69747
R18942 vdd.n1629 vdd.n1614 9.69747
R18943 vdd.n1477 vdd.n1462 9.69747
R18944 vdd.n1532 vdd.n1517 9.69747
R18945 vdd.n2232 vdd.n2231 9.67831
R18946 vdd.n2943 vdd.n2942 9.67831
R18947 vdd.n3010 vdd.n3009 9.67831
R18948 vdd.n2256 vdd.n2255 9.67831
R18949 vdd.t140 vdd.n1398 9.63654
R18950 vdd.n3236 vdd.t153 9.63654
R18951 vdd.n319 vdd.n318 9.45567
R18952 vdd.n264 vdd.n263 9.45567
R18953 vdd.n221 vdd.n220 9.45567
R18954 vdd.n166 vdd.n165 9.45567
R18955 vdd.n124 vdd.n123 9.45567
R18956 vdd.n69 vdd.n68 9.45567
R18957 vdd.n1688 vdd.n1687 9.45567
R18958 vdd.n1743 vdd.n1742 9.45567
R18959 vdd.n1590 vdd.n1589 9.45567
R18960 vdd.n1645 vdd.n1644 9.45567
R18961 vdd.n1493 vdd.n1492 9.45567
R18962 vdd.n1548 vdd.n1547 9.45567
R18963 vdd.n1992 vdd.n1846 9.3005
R18964 vdd.n1991 vdd.n1990 9.3005
R18965 vdd.n1852 vdd.n1851 9.3005
R18966 vdd.n1985 vdd.n1856 9.3005
R18967 vdd.n1984 vdd.n1857 9.3005
R18968 vdd.n1983 vdd.n1858 9.3005
R18969 vdd.n1862 vdd.n1859 9.3005
R18970 vdd.n1978 vdd.n1863 9.3005
R18971 vdd.n1977 vdd.n1864 9.3005
R18972 vdd.n1976 vdd.n1865 9.3005
R18973 vdd.n1869 vdd.n1866 9.3005
R18974 vdd.n1971 vdd.n1870 9.3005
R18975 vdd.n1970 vdd.n1871 9.3005
R18976 vdd.n1969 vdd.n1872 9.3005
R18977 vdd.n1876 vdd.n1873 9.3005
R18978 vdd.n1964 vdd.n1877 9.3005
R18979 vdd.n1963 vdd.n1878 9.3005
R18980 vdd.n1962 vdd.n1879 9.3005
R18981 vdd.n1883 vdd.n1880 9.3005
R18982 vdd.n1957 vdd.n1884 9.3005
R18983 vdd.n1956 vdd.n1885 9.3005
R18984 vdd.n1955 vdd.n1954 9.3005
R18985 vdd.n1953 vdd.n1886 9.3005
R18986 vdd.n1952 vdd.n1951 9.3005
R18987 vdd.n1892 vdd.n1891 9.3005
R18988 vdd.n1946 vdd.n1896 9.3005
R18989 vdd.n1945 vdd.n1897 9.3005
R18990 vdd.n1944 vdd.n1898 9.3005
R18991 vdd.n1902 vdd.n1899 9.3005
R18992 vdd.n1939 vdd.n1903 9.3005
R18993 vdd.n1938 vdd.n1904 9.3005
R18994 vdd.n1937 vdd.n1905 9.3005
R18995 vdd.n1909 vdd.n1906 9.3005
R18996 vdd.n1932 vdd.n1910 9.3005
R18997 vdd.n1931 vdd.n1911 9.3005
R18998 vdd.n1930 vdd.n1912 9.3005
R18999 vdd.n1914 vdd.n1913 9.3005
R19000 vdd.n1925 vdd.n1035 9.3005
R19001 vdd.n1994 vdd.n1993 9.3005
R19002 vdd.n2018 vdd.n2017 9.3005
R19003 vdd.n1824 vdd.n1823 9.3005
R19004 vdd.n1829 vdd.n1827 9.3005
R19005 vdd.n2010 vdd.n1830 9.3005
R19006 vdd.n2009 vdd.n1831 9.3005
R19007 vdd.n2008 vdd.n1832 9.3005
R19008 vdd.n1836 vdd.n1833 9.3005
R19009 vdd.n2003 vdd.n1837 9.3005
R19010 vdd.n2002 vdd.n1838 9.3005
R19011 vdd.n2001 vdd.n1839 9.3005
R19012 vdd.n1843 vdd.n1840 9.3005
R19013 vdd.n1996 vdd.n1844 9.3005
R19014 vdd.n1995 vdd.n1845 9.3005
R19015 vdd.n2240 vdd.n1817 9.3005
R19016 vdd.n2242 vdd.n2241 9.3005
R19017 vdd.n1748 vdd.n1094 9.3005
R19018 vdd.n1750 vdd.n1749 9.3005
R19019 vdd.n1085 vdd.n1084 9.3005
R19020 vdd.n1763 vdd.n1762 9.3005
R19021 vdd.n1764 vdd.n1083 9.3005
R19022 vdd.n1766 vdd.n1765 9.3005
R19023 vdd.n1073 vdd.n1072 9.3005
R19024 vdd.n1780 vdd.n1779 9.3005
R19025 vdd.n1781 vdd.n1071 9.3005
R19026 vdd.n1783 vdd.n1782 9.3005
R19027 vdd.n1062 vdd.n1061 9.3005
R19028 vdd.n1797 vdd.n1796 9.3005
R19029 vdd.n1798 vdd.n1060 9.3005
R19030 vdd.n1800 vdd.n1799 9.3005
R19031 vdd.n1050 vdd.n1049 9.3005
R19032 vdd.n1815 vdd.n1814 9.3005
R19033 vdd.n1816 vdd.n1048 9.3005
R19034 vdd.n2244 vdd.n2243 9.3005
R19035 vdd.n295 vdd.n294 9.3005
R19036 vdd.n290 vdd.n289 9.3005
R19037 vdd.n301 vdd.n300 9.3005
R19038 vdd.n303 vdd.n302 9.3005
R19039 vdd.n286 vdd.n285 9.3005
R19040 vdd.n309 vdd.n308 9.3005
R19041 vdd.n311 vdd.n310 9.3005
R19042 vdd.n283 vdd.n280 9.3005
R19043 vdd.n318 vdd.n317 9.3005
R19044 vdd.n240 vdd.n239 9.3005
R19045 vdd.n235 vdd.n234 9.3005
R19046 vdd.n246 vdd.n245 9.3005
R19047 vdd.n248 vdd.n247 9.3005
R19048 vdd.n231 vdd.n230 9.3005
R19049 vdd.n254 vdd.n253 9.3005
R19050 vdd.n256 vdd.n255 9.3005
R19051 vdd.n228 vdd.n225 9.3005
R19052 vdd.n263 vdd.n262 9.3005
R19053 vdd.n197 vdd.n196 9.3005
R19054 vdd.n192 vdd.n191 9.3005
R19055 vdd.n203 vdd.n202 9.3005
R19056 vdd.n205 vdd.n204 9.3005
R19057 vdd.n188 vdd.n187 9.3005
R19058 vdd.n211 vdd.n210 9.3005
R19059 vdd.n213 vdd.n212 9.3005
R19060 vdd.n185 vdd.n182 9.3005
R19061 vdd.n220 vdd.n219 9.3005
R19062 vdd.n142 vdd.n141 9.3005
R19063 vdd.n137 vdd.n136 9.3005
R19064 vdd.n148 vdd.n147 9.3005
R19065 vdd.n150 vdd.n149 9.3005
R19066 vdd.n133 vdd.n132 9.3005
R19067 vdd.n156 vdd.n155 9.3005
R19068 vdd.n158 vdd.n157 9.3005
R19069 vdd.n130 vdd.n127 9.3005
R19070 vdd.n165 vdd.n164 9.3005
R19071 vdd.n100 vdd.n99 9.3005
R19072 vdd.n95 vdd.n94 9.3005
R19073 vdd.n106 vdd.n105 9.3005
R19074 vdd.n108 vdd.n107 9.3005
R19075 vdd.n91 vdd.n90 9.3005
R19076 vdd.n114 vdd.n113 9.3005
R19077 vdd.n116 vdd.n115 9.3005
R19078 vdd.n88 vdd.n85 9.3005
R19079 vdd.n123 vdd.n122 9.3005
R19080 vdd.n45 vdd.n44 9.3005
R19081 vdd.n40 vdd.n39 9.3005
R19082 vdd.n51 vdd.n50 9.3005
R19083 vdd.n53 vdd.n52 9.3005
R19084 vdd.n36 vdd.n35 9.3005
R19085 vdd.n59 vdd.n58 9.3005
R19086 vdd.n61 vdd.n60 9.3005
R19087 vdd.n33 vdd.n30 9.3005
R19088 vdd.n68 vdd.n67 9.3005
R19089 vdd.n3059 vdd.n3058 9.3005
R19090 vdd.n3060 vdd.n721 9.3005
R19091 vdd.n720 vdd.n718 9.3005
R19092 vdd.n3066 vdd.n717 9.3005
R19093 vdd.n3067 vdd.n716 9.3005
R19094 vdd.n3068 vdd.n715 9.3005
R19095 vdd.n714 vdd.n712 9.3005
R19096 vdd.n3074 vdd.n711 9.3005
R19097 vdd.n3075 vdd.n710 9.3005
R19098 vdd.n3076 vdd.n709 9.3005
R19099 vdd.n708 vdd.n706 9.3005
R19100 vdd.n3082 vdd.n705 9.3005
R19101 vdd.n3083 vdd.n704 9.3005
R19102 vdd.n3084 vdd.n703 9.3005
R19103 vdd.n702 vdd.n700 9.3005
R19104 vdd.n3090 vdd.n699 9.3005
R19105 vdd.n3091 vdd.n698 9.3005
R19106 vdd.n3092 vdd.n697 9.3005
R19107 vdd.n696 vdd.n694 9.3005
R19108 vdd.n3098 vdd.n693 9.3005
R19109 vdd.n3099 vdd.n692 9.3005
R19110 vdd.n3100 vdd.n691 9.3005
R19111 vdd.n690 vdd.n688 9.3005
R19112 vdd.n3106 vdd.n685 9.3005
R19113 vdd.n3107 vdd.n684 9.3005
R19114 vdd.n3108 vdd.n683 9.3005
R19115 vdd.n682 vdd.n680 9.3005
R19116 vdd.n3114 vdd.n679 9.3005
R19117 vdd.n3115 vdd.n678 9.3005
R19118 vdd.n3116 vdd.n677 9.3005
R19119 vdd.n676 vdd.n674 9.3005
R19120 vdd.n3122 vdd.n673 9.3005
R19121 vdd.n3123 vdd.n672 9.3005
R19122 vdd.n3124 vdd.n671 9.3005
R19123 vdd.n670 vdd.n668 9.3005
R19124 vdd.n3129 vdd.n667 9.3005
R19125 vdd.n3139 vdd.n661 9.3005
R19126 vdd.n3141 vdd.n3140 9.3005
R19127 vdd.n652 vdd.n651 9.3005
R19128 vdd.n3156 vdd.n3155 9.3005
R19129 vdd.n3157 vdd.n650 9.3005
R19130 vdd.n3159 vdd.n3158 9.3005
R19131 vdd.n640 vdd.n639 9.3005
R19132 vdd.n3172 vdd.n3171 9.3005
R19133 vdd.n3173 vdd.n638 9.3005
R19134 vdd.n3175 vdd.n3174 9.3005
R19135 vdd.n628 vdd.n627 9.3005
R19136 vdd.n3189 vdd.n3188 9.3005
R19137 vdd.n3190 vdd.n626 9.3005
R19138 vdd.n3192 vdd.n3191 9.3005
R19139 vdd.n617 vdd.n616 9.3005
R19140 vdd.n3208 vdd.n3207 9.3005
R19141 vdd.n3209 vdd.n615 9.3005
R19142 vdd.n3211 vdd.n3210 9.3005
R19143 vdd.n324 vdd.n322 9.3005
R19144 vdd.n3143 vdd.n3142 9.3005
R19145 vdd.n3290 vdd.n3289 9.3005
R19146 vdd.n325 vdd.n323 9.3005
R19147 vdd.n3283 vdd.n334 9.3005
R19148 vdd.n3282 vdd.n335 9.3005
R19149 vdd.n3281 vdd.n336 9.3005
R19150 vdd.n343 vdd.n337 9.3005
R19151 vdd.n3275 vdd.n344 9.3005
R19152 vdd.n3274 vdd.n345 9.3005
R19153 vdd.n3273 vdd.n346 9.3005
R19154 vdd.n354 vdd.n347 9.3005
R19155 vdd.n3267 vdd.n355 9.3005
R19156 vdd.n3266 vdd.n356 9.3005
R19157 vdd.n3265 vdd.n357 9.3005
R19158 vdd.n365 vdd.n358 9.3005
R19159 vdd.n3259 vdd.n366 9.3005
R19160 vdd.n3258 vdd.n367 9.3005
R19161 vdd.n3257 vdd.n368 9.3005
R19162 vdd.n443 vdd.n369 9.3005
R19163 vdd.n447 vdd.n442 9.3005
R19164 vdd.n451 vdd.n450 9.3005
R19165 vdd.n452 vdd.n441 9.3005
R19166 vdd.n456 vdd.n453 9.3005
R19167 vdd.n457 vdd.n440 9.3005
R19168 vdd.n461 vdd.n460 9.3005
R19169 vdd.n462 vdd.n439 9.3005
R19170 vdd.n466 vdd.n463 9.3005
R19171 vdd.n467 vdd.n438 9.3005
R19172 vdd.n471 vdd.n470 9.3005
R19173 vdd.n472 vdd.n437 9.3005
R19174 vdd.n476 vdd.n473 9.3005
R19175 vdd.n477 vdd.n436 9.3005
R19176 vdd.n481 vdd.n480 9.3005
R19177 vdd.n482 vdd.n435 9.3005
R19178 vdd.n486 vdd.n483 9.3005
R19179 vdd.n487 vdd.n434 9.3005
R19180 vdd.n491 vdd.n490 9.3005
R19181 vdd.n492 vdd.n433 9.3005
R19182 vdd.n496 vdd.n493 9.3005
R19183 vdd.n497 vdd.n430 9.3005
R19184 vdd.n501 vdd.n500 9.3005
R19185 vdd.n502 vdd.n429 9.3005
R19186 vdd.n506 vdd.n503 9.3005
R19187 vdd.n507 vdd.n428 9.3005
R19188 vdd.n511 vdd.n510 9.3005
R19189 vdd.n512 vdd.n427 9.3005
R19190 vdd.n516 vdd.n513 9.3005
R19191 vdd.n517 vdd.n426 9.3005
R19192 vdd.n521 vdd.n520 9.3005
R19193 vdd.n522 vdd.n425 9.3005
R19194 vdd.n526 vdd.n523 9.3005
R19195 vdd.n527 vdd.n424 9.3005
R19196 vdd.n531 vdd.n530 9.3005
R19197 vdd.n532 vdd.n423 9.3005
R19198 vdd.n536 vdd.n533 9.3005
R19199 vdd.n537 vdd.n422 9.3005
R19200 vdd.n541 vdd.n540 9.3005
R19201 vdd.n542 vdd.n421 9.3005
R19202 vdd.n546 vdd.n543 9.3005
R19203 vdd.n547 vdd.n418 9.3005
R19204 vdd.n551 vdd.n550 9.3005
R19205 vdd.n552 vdd.n417 9.3005
R19206 vdd.n556 vdd.n553 9.3005
R19207 vdd.n557 vdd.n416 9.3005
R19208 vdd.n561 vdd.n560 9.3005
R19209 vdd.n562 vdd.n415 9.3005
R19210 vdd.n566 vdd.n563 9.3005
R19211 vdd.n567 vdd.n414 9.3005
R19212 vdd.n571 vdd.n570 9.3005
R19213 vdd.n572 vdd.n413 9.3005
R19214 vdd.n576 vdd.n573 9.3005
R19215 vdd.n577 vdd.n412 9.3005
R19216 vdd.n581 vdd.n580 9.3005
R19217 vdd.n582 vdd.n411 9.3005
R19218 vdd.n586 vdd.n583 9.3005
R19219 vdd.n587 vdd.n410 9.3005
R19220 vdd.n591 vdd.n590 9.3005
R19221 vdd.n592 vdd.n409 9.3005
R19222 vdd.n596 vdd.n593 9.3005
R19223 vdd.n598 vdd.n408 9.3005
R19224 vdd.n600 vdd.n599 9.3005
R19225 vdd.n3250 vdd.n3249 9.3005
R19226 vdd.n446 vdd.n444 9.3005
R19227 vdd.n3149 vdd.n655 9.3005
R19228 vdd.n3151 vdd.n3150 9.3005
R19229 vdd.n646 vdd.n645 9.3005
R19230 vdd.n3164 vdd.n3163 9.3005
R19231 vdd.n3165 vdd.n644 9.3005
R19232 vdd.n3167 vdd.n3166 9.3005
R19233 vdd.n633 vdd.n632 9.3005
R19234 vdd.n3180 vdd.n3179 9.3005
R19235 vdd.n3181 vdd.n631 9.3005
R19236 vdd.n3183 vdd.n3182 9.3005
R19237 vdd.n622 vdd.n621 9.3005
R19238 vdd.n3197 vdd.n3196 9.3005
R19239 vdd.n3198 vdd.n620 9.3005
R19240 vdd.n3203 vdd.n3199 9.3005
R19241 vdd.n3202 vdd.n3201 9.3005
R19242 vdd.n3200 vdd.n610 9.3005
R19243 vdd.n3216 vdd.n611 9.3005
R19244 vdd.n3217 vdd.n609 9.3005
R19245 vdd.n3219 vdd.n3218 9.3005
R19246 vdd.n3220 vdd.n608 9.3005
R19247 vdd.n3223 vdd.n3221 9.3005
R19248 vdd.n3224 vdd.n607 9.3005
R19249 vdd.n3226 vdd.n3225 9.3005
R19250 vdd.n3227 vdd.n606 9.3005
R19251 vdd.n3230 vdd.n3228 9.3005
R19252 vdd.n3231 vdd.n605 9.3005
R19253 vdd.n3233 vdd.n3232 9.3005
R19254 vdd.n3234 vdd.n604 9.3005
R19255 vdd.n3238 vdd.n3235 9.3005
R19256 vdd.n3239 vdd.n603 9.3005
R19257 vdd.n3241 vdd.n3240 9.3005
R19258 vdd.n3242 vdd.n602 9.3005
R19259 vdd.n3245 vdd.n3243 9.3005
R19260 vdd.n3246 vdd.n601 9.3005
R19261 vdd.n3248 vdd.n3247 9.3005
R19262 vdd.n3148 vdd.n3147 9.3005
R19263 vdd.n3012 vdd.n656 9.3005
R19264 vdd.n3017 vdd.n3011 9.3005
R19265 vdd.n3027 vdd.n748 9.3005
R19266 vdd.n3028 vdd.n747 9.3005
R19267 vdd.n746 vdd.n744 9.3005
R19268 vdd.n3034 vdd.n743 9.3005
R19269 vdd.n3035 vdd.n742 9.3005
R19270 vdd.n3036 vdd.n741 9.3005
R19271 vdd.n740 vdd.n738 9.3005
R19272 vdd.n3042 vdd.n737 9.3005
R19273 vdd.n3043 vdd.n736 9.3005
R19274 vdd.n3044 vdd.n735 9.3005
R19275 vdd.n734 vdd.n732 9.3005
R19276 vdd.n3049 vdd.n731 9.3005
R19277 vdd.n3050 vdd.n730 9.3005
R19278 vdd.n726 vdd.n725 9.3005
R19279 vdd.n3056 vdd.n3055 9.3005
R19280 vdd.n3057 vdd.n722 9.3005
R19281 vdd.n2254 vdd.n2253 9.3005
R19282 vdd.n2249 vdd.n1038 9.3005
R19283 vdd.n1380 vdd.n1379 9.3005
R19284 vdd.n1136 vdd.n1135 9.3005
R19285 vdd.n1393 vdd.n1392 9.3005
R19286 vdd.n1394 vdd.n1134 9.3005
R19287 vdd.n1396 vdd.n1395 9.3005
R19288 vdd.n1124 vdd.n1123 9.3005
R19289 vdd.n1410 vdd.n1409 9.3005
R19290 vdd.n1411 vdd.n1122 9.3005
R19291 vdd.n1413 vdd.n1412 9.3005
R19292 vdd.n1114 vdd.n1113 9.3005
R19293 vdd.n1427 vdd.n1426 9.3005
R19294 vdd.n1428 vdd.n1112 9.3005
R19295 vdd.n1430 vdd.n1429 9.3005
R19296 vdd.n1101 vdd.n1100 9.3005
R19297 vdd.n1443 vdd.n1442 9.3005
R19298 vdd.n1444 vdd.n1099 9.3005
R19299 vdd.n1446 vdd.n1445 9.3005
R19300 vdd.n1090 vdd.n1089 9.3005
R19301 vdd.n1755 vdd.n1754 9.3005
R19302 vdd.n1756 vdd.n1088 9.3005
R19303 vdd.n1758 vdd.n1757 9.3005
R19304 vdd.n1079 vdd.n1078 9.3005
R19305 vdd.n1771 vdd.n1770 9.3005
R19306 vdd.n1772 vdd.n1077 9.3005
R19307 vdd.n1774 vdd.n1773 9.3005
R19308 vdd.n1067 vdd.n1066 9.3005
R19309 vdd.n1788 vdd.n1787 9.3005
R19310 vdd.n1789 vdd.n1065 9.3005
R19311 vdd.n1791 vdd.n1790 9.3005
R19312 vdd.n1057 vdd.n1056 9.3005
R19313 vdd.n1805 vdd.n1804 9.3005
R19314 vdd.n1806 vdd.n1054 9.3005
R19315 vdd.n1810 vdd.n1809 9.3005
R19316 vdd.n1808 vdd.n1055 9.3005
R19317 vdd.n1807 vdd.n1043 9.3005
R19318 vdd.n1378 vdd.n1146 9.3005
R19319 vdd.n1271 vdd.n1147 9.3005
R19320 vdd.n1273 vdd.n1272 9.3005
R19321 vdd.n1274 vdd.n1266 9.3005
R19322 vdd.n1276 vdd.n1275 9.3005
R19323 vdd.n1277 vdd.n1265 9.3005
R19324 vdd.n1279 vdd.n1278 9.3005
R19325 vdd.n1280 vdd.n1260 9.3005
R19326 vdd.n1282 vdd.n1281 9.3005
R19327 vdd.n1283 vdd.n1259 9.3005
R19328 vdd.n1285 vdd.n1284 9.3005
R19329 vdd.n1286 vdd.n1254 9.3005
R19330 vdd.n1288 vdd.n1287 9.3005
R19331 vdd.n1289 vdd.n1253 9.3005
R19332 vdd.n1291 vdd.n1290 9.3005
R19333 vdd.n1292 vdd.n1248 9.3005
R19334 vdd.n1294 vdd.n1293 9.3005
R19335 vdd.n1295 vdd.n1247 9.3005
R19336 vdd.n1297 vdd.n1296 9.3005
R19337 vdd.n1298 vdd.n1242 9.3005
R19338 vdd.n1300 vdd.n1299 9.3005
R19339 vdd.n1301 vdd.n1241 9.3005
R19340 vdd.n1306 vdd.n1302 9.3005
R19341 vdd.n1307 vdd.n1237 9.3005
R19342 vdd.n1309 vdd.n1308 9.3005
R19343 vdd.n1310 vdd.n1236 9.3005
R19344 vdd.n1312 vdd.n1311 9.3005
R19345 vdd.n1313 vdd.n1231 9.3005
R19346 vdd.n1315 vdd.n1314 9.3005
R19347 vdd.n1316 vdd.n1230 9.3005
R19348 vdd.n1318 vdd.n1317 9.3005
R19349 vdd.n1319 vdd.n1225 9.3005
R19350 vdd.n1321 vdd.n1320 9.3005
R19351 vdd.n1322 vdd.n1224 9.3005
R19352 vdd.n1324 vdd.n1323 9.3005
R19353 vdd.n1325 vdd.n1219 9.3005
R19354 vdd.n1327 vdd.n1326 9.3005
R19355 vdd.n1328 vdd.n1218 9.3005
R19356 vdd.n1330 vdd.n1329 9.3005
R19357 vdd.n1331 vdd.n1213 9.3005
R19358 vdd.n1333 vdd.n1332 9.3005
R19359 vdd.n1334 vdd.n1212 9.3005
R19360 vdd.n1336 vdd.n1335 9.3005
R19361 vdd.n1337 vdd.n1209 9.3005
R19362 vdd.n1343 vdd.n1342 9.3005
R19363 vdd.n1344 vdd.n1208 9.3005
R19364 vdd.n1346 vdd.n1345 9.3005
R19365 vdd.n1347 vdd.n1203 9.3005
R19366 vdd.n1349 vdd.n1348 9.3005
R19367 vdd.n1350 vdd.n1202 9.3005
R19368 vdd.n1352 vdd.n1351 9.3005
R19369 vdd.n1353 vdd.n1197 9.3005
R19370 vdd.n1355 vdd.n1354 9.3005
R19371 vdd.n1356 vdd.n1196 9.3005
R19372 vdd.n1358 vdd.n1357 9.3005
R19373 vdd.n1359 vdd.n1191 9.3005
R19374 vdd.n1361 vdd.n1360 9.3005
R19375 vdd.n1362 vdd.n1190 9.3005
R19376 vdd.n1364 vdd.n1363 9.3005
R19377 vdd.n1365 vdd.n1186 9.3005
R19378 vdd.n1367 vdd.n1366 9.3005
R19379 vdd.n1368 vdd.n1185 9.3005
R19380 vdd.n1370 vdd.n1369 9.3005
R19381 vdd.n1371 vdd.n1184 9.3005
R19382 vdd.n1377 vdd.n1376 9.3005
R19383 vdd.n1385 vdd.n1384 9.3005
R19384 vdd.n1386 vdd.n1140 9.3005
R19385 vdd.n1388 vdd.n1387 9.3005
R19386 vdd.n1130 vdd.n1129 9.3005
R19387 vdd.n1402 vdd.n1401 9.3005
R19388 vdd.n1403 vdd.n1128 9.3005
R19389 vdd.n1405 vdd.n1404 9.3005
R19390 vdd.n1119 vdd.n1118 9.3005
R19391 vdd.n1419 vdd.n1418 9.3005
R19392 vdd.n1420 vdd.n1117 9.3005
R19393 vdd.n1422 vdd.n1421 9.3005
R19394 vdd.n1108 vdd.n1107 9.3005
R19395 vdd.n1435 vdd.n1434 9.3005
R19396 vdd.n1436 vdd.n1106 9.3005
R19397 vdd.n1438 vdd.n1437 9.3005
R19398 vdd.n1096 vdd.n1095 9.3005
R19399 vdd.n1452 vdd.n1451 9.3005
R19400 vdd.n1142 vdd.n1141 9.3005
R19401 vdd.n1664 vdd.n1663 9.3005
R19402 vdd.n1659 vdd.n1658 9.3005
R19403 vdd.n1670 vdd.n1669 9.3005
R19404 vdd.n1672 vdd.n1671 9.3005
R19405 vdd.n1655 vdd.n1654 9.3005
R19406 vdd.n1678 vdd.n1677 9.3005
R19407 vdd.n1680 vdd.n1679 9.3005
R19408 vdd.n1652 vdd.n1649 9.3005
R19409 vdd.n1687 vdd.n1686 9.3005
R19410 vdd.n1719 vdd.n1718 9.3005
R19411 vdd.n1714 vdd.n1713 9.3005
R19412 vdd.n1725 vdd.n1724 9.3005
R19413 vdd.n1727 vdd.n1726 9.3005
R19414 vdd.n1710 vdd.n1709 9.3005
R19415 vdd.n1733 vdd.n1732 9.3005
R19416 vdd.n1735 vdd.n1734 9.3005
R19417 vdd.n1707 vdd.n1704 9.3005
R19418 vdd.n1742 vdd.n1741 9.3005
R19419 vdd.n1566 vdd.n1565 9.3005
R19420 vdd.n1561 vdd.n1560 9.3005
R19421 vdd.n1572 vdd.n1571 9.3005
R19422 vdd.n1574 vdd.n1573 9.3005
R19423 vdd.n1557 vdd.n1556 9.3005
R19424 vdd.n1580 vdd.n1579 9.3005
R19425 vdd.n1582 vdd.n1581 9.3005
R19426 vdd.n1554 vdd.n1551 9.3005
R19427 vdd.n1589 vdd.n1588 9.3005
R19428 vdd.n1621 vdd.n1620 9.3005
R19429 vdd.n1616 vdd.n1615 9.3005
R19430 vdd.n1627 vdd.n1626 9.3005
R19431 vdd.n1629 vdd.n1628 9.3005
R19432 vdd.n1612 vdd.n1611 9.3005
R19433 vdd.n1635 vdd.n1634 9.3005
R19434 vdd.n1637 vdd.n1636 9.3005
R19435 vdd.n1609 vdd.n1606 9.3005
R19436 vdd.n1644 vdd.n1643 9.3005
R19437 vdd.n1469 vdd.n1468 9.3005
R19438 vdd.n1464 vdd.n1463 9.3005
R19439 vdd.n1475 vdd.n1474 9.3005
R19440 vdd.n1477 vdd.n1476 9.3005
R19441 vdd.n1460 vdd.n1459 9.3005
R19442 vdd.n1483 vdd.n1482 9.3005
R19443 vdd.n1485 vdd.n1484 9.3005
R19444 vdd.n1457 vdd.n1454 9.3005
R19445 vdd.n1492 vdd.n1491 9.3005
R19446 vdd.n1524 vdd.n1523 9.3005
R19447 vdd.n1519 vdd.n1518 9.3005
R19448 vdd.n1530 vdd.n1529 9.3005
R19449 vdd.n1532 vdd.n1531 9.3005
R19450 vdd.n1515 vdd.n1514 9.3005
R19451 vdd.n1538 vdd.n1537 9.3005
R19452 vdd.n1540 vdd.n1539 9.3005
R19453 vdd.n1512 vdd.n1509 9.3005
R19454 vdd.n1547 vdd.n1546 9.3005
R19455 vdd.n1398 vdd.t202 9.18308
R19456 vdd.n3236 vdd.t146 9.18308
R19457 vdd.n1424 vdd.t150 8.95635
R19458 vdd.t148 vdd.n3277 8.95635
R19459 vdd.n300 vdd.n299 8.92171
R19460 vdd.n245 vdd.n244 8.92171
R19461 vdd.n202 vdd.n201 8.92171
R19462 vdd.n147 vdd.n146 8.92171
R19463 vdd.n105 vdd.n104 8.92171
R19464 vdd.n50 vdd.n49 8.92171
R19465 vdd.n1669 vdd.n1668 8.92171
R19466 vdd.n1724 vdd.n1723 8.92171
R19467 vdd.n1571 vdd.n1570 8.92171
R19468 vdd.n1626 vdd.n1625 8.92171
R19469 vdd.n1474 vdd.n1473 8.92171
R19470 vdd.n1529 vdd.n1528 8.92171
R19471 vdd.n223 vdd.n125 8.81535
R19472 vdd.n1647 vdd.n1549 8.81535
R19473 vdd.n1104 vdd.t206 8.72962
R19474 vdd.t175 vdd.n3286 8.72962
R19475 vdd.n1760 vdd.t138 8.50289
R19476 vdd.n3205 vdd.t218 8.50289
R19477 vdd.n28 vdd.n14 8.42249
R19478 vdd.n1776 vdd.t144 8.27616
R19479 vdd.t191 vdd.n636 8.27616
R19480 vdd.n3292 vdd.n3291 8.16225
R19481 vdd.n1747 vdd.n1746 8.16225
R19482 vdd.n296 vdd.n290 8.14595
R19483 vdd.n241 vdd.n235 8.14595
R19484 vdd.n198 vdd.n192 8.14595
R19485 vdd.n143 vdd.n137 8.14595
R19486 vdd.n101 vdd.n95 8.14595
R19487 vdd.n46 vdd.n40 8.14595
R19488 vdd.n1665 vdd.n1659 8.14595
R19489 vdd.n1720 vdd.n1714 8.14595
R19490 vdd.n1567 vdd.n1561 8.14595
R19491 vdd.n1622 vdd.n1616 8.14595
R19492 vdd.n1470 vdd.n1464 8.14595
R19493 vdd.n1525 vdd.n1519 8.14595
R19494 vdd.n2840 vdd.n820 8.11757
R19495 vdd.n2314 vdd.n2313 8.11757
R19496 vdd.t36 vdd.n1138 7.8227
R19497 vdd.t32 vdd.n363 7.8227
R19498 vdd.n2292 vdd.n1014 7.70933
R19499 vdd.n2298 vdd.n1014 7.70933
R19500 vdd.n2304 vdd.n1008 7.70933
R19501 vdd.n2304 vdd.n1001 7.70933
R19502 vdd.n2310 vdd.n1001 7.70933
R19503 vdd.n2310 vdd.n1004 7.70933
R19504 vdd.n2317 vdd.n989 7.70933
R19505 vdd.n2323 vdd.n989 7.70933
R19506 vdd.n2329 vdd.n983 7.70933
R19507 vdd.n2335 vdd.n979 7.70933
R19508 vdd.n2341 vdd.n973 7.70933
R19509 vdd.n2353 vdd.n960 7.70933
R19510 vdd.n2359 vdd.n954 7.70933
R19511 vdd.n2359 vdd.n947 7.70933
R19512 vdd.n2367 vdd.n947 7.70933
R19513 vdd.n2374 vdd.t256 7.70933
R19514 vdd.n2449 vdd.t256 7.70933
R19515 vdd.n2781 vdd.t260 7.70933
R19516 vdd.n2787 vdd.t260 7.70933
R19517 vdd.n2793 vdd.n868 7.70933
R19518 vdd.n2799 vdd.n868 7.70933
R19519 vdd.n2799 vdd.n871 7.70933
R19520 vdd.n2805 vdd.n864 7.70933
R19521 vdd.n2817 vdd.n851 7.70933
R19522 vdd.n2823 vdd.n845 7.70933
R19523 vdd.n2829 vdd.n841 7.70933
R19524 vdd.n2835 vdd.n828 7.70933
R19525 vdd.n2843 vdd.n828 7.70933
R19526 vdd.n2849 vdd.n822 7.70933
R19527 vdd.n2849 vdd.n814 7.70933
R19528 vdd.n2900 vdd.n814 7.70933
R19529 vdd.n2900 vdd.n817 7.70933
R19530 vdd.n2906 vdd.n774 7.70933
R19531 vdd.n2976 vdd.n774 7.70933
R19532 vdd.n295 vdd.n292 7.3702
R19533 vdd.n240 vdd.n237 7.3702
R19534 vdd.n197 vdd.n194 7.3702
R19535 vdd.n142 vdd.n139 7.3702
R19536 vdd.n100 vdd.n97 7.3702
R19537 vdd.n45 vdd.n42 7.3702
R19538 vdd.n1664 vdd.n1661 7.3702
R19539 vdd.n1719 vdd.n1716 7.3702
R19540 vdd.n1566 vdd.n1563 7.3702
R19541 vdd.n1621 vdd.n1618 7.3702
R19542 vdd.n1469 vdd.n1466 7.3702
R19543 vdd.n1524 vdd.n1521 7.3702
R19544 vdd.n1307 vdd.n1306 6.98232
R19545 vdd.n1956 vdd.n1955 6.98232
R19546 vdd.n547 vdd.n546 6.98232
R19547 vdd.n3060 vdd.n3059 6.98232
R19548 vdd.n1794 vdd.t236 6.91577
R19549 vdd.n3169 vdd.t198 6.91577
R19550 vdd.t165 vdd.n1075 6.68904
R19551 vdd.n3185 vdd.t163 6.68904
R19552 vdd.n1752 vdd.t214 6.46231
R19553 vdd.n3213 vdd.t173 6.46231
R19554 vdd.n3292 vdd.n321 6.32949
R19555 vdd.n1746 vdd.n1745 6.32949
R19556 vdd.t178 vdd.n1103 6.23558
R19557 vdd.t168 vdd.n332 6.23558
R19558 vdd.n1416 vdd.t200 6.00885
R19559 vdd.n2329 vdd.t12 6.00885
R19560 vdd.n2829 vdd.t22 6.00885
R19561 vdd.n3271 vdd.t171 6.00885
R19562 vdd.n1004 vdd.t81 5.89549
R19563 vdd.t50 vdd.n822 5.89549
R19564 vdd.n296 vdd.n295 5.81868
R19565 vdd.n241 vdd.n240 5.81868
R19566 vdd.n198 vdd.n197 5.81868
R19567 vdd.n143 vdd.n142 5.81868
R19568 vdd.n101 vdd.n100 5.81868
R19569 vdd.n46 vdd.n45 5.81868
R19570 vdd.n1665 vdd.n1664 5.81868
R19571 vdd.n1720 vdd.n1719 5.81868
R19572 vdd.n1567 vdd.n1566 5.81868
R19573 vdd.n1622 vdd.n1621 5.81868
R19574 vdd.n1470 vdd.n1469 5.81868
R19575 vdd.n1525 vdd.n1524 5.81868
R19576 vdd.t24 vdd.n1008 5.78212
R19577 vdd.n2073 vdd.t63 5.78212
R19578 vdd.n2698 vdd.t71 5.78212
R19579 vdd.n817 vdd.t67 5.78212
R19580 vdd.n2457 vdd.n2456 5.77611
R19581 vdd.n2200 vdd.n2070 5.77611
R19582 vdd.n2711 vdd.n2710 5.77611
R19583 vdd.n2915 vdd.n806 5.77611
R19584 vdd.n2981 vdd.n770 5.77611
R19585 vdd.n2621 vdd.n2561 5.77611
R19586 vdd.n2382 vdd.n938 5.77611
R19587 vdd.n2130 vdd.n2129 5.77611
R19588 vdd.n1376 vdd.n1150 5.62474
R19589 vdd.n2252 vdd.n2249 5.62474
R19590 vdd.n3250 vdd.n407 5.62474
R19591 vdd.n3015 vdd.n3012 5.62474
R19592 vdd.t2 vdd.n960 5.44203
R19593 vdd.n864 vdd.t103 5.44203
R19594 vdd.n1126 vdd.t200 5.32866
R19595 vdd.t171 vdd.n3270 5.32866
R19596 vdd.n1432 vdd.t178 5.10193
R19597 vdd.t100 vdd.n983 5.10193
R19598 vdd.n973 vdd.t7 5.10193
R19599 vdd.t8 vdd.n851 5.10193
R19600 vdd.n841 vdd.t99 5.10193
R19601 vdd.n3279 vdd.t168 5.10193
R19602 vdd.n299 vdd.n290 5.04292
R19603 vdd.n244 vdd.n235 5.04292
R19604 vdd.n201 vdd.n192 5.04292
R19605 vdd.n146 vdd.n137 5.04292
R19606 vdd.n104 vdd.n95 5.04292
R19607 vdd.n49 vdd.n40 5.04292
R19608 vdd.n1668 vdd.n1659 5.04292
R19609 vdd.n1723 vdd.n1714 5.04292
R19610 vdd.n1570 vdd.n1561 5.04292
R19611 vdd.n1625 vdd.n1616 5.04292
R19612 vdd.n1473 vdd.n1464 5.04292
R19613 vdd.n1528 vdd.n1519 5.04292
R19614 vdd.n1448 vdd.t214 4.8752
R19615 vdd.t6 vdd.t101 4.8752
R19616 vdd.t0 vdd.t4 4.8752
R19617 vdd.t10 vdd.t105 4.8752
R19618 vdd.t117 vdd.t108 4.8752
R19619 vdd.t173 vdd.n328 4.8752
R19620 vdd.n2458 vdd.n2457 4.83952
R19621 vdd.n2070 vdd.n2066 4.83952
R19622 vdd.n2712 vdd.n2711 4.83952
R19623 vdd.n806 vdd.n801 4.83952
R19624 vdd.n770 vdd.n765 4.83952
R19625 vdd.n2618 vdd.n2561 4.83952
R19626 vdd.n2385 vdd.n938 4.83952
R19627 vdd.n2129 vdd.n2128 4.83952
R19628 vdd.n1924 vdd.n1036 4.74817
R19629 vdd.n1919 vdd.n1037 4.74817
R19630 vdd.n1821 vdd.n1818 4.74817
R19631 vdd.n2233 vdd.n1822 4.74817
R19632 vdd.n2235 vdd.n1821 4.74817
R19633 vdd.n2234 vdd.n2233 4.74817
R19634 vdd.n664 vdd.n662 4.74817
R19635 vdd.n3130 vdd.n665 4.74817
R19636 vdd.n3133 vdd.n665 4.74817
R19637 vdd.n3134 vdd.n664 4.74817
R19638 vdd.n3022 vdd.n749 4.74817
R19639 vdd.n3018 vdd.n751 4.74817
R19640 vdd.n3021 vdd.n751 4.74817
R19641 vdd.n3026 vdd.n749 4.74817
R19642 vdd.n1920 vdd.n1036 4.74817
R19643 vdd.n1039 vdd.n1037 4.74817
R19644 vdd.n321 vdd.n320 4.7074
R19645 vdd.n223 vdd.n222 4.7074
R19646 vdd.n1745 vdd.n1744 4.7074
R19647 vdd.n1647 vdd.n1646 4.7074
R19648 vdd.n1768 vdd.t165 4.64847
R19649 vdd.n3194 vdd.t163 4.64847
R19650 vdd.n2335 vdd.t258 4.53511
R19651 vdd.n2823 vdd.t121 4.53511
R19652 vdd.n1069 vdd.t236 4.42174
R19653 vdd.t198 vdd.n635 4.42174
R19654 vdd.n2367 vdd.t115 4.30838
R19655 vdd.n2793 vdd.t119 4.30838
R19656 vdd.n300 vdd.n288 4.26717
R19657 vdd.n245 vdd.n233 4.26717
R19658 vdd.n202 vdd.n190 4.26717
R19659 vdd.n147 vdd.n135 4.26717
R19660 vdd.n105 vdd.n93 4.26717
R19661 vdd.n50 vdd.n38 4.26717
R19662 vdd.n1669 vdd.n1657 4.26717
R19663 vdd.n1724 vdd.n1712 4.26717
R19664 vdd.n1571 vdd.n1559 4.26717
R19665 vdd.n1626 vdd.n1614 4.26717
R19666 vdd.n1474 vdd.n1462 4.26717
R19667 vdd.n1529 vdd.n1517 4.26717
R19668 vdd.n321 vdd.n223 4.10845
R19669 vdd.n1745 vdd.n1647 4.10845
R19670 vdd.n277 vdd.t251 4.06363
R19671 vdd.n277 vdd.t162 4.06363
R19672 vdd.n275 vdd.t183 4.06363
R19673 vdd.n275 vdd.t250 4.06363
R19674 vdd.n273 vdd.t252 4.06363
R19675 vdd.n273 vdd.t182 4.06363
R19676 vdd.n271 vdd.t188 4.06363
R19677 vdd.n271 vdd.t190 4.06363
R19678 vdd.n269 vdd.t230 4.06363
R19679 vdd.n269 vdd.t152 4.06363
R19680 vdd.n267 vdd.t157 4.06363
R19681 vdd.n267 vdd.t208 4.06363
R19682 vdd.n265 vdd.t209 4.06363
R19683 vdd.n265 vdd.t235 4.06363
R19684 vdd.n179 vdd.t241 4.06363
R19685 vdd.n179 vdd.t147 4.06363
R19686 vdd.n177 vdd.t170 4.06363
R19687 vdd.n177 vdd.t240 4.06363
R19688 vdd.n175 vdd.t227 4.06363
R19689 vdd.n175 vdd.t169 4.06363
R19690 vdd.n173 vdd.t174 4.06363
R19691 vdd.n173 vdd.t176 4.06363
R19692 vdd.n171 vdd.t219 4.06363
R19693 vdd.n171 vdd.t129 4.06363
R19694 vdd.n169 vdd.t131 4.06363
R19695 vdd.n169 vdd.t185 4.06363
R19696 vdd.n167 vdd.t199 4.06363
R19697 vdd.n167 vdd.t221 4.06363
R19698 vdd.n82 vdd.t172 4.06363
R19699 vdd.n82 vdd.t238 4.06363
R19700 vdd.n80 vdd.t149 4.06363
R19701 vdd.n80 vdd.t195 4.06363
R19702 vdd.n78 vdd.t133 4.06363
R19703 vdd.n78 vdd.t177 4.06363
R19704 vdd.n76 vdd.t248 4.06363
R19705 vdd.n76 vdd.t226 4.06363
R19706 vdd.n74 vdd.t231 4.06363
R19707 vdd.n74 vdd.t184 4.06363
R19708 vdd.n72 vdd.t253 4.06363
R19709 vdd.n72 vdd.t164 4.06363
R19710 vdd.n70 vdd.t242 4.06363
R19711 vdd.n70 vdd.t192 4.06363
R19712 vdd.n1689 vdd.t159 4.06363
R19713 vdd.n1689 vdd.t247 4.06363
R19714 vdd.n1691 vdd.t244 4.06363
R19715 vdd.n1691 vdd.t229 4.06363
R19716 vdd.n1693 vdd.t204 4.06363
R19717 vdd.n1693 vdd.t156 4.06363
R19718 vdd.n1695 vdd.t255 4.06363
R19719 vdd.n1695 vdd.t225 4.06363
R19720 vdd.n1697 vdd.t222 4.06363
R19721 vdd.n1697 vdd.t181 4.06363
R19722 vdd.n1699 vdd.t180 4.06363
R19723 vdd.n1699 vdd.t223 4.06363
R19724 vdd.n1701 vdd.t211 4.06363
R19725 vdd.n1701 vdd.t210 4.06363
R19726 vdd.n1591 vdd.t145 4.06363
R19727 vdd.n1591 vdd.t237 4.06363
R19728 vdd.n1593 vdd.t228 4.06363
R19729 vdd.n1593 vdd.t217 4.06363
R19730 vdd.n1595 vdd.t189 4.06363
R19731 vdd.n1595 vdd.t139 4.06363
R19732 vdd.n1597 vdd.t245 4.06363
R19733 vdd.n1597 vdd.t215 4.06363
R19734 vdd.n1599 vdd.t212 4.06363
R19735 vdd.n1599 vdd.t167 4.06363
R19736 vdd.n1601 vdd.t161 4.06363
R19737 vdd.n1601 vdd.t213 4.06363
R19738 vdd.n1603 vdd.t203 4.06363
R19739 vdd.n1603 vdd.t201 4.06363
R19740 vdd.n1494 vdd.t193 4.06363
R19741 vdd.n1494 vdd.t243 4.06363
R19742 vdd.n1496 vdd.t166 4.06363
R19743 vdd.n1496 vdd.t224 4.06363
R19744 vdd.n1498 vdd.t187 4.06363
R19745 vdd.n1498 vdd.t232 4.06363
R19746 vdd.n1500 vdd.t207 4.06363
R19747 vdd.n1500 vdd.t249 4.06363
R19748 vdd.n1502 vdd.t179 4.06363
R19749 vdd.n1502 vdd.t143 4.06363
R19750 vdd.n1504 vdd.t196 4.06363
R19751 vdd.n1504 vdd.t151 4.06363
R19752 vdd.n1506 vdd.t239 4.06363
R19753 vdd.n1506 vdd.t254 4.06363
R19754 vdd.n26 vdd.t125 3.9605
R19755 vdd.n26 vdd.t16 3.9605
R19756 vdd.n23 vdd.t19 3.9605
R19757 vdd.n23 vdd.t20 3.9605
R19758 vdd.n21 vdd.t15 3.9605
R19759 vdd.n21 vdd.t112 3.9605
R19760 vdd.n20 vdd.t21 3.9605
R19761 vdd.n20 vdd.t124 3.9605
R19762 vdd.n15 vdd.t114 3.9605
R19763 vdd.n15 vdd.t126 3.9605
R19764 vdd.n16 vdd.t18 3.9605
R19765 vdd.n16 vdd.t123 3.9605
R19766 vdd.n18 vdd.t17 3.9605
R19767 vdd.n18 vdd.t127 3.9605
R19768 vdd.n25 vdd.t113 3.9605
R19769 vdd.n25 vdd.t111 3.9605
R19770 vdd.n7 vdd.t118 3.61217
R19771 vdd.n7 vdd.t122 3.61217
R19772 vdd.n8 vdd.t11 3.61217
R19773 vdd.n8 vdd.t104 3.61217
R19774 vdd.n10 vdd.t261 3.61217
R19775 vdd.n10 vdd.t120 3.61217
R19776 vdd.n12 vdd.t263 3.61217
R19777 vdd.n12 vdd.t107 3.61217
R19778 vdd.n5 vdd.t110 3.61217
R19779 vdd.n5 vdd.t14 3.61217
R19780 vdd.n3 vdd.t116 3.61217
R19781 vdd.n3 vdd.t257 3.61217
R19782 vdd.n1 vdd.t3 3.61217
R19783 vdd.n1 vdd.t5 3.61217
R19784 vdd.n0 vdd.t259 3.61217
R19785 vdd.n0 vdd.t102 3.61217
R19786 vdd.n1382 vdd.t36 3.51482
R19787 vdd.n3255 vdd.t32 3.51482
R19788 vdd.n304 vdd.n303 3.49141
R19789 vdd.n249 vdd.n248 3.49141
R19790 vdd.n206 vdd.n205 3.49141
R19791 vdd.n151 vdd.n150 3.49141
R19792 vdd.n109 vdd.n108 3.49141
R19793 vdd.n54 vdd.n53 3.49141
R19794 vdd.n1673 vdd.n1672 3.49141
R19795 vdd.n1728 vdd.n1727 3.49141
R19796 vdd.n1575 vdd.n1574 3.49141
R19797 vdd.n1630 vdd.n1629 3.49141
R19798 vdd.n1478 vdd.n1477 3.49141
R19799 vdd.n1533 vdd.n1532 3.49141
R19800 vdd.n2073 vdd.t115 3.40145
R19801 vdd.n2521 vdd.t109 3.40145
R19802 vdd.n2774 vdd.t106 3.40145
R19803 vdd.n2698 vdd.t119 3.40145
R19804 vdd.n2174 vdd.t258 3.17472
R19805 vdd.n2677 vdd.t121 3.17472
R19806 vdd.n1785 vdd.t144 3.06136
R19807 vdd.n3177 vdd.t191 3.06136
R19808 vdd.t138 vdd.n1081 2.83463
R19809 vdd.n624 vdd.t218 2.83463
R19810 vdd.n307 vdd.n286 2.71565
R19811 vdd.n252 vdd.n231 2.71565
R19812 vdd.n209 vdd.n188 2.71565
R19813 vdd.n154 vdd.n133 2.71565
R19814 vdd.n112 vdd.n91 2.71565
R19815 vdd.n57 vdd.n36 2.71565
R19816 vdd.n1676 vdd.n1655 2.71565
R19817 vdd.n1731 vdd.n1710 2.71565
R19818 vdd.n1578 vdd.n1557 2.71565
R19819 vdd.n1633 vdd.n1612 2.71565
R19820 vdd.n1481 vdd.n1460 2.71565
R19821 vdd.n1536 vdd.n1515 2.71565
R19822 vdd.n1449 vdd.t206 2.6079
R19823 vdd.n2323 vdd.t100 2.6079
R19824 vdd.n2347 vdd.t7 2.6079
R19825 vdd.n2811 vdd.t8 2.6079
R19826 vdd.n2835 vdd.t99 2.6079
R19827 vdd.n3287 vdd.t175 2.6079
R19828 vdd.n2841 vdd.n2840 2.49806
R19829 vdd.n2315 vdd.n2314 2.49806
R19830 vdd.n294 vdd.n293 2.4129
R19831 vdd.n239 vdd.n238 2.4129
R19832 vdd.n196 vdd.n195 2.4129
R19833 vdd.n141 vdd.n140 2.4129
R19834 vdd.n99 vdd.n98 2.4129
R19835 vdd.n44 vdd.n43 2.4129
R19836 vdd.n1663 vdd.n1662 2.4129
R19837 vdd.n1718 vdd.n1717 2.4129
R19838 vdd.n1565 vdd.n1564 2.4129
R19839 vdd.n1620 vdd.n1619 2.4129
R19840 vdd.n1468 vdd.n1467 2.4129
R19841 vdd.n1523 vdd.n1522 2.4129
R19842 vdd.t150 vdd.n1110 2.38117
R19843 vdd.n3278 vdd.t148 2.38117
R19844 vdd.n2232 vdd.n1821 2.27742
R19845 vdd.n2233 vdd.n2232 2.27742
R19846 vdd.n2942 vdd.n665 2.27742
R19847 vdd.n2942 vdd.n664 2.27742
R19848 vdd.n3010 vdd.n751 2.27742
R19849 vdd.n3010 vdd.n749 2.27742
R19850 vdd.n2255 vdd.n1036 2.27742
R19851 vdd.n2255 vdd.n1037 2.27742
R19852 vdd.n2347 vdd.t2 2.2678
R19853 vdd.n2811 vdd.t103 2.2678
R19854 vdd.n1407 vdd.t202 2.15444
R19855 vdd.n3269 vdd.t146 2.15444
R19856 vdd.t4 vdd.n954 2.04107
R19857 vdd.n871 vdd.t10 2.04107
R19858 vdd.n308 vdd.n284 1.93989
R19859 vdd.n253 vdd.n229 1.93989
R19860 vdd.n210 vdd.n186 1.93989
R19861 vdd.n155 vdd.n131 1.93989
R19862 vdd.n113 vdd.n89 1.93989
R19863 vdd.n58 vdd.n34 1.93989
R19864 vdd.n1677 vdd.n1653 1.93989
R19865 vdd.n1732 vdd.n1708 1.93989
R19866 vdd.n1579 vdd.n1555 1.93989
R19867 vdd.n1634 vdd.n1610 1.93989
R19868 vdd.n1482 vdd.n1458 1.93989
R19869 vdd.n1537 vdd.n1513 1.93989
R19870 vdd.n2298 vdd.t24 1.92771
R19871 vdd.n2374 vdd.t63 1.92771
R19872 vdd.n2787 vdd.t71 1.92771
R19873 vdd.n2906 vdd.t67 1.92771
R19874 vdd.n1399 vdd.t140 1.70098
R19875 vdd.n2174 vdd.t12 1.70098
R19876 vdd.n979 vdd.t6 1.70098
R19877 vdd.t108 vdd.n845 1.70098
R19878 vdd.n2677 vdd.t22 1.70098
R19879 vdd.n3263 vdd.t153 1.70098
R19880 vdd.n1415 vdd.t160 1.47425
R19881 vdd.n349 vdd.t194 1.47425
R19882 vdd.n1440 vdd.t142 1.24752
R19883 vdd.t43 vdd.n1044 1.24752
R19884 vdd.n659 vdd.t28 1.24752
R19885 vdd.t132 vdd.n3285 1.24752
R19886 vdd.n319 vdd.n279 1.16414
R19887 vdd.n312 vdd.n311 1.16414
R19888 vdd.n264 vdd.n224 1.16414
R19889 vdd.n257 vdd.n256 1.16414
R19890 vdd.n221 vdd.n181 1.16414
R19891 vdd.n214 vdd.n213 1.16414
R19892 vdd.n166 vdd.n126 1.16414
R19893 vdd.n159 vdd.n158 1.16414
R19894 vdd.n124 vdd.n84 1.16414
R19895 vdd.n117 vdd.n116 1.16414
R19896 vdd.n69 vdd.n29 1.16414
R19897 vdd.n62 vdd.n61 1.16414
R19898 vdd.n1688 vdd.n1648 1.16414
R19899 vdd.n1681 vdd.n1680 1.16414
R19900 vdd.n1743 vdd.n1703 1.16414
R19901 vdd.n1736 vdd.n1735 1.16414
R19902 vdd.n1590 vdd.n1550 1.16414
R19903 vdd.n1583 vdd.n1582 1.16414
R19904 vdd.n1645 vdd.n1605 1.16414
R19905 vdd.n1638 vdd.n1637 1.16414
R19906 vdd.n1493 vdd.n1453 1.16414
R19907 vdd.n1486 vdd.n1485 1.16414
R19908 vdd.n1548 vdd.n1508 1.16414
R19909 vdd.n1541 vdd.n1540 1.16414
R19910 vdd.n2341 vdd.t101 1.13415
R19911 vdd.n2817 vdd.t117 1.13415
R19912 vdd.n1092 vdd.t186 1.02079
R19913 vdd.t81 vdd.t1 1.02079
R19914 vdd.t9 vdd.t50 1.02079
R19915 vdd.t128 vdd.n613 1.02079
R19916 vdd.n1271 vdd.n1150 0.970197
R19917 vdd.n2253 vdd.n2252 0.970197
R19918 vdd.n599 vdd.n407 0.970197
R19919 vdd.n3017 vdd.n3015 0.970197
R19920 vdd.n1746 vdd.n28 0.852297
R19921 vdd vdd.n3292 0.844463
R19922 vdd.n1777 vdd.t216 0.794056
R19923 vdd.n2317 vdd.t1 0.794056
R19924 vdd.n2353 vdd.t0 0.794056
R19925 vdd.n2805 vdd.t105 0.794056
R19926 vdd.n2843 vdd.t9 0.794056
R19927 vdd.n3186 vdd.t130 0.794056
R19928 vdd.n1793 vdd.t136 0.567326
R19929 vdd.t134 vdd.n642 0.567326
R19930 vdd.n2243 vdd.n2242 0.482207
R19931 vdd.n3142 vdd.n3141 0.482207
R19932 vdd.n444 vdd.n443 0.482207
R19933 vdd.n3249 vdd.n3248 0.482207
R19934 vdd.n3148 vdd.n656 0.482207
R19935 vdd.n1807 vdd.n1038 0.482207
R19936 vdd.n1378 vdd.n1377 0.482207
R19937 vdd.n1184 vdd.n1141 0.482207
R19938 vdd.n4 vdd.n2 0.459552
R19939 vdd.n11 vdd.n9 0.459552
R19940 vdd.n317 vdd.n316 0.388379
R19941 vdd.n283 vdd.n281 0.388379
R19942 vdd.n262 vdd.n261 0.388379
R19943 vdd.n228 vdd.n226 0.388379
R19944 vdd.n219 vdd.n218 0.388379
R19945 vdd.n185 vdd.n183 0.388379
R19946 vdd.n164 vdd.n163 0.388379
R19947 vdd.n130 vdd.n128 0.388379
R19948 vdd.n122 vdd.n121 0.388379
R19949 vdd.n88 vdd.n86 0.388379
R19950 vdd.n67 vdd.n66 0.388379
R19951 vdd.n33 vdd.n31 0.388379
R19952 vdd.n1686 vdd.n1685 0.388379
R19953 vdd.n1652 vdd.n1650 0.388379
R19954 vdd.n1741 vdd.n1740 0.388379
R19955 vdd.n1707 vdd.n1705 0.388379
R19956 vdd.n1588 vdd.n1587 0.388379
R19957 vdd.n1554 vdd.n1552 0.388379
R19958 vdd.n1643 vdd.n1642 0.388379
R19959 vdd.n1609 vdd.n1607 0.388379
R19960 vdd.n1491 vdd.n1490 0.388379
R19961 vdd.n1457 vdd.n1455 0.388379
R19962 vdd.n1546 vdd.n1545 0.388379
R19963 vdd.n1512 vdd.n1510 0.388379
R19964 vdd.n19 vdd.n17 0.387128
R19965 vdd.n24 vdd.n22 0.387128
R19966 vdd.n6 vdd.n4 0.358259
R19967 vdd.n13 vdd.n11 0.358259
R19968 vdd.n268 vdd.n266 0.358259
R19969 vdd.n270 vdd.n268 0.358259
R19970 vdd.n272 vdd.n270 0.358259
R19971 vdd.n274 vdd.n272 0.358259
R19972 vdd.n276 vdd.n274 0.358259
R19973 vdd.n278 vdd.n276 0.358259
R19974 vdd.n320 vdd.n278 0.358259
R19975 vdd.n170 vdd.n168 0.358259
R19976 vdd.n172 vdd.n170 0.358259
R19977 vdd.n174 vdd.n172 0.358259
R19978 vdd.n176 vdd.n174 0.358259
R19979 vdd.n178 vdd.n176 0.358259
R19980 vdd.n180 vdd.n178 0.358259
R19981 vdd.n222 vdd.n180 0.358259
R19982 vdd.n73 vdd.n71 0.358259
R19983 vdd.n75 vdd.n73 0.358259
R19984 vdd.n77 vdd.n75 0.358259
R19985 vdd.n79 vdd.n77 0.358259
R19986 vdd.n81 vdd.n79 0.358259
R19987 vdd.n83 vdd.n81 0.358259
R19988 vdd.n125 vdd.n83 0.358259
R19989 vdd.n1744 vdd.n1702 0.358259
R19990 vdd.n1702 vdd.n1700 0.358259
R19991 vdd.n1700 vdd.n1698 0.358259
R19992 vdd.n1698 vdd.n1696 0.358259
R19993 vdd.n1696 vdd.n1694 0.358259
R19994 vdd.n1694 vdd.n1692 0.358259
R19995 vdd.n1692 vdd.n1690 0.358259
R19996 vdd.n1646 vdd.n1604 0.358259
R19997 vdd.n1604 vdd.n1602 0.358259
R19998 vdd.n1602 vdd.n1600 0.358259
R19999 vdd.n1600 vdd.n1598 0.358259
R20000 vdd.n1598 vdd.n1596 0.358259
R20001 vdd.n1596 vdd.n1594 0.358259
R20002 vdd.n1594 vdd.n1592 0.358259
R20003 vdd.n1549 vdd.n1507 0.358259
R20004 vdd.n1507 vdd.n1505 0.358259
R20005 vdd.n1505 vdd.n1503 0.358259
R20006 vdd.n1503 vdd.n1501 0.358259
R20007 vdd.n1501 vdd.n1499 0.358259
R20008 vdd.n1499 vdd.n1497 0.358259
R20009 vdd.n1497 vdd.n1495 0.358259
R20010 vdd.n14 vdd.n6 0.334552
R20011 vdd.n14 vdd.n13 0.334552
R20012 vdd.n27 vdd.n19 0.21707
R20013 vdd.n27 vdd.n24 0.21707
R20014 vdd.n318 vdd.n280 0.155672
R20015 vdd.n310 vdd.n280 0.155672
R20016 vdd.n310 vdd.n309 0.155672
R20017 vdd.n309 vdd.n285 0.155672
R20018 vdd.n302 vdd.n285 0.155672
R20019 vdd.n302 vdd.n301 0.155672
R20020 vdd.n301 vdd.n289 0.155672
R20021 vdd.n294 vdd.n289 0.155672
R20022 vdd.n263 vdd.n225 0.155672
R20023 vdd.n255 vdd.n225 0.155672
R20024 vdd.n255 vdd.n254 0.155672
R20025 vdd.n254 vdd.n230 0.155672
R20026 vdd.n247 vdd.n230 0.155672
R20027 vdd.n247 vdd.n246 0.155672
R20028 vdd.n246 vdd.n234 0.155672
R20029 vdd.n239 vdd.n234 0.155672
R20030 vdd.n220 vdd.n182 0.155672
R20031 vdd.n212 vdd.n182 0.155672
R20032 vdd.n212 vdd.n211 0.155672
R20033 vdd.n211 vdd.n187 0.155672
R20034 vdd.n204 vdd.n187 0.155672
R20035 vdd.n204 vdd.n203 0.155672
R20036 vdd.n203 vdd.n191 0.155672
R20037 vdd.n196 vdd.n191 0.155672
R20038 vdd.n165 vdd.n127 0.155672
R20039 vdd.n157 vdd.n127 0.155672
R20040 vdd.n157 vdd.n156 0.155672
R20041 vdd.n156 vdd.n132 0.155672
R20042 vdd.n149 vdd.n132 0.155672
R20043 vdd.n149 vdd.n148 0.155672
R20044 vdd.n148 vdd.n136 0.155672
R20045 vdd.n141 vdd.n136 0.155672
R20046 vdd.n123 vdd.n85 0.155672
R20047 vdd.n115 vdd.n85 0.155672
R20048 vdd.n115 vdd.n114 0.155672
R20049 vdd.n114 vdd.n90 0.155672
R20050 vdd.n107 vdd.n90 0.155672
R20051 vdd.n107 vdd.n106 0.155672
R20052 vdd.n106 vdd.n94 0.155672
R20053 vdd.n99 vdd.n94 0.155672
R20054 vdd.n68 vdd.n30 0.155672
R20055 vdd.n60 vdd.n30 0.155672
R20056 vdd.n60 vdd.n59 0.155672
R20057 vdd.n59 vdd.n35 0.155672
R20058 vdd.n52 vdd.n35 0.155672
R20059 vdd.n52 vdd.n51 0.155672
R20060 vdd.n51 vdd.n39 0.155672
R20061 vdd.n44 vdd.n39 0.155672
R20062 vdd.n1687 vdd.n1649 0.155672
R20063 vdd.n1679 vdd.n1649 0.155672
R20064 vdd.n1679 vdd.n1678 0.155672
R20065 vdd.n1678 vdd.n1654 0.155672
R20066 vdd.n1671 vdd.n1654 0.155672
R20067 vdd.n1671 vdd.n1670 0.155672
R20068 vdd.n1670 vdd.n1658 0.155672
R20069 vdd.n1663 vdd.n1658 0.155672
R20070 vdd.n1742 vdd.n1704 0.155672
R20071 vdd.n1734 vdd.n1704 0.155672
R20072 vdd.n1734 vdd.n1733 0.155672
R20073 vdd.n1733 vdd.n1709 0.155672
R20074 vdd.n1726 vdd.n1709 0.155672
R20075 vdd.n1726 vdd.n1725 0.155672
R20076 vdd.n1725 vdd.n1713 0.155672
R20077 vdd.n1718 vdd.n1713 0.155672
R20078 vdd.n1589 vdd.n1551 0.155672
R20079 vdd.n1581 vdd.n1551 0.155672
R20080 vdd.n1581 vdd.n1580 0.155672
R20081 vdd.n1580 vdd.n1556 0.155672
R20082 vdd.n1573 vdd.n1556 0.155672
R20083 vdd.n1573 vdd.n1572 0.155672
R20084 vdd.n1572 vdd.n1560 0.155672
R20085 vdd.n1565 vdd.n1560 0.155672
R20086 vdd.n1644 vdd.n1606 0.155672
R20087 vdd.n1636 vdd.n1606 0.155672
R20088 vdd.n1636 vdd.n1635 0.155672
R20089 vdd.n1635 vdd.n1611 0.155672
R20090 vdd.n1628 vdd.n1611 0.155672
R20091 vdd.n1628 vdd.n1627 0.155672
R20092 vdd.n1627 vdd.n1615 0.155672
R20093 vdd.n1620 vdd.n1615 0.155672
R20094 vdd.n1492 vdd.n1454 0.155672
R20095 vdd.n1484 vdd.n1454 0.155672
R20096 vdd.n1484 vdd.n1483 0.155672
R20097 vdd.n1483 vdd.n1459 0.155672
R20098 vdd.n1476 vdd.n1459 0.155672
R20099 vdd.n1476 vdd.n1475 0.155672
R20100 vdd.n1475 vdd.n1463 0.155672
R20101 vdd.n1468 vdd.n1463 0.155672
R20102 vdd.n1547 vdd.n1509 0.155672
R20103 vdd.n1539 vdd.n1509 0.155672
R20104 vdd.n1539 vdd.n1538 0.155672
R20105 vdd.n1538 vdd.n1514 0.155672
R20106 vdd.n1531 vdd.n1514 0.155672
R20107 vdd.n1531 vdd.n1530 0.155672
R20108 vdd.n1530 vdd.n1518 0.155672
R20109 vdd.n1523 vdd.n1518 0.155672
R20110 vdd.n2018 vdd.n1823 0.152939
R20111 vdd.n1829 vdd.n1823 0.152939
R20112 vdd.n1830 vdd.n1829 0.152939
R20113 vdd.n1831 vdd.n1830 0.152939
R20114 vdd.n1832 vdd.n1831 0.152939
R20115 vdd.n1836 vdd.n1832 0.152939
R20116 vdd.n1837 vdd.n1836 0.152939
R20117 vdd.n1838 vdd.n1837 0.152939
R20118 vdd.n1839 vdd.n1838 0.152939
R20119 vdd.n1843 vdd.n1839 0.152939
R20120 vdd.n1844 vdd.n1843 0.152939
R20121 vdd.n1845 vdd.n1844 0.152939
R20122 vdd.n1993 vdd.n1845 0.152939
R20123 vdd.n1993 vdd.n1992 0.152939
R20124 vdd.n1992 vdd.n1991 0.152939
R20125 vdd.n1991 vdd.n1851 0.152939
R20126 vdd.n1856 vdd.n1851 0.152939
R20127 vdd.n1857 vdd.n1856 0.152939
R20128 vdd.n1858 vdd.n1857 0.152939
R20129 vdd.n1862 vdd.n1858 0.152939
R20130 vdd.n1863 vdd.n1862 0.152939
R20131 vdd.n1864 vdd.n1863 0.152939
R20132 vdd.n1865 vdd.n1864 0.152939
R20133 vdd.n1869 vdd.n1865 0.152939
R20134 vdd.n1870 vdd.n1869 0.152939
R20135 vdd.n1871 vdd.n1870 0.152939
R20136 vdd.n1872 vdd.n1871 0.152939
R20137 vdd.n1876 vdd.n1872 0.152939
R20138 vdd.n1877 vdd.n1876 0.152939
R20139 vdd.n1878 vdd.n1877 0.152939
R20140 vdd.n1879 vdd.n1878 0.152939
R20141 vdd.n1883 vdd.n1879 0.152939
R20142 vdd.n1884 vdd.n1883 0.152939
R20143 vdd.n1885 vdd.n1884 0.152939
R20144 vdd.n1954 vdd.n1885 0.152939
R20145 vdd.n1954 vdd.n1953 0.152939
R20146 vdd.n1953 vdd.n1952 0.152939
R20147 vdd.n1952 vdd.n1891 0.152939
R20148 vdd.n1896 vdd.n1891 0.152939
R20149 vdd.n1897 vdd.n1896 0.152939
R20150 vdd.n1898 vdd.n1897 0.152939
R20151 vdd.n1902 vdd.n1898 0.152939
R20152 vdd.n1903 vdd.n1902 0.152939
R20153 vdd.n1904 vdd.n1903 0.152939
R20154 vdd.n1905 vdd.n1904 0.152939
R20155 vdd.n1909 vdd.n1905 0.152939
R20156 vdd.n1910 vdd.n1909 0.152939
R20157 vdd.n1911 vdd.n1910 0.152939
R20158 vdd.n1912 vdd.n1911 0.152939
R20159 vdd.n1913 vdd.n1912 0.152939
R20160 vdd.n1913 vdd.n1035 0.152939
R20161 vdd.n2242 vdd.n1817 0.152939
R20162 vdd.n1749 vdd.n1748 0.152939
R20163 vdd.n1749 vdd.n1084 0.152939
R20164 vdd.n1763 vdd.n1084 0.152939
R20165 vdd.n1764 vdd.n1763 0.152939
R20166 vdd.n1765 vdd.n1764 0.152939
R20167 vdd.n1765 vdd.n1072 0.152939
R20168 vdd.n1780 vdd.n1072 0.152939
R20169 vdd.n1781 vdd.n1780 0.152939
R20170 vdd.n1782 vdd.n1781 0.152939
R20171 vdd.n1782 vdd.n1061 0.152939
R20172 vdd.n1797 vdd.n1061 0.152939
R20173 vdd.n1798 vdd.n1797 0.152939
R20174 vdd.n1799 vdd.n1798 0.152939
R20175 vdd.n1799 vdd.n1049 0.152939
R20176 vdd.n1815 vdd.n1049 0.152939
R20177 vdd.n1816 vdd.n1815 0.152939
R20178 vdd.n2243 vdd.n1816 0.152939
R20179 vdd.n670 vdd.n667 0.152939
R20180 vdd.n671 vdd.n670 0.152939
R20181 vdd.n672 vdd.n671 0.152939
R20182 vdd.n673 vdd.n672 0.152939
R20183 vdd.n676 vdd.n673 0.152939
R20184 vdd.n677 vdd.n676 0.152939
R20185 vdd.n678 vdd.n677 0.152939
R20186 vdd.n679 vdd.n678 0.152939
R20187 vdd.n682 vdd.n679 0.152939
R20188 vdd.n683 vdd.n682 0.152939
R20189 vdd.n684 vdd.n683 0.152939
R20190 vdd.n685 vdd.n684 0.152939
R20191 vdd.n690 vdd.n685 0.152939
R20192 vdd.n691 vdd.n690 0.152939
R20193 vdd.n692 vdd.n691 0.152939
R20194 vdd.n693 vdd.n692 0.152939
R20195 vdd.n696 vdd.n693 0.152939
R20196 vdd.n697 vdd.n696 0.152939
R20197 vdd.n698 vdd.n697 0.152939
R20198 vdd.n699 vdd.n698 0.152939
R20199 vdd.n702 vdd.n699 0.152939
R20200 vdd.n703 vdd.n702 0.152939
R20201 vdd.n704 vdd.n703 0.152939
R20202 vdd.n705 vdd.n704 0.152939
R20203 vdd.n708 vdd.n705 0.152939
R20204 vdd.n709 vdd.n708 0.152939
R20205 vdd.n710 vdd.n709 0.152939
R20206 vdd.n711 vdd.n710 0.152939
R20207 vdd.n714 vdd.n711 0.152939
R20208 vdd.n715 vdd.n714 0.152939
R20209 vdd.n716 vdd.n715 0.152939
R20210 vdd.n717 vdd.n716 0.152939
R20211 vdd.n720 vdd.n717 0.152939
R20212 vdd.n721 vdd.n720 0.152939
R20213 vdd.n3058 vdd.n721 0.152939
R20214 vdd.n3058 vdd.n3057 0.152939
R20215 vdd.n3057 vdd.n3056 0.152939
R20216 vdd.n3056 vdd.n725 0.152939
R20217 vdd.n730 vdd.n725 0.152939
R20218 vdd.n731 vdd.n730 0.152939
R20219 vdd.n734 vdd.n731 0.152939
R20220 vdd.n735 vdd.n734 0.152939
R20221 vdd.n736 vdd.n735 0.152939
R20222 vdd.n737 vdd.n736 0.152939
R20223 vdd.n740 vdd.n737 0.152939
R20224 vdd.n741 vdd.n740 0.152939
R20225 vdd.n742 vdd.n741 0.152939
R20226 vdd.n743 vdd.n742 0.152939
R20227 vdd.n746 vdd.n743 0.152939
R20228 vdd.n747 vdd.n746 0.152939
R20229 vdd.n748 vdd.n747 0.152939
R20230 vdd.n3141 vdd.n661 0.152939
R20231 vdd.n3142 vdd.n651 0.152939
R20232 vdd.n3156 vdd.n651 0.152939
R20233 vdd.n3157 vdd.n3156 0.152939
R20234 vdd.n3158 vdd.n3157 0.152939
R20235 vdd.n3158 vdd.n639 0.152939
R20236 vdd.n3172 vdd.n639 0.152939
R20237 vdd.n3173 vdd.n3172 0.152939
R20238 vdd.n3174 vdd.n3173 0.152939
R20239 vdd.n3174 vdd.n627 0.152939
R20240 vdd.n3189 vdd.n627 0.152939
R20241 vdd.n3190 vdd.n3189 0.152939
R20242 vdd.n3191 vdd.n3190 0.152939
R20243 vdd.n3191 vdd.n616 0.152939
R20244 vdd.n3208 vdd.n616 0.152939
R20245 vdd.n3209 vdd.n3208 0.152939
R20246 vdd.n3210 vdd.n3209 0.152939
R20247 vdd.n3210 vdd.n322 0.152939
R20248 vdd.n3290 vdd.n323 0.152939
R20249 vdd.n334 vdd.n323 0.152939
R20250 vdd.n335 vdd.n334 0.152939
R20251 vdd.n336 vdd.n335 0.152939
R20252 vdd.n343 vdd.n336 0.152939
R20253 vdd.n344 vdd.n343 0.152939
R20254 vdd.n345 vdd.n344 0.152939
R20255 vdd.n346 vdd.n345 0.152939
R20256 vdd.n354 vdd.n346 0.152939
R20257 vdd.n355 vdd.n354 0.152939
R20258 vdd.n356 vdd.n355 0.152939
R20259 vdd.n357 vdd.n356 0.152939
R20260 vdd.n365 vdd.n357 0.152939
R20261 vdd.n366 vdd.n365 0.152939
R20262 vdd.n367 vdd.n366 0.152939
R20263 vdd.n368 vdd.n367 0.152939
R20264 vdd.n443 vdd.n368 0.152939
R20265 vdd.n444 vdd.n442 0.152939
R20266 vdd.n451 vdd.n442 0.152939
R20267 vdd.n452 vdd.n451 0.152939
R20268 vdd.n453 vdd.n452 0.152939
R20269 vdd.n453 vdd.n440 0.152939
R20270 vdd.n461 vdd.n440 0.152939
R20271 vdd.n462 vdd.n461 0.152939
R20272 vdd.n463 vdd.n462 0.152939
R20273 vdd.n463 vdd.n438 0.152939
R20274 vdd.n471 vdd.n438 0.152939
R20275 vdd.n472 vdd.n471 0.152939
R20276 vdd.n473 vdd.n472 0.152939
R20277 vdd.n473 vdd.n436 0.152939
R20278 vdd.n481 vdd.n436 0.152939
R20279 vdd.n482 vdd.n481 0.152939
R20280 vdd.n483 vdd.n482 0.152939
R20281 vdd.n483 vdd.n434 0.152939
R20282 vdd.n491 vdd.n434 0.152939
R20283 vdd.n492 vdd.n491 0.152939
R20284 vdd.n493 vdd.n492 0.152939
R20285 vdd.n493 vdd.n430 0.152939
R20286 vdd.n501 vdd.n430 0.152939
R20287 vdd.n502 vdd.n501 0.152939
R20288 vdd.n503 vdd.n502 0.152939
R20289 vdd.n503 vdd.n428 0.152939
R20290 vdd.n511 vdd.n428 0.152939
R20291 vdd.n512 vdd.n511 0.152939
R20292 vdd.n513 vdd.n512 0.152939
R20293 vdd.n513 vdd.n426 0.152939
R20294 vdd.n521 vdd.n426 0.152939
R20295 vdd.n522 vdd.n521 0.152939
R20296 vdd.n523 vdd.n522 0.152939
R20297 vdd.n523 vdd.n424 0.152939
R20298 vdd.n531 vdd.n424 0.152939
R20299 vdd.n532 vdd.n531 0.152939
R20300 vdd.n533 vdd.n532 0.152939
R20301 vdd.n533 vdd.n422 0.152939
R20302 vdd.n541 vdd.n422 0.152939
R20303 vdd.n542 vdd.n541 0.152939
R20304 vdd.n543 vdd.n542 0.152939
R20305 vdd.n543 vdd.n418 0.152939
R20306 vdd.n551 vdd.n418 0.152939
R20307 vdd.n552 vdd.n551 0.152939
R20308 vdd.n553 vdd.n552 0.152939
R20309 vdd.n553 vdd.n416 0.152939
R20310 vdd.n561 vdd.n416 0.152939
R20311 vdd.n562 vdd.n561 0.152939
R20312 vdd.n563 vdd.n562 0.152939
R20313 vdd.n563 vdd.n414 0.152939
R20314 vdd.n571 vdd.n414 0.152939
R20315 vdd.n572 vdd.n571 0.152939
R20316 vdd.n573 vdd.n572 0.152939
R20317 vdd.n573 vdd.n412 0.152939
R20318 vdd.n581 vdd.n412 0.152939
R20319 vdd.n582 vdd.n581 0.152939
R20320 vdd.n583 vdd.n582 0.152939
R20321 vdd.n583 vdd.n410 0.152939
R20322 vdd.n591 vdd.n410 0.152939
R20323 vdd.n592 vdd.n591 0.152939
R20324 vdd.n593 vdd.n592 0.152939
R20325 vdd.n593 vdd.n408 0.152939
R20326 vdd.n600 vdd.n408 0.152939
R20327 vdd.n3249 vdd.n600 0.152939
R20328 vdd.n3149 vdd.n3148 0.152939
R20329 vdd.n3150 vdd.n3149 0.152939
R20330 vdd.n3150 vdd.n645 0.152939
R20331 vdd.n3164 vdd.n645 0.152939
R20332 vdd.n3165 vdd.n3164 0.152939
R20333 vdd.n3166 vdd.n3165 0.152939
R20334 vdd.n3166 vdd.n632 0.152939
R20335 vdd.n3180 vdd.n632 0.152939
R20336 vdd.n3181 vdd.n3180 0.152939
R20337 vdd.n3182 vdd.n3181 0.152939
R20338 vdd.n3182 vdd.n621 0.152939
R20339 vdd.n3197 vdd.n621 0.152939
R20340 vdd.n3198 vdd.n3197 0.152939
R20341 vdd.n3199 vdd.n3198 0.152939
R20342 vdd.n3201 vdd.n3199 0.152939
R20343 vdd.n3201 vdd.n3200 0.152939
R20344 vdd.n3200 vdd.n611 0.152939
R20345 vdd.n611 vdd.n609 0.152939
R20346 vdd.n3219 vdd.n609 0.152939
R20347 vdd.n3220 vdd.n3219 0.152939
R20348 vdd.n3221 vdd.n3220 0.152939
R20349 vdd.n3221 vdd.n607 0.152939
R20350 vdd.n3226 vdd.n607 0.152939
R20351 vdd.n3227 vdd.n3226 0.152939
R20352 vdd.n3228 vdd.n3227 0.152939
R20353 vdd.n3228 vdd.n605 0.152939
R20354 vdd.n3233 vdd.n605 0.152939
R20355 vdd.n3234 vdd.n3233 0.152939
R20356 vdd.n3235 vdd.n3234 0.152939
R20357 vdd.n3235 vdd.n603 0.152939
R20358 vdd.n3241 vdd.n603 0.152939
R20359 vdd.n3242 vdd.n3241 0.152939
R20360 vdd.n3243 vdd.n3242 0.152939
R20361 vdd.n3243 vdd.n601 0.152939
R20362 vdd.n3248 vdd.n601 0.152939
R20363 vdd.n3011 vdd.n656 0.152939
R20364 vdd.n2254 vdd.n1038 0.152939
R20365 vdd.n1379 vdd.n1378 0.152939
R20366 vdd.n1379 vdd.n1135 0.152939
R20367 vdd.n1393 vdd.n1135 0.152939
R20368 vdd.n1394 vdd.n1393 0.152939
R20369 vdd.n1395 vdd.n1394 0.152939
R20370 vdd.n1395 vdd.n1123 0.152939
R20371 vdd.n1410 vdd.n1123 0.152939
R20372 vdd.n1411 vdd.n1410 0.152939
R20373 vdd.n1412 vdd.n1411 0.152939
R20374 vdd.n1412 vdd.n1113 0.152939
R20375 vdd.n1427 vdd.n1113 0.152939
R20376 vdd.n1428 vdd.n1427 0.152939
R20377 vdd.n1429 vdd.n1428 0.152939
R20378 vdd.n1429 vdd.n1100 0.152939
R20379 vdd.n1443 vdd.n1100 0.152939
R20380 vdd.n1444 vdd.n1443 0.152939
R20381 vdd.n1445 vdd.n1444 0.152939
R20382 vdd.n1445 vdd.n1089 0.152939
R20383 vdd.n1755 vdd.n1089 0.152939
R20384 vdd.n1756 vdd.n1755 0.152939
R20385 vdd.n1757 vdd.n1756 0.152939
R20386 vdd.n1757 vdd.n1078 0.152939
R20387 vdd.n1771 vdd.n1078 0.152939
R20388 vdd.n1772 vdd.n1771 0.152939
R20389 vdd.n1773 vdd.n1772 0.152939
R20390 vdd.n1773 vdd.n1066 0.152939
R20391 vdd.n1788 vdd.n1066 0.152939
R20392 vdd.n1789 vdd.n1788 0.152939
R20393 vdd.n1790 vdd.n1789 0.152939
R20394 vdd.n1790 vdd.n1056 0.152939
R20395 vdd.n1805 vdd.n1056 0.152939
R20396 vdd.n1806 vdd.n1805 0.152939
R20397 vdd.n1809 vdd.n1806 0.152939
R20398 vdd.n1809 vdd.n1808 0.152939
R20399 vdd.n1808 vdd.n1807 0.152939
R20400 vdd.n1369 vdd.n1184 0.152939
R20401 vdd.n1369 vdd.n1368 0.152939
R20402 vdd.n1368 vdd.n1367 0.152939
R20403 vdd.n1367 vdd.n1186 0.152939
R20404 vdd.n1363 vdd.n1186 0.152939
R20405 vdd.n1363 vdd.n1362 0.152939
R20406 vdd.n1362 vdd.n1361 0.152939
R20407 vdd.n1361 vdd.n1191 0.152939
R20408 vdd.n1357 vdd.n1191 0.152939
R20409 vdd.n1357 vdd.n1356 0.152939
R20410 vdd.n1356 vdd.n1355 0.152939
R20411 vdd.n1355 vdd.n1197 0.152939
R20412 vdd.n1351 vdd.n1197 0.152939
R20413 vdd.n1351 vdd.n1350 0.152939
R20414 vdd.n1350 vdd.n1349 0.152939
R20415 vdd.n1349 vdd.n1203 0.152939
R20416 vdd.n1345 vdd.n1203 0.152939
R20417 vdd.n1345 vdd.n1344 0.152939
R20418 vdd.n1344 vdd.n1343 0.152939
R20419 vdd.n1343 vdd.n1209 0.152939
R20420 vdd.n1335 vdd.n1209 0.152939
R20421 vdd.n1335 vdd.n1334 0.152939
R20422 vdd.n1334 vdd.n1333 0.152939
R20423 vdd.n1333 vdd.n1213 0.152939
R20424 vdd.n1329 vdd.n1213 0.152939
R20425 vdd.n1329 vdd.n1328 0.152939
R20426 vdd.n1328 vdd.n1327 0.152939
R20427 vdd.n1327 vdd.n1219 0.152939
R20428 vdd.n1323 vdd.n1219 0.152939
R20429 vdd.n1323 vdd.n1322 0.152939
R20430 vdd.n1322 vdd.n1321 0.152939
R20431 vdd.n1321 vdd.n1225 0.152939
R20432 vdd.n1317 vdd.n1225 0.152939
R20433 vdd.n1317 vdd.n1316 0.152939
R20434 vdd.n1316 vdd.n1315 0.152939
R20435 vdd.n1315 vdd.n1231 0.152939
R20436 vdd.n1311 vdd.n1231 0.152939
R20437 vdd.n1311 vdd.n1310 0.152939
R20438 vdd.n1310 vdd.n1309 0.152939
R20439 vdd.n1309 vdd.n1237 0.152939
R20440 vdd.n1302 vdd.n1237 0.152939
R20441 vdd.n1302 vdd.n1301 0.152939
R20442 vdd.n1301 vdd.n1300 0.152939
R20443 vdd.n1300 vdd.n1242 0.152939
R20444 vdd.n1296 vdd.n1242 0.152939
R20445 vdd.n1296 vdd.n1295 0.152939
R20446 vdd.n1295 vdd.n1294 0.152939
R20447 vdd.n1294 vdd.n1248 0.152939
R20448 vdd.n1290 vdd.n1248 0.152939
R20449 vdd.n1290 vdd.n1289 0.152939
R20450 vdd.n1289 vdd.n1288 0.152939
R20451 vdd.n1288 vdd.n1254 0.152939
R20452 vdd.n1284 vdd.n1254 0.152939
R20453 vdd.n1284 vdd.n1283 0.152939
R20454 vdd.n1283 vdd.n1282 0.152939
R20455 vdd.n1282 vdd.n1260 0.152939
R20456 vdd.n1278 vdd.n1260 0.152939
R20457 vdd.n1278 vdd.n1277 0.152939
R20458 vdd.n1277 vdd.n1276 0.152939
R20459 vdd.n1276 vdd.n1266 0.152939
R20460 vdd.n1272 vdd.n1266 0.152939
R20461 vdd.n1272 vdd.n1147 0.152939
R20462 vdd.n1377 vdd.n1147 0.152939
R20463 vdd.n1385 vdd.n1141 0.152939
R20464 vdd.n1386 vdd.n1385 0.152939
R20465 vdd.n1387 vdd.n1386 0.152939
R20466 vdd.n1387 vdd.n1129 0.152939
R20467 vdd.n1402 vdd.n1129 0.152939
R20468 vdd.n1403 vdd.n1402 0.152939
R20469 vdd.n1404 vdd.n1403 0.152939
R20470 vdd.n1404 vdd.n1118 0.152939
R20471 vdd.n1419 vdd.n1118 0.152939
R20472 vdd.n1420 vdd.n1419 0.152939
R20473 vdd.n1421 vdd.n1420 0.152939
R20474 vdd.n1421 vdd.n1107 0.152939
R20475 vdd.n1435 vdd.n1107 0.152939
R20476 vdd.n1436 vdd.n1435 0.152939
R20477 vdd.n1437 vdd.n1436 0.152939
R20478 vdd.n1437 vdd.n1095 0.152939
R20479 vdd.n1452 vdd.n1095 0.152939
R20480 vdd.n2232 vdd.n1817 0.110256
R20481 vdd.n2942 vdd.n661 0.110256
R20482 vdd.n3011 vdd.n3010 0.110256
R20483 vdd.n2255 vdd.n2254 0.110256
R20484 vdd.n1748 vdd.n1747 0.0695946
R20485 vdd.n3291 vdd.n322 0.0695946
R20486 vdd.n3291 vdd.n3290 0.0695946
R20487 vdd.n1747 vdd.n1452 0.0695946
R20488 vdd.n2232 vdd.n2018 0.0431829
R20489 vdd.n2255 vdd.n1035 0.0431829
R20490 vdd.n2942 vdd.n667 0.0431829
R20491 vdd.n3010 vdd.n748 0.0431829
R20492 vdd vdd.n28 0.00833333
R20493 CSoutput.n19 CSoutput.t180 184.661
R20494 CSoutput.n78 CSoutput.n77 165.8
R20495 CSoutput.n76 CSoutput.n0 165.8
R20496 CSoutput.n75 CSoutput.n74 165.8
R20497 CSoutput.n73 CSoutput.n72 165.8
R20498 CSoutput.n71 CSoutput.n2 165.8
R20499 CSoutput.n69 CSoutput.n68 165.8
R20500 CSoutput.n67 CSoutput.n3 165.8
R20501 CSoutput.n66 CSoutput.n65 165.8
R20502 CSoutput.n63 CSoutput.n4 165.8
R20503 CSoutput.n61 CSoutput.n60 165.8
R20504 CSoutput.n59 CSoutput.n5 165.8
R20505 CSoutput.n58 CSoutput.n57 165.8
R20506 CSoutput.n55 CSoutput.n6 165.8
R20507 CSoutput.n54 CSoutput.n53 165.8
R20508 CSoutput.n52 CSoutput.n51 165.8
R20509 CSoutput.n50 CSoutput.n8 165.8
R20510 CSoutput.n48 CSoutput.n47 165.8
R20511 CSoutput.n46 CSoutput.n9 165.8
R20512 CSoutput.n45 CSoutput.n44 165.8
R20513 CSoutput.n42 CSoutput.n10 165.8
R20514 CSoutput.n41 CSoutput.n40 165.8
R20515 CSoutput.n39 CSoutput.n38 165.8
R20516 CSoutput.n37 CSoutput.n12 165.8
R20517 CSoutput.n35 CSoutput.n34 165.8
R20518 CSoutput.n33 CSoutput.n13 165.8
R20519 CSoutput.n32 CSoutput.n31 165.8
R20520 CSoutput.n29 CSoutput.n14 165.8
R20521 CSoutput.n28 CSoutput.n27 165.8
R20522 CSoutput.n26 CSoutput.n25 165.8
R20523 CSoutput.n24 CSoutput.n16 165.8
R20524 CSoutput.n22 CSoutput.n21 165.8
R20525 CSoutput.n20 CSoutput.n17 165.8
R20526 CSoutput.n77 CSoutput.t183 162.194
R20527 CSoutput.n18 CSoutput.t177 120.501
R20528 CSoutput.n23 CSoutput.t194 120.501
R20529 CSoutput.n15 CSoutput.t189 120.501
R20530 CSoutput.n30 CSoutput.t178 120.501
R20531 CSoutput.n36 CSoutput.t179 120.501
R20532 CSoutput.n11 CSoutput.t191 120.501
R20533 CSoutput.n43 CSoutput.t188 120.501
R20534 CSoutput.n49 CSoutput.t182 120.501
R20535 CSoutput.n7 CSoutput.t195 120.501
R20536 CSoutput.n56 CSoutput.t196 120.501
R20537 CSoutput.n62 CSoutput.t185 120.501
R20538 CSoutput.n64 CSoutput.t197 120.501
R20539 CSoutput.n70 CSoutput.t176 120.501
R20540 CSoutput.n1 CSoutput.t193 120.501
R20541 CSoutput.n310 CSoutput.n308 103.469
R20542 CSoutput.n294 CSoutput.n292 103.469
R20543 CSoutput.n279 CSoutput.n277 103.469
R20544 CSoutput.n112 CSoutput.n110 103.469
R20545 CSoutput.n96 CSoutput.n94 103.469
R20546 CSoutput.n81 CSoutput.n79 103.469
R20547 CSoutput.n320 CSoutput.n319 103.111
R20548 CSoutput.n318 CSoutput.n317 103.111
R20549 CSoutput.n316 CSoutput.n315 103.111
R20550 CSoutput.n314 CSoutput.n313 103.111
R20551 CSoutput.n312 CSoutput.n311 103.111
R20552 CSoutput.n310 CSoutput.n309 103.111
R20553 CSoutput.n306 CSoutput.n305 103.111
R20554 CSoutput.n304 CSoutput.n303 103.111
R20555 CSoutput.n302 CSoutput.n301 103.111
R20556 CSoutput.n300 CSoutput.n299 103.111
R20557 CSoutput.n298 CSoutput.n297 103.111
R20558 CSoutput.n296 CSoutput.n295 103.111
R20559 CSoutput.n294 CSoutput.n293 103.111
R20560 CSoutput.n291 CSoutput.n290 103.111
R20561 CSoutput.n289 CSoutput.n288 103.111
R20562 CSoutput.n287 CSoutput.n286 103.111
R20563 CSoutput.n285 CSoutput.n284 103.111
R20564 CSoutput.n283 CSoutput.n282 103.111
R20565 CSoutput.n281 CSoutput.n280 103.111
R20566 CSoutput.n279 CSoutput.n278 103.111
R20567 CSoutput.n112 CSoutput.n111 103.111
R20568 CSoutput.n114 CSoutput.n113 103.111
R20569 CSoutput.n116 CSoutput.n115 103.111
R20570 CSoutput.n118 CSoutput.n117 103.111
R20571 CSoutput.n120 CSoutput.n119 103.111
R20572 CSoutput.n122 CSoutput.n121 103.111
R20573 CSoutput.n124 CSoutput.n123 103.111
R20574 CSoutput.n96 CSoutput.n95 103.111
R20575 CSoutput.n98 CSoutput.n97 103.111
R20576 CSoutput.n100 CSoutput.n99 103.111
R20577 CSoutput.n102 CSoutput.n101 103.111
R20578 CSoutput.n104 CSoutput.n103 103.111
R20579 CSoutput.n106 CSoutput.n105 103.111
R20580 CSoutput.n108 CSoutput.n107 103.111
R20581 CSoutput.n81 CSoutput.n80 103.111
R20582 CSoutput.n83 CSoutput.n82 103.111
R20583 CSoutput.n85 CSoutput.n84 103.111
R20584 CSoutput.n87 CSoutput.n86 103.111
R20585 CSoutput.n89 CSoutput.n88 103.111
R20586 CSoutput.n91 CSoutput.n90 103.111
R20587 CSoutput.n93 CSoutput.n92 103.111
R20588 CSoutput.n322 CSoutput.n321 103.111
R20589 CSoutput.n346 CSoutput.n344 81.5057
R20590 CSoutput.n327 CSoutput.n325 81.5057
R20591 CSoutput.n386 CSoutput.n384 81.5057
R20592 CSoutput.n367 CSoutput.n365 81.5057
R20593 CSoutput.n362 CSoutput.n361 80.9324
R20594 CSoutput.n360 CSoutput.n359 80.9324
R20595 CSoutput.n358 CSoutput.n357 80.9324
R20596 CSoutput.n356 CSoutput.n355 80.9324
R20597 CSoutput.n354 CSoutput.n353 80.9324
R20598 CSoutput.n352 CSoutput.n351 80.9324
R20599 CSoutput.n350 CSoutput.n349 80.9324
R20600 CSoutput.n348 CSoutput.n347 80.9324
R20601 CSoutput.n346 CSoutput.n345 80.9324
R20602 CSoutput.n343 CSoutput.n342 80.9324
R20603 CSoutput.n341 CSoutput.n340 80.9324
R20604 CSoutput.n339 CSoutput.n338 80.9324
R20605 CSoutput.n337 CSoutput.n336 80.9324
R20606 CSoutput.n335 CSoutput.n334 80.9324
R20607 CSoutput.n333 CSoutput.n332 80.9324
R20608 CSoutput.n331 CSoutput.n330 80.9324
R20609 CSoutput.n329 CSoutput.n328 80.9324
R20610 CSoutput.n327 CSoutput.n326 80.9324
R20611 CSoutput.n386 CSoutput.n385 80.9324
R20612 CSoutput.n388 CSoutput.n387 80.9324
R20613 CSoutput.n390 CSoutput.n389 80.9324
R20614 CSoutput.n392 CSoutput.n391 80.9324
R20615 CSoutput.n394 CSoutput.n393 80.9324
R20616 CSoutput.n396 CSoutput.n395 80.9324
R20617 CSoutput.n398 CSoutput.n397 80.9324
R20618 CSoutput.n400 CSoutput.n399 80.9324
R20619 CSoutput.n402 CSoutput.n401 80.9324
R20620 CSoutput.n367 CSoutput.n366 80.9324
R20621 CSoutput.n369 CSoutput.n368 80.9324
R20622 CSoutput.n371 CSoutput.n370 80.9324
R20623 CSoutput.n373 CSoutput.n372 80.9324
R20624 CSoutput.n375 CSoutput.n374 80.9324
R20625 CSoutput.n377 CSoutput.n376 80.9324
R20626 CSoutput.n379 CSoutput.n378 80.9324
R20627 CSoutput.n381 CSoutput.n380 80.9324
R20628 CSoutput.n383 CSoutput.n382 80.9324
R20629 CSoutput.n25 CSoutput.n24 48.1486
R20630 CSoutput.n69 CSoutput.n3 48.1486
R20631 CSoutput.n38 CSoutput.n37 48.1486
R20632 CSoutput.n42 CSoutput.n41 48.1486
R20633 CSoutput.n51 CSoutput.n50 48.1486
R20634 CSoutput.n55 CSoutput.n54 48.1486
R20635 CSoutput.n22 CSoutput.n17 46.462
R20636 CSoutput.n72 CSoutput.n71 46.462
R20637 CSoutput.n20 CSoutput.n19 44.9055
R20638 CSoutput.n29 CSoutput.n28 43.7635
R20639 CSoutput.n65 CSoutput.n63 43.7635
R20640 CSoutput.n35 CSoutput.n13 41.7396
R20641 CSoutput.n57 CSoutput.n5 41.7396
R20642 CSoutput.n44 CSoutput.n9 37.0171
R20643 CSoutput.n48 CSoutput.n9 37.0171
R20644 CSoutput.n76 CSoutput.n75 34.9932
R20645 CSoutput.n31 CSoutput.n13 32.2947
R20646 CSoutput.n61 CSoutput.n5 32.2947
R20647 CSoutput.n30 CSoutput.n29 29.6014
R20648 CSoutput.n63 CSoutput.n62 29.6014
R20649 CSoutput.n19 CSoutput.n18 28.4085
R20650 CSoutput.n18 CSoutput.n17 25.1176
R20651 CSoutput.n72 CSoutput.n1 25.1176
R20652 CSoutput.n43 CSoutput.n42 22.0922
R20653 CSoutput.n50 CSoutput.n49 22.0922
R20654 CSoutput.n77 CSoutput.n76 21.8586
R20655 CSoutput.n37 CSoutput.n36 18.9681
R20656 CSoutput.n56 CSoutput.n55 18.9681
R20657 CSoutput.n25 CSoutput.n15 17.6292
R20658 CSoutput.n64 CSoutput.n3 17.6292
R20659 CSoutput.n24 CSoutput.n23 15.844
R20660 CSoutput.n70 CSoutput.n69 15.844
R20661 CSoutput.n38 CSoutput.n11 14.5051
R20662 CSoutput.n54 CSoutput.n7 14.5051
R20663 CSoutput.n405 CSoutput.n78 11.6139
R20664 CSoutput.n41 CSoutput.n11 11.3811
R20665 CSoutput.n51 CSoutput.n7 11.3811
R20666 CSoutput.n23 CSoutput.n22 10.0422
R20667 CSoutput.n71 CSoutput.n70 10.0422
R20668 CSoutput.n307 CSoutput.n291 9.25285
R20669 CSoutput.n109 CSoutput.n93 9.25285
R20670 CSoutput.n364 CSoutput.n324 9.1987
R20671 CSoutput.n363 CSoutput.n343 8.97993
R20672 CSoutput.n403 CSoutput.n383 8.97993
R20673 CSoutput.n28 CSoutput.n15 8.25698
R20674 CSoutput.n65 CSoutput.n64 8.25698
R20675 CSoutput.n364 CSoutput.n363 7.89345
R20676 CSoutput.n404 CSoutput.n403 7.89345
R20677 CSoutput.n324 CSoutput.n323 7.12641
R20678 CSoutput.n126 CSoutput.n125 7.12641
R20679 CSoutput.n36 CSoutput.n35 6.91809
R20680 CSoutput.n57 CSoutput.n56 6.91809
R20681 CSoutput.n405 CSoutput.n126 5.60626
R20682 CSoutput.n363 CSoutput.n362 5.25266
R20683 CSoutput.n403 CSoutput.n402 5.25266
R20684 CSoutput.n323 CSoutput.n322 5.1449
R20685 CSoutput.n307 CSoutput.n306 5.1449
R20686 CSoutput.n125 CSoutput.n124 5.1449
R20687 CSoutput.n109 CSoutput.n108 5.1449
R20688 CSoutput.n217 CSoutput.n170 4.5005
R20689 CSoutput.n186 CSoutput.n170 4.5005
R20690 CSoutput.n181 CSoutput.n165 4.5005
R20691 CSoutput.n181 CSoutput.n167 4.5005
R20692 CSoutput.n181 CSoutput.n164 4.5005
R20693 CSoutput.n181 CSoutput.n168 4.5005
R20694 CSoutput.n181 CSoutput.n163 4.5005
R20695 CSoutput.n181 CSoutput.t184 4.5005
R20696 CSoutput.n181 CSoutput.n162 4.5005
R20697 CSoutput.n181 CSoutput.n169 4.5005
R20698 CSoutput.n181 CSoutput.n170 4.5005
R20699 CSoutput.n179 CSoutput.n165 4.5005
R20700 CSoutput.n179 CSoutput.n167 4.5005
R20701 CSoutput.n179 CSoutput.n164 4.5005
R20702 CSoutput.n179 CSoutput.n168 4.5005
R20703 CSoutput.n179 CSoutput.n163 4.5005
R20704 CSoutput.n179 CSoutput.t184 4.5005
R20705 CSoutput.n179 CSoutput.n162 4.5005
R20706 CSoutput.n179 CSoutput.n169 4.5005
R20707 CSoutput.n179 CSoutput.n170 4.5005
R20708 CSoutput.n178 CSoutput.n165 4.5005
R20709 CSoutput.n178 CSoutput.n167 4.5005
R20710 CSoutput.n178 CSoutput.n164 4.5005
R20711 CSoutput.n178 CSoutput.n168 4.5005
R20712 CSoutput.n178 CSoutput.n163 4.5005
R20713 CSoutput.n178 CSoutput.t184 4.5005
R20714 CSoutput.n178 CSoutput.n162 4.5005
R20715 CSoutput.n178 CSoutput.n169 4.5005
R20716 CSoutput.n178 CSoutput.n170 4.5005
R20717 CSoutput.n263 CSoutput.n165 4.5005
R20718 CSoutput.n263 CSoutput.n167 4.5005
R20719 CSoutput.n263 CSoutput.n164 4.5005
R20720 CSoutput.n263 CSoutput.n168 4.5005
R20721 CSoutput.n263 CSoutput.n163 4.5005
R20722 CSoutput.n263 CSoutput.t184 4.5005
R20723 CSoutput.n263 CSoutput.n162 4.5005
R20724 CSoutput.n263 CSoutput.n169 4.5005
R20725 CSoutput.n263 CSoutput.n170 4.5005
R20726 CSoutput.n261 CSoutput.n165 4.5005
R20727 CSoutput.n261 CSoutput.n167 4.5005
R20728 CSoutput.n261 CSoutput.n164 4.5005
R20729 CSoutput.n261 CSoutput.n168 4.5005
R20730 CSoutput.n261 CSoutput.n163 4.5005
R20731 CSoutput.n261 CSoutput.t184 4.5005
R20732 CSoutput.n261 CSoutput.n162 4.5005
R20733 CSoutput.n261 CSoutput.n169 4.5005
R20734 CSoutput.n259 CSoutput.n165 4.5005
R20735 CSoutput.n259 CSoutput.n167 4.5005
R20736 CSoutput.n259 CSoutput.n164 4.5005
R20737 CSoutput.n259 CSoutput.n168 4.5005
R20738 CSoutput.n259 CSoutput.n163 4.5005
R20739 CSoutput.n259 CSoutput.t184 4.5005
R20740 CSoutput.n259 CSoutput.n162 4.5005
R20741 CSoutput.n259 CSoutput.n169 4.5005
R20742 CSoutput.n189 CSoutput.n165 4.5005
R20743 CSoutput.n189 CSoutput.n167 4.5005
R20744 CSoutput.n189 CSoutput.n164 4.5005
R20745 CSoutput.n189 CSoutput.n168 4.5005
R20746 CSoutput.n189 CSoutput.n163 4.5005
R20747 CSoutput.n189 CSoutput.t184 4.5005
R20748 CSoutput.n189 CSoutput.n162 4.5005
R20749 CSoutput.n189 CSoutput.n169 4.5005
R20750 CSoutput.n189 CSoutput.n170 4.5005
R20751 CSoutput.n188 CSoutput.n165 4.5005
R20752 CSoutput.n188 CSoutput.n167 4.5005
R20753 CSoutput.n188 CSoutput.n164 4.5005
R20754 CSoutput.n188 CSoutput.n168 4.5005
R20755 CSoutput.n188 CSoutput.n163 4.5005
R20756 CSoutput.n188 CSoutput.t184 4.5005
R20757 CSoutput.n188 CSoutput.n162 4.5005
R20758 CSoutput.n188 CSoutput.n169 4.5005
R20759 CSoutput.n188 CSoutput.n170 4.5005
R20760 CSoutput.n192 CSoutput.n165 4.5005
R20761 CSoutput.n192 CSoutput.n167 4.5005
R20762 CSoutput.n192 CSoutput.n164 4.5005
R20763 CSoutput.n192 CSoutput.n168 4.5005
R20764 CSoutput.n192 CSoutput.n163 4.5005
R20765 CSoutput.n192 CSoutput.t184 4.5005
R20766 CSoutput.n192 CSoutput.n162 4.5005
R20767 CSoutput.n192 CSoutput.n169 4.5005
R20768 CSoutput.n192 CSoutput.n170 4.5005
R20769 CSoutput.n191 CSoutput.n165 4.5005
R20770 CSoutput.n191 CSoutput.n167 4.5005
R20771 CSoutput.n191 CSoutput.n164 4.5005
R20772 CSoutput.n191 CSoutput.n168 4.5005
R20773 CSoutput.n191 CSoutput.n163 4.5005
R20774 CSoutput.n191 CSoutput.t184 4.5005
R20775 CSoutput.n191 CSoutput.n162 4.5005
R20776 CSoutput.n191 CSoutput.n169 4.5005
R20777 CSoutput.n191 CSoutput.n170 4.5005
R20778 CSoutput.n174 CSoutput.n165 4.5005
R20779 CSoutput.n174 CSoutput.n167 4.5005
R20780 CSoutput.n174 CSoutput.n164 4.5005
R20781 CSoutput.n174 CSoutput.n168 4.5005
R20782 CSoutput.n174 CSoutput.n163 4.5005
R20783 CSoutput.n174 CSoutput.t184 4.5005
R20784 CSoutput.n174 CSoutput.n162 4.5005
R20785 CSoutput.n174 CSoutput.n169 4.5005
R20786 CSoutput.n174 CSoutput.n170 4.5005
R20787 CSoutput.n266 CSoutput.n165 4.5005
R20788 CSoutput.n266 CSoutput.n167 4.5005
R20789 CSoutput.n266 CSoutput.n164 4.5005
R20790 CSoutput.n266 CSoutput.n168 4.5005
R20791 CSoutput.n266 CSoutput.n163 4.5005
R20792 CSoutput.n266 CSoutput.t184 4.5005
R20793 CSoutput.n266 CSoutput.n162 4.5005
R20794 CSoutput.n266 CSoutput.n169 4.5005
R20795 CSoutput.n266 CSoutput.n170 4.5005
R20796 CSoutput.n253 CSoutput.n224 4.5005
R20797 CSoutput.n253 CSoutput.n230 4.5005
R20798 CSoutput.n211 CSoutput.n200 4.5005
R20799 CSoutput.n211 CSoutput.n202 4.5005
R20800 CSoutput.n211 CSoutput.n199 4.5005
R20801 CSoutput.n211 CSoutput.n203 4.5005
R20802 CSoutput.n211 CSoutput.n198 4.5005
R20803 CSoutput.n211 CSoutput.t186 4.5005
R20804 CSoutput.n211 CSoutput.n197 4.5005
R20805 CSoutput.n211 CSoutput.n204 4.5005
R20806 CSoutput.n253 CSoutput.n211 4.5005
R20807 CSoutput.n232 CSoutput.n200 4.5005
R20808 CSoutput.n232 CSoutput.n202 4.5005
R20809 CSoutput.n232 CSoutput.n199 4.5005
R20810 CSoutput.n232 CSoutput.n203 4.5005
R20811 CSoutput.n232 CSoutput.n198 4.5005
R20812 CSoutput.n232 CSoutput.t186 4.5005
R20813 CSoutput.n232 CSoutput.n197 4.5005
R20814 CSoutput.n232 CSoutput.n204 4.5005
R20815 CSoutput.n253 CSoutput.n232 4.5005
R20816 CSoutput.n210 CSoutput.n200 4.5005
R20817 CSoutput.n210 CSoutput.n202 4.5005
R20818 CSoutput.n210 CSoutput.n199 4.5005
R20819 CSoutput.n210 CSoutput.n203 4.5005
R20820 CSoutput.n210 CSoutput.n198 4.5005
R20821 CSoutput.n210 CSoutput.t186 4.5005
R20822 CSoutput.n210 CSoutput.n197 4.5005
R20823 CSoutput.n210 CSoutput.n204 4.5005
R20824 CSoutput.n253 CSoutput.n210 4.5005
R20825 CSoutput.n234 CSoutput.n200 4.5005
R20826 CSoutput.n234 CSoutput.n202 4.5005
R20827 CSoutput.n234 CSoutput.n199 4.5005
R20828 CSoutput.n234 CSoutput.n203 4.5005
R20829 CSoutput.n234 CSoutput.n198 4.5005
R20830 CSoutput.n234 CSoutput.t186 4.5005
R20831 CSoutput.n234 CSoutput.n197 4.5005
R20832 CSoutput.n234 CSoutput.n204 4.5005
R20833 CSoutput.n253 CSoutput.n234 4.5005
R20834 CSoutput.n200 CSoutput.n195 4.5005
R20835 CSoutput.n202 CSoutput.n195 4.5005
R20836 CSoutput.n199 CSoutput.n195 4.5005
R20837 CSoutput.n203 CSoutput.n195 4.5005
R20838 CSoutput.n198 CSoutput.n195 4.5005
R20839 CSoutput.t186 CSoutput.n195 4.5005
R20840 CSoutput.n197 CSoutput.n195 4.5005
R20841 CSoutput.n204 CSoutput.n195 4.5005
R20842 CSoutput.n256 CSoutput.n200 4.5005
R20843 CSoutput.n256 CSoutput.n202 4.5005
R20844 CSoutput.n256 CSoutput.n199 4.5005
R20845 CSoutput.n256 CSoutput.n203 4.5005
R20846 CSoutput.n256 CSoutput.n198 4.5005
R20847 CSoutput.n256 CSoutput.t186 4.5005
R20848 CSoutput.n256 CSoutput.n197 4.5005
R20849 CSoutput.n256 CSoutput.n204 4.5005
R20850 CSoutput.n254 CSoutput.n200 4.5005
R20851 CSoutput.n254 CSoutput.n202 4.5005
R20852 CSoutput.n254 CSoutput.n199 4.5005
R20853 CSoutput.n254 CSoutput.n203 4.5005
R20854 CSoutput.n254 CSoutput.n198 4.5005
R20855 CSoutput.n254 CSoutput.t186 4.5005
R20856 CSoutput.n254 CSoutput.n197 4.5005
R20857 CSoutput.n254 CSoutput.n204 4.5005
R20858 CSoutput.n254 CSoutput.n253 4.5005
R20859 CSoutput.n236 CSoutput.n200 4.5005
R20860 CSoutput.n236 CSoutput.n202 4.5005
R20861 CSoutput.n236 CSoutput.n199 4.5005
R20862 CSoutput.n236 CSoutput.n203 4.5005
R20863 CSoutput.n236 CSoutput.n198 4.5005
R20864 CSoutput.n236 CSoutput.t186 4.5005
R20865 CSoutput.n236 CSoutput.n197 4.5005
R20866 CSoutput.n236 CSoutput.n204 4.5005
R20867 CSoutput.n253 CSoutput.n236 4.5005
R20868 CSoutput.n208 CSoutput.n200 4.5005
R20869 CSoutput.n208 CSoutput.n202 4.5005
R20870 CSoutput.n208 CSoutput.n199 4.5005
R20871 CSoutput.n208 CSoutput.n203 4.5005
R20872 CSoutput.n208 CSoutput.n198 4.5005
R20873 CSoutput.n208 CSoutput.t186 4.5005
R20874 CSoutput.n208 CSoutput.n197 4.5005
R20875 CSoutput.n208 CSoutput.n204 4.5005
R20876 CSoutput.n253 CSoutput.n208 4.5005
R20877 CSoutput.n238 CSoutput.n200 4.5005
R20878 CSoutput.n238 CSoutput.n202 4.5005
R20879 CSoutput.n238 CSoutput.n199 4.5005
R20880 CSoutput.n238 CSoutput.n203 4.5005
R20881 CSoutput.n238 CSoutput.n198 4.5005
R20882 CSoutput.n238 CSoutput.t186 4.5005
R20883 CSoutput.n238 CSoutput.n197 4.5005
R20884 CSoutput.n238 CSoutput.n204 4.5005
R20885 CSoutput.n253 CSoutput.n238 4.5005
R20886 CSoutput.n207 CSoutput.n200 4.5005
R20887 CSoutput.n207 CSoutput.n202 4.5005
R20888 CSoutput.n207 CSoutput.n199 4.5005
R20889 CSoutput.n207 CSoutput.n203 4.5005
R20890 CSoutput.n207 CSoutput.n198 4.5005
R20891 CSoutput.n207 CSoutput.t186 4.5005
R20892 CSoutput.n207 CSoutput.n197 4.5005
R20893 CSoutput.n207 CSoutput.n204 4.5005
R20894 CSoutput.n253 CSoutput.n207 4.5005
R20895 CSoutput.n252 CSoutput.n200 4.5005
R20896 CSoutput.n252 CSoutput.n202 4.5005
R20897 CSoutput.n252 CSoutput.n199 4.5005
R20898 CSoutput.n252 CSoutput.n203 4.5005
R20899 CSoutput.n252 CSoutput.n198 4.5005
R20900 CSoutput.n252 CSoutput.t186 4.5005
R20901 CSoutput.n252 CSoutput.n197 4.5005
R20902 CSoutput.n252 CSoutput.n204 4.5005
R20903 CSoutput.n253 CSoutput.n252 4.5005
R20904 CSoutput.n251 CSoutput.n136 4.5005
R20905 CSoutput.n152 CSoutput.n136 4.5005
R20906 CSoutput.n147 CSoutput.n131 4.5005
R20907 CSoutput.n147 CSoutput.n133 4.5005
R20908 CSoutput.n147 CSoutput.n130 4.5005
R20909 CSoutput.n147 CSoutput.n134 4.5005
R20910 CSoutput.n147 CSoutput.n129 4.5005
R20911 CSoutput.n147 CSoutput.t187 4.5005
R20912 CSoutput.n147 CSoutput.n128 4.5005
R20913 CSoutput.n147 CSoutput.n135 4.5005
R20914 CSoutput.n147 CSoutput.n136 4.5005
R20915 CSoutput.n145 CSoutput.n131 4.5005
R20916 CSoutput.n145 CSoutput.n133 4.5005
R20917 CSoutput.n145 CSoutput.n130 4.5005
R20918 CSoutput.n145 CSoutput.n134 4.5005
R20919 CSoutput.n145 CSoutput.n129 4.5005
R20920 CSoutput.n145 CSoutput.t187 4.5005
R20921 CSoutput.n145 CSoutput.n128 4.5005
R20922 CSoutput.n145 CSoutput.n135 4.5005
R20923 CSoutput.n145 CSoutput.n136 4.5005
R20924 CSoutput.n144 CSoutput.n131 4.5005
R20925 CSoutput.n144 CSoutput.n133 4.5005
R20926 CSoutput.n144 CSoutput.n130 4.5005
R20927 CSoutput.n144 CSoutput.n134 4.5005
R20928 CSoutput.n144 CSoutput.n129 4.5005
R20929 CSoutput.n144 CSoutput.t187 4.5005
R20930 CSoutput.n144 CSoutput.n128 4.5005
R20931 CSoutput.n144 CSoutput.n135 4.5005
R20932 CSoutput.n144 CSoutput.n136 4.5005
R20933 CSoutput.n273 CSoutput.n131 4.5005
R20934 CSoutput.n273 CSoutput.n133 4.5005
R20935 CSoutput.n273 CSoutput.n130 4.5005
R20936 CSoutput.n273 CSoutput.n134 4.5005
R20937 CSoutput.n273 CSoutput.n129 4.5005
R20938 CSoutput.n273 CSoutput.t187 4.5005
R20939 CSoutput.n273 CSoutput.n128 4.5005
R20940 CSoutput.n273 CSoutput.n135 4.5005
R20941 CSoutput.n273 CSoutput.n136 4.5005
R20942 CSoutput.n271 CSoutput.n131 4.5005
R20943 CSoutput.n271 CSoutput.n133 4.5005
R20944 CSoutput.n271 CSoutput.n130 4.5005
R20945 CSoutput.n271 CSoutput.n134 4.5005
R20946 CSoutput.n271 CSoutput.n129 4.5005
R20947 CSoutput.n271 CSoutput.t187 4.5005
R20948 CSoutput.n271 CSoutput.n128 4.5005
R20949 CSoutput.n271 CSoutput.n135 4.5005
R20950 CSoutput.n269 CSoutput.n131 4.5005
R20951 CSoutput.n269 CSoutput.n133 4.5005
R20952 CSoutput.n269 CSoutput.n130 4.5005
R20953 CSoutput.n269 CSoutput.n134 4.5005
R20954 CSoutput.n269 CSoutput.n129 4.5005
R20955 CSoutput.n269 CSoutput.t187 4.5005
R20956 CSoutput.n269 CSoutput.n128 4.5005
R20957 CSoutput.n269 CSoutput.n135 4.5005
R20958 CSoutput.n155 CSoutput.n131 4.5005
R20959 CSoutput.n155 CSoutput.n133 4.5005
R20960 CSoutput.n155 CSoutput.n130 4.5005
R20961 CSoutput.n155 CSoutput.n134 4.5005
R20962 CSoutput.n155 CSoutput.n129 4.5005
R20963 CSoutput.n155 CSoutput.t187 4.5005
R20964 CSoutput.n155 CSoutput.n128 4.5005
R20965 CSoutput.n155 CSoutput.n135 4.5005
R20966 CSoutput.n155 CSoutput.n136 4.5005
R20967 CSoutput.n154 CSoutput.n131 4.5005
R20968 CSoutput.n154 CSoutput.n133 4.5005
R20969 CSoutput.n154 CSoutput.n130 4.5005
R20970 CSoutput.n154 CSoutput.n134 4.5005
R20971 CSoutput.n154 CSoutput.n129 4.5005
R20972 CSoutput.n154 CSoutput.t187 4.5005
R20973 CSoutput.n154 CSoutput.n128 4.5005
R20974 CSoutput.n154 CSoutput.n135 4.5005
R20975 CSoutput.n154 CSoutput.n136 4.5005
R20976 CSoutput.n158 CSoutput.n131 4.5005
R20977 CSoutput.n158 CSoutput.n133 4.5005
R20978 CSoutput.n158 CSoutput.n130 4.5005
R20979 CSoutput.n158 CSoutput.n134 4.5005
R20980 CSoutput.n158 CSoutput.n129 4.5005
R20981 CSoutput.n158 CSoutput.t187 4.5005
R20982 CSoutput.n158 CSoutput.n128 4.5005
R20983 CSoutput.n158 CSoutput.n135 4.5005
R20984 CSoutput.n158 CSoutput.n136 4.5005
R20985 CSoutput.n157 CSoutput.n131 4.5005
R20986 CSoutput.n157 CSoutput.n133 4.5005
R20987 CSoutput.n157 CSoutput.n130 4.5005
R20988 CSoutput.n157 CSoutput.n134 4.5005
R20989 CSoutput.n157 CSoutput.n129 4.5005
R20990 CSoutput.n157 CSoutput.t187 4.5005
R20991 CSoutput.n157 CSoutput.n128 4.5005
R20992 CSoutput.n157 CSoutput.n135 4.5005
R20993 CSoutput.n157 CSoutput.n136 4.5005
R20994 CSoutput.n140 CSoutput.n131 4.5005
R20995 CSoutput.n140 CSoutput.n133 4.5005
R20996 CSoutput.n140 CSoutput.n130 4.5005
R20997 CSoutput.n140 CSoutput.n134 4.5005
R20998 CSoutput.n140 CSoutput.n129 4.5005
R20999 CSoutput.n140 CSoutput.t187 4.5005
R21000 CSoutput.n140 CSoutput.n128 4.5005
R21001 CSoutput.n140 CSoutput.n135 4.5005
R21002 CSoutput.n140 CSoutput.n136 4.5005
R21003 CSoutput.n276 CSoutput.n131 4.5005
R21004 CSoutput.n276 CSoutput.n133 4.5005
R21005 CSoutput.n276 CSoutput.n130 4.5005
R21006 CSoutput.n276 CSoutput.n134 4.5005
R21007 CSoutput.n276 CSoutput.n129 4.5005
R21008 CSoutput.n276 CSoutput.t187 4.5005
R21009 CSoutput.n276 CSoutput.n128 4.5005
R21010 CSoutput.n276 CSoutput.n135 4.5005
R21011 CSoutput.n276 CSoutput.n136 4.5005
R21012 CSoutput.n323 CSoutput.n307 4.10845
R21013 CSoutput.n125 CSoutput.n109 4.10845
R21014 CSoutput.n321 CSoutput.t66 4.06363
R21015 CSoutput.n321 CSoutput.t119 4.06363
R21016 CSoutput.n319 CSoutput.t136 4.06363
R21017 CSoutput.n319 CSoutput.t137 4.06363
R21018 CSoutput.n317 CSoutput.t79 4.06363
R21019 CSoutput.n317 CSoutput.t80 4.06363
R21020 CSoutput.n315 CSoutput.t85 4.06363
R21021 CSoutput.n315 CSoutput.t138 4.06363
R21022 CSoutput.n313 CSoutput.t58 4.06363
R21023 CSoutput.n313 CSoutput.t83 4.06363
R21024 CSoutput.n311 CSoutput.t97 4.06363
R21025 CSoutput.n311 CSoutput.t115 4.06363
R21026 CSoutput.n309 CSoutput.t121 4.06363
R21027 CSoutput.n309 CSoutput.t62 4.06363
R21028 CSoutput.n308 CSoutput.t98 4.06363
R21029 CSoutput.n308 CSoutput.t99 4.06363
R21030 CSoutput.n305 CSoutput.t55 4.06363
R21031 CSoutput.n305 CSoutput.t107 4.06363
R21032 CSoutput.n303 CSoutput.t125 4.06363
R21033 CSoutput.n303 CSoutput.t126 4.06363
R21034 CSoutput.n301 CSoutput.t70 4.06363
R21035 CSoutput.n301 CSoutput.t71 4.06363
R21036 CSoutput.n299 CSoutput.t74 4.06363
R21037 CSoutput.n299 CSoutput.t129 4.06363
R21038 CSoutput.n297 CSoutput.t46 4.06363
R21039 CSoutput.n297 CSoutput.t73 4.06363
R21040 CSoutput.n295 CSoutput.t86 4.06363
R21041 CSoutput.n295 CSoutput.t106 4.06363
R21042 CSoutput.n293 CSoutput.t108 4.06363
R21043 CSoutput.n293 CSoutput.t50 4.06363
R21044 CSoutput.n292 CSoutput.t91 4.06363
R21045 CSoutput.n292 CSoutput.t92 4.06363
R21046 CSoutput.n290 CSoutput.t123 4.06363
R21047 CSoutput.n290 CSoutput.t59 4.06363
R21048 CSoutput.n288 CSoutput.t89 4.06363
R21049 CSoutput.n288 CSoutput.t72 4.06363
R21050 CSoutput.n286 CSoutput.t75 4.06363
R21051 CSoutput.n286 CSoutput.t56 4.06363
R21052 CSoutput.n284 CSoutput.t113 4.06363
R21053 CSoutput.n284 CSoutput.t51 4.06363
R21054 CSoutput.n282 CSoutput.t81 4.06363
R21055 CSoutput.n282 CSoutput.t134 4.06363
R21056 CSoutput.n280 CSoutput.t67 4.06363
R21057 CSoutput.n280 CSoutput.t117 4.06363
R21058 CSoutput.n278 CSoutput.t87 4.06363
R21059 CSoutput.n278 CSoutput.t139 4.06363
R21060 CSoutput.n277 CSoutput.t47 4.06363
R21061 CSoutput.n277 CSoutput.t127 4.06363
R21062 CSoutput.n110 CSoutput.t133 4.06363
R21063 CSoutput.n110 CSoutput.t132 4.06363
R21064 CSoutput.n111 CSoutput.t114 4.06363
R21065 CSoutput.n111 CSoutput.t64 4.06363
R21066 CSoutput.n113 CSoutput.t61 4.06363
R21067 CSoutput.n113 CSoutput.t130 4.06363
R21068 CSoutput.n115 CSoutput.t112 4.06363
R21069 CSoutput.n115 CSoutput.t95 4.06363
R21070 CSoutput.n117 CSoutput.t78 4.06363
R21071 CSoutput.n117 CSoutput.t141 4.06363
R21072 CSoutput.n119 CSoutput.t110 4.06363
R21073 CSoutput.n119 CSoutput.t109 4.06363
R21074 CSoutput.n121 CSoutput.t100 4.06363
R21075 CSoutput.n121 CSoutput.t77 4.06363
R21076 CSoutput.n123 CSoutput.t63 4.06363
R21077 CSoutput.n123 CSoutput.t101 4.06363
R21078 CSoutput.n94 CSoutput.t122 4.06363
R21079 CSoutput.n94 CSoutput.t120 4.06363
R21080 CSoutput.n95 CSoutput.t105 4.06363
R21081 CSoutput.n95 CSoutput.t54 4.06363
R21082 CSoutput.n97 CSoutput.t49 4.06363
R21083 CSoutput.n97 CSoutput.t116 4.06363
R21084 CSoutput.n99 CSoutput.t104 4.06363
R21085 CSoutput.n99 CSoutput.t84 4.06363
R21086 CSoutput.n101 CSoutput.t69 4.06363
R21087 CSoutput.n101 CSoutput.t131 4.06363
R21088 CSoutput.n103 CSoutput.t103 4.06363
R21089 CSoutput.n103 CSoutput.t102 4.06363
R21090 CSoutput.n105 CSoutput.t93 4.06363
R21091 CSoutput.n105 CSoutput.t65 4.06363
R21092 CSoutput.n107 CSoutput.t52 4.06363
R21093 CSoutput.n107 CSoutput.t94 4.06363
R21094 CSoutput.n79 CSoutput.t128 4.06363
R21095 CSoutput.n79 CSoutput.t48 4.06363
R21096 CSoutput.n80 CSoutput.t111 4.06363
R21097 CSoutput.n80 CSoutput.t88 4.06363
R21098 CSoutput.n82 CSoutput.t118 4.06363
R21099 CSoutput.n82 CSoutput.t68 4.06363
R21100 CSoutput.n84 CSoutput.t135 4.06363
R21101 CSoutput.n84 CSoutput.t82 4.06363
R21102 CSoutput.n86 CSoutput.t53 4.06363
R21103 CSoutput.n86 CSoutput.t96 4.06363
R21104 CSoutput.n88 CSoutput.t57 4.06363
R21105 CSoutput.n88 CSoutput.t76 4.06363
R21106 CSoutput.n90 CSoutput.t140 4.06363
R21107 CSoutput.n90 CSoutput.t90 4.06363
R21108 CSoutput.n92 CSoutput.t60 4.06363
R21109 CSoutput.n92 CSoutput.t124 4.06363
R21110 CSoutput.n44 CSoutput.n43 3.79402
R21111 CSoutput.n49 CSoutput.n48 3.79402
R21112 CSoutput.n404 CSoutput.n364 3.71319
R21113 CSoutput.n405 CSoutput.n404 3.57343
R21114 CSoutput.n361 CSoutput.t26 2.82907
R21115 CSoutput.n361 CSoutput.t174 2.82907
R21116 CSoutput.n359 CSoutput.t10 2.82907
R21117 CSoutput.n359 CSoutput.t165 2.82907
R21118 CSoutput.n357 CSoutput.t12 2.82907
R21119 CSoutput.n357 CSoutput.t170 2.82907
R21120 CSoutput.n355 CSoutput.t8 2.82907
R21121 CSoutput.n355 CSoutput.t38 2.82907
R21122 CSoutput.n353 CSoutput.t3 2.82907
R21123 CSoutput.n353 CSoutput.t5 2.82907
R21124 CSoutput.n351 CSoutput.t39 2.82907
R21125 CSoutput.n351 CSoutput.t16 2.82907
R21126 CSoutput.n349 CSoutput.t25 2.82907
R21127 CSoutput.n349 CSoutput.t152 2.82907
R21128 CSoutput.n347 CSoutput.t147 2.82907
R21129 CSoutput.n347 CSoutput.t162 2.82907
R21130 CSoutput.n345 CSoutput.t20 2.82907
R21131 CSoutput.n345 CSoutput.t169 2.82907
R21132 CSoutput.n344 CSoutput.t173 2.82907
R21133 CSoutput.n344 CSoutput.t146 2.82907
R21134 CSoutput.n342 CSoutput.t24 2.82907
R21135 CSoutput.n342 CSoutput.t31 2.82907
R21136 CSoutput.n340 CSoutput.t166 2.82907
R21137 CSoutput.n340 CSoutput.t175 2.82907
R21138 CSoutput.n338 CSoutput.t160 2.82907
R21139 CSoutput.n338 CSoutput.t148 2.82907
R21140 CSoutput.n336 CSoutput.t145 2.82907
R21141 CSoutput.n336 CSoutput.t44 2.82907
R21142 CSoutput.n334 CSoutput.t149 2.82907
R21143 CSoutput.n334 CSoutput.t168 2.82907
R21144 CSoutput.n332 CSoutput.t21 2.82907
R21145 CSoutput.n332 CSoutput.t4 2.82907
R21146 CSoutput.n330 CSoutput.t23 2.82907
R21147 CSoutput.n330 CSoutput.t11 2.82907
R21148 CSoutput.n328 CSoutput.t167 2.82907
R21149 CSoutput.n328 CSoutput.t153 2.82907
R21150 CSoutput.n326 CSoutput.t33 2.82907
R21151 CSoutput.n326 CSoutput.t32 2.82907
R21152 CSoutput.n325 CSoutput.t7 2.82907
R21153 CSoutput.n325 CSoutput.t17 2.82907
R21154 CSoutput.n384 CSoutput.t155 2.82907
R21155 CSoutput.n384 CSoutput.t37 2.82907
R21156 CSoutput.n385 CSoutput.t0 2.82907
R21157 CSoutput.n385 CSoutput.t6 2.82907
R21158 CSoutput.n387 CSoutput.t34 2.82907
R21159 CSoutput.n387 CSoutput.t163 2.82907
R21160 CSoutput.n389 CSoutput.t2 2.82907
R21161 CSoutput.n389 CSoutput.t28 2.82907
R21162 CSoutput.n391 CSoutput.t19 2.82907
R21163 CSoutput.n391 CSoutput.t41 2.82907
R21164 CSoutput.n393 CSoutput.t43 2.82907
R21165 CSoutput.n393 CSoutput.t30 2.82907
R21166 CSoutput.n395 CSoutput.t171 2.82907
R21167 CSoutput.n395 CSoutput.t35 2.82907
R21168 CSoutput.n397 CSoutput.t1 2.82907
R21169 CSoutput.n397 CSoutput.t157 2.82907
R21170 CSoutput.n399 CSoutput.t18 2.82907
R21171 CSoutput.n399 CSoutput.t143 2.82907
R21172 CSoutput.n401 CSoutput.t161 2.82907
R21173 CSoutput.n401 CSoutput.t156 2.82907
R21174 CSoutput.n365 CSoutput.t29 2.82907
R21175 CSoutput.n365 CSoutput.t45 2.82907
R21176 CSoutput.n366 CSoutput.t164 2.82907
R21177 CSoutput.n366 CSoutput.t158 2.82907
R21178 CSoutput.n368 CSoutput.t27 2.82907
R21179 CSoutput.n368 CSoutput.t42 2.82907
R21180 CSoutput.n370 CSoutput.t40 2.82907
R21181 CSoutput.n370 CSoutput.t150 2.82907
R21182 CSoutput.n372 CSoutput.t159 2.82907
R21183 CSoutput.n372 CSoutput.t14 2.82907
R21184 CSoutput.n374 CSoutput.t142 2.82907
R21185 CSoutput.n374 CSoutput.t151 2.82907
R21186 CSoutput.n376 CSoutput.t13 2.82907
R21187 CSoutput.n376 CSoutput.t154 2.82907
R21188 CSoutput.n378 CSoutput.t172 2.82907
R21189 CSoutput.n378 CSoutput.t144 2.82907
R21190 CSoutput.n380 CSoutput.t15 2.82907
R21191 CSoutput.n380 CSoutput.t22 2.82907
R21192 CSoutput.n382 CSoutput.t36 2.82907
R21193 CSoutput.n382 CSoutput.t9 2.82907
R21194 CSoutput.n75 CSoutput.n1 2.45513
R21195 CSoutput.n324 CSoutput.n126 2.36742
R21196 CSoutput.n217 CSoutput.n215 2.251
R21197 CSoutput.n217 CSoutput.n214 2.251
R21198 CSoutput.n217 CSoutput.n213 2.251
R21199 CSoutput.n217 CSoutput.n212 2.251
R21200 CSoutput.n186 CSoutput.n185 2.251
R21201 CSoutput.n186 CSoutput.n184 2.251
R21202 CSoutput.n186 CSoutput.n183 2.251
R21203 CSoutput.n186 CSoutput.n182 2.251
R21204 CSoutput.n259 CSoutput.n258 2.251
R21205 CSoutput.n224 CSoutput.n222 2.251
R21206 CSoutput.n224 CSoutput.n221 2.251
R21207 CSoutput.n224 CSoutput.n220 2.251
R21208 CSoutput.n242 CSoutput.n224 2.251
R21209 CSoutput.n230 CSoutput.n229 2.251
R21210 CSoutput.n230 CSoutput.n228 2.251
R21211 CSoutput.n230 CSoutput.n227 2.251
R21212 CSoutput.n230 CSoutput.n226 2.251
R21213 CSoutput.n256 CSoutput.n196 2.251
R21214 CSoutput.n251 CSoutput.n249 2.251
R21215 CSoutput.n251 CSoutput.n248 2.251
R21216 CSoutput.n251 CSoutput.n247 2.251
R21217 CSoutput.n251 CSoutput.n246 2.251
R21218 CSoutput.n152 CSoutput.n151 2.251
R21219 CSoutput.n152 CSoutput.n150 2.251
R21220 CSoutput.n152 CSoutput.n149 2.251
R21221 CSoutput.n152 CSoutput.n148 2.251
R21222 CSoutput.n269 CSoutput.n268 2.251
R21223 CSoutput.n186 CSoutput.n166 2.2505
R21224 CSoutput.n181 CSoutput.n166 2.2505
R21225 CSoutput.n179 CSoutput.n166 2.2505
R21226 CSoutput.n178 CSoutput.n166 2.2505
R21227 CSoutput.n263 CSoutput.n166 2.2505
R21228 CSoutput.n261 CSoutput.n166 2.2505
R21229 CSoutput.n259 CSoutput.n166 2.2505
R21230 CSoutput.n189 CSoutput.n166 2.2505
R21231 CSoutput.n188 CSoutput.n166 2.2505
R21232 CSoutput.n192 CSoutput.n166 2.2505
R21233 CSoutput.n191 CSoutput.n166 2.2505
R21234 CSoutput.n174 CSoutput.n166 2.2505
R21235 CSoutput.n266 CSoutput.n166 2.2505
R21236 CSoutput.n266 CSoutput.n265 2.2505
R21237 CSoutput.n230 CSoutput.n201 2.2505
R21238 CSoutput.n211 CSoutput.n201 2.2505
R21239 CSoutput.n232 CSoutput.n201 2.2505
R21240 CSoutput.n210 CSoutput.n201 2.2505
R21241 CSoutput.n234 CSoutput.n201 2.2505
R21242 CSoutput.n201 CSoutput.n195 2.2505
R21243 CSoutput.n256 CSoutput.n201 2.2505
R21244 CSoutput.n254 CSoutput.n201 2.2505
R21245 CSoutput.n236 CSoutput.n201 2.2505
R21246 CSoutput.n208 CSoutput.n201 2.2505
R21247 CSoutput.n238 CSoutput.n201 2.2505
R21248 CSoutput.n207 CSoutput.n201 2.2505
R21249 CSoutput.n252 CSoutput.n201 2.2505
R21250 CSoutput.n252 CSoutput.n205 2.2505
R21251 CSoutput.n152 CSoutput.n132 2.2505
R21252 CSoutput.n147 CSoutput.n132 2.2505
R21253 CSoutput.n145 CSoutput.n132 2.2505
R21254 CSoutput.n144 CSoutput.n132 2.2505
R21255 CSoutput.n273 CSoutput.n132 2.2505
R21256 CSoutput.n271 CSoutput.n132 2.2505
R21257 CSoutput.n269 CSoutput.n132 2.2505
R21258 CSoutput.n155 CSoutput.n132 2.2505
R21259 CSoutput.n154 CSoutput.n132 2.2505
R21260 CSoutput.n158 CSoutput.n132 2.2505
R21261 CSoutput.n157 CSoutput.n132 2.2505
R21262 CSoutput.n140 CSoutput.n132 2.2505
R21263 CSoutput.n276 CSoutput.n132 2.2505
R21264 CSoutput.n276 CSoutput.n275 2.2505
R21265 CSoutput.n194 CSoutput.n187 2.25024
R21266 CSoutput.n194 CSoutput.n180 2.25024
R21267 CSoutput.n262 CSoutput.n194 2.25024
R21268 CSoutput.n194 CSoutput.n190 2.25024
R21269 CSoutput.n194 CSoutput.n193 2.25024
R21270 CSoutput.n194 CSoutput.n161 2.25024
R21271 CSoutput.n244 CSoutput.n241 2.25024
R21272 CSoutput.n244 CSoutput.n240 2.25024
R21273 CSoutput.n244 CSoutput.n239 2.25024
R21274 CSoutput.n244 CSoutput.n206 2.25024
R21275 CSoutput.n244 CSoutput.n243 2.25024
R21276 CSoutput.n245 CSoutput.n244 2.25024
R21277 CSoutput.n160 CSoutput.n153 2.25024
R21278 CSoutput.n160 CSoutput.n146 2.25024
R21279 CSoutput.n272 CSoutput.n160 2.25024
R21280 CSoutput.n160 CSoutput.n156 2.25024
R21281 CSoutput.n160 CSoutput.n159 2.25024
R21282 CSoutput.n160 CSoutput.n127 2.25024
R21283 CSoutput.n261 CSoutput.n171 1.50111
R21284 CSoutput.n209 CSoutput.n195 1.50111
R21285 CSoutput.n271 CSoutput.n137 1.50111
R21286 CSoutput.n217 CSoutput.n216 1.501
R21287 CSoutput.n224 CSoutput.n223 1.501
R21288 CSoutput.n251 CSoutput.n250 1.501
R21289 CSoutput.n265 CSoutput.n176 1.12536
R21290 CSoutput.n265 CSoutput.n177 1.12536
R21291 CSoutput.n265 CSoutput.n264 1.12536
R21292 CSoutput.n225 CSoutput.n205 1.12536
R21293 CSoutput.n231 CSoutput.n205 1.12536
R21294 CSoutput.n233 CSoutput.n205 1.12536
R21295 CSoutput.n275 CSoutput.n142 1.12536
R21296 CSoutput.n275 CSoutput.n143 1.12536
R21297 CSoutput.n275 CSoutput.n274 1.12536
R21298 CSoutput.n265 CSoutput.n172 1.12536
R21299 CSoutput.n265 CSoutput.n173 1.12536
R21300 CSoutput.n265 CSoutput.n175 1.12536
R21301 CSoutput.n255 CSoutput.n205 1.12536
R21302 CSoutput.n235 CSoutput.n205 1.12536
R21303 CSoutput.n237 CSoutput.n205 1.12536
R21304 CSoutput.n275 CSoutput.n138 1.12536
R21305 CSoutput.n275 CSoutput.n139 1.12536
R21306 CSoutput.n275 CSoutput.n141 1.12536
R21307 CSoutput.n31 CSoutput.n30 0.669944
R21308 CSoutput.n62 CSoutput.n61 0.669944
R21309 CSoutput.n348 CSoutput.n346 0.573776
R21310 CSoutput.n350 CSoutput.n348 0.573776
R21311 CSoutput.n352 CSoutput.n350 0.573776
R21312 CSoutput.n354 CSoutput.n352 0.573776
R21313 CSoutput.n356 CSoutput.n354 0.573776
R21314 CSoutput.n358 CSoutput.n356 0.573776
R21315 CSoutput.n360 CSoutput.n358 0.573776
R21316 CSoutput.n362 CSoutput.n360 0.573776
R21317 CSoutput.n329 CSoutput.n327 0.573776
R21318 CSoutput.n331 CSoutput.n329 0.573776
R21319 CSoutput.n333 CSoutput.n331 0.573776
R21320 CSoutput.n335 CSoutput.n333 0.573776
R21321 CSoutput.n337 CSoutput.n335 0.573776
R21322 CSoutput.n339 CSoutput.n337 0.573776
R21323 CSoutput.n341 CSoutput.n339 0.573776
R21324 CSoutput.n343 CSoutput.n341 0.573776
R21325 CSoutput.n402 CSoutput.n400 0.573776
R21326 CSoutput.n400 CSoutput.n398 0.573776
R21327 CSoutput.n398 CSoutput.n396 0.573776
R21328 CSoutput.n396 CSoutput.n394 0.573776
R21329 CSoutput.n394 CSoutput.n392 0.573776
R21330 CSoutput.n392 CSoutput.n390 0.573776
R21331 CSoutput.n390 CSoutput.n388 0.573776
R21332 CSoutput.n388 CSoutput.n386 0.573776
R21333 CSoutput.n383 CSoutput.n381 0.573776
R21334 CSoutput.n381 CSoutput.n379 0.573776
R21335 CSoutput.n379 CSoutput.n377 0.573776
R21336 CSoutput.n377 CSoutput.n375 0.573776
R21337 CSoutput.n375 CSoutput.n373 0.573776
R21338 CSoutput.n373 CSoutput.n371 0.573776
R21339 CSoutput.n371 CSoutput.n369 0.573776
R21340 CSoutput.n369 CSoutput.n367 0.573776
R21341 CSoutput.n405 CSoutput.n276 0.53442
R21342 CSoutput.n312 CSoutput.n310 0.358259
R21343 CSoutput.n314 CSoutput.n312 0.358259
R21344 CSoutput.n316 CSoutput.n314 0.358259
R21345 CSoutput.n318 CSoutput.n316 0.358259
R21346 CSoutput.n320 CSoutput.n318 0.358259
R21347 CSoutput.n322 CSoutput.n320 0.358259
R21348 CSoutput.n296 CSoutput.n294 0.358259
R21349 CSoutput.n298 CSoutput.n296 0.358259
R21350 CSoutput.n300 CSoutput.n298 0.358259
R21351 CSoutput.n302 CSoutput.n300 0.358259
R21352 CSoutput.n304 CSoutput.n302 0.358259
R21353 CSoutput.n306 CSoutput.n304 0.358259
R21354 CSoutput.n281 CSoutput.n279 0.358259
R21355 CSoutput.n283 CSoutput.n281 0.358259
R21356 CSoutput.n285 CSoutput.n283 0.358259
R21357 CSoutput.n287 CSoutput.n285 0.358259
R21358 CSoutput.n289 CSoutput.n287 0.358259
R21359 CSoutput.n291 CSoutput.n289 0.358259
R21360 CSoutput.n124 CSoutput.n122 0.358259
R21361 CSoutput.n122 CSoutput.n120 0.358259
R21362 CSoutput.n120 CSoutput.n118 0.358259
R21363 CSoutput.n118 CSoutput.n116 0.358259
R21364 CSoutput.n116 CSoutput.n114 0.358259
R21365 CSoutput.n114 CSoutput.n112 0.358259
R21366 CSoutput.n108 CSoutput.n106 0.358259
R21367 CSoutput.n106 CSoutput.n104 0.358259
R21368 CSoutput.n104 CSoutput.n102 0.358259
R21369 CSoutput.n102 CSoutput.n100 0.358259
R21370 CSoutput.n100 CSoutput.n98 0.358259
R21371 CSoutput.n98 CSoutput.n96 0.358259
R21372 CSoutput.n93 CSoutput.n91 0.358259
R21373 CSoutput.n91 CSoutput.n89 0.358259
R21374 CSoutput.n89 CSoutput.n87 0.358259
R21375 CSoutput.n87 CSoutput.n85 0.358259
R21376 CSoutput.n85 CSoutput.n83 0.358259
R21377 CSoutput.n83 CSoutput.n81 0.358259
R21378 CSoutput.n21 CSoutput.n20 0.169105
R21379 CSoutput.n21 CSoutput.n16 0.169105
R21380 CSoutput.n26 CSoutput.n16 0.169105
R21381 CSoutput.n27 CSoutput.n26 0.169105
R21382 CSoutput.n27 CSoutput.n14 0.169105
R21383 CSoutput.n32 CSoutput.n14 0.169105
R21384 CSoutput.n33 CSoutput.n32 0.169105
R21385 CSoutput.n34 CSoutput.n33 0.169105
R21386 CSoutput.n34 CSoutput.n12 0.169105
R21387 CSoutput.n39 CSoutput.n12 0.169105
R21388 CSoutput.n40 CSoutput.n39 0.169105
R21389 CSoutput.n40 CSoutput.n10 0.169105
R21390 CSoutput.n45 CSoutput.n10 0.169105
R21391 CSoutput.n46 CSoutput.n45 0.169105
R21392 CSoutput.n47 CSoutput.n46 0.169105
R21393 CSoutput.n47 CSoutput.n8 0.169105
R21394 CSoutput.n52 CSoutput.n8 0.169105
R21395 CSoutput.n53 CSoutput.n52 0.169105
R21396 CSoutput.n53 CSoutput.n6 0.169105
R21397 CSoutput.n58 CSoutput.n6 0.169105
R21398 CSoutput.n59 CSoutput.n58 0.169105
R21399 CSoutput.n60 CSoutput.n59 0.169105
R21400 CSoutput.n60 CSoutput.n4 0.169105
R21401 CSoutput.n66 CSoutput.n4 0.169105
R21402 CSoutput.n67 CSoutput.n66 0.169105
R21403 CSoutput.n68 CSoutput.n67 0.169105
R21404 CSoutput.n68 CSoutput.n2 0.169105
R21405 CSoutput.n73 CSoutput.n2 0.169105
R21406 CSoutput.n74 CSoutput.n73 0.169105
R21407 CSoutput.n74 CSoutput.n0 0.169105
R21408 CSoutput.n78 CSoutput.n0 0.169105
R21409 CSoutput.n219 CSoutput.n218 0.0910737
R21410 CSoutput.n270 CSoutput.n267 0.0723685
R21411 CSoutput.n224 CSoutput.n219 0.0522944
R21412 CSoutput.n267 CSoutput.n266 0.0499135
R21413 CSoutput.n218 CSoutput.n217 0.0499135
R21414 CSoutput.n252 CSoutput.n251 0.0464294
R21415 CSoutput.n260 CSoutput.n257 0.0391444
R21416 CSoutput.n219 CSoutput.t192 0.023435
R21417 CSoutput.n267 CSoutput.t181 0.02262
R21418 CSoutput.n218 CSoutput.t190 0.02262
R21419 CSoutput CSoutput.n405 0.0052
R21420 CSoutput.n189 CSoutput.n172 0.00365111
R21421 CSoutput.n192 CSoutput.n173 0.00365111
R21422 CSoutput.n175 CSoutput.n174 0.00365111
R21423 CSoutput.n217 CSoutput.n176 0.00365111
R21424 CSoutput.n181 CSoutput.n177 0.00365111
R21425 CSoutput.n264 CSoutput.n178 0.00365111
R21426 CSoutput.n255 CSoutput.n254 0.00365111
R21427 CSoutput.n235 CSoutput.n208 0.00365111
R21428 CSoutput.n237 CSoutput.n207 0.00365111
R21429 CSoutput.n225 CSoutput.n224 0.00365111
R21430 CSoutput.n231 CSoutput.n211 0.00365111
R21431 CSoutput.n233 CSoutput.n210 0.00365111
R21432 CSoutput.n155 CSoutput.n138 0.00365111
R21433 CSoutput.n158 CSoutput.n139 0.00365111
R21434 CSoutput.n141 CSoutput.n140 0.00365111
R21435 CSoutput.n251 CSoutput.n142 0.00365111
R21436 CSoutput.n147 CSoutput.n143 0.00365111
R21437 CSoutput.n274 CSoutput.n144 0.00365111
R21438 CSoutput.n186 CSoutput.n176 0.00340054
R21439 CSoutput.n179 CSoutput.n177 0.00340054
R21440 CSoutput.n264 CSoutput.n263 0.00340054
R21441 CSoutput.n259 CSoutput.n172 0.00340054
R21442 CSoutput.n188 CSoutput.n173 0.00340054
R21443 CSoutput.n191 CSoutput.n175 0.00340054
R21444 CSoutput.n230 CSoutput.n225 0.00340054
R21445 CSoutput.n232 CSoutput.n231 0.00340054
R21446 CSoutput.n234 CSoutput.n233 0.00340054
R21447 CSoutput.n256 CSoutput.n255 0.00340054
R21448 CSoutput.n236 CSoutput.n235 0.00340054
R21449 CSoutput.n238 CSoutput.n237 0.00340054
R21450 CSoutput.n152 CSoutput.n142 0.00340054
R21451 CSoutput.n145 CSoutput.n143 0.00340054
R21452 CSoutput.n274 CSoutput.n273 0.00340054
R21453 CSoutput.n269 CSoutput.n138 0.00340054
R21454 CSoutput.n154 CSoutput.n139 0.00340054
R21455 CSoutput.n157 CSoutput.n141 0.00340054
R21456 CSoutput.n187 CSoutput.n181 0.00252698
R21457 CSoutput.n180 CSoutput.n178 0.00252698
R21458 CSoutput.n262 CSoutput.n261 0.00252698
R21459 CSoutput.n190 CSoutput.n188 0.00252698
R21460 CSoutput.n193 CSoutput.n191 0.00252698
R21461 CSoutput.n266 CSoutput.n161 0.00252698
R21462 CSoutput.n187 CSoutput.n186 0.00252698
R21463 CSoutput.n180 CSoutput.n179 0.00252698
R21464 CSoutput.n263 CSoutput.n262 0.00252698
R21465 CSoutput.n190 CSoutput.n189 0.00252698
R21466 CSoutput.n193 CSoutput.n192 0.00252698
R21467 CSoutput.n174 CSoutput.n161 0.00252698
R21468 CSoutput.n241 CSoutput.n211 0.00252698
R21469 CSoutput.n240 CSoutput.n210 0.00252698
R21470 CSoutput.n239 CSoutput.n195 0.00252698
R21471 CSoutput.n236 CSoutput.n206 0.00252698
R21472 CSoutput.n243 CSoutput.n238 0.00252698
R21473 CSoutput.n252 CSoutput.n245 0.00252698
R21474 CSoutput.n241 CSoutput.n230 0.00252698
R21475 CSoutput.n240 CSoutput.n232 0.00252698
R21476 CSoutput.n239 CSoutput.n234 0.00252698
R21477 CSoutput.n254 CSoutput.n206 0.00252698
R21478 CSoutput.n243 CSoutput.n208 0.00252698
R21479 CSoutput.n245 CSoutput.n207 0.00252698
R21480 CSoutput.n153 CSoutput.n147 0.00252698
R21481 CSoutput.n146 CSoutput.n144 0.00252698
R21482 CSoutput.n272 CSoutput.n271 0.00252698
R21483 CSoutput.n156 CSoutput.n154 0.00252698
R21484 CSoutput.n159 CSoutput.n157 0.00252698
R21485 CSoutput.n276 CSoutput.n127 0.00252698
R21486 CSoutput.n153 CSoutput.n152 0.00252698
R21487 CSoutput.n146 CSoutput.n145 0.00252698
R21488 CSoutput.n273 CSoutput.n272 0.00252698
R21489 CSoutput.n156 CSoutput.n155 0.00252698
R21490 CSoutput.n159 CSoutput.n158 0.00252698
R21491 CSoutput.n140 CSoutput.n127 0.00252698
R21492 CSoutput.n261 CSoutput.n260 0.0020275
R21493 CSoutput.n260 CSoutput.n259 0.0020275
R21494 CSoutput.n257 CSoutput.n195 0.0020275
R21495 CSoutput.n257 CSoutput.n256 0.0020275
R21496 CSoutput.n271 CSoutput.n270 0.0020275
R21497 CSoutput.n270 CSoutput.n269 0.0020275
R21498 CSoutput.n171 CSoutput.n170 0.00166668
R21499 CSoutput.n253 CSoutput.n209 0.00166668
R21500 CSoutput.n137 CSoutput.n136 0.00166668
R21501 CSoutput.n275 CSoutput.n137 0.00133328
R21502 CSoutput.n209 CSoutput.n205 0.00133328
R21503 CSoutput.n265 CSoutput.n171 0.00133328
R21504 CSoutput.n268 CSoutput.n160 0.001
R21505 CSoutput.n246 CSoutput.n160 0.001
R21506 CSoutput.n148 CSoutput.n128 0.001
R21507 CSoutput.n247 CSoutput.n128 0.001
R21508 CSoutput.n149 CSoutput.n129 0.001
R21509 CSoutput.n248 CSoutput.n129 0.001
R21510 CSoutput.n150 CSoutput.n130 0.001
R21511 CSoutput.n249 CSoutput.n130 0.001
R21512 CSoutput.n151 CSoutput.n131 0.001
R21513 CSoutput.n250 CSoutput.n131 0.001
R21514 CSoutput.n244 CSoutput.n196 0.001
R21515 CSoutput.n244 CSoutput.n242 0.001
R21516 CSoutput.n226 CSoutput.n197 0.001
R21517 CSoutput.n220 CSoutput.n197 0.001
R21518 CSoutput.n227 CSoutput.n198 0.001
R21519 CSoutput.n221 CSoutput.n198 0.001
R21520 CSoutput.n228 CSoutput.n199 0.001
R21521 CSoutput.n222 CSoutput.n199 0.001
R21522 CSoutput.n229 CSoutput.n200 0.001
R21523 CSoutput.n223 CSoutput.n200 0.001
R21524 CSoutput.n258 CSoutput.n194 0.001
R21525 CSoutput.n212 CSoutput.n194 0.001
R21526 CSoutput.n182 CSoutput.n162 0.001
R21527 CSoutput.n213 CSoutput.n162 0.001
R21528 CSoutput.n183 CSoutput.n163 0.001
R21529 CSoutput.n214 CSoutput.n163 0.001
R21530 CSoutput.n184 CSoutput.n164 0.001
R21531 CSoutput.n215 CSoutput.n164 0.001
R21532 CSoutput.n185 CSoutput.n165 0.001
R21533 CSoutput.n216 CSoutput.n165 0.001
R21534 CSoutput.n216 CSoutput.n166 0.001
R21535 CSoutput.n215 CSoutput.n167 0.001
R21536 CSoutput.n214 CSoutput.n168 0.001
R21537 CSoutput.n213 CSoutput.t184 0.001
R21538 CSoutput.n212 CSoutput.n169 0.001
R21539 CSoutput.n185 CSoutput.n167 0.001
R21540 CSoutput.n184 CSoutput.n168 0.001
R21541 CSoutput.n183 CSoutput.t184 0.001
R21542 CSoutput.n182 CSoutput.n169 0.001
R21543 CSoutput.n258 CSoutput.n170 0.001
R21544 CSoutput.n223 CSoutput.n201 0.001
R21545 CSoutput.n222 CSoutput.n202 0.001
R21546 CSoutput.n221 CSoutput.n203 0.001
R21547 CSoutput.n220 CSoutput.t186 0.001
R21548 CSoutput.n242 CSoutput.n204 0.001
R21549 CSoutput.n229 CSoutput.n202 0.001
R21550 CSoutput.n228 CSoutput.n203 0.001
R21551 CSoutput.n227 CSoutput.t186 0.001
R21552 CSoutput.n226 CSoutput.n204 0.001
R21553 CSoutput.n253 CSoutput.n196 0.001
R21554 CSoutput.n250 CSoutput.n132 0.001
R21555 CSoutput.n249 CSoutput.n133 0.001
R21556 CSoutput.n248 CSoutput.n134 0.001
R21557 CSoutput.n247 CSoutput.t187 0.001
R21558 CSoutput.n246 CSoutput.n135 0.001
R21559 CSoutput.n151 CSoutput.n133 0.001
R21560 CSoutput.n150 CSoutput.n134 0.001
R21561 CSoutput.n149 CSoutput.t187 0.001
R21562 CSoutput.n148 CSoutput.n135 0.001
R21563 CSoutput.n268 CSoutput.n136 0.001
R21564 a_n1996_n452.n86 a_n1996_n452.t59 512.366
R21565 a_n1996_n452.n76 a_n1996_n452.t50 512.366
R21566 a_n1996_n452.n87 a_n1996_n452.t44 512.366
R21567 a_n1996_n452.n84 a_n1996_n452.t67 512.366
R21568 a_n1996_n452.n77 a_n1996_n452.t56 512.366
R21569 a_n1996_n452.n85 a_n1996_n452.t55 512.366
R21570 a_n1996_n452.n82 a_n1996_n452.t63 512.366
R21571 a_n1996_n452.n78 a_n1996_n452.t48 512.366
R21572 a_n1996_n452.n83 a_n1996_n452.t49 512.366
R21573 a_n1996_n452.n80 a_n1996_n452.t51 512.366
R21574 a_n1996_n452.n79 a_n1996_n452.t60 512.366
R21575 a_n1996_n452.n81 a_n1996_n452.t71 512.366
R21576 a_n1996_n452.n24 a_n1996_n452.t70 539.01
R21577 a_n1996_n452.n91 a_n1996_n452.t53 512.366
R21578 a_n1996_n452.n90 a_n1996_n452.t57 512.366
R21579 a_n1996_n452.n64 a_n1996_n452.t47 512.366
R21580 a_n1996_n452.n89 a_n1996_n452.t62 512.366
R21581 a_n1996_n452.n52 a_n1996_n452.t31 533.058
R21582 a_n1996_n452.n26 a_n1996_n452.t21 539.01
R21583 a_n1996_n452.n94 a_n1996_n452.t19 512.366
R21584 a_n1996_n452.n93 a_n1996_n452.t33 512.366
R21585 a_n1996_n452.n53 a_n1996_n452.t29 512.366
R21586 a_n1996_n452.n92 a_n1996_n452.t25 512.366
R21587 a_n1996_n452.n16 a_n1996_n452.t23 539.01
R21588 a_n1996_n452.n72 a_n1996_n452.t37 512.366
R21589 a_n1996_n452.n73 a_n1996_n452.t41 512.366
R21590 a_n1996_n452.n67 a_n1996_n452.t35 512.366
R21591 a_n1996_n452.n74 a_n1996_n452.t39 512.366
R21592 a_n1996_n452.n20 a_n1996_n452.t65 539.01
R21593 a_n1996_n452.n69 a_n1996_n452.t66 512.366
R21594 a_n1996_n452.n70 a_n1996_n452.t45 512.366
R21595 a_n1996_n452.n68 a_n1996_n452.t52 512.366
R21596 a_n1996_n452.n71 a_n1996_n452.t61 512.366
R21597 a_n1996_n452.n4 a_n1996_n452.n51 70.1674
R21598 a_n1996_n452.n6 a_n1996_n452.n49 70.1674
R21599 a_n1996_n452.n8 a_n1996_n452.n47 70.1674
R21600 a_n1996_n452.n11 a_n1996_n452.n45 70.1674
R21601 a_n1996_n452.n37 a_n1996_n452.n22 70.3058
R21602 a_n1996_n452.n31 a_n1996_n452.n34 70.1674
R21603 a_n1996_n452.n34 a_n1996_n452.n53 20.9683
R21604 a_n1996_n452.n33 a_n1996_n452.n32 75.0448
R21605 a_n1996_n452.n93 a_n1996_n452.n33 11.2134
R21606 a_n1996_n452.n25 a_n1996_n452.n26 44.8194
R21607 a_n1996_n452.n52 a_n1996_n452.n31 70.3058
R21608 a_n1996_n452.n23 a_n1996_n452.n36 70.1674
R21609 a_n1996_n452.n36 a_n1996_n452.n64 20.9683
R21610 a_n1996_n452.n35 a_n1996_n452.n23 75.0448
R21611 a_n1996_n452.n90 a_n1996_n452.n35 11.2134
R21612 a_n1996_n452.n21 a_n1996_n452.n24 44.8194
R21613 a_n1996_n452.n13 a_n1996_n452.n43 70.3058
R21614 a_n1996_n452.n17 a_n1996_n452.n40 70.3058
R21615 a_n1996_n452.n39 a_n1996_n452.n18 70.1674
R21616 a_n1996_n452.n39 a_n1996_n452.n68 20.9683
R21617 a_n1996_n452.n18 a_n1996_n452.n38 75.0448
R21618 a_n1996_n452.n70 a_n1996_n452.n38 11.2134
R21619 a_n1996_n452.n19 a_n1996_n452.n20 44.8194
R21620 a_n1996_n452.n42 a_n1996_n452.n14 70.1674
R21621 a_n1996_n452.n42 a_n1996_n452.n67 20.9683
R21622 a_n1996_n452.n14 a_n1996_n452.n41 75.0448
R21623 a_n1996_n452.n73 a_n1996_n452.n41 11.2134
R21624 a_n1996_n452.n15 a_n1996_n452.n16 44.8194
R21625 a_n1996_n452.n81 a_n1996_n452.n45 20.9683
R21626 a_n1996_n452.n44 a_n1996_n452.n12 75.0448
R21627 a_n1996_n452.n44 a_n1996_n452.n79 11.2134
R21628 a_n1996_n452.n12 a_n1996_n452.n80 161.3
R21629 a_n1996_n452.n83 a_n1996_n452.n47 20.9683
R21630 a_n1996_n452.n46 a_n1996_n452.n9 75.0448
R21631 a_n1996_n452.n46 a_n1996_n452.n78 11.2134
R21632 a_n1996_n452.n9 a_n1996_n452.n82 161.3
R21633 a_n1996_n452.n85 a_n1996_n452.n49 20.9683
R21634 a_n1996_n452.n48 a_n1996_n452.n7 75.0448
R21635 a_n1996_n452.n48 a_n1996_n452.n77 11.2134
R21636 a_n1996_n452.n7 a_n1996_n452.n84 161.3
R21637 a_n1996_n452.n87 a_n1996_n452.n51 20.9683
R21638 a_n1996_n452.n50 a_n1996_n452.n5 75.0448
R21639 a_n1996_n452.n50 a_n1996_n452.n76 11.2134
R21640 a_n1996_n452.n5 a_n1996_n452.n86 161.3
R21641 a_n1996_n452.n3 a_n1996_n452.n62 81.3764
R21642 a_n1996_n452.n1 a_n1996_n452.n57 81.3764
R21643 a_n1996_n452.n0 a_n1996_n452.n54 81.3764
R21644 a_n1996_n452.n3 a_n1996_n452.n63 80.9324
R21645 a_n1996_n452.n3 a_n1996_n452.n61 80.9324
R21646 a_n1996_n452.n2 a_n1996_n452.n60 80.9324
R21647 a_n1996_n452.n2 a_n1996_n452.n59 80.9324
R21648 a_n1996_n452.n1 a_n1996_n452.n58 80.9324
R21649 a_n1996_n452.n1 a_n1996_n452.n56 80.9324
R21650 a_n1996_n452.n0 a_n1996_n452.n55 80.9324
R21651 a_n1996_n452.n30 a_n1996_n452.t32 74.6477
R21652 a_n1996_n452.n27 a_n1996_n452.t24 74.6477
R21653 a_n1996_n452.n29 a_n1996_n452.t22 74.2899
R21654 a_n1996_n452.n28 a_n1996_n452.t28 74.2897
R21655 a_n1996_n452.n30 a_n1996_n452.n96 70.6783
R21656 a_n1996_n452.n28 a_n1996_n452.n66 70.6783
R21657 a_n1996_n452.n27 a_n1996_n452.n65 70.6783
R21658 a_n1996_n452.n97 a_n1996_n452.n30 70.6782
R21659 a_n1996_n452.n86 a_n1996_n452.n76 48.2005
R21660 a_n1996_n452.t64 a_n1996_n452.n51 533.335
R21661 a_n1996_n452.n84 a_n1996_n452.n77 48.2005
R21662 a_n1996_n452.t69 a_n1996_n452.n49 533.335
R21663 a_n1996_n452.n82 a_n1996_n452.n78 48.2005
R21664 a_n1996_n452.t58 a_n1996_n452.n47 533.335
R21665 a_n1996_n452.n80 a_n1996_n452.n79 48.2005
R21666 a_n1996_n452.t54 a_n1996_n452.n45 533.335
R21667 a_n1996_n452.n91 a_n1996_n452.n90 48.2005
R21668 a_n1996_n452.n89 a_n1996_n452.n36 20.9683
R21669 a_n1996_n452.n94 a_n1996_n452.n93 48.2005
R21670 a_n1996_n452.n92 a_n1996_n452.n34 20.9683
R21671 a_n1996_n452.n73 a_n1996_n452.n72 48.2005
R21672 a_n1996_n452.n74 a_n1996_n452.n42 20.9683
R21673 a_n1996_n452.n70 a_n1996_n452.n69 48.2005
R21674 a_n1996_n452.n71 a_n1996_n452.n39 20.9683
R21675 a_n1996_n452.n37 a_n1996_n452.t68 533.058
R21676 a_n1996_n452.t27 a_n1996_n452.n43 533.058
R21677 a_n1996_n452.t46 a_n1996_n452.n40 533.058
R21678 a_n1996_n452.n2 a_n1996_n452.n1 32.0139
R21679 a_n1996_n452.n87 a_n1996_n452.n50 35.3134
R21680 a_n1996_n452.n85 a_n1996_n452.n48 35.3134
R21681 a_n1996_n452.n83 a_n1996_n452.n46 35.3134
R21682 a_n1996_n452.n81 a_n1996_n452.n44 35.3134
R21683 a_n1996_n452.n35 a_n1996_n452.n64 35.3134
R21684 a_n1996_n452.n33 a_n1996_n452.n53 35.3134
R21685 a_n1996_n452.n67 a_n1996_n452.n41 35.3134
R21686 a_n1996_n452.n68 a_n1996_n452.n38 35.3134
R21687 a_n1996_n452.n31 a_n1996_n452.n3 23.891
R21688 a_n1996_n452.n19 a_n1996_n452.n10 12.046
R21689 a_n1996_n452.n22 a_n1996_n452.n88 11.8414
R21690 a_n1996_n452.n95 a_n1996_n452.n25 10.5365
R21691 a_n1996_n452.n75 a_n1996_n452.n28 9.50122
R21692 a_n1996_n452.n88 a_n1996_n452.n4 7.47588
R21693 a_n1996_n452.n12 a_n1996_n452.n10 7.47588
R21694 a_n1996_n452.n75 a_n1996_n452.n13 6.70126
R21695 a_n1996_n452.n29 a_n1996_n452.n95 5.65783
R21696 a_n1996_n452.n88 a_n1996_n452.n75 5.3452
R21697 a_n1996_n452.n31 a_n1996_n452.n21 3.95126
R21698 a_n1996_n452.n15 a_n1996_n452.n17 3.95126
R21699 a_n1996_n452.n96 a_n1996_n452.t30 3.61217
R21700 a_n1996_n452.n96 a_n1996_n452.t26 3.61217
R21701 a_n1996_n452.n66 a_n1996_n452.t36 3.61217
R21702 a_n1996_n452.n66 a_n1996_n452.t40 3.61217
R21703 a_n1996_n452.n65 a_n1996_n452.t38 3.61217
R21704 a_n1996_n452.n65 a_n1996_n452.t42 3.61217
R21705 a_n1996_n452.t20 a_n1996_n452.n97 3.61217
R21706 a_n1996_n452.n97 a_n1996_n452.t34 3.61217
R21707 a_n1996_n452.n62 a_n1996_n452.t13 2.82907
R21708 a_n1996_n452.n62 a_n1996_n452.t12 2.82907
R21709 a_n1996_n452.n63 a_n1996_n452.t10 2.82907
R21710 a_n1996_n452.n63 a_n1996_n452.t2 2.82907
R21711 a_n1996_n452.n61 a_n1996_n452.t1 2.82907
R21712 a_n1996_n452.n61 a_n1996_n452.t17 2.82907
R21713 a_n1996_n452.n60 a_n1996_n452.t14 2.82907
R21714 a_n1996_n452.n60 a_n1996_n452.t11 2.82907
R21715 a_n1996_n452.n59 a_n1996_n452.t43 2.82907
R21716 a_n1996_n452.n59 a_n1996_n452.t7 2.82907
R21717 a_n1996_n452.n57 a_n1996_n452.t3 2.82907
R21718 a_n1996_n452.n57 a_n1996_n452.t4 2.82907
R21719 a_n1996_n452.n58 a_n1996_n452.t9 2.82907
R21720 a_n1996_n452.n58 a_n1996_n452.t0 2.82907
R21721 a_n1996_n452.n56 a_n1996_n452.t18 2.82907
R21722 a_n1996_n452.n56 a_n1996_n452.t15 2.82907
R21723 a_n1996_n452.n55 a_n1996_n452.t8 2.82907
R21724 a_n1996_n452.n55 a_n1996_n452.t5 2.82907
R21725 a_n1996_n452.n54 a_n1996_n452.t16 2.82907
R21726 a_n1996_n452.n54 a_n1996_n452.t6 2.82907
R21727 a_n1996_n452.n95 a_n1996_n452.n10 1.30542
R21728 a_n1996_n452.n7 a_n1996_n452.n8 1.04595
R21729 a_n1996_n452.n24 a_n1996_n452.n91 13.657
R21730 a_n1996_n452.n89 a_n1996_n452.n37 21.4216
R21731 a_n1996_n452.n26 a_n1996_n452.n94 13.657
R21732 a_n1996_n452.n92 a_n1996_n452.n52 21.4216
R21733 a_n1996_n452.n72 a_n1996_n452.n16 13.657
R21734 a_n1996_n452.n43 a_n1996_n452.n74 21.4216
R21735 a_n1996_n452.n69 a_n1996_n452.n20 13.657
R21736 a_n1996_n452.n40 a_n1996_n452.n71 21.4216
R21737 a_n1996_n452.n3 a_n1996_n452.n2 1.3324
R21738 a_n1996_n452.n1 a_n1996_n452.n0 0.888431
R21739 a_n1996_n452.n32 a_n1996_n452.n25 0.758076
R21740 a_n1996_n452.n23 a_n1996_n452.n21 0.758076
R21741 a_n1996_n452.n23 a_n1996_n452.n22 0.758076
R21742 a_n1996_n452.n19 a_n1996_n452.n18 0.758076
R21743 a_n1996_n452.n18 a_n1996_n452.n17 0.758076
R21744 a_n1996_n452.n15 a_n1996_n452.n14 0.758076
R21745 a_n1996_n452.n14 a_n1996_n452.n13 0.758076
R21746 a_n1996_n452.n12 a_n1996_n452.n11 0.758076
R21747 a_n1996_n452.n9 a_n1996_n452.n8 0.758076
R21748 a_n1996_n452.n7 a_n1996_n452.n6 0.758076
R21749 a_n1996_n452.n5 a_n1996_n452.n4 0.758076
R21750 a_n1996_n452.n32 a_n1996_n452.n31 0.720197
R21751 a_n1996_n452.n30 a_n1996_n452.n29 0.716017
R21752 a_n1996_n452.n28 a_n1996_n452.n27 0.716017
R21753 a_n1996_n452.n9 a_n1996_n452.n11 0.67853
R21754 a_n1996_n452.n5 a_n1996_n452.n6 0.67853
R21755 a_n1808_13878.n2 a_n1808_13878.n0 98.9633
R21756 a_n1808_13878.n5 a_n1808_13878.n3 98.7517
R21757 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R21758 a_n1808_13878.n7 a_n1808_13878.n6 98.6055
R21759 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R21760 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R21761 a_n1808_13878.n9 a_n1808_13878.t1 74.6477
R21762 a_n1808_13878.n14 a_n1808_13878.t2 74.2899
R21763 a_n1808_13878.n11 a_n1808_13878.t3 74.2899
R21764 a_n1808_13878.n10 a_n1808_13878.t0 74.2899
R21765 a_n1808_13878.n13 a_n1808_13878.n12 70.6783
R21766 a_n1808_13878.n9 a_n1808_13878.n8 70.6783
R21767 a_n1808_13878.n15 a_n1808_13878.n7 13.5694
R21768 a_n1808_13878.n16 a_n1808_13878.n15 11.5762
R21769 a_n1808_13878.n15 a_n1808_13878.n14 6.2408
R21770 a_n1808_13878.n1 a_n1808_13878.t8 3.61217
R21771 a_n1808_13878.n1 a_n1808_13878.t13 3.61217
R21772 a_n1808_13878.n0 a_n1808_13878.t15 3.61217
R21773 a_n1808_13878.n0 a_n1808_13878.t19 3.61217
R21774 a_n1808_13878.n12 a_n1808_13878.t6 3.61217
R21775 a_n1808_13878.n12 a_n1808_13878.t7 3.61217
R21776 a_n1808_13878.n8 a_n1808_13878.t4 3.61217
R21777 a_n1808_13878.n8 a_n1808_13878.t5 3.61217
R21778 a_n1808_13878.n6 a_n1808_13878.t14 3.61217
R21779 a_n1808_13878.n6 a_n1808_13878.t9 3.61217
R21780 a_n1808_13878.n4 a_n1808_13878.t16 3.61217
R21781 a_n1808_13878.n4 a_n1808_13878.t11 3.61217
R21782 a_n1808_13878.n3 a_n1808_13878.t10 3.61217
R21783 a_n1808_13878.n3 a_n1808_13878.t12 3.61217
R21784 a_n1808_13878.n17 a_n1808_13878.t17 3.61217
R21785 a_n1808_13878.t18 a_n1808_13878.n17 3.61217
R21786 a_n1808_13878.n10 a_n1808_13878.n9 0.358259
R21787 a_n1808_13878.n13 a_n1808_13878.n11 0.358259
R21788 a_n1808_13878.n14 a_n1808_13878.n13 0.358259
R21789 a_n1808_13878.n16 a_n1808_13878.n2 0.358259
R21790 a_n1808_13878.n7 a_n1808_13878.n5 0.146627
R21791 a_n1808_13878.n11 a_n1808_13878.n10 0.101793
R21792 outputibias.n27 outputibias.n1 289.615
R21793 outputibias.n58 outputibias.n32 289.615
R21794 outputibias.n90 outputibias.n64 289.615
R21795 outputibias.n122 outputibias.n96 289.615
R21796 outputibias.n28 outputibias.n27 185
R21797 outputibias.n26 outputibias.n25 185
R21798 outputibias.n5 outputibias.n4 185
R21799 outputibias.n20 outputibias.n19 185
R21800 outputibias.n18 outputibias.n17 185
R21801 outputibias.n9 outputibias.n8 185
R21802 outputibias.n12 outputibias.n11 185
R21803 outputibias.n59 outputibias.n58 185
R21804 outputibias.n57 outputibias.n56 185
R21805 outputibias.n36 outputibias.n35 185
R21806 outputibias.n51 outputibias.n50 185
R21807 outputibias.n49 outputibias.n48 185
R21808 outputibias.n40 outputibias.n39 185
R21809 outputibias.n43 outputibias.n42 185
R21810 outputibias.n91 outputibias.n90 185
R21811 outputibias.n89 outputibias.n88 185
R21812 outputibias.n68 outputibias.n67 185
R21813 outputibias.n83 outputibias.n82 185
R21814 outputibias.n81 outputibias.n80 185
R21815 outputibias.n72 outputibias.n71 185
R21816 outputibias.n75 outputibias.n74 185
R21817 outputibias.n123 outputibias.n122 185
R21818 outputibias.n121 outputibias.n120 185
R21819 outputibias.n100 outputibias.n99 185
R21820 outputibias.n115 outputibias.n114 185
R21821 outputibias.n113 outputibias.n112 185
R21822 outputibias.n104 outputibias.n103 185
R21823 outputibias.n107 outputibias.n106 185
R21824 outputibias.n0 outputibias.t8 178.945
R21825 outputibias.n133 outputibias.t9 177.018
R21826 outputibias.n132 outputibias.t11 177.018
R21827 outputibias.n0 outputibias.t10 177.018
R21828 outputibias.t5 outputibias.n10 147.661
R21829 outputibias.t3 outputibias.n41 147.661
R21830 outputibias.t1 outputibias.n73 147.661
R21831 outputibias.t7 outputibias.n105 147.661
R21832 outputibias.n128 outputibias.t4 132.363
R21833 outputibias.n128 outputibias.t2 130.436
R21834 outputibias.n129 outputibias.t0 130.436
R21835 outputibias.n130 outputibias.t6 130.436
R21836 outputibias.n27 outputibias.n26 104.615
R21837 outputibias.n26 outputibias.n4 104.615
R21838 outputibias.n19 outputibias.n4 104.615
R21839 outputibias.n19 outputibias.n18 104.615
R21840 outputibias.n18 outputibias.n8 104.615
R21841 outputibias.n11 outputibias.n8 104.615
R21842 outputibias.n58 outputibias.n57 104.615
R21843 outputibias.n57 outputibias.n35 104.615
R21844 outputibias.n50 outputibias.n35 104.615
R21845 outputibias.n50 outputibias.n49 104.615
R21846 outputibias.n49 outputibias.n39 104.615
R21847 outputibias.n42 outputibias.n39 104.615
R21848 outputibias.n90 outputibias.n89 104.615
R21849 outputibias.n89 outputibias.n67 104.615
R21850 outputibias.n82 outputibias.n67 104.615
R21851 outputibias.n82 outputibias.n81 104.615
R21852 outputibias.n81 outputibias.n71 104.615
R21853 outputibias.n74 outputibias.n71 104.615
R21854 outputibias.n122 outputibias.n121 104.615
R21855 outputibias.n121 outputibias.n99 104.615
R21856 outputibias.n114 outputibias.n99 104.615
R21857 outputibias.n114 outputibias.n113 104.615
R21858 outputibias.n113 outputibias.n103 104.615
R21859 outputibias.n106 outputibias.n103 104.615
R21860 outputibias.n63 outputibias.n31 95.6354
R21861 outputibias.n63 outputibias.n62 94.6732
R21862 outputibias.n95 outputibias.n94 94.6732
R21863 outputibias.n127 outputibias.n126 94.6732
R21864 outputibias.n11 outputibias.t5 52.3082
R21865 outputibias.n42 outputibias.t3 52.3082
R21866 outputibias.n74 outputibias.t1 52.3082
R21867 outputibias.n106 outputibias.t7 52.3082
R21868 outputibias.n12 outputibias.n10 15.6674
R21869 outputibias.n43 outputibias.n41 15.6674
R21870 outputibias.n75 outputibias.n73 15.6674
R21871 outputibias.n107 outputibias.n105 15.6674
R21872 outputibias.n13 outputibias.n9 12.8005
R21873 outputibias.n44 outputibias.n40 12.8005
R21874 outputibias.n76 outputibias.n72 12.8005
R21875 outputibias.n108 outputibias.n104 12.8005
R21876 outputibias.n17 outputibias.n16 12.0247
R21877 outputibias.n48 outputibias.n47 12.0247
R21878 outputibias.n80 outputibias.n79 12.0247
R21879 outputibias.n112 outputibias.n111 12.0247
R21880 outputibias.n20 outputibias.n7 11.249
R21881 outputibias.n51 outputibias.n38 11.249
R21882 outputibias.n83 outputibias.n70 11.249
R21883 outputibias.n115 outputibias.n102 11.249
R21884 outputibias.n21 outputibias.n5 10.4732
R21885 outputibias.n52 outputibias.n36 10.4732
R21886 outputibias.n84 outputibias.n68 10.4732
R21887 outputibias.n116 outputibias.n100 10.4732
R21888 outputibias.n25 outputibias.n24 9.69747
R21889 outputibias.n56 outputibias.n55 9.69747
R21890 outputibias.n88 outputibias.n87 9.69747
R21891 outputibias.n120 outputibias.n119 9.69747
R21892 outputibias.n31 outputibias.n30 9.45567
R21893 outputibias.n62 outputibias.n61 9.45567
R21894 outputibias.n94 outputibias.n93 9.45567
R21895 outputibias.n126 outputibias.n125 9.45567
R21896 outputibias.n30 outputibias.n29 9.3005
R21897 outputibias.n3 outputibias.n2 9.3005
R21898 outputibias.n24 outputibias.n23 9.3005
R21899 outputibias.n22 outputibias.n21 9.3005
R21900 outputibias.n7 outputibias.n6 9.3005
R21901 outputibias.n16 outputibias.n15 9.3005
R21902 outputibias.n14 outputibias.n13 9.3005
R21903 outputibias.n61 outputibias.n60 9.3005
R21904 outputibias.n34 outputibias.n33 9.3005
R21905 outputibias.n55 outputibias.n54 9.3005
R21906 outputibias.n53 outputibias.n52 9.3005
R21907 outputibias.n38 outputibias.n37 9.3005
R21908 outputibias.n47 outputibias.n46 9.3005
R21909 outputibias.n45 outputibias.n44 9.3005
R21910 outputibias.n93 outputibias.n92 9.3005
R21911 outputibias.n66 outputibias.n65 9.3005
R21912 outputibias.n87 outputibias.n86 9.3005
R21913 outputibias.n85 outputibias.n84 9.3005
R21914 outputibias.n70 outputibias.n69 9.3005
R21915 outputibias.n79 outputibias.n78 9.3005
R21916 outputibias.n77 outputibias.n76 9.3005
R21917 outputibias.n125 outputibias.n124 9.3005
R21918 outputibias.n98 outputibias.n97 9.3005
R21919 outputibias.n119 outputibias.n118 9.3005
R21920 outputibias.n117 outputibias.n116 9.3005
R21921 outputibias.n102 outputibias.n101 9.3005
R21922 outputibias.n111 outputibias.n110 9.3005
R21923 outputibias.n109 outputibias.n108 9.3005
R21924 outputibias.n28 outputibias.n3 8.92171
R21925 outputibias.n59 outputibias.n34 8.92171
R21926 outputibias.n91 outputibias.n66 8.92171
R21927 outputibias.n123 outputibias.n98 8.92171
R21928 outputibias.n29 outputibias.n1 8.14595
R21929 outputibias.n60 outputibias.n32 8.14595
R21930 outputibias.n92 outputibias.n64 8.14595
R21931 outputibias.n124 outputibias.n96 8.14595
R21932 outputibias.n31 outputibias.n1 5.81868
R21933 outputibias.n62 outputibias.n32 5.81868
R21934 outputibias.n94 outputibias.n64 5.81868
R21935 outputibias.n126 outputibias.n96 5.81868
R21936 outputibias.n131 outputibias.n130 5.20947
R21937 outputibias.n29 outputibias.n28 5.04292
R21938 outputibias.n60 outputibias.n59 5.04292
R21939 outputibias.n92 outputibias.n91 5.04292
R21940 outputibias.n124 outputibias.n123 5.04292
R21941 outputibias.n131 outputibias.n127 4.42209
R21942 outputibias.n14 outputibias.n10 4.38594
R21943 outputibias.n45 outputibias.n41 4.38594
R21944 outputibias.n77 outputibias.n73 4.38594
R21945 outputibias.n109 outputibias.n105 4.38594
R21946 outputibias.n132 outputibias.n131 4.28454
R21947 outputibias.n25 outputibias.n3 4.26717
R21948 outputibias.n56 outputibias.n34 4.26717
R21949 outputibias.n88 outputibias.n66 4.26717
R21950 outputibias.n120 outputibias.n98 4.26717
R21951 outputibias.n24 outputibias.n5 3.49141
R21952 outputibias.n55 outputibias.n36 3.49141
R21953 outputibias.n87 outputibias.n68 3.49141
R21954 outputibias.n119 outputibias.n100 3.49141
R21955 outputibias.n21 outputibias.n20 2.71565
R21956 outputibias.n52 outputibias.n51 2.71565
R21957 outputibias.n84 outputibias.n83 2.71565
R21958 outputibias.n116 outputibias.n115 2.71565
R21959 outputibias.n17 outputibias.n7 1.93989
R21960 outputibias.n48 outputibias.n38 1.93989
R21961 outputibias.n80 outputibias.n70 1.93989
R21962 outputibias.n112 outputibias.n102 1.93989
R21963 outputibias.n130 outputibias.n129 1.9266
R21964 outputibias.n129 outputibias.n128 1.9266
R21965 outputibias.n133 outputibias.n132 1.92658
R21966 outputibias.n134 outputibias.n133 1.29913
R21967 outputibias.n16 outputibias.n9 1.16414
R21968 outputibias.n47 outputibias.n40 1.16414
R21969 outputibias.n79 outputibias.n72 1.16414
R21970 outputibias.n111 outputibias.n104 1.16414
R21971 outputibias.n127 outputibias.n95 0.962709
R21972 outputibias.n95 outputibias.n63 0.962709
R21973 outputibias.n13 outputibias.n12 0.388379
R21974 outputibias.n44 outputibias.n43 0.388379
R21975 outputibias.n76 outputibias.n75 0.388379
R21976 outputibias.n108 outputibias.n107 0.388379
R21977 outputibias.n134 outputibias.n0 0.337251
R21978 outputibias outputibias.n134 0.302375
R21979 outputibias.n30 outputibias.n2 0.155672
R21980 outputibias.n23 outputibias.n2 0.155672
R21981 outputibias.n23 outputibias.n22 0.155672
R21982 outputibias.n22 outputibias.n6 0.155672
R21983 outputibias.n15 outputibias.n6 0.155672
R21984 outputibias.n15 outputibias.n14 0.155672
R21985 outputibias.n61 outputibias.n33 0.155672
R21986 outputibias.n54 outputibias.n33 0.155672
R21987 outputibias.n54 outputibias.n53 0.155672
R21988 outputibias.n53 outputibias.n37 0.155672
R21989 outputibias.n46 outputibias.n37 0.155672
R21990 outputibias.n46 outputibias.n45 0.155672
R21991 outputibias.n93 outputibias.n65 0.155672
R21992 outputibias.n86 outputibias.n65 0.155672
R21993 outputibias.n86 outputibias.n85 0.155672
R21994 outputibias.n85 outputibias.n69 0.155672
R21995 outputibias.n78 outputibias.n69 0.155672
R21996 outputibias.n78 outputibias.n77 0.155672
R21997 outputibias.n125 outputibias.n97 0.155672
R21998 outputibias.n118 outputibias.n97 0.155672
R21999 outputibias.n118 outputibias.n117 0.155672
R22000 outputibias.n117 outputibias.n101 0.155672
R22001 outputibias.n110 outputibias.n101 0.155672
R22002 outputibias.n110 outputibias.n109 0.155672
R22003 diffpairibias.n0 diffpairibias.t27 436.822
R22004 diffpairibias.n27 diffpairibias.t24 435.479
R22005 diffpairibias.n26 diffpairibias.t21 435.479
R22006 diffpairibias.n25 diffpairibias.t22 435.479
R22007 diffpairibias.n24 diffpairibias.t26 435.479
R22008 diffpairibias.n23 diffpairibias.t20 435.479
R22009 diffpairibias.n0 diffpairibias.t23 435.479
R22010 diffpairibias.n1 diffpairibias.t28 435.479
R22011 diffpairibias.n2 diffpairibias.t25 435.479
R22012 diffpairibias.n3 diffpairibias.t29 435.479
R22013 diffpairibias.n13 diffpairibias.t14 377.536
R22014 diffpairibias.n13 diffpairibias.t0 376.193
R22015 diffpairibias.n14 diffpairibias.t10 376.193
R22016 diffpairibias.n15 diffpairibias.t12 376.193
R22017 diffpairibias.n16 diffpairibias.t6 376.193
R22018 diffpairibias.n17 diffpairibias.t2 376.193
R22019 diffpairibias.n18 diffpairibias.t16 376.193
R22020 diffpairibias.n19 diffpairibias.t4 376.193
R22021 diffpairibias.n20 diffpairibias.t18 376.193
R22022 diffpairibias.n21 diffpairibias.t8 376.193
R22023 diffpairibias.n4 diffpairibias.t15 113.368
R22024 diffpairibias.n4 diffpairibias.t1 112.698
R22025 diffpairibias.n5 diffpairibias.t11 112.698
R22026 diffpairibias.n6 diffpairibias.t13 112.698
R22027 diffpairibias.n7 diffpairibias.t7 112.698
R22028 diffpairibias.n8 diffpairibias.t3 112.698
R22029 diffpairibias.n9 diffpairibias.t17 112.698
R22030 diffpairibias.n10 diffpairibias.t5 112.698
R22031 diffpairibias.n11 diffpairibias.t19 112.698
R22032 diffpairibias.n12 diffpairibias.t9 112.698
R22033 diffpairibias.n22 diffpairibias.n21 4.77242
R22034 diffpairibias.n22 diffpairibias.n12 4.30807
R22035 diffpairibias.n23 diffpairibias.n22 4.13945
R22036 diffpairibias.n21 diffpairibias.n20 1.34352
R22037 diffpairibias.n20 diffpairibias.n19 1.34352
R22038 diffpairibias.n19 diffpairibias.n18 1.34352
R22039 diffpairibias.n18 diffpairibias.n17 1.34352
R22040 diffpairibias.n17 diffpairibias.n16 1.34352
R22041 diffpairibias.n16 diffpairibias.n15 1.34352
R22042 diffpairibias.n15 diffpairibias.n14 1.34352
R22043 diffpairibias.n14 diffpairibias.n13 1.34352
R22044 diffpairibias.n3 diffpairibias.n2 1.34352
R22045 diffpairibias.n2 diffpairibias.n1 1.34352
R22046 diffpairibias.n1 diffpairibias.n0 1.34352
R22047 diffpairibias.n24 diffpairibias.n23 1.34352
R22048 diffpairibias.n25 diffpairibias.n24 1.34352
R22049 diffpairibias.n26 diffpairibias.n25 1.34352
R22050 diffpairibias.n27 diffpairibias.n26 1.34352
R22051 diffpairibias.n28 diffpairibias.n27 0.862419
R22052 diffpairibias diffpairibias.n28 0.684875
R22053 diffpairibias.n12 diffpairibias.n11 0.672012
R22054 diffpairibias.n11 diffpairibias.n10 0.672012
R22055 diffpairibias.n10 diffpairibias.n9 0.672012
R22056 diffpairibias.n9 diffpairibias.n8 0.672012
R22057 diffpairibias.n8 diffpairibias.n7 0.672012
R22058 diffpairibias.n7 diffpairibias.n6 0.672012
R22059 diffpairibias.n6 diffpairibias.n5 0.672012
R22060 diffpairibias.n5 diffpairibias.n4 0.672012
R22061 diffpairibias.n28 diffpairibias.n3 0.190907
R22062 commonsourceibias.n281 commonsourceibias.t101 222.032
R22063 commonsourceibias.n44 commonsourceibias.t78 222.032
R22064 commonsourceibias.n166 commonsourceibias.t117 222.032
R22065 commonsourceibias.n643 commonsourceibias.t106 222.032
R22066 commonsourceibias.n413 commonsourceibias.t28 222.032
R22067 commonsourceibias.n529 commonsourceibias.t123 222.032
R22068 commonsourceibias.n364 commonsourceibias.t100 207.983
R22069 commonsourceibias.n127 commonsourceibias.t74 207.983
R22070 commonsourceibias.n249 commonsourceibias.t115 207.983
R22071 commonsourceibias.n731 commonsourceibias.t122 207.983
R22072 commonsourceibias.n501 commonsourceibias.t14 207.983
R22073 commonsourceibias.n616 commonsourceibias.t140 207.983
R22074 commonsourceibias.n280 commonsourceibias.t87 168.701
R22075 commonsourceibias.n286 commonsourceibias.t129 168.701
R22076 commonsourceibias.n292 commonsourceibias.t110 168.701
R22077 commonsourceibias.n276 commonsourceibias.t93 168.701
R22078 commonsourceibias.n300 commonsourceibias.t95 168.701
R22079 commonsourceibias.n306 commonsourceibias.t121 168.701
R22080 commonsourceibias.n271 commonsourceibias.t102 168.701
R22081 commonsourceibias.n314 commonsourceibias.t108 168.701
R22082 commonsourceibias.n320 commonsourceibias.t159 168.701
R22083 commonsourceibias.n266 commonsourceibias.t138 168.701
R22084 commonsourceibias.n328 commonsourceibias.t118 168.701
R22085 commonsourceibias.n334 commonsourceibias.t83 168.701
R22086 commonsourceibias.n261 commonsourceibias.t86 168.701
R22087 commonsourceibias.n342 commonsourceibias.t128 168.701
R22088 commonsourceibias.n348 commonsourceibias.t109 168.701
R22089 commonsourceibias.n256 commonsourceibias.t92 168.701
R22090 commonsourceibias.n356 commonsourceibias.t137 168.701
R22091 commonsourceibias.n362 commonsourceibias.t119 168.701
R22092 commonsourceibias.n125 commonsourceibias.t20 168.701
R22093 commonsourceibias.n119 commonsourceibias.t50 168.701
R22094 commonsourceibias.n19 commonsourceibias.t8 168.701
R22095 commonsourceibias.n111 commonsourceibias.t36 168.701
R22096 commonsourceibias.n105 commonsourceibias.t76 168.701
R22097 commonsourceibias.n24 commonsourceibias.t24 168.701
R22098 commonsourceibias.n97 commonsourceibias.t34 168.701
R22099 commonsourceibias.n91 commonsourceibias.t10 168.701
R22100 commonsourceibias.n29 commonsourceibias.t40 168.701
R22101 commonsourceibias.n83 commonsourceibias.t56 168.701
R22102 commonsourceibias.n77 commonsourceibias.t26 168.701
R22103 commonsourceibias.n34 commonsourceibias.t38 168.701
R22104 commonsourceibias.n69 commonsourceibias.t70 168.701
R22105 commonsourceibias.n63 commonsourceibias.t18 168.701
R22106 commonsourceibias.n39 commonsourceibias.t22 168.701
R22107 commonsourceibias.n55 commonsourceibias.t54 168.701
R22108 commonsourceibias.n49 commonsourceibias.t4 168.701
R22109 commonsourceibias.n43 commonsourceibias.t46 168.701
R22110 commonsourceibias.n247 commonsourceibias.t136 168.701
R22111 commonsourceibias.n241 commonsourceibias.t151 168.701
R22112 commonsourceibias.n5 commonsourceibias.t105 168.701
R22113 commonsourceibias.n233 commonsourceibias.t126 168.701
R22114 commonsourceibias.n227 commonsourceibias.t144 168.701
R22115 commonsourceibias.n10 commonsourceibias.t98 168.701
R22116 commonsourceibias.n219 commonsourceibias.t94 168.701
R22117 commonsourceibias.n213 commonsourceibias.t135 168.701
R22118 commonsourceibias.n150 commonsourceibias.t153 168.701
R22119 commonsourceibias.n151 commonsourceibias.t88 168.701
R22120 commonsourceibias.n153 commonsourceibias.t125 168.701
R22121 commonsourceibias.n155 commonsourceibias.t120 168.701
R22122 commonsourceibias.n191 commonsourceibias.t139 168.701
R22123 commonsourceibias.n185 commonsourceibias.t112 168.701
R22124 commonsourceibias.n161 commonsourceibias.t107 168.701
R22125 commonsourceibias.n177 commonsourceibias.t127 168.701
R22126 commonsourceibias.n171 commonsourceibias.t146 168.701
R22127 commonsourceibias.n165 commonsourceibias.t99 168.701
R22128 commonsourceibias.n642 commonsourceibias.t90 168.701
R22129 commonsourceibias.n648 commonsourceibias.t134 168.701
R22130 commonsourceibias.n654 commonsourceibias.t116 168.701
R22131 commonsourceibias.n656 commonsourceibias.t96 168.701
R22132 commonsourceibias.n663 commonsourceibias.t91 168.701
R22133 commonsourceibias.n669 commonsourceibias.t145 168.701
R22134 commonsourceibias.n671 commonsourceibias.t124 168.701
R22135 commonsourceibias.n678 commonsourceibias.t131 168.701
R22136 commonsourceibias.n684 commonsourceibias.t152 168.701
R22137 commonsourceibias.n686 commonsourceibias.t157 168.701
R22138 commonsourceibias.n693 commonsourceibias.t141 168.701
R22139 commonsourceibias.n699 commonsourceibias.t97 168.701
R22140 commonsourceibias.n701 commonsourceibias.t81 168.701
R22141 commonsourceibias.n708 commonsourceibias.t149 168.701
R22142 commonsourceibias.n714 commonsourceibias.t132 168.701
R22143 commonsourceibias.n716 commonsourceibias.t111 168.701
R22144 commonsourceibias.n723 commonsourceibias.t156 168.701
R22145 commonsourceibias.n729 commonsourceibias.t142 168.701
R22146 commonsourceibias.n412 commonsourceibias.t2 168.701
R22147 commonsourceibias.n418 commonsourceibias.t48 168.701
R22148 commonsourceibias.n424 commonsourceibias.t12 168.701
R22149 commonsourceibias.n426 commonsourceibias.t68 168.701
R22150 commonsourceibias.n433 commonsourceibias.t66 168.701
R22151 commonsourceibias.n439 commonsourceibias.t6 168.701
R22152 commonsourceibias.n441 commonsourceibias.t62 168.701
R22153 commonsourceibias.n448 commonsourceibias.t52 168.701
R22154 commonsourceibias.n454 commonsourceibias.t72 168.701
R22155 commonsourceibias.n456 commonsourceibias.t64 168.701
R22156 commonsourceibias.n463 commonsourceibias.t32 168.701
R22157 commonsourceibias.n469 commonsourceibias.t58 168.701
R22158 commonsourceibias.n471 commonsourceibias.t44 168.701
R22159 commonsourceibias.n478 commonsourceibias.t16 168.701
R22160 commonsourceibias.n484 commonsourceibias.t60 168.701
R22161 commonsourceibias.n486 commonsourceibias.t30 168.701
R22162 commonsourceibias.n493 commonsourceibias.t0 168.701
R22163 commonsourceibias.n499 commonsourceibias.t42 168.701
R22164 commonsourceibias.n614 commonsourceibias.t155 168.701
R22165 commonsourceibias.n608 commonsourceibias.t84 168.701
R22166 commonsourceibias.n601 commonsourceibias.t130 168.701
R22167 commonsourceibias.n599 commonsourceibias.t148 168.701
R22168 commonsourceibias.n593 commonsourceibias.t80 168.701
R22169 commonsourceibias.n586 commonsourceibias.t89 168.701
R22170 commonsourceibias.n584 commonsourceibias.t113 168.701
R22171 commonsourceibias.n578 commonsourceibias.t154 168.701
R22172 commonsourceibias.n571 commonsourceibias.t85 168.701
R22173 commonsourceibias.n528 commonsourceibias.t103 168.701
R22174 commonsourceibias.n534 commonsourceibias.t150 168.701
R22175 commonsourceibias.n540 commonsourceibias.t133 168.701
R22176 commonsourceibias.n542 commonsourceibias.t114 168.701
R22177 commonsourceibias.n549 commonsourceibias.t104 168.701
R22178 commonsourceibias.n555 commonsourceibias.t158 168.701
R22179 commonsourceibias.n519 commonsourceibias.t143 168.701
R22180 commonsourceibias.n517 commonsourceibias.t147 168.701
R22181 commonsourceibias.n515 commonsourceibias.t82 168.701
R22182 commonsourceibias.n363 commonsourceibias.n251 161.3
R22183 commonsourceibias.n361 commonsourceibias.n360 161.3
R22184 commonsourceibias.n359 commonsourceibias.n252 161.3
R22185 commonsourceibias.n358 commonsourceibias.n357 161.3
R22186 commonsourceibias.n355 commonsourceibias.n253 161.3
R22187 commonsourceibias.n354 commonsourceibias.n353 161.3
R22188 commonsourceibias.n352 commonsourceibias.n254 161.3
R22189 commonsourceibias.n351 commonsourceibias.n350 161.3
R22190 commonsourceibias.n349 commonsourceibias.n255 161.3
R22191 commonsourceibias.n347 commonsourceibias.n346 161.3
R22192 commonsourceibias.n345 commonsourceibias.n257 161.3
R22193 commonsourceibias.n344 commonsourceibias.n343 161.3
R22194 commonsourceibias.n341 commonsourceibias.n258 161.3
R22195 commonsourceibias.n340 commonsourceibias.n339 161.3
R22196 commonsourceibias.n338 commonsourceibias.n259 161.3
R22197 commonsourceibias.n337 commonsourceibias.n336 161.3
R22198 commonsourceibias.n335 commonsourceibias.n260 161.3
R22199 commonsourceibias.n333 commonsourceibias.n332 161.3
R22200 commonsourceibias.n331 commonsourceibias.n262 161.3
R22201 commonsourceibias.n330 commonsourceibias.n329 161.3
R22202 commonsourceibias.n327 commonsourceibias.n263 161.3
R22203 commonsourceibias.n326 commonsourceibias.n325 161.3
R22204 commonsourceibias.n324 commonsourceibias.n264 161.3
R22205 commonsourceibias.n323 commonsourceibias.n322 161.3
R22206 commonsourceibias.n321 commonsourceibias.n265 161.3
R22207 commonsourceibias.n319 commonsourceibias.n318 161.3
R22208 commonsourceibias.n317 commonsourceibias.n267 161.3
R22209 commonsourceibias.n316 commonsourceibias.n315 161.3
R22210 commonsourceibias.n313 commonsourceibias.n268 161.3
R22211 commonsourceibias.n312 commonsourceibias.n311 161.3
R22212 commonsourceibias.n310 commonsourceibias.n269 161.3
R22213 commonsourceibias.n309 commonsourceibias.n308 161.3
R22214 commonsourceibias.n307 commonsourceibias.n270 161.3
R22215 commonsourceibias.n305 commonsourceibias.n304 161.3
R22216 commonsourceibias.n303 commonsourceibias.n272 161.3
R22217 commonsourceibias.n302 commonsourceibias.n301 161.3
R22218 commonsourceibias.n299 commonsourceibias.n273 161.3
R22219 commonsourceibias.n298 commonsourceibias.n297 161.3
R22220 commonsourceibias.n296 commonsourceibias.n274 161.3
R22221 commonsourceibias.n295 commonsourceibias.n294 161.3
R22222 commonsourceibias.n293 commonsourceibias.n275 161.3
R22223 commonsourceibias.n291 commonsourceibias.n290 161.3
R22224 commonsourceibias.n289 commonsourceibias.n277 161.3
R22225 commonsourceibias.n288 commonsourceibias.n287 161.3
R22226 commonsourceibias.n285 commonsourceibias.n278 161.3
R22227 commonsourceibias.n284 commonsourceibias.n283 161.3
R22228 commonsourceibias.n282 commonsourceibias.n279 161.3
R22229 commonsourceibias.n45 commonsourceibias.n42 161.3
R22230 commonsourceibias.n47 commonsourceibias.n46 161.3
R22231 commonsourceibias.n48 commonsourceibias.n41 161.3
R22232 commonsourceibias.n51 commonsourceibias.n50 161.3
R22233 commonsourceibias.n52 commonsourceibias.n40 161.3
R22234 commonsourceibias.n54 commonsourceibias.n53 161.3
R22235 commonsourceibias.n56 commonsourceibias.n38 161.3
R22236 commonsourceibias.n58 commonsourceibias.n57 161.3
R22237 commonsourceibias.n59 commonsourceibias.n37 161.3
R22238 commonsourceibias.n61 commonsourceibias.n60 161.3
R22239 commonsourceibias.n62 commonsourceibias.n36 161.3
R22240 commonsourceibias.n65 commonsourceibias.n64 161.3
R22241 commonsourceibias.n66 commonsourceibias.n35 161.3
R22242 commonsourceibias.n68 commonsourceibias.n67 161.3
R22243 commonsourceibias.n70 commonsourceibias.n33 161.3
R22244 commonsourceibias.n72 commonsourceibias.n71 161.3
R22245 commonsourceibias.n73 commonsourceibias.n32 161.3
R22246 commonsourceibias.n75 commonsourceibias.n74 161.3
R22247 commonsourceibias.n76 commonsourceibias.n31 161.3
R22248 commonsourceibias.n79 commonsourceibias.n78 161.3
R22249 commonsourceibias.n80 commonsourceibias.n30 161.3
R22250 commonsourceibias.n82 commonsourceibias.n81 161.3
R22251 commonsourceibias.n84 commonsourceibias.n28 161.3
R22252 commonsourceibias.n86 commonsourceibias.n85 161.3
R22253 commonsourceibias.n87 commonsourceibias.n27 161.3
R22254 commonsourceibias.n89 commonsourceibias.n88 161.3
R22255 commonsourceibias.n90 commonsourceibias.n26 161.3
R22256 commonsourceibias.n93 commonsourceibias.n92 161.3
R22257 commonsourceibias.n94 commonsourceibias.n25 161.3
R22258 commonsourceibias.n96 commonsourceibias.n95 161.3
R22259 commonsourceibias.n98 commonsourceibias.n23 161.3
R22260 commonsourceibias.n100 commonsourceibias.n99 161.3
R22261 commonsourceibias.n101 commonsourceibias.n22 161.3
R22262 commonsourceibias.n103 commonsourceibias.n102 161.3
R22263 commonsourceibias.n104 commonsourceibias.n21 161.3
R22264 commonsourceibias.n107 commonsourceibias.n106 161.3
R22265 commonsourceibias.n108 commonsourceibias.n20 161.3
R22266 commonsourceibias.n110 commonsourceibias.n109 161.3
R22267 commonsourceibias.n112 commonsourceibias.n18 161.3
R22268 commonsourceibias.n114 commonsourceibias.n113 161.3
R22269 commonsourceibias.n115 commonsourceibias.n17 161.3
R22270 commonsourceibias.n117 commonsourceibias.n116 161.3
R22271 commonsourceibias.n118 commonsourceibias.n16 161.3
R22272 commonsourceibias.n121 commonsourceibias.n120 161.3
R22273 commonsourceibias.n122 commonsourceibias.n15 161.3
R22274 commonsourceibias.n124 commonsourceibias.n123 161.3
R22275 commonsourceibias.n126 commonsourceibias.n14 161.3
R22276 commonsourceibias.n167 commonsourceibias.n164 161.3
R22277 commonsourceibias.n169 commonsourceibias.n168 161.3
R22278 commonsourceibias.n170 commonsourceibias.n163 161.3
R22279 commonsourceibias.n173 commonsourceibias.n172 161.3
R22280 commonsourceibias.n174 commonsourceibias.n162 161.3
R22281 commonsourceibias.n176 commonsourceibias.n175 161.3
R22282 commonsourceibias.n178 commonsourceibias.n160 161.3
R22283 commonsourceibias.n180 commonsourceibias.n179 161.3
R22284 commonsourceibias.n181 commonsourceibias.n159 161.3
R22285 commonsourceibias.n183 commonsourceibias.n182 161.3
R22286 commonsourceibias.n184 commonsourceibias.n158 161.3
R22287 commonsourceibias.n187 commonsourceibias.n186 161.3
R22288 commonsourceibias.n188 commonsourceibias.n157 161.3
R22289 commonsourceibias.n190 commonsourceibias.n189 161.3
R22290 commonsourceibias.n192 commonsourceibias.n156 161.3
R22291 commonsourceibias.n194 commonsourceibias.n193 161.3
R22292 commonsourceibias.n196 commonsourceibias.n195 161.3
R22293 commonsourceibias.n197 commonsourceibias.n154 161.3
R22294 commonsourceibias.n199 commonsourceibias.n198 161.3
R22295 commonsourceibias.n201 commonsourceibias.n200 161.3
R22296 commonsourceibias.n202 commonsourceibias.n152 161.3
R22297 commonsourceibias.n204 commonsourceibias.n203 161.3
R22298 commonsourceibias.n206 commonsourceibias.n205 161.3
R22299 commonsourceibias.n208 commonsourceibias.n207 161.3
R22300 commonsourceibias.n209 commonsourceibias.n13 161.3
R22301 commonsourceibias.n211 commonsourceibias.n210 161.3
R22302 commonsourceibias.n212 commonsourceibias.n12 161.3
R22303 commonsourceibias.n215 commonsourceibias.n214 161.3
R22304 commonsourceibias.n216 commonsourceibias.n11 161.3
R22305 commonsourceibias.n218 commonsourceibias.n217 161.3
R22306 commonsourceibias.n220 commonsourceibias.n9 161.3
R22307 commonsourceibias.n222 commonsourceibias.n221 161.3
R22308 commonsourceibias.n223 commonsourceibias.n8 161.3
R22309 commonsourceibias.n225 commonsourceibias.n224 161.3
R22310 commonsourceibias.n226 commonsourceibias.n7 161.3
R22311 commonsourceibias.n229 commonsourceibias.n228 161.3
R22312 commonsourceibias.n230 commonsourceibias.n6 161.3
R22313 commonsourceibias.n232 commonsourceibias.n231 161.3
R22314 commonsourceibias.n234 commonsourceibias.n4 161.3
R22315 commonsourceibias.n236 commonsourceibias.n235 161.3
R22316 commonsourceibias.n237 commonsourceibias.n3 161.3
R22317 commonsourceibias.n239 commonsourceibias.n238 161.3
R22318 commonsourceibias.n240 commonsourceibias.n2 161.3
R22319 commonsourceibias.n243 commonsourceibias.n242 161.3
R22320 commonsourceibias.n244 commonsourceibias.n1 161.3
R22321 commonsourceibias.n246 commonsourceibias.n245 161.3
R22322 commonsourceibias.n248 commonsourceibias.n0 161.3
R22323 commonsourceibias.n730 commonsourceibias.n618 161.3
R22324 commonsourceibias.n728 commonsourceibias.n727 161.3
R22325 commonsourceibias.n726 commonsourceibias.n619 161.3
R22326 commonsourceibias.n725 commonsourceibias.n724 161.3
R22327 commonsourceibias.n722 commonsourceibias.n620 161.3
R22328 commonsourceibias.n721 commonsourceibias.n720 161.3
R22329 commonsourceibias.n719 commonsourceibias.n621 161.3
R22330 commonsourceibias.n718 commonsourceibias.n717 161.3
R22331 commonsourceibias.n715 commonsourceibias.n622 161.3
R22332 commonsourceibias.n713 commonsourceibias.n712 161.3
R22333 commonsourceibias.n711 commonsourceibias.n623 161.3
R22334 commonsourceibias.n710 commonsourceibias.n709 161.3
R22335 commonsourceibias.n707 commonsourceibias.n624 161.3
R22336 commonsourceibias.n706 commonsourceibias.n705 161.3
R22337 commonsourceibias.n704 commonsourceibias.n625 161.3
R22338 commonsourceibias.n703 commonsourceibias.n702 161.3
R22339 commonsourceibias.n700 commonsourceibias.n626 161.3
R22340 commonsourceibias.n698 commonsourceibias.n697 161.3
R22341 commonsourceibias.n696 commonsourceibias.n627 161.3
R22342 commonsourceibias.n695 commonsourceibias.n694 161.3
R22343 commonsourceibias.n692 commonsourceibias.n628 161.3
R22344 commonsourceibias.n691 commonsourceibias.n690 161.3
R22345 commonsourceibias.n689 commonsourceibias.n629 161.3
R22346 commonsourceibias.n688 commonsourceibias.n687 161.3
R22347 commonsourceibias.n685 commonsourceibias.n630 161.3
R22348 commonsourceibias.n683 commonsourceibias.n682 161.3
R22349 commonsourceibias.n681 commonsourceibias.n631 161.3
R22350 commonsourceibias.n680 commonsourceibias.n679 161.3
R22351 commonsourceibias.n677 commonsourceibias.n632 161.3
R22352 commonsourceibias.n676 commonsourceibias.n675 161.3
R22353 commonsourceibias.n674 commonsourceibias.n633 161.3
R22354 commonsourceibias.n673 commonsourceibias.n672 161.3
R22355 commonsourceibias.n670 commonsourceibias.n634 161.3
R22356 commonsourceibias.n668 commonsourceibias.n667 161.3
R22357 commonsourceibias.n666 commonsourceibias.n635 161.3
R22358 commonsourceibias.n665 commonsourceibias.n664 161.3
R22359 commonsourceibias.n662 commonsourceibias.n636 161.3
R22360 commonsourceibias.n661 commonsourceibias.n660 161.3
R22361 commonsourceibias.n659 commonsourceibias.n637 161.3
R22362 commonsourceibias.n658 commonsourceibias.n657 161.3
R22363 commonsourceibias.n655 commonsourceibias.n638 161.3
R22364 commonsourceibias.n653 commonsourceibias.n652 161.3
R22365 commonsourceibias.n651 commonsourceibias.n639 161.3
R22366 commonsourceibias.n650 commonsourceibias.n649 161.3
R22367 commonsourceibias.n647 commonsourceibias.n640 161.3
R22368 commonsourceibias.n646 commonsourceibias.n645 161.3
R22369 commonsourceibias.n644 commonsourceibias.n641 161.3
R22370 commonsourceibias.n500 commonsourceibias.n388 161.3
R22371 commonsourceibias.n498 commonsourceibias.n497 161.3
R22372 commonsourceibias.n496 commonsourceibias.n389 161.3
R22373 commonsourceibias.n495 commonsourceibias.n494 161.3
R22374 commonsourceibias.n492 commonsourceibias.n390 161.3
R22375 commonsourceibias.n491 commonsourceibias.n490 161.3
R22376 commonsourceibias.n489 commonsourceibias.n391 161.3
R22377 commonsourceibias.n488 commonsourceibias.n487 161.3
R22378 commonsourceibias.n485 commonsourceibias.n392 161.3
R22379 commonsourceibias.n483 commonsourceibias.n482 161.3
R22380 commonsourceibias.n481 commonsourceibias.n393 161.3
R22381 commonsourceibias.n480 commonsourceibias.n479 161.3
R22382 commonsourceibias.n477 commonsourceibias.n394 161.3
R22383 commonsourceibias.n476 commonsourceibias.n475 161.3
R22384 commonsourceibias.n474 commonsourceibias.n395 161.3
R22385 commonsourceibias.n473 commonsourceibias.n472 161.3
R22386 commonsourceibias.n470 commonsourceibias.n396 161.3
R22387 commonsourceibias.n468 commonsourceibias.n467 161.3
R22388 commonsourceibias.n466 commonsourceibias.n397 161.3
R22389 commonsourceibias.n465 commonsourceibias.n464 161.3
R22390 commonsourceibias.n462 commonsourceibias.n398 161.3
R22391 commonsourceibias.n461 commonsourceibias.n460 161.3
R22392 commonsourceibias.n459 commonsourceibias.n399 161.3
R22393 commonsourceibias.n458 commonsourceibias.n457 161.3
R22394 commonsourceibias.n455 commonsourceibias.n400 161.3
R22395 commonsourceibias.n453 commonsourceibias.n452 161.3
R22396 commonsourceibias.n451 commonsourceibias.n401 161.3
R22397 commonsourceibias.n450 commonsourceibias.n449 161.3
R22398 commonsourceibias.n447 commonsourceibias.n402 161.3
R22399 commonsourceibias.n446 commonsourceibias.n445 161.3
R22400 commonsourceibias.n444 commonsourceibias.n403 161.3
R22401 commonsourceibias.n443 commonsourceibias.n442 161.3
R22402 commonsourceibias.n440 commonsourceibias.n404 161.3
R22403 commonsourceibias.n438 commonsourceibias.n437 161.3
R22404 commonsourceibias.n436 commonsourceibias.n405 161.3
R22405 commonsourceibias.n435 commonsourceibias.n434 161.3
R22406 commonsourceibias.n432 commonsourceibias.n406 161.3
R22407 commonsourceibias.n431 commonsourceibias.n430 161.3
R22408 commonsourceibias.n429 commonsourceibias.n407 161.3
R22409 commonsourceibias.n428 commonsourceibias.n427 161.3
R22410 commonsourceibias.n425 commonsourceibias.n408 161.3
R22411 commonsourceibias.n423 commonsourceibias.n422 161.3
R22412 commonsourceibias.n421 commonsourceibias.n409 161.3
R22413 commonsourceibias.n420 commonsourceibias.n419 161.3
R22414 commonsourceibias.n417 commonsourceibias.n410 161.3
R22415 commonsourceibias.n416 commonsourceibias.n415 161.3
R22416 commonsourceibias.n414 commonsourceibias.n411 161.3
R22417 commonsourceibias.n570 commonsourceibias.n569 161.3
R22418 commonsourceibias.n568 commonsourceibias.n567 161.3
R22419 commonsourceibias.n566 commonsourceibias.n516 161.3
R22420 commonsourceibias.n565 commonsourceibias.n564 161.3
R22421 commonsourceibias.n563 commonsourceibias.n562 161.3
R22422 commonsourceibias.n561 commonsourceibias.n518 161.3
R22423 commonsourceibias.n560 commonsourceibias.n559 161.3
R22424 commonsourceibias.n558 commonsourceibias.n557 161.3
R22425 commonsourceibias.n556 commonsourceibias.n520 161.3
R22426 commonsourceibias.n554 commonsourceibias.n553 161.3
R22427 commonsourceibias.n552 commonsourceibias.n521 161.3
R22428 commonsourceibias.n551 commonsourceibias.n550 161.3
R22429 commonsourceibias.n548 commonsourceibias.n522 161.3
R22430 commonsourceibias.n547 commonsourceibias.n546 161.3
R22431 commonsourceibias.n545 commonsourceibias.n523 161.3
R22432 commonsourceibias.n544 commonsourceibias.n543 161.3
R22433 commonsourceibias.n541 commonsourceibias.n524 161.3
R22434 commonsourceibias.n539 commonsourceibias.n538 161.3
R22435 commonsourceibias.n537 commonsourceibias.n525 161.3
R22436 commonsourceibias.n536 commonsourceibias.n535 161.3
R22437 commonsourceibias.n533 commonsourceibias.n526 161.3
R22438 commonsourceibias.n532 commonsourceibias.n531 161.3
R22439 commonsourceibias.n530 commonsourceibias.n527 161.3
R22440 commonsourceibias.n615 commonsourceibias.n367 161.3
R22441 commonsourceibias.n613 commonsourceibias.n612 161.3
R22442 commonsourceibias.n611 commonsourceibias.n368 161.3
R22443 commonsourceibias.n610 commonsourceibias.n609 161.3
R22444 commonsourceibias.n607 commonsourceibias.n369 161.3
R22445 commonsourceibias.n606 commonsourceibias.n605 161.3
R22446 commonsourceibias.n604 commonsourceibias.n370 161.3
R22447 commonsourceibias.n603 commonsourceibias.n602 161.3
R22448 commonsourceibias.n600 commonsourceibias.n371 161.3
R22449 commonsourceibias.n598 commonsourceibias.n597 161.3
R22450 commonsourceibias.n596 commonsourceibias.n372 161.3
R22451 commonsourceibias.n595 commonsourceibias.n594 161.3
R22452 commonsourceibias.n592 commonsourceibias.n373 161.3
R22453 commonsourceibias.n591 commonsourceibias.n590 161.3
R22454 commonsourceibias.n589 commonsourceibias.n374 161.3
R22455 commonsourceibias.n588 commonsourceibias.n587 161.3
R22456 commonsourceibias.n585 commonsourceibias.n375 161.3
R22457 commonsourceibias.n583 commonsourceibias.n582 161.3
R22458 commonsourceibias.n581 commonsourceibias.n376 161.3
R22459 commonsourceibias.n580 commonsourceibias.n579 161.3
R22460 commonsourceibias.n577 commonsourceibias.n377 161.3
R22461 commonsourceibias.n576 commonsourceibias.n575 161.3
R22462 commonsourceibias.n574 commonsourceibias.n378 161.3
R22463 commonsourceibias.n573 commonsourceibias.n572 161.3
R22464 commonsourceibias.n141 commonsourceibias.n139 81.5057
R22465 commonsourceibias.n381 commonsourceibias.n379 81.5057
R22466 commonsourceibias.n141 commonsourceibias.n140 80.9324
R22467 commonsourceibias.n143 commonsourceibias.n142 80.9324
R22468 commonsourceibias.n145 commonsourceibias.n144 80.9324
R22469 commonsourceibias.n147 commonsourceibias.n146 80.9324
R22470 commonsourceibias.n138 commonsourceibias.n137 80.9324
R22471 commonsourceibias.n136 commonsourceibias.n135 80.9324
R22472 commonsourceibias.n134 commonsourceibias.n133 80.9324
R22473 commonsourceibias.n132 commonsourceibias.n131 80.9324
R22474 commonsourceibias.n130 commonsourceibias.n129 80.9324
R22475 commonsourceibias.n504 commonsourceibias.n503 80.9324
R22476 commonsourceibias.n506 commonsourceibias.n505 80.9324
R22477 commonsourceibias.n508 commonsourceibias.n507 80.9324
R22478 commonsourceibias.n510 commonsourceibias.n509 80.9324
R22479 commonsourceibias.n512 commonsourceibias.n511 80.9324
R22480 commonsourceibias.n387 commonsourceibias.n386 80.9324
R22481 commonsourceibias.n385 commonsourceibias.n384 80.9324
R22482 commonsourceibias.n383 commonsourceibias.n382 80.9324
R22483 commonsourceibias.n381 commonsourceibias.n380 80.9324
R22484 commonsourceibias.n365 commonsourceibias.n364 80.6037
R22485 commonsourceibias.n128 commonsourceibias.n127 80.6037
R22486 commonsourceibias.n250 commonsourceibias.n249 80.6037
R22487 commonsourceibias.n732 commonsourceibias.n731 80.6037
R22488 commonsourceibias.n502 commonsourceibias.n501 80.6037
R22489 commonsourceibias.n617 commonsourceibias.n616 80.6037
R22490 commonsourceibias.n322 commonsourceibias.n321 56.5617
R22491 commonsourceibias.n336 commonsourceibias.n335 56.5617
R22492 commonsourceibias.n85 commonsourceibias.n84 56.5617
R22493 commonsourceibias.n71 commonsourceibias.n70 56.5617
R22494 commonsourceibias.n207 commonsourceibias.n206 56.5617
R22495 commonsourceibias.n193 commonsourceibias.n192 56.5617
R22496 commonsourceibias.n687 commonsourceibias.n685 56.5617
R22497 commonsourceibias.n702 commonsourceibias.n700 56.5617
R22498 commonsourceibias.n457 commonsourceibias.n455 56.5617
R22499 commonsourceibias.n472 commonsourceibias.n470 56.5617
R22500 commonsourceibias.n572 commonsourceibias.n570 56.5617
R22501 commonsourceibias.n294 commonsourceibias.n293 56.5617
R22502 commonsourceibias.n308 commonsourceibias.n307 56.5617
R22503 commonsourceibias.n350 commonsourceibias.n349 56.5617
R22504 commonsourceibias.n113 commonsourceibias.n112 56.5617
R22505 commonsourceibias.n99 commonsourceibias.n98 56.5617
R22506 commonsourceibias.n57 commonsourceibias.n56 56.5617
R22507 commonsourceibias.n235 commonsourceibias.n234 56.5617
R22508 commonsourceibias.n221 commonsourceibias.n220 56.5617
R22509 commonsourceibias.n179 commonsourceibias.n178 56.5617
R22510 commonsourceibias.n657 commonsourceibias.n655 56.5617
R22511 commonsourceibias.n672 commonsourceibias.n670 56.5617
R22512 commonsourceibias.n717 commonsourceibias.n715 56.5617
R22513 commonsourceibias.n427 commonsourceibias.n425 56.5617
R22514 commonsourceibias.n442 commonsourceibias.n440 56.5617
R22515 commonsourceibias.n487 commonsourceibias.n485 56.5617
R22516 commonsourceibias.n602 commonsourceibias.n600 56.5617
R22517 commonsourceibias.n587 commonsourceibias.n585 56.5617
R22518 commonsourceibias.n543 commonsourceibias.n541 56.5617
R22519 commonsourceibias.n557 commonsourceibias.n556 56.5617
R22520 commonsourceibias.n285 commonsourceibias.n284 51.2335
R22521 commonsourceibias.n357 commonsourceibias.n252 51.2335
R22522 commonsourceibias.n120 commonsourceibias.n15 51.2335
R22523 commonsourceibias.n48 commonsourceibias.n47 51.2335
R22524 commonsourceibias.n242 commonsourceibias.n1 51.2335
R22525 commonsourceibias.n170 commonsourceibias.n169 51.2335
R22526 commonsourceibias.n647 commonsourceibias.n646 51.2335
R22527 commonsourceibias.n724 commonsourceibias.n619 51.2335
R22528 commonsourceibias.n417 commonsourceibias.n416 51.2335
R22529 commonsourceibias.n494 commonsourceibias.n389 51.2335
R22530 commonsourceibias.n609 commonsourceibias.n368 51.2335
R22531 commonsourceibias.n533 commonsourceibias.n532 51.2335
R22532 commonsourceibias.n364 commonsourceibias.n363 50.9056
R22533 commonsourceibias.n127 commonsourceibias.n126 50.9056
R22534 commonsourceibias.n249 commonsourceibias.n248 50.9056
R22535 commonsourceibias.n731 commonsourceibias.n730 50.9056
R22536 commonsourceibias.n501 commonsourceibias.n500 50.9056
R22537 commonsourceibias.n616 commonsourceibias.n615 50.9056
R22538 commonsourceibias.n299 commonsourceibias.n298 50.2647
R22539 commonsourceibias.n343 commonsourceibias.n257 50.2647
R22540 commonsourceibias.n106 commonsourceibias.n20 50.2647
R22541 commonsourceibias.n62 commonsourceibias.n61 50.2647
R22542 commonsourceibias.n228 commonsourceibias.n6 50.2647
R22543 commonsourceibias.n184 commonsourceibias.n183 50.2647
R22544 commonsourceibias.n662 commonsourceibias.n661 50.2647
R22545 commonsourceibias.n709 commonsourceibias.n623 50.2647
R22546 commonsourceibias.n432 commonsourceibias.n431 50.2647
R22547 commonsourceibias.n479 commonsourceibias.n393 50.2647
R22548 commonsourceibias.n594 commonsourceibias.n372 50.2647
R22549 commonsourceibias.n548 commonsourceibias.n547 50.2647
R22550 commonsourceibias.n281 commonsourceibias.n280 49.9027
R22551 commonsourceibias.n44 commonsourceibias.n43 49.9027
R22552 commonsourceibias.n166 commonsourceibias.n165 49.9027
R22553 commonsourceibias.n643 commonsourceibias.n642 49.9027
R22554 commonsourceibias.n413 commonsourceibias.n412 49.9027
R22555 commonsourceibias.n529 commonsourceibias.n528 49.9027
R22556 commonsourceibias.n313 commonsourceibias.n312 49.296
R22557 commonsourceibias.n329 commonsourceibias.n262 49.296
R22558 commonsourceibias.n92 commonsourceibias.n25 49.296
R22559 commonsourceibias.n76 commonsourceibias.n75 49.296
R22560 commonsourceibias.n214 commonsourceibias.n11 49.296
R22561 commonsourceibias.n198 commonsourceibias.n197 49.296
R22562 commonsourceibias.n677 commonsourceibias.n676 49.296
R22563 commonsourceibias.n694 commonsourceibias.n627 49.296
R22564 commonsourceibias.n447 commonsourceibias.n446 49.296
R22565 commonsourceibias.n464 commonsourceibias.n397 49.296
R22566 commonsourceibias.n579 commonsourceibias.n376 49.296
R22567 commonsourceibias.n562 commonsourceibias.n561 49.296
R22568 commonsourceibias.n315 commonsourceibias.n267 48.3272
R22569 commonsourceibias.n327 commonsourceibias.n326 48.3272
R22570 commonsourceibias.n90 commonsourceibias.n89 48.3272
R22571 commonsourceibias.n78 commonsourceibias.n30 48.3272
R22572 commonsourceibias.n212 commonsourceibias.n211 48.3272
R22573 commonsourceibias.n202 commonsourceibias.n201 48.3272
R22574 commonsourceibias.n679 commonsourceibias.n631 48.3272
R22575 commonsourceibias.n692 commonsourceibias.n691 48.3272
R22576 commonsourceibias.n449 commonsourceibias.n401 48.3272
R22577 commonsourceibias.n462 commonsourceibias.n461 48.3272
R22578 commonsourceibias.n577 commonsourceibias.n576 48.3272
R22579 commonsourceibias.n566 commonsourceibias.n565 48.3272
R22580 commonsourceibias.n301 commonsourceibias.n272 47.3584
R22581 commonsourceibias.n341 commonsourceibias.n340 47.3584
R22582 commonsourceibias.n104 commonsourceibias.n103 47.3584
R22583 commonsourceibias.n64 commonsourceibias.n35 47.3584
R22584 commonsourceibias.n226 commonsourceibias.n225 47.3584
R22585 commonsourceibias.n186 commonsourceibias.n157 47.3584
R22586 commonsourceibias.n664 commonsourceibias.n635 47.3584
R22587 commonsourceibias.n707 commonsourceibias.n706 47.3584
R22588 commonsourceibias.n434 commonsourceibias.n405 47.3584
R22589 commonsourceibias.n477 commonsourceibias.n476 47.3584
R22590 commonsourceibias.n592 commonsourceibias.n591 47.3584
R22591 commonsourceibias.n550 commonsourceibias.n521 47.3584
R22592 commonsourceibias.n287 commonsourceibias.n277 46.3896
R22593 commonsourceibias.n355 commonsourceibias.n354 46.3896
R22594 commonsourceibias.n118 commonsourceibias.n117 46.3896
R22595 commonsourceibias.n50 commonsourceibias.n40 46.3896
R22596 commonsourceibias.n240 commonsourceibias.n239 46.3896
R22597 commonsourceibias.n172 commonsourceibias.n162 46.3896
R22598 commonsourceibias.n649 commonsourceibias.n639 46.3896
R22599 commonsourceibias.n722 commonsourceibias.n721 46.3896
R22600 commonsourceibias.n419 commonsourceibias.n409 46.3896
R22601 commonsourceibias.n492 commonsourceibias.n491 46.3896
R22602 commonsourceibias.n607 commonsourceibias.n606 46.3896
R22603 commonsourceibias.n535 commonsourceibias.n525 46.3896
R22604 commonsourceibias.n282 commonsourceibias.n281 44.7059
R22605 commonsourceibias.n644 commonsourceibias.n643 44.7059
R22606 commonsourceibias.n414 commonsourceibias.n413 44.7059
R22607 commonsourceibias.n530 commonsourceibias.n529 44.7059
R22608 commonsourceibias.n45 commonsourceibias.n44 44.7059
R22609 commonsourceibias.n167 commonsourceibias.n166 44.7059
R22610 commonsourceibias.n291 commonsourceibias.n277 34.7644
R22611 commonsourceibias.n354 commonsourceibias.n254 34.7644
R22612 commonsourceibias.n117 commonsourceibias.n17 34.7644
R22613 commonsourceibias.n54 commonsourceibias.n40 34.7644
R22614 commonsourceibias.n239 commonsourceibias.n3 34.7644
R22615 commonsourceibias.n176 commonsourceibias.n162 34.7644
R22616 commonsourceibias.n653 commonsourceibias.n639 34.7644
R22617 commonsourceibias.n721 commonsourceibias.n621 34.7644
R22618 commonsourceibias.n423 commonsourceibias.n409 34.7644
R22619 commonsourceibias.n491 commonsourceibias.n391 34.7644
R22620 commonsourceibias.n606 commonsourceibias.n370 34.7644
R22621 commonsourceibias.n539 commonsourceibias.n525 34.7644
R22622 commonsourceibias.n305 commonsourceibias.n272 33.7956
R22623 commonsourceibias.n340 commonsourceibias.n259 33.7956
R22624 commonsourceibias.n103 commonsourceibias.n22 33.7956
R22625 commonsourceibias.n68 commonsourceibias.n35 33.7956
R22626 commonsourceibias.n225 commonsourceibias.n8 33.7956
R22627 commonsourceibias.n190 commonsourceibias.n157 33.7956
R22628 commonsourceibias.n668 commonsourceibias.n635 33.7956
R22629 commonsourceibias.n706 commonsourceibias.n625 33.7956
R22630 commonsourceibias.n438 commonsourceibias.n405 33.7956
R22631 commonsourceibias.n476 commonsourceibias.n395 33.7956
R22632 commonsourceibias.n591 commonsourceibias.n374 33.7956
R22633 commonsourceibias.n554 commonsourceibias.n521 33.7956
R22634 commonsourceibias.n319 commonsourceibias.n267 32.8269
R22635 commonsourceibias.n326 commonsourceibias.n264 32.8269
R22636 commonsourceibias.n89 commonsourceibias.n27 32.8269
R22637 commonsourceibias.n82 commonsourceibias.n30 32.8269
R22638 commonsourceibias.n211 commonsourceibias.n13 32.8269
R22639 commonsourceibias.n203 commonsourceibias.n202 32.8269
R22640 commonsourceibias.n683 commonsourceibias.n631 32.8269
R22641 commonsourceibias.n691 commonsourceibias.n629 32.8269
R22642 commonsourceibias.n453 commonsourceibias.n401 32.8269
R22643 commonsourceibias.n461 commonsourceibias.n399 32.8269
R22644 commonsourceibias.n576 commonsourceibias.n378 32.8269
R22645 commonsourceibias.n567 commonsourceibias.n566 32.8269
R22646 commonsourceibias.n312 commonsourceibias.n269 31.8581
R22647 commonsourceibias.n333 commonsourceibias.n262 31.8581
R22648 commonsourceibias.n96 commonsourceibias.n25 31.8581
R22649 commonsourceibias.n75 commonsourceibias.n32 31.8581
R22650 commonsourceibias.n218 commonsourceibias.n11 31.8581
R22651 commonsourceibias.n197 commonsourceibias.n196 31.8581
R22652 commonsourceibias.n676 commonsourceibias.n633 31.8581
R22653 commonsourceibias.n698 commonsourceibias.n627 31.8581
R22654 commonsourceibias.n446 commonsourceibias.n403 31.8581
R22655 commonsourceibias.n468 commonsourceibias.n397 31.8581
R22656 commonsourceibias.n583 commonsourceibias.n376 31.8581
R22657 commonsourceibias.n561 commonsourceibias.n560 31.8581
R22658 commonsourceibias.n298 commonsourceibias.n274 30.8893
R22659 commonsourceibias.n347 commonsourceibias.n257 30.8893
R22660 commonsourceibias.n110 commonsourceibias.n20 30.8893
R22661 commonsourceibias.n61 commonsourceibias.n37 30.8893
R22662 commonsourceibias.n232 commonsourceibias.n6 30.8893
R22663 commonsourceibias.n183 commonsourceibias.n159 30.8893
R22664 commonsourceibias.n661 commonsourceibias.n637 30.8893
R22665 commonsourceibias.n713 commonsourceibias.n623 30.8893
R22666 commonsourceibias.n431 commonsourceibias.n407 30.8893
R22667 commonsourceibias.n483 commonsourceibias.n393 30.8893
R22668 commonsourceibias.n598 commonsourceibias.n372 30.8893
R22669 commonsourceibias.n547 commonsourceibias.n523 30.8893
R22670 commonsourceibias.n284 commonsourceibias.n279 29.9206
R22671 commonsourceibias.n361 commonsourceibias.n252 29.9206
R22672 commonsourceibias.n124 commonsourceibias.n15 29.9206
R22673 commonsourceibias.n47 commonsourceibias.n42 29.9206
R22674 commonsourceibias.n246 commonsourceibias.n1 29.9206
R22675 commonsourceibias.n169 commonsourceibias.n164 29.9206
R22676 commonsourceibias.n646 commonsourceibias.n641 29.9206
R22677 commonsourceibias.n728 commonsourceibias.n619 29.9206
R22678 commonsourceibias.n416 commonsourceibias.n411 29.9206
R22679 commonsourceibias.n498 commonsourceibias.n389 29.9206
R22680 commonsourceibias.n613 commonsourceibias.n368 29.9206
R22681 commonsourceibias.n532 commonsourceibias.n527 29.9206
R22682 commonsourceibias.n363 commonsourceibias.n362 21.8872
R22683 commonsourceibias.n126 commonsourceibias.n125 21.8872
R22684 commonsourceibias.n248 commonsourceibias.n247 21.8872
R22685 commonsourceibias.n730 commonsourceibias.n729 21.8872
R22686 commonsourceibias.n500 commonsourceibias.n499 21.8872
R22687 commonsourceibias.n615 commonsourceibias.n614 21.8872
R22688 commonsourceibias.n294 commonsourceibias.n276 21.3954
R22689 commonsourceibias.n349 commonsourceibias.n348 21.3954
R22690 commonsourceibias.n112 commonsourceibias.n111 21.3954
R22691 commonsourceibias.n57 commonsourceibias.n39 21.3954
R22692 commonsourceibias.n234 commonsourceibias.n233 21.3954
R22693 commonsourceibias.n179 commonsourceibias.n161 21.3954
R22694 commonsourceibias.n657 commonsourceibias.n656 21.3954
R22695 commonsourceibias.n715 commonsourceibias.n714 21.3954
R22696 commonsourceibias.n427 commonsourceibias.n426 21.3954
R22697 commonsourceibias.n485 commonsourceibias.n484 21.3954
R22698 commonsourceibias.n600 commonsourceibias.n599 21.3954
R22699 commonsourceibias.n543 commonsourceibias.n542 21.3954
R22700 commonsourceibias.n308 commonsourceibias.n271 20.9036
R22701 commonsourceibias.n335 commonsourceibias.n334 20.9036
R22702 commonsourceibias.n98 commonsourceibias.n97 20.9036
R22703 commonsourceibias.n71 commonsourceibias.n34 20.9036
R22704 commonsourceibias.n220 commonsourceibias.n219 20.9036
R22705 commonsourceibias.n193 commonsourceibias.n155 20.9036
R22706 commonsourceibias.n672 commonsourceibias.n671 20.9036
R22707 commonsourceibias.n700 commonsourceibias.n699 20.9036
R22708 commonsourceibias.n442 commonsourceibias.n441 20.9036
R22709 commonsourceibias.n470 commonsourceibias.n469 20.9036
R22710 commonsourceibias.n585 commonsourceibias.n584 20.9036
R22711 commonsourceibias.n557 commonsourceibias.n519 20.9036
R22712 commonsourceibias.n321 commonsourceibias.n320 20.4117
R22713 commonsourceibias.n322 commonsourceibias.n266 20.4117
R22714 commonsourceibias.n85 commonsourceibias.n29 20.4117
R22715 commonsourceibias.n84 commonsourceibias.n83 20.4117
R22716 commonsourceibias.n207 commonsourceibias.n150 20.4117
R22717 commonsourceibias.n206 commonsourceibias.n151 20.4117
R22718 commonsourceibias.n685 commonsourceibias.n684 20.4117
R22719 commonsourceibias.n687 commonsourceibias.n686 20.4117
R22720 commonsourceibias.n455 commonsourceibias.n454 20.4117
R22721 commonsourceibias.n457 commonsourceibias.n456 20.4117
R22722 commonsourceibias.n572 commonsourceibias.n571 20.4117
R22723 commonsourceibias.n570 commonsourceibias.n515 20.4117
R22724 commonsourceibias.n307 commonsourceibias.n306 19.9199
R22725 commonsourceibias.n336 commonsourceibias.n261 19.9199
R22726 commonsourceibias.n99 commonsourceibias.n24 19.9199
R22727 commonsourceibias.n70 commonsourceibias.n69 19.9199
R22728 commonsourceibias.n221 commonsourceibias.n10 19.9199
R22729 commonsourceibias.n192 commonsourceibias.n191 19.9199
R22730 commonsourceibias.n670 commonsourceibias.n669 19.9199
R22731 commonsourceibias.n702 commonsourceibias.n701 19.9199
R22732 commonsourceibias.n440 commonsourceibias.n439 19.9199
R22733 commonsourceibias.n472 commonsourceibias.n471 19.9199
R22734 commonsourceibias.n587 commonsourceibias.n586 19.9199
R22735 commonsourceibias.n556 commonsourceibias.n555 19.9199
R22736 commonsourceibias.n293 commonsourceibias.n292 19.4281
R22737 commonsourceibias.n350 commonsourceibias.n256 19.4281
R22738 commonsourceibias.n113 commonsourceibias.n19 19.4281
R22739 commonsourceibias.n56 commonsourceibias.n55 19.4281
R22740 commonsourceibias.n235 commonsourceibias.n5 19.4281
R22741 commonsourceibias.n178 commonsourceibias.n177 19.4281
R22742 commonsourceibias.n655 commonsourceibias.n654 19.4281
R22743 commonsourceibias.n717 commonsourceibias.n716 19.4281
R22744 commonsourceibias.n425 commonsourceibias.n424 19.4281
R22745 commonsourceibias.n487 commonsourceibias.n486 19.4281
R22746 commonsourceibias.n602 commonsourceibias.n601 19.4281
R22747 commonsourceibias.n541 commonsourceibias.n540 19.4281
R22748 commonsourceibias.n286 commonsourceibias.n285 13.526
R22749 commonsourceibias.n357 commonsourceibias.n356 13.526
R22750 commonsourceibias.n120 commonsourceibias.n119 13.526
R22751 commonsourceibias.n49 commonsourceibias.n48 13.526
R22752 commonsourceibias.n242 commonsourceibias.n241 13.526
R22753 commonsourceibias.n171 commonsourceibias.n170 13.526
R22754 commonsourceibias.n648 commonsourceibias.n647 13.526
R22755 commonsourceibias.n724 commonsourceibias.n723 13.526
R22756 commonsourceibias.n418 commonsourceibias.n417 13.526
R22757 commonsourceibias.n494 commonsourceibias.n493 13.526
R22758 commonsourceibias.n609 commonsourceibias.n608 13.526
R22759 commonsourceibias.n534 commonsourceibias.n533 13.526
R22760 commonsourceibias.n130 commonsourceibias.n128 13.2322
R22761 commonsourceibias.n504 commonsourceibias.n502 13.2322
R22762 commonsourceibias.n300 commonsourceibias.n299 13.0342
R22763 commonsourceibias.n343 commonsourceibias.n342 13.0342
R22764 commonsourceibias.n106 commonsourceibias.n105 13.0342
R22765 commonsourceibias.n63 commonsourceibias.n62 13.0342
R22766 commonsourceibias.n228 commonsourceibias.n227 13.0342
R22767 commonsourceibias.n185 commonsourceibias.n184 13.0342
R22768 commonsourceibias.n663 commonsourceibias.n662 13.0342
R22769 commonsourceibias.n709 commonsourceibias.n708 13.0342
R22770 commonsourceibias.n433 commonsourceibias.n432 13.0342
R22771 commonsourceibias.n479 commonsourceibias.n478 13.0342
R22772 commonsourceibias.n594 commonsourceibias.n593 13.0342
R22773 commonsourceibias.n549 commonsourceibias.n548 13.0342
R22774 commonsourceibias.n314 commonsourceibias.n313 12.5423
R22775 commonsourceibias.n329 commonsourceibias.n328 12.5423
R22776 commonsourceibias.n92 commonsourceibias.n91 12.5423
R22777 commonsourceibias.n77 commonsourceibias.n76 12.5423
R22778 commonsourceibias.n214 commonsourceibias.n213 12.5423
R22779 commonsourceibias.n198 commonsourceibias.n153 12.5423
R22780 commonsourceibias.n678 commonsourceibias.n677 12.5423
R22781 commonsourceibias.n694 commonsourceibias.n693 12.5423
R22782 commonsourceibias.n448 commonsourceibias.n447 12.5423
R22783 commonsourceibias.n464 commonsourceibias.n463 12.5423
R22784 commonsourceibias.n579 commonsourceibias.n578 12.5423
R22785 commonsourceibias.n562 commonsourceibias.n517 12.5423
R22786 commonsourceibias.n734 commonsourceibias.n366 12.2777
R22787 commonsourceibias.n315 commonsourceibias.n314 12.0505
R22788 commonsourceibias.n328 commonsourceibias.n327 12.0505
R22789 commonsourceibias.n91 commonsourceibias.n90 12.0505
R22790 commonsourceibias.n78 commonsourceibias.n77 12.0505
R22791 commonsourceibias.n213 commonsourceibias.n212 12.0505
R22792 commonsourceibias.n201 commonsourceibias.n153 12.0505
R22793 commonsourceibias.n679 commonsourceibias.n678 12.0505
R22794 commonsourceibias.n693 commonsourceibias.n692 12.0505
R22795 commonsourceibias.n449 commonsourceibias.n448 12.0505
R22796 commonsourceibias.n463 commonsourceibias.n462 12.0505
R22797 commonsourceibias.n578 commonsourceibias.n577 12.0505
R22798 commonsourceibias.n565 commonsourceibias.n517 12.0505
R22799 commonsourceibias.n301 commonsourceibias.n300 11.5587
R22800 commonsourceibias.n342 commonsourceibias.n341 11.5587
R22801 commonsourceibias.n105 commonsourceibias.n104 11.5587
R22802 commonsourceibias.n64 commonsourceibias.n63 11.5587
R22803 commonsourceibias.n227 commonsourceibias.n226 11.5587
R22804 commonsourceibias.n186 commonsourceibias.n185 11.5587
R22805 commonsourceibias.n664 commonsourceibias.n663 11.5587
R22806 commonsourceibias.n708 commonsourceibias.n707 11.5587
R22807 commonsourceibias.n434 commonsourceibias.n433 11.5587
R22808 commonsourceibias.n478 commonsourceibias.n477 11.5587
R22809 commonsourceibias.n593 commonsourceibias.n592 11.5587
R22810 commonsourceibias.n550 commonsourceibias.n549 11.5587
R22811 commonsourceibias.n287 commonsourceibias.n286 11.0668
R22812 commonsourceibias.n356 commonsourceibias.n355 11.0668
R22813 commonsourceibias.n119 commonsourceibias.n118 11.0668
R22814 commonsourceibias.n50 commonsourceibias.n49 11.0668
R22815 commonsourceibias.n241 commonsourceibias.n240 11.0668
R22816 commonsourceibias.n172 commonsourceibias.n171 11.0668
R22817 commonsourceibias.n649 commonsourceibias.n648 11.0668
R22818 commonsourceibias.n723 commonsourceibias.n722 11.0668
R22819 commonsourceibias.n419 commonsourceibias.n418 11.0668
R22820 commonsourceibias.n493 commonsourceibias.n492 11.0668
R22821 commonsourceibias.n608 commonsourceibias.n607 11.0668
R22822 commonsourceibias.n535 commonsourceibias.n534 11.0668
R22823 commonsourceibias.n734 commonsourceibias.n733 10.3347
R22824 commonsourceibias.n149 commonsourceibias.n148 9.50363
R22825 commonsourceibias.n514 commonsourceibias.n513 9.50363
R22826 commonsourceibias.n366 commonsourceibias.n250 8.75852
R22827 commonsourceibias.n733 commonsourceibias.n617 8.75852
R22828 commonsourceibias.n292 commonsourceibias.n291 5.16479
R22829 commonsourceibias.n256 commonsourceibias.n254 5.16479
R22830 commonsourceibias.n19 commonsourceibias.n17 5.16479
R22831 commonsourceibias.n55 commonsourceibias.n54 5.16479
R22832 commonsourceibias.n5 commonsourceibias.n3 5.16479
R22833 commonsourceibias.n177 commonsourceibias.n176 5.16479
R22834 commonsourceibias.n654 commonsourceibias.n653 5.16479
R22835 commonsourceibias.n716 commonsourceibias.n621 5.16479
R22836 commonsourceibias.n424 commonsourceibias.n423 5.16479
R22837 commonsourceibias.n486 commonsourceibias.n391 5.16479
R22838 commonsourceibias.n601 commonsourceibias.n370 5.16479
R22839 commonsourceibias.n540 commonsourceibias.n539 5.16479
R22840 commonsourceibias.n366 commonsourceibias.n365 5.03125
R22841 commonsourceibias.n733 commonsourceibias.n732 5.03125
R22842 commonsourceibias.n306 commonsourceibias.n305 4.67295
R22843 commonsourceibias.n261 commonsourceibias.n259 4.67295
R22844 commonsourceibias.n24 commonsourceibias.n22 4.67295
R22845 commonsourceibias.n69 commonsourceibias.n68 4.67295
R22846 commonsourceibias.n10 commonsourceibias.n8 4.67295
R22847 commonsourceibias.n191 commonsourceibias.n190 4.67295
R22848 commonsourceibias.n669 commonsourceibias.n668 4.67295
R22849 commonsourceibias.n701 commonsourceibias.n625 4.67295
R22850 commonsourceibias.n439 commonsourceibias.n438 4.67295
R22851 commonsourceibias.n471 commonsourceibias.n395 4.67295
R22852 commonsourceibias.n586 commonsourceibias.n374 4.67295
R22853 commonsourceibias.n555 commonsourceibias.n554 4.67295
R22854 commonsourceibias commonsourceibias.n734 4.20978
R22855 commonsourceibias.n320 commonsourceibias.n319 4.18111
R22856 commonsourceibias.n266 commonsourceibias.n264 4.18111
R22857 commonsourceibias.n29 commonsourceibias.n27 4.18111
R22858 commonsourceibias.n83 commonsourceibias.n82 4.18111
R22859 commonsourceibias.n150 commonsourceibias.n13 4.18111
R22860 commonsourceibias.n203 commonsourceibias.n151 4.18111
R22861 commonsourceibias.n684 commonsourceibias.n683 4.18111
R22862 commonsourceibias.n686 commonsourceibias.n629 4.18111
R22863 commonsourceibias.n454 commonsourceibias.n453 4.18111
R22864 commonsourceibias.n456 commonsourceibias.n399 4.18111
R22865 commonsourceibias.n571 commonsourceibias.n378 4.18111
R22866 commonsourceibias.n567 commonsourceibias.n515 4.18111
R22867 commonsourceibias.n271 commonsourceibias.n269 3.68928
R22868 commonsourceibias.n334 commonsourceibias.n333 3.68928
R22869 commonsourceibias.n97 commonsourceibias.n96 3.68928
R22870 commonsourceibias.n34 commonsourceibias.n32 3.68928
R22871 commonsourceibias.n219 commonsourceibias.n218 3.68928
R22872 commonsourceibias.n196 commonsourceibias.n155 3.68928
R22873 commonsourceibias.n671 commonsourceibias.n633 3.68928
R22874 commonsourceibias.n699 commonsourceibias.n698 3.68928
R22875 commonsourceibias.n441 commonsourceibias.n403 3.68928
R22876 commonsourceibias.n469 commonsourceibias.n468 3.68928
R22877 commonsourceibias.n584 commonsourceibias.n583 3.68928
R22878 commonsourceibias.n560 commonsourceibias.n519 3.68928
R22879 commonsourceibias.n276 commonsourceibias.n274 3.19744
R22880 commonsourceibias.n348 commonsourceibias.n347 3.19744
R22881 commonsourceibias.n111 commonsourceibias.n110 3.19744
R22882 commonsourceibias.n39 commonsourceibias.n37 3.19744
R22883 commonsourceibias.n233 commonsourceibias.n232 3.19744
R22884 commonsourceibias.n161 commonsourceibias.n159 3.19744
R22885 commonsourceibias.n656 commonsourceibias.n637 3.19744
R22886 commonsourceibias.n714 commonsourceibias.n713 3.19744
R22887 commonsourceibias.n426 commonsourceibias.n407 3.19744
R22888 commonsourceibias.n484 commonsourceibias.n483 3.19744
R22889 commonsourceibias.n599 commonsourceibias.n598 3.19744
R22890 commonsourceibias.n542 commonsourceibias.n523 3.19744
R22891 commonsourceibias.n139 commonsourceibias.t47 2.82907
R22892 commonsourceibias.n139 commonsourceibias.t79 2.82907
R22893 commonsourceibias.n140 commonsourceibias.t55 2.82907
R22894 commonsourceibias.n140 commonsourceibias.t5 2.82907
R22895 commonsourceibias.n142 commonsourceibias.t19 2.82907
R22896 commonsourceibias.n142 commonsourceibias.t23 2.82907
R22897 commonsourceibias.n144 commonsourceibias.t39 2.82907
R22898 commonsourceibias.n144 commonsourceibias.t71 2.82907
R22899 commonsourceibias.n146 commonsourceibias.t57 2.82907
R22900 commonsourceibias.n146 commonsourceibias.t27 2.82907
R22901 commonsourceibias.n137 commonsourceibias.t11 2.82907
R22902 commonsourceibias.n137 commonsourceibias.t41 2.82907
R22903 commonsourceibias.n135 commonsourceibias.t25 2.82907
R22904 commonsourceibias.n135 commonsourceibias.t35 2.82907
R22905 commonsourceibias.n133 commonsourceibias.t37 2.82907
R22906 commonsourceibias.n133 commonsourceibias.t77 2.82907
R22907 commonsourceibias.n131 commonsourceibias.t51 2.82907
R22908 commonsourceibias.n131 commonsourceibias.t9 2.82907
R22909 commonsourceibias.n129 commonsourceibias.t75 2.82907
R22910 commonsourceibias.n129 commonsourceibias.t21 2.82907
R22911 commonsourceibias.n503 commonsourceibias.t43 2.82907
R22912 commonsourceibias.n503 commonsourceibias.t15 2.82907
R22913 commonsourceibias.n505 commonsourceibias.t31 2.82907
R22914 commonsourceibias.n505 commonsourceibias.t1 2.82907
R22915 commonsourceibias.n507 commonsourceibias.t17 2.82907
R22916 commonsourceibias.n507 commonsourceibias.t61 2.82907
R22917 commonsourceibias.n509 commonsourceibias.t59 2.82907
R22918 commonsourceibias.n509 commonsourceibias.t45 2.82907
R22919 commonsourceibias.n511 commonsourceibias.t65 2.82907
R22920 commonsourceibias.n511 commonsourceibias.t33 2.82907
R22921 commonsourceibias.n386 commonsourceibias.t53 2.82907
R22922 commonsourceibias.n386 commonsourceibias.t73 2.82907
R22923 commonsourceibias.n384 commonsourceibias.t7 2.82907
R22924 commonsourceibias.n384 commonsourceibias.t63 2.82907
R22925 commonsourceibias.n382 commonsourceibias.t69 2.82907
R22926 commonsourceibias.n382 commonsourceibias.t67 2.82907
R22927 commonsourceibias.n380 commonsourceibias.t49 2.82907
R22928 commonsourceibias.n380 commonsourceibias.t13 2.82907
R22929 commonsourceibias.n379 commonsourceibias.t29 2.82907
R22930 commonsourceibias.n379 commonsourceibias.t3 2.82907
R22931 commonsourceibias.n280 commonsourceibias.n279 2.7056
R22932 commonsourceibias.n362 commonsourceibias.n361 2.7056
R22933 commonsourceibias.n125 commonsourceibias.n124 2.7056
R22934 commonsourceibias.n43 commonsourceibias.n42 2.7056
R22935 commonsourceibias.n247 commonsourceibias.n246 2.7056
R22936 commonsourceibias.n165 commonsourceibias.n164 2.7056
R22937 commonsourceibias.n642 commonsourceibias.n641 2.7056
R22938 commonsourceibias.n729 commonsourceibias.n728 2.7056
R22939 commonsourceibias.n412 commonsourceibias.n411 2.7056
R22940 commonsourceibias.n499 commonsourceibias.n498 2.7056
R22941 commonsourceibias.n614 commonsourceibias.n613 2.7056
R22942 commonsourceibias.n528 commonsourceibias.n527 2.7056
R22943 commonsourceibias.n132 commonsourceibias.n130 0.573776
R22944 commonsourceibias.n134 commonsourceibias.n132 0.573776
R22945 commonsourceibias.n136 commonsourceibias.n134 0.573776
R22946 commonsourceibias.n138 commonsourceibias.n136 0.573776
R22947 commonsourceibias.n147 commonsourceibias.n145 0.573776
R22948 commonsourceibias.n145 commonsourceibias.n143 0.573776
R22949 commonsourceibias.n143 commonsourceibias.n141 0.573776
R22950 commonsourceibias.n383 commonsourceibias.n381 0.573776
R22951 commonsourceibias.n385 commonsourceibias.n383 0.573776
R22952 commonsourceibias.n387 commonsourceibias.n385 0.573776
R22953 commonsourceibias.n512 commonsourceibias.n510 0.573776
R22954 commonsourceibias.n510 commonsourceibias.n508 0.573776
R22955 commonsourceibias.n508 commonsourceibias.n506 0.573776
R22956 commonsourceibias.n506 commonsourceibias.n504 0.573776
R22957 commonsourceibias.n148 commonsourceibias.n138 0.287138
R22958 commonsourceibias.n148 commonsourceibias.n147 0.287138
R22959 commonsourceibias.n513 commonsourceibias.n387 0.287138
R22960 commonsourceibias.n513 commonsourceibias.n512 0.287138
R22961 commonsourceibias.n365 commonsourceibias.n251 0.285035
R22962 commonsourceibias.n128 commonsourceibias.n14 0.285035
R22963 commonsourceibias.n250 commonsourceibias.n0 0.285035
R22964 commonsourceibias.n732 commonsourceibias.n618 0.285035
R22965 commonsourceibias.n502 commonsourceibias.n388 0.285035
R22966 commonsourceibias.n617 commonsourceibias.n367 0.285035
R22967 commonsourceibias.n360 commonsourceibias.n251 0.189894
R22968 commonsourceibias.n360 commonsourceibias.n359 0.189894
R22969 commonsourceibias.n359 commonsourceibias.n358 0.189894
R22970 commonsourceibias.n358 commonsourceibias.n253 0.189894
R22971 commonsourceibias.n353 commonsourceibias.n253 0.189894
R22972 commonsourceibias.n353 commonsourceibias.n352 0.189894
R22973 commonsourceibias.n352 commonsourceibias.n351 0.189894
R22974 commonsourceibias.n351 commonsourceibias.n255 0.189894
R22975 commonsourceibias.n346 commonsourceibias.n255 0.189894
R22976 commonsourceibias.n346 commonsourceibias.n345 0.189894
R22977 commonsourceibias.n345 commonsourceibias.n344 0.189894
R22978 commonsourceibias.n344 commonsourceibias.n258 0.189894
R22979 commonsourceibias.n339 commonsourceibias.n258 0.189894
R22980 commonsourceibias.n339 commonsourceibias.n338 0.189894
R22981 commonsourceibias.n338 commonsourceibias.n337 0.189894
R22982 commonsourceibias.n337 commonsourceibias.n260 0.189894
R22983 commonsourceibias.n332 commonsourceibias.n260 0.189894
R22984 commonsourceibias.n332 commonsourceibias.n331 0.189894
R22985 commonsourceibias.n331 commonsourceibias.n330 0.189894
R22986 commonsourceibias.n330 commonsourceibias.n263 0.189894
R22987 commonsourceibias.n325 commonsourceibias.n263 0.189894
R22988 commonsourceibias.n325 commonsourceibias.n324 0.189894
R22989 commonsourceibias.n324 commonsourceibias.n323 0.189894
R22990 commonsourceibias.n323 commonsourceibias.n265 0.189894
R22991 commonsourceibias.n318 commonsourceibias.n265 0.189894
R22992 commonsourceibias.n318 commonsourceibias.n317 0.189894
R22993 commonsourceibias.n317 commonsourceibias.n316 0.189894
R22994 commonsourceibias.n316 commonsourceibias.n268 0.189894
R22995 commonsourceibias.n311 commonsourceibias.n268 0.189894
R22996 commonsourceibias.n311 commonsourceibias.n310 0.189894
R22997 commonsourceibias.n310 commonsourceibias.n309 0.189894
R22998 commonsourceibias.n309 commonsourceibias.n270 0.189894
R22999 commonsourceibias.n304 commonsourceibias.n270 0.189894
R23000 commonsourceibias.n304 commonsourceibias.n303 0.189894
R23001 commonsourceibias.n303 commonsourceibias.n302 0.189894
R23002 commonsourceibias.n302 commonsourceibias.n273 0.189894
R23003 commonsourceibias.n297 commonsourceibias.n273 0.189894
R23004 commonsourceibias.n297 commonsourceibias.n296 0.189894
R23005 commonsourceibias.n296 commonsourceibias.n295 0.189894
R23006 commonsourceibias.n295 commonsourceibias.n275 0.189894
R23007 commonsourceibias.n290 commonsourceibias.n275 0.189894
R23008 commonsourceibias.n290 commonsourceibias.n289 0.189894
R23009 commonsourceibias.n289 commonsourceibias.n288 0.189894
R23010 commonsourceibias.n288 commonsourceibias.n278 0.189894
R23011 commonsourceibias.n283 commonsourceibias.n278 0.189894
R23012 commonsourceibias.n283 commonsourceibias.n282 0.189894
R23013 commonsourceibias.n123 commonsourceibias.n14 0.189894
R23014 commonsourceibias.n123 commonsourceibias.n122 0.189894
R23015 commonsourceibias.n122 commonsourceibias.n121 0.189894
R23016 commonsourceibias.n121 commonsourceibias.n16 0.189894
R23017 commonsourceibias.n116 commonsourceibias.n16 0.189894
R23018 commonsourceibias.n116 commonsourceibias.n115 0.189894
R23019 commonsourceibias.n115 commonsourceibias.n114 0.189894
R23020 commonsourceibias.n114 commonsourceibias.n18 0.189894
R23021 commonsourceibias.n109 commonsourceibias.n18 0.189894
R23022 commonsourceibias.n109 commonsourceibias.n108 0.189894
R23023 commonsourceibias.n108 commonsourceibias.n107 0.189894
R23024 commonsourceibias.n107 commonsourceibias.n21 0.189894
R23025 commonsourceibias.n102 commonsourceibias.n21 0.189894
R23026 commonsourceibias.n102 commonsourceibias.n101 0.189894
R23027 commonsourceibias.n101 commonsourceibias.n100 0.189894
R23028 commonsourceibias.n100 commonsourceibias.n23 0.189894
R23029 commonsourceibias.n95 commonsourceibias.n23 0.189894
R23030 commonsourceibias.n95 commonsourceibias.n94 0.189894
R23031 commonsourceibias.n94 commonsourceibias.n93 0.189894
R23032 commonsourceibias.n93 commonsourceibias.n26 0.189894
R23033 commonsourceibias.n88 commonsourceibias.n26 0.189894
R23034 commonsourceibias.n88 commonsourceibias.n87 0.189894
R23035 commonsourceibias.n87 commonsourceibias.n86 0.189894
R23036 commonsourceibias.n86 commonsourceibias.n28 0.189894
R23037 commonsourceibias.n81 commonsourceibias.n28 0.189894
R23038 commonsourceibias.n81 commonsourceibias.n80 0.189894
R23039 commonsourceibias.n80 commonsourceibias.n79 0.189894
R23040 commonsourceibias.n79 commonsourceibias.n31 0.189894
R23041 commonsourceibias.n74 commonsourceibias.n31 0.189894
R23042 commonsourceibias.n74 commonsourceibias.n73 0.189894
R23043 commonsourceibias.n73 commonsourceibias.n72 0.189894
R23044 commonsourceibias.n72 commonsourceibias.n33 0.189894
R23045 commonsourceibias.n67 commonsourceibias.n33 0.189894
R23046 commonsourceibias.n67 commonsourceibias.n66 0.189894
R23047 commonsourceibias.n66 commonsourceibias.n65 0.189894
R23048 commonsourceibias.n65 commonsourceibias.n36 0.189894
R23049 commonsourceibias.n60 commonsourceibias.n36 0.189894
R23050 commonsourceibias.n60 commonsourceibias.n59 0.189894
R23051 commonsourceibias.n59 commonsourceibias.n58 0.189894
R23052 commonsourceibias.n58 commonsourceibias.n38 0.189894
R23053 commonsourceibias.n53 commonsourceibias.n38 0.189894
R23054 commonsourceibias.n53 commonsourceibias.n52 0.189894
R23055 commonsourceibias.n52 commonsourceibias.n51 0.189894
R23056 commonsourceibias.n51 commonsourceibias.n41 0.189894
R23057 commonsourceibias.n46 commonsourceibias.n41 0.189894
R23058 commonsourceibias.n46 commonsourceibias.n45 0.189894
R23059 commonsourceibias.n205 commonsourceibias.n204 0.189894
R23060 commonsourceibias.n204 commonsourceibias.n152 0.189894
R23061 commonsourceibias.n200 commonsourceibias.n152 0.189894
R23062 commonsourceibias.n200 commonsourceibias.n199 0.189894
R23063 commonsourceibias.n199 commonsourceibias.n154 0.189894
R23064 commonsourceibias.n195 commonsourceibias.n154 0.189894
R23065 commonsourceibias.n195 commonsourceibias.n194 0.189894
R23066 commonsourceibias.n194 commonsourceibias.n156 0.189894
R23067 commonsourceibias.n189 commonsourceibias.n156 0.189894
R23068 commonsourceibias.n189 commonsourceibias.n188 0.189894
R23069 commonsourceibias.n188 commonsourceibias.n187 0.189894
R23070 commonsourceibias.n187 commonsourceibias.n158 0.189894
R23071 commonsourceibias.n182 commonsourceibias.n158 0.189894
R23072 commonsourceibias.n182 commonsourceibias.n181 0.189894
R23073 commonsourceibias.n181 commonsourceibias.n180 0.189894
R23074 commonsourceibias.n180 commonsourceibias.n160 0.189894
R23075 commonsourceibias.n175 commonsourceibias.n160 0.189894
R23076 commonsourceibias.n175 commonsourceibias.n174 0.189894
R23077 commonsourceibias.n174 commonsourceibias.n173 0.189894
R23078 commonsourceibias.n173 commonsourceibias.n163 0.189894
R23079 commonsourceibias.n168 commonsourceibias.n163 0.189894
R23080 commonsourceibias.n168 commonsourceibias.n167 0.189894
R23081 commonsourceibias.n245 commonsourceibias.n0 0.189894
R23082 commonsourceibias.n245 commonsourceibias.n244 0.189894
R23083 commonsourceibias.n244 commonsourceibias.n243 0.189894
R23084 commonsourceibias.n243 commonsourceibias.n2 0.189894
R23085 commonsourceibias.n238 commonsourceibias.n2 0.189894
R23086 commonsourceibias.n238 commonsourceibias.n237 0.189894
R23087 commonsourceibias.n237 commonsourceibias.n236 0.189894
R23088 commonsourceibias.n236 commonsourceibias.n4 0.189894
R23089 commonsourceibias.n231 commonsourceibias.n4 0.189894
R23090 commonsourceibias.n231 commonsourceibias.n230 0.189894
R23091 commonsourceibias.n230 commonsourceibias.n229 0.189894
R23092 commonsourceibias.n229 commonsourceibias.n7 0.189894
R23093 commonsourceibias.n224 commonsourceibias.n7 0.189894
R23094 commonsourceibias.n224 commonsourceibias.n223 0.189894
R23095 commonsourceibias.n223 commonsourceibias.n222 0.189894
R23096 commonsourceibias.n222 commonsourceibias.n9 0.189894
R23097 commonsourceibias.n217 commonsourceibias.n9 0.189894
R23098 commonsourceibias.n217 commonsourceibias.n216 0.189894
R23099 commonsourceibias.n216 commonsourceibias.n215 0.189894
R23100 commonsourceibias.n215 commonsourceibias.n12 0.189894
R23101 commonsourceibias.n210 commonsourceibias.n12 0.189894
R23102 commonsourceibias.n210 commonsourceibias.n209 0.189894
R23103 commonsourceibias.n209 commonsourceibias.n208 0.189894
R23104 commonsourceibias.n645 commonsourceibias.n644 0.189894
R23105 commonsourceibias.n645 commonsourceibias.n640 0.189894
R23106 commonsourceibias.n650 commonsourceibias.n640 0.189894
R23107 commonsourceibias.n651 commonsourceibias.n650 0.189894
R23108 commonsourceibias.n652 commonsourceibias.n651 0.189894
R23109 commonsourceibias.n652 commonsourceibias.n638 0.189894
R23110 commonsourceibias.n658 commonsourceibias.n638 0.189894
R23111 commonsourceibias.n659 commonsourceibias.n658 0.189894
R23112 commonsourceibias.n660 commonsourceibias.n659 0.189894
R23113 commonsourceibias.n660 commonsourceibias.n636 0.189894
R23114 commonsourceibias.n665 commonsourceibias.n636 0.189894
R23115 commonsourceibias.n666 commonsourceibias.n665 0.189894
R23116 commonsourceibias.n667 commonsourceibias.n666 0.189894
R23117 commonsourceibias.n667 commonsourceibias.n634 0.189894
R23118 commonsourceibias.n673 commonsourceibias.n634 0.189894
R23119 commonsourceibias.n674 commonsourceibias.n673 0.189894
R23120 commonsourceibias.n675 commonsourceibias.n674 0.189894
R23121 commonsourceibias.n675 commonsourceibias.n632 0.189894
R23122 commonsourceibias.n680 commonsourceibias.n632 0.189894
R23123 commonsourceibias.n681 commonsourceibias.n680 0.189894
R23124 commonsourceibias.n682 commonsourceibias.n681 0.189894
R23125 commonsourceibias.n682 commonsourceibias.n630 0.189894
R23126 commonsourceibias.n688 commonsourceibias.n630 0.189894
R23127 commonsourceibias.n689 commonsourceibias.n688 0.189894
R23128 commonsourceibias.n690 commonsourceibias.n689 0.189894
R23129 commonsourceibias.n690 commonsourceibias.n628 0.189894
R23130 commonsourceibias.n695 commonsourceibias.n628 0.189894
R23131 commonsourceibias.n696 commonsourceibias.n695 0.189894
R23132 commonsourceibias.n697 commonsourceibias.n696 0.189894
R23133 commonsourceibias.n697 commonsourceibias.n626 0.189894
R23134 commonsourceibias.n703 commonsourceibias.n626 0.189894
R23135 commonsourceibias.n704 commonsourceibias.n703 0.189894
R23136 commonsourceibias.n705 commonsourceibias.n704 0.189894
R23137 commonsourceibias.n705 commonsourceibias.n624 0.189894
R23138 commonsourceibias.n710 commonsourceibias.n624 0.189894
R23139 commonsourceibias.n711 commonsourceibias.n710 0.189894
R23140 commonsourceibias.n712 commonsourceibias.n711 0.189894
R23141 commonsourceibias.n712 commonsourceibias.n622 0.189894
R23142 commonsourceibias.n718 commonsourceibias.n622 0.189894
R23143 commonsourceibias.n719 commonsourceibias.n718 0.189894
R23144 commonsourceibias.n720 commonsourceibias.n719 0.189894
R23145 commonsourceibias.n720 commonsourceibias.n620 0.189894
R23146 commonsourceibias.n725 commonsourceibias.n620 0.189894
R23147 commonsourceibias.n726 commonsourceibias.n725 0.189894
R23148 commonsourceibias.n727 commonsourceibias.n726 0.189894
R23149 commonsourceibias.n727 commonsourceibias.n618 0.189894
R23150 commonsourceibias.n415 commonsourceibias.n414 0.189894
R23151 commonsourceibias.n415 commonsourceibias.n410 0.189894
R23152 commonsourceibias.n420 commonsourceibias.n410 0.189894
R23153 commonsourceibias.n421 commonsourceibias.n420 0.189894
R23154 commonsourceibias.n422 commonsourceibias.n421 0.189894
R23155 commonsourceibias.n422 commonsourceibias.n408 0.189894
R23156 commonsourceibias.n428 commonsourceibias.n408 0.189894
R23157 commonsourceibias.n429 commonsourceibias.n428 0.189894
R23158 commonsourceibias.n430 commonsourceibias.n429 0.189894
R23159 commonsourceibias.n430 commonsourceibias.n406 0.189894
R23160 commonsourceibias.n435 commonsourceibias.n406 0.189894
R23161 commonsourceibias.n436 commonsourceibias.n435 0.189894
R23162 commonsourceibias.n437 commonsourceibias.n436 0.189894
R23163 commonsourceibias.n437 commonsourceibias.n404 0.189894
R23164 commonsourceibias.n443 commonsourceibias.n404 0.189894
R23165 commonsourceibias.n444 commonsourceibias.n443 0.189894
R23166 commonsourceibias.n445 commonsourceibias.n444 0.189894
R23167 commonsourceibias.n445 commonsourceibias.n402 0.189894
R23168 commonsourceibias.n450 commonsourceibias.n402 0.189894
R23169 commonsourceibias.n451 commonsourceibias.n450 0.189894
R23170 commonsourceibias.n452 commonsourceibias.n451 0.189894
R23171 commonsourceibias.n452 commonsourceibias.n400 0.189894
R23172 commonsourceibias.n458 commonsourceibias.n400 0.189894
R23173 commonsourceibias.n459 commonsourceibias.n458 0.189894
R23174 commonsourceibias.n460 commonsourceibias.n459 0.189894
R23175 commonsourceibias.n460 commonsourceibias.n398 0.189894
R23176 commonsourceibias.n465 commonsourceibias.n398 0.189894
R23177 commonsourceibias.n466 commonsourceibias.n465 0.189894
R23178 commonsourceibias.n467 commonsourceibias.n466 0.189894
R23179 commonsourceibias.n467 commonsourceibias.n396 0.189894
R23180 commonsourceibias.n473 commonsourceibias.n396 0.189894
R23181 commonsourceibias.n474 commonsourceibias.n473 0.189894
R23182 commonsourceibias.n475 commonsourceibias.n474 0.189894
R23183 commonsourceibias.n475 commonsourceibias.n394 0.189894
R23184 commonsourceibias.n480 commonsourceibias.n394 0.189894
R23185 commonsourceibias.n481 commonsourceibias.n480 0.189894
R23186 commonsourceibias.n482 commonsourceibias.n481 0.189894
R23187 commonsourceibias.n482 commonsourceibias.n392 0.189894
R23188 commonsourceibias.n488 commonsourceibias.n392 0.189894
R23189 commonsourceibias.n489 commonsourceibias.n488 0.189894
R23190 commonsourceibias.n490 commonsourceibias.n489 0.189894
R23191 commonsourceibias.n490 commonsourceibias.n390 0.189894
R23192 commonsourceibias.n495 commonsourceibias.n390 0.189894
R23193 commonsourceibias.n496 commonsourceibias.n495 0.189894
R23194 commonsourceibias.n497 commonsourceibias.n496 0.189894
R23195 commonsourceibias.n497 commonsourceibias.n388 0.189894
R23196 commonsourceibias.n531 commonsourceibias.n530 0.189894
R23197 commonsourceibias.n531 commonsourceibias.n526 0.189894
R23198 commonsourceibias.n536 commonsourceibias.n526 0.189894
R23199 commonsourceibias.n537 commonsourceibias.n536 0.189894
R23200 commonsourceibias.n538 commonsourceibias.n537 0.189894
R23201 commonsourceibias.n538 commonsourceibias.n524 0.189894
R23202 commonsourceibias.n544 commonsourceibias.n524 0.189894
R23203 commonsourceibias.n545 commonsourceibias.n544 0.189894
R23204 commonsourceibias.n546 commonsourceibias.n545 0.189894
R23205 commonsourceibias.n546 commonsourceibias.n522 0.189894
R23206 commonsourceibias.n551 commonsourceibias.n522 0.189894
R23207 commonsourceibias.n552 commonsourceibias.n551 0.189894
R23208 commonsourceibias.n553 commonsourceibias.n552 0.189894
R23209 commonsourceibias.n553 commonsourceibias.n520 0.189894
R23210 commonsourceibias.n558 commonsourceibias.n520 0.189894
R23211 commonsourceibias.n559 commonsourceibias.n558 0.189894
R23212 commonsourceibias.n559 commonsourceibias.n518 0.189894
R23213 commonsourceibias.n563 commonsourceibias.n518 0.189894
R23214 commonsourceibias.n564 commonsourceibias.n563 0.189894
R23215 commonsourceibias.n564 commonsourceibias.n516 0.189894
R23216 commonsourceibias.n568 commonsourceibias.n516 0.189894
R23217 commonsourceibias.n569 commonsourceibias.n568 0.189894
R23218 commonsourceibias.n574 commonsourceibias.n573 0.189894
R23219 commonsourceibias.n575 commonsourceibias.n574 0.189894
R23220 commonsourceibias.n575 commonsourceibias.n377 0.189894
R23221 commonsourceibias.n580 commonsourceibias.n377 0.189894
R23222 commonsourceibias.n581 commonsourceibias.n580 0.189894
R23223 commonsourceibias.n582 commonsourceibias.n581 0.189894
R23224 commonsourceibias.n582 commonsourceibias.n375 0.189894
R23225 commonsourceibias.n588 commonsourceibias.n375 0.189894
R23226 commonsourceibias.n589 commonsourceibias.n588 0.189894
R23227 commonsourceibias.n590 commonsourceibias.n589 0.189894
R23228 commonsourceibias.n590 commonsourceibias.n373 0.189894
R23229 commonsourceibias.n595 commonsourceibias.n373 0.189894
R23230 commonsourceibias.n596 commonsourceibias.n595 0.189894
R23231 commonsourceibias.n597 commonsourceibias.n596 0.189894
R23232 commonsourceibias.n597 commonsourceibias.n371 0.189894
R23233 commonsourceibias.n603 commonsourceibias.n371 0.189894
R23234 commonsourceibias.n604 commonsourceibias.n603 0.189894
R23235 commonsourceibias.n605 commonsourceibias.n604 0.189894
R23236 commonsourceibias.n605 commonsourceibias.n369 0.189894
R23237 commonsourceibias.n610 commonsourceibias.n369 0.189894
R23238 commonsourceibias.n611 commonsourceibias.n610 0.189894
R23239 commonsourceibias.n612 commonsourceibias.n611 0.189894
R23240 commonsourceibias.n612 commonsourceibias.n367 0.189894
R23241 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R23242 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R23243 commonsourceibias.n569 commonsourceibias.n514 0.0762576
R23244 commonsourceibias.n573 commonsourceibias.n514 0.0762576
R23245 minus.n43 minus.t24 322.512
R23246 minus.n9 minus.t8 322.512
R23247 minus.n66 minus.t5 297.12
R23248 minus.n64 minus.t6 297.12
R23249 minus.n36 minus.t22 297.12
R23250 minus.n58 minus.t18 297.12
R23251 minus.n38 minus.t19 297.12
R23252 minus.n52 minus.t14 297.12
R23253 minus.n40 minus.t15 297.12
R23254 minus.n46 minus.t9 297.12
R23255 minus.n42 minus.t23 297.12
R23256 minus.n8 minus.t7 297.12
R23257 minus.n12 minus.t11 297.12
R23258 minus.n14 minus.t10 297.12
R23259 minus.n18 minus.t12 297.12
R23260 minus.n20 minus.t17 297.12
R23261 minus.n24 minus.t16 297.12
R23262 minus.n26 minus.t21 297.12
R23263 minus.n30 minus.t20 297.12
R23264 minus.n32 minus.t13 297.12
R23265 minus.n72 minus.t4 243.255
R23266 minus.n71 minus.n69 224.169
R23267 minus.n71 minus.n70 223.454
R23268 minus.n45 minus.n44 161.3
R23269 minus.n46 minus.n41 161.3
R23270 minus.n48 minus.n47 161.3
R23271 minus.n49 minus.n40 161.3
R23272 minus.n51 minus.n50 161.3
R23273 minus.n52 minus.n39 161.3
R23274 minus.n54 minus.n53 161.3
R23275 minus.n55 minus.n38 161.3
R23276 minus.n57 minus.n56 161.3
R23277 minus.n58 minus.n37 161.3
R23278 minus.n60 minus.n59 161.3
R23279 minus.n61 minus.n36 161.3
R23280 minus.n63 minus.n62 161.3
R23281 minus.n64 minus.n35 161.3
R23282 minus.n65 minus.n34 161.3
R23283 minus.n67 minus.n66 161.3
R23284 minus.n33 minus.n32 161.3
R23285 minus.n31 minus.n0 161.3
R23286 minus.n30 minus.n29 161.3
R23287 minus.n28 minus.n1 161.3
R23288 minus.n27 minus.n26 161.3
R23289 minus.n25 minus.n2 161.3
R23290 minus.n24 minus.n23 161.3
R23291 minus.n22 minus.n3 161.3
R23292 minus.n21 minus.n20 161.3
R23293 minus.n19 minus.n4 161.3
R23294 minus.n18 minus.n17 161.3
R23295 minus.n16 minus.n5 161.3
R23296 minus.n15 minus.n14 161.3
R23297 minus.n13 minus.n6 161.3
R23298 minus.n12 minus.n11 161.3
R23299 minus.n10 minus.n7 161.3
R23300 minus.n44 minus.n43 45.0031
R23301 minus.n10 minus.n9 45.0031
R23302 minus.n66 minus.n65 41.6278
R23303 minus.n32 minus.n31 41.6278
R23304 minus.n64 minus.n63 37.246
R23305 minus.n45 minus.n42 37.246
R23306 minus.n8 minus.n7 37.246
R23307 minus.n30 minus.n1 37.246
R23308 minus.n59 minus.n36 32.8641
R23309 minus.n47 minus.n46 32.8641
R23310 minus.n13 minus.n12 32.8641
R23311 minus.n26 minus.n25 32.8641
R23312 minus.n68 minus.n67 31.8206
R23313 minus.n58 minus.n57 28.4823
R23314 minus.n51 minus.n40 28.4823
R23315 minus.n14 minus.n5 28.4823
R23316 minus.n24 minus.n3 28.4823
R23317 minus.n53 minus.n38 24.1005
R23318 minus.n53 minus.n52 24.1005
R23319 minus.n19 minus.n18 24.1005
R23320 minus.n20 minus.n19 24.1005
R23321 minus.n70 minus.t3 19.8005
R23322 minus.n70 minus.t1 19.8005
R23323 minus.n69 minus.t2 19.8005
R23324 minus.n69 minus.t0 19.8005
R23325 minus.n57 minus.n38 19.7187
R23326 minus.n52 minus.n51 19.7187
R23327 minus.n18 minus.n5 19.7187
R23328 minus.n20 minus.n3 19.7187
R23329 minus.n43 minus.n42 15.6319
R23330 minus.n9 minus.n8 15.6319
R23331 minus.n59 minus.n58 15.3369
R23332 minus.n47 minus.n40 15.3369
R23333 minus.n14 minus.n13 15.3369
R23334 minus.n25 minus.n24 15.3369
R23335 minus minus.n73 12.1618
R23336 minus.n68 minus.n33 12.0819
R23337 minus.n63 minus.n36 10.955
R23338 minus.n46 minus.n45 10.955
R23339 minus.n12 minus.n7 10.955
R23340 minus.n26 minus.n1 10.955
R23341 minus.n65 minus.n64 6.57323
R23342 minus.n31 minus.n30 6.57323
R23343 minus.n73 minus.n72 4.80222
R23344 minus.n73 minus.n68 0.972091
R23345 minus.n72 minus.n71 0.716017
R23346 minus.n67 minus.n34 0.189894
R23347 minus.n35 minus.n34 0.189894
R23348 minus.n62 minus.n35 0.189894
R23349 minus.n62 minus.n61 0.189894
R23350 minus.n61 minus.n60 0.189894
R23351 minus.n60 minus.n37 0.189894
R23352 minus.n56 minus.n37 0.189894
R23353 minus.n56 minus.n55 0.189894
R23354 minus.n55 minus.n54 0.189894
R23355 minus.n54 minus.n39 0.189894
R23356 minus.n50 minus.n39 0.189894
R23357 minus.n50 minus.n49 0.189894
R23358 minus.n49 minus.n48 0.189894
R23359 minus.n48 minus.n41 0.189894
R23360 minus.n44 minus.n41 0.189894
R23361 minus.n11 minus.n10 0.189894
R23362 minus.n11 minus.n6 0.189894
R23363 minus.n15 minus.n6 0.189894
R23364 minus.n16 minus.n15 0.189894
R23365 minus.n17 minus.n16 0.189894
R23366 minus.n17 minus.n4 0.189894
R23367 minus.n21 minus.n4 0.189894
R23368 minus.n22 minus.n21 0.189894
R23369 minus.n23 minus.n22 0.189894
R23370 minus.n23 minus.n2 0.189894
R23371 minus.n27 minus.n2 0.189894
R23372 minus.n28 minus.n27 0.189894
R23373 minus.n29 minus.n28 0.189894
R23374 minus.n29 minus.n0 0.189894
R23375 minus.n33 minus.n0 0.189894
R23376 output.n41 output.n15 289.615
R23377 output.n72 output.n46 289.615
R23378 output.n104 output.n78 289.615
R23379 output.n136 output.n110 289.615
R23380 output.n77 output.n45 197.26
R23381 output.n77 output.n76 196.298
R23382 output.n109 output.n108 196.298
R23383 output.n141 output.n140 196.298
R23384 output.n42 output.n41 185
R23385 output.n40 output.n39 185
R23386 output.n19 output.n18 185
R23387 output.n34 output.n33 185
R23388 output.n32 output.n31 185
R23389 output.n23 output.n22 185
R23390 output.n26 output.n25 185
R23391 output.n73 output.n72 185
R23392 output.n71 output.n70 185
R23393 output.n50 output.n49 185
R23394 output.n65 output.n64 185
R23395 output.n63 output.n62 185
R23396 output.n54 output.n53 185
R23397 output.n57 output.n56 185
R23398 output.n105 output.n104 185
R23399 output.n103 output.n102 185
R23400 output.n82 output.n81 185
R23401 output.n97 output.n96 185
R23402 output.n95 output.n94 185
R23403 output.n86 output.n85 185
R23404 output.n89 output.n88 185
R23405 output.n137 output.n136 185
R23406 output.n135 output.n134 185
R23407 output.n114 output.n113 185
R23408 output.n129 output.n128 185
R23409 output.n127 output.n126 185
R23410 output.n118 output.n117 185
R23411 output.n121 output.n120 185
R23412 output.t19 output.n24 147.661
R23413 output.t17 output.n55 147.661
R23414 output.t18 output.n87 147.661
R23415 output.t16 output.n119 147.661
R23416 output.n41 output.n40 104.615
R23417 output.n40 output.n18 104.615
R23418 output.n33 output.n18 104.615
R23419 output.n33 output.n32 104.615
R23420 output.n32 output.n22 104.615
R23421 output.n25 output.n22 104.615
R23422 output.n72 output.n71 104.615
R23423 output.n71 output.n49 104.615
R23424 output.n64 output.n49 104.615
R23425 output.n64 output.n63 104.615
R23426 output.n63 output.n53 104.615
R23427 output.n56 output.n53 104.615
R23428 output.n104 output.n103 104.615
R23429 output.n103 output.n81 104.615
R23430 output.n96 output.n81 104.615
R23431 output.n96 output.n95 104.615
R23432 output.n95 output.n85 104.615
R23433 output.n88 output.n85 104.615
R23434 output.n136 output.n135 104.615
R23435 output.n135 output.n113 104.615
R23436 output.n128 output.n113 104.615
R23437 output.n128 output.n127 104.615
R23438 output.n127 output.n117 104.615
R23439 output.n120 output.n117 104.615
R23440 output.n1 output.t9 77.056
R23441 output.n14 output.t11 76.6694
R23442 output.n1 output.n0 72.7095
R23443 output.n3 output.n2 72.7095
R23444 output.n5 output.n4 72.7095
R23445 output.n7 output.n6 72.7095
R23446 output.n9 output.n8 72.7095
R23447 output.n11 output.n10 72.7095
R23448 output.n13 output.n12 72.7095
R23449 output.n25 output.t19 52.3082
R23450 output.n56 output.t17 52.3082
R23451 output.n88 output.t18 52.3082
R23452 output.n120 output.t16 52.3082
R23453 output.n26 output.n24 15.6674
R23454 output.n57 output.n55 15.6674
R23455 output.n89 output.n87 15.6674
R23456 output.n121 output.n119 15.6674
R23457 output.n27 output.n23 12.8005
R23458 output.n58 output.n54 12.8005
R23459 output.n90 output.n86 12.8005
R23460 output.n122 output.n118 12.8005
R23461 output.n31 output.n30 12.0247
R23462 output.n62 output.n61 12.0247
R23463 output.n94 output.n93 12.0247
R23464 output.n126 output.n125 12.0247
R23465 output.n34 output.n21 11.249
R23466 output.n65 output.n52 11.249
R23467 output.n97 output.n84 11.249
R23468 output.n129 output.n116 11.249
R23469 output.n35 output.n19 10.4732
R23470 output.n66 output.n50 10.4732
R23471 output.n98 output.n82 10.4732
R23472 output.n130 output.n114 10.4732
R23473 output.n39 output.n38 9.69747
R23474 output.n70 output.n69 9.69747
R23475 output.n102 output.n101 9.69747
R23476 output.n134 output.n133 9.69747
R23477 output.n45 output.n44 9.45567
R23478 output.n76 output.n75 9.45567
R23479 output.n108 output.n107 9.45567
R23480 output.n140 output.n139 9.45567
R23481 output.n44 output.n43 9.3005
R23482 output.n17 output.n16 9.3005
R23483 output.n38 output.n37 9.3005
R23484 output.n36 output.n35 9.3005
R23485 output.n21 output.n20 9.3005
R23486 output.n30 output.n29 9.3005
R23487 output.n28 output.n27 9.3005
R23488 output.n75 output.n74 9.3005
R23489 output.n48 output.n47 9.3005
R23490 output.n69 output.n68 9.3005
R23491 output.n67 output.n66 9.3005
R23492 output.n52 output.n51 9.3005
R23493 output.n61 output.n60 9.3005
R23494 output.n59 output.n58 9.3005
R23495 output.n107 output.n106 9.3005
R23496 output.n80 output.n79 9.3005
R23497 output.n101 output.n100 9.3005
R23498 output.n99 output.n98 9.3005
R23499 output.n84 output.n83 9.3005
R23500 output.n93 output.n92 9.3005
R23501 output.n91 output.n90 9.3005
R23502 output.n139 output.n138 9.3005
R23503 output.n112 output.n111 9.3005
R23504 output.n133 output.n132 9.3005
R23505 output.n131 output.n130 9.3005
R23506 output.n116 output.n115 9.3005
R23507 output.n125 output.n124 9.3005
R23508 output.n123 output.n122 9.3005
R23509 output.n42 output.n17 8.92171
R23510 output.n73 output.n48 8.92171
R23511 output.n105 output.n80 8.92171
R23512 output.n137 output.n112 8.92171
R23513 output output.n141 8.15037
R23514 output.n43 output.n15 8.14595
R23515 output.n74 output.n46 8.14595
R23516 output.n106 output.n78 8.14595
R23517 output.n138 output.n110 8.14595
R23518 output.n45 output.n15 5.81868
R23519 output.n76 output.n46 5.81868
R23520 output.n108 output.n78 5.81868
R23521 output.n140 output.n110 5.81868
R23522 output.n43 output.n42 5.04292
R23523 output.n74 output.n73 5.04292
R23524 output.n106 output.n105 5.04292
R23525 output.n138 output.n137 5.04292
R23526 output.n28 output.n24 4.38594
R23527 output.n59 output.n55 4.38594
R23528 output.n91 output.n87 4.38594
R23529 output.n123 output.n119 4.38594
R23530 output.n39 output.n17 4.26717
R23531 output.n70 output.n48 4.26717
R23532 output.n102 output.n80 4.26717
R23533 output.n134 output.n112 4.26717
R23534 output.n0 output.t15 3.9605
R23535 output.n0 output.t4 3.9605
R23536 output.n2 output.t8 3.9605
R23537 output.n2 output.t0 3.9605
R23538 output.n4 output.t2 3.9605
R23539 output.n4 output.t1 3.9605
R23540 output.n6 output.t7 3.9605
R23541 output.n6 output.t10 3.9605
R23542 output.n8 output.t12 3.9605
R23543 output.n8 output.t5 3.9605
R23544 output.n10 output.t6 3.9605
R23545 output.n10 output.t13 3.9605
R23546 output.n12 output.t14 3.9605
R23547 output.n12 output.t3 3.9605
R23548 output.n38 output.n19 3.49141
R23549 output.n69 output.n50 3.49141
R23550 output.n101 output.n82 3.49141
R23551 output.n133 output.n114 3.49141
R23552 output.n35 output.n34 2.71565
R23553 output.n66 output.n65 2.71565
R23554 output.n98 output.n97 2.71565
R23555 output.n130 output.n129 2.71565
R23556 output.n31 output.n21 1.93989
R23557 output.n62 output.n52 1.93989
R23558 output.n94 output.n84 1.93989
R23559 output.n126 output.n116 1.93989
R23560 output.n30 output.n23 1.16414
R23561 output.n61 output.n54 1.16414
R23562 output.n93 output.n86 1.16414
R23563 output.n125 output.n118 1.16414
R23564 output.n141 output.n109 0.962709
R23565 output.n109 output.n77 0.962709
R23566 output.n27 output.n26 0.388379
R23567 output.n58 output.n57 0.388379
R23568 output.n90 output.n89 0.388379
R23569 output.n122 output.n121 0.388379
R23570 output.n14 output.n13 0.387128
R23571 output.n13 output.n11 0.387128
R23572 output.n11 output.n9 0.387128
R23573 output.n9 output.n7 0.387128
R23574 output.n7 output.n5 0.387128
R23575 output.n5 output.n3 0.387128
R23576 output.n3 output.n1 0.387128
R23577 output.n44 output.n16 0.155672
R23578 output.n37 output.n16 0.155672
R23579 output.n37 output.n36 0.155672
R23580 output.n36 output.n20 0.155672
R23581 output.n29 output.n20 0.155672
R23582 output.n29 output.n28 0.155672
R23583 output.n75 output.n47 0.155672
R23584 output.n68 output.n47 0.155672
R23585 output.n68 output.n67 0.155672
R23586 output.n67 output.n51 0.155672
R23587 output.n60 output.n51 0.155672
R23588 output.n60 output.n59 0.155672
R23589 output.n107 output.n79 0.155672
R23590 output.n100 output.n79 0.155672
R23591 output.n100 output.n99 0.155672
R23592 output.n99 output.n83 0.155672
R23593 output.n92 output.n83 0.155672
R23594 output.n92 output.n91 0.155672
R23595 output.n139 output.n111 0.155672
R23596 output.n132 output.n111 0.155672
R23597 output.n132 output.n131 0.155672
R23598 output.n131 output.n115 0.155672
R23599 output.n124 output.n115 0.155672
R23600 output.n124 output.n123 0.155672
R23601 output output.n14 0.126227
R23602 a_n1986_8322.n6 a_n1986_8322.t5 74.6477
R23603 a_n1986_8322.n1 a_n1986_8322.t11 74.6477
R23604 a_n1986_8322.t20 a_n1986_8322.n18 74.6476
R23605 a_n1986_8322.n14 a_n1986_8322.t13 74.2899
R23606 a_n1986_8322.n7 a_n1986_8322.t3 74.2899
R23607 a_n1986_8322.n8 a_n1986_8322.t6 74.2899
R23608 a_n1986_8322.n11 a_n1986_8322.t7 74.2899
R23609 a_n1986_8322.n4 a_n1986_8322.t10 74.2899
R23610 a_n1986_8322.n18 a_n1986_8322.n17 70.6783
R23611 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R23612 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R23613 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R23614 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R23615 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R23616 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R23617 a_n1986_8322.n13 a_n1986_8322.t0 10.2757
R23618 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R23619 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R23620 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R23621 a_n1986_8322.n17 a_n1986_8322.t18 3.61217
R23622 a_n1986_8322.n17 a_n1986_8322.t15 3.61217
R23623 a_n1986_8322.n15 a_n1986_8322.t12 3.61217
R23624 a_n1986_8322.n15 a_n1986_8322.t21 3.61217
R23625 a_n1986_8322.n5 a_n1986_8322.t9 3.61217
R23626 a_n1986_8322.n5 a_n1986_8322.t8 3.61217
R23627 a_n1986_8322.n9 a_n1986_8322.t4 3.61217
R23628 a_n1986_8322.n9 a_n1986_8322.t2 3.61217
R23629 a_n1986_8322.n0 a_n1986_8322.t19 3.61217
R23630 a_n1986_8322.n0 a_n1986_8322.t14 3.61217
R23631 a_n1986_8322.n2 a_n1986_8322.t17 3.61217
R23632 a_n1986_8322.n2 a_n1986_8322.t16 3.61217
R23633 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R23634 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R23635 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R23636 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R23637 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R23638 a_n1986_8322.n16 a_n1986_8322.n14 0.358259
R23639 a_n1986_8322.n18 a_n1986_8322.n16 0.358259
R23640 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R23641 a_n1986_8322.t0 a_n1986_8322.t1 0.057021
C0 CSoutput output 6.13571f
C1 CSoutput outputibias 0.032386f
C2 vdd CSoutput 0.116309p
C3 minus diffpairibias 3.4e-19
C4 commonsourceibias output 0.006808f
C5 CSoutput minus 3.2739f
C6 vdd plus 0.081925f
C7 commonsourceibias outputibias 0.003832f
C8 plus diffpairibias 3.42e-19
C9 vdd commonsourceibias 0.004218f
C10 CSoutput plus 0.896085f
C11 commonsourceibias diffpairibias 0.052527f
C12 CSoutput commonsourceibias 45.462303f
C13 minus plus 9.93573f
C14 minus commonsourceibias 0.332601f
C15 plus commonsourceibias 0.278362f
C16 output outputibias 2.34152f
C17 vdd output 7.23429f
C18 diffpairibias gnd 59.99123f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.182005p
C22 plus gnd 35.1216f
C23 minus gnd 29.926321f
C24 CSoutput gnd 0.115858p
C25 vdd gnd 0.409034p
C26 a_n1986_8322.t1 gnd 49.329998f
C27 a_n1986_8322.t0 gnd 76.771f
C28 a_n1986_8322.t11 gnd 0.875297f
C29 a_n1986_8322.t19 gnd 0.09348f
C30 a_n1986_8322.t14 gnd 0.09348f
C31 a_n1986_8322.n0 gnd 0.658471f
C32 a_n1986_8322.n1 gnd 0.735745f
C33 a_n1986_8322.t17 gnd 0.09348f
C34 a_n1986_8322.t16 gnd 0.09348f
C35 a_n1986_8322.n2 gnd 0.658471f
C36 a_n1986_8322.n3 gnd 0.373822f
C37 a_n1986_8322.t10 gnd 0.873554f
C38 a_n1986_8322.n4 gnd 1.39817f
C39 a_n1986_8322.t5 gnd 0.875297f
C40 a_n1986_8322.t9 gnd 0.09348f
C41 a_n1986_8322.t8 gnd 0.09348f
C42 a_n1986_8322.n5 gnd 0.658471f
C43 a_n1986_8322.n6 gnd 0.735745f
C44 a_n1986_8322.t3 gnd 0.873554f
C45 a_n1986_8322.n7 gnd 0.370237f
C46 a_n1986_8322.t6 gnd 0.873554f
C47 a_n1986_8322.n8 gnd 0.370237f
C48 a_n1986_8322.t4 gnd 0.09348f
C49 a_n1986_8322.t2 gnd 0.09348f
C50 a_n1986_8322.n9 gnd 0.658471f
C51 a_n1986_8322.n10 gnd 0.373822f
C52 a_n1986_8322.t7 gnd 0.873554f
C53 a_n1986_8322.n11 gnd 0.871824f
C54 a_n1986_8322.n12 gnd 1.58981f
C55 a_n1986_8322.n13 gnd 4.0376f
C56 a_n1986_8322.t13 gnd 0.873554f
C57 a_n1986_8322.n14 gnd 0.766087f
C58 a_n1986_8322.t12 gnd 0.09348f
C59 a_n1986_8322.t21 gnd 0.09348f
C60 a_n1986_8322.n15 gnd 0.658471f
C61 a_n1986_8322.n16 gnd 0.373822f
C62 a_n1986_8322.t18 gnd 0.09348f
C63 a_n1986_8322.t15 gnd 0.09348f
C64 a_n1986_8322.n17 gnd 0.658471f
C65 a_n1986_8322.n18 gnd 0.735743f
C66 a_n1986_8322.t20 gnd 0.875299f
C67 output.t9 gnd 0.464308f
C68 output.t15 gnd 0.044422f
C69 output.t4 gnd 0.044422f
C70 output.n0 gnd 0.364624f
C71 output.n1 gnd 0.614102f
C72 output.t8 gnd 0.044422f
C73 output.t0 gnd 0.044422f
C74 output.n2 gnd 0.364624f
C75 output.n3 gnd 0.350265f
C76 output.t2 gnd 0.044422f
C77 output.t1 gnd 0.044422f
C78 output.n4 gnd 0.364624f
C79 output.n5 gnd 0.350265f
C80 output.t7 gnd 0.044422f
C81 output.t10 gnd 0.044422f
C82 output.n6 gnd 0.364624f
C83 output.n7 gnd 0.350265f
C84 output.t12 gnd 0.044422f
C85 output.t5 gnd 0.044422f
C86 output.n8 gnd 0.364624f
C87 output.n9 gnd 0.350265f
C88 output.t6 gnd 0.044422f
C89 output.t13 gnd 0.044422f
C90 output.n10 gnd 0.364624f
C91 output.n11 gnd 0.350265f
C92 output.t14 gnd 0.044422f
C93 output.t3 gnd 0.044422f
C94 output.n12 gnd 0.364624f
C95 output.n13 gnd 0.350265f
C96 output.t11 gnd 0.462979f
C97 output.n14 gnd 0.28994f
C98 output.n15 gnd 0.015803f
C99 output.n16 gnd 0.011243f
C100 output.n17 gnd 0.006041f
C101 output.n18 gnd 0.01428f
C102 output.n19 gnd 0.006397f
C103 output.n20 gnd 0.011243f
C104 output.n21 gnd 0.006041f
C105 output.n22 gnd 0.01428f
C106 output.n23 gnd 0.006397f
C107 output.n24 gnd 0.048111f
C108 output.t19 gnd 0.023274f
C109 output.n25 gnd 0.01071f
C110 output.n26 gnd 0.008435f
C111 output.n27 gnd 0.006041f
C112 output.n28 gnd 0.267512f
C113 output.n29 gnd 0.011243f
C114 output.n30 gnd 0.006041f
C115 output.n31 gnd 0.006397f
C116 output.n32 gnd 0.01428f
C117 output.n33 gnd 0.01428f
C118 output.n34 gnd 0.006397f
C119 output.n35 gnd 0.006041f
C120 output.n36 gnd 0.011243f
C121 output.n37 gnd 0.011243f
C122 output.n38 gnd 0.006041f
C123 output.n39 gnd 0.006397f
C124 output.n40 gnd 0.01428f
C125 output.n41 gnd 0.030913f
C126 output.n42 gnd 0.006397f
C127 output.n43 gnd 0.006041f
C128 output.n44 gnd 0.025987f
C129 output.n45 gnd 0.097665f
C130 output.n46 gnd 0.015803f
C131 output.n47 gnd 0.011243f
C132 output.n48 gnd 0.006041f
C133 output.n49 gnd 0.01428f
C134 output.n50 gnd 0.006397f
C135 output.n51 gnd 0.011243f
C136 output.n52 gnd 0.006041f
C137 output.n53 gnd 0.01428f
C138 output.n54 gnd 0.006397f
C139 output.n55 gnd 0.048111f
C140 output.t17 gnd 0.023274f
C141 output.n56 gnd 0.01071f
C142 output.n57 gnd 0.008435f
C143 output.n58 gnd 0.006041f
C144 output.n59 gnd 0.267512f
C145 output.n60 gnd 0.011243f
C146 output.n61 gnd 0.006041f
C147 output.n62 gnd 0.006397f
C148 output.n63 gnd 0.01428f
C149 output.n64 gnd 0.01428f
C150 output.n65 gnd 0.006397f
C151 output.n66 gnd 0.006041f
C152 output.n67 gnd 0.011243f
C153 output.n68 gnd 0.011243f
C154 output.n69 gnd 0.006041f
C155 output.n70 gnd 0.006397f
C156 output.n71 gnd 0.01428f
C157 output.n72 gnd 0.030913f
C158 output.n73 gnd 0.006397f
C159 output.n74 gnd 0.006041f
C160 output.n75 gnd 0.025987f
C161 output.n76 gnd 0.09306f
C162 output.n77 gnd 1.65264f
C163 output.n78 gnd 0.015803f
C164 output.n79 gnd 0.011243f
C165 output.n80 gnd 0.006041f
C166 output.n81 gnd 0.01428f
C167 output.n82 gnd 0.006397f
C168 output.n83 gnd 0.011243f
C169 output.n84 gnd 0.006041f
C170 output.n85 gnd 0.01428f
C171 output.n86 gnd 0.006397f
C172 output.n87 gnd 0.048111f
C173 output.t18 gnd 0.023274f
C174 output.n88 gnd 0.01071f
C175 output.n89 gnd 0.008435f
C176 output.n90 gnd 0.006041f
C177 output.n91 gnd 0.267512f
C178 output.n92 gnd 0.011243f
C179 output.n93 gnd 0.006041f
C180 output.n94 gnd 0.006397f
C181 output.n95 gnd 0.01428f
C182 output.n96 gnd 0.01428f
C183 output.n97 gnd 0.006397f
C184 output.n98 gnd 0.006041f
C185 output.n99 gnd 0.011243f
C186 output.n100 gnd 0.011243f
C187 output.n101 gnd 0.006041f
C188 output.n102 gnd 0.006397f
C189 output.n103 gnd 0.01428f
C190 output.n104 gnd 0.030913f
C191 output.n105 gnd 0.006397f
C192 output.n106 gnd 0.006041f
C193 output.n107 gnd 0.025987f
C194 output.n108 gnd 0.09306f
C195 output.n109 gnd 0.713089f
C196 output.n110 gnd 0.015803f
C197 output.n111 gnd 0.011243f
C198 output.n112 gnd 0.006041f
C199 output.n113 gnd 0.01428f
C200 output.n114 gnd 0.006397f
C201 output.n115 gnd 0.011243f
C202 output.n116 gnd 0.006041f
C203 output.n117 gnd 0.01428f
C204 output.n118 gnd 0.006397f
C205 output.n119 gnd 0.048111f
C206 output.t16 gnd 0.023274f
C207 output.n120 gnd 0.01071f
C208 output.n121 gnd 0.008435f
C209 output.n122 gnd 0.006041f
C210 output.n123 gnd 0.267512f
C211 output.n124 gnd 0.011243f
C212 output.n125 gnd 0.006041f
C213 output.n126 gnd 0.006397f
C214 output.n127 gnd 0.01428f
C215 output.n128 gnd 0.01428f
C216 output.n129 gnd 0.006397f
C217 output.n130 gnd 0.006041f
C218 output.n131 gnd 0.011243f
C219 output.n132 gnd 0.011243f
C220 output.n133 gnd 0.006041f
C221 output.n134 gnd 0.006397f
C222 output.n135 gnd 0.01428f
C223 output.n136 gnd 0.030913f
C224 output.n137 gnd 0.006397f
C225 output.n138 gnd 0.006041f
C226 output.n139 gnd 0.025987f
C227 output.n140 gnd 0.09306f
C228 output.n141 gnd 1.67353f
C229 minus.n0 gnd 0.030538f
C230 minus.n1 gnd 0.00693f
C231 minus.n2 gnd 0.030538f
C232 minus.n3 gnd 0.00693f
C233 minus.n4 gnd 0.030538f
C234 minus.n5 gnd 0.00693f
C235 minus.n6 gnd 0.030538f
C236 minus.n7 gnd 0.00693f
C237 minus.t8 gnd 0.447069f
C238 minus.t7 gnd 0.431937f
C239 minus.n8 gnd 0.196988f
C240 minus.n9 gnd 0.17894f
C241 minus.n10 gnd 0.13035f
C242 minus.n11 gnd 0.030538f
C243 minus.t11 gnd 0.431937f
C244 minus.n12 gnd 0.19188f
C245 minus.n13 gnd 0.00693f
C246 minus.t10 gnd 0.431937f
C247 minus.n14 gnd 0.19188f
C248 minus.n15 gnd 0.030538f
C249 minus.n16 gnd 0.030538f
C250 minus.n17 gnd 0.030538f
C251 minus.t12 gnd 0.431937f
C252 minus.n18 gnd 0.19188f
C253 minus.n19 gnd 0.00693f
C254 minus.t17 gnd 0.431937f
C255 minus.n20 gnd 0.19188f
C256 minus.n21 gnd 0.030538f
C257 minus.n22 gnd 0.030538f
C258 minus.n23 gnd 0.030538f
C259 minus.t16 gnd 0.431937f
C260 minus.n24 gnd 0.19188f
C261 minus.n25 gnd 0.00693f
C262 minus.t21 gnd 0.431937f
C263 minus.n26 gnd 0.19188f
C264 minus.n27 gnd 0.030538f
C265 minus.n28 gnd 0.030538f
C266 minus.n29 gnd 0.030538f
C267 minus.t20 gnd 0.431937f
C268 minus.n30 gnd 0.19188f
C269 minus.n31 gnd 0.00693f
C270 minus.t13 gnd 0.431937f
C271 minus.n32 gnd 0.191598f
C272 minus.n33 gnd 0.352847f
C273 minus.n34 gnd 0.030538f
C274 minus.t5 gnd 0.431937f
C275 minus.t6 gnd 0.431937f
C276 minus.n35 gnd 0.030538f
C277 minus.t22 gnd 0.431937f
C278 minus.n36 gnd 0.19188f
C279 minus.n37 gnd 0.030538f
C280 minus.t18 gnd 0.431937f
C281 minus.t19 gnd 0.431937f
C282 minus.n38 gnd 0.19188f
C283 minus.n39 gnd 0.030538f
C284 minus.t14 gnd 0.431937f
C285 minus.t15 gnd 0.431937f
C286 minus.n40 gnd 0.19188f
C287 minus.n41 gnd 0.030538f
C288 minus.t9 gnd 0.431937f
C289 minus.t23 gnd 0.431937f
C290 minus.n42 gnd 0.196988f
C291 minus.t24 gnd 0.447069f
C292 minus.n43 gnd 0.17894f
C293 minus.n44 gnd 0.13035f
C294 minus.n45 gnd 0.00693f
C295 minus.n46 gnd 0.19188f
C296 minus.n47 gnd 0.00693f
C297 minus.n48 gnd 0.030538f
C298 minus.n49 gnd 0.030538f
C299 minus.n50 gnd 0.030538f
C300 minus.n51 gnd 0.00693f
C301 minus.n52 gnd 0.19188f
C302 minus.n53 gnd 0.00693f
C303 minus.n54 gnd 0.030538f
C304 minus.n55 gnd 0.030538f
C305 minus.n56 gnd 0.030538f
C306 minus.n57 gnd 0.00693f
C307 minus.n58 gnd 0.19188f
C308 minus.n59 gnd 0.00693f
C309 minus.n60 gnd 0.030538f
C310 minus.n61 gnd 0.030538f
C311 minus.n62 gnd 0.030538f
C312 minus.n63 gnd 0.00693f
C313 minus.n64 gnd 0.19188f
C314 minus.n65 gnd 0.00693f
C315 minus.n66 gnd 0.191598f
C316 minus.n67 gnd 0.954237f
C317 minus.n68 gnd 1.43659f
C318 minus.t2 gnd 0.009414f
C319 minus.t0 gnd 0.009414f
C320 minus.n69 gnd 0.030956f
C321 minus.t3 gnd 0.009414f
C322 minus.t1 gnd 0.009414f
C323 minus.n70 gnd 0.030532f
C324 minus.n71 gnd 0.260573f
C325 minus.t4 gnd 0.052398f
C326 minus.n72 gnd 0.142192f
C327 minus.n73 gnd 2.36188f
C328 commonsourceibias.n0 gnd 0.010724f
C329 commonsourceibias.t115 gnd 0.162395f
C330 commonsourceibias.t136 gnd 0.150157f
C331 commonsourceibias.n1 gnd 0.007823f
C332 commonsourceibias.n2 gnd 0.008037f
C333 commonsourceibias.t151 gnd 0.150157f
C334 commonsourceibias.n3 gnd 0.01034f
C335 commonsourceibias.n4 gnd 0.008037f
C336 commonsourceibias.t105 gnd 0.150157f
C337 commonsourceibias.n5 gnd 0.059912f
C338 commonsourceibias.t126 gnd 0.150157f
C339 commonsourceibias.n6 gnd 0.007578f
C340 commonsourceibias.n7 gnd 0.008037f
C341 commonsourceibias.t144 gnd 0.150157f
C342 commonsourceibias.n8 gnd 0.010186f
C343 commonsourceibias.n9 gnd 0.008037f
C344 commonsourceibias.t98 gnd 0.150157f
C345 commonsourceibias.n10 gnd 0.059912f
C346 commonsourceibias.t94 gnd 0.150157f
C347 commonsourceibias.n11 gnd 0.007361f
C348 commonsourceibias.n12 gnd 0.008037f
C349 commonsourceibias.t135 gnd 0.150157f
C350 commonsourceibias.n13 gnd 0.010015f
C351 commonsourceibias.n14 gnd 0.010724f
C352 commonsourceibias.t74 gnd 0.162395f
C353 commonsourceibias.t20 gnd 0.150157f
C354 commonsourceibias.n15 gnd 0.007823f
C355 commonsourceibias.n16 gnd 0.008037f
C356 commonsourceibias.t50 gnd 0.150157f
C357 commonsourceibias.n17 gnd 0.01034f
C358 commonsourceibias.n18 gnd 0.008037f
C359 commonsourceibias.t8 gnd 0.150157f
C360 commonsourceibias.n19 gnd 0.059912f
C361 commonsourceibias.t36 gnd 0.150157f
C362 commonsourceibias.n20 gnd 0.007578f
C363 commonsourceibias.n21 gnd 0.008037f
C364 commonsourceibias.t76 gnd 0.150157f
C365 commonsourceibias.n22 gnd 0.010186f
C366 commonsourceibias.n23 gnd 0.008037f
C367 commonsourceibias.t24 gnd 0.150157f
C368 commonsourceibias.n24 gnd 0.059912f
C369 commonsourceibias.t34 gnd 0.150157f
C370 commonsourceibias.n25 gnd 0.007361f
C371 commonsourceibias.n26 gnd 0.008037f
C372 commonsourceibias.t10 gnd 0.150157f
C373 commonsourceibias.n27 gnd 0.010015f
C374 commonsourceibias.n28 gnd 0.008037f
C375 commonsourceibias.t40 gnd 0.150157f
C376 commonsourceibias.n29 gnd 0.059912f
C377 commonsourceibias.t56 gnd 0.150157f
C378 commonsourceibias.n30 gnd 0.007172f
C379 commonsourceibias.n31 gnd 0.008037f
C380 commonsourceibias.t26 gnd 0.150157f
C381 commonsourceibias.n32 gnd 0.009825f
C382 commonsourceibias.n33 gnd 0.008037f
C383 commonsourceibias.t38 gnd 0.150157f
C384 commonsourceibias.n34 gnd 0.059912f
C385 commonsourceibias.t70 gnd 0.150157f
C386 commonsourceibias.n35 gnd 0.007008f
C387 commonsourceibias.n36 gnd 0.008037f
C388 commonsourceibias.t18 gnd 0.150157f
C389 commonsourceibias.n37 gnd 0.009613f
C390 commonsourceibias.n38 gnd 0.008037f
C391 commonsourceibias.t22 gnd 0.150157f
C392 commonsourceibias.n39 gnd 0.059912f
C393 commonsourceibias.t54 gnd 0.150157f
C394 commonsourceibias.n40 gnd 0.006868f
C395 commonsourceibias.n41 gnd 0.008037f
C396 commonsourceibias.t4 gnd 0.150157f
C397 commonsourceibias.n42 gnd 0.009378f
C398 commonsourceibias.t78 gnd 0.166947f
C399 commonsourceibias.t46 gnd 0.150157f
C400 commonsourceibias.n43 gnd 0.065449f
C401 commonsourceibias.n44 gnd 0.071822f
C402 commonsourceibias.n45 gnd 0.033327f
C403 commonsourceibias.n46 gnd 0.008037f
C404 commonsourceibias.n47 gnd 0.007823f
C405 commonsourceibias.n48 gnd 0.01121f
C406 commonsourceibias.n49 gnd 0.059912f
C407 commonsourceibias.n50 gnd 0.011203f
C408 commonsourceibias.n51 gnd 0.008037f
C409 commonsourceibias.n52 gnd 0.008037f
C410 commonsourceibias.n53 gnd 0.008037f
C411 commonsourceibias.n54 gnd 0.01034f
C412 commonsourceibias.n55 gnd 0.059912f
C413 commonsourceibias.n56 gnd 0.010583f
C414 commonsourceibias.n57 gnd 0.010282f
C415 commonsourceibias.n58 gnd 0.008037f
C416 commonsourceibias.n59 gnd 0.008037f
C417 commonsourceibias.n60 gnd 0.008037f
C418 commonsourceibias.n61 gnd 0.007578f
C419 commonsourceibias.n62 gnd 0.01122f
C420 commonsourceibias.n63 gnd 0.059912f
C421 commonsourceibias.n64 gnd 0.011217f
C422 commonsourceibias.n65 gnd 0.008037f
C423 commonsourceibias.n66 gnd 0.008037f
C424 commonsourceibias.n67 gnd 0.008037f
C425 commonsourceibias.n68 gnd 0.010186f
C426 commonsourceibias.n69 gnd 0.059912f
C427 commonsourceibias.n70 gnd 0.010507f
C428 commonsourceibias.n71 gnd 0.010357f
C429 commonsourceibias.n72 gnd 0.008037f
C430 commonsourceibias.n73 gnd 0.008037f
C431 commonsourceibias.n74 gnd 0.008037f
C432 commonsourceibias.n75 gnd 0.007361f
C433 commonsourceibias.n76 gnd 0.011225f
C434 commonsourceibias.n77 gnd 0.059912f
C435 commonsourceibias.n78 gnd 0.011224f
C436 commonsourceibias.n79 gnd 0.008037f
C437 commonsourceibias.n80 gnd 0.008037f
C438 commonsourceibias.n81 gnd 0.008037f
C439 commonsourceibias.n82 gnd 0.010015f
C440 commonsourceibias.n83 gnd 0.059912f
C441 commonsourceibias.n84 gnd 0.010432f
C442 commonsourceibias.n85 gnd 0.010432f
C443 commonsourceibias.n86 gnd 0.008037f
C444 commonsourceibias.n87 gnd 0.008037f
C445 commonsourceibias.n88 gnd 0.008037f
C446 commonsourceibias.n89 gnd 0.007172f
C447 commonsourceibias.n90 gnd 0.011224f
C448 commonsourceibias.n91 gnd 0.059912f
C449 commonsourceibias.n92 gnd 0.011225f
C450 commonsourceibias.n93 gnd 0.008037f
C451 commonsourceibias.n94 gnd 0.008037f
C452 commonsourceibias.n95 gnd 0.008037f
C453 commonsourceibias.n96 gnd 0.009825f
C454 commonsourceibias.n97 gnd 0.059912f
C455 commonsourceibias.n98 gnd 0.010357f
C456 commonsourceibias.n99 gnd 0.010507f
C457 commonsourceibias.n100 gnd 0.008037f
C458 commonsourceibias.n101 gnd 0.008037f
C459 commonsourceibias.n102 gnd 0.008037f
C460 commonsourceibias.n103 gnd 0.007008f
C461 commonsourceibias.n104 gnd 0.011217f
C462 commonsourceibias.n105 gnd 0.059912f
C463 commonsourceibias.n106 gnd 0.01122f
C464 commonsourceibias.n107 gnd 0.008037f
C465 commonsourceibias.n108 gnd 0.008037f
C466 commonsourceibias.n109 gnd 0.008037f
C467 commonsourceibias.n110 gnd 0.009613f
C468 commonsourceibias.n111 gnd 0.059912f
C469 commonsourceibias.n112 gnd 0.010282f
C470 commonsourceibias.n113 gnd 0.010583f
C471 commonsourceibias.n114 gnd 0.008037f
C472 commonsourceibias.n115 gnd 0.008037f
C473 commonsourceibias.n116 gnd 0.008037f
C474 commonsourceibias.n117 gnd 0.006868f
C475 commonsourceibias.n118 gnd 0.011203f
C476 commonsourceibias.n119 gnd 0.059912f
C477 commonsourceibias.n120 gnd 0.01121f
C478 commonsourceibias.n121 gnd 0.008037f
C479 commonsourceibias.n122 gnd 0.008037f
C480 commonsourceibias.n123 gnd 0.008037f
C481 commonsourceibias.n124 gnd 0.009378f
C482 commonsourceibias.n125 gnd 0.059912f
C483 commonsourceibias.n126 gnd 0.009861f
C484 commonsourceibias.n127 gnd 0.07189f
C485 commonsourceibias.n128 gnd 0.080075f
C486 commonsourceibias.t75 gnd 0.017343f
C487 commonsourceibias.t21 gnd 0.017343f
C488 commonsourceibias.n129 gnd 0.15325f
C489 commonsourceibias.n130 gnd 0.132562f
C490 commonsourceibias.t51 gnd 0.017343f
C491 commonsourceibias.t9 gnd 0.017343f
C492 commonsourceibias.n131 gnd 0.15325f
C493 commonsourceibias.n132 gnd 0.070394f
C494 commonsourceibias.t37 gnd 0.017343f
C495 commonsourceibias.t77 gnd 0.017343f
C496 commonsourceibias.n133 gnd 0.15325f
C497 commonsourceibias.n134 gnd 0.070394f
C498 commonsourceibias.t25 gnd 0.017343f
C499 commonsourceibias.t35 gnd 0.017343f
C500 commonsourceibias.n135 gnd 0.15325f
C501 commonsourceibias.n136 gnd 0.070394f
C502 commonsourceibias.t11 gnd 0.017343f
C503 commonsourceibias.t41 gnd 0.017343f
C504 commonsourceibias.n137 gnd 0.15325f
C505 commonsourceibias.n138 gnd 0.058811f
C506 commonsourceibias.t47 gnd 0.017343f
C507 commonsourceibias.t79 gnd 0.017343f
C508 commonsourceibias.n139 gnd 0.153763f
C509 commonsourceibias.t55 gnd 0.017343f
C510 commonsourceibias.t5 gnd 0.017343f
C511 commonsourceibias.n140 gnd 0.15325f
C512 commonsourceibias.n141 gnd 0.1428f
C513 commonsourceibias.t19 gnd 0.017343f
C514 commonsourceibias.t23 gnd 0.017343f
C515 commonsourceibias.n142 gnd 0.15325f
C516 commonsourceibias.n143 gnd 0.070394f
C517 commonsourceibias.t39 gnd 0.017343f
C518 commonsourceibias.t71 gnd 0.017343f
C519 commonsourceibias.n144 gnd 0.15325f
C520 commonsourceibias.n145 gnd 0.070394f
C521 commonsourceibias.t57 gnd 0.017343f
C522 commonsourceibias.t27 gnd 0.017343f
C523 commonsourceibias.n146 gnd 0.15325f
C524 commonsourceibias.n147 gnd 0.058811f
C525 commonsourceibias.n148 gnd 0.071213f
C526 commonsourceibias.n149 gnd 0.052016f
C527 commonsourceibias.t153 gnd 0.150157f
C528 commonsourceibias.n150 gnd 0.059912f
C529 commonsourceibias.t88 gnd 0.150157f
C530 commonsourceibias.n151 gnd 0.059912f
C531 commonsourceibias.n152 gnd 0.008037f
C532 commonsourceibias.t125 gnd 0.150157f
C533 commonsourceibias.n153 gnd 0.059912f
C534 commonsourceibias.n154 gnd 0.008037f
C535 commonsourceibias.t120 gnd 0.150157f
C536 commonsourceibias.n155 gnd 0.059912f
C537 commonsourceibias.n156 gnd 0.008037f
C538 commonsourceibias.t139 gnd 0.150157f
C539 commonsourceibias.n157 gnd 0.007008f
C540 commonsourceibias.n158 gnd 0.008037f
C541 commonsourceibias.t112 gnd 0.150157f
C542 commonsourceibias.n159 gnd 0.009613f
C543 commonsourceibias.n160 gnd 0.008037f
C544 commonsourceibias.t107 gnd 0.150157f
C545 commonsourceibias.n161 gnd 0.059912f
C546 commonsourceibias.t127 gnd 0.150157f
C547 commonsourceibias.n162 gnd 0.006868f
C548 commonsourceibias.n163 gnd 0.008037f
C549 commonsourceibias.t146 gnd 0.150157f
C550 commonsourceibias.n164 gnd 0.009378f
C551 commonsourceibias.t117 gnd 0.166947f
C552 commonsourceibias.t99 gnd 0.150157f
C553 commonsourceibias.n165 gnd 0.065449f
C554 commonsourceibias.n166 gnd 0.071822f
C555 commonsourceibias.n167 gnd 0.033327f
C556 commonsourceibias.n168 gnd 0.008037f
C557 commonsourceibias.n169 gnd 0.007823f
C558 commonsourceibias.n170 gnd 0.01121f
C559 commonsourceibias.n171 gnd 0.059912f
C560 commonsourceibias.n172 gnd 0.011203f
C561 commonsourceibias.n173 gnd 0.008037f
C562 commonsourceibias.n174 gnd 0.008037f
C563 commonsourceibias.n175 gnd 0.008037f
C564 commonsourceibias.n176 gnd 0.01034f
C565 commonsourceibias.n177 gnd 0.059912f
C566 commonsourceibias.n178 gnd 0.010583f
C567 commonsourceibias.n179 gnd 0.010282f
C568 commonsourceibias.n180 gnd 0.008037f
C569 commonsourceibias.n181 gnd 0.008037f
C570 commonsourceibias.n182 gnd 0.008037f
C571 commonsourceibias.n183 gnd 0.007578f
C572 commonsourceibias.n184 gnd 0.01122f
C573 commonsourceibias.n185 gnd 0.059912f
C574 commonsourceibias.n186 gnd 0.011217f
C575 commonsourceibias.n187 gnd 0.008037f
C576 commonsourceibias.n188 gnd 0.008037f
C577 commonsourceibias.n189 gnd 0.008037f
C578 commonsourceibias.n190 gnd 0.010186f
C579 commonsourceibias.n191 gnd 0.059912f
C580 commonsourceibias.n192 gnd 0.010507f
C581 commonsourceibias.n193 gnd 0.010357f
C582 commonsourceibias.n194 gnd 0.008037f
C583 commonsourceibias.n195 gnd 0.008037f
C584 commonsourceibias.n196 gnd 0.009825f
C585 commonsourceibias.n197 gnd 0.007361f
C586 commonsourceibias.n198 gnd 0.011225f
C587 commonsourceibias.n199 gnd 0.008037f
C588 commonsourceibias.n200 gnd 0.008037f
C589 commonsourceibias.n201 gnd 0.011224f
C590 commonsourceibias.n202 gnd 0.007172f
C591 commonsourceibias.n203 gnd 0.010015f
C592 commonsourceibias.n204 gnd 0.008037f
C593 commonsourceibias.n205 gnd 0.007021f
C594 commonsourceibias.n206 gnd 0.010432f
C595 commonsourceibias.n207 gnd 0.010432f
C596 commonsourceibias.n208 gnd 0.007021f
C597 commonsourceibias.n209 gnd 0.008037f
C598 commonsourceibias.n210 gnd 0.008037f
C599 commonsourceibias.n211 gnd 0.007172f
C600 commonsourceibias.n212 gnd 0.011224f
C601 commonsourceibias.n213 gnd 0.059912f
C602 commonsourceibias.n214 gnd 0.011225f
C603 commonsourceibias.n215 gnd 0.008037f
C604 commonsourceibias.n216 gnd 0.008037f
C605 commonsourceibias.n217 gnd 0.008037f
C606 commonsourceibias.n218 gnd 0.009825f
C607 commonsourceibias.n219 gnd 0.059912f
C608 commonsourceibias.n220 gnd 0.010357f
C609 commonsourceibias.n221 gnd 0.010507f
C610 commonsourceibias.n222 gnd 0.008037f
C611 commonsourceibias.n223 gnd 0.008037f
C612 commonsourceibias.n224 gnd 0.008037f
C613 commonsourceibias.n225 gnd 0.007008f
C614 commonsourceibias.n226 gnd 0.011217f
C615 commonsourceibias.n227 gnd 0.059912f
C616 commonsourceibias.n228 gnd 0.01122f
C617 commonsourceibias.n229 gnd 0.008037f
C618 commonsourceibias.n230 gnd 0.008037f
C619 commonsourceibias.n231 gnd 0.008037f
C620 commonsourceibias.n232 gnd 0.009613f
C621 commonsourceibias.n233 gnd 0.059912f
C622 commonsourceibias.n234 gnd 0.010282f
C623 commonsourceibias.n235 gnd 0.010583f
C624 commonsourceibias.n236 gnd 0.008037f
C625 commonsourceibias.n237 gnd 0.008037f
C626 commonsourceibias.n238 gnd 0.008037f
C627 commonsourceibias.n239 gnd 0.006868f
C628 commonsourceibias.n240 gnd 0.011203f
C629 commonsourceibias.n241 gnd 0.059912f
C630 commonsourceibias.n242 gnd 0.01121f
C631 commonsourceibias.n243 gnd 0.008037f
C632 commonsourceibias.n244 gnd 0.008037f
C633 commonsourceibias.n245 gnd 0.008037f
C634 commonsourceibias.n246 gnd 0.009378f
C635 commonsourceibias.n247 gnd 0.059912f
C636 commonsourceibias.n248 gnd 0.009861f
C637 commonsourceibias.n249 gnd 0.07189f
C638 commonsourceibias.n250 gnd 0.04697f
C639 commonsourceibias.n251 gnd 0.010724f
C640 commonsourceibias.t119 gnd 0.150157f
C641 commonsourceibias.n252 gnd 0.007823f
C642 commonsourceibias.n253 gnd 0.008037f
C643 commonsourceibias.t137 gnd 0.150157f
C644 commonsourceibias.n254 gnd 0.01034f
C645 commonsourceibias.n255 gnd 0.008037f
C646 commonsourceibias.t92 gnd 0.150157f
C647 commonsourceibias.n256 gnd 0.059912f
C648 commonsourceibias.t109 gnd 0.150157f
C649 commonsourceibias.n257 gnd 0.007578f
C650 commonsourceibias.n258 gnd 0.008037f
C651 commonsourceibias.t128 gnd 0.150157f
C652 commonsourceibias.n259 gnd 0.010186f
C653 commonsourceibias.n260 gnd 0.008037f
C654 commonsourceibias.t86 gnd 0.150157f
C655 commonsourceibias.n261 gnd 0.059912f
C656 commonsourceibias.t83 gnd 0.150157f
C657 commonsourceibias.n262 gnd 0.007361f
C658 commonsourceibias.n263 gnd 0.008037f
C659 commonsourceibias.t118 gnd 0.150157f
C660 commonsourceibias.n264 gnd 0.010015f
C661 commonsourceibias.n265 gnd 0.008037f
C662 commonsourceibias.t138 gnd 0.150157f
C663 commonsourceibias.n266 gnd 0.059912f
C664 commonsourceibias.t159 gnd 0.150157f
C665 commonsourceibias.n267 gnd 0.007172f
C666 commonsourceibias.n268 gnd 0.008037f
C667 commonsourceibias.t108 gnd 0.150157f
C668 commonsourceibias.n269 gnd 0.009825f
C669 commonsourceibias.n270 gnd 0.008037f
C670 commonsourceibias.t102 gnd 0.150157f
C671 commonsourceibias.n271 gnd 0.059912f
C672 commonsourceibias.t121 gnd 0.150157f
C673 commonsourceibias.n272 gnd 0.007008f
C674 commonsourceibias.n273 gnd 0.008037f
C675 commonsourceibias.t95 gnd 0.150157f
C676 commonsourceibias.n274 gnd 0.009613f
C677 commonsourceibias.n275 gnd 0.008037f
C678 commonsourceibias.t93 gnd 0.150157f
C679 commonsourceibias.n276 gnd 0.059912f
C680 commonsourceibias.t110 gnd 0.150157f
C681 commonsourceibias.n277 gnd 0.006868f
C682 commonsourceibias.n278 gnd 0.008037f
C683 commonsourceibias.t129 gnd 0.150157f
C684 commonsourceibias.n279 gnd 0.009378f
C685 commonsourceibias.t101 gnd 0.166947f
C686 commonsourceibias.t87 gnd 0.150157f
C687 commonsourceibias.n280 gnd 0.065449f
C688 commonsourceibias.n281 gnd 0.071822f
C689 commonsourceibias.n282 gnd 0.033327f
C690 commonsourceibias.n283 gnd 0.008037f
C691 commonsourceibias.n284 gnd 0.007823f
C692 commonsourceibias.n285 gnd 0.01121f
C693 commonsourceibias.n286 gnd 0.059912f
C694 commonsourceibias.n287 gnd 0.011203f
C695 commonsourceibias.n288 gnd 0.008037f
C696 commonsourceibias.n289 gnd 0.008037f
C697 commonsourceibias.n290 gnd 0.008037f
C698 commonsourceibias.n291 gnd 0.01034f
C699 commonsourceibias.n292 gnd 0.059912f
C700 commonsourceibias.n293 gnd 0.010583f
C701 commonsourceibias.n294 gnd 0.010282f
C702 commonsourceibias.n295 gnd 0.008037f
C703 commonsourceibias.n296 gnd 0.008037f
C704 commonsourceibias.n297 gnd 0.008037f
C705 commonsourceibias.n298 gnd 0.007578f
C706 commonsourceibias.n299 gnd 0.01122f
C707 commonsourceibias.n300 gnd 0.059912f
C708 commonsourceibias.n301 gnd 0.011217f
C709 commonsourceibias.n302 gnd 0.008037f
C710 commonsourceibias.n303 gnd 0.008037f
C711 commonsourceibias.n304 gnd 0.008037f
C712 commonsourceibias.n305 gnd 0.010186f
C713 commonsourceibias.n306 gnd 0.059912f
C714 commonsourceibias.n307 gnd 0.010507f
C715 commonsourceibias.n308 gnd 0.010357f
C716 commonsourceibias.n309 gnd 0.008037f
C717 commonsourceibias.n310 gnd 0.008037f
C718 commonsourceibias.n311 gnd 0.008037f
C719 commonsourceibias.n312 gnd 0.007361f
C720 commonsourceibias.n313 gnd 0.011225f
C721 commonsourceibias.n314 gnd 0.059912f
C722 commonsourceibias.n315 gnd 0.011224f
C723 commonsourceibias.n316 gnd 0.008037f
C724 commonsourceibias.n317 gnd 0.008037f
C725 commonsourceibias.n318 gnd 0.008037f
C726 commonsourceibias.n319 gnd 0.010015f
C727 commonsourceibias.n320 gnd 0.059912f
C728 commonsourceibias.n321 gnd 0.010432f
C729 commonsourceibias.n322 gnd 0.010432f
C730 commonsourceibias.n323 gnd 0.008037f
C731 commonsourceibias.n324 gnd 0.008037f
C732 commonsourceibias.n325 gnd 0.008037f
C733 commonsourceibias.n326 gnd 0.007172f
C734 commonsourceibias.n327 gnd 0.011224f
C735 commonsourceibias.n328 gnd 0.059912f
C736 commonsourceibias.n329 gnd 0.011225f
C737 commonsourceibias.n330 gnd 0.008037f
C738 commonsourceibias.n331 gnd 0.008037f
C739 commonsourceibias.n332 gnd 0.008037f
C740 commonsourceibias.n333 gnd 0.009825f
C741 commonsourceibias.n334 gnd 0.059912f
C742 commonsourceibias.n335 gnd 0.010357f
C743 commonsourceibias.n336 gnd 0.010507f
C744 commonsourceibias.n337 gnd 0.008037f
C745 commonsourceibias.n338 gnd 0.008037f
C746 commonsourceibias.n339 gnd 0.008037f
C747 commonsourceibias.n340 gnd 0.007008f
C748 commonsourceibias.n341 gnd 0.011217f
C749 commonsourceibias.n342 gnd 0.059912f
C750 commonsourceibias.n343 gnd 0.01122f
C751 commonsourceibias.n344 gnd 0.008037f
C752 commonsourceibias.n345 gnd 0.008037f
C753 commonsourceibias.n346 gnd 0.008037f
C754 commonsourceibias.n347 gnd 0.009613f
C755 commonsourceibias.n348 gnd 0.059912f
C756 commonsourceibias.n349 gnd 0.010282f
C757 commonsourceibias.n350 gnd 0.010583f
C758 commonsourceibias.n351 gnd 0.008037f
C759 commonsourceibias.n352 gnd 0.008037f
C760 commonsourceibias.n353 gnd 0.008037f
C761 commonsourceibias.n354 gnd 0.006868f
C762 commonsourceibias.n355 gnd 0.011203f
C763 commonsourceibias.n356 gnd 0.059912f
C764 commonsourceibias.n357 gnd 0.01121f
C765 commonsourceibias.n358 gnd 0.008037f
C766 commonsourceibias.n359 gnd 0.008037f
C767 commonsourceibias.n360 gnd 0.008037f
C768 commonsourceibias.n361 gnd 0.009378f
C769 commonsourceibias.n362 gnd 0.059912f
C770 commonsourceibias.n363 gnd 0.009861f
C771 commonsourceibias.t100 gnd 0.162395f
C772 commonsourceibias.n364 gnd 0.07189f
C773 commonsourceibias.n365 gnd 0.025003f
C774 commonsourceibias.n366 gnd 0.464917f
C775 commonsourceibias.n367 gnd 0.010724f
C776 commonsourceibias.t140 gnd 0.162395f
C777 commonsourceibias.t155 gnd 0.150157f
C778 commonsourceibias.n368 gnd 0.007823f
C779 commonsourceibias.n369 gnd 0.008037f
C780 commonsourceibias.t84 gnd 0.150157f
C781 commonsourceibias.n370 gnd 0.01034f
C782 commonsourceibias.n371 gnd 0.008037f
C783 commonsourceibias.t148 gnd 0.150157f
C784 commonsourceibias.n372 gnd 0.007578f
C785 commonsourceibias.n373 gnd 0.008037f
C786 commonsourceibias.t80 gnd 0.150157f
C787 commonsourceibias.n374 gnd 0.010186f
C788 commonsourceibias.n375 gnd 0.008037f
C789 commonsourceibias.t113 gnd 0.150157f
C790 commonsourceibias.n376 gnd 0.007361f
C791 commonsourceibias.n377 gnd 0.008037f
C792 commonsourceibias.t154 gnd 0.150157f
C793 commonsourceibias.n378 gnd 0.010015f
C794 commonsourceibias.t29 gnd 0.017343f
C795 commonsourceibias.t3 gnd 0.017343f
C796 commonsourceibias.n379 gnd 0.153763f
C797 commonsourceibias.t49 gnd 0.017343f
C798 commonsourceibias.t13 gnd 0.017343f
C799 commonsourceibias.n380 gnd 0.15325f
C800 commonsourceibias.n381 gnd 0.1428f
C801 commonsourceibias.t69 gnd 0.017343f
C802 commonsourceibias.t67 gnd 0.017343f
C803 commonsourceibias.n382 gnd 0.15325f
C804 commonsourceibias.n383 gnd 0.070394f
C805 commonsourceibias.t7 gnd 0.017343f
C806 commonsourceibias.t63 gnd 0.017343f
C807 commonsourceibias.n384 gnd 0.15325f
C808 commonsourceibias.n385 gnd 0.070394f
C809 commonsourceibias.t53 gnd 0.017343f
C810 commonsourceibias.t73 gnd 0.017343f
C811 commonsourceibias.n386 gnd 0.15325f
C812 commonsourceibias.n387 gnd 0.058811f
C813 commonsourceibias.n388 gnd 0.010724f
C814 commonsourceibias.t42 gnd 0.150157f
C815 commonsourceibias.n389 gnd 0.007823f
C816 commonsourceibias.n390 gnd 0.008037f
C817 commonsourceibias.t0 gnd 0.150157f
C818 commonsourceibias.n391 gnd 0.01034f
C819 commonsourceibias.n392 gnd 0.008037f
C820 commonsourceibias.t60 gnd 0.150157f
C821 commonsourceibias.n393 gnd 0.007578f
C822 commonsourceibias.n394 gnd 0.008037f
C823 commonsourceibias.t16 gnd 0.150157f
C824 commonsourceibias.n395 gnd 0.010186f
C825 commonsourceibias.n396 gnd 0.008037f
C826 commonsourceibias.t58 gnd 0.150157f
C827 commonsourceibias.n397 gnd 0.007361f
C828 commonsourceibias.n398 gnd 0.008037f
C829 commonsourceibias.t32 gnd 0.150157f
C830 commonsourceibias.n399 gnd 0.010015f
C831 commonsourceibias.n400 gnd 0.008037f
C832 commonsourceibias.t72 gnd 0.150157f
C833 commonsourceibias.n401 gnd 0.007172f
C834 commonsourceibias.n402 gnd 0.008037f
C835 commonsourceibias.t52 gnd 0.150157f
C836 commonsourceibias.n403 gnd 0.009825f
C837 commonsourceibias.n404 gnd 0.008037f
C838 commonsourceibias.t6 gnd 0.150157f
C839 commonsourceibias.n405 gnd 0.007008f
C840 commonsourceibias.n406 gnd 0.008037f
C841 commonsourceibias.t66 gnd 0.150157f
C842 commonsourceibias.n407 gnd 0.009613f
C843 commonsourceibias.n408 gnd 0.008037f
C844 commonsourceibias.t12 gnd 0.150157f
C845 commonsourceibias.n409 gnd 0.006868f
C846 commonsourceibias.n410 gnd 0.008037f
C847 commonsourceibias.t48 gnd 0.150157f
C848 commonsourceibias.n411 gnd 0.009378f
C849 commonsourceibias.t28 gnd 0.166947f
C850 commonsourceibias.t2 gnd 0.150157f
C851 commonsourceibias.n412 gnd 0.065449f
C852 commonsourceibias.n413 gnd 0.071822f
C853 commonsourceibias.n414 gnd 0.033327f
C854 commonsourceibias.n415 gnd 0.008037f
C855 commonsourceibias.n416 gnd 0.007823f
C856 commonsourceibias.n417 gnd 0.01121f
C857 commonsourceibias.n418 gnd 0.059912f
C858 commonsourceibias.n419 gnd 0.011203f
C859 commonsourceibias.n420 gnd 0.008037f
C860 commonsourceibias.n421 gnd 0.008037f
C861 commonsourceibias.n422 gnd 0.008037f
C862 commonsourceibias.n423 gnd 0.01034f
C863 commonsourceibias.n424 gnd 0.059912f
C864 commonsourceibias.n425 gnd 0.010583f
C865 commonsourceibias.t68 gnd 0.150157f
C866 commonsourceibias.n426 gnd 0.059912f
C867 commonsourceibias.n427 gnd 0.010282f
C868 commonsourceibias.n428 gnd 0.008037f
C869 commonsourceibias.n429 gnd 0.008037f
C870 commonsourceibias.n430 gnd 0.008037f
C871 commonsourceibias.n431 gnd 0.007578f
C872 commonsourceibias.n432 gnd 0.01122f
C873 commonsourceibias.n433 gnd 0.059912f
C874 commonsourceibias.n434 gnd 0.011217f
C875 commonsourceibias.n435 gnd 0.008037f
C876 commonsourceibias.n436 gnd 0.008037f
C877 commonsourceibias.n437 gnd 0.008037f
C878 commonsourceibias.n438 gnd 0.010186f
C879 commonsourceibias.n439 gnd 0.059912f
C880 commonsourceibias.n440 gnd 0.010507f
C881 commonsourceibias.t62 gnd 0.150157f
C882 commonsourceibias.n441 gnd 0.059912f
C883 commonsourceibias.n442 gnd 0.010357f
C884 commonsourceibias.n443 gnd 0.008037f
C885 commonsourceibias.n444 gnd 0.008037f
C886 commonsourceibias.n445 gnd 0.008037f
C887 commonsourceibias.n446 gnd 0.007361f
C888 commonsourceibias.n447 gnd 0.011225f
C889 commonsourceibias.n448 gnd 0.059912f
C890 commonsourceibias.n449 gnd 0.011224f
C891 commonsourceibias.n450 gnd 0.008037f
C892 commonsourceibias.n451 gnd 0.008037f
C893 commonsourceibias.n452 gnd 0.008037f
C894 commonsourceibias.n453 gnd 0.010015f
C895 commonsourceibias.n454 gnd 0.059912f
C896 commonsourceibias.n455 gnd 0.010432f
C897 commonsourceibias.t64 gnd 0.150157f
C898 commonsourceibias.n456 gnd 0.059912f
C899 commonsourceibias.n457 gnd 0.010432f
C900 commonsourceibias.n458 gnd 0.008037f
C901 commonsourceibias.n459 gnd 0.008037f
C902 commonsourceibias.n460 gnd 0.008037f
C903 commonsourceibias.n461 gnd 0.007172f
C904 commonsourceibias.n462 gnd 0.011224f
C905 commonsourceibias.n463 gnd 0.059912f
C906 commonsourceibias.n464 gnd 0.011225f
C907 commonsourceibias.n465 gnd 0.008037f
C908 commonsourceibias.n466 gnd 0.008037f
C909 commonsourceibias.n467 gnd 0.008037f
C910 commonsourceibias.n468 gnd 0.009825f
C911 commonsourceibias.n469 gnd 0.059912f
C912 commonsourceibias.n470 gnd 0.010357f
C913 commonsourceibias.t44 gnd 0.150157f
C914 commonsourceibias.n471 gnd 0.059912f
C915 commonsourceibias.n472 gnd 0.010507f
C916 commonsourceibias.n473 gnd 0.008037f
C917 commonsourceibias.n474 gnd 0.008037f
C918 commonsourceibias.n475 gnd 0.008037f
C919 commonsourceibias.n476 gnd 0.007008f
C920 commonsourceibias.n477 gnd 0.011217f
C921 commonsourceibias.n478 gnd 0.059912f
C922 commonsourceibias.n479 gnd 0.01122f
C923 commonsourceibias.n480 gnd 0.008037f
C924 commonsourceibias.n481 gnd 0.008037f
C925 commonsourceibias.n482 gnd 0.008037f
C926 commonsourceibias.n483 gnd 0.009613f
C927 commonsourceibias.n484 gnd 0.059912f
C928 commonsourceibias.n485 gnd 0.010282f
C929 commonsourceibias.t30 gnd 0.150157f
C930 commonsourceibias.n486 gnd 0.059912f
C931 commonsourceibias.n487 gnd 0.010583f
C932 commonsourceibias.n488 gnd 0.008037f
C933 commonsourceibias.n489 gnd 0.008037f
C934 commonsourceibias.n490 gnd 0.008037f
C935 commonsourceibias.n491 gnd 0.006868f
C936 commonsourceibias.n492 gnd 0.011203f
C937 commonsourceibias.n493 gnd 0.059912f
C938 commonsourceibias.n494 gnd 0.01121f
C939 commonsourceibias.n495 gnd 0.008037f
C940 commonsourceibias.n496 gnd 0.008037f
C941 commonsourceibias.n497 gnd 0.008037f
C942 commonsourceibias.n498 gnd 0.009378f
C943 commonsourceibias.n499 gnd 0.059912f
C944 commonsourceibias.n500 gnd 0.009861f
C945 commonsourceibias.t14 gnd 0.162395f
C946 commonsourceibias.n501 gnd 0.07189f
C947 commonsourceibias.n502 gnd 0.080075f
C948 commonsourceibias.t43 gnd 0.017343f
C949 commonsourceibias.t15 gnd 0.017343f
C950 commonsourceibias.n503 gnd 0.15325f
C951 commonsourceibias.n504 gnd 0.132562f
C952 commonsourceibias.t31 gnd 0.017343f
C953 commonsourceibias.t1 gnd 0.017343f
C954 commonsourceibias.n505 gnd 0.15325f
C955 commonsourceibias.n506 gnd 0.070394f
C956 commonsourceibias.t17 gnd 0.017343f
C957 commonsourceibias.t61 gnd 0.017343f
C958 commonsourceibias.n507 gnd 0.15325f
C959 commonsourceibias.n508 gnd 0.070394f
C960 commonsourceibias.t59 gnd 0.017343f
C961 commonsourceibias.t45 gnd 0.017343f
C962 commonsourceibias.n509 gnd 0.15325f
C963 commonsourceibias.n510 gnd 0.070394f
C964 commonsourceibias.t65 gnd 0.017343f
C965 commonsourceibias.t33 gnd 0.017343f
C966 commonsourceibias.n511 gnd 0.15325f
C967 commonsourceibias.n512 gnd 0.058811f
C968 commonsourceibias.n513 gnd 0.071213f
C969 commonsourceibias.n514 gnd 0.052016f
C970 commonsourceibias.t82 gnd 0.150157f
C971 commonsourceibias.n515 gnd 0.059912f
C972 commonsourceibias.n516 gnd 0.008037f
C973 commonsourceibias.t147 gnd 0.150157f
C974 commonsourceibias.n517 gnd 0.059912f
C975 commonsourceibias.n518 gnd 0.008037f
C976 commonsourceibias.t143 gnd 0.150157f
C977 commonsourceibias.n519 gnd 0.059912f
C978 commonsourceibias.n520 gnd 0.008037f
C979 commonsourceibias.t158 gnd 0.150157f
C980 commonsourceibias.n521 gnd 0.007008f
C981 commonsourceibias.n522 gnd 0.008037f
C982 commonsourceibias.t104 gnd 0.150157f
C983 commonsourceibias.n523 gnd 0.009613f
C984 commonsourceibias.n524 gnd 0.008037f
C985 commonsourceibias.t133 gnd 0.150157f
C986 commonsourceibias.n525 gnd 0.006868f
C987 commonsourceibias.n526 gnd 0.008037f
C988 commonsourceibias.t150 gnd 0.150157f
C989 commonsourceibias.n527 gnd 0.009378f
C990 commonsourceibias.t123 gnd 0.166947f
C991 commonsourceibias.t103 gnd 0.150157f
C992 commonsourceibias.n528 gnd 0.065449f
C993 commonsourceibias.n529 gnd 0.071822f
C994 commonsourceibias.n530 gnd 0.033327f
C995 commonsourceibias.n531 gnd 0.008037f
C996 commonsourceibias.n532 gnd 0.007823f
C997 commonsourceibias.n533 gnd 0.01121f
C998 commonsourceibias.n534 gnd 0.059912f
C999 commonsourceibias.n535 gnd 0.011203f
C1000 commonsourceibias.n536 gnd 0.008037f
C1001 commonsourceibias.n537 gnd 0.008037f
C1002 commonsourceibias.n538 gnd 0.008037f
C1003 commonsourceibias.n539 gnd 0.01034f
C1004 commonsourceibias.n540 gnd 0.059912f
C1005 commonsourceibias.n541 gnd 0.010583f
C1006 commonsourceibias.t114 gnd 0.150157f
C1007 commonsourceibias.n542 gnd 0.059912f
C1008 commonsourceibias.n543 gnd 0.010282f
C1009 commonsourceibias.n544 gnd 0.008037f
C1010 commonsourceibias.n545 gnd 0.008037f
C1011 commonsourceibias.n546 gnd 0.008037f
C1012 commonsourceibias.n547 gnd 0.007578f
C1013 commonsourceibias.n548 gnd 0.01122f
C1014 commonsourceibias.n549 gnd 0.059912f
C1015 commonsourceibias.n550 gnd 0.011217f
C1016 commonsourceibias.n551 gnd 0.008037f
C1017 commonsourceibias.n552 gnd 0.008037f
C1018 commonsourceibias.n553 gnd 0.008037f
C1019 commonsourceibias.n554 gnd 0.010186f
C1020 commonsourceibias.n555 gnd 0.059912f
C1021 commonsourceibias.n556 gnd 0.010507f
C1022 commonsourceibias.n557 gnd 0.010357f
C1023 commonsourceibias.n558 gnd 0.008037f
C1024 commonsourceibias.n559 gnd 0.008037f
C1025 commonsourceibias.n560 gnd 0.009825f
C1026 commonsourceibias.n561 gnd 0.007361f
C1027 commonsourceibias.n562 gnd 0.011225f
C1028 commonsourceibias.n563 gnd 0.008037f
C1029 commonsourceibias.n564 gnd 0.008037f
C1030 commonsourceibias.n565 gnd 0.011224f
C1031 commonsourceibias.n566 gnd 0.007172f
C1032 commonsourceibias.n567 gnd 0.010015f
C1033 commonsourceibias.n568 gnd 0.008037f
C1034 commonsourceibias.n569 gnd 0.007021f
C1035 commonsourceibias.n570 gnd 0.010432f
C1036 commonsourceibias.t85 gnd 0.150157f
C1037 commonsourceibias.n571 gnd 0.059912f
C1038 commonsourceibias.n572 gnd 0.010432f
C1039 commonsourceibias.n573 gnd 0.007021f
C1040 commonsourceibias.n574 gnd 0.008037f
C1041 commonsourceibias.n575 gnd 0.008037f
C1042 commonsourceibias.n576 gnd 0.007172f
C1043 commonsourceibias.n577 gnd 0.011224f
C1044 commonsourceibias.n578 gnd 0.059912f
C1045 commonsourceibias.n579 gnd 0.011225f
C1046 commonsourceibias.n580 gnd 0.008037f
C1047 commonsourceibias.n581 gnd 0.008037f
C1048 commonsourceibias.n582 gnd 0.008037f
C1049 commonsourceibias.n583 gnd 0.009825f
C1050 commonsourceibias.n584 gnd 0.059912f
C1051 commonsourceibias.n585 gnd 0.010357f
C1052 commonsourceibias.t89 gnd 0.150157f
C1053 commonsourceibias.n586 gnd 0.059912f
C1054 commonsourceibias.n587 gnd 0.010507f
C1055 commonsourceibias.n588 gnd 0.008037f
C1056 commonsourceibias.n589 gnd 0.008037f
C1057 commonsourceibias.n590 gnd 0.008037f
C1058 commonsourceibias.n591 gnd 0.007008f
C1059 commonsourceibias.n592 gnd 0.011217f
C1060 commonsourceibias.n593 gnd 0.059912f
C1061 commonsourceibias.n594 gnd 0.01122f
C1062 commonsourceibias.n595 gnd 0.008037f
C1063 commonsourceibias.n596 gnd 0.008037f
C1064 commonsourceibias.n597 gnd 0.008037f
C1065 commonsourceibias.n598 gnd 0.009613f
C1066 commonsourceibias.n599 gnd 0.059912f
C1067 commonsourceibias.n600 gnd 0.010282f
C1068 commonsourceibias.t130 gnd 0.150157f
C1069 commonsourceibias.n601 gnd 0.059912f
C1070 commonsourceibias.n602 gnd 0.010583f
C1071 commonsourceibias.n603 gnd 0.008037f
C1072 commonsourceibias.n604 gnd 0.008037f
C1073 commonsourceibias.n605 gnd 0.008037f
C1074 commonsourceibias.n606 gnd 0.006868f
C1075 commonsourceibias.n607 gnd 0.011203f
C1076 commonsourceibias.n608 gnd 0.059912f
C1077 commonsourceibias.n609 gnd 0.01121f
C1078 commonsourceibias.n610 gnd 0.008037f
C1079 commonsourceibias.n611 gnd 0.008037f
C1080 commonsourceibias.n612 gnd 0.008037f
C1081 commonsourceibias.n613 gnd 0.009378f
C1082 commonsourceibias.n614 gnd 0.059912f
C1083 commonsourceibias.n615 gnd 0.009861f
C1084 commonsourceibias.n616 gnd 0.07189f
C1085 commonsourceibias.n617 gnd 0.04697f
C1086 commonsourceibias.n618 gnd 0.010724f
C1087 commonsourceibias.t142 gnd 0.150157f
C1088 commonsourceibias.n619 gnd 0.007823f
C1089 commonsourceibias.n620 gnd 0.008037f
C1090 commonsourceibias.t156 gnd 0.150157f
C1091 commonsourceibias.n621 gnd 0.01034f
C1092 commonsourceibias.n622 gnd 0.008037f
C1093 commonsourceibias.t132 gnd 0.150157f
C1094 commonsourceibias.n623 gnd 0.007578f
C1095 commonsourceibias.n624 gnd 0.008037f
C1096 commonsourceibias.t149 gnd 0.150157f
C1097 commonsourceibias.n625 gnd 0.010186f
C1098 commonsourceibias.n626 gnd 0.008037f
C1099 commonsourceibias.t97 gnd 0.150157f
C1100 commonsourceibias.n627 gnd 0.007361f
C1101 commonsourceibias.n628 gnd 0.008037f
C1102 commonsourceibias.t141 gnd 0.150157f
C1103 commonsourceibias.n629 gnd 0.010015f
C1104 commonsourceibias.n630 gnd 0.008037f
C1105 commonsourceibias.t152 gnd 0.150157f
C1106 commonsourceibias.n631 gnd 0.007172f
C1107 commonsourceibias.n632 gnd 0.008037f
C1108 commonsourceibias.t131 gnd 0.150157f
C1109 commonsourceibias.n633 gnd 0.009825f
C1110 commonsourceibias.n634 gnd 0.008037f
C1111 commonsourceibias.t145 gnd 0.150157f
C1112 commonsourceibias.n635 gnd 0.007008f
C1113 commonsourceibias.n636 gnd 0.008037f
C1114 commonsourceibias.t91 gnd 0.150157f
C1115 commonsourceibias.n637 gnd 0.009613f
C1116 commonsourceibias.n638 gnd 0.008037f
C1117 commonsourceibias.t116 gnd 0.150157f
C1118 commonsourceibias.n639 gnd 0.006868f
C1119 commonsourceibias.n640 gnd 0.008037f
C1120 commonsourceibias.t134 gnd 0.150157f
C1121 commonsourceibias.n641 gnd 0.009378f
C1122 commonsourceibias.t106 gnd 0.166947f
C1123 commonsourceibias.t90 gnd 0.150157f
C1124 commonsourceibias.n642 gnd 0.065449f
C1125 commonsourceibias.n643 gnd 0.071822f
C1126 commonsourceibias.n644 gnd 0.033327f
C1127 commonsourceibias.n645 gnd 0.008037f
C1128 commonsourceibias.n646 gnd 0.007823f
C1129 commonsourceibias.n647 gnd 0.01121f
C1130 commonsourceibias.n648 gnd 0.059912f
C1131 commonsourceibias.n649 gnd 0.011203f
C1132 commonsourceibias.n650 gnd 0.008037f
C1133 commonsourceibias.n651 gnd 0.008037f
C1134 commonsourceibias.n652 gnd 0.008037f
C1135 commonsourceibias.n653 gnd 0.01034f
C1136 commonsourceibias.n654 gnd 0.059912f
C1137 commonsourceibias.n655 gnd 0.010583f
C1138 commonsourceibias.t96 gnd 0.150157f
C1139 commonsourceibias.n656 gnd 0.059912f
C1140 commonsourceibias.n657 gnd 0.010282f
C1141 commonsourceibias.n658 gnd 0.008037f
C1142 commonsourceibias.n659 gnd 0.008037f
C1143 commonsourceibias.n660 gnd 0.008037f
C1144 commonsourceibias.n661 gnd 0.007578f
C1145 commonsourceibias.n662 gnd 0.01122f
C1146 commonsourceibias.n663 gnd 0.059912f
C1147 commonsourceibias.n664 gnd 0.011217f
C1148 commonsourceibias.n665 gnd 0.008037f
C1149 commonsourceibias.n666 gnd 0.008037f
C1150 commonsourceibias.n667 gnd 0.008037f
C1151 commonsourceibias.n668 gnd 0.010186f
C1152 commonsourceibias.n669 gnd 0.059912f
C1153 commonsourceibias.n670 gnd 0.010507f
C1154 commonsourceibias.t124 gnd 0.150157f
C1155 commonsourceibias.n671 gnd 0.059912f
C1156 commonsourceibias.n672 gnd 0.010357f
C1157 commonsourceibias.n673 gnd 0.008037f
C1158 commonsourceibias.n674 gnd 0.008037f
C1159 commonsourceibias.n675 gnd 0.008037f
C1160 commonsourceibias.n676 gnd 0.007361f
C1161 commonsourceibias.n677 gnd 0.011225f
C1162 commonsourceibias.n678 gnd 0.059912f
C1163 commonsourceibias.n679 gnd 0.011224f
C1164 commonsourceibias.n680 gnd 0.008037f
C1165 commonsourceibias.n681 gnd 0.008037f
C1166 commonsourceibias.n682 gnd 0.008037f
C1167 commonsourceibias.n683 gnd 0.010015f
C1168 commonsourceibias.n684 gnd 0.059912f
C1169 commonsourceibias.n685 gnd 0.010432f
C1170 commonsourceibias.t157 gnd 0.150157f
C1171 commonsourceibias.n686 gnd 0.059912f
C1172 commonsourceibias.n687 gnd 0.010432f
C1173 commonsourceibias.n688 gnd 0.008037f
C1174 commonsourceibias.n689 gnd 0.008037f
C1175 commonsourceibias.n690 gnd 0.008037f
C1176 commonsourceibias.n691 gnd 0.007172f
C1177 commonsourceibias.n692 gnd 0.011224f
C1178 commonsourceibias.n693 gnd 0.059912f
C1179 commonsourceibias.n694 gnd 0.011225f
C1180 commonsourceibias.n695 gnd 0.008037f
C1181 commonsourceibias.n696 gnd 0.008037f
C1182 commonsourceibias.n697 gnd 0.008037f
C1183 commonsourceibias.n698 gnd 0.009825f
C1184 commonsourceibias.n699 gnd 0.059912f
C1185 commonsourceibias.n700 gnd 0.010357f
C1186 commonsourceibias.t81 gnd 0.150157f
C1187 commonsourceibias.n701 gnd 0.059912f
C1188 commonsourceibias.n702 gnd 0.010507f
C1189 commonsourceibias.n703 gnd 0.008037f
C1190 commonsourceibias.n704 gnd 0.008037f
C1191 commonsourceibias.n705 gnd 0.008037f
C1192 commonsourceibias.n706 gnd 0.007008f
C1193 commonsourceibias.n707 gnd 0.011217f
C1194 commonsourceibias.n708 gnd 0.059912f
C1195 commonsourceibias.n709 gnd 0.01122f
C1196 commonsourceibias.n710 gnd 0.008037f
C1197 commonsourceibias.n711 gnd 0.008037f
C1198 commonsourceibias.n712 gnd 0.008037f
C1199 commonsourceibias.n713 gnd 0.009613f
C1200 commonsourceibias.n714 gnd 0.059912f
C1201 commonsourceibias.n715 gnd 0.010282f
C1202 commonsourceibias.t111 gnd 0.150157f
C1203 commonsourceibias.n716 gnd 0.059912f
C1204 commonsourceibias.n717 gnd 0.010583f
C1205 commonsourceibias.n718 gnd 0.008037f
C1206 commonsourceibias.n719 gnd 0.008037f
C1207 commonsourceibias.n720 gnd 0.008037f
C1208 commonsourceibias.n721 gnd 0.006868f
C1209 commonsourceibias.n722 gnd 0.011203f
C1210 commonsourceibias.n723 gnd 0.059912f
C1211 commonsourceibias.n724 gnd 0.01121f
C1212 commonsourceibias.n725 gnd 0.008037f
C1213 commonsourceibias.n726 gnd 0.008037f
C1214 commonsourceibias.n727 gnd 0.008037f
C1215 commonsourceibias.n728 gnd 0.009378f
C1216 commonsourceibias.n729 gnd 0.059912f
C1217 commonsourceibias.n730 gnd 0.009861f
C1218 commonsourceibias.t122 gnd 0.162395f
C1219 commonsourceibias.n731 gnd 0.07189f
C1220 commonsourceibias.n732 gnd 0.025003f
C1221 commonsourceibias.n733 gnd 0.221951f
C1222 commonsourceibias.n734 gnd 4.85761f
C1223 diffpairibias.t27 gnd 0.090128f
C1224 diffpairibias.t23 gnd 0.08996f
C1225 diffpairibias.n0 gnd 0.105991f
C1226 diffpairibias.t28 gnd 0.08996f
C1227 diffpairibias.n1 gnd 0.051736f
C1228 diffpairibias.t25 gnd 0.08996f
C1229 diffpairibias.n2 gnd 0.051736f
C1230 diffpairibias.t29 gnd 0.08996f
C1231 diffpairibias.n3 gnd 0.041084f
C1232 diffpairibias.t15 gnd 0.086371f
C1233 diffpairibias.t1 gnd 0.085993f
C1234 diffpairibias.n4 gnd 0.13579f
C1235 diffpairibias.t11 gnd 0.085993f
C1236 diffpairibias.n5 gnd 0.072463f
C1237 diffpairibias.t13 gnd 0.085993f
C1238 diffpairibias.n6 gnd 0.072463f
C1239 diffpairibias.t7 gnd 0.085993f
C1240 diffpairibias.n7 gnd 0.072463f
C1241 diffpairibias.t3 gnd 0.085993f
C1242 diffpairibias.n8 gnd 0.072463f
C1243 diffpairibias.t17 gnd 0.085993f
C1244 diffpairibias.n9 gnd 0.072463f
C1245 diffpairibias.t5 gnd 0.085993f
C1246 diffpairibias.n10 gnd 0.072463f
C1247 diffpairibias.t19 gnd 0.085993f
C1248 diffpairibias.n11 gnd 0.072463f
C1249 diffpairibias.t9 gnd 0.085993f
C1250 diffpairibias.n12 gnd 0.102883f
C1251 diffpairibias.t14 gnd 0.086899f
C1252 diffpairibias.t0 gnd 0.086748f
C1253 diffpairibias.n13 gnd 0.094648f
C1254 diffpairibias.t10 gnd 0.086748f
C1255 diffpairibias.n14 gnd 0.052262f
C1256 diffpairibias.t12 gnd 0.086748f
C1257 diffpairibias.n15 gnd 0.052262f
C1258 diffpairibias.t6 gnd 0.086748f
C1259 diffpairibias.n16 gnd 0.052262f
C1260 diffpairibias.t2 gnd 0.086748f
C1261 diffpairibias.n17 gnd 0.052262f
C1262 diffpairibias.t16 gnd 0.086748f
C1263 diffpairibias.n18 gnd 0.052262f
C1264 diffpairibias.t4 gnd 0.086748f
C1265 diffpairibias.n19 gnd 0.052262f
C1266 diffpairibias.t18 gnd 0.086748f
C1267 diffpairibias.n20 gnd 0.052262f
C1268 diffpairibias.t8 gnd 0.086748f
C1269 diffpairibias.n21 gnd 0.061849f
C1270 diffpairibias.n22 gnd 0.233513f
C1271 diffpairibias.t20 gnd 0.08996f
C1272 diffpairibias.n23 gnd 0.051747f
C1273 diffpairibias.t26 gnd 0.08996f
C1274 diffpairibias.n24 gnd 0.051736f
C1275 diffpairibias.t22 gnd 0.08996f
C1276 diffpairibias.n25 gnd 0.051736f
C1277 diffpairibias.t21 gnd 0.08996f
C1278 diffpairibias.n26 gnd 0.051736f
C1279 diffpairibias.t24 gnd 0.08996f
C1280 diffpairibias.n27 gnd 0.04729f
C1281 diffpairibias.n28 gnd 0.047711f
C1282 outputibias.t10 gnd 0.11477f
C1283 outputibias.t8 gnd 0.115567f
C1284 outputibias.n0 gnd 0.130108f
C1285 outputibias.n1 gnd 0.001372f
C1286 outputibias.n2 gnd 9.76e-19
C1287 outputibias.n3 gnd 5.24e-19
C1288 outputibias.n4 gnd 0.001239f
C1289 outputibias.n5 gnd 5.55e-19
C1290 outputibias.n6 gnd 9.76e-19
C1291 outputibias.n7 gnd 5.24e-19
C1292 outputibias.n8 gnd 0.001239f
C1293 outputibias.n9 gnd 5.55e-19
C1294 outputibias.n10 gnd 0.004176f
C1295 outputibias.t5 gnd 0.00202f
C1296 outputibias.n11 gnd 9.3e-19
C1297 outputibias.n12 gnd 7.32e-19
C1298 outputibias.n13 gnd 5.24e-19
C1299 outputibias.n14 gnd 0.02322f
C1300 outputibias.n15 gnd 9.76e-19
C1301 outputibias.n16 gnd 5.24e-19
C1302 outputibias.n17 gnd 5.55e-19
C1303 outputibias.n18 gnd 0.001239f
C1304 outputibias.n19 gnd 0.001239f
C1305 outputibias.n20 gnd 5.55e-19
C1306 outputibias.n21 gnd 5.24e-19
C1307 outputibias.n22 gnd 9.76e-19
C1308 outputibias.n23 gnd 9.76e-19
C1309 outputibias.n24 gnd 5.24e-19
C1310 outputibias.n25 gnd 5.55e-19
C1311 outputibias.n26 gnd 0.001239f
C1312 outputibias.n27 gnd 0.002683f
C1313 outputibias.n28 gnd 5.55e-19
C1314 outputibias.n29 gnd 5.24e-19
C1315 outputibias.n30 gnd 0.002256f
C1316 outputibias.n31 gnd 0.005781f
C1317 outputibias.n32 gnd 0.001372f
C1318 outputibias.n33 gnd 9.76e-19
C1319 outputibias.n34 gnd 5.24e-19
C1320 outputibias.n35 gnd 0.001239f
C1321 outputibias.n36 gnd 5.55e-19
C1322 outputibias.n37 gnd 9.76e-19
C1323 outputibias.n38 gnd 5.24e-19
C1324 outputibias.n39 gnd 0.001239f
C1325 outputibias.n40 gnd 5.55e-19
C1326 outputibias.n41 gnd 0.004176f
C1327 outputibias.t3 gnd 0.00202f
C1328 outputibias.n42 gnd 9.3e-19
C1329 outputibias.n43 gnd 7.32e-19
C1330 outputibias.n44 gnd 5.24e-19
C1331 outputibias.n45 gnd 0.02322f
C1332 outputibias.n46 gnd 9.76e-19
C1333 outputibias.n47 gnd 5.24e-19
C1334 outputibias.n48 gnd 5.55e-19
C1335 outputibias.n49 gnd 0.001239f
C1336 outputibias.n50 gnd 0.001239f
C1337 outputibias.n51 gnd 5.55e-19
C1338 outputibias.n52 gnd 5.24e-19
C1339 outputibias.n53 gnd 9.76e-19
C1340 outputibias.n54 gnd 9.76e-19
C1341 outputibias.n55 gnd 5.24e-19
C1342 outputibias.n56 gnd 5.55e-19
C1343 outputibias.n57 gnd 0.001239f
C1344 outputibias.n58 gnd 0.002683f
C1345 outputibias.n59 gnd 5.55e-19
C1346 outputibias.n60 gnd 5.24e-19
C1347 outputibias.n61 gnd 0.002256f
C1348 outputibias.n62 gnd 0.005197f
C1349 outputibias.n63 gnd 0.121892f
C1350 outputibias.n64 gnd 0.001372f
C1351 outputibias.n65 gnd 9.76e-19
C1352 outputibias.n66 gnd 5.24e-19
C1353 outputibias.n67 gnd 0.001239f
C1354 outputibias.n68 gnd 5.55e-19
C1355 outputibias.n69 gnd 9.76e-19
C1356 outputibias.n70 gnd 5.24e-19
C1357 outputibias.n71 gnd 0.001239f
C1358 outputibias.n72 gnd 5.55e-19
C1359 outputibias.n73 gnd 0.004176f
C1360 outputibias.t1 gnd 0.00202f
C1361 outputibias.n74 gnd 9.3e-19
C1362 outputibias.n75 gnd 7.32e-19
C1363 outputibias.n76 gnd 5.24e-19
C1364 outputibias.n77 gnd 0.02322f
C1365 outputibias.n78 gnd 9.76e-19
C1366 outputibias.n79 gnd 5.24e-19
C1367 outputibias.n80 gnd 5.55e-19
C1368 outputibias.n81 gnd 0.001239f
C1369 outputibias.n82 gnd 0.001239f
C1370 outputibias.n83 gnd 5.55e-19
C1371 outputibias.n84 gnd 5.24e-19
C1372 outputibias.n85 gnd 9.76e-19
C1373 outputibias.n86 gnd 9.76e-19
C1374 outputibias.n87 gnd 5.24e-19
C1375 outputibias.n88 gnd 5.55e-19
C1376 outputibias.n89 gnd 0.001239f
C1377 outputibias.n90 gnd 0.002683f
C1378 outputibias.n91 gnd 5.55e-19
C1379 outputibias.n92 gnd 5.24e-19
C1380 outputibias.n93 gnd 0.002256f
C1381 outputibias.n94 gnd 0.005197f
C1382 outputibias.n95 gnd 0.064513f
C1383 outputibias.n96 gnd 0.001372f
C1384 outputibias.n97 gnd 9.76e-19
C1385 outputibias.n98 gnd 5.24e-19
C1386 outputibias.n99 gnd 0.001239f
C1387 outputibias.n100 gnd 5.55e-19
C1388 outputibias.n101 gnd 9.76e-19
C1389 outputibias.n102 gnd 5.24e-19
C1390 outputibias.n103 gnd 0.001239f
C1391 outputibias.n104 gnd 5.55e-19
C1392 outputibias.n105 gnd 0.004176f
C1393 outputibias.t7 gnd 0.00202f
C1394 outputibias.n106 gnd 9.3e-19
C1395 outputibias.n107 gnd 7.32e-19
C1396 outputibias.n108 gnd 5.24e-19
C1397 outputibias.n109 gnd 0.02322f
C1398 outputibias.n110 gnd 9.76e-19
C1399 outputibias.n111 gnd 5.24e-19
C1400 outputibias.n112 gnd 5.55e-19
C1401 outputibias.n113 gnd 0.001239f
C1402 outputibias.n114 gnd 0.001239f
C1403 outputibias.n115 gnd 5.55e-19
C1404 outputibias.n116 gnd 5.24e-19
C1405 outputibias.n117 gnd 9.76e-19
C1406 outputibias.n118 gnd 9.76e-19
C1407 outputibias.n119 gnd 5.24e-19
C1408 outputibias.n120 gnd 5.55e-19
C1409 outputibias.n121 gnd 0.001239f
C1410 outputibias.n122 gnd 0.002683f
C1411 outputibias.n123 gnd 5.55e-19
C1412 outputibias.n124 gnd 5.24e-19
C1413 outputibias.n125 gnd 0.002256f
C1414 outputibias.n126 gnd 0.005197f
C1415 outputibias.n127 gnd 0.084814f
C1416 outputibias.t6 gnd 0.108319f
C1417 outputibias.t0 gnd 0.108319f
C1418 outputibias.t2 gnd 0.108319f
C1419 outputibias.t4 gnd 0.109238f
C1420 outputibias.n128 gnd 0.134674f
C1421 outputibias.n129 gnd 0.07244f
C1422 outputibias.n130 gnd 0.079818f
C1423 outputibias.n131 gnd 0.164901f
C1424 outputibias.t11 gnd 0.11477f
C1425 outputibias.n132 gnd 0.067481f
C1426 outputibias.t9 gnd 0.11477f
C1427 outputibias.n133 gnd 0.065115f
C1428 outputibias.n134 gnd 0.029159f
C1429 a_n1808_13878.t17 gnd 0.185195f
C1430 a_n1808_13878.t15 gnd 0.185195f
C1431 a_n1808_13878.t19 gnd 0.185195f
C1432 a_n1808_13878.n0 gnd 1.46067f
C1433 a_n1808_13878.t8 gnd 0.185195f
C1434 a_n1808_13878.t13 gnd 0.185195f
C1435 a_n1808_13878.n1 gnd 1.45825f
C1436 a_n1808_13878.n2 gnd 1.31079f
C1437 a_n1808_13878.t10 gnd 0.185195f
C1438 a_n1808_13878.t12 gnd 0.185195f
C1439 a_n1808_13878.n3 gnd 1.4598f
C1440 a_n1808_13878.t16 gnd 0.185195f
C1441 a_n1808_13878.t11 gnd 0.185195f
C1442 a_n1808_13878.n4 gnd 1.45825f
C1443 a_n1808_13878.n5 gnd 2.03762f
C1444 a_n1808_13878.t14 gnd 0.185195f
C1445 a_n1808_13878.t9 gnd 0.185195f
C1446 a_n1808_13878.n6 gnd 1.45825f
C1447 a_n1808_13878.n7 gnd 3.69301f
C1448 a_n1808_13878.t1 gnd 1.73408f
C1449 a_n1808_13878.t4 gnd 0.185195f
C1450 a_n1808_13878.t5 gnd 0.185195f
C1451 a_n1808_13878.n8 gnd 1.30452f
C1452 a_n1808_13878.n9 gnd 1.4576f
C1453 a_n1808_13878.t0 gnd 1.73062f
C1454 a_n1808_13878.n10 gnd 0.733487f
C1455 a_n1808_13878.t3 gnd 1.73062f
C1456 a_n1808_13878.n11 gnd 0.733487f
C1457 a_n1808_13878.t6 gnd 0.185195f
C1458 a_n1808_13878.t7 gnd 0.185195f
C1459 a_n1808_13878.n12 gnd 1.30452f
C1460 a_n1808_13878.n13 gnd 0.74059f
C1461 a_n1808_13878.t2 gnd 1.73062f
C1462 a_n1808_13878.n14 gnd 1.7272f
C1463 a_n1808_13878.n15 gnd 2.51438f
C1464 a_n1808_13878.n16 gnd 1.80025f
C1465 a_n1808_13878.n17 gnd 1.45826f
C1466 a_n1808_13878.t18 gnd 0.185195f
C1467 a_n1996_n452.n0 gnd 0.822727f
C1468 a_n1996_n452.n1 gnd 3.34433f
C1469 a_n1996_n452.n2 gnd 3.17111f
C1470 a_n1996_n452.n3 gnd 3.91594f
C1471 a_n1996_n452.n4 gnd 0.527811f
C1472 a_n1996_n452.n5 gnd 0.205584f
C1473 a_n1996_n452.n6 gnd 0.151417f
C1474 a_n1996_n452.n7 gnd 0.237979f
C1475 a_n1996_n452.n8 gnd 0.183812f
C1476 a_n1996_n452.n9 gnd 0.205584f
C1477 a_n1996_n452.n10 gnd 1.00969f
C1478 a_n1996_n452.n11 gnd 0.151417f
C1479 a_n1996_n452.n12 gnd 0.581979f
C1480 a_n1996_n452.n13 gnd 0.433746f
C1481 a_n1996_n452.n14 gnd 0.21667f
C1482 a_n1996_n452.n15 gnd 0.494132f
C1483 a_n1996_n452.n16 gnd 0.283464f
C1484 a_n1996_n452.n17 gnd 0.439964f
C1485 a_n1996_n452.n18 gnd 0.21667f
C1486 a_n1996_n452.n19 gnd 0.734001f
C1487 a_n1996_n452.n20 gnd 0.283464f
C1488 a_n1996_n452.n21 gnd 0.494132f
C1489 a_n1996_n452.n22 gnd 0.666675f
C1490 a_n1996_n452.n23 gnd 0.21667f
C1491 a_n1996_n452.n24 gnd 0.283464f
C1492 a_n1996_n452.n25 gnd 0.641354f
C1493 a_n1996_n452.n26 gnd 0.283464f
C1494 a_n1996_n452.n27 gnd 1.18284f
C1495 a_n1996_n452.n28 gnd 1.92214f
C1496 a_n1996_n452.n29 gnd 1.14844f
C1497 a_n1996_n452.n30 gnd 1.78382f
C1498 a_n1996_n452.n31 gnd 3.22512f
C1499 a_n1996_n452.n32 gnd 0.108335f
C1500 a_n1996_n452.n33 gnd 0.008389f
C1501 a_n1996_n452.n35 gnd 0.008389f
C1502 a_n1996_n452.n37 gnd 0.286629f
C1503 a_n1996_n452.n38 gnd 0.008389f
C1504 a_n1996_n452.n40 gnd 0.286629f
C1505 a_n1996_n452.n41 gnd 0.008389f
C1506 a_n1996_n452.n43 gnd 0.286629f
C1507 a_n1996_n452.n44 gnd 0.008389f
C1508 a_n1996_n452.n45 gnd 0.286221f
C1509 a_n1996_n452.n46 gnd 0.008389f
C1510 a_n1996_n452.n47 gnd 0.286221f
C1511 a_n1996_n452.n48 gnd 0.008389f
C1512 a_n1996_n452.n49 gnd 0.286221f
C1513 a_n1996_n452.n50 gnd 0.008389f
C1514 a_n1996_n452.n51 gnd 0.286221f
C1515 a_n1996_n452.n52 gnd 0.286629f
C1516 a_n1996_n452.t34 gnd 0.150285f
C1517 a_n1996_n452.t21 gnd 0.713776f
C1518 a_n1996_n452.t19 gnd 0.699053f
C1519 a_n1996_n452.t33 gnd 0.699053f
C1520 a_n1996_n452.t29 gnd 0.699053f
C1521 a_n1996_n452.n53 gnd 0.307348f
C1522 a_n1996_n452.t31 gnd 0.710611f
C1523 a_n1996_n452.t16 gnd 0.116888f
C1524 a_n1996_n452.t6 gnd 0.116888f
C1525 a_n1996_n452.n54 gnd 1.03516f
C1526 a_n1996_n452.t8 gnd 0.116888f
C1527 a_n1996_n452.t5 gnd 0.116888f
C1528 a_n1996_n452.n55 gnd 1.03287f
C1529 a_n1996_n452.t18 gnd 0.116888f
C1530 a_n1996_n452.t15 gnd 0.116888f
C1531 a_n1996_n452.n56 gnd 1.03287f
C1532 a_n1996_n452.t3 gnd 0.116888f
C1533 a_n1996_n452.t4 gnd 0.116888f
C1534 a_n1996_n452.n57 gnd 1.03516f
C1535 a_n1996_n452.t9 gnd 0.116888f
C1536 a_n1996_n452.t0 gnd 0.116888f
C1537 a_n1996_n452.n58 gnd 1.03287f
C1538 a_n1996_n452.t43 gnd 0.116888f
C1539 a_n1996_n452.t7 gnd 0.116888f
C1540 a_n1996_n452.n59 gnd 1.03287f
C1541 a_n1996_n452.t14 gnd 0.116888f
C1542 a_n1996_n452.t11 gnd 0.116888f
C1543 a_n1996_n452.n60 gnd 1.03287f
C1544 a_n1996_n452.t1 gnd 0.116888f
C1545 a_n1996_n452.t17 gnd 0.116888f
C1546 a_n1996_n452.n61 gnd 1.03287f
C1547 a_n1996_n452.t13 gnd 0.116888f
C1548 a_n1996_n452.t12 gnd 0.116888f
C1549 a_n1996_n452.n62 gnd 1.03516f
C1550 a_n1996_n452.t10 gnd 0.116888f
C1551 a_n1996_n452.t2 gnd 0.116888f
C1552 a_n1996_n452.n63 gnd 1.03287f
C1553 a_n1996_n452.t70 gnd 0.713776f
C1554 a_n1996_n452.t53 gnd 0.699053f
C1555 a_n1996_n452.t57 gnd 0.699053f
C1556 a_n1996_n452.t47 gnd 0.699053f
C1557 a_n1996_n452.n64 gnd 0.307348f
C1558 a_n1996_n452.t62 gnd 0.699053f
C1559 a_n1996_n452.t68 gnd 0.710611f
C1560 a_n1996_n452.t24 gnd 1.40719f
C1561 a_n1996_n452.t38 gnd 0.150285f
C1562 a_n1996_n452.t42 gnd 0.150285f
C1563 a_n1996_n452.n65 gnd 1.05861f
C1564 a_n1996_n452.t36 gnd 0.150285f
C1565 a_n1996_n452.t40 gnd 0.150285f
C1566 a_n1996_n452.n66 gnd 1.05861f
C1567 a_n1996_n452.t28 gnd 1.40439f
C1568 a_n1996_n452.t35 gnd 0.699053f
C1569 a_n1996_n452.n67 gnd 0.307348f
C1570 a_n1996_n452.t39 gnd 0.699053f
C1571 a_n1996_n452.t37 gnd 0.699053f
C1572 a_n1996_n452.t52 gnd 0.699053f
C1573 a_n1996_n452.n68 gnd 0.307348f
C1574 a_n1996_n452.t61 gnd 0.699053f
C1575 a_n1996_n452.t66 gnd 0.699053f
C1576 a_n1996_n452.t65 gnd 0.713776f
C1577 a_n1996_n452.n69 gnd 0.309974f
C1578 a_n1996_n452.t45 gnd 0.699053f
C1579 a_n1996_n452.n70 gnd 0.303445f
C1580 a_n1996_n452.n71 gnd 0.309974f
C1581 a_n1996_n452.t46 gnd 0.710611f
C1582 a_n1996_n452.t23 gnd 0.713776f
C1583 a_n1996_n452.n72 gnd 0.309974f
C1584 a_n1996_n452.t41 gnd 0.699053f
C1585 a_n1996_n452.n73 gnd 0.303445f
C1586 a_n1996_n452.n74 gnd 0.309974f
C1587 a_n1996_n452.t27 gnd 0.710611f
C1588 a_n1996_n452.n75 gnd 1.13585f
C1589 a_n1996_n452.t50 gnd 0.699053f
C1590 a_n1996_n452.n76 gnd 0.303445f
C1591 a_n1996_n452.t56 gnd 0.699053f
C1592 a_n1996_n452.n77 gnd 0.303445f
C1593 a_n1996_n452.t48 gnd 0.699053f
C1594 a_n1996_n452.n78 gnd 0.303445f
C1595 a_n1996_n452.t60 gnd 0.699053f
C1596 a_n1996_n452.n79 gnd 0.303445f
C1597 a_n1996_n452.t51 gnd 0.699053f
C1598 a_n1996_n452.n80 gnd 0.297934f
C1599 a_n1996_n452.t71 gnd 0.699053f
C1600 a_n1996_n452.n81 gnd 0.307348f
C1601 a_n1996_n452.t54 gnd 0.710766f
C1602 a_n1996_n452.t63 gnd 0.699053f
C1603 a_n1996_n452.n82 gnd 0.297934f
C1604 a_n1996_n452.t49 gnd 0.699053f
C1605 a_n1996_n452.n83 gnd 0.307348f
C1606 a_n1996_n452.t58 gnd 0.710766f
C1607 a_n1996_n452.t67 gnd 0.699053f
C1608 a_n1996_n452.n84 gnd 0.297934f
C1609 a_n1996_n452.t55 gnd 0.699053f
C1610 a_n1996_n452.n85 gnd 0.307348f
C1611 a_n1996_n452.t69 gnd 0.710766f
C1612 a_n1996_n452.t59 gnd 0.699053f
C1613 a_n1996_n452.n86 gnd 0.297934f
C1614 a_n1996_n452.t44 gnd 0.699053f
C1615 a_n1996_n452.n87 gnd 0.307348f
C1616 a_n1996_n452.t64 gnd 0.710766f
C1617 a_n1996_n452.n88 gnd 1.34296f
C1618 a_n1996_n452.n89 gnd 0.309974f
C1619 a_n1996_n452.n90 gnd 0.303445f
C1620 a_n1996_n452.n91 gnd 0.309974f
C1621 a_n1996_n452.t25 gnd 0.699053f
C1622 a_n1996_n452.n92 gnd 0.309974f
C1623 a_n1996_n452.n93 gnd 0.303445f
C1624 a_n1996_n452.n94 gnd 0.309974f
C1625 a_n1996_n452.n95 gnd 0.789588f
C1626 a_n1996_n452.t22 gnd 1.40439f
C1627 a_n1996_n452.t32 gnd 1.40719f
C1628 a_n1996_n452.t30 gnd 0.150285f
C1629 a_n1996_n452.t26 gnd 0.150285f
C1630 a_n1996_n452.n96 gnd 1.05861f
C1631 a_n1996_n452.n97 gnd 1.05861f
C1632 a_n1996_n452.t20 gnd 0.150285f
C1633 CSoutput.n0 gnd 0.044617f
C1634 CSoutput.t193 gnd 0.295134f
C1635 CSoutput.n1 gnd 0.133268f
C1636 CSoutput.n2 gnd 0.044617f
C1637 CSoutput.t176 gnd 0.295134f
C1638 CSoutput.n3 gnd 0.035363f
C1639 CSoutput.n4 gnd 0.044617f
C1640 CSoutput.t185 gnd 0.295134f
C1641 CSoutput.n5 gnd 0.030494f
C1642 CSoutput.n6 gnd 0.044617f
C1643 CSoutput.t196 gnd 0.295134f
C1644 CSoutput.t195 gnd 0.295134f
C1645 CSoutput.n7 gnd 0.131815f
C1646 CSoutput.n8 gnd 0.044617f
C1647 CSoutput.t182 gnd 0.295134f
C1648 CSoutput.n9 gnd 0.029074f
C1649 CSoutput.n10 gnd 0.044617f
C1650 CSoutput.t188 gnd 0.295134f
C1651 CSoutput.t191 gnd 0.295134f
C1652 CSoutput.n11 gnd 0.131815f
C1653 CSoutput.n12 gnd 0.044617f
C1654 CSoutput.t179 gnd 0.295134f
C1655 CSoutput.n13 gnd 0.030494f
C1656 CSoutput.n14 gnd 0.044617f
C1657 CSoutput.t178 gnd 0.295134f
C1658 CSoutput.t189 gnd 0.295134f
C1659 CSoutput.n15 gnd 0.131815f
C1660 CSoutput.n16 gnd 0.044617f
C1661 CSoutput.t194 gnd 0.295134f
C1662 CSoutput.n17 gnd 0.032569f
C1663 CSoutput.t180 gnd 0.352693f
C1664 CSoutput.t177 gnd 0.295134f
C1665 CSoutput.n18 gnd 0.168277f
C1666 CSoutput.n19 gnd 0.163287f
C1667 CSoutput.n20 gnd 0.189432f
C1668 CSoutput.n21 gnd 0.044617f
C1669 CSoutput.n22 gnd 0.037238f
C1670 CSoutput.n23 gnd 0.131815f
C1671 CSoutput.n24 gnd 0.035896f
C1672 CSoutput.n25 gnd 0.035363f
C1673 CSoutput.n26 gnd 0.044617f
C1674 CSoutput.n27 gnd 0.044617f
C1675 CSoutput.n28 gnd 0.036952f
C1676 CSoutput.n29 gnd 0.031373f
C1677 CSoutput.n30 gnd 0.13475f
C1678 CSoutput.n31 gnd 0.031805f
C1679 CSoutput.n32 gnd 0.044617f
C1680 CSoutput.n33 gnd 0.044617f
C1681 CSoutput.n34 gnd 0.044617f
C1682 CSoutput.n35 gnd 0.036558f
C1683 CSoutput.n36 gnd 0.131815f
C1684 CSoutput.n37 gnd 0.034963f
C1685 CSoutput.n38 gnd 0.036297f
C1686 CSoutput.n39 gnd 0.044617f
C1687 CSoutput.n40 gnd 0.044617f
C1688 CSoutput.n41 gnd 0.03723f
C1689 CSoutput.n42 gnd 0.034029f
C1690 CSoutput.n43 gnd 0.131815f
C1691 CSoutput.n44 gnd 0.034891f
C1692 CSoutput.n45 gnd 0.044617f
C1693 CSoutput.n46 gnd 0.044617f
C1694 CSoutput.n47 gnd 0.044617f
C1695 CSoutput.n48 gnd 0.034891f
C1696 CSoutput.n49 gnd 0.131815f
C1697 CSoutput.n50 gnd 0.034029f
C1698 CSoutput.n51 gnd 0.03723f
C1699 CSoutput.n52 gnd 0.044617f
C1700 CSoutput.n53 gnd 0.044617f
C1701 CSoutput.n54 gnd 0.036297f
C1702 CSoutput.n55 gnd 0.034963f
C1703 CSoutput.n56 gnd 0.131815f
C1704 CSoutput.n57 gnd 0.036558f
C1705 CSoutput.n58 gnd 0.044617f
C1706 CSoutput.n59 gnd 0.044617f
C1707 CSoutput.n60 gnd 0.044617f
C1708 CSoutput.n61 gnd 0.031805f
C1709 CSoutput.n62 gnd 0.13475f
C1710 CSoutput.n63 gnd 0.031373f
C1711 CSoutput.t197 gnd 0.295134f
C1712 CSoutput.n64 gnd 0.131815f
C1713 CSoutput.n65 gnd 0.036952f
C1714 CSoutput.n66 gnd 0.044617f
C1715 CSoutput.n67 gnd 0.044617f
C1716 CSoutput.n68 gnd 0.044617f
C1717 CSoutput.n69 gnd 0.035896f
C1718 CSoutput.n70 gnd 0.131815f
C1719 CSoutput.n71 gnd 0.037238f
C1720 CSoutput.n72 gnd 0.032569f
C1721 CSoutput.n73 gnd 0.044617f
C1722 CSoutput.n74 gnd 0.044617f
C1723 CSoutput.n75 gnd 0.033776f
C1724 CSoutput.n76 gnd 0.02006f
C1725 CSoutput.t183 gnd 0.331604f
C1726 CSoutput.n77 gnd 0.164727f
C1727 CSoutput.n78 gnd 0.704854f
C1728 CSoutput.t128 gnd 0.055654f
C1729 CSoutput.t48 gnd 0.055654f
C1730 CSoutput.n79 gnd 0.43089f
C1731 CSoutput.t111 gnd 0.055654f
C1732 CSoutput.t88 gnd 0.055654f
C1733 CSoutput.n80 gnd 0.430122f
C1734 CSoutput.n81 gnd 0.436573f
C1735 CSoutput.t118 gnd 0.055654f
C1736 CSoutput.t68 gnd 0.055654f
C1737 CSoutput.n82 gnd 0.430122f
C1738 CSoutput.n83 gnd 0.215125f
C1739 CSoutput.t135 gnd 0.055654f
C1740 CSoutput.t82 gnd 0.055654f
C1741 CSoutput.n84 gnd 0.430122f
C1742 CSoutput.n85 gnd 0.215125f
C1743 CSoutput.t53 gnd 0.055654f
C1744 CSoutput.t96 gnd 0.055654f
C1745 CSoutput.n86 gnd 0.430122f
C1746 CSoutput.n87 gnd 0.215125f
C1747 CSoutput.t57 gnd 0.055654f
C1748 CSoutput.t76 gnd 0.055654f
C1749 CSoutput.n88 gnd 0.430122f
C1750 CSoutput.n89 gnd 0.215125f
C1751 CSoutput.t140 gnd 0.055654f
C1752 CSoutput.t90 gnd 0.055654f
C1753 CSoutput.n90 gnd 0.430122f
C1754 CSoutput.n91 gnd 0.215125f
C1755 CSoutput.t60 gnd 0.055654f
C1756 CSoutput.t124 gnd 0.055654f
C1757 CSoutput.n92 gnd 0.430122f
C1758 CSoutput.n93 gnd 0.394489f
C1759 CSoutput.t122 gnd 0.055654f
C1760 CSoutput.t120 gnd 0.055654f
C1761 CSoutput.n94 gnd 0.43089f
C1762 CSoutput.t105 gnd 0.055654f
C1763 CSoutput.t54 gnd 0.055654f
C1764 CSoutput.n95 gnd 0.430122f
C1765 CSoutput.n96 gnd 0.436573f
C1766 CSoutput.t49 gnd 0.055654f
C1767 CSoutput.t116 gnd 0.055654f
C1768 CSoutput.n97 gnd 0.430122f
C1769 CSoutput.n98 gnd 0.215125f
C1770 CSoutput.t104 gnd 0.055654f
C1771 CSoutput.t84 gnd 0.055654f
C1772 CSoutput.n99 gnd 0.430122f
C1773 CSoutput.n100 gnd 0.215125f
C1774 CSoutput.t69 gnd 0.055654f
C1775 CSoutput.t131 gnd 0.055654f
C1776 CSoutput.n101 gnd 0.430122f
C1777 CSoutput.n102 gnd 0.215125f
C1778 CSoutput.t103 gnd 0.055654f
C1779 CSoutput.t102 gnd 0.055654f
C1780 CSoutput.n103 gnd 0.430122f
C1781 CSoutput.n104 gnd 0.215125f
C1782 CSoutput.t93 gnd 0.055654f
C1783 CSoutput.t65 gnd 0.055654f
C1784 CSoutput.n105 gnd 0.430122f
C1785 CSoutput.n106 gnd 0.215125f
C1786 CSoutput.t52 gnd 0.055654f
C1787 CSoutput.t94 gnd 0.055654f
C1788 CSoutput.n107 gnd 0.430122f
C1789 CSoutput.n108 gnd 0.320805f
C1790 CSoutput.n109 gnd 0.404533f
C1791 CSoutput.t133 gnd 0.055654f
C1792 CSoutput.t132 gnd 0.055654f
C1793 CSoutput.n110 gnd 0.43089f
C1794 CSoutput.t114 gnd 0.055654f
C1795 CSoutput.t64 gnd 0.055654f
C1796 CSoutput.n111 gnd 0.430122f
C1797 CSoutput.n112 gnd 0.436573f
C1798 CSoutput.t61 gnd 0.055654f
C1799 CSoutput.t130 gnd 0.055654f
C1800 CSoutput.n113 gnd 0.430122f
C1801 CSoutput.n114 gnd 0.215125f
C1802 CSoutput.t112 gnd 0.055654f
C1803 CSoutput.t95 gnd 0.055654f
C1804 CSoutput.n115 gnd 0.430122f
C1805 CSoutput.n116 gnd 0.215125f
C1806 CSoutput.t78 gnd 0.055654f
C1807 CSoutput.t141 gnd 0.055654f
C1808 CSoutput.n117 gnd 0.430122f
C1809 CSoutput.n118 gnd 0.215125f
C1810 CSoutput.t110 gnd 0.055654f
C1811 CSoutput.t109 gnd 0.055654f
C1812 CSoutput.n119 gnd 0.430122f
C1813 CSoutput.n120 gnd 0.215125f
C1814 CSoutput.t100 gnd 0.055654f
C1815 CSoutput.t77 gnd 0.055654f
C1816 CSoutput.n121 gnd 0.430122f
C1817 CSoutput.n122 gnd 0.215125f
C1818 CSoutput.t63 gnd 0.055654f
C1819 CSoutput.t101 gnd 0.055654f
C1820 CSoutput.n123 gnd 0.430122f
C1821 CSoutput.n124 gnd 0.320805f
C1822 CSoutput.n125 gnd 0.452165f
C1823 CSoutput.n126 gnd 9.338679f
C1824 CSoutput.n128 gnd 0.789272f
C1825 CSoutput.n129 gnd 0.591954f
C1826 CSoutput.n130 gnd 0.789272f
C1827 CSoutput.n131 gnd 0.789272f
C1828 CSoutput.n132 gnd 2.12496f
C1829 CSoutput.n133 gnd 0.789272f
C1830 CSoutput.n134 gnd 0.789272f
C1831 CSoutput.t187 gnd 0.98659f
C1832 CSoutput.n135 gnd 0.789272f
C1833 CSoutput.n136 gnd 0.789272f
C1834 CSoutput.n140 gnd 0.789272f
C1835 CSoutput.n144 gnd 0.789272f
C1836 CSoutput.n145 gnd 0.789272f
C1837 CSoutput.n147 gnd 0.789272f
C1838 CSoutput.n152 gnd 0.789272f
C1839 CSoutput.n154 gnd 0.789272f
C1840 CSoutput.n155 gnd 0.789272f
C1841 CSoutput.n157 gnd 0.789272f
C1842 CSoutput.n158 gnd 0.789272f
C1843 CSoutput.n160 gnd 0.789272f
C1844 CSoutput.t181 gnd 13.1886f
C1845 CSoutput.n162 gnd 0.789272f
C1846 CSoutput.n163 gnd 0.591954f
C1847 CSoutput.n164 gnd 0.789272f
C1848 CSoutput.n165 gnd 0.789272f
C1849 CSoutput.n166 gnd 2.12496f
C1850 CSoutput.n167 gnd 0.789272f
C1851 CSoutput.n168 gnd 0.789272f
C1852 CSoutput.t184 gnd 0.98659f
C1853 CSoutput.n169 gnd 0.789272f
C1854 CSoutput.n170 gnd 0.789272f
C1855 CSoutput.n174 gnd 0.789272f
C1856 CSoutput.n178 gnd 0.789272f
C1857 CSoutput.n179 gnd 0.789272f
C1858 CSoutput.n181 gnd 0.789272f
C1859 CSoutput.n186 gnd 0.789272f
C1860 CSoutput.n188 gnd 0.789272f
C1861 CSoutput.n189 gnd 0.789272f
C1862 CSoutput.n191 gnd 0.789272f
C1863 CSoutput.n192 gnd 0.789272f
C1864 CSoutput.n194 gnd 0.789272f
C1865 CSoutput.n195 gnd 0.591954f
C1866 CSoutput.n197 gnd 0.789272f
C1867 CSoutput.n198 gnd 0.591954f
C1868 CSoutput.n199 gnd 0.789272f
C1869 CSoutput.n200 gnd 0.789272f
C1870 CSoutput.n201 gnd 2.12496f
C1871 CSoutput.n202 gnd 0.789272f
C1872 CSoutput.n203 gnd 0.789272f
C1873 CSoutput.t186 gnd 0.98659f
C1874 CSoutput.n204 gnd 0.789272f
C1875 CSoutput.n205 gnd 2.12496f
C1876 CSoutput.n207 gnd 0.789272f
C1877 CSoutput.n208 gnd 0.789272f
C1878 CSoutput.n210 gnd 0.789272f
C1879 CSoutput.n211 gnd 0.789272f
C1880 CSoutput.t192 gnd 12.973701f
C1881 CSoutput.t190 gnd 13.1886f
C1882 CSoutput.n217 gnd 2.47606f
C1883 CSoutput.n218 gnd 10.086599f
C1884 CSoutput.n219 gnd 10.5086f
C1885 CSoutput.n224 gnd 2.68224f
C1886 CSoutput.n230 gnd 0.789272f
C1887 CSoutput.n232 gnd 0.789272f
C1888 CSoutput.n234 gnd 0.789272f
C1889 CSoutput.n236 gnd 0.789272f
C1890 CSoutput.n238 gnd 0.789272f
C1891 CSoutput.n244 gnd 0.789272f
C1892 CSoutput.n251 gnd 1.44801f
C1893 CSoutput.n252 gnd 1.44801f
C1894 CSoutput.n253 gnd 0.789272f
C1895 CSoutput.n254 gnd 0.789272f
C1896 CSoutput.n256 gnd 0.591954f
C1897 CSoutput.n257 gnd 0.506956f
C1898 CSoutput.n259 gnd 0.591954f
C1899 CSoutput.n260 gnd 0.506956f
C1900 CSoutput.n261 gnd 0.591954f
C1901 CSoutput.n263 gnd 0.789272f
C1902 CSoutput.n265 gnd 2.12496f
C1903 CSoutput.n266 gnd 2.47606f
C1904 CSoutput.n267 gnd 9.27706f
C1905 CSoutput.n269 gnd 0.591954f
C1906 CSoutput.n270 gnd 1.52313f
C1907 CSoutput.n271 gnd 0.591954f
C1908 CSoutput.n273 gnd 0.789272f
C1909 CSoutput.n275 gnd 2.12496f
C1910 CSoutput.n276 gnd 4.62851f
C1911 CSoutput.t47 gnd 0.055654f
C1912 CSoutput.t127 gnd 0.055654f
C1913 CSoutput.n277 gnd 0.43089f
C1914 CSoutput.t87 gnd 0.055654f
C1915 CSoutput.t139 gnd 0.055654f
C1916 CSoutput.n278 gnd 0.430122f
C1917 CSoutput.n279 gnd 0.436573f
C1918 CSoutput.t67 gnd 0.055654f
C1919 CSoutput.t117 gnd 0.055654f
C1920 CSoutput.n280 gnd 0.430122f
C1921 CSoutput.n281 gnd 0.215125f
C1922 CSoutput.t81 gnd 0.055654f
C1923 CSoutput.t134 gnd 0.055654f
C1924 CSoutput.n282 gnd 0.430122f
C1925 CSoutput.n283 gnd 0.215125f
C1926 CSoutput.t113 gnd 0.055654f
C1927 CSoutput.t51 gnd 0.055654f
C1928 CSoutput.n284 gnd 0.430122f
C1929 CSoutput.n285 gnd 0.215125f
C1930 CSoutput.t75 gnd 0.055654f
C1931 CSoutput.t56 gnd 0.055654f
C1932 CSoutput.n286 gnd 0.430122f
C1933 CSoutput.n287 gnd 0.215125f
C1934 CSoutput.t89 gnd 0.055654f
C1935 CSoutput.t72 gnd 0.055654f
C1936 CSoutput.n288 gnd 0.430122f
C1937 CSoutput.n289 gnd 0.215125f
C1938 CSoutput.t123 gnd 0.055654f
C1939 CSoutput.t59 gnd 0.055654f
C1940 CSoutput.n290 gnd 0.430122f
C1941 CSoutput.n291 gnd 0.394489f
C1942 CSoutput.t91 gnd 0.055654f
C1943 CSoutput.t92 gnd 0.055654f
C1944 CSoutput.n292 gnd 0.43089f
C1945 CSoutput.t108 gnd 0.055654f
C1946 CSoutput.t50 gnd 0.055654f
C1947 CSoutput.n293 gnd 0.430122f
C1948 CSoutput.n294 gnd 0.436573f
C1949 CSoutput.t86 gnd 0.055654f
C1950 CSoutput.t106 gnd 0.055654f
C1951 CSoutput.n295 gnd 0.430122f
C1952 CSoutput.n296 gnd 0.215125f
C1953 CSoutput.t46 gnd 0.055654f
C1954 CSoutput.t73 gnd 0.055654f
C1955 CSoutput.n297 gnd 0.430122f
C1956 CSoutput.n298 gnd 0.215125f
C1957 CSoutput.t74 gnd 0.055654f
C1958 CSoutput.t129 gnd 0.055654f
C1959 CSoutput.n299 gnd 0.430122f
C1960 CSoutput.n300 gnd 0.215125f
C1961 CSoutput.t70 gnd 0.055654f
C1962 CSoutput.t71 gnd 0.055654f
C1963 CSoutput.n301 gnd 0.430122f
C1964 CSoutput.n302 gnd 0.215125f
C1965 CSoutput.t125 gnd 0.055654f
C1966 CSoutput.t126 gnd 0.055654f
C1967 CSoutput.n303 gnd 0.430122f
C1968 CSoutput.n304 gnd 0.215125f
C1969 CSoutput.t55 gnd 0.055654f
C1970 CSoutput.t107 gnd 0.055654f
C1971 CSoutput.n305 gnd 0.430122f
C1972 CSoutput.n306 gnd 0.320805f
C1973 CSoutput.n307 gnd 0.404533f
C1974 CSoutput.t98 gnd 0.055654f
C1975 CSoutput.t99 gnd 0.055654f
C1976 CSoutput.n308 gnd 0.43089f
C1977 CSoutput.t121 gnd 0.055654f
C1978 CSoutput.t62 gnd 0.055654f
C1979 CSoutput.n309 gnd 0.430122f
C1980 CSoutput.n310 gnd 0.436573f
C1981 CSoutput.t97 gnd 0.055654f
C1982 CSoutput.t115 gnd 0.055654f
C1983 CSoutput.n311 gnd 0.430122f
C1984 CSoutput.n312 gnd 0.215125f
C1985 CSoutput.t58 gnd 0.055654f
C1986 CSoutput.t83 gnd 0.055654f
C1987 CSoutput.n313 gnd 0.430122f
C1988 CSoutput.n314 gnd 0.215125f
C1989 CSoutput.t85 gnd 0.055654f
C1990 CSoutput.t138 gnd 0.055654f
C1991 CSoutput.n315 gnd 0.430122f
C1992 CSoutput.n316 gnd 0.215125f
C1993 CSoutput.t79 gnd 0.055654f
C1994 CSoutput.t80 gnd 0.055654f
C1995 CSoutput.n317 gnd 0.430122f
C1996 CSoutput.n318 gnd 0.215125f
C1997 CSoutput.t136 gnd 0.055654f
C1998 CSoutput.t137 gnd 0.055654f
C1999 CSoutput.n319 gnd 0.430122f
C2000 CSoutput.n320 gnd 0.215125f
C2001 CSoutput.t66 gnd 0.055654f
C2002 CSoutput.t119 gnd 0.055654f
C2003 CSoutput.n321 gnd 0.43012f
C2004 CSoutput.n322 gnd 0.320807f
C2005 CSoutput.n323 gnd 0.452165f
C2006 CSoutput.n324 gnd 12.8735f
C2007 CSoutput.t7 gnd 0.048697f
C2008 CSoutput.t17 gnd 0.048697f
C2009 CSoutput.n325 gnd 0.431745f
C2010 CSoutput.t33 gnd 0.048697f
C2011 CSoutput.t32 gnd 0.048697f
C2012 CSoutput.n326 gnd 0.430304f
C2013 CSoutput.n327 gnd 0.400963f
C2014 CSoutput.t167 gnd 0.048697f
C2015 CSoutput.t153 gnd 0.048697f
C2016 CSoutput.n328 gnd 0.430304f
C2017 CSoutput.n329 gnd 0.197656f
C2018 CSoutput.t23 gnd 0.048697f
C2019 CSoutput.t11 gnd 0.048697f
C2020 CSoutput.n330 gnd 0.430304f
C2021 CSoutput.n331 gnd 0.197656f
C2022 CSoutput.t21 gnd 0.048697f
C2023 CSoutput.t4 gnd 0.048697f
C2024 CSoutput.n332 gnd 0.430304f
C2025 CSoutput.n333 gnd 0.197656f
C2026 CSoutput.t149 gnd 0.048697f
C2027 CSoutput.t168 gnd 0.048697f
C2028 CSoutput.n334 gnd 0.430304f
C2029 CSoutput.n335 gnd 0.197656f
C2030 CSoutput.t145 gnd 0.048697f
C2031 CSoutput.t44 gnd 0.048697f
C2032 CSoutput.n336 gnd 0.430304f
C2033 CSoutput.n337 gnd 0.197656f
C2034 CSoutput.t160 gnd 0.048697f
C2035 CSoutput.t148 gnd 0.048697f
C2036 CSoutput.n338 gnd 0.430304f
C2037 CSoutput.n339 gnd 0.197656f
C2038 CSoutput.t166 gnd 0.048697f
C2039 CSoutput.t175 gnd 0.048697f
C2040 CSoutput.n340 gnd 0.430304f
C2041 CSoutput.n341 gnd 0.197656f
C2042 CSoutput.t24 gnd 0.048697f
C2043 CSoutput.t31 gnd 0.048697f
C2044 CSoutput.n342 gnd 0.430304f
C2045 CSoutput.n343 gnd 0.364518f
C2046 CSoutput.t173 gnd 0.048697f
C2047 CSoutput.t146 gnd 0.048697f
C2048 CSoutput.n344 gnd 0.431745f
C2049 CSoutput.t20 gnd 0.048697f
C2050 CSoutput.t169 gnd 0.048697f
C2051 CSoutput.n345 gnd 0.430304f
C2052 CSoutput.n346 gnd 0.400963f
C2053 CSoutput.t147 gnd 0.048697f
C2054 CSoutput.t162 gnd 0.048697f
C2055 CSoutput.n347 gnd 0.430304f
C2056 CSoutput.n348 gnd 0.197656f
C2057 CSoutput.t25 gnd 0.048697f
C2058 CSoutput.t152 gnd 0.048697f
C2059 CSoutput.n349 gnd 0.430304f
C2060 CSoutput.n350 gnd 0.197656f
C2061 CSoutput.t39 gnd 0.048697f
C2062 CSoutput.t16 gnd 0.048697f
C2063 CSoutput.n351 gnd 0.430304f
C2064 CSoutput.n352 gnd 0.197656f
C2065 CSoutput.t3 gnd 0.048697f
C2066 CSoutput.t5 gnd 0.048697f
C2067 CSoutput.n353 gnd 0.430304f
C2068 CSoutput.n354 gnd 0.197656f
C2069 CSoutput.t8 gnd 0.048697f
C2070 CSoutput.t38 gnd 0.048697f
C2071 CSoutput.n355 gnd 0.430304f
C2072 CSoutput.n356 gnd 0.197656f
C2073 CSoutput.t12 gnd 0.048697f
C2074 CSoutput.t170 gnd 0.048697f
C2075 CSoutput.n357 gnd 0.430304f
C2076 CSoutput.n358 gnd 0.197656f
C2077 CSoutput.t10 gnd 0.048697f
C2078 CSoutput.t165 gnd 0.048697f
C2079 CSoutput.n359 gnd 0.430304f
C2080 CSoutput.n360 gnd 0.197656f
C2081 CSoutput.t26 gnd 0.048697f
C2082 CSoutput.t174 gnd 0.048697f
C2083 CSoutput.n361 gnd 0.430304f
C2084 CSoutput.n362 gnd 0.300084f
C2085 CSoutput.n363 gnd 0.557579f
C2086 CSoutput.n364 gnd 13.9417f
C2087 CSoutput.t29 gnd 0.048697f
C2088 CSoutput.t45 gnd 0.048697f
C2089 CSoutput.n365 gnd 0.431745f
C2090 CSoutput.t164 gnd 0.048697f
C2091 CSoutput.t158 gnd 0.048697f
C2092 CSoutput.n366 gnd 0.430304f
C2093 CSoutput.n367 gnd 0.400963f
C2094 CSoutput.t27 gnd 0.048697f
C2095 CSoutput.t42 gnd 0.048697f
C2096 CSoutput.n368 gnd 0.430304f
C2097 CSoutput.n369 gnd 0.197656f
C2098 CSoutput.t40 gnd 0.048697f
C2099 CSoutput.t150 gnd 0.048697f
C2100 CSoutput.n370 gnd 0.430304f
C2101 CSoutput.n371 gnd 0.197656f
C2102 CSoutput.t159 gnd 0.048697f
C2103 CSoutput.t14 gnd 0.048697f
C2104 CSoutput.n372 gnd 0.430304f
C2105 CSoutput.n373 gnd 0.197656f
C2106 CSoutput.t142 gnd 0.048697f
C2107 CSoutput.t151 gnd 0.048697f
C2108 CSoutput.n374 gnd 0.430304f
C2109 CSoutput.n375 gnd 0.197656f
C2110 CSoutput.t13 gnd 0.048697f
C2111 CSoutput.t154 gnd 0.048697f
C2112 CSoutput.n376 gnd 0.430304f
C2113 CSoutput.n377 gnd 0.197656f
C2114 CSoutput.t172 gnd 0.048697f
C2115 CSoutput.t144 gnd 0.048697f
C2116 CSoutput.n378 gnd 0.430304f
C2117 CSoutput.n379 gnd 0.197656f
C2118 CSoutput.t15 gnd 0.048697f
C2119 CSoutput.t22 gnd 0.048697f
C2120 CSoutput.n380 gnd 0.430304f
C2121 CSoutput.n381 gnd 0.197656f
C2122 CSoutput.t36 gnd 0.048697f
C2123 CSoutput.t9 gnd 0.048697f
C2124 CSoutput.n382 gnd 0.430304f
C2125 CSoutput.n383 gnd 0.364518f
C2126 CSoutput.t155 gnd 0.048697f
C2127 CSoutput.t37 gnd 0.048697f
C2128 CSoutput.n384 gnd 0.431745f
C2129 CSoutput.t0 gnd 0.048697f
C2130 CSoutput.t6 gnd 0.048697f
C2131 CSoutput.n385 gnd 0.430304f
C2132 CSoutput.n386 gnd 0.400963f
C2133 CSoutput.t34 gnd 0.048697f
C2134 CSoutput.t163 gnd 0.048697f
C2135 CSoutput.n387 gnd 0.430304f
C2136 CSoutput.n388 gnd 0.197656f
C2137 CSoutput.t2 gnd 0.048697f
C2138 CSoutput.t28 gnd 0.048697f
C2139 CSoutput.n389 gnd 0.430304f
C2140 CSoutput.n390 gnd 0.197656f
C2141 CSoutput.t19 gnd 0.048697f
C2142 CSoutput.t41 gnd 0.048697f
C2143 CSoutput.n391 gnd 0.430304f
C2144 CSoutput.n392 gnd 0.197656f
C2145 CSoutput.t43 gnd 0.048697f
C2146 CSoutput.t30 gnd 0.048697f
C2147 CSoutput.n393 gnd 0.430304f
C2148 CSoutput.n394 gnd 0.197656f
C2149 CSoutput.t171 gnd 0.048697f
C2150 CSoutput.t35 gnd 0.048697f
C2151 CSoutput.n395 gnd 0.430304f
C2152 CSoutput.n396 gnd 0.197656f
C2153 CSoutput.t1 gnd 0.048697f
C2154 CSoutput.t157 gnd 0.048697f
C2155 CSoutput.n397 gnd 0.430304f
C2156 CSoutput.n398 gnd 0.197656f
C2157 CSoutput.t18 gnd 0.048697f
C2158 CSoutput.t143 gnd 0.048697f
C2159 CSoutput.n399 gnd 0.430304f
C2160 CSoutput.n400 gnd 0.197656f
C2161 CSoutput.t161 gnd 0.048697f
C2162 CSoutput.t156 gnd 0.048697f
C2163 CSoutput.n401 gnd 0.430304f
C2164 CSoutput.n402 gnd 0.300084f
C2165 CSoutput.n403 gnd 0.557579f
C2166 CSoutput.n404 gnd 8.42525f
C2167 CSoutput.n405 gnd 14.623501f
C2168 vdd.t259 gnd 0.038369f
C2169 vdd.t102 gnd 0.038369f
C2170 vdd.n0 gnd 0.302625f
C2171 vdd.t3 gnd 0.038369f
C2172 vdd.t5 gnd 0.038369f
C2173 vdd.n1 gnd 0.302125f
C2174 vdd.n2 gnd 0.278617f
C2175 vdd.t116 gnd 0.038369f
C2176 vdd.t257 gnd 0.038369f
C2177 vdd.n3 gnd 0.302125f
C2178 vdd.n4 gnd 0.140907f
C2179 vdd.t110 gnd 0.038369f
C2180 vdd.t14 gnd 0.038369f
C2181 vdd.n5 gnd 0.302125f
C2182 vdd.n6 gnd 0.132215f
C2183 vdd.t118 gnd 0.038369f
C2184 vdd.t122 gnd 0.038369f
C2185 vdd.n7 gnd 0.302625f
C2186 vdd.t11 gnd 0.038369f
C2187 vdd.t104 gnd 0.038369f
C2188 vdd.n8 gnd 0.302125f
C2189 vdd.n9 gnd 0.278617f
C2190 vdd.t261 gnd 0.038369f
C2191 vdd.t120 gnd 0.038369f
C2192 vdd.n10 gnd 0.302125f
C2193 vdd.n11 gnd 0.140907f
C2194 vdd.t263 gnd 0.038369f
C2195 vdd.t107 gnd 0.038369f
C2196 vdd.n12 gnd 0.302125f
C2197 vdd.n13 gnd 0.132215f
C2198 vdd.n14 gnd 0.093474f
C2199 vdd.t114 gnd 0.021316f
C2200 vdd.t126 gnd 0.021316f
C2201 vdd.n15 gnd 0.196207f
C2202 vdd.t18 gnd 0.021316f
C2203 vdd.t123 gnd 0.021316f
C2204 vdd.n16 gnd 0.195633f
C2205 vdd.n17 gnd 0.340462f
C2206 vdd.t17 gnd 0.021316f
C2207 vdd.t127 gnd 0.021316f
C2208 vdd.n18 gnd 0.195633f
C2209 vdd.n19 gnd 0.140854f
C2210 vdd.t21 gnd 0.021316f
C2211 vdd.t124 gnd 0.021316f
C2212 vdd.n20 gnd 0.196207f
C2213 vdd.t15 gnd 0.021316f
C2214 vdd.t112 gnd 0.021316f
C2215 vdd.n21 gnd 0.195633f
C2216 vdd.n22 gnd 0.340462f
C2217 vdd.t19 gnd 0.021316f
C2218 vdd.t20 gnd 0.021316f
C2219 vdd.n23 gnd 0.195633f
C2220 vdd.n24 gnd 0.140854f
C2221 vdd.t113 gnd 0.021316f
C2222 vdd.t111 gnd 0.021316f
C2223 vdd.n25 gnd 0.195633f
C2224 vdd.t125 gnd 0.021316f
C2225 vdd.t16 gnd 0.021316f
C2226 vdd.n26 gnd 0.195633f
C2227 vdd.n27 gnd 22.976099f
C2228 vdd.n28 gnd 8.6566f
C2229 vdd.n29 gnd 0.005814f
C2230 vdd.n30 gnd 0.005395f
C2231 vdd.n31 gnd 0.002984f
C2232 vdd.n32 gnd 0.006852f
C2233 vdd.n33 gnd 0.002899f
C2234 vdd.n34 gnd 0.00307f
C2235 vdd.n35 gnd 0.005395f
C2236 vdd.n36 gnd 0.002899f
C2237 vdd.n37 gnd 0.006852f
C2238 vdd.n38 gnd 0.00307f
C2239 vdd.n39 gnd 0.005395f
C2240 vdd.n40 gnd 0.002899f
C2241 vdd.n41 gnd 0.005139f
C2242 vdd.n42 gnd 0.005155f
C2243 vdd.t135 gnd 0.014721f
C2244 vdd.n43 gnd 0.032755f
C2245 vdd.n44 gnd 0.170464f
C2246 vdd.n45 gnd 0.002899f
C2247 vdd.n46 gnd 0.00307f
C2248 vdd.n47 gnd 0.006852f
C2249 vdd.n48 gnd 0.006852f
C2250 vdd.n49 gnd 0.00307f
C2251 vdd.n50 gnd 0.002899f
C2252 vdd.n51 gnd 0.005395f
C2253 vdd.n52 gnd 0.005395f
C2254 vdd.n53 gnd 0.002899f
C2255 vdd.n54 gnd 0.00307f
C2256 vdd.n55 gnd 0.006852f
C2257 vdd.n56 gnd 0.006852f
C2258 vdd.n57 gnd 0.00307f
C2259 vdd.n58 gnd 0.002899f
C2260 vdd.n59 gnd 0.005395f
C2261 vdd.n60 gnd 0.005395f
C2262 vdd.n61 gnd 0.002899f
C2263 vdd.n62 gnd 0.00307f
C2264 vdd.n63 gnd 0.006852f
C2265 vdd.n64 gnd 0.006852f
C2266 vdd.n65 gnd 0.0162f
C2267 vdd.n66 gnd 0.002984f
C2268 vdd.n67 gnd 0.002899f
C2269 vdd.n68 gnd 0.013944f
C2270 vdd.n69 gnd 0.009735f
C2271 vdd.t242 gnd 0.034106f
C2272 vdd.t192 gnd 0.034106f
C2273 vdd.n70 gnd 0.2344f
C2274 vdd.n71 gnd 0.18432f
C2275 vdd.t253 gnd 0.034106f
C2276 vdd.t164 gnd 0.034106f
C2277 vdd.n72 gnd 0.2344f
C2278 vdd.n73 gnd 0.148745f
C2279 vdd.t231 gnd 0.034106f
C2280 vdd.t184 gnd 0.034106f
C2281 vdd.n74 gnd 0.2344f
C2282 vdd.n75 gnd 0.148745f
C2283 vdd.t248 gnd 0.034106f
C2284 vdd.t226 gnd 0.034106f
C2285 vdd.n76 gnd 0.2344f
C2286 vdd.n77 gnd 0.148745f
C2287 vdd.t133 gnd 0.034106f
C2288 vdd.t177 gnd 0.034106f
C2289 vdd.n78 gnd 0.2344f
C2290 vdd.n79 gnd 0.148745f
C2291 vdd.t149 gnd 0.034106f
C2292 vdd.t195 gnd 0.034106f
C2293 vdd.n80 gnd 0.2344f
C2294 vdd.n81 gnd 0.148745f
C2295 vdd.t172 gnd 0.034106f
C2296 vdd.t238 gnd 0.034106f
C2297 vdd.n82 gnd 0.2344f
C2298 vdd.n83 gnd 0.148745f
C2299 vdd.n84 gnd 0.005814f
C2300 vdd.n85 gnd 0.005395f
C2301 vdd.n86 gnd 0.002984f
C2302 vdd.n87 gnd 0.006852f
C2303 vdd.n88 gnd 0.002899f
C2304 vdd.n89 gnd 0.00307f
C2305 vdd.n90 gnd 0.005395f
C2306 vdd.n91 gnd 0.002899f
C2307 vdd.n92 gnd 0.006852f
C2308 vdd.n93 gnd 0.00307f
C2309 vdd.n94 gnd 0.005395f
C2310 vdd.n95 gnd 0.002899f
C2311 vdd.n96 gnd 0.005139f
C2312 vdd.n97 gnd 0.005155f
C2313 vdd.t154 gnd 0.014721f
C2314 vdd.n98 gnd 0.032755f
C2315 vdd.n99 gnd 0.170464f
C2316 vdd.n100 gnd 0.002899f
C2317 vdd.n101 gnd 0.00307f
C2318 vdd.n102 gnd 0.006852f
C2319 vdd.n103 gnd 0.006852f
C2320 vdd.n104 gnd 0.00307f
C2321 vdd.n105 gnd 0.002899f
C2322 vdd.n106 gnd 0.005395f
C2323 vdd.n107 gnd 0.005395f
C2324 vdd.n108 gnd 0.002899f
C2325 vdd.n109 gnd 0.00307f
C2326 vdd.n110 gnd 0.006852f
C2327 vdd.n111 gnd 0.006852f
C2328 vdd.n112 gnd 0.00307f
C2329 vdd.n113 gnd 0.002899f
C2330 vdd.n114 gnd 0.005395f
C2331 vdd.n115 gnd 0.005395f
C2332 vdd.n116 gnd 0.002899f
C2333 vdd.n117 gnd 0.00307f
C2334 vdd.n118 gnd 0.006852f
C2335 vdd.n119 gnd 0.006852f
C2336 vdd.n120 gnd 0.0162f
C2337 vdd.n121 gnd 0.002984f
C2338 vdd.n122 gnd 0.002899f
C2339 vdd.n123 gnd 0.013944f
C2340 vdd.n124 gnd 0.00943f
C2341 vdd.n125 gnd 0.110667f
C2342 vdd.n126 gnd 0.005814f
C2343 vdd.n127 gnd 0.005395f
C2344 vdd.n128 gnd 0.002984f
C2345 vdd.n129 gnd 0.006852f
C2346 vdd.n130 gnd 0.002899f
C2347 vdd.n131 gnd 0.00307f
C2348 vdd.n132 gnd 0.005395f
C2349 vdd.n133 gnd 0.002899f
C2350 vdd.n134 gnd 0.006852f
C2351 vdd.n135 gnd 0.00307f
C2352 vdd.n136 gnd 0.005395f
C2353 vdd.n137 gnd 0.002899f
C2354 vdd.n138 gnd 0.005139f
C2355 vdd.n139 gnd 0.005155f
C2356 vdd.t197 gnd 0.014721f
C2357 vdd.n140 gnd 0.032755f
C2358 vdd.n141 gnd 0.170464f
C2359 vdd.n142 gnd 0.002899f
C2360 vdd.n143 gnd 0.00307f
C2361 vdd.n144 gnd 0.006852f
C2362 vdd.n145 gnd 0.006852f
C2363 vdd.n146 gnd 0.00307f
C2364 vdd.n147 gnd 0.002899f
C2365 vdd.n148 gnd 0.005395f
C2366 vdd.n149 gnd 0.005395f
C2367 vdd.n150 gnd 0.002899f
C2368 vdd.n151 gnd 0.00307f
C2369 vdd.n152 gnd 0.006852f
C2370 vdd.n153 gnd 0.006852f
C2371 vdd.n154 gnd 0.00307f
C2372 vdd.n155 gnd 0.002899f
C2373 vdd.n156 gnd 0.005395f
C2374 vdd.n157 gnd 0.005395f
C2375 vdd.n158 gnd 0.002899f
C2376 vdd.n159 gnd 0.00307f
C2377 vdd.n160 gnd 0.006852f
C2378 vdd.n161 gnd 0.006852f
C2379 vdd.n162 gnd 0.0162f
C2380 vdd.n163 gnd 0.002984f
C2381 vdd.n164 gnd 0.002899f
C2382 vdd.n165 gnd 0.013944f
C2383 vdd.n166 gnd 0.009735f
C2384 vdd.t199 gnd 0.034106f
C2385 vdd.t221 gnd 0.034106f
C2386 vdd.n167 gnd 0.2344f
C2387 vdd.n168 gnd 0.18432f
C2388 vdd.t131 gnd 0.034106f
C2389 vdd.t185 gnd 0.034106f
C2390 vdd.n169 gnd 0.2344f
C2391 vdd.n170 gnd 0.148745f
C2392 vdd.t219 gnd 0.034106f
C2393 vdd.t129 gnd 0.034106f
C2394 vdd.n171 gnd 0.2344f
C2395 vdd.n172 gnd 0.148745f
C2396 vdd.t174 gnd 0.034106f
C2397 vdd.t176 gnd 0.034106f
C2398 vdd.n173 gnd 0.2344f
C2399 vdd.n174 gnd 0.148745f
C2400 vdd.t227 gnd 0.034106f
C2401 vdd.t169 gnd 0.034106f
C2402 vdd.n175 gnd 0.2344f
C2403 vdd.n176 gnd 0.148745f
C2404 vdd.t170 gnd 0.034106f
C2405 vdd.t240 gnd 0.034106f
C2406 vdd.n177 gnd 0.2344f
C2407 vdd.n178 gnd 0.148745f
C2408 vdd.t241 gnd 0.034106f
C2409 vdd.t147 gnd 0.034106f
C2410 vdd.n179 gnd 0.2344f
C2411 vdd.n180 gnd 0.148745f
C2412 vdd.n181 gnd 0.005814f
C2413 vdd.n182 gnd 0.005395f
C2414 vdd.n183 gnd 0.002984f
C2415 vdd.n184 gnd 0.006852f
C2416 vdd.n185 gnd 0.002899f
C2417 vdd.n186 gnd 0.00307f
C2418 vdd.n187 gnd 0.005395f
C2419 vdd.n188 gnd 0.002899f
C2420 vdd.n189 gnd 0.006852f
C2421 vdd.n190 gnd 0.00307f
C2422 vdd.n191 gnd 0.005395f
C2423 vdd.n192 gnd 0.002899f
C2424 vdd.n193 gnd 0.005139f
C2425 vdd.n194 gnd 0.005155f
C2426 vdd.t220 gnd 0.014721f
C2427 vdd.n195 gnd 0.032755f
C2428 vdd.n196 gnd 0.170464f
C2429 vdd.n197 gnd 0.002899f
C2430 vdd.n198 gnd 0.00307f
C2431 vdd.n199 gnd 0.006852f
C2432 vdd.n200 gnd 0.006852f
C2433 vdd.n201 gnd 0.00307f
C2434 vdd.n202 gnd 0.002899f
C2435 vdd.n203 gnd 0.005395f
C2436 vdd.n204 gnd 0.005395f
C2437 vdd.n205 gnd 0.002899f
C2438 vdd.n206 gnd 0.00307f
C2439 vdd.n207 gnd 0.006852f
C2440 vdd.n208 gnd 0.006852f
C2441 vdd.n209 gnd 0.00307f
C2442 vdd.n210 gnd 0.002899f
C2443 vdd.n211 gnd 0.005395f
C2444 vdd.n212 gnd 0.005395f
C2445 vdd.n213 gnd 0.002899f
C2446 vdd.n214 gnd 0.00307f
C2447 vdd.n215 gnd 0.006852f
C2448 vdd.n216 gnd 0.006852f
C2449 vdd.n217 gnd 0.0162f
C2450 vdd.n218 gnd 0.002984f
C2451 vdd.n219 gnd 0.002899f
C2452 vdd.n220 gnd 0.013944f
C2453 vdd.n221 gnd 0.00943f
C2454 vdd.n222 gnd 0.065836f
C2455 vdd.n223 gnd 0.237223f
C2456 vdd.n224 gnd 0.005814f
C2457 vdd.n225 gnd 0.005395f
C2458 vdd.n226 gnd 0.002984f
C2459 vdd.n227 gnd 0.006852f
C2460 vdd.n228 gnd 0.002899f
C2461 vdd.n229 gnd 0.00307f
C2462 vdd.n230 gnd 0.005395f
C2463 vdd.n231 gnd 0.002899f
C2464 vdd.n232 gnd 0.006852f
C2465 vdd.n233 gnd 0.00307f
C2466 vdd.n234 gnd 0.005395f
C2467 vdd.n235 gnd 0.002899f
C2468 vdd.n236 gnd 0.005139f
C2469 vdd.n237 gnd 0.005155f
C2470 vdd.t205 gnd 0.014721f
C2471 vdd.n238 gnd 0.032755f
C2472 vdd.n239 gnd 0.170464f
C2473 vdd.n240 gnd 0.002899f
C2474 vdd.n241 gnd 0.00307f
C2475 vdd.n242 gnd 0.006852f
C2476 vdd.n243 gnd 0.006852f
C2477 vdd.n244 gnd 0.00307f
C2478 vdd.n245 gnd 0.002899f
C2479 vdd.n246 gnd 0.005395f
C2480 vdd.n247 gnd 0.005395f
C2481 vdd.n248 gnd 0.002899f
C2482 vdd.n249 gnd 0.00307f
C2483 vdd.n250 gnd 0.006852f
C2484 vdd.n251 gnd 0.006852f
C2485 vdd.n252 gnd 0.00307f
C2486 vdd.n253 gnd 0.002899f
C2487 vdd.n254 gnd 0.005395f
C2488 vdd.n255 gnd 0.005395f
C2489 vdd.n256 gnd 0.002899f
C2490 vdd.n257 gnd 0.00307f
C2491 vdd.n258 gnd 0.006852f
C2492 vdd.n259 gnd 0.006852f
C2493 vdd.n260 gnd 0.0162f
C2494 vdd.n261 gnd 0.002984f
C2495 vdd.n262 gnd 0.002899f
C2496 vdd.n263 gnd 0.013944f
C2497 vdd.n264 gnd 0.009735f
C2498 vdd.t209 gnd 0.034106f
C2499 vdd.t235 gnd 0.034106f
C2500 vdd.n265 gnd 0.2344f
C2501 vdd.n266 gnd 0.18432f
C2502 vdd.t157 gnd 0.034106f
C2503 vdd.t208 gnd 0.034106f
C2504 vdd.n267 gnd 0.2344f
C2505 vdd.n268 gnd 0.148745f
C2506 vdd.t230 gnd 0.034106f
C2507 vdd.t152 gnd 0.034106f
C2508 vdd.n269 gnd 0.2344f
C2509 vdd.n270 gnd 0.148745f
C2510 vdd.t188 gnd 0.034106f
C2511 vdd.t190 gnd 0.034106f
C2512 vdd.n271 gnd 0.2344f
C2513 vdd.n272 gnd 0.148745f
C2514 vdd.t252 gnd 0.034106f
C2515 vdd.t182 gnd 0.034106f
C2516 vdd.n273 gnd 0.2344f
C2517 vdd.n274 gnd 0.148745f
C2518 vdd.t183 gnd 0.034106f
C2519 vdd.t250 gnd 0.034106f
C2520 vdd.n275 gnd 0.2344f
C2521 vdd.n276 gnd 0.148745f
C2522 vdd.t251 gnd 0.034106f
C2523 vdd.t162 gnd 0.034106f
C2524 vdd.n277 gnd 0.2344f
C2525 vdd.n278 gnd 0.148745f
C2526 vdd.n279 gnd 0.005814f
C2527 vdd.n280 gnd 0.005395f
C2528 vdd.n281 gnd 0.002984f
C2529 vdd.n282 gnd 0.006852f
C2530 vdd.n283 gnd 0.002899f
C2531 vdd.n284 gnd 0.00307f
C2532 vdd.n285 gnd 0.005395f
C2533 vdd.n286 gnd 0.002899f
C2534 vdd.n287 gnd 0.006852f
C2535 vdd.n288 gnd 0.00307f
C2536 vdd.n289 gnd 0.005395f
C2537 vdd.n290 gnd 0.002899f
C2538 vdd.n291 gnd 0.005139f
C2539 vdd.n292 gnd 0.005155f
C2540 vdd.t233 gnd 0.014721f
C2541 vdd.n293 gnd 0.032755f
C2542 vdd.n294 gnd 0.170464f
C2543 vdd.n295 gnd 0.002899f
C2544 vdd.n296 gnd 0.00307f
C2545 vdd.n297 gnd 0.006852f
C2546 vdd.n298 gnd 0.006852f
C2547 vdd.n299 gnd 0.00307f
C2548 vdd.n300 gnd 0.002899f
C2549 vdd.n301 gnd 0.005395f
C2550 vdd.n302 gnd 0.005395f
C2551 vdd.n303 gnd 0.002899f
C2552 vdd.n304 gnd 0.00307f
C2553 vdd.n305 gnd 0.006852f
C2554 vdd.n306 gnd 0.006852f
C2555 vdd.n307 gnd 0.00307f
C2556 vdd.n308 gnd 0.002899f
C2557 vdd.n309 gnd 0.005395f
C2558 vdd.n310 gnd 0.005395f
C2559 vdd.n311 gnd 0.002899f
C2560 vdd.n312 gnd 0.00307f
C2561 vdd.n313 gnd 0.006852f
C2562 vdd.n314 gnd 0.006852f
C2563 vdd.n315 gnd 0.0162f
C2564 vdd.n316 gnd 0.002984f
C2565 vdd.n317 gnd 0.002899f
C2566 vdd.n318 gnd 0.013944f
C2567 vdd.n319 gnd 0.00943f
C2568 vdd.n320 gnd 0.065836f
C2569 vdd.n321 gnd 0.265659f
C2570 vdd.n322 gnd 0.008142f
C2571 vdd.n323 gnd 0.010593f
C2572 vdd.n324 gnd 0.008527f
C2573 vdd.n325 gnd 0.008527f
C2574 vdd.n326 gnd 0.010593f
C2575 vdd.n327 gnd 0.010593f
C2576 vdd.n328 gnd 0.774064f
C2577 vdd.n329 gnd 0.010593f
C2578 vdd.n330 gnd 0.010593f
C2579 vdd.n331 gnd 0.010593f
C2580 vdd.n332 gnd 0.839021f
C2581 vdd.n333 gnd 0.010593f
C2582 vdd.n334 gnd 0.010593f
C2583 vdd.n335 gnd 0.010593f
C2584 vdd.n336 gnd 0.010593f
C2585 vdd.n337 gnd 0.008527f
C2586 vdd.n338 gnd 0.010593f
C2587 vdd.t168 gnd 0.541304f
C2588 vdd.n339 gnd 0.010593f
C2589 vdd.n340 gnd 0.010593f
C2590 vdd.n341 gnd 0.010593f
C2591 vdd.t194 gnd 0.541304f
C2592 vdd.n342 gnd 0.010593f
C2593 vdd.n343 gnd 0.010593f
C2594 vdd.n344 gnd 0.010593f
C2595 vdd.n345 gnd 0.010593f
C2596 vdd.n346 gnd 0.010593f
C2597 vdd.n347 gnd 0.008527f
C2598 vdd.n348 gnd 0.010593f
C2599 vdd.n349 gnd 0.611673f
C2600 vdd.n350 gnd 0.010593f
C2601 vdd.n351 gnd 0.010593f
C2602 vdd.n352 gnd 0.010593f
C2603 vdd.t146 gnd 0.541304f
C2604 vdd.n353 gnd 0.010593f
C2605 vdd.n354 gnd 0.010593f
C2606 vdd.n355 gnd 0.010593f
C2607 vdd.n356 gnd 0.010593f
C2608 vdd.n357 gnd 0.010593f
C2609 vdd.n358 gnd 0.008527f
C2610 vdd.n359 gnd 0.010593f
C2611 vdd.t153 gnd 0.541304f
C2612 vdd.n360 gnd 0.010593f
C2613 vdd.n361 gnd 0.010593f
C2614 vdd.n362 gnd 0.010593f
C2615 vdd.n363 gnd 0.914803f
C2616 vdd.n364 gnd 0.010593f
C2617 vdd.n365 gnd 0.010593f
C2618 vdd.n366 gnd 0.010593f
C2619 vdd.n367 gnd 0.010593f
C2620 vdd.n368 gnd 0.010593f
C2621 vdd.n369 gnd 0.007077f
C2622 vdd.n370 gnd 0.024124f
C2623 vdd.t32 gnd 0.541304f
C2624 vdd.n371 gnd 0.010593f
C2625 vdd.n372 gnd 0.024124f
C2626 vdd.n404 gnd 0.010593f
C2627 vdd.t34 gnd 0.130328f
C2628 vdd.t33 gnd 0.139285f
C2629 vdd.t31 gnd 0.170207f
C2630 vdd.n405 gnd 0.218181f
C2631 vdd.n406 gnd 0.184164f
C2632 vdd.n407 gnd 0.013984f
C2633 vdd.n408 gnd 0.010593f
C2634 vdd.n409 gnd 0.008527f
C2635 vdd.n410 gnd 0.010593f
C2636 vdd.n411 gnd 0.008527f
C2637 vdd.n412 gnd 0.010593f
C2638 vdd.n413 gnd 0.008527f
C2639 vdd.n414 gnd 0.010593f
C2640 vdd.n415 gnd 0.008527f
C2641 vdd.n416 gnd 0.010593f
C2642 vdd.n417 gnd 0.008527f
C2643 vdd.n418 gnd 0.010593f
C2644 vdd.t92 gnd 0.130328f
C2645 vdd.t91 gnd 0.139285f
C2646 vdd.t90 gnd 0.170207f
C2647 vdd.n419 gnd 0.218181f
C2648 vdd.n420 gnd 0.184164f
C2649 vdd.n421 gnd 0.008527f
C2650 vdd.n422 gnd 0.010593f
C2651 vdd.n423 gnd 0.008527f
C2652 vdd.n424 gnd 0.010593f
C2653 vdd.n425 gnd 0.008527f
C2654 vdd.n426 gnd 0.010593f
C2655 vdd.n427 gnd 0.008527f
C2656 vdd.n428 gnd 0.010593f
C2657 vdd.n429 gnd 0.008527f
C2658 vdd.n430 gnd 0.010593f
C2659 vdd.t98 gnd 0.130328f
C2660 vdd.t97 gnd 0.139285f
C2661 vdd.t96 gnd 0.170207f
C2662 vdd.n431 gnd 0.218181f
C2663 vdd.n432 gnd 0.184164f
C2664 vdd.n433 gnd 0.018247f
C2665 vdd.n434 gnd 0.010593f
C2666 vdd.n435 gnd 0.008527f
C2667 vdd.n436 gnd 0.010593f
C2668 vdd.n437 gnd 0.008527f
C2669 vdd.n438 gnd 0.010593f
C2670 vdd.n439 gnd 0.008527f
C2671 vdd.n440 gnd 0.010593f
C2672 vdd.n441 gnd 0.008527f
C2673 vdd.n442 gnd 0.010593f
C2674 vdd.n443 gnd 0.024124f
C2675 vdd.n444 gnd 0.024289f
C2676 vdd.n445 gnd 0.024289f
C2677 vdd.n446 gnd 0.007077f
C2678 vdd.n447 gnd 0.008527f
C2679 vdd.n448 gnd 0.010593f
C2680 vdd.n449 gnd 0.010593f
C2681 vdd.n450 gnd 0.008527f
C2682 vdd.n451 gnd 0.010593f
C2683 vdd.n452 gnd 0.010593f
C2684 vdd.n453 gnd 0.010593f
C2685 vdd.n454 gnd 0.010593f
C2686 vdd.n455 gnd 0.010593f
C2687 vdd.n456 gnd 0.008527f
C2688 vdd.n457 gnd 0.008527f
C2689 vdd.n458 gnd 0.010593f
C2690 vdd.n459 gnd 0.010593f
C2691 vdd.n460 gnd 0.008527f
C2692 vdd.n461 gnd 0.010593f
C2693 vdd.n462 gnd 0.010593f
C2694 vdd.n463 gnd 0.010593f
C2695 vdd.n464 gnd 0.010593f
C2696 vdd.n465 gnd 0.010593f
C2697 vdd.n466 gnd 0.008527f
C2698 vdd.n467 gnd 0.008527f
C2699 vdd.n468 gnd 0.010593f
C2700 vdd.n469 gnd 0.010593f
C2701 vdd.n470 gnd 0.008527f
C2702 vdd.n471 gnd 0.010593f
C2703 vdd.n472 gnd 0.010593f
C2704 vdd.n473 gnd 0.010593f
C2705 vdd.n474 gnd 0.010593f
C2706 vdd.n475 gnd 0.010593f
C2707 vdd.n476 gnd 0.008527f
C2708 vdd.n477 gnd 0.008527f
C2709 vdd.n478 gnd 0.010593f
C2710 vdd.n479 gnd 0.010593f
C2711 vdd.n480 gnd 0.008527f
C2712 vdd.n481 gnd 0.010593f
C2713 vdd.n482 gnd 0.010593f
C2714 vdd.n483 gnd 0.010593f
C2715 vdd.n484 gnd 0.010593f
C2716 vdd.n485 gnd 0.010593f
C2717 vdd.n486 gnd 0.008527f
C2718 vdd.n487 gnd 0.008527f
C2719 vdd.n488 gnd 0.010593f
C2720 vdd.n489 gnd 0.010593f
C2721 vdd.n490 gnd 0.00712f
C2722 vdd.n491 gnd 0.010593f
C2723 vdd.n492 gnd 0.010593f
C2724 vdd.n493 gnd 0.010593f
C2725 vdd.n494 gnd 0.010593f
C2726 vdd.n495 gnd 0.010593f
C2727 vdd.n496 gnd 0.00712f
C2728 vdd.n497 gnd 0.008527f
C2729 vdd.n498 gnd 0.010593f
C2730 vdd.n499 gnd 0.010593f
C2731 vdd.n500 gnd 0.008527f
C2732 vdd.n501 gnd 0.010593f
C2733 vdd.n502 gnd 0.010593f
C2734 vdd.n503 gnd 0.010593f
C2735 vdd.n504 gnd 0.010593f
C2736 vdd.n505 gnd 0.010593f
C2737 vdd.n506 gnd 0.008527f
C2738 vdd.n507 gnd 0.008527f
C2739 vdd.n508 gnd 0.010593f
C2740 vdd.n509 gnd 0.010593f
C2741 vdd.n510 gnd 0.008527f
C2742 vdd.n511 gnd 0.010593f
C2743 vdd.n512 gnd 0.010593f
C2744 vdd.n513 gnd 0.010593f
C2745 vdd.n514 gnd 0.010593f
C2746 vdd.n515 gnd 0.010593f
C2747 vdd.n516 gnd 0.008527f
C2748 vdd.n517 gnd 0.008527f
C2749 vdd.n518 gnd 0.010593f
C2750 vdd.n519 gnd 0.010593f
C2751 vdd.n520 gnd 0.008527f
C2752 vdd.n521 gnd 0.010593f
C2753 vdd.n522 gnd 0.010593f
C2754 vdd.n523 gnd 0.010593f
C2755 vdd.n524 gnd 0.010593f
C2756 vdd.n525 gnd 0.010593f
C2757 vdd.n526 gnd 0.008527f
C2758 vdd.n527 gnd 0.008527f
C2759 vdd.n528 gnd 0.010593f
C2760 vdd.n529 gnd 0.010593f
C2761 vdd.n530 gnd 0.008527f
C2762 vdd.n531 gnd 0.010593f
C2763 vdd.n532 gnd 0.010593f
C2764 vdd.n533 gnd 0.010593f
C2765 vdd.n534 gnd 0.010593f
C2766 vdd.n535 gnd 0.010593f
C2767 vdd.n536 gnd 0.008527f
C2768 vdd.n537 gnd 0.008527f
C2769 vdd.n538 gnd 0.010593f
C2770 vdd.n539 gnd 0.010593f
C2771 vdd.n540 gnd 0.008527f
C2772 vdd.n541 gnd 0.010593f
C2773 vdd.n542 gnd 0.010593f
C2774 vdd.n543 gnd 0.010593f
C2775 vdd.n544 gnd 0.010593f
C2776 vdd.n545 gnd 0.010593f
C2777 vdd.n546 gnd 0.005798f
C2778 vdd.n547 gnd 0.018247f
C2779 vdd.n548 gnd 0.010593f
C2780 vdd.n549 gnd 0.010593f
C2781 vdd.n550 gnd 0.008441f
C2782 vdd.n551 gnd 0.010593f
C2783 vdd.n552 gnd 0.010593f
C2784 vdd.n553 gnd 0.010593f
C2785 vdd.n554 gnd 0.010593f
C2786 vdd.n555 gnd 0.010593f
C2787 vdd.n556 gnd 0.008527f
C2788 vdd.n557 gnd 0.008527f
C2789 vdd.n558 gnd 0.010593f
C2790 vdd.n559 gnd 0.010593f
C2791 vdd.n560 gnd 0.008527f
C2792 vdd.n561 gnd 0.010593f
C2793 vdd.n562 gnd 0.010593f
C2794 vdd.n563 gnd 0.010593f
C2795 vdd.n564 gnd 0.010593f
C2796 vdd.n565 gnd 0.010593f
C2797 vdd.n566 gnd 0.008527f
C2798 vdd.n567 gnd 0.008527f
C2799 vdd.n568 gnd 0.010593f
C2800 vdd.n569 gnd 0.010593f
C2801 vdd.n570 gnd 0.008527f
C2802 vdd.n571 gnd 0.010593f
C2803 vdd.n572 gnd 0.010593f
C2804 vdd.n573 gnd 0.010593f
C2805 vdd.n574 gnd 0.010593f
C2806 vdd.n575 gnd 0.010593f
C2807 vdd.n576 gnd 0.008527f
C2808 vdd.n577 gnd 0.008527f
C2809 vdd.n578 gnd 0.010593f
C2810 vdd.n579 gnd 0.010593f
C2811 vdd.n580 gnd 0.008527f
C2812 vdd.n581 gnd 0.010593f
C2813 vdd.n582 gnd 0.010593f
C2814 vdd.n583 gnd 0.010593f
C2815 vdd.n584 gnd 0.010593f
C2816 vdd.n585 gnd 0.010593f
C2817 vdd.n586 gnd 0.008527f
C2818 vdd.n587 gnd 0.008527f
C2819 vdd.n588 gnd 0.010593f
C2820 vdd.n589 gnd 0.010593f
C2821 vdd.n590 gnd 0.008527f
C2822 vdd.n591 gnd 0.010593f
C2823 vdd.n592 gnd 0.010593f
C2824 vdd.n593 gnd 0.010593f
C2825 vdd.n594 gnd 0.010593f
C2826 vdd.n595 gnd 0.010593f
C2827 vdd.n596 gnd 0.008527f
C2828 vdd.n597 gnd 0.010593f
C2829 vdd.n598 gnd 0.008527f
C2830 vdd.n599 gnd 0.004476f
C2831 vdd.n600 gnd 0.010593f
C2832 vdd.n601 gnd 0.010593f
C2833 vdd.n602 gnd 0.008527f
C2834 vdd.n603 gnd 0.010593f
C2835 vdd.n604 gnd 0.008527f
C2836 vdd.n605 gnd 0.010593f
C2837 vdd.n606 gnd 0.008527f
C2838 vdd.n607 gnd 0.010593f
C2839 vdd.n608 gnd 0.008527f
C2840 vdd.n609 gnd 0.010593f
C2841 vdd.n610 gnd 0.008527f
C2842 vdd.n611 gnd 0.010593f
C2843 vdd.n612 gnd 0.010593f
C2844 vdd.n613 gnd 0.590021f
C2845 vdd.t173 gnd 0.541304f
C2846 vdd.n614 gnd 0.010593f
C2847 vdd.n615 gnd 0.008527f
C2848 vdd.n616 gnd 0.010593f
C2849 vdd.n617 gnd 0.008527f
C2850 vdd.n618 gnd 0.010593f
C2851 vdd.t218 gnd 0.541304f
C2852 vdd.n619 gnd 0.010593f
C2853 vdd.n620 gnd 0.008527f
C2854 vdd.n621 gnd 0.010593f
C2855 vdd.n622 gnd 0.008527f
C2856 vdd.n623 gnd 0.010593f
C2857 vdd.t163 gnd 0.541304f
C2858 vdd.n624 gnd 0.67663f
C2859 vdd.n625 gnd 0.010593f
C2860 vdd.n626 gnd 0.008527f
C2861 vdd.n627 gnd 0.010593f
C2862 vdd.n628 gnd 0.008527f
C2863 vdd.n629 gnd 0.010593f
C2864 vdd.t130 gnd 0.541304f
C2865 vdd.n630 gnd 0.010593f
C2866 vdd.n631 gnd 0.008527f
C2867 vdd.n632 gnd 0.010593f
C2868 vdd.n633 gnd 0.008527f
C2869 vdd.n634 gnd 0.010593f
C2870 vdd.n635 gnd 0.752412f
C2871 vdd.n636 gnd 0.898564f
C2872 vdd.t191 gnd 0.541304f
C2873 vdd.n637 gnd 0.010593f
C2874 vdd.n638 gnd 0.008527f
C2875 vdd.n639 gnd 0.010593f
C2876 vdd.n640 gnd 0.008527f
C2877 vdd.n641 gnd 0.010593f
C2878 vdd.n642 gnd 0.568369f
C2879 vdd.n643 gnd 0.010593f
C2880 vdd.n644 gnd 0.008527f
C2881 vdd.n645 gnd 0.010593f
C2882 vdd.n646 gnd 0.008527f
C2883 vdd.n647 gnd 0.010593f
C2884 vdd.n648 gnd 1.08261f
C2885 vdd.t134 gnd 0.541304f
C2886 vdd.n649 gnd 0.010593f
C2887 vdd.n650 gnd 0.008527f
C2888 vdd.n651 gnd 0.010593f
C2889 vdd.n652 gnd 0.008527f
C2890 vdd.n653 gnd 0.010593f
C2891 vdd.t28 gnd 0.541304f
C2892 vdd.n654 gnd 0.010593f
C2893 vdd.n655 gnd 0.008527f
C2894 vdd.n656 gnd 0.024289f
C2895 vdd.n657 gnd 0.024289f
C2896 vdd.n658 gnd 7.65404f
C2897 vdd.n659 gnd 0.600847f
C2898 vdd.n660 gnd 0.024289f
C2899 vdd.n661 gnd 0.00911f
C2900 vdd.n662 gnd 0.008527f
C2901 vdd.n667 gnd 0.00678f
C2902 vdd.n668 gnd 0.008527f
C2903 vdd.n669 gnd 0.010593f
C2904 vdd.n670 gnd 0.010593f
C2905 vdd.n671 gnd 0.010593f
C2906 vdd.n672 gnd 0.010593f
C2907 vdd.n673 gnd 0.010593f
C2908 vdd.n674 gnd 0.008527f
C2909 vdd.n675 gnd 0.010593f
C2910 vdd.n676 gnd 0.010593f
C2911 vdd.n677 gnd 0.010593f
C2912 vdd.n678 gnd 0.010593f
C2913 vdd.n679 gnd 0.010593f
C2914 vdd.n680 gnd 0.008527f
C2915 vdd.n681 gnd 0.010593f
C2916 vdd.n682 gnd 0.010593f
C2917 vdd.n683 gnd 0.010593f
C2918 vdd.n684 gnd 0.010593f
C2919 vdd.n685 gnd 0.010593f
C2920 vdd.t40 gnd 0.130328f
C2921 vdd.t41 gnd 0.139285f
C2922 vdd.t39 gnd 0.170207f
C2923 vdd.n686 gnd 0.218181f
C2924 vdd.n687 gnd 0.183312f
C2925 vdd.n688 gnd 0.017394f
C2926 vdd.n689 gnd 0.010593f
C2927 vdd.n690 gnd 0.010593f
C2928 vdd.n691 gnd 0.010593f
C2929 vdd.n692 gnd 0.010593f
C2930 vdd.n693 gnd 0.010593f
C2931 vdd.n694 gnd 0.008527f
C2932 vdd.n695 gnd 0.010593f
C2933 vdd.n696 gnd 0.010593f
C2934 vdd.n697 gnd 0.010593f
C2935 vdd.n698 gnd 0.010593f
C2936 vdd.n699 gnd 0.010593f
C2937 vdd.n700 gnd 0.008527f
C2938 vdd.n701 gnd 0.010593f
C2939 vdd.n702 gnd 0.010593f
C2940 vdd.n703 gnd 0.010593f
C2941 vdd.n704 gnd 0.010593f
C2942 vdd.n705 gnd 0.010593f
C2943 vdd.n706 gnd 0.008527f
C2944 vdd.n707 gnd 0.010593f
C2945 vdd.n708 gnd 0.010593f
C2946 vdd.n709 gnd 0.010593f
C2947 vdd.n710 gnd 0.010593f
C2948 vdd.n711 gnd 0.010593f
C2949 vdd.n712 gnd 0.008527f
C2950 vdd.n713 gnd 0.010593f
C2951 vdd.n714 gnd 0.010593f
C2952 vdd.n715 gnd 0.010593f
C2953 vdd.n716 gnd 0.010593f
C2954 vdd.n717 gnd 0.010593f
C2955 vdd.n718 gnd 0.008527f
C2956 vdd.n719 gnd 0.010593f
C2957 vdd.n720 gnd 0.010593f
C2958 vdd.n721 gnd 0.010593f
C2959 vdd.n722 gnd 0.008441f
C2960 vdd.t29 gnd 0.130328f
C2961 vdd.t30 gnd 0.139285f
C2962 vdd.t27 gnd 0.170207f
C2963 vdd.n723 gnd 0.218181f
C2964 vdd.n724 gnd 0.183312f
C2965 vdd.n725 gnd 0.010593f
C2966 vdd.n726 gnd 0.008527f
C2967 vdd.n728 gnd 0.010593f
C2968 vdd.n730 gnd 0.010593f
C2969 vdd.n731 gnd 0.010593f
C2970 vdd.n732 gnd 0.008527f
C2971 vdd.n733 gnd 0.010593f
C2972 vdd.n734 gnd 0.010593f
C2973 vdd.n735 gnd 0.010593f
C2974 vdd.n736 gnd 0.010593f
C2975 vdd.n737 gnd 0.010593f
C2976 vdd.n738 gnd 0.008527f
C2977 vdd.n739 gnd 0.010593f
C2978 vdd.n740 gnd 0.010593f
C2979 vdd.n741 gnd 0.010593f
C2980 vdd.n742 gnd 0.010593f
C2981 vdd.n743 gnd 0.010593f
C2982 vdd.n744 gnd 0.008527f
C2983 vdd.n745 gnd 0.010593f
C2984 vdd.n746 gnd 0.010593f
C2985 vdd.n747 gnd 0.010593f
C2986 vdd.n748 gnd 0.00678f
C2987 vdd.n753 gnd 0.007204f
C2988 vdd.n754 gnd 0.007204f
C2989 vdd.n755 gnd 0.007204f
C2990 vdd.n756 gnd 7.45917f
C2991 vdd.n757 gnd 0.007204f
C2992 vdd.n758 gnd 0.007204f
C2993 vdd.n759 gnd 0.007204f
C2994 vdd.n761 gnd 0.007204f
C2995 vdd.n762 gnd 0.007204f
C2996 vdd.n764 gnd 0.007204f
C2997 vdd.n765 gnd 0.005244f
C2998 vdd.n767 gnd 0.007204f
C2999 vdd.t76 gnd 0.291096f
C3000 vdd.t75 gnd 0.297973f
C3001 vdd.t74 gnd 0.190039f
C3002 vdd.n768 gnd 0.102706f
C3003 vdd.n769 gnd 0.058258f
C3004 vdd.n770 gnd 0.010295f
C3005 vdd.n771 gnd 0.016836f
C3006 vdd.n773 gnd 0.007204f
C3007 vdd.n774 gnd 0.736173f
C3008 vdd.n775 gnd 0.015959f
C3009 vdd.n776 gnd 0.015959f
C3010 vdd.n777 gnd 0.007204f
C3011 vdd.n778 gnd 0.017093f
C3012 vdd.n779 gnd 0.007204f
C3013 vdd.n780 gnd 0.007204f
C3014 vdd.n781 gnd 0.007204f
C3015 vdd.n782 gnd 0.007204f
C3016 vdd.n783 gnd 0.007204f
C3017 vdd.n785 gnd 0.007204f
C3018 vdd.n786 gnd 0.007204f
C3019 vdd.n788 gnd 0.007204f
C3020 vdd.n789 gnd 0.007204f
C3021 vdd.n791 gnd 0.007204f
C3022 vdd.n792 gnd 0.007204f
C3023 vdd.n794 gnd 0.007204f
C3024 vdd.n795 gnd 0.007204f
C3025 vdd.n797 gnd 0.007204f
C3026 vdd.n798 gnd 0.007204f
C3027 vdd.n800 gnd 0.007204f
C3028 vdd.n801 gnd 0.005244f
C3029 vdd.n803 gnd 0.007204f
C3030 vdd.t69 gnd 0.291096f
C3031 vdd.t68 gnd 0.297973f
C3032 vdd.t66 gnd 0.190039f
C3033 vdd.n804 gnd 0.102706f
C3034 vdd.n805 gnd 0.058258f
C3035 vdd.n806 gnd 0.010295f
C3036 vdd.n807 gnd 0.007204f
C3037 vdd.n808 gnd 0.007204f
C3038 vdd.t67 gnd 0.368087f
C3039 vdd.n809 gnd 0.007204f
C3040 vdd.n810 gnd 0.007204f
C3041 vdd.n811 gnd 0.007204f
C3042 vdd.n812 gnd 0.007204f
C3043 vdd.n813 gnd 0.007204f
C3044 vdd.n814 gnd 0.736173f
C3045 vdd.n815 gnd 0.007204f
C3046 vdd.n816 gnd 0.007204f
C3047 vdd.n817 gnd 0.644151f
C3048 vdd.n818 gnd 0.007204f
C3049 vdd.n819 gnd 0.007204f
C3050 vdd.n820 gnd 0.006356f
C3051 vdd.n821 gnd 0.007204f
C3052 vdd.n822 gnd 0.649565f
C3053 vdd.n823 gnd 0.007204f
C3054 vdd.n824 gnd 0.007204f
C3055 vdd.n825 gnd 0.007204f
C3056 vdd.n826 gnd 0.007204f
C3057 vdd.n827 gnd 0.007204f
C3058 vdd.n828 gnd 0.736173f
C3059 vdd.n829 gnd 0.007204f
C3060 vdd.n830 gnd 0.007204f
C3061 vdd.t50 gnd 0.330195f
C3062 vdd.t9 gnd 0.086609f
C3063 vdd.n831 gnd 0.007204f
C3064 vdd.n832 gnd 0.007204f
C3065 vdd.n833 gnd 0.007204f
C3066 vdd.t99 gnd 0.368087f
C3067 vdd.n834 gnd 0.007204f
C3068 vdd.n835 gnd 0.007204f
C3069 vdd.n836 gnd 0.007204f
C3070 vdd.n837 gnd 0.007204f
C3071 vdd.n838 gnd 0.007204f
C3072 vdd.t22 gnd 0.368087f
C3073 vdd.n839 gnd 0.007204f
C3074 vdd.n840 gnd 0.007204f
C3075 vdd.n841 gnd 0.611673f
C3076 vdd.n842 gnd 0.007204f
C3077 vdd.n843 gnd 0.007204f
C3078 vdd.n844 gnd 0.007204f
C3079 vdd.n845 gnd 0.449282f
C3080 vdd.n846 gnd 0.007204f
C3081 vdd.n847 gnd 0.007204f
C3082 vdd.t121 gnd 0.368087f
C3083 vdd.n848 gnd 0.007204f
C3084 vdd.n849 gnd 0.007204f
C3085 vdd.n850 gnd 0.007204f
C3086 vdd.n851 gnd 0.611673f
C3087 vdd.n852 gnd 0.007204f
C3088 vdd.n853 gnd 0.007204f
C3089 vdd.t108 gnd 0.313956f
C3090 vdd.t117 gnd 0.286891f
C3091 vdd.n854 gnd 0.007204f
C3092 vdd.n855 gnd 0.007204f
C3093 vdd.n856 gnd 0.007204f
C3094 vdd.t103 gnd 0.368087f
C3095 vdd.n857 gnd 0.007204f
C3096 vdd.n858 gnd 0.007204f
C3097 vdd.t8 gnd 0.368087f
C3098 vdd.n859 gnd 0.007204f
C3099 vdd.n860 gnd 0.007204f
C3100 vdd.n861 gnd 0.007204f
C3101 vdd.t105 gnd 0.270652f
C3102 vdd.n862 gnd 0.007204f
C3103 vdd.n863 gnd 0.007204f
C3104 vdd.n864 gnd 0.627912f
C3105 vdd.n865 gnd 0.007204f
C3106 vdd.n866 gnd 0.007204f
C3107 vdd.n867 gnd 0.007204f
C3108 vdd.n868 gnd 0.736173f
C3109 vdd.n869 gnd 0.007204f
C3110 vdd.n870 gnd 0.007204f
C3111 vdd.t10 gnd 0.330195f
C3112 vdd.n871 gnd 0.465521f
C3113 vdd.n872 gnd 0.007204f
C3114 vdd.n873 gnd 0.007204f
C3115 vdd.n874 gnd 0.007204f
C3116 vdd.t119 gnd 0.368087f
C3117 vdd.n875 gnd 0.007204f
C3118 vdd.n876 gnd 0.007204f
C3119 vdd.n877 gnd 0.007204f
C3120 vdd.n878 gnd 0.007204f
C3121 vdd.n879 gnd 0.007204f
C3122 vdd.t260 gnd 0.736173f
C3123 vdd.n880 gnd 0.007204f
C3124 vdd.n881 gnd 0.007204f
C3125 vdd.t71 gnd 0.368087f
C3126 vdd.n882 gnd 0.007204f
C3127 vdd.n883 gnd 0.017093f
C3128 vdd.n884 gnd 0.017093f
C3129 vdd.t106 gnd 0.692869f
C3130 vdd.n885 gnd 0.015959f
C3131 vdd.n886 gnd 0.015959f
C3132 vdd.n887 gnd 0.017093f
C3133 vdd.n888 gnd 0.007204f
C3134 vdd.n889 gnd 0.007204f
C3135 vdd.t109 gnd 0.692869f
C3136 vdd.n907 gnd 0.017093f
C3137 vdd.n925 gnd 0.015959f
C3138 vdd.n926 gnd 0.007204f
C3139 vdd.n927 gnd 0.015959f
C3140 vdd.t89 gnd 0.291096f
C3141 vdd.t88 gnd 0.297973f
C3142 vdd.t87 gnd 0.190039f
C3143 vdd.n928 gnd 0.102706f
C3144 vdd.n929 gnd 0.058258f
C3145 vdd.n930 gnd 0.016836f
C3146 vdd.n931 gnd 0.007204f
C3147 vdd.t256 gnd 0.736173f
C3148 vdd.n932 gnd 0.015959f
C3149 vdd.n933 gnd 0.007204f
C3150 vdd.n934 gnd 0.017093f
C3151 vdd.n935 gnd 0.007204f
C3152 vdd.t65 gnd 0.291096f
C3153 vdd.t64 gnd 0.297973f
C3154 vdd.t62 gnd 0.190039f
C3155 vdd.n936 gnd 0.102706f
C3156 vdd.n937 gnd 0.058258f
C3157 vdd.n938 gnd 0.010295f
C3158 vdd.n939 gnd 0.007204f
C3159 vdd.n940 gnd 0.007204f
C3160 vdd.t63 gnd 0.368087f
C3161 vdd.n941 gnd 0.007204f
C3162 vdd.n942 gnd 0.007204f
C3163 vdd.n943 gnd 0.007204f
C3164 vdd.n944 gnd 0.007204f
C3165 vdd.n945 gnd 0.007204f
C3166 vdd.n946 gnd 0.007204f
C3167 vdd.n947 gnd 0.736173f
C3168 vdd.n948 gnd 0.007204f
C3169 vdd.n949 gnd 0.007204f
C3170 vdd.t115 gnd 0.368087f
C3171 vdd.n950 gnd 0.007204f
C3172 vdd.n951 gnd 0.007204f
C3173 vdd.n952 gnd 0.007204f
C3174 vdd.n953 gnd 0.007204f
C3175 vdd.n954 gnd 0.465521f
C3176 vdd.n955 gnd 0.007204f
C3177 vdd.n956 gnd 0.007204f
C3178 vdd.n957 gnd 0.007204f
C3179 vdd.n958 gnd 0.007204f
C3180 vdd.n959 gnd 0.007204f
C3181 vdd.n960 gnd 0.627912f
C3182 vdd.n961 gnd 0.007204f
C3183 vdd.n962 gnd 0.007204f
C3184 vdd.t4 gnd 0.330195f
C3185 vdd.t0 gnd 0.270652f
C3186 vdd.n963 gnd 0.007204f
C3187 vdd.n964 gnd 0.007204f
C3188 vdd.n965 gnd 0.007204f
C3189 vdd.t7 gnd 0.368087f
C3190 vdd.n966 gnd 0.007204f
C3191 vdd.n967 gnd 0.007204f
C3192 vdd.t2 gnd 0.368087f
C3193 vdd.n968 gnd 0.007204f
C3194 vdd.n969 gnd 0.007204f
C3195 vdd.n970 gnd 0.007204f
C3196 vdd.t101 gnd 0.286891f
C3197 vdd.n971 gnd 0.007204f
C3198 vdd.n972 gnd 0.007204f
C3199 vdd.n973 gnd 0.611673f
C3200 vdd.n974 gnd 0.007204f
C3201 vdd.n975 gnd 0.007204f
C3202 vdd.n976 gnd 0.007204f
C3203 vdd.t258 gnd 0.368087f
C3204 vdd.n977 gnd 0.007204f
C3205 vdd.n978 gnd 0.007204f
C3206 vdd.t6 gnd 0.313956f
C3207 vdd.n979 gnd 0.449282f
C3208 vdd.n980 gnd 0.007204f
C3209 vdd.n981 gnd 0.007204f
C3210 vdd.n982 gnd 0.007204f
C3211 vdd.n983 gnd 0.611673f
C3212 vdd.n984 gnd 0.007204f
C3213 vdd.n985 gnd 0.007204f
C3214 vdd.t12 gnd 0.368087f
C3215 vdd.n986 gnd 0.007204f
C3216 vdd.n987 gnd 0.007204f
C3217 vdd.n988 gnd 0.007204f
C3218 vdd.n989 gnd 0.736173f
C3219 vdd.n990 gnd 0.007204f
C3220 vdd.n991 gnd 0.007204f
C3221 vdd.t100 gnd 0.368087f
C3222 vdd.n992 gnd 0.007204f
C3223 vdd.n993 gnd 0.007204f
C3224 vdd.n994 gnd 0.007204f
C3225 vdd.t1 gnd 0.086609f
C3226 vdd.n995 gnd 0.007204f
C3227 vdd.n996 gnd 0.007204f
C3228 vdd.n997 gnd 0.007204f
C3229 vdd.t82 gnd 0.297973f
C3230 vdd.t80 gnd 0.190039f
C3231 vdd.t83 gnd 0.297973f
C3232 vdd.n998 gnd 0.167473f
C3233 vdd.n999 gnd 0.007204f
C3234 vdd.n1000 gnd 0.007204f
C3235 vdd.n1001 gnd 0.736173f
C3236 vdd.n1002 gnd 0.007204f
C3237 vdd.n1003 gnd 0.007204f
C3238 vdd.t81 gnd 0.330195f
C3239 vdd.n1004 gnd 0.649565f
C3240 vdd.n1005 gnd 0.007204f
C3241 vdd.n1006 gnd 0.007204f
C3242 vdd.n1007 gnd 0.007204f
C3243 vdd.n1008 gnd 0.644151f
C3244 vdd.n1009 gnd 0.007204f
C3245 vdd.n1010 gnd 0.007204f
C3246 vdd.n1011 gnd 0.007204f
C3247 vdd.n1012 gnd 0.007204f
C3248 vdd.n1013 gnd 0.007204f
C3249 vdd.n1014 gnd 0.736173f
C3250 vdd.n1015 gnd 0.007204f
C3251 vdd.n1016 gnd 0.007204f
C3252 vdd.t24 gnd 0.368087f
C3253 vdd.n1017 gnd 0.007204f
C3254 vdd.n1018 gnd 0.017093f
C3255 vdd.n1019 gnd 0.017093f
C3256 vdd.n1020 gnd 7.45917f
C3257 vdd.n1021 gnd 0.015959f
C3258 vdd.n1022 gnd 0.015959f
C3259 vdd.n1023 gnd 0.017093f
C3260 vdd.n1024 gnd 0.007204f
C3261 vdd.n1025 gnd 0.007204f
C3262 vdd.n1026 gnd 0.007204f
C3263 vdd.n1027 gnd 0.007204f
C3264 vdd.n1028 gnd 0.007204f
C3265 vdd.n1029 gnd 0.007204f
C3266 vdd.n1030 gnd 0.007204f
C3267 vdd.n1031 gnd 0.007204f
C3268 vdd.n1033 gnd 0.007204f
C3269 vdd.n1034 gnd 0.007204f
C3270 vdd.n1035 gnd 0.00678f
C3271 vdd.n1038 gnd 0.024289f
C3272 vdd.n1039 gnd 0.008527f
C3273 vdd.n1040 gnd 0.010593f
C3274 vdd.n1042 gnd 0.010593f
C3275 vdd.n1043 gnd 0.007077f
C3276 vdd.n1044 gnd 0.600847f
C3277 vdd.n1045 gnd 7.65404f
C3278 vdd.n1046 gnd 0.010593f
C3279 vdd.n1047 gnd 0.024289f
C3280 vdd.n1048 gnd 0.008527f
C3281 vdd.n1049 gnd 0.010593f
C3282 vdd.n1050 gnd 0.008527f
C3283 vdd.n1051 gnd 0.010593f
C3284 vdd.n1052 gnd 1.08261f
C3285 vdd.n1053 gnd 0.010593f
C3286 vdd.n1054 gnd 0.008527f
C3287 vdd.n1055 gnd 0.008527f
C3288 vdd.n1056 gnd 0.010593f
C3289 vdd.n1057 gnd 0.008527f
C3290 vdd.n1058 gnd 0.010593f
C3291 vdd.t136 gnd 0.541304f
C3292 vdd.n1059 gnd 0.010593f
C3293 vdd.n1060 gnd 0.008527f
C3294 vdd.n1061 gnd 0.010593f
C3295 vdd.n1062 gnd 0.008527f
C3296 vdd.n1063 gnd 0.010593f
C3297 vdd.t236 gnd 0.541304f
C3298 vdd.n1064 gnd 0.010593f
C3299 vdd.n1065 gnd 0.008527f
C3300 vdd.n1066 gnd 0.010593f
C3301 vdd.n1067 gnd 0.008527f
C3302 vdd.n1068 gnd 0.010593f
C3303 vdd.t144 gnd 0.541304f
C3304 vdd.n1069 gnd 0.752412f
C3305 vdd.n1070 gnd 0.010593f
C3306 vdd.n1071 gnd 0.008527f
C3307 vdd.n1072 gnd 0.010593f
C3308 vdd.n1073 gnd 0.008527f
C3309 vdd.n1074 gnd 0.010593f
C3310 vdd.n1075 gnd 0.860673f
C3311 vdd.n1076 gnd 0.010593f
C3312 vdd.n1077 gnd 0.008527f
C3313 vdd.n1078 gnd 0.010593f
C3314 vdd.n1079 gnd 0.008527f
C3315 vdd.n1080 gnd 0.010593f
C3316 vdd.n1081 gnd 0.67663f
C3317 vdd.t165 gnd 0.541304f
C3318 vdd.n1082 gnd 0.010593f
C3319 vdd.n1083 gnd 0.008527f
C3320 vdd.n1084 gnd 0.010593f
C3321 vdd.n1085 gnd 0.008527f
C3322 vdd.n1086 gnd 0.010593f
C3323 vdd.t186 gnd 0.541304f
C3324 vdd.n1087 gnd 0.010593f
C3325 vdd.n1088 gnd 0.008527f
C3326 vdd.n1089 gnd 0.010593f
C3327 vdd.n1090 gnd 0.008527f
C3328 vdd.n1091 gnd 0.010593f
C3329 vdd.t214 gnd 0.541304f
C3330 vdd.n1092 gnd 0.590021f
C3331 vdd.n1093 gnd 0.010593f
C3332 vdd.n1094 gnd 0.008527f
C3333 vdd.n1095 gnd 0.010593f
C3334 vdd.n1096 gnd 0.008527f
C3335 vdd.n1097 gnd 0.010593f
C3336 vdd.t206 gnd 0.541304f
C3337 vdd.n1098 gnd 0.010593f
C3338 vdd.n1099 gnd 0.008527f
C3339 vdd.n1100 gnd 0.010593f
C3340 vdd.n1101 gnd 0.008527f
C3341 vdd.n1102 gnd 0.010593f
C3342 vdd.n1103 gnd 0.839021f
C3343 vdd.n1104 gnd 0.898564f
C3344 vdd.t142 gnd 0.541304f
C3345 vdd.n1105 gnd 0.010593f
C3346 vdd.n1106 gnd 0.008527f
C3347 vdd.n1107 gnd 0.010593f
C3348 vdd.n1108 gnd 0.008527f
C3349 vdd.n1109 gnd 0.010593f
C3350 vdd.n1110 gnd 0.654978f
C3351 vdd.n1111 gnd 0.010593f
C3352 vdd.n1112 gnd 0.008527f
C3353 vdd.n1113 gnd 0.010593f
C3354 vdd.n1114 gnd 0.008527f
C3355 vdd.n1115 gnd 0.010593f
C3356 vdd.t160 gnd 0.541304f
C3357 vdd.t150 gnd 0.541304f
C3358 vdd.n1116 gnd 0.010593f
C3359 vdd.n1117 gnd 0.008527f
C3360 vdd.n1118 gnd 0.010593f
C3361 vdd.n1119 gnd 0.008527f
C3362 vdd.n1120 gnd 0.010593f
C3363 vdd.t200 gnd 0.541304f
C3364 vdd.n1121 gnd 0.010593f
C3365 vdd.n1122 gnd 0.008527f
C3366 vdd.n1123 gnd 0.010593f
C3367 vdd.n1124 gnd 0.008527f
C3368 vdd.n1125 gnd 0.010593f
C3369 vdd.t202 gnd 0.541304f
C3370 vdd.n1126 gnd 0.795717f
C3371 vdd.n1127 gnd 0.010593f
C3372 vdd.n1128 gnd 0.008527f
C3373 vdd.n1129 gnd 0.010593f
C3374 vdd.n1130 gnd 0.008527f
C3375 vdd.n1131 gnd 0.010593f
C3376 vdd.n1132 gnd 1.08261f
C3377 vdd.n1133 gnd 0.010593f
C3378 vdd.n1134 gnd 0.008527f
C3379 vdd.n1135 gnd 0.010593f
C3380 vdd.n1136 gnd 0.008527f
C3381 vdd.n1137 gnd 0.010593f
C3382 vdd.n1138 gnd 0.914803f
C3383 vdd.n1139 gnd 0.010593f
C3384 vdd.n1140 gnd 0.008527f
C3385 vdd.n1141 gnd 0.024124f
C3386 vdd.n1142 gnd 0.007077f
C3387 vdd.n1143 gnd 0.024124f
C3388 vdd.n1144 gnd 1.42904f
C3389 vdd.n1145 gnd 0.024124f
C3390 vdd.n1146 gnd 0.007077f
C3391 vdd.n1147 gnd 0.010593f
C3392 vdd.t37 gnd 0.130328f
C3393 vdd.t38 gnd 0.139285f
C3394 vdd.t35 gnd 0.170207f
C3395 vdd.n1148 gnd 0.218181f
C3396 vdd.n1149 gnd 0.184164f
C3397 vdd.n1150 gnd 0.013984f
C3398 vdd.n1151 gnd 0.010593f
C3399 vdd.n1182 gnd 0.010593f
C3400 vdd.n1183 gnd 0.010593f
C3401 vdd.n1184 gnd 0.024289f
C3402 vdd.n1185 gnd 0.008527f
C3403 vdd.n1186 gnd 0.010593f
C3404 vdd.n1187 gnd 0.010593f
C3405 vdd.n1188 gnd 0.010593f
C3406 vdd.n1189 gnd 0.010593f
C3407 vdd.n1190 gnd 0.008527f
C3408 vdd.n1191 gnd 0.010593f
C3409 vdd.n1192 gnd 0.010593f
C3410 vdd.n1193 gnd 0.010593f
C3411 vdd.n1194 gnd 0.010593f
C3412 vdd.n1195 gnd 0.010593f
C3413 vdd.n1196 gnd 0.008527f
C3414 vdd.n1197 gnd 0.010593f
C3415 vdd.n1198 gnd 0.010593f
C3416 vdd.n1199 gnd 0.010593f
C3417 vdd.n1200 gnd 0.010593f
C3418 vdd.n1201 gnd 0.010593f
C3419 vdd.n1202 gnd 0.008527f
C3420 vdd.n1203 gnd 0.010593f
C3421 vdd.n1204 gnd 0.010593f
C3422 vdd.n1205 gnd 0.010593f
C3423 vdd.n1206 gnd 0.010593f
C3424 vdd.n1207 gnd 0.010593f
C3425 vdd.n1208 gnd 0.00712f
C3426 vdd.n1209 gnd 0.010593f
C3427 vdd.n1210 gnd 0.010593f
C3428 vdd.n1211 gnd 0.010593f
C3429 vdd.n1212 gnd 0.008527f
C3430 vdd.n1213 gnd 0.010593f
C3431 vdd.n1214 gnd 0.010593f
C3432 vdd.n1215 gnd 0.010593f
C3433 vdd.n1216 gnd 0.010593f
C3434 vdd.n1217 gnd 0.010593f
C3435 vdd.n1218 gnd 0.008527f
C3436 vdd.n1219 gnd 0.010593f
C3437 vdd.n1220 gnd 0.010593f
C3438 vdd.n1221 gnd 0.010593f
C3439 vdd.n1222 gnd 0.010593f
C3440 vdd.n1223 gnd 0.010593f
C3441 vdd.n1224 gnd 0.008527f
C3442 vdd.n1225 gnd 0.010593f
C3443 vdd.n1226 gnd 0.010593f
C3444 vdd.n1227 gnd 0.010593f
C3445 vdd.n1228 gnd 0.010593f
C3446 vdd.n1229 gnd 0.010593f
C3447 vdd.n1230 gnd 0.008527f
C3448 vdd.n1231 gnd 0.010593f
C3449 vdd.n1232 gnd 0.010593f
C3450 vdd.n1233 gnd 0.010593f
C3451 vdd.n1234 gnd 0.010593f
C3452 vdd.n1235 gnd 0.010593f
C3453 vdd.n1236 gnd 0.008527f
C3454 vdd.n1237 gnd 0.010593f
C3455 vdd.n1238 gnd 0.010593f
C3456 vdd.n1239 gnd 0.010593f
C3457 vdd.n1240 gnd 0.010593f
C3458 vdd.n1241 gnd 0.008441f
C3459 vdd.n1242 gnd 0.010593f
C3460 vdd.n1243 gnd 0.010593f
C3461 vdd.n1244 gnd 0.010593f
C3462 vdd.n1245 gnd 0.010593f
C3463 vdd.n1246 gnd 0.010593f
C3464 vdd.n1247 gnd 0.008527f
C3465 vdd.n1248 gnd 0.010593f
C3466 vdd.n1249 gnd 0.010593f
C3467 vdd.n1250 gnd 0.010593f
C3468 vdd.n1251 gnd 0.010593f
C3469 vdd.n1252 gnd 0.010593f
C3470 vdd.n1253 gnd 0.008527f
C3471 vdd.n1254 gnd 0.010593f
C3472 vdd.n1255 gnd 0.010593f
C3473 vdd.n1256 gnd 0.010593f
C3474 vdd.n1257 gnd 0.010593f
C3475 vdd.n1258 gnd 0.010593f
C3476 vdd.n1259 gnd 0.008527f
C3477 vdd.n1260 gnd 0.010593f
C3478 vdd.n1261 gnd 0.010593f
C3479 vdd.n1262 gnd 0.010593f
C3480 vdd.n1263 gnd 0.010593f
C3481 vdd.n1264 gnd 0.010593f
C3482 vdd.n1265 gnd 0.008527f
C3483 vdd.n1266 gnd 0.010593f
C3484 vdd.n1267 gnd 0.010593f
C3485 vdd.n1268 gnd 0.010593f
C3486 vdd.n1269 gnd 0.010593f
C3487 vdd.n1270 gnd 0.010593f
C3488 vdd.n1271 gnd 0.004476f
C3489 vdd.n1272 gnd 0.010593f
C3490 vdd.n1273 gnd 0.008527f
C3491 vdd.n1274 gnd 0.008527f
C3492 vdd.n1275 gnd 0.008527f
C3493 vdd.n1276 gnd 0.010593f
C3494 vdd.n1277 gnd 0.010593f
C3495 vdd.n1278 gnd 0.010593f
C3496 vdd.n1279 gnd 0.008527f
C3497 vdd.n1280 gnd 0.008527f
C3498 vdd.n1281 gnd 0.008527f
C3499 vdd.n1282 gnd 0.010593f
C3500 vdd.n1283 gnd 0.010593f
C3501 vdd.n1284 gnd 0.010593f
C3502 vdd.n1285 gnd 0.008527f
C3503 vdd.n1286 gnd 0.008527f
C3504 vdd.n1287 gnd 0.008527f
C3505 vdd.n1288 gnd 0.010593f
C3506 vdd.n1289 gnd 0.010593f
C3507 vdd.n1290 gnd 0.010593f
C3508 vdd.n1291 gnd 0.008527f
C3509 vdd.n1292 gnd 0.008527f
C3510 vdd.n1293 gnd 0.008527f
C3511 vdd.n1294 gnd 0.010593f
C3512 vdd.n1295 gnd 0.010593f
C3513 vdd.n1296 gnd 0.010593f
C3514 vdd.n1297 gnd 0.008527f
C3515 vdd.n1298 gnd 0.008527f
C3516 vdd.n1299 gnd 0.008527f
C3517 vdd.n1300 gnd 0.010593f
C3518 vdd.n1301 gnd 0.010593f
C3519 vdd.n1302 gnd 0.010593f
C3520 vdd.n1303 gnd 0.010593f
C3521 vdd.t47 gnd 0.130328f
C3522 vdd.t48 gnd 0.139285f
C3523 vdd.t46 gnd 0.170207f
C3524 vdd.n1304 gnd 0.218181f
C3525 vdd.n1305 gnd 0.184164f
C3526 vdd.n1306 gnd 0.018247f
C3527 vdd.n1307 gnd 0.005798f
C3528 vdd.n1308 gnd 0.008527f
C3529 vdd.n1309 gnd 0.010593f
C3530 vdd.n1310 gnd 0.010593f
C3531 vdd.n1311 gnd 0.010593f
C3532 vdd.n1312 gnd 0.008527f
C3533 vdd.n1313 gnd 0.008527f
C3534 vdd.n1314 gnd 0.008527f
C3535 vdd.n1315 gnd 0.010593f
C3536 vdd.n1316 gnd 0.010593f
C3537 vdd.n1317 gnd 0.010593f
C3538 vdd.n1318 gnd 0.008527f
C3539 vdd.n1319 gnd 0.008527f
C3540 vdd.n1320 gnd 0.008527f
C3541 vdd.n1321 gnd 0.010593f
C3542 vdd.n1322 gnd 0.010593f
C3543 vdd.n1323 gnd 0.010593f
C3544 vdd.n1324 gnd 0.008527f
C3545 vdd.n1325 gnd 0.008527f
C3546 vdd.n1326 gnd 0.008527f
C3547 vdd.n1327 gnd 0.010593f
C3548 vdd.n1328 gnd 0.010593f
C3549 vdd.n1329 gnd 0.010593f
C3550 vdd.n1330 gnd 0.008527f
C3551 vdd.n1331 gnd 0.008527f
C3552 vdd.n1332 gnd 0.008527f
C3553 vdd.n1333 gnd 0.010593f
C3554 vdd.n1334 gnd 0.010593f
C3555 vdd.n1335 gnd 0.010593f
C3556 vdd.n1336 gnd 0.008527f
C3557 vdd.n1337 gnd 0.00712f
C3558 vdd.n1338 gnd 0.010593f
C3559 vdd.n1339 gnd 0.010593f
C3560 vdd.t54 gnd 0.130328f
C3561 vdd.t55 gnd 0.139285f
C3562 vdd.t53 gnd 0.170207f
C3563 vdd.n1340 gnd 0.218181f
C3564 vdd.n1341 gnd 0.184164f
C3565 vdd.n1342 gnd 0.018247f
C3566 vdd.n1343 gnd 0.010593f
C3567 vdd.n1344 gnd 0.010593f
C3568 vdd.n1345 gnd 0.010593f
C3569 vdd.n1346 gnd 0.008527f
C3570 vdd.n1347 gnd 0.008527f
C3571 vdd.n1348 gnd 0.008527f
C3572 vdd.n1349 gnd 0.010593f
C3573 vdd.n1350 gnd 0.010593f
C3574 vdd.n1351 gnd 0.010593f
C3575 vdd.n1352 gnd 0.008527f
C3576 vdd.n1353 gnd 0.008527f
C3577 vdd.n1354 gnd 0.008527f
C3578 vdd.n1355 gnd 0.010593f
C3579 vdd.n1356 gnd 0.010593f
C3580 vdd.n1357 gnd 0.010593f
C3581 vdd.n1358 gnd 0.008527f
C3582 vdd.n1359 gnd 0.008527f
C3583 vdd.n1360 gnd 0.008527f
C3584 vdd.n1361 gnd 0.010593f
C3585 vdd.n1362 gnd 0.010593f
C3586 vdd.n1363 gnd 0.010593f
C3587 vdd.n1364 gnd 0.008527f
C3588 vdd.n1365 gnd 0.008527f
C3589 vdd.n1366 gnd 0.008527f
C3590 vdd.n1367 gnd 0.010593f
C3591 vdd.n1368 gnd 0.010593f
C3592 vdd.n1369 gnd 0.010593f
C3593 vdd.n1370 gnd 0.008527f
C3594 vdd.n1371 gnd 0.007077f
C3595 vdd.n1372 gnd 0.024289f
C3596 vdd.n1374 gnd 2.39256f
C3597 vdd.n1375 gnd 0.024289f
C3598 vdd.n1376 gnd 0.00405f
C3599 vdd.n1377 gnd 0.024289f
C3600 vdd.n1378 gnd 0.024124f
C3601 vdd.n1379 gnd 0.010593f
C3602 vdd.n1380 gnd 0.008527f
C3603 vdd.n1381 gnd 0.010593f
C3604 vdd.t36 gnd 0.541304f
C3605 vdd.n1382 gnd 0.709108f
C3606 vdd.n1383 gnd 0.010593f
C3607 vdd.n1384 gnd 0.008527f
C3608 vdd.n1385 gnd 0.010593f
C3609 vdd.n1386 gnd 0.010593f
C3610 vdd.n1387 gnd 0.010593f
C3611 vdd.n1388 gnd 0.008527f
C3612 vdd.n1389 gnd 0.010593f
C3613 vdd.n1390 gnd 1.08261f
C3614 vdd.n1391 gnd 0.010593f
C3615 vdd.n1392 gnd 0.008527f
C3616 vdd.n1393 gnd 0.010593f
C3617 vdd.n1394 gnd 0.010593f
C3618 vdd.n1395 gnd 0.010593f
C3619 vdd.n1396 gnd 0.008527f
C3620 vdd.n1397 gnd 0.010593f
C3621 vdd.n1398 gnd 0.898564f
C3622 vdd.t140 gnd 0.541304f
C3623 vdd.n1399 gnd 0.622499f
C3624 vdd.n1400 gnd 0.010593f
C3625 vdd.n1401 gnd 0.008527f
C3626 vdd.n1402 gnd 0.010593f
C3627 vdd.n1403 gnd 0.010593f
C3628 vdd.n1404 gnd 0.010593f
C3629 vdd.n1405 gnd 0.008527f
C3630 vdd.n1406 gnd 0.010593f
C3631 vdd.n1407 gnd 0.644151f
C3632 vdd.n1408 gnd 0.010593f
C3633 vdd.n1409 gnd 0.008527f
C3634 vdd.n1410 gnd 0.010593f
C3635 vdd.n1411 gnd 0.010593f
C3636 vdd.n1412 gnd 0.010593f
C3637 vdd.n1413 gnd 0.008527f
C3638 vdd.n1414 gnd 0.010593f
C3639 vdd.n1415 gnd 0.611673f
C3640 vdd.n1416 gnd 0.828195f
C3641 vdd.n1417 gnd 0.010593f
C3642 vdd.n1418 gnd 0.008527f
C3643 vdd.n1419 gnd 0.010593f
C3644 vdd.n1420 gnd 0.010593f
C3645 vdd.n1421 gnd 0.010593f
C3646 vdd.n1422 gnd 0.008527f
C3647 vdd.n1423 gnd 0.010593f
C3648 vdd.n1424 gnd 0.898564f
C3649 vdd.n1425 gnd 0.010593f
C3650 vdd.n1426 gnd 0.008527f
C3651 vdd.n1427 gnd 0.010593f
C3652 vdd.n1428 gnd 0.010593f
C3653 vdd.n1429 gnd 0.010593f
C3654 vdd.n1430 gnd 0.008527f
C3655 vdd.n1431 gnd 0.010593f
C3656 vdd.t178 gnd 0.541304f
C3657 vdd.n1432 gnd 0.784891f
C3658 vdd.n1433 gnd 0.010593f
C3659 vdd.n1434 gnd 0.008527f
C3660 vdd.n1435 gnd 0.010593f
C3661 vdd.n1436 gnd 0.010593f
C3662 vdd.n1437 gnd 0.010593f
C3663 vdd.n1438 gnd 0.008527f
C3664 vdd.n1439 gnd 0.010593f
C3665 vdd.n1440 gnd 0.600847f
C3666 vdd.n1441 gnd 0.010593f
C3667 vdd.n1442 gnd 0.008527f
C3668 vdd.n1443 gnd 0.010593f
C3669 vdd.n1444 gnd 0.010593f
C3670 vdd.n1445 gnd 0.010593f
C3671 vdd.n1446 gnd 0.008527f
C3672 vdd.n1447 gnd 0.010593f
C3673 vdd.n1448 gnd 0.774064f
C3674 vdd.n1449 gnd 0.665804f
C3675 vdd.n1450 gnd 0.010593f
C3676 vdd.n1451 gnd 0.008527f
C3677 vdd.n1452 gnd 0.008142f
C3678 vdd.n1453 gnd 0.005814f
C3679 vdd.n1454 gnd 0.005395f
C3680 vdd.n1455 gnd 0.002984f
C3681 vdd.n1456 gnd 0.006852f
C3682 vdd.n1457 gnd 0.002899f
C3683 vdd.n1458 gnd 0.00307f
C3684 vdd.n1459 gnd 0.005395f
C3685 vdd.n1460 gnd 0.002899f
C3686 vdd.n1461 gnd 0.006852f
C3687 vdd.n1462 gnd 0.00307f
C3688 vdd.n1463 gnd 0.005395f
C3689 vdd.n1464 gnd 0.002899f
C3690 vdd.n1465 gnd 0.005139f
C3691 vdd.n1466 gnd 0.005155f
C3692 vdd.t137 gnd 0.014721f
C3693 vdd.n1467 gnd 0.032755f
C3694 vdd.n1468 gnd 0.170464f
C3695 vdd.n1469 gnd 0.002899f
C3696 vdd.n1470 gnd 0.00307f
C3697 vdd.n1471 gnd 0.006852f
C3698 vdd.n1472 gnd 0.006852f
C3699 vdd.n1473 gnd 0.00307f
C3700 vdd.n1474 gnd 0.002899f
C3701 vdd.n1475 gnd 0.005395f
C3702 vdd.n1476 gnd 0.005395f
C3703 vdd.n1477 gnd 0.002899f
C3704 vdd.n1478 gnd 0.00307f
C3705 vdd.n1479 gnd 0.006852f
C3706 vdd.n1480 gnd 0.006852f
C3707 vdd.n1481 gnd 0.00307f
C3708 vdd.n1482 gnd 0.002899f
C3709 vdd.n1483 gnd 0.005395f
C3710 vdd.n1484 gnd 0.005395f
C3711 vdd.n1485 gnd 0.002899f
C3712 vdd.n1486 gnd 0.00307f
C3713 vdd.n1487 gnd 0.006852f
C3714 vdd.n1488 gnd 0.006852f
C3715 vdd.n1489 gnd 0.0162f
C3716 vdd.n1490 gnd 0.002984f
C3717 vdd.n1491 gnd 0.002899f
C3718 vdd.n1492 gnd 0.013944f
C3719 vdd.n1493 gnd 0.009735f
C3720 vdd.t193 gnd 0.034106f
C3721 vdd.t243 gnd 0.034106f
C3722 vdd.n1494 gnd 0.2344f
C3723 vdd.n1495 gnd 0.18432f
C3724 vdd.t166 gnd 0.034106f
C3725 vdd.t224 gnd 0.034106f
C3726 vdd.n1496 gnd 0.2344f
C3727 vdd.n1497 gnd 0.148745f
C3728 vdd.t187 gnd 0.034106f
C3729 vdd.t232 gnd 0.034106f
C3730 vdd.n1498 gnd 0.2344f
C3731 vdd.n1499 gnd 0.148745f
C3732 vdd.t207 gnd 0.034106f
C3733 vdd.t249 gnd 0.034106f
C3734 vdd.n1500 gnd 0.2344f
C3735 vdd.n1501 gnd 0.148745f
C3736 vdd.t179 gnd 0.034106f
C3737 vdd.t143 gnd 0.034106f
C3738 vdd.n1502 gnd 0.2344f
C3739 vdd.n1503 gnd 0.148745f
C3740 vdd.t196 gnd 0.034106f
C3741 vdd.t151 gnd 0.034106f
C3742 vdd.n1504 gnd 0.2344f
C3743 vdd.n1505 gnd 0.148745f
C3744 vdd.t239 gnd 0.034106f
C3745 vdd.t254 gnd 0.034106f
C3746 vdd.n1506 gnd 0.2344f
C3747 vdd.n1507 gnd 0.148745f
C3748 vdd.n1508 gnd 0.005814f
C3749 vdd.n1509 gnd 0.005395f
C3750 vdd.n1510 gnd 0.002984f
C3751 vdd.n1511 gnd 0.006852f
C3752 vdd.n1512 gnd 0.002899f
C3753 vdd.n1513 gnd 0.00307f
C3754 vdd.n1514 gnd 0.005395f
C3755 vdd.n1515 gnd 0.002899f
C3756 vdd.n1516 gnd 0.006852f
C3757 vdd.n1517 gnd 0.00307f
C3758 vdd.n1518 gnd 0.005395f
C3759 vdd.n1519 gnd 0.002899f
C3760 vdd.n1520 gnd 0.005139f
C3761 vdd.n1521 gnd 0.005155f
C3762 vdd.t155 gnd 0.014721f
C3763 vdd.n1522 gnd 0.032755f
C3764 vdd.n1523 gnd 0.170464f
C3765 vdd.n1524 gnd 0.002899f
C3766 vdd.n1525 gnd 0.00307f
C3767 vdd.n1526 gnd 0.006852f
C3768 vdd.n1527 gnd 0.006852f
C3769 vdd.n1528 gnd 0.00307f
C3770 vdd.n1529 gnd 0.002899f
C3771 vdd.n1530 gnd 0.005395f
C3772 vdd.n1531 gnd 0.005395f
C3773 vdd.n1532 gnd 0.002899f
C3774 vdd.n1533 gnd 0.00307f
C3775 vdd.n1534 gnd 0.006852f
C3776 vdd.n1535 gnd 0.006852f
C3777 vdd.n1536 gnd 0.00307f
C3778 vdd.n1537 gnd 0.002899f
C3779 vdd.n1538 gnd 0.005395f
C3780 vdd.n1539 gnd 0.005395f
C3781 vdd.n1540 gnd 0.002899f
C3782 vdd.n1541 gnd 0.00307f
C3783 vdd.n1542 gnd 0.006852f
C3784 vdd.n1543 gnd 0.006852f
C3785 vdd.n1544 gnd 0.0162f
C3786 vdd.n1545 gnd 0.002984f
C3787 vdd.n1546 gnd 0.002899f
C3788 vdd.n1547 gnd 0.013944f
C3789 vdd.n1548 gnd 0.00943f
C3790 vdd.n1549 gnd 0.110667f
C3791 vdd.n1550 gnd 0.005814f
C3792 vdd.n1551 gnd 0.005395f
C3793 vdd.n1552 gnd 0.002984f
C3794 vdd.n1553 gnd 0.006852f
C3795 vdd.n1554 gnd 0.002899f
C3796 vdd.n1555 gnd 0.00307f
C3797 vdd.n1556 gnd 0.005395f
C3798 vdd.n1557 gnd 0.002899f
C3799 vdd.n1558 gnd 0.006852f
C3800 vdd.n1559 gnd 0.00307f
C3801 vdd.n1560 gnd 0.005395f
C3802 vdd.n1561 gnd 0.002899f
C3803 vdd.n1562 gnd 0.005139f
C3804 vdd.n1563 gnd 0.005155f
C3805 vdd.t234 gnd 0.014721f
C3806 vdd.n1564 gnd 0.032755f
C3807 vdd.n1565 gnd 0.170464f
C3808 vdd.n1566 gnd 0.002899f
C3809 vdd.n1567 gnd 0.00307f
C3810 vdd.n1568 gnd 0.006852f
C3811 vdd.n1569 gnd 0.006852f
C3812 vdd.n1570 gnd 0.00307f
C3813 vdd.n1571 gnd 0.002899f
C3814 vdd.n1572 gnd 0.005395f
C3815 vdd.n1573 gnd 0.005395f
C3816 vdd.n1574 gnd 0.002899f
C3817 vdd.n1575 gnd 0.00307f
C3818 vdd.n1576 gnd 0.006852f
C3819 vdd.n1577 gnd 0.006852f
C3820 vdd.n1578 gnd 0.00307f
C3821 vdd.n1579 gnd 0.002899f
C3822 vdd.n1580 gnd 0.005395f
C3823 vdd.n1581 gnd 0.005395f
C3824 vdd.n1582 gnd 0.002899f
C3825 vdd.n1583 gnd 0.00307f
C3826 vdd.n1584 gnd 0.006852f
C3827 vdd.n1585 gnd 0.006852f
C3828 vdd.n1586 gnd 0.0162f
C3829 vdd.n1587 gnd 0.002984f
C3830 vdd.n1588 gnd 0.002899f
C3831 vdd.n1589 gnd 0.013944f
C3832 vdd.n1590 gnd 0.009735f
C3833 vdd.t145 gnd 0.034106f
C3834 vdd.t237 gnd 0.034106f
C3835 vdd.n1591 gnd 0.2344f
C3836 vdd.n1592 gnd 0.18432f
C3837 vdd.t228 gnd 0.034106f
C3838 vdd.t217 gnd 0.034106f
C3839 vdd.n1593 gnd 0.2344f
C3840 vdd.n1594 gnd 0.148745f
C3841 vdd.t189 gnd 0.034106f
C3842 vdd.t139 gnd 0.034106f
C3843 vdd.n1595 gnd 0.2344f
C3844 vdd.n1596 gnd 0.148745f
C3845 vdd.t245 gnd 0.034106f
C3846 vdd.t215 gnd 0.034106f
C3847 vdd.n1597 gnd 0.2344f
C3848 vdd.n1598 gnd 0.148745f
C3849 vdd.t212 gnd 0.034106f
C3850 vdd.t167 gnd 0.034106f
C3851 vdd.n1599 gnd 0.2344f
C3852 vdd.n1600 gnd 0.148745f
C3853 vdd.t161 gnd 0.034106f
C3854 vdd.t213 gnd 0.034106f
C3855 vdd.n1601 gnd 0.2344f
C3856 vdd.n1602 gnd 0.148745f
C3857 vdd.t203 gnd 0.034106f
C3858 vdd.t201 gnd 0.034106f
C3859 vdd.n1603 gnd 0.2344f
C3860 vdd.n1604 gnd 0.148745f
C3861 vdd.n1605 gnd 0.005814f
C3862 vdd.n1606 gnd 0.005395f
C3863 vdd.n1607 gnd 0.002984f
C3864 vdd.n1608 gnd 0.006852f
C3865 vdd.n1609 gnd 0.002899f
C3866 vdd.n1610 gnd 0.00307f
C3867 vdd.n1611 gnd 0.005395f
C3868 vdd.n1612 gnd 0.002899f
C3869 vdd.n1613 gnd 0.006852f
C3870 vdd.n1614 gnd 0.00307f
C3871 vdd.n1615 gnd 0.005395f
C3872 vdd.n1616 gnd 0.002899f
C3873 vdd.n1617 gnd 0.005139f
C3874 vdd.n1618 gnd 0.005155f
C3875 vdd.t141 gnd 0.014721f
C3876 vdd.n1619 gnd 0.032755f
C3877 vdd.n1620 gnd 0.170464f
C3878 vdd.n1621 gnd 0.002899f
C3879 vdd.n1622 gnd 0.00307f
C3880 vdd.n1623 gnd 0.006852f
C3881 vdd.n1624 gnd 0.006852f
C3882 vdd.n1625 gnd 0.00307f
C3883 vdd.n1626 gnd 0.002899f
C3884 vdd.n1627 gnd 0.005395f
C3885 vdd.n1628 gnd 0.005395f
C3886 vdd.n1629 gnd 0.002899f
C3887 vdd.n1630 gnd 0.00307f
C3888 vdd.n1631 gnd 0.006852f
C3889 vdd.n1632 gnd 0.006852f
C3890 vdd.n1633 gnd 0.00307f
C3891 vdd.n1634 gnd 0.002899f
C3892 vdd.n1635 gnd 0.005395f
C3893 vdd.n1636 gnd 0.005395f
C3894 vdd.n1637 gnd 0.002899f
C3895 vdd.n1638 gnd 0.00307f
C3896 vdd.n1639 gnd 0.006852f
C3897 vdd.n1640 gnd 0.006852f
C3898 vdd.n1641 gnd 0.0162f
C3899 vdd.n1642 gnd 0.002984f
C3900 vdd.n1643 gnd 0.002899f
C3901 vdd.n1644 gnd 0.013944f
C3902 vdd.n1645 gnd 0.00943f
C3903 vdd.n1646 gnd 0.065836f
C3904 vdd.n1647 gnd 0.237223f
C3905 vdd.n1648 gnd 0.005814f
C3906 vdd.n1649 gnd 0.005395f
C3907 vdd.n1650 gnd 0.002984f
C3908 vdd.n1651 gnd 0.006852f
C3909 vdd.n1652 gnd 0.002899f
C3910 vdd.n1653 gnd 0.00307f
C3911 vdd.n1654 gnd 0.005395f
C3912 vdd.n1655 gnd 0.002899f
C3913 vdd.n1656 gnd 0.006852f
C3914 vdd.n1657 gnd 0.00307f
C3915 vdd.n1658 gnd 0.005395f
C3916 vdd.n1659 gnd 0.002899f
C3917 vdd.n1660 gnd 0.005139f
C3918 vdd.n1661 gnd 0.005155f
C3919 vdd.t246 gnd 0.014721f
C3920 vdd.n1662 gnd 0.032755f
C3921 vdd.n1663 gnd 0.170464f
C3922 vdd.n1664 gnd 0.002899f
C3923 vdd.n1665 gnd 0.00307f
C3924 vdd.n1666 gnd 0.006852f
C3925 vdd.n1667 gnd 0.006852f
C3926 vdd.n1668 gnd 0.00307f
C3927 vdd.n1669 gnd 0.002899f
C3928 vdd.n1670 gnd 0.005395f
C3929 vdd.n1671 gnd 0.005395f
C3930 vdd.n1672 gnd 0.002899f
C3931 vdd.n1673 gnd 0.00307f
C3932 vdd.n1674 gnd 0.006852f
C3933 vdd.n1675 gnd 0.006852f
C3934 vdd.n1676 gnd 0.00307f
C3935 vdd.n1677 gnd 0.002899f
C3936 vdd.n1678 gnd 0.005395f
C3937 vdd.n1679 gnd 0.005395f
C3938 vdd.n1680 gnd 0.002899f
C3939 vdd.n1681 gnd 0.00307f
C3940 vdd.n1682 gnd 0.006852f
C3941 vdd.n1683 gnd 0.006852f
C3942 vdd.n1684 gnd 0.0162f
C3943 vdd.n1685 gnd 0.002984f
C3944 vdd.n1686 gnd 0.002899f
C3945 vdd.n1687 gnd 0.013944f
C3946 vdd.n1688 gnd 0.009735f
C3947 vdd.t159 gnd 0.034106f
C3948 vdd.t247 gnd 0.034106f
C3949 vdd.n1689 gnd 0.2344f
C3950 vdd.n1690 gnd 0.18432f
C3951 vdd.t244 gnd 0.034106f
C3952 vdd.t229 gnd 0.034106f
C3953 vdd.n1691 gnd 0.2344f
C3954 vdd.n1692 gnd 0.148745f
C3955 vdd.t204 gnd 0.034106f
C3956 vdd.t156 gnd 0.034106f
C3957 vdd.n1693 gnd 0.2344f
C3958 vdd.n1694 gnd 0.148745f
C3959 vdd.t255 gnd 0.034106f
C3960 vdd.t225 gnd 0.034106f
C3961 vdd.n1695 gnd 0.2344f
C3962 vdd.n1696 gnd 0.148745f
C3963 vdd.t222 gnd 0.034106f
C3964 vdd.t181 gnd 0.034106f
C3965 vdd.n1697 gnd 0.2344f
C3966 vdd.n1698 gnd 0.148745f
C3967 vdd.t180 gnd 0.034106f
C3968 vdd.t223 gnd 0.034106f
C3969 vdd.n1699 gnd 0.2344f
C3970 vdd.n1700 gnd 0.148745f
C3971 vdd.t211 gnd 0.034106f
C3972 vdd.t210 gnd 0.034106f
C3973 vdd.n1701 gnd 0.2344f
C3974 vdd.n1702 gnd 0.148745f
C3975 vdd.n1703 gnd 0.005814f
C3976 vdd.n1704 gnd 0.005395f
C3977 vdd.n1705 gnd 0.002984f
C3978 vdd.n1706 gnd 0.006852f
C3979 vdd.n1707 gnd 0.002899f
C3980 vdd.n1708 gnd 0.00307f
C3981 vdd.n1709 gnd 0.005395f
C3982 vdd.n1710 gnd 0.002899f
C3983 vdd.n1711 gnd 0.006852f
C3984 vdd.n1712 gnd 0.00307f
C3985 vdd.n1713 gnd 0.005395f
C3986 vdd.n1714 gnd 0.002899f
C3987 vdd.n1715 gnd 0.005139f
C3988 vdd.n1716 gnd 0.005155f
C3989 vdd.t158 gnd 0.014721f
C3990 vdd.n1717 gnd 0.032755f
C3991 vdd.n1718 gnd 0.170464f
C3992 vdd.n1719 gnd 0.002899f
C3993 vdd.n1720 gnd 0.00307f
C3994 vdd.n1721 gnd 0.006852f
C3995 vdd.n1722 gnd 0.006852f
C3996 vdd.n1723 gnd 0.00307f
C3997 vdd.n1724 gnd 0.002899f
C3998 vdd.n1725 gnd 0.005395f
C3999 vdd.n1726 gnd 0.005395f
C4000 vdd.n1727 gnd 0.002899f
C4001 vdd.n1728 gnd 0.00307f
C4002 vdd.n1729 gnd 0.006852f
C4003 vdd.n1730 gnd 0.006852f
C4004 vdd.n1731 gnd 0.00307f
C4005 vdd.n1732 gnd 0.002899f
C4006 vdd.n1733 gnd 0.005395f
C4007 vdd.n1734 gnd 0.005395f
C4008 vdd.n1735 gnd 0.002899f
C4009 vdd.n1736 gnd 0.00307f
C4010 vdd.n1737 gnd 0.006852f
C4011 vdd.n1738 gnd 0.006852f
C4012 vdd.n1739 gnd 0.0162f
C4013 vdd.n1740 gnd 0.002984f
C4014 vdd.n1741 gnd 0.002899f
C4015 vdd.n1742 gnd 0.013944f
C4016 vdd.n1743 gnd 0.00943f
C4017 vdd.n1744 gnd 0.065836f
C4018 vdd.n1745 gnd 0.265659f
C4019 vdd.n1746 gnd 2.53412f
C4020 vdd.n1747 gnd 0.624846f
C4021 vdd.n1748 gnd 0.008142f
C4022 vdd.n1749 gnd 0.010593f
C4023 vdd.n1750 gnd 0.008527f
C4024 vdd.n1751 gnd 0.010593f
C4025 vdd.n1752 gnd 0.849847f
C4026 vdd.n1753 gnd 0.010593f
C4027 vdd.n1754 gnd 0.008527f
C4028 vdd.n1755 gnd 0.010593f
C4029 vdd.n1756 gnd 0.010593f
C4030 vdd.n1757 gnd 0.010593f
C4031 vdd.n1758 gnd 0.008527f
C4032 vdd.n1759 gnd 0.010593f
C4033 vdd.t138 gnd 0.541304f
C4034 vdd.n1760 gnd 0.898564f
C4035 vdd.n1761 gnd 0.010593f
C4036 vdd.n1762 gnd 0.008527f
C4037 vdd.n1763 gnd 0.010593f
C4038 vdd.n1764 gnd 0.010593f
C4039 vdd.n1765 gnd 0.010593f
C4040 vdd.n1766 gnd 0.008527f
C4041 vdd.n1767 gnd 0.010593f
C4042 vdd.n1768 gnd 0.763238f
C4043 vdd.n1769 gnd 0.010593f
C4044 vdd.n1770 gnd 0.008527f
C4045 vdd.n1771 gnd 0.010593f
C4046 vdd.n1772 gnd 0.010593f
C4047 vdd.n1773 gnd 0.010593f
C4048 vdd.n1774 gnd 0.008527f
C4049 vdd.n1775 gnd 0.010593f
C4050 vdd.n1776 gnd 0.898564f
C4051 vdd.t216 gnd 0.541304f
C4052 vdd.n1777 gnd 0.579195f
C4053 vdd.n1778 gnd 0.010593f
C4054 vdd.n1779 gnd 0.008527f
C4055 vdd.n1780 gnd 0.010593f
C4056 vdd.n1781 gnd 0.010593f
C4057 vdd.n1782 gnd 0.010593f
C4058 vdd.n1783 gnd 0.008527f
C4059 vdd.n1784 gnd 0.010593f
C4060 vdd.n1785 gnd 0.687456f
C4061 vdd.n1786 gnd 0.010593f
C4062 vdd.n1787 gnd 0.008527f
C4063 vdd.n1788 gnd 0.010593f
C4064 vdd.n1789 gnd 0.010593f
C4065 vdd.n1790 gnd 0.010593f
C4066 vdd.n1791 gnd 0.008527f
C4067 vdd.n1792 gnd 0.010593f
C4068 vdd.n1793 gnd 0.568369f
C4069 vdd.n1794 gnd 0.871499f
C4070 vdd.n1795 gnd 0.010593f
C4071 vdd.n1796 gnd 0.008527f
C4072 vdd.n1797 gnd 0.010593f
C4073 vdd.n1798 gnd 0.010593f
C4074 vdd.n1799 gnd 0.010593f
C4075 vdd.n1800 gnd 0.008527f
C4076 vdd.n1801 gnd 0.010593f
C4077 vdd.n1802 gnd 1.05554f
C4078 vdd.n1803 gnd 0.010593f
C4079 vdd.n1804 gnd 0.008527f
C4080 vdd.n1805 gnd 0.010593f
C4081 vdd.n1806 gnd 0.010593f
C4082 vdd.n1807 gnd 0.024124f
C4083 vdd.n1808 gnd 0.010593f
C4084 vdd.n1809 gnd 0.010593f
C4085 vdd.n1810 gnd 0.008527f
C4086 vdd.n1811 gnd 0.010593f
C4087 vdd.t43 gnd 0.541304f
C4088 vdd.n1812 gnd 1.02306f
C4089 vdd.n1813 gnd 0.010593f
C4090 vdd.n1814 gnd 0.008527f
C4091 vdd.n1815 gnd 0.010593f
C4092 vdd.n1816 gnd 0.010593f
C4093 vdd.n1817 gnd 0.00911f
C4094 vdd.n1818 gnd 0.008527f
C4095 vdd.n1820 gnd 0.010593f
C4096 vdd.n1822 gnd 0.008527f
C4097 vdd.n1823 gnd 0.010593f
C4098 vdd.n1824 gnd 0.008527f
C4099 vdd.n1826 gnd 0.010593f
C4100 vdd.n1827 gnd 0.008527f
C4101 vdd.n1828 gnd 0.010593f
C4102 vdd.n1829 gnd 0.010593f
C4103 vdd.n1830 gnd 0.010593f
C4104 vdd.n1831 gnd 0.010593f
C4105 vdd.n1832 gnd 0.010593f
C4106 vdd.n1833 gnd 0.008527f
C4107 vdd.n1835 gnd 0.010593f
C4108 vdd.n1836 gnd 0.010593f
C4109 vdd.n1837 gnd 0.010593f
C4110 vdd.n1838 gnd 0.010593f
C4111 vdd.n1839 gnd 0.010593f
C4112 vdd.n1840 gnd 0.008527f
C4113 vdd.n1842 gnd 0.010593f
C4114 vdd.n1843 gnd 0.010593f
C4115 vdd.n1844 gnd 0.010593f
C4116 vdd.n1845 gnd 0.010593f
C4117 vdd.n1846 gnd 0.00712f
C4118 vdd.t61 gnd 0.130328f
C4119 vdd.t60 gnd 0.139285f
C4120 vdd.t59 gnd 0.170207f
C4121 vdd.n1847 gnd 0.218181f
C4122 vdd.n1848 gnd 0.183312f
C4123 vdd.n1850 gnd 0.010593f
C4124 vdd.n1851 gnd 0.010593f
C4125 vdd.n1852 gnd 0.008527f
C4126 vdd.n1853 gnd 0.010593f
C4127 vdd.n1855 gnd 0.010593f
C4128 vdd.n1856 gnd 0.010593f
C4129 vdd.n1857 gnd 0.010593f
C4130 vdd.n1858 gnd 0.010593f
C4131 vdd.n1859 gnd 0.008527f
C4132 vdd.n1861 gnd 0.010593f
C4133 vdd.n1862 gnd 0.010593f
C4134 vdd.n1863 gnd 0.010593f
C4135 vdd.n1864 gnd 0.010593f
C4136 vdd.n1865 gnd 0.010593f
C4137 vdd.n1866 gnd 0.008527f
C4138 vdd.n1868 gnd 0.010593f
C4139 vdd.n1869 gnd 0.010593f
C4140 vdd.n1870 gnd 0.010593f
C4141 vdd.n1871 gnd 0.010593f
C4142 vdd.n1872 gnd 0.010593f
C4143 vdd.n1873 gnd 0.008527f
C4144 vdd.n1875 gnd 0.010593f
C4145 vdd.n1876 gnd 0.010593f
C4146 vdd.n1877 gnd 0.010593f
C4147 vdd.n1878 gnd 0.010593f
C4148 vdd.n1879 gnd 0.010593f
C4149 vdd.n1880 gnd 0.008527f
C4150 vdd.n1882 gnd 0.010593f
C4151 vdd.n1883 gnd 0.010593f
C4152 vdd.n1884 gnd 0.010593f
C4153 vdd.n1885 gnd 0.010593f
C4154 vdd.n1886 gnd 0.008441f
C4155 vdd.t58 gnd 0.130328f
C4156 vdd.t57 gnd 0.139285f
C4157 vdd.t56 gnd 0.170207f
C4158 vdd.n1887 gnd 0.218181f
C4159 vdd.n1888 gnd 0.183312f
C4160 vdd.n1890 gnd 0.010593f
C4161 vdd.n1891 gnd 0.010593f
C4162 vdd.n1892 gnd 0.008527f
C4163 vdd.n1893 gnd 0.010593f
C4164 vdd.n1895 gnd 0.010593f
C4165 vdd.n1896 gnd 0.010593f
C4166 vdd.n1897 gnd 0.010593f
C4167 vdd.n1898 gnd 0.010593f
C4168 vdd.n1899 gnd 0.008527f
C4169 vdd.n1901 gnd 0.010593f
C4170 vdd.n1902 gnd 0.010593f
C4171 vdd.n1903 gnd 0.010593f
C4172 vdd.n1904 gnd 0.010593f
C4173 vdd.n1905 gnd 0.010593f
C4174 vdd.n1906 gnd 0.008527f
C4175 vdd.n1908 gnd 0.010593f
C4176 vdd.n1909 gnd 0.010593f
C4177 vdd.n1910 gnd 0.010593f
C4178 vdd.n1911 gnd 0.010593f
C4179 vdd.n1912 gnd 0.010593f
C4180 vdd.n1913 gnd 0.010593f
C4181 vdd.n1914 gnd 0.008527f
C4182 vdd.n1916 gnd 0.010593f
C4183 vdd.n1918 gnd 0.010593f
C4184 vdd.n1919 gnd 0.008527f
C4185 vdd.n1920 gnd 0.008527f
C4186 vdd.n1921 gnd 0.010593f
C4187 vdd.n1923 gnd 0.010593f
C4188 vdd.n1924 gnd 0.008527f
C4189 vdd.n1925 gnd 0.008527f
C4190 vdd.n1926 gnd 0.010593f
C4191 vdd.n1928 gnd 0.010593f
C4192 vdd.n1929 gnd 0.010593f
C4193 vdd.n1930 gnd 0.008527f
C4194 vdd.n1931 gnd 0.008527f
C4195 vdd.n1932 gnd 0.008527f
C4196 vdd.n1933 gnd 0.010593f
C4197 vdd.n1935 gnd 0.010593f
C4198 vdd.n1936 gnd 0.010593f
C4199 vdd.n1937 gnd 0.008527f
C4200 vdd.n1938 gnd 0.008527f
C4201 vdd.n1939 gnd 0.008527f
C4202 vdd.n1940 gnd 0.010593f
C4203 vdd.n1942 gnd 0.010593f
C4204 vdd.n1943 gnd 0.010593f
C4205 vdd.n1944 gnd 0.008527f
C4206 vdd.n1945 gnd 0.008527f
C4207 vdd.n1946 gnd 0.008527f
C4208 vdd.n1947 gnd 0.010593f
C4209 vdd.n1949 gnd 0.010593f
C4210 vdd.n1950 gnd 0.010593f
C4211 vdd.n1951 gnd 0.008527f
C4212 vdd.n1952 gnd 0.010593f
C4213 vdd.n1953 gnd 0.010593f
C4214 vdd.n1954 gnd 0.010593f
C4215 vdd.n1955 gnd 0.017394f
C4216 vdd.n1956 gnd 0.005798f
C4217 vdd.n1957 gnd 0.008527f
C4218 vdd.n1958 gnd 0.010593f
C4219 vdd.n1960 gnd 0.010593f
C4220 vdd.n1961 gnd 0.010593f
C4221 vdd.n1962 gnd 0.008527f
C4222 vdd.n1963 gnd 0.008527f
C4223 vdd.n1964 gnd 0.008527f
C4224 vdd.n1965 gnd 0.010593f
C4225 vdd.n1967 gnd 0.010593f
C4226 vdd.n1968 gnd 0.010593f
C4227 vdd.n1969 gnd 0.008527f
C4228 vdd.n1970 gnd 0.008527f
C4229 vdd.n1971 gnd 0.008527f
C4230 vdd.n1972 gnd 0.010593f
C4231 vdd.n1974 gnd 0.010593f
C4232 vdd.n1975 gnd 0.010593f
C4233 vdd.n1976 gnd 0.008527f
C4234 vdd.n1977 gnd 0.008527f
C4235 vdd.n1978 gnd 0.008527f
C4236 vdd.n1979 gnd 0.010593f
C4237 vdd.n1981 gnd 0.010593f
C4238 vdd.n1982 gnd 0.010593f
C4239 vdd.n1983 gnd 0.008527f
C4240 vdd.n1984 gnd 0.008527f
C4241 vdd.n1985 gnd 0.008527f
C4242 vdd.n1986 gnd 0.010593f
C4243 vdd.n1988 gnd 0.010593f
C4244 vdd.n1989 gnd 0.010593f
C4245 vdd.n1990 gnd 0.008527f
C4246 vdd.n1991 gnd 0.010593f
C4247 vdd.n1992 gnd 0.010593f
C4248 vdd.n1993 gnd 0.010593f
C4249 vdd.n1994 gnd 0.017394f
C4250 vdd.n1995 gnd 0.00712f
C4251 vdd.n1996 gnd 0.008527f
C4252 vdd.n1997 gnd 0.010593f
C4253 vdd.n1999 gnd 0.010593f
C4254 vdd.n2000 gnd 0.010593f
C4255 vdd.n2001 gnd 0.008527f
C4256 vdd.n2002 gnd 0.008527f
C4257 vdd.n2003 gnd 0.008527f
C4258 vdd.n2004 gnd 0.010593f
C4259 vdd.n2006 gnd 0.010593f
C4260 vdd.n2007 gnd 0.010593f
C4261 vdd.n2008 gnd 0.008527f
C4262 vdd.n2009 gnd 0.008527f
C4263 vdd.n2010 gnd 0.008527f
C4264 vdd.n2011 gnd 0.010593f
C4265 vdd.n2013 gnd 0.010593f
C4266 vdd.n2014 gnd 0.010593f
C4267 vdd.n2016 gnd 0.010593f
C4268 vdd.n2017 gnd 0.008527f
C4269 vdd.n2018 gnd 0.00678f
C4270 vdd.n2019 gnd 0.007204f
C4271 vdd.n2020 gnd 0.007204f
C4272 vdd.n2021 gnd 0.007204f
C4273 vdd.n2022 gnd 0.007204f
C4274 vdd.n2023 gnd 0.007204f
C4275 vdd.n2024 gnd 0.007204f
C4276 vdd.n2025 gnd 0.007204f
C4277 vdd.n2026 gnd 0.007204f
C4278 vdd.n2028 gnd 0.007204f
C4279 vdd.n2029 gnd 0.007204f
C4280 vdd.n2030 gnd 0.007204f
C4281 vdd.n2031 gnd 0.007204f
C4282 vdd.n2032 gnd 0.007204f
C4283 vdd.n2034 gnd 0.007204f
C4284 vdd.n2036 gnd 0.007204f
C4285 vdd.n2037 gnd 0.007204f
C4286 vdd.n2038 gnd 0.007204f
C4287 vdd.n2039 gnd 0.007204f
C4288 vdd.n2040 gnd 0.007204f
C4289 vdd.n2042 gnd 0.007204f
C4290 vdd.n2044 gnd 0.007204f
C4291 vdd.n2045 gnd 0.007204f
C4292 vdd.n2046 gnd 0.007204f
C4293 vdd.n2047 gnd 0.007204f
C4294 vdd.n2048 gnd 0.007204f
C4295 vdd.n2050 gnd 0.007204f
C4296 vdd.n2052 gnd 0.007204f
C4297 vdd.n2053 gnd 0.007204f
C4298 vdd.n2054 gnd 0.007204f
C4299 vdd.n2055 gnd 0.007204f
C4300 vdd.n2056 gnd 0.007204f
C4301 vdd.n2058 gnd 0.007204f
C4302 vdd.n2059 gnd 0.007204f
C4303 vdd.n2060 gnd 0.007204f
C4304 vdd.n2061 gnd 0.007204f
C4305 vdd.n2062 gnd 0.007204f
C4306 vdd.n2063 gnd 0.007204f
C4307 vdd.n2064 gnd 0.007204f
C4308 vdd.n2065 gnd 0.007204f
C4309 vdd.n2066 gnd 0.005244f
C4310 vdd.n2067 gnd 0.007204f
C4311 vdd.t25 gnd 0.291096f
C4312 vdd.t26 gnd 0.297973f
C4313 vdd.t23 gnd 0.190039f
C4314 vdd.n2068 gnd 0.102706f
C4315 vdd.n2069 gnd 0.058258f
C4316 vdd.n2070 gnd 0.010295f
C4317 vdd.n2071 gnd 0.007204f
C4318 vdd.n2072 gnd 0.007204f
C4319 vdd.n2073 gnd 0.438456f
C4320 vdd.n2074 gnd 0.007204f
C4321 vdd.n2075 gnd 0.007204f
C4322 vdd.n2076 gnd 0.007204f
C4323 vdd.n2077 gnd 0.007204f
C4324 vdd.n2078 gnd 0.007204f
C4325 vdd.n2079 gnd 0.007204f
C4326 vdd.n2080 gnd 0.007204f
C4327 vdd.n2081 gnd 0.007204f
C4328 vdd.n2082 gnd 0.007204f
C4329 vdd.n2083 gnd 0.007204f
C4330 vdd.n2084 gnd 0.007204f
C4331 vdd.n2085 gnd 0.007204f
C4332 vdd.n2086 gnd 0.007204f
C4333 vdd.n2087 gnd 0.007204f
C4334 vdd.n2088 gnd 0.007204f
C4335 vdd.n2089 gnd 0.007204f
C4336 vdd.n2090 gnd 0.007204f
C4337 vdd.n2091 gnd 0.007204f
C4338 vdd.n2092 gnd 0.007204f
C4339 vdd.n2093 gnd 0.007204f
C4340 vdd.t78 gnd 0.291096f
C4341 vdd.t79 gnd 0.297973f
C4342 vdd.t77 gnd 0.190039f
C4343 vdd.n2094 gnd 0.102706f
C4344 vdd.n2095 gnd 0.058258f
C4345 vdd.n2096 gnd 0.007204f
C4346 vdd.n2097 gnd 0.007204f
C4347 vdd.n2098 gnd 0.007204f
C4348 vdd.n2099 gnd 0.007204f
C4349 vdd.n2100 gnd 0.007204f
C4350 vdd.n2101 gnd 0.007204f
C4351 vdd.n2103 gnd 0.007204f
C4352 vdd.n2104 gnd 0.007204f
C4353 vdd.n2105 gnd 0.007204f
C4354 vdd.n2106 gnd 0.007204f
C4355 vdd.n2108 gnd 0.007204f
C4356 vdd.n2110 gnd 0.007204f
C4357 vdd.n2111 gnd 0.007204f
C4358 vdd.n2112 gnd 0.007204f
C4359 vdd.n2113 gnd 0.007204f
C4360 vdd.n2114 gnd 0.007204f
C4361 vdd.n2116 gnd 0.007204f
C4362 vdd.n2118 gnd 0.007204f
C4363 vdd.n2119 gnd 0.007204f
C4364 vdd.n2120 gnd 0.007204f
C4365 vdd.n2121 gnd 0.007204f
C4366 vdd.n2122 gnd 0.007204f
C4367 vdd.n2124 gnd 0.007204f
C4368 vdd.n2126 gnd 0.007204f
C4369 vdd.n2127 gnd 0.007204f
C4370 vdd.n2128 gnd 0.005244f
C4371 vdd.n2129 gnd 0.010295f
C4372 vdd.n2130 gnd 0.005562f
C4373 vdd.n2131 gnd 0.007204f
C4374 vdd.n2133 gnd 0.007204f
C4375 vdd.n2134 gnd 0.017093f
C4376 vdd.n2135 gnd 0.017093f
C4377 vdd.n2136 gnd 0.015959f
C4378 vdd.n2137 gnd 0.007204f
C4379 vdd.n2138 gnd 0.007204f
C4380 vdd.n2139 gnd 0.007204f
C4381 vdd.n2140 gnd 0.007204f
C4382 vdd.n2141 gnd 0.007204f
C4383 vdd.n2142 gnd 0.007204f
C4384 vdd.n2143 gnd 0.007204f
C4385 vdd.n2144 gnd 0.007204f
C4386 vdd.n2145 gnd 0.007204f
C4387 vdd.n2146 gnd 0.007204f
C4388 vdd.n2147 gnd 0.007204f
C4389 vdd.n2148 gnd 0.007204f
C4390 vdd.n2149 gnd 0.007204f
C4391 vdd.n2150 gnd 0.007204f
C4392 vdd.n2151 gnd 0.007204f
C4393 vdd.n2152 gnd 0.007204f
C4394 vdd.n2153 gnd 0.007204f
C4395 vdd.n2154 gnd 0.007204f
C4396 vdd.n2155 gnd 0.007204f
C4397 vdd.n2156 gnd 0.007204f
C4398 vdd.n2157 gnd 0.007204f
C4399 vdd.n2158 gnd 0.007204f
C4400 vdd.n2159 gnd 0.007204f
C4401 vdd.n2160 gnd 0.007204f
C4402 vdd.n2161 gnd 0.007204f
C4403 vdd.n2162 gnd 0.007204f
C4404 vdd.n2163 gnd 0.007204f
C4405 vdd.n2164 gnd 0.007204f
C4406 vdd.n2165 gnd 0.007204f
C4407 vdd.n2166 gnd 0.007204f
C4408 vdd.n2167 gnd 0.007204f
C4409 vdd.n2168 gnd 0.007204f
C4410 vdd.n2169 gnd 0.007204f
C4411 vdd.n2170 gnd 0.007204f
C4412 vdd.n2171 gnd 0.007204f
C4413 vdd.n2172 gnd 0.007204f
C4414 vdd.n2173 gnd 0.007204f
C4415 vdd.n2174 gnd 0.232761f
C4416 vdd.n2175 gnd 0.007204f
C4417 vdd.n2176 gnd 0.007204f
C4418 vdd.n2177 gnd 0.007204f
C4419 vdd.n2178 gnd 0.007204f
C4420 vdd.n2179 gnd 0.007204f
C4421 vdd.n2180 gnd 0.007204f
C4422 vdd.n2181 gnd 0.007204f
C4423 vdd.n2182 gnd 0.007204f
C4424 vdd.n2183 gnd 0.007204f
C4425 vdd.n2184 gnd 0.007204f
C4426 vdd.n2185 gnd 0.007204f
C4427 vdd.n2186 gnd 0.007204f
C4428 vdd.n2187 gnd 0.007204f
C4429 vdd.n2188 gnd 0.007204f
C4430 vdd.n2189 gnd 0.007204f
C4431 vdd.n2190 gnd 0.007204f
C4432 vdd.n2191 gnd 0.007204f
C4433 vdd.n2192 gnd 0.007204f
C4434 vdd.n2193 gnd 0.007204f
C4435 vdd.n2194 gnd 0.007204f
C4436 vdd.n2195 gnd 0.015959f
C4437 vdd.n2197 gnd 0.017093f
C4438 vdd.n2198 gnd 0.017093f
C4439 vdd.n2199 gnd 0.007204f
C4440 vdd.n2200 gnd 0.005562f
C4441 vdd.n2201 gnd 0.007204f
C4442 vdd.n2203 gnd 0.007204f
C4443 vdd.n2205 gnd 0.007204f
C4444 vdd.n2206 gnd 0.007204f
C4445 vdd.n2207 gnd 0.007204f
C4446 vdd.n2208 gnd 0.007204f
C4447 vdd.n2209 gnd 0.007204f
C4448 vdd.n2211 gnd 0.007204f
C4449 vdd.n2213 gnd 0.007204f
C4450 vdd.n2214 gnd 0.007204f
C4451 vdd.n2215 gnd 0.007204f
C4452 vdd.n2216 gnd 0.007204f
C4453 vdd.n2217 gnd 0.007204f
C4454 vdd.n2219 gnd 0.007204f
C4455 vdd.n2221 gnd 0.007204f
C4456 vdd.n2222 gnd 0.007204f
C4457 vdd.n2223 gnd 0.007204f
C4458 vdd.n2224 gnd 0.007204f
C4459 vdd.n2225 gnd 0.007204f
C4460 vdd.n2227 gnd 0.007204f
C4461 vdd.n2229 gnd 0.007204f
C4462 vdd.n2230 gnd 0.007204f
C4463 vdd.n2231 gnd 0.021487f
C4464 vdd.n2232 gnd 0.636961f
C4465 vdd.n2234 gnd 0.008527f
C4466 vdd.n2235 gnd 0.008527f
C4467 vdd.n2236 gnd 0.010593f
C4468 vdd.n2238 gnd 0.010593f
C4469 vdd.n2239 gnd 0.010593f
C4470 vdd.n2240 gnd 0.008527f
C4471 vdd.n2241 gnd 0.007077f
C4472 vdd.n2242 gnd 0.024289f
C4473 vdd.n2243 gnd 0.024124f
C4474 vdd.n2244 gnd 0.007077f
C4475 vdd.n2245 gnd 0.024124f
C4476 vdd.n2246 gnd 1.42904f
C4477 vdd.n2247 gnd 0.024124f
C4478 vdd.n2248 gnd 0.024289f
C4479 vdd.n2249 gnd 0.00405f
C4480 vdd.t45 gnd 0.130328f
C4481 vdd.t44 gnd 0.139285f
C4482 vdd.t42 gnd 0.170207f
C4483 vdd.n2250 gnd 0.218181f
C4484 vdd.n2251 gnd 0.183312f
C4485 vdd.n2252 gnd 0.013131f
C4486 vdd.n2253 gnd 0.004476f
C4487 vdd.n2254 gnd 0.00911f
C4488 vdd.n2255 gnd 0.636961f
C4489 vdd.n2256 gnd 0.021487f
C4490 vdd.n2257 gnd 0.007204f
C4491 vdd.n2258 gnd 0.007204f
C4492 vdd.n2259 gnd 0.007204f
C4493 vdd.n2261 gnd 0.007204f
C4494 vdd.n2263 gnd 0.007204f
C4495 vdd.n2264 gnd 0.007204f
C4496 vdd.n2265 gnd 0.007204f
C4497 vdd.n2266 gnd 0.007204f
C4498 vdd.n2267 gnd 0.007204f
C4499 vdd.n2269 gnd 0.007204f
C4500 vdd.n2271 gnd 0.007204f
C4501 vdd.n2272 gnd 0.007204f
C4502 vdd.n2273 gnd 0.007204f
C4503 vdd.n2274 gnd 0.007204f
C4504 vdd.n2275 gnd 0.007204f
C4505 vdd.n2277 gnd 0.007204f
C4506 vdd.n2279 gnd 0.007204f
C4507 vdd.n2280 gnd 0.007204f
C4508 vdd.n2281 gnd 0.007204f
C4509 vdd.n2282 gnd 0.007204f
C4510 vdd.n2283 gnd 0.007204f
C4511 vdd.n2285 gnd 0.007204f
C4512 vdd.n2287 gnd 0.007204f
C4513 vdd.n2288 gnd 0.007204f
C4514 vdd.n2289 gnd 0.017093f
C4515 vdd.n2290 gnd 0.015959f
C4516 vdd.n2291 gnd 0.015959f
C4517 vdd.n2292 gnd 1.06096f
C4518 vdd.n2293 gnd 0.015959f
C4519 vdd.n2294 gnd 0.015959f
C4520 vdd.n2295 gnd 0.007204f
C4521 vdd.n2296 gnd 0.007204f
C4522 vdd.n2297 gnd 0.007204f
C4523 vdd.n2298 gnd 0.460108f
C4524 vdd.n2299 gnd 0.007204f
C4525 vdd.n2300 gnd 0.007204f
C4526 vdd.n2301 gnd 0.007204f
C4527 vdd.n2302 gnd 0.007204f
C4528 vdd.n2303 gnd 0.007204f
C4529 vdd.n2304 gnd 0.736173f
C4530 vdd.n2305 gnd 0.007204f
C4531 vdd.n2306 gnd 0.007204f
C4532 vdd.n2307 gnd 0.007204f
C4533 vdd.n2308 gnd 0.007204f
C4534 vdd.n2309 gnd 0.007204f
C4535 vdd.n2310 gnd 0.736173f
C4536 vdd.n2311 gnd 0.007204f
C4537 vdd.n2312 gnd 0.007204f
C4538 vdd.n2313 gnd 0.006356f
C4539 vdd.n2314 gnd 0.020868f
C4540 vdd.n2315 gnd 0.004449f
C4541 vdd.n2316 gnd 0.007204f
C4542 vdd.n2317 gnd 0.405978f
C4543 vdd.n2318 gnd 0.007204f
C4544 vdd.n2319 gnd 0.007204f
C4545 vdd.n2320 gnd 0.007204f
C4546 vdd.n2321 gnd 0.007204f
C4547 vdd.n2322 gnd 0.007204f
C4548 vdd.n2323 gnd 0.492586f
C4549 vdd.n2324 gnd 0.007204f
C4550 vdd.n2325 gnd 0.007204f
C4551 vdd.n2326 gnd 0.007204f
C4552 vdd.n2327 gnd 0.007204f
C4553 vdd.n2328 gnd 0.007204f
C4554 vdd.n2329 gnd 0.654978f
C4555 vdd.n2330 gnd 0.007204f
C4556 vdd.n2331 gnd 0.007204f
C4557 vdd.n2332 gnd 0.007204f
C4558 vdd.n2333 gnd 0.007204f
C4559 vdd.n2334 gnd 0.007204f
C4560 vdd.n2335 gnd 0.584608f
C4561 vdd.n2336 gnd 0.007204f
C4562 vdd.n2337 gnd 0.007204f
C4563 vdd.n2338 gnd 0.007204f
C4564 vdd.n2339 gnd 0.007204f
C4565 vdd.n2340 gnd 0.007204f
C4566 vdd.n2341 gnd 0.422217f
C4567 vdd.n2342 gnd 0.007204f
C4568 vdd.n2343 gnd 0.007204f
C4569 vdd.n2344 gnd 0.007204f
C4570 vdd.n2345 gnd 0.007204f
C4571 vdd.n2346 gnd 0.007204f
C4572 vdd.n2347 gnd 0.232761f
C4573 vdd.n2348 gnd 0.007204f
C4574 vdd.n2349 gnd 0.007204f
C4575 vdd.n2350 gnd 0.007204f
C4576 vdd.n2351 gnd 0.007204f
C4577 vdd.n2352 gnd 0.007204f
C4578 vdd.n2353 gnd 0.405978f
C4579 vdd.n2354 gnd 0.007204f
C4580 vdd.n2355 gnd 0.007204f
C4581 vdd.n2356 gnd 0.007204f
C4582 vdd.n2357 gnd 0.007204f
C4583 vdd.n2358 gnd 0.007204f
C4584 vdd.n2359 gnd 0.736173f
C4585 vdd.n2360 gnd 0.007204f
C4586 vdd.n2361 gnd 0.007204f
C4587 vdd.n2362 gnd 0.007204f
C4588 vdd.n2363 gnd 0.007204f
C4589 vdd.n2364 gnd 0.007204f
C4590 vdd.n2365 gnd 0.007204f
C4591 vdd.n2366 gnd 0.007204f
C4592 vdd.n2367 gnd 0.573782f
C4593 vdd.n2368 gnd 0.007204f
C4594 vdd.n2369 gnd 0.007204f
C4595 vdd.n2370 gnd 0.007204f
C4596 vdd.n2371 gnd 0.007204f
C4597 vdd.n2372 gnd 0.007204f
C4598 vdd.n2373 gnd 0.007204f
C4599 vdd.n2374 gnd 0.460108f
C4600 vdd.n2375 gnd 0.007204f
C4601 vdd.n2376 gnd 0.007204f
C4602 vdd.n2377 gnd 0.007204f
C4603 vdd.n2378 gnd 0.016836f
C4604 vdd.n2379 gnd 0.016216f
C4605 vdd.n2380 gnd 0.007204f
C4606 vdd.n2381 gnd 0.007204f
C4607 vdd.n2382 gnd 0.005562f
C4608 vdd.n2383 gnd 0.007204f
C4609 vdd.n2384 gnd 0.007204f
C4610 vdd.n2385 gnd 0.005244f
C4611 vdd.n2386 gnd 0.007204f
C4612 vdd.n2387 gnd 0.007204f
C4613 vdd.n2388 gnd 0.007204f
C4614 vdd.n2389 gnd 0.007204f
C4615 vdd.n2390 gnd 0.007204f
C4616 vdd.n2391 gnd 0.007204f
C4617 vdd.n2392 gnd 0.007204f
C4618 vdd.n2393 gnd 0.007204f
C4619 vdd.n2394 gnd 0.007204f
C4620 vdd.n2395 gnd 0.007204f
C4621 vdd.n2396 gnd 0.007204f
C4622 vdd.n2397 gnd 0.007204f
C4623 vdd.n2398 gnd 0.007204f
C4624 vdd.n2399 gnd 0.007204f
C4625 vdd.n2400 gnd 0.007204f
C4626 vdd.n2401 gnd 0.007204f
C4627 vdd.n2402 gnd 0.007204f
C4628 vdd.n2403 gnd 0.007204f
C4629 vdd.n2404 gnd 0.007204f
C4630 vdd.n2405 gnd 0.007204f
C4631 vdd.n2406 gnd 0.007204f
C4632 vdd.n2407 gnd 0.007204f
C4633 vdd.n2408 gnd 0.007204f
C4634 vdd.n2409 gnd 0.007204f
C4635 vdd.n2410 gnd 0.007204f
C4636 vdd.n2411 gnd 0.007204f
C4637 vdd.n2412 gnd 0.007204f
C4638 vdd.n2413 gnd 0.007204f
C4639 vdd.n2414 gnd 0.007204f
C4640 vdd.n2415 gnd 0.007204f
C4641 vdd.n2416 gnd 0.007204f
C4642 vdd.n2417 gnd 0.007204f
C4643 vdd.n2418 gnd 0.007204f
C4644 vdd.n2419 gnd 0.007204f
C4645 vdd.n2420 gnd 0.007204f
C4646 vdd.n2421 gnd 0.007204f
C4647 vdd.n2422 gnd 0.007204f
C4648 vdd.n2423 gnd 0.007204f
C4649 vdd.n2424 gnd 0.007204f
C4650 vdd.n2425 gnd 0.007204f
C4651 vdd.n2426 gnd 0.007204f
C4652 vdd.n2427 gnd 0.007204f
C4653 vdd.n2428 gnd 0.007204f
C4654 vdd.n2429 gnd 0.007204f
C4655 vdd.n2430 gnd 0.007204f
C4656 vdd.n2431 gnd 0.007204f
C4657 vdd.n2432 gnd 0.007204f
C4658 vdd.n2433 gnd 0.007204f
C4659 vdd.n2434 gnd 0.007204f
C4660 vdd.n2435 gnd 0.007204f
C4661 vdd.n2436 gnd 0.007204f
C4662 vdd.n2437 gnd 0.007204f
C4663 vdd.n2438 gnd 0.007204f
C4664 vdd.n2439 gnd 0.007204f
C4665 vdd.n2440 gnd 0.007204f
C4666 vdd.n2441 gnd 0.007204f
C4667 vdd.n2442 gnd 0.007204f
C4668 vdd.n2443 gnd 0.007204f
C4669 vdd.n2444 gnd 0.007204f
C4670 vdd.n2445 gnd 0.007204f
C4671 vdd.n2446 gnd 0.017093f
C4672 vdd.n2447 gnd 0.015959f
C4673 vdd.n2448 gnd 0.015959f
C4674 vdd.n2449 gnd 0.898564f
C4675 vdd.n2450 gnd 0.015959f
C4676 vdd.n2451 gnd 0.017093f
C4677 vdd.n2452 gnd 0.016216f
C4678 vdd.n2453 gnd 0.007204f
C4679 vdd.n2454 gnd 0.007204f
C4680 vdd.n2455 gnd 0.007204f
C4681 vdd.n2456 gnd 0.005562f
C4682 vdd.n2457 gnd 0.010295f
C4683 vdd.n2458 gnd 0.005244f
C4684 vdd.n2459 gnd 0.007204f
C4685 vdd.n2460 gnd 0.007204f
C4686 vdd.n2461 gnd 0.007204f
C4687 vdd.n2462 gnd 0.007204f
C4688 vdd.n2463 gnd 0.007204f
C4689 vdd.n2464 gnd 0.007204f
C4690 vdd.n2465 gnd 0.007204f
C4691 vdd.n2466 gnd 0.007204f
C4692 vdd.n2467 gnd 0.007204f
C4693 vdd.n2468 gnd 0.007204f
C4694 vdd.n2469 gnd 0.007204f
C4695 vdd.n2470 gnd 0.007204f
C4696 vdd.n2471 gnd 0.007204f
C4697 vdd.n2472 gnd 0.007204f
C4698 vdd.n2473 gnd 0.007204f
C4699 vdd.n2474 gnd 0.007204f
C4700 vdd.n2475 gnd 0.007204f
C4701 vdd.n2476 gnd 0.007204f
C4702 vdd.n2477 gnd 0.007204f
C4703 vdd.n2478 gnd 0.007204f
C4704 vdd.n2479 gnd 0.007204f
C4705 vdd.n2480 gnd 0.007204f
C4706 vdd.n2481 gnd 0.007204f
C4707 vdd.n2482 gnd 0.007204f
C4708 vdd.n2483 gnd 0.007204f
C4709 vdd.n2484 gnd 0.007204f
C4710 vdd.n2485 gnd 0.007204f
C4711 vdd.n2486 gnd 0.007204f
C4712 vdd.n2487 gnd 0.007204f
C4713 vdd.n2488 gnd 0.007204f
C4714 vdd.n2489 gnd 0.007204f
C4715 vdd.n2490 gnd 0.007204f
C4716 vdd.n2491 gnd 0.007204f
C4717 vdd.n2492 gnd 0.007204f
C4718 vdd.n2493 gnd 0.007204f
C4719 vdd.n2494 gnd 0.007204f
C4720 vdd.n2495 gnd 0.007204f
C4721 vdd.n2496 gnd 0.007204f
C4722 vdd.n2497 gnd 0.007204f
C4723 vdd.n2498 gnd 0.007204f
C4724 vdd.n2499 gnd 0.007204f
C4725 vdd.n2500 gnd 0.007204f
C4726 vdd.n2501 gnd 0.007204f
C4727 vdd.n2502 gnd 0.007204f
C4728 vdd.n2503 gnd 0.007204f
C4729 vdd.n2504 gnd 0.007204f
C4730 vdd.n2505 gnd 0.007204f
C4731 vdd.n2506 gnd 0.007204f
C4732 vdd.n2507 gnd 0.007204f
C4733 vdd.n2508 gnd 0.007204f
C4734 vdd.n2509 gnd 0.007204f
C4735 vdd.n2510 gnd 0.007204f
C4736 vdd.n2511 gnd 0.007204f
C4737 vdd.n2512 gnd 0.007204f
C4738 vdd.n2513 gnd 0.007204f
C4739 vdd.n2514 gnd 0.007204f
C4740 vdd.n2515 gnd 0.007204f
C4741 vdd.n2516 gnd 0.007204f
C4742 vdd.n2517 gnd 0.007204f
C4743 vdd.n2518 gnd 0.007204f
C4744 vdd.n2519 gnd 0.017093f
C4745 vdd.n2520 gnd 0.017093f
C4746 vdd.n2521 gnd 0.898564f
C4747 vdd.t13 gnd 3.19369f
C4748 vdd.t262 gnd 3.19369f
C4749 vdd.n2554 gnd 0.017093f
C4750 vdd.n2555 gnd 0.007204f
C4751 vdd.t72 gnd 0.291096f
C4752 vdd.t73 gnd 0.297973f
C4753 vdd.t70 gnd 0.190039f
C4754 vdd.n2556 gnd 0.102706f
C4755 vdd.n2557 gnd 0.058258f
C4756 vdd.n2558 gnd 0.007204f
C4757 vdd.t85 gnd 0.291096f
C4758 vdd.t86 gnd 0.297973f
C4759 vdd.t84 gnd 0.190039f
C4760 vdd.n2559 gnd 0.102706f
C4761 vdd.n2560 gnd 0.058258f
C4762 vdd.n2561 gnd 0.010295f
C4763 vdd.n2562 gnd 0.007204f
C4764 vdd.n2563 gnd 0.007204f
C4765 vdd.n2564 gnd 0.007204f
C4766 vdd.n2565 gnd 0.007204f
C4767 vdd.n2566 gnd 0.007204f
C4768 vdd.n2567 gnd 0.007204f
C4769 vdd.n2568 gnd 0.007204f
C4770 vdd.n2569 gnd 0.007204f
C4771 vdd.n2570 gnd 0.007204f
C4772 vdd.n2571 gnd 0.007204f
C4773 vdd.n2572 gnd 0.007204f
C4774 vdd.n2573 gnd 0.007204f
C4775 vdd.n2574 gnd 0.007204f
C4776 vdd.n2575 gnd 0.007204f
C4777 vdd.n2576 gnd 0.007204f
C4778 vdd.n2577 gnd 0.007204f
C4779 vdd.n2578 gnd 0.007204f
C4780 vdd.n2579 gnd 0.007204f
C4781 vdd.n2580 gnd 0.007204f
C4782 vdd.n2581 gnd 0.007204f
C4783 vdd.n2582 gnd 0.007204f
C4784 vdd.n2583 gnd 0.007204f
C4785 vdd.n2584 gnd 0.007204f
C4786 vdd.n2585 gnd 0.007204f
C4787 vdd.n2586 gnd 0.007204f
C4788 vdd.n2587 gnd 0.007204f
C4789 vdd.n2588 gnd 0.007204f
C4790 vdd.n2589 gnd 0.007204f
C4791 vdd.n2590 gnd 0.007204f
C4792 vdd.n2591 gnd 0.007204f
C4793 vdd.n2592 gnd 0.007204f
C4794 vdd.n2593 gnd 0.007204f
C4795 vdd.n2594 gnd 0.007204f
C4796 vdd.n2595 gnd 0.007204f
C4797 vdd.n2596 gnd 0.007204f
C4798 vdd.n2597 gnd 0.007204f
C4799 vdd.n2598 gnd 0.007204f
C4800 vdd.n2599 gnd 0.007204f
C4801 vdd.n2600 gnd 0.007204f
C4802 vdd.n2601 gnd 0.007204f
C4803 vdd.n2602 gnd 0.007204f
C4804 vdd.n2603 gnd 0.007204f
C4805 vdd.n2604 gnd 0.007204f
C4806 vdd.n2605 gnd 0.007204f
C4807 vdd.n2606 gnd 0.007204f
C4808 vdd.n2607 gnd 0.007204f
C4809 vdd.n2608 gnd 0.007204f
C4810 vdd.n2609 gnd 0.007204f
C4811 vdd.n2610 gnd 0.007204f
C4812 vdd.n2611 gnd 0.007204f
C4813 vdd.n2612 gnd 0.007204f
C4814 vdd.n2613 gnd 0.007204f
C4815 vdd.n2614 gnd 0.007204f
C4816 vdd.n2615 gnd 0.007204f
C4817 vdd.n2616 gnd 0.007204f
C4818 vdd.n2617 gnd 0.007204f
C4819 vdd.n2618 gnd 0.005244f
C4820 vdd.n2619 gnd 0.007204f
C4821 vdd.n2620 gnd 0.007204f
C4822 vdd.n2621 gnd 0.005562f
C4823 vdd.n2622 gnd 0.007204f
C4824 vdd.n2623 gnd 0.007204f
C4825 vdd.n2624 gnd 0.017093f
C4826 vdd.n2625 gnd 0.015959f
C4827 vdd.n2626 gnd 0.007204f
C4828 vdd.n2627 gnd 0.007204f
C4829 vdd.n2628 gnd 0.007204f
C4830 vdd.n2629 gnd 0.007204f
C4831 vdd.n2630 gnd 0.007204f
C4832 vdd.n2631 gnd 0.007204f
C4833 vdd.n2632 gnd 0.007204f
C4834 vdd.n2633 gnd 0.007204f
C4835 vdd.n2634 gnd 0.007204f
C4836 vdd.n2635 gnd 0.007204f
C4837 vdd.n2636 gnd 0.007204f
C4838 vdd.n2637 gnd 0.007204f
C4839 vdd.n2638 gnd 0.007204f
C4840 vdd.n2639 gnd 0.007204f
C4841 vdd.n2640 gnd 0.007204f
C4842 vdd.n2641 gnd 0.007204f
C4843 vdd.n2642 gnd 0.007204f
C4844 vdd.n2643 gnd 0.007204f
C4845 vdd.n2644 gnd 0.007204f
C4846 vdd.n2645 gnd 0.007204f
C4847 vdd.n2646 gnd 0.007204f
C4848 vdd.n2647 gnd 0.007204f
C4849 vdd.n2648 gnd 0.007204f
C4850 vdd.n2649 gnd 0.007204f
C4851 vdd.n2650 gnd 0.007204f
C4852 vdd.n2651 gnd 0.007204f
C4853 vdd.n2652 gnd 0.007204f
C4854 vdd.n2653 gnd 0.007204f
C4855 vdd.n2654 gnd 0.007204f
C4856 vdd.n2655 gnd 0.007204f
C4857 vdd.n2656 gnd 0.007204f
C4858 vdd.n2657 gnd 0.007204f
C4859 vdd.n2658 gnd 0.007204f
C4860 vdd.n2659 gnd 0.007204f
C4861 vdd.n2660 gnd 0.007204f
C4862 vdd.n2661 gnd 0.007204f
C4863 vdd.n2662 gnd 0.007204f
C4864 vdd.n2663 gnd 0.007204f
C4865 vdd.n2664 gnd 0.007204f
C4866 vdd.n2665 gnd 0.007204f
C4867 vdd.n2666 gnd 0.007204f
C4868 vdd.n2667 gnd 0.007204f
C4869 vdd.n2668 gnd 0.007204f
C4870 vdd.n2669 gnd 0.007204f
C4871 vdd.n2670 gnd 0.007204f
C4872 vdd.n2671 gnd 0.007204f
C4873 vdd.n2672 gnd 0.007204f
C4874 vdd.n2673 gnd 0.007204f
C4875 vdd.n2674 gnd 0.007204f
C4876 vdd.n2675 gnd 0.007204f
C4877 vdd.n2676 gnd 0.007204f
C4878 vdd.n2677 gnd 0.232761f
C4879 vdd.n2678 gnd 0.007204f
C4880 vdd.n2679 gnd 0.007204f
C4881 vdd.n2680 gnd 0.007204f
C4882 vdd.n2681 gnd 0.007204f
C4883 vdd.n2682 gnd 0.007204f
C4884 vdd.n2683 gnd 0.007204f
C4885 vdd.n2684 gnd 0.007204f
C4886 vdd.n2685 gnd 0.007204f
C4887 vdd.n2686 gnd 0.007204f
C4888 vdd.n2687 gnd 0.007204f
C4889 vdd.n2688 gnd 0.007204f
C4890 vdd.n2689 gnd 0.007204f
C4891 vdd.n2690 gnd 0.007204f
C4892 vdd.n2691 gnd 0.007204f
C4893 vdd.n2692 gnd 0.007204f
C4894 vdd.n2693 gnd 0.007204f
C4895 vdd.n2694 gnd 0.007204f
C4896 vdd.n2695 gnd 0.007204f
C4897 vdd.n2696 gnd 0.007204f
C4898 vdd.n2697 gnd 0.007204f
C4899 vdd.n2698 gnd 0.438456f
C4900 vdd.n2699 gnd 0.007204f
C4901 vdd.n2700 gnd 0.007204f
C4902 vdd.n2701 gnd 0.007204f
C4903 vdd.n2702 gnd 0.007204f
C4904 vdd.n2703 gnd 0.007204f
C4905 vdd.n2704 gnd 0.015959f
C4906 vdd.n2705 gnd 0.017093f
C4907 vdd.n2706 gnd 0.017093f
C4908 vdd.n2707 gnd 0.007204f
C4909 vdd.n2708 gnd 0.007204f
C4910 vdd.n2709 gnd 0.007204f
C4911 vdd.n2710 gnd 0.005562f
C4912 vdd.n2711 gnd 0.010295f
C4913 vdd.n2712 gnd 0.005244f
C4914 vdd.n2713 gnd 0.007204f
C4915 vdd.n2714 gnd 0.007204f
C4916 vdd.n2715 gnd 0.007204f
C4917 vdd.n2716 gnd 0.007204f
C4918 vdd.n2717 gnd 0.007204f
C4919 vdd.n2718 gnd 0.007204f
C4920 vdd.n2719 gnd 0.007204f
C4921 vdd.n2720 gnd 0.007204f
C4922 vdd.n2721 gnd 0.007204f
C4923 vdd.n2722 gnd 0.007204f
C4924 vdd.n2723 gnd 0.007204f
C4925 vdd.n2724 gnd 0.007204f
C4926 vdd.n2725 gnd 0.007204f
C4927 vdd.n2726 gnd 0.007204f
C4928 vdd.n2727 gnd 0.007204f
C4929 vdd.n2728 gnd 0.007204f
C4930 vdd.n2729 gnd 0.007204f
C4931 vdd.n2730 gnd 0.007204f
C4932 vdd.n2731 gnd 0.007204f
C4933 vdd.n2732 gnd 0.007204f
C4934 vdd.n2733 gnd 0.007204f
C4935 vdd.n2734 gnd 0.007204f
C4936 vdd.n2735 gnd 0.007204f
C4937 vdd.n2736 gnd 0.007204f
C4938 vdd.n2737 gnd 0.007204f
C4939 vdd.n2738 gnd 0.007204f
C4940 vdd.n2739 gnd 0.007204f
C4941 vdd.n2740 gnd 0.007204f
C4942 vdd.n2741 gnd 0.007204f
C4943 vdd.n2742 gnd 0.007204f
C4944 vdd.n2743 gnd 0.007204f
C4945 vdd.n2744 gnd 0.007204f
C4946 vdd.n2745 gnd 0.007204f
C4947 vdd.n2746 gnd 0.007204f
C4948 vdd.n2747 gnd 0.007204f
C4949 vdd.n2748 gnd 0.007204f
C4950 vdd.n2749 gnd 0.007204f
C4951 vdd.n2750 gnd 0.007204f
C4952 vdd.n2751 gnd 0.007204f
C4953 vdd.n2752 gnd 0.007204f
C4954 vdd.n2753 gnd 0.007204f
C4955 vdd.n2754 gnd 0.007204f
C4956 vdd.n2755 gnd 0.007204f
C4957 vdd.n2756 gnd 0.007204f
C4958 vdd.n2757 gnd 0.007204f
C4959 vdd.n2758 gnd 0.007204f
C4960 vdd.n2759 gnd 0.007204f
C4961 vdd.n2760 gnd 0.007204f
C4962 vdd.n2761 gnd 0.007204f
C4963 vdd.n2762 gnd 0.007204f
C4964 vdd.n2763 gnd 0.007204f
C4965 vdd.n2764 gnd 0.007204f
C4966 vdd.n2765 gnd 0.007204f
C4967 vdd.n2766 gnd 0.007204f
C4968 vdd.n2767 gnd 0.007204f
C4969 vdd.n2768 gnd 0.007204f
C4970 vdd.n2769 gnd 0.007204f
C4971 vdd.n2770 gnd 0.007204f
C4972 vdd.n2771 gnd 0.007204f
C4973 vdd.n2772 gnd 0.007204f
C4974 vdd.n2774 gnd 0.898564f
C4975 vdd.n2776 gnd 0.007204f
C4976 vdd.n2777 gnd 0.007204f
C4977 vdd.n2778 gnd 0.017093f
C4978 vdd.n2779 gnd 0.015959f
C4979 vdd.n2780 gnd 0.015959f
C4980 vdd.n2781 gnd 0.898564f
C4981 vdd.n2782 gnd 0.015959f
C4982 vdd.n2783 gnd 0.015959f
C4983 vdd.n2784 gnd 0.007204f
C4984 vdd.n2785 gnd 0.007204f
C4985 vdd.n2786 gnd 0.007204f
C4986 vdd.n2787 gnd 0.460108f
C4987 vdd.n2788 gnd 0.007204f
C4988 vdd.n2789 gnd 0.007204f
C4989 vdd.n2790 gnd 0.007204f
C4990 vdd.n2791 gnd 0.007204f
C4991 vdd.n2792 gnd 0.007204f
C4992 vdd.n2793 gnd 0.573782f
C4993 vdd.n2794 gnd 0.007204f
C4994 vdd.n2795 gnd 0.007204f
C4995 vdd.n2796 gnd 0.007204f
C4996 vdd.n2797 gnd 0.007204f
C4997 vdd.n2798 gnd 0.007204f
C4998 vdd.n2799 gnd 0.736173f
C4999 vdd.n2800 gnd 0.007204f
C5000 vdd.n2801 gnd 0.007204f
C5001 vdd.n2802 gnd 0.007204f
C5002 vdd.n2803 gnd 0.007204f
C5003 vdd.n2804 gnd 0.007204f
C5004 vdd.n2805 gnd 0.405978f
C5005 vdd.n2806 gnd 0.007204f
C5006 vdd.n2807 gnd 0.007204f
C5007 vdd.n2808 gnd 0.007204f
C5008 vdd.n2809 gnd 0.007204f
C5009 vdd.n2810 gnd 0.007204f
C5010 vdd.n2811 gnd 0.232761f
C5011 vdd.n2812 gnd 0.007204f
C5012 vdd.n2813 gnd 0.007204f
C5013 vdd.n2814 gnd 0.007204f
C5014 vdd.n2815 gnd 0.007204f
C5015 vdd.n2816 gnd 0.007204f
C5016 vdd.n2817 gnd 0.422217f
C5017 vdd.n2818 gnd 0.007204f
C5018 vdd.n2819 gnd 0.007204f
C5019 vdd.n2820 gnd 0.007204f
C5020 vdd.n2821 gnd 0.007204f
C5021 vdd.n2822 gnd 0.007204f
C5022 vdd.n2823 gnd 0.584608f
C5023 vdd.n2824 gnd 0.007204f
C5024 vdd.n2825 gnd 0.007204f
C5025 vdd.n2826 gnd 0.007204f
C5026 vdd.n2827 gnd 0.007204f
C5027 vdd.n2828 gnd 0.007204f
C5028 vdd.n2829 gnd 0.654978f
C5029 vdd.n2830 gnd 0.007204f
C5030 vdd.n2831 gnd 0.007204f
C5031 vdd.n2832 gnd 0.007204f
C5032 vdd.n2833 gnd 0.007204f
C5033 vdd.n2834 gnd 0.007204f
C5034 vdd.n2835 gnd 0.492586f
C5035 vdd.n2836 gnd 0.007204f
C5036 vdd.n2837 gnd 0.007204f
C5037 vdd.n2838 gnd 0.007204f
C5038 vdd.t51 gnd 0.297973f
C5039 vdd.t49 gnd 0.190039f
C5040 vdd.t52 gnd 0.297973f
C5041 vdd.n2839 gnd 0.167473f
C5042 vdd.n2840 gnd 0.020868f
C5043 vdd.n2841 gnd 0.004449f
C5044 vdd.n2842 gnd 0.007204f
C5045 vdd.n2843 gnd 0.405978f
C5046 vdd.n2844 gnd 0.007204f
C5047 vdd.n2845 gnd 0.007204f
C5048 vdd.n2846 gnd 0.007204f
C5049 vdd.n2847 gnd 0.007204f
C5050 vdd.n2848 gnd 0.007204f
C5051 vdd.n2849 gnd 0.736173f
C5052 vdd.n2850 gnd 0.007204f
C5053 vdd.n2851 gnd 0.007204f
C5054 vdd.n2852 gnd 0.007204f
C5055 vdd.n2853 gnd 0.007204f
C5056 vdd.n2854 gnd 0.007204f
C5057 vdd.n2855 gnd 0.007204f
C5058 vdd.n2857 gnd 0.007204f
C5059 vdd.n2858 gnd 0.007204f
C5060 vdd.n2860 gnd 0.007204f
C5061 vdd.n2861 gnd 0.007204f
C5062 vdd.n2864 gnd 0.007204f
C5063 vdd.n2865 gnd 0.007204f
C5064 vdd.n2866 gnd 0.007204f
C5065 vdd.n2867 gnd 0.007204f
C5066 vdd.n2869 gnd 0.007204f
C5067 vdd.n2870 gnd 0.007204f
C5068 vdd.n2871 gnd 0.007204f
C5069 vdd.n2872 gnd 0.007204f
C5070 vdd.n2873 gnd 0.007204f
C5071 vdd.n2874 gnd 0.007204f
C5072 vdd.n2876 gnd 0.007204f
C5073 vdd.n2877 gnd 0.007204f
C5074 vdd.n2878 gnd 0.007204f
C5075 vdd.n2879 gnd 0.007204f
C5076 vdd.n2880 gnd 0.007204f
C5077 vdd.n2881 gnd 0.007204f
C5078 vdd.n2883 gnd 0.007204f
C5079 vdd.n2884 gnd 0.007204f
C5080 vdd.n2885 gnd 0.007204f
C5081 vdd.n2886 gnd 0.007204f
C5082 vdd.n2887 gnd 0.007204f
C5083 vdd.n2888 gnd 0.007204f
C5084 vdd.n2890 gnd 0.007204f
C5085 vdd.n2891 gnd 0.017093f
C5086 vdd.n2892 gnd 0.017093f
C5087 vdd.n2893 gnd 0.015959f
C5088 vdd.n2894 gnd 0.007204f
C5089 vdd.n2895 gnd 0.007204f
C5090 vdd.n2896 gnd 0.007204f
C5091 vdd.n2897 gnd 0.007204f
C5092 vdd.n2898 gnd 0.007204f
C5093 vdd.n2899 gnd 0.007204f
C5094 vdd.n2900 gnd 0.736173f
C5095 vdd.n2901 gnd 0.007204f
C5096 vdd.n2902 gnd 0.007204f
C5097 vdd.n2903 gnd 0.007204f
C5098 vdd.n2904 gnd 0.007204f
C5099 vdd.n2905 gnd 0.007204f
C5100 vdd.n2906 gnd 0.460108f
C5101 vdd.n2907 gnd 0.007204f
C5102 vdd.n2908 gnd 0.007204f
C5103 vdd.n2909 gnd 0.007204f
C5104 vdd.n2910 gnd 0.016836f
C5105 vdd.n2912 gnd 0.017093f
C5106 vdd.n2913 gnd 0.016216f
C5107 vdd.n2914 gnd 0.007204f
C5108 vdd.n2915 gnd 0.005562f
C5109 vdd.n2916 gnd 0.007204f
C5110 vdd.n2918 gnd 0.007204f
C5111 vdd.n2919 gnd 0.007204f
C5112 vdd.n2920 gnd 0.007204f
C5113 vdd.n2921 gnd 0.007204f
C5114 vdd.n2922 gnd 0.007204f
C5115 vdd.n2923 gnd 0.007204f
C5116 vdd.n2925 gnd 0.007204f
C5117 vdd.n2926 gnd 0.007204f
C5118 vdd.n2927 gnd 0.007204f
C5119 vdd.n2928 gnd 0.007204f
C5120 vdd.n2929 gnd 0.007204f
C5121 vdd.n2930 gnd 0.007204f
C5122 vdd.n2932 gnd 0.007204f
C5123 vdd.n2933 gnd 0.007204f
C5124 vdd.n2934 gnd 0.007204f
C5125 vdd.n2935 gnd 0.007204f
C5126 vdd.n2936 gnd 0.007204f
C5127 vdd.n2937 gnd 0.007204f
C5128 vdd.n2939 gnd 0.007204f
C5129 vdd.n2940 gnd 0.007204f
C5130 vdd.n2941 gnd 0.007204f
C5131 vdd.n2942 gnd 0.641137f
C5132 vdd.n2943 gnd 0.017311f
C5133 vdd.n2944 gnd 0.007204f
C5134 vdd.n2945 gnd 0.007204f
C5135 vdd.n2947 gnd 0.007204f
C5136 vdd.n2948 gnd 0.007204f
C5137 vdd.n2949 gnd 0.007204f
C5138 vdd.n2950 gnd 0.007204f
C5139 vdd.n2951 gnd 0.007204f
C5140 vdd.n2952 gnd 0.007204f
C5141 vdd.n2954 gnd 0.007204f
C5142 vdd.n2955 gnd 0.007204f
C5143 vdd.n2956 gnd 0.007204f
C5144 vdd.n2957 gnd 0.007204f
C5145 vdd.n2958 gnd 0.007204f
C5146 vdd.n2959 gnd 0.007204f
C5147 vdd.n2961 gnd 0.007204f
C5148 vdd.n2962 gnd 0.007204f
C5149 vdd.n2963 gnd 0.007204f
C5150 vdd.n2964 gnd 0.007204f
C5151 vdd.n2965 gnd 0.007204f
C5152 vdd.n2966 gnd 0.007204f
C5153 vdd.n2968 gnd 0.007204f
C5154 vdd.n2969 gnd 0.007204f
C5155 vdd.n2971 gnd 0.007204f
C5156 vdd.n2972 gnd 0.007204f
C5157 vdd.n2973 gnd 0.017093f
C5158 vdd.n2974 gnd 0.015959f
C5159 vdd.n2975 gnd 0.015959f
C5160 vdd.n2976 gnd 1.06096f
C5161 vdd.n2977 gnd 0.015959f
C5162 vdd.n2978 gnd 0.017093f
C5163 vdd.n2979 gnd 0.016216f
C5164 vdd.n2980 gnd 0.007204f
C5165 vdd.n2981 gnd 0.005562f
C5166 vdd.n2982 gnd 0.007204f
C5167 vdd.n2984 gnd 0.007204f
C5168 vdd.n2985 gnd 0.007204f
C5169 vdd.n2986 gnd 0.007204f
C5170 vdd.n2987 gnd 0.007204f
C5171 vdd.n2988 gnd 0.007204f
C5172 vdd.n2989 gnd 0.007204f
C5173 vdd.n2991 gnd 0.007204f
C5174 vdd.n2992 gnd 0.007204f
C5175 vdd.n2993 gnd 0.007204f
C5176 vdd.n2994 gnd 0.007204f
C5177 vdd.n2995 gnd 0.007204f
C5178 vdd.n2996 gnd 0.007204f
C5179 vdd.n2998 gnd 0.007204f
C5180 vdd.n2999 gnd 0.007204f
C5181 vdd.n3000 gnd 0.007204f
C5182 vdd.n3001 gnd 0.007204f
C5183 vdd.n3002 gnd 0.007204f
C5184 vdd.n3003 gnd 0.007204f
C5185 vdd.n3005 gnd 0.007204f
C5186 vdd.n3006 gnd 0.007204f
C5187 vdd.n3008 gnd 0.007204f
C5188 vdd.n3009 gnd 0.017311f
C5189 vdd.n3010 gnd 0.641137f
C5190 vdd.n3011 gnd 0.00911f
C5191 vdd.n3012 gnd 0.00405f
C5192 vdd.t94 gnd 0.130328f
C5193 vdd.t95 gnd 0.139285f
C5194 vdd.t93 gnd 0.170207f
C5195 vdd.n3013 gnd 0.218181f
C5196 vdd.n3014 gnd 0.183312f
C5197 vdd.n3015 gnd 0.013131f
C5198 vdd.n3016 gnd 0.010593f
C5199 vdd.n3017 gnd 0.004476f
C5200 vdd.n3018 gnd 0.008527f
C5201 vdd.n3019 gnd 0.010593f
C5202 vdd.n3020 gnd 0.010593f
C5203 vdd.n3021 gnd 0.008527f
C5204 vdd.n3022 gnd 0.008527f
C5205 vdd.n3023 gnd 0.010593f
C5206 vdd.n3025 gnd 0.010593f
C5207 vdd.n3026 gnd 0.008527f
C5208 vdd.n3027 gnd 0.008527f
C5209 vdd.n3028 gnd 0.008527f
C5210 vdd.n3029 gnd 0.010593f
C5211 vdd.n3031 gnd 0.010593f
C5212 vdd.n3033 gnd 0.010593f
C5213 vdd.n3034 gnd 0.008527f
C5214 vdd.n3035 gnd 0.008527f
C5215 vdd.n3036 gnd 0.008527f
C5216 vdd.n3037 gnd 0.010593f
C5217 vdd.n3039 gnd 0.010593f
C5218 vdd.n3041 gnd 0.010593f
C5219 vdd.n3042 gnd 0.008527f
C5220 vdd.n3043 gnd 0.008527f
C5221 vdd.n3044 gnd 0.008527f
C5222 vdd.n3045 gnd 0.010593f
C5223 vdd.n3047 gnd 0.010593f
C5224 vdd.n3048 gnd 0.010593f
C5225 vdd.n3049 gnd 0.008527f
C5226 vdd.n3050 gnd 0.008527f
C5227 vdd.n3051 gnd 0.010593f
C5228 vdd.n3052 gnd 0.010593f
C5229 vdd.n3054 gnd 0.010593f
C5230 vdd.n3055 gnd 0.008527f
C5231 vdd.n3056 gnd 0.010593f
C5232 vdd.n3057 gnd 0.010593f
C5233 vdd.n3058 gnd 0.010593f
C5234 vdd.n3059 gnd 0.017394f
C5235 vdd.n3060 gnd 0.005798f
C5236 vdd.n3061 gnd 0.010593f
C5237 vdd.n3063 gnd 0.010593f
C5238 vdd.n3065 gnd 0.010593f
C5239 vdd.n3066 gnd 0.008527f
C5240 vdd.n3067 gnd 0.008527f
C5241 vdd.n3068 gnd 0.008527f
C5242 vdd.n3069 gnd 0.010593f
C5243 vdd.n3071 gnd 0.010593f
C5244 vdd.n3073 gnd 0.010593f
C5245 vdd.n3074 gnd 0.008527f
C5246 vdd.n3075 gnd 0.008527f
C5247 vdd.n3076 gnd 0.008527f
C5248 vdd.n3077 gnd 0.010593f
C5249 vdd.n3079 gnd 0.010593f
C5250 vdd.n3081 gnd 0.010593f
C5251 vdd.n3082 gnd 0.008527f
C5252 vdd.n3083 gnd 0.008527f
C5253 vdd.n3084 gnd 0.008527f
C5254 vdd.n3085 gnd 0.010593f
C5255 vdd.n3087 gnd 0.010593f
C5256 vdd.n3089 gnd 0.010593f
C5257 vdd.n3090 gnd 0.008527f
C5258 vdd.n3091 gnd 0.008527f
C5259 vdd.n3092 gnd 0.008527f
C5260 vdd.n3093 gnd 0.010593f
C5261 vdd.n3095 gnd 0.010593f
C5262 vdd.n3097 gnd 0.010593f
C5263 vdd.n3098 gnd 0.008527f
C5264 vdd.n3099 gnd 0.008527f
C5265 vdd.n3100 gnd 0.00712f
C5266 vdd.n3101 gnd 0.010593f
C5267 vdd.n3103 gnd 0.010593f
C5268 vdd.n3105 gnd 0.010593f
C5269 vdd.n3106 gnd 0.00712f
C5270 vdd.n3107 gnd 0.008527f
C5271 vdd.n3108 gnd 0.008527f
C5272 vdd.n3109 gnd 0.010593f
C5273 vdd.n3111 gnd 0.010593f
C5274 vdd.n3113 gnd 0.010593f
C5275 vdd.n3114 gnd 0.008527f
C5276 vdd.n3115 gnd 0.008527f
C5277 vdd.n3116 gnd 0.008527f
C5278 vdd.n3117 gnd 0.010593f
C5279 vdd.n3119 gnd 0.010593f
C5280 vdd.n3121 gnd 0.010593f
C5281 vdd.n3122 gnd 0.008527f
C5282 vdd.n3123 gnd 0.008527f
C5283 vdd.n3124 gnd 0.008527f
C5284 vdd.n3125 gnd 0.010593f
C5285 vdd.n3127 gnd 0.010593f
C5286 vdd.n3128 gnd 0.010593f
C5287 vdd.n3129 gnd 0.008527f
C5288 vdd.n3130 gnd 0.008527f
C5289 vdd.n3131 gnd 0.010593f
C5290 vdd.n3132 gnd 0.010593f
C5291 vdd.n3133 gnd 0.008527f
C5292 vdd.n3134 gnd 0.008527f
C5293 vdd.n3135 gnd 0.010593f
C5294 vdd.n3136 gnd 0.010593f
C5295 vdd.n3138 gnd 0.010593f
C5296 vdd.n3139 gnd 0.008527f
C5297 vdd.n3140 gnd 0.007077f
C5298 vdd.n3141 gnd 0.024289f
C5299 vdd.n3142 gnd 0.024124f
C5300 vdd.n3143 gnd 0.007077f
C5301 vdd.n3144 gnd 0.024124f
C5302 vdd.n3145 gnd 1.42904f
C5303 vdd.n3146 gnd 0.024124f
C5304 vdd.n3147 gnd 0.007077f
C5305 vdd.n3148 gnd 0.024124f
C5306 vdd.n3149 gnd 0.010593f
C5307 vdd.n3150 gnd 0.010593f
C5308 vdd.n3151 gnd 0.008527f
C5309 vdd.n3152 gnd 0.010593f
C5310 vdd.n3153 gnd 1.02306f
C5311 vdd.n3154 gnd 0.010593f
C5312 vdd.n3155 gnd 0.008527f
C5313 vdd.n3156 gnd 0.010593f
C5314 vdd.n3157 gnd 0.010593f
C5315 vdd.n3158 gnd 0.010593f
C5316 vdd.n3159 gnd 0.008527f
C5317 vdd.n3160 gnd 0.010593f
C5318 vdd.n3161 gnd 1.05554f
C5319 vdd.n3162 gnd 0.010593f
C5320 vdd.n3163 gnd 0.008527f
C5321 vdd.n3164 gnd 0.010593f
C5322 vdd.n3165 gnd 0.010593f
C5323 vdd.n3166 gnd 0.010593f
C5324 vdd.n3167 gnd 0.008527f
C5325 vdd.n3168 gnd 0.010593f
C5326 vdd.t198 gnd 0.541304f
C5327 vdd.n3169 gnd 0.871499f
C5328 vdd.n3170 gnd 0.010593f
C5329 vdd.n3171 gnd 0.008527f
C5330 vdd.n3172 gnd 0.010593f
C5331 vdd.n3173 gnd 0.010593f
C5332 vdd.n3174 gnd 0.010593f
C5333 vdd.n3175 gnd 0.008527f
C5334 vdd.n3176 gnd 0.010593f
C5335 vdd.n3177 gnd 0.687456f
C5336 vdd.n3178 gnd 0.010593f
C5337 vdd.n3179 gnd 0.008527f
C5338 vdd.n3180 gnd 0.010593f
C5339 vdd.n3181 gnd 0.010593f
C5340 vdd.n3182 gnd 0.010593f
C5341 vdd.n3183 gnd 0.008527f
C5342 vdd.n3184 gnd 0.010593f
C5343 vdd.n3185 gnd 0.860673f
C5344 vdd.n3186 gnd 0.579195f
C5345 vdd.n3187 gnd 0.010593f
C5346 vdd.n3188 gnd 0.008527f
C5347 vdd.n3189 gnd 0.010593f
C5348 vdd.n3190 gnd 0.010593f
C5349 vdd.n3191 gnd 0.010593f
C5350 vdd.n3192 gnd 0.008527f
C5351 vdd.n3193 gnd 0.010593f
C5352 vdd.n3194 gnd 0.763238f
C5353 vdd.n3195 gnd 0.010593f
C5354 vdd.n3196 gnd 0.008527f
C5355 vdd.n3197 gnd 0.010593f
C5356 vdd.n3198 gnd 0.010593f
C5357 vdd.n3199 gnd 0.010593f
C5358 vdd.n3200 gnd 0.010593f
C5359 vdd.n3201 gnd 0.010593f
C5360 vdd.n3202 gnd 0.008527f
C5361 vdd.n3203 gnd 0.008527f
C5362 vdd.n3204 gnd 0.010593f
C5363 vdd.t128 gnd 0.541304f
C5364 vdd.n3205 gnd 0.898564f
C5365 vdd.n3206 gnd 0.010593f
C5366 vdd.n3207 gnd 0.008527f
C5367 vdd.n3208 gnd 0.010593f
C5368 vdd.n3209 gnd 0.010593f
C5369 vdd.n3210 gnd 0.010593f
C5370 vdd.n3211 gnd 0.008527f
C5371 vdd.n3212 gnd 0.010593f
C5372 vdd.n3213 gnd 0.849847f
C5373 vdd.n3214 gnd 0.010593f
C5374 vdd.n3215 gnd 0.010593f
C5375 vdd.n3216 gnd 0.008527f
C5376 vdd.n3217 gnd 0.008527f
C5377 vdd.n3218 gnd 0.008527f
C5378 vdd.n3219 gnd 0.010593f
C5379 vdd.n3220 gnd 0.010593f
C5380 vdd.n3221 gnd 0.010593f
C5381 vdd.n3222 gnd 0.010593f
C5382 vdd.n3223 gnd 0.008527f
C5383 vdd.n3224 gnd 0.008527f
C5384 vdd.n3225 gnd 0.008527f
C5385 vdd.n3226 gnd 0.010593f
C5386 vdd.n3227 gnd 0.010593f
C5387 vdd.n3228 gnd 0.010593f
C5388 vdd.n3229 gnd 0.010593f
C5389 vdd.n3230 gnd 0.008527f
C5390 vdd.n3231 gnd 0.008527f
C5391 vdd.n3232 gnd 0.008527f
C5392 vdd.n3233 gnd 0.010593f
C5393 vdd.n3234 gnd 0.010593f
C5394 vdd.n3235 gnd 0.010593f
C5395 vdd.n3236 gnd 0.898564f
C5396 vdd.n3237 gnd 0.010593f
C5397 vdd.n3238 gnd 0.008527f
C5398 vdd.n3239 gnd 0.008527f
C5399 vdd.n3240 gnd 0.008527f
C5400 vdd.n3241 gnd 0.010593f
C5401 vdd.n3242 gnd 0.010593f
C5402 vdd.n3243 gnd 0.010593f
C5403 vdd.n3244 gnd 0.010593f
C5404 vdd.n3245 gnd 0.008527f
C5405 vdd.n3246 gnd 0.008527f
C5406 vdd.n3247 gnd 0.007077f
C5407 vdd.n3248 gnd 0.024124f
C5408 vdd.n3249 gnd 0.024289f
C5409 vdd.n3250 gnd 0.00405f
C5410 vdd.n3251 gnd 0.024289f
C5411 vdd.n3253 gnd 2.39256f
C5412 vdd.n3254 gnd 1.42904f
C5413 vdd.n3255 gnd 0.709108f
C5414 vdd.n3256 gnd 0.010593f
C5415 vdd.n3257 gnd 0.008527f
C5416 vdd.n3258 gnd 0.008527f
C5417 vdd.n3259 gnd 0.008527f
C5418 vdd.n3260 gnd 0.010593f
C5419 vdd.n3261 gnd 1.08261f
C5420 vdd.n3262 gnd 1.08261f
C5421 vdd.n3263 gnd 0.622499f
C5422 vdd.n3264 gnd 0.010593f
C5423 vdd.n3265 gnd 0.008527f
C5424 vdd.n3266 gnd 0.008527f
C5425 vdd.n3267 gnd 0.008527f
C5426 vdd.n3268 gnd 0.010593f
C5427 vdd.n3269 gnd 0.644151f
C5428 vdd.n3270 gnd 0.795717f
C5429 vdd.t171 gnd 0.541304f
C5430 vdd.n3271 gnd 0.828195f
C5431 vdd.n3272 gnd 0.010593f
C5432 vdd.n3273 gnd 0.008527f
C5433 vdd.n3274 gnd 0.008527f
C5434 vdd.n3275 gnd 0.008527f
C5435 vdd.n3276 gnd 0.010593f
C5436 vdd.n3277 gnd 0.898564f
C5437 vdd.t148 gnd 0.541304f
C5438 vdd.n3278 gnd 0.654978f
C5439 vdd.n3279 gnd 0.784891f
C5440 vdd.n3280 gnd 0.010593f
C5441 vdd.n3281 gnd 0.008527f
C5442 vdd.n3282 gnd 0.008527f
C5443 vdd.n3283 gnd 0.008527f
C5444 vdd.n3284 gnd 0.010593f
C5445 vdd.n3285 gnd 0.600847f
C5446 vdd.t132 gnd 0.541304f
C5447 vdd.n3286 gnd 0.898564f
C5448 vdd.t175 gnd 0.541304f
C5449 vdd.n3287 gnd 0.665804f
C5450 vdd.n3288 gnd 0.010593f
C5451 vdd.n3289 gnd 0.008527f
C5452 vdd.n3290 gnd 0.008142f
C5453 vdd.n3291 gnd 0.624846f
C5454 vdd.n3292 gnd 2.52207f
C5455 a_n6972_8799.t26 gnd 0.112027f
C5456 a_n6972_8799.t21 gnd 0.112027f
C5457 a_n6972_8799.t20 gnd 0.112027f
C5458 a_n6972_8799.n0 gnd 0.992109f
C5459 a_n6972_8799.t1 gnd 0.144034f
C5460 a_n6972_8799.t3 gnd 0.144034f
C5461 a_n6972_8799.n1 gnd 1.13602f
C5462 a_n6972_8799.t4 gnd 0.144034f
C5463 a_n6972_8799.t6 gnd 0.144034f
C5464 a_n6972_8799.n2 gnd 1.13415f
C5465 a_n6972_8799.n3 gnd 1.01946f
C5466 a_n6972_8799.t0 gnd 0.144034f
C5467 a_n6972_8799.t8 gnd 0.144034f
C5468 a_n6972_8799.n4 gnd 1.13415f
C5469 a_n6972_8799.n5 gnd 2.95084f
C5470 a_n6972_8799.t31 gnd 0.144034f
C5471 a_n6972_8799.t2 gnd 0.144034f
C5472 a_n6972_8799.n6 gnd 1.13602f
C5473 a_n6972_8799.t9 gnd 0.144034f
C5474 a_n6972_8799.t5 gnd 0.144034f
C5475 a_n6972_8799.n7 gnd 1.13415f
C5476 a_n6972_8799.n8 gnd 1.01946f
C5477 a_n6972_8799.t7 gnd 0.144034f
C5478 a_n6972_8799.t10 gnd 0.144034f
C5479 a_n6972_8799.n9 gnd 1.13415f
C5480 a_n6972_8799.n10 gnd 1.81107f
C5481 a_n6972_8799.n11 gnd 5.68596f
C5482 a_n6972_8799.n12 gnd 0.051915f
C5483 a_n6972_8799.t109 gnd 0.597234f
C5484 a_n6972_8799.n13 gnd 0.266736f
C5485 a_n6972_8799.n14 gnd 0.051915f
C5486 a_n6972_8799.n15 gnd 0.011781f
C5487 a_n6972_8799.t43 gnd 0.597234f
C5488 a_n6972_8799.n16 gnd 0.051915f
C5489 a_n6972_8799.t61 gnd 0.597234f
C5490 a_n6972_8799.n17 gnd 0.266576f
C5491 a_n6972_8799.t78 gnd 0.597234f
C5492 a_n6972_8799.n18 gnd 0.051915f
C5493 a_n6972_8799.n19 gnd 0.011781f
C5494 a_n6972_8799.t95 gnd 0.597234f
C5495 a_n6972_8799.n20 gnd 0.051915f
C5496 a_n6972_8799.t96 gnd 0.597234f
C5497 a_n6972_8799.n21 gnd 0.261775f
C5498 a_n6972_8799.t63 gnd 0.597234f
C5499 a_n6972_8799.n22 gnd 0.051915f
C5500 a_n6972_8799.t72 gnd 0.597234f
C5501 a_n6972_8799.n23 gnd 0.265936f
C5502 a_n6972_8799.t110 gnd 0.608538f
C5503 a_n6972_8799.n24 gnd 0.250387f
C5504 a_n6972_8799.n25 gnd 0.169752f
C5505 a_n6972_8799.n26 gnd 0.011781f
C5506 a_n6972_8799.t73 gnd 0.597234f
C5507 a_n6972_8799.n27 gnd 0.266736f
C5508 a_n6972_8799.n28 gnd 0.011781f
C5509 a_n6972_8799.n29 gnd 0.051915f
C5510 a_n6972_8799.n30 gnd 0.051915f
C5511 a_n6972_8799.n31 gnd 0.051915f
C5512 a_n6972_8799.n32 gnd 0.266256f
C5513 a_n6972_8799.n33 gnd 0.011781f
C5514 a_n6972_8799.t64 gnd 0.597234f
C5515 a_n6972_8799.n34 gnd 0.266736f
C5516 a_n6972_8799.n35 gnd 0.051915f
C5517 a_n6972_8799.n36 gnd 0.051915f
C5518 a_n6972_8799.n37 gnd 0.051915f
C5519 a_n6972_8799.n38 gnd 0.261455f
C5520 a_n6972_8799.t32 gnd 0.597234f
C5521 a_n6972_8799.n39 gnd 0.266576f
C5522 a_n6972_8799.n40 gnd 0.011781f
C5523 a_n6972_8799.n41 gnd 0.051915f
C5524 a_n6972_8799.n42 gnd 0.051915f
C5525 a_n6972_8799.n43 gnd 0.051915f
C5526 a_n6972_8799.n44 gnd 0.261455f
C5527 a_n6972_8799.n45 gnd 0.011781f
C5528 a_n6972_8799.t112 gnd 0.597234f
C5529 a_n6972_8799.n46 gnd 0.266736f
C5530 a_n6972_8799.n47 gnd 0.051915f
C5531 a_n6972_8799.n48 gnd 0.051915f
C5532 a_n6972_8799.n49 gnd 0.051915f
C5533 a_n6972_8799.n50 gnd 0.266256f
C5534 a_n6972_8799.t59 gnd 0.597234f
C5535 a_n6972_8799.n51 gnd 0.261775f
C5536 a_n6972_8799.n52 gnd 0.011781f
C5537 a_n6972_8799.n53 gnd 0.051915f
C5538 a_n6972_8799.n54 gnd 0.051915f
C5539 a_n6972_8799.n55 gnd 0.051915f
C5540 a_n6972_8799.n56 gnd 0.011781f
C5541 a_n6972_8799.t40 gnd 0.597234f
C5542 a_n6972_8799.n57 gnd 0.265936f
C5543 a_n6972_8799.t41 gnd 0.597234f
C5544 a_n6972_8799.n58 gnd 0.261295f
C5545 a_n6972_8799.n59 gnd 0.299123f
C5546 a_n6972_8799.n60 gnd 0.051915f
C5547 a_n6972_8799.t119 gnd 0.597234f
C5548 a_n6972_8799.n61 gnd 0.266736f
C5549 a_n6972_8799.n62 gnd 0.051915f
C5550 a_n6972_8799.n63 gnd 0.011781f
C5551 a_n6972_8799.t57 gnd 0.597234f
C5552 a_n6972_8799.n64 gnd 0.051915f
C5553 a_n6972_8799.t69 gnd 0.597234f
C5554 a_n6972_8799.n65 gnd 0.266576f
C5555 a_n6972_8799.t89 gnd 0.597234f
C5556 a_n6972_8799.n66 gnd 0.051915f
C5557 a_n6972_8799.n67 gnd 0.011781f
C5558 a_n6972_8799.t104 gnd 0.597234f
C5559 a_n6972_8799.n68 gnd 0.051915f
C5560 a_n6972_8799.t108 gnd 0.597234f
C5561 a_n6972_8799.n69 gnd 0.261775f
C5562 a_n6972_8799.t70 gnd 0.597234f
C5563 a_n6972_8799.n70 gnd 0.051915f
C5564 a_n6972_8799.t79 gnd 0.597234f
C5565 a_n6972_8799.n71 gnd 0.265936f
C5566 a_n6972_8799.t121 gnd 0.608538f
C5567 a_n6972_8799.n72 gnd 0.250387f
C5568 a_n6972_8799.n73 gnd 0.169752f
C5569 a_n6972_8799.n74 gnd 0.011781f
C5570 a_n6972_8799.t80 gnd 0.597234f
C5571 a_n6972_8799.n75 gnd 0.266736f
C5572 a_n6972_8799.n76 gnd 0.011781f
C5573 a_n6972_8799.n77 gnd 0.051915f
C5574 a_n6972_8799.n78 gnd 0.051915f
C5575 a_n6972_8799.n79 gnd 0.051915f
C5576 a_n6972_8799.n80 gnd 0.266256f
C5577 a_n6972_8799.n81 gnd 0.011781f
C5578 a_n6972_8799.t71 gnd 0.597234f
C5579 a_n6972_8799.n82 gnd 0.266736f
C5580 a_n6972_8799.n83 gnd 0.051915f
C5581 a_n6972_8799.n84 gnd 0.051915f
C5582 a_n6972_8799.n85 gnd 0.051915f
C5583 a_n6972_8799.n86 gnd 0.261455f
C5584 a_n6972_8799.t42 gnd 0.597234f
C5585 a_n6972_8799.n87 gnd 0.266576f
C5586 a_n6972_8799.n88 gnd 0.011781f
C5587 a_n6972_8799.n89 gnd 0.051915f
C5588 a_n6972_8799.n90 gnd 0.051915f
C5589 a_n6972_8799.n91 gnd 0.051915f
C5590 a_n6972_8799.n92 gnd 0.261455f
C5591 a_n6972_8799.n93 gnd 0.011781f
C5592 a_n6972_8799.t124 gnd 0.597234f
C5593 a_n6972_8799.n94 gnd 0.266736f
C5594 a_n6972_8799.n95 gnd 0.051915f
C5595 a_n6972_8799.n96 gnd 0.051915f
C5596 a_n6972_8799.n97 gnd 0.051915f
C5597 a_n6972_8799.n98 gnd 0.266256f
C5598 a_n6972_8799.t68 gnd 0.597234f
C5599 a_n6972_8799.n99 gnd 0.261775f
C5600 a_n6972_8799.n100 gnd 0.011781f
C5601 a_n6972_8799.n101 gnd 0.051915f
C5602 a_n6972_8799.n102 gnd 0.051915f
C5603 a_n6972_8799.n103 gnd 0.051915f
C5604 a_n6972_8799.n104 gnd 0.011781f
C5605 a_n6972_8799.t51 gnd 0.597234f
C5606 a_n6972_8799.n105 gnd 0.265936f
C5607 a_n6972_8799.t53 gnd 0.597234f
C5608 a_n6972_8799.n106 gnd 0.261295f
C5609 a_n6972_8799.n107 gnd 0.134499f
C5610 a_n6972_8799.n108 gnd 0.8995f
C5611 a_n6972_8799.n109 gnd 0.051915f
C5612 a_n6972_8799.t85 gnd 0.597234f
C5613 a_n6972_8799.n110 gnd 0.266736f
C5614 a_n6972_8799.n111 gnd 0.051915f
C5615 a_n6972_8799.n112 gnd 0.011781f
C5616 a_n6972_8799.t105 gnd 0.597234f
C5617 a_n6972_8799.n113 gnd 0.051915f
C5618 a_n6972_8799.t38 gnd 0.597234f
C5619 a_n6972_8799.n114 gnd 0.266576f
C5620 a_n6972_8799.t91 gnd 0.597234f
C5621 a_n6972_8799.n115 gnd 0.051915f
C5622 a_n6972_8799.n116 gnd 0.011781f
C5623 a_n6972_8799.t120 gnd 0.597234f
C5624 a_n6972_8799.n117 gnd 0.051915f
C5625 a_n6972_8799.t83 gnd 0.597234f
C5626 a_n6972_8799.n118 gnd 0.261775f
C5627 a_n6972_8799.t116 gnd 0.597234f
C5628 a_n6972_8799.n119 gnd 0.051915f
C5629 a_n6972_8799.t49 gnd 0.597234f
C5630 a_n6972_8799.n120 gnd 0.265936f
C5631 a_n6972_8799.t113 gnd 0.608538f
C5632 a_n6972_8799.n121 gnd 0.250387f
C5633 a_n6972_8799.n122 gnd 0.169752f
C5634 a_n6972_8799.n123 gnd 0.011781f
C5635 a_n6972_8799.t33 gnd 0.597234f
C5636 a_n6972_8799.n124 gnd 0.266736f
C5637 a_n6972_8799.n125 gnd 0.011781f
C5638 a_n6972_8799.n126 gnd 0.051915f
C5639 a_n6972_8799.n127 gnd 0.051915f
C5640 a_n6972_8799.n128 gnd 0.051915f
C5641 a_n6972_8799.n129 gnd 0.266256f
C5642 a_n6972_8799.n130 gnd 0.011781f
C5643 a_n6972_8799.t97 gnd 0.597234f
C5644 a_n6972_8799.n131 gnd 0.266736f
C5645 a_n6972_8799.n132 gnd 0.051915f
C5646 a_n6972_8799.n133 gnd 0.051915f
C5647 a_n6972_8799.n134 gnd 0.051915f
C5648 a_n6972_8799.n135 gnd 0.261455f
C5649 a_n6972_8799.t77 gnd 0.597234f
C5650 a_n6972_8799.n136 gnd 0.266576f
C5651 a_n6972_8799.n137 gnd 0.011781f
C5652 a_n6972_8799.n138 gnd 0.051915f
C5653 a_n6972_8799.n139 gnd 0.051915f
C5654 a_n6972_8799.n140 gnd 0.051915f
C5655 a_n6972_8799.n141 gnd 0.261455f
C5656 a_n6972_8799.n142 gnd 0.011781f
C5657 a_n6972_8799.t55 gnd 0.597234f
C5658 a_n6972_8799.n143 gnd 0.266736f
C5659 a_n6972_8799.n144 gnd 0.051915f
C5660 a_n6972_8799.n145 gnd 0.051915f
C5661 a_n6972_8799.n146 gnd 0.051915f
C5662 a_n6972_8799.n147 gnd 0.266256f
C5663 a_n6972_8799.t62 gnd 0.597234f
C5664 a_n6972_8799.n148 gnd 0.261775f
C5665 a_n6972_8799.n149 gnd 0.011781f
C5666 a_n6972_8799.n150 gnd 0.051915f
C5667 a_n6972_8799.n151 gnd 0.051915f
C5668 a_n6972_8799.n152 gnd 0.051915f
C5669 a_n6972_8799.n153 gnd 0.011781f
C5670 a_n6972_8799.t45 gnd 0.597234f
C5671 a_n6972_8799.n154 gnd 0.265936f
C5672 a_n6972_8799.t125 gnd 0.597234f
C5673 a_n6972_8799.n155 gnd 0.261295f
C5674 a_n6972_8799.n156 gnd 0.134499f
C5675 a_n6972_8799.n157 gnd 1.45854f
C5676 a_n6972_8799.n158 gnd 0.051915f
C5677 a_n6972_8799.t75 gnd 0.597234f
C5678 a_n6972_8799.t74 gnd 0.597234f
C5679 a_n6972_8799.t52 gnd 0.597234f
C5680 a_n6972_8799.n159 gnd 0.266736f
C5681 a_n6972_8799.n160 gnd 0.051915f
C5682 a_n6972_8799.t111 gnd 0.597234f
C5683 a_n6972_8799.t76 gnd 0.597234f
C5684 a_n6972_8799.n161 gnd 0.051915f
C5685 a_n6972_8799.t58 gnd 0.597234f
C5686 a_n6972_8799.n162 gnd 0.266736f
C5687 a_n6972_8799.n163 gnd 0.051915f
C5688 a_n6972_8799.t115 gnd 0.597234f
C5689 a_n6972_8799.t90 gnd 0.597234f
C5690 a_n6972_8799.n164 gnd 0.051915f
C5691 a_n6972_8799.t88 gnd 0.597234f
C5692 a_n6972_8799.n165 gnd 0.266576f
C5693 a_n6972_8799.n166 gnd 0.051915f
C5694 a_n6972_8799.t35 gnd 0.597234f
C5695 a_n6972_8799.t94 gnd 0.597234f
C5696 a_n6972_8799.n167 gnd 0.051915f
C5697 a_n6972_8799.t93 gnd 0.597234f
C5698 a_n6972_8799.n168 gnd 0.266256f
C5699 a_n6972_8799.n169 gnd 0.051915f
C5700 a_n6972_8799.t37 gnd 0.597234f
C5701 a_n6972_8799.t36 gnd 0.597234f
C5702 a_n6972_8799.n170 gnd 0.051915f
C5703 a_n6972_8799.t107 gnd 0.597234f
C5704 a_n6972_8799.n171 gnd 0.265936f
C5705 a_n6972_8799.t54 gnd 0.608538f
C5706 a_n6972_8799.n172 gnd 0.250387f
C5707 a_n6972_8799.n173 gnd 0.169752f
C5708 a_n6972_8799.n174 gnd 0.011781f
C5709 a_n6972_8799.n175 gnd 0.266736f
C5710 a_n6972_8799.n176 gnd 0.011781f
C5711 a_n6972_8799.n177 gnd 0.261775f
C5712 a_n6972_8799.n178 gnd 0.051915f
C5713 a_n6972_8799.n179 gnd 0.051915f
C5714 a_n6972_8799.n180 gnd 0.051915f
C5715 a_n6972_8799.n181 gnd 0.011781f
C5716 a_n6972_8799.n182 gnd 0.266736f
C5717 a_n6972_8799.n183 gnd 0.011781f
C5718 a_n6972_8799.n184 gnd 0.261455f
C5719 a_n6972_8799.n185 gnd 0.051915f
C5720 a_n6972_8799.n186 gnd 0.051915f
C5721 a_n6972_8799.n187 gnd 0.051915f
C5722 a_n6972_8799.n188 gnd 0.011781f
C5723 a_n6972_8799.n189 gnd 0.266576f
C5724 a_n6972_8799.n190 gnd 0.261455f
C5725 a_n6972_8799.n191 gnd 0.011781f
C5726 a_n6972_8799.n192 gnd 0.051915f
C5727 a_n6972_8799.n193 gnd 0.051915f
C5728 a_n6972_8799.n194 gnd 0.051915f
C5729 a_n6972_8799.n195 gnd 0.011781f
C5730 a_n6972_8799.n196 gnd 0.266256f
C5731 a_n6972_8799.n197 gnd 0.261775f
C5732 a_n6972_8799.n198 gnd 0.011781f
C5733 a_n6972_8799.n199 gnd 0.051915f
C5734 a_n6972_8799.n200 gnd 0.051915f
C5735 a_n6972_8799.n201 gnd 0.051915f
C5736 a_n6972_8799.n202 gnd 0.011781f
C5737 a_n6972_8799.n203 gnd 0.265936f
C5738 a_n6972_8799.n204 gnd 0.261295f
C5739 a_n6972_8799.n205 gnd 0.299123f
C5740 a_n6972_8799.n206 gnd 0.051915f
C5741 a_n6972_8799.t82 gnd 0.597234f
C5742 a_n6972_8799.t81 gnd 0.597234f
C5743 a_n6972_8799.t65 gnd 0.597234f
C5744 a_n6972_8799.n207 gnd 0.266736f
C5745 a_n6972_8799.n208 gnd 0.051915f
C5746 a_n6972_8799.t123 gnd 0.597234f
C5747 a_n6972_8799.t87 gnd 0.597234f
C5748 a_n6972_8799.n209 gnd 0.051915f
C5749 a_n6972_8799.t67 gnd 0.597234f
C5750 a_n6972_8799.n210 gnd 0.266736f
C5751 a_n6972_8799.n211 gnd 0.051915f
C5752 a_n6972_8799.t127 gnd 0.597234f
C5753 a_n6972_8799.t100 gnd 0.597234f
C5754 a_n6972_8799.n212 gnd 0.051915f
C5755 a_n6972_8799.t99 gnd 0.597234f
C5756 a_n6972_8799.n213 gnd 0.266576f
C5757 a_n6972_8799.n214 gnd 0.051915f
C5758 a_n6972_8799.t44 gnd 0.597234f
C5759 a_n6972_8799.t103 gnd 0.597234f
C5760 a_n6972_8799.n215 gnd 0.051915f
C5761 a_n6972_8799.t102 gnd 0.597234f
C5762 a_n6972_8799.n216 gnd 0.266256f
C5763 a_n6972_8799.n217 gnd 0.051915f
C5764 a_n6972_8799.t48 gnd 0.597234f
C5765 a_n6972_8799.t47 gnd 0.597234f
C5766 a_n6972_8799.n218 gnd 0.051915f
C5767 a_n6972_8799.t118 gnd 0.597234f
C5768 a_n6972_8799.n219 gnd 0.265936f
C5769 a_n6972_8799.t66 gnd 0.608538f
C5770 a_n6972_8799.n220 gnd 0.250387f
C5771 a_n6972_8799.n221 gnd 0.169752f
C5772 a_n6972_8799.n222 gnd 0.011781f
C5773 a_n6972_8799.n223 gnd 0.266736f
C5774 a_n6972_8799.n224 gnd 0.011781f
C5775 a_n6972_8799.n225 gnd 0.261775f
C5776 a_n6972_8799.n226 gnd 0.051915f
C5777 a_n6972_8799.n227 gnd 0.051915f
C5778 a_n6972_8799.n228 gnd 0.051915f
C5779 a_n6972_8799.n229 gnd 0.011781f
C5780 a_n6972_8799.n230 gnd 0.266736f
C5781 a_n6972_8799.n231 gnd 0.011781f
C5782 a_n6972_8799.n232 gnd 0.261455f
C5783 a_n6972_8799.n233 gnd 0.051915f
C5784 a_n6972_8799.n234 gnd 0.051915f
C5785 a_n6972_8799.n235 gnd 0.051915f
C5786 a_n6972_8799.n236 gnd 0.011781f
C5787 a_n6972_8799.n237 gnd 0.266576f
C5788 a_n6972_8799.n238 gnd 0.261455f
C5789 a_n6972_8799.n239 gnd 0.011781f
C5790 a_n6972_8799.n240 gnd 0.051915f
C5791 a_n6972_8799.n241 gnd 0.051915f
C5792 a_n6972_8799.n242 gnd 0.051915f
C5793 a_n6972_8799.n243 gnd 0.011781f
C5794 a_n6972_8799.n244 gnd 0.266256f
C5795 a_n6972_8799.n245 gnd 0.261775f
C5796 a_n6972_8799.n246 gnd 0.011781f
C5797 a_n6972_8799.n247 gnd 0.051915f
C5798 a_n6972_8799.n248 gnd 0.051915f
C5799 a_n6972_8799.n249 gnd 0.051915f
C5800 a_n6972_8799.n250 gnd 0.011781f
C5801 a_n6972_8799.n251 gnd 0.265936f
C5802 a_n6972_8799.n252 gnd 0.261295f
C5803 a_n6972_8799.n253 gnd 0.134499f
C5804 a_n6972_8799.n254 gnd 0.8995f
C5805 a_n6972_8799.n255 gnd 0.051915f
C5806 a_n6972_8799.t126 gnd 0.597234f
C5807 a_n6972_8799.t46 gnd 0.597234f
C5808 a_n6972_8799.t86 gnd 0.597234f
C5809 a_n6972_8799.n256 gnd 0.266736f
C5810 a_n6972_8799.n257 gnd 0.051915f
C5811 a_n6972_8799.t34 gnd 0.597234f
C5812 a_n6972_8799.t106 gnd 0.597234f
C5813 a_n6972_8799.n258 gnd 0.051915f
C5814 a_n6972_8799.t56 gnd 0.597234f
C5815 a_n6972_8799.n259 gnd 0.266736f
C5816 a_n6972_8799.n260 gnd 0.051915f
C5817 a_n6972_8799.t92 gnd 0.597234f
C5818 a_n6972_8799.t39 gnd 0.597234f
C5819 a_n6972_8799.n261 gnd 0.051915f
C5820 a_n6972_8799.t60 gnd 0.597234f
C5821 a_n6972_8799.n262 gnd 0.266576f
C5822 a_n6972_8799.n263 gnd 0.051915f
C5823 a_n6972_8799.t122 gnd 0.597234f
C5824 a_n6972_8799.t98 gnd 0.597234f
C5825 a_n6972_8799.n264 gnd 0.051915f
C5826 a_n6972_8799.t117 gnd 0.597234f
C5827 a_n6972_8799.n265 gnd 0.266256f
C5828 a_n6972_8799.n266 gnd 0.051915f
C5829 a_n6972_8799.t84 gnd 0.597234f
C5830 a_n6972_8799.t101 gnd 0.597234f
C5831 a_n6972_8799.n267 gnd 0.051915f
C5832 a_n6972_8799.t50 gnd 0.597234f
C5833 a_n6972_8799.n268 gnd 0.265936f
C5834 a_n6972_8799.t114 gnd 0.608538f
C5835 a_n6972_8799.n269 gnd 0.250387f
C5836 a_n6972_8799.n270 gnd 0.169752f
C5837 a_n6972_8799.n271 gnd 0.011781f
C5838 a_n6972_8799.n272 gnd 0.266736f
C5839 a_n6972_8799.n273 gnd 0.011781f
C5840 a_n6972_8799.n274 gnd 0.261775f
C5841 a_n6972_8799.n275 gnd 0.051915f
C5842 a_n6972_8799.n276 gnd 0.051915f
C5843 a_n6972_8799.n277 gnd 0.051915f
C5844 a_n6972_8799.n278 gnd 0.011781f
C5845 a_n6972_8799.n279 gnd 0.266736f
C5846 a_n6972_8799.n280 gnd 0.011781f
C5847 a_n6972_8799.n281 gnd 0.261455f
C5848 a_n6972_8799.n282 gnd 0.051915f
C5849 a_n6972_8799.n283 gnd 0.051915f
C5850 a_n6972_8799.n284 gnd 0.051915f
C5851 a_n6972_8799.n285 gnd 0.011781f
C5852 a_n6972_8799.n286 gnd 0.266576f
C5853 a_n6972_8799.n287 gnd 0.261455f
C5854 a_n6972_8799.n288 gnd 0.011781f
C5855 a_n6972_8799.n289 gnd 0.051915f
C5856 a_n6972_8799.n290 gnd 0.051915f
C5857 a_n6972_8799.n291 gnd 0.051915f
C5858 a_n6972_8799.n292 gnd 0.011781f
C5859 a_n6972_8799.n293 gnd 0.266256f
C5860 a_n6972_8799.n294 gnd 0.261775f
C5861 a_n6972_8799.n295 gnd 0.011781f
C5862 a_n6972_8799.n296 gnd 0.051915f
C5863 a_n6972_8799.n297 gnd 0.051915f
C5864 a_n6972_8799.n298 gnd 0.051915f
C5865 a_n6972_8799.n299 gnd 0.011781f
C5866 a_n6972_8799.n300 gnd 0.265936f
C5867 a_n6972_8799.n301 gnd 0.261295f
C5868 a_n6972_8799.n302 gnd 0.134499f
C5869 a_n6972_8799.n303 gnd 1.13233f
C5870 a_n6972_8799.n304 gnd 12.2315f
C5871 a_n6972_8799.n305 gnd 4.37088f
C5872 a_n6972_8799.t17 gnd 0.112027f
C5873 a_n6972_8799.t18 gnd 0.112027f
C5874 a_n6972_8799.n306 gnd 0.992109f
C5875 a_n6972_8799.t13 gnd 0.112027f
C5876 a_n6972_8799.t14 gnd 0.112027f
C5877 a_n6972_8799.n307 gnd 0.989908f
C5878 a_n6972_8799.n308 gnd 0.788507f
C5879 a_n6972_8799.t12 gnd 0.112027f
C5880 a_n6972_8799.t27 gnd 0.112027f
C5881 a_n6972_8799.n309 gnd 0.989908f
C5882 a_n6972_8799.n310 gnd 0.741378f
C5883 a_n6972_8799.t28 gnd 0.112027f
C5884 a_n6972_8799.t23 gnd 0.112027f
C5885 a_n6972_8799.n311 gnd 0.989908f
C5886 a_n6972_8799.n312 gnd 0.387197f
C5887 a_n6972_8799.t25 gnd 0.112027f
C5888 a_n6972_8799.t11 gnd 0.112027f
C5889 a_n6972_8799.n313 gnd 0.989908f
C5890 a_n6972_8799.n314 gnd 2.70813f
C5891 a_n6972_8799.t24 gnd 0.112027f
C5892 a_n6972_8799.t22 gnd 0.112027f
C5893 a_n6972_8799.n315 gnd 0.992109f
C5894 a_n6972_8799.t15 gnd 0.112027f
C5895 a_n6972_8799.t19 gnd 0.112027f
C5896 a_n6972_8799.n316 gnd 0.989907f
C5897 a_n6972_8799.n317 gnd 0.788509f
C5898 a_n6972_8799.t29 gnd 0.112027f
C5899 a_n6972_8799.t16 gnd 0.112027f
C5900 a_n6972_8799.n318 gnd 0.989907f
C5901 a_n6972_8799.n319 gnd 2.4653f
C5902 a_n6972_8799.n320 gnd 0.788511f
C5903 a_n6972_8799.n321 gnd 0.989904f
C5904 a_n6972_8799.t30 gnd 0.112027f
C5905 a_n3827_n3924.n0 gnd 1.70953f
C5906 a_n3827_n3924.n1 gnd 0.682769f
C5907 a_n3827_n3924.n2 gnd 1.24153f
C5908 a_n3827_n3924.n3 gnd 1.20073f
C5909 a_n3827_n3924.n4 gnd 1.70952f
C5910 a_n3827_n3924.n5 gnd 0.682766f
C5911 a_n3827_n3924.n6 gnd 1.54211f
C5912 a_n3827_n3924.n7 gnd 2.34829f
C5913 a_n3827_n3924.n8 gnd 1.67197f
C5914 a_n3827_n3924.n9 gnd 1.67197f
C5915 a_n3827_n3924.n10 gnd 2.84498f
C5916 a_n3827_n3924.n11 gnd 0.900148f
C5917 a_n3827_n3924.t19 gnd 0.091917f
C5918 a_n3827_n3924.t11 gnd 0.091917f
C5919 a_n3827_n3924.n12 gnd 0.750696f
C5920 a_n3827_n3924.t29 gnd 0.955301f
C5921 a_n3827_n3924.t39 gnd 0.091917f
C5922 a_n3827_n3924.t28 gnd 0.091917f
C5923 a_n3827_n3924.n13 gnd 0.750697f
C5924 a_n3827_n3924.t42 gnd 0.091917f
C5925 a_n3827_n3924.t41 gnd 0.091917f
C5926 a_n3827_n3924.n14 gnd 0.750697f
C5927 a_n3827_n3924.t27 gnd 0.091917f
C5928 a_n3827_n3924.t37 gnd 0.091917f
C5929 a_n3827_n3924.n15 gnd 0.750697f
C5930 a_n3827_n3924.t38 gnd 0.091917f
C5931 a_n3827_n3924.t45 gnd 0.091917f
C5932 a_n3827_n3924.n16 gnd 0.750697f
C5933 a_n3827_n3924.t40 gnd 0.955305f
C5934 a_n3827_n3924.t16 gnd 0.955305f
C5935 a_n3827_n3924.t2 gnd 0.091917f
C5936 a_n3827_n3924.t17 gnd 0.091917f
C5937 a_n3827_n3924.n17 gnd 0.750697f
C5938 a_n3827_n3924.t23 gnd 0.091917f
C5939 a_n3827_n3924.t12 gnd 0.091917f
C5940 a_n3827_n3924.n18 gnd 0.750697f
C5941 a_n3827_n3924.t14 gnd 0.091917f
C5942 a_n3827_n3924.t1 gnd 0.091917f
C5943 a_n3827_n3924.n19 gnd 0.750697f
C5944 a_n3827_n3924.t8 gnd 0.091917f
C5945 a_n3827_n3924.t18 gnd 0.091917f
C5946 a_n3827_n3924.n20 gnd 0.750697f
C5947 a_n3827_n3924.t46 gnd 0.955305f
C5948 a_n3827_n3924.t5 gnd 0.091917f
C5949 a_n3827_n3924.t24 gnd 0.091917f
C5950 a_n3827_n3924.n21 gnd 0.750696f
C5951 a_n3827_n3924.t6 gnd 0.091917f
C5952 a_n3827_n3924.t9 gnd 0.091917f
C5953 a_n3827_n3924.n22 gnd 0.750696f
C5954 a_n3827_n3924.t22 gnd 0.955301f
C5955 a_n3827_n3924.t30 gnd 0.955301f
C5956 a_n3827_n3924.t36 gnd 0.091917f
C5957 a_n3827_n3924.t32 gnd 0.091917f
C5958 a_n3827_n3924.n23 gnd 0.750696f
C5959 a_n3827_n3924.t35 gnd 0.091917f
C5960 a_n3827_n3924.t44 gnd 0.091917f
C5961 a_n3827_n3924.n24 gnd 0.750696f
C5962 a_n3827_n3924.t33 gnd 0.091917f
C5963 a_n3827_n3924.t26 gnd 0.091917f
C5964 a_n3827_n3924.n25 gnd 0.750696f
C5965 a_n3827_n3924.t34 gnd 0.091917f
C5966 a_n3827_n3924.t43 gnd 0.091917f
C5967 a_n3827_n3924.n26 gnd 0.750696f
C5968 a_n3827_n3924.t31 gnd 0.955301f
C5969 a_n3827_n3924.n27 gnd 0.862207f
C5970 a_n3827_n3924.t20 gnd 1.18864f
C5971 a_n3827_n3924.t49 gnd 1.18694f
C5972 a_n3827_n3924.t10 gnd 1.18694f
C5973 a_n3827_n3924.t25 gnd 1.18694f
C5974 a_n3827_n3924.t47 gnd 1.18694f
C5975 a_n3827_n3924.t21 gnd 1.18694f
C5976 a_n3827_n3924.t7 gnd 1.18694f
C5977 a_n3827_n3924.t15 gnd 1.18694f
C5978 a_n3827_n3924.t13 gnd 1.19019f
C5979 a_n3827_n3924.t48 gnd 1.18694f
C5980 a_n3827_n3924.n28 gnd 0.862207f
C5981 a_n3827_n3924.t4 gnd 0.955301f
C5982 a_n3827_n3924.t3 gnd 0.091917f
C5983 a_n3827_n3924.n29 gnd 0.750693f
C5984 a_n3827_n3924.t0 gnd 0.091917f
C5985 plus.n0 gnd 0.022293f
C5986 plus.t14 gnd 0.315318f
C5987 plus.n1 gnd 0.022293f
C5988 plus.t15 gnd 0.315318f
C5989 plus.t9 gnd 0.315318f
C5990 plus.n2 gnd 0.140074f
C5991 plus.n3 gnd 0.022293f
C5992 plus.t5 gnd 0.315318f
C5993 plus.t6 gnd 0.315318f
C5994 plus.n4 gnd 0.140074f
C5995 plus.n5 gnd 0.022293f
C5996 plus.t19 gnd 0.315318f
C5997 plus.t20 gnd 0.315318f
C5998 plus.n6 gnd 0.140074f
C5999 plus.n7 gnd 0.022293f
C6000 plus.t16 gnd 0.315318f
C6001 plus.t11 gnd 0.315318f
C6002 plus.n8 gnd 0.143803f
C6003 plus.t13 gnd 0.326365f
C6004 plus.n9 gnd 0.130628f
C6005 plus.n10 gnd 0.095157f
C6006 plus.n11 gnd 0.005059f
C6007 plus.n12 gnd 0.140074f
C6008 plus.n13 gnd 0.005059f
C6009 plus.n14 gnd 0.022293f
C6010 plus.n15 gnd 0.022293f
C6011 plus.n16 gnd 0.022293f
C6012 plus.n17 gnd 0.005059f
C6013 plus.n18 gnd 0.140074f
C6014 plus.n19 gnd 0.005059f
C6015 plus.n20 gnd 0.022293f
C6016 plus.n21 gnd 0.022293f
C6017 plus.n22 gnd 0.022293f
C6018 plus.n23 gnd 0.005059f
C6019 plus.n24 gnd 0.140074f
C6020 plus.n25 gnd 0.005059f
C6021 plus.n26 gnd 0.022293f
C6022 plus.n27 gnd 0.022293f
C6023 plus.n28 gnd 0.022293f
C6024 plus.n29 gnd 0.005059f
C6025 plus.n30 gnd 0.140074f
C6026 plus.n31 gnd 0.005059f
C6027 plus.n32 gnd 0.139868f
C6028 plus.n33 gnd 0.251839f
C6029 plus.n34 gnd 0.022293f
C6030 plus.n35 gnd 0.005059f
C6031 plus.t10 gnd 0.315318f
C6032 plus.n36 gnd 0.022293f
C6033 plus.n37 gnd 0.005059f
C6034 plus.t7 gnd 0.315318f
C6035 plus.n38 gnd 0.022293f
C6036 plus.n39 gnd 0.005059f
C6037 plus.t23 gnd 0.315318f
C6038 plus.n40 gnd 0.022293f
C6039 plus.n41 gnd 0.005059f
C6040 plus.t22 gnd 0.315318f
C6041 plus.t18 gnd 0.326365f
C6042 plus.t17 gnd 0.315318f
C6043 plus.n42 gnd 0.143803f
C6044 plus.n43 gnd 0.130628f
C6045 plus.n44 gnd 0.095157f
C6046 plus.n45 gnd 0.022293f
C6047 plus.n46 gnd 0.140074f
C6048 plus.n47 gnd 0.005059f
C6049 plus.t21 gnd 0.315318f
C6050 plus.n48 gnd 0.140074f
C6051 plus.n49 gnd 0.022293f
C6052 plus.n50 gnd 0.022293f
C6053 plus.n51 gnd 0.022293f
C6054 plus.n52 gnd 0.140074f
C6055 plus.n53 gnd 0.005059f
C6056 plus.t8 gnd 0.315318f
C6057 plus.n54 gnd 0.140074f
C6058 plus.n55 gnd 0.022293f
C6059 plus.n56 gnd 0.022293f
C6060 plus.n57 gnd 0.022293f
C6061 plus.n58 gnd 0.140074f
C6062 plus.n59 gnd 0.005059f
C6063 plus.t12 gnd 0.315318f
C6064 plus.n60 gnd 0.140074f
C6065 plus.n61 gnd 0.022293f
C6066 plus.n62 gnd 0.022293f
C6067 plus.n63 gnd 0.022293f
C6068 plus.n64 gnd 0.140074f
C6069 plus.n65 gnd 0.005059f
C6070 plus.t24 gnd 0.315318f
C6071 plus.n66 gnd 0.139868f
C6072 plus.n67 gnd 0.687659f
C6073 plus.n68 gnd 1.03991f
C6074 plus.t3 gnd 0.038485f
C6075 plus.t1 gnd 0.006872f
C6076 plus.t2 gnd 0.006872f
C6077 plus.n69 gnd 0.022288f
C6078 plus.n70 gnd 0.173026f
C6079 plus.t4 gnd 0.006872f
C6080 plus.t0 gnd 0.006872f
C6081 plus.n71 gnd 0.022288f
C6082 plus.n72 gnd 0.129877f
C6083 plus.n73 gnd 2.95718f
.ends

