* NGSPICE file created from opamp154.ext - technology: sky130A

.subckt opamp154 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 CSoutput.t192 a_n7636_8799.t32 vdd.t290 vdd.t230 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X1 gnd.t341 commonsourceibias.t24 commonsourceibias.t25 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X2 a_n7636_8799.t18 plus.t5 a_n3827_n3924.t21 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X3 a_n1808_13878.t19 a_n1996_n452.t36 a_n1996_n452.t37 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 a_n1808_13878.t7 a_n1996_n452.t44 vdd.t123 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 CSoutput.t42 commonsourceibias.t64 gnd.t340 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X6 vdd.t289 a_n7636_8799.t33 CSoutput.t191 vdd.t224 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X7 CSoutput.t190 a_n7636_8799.t34 vdd.t288 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X8 commonsourceibias.t23 commonsourceibias.t22 gnd.t339 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 gnd.t338 commonsourceibias.t65 CSoutput.t43 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 gnd.t130 gnd.t128 plus.t4 gnd.t129 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X11 gnd.t337 commonsourceibias.t20 commonsourceibias.t21 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X12 a_n3827_n3924.t0 diffpairibias.t20 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X13 CSoutput.t189 a_n7636_8799.t35 vdd.t287 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X14 a_n3827_n3924.t20 plus.t6 a_n7636_8799.t26 gnd.t161 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X15 gnd.t336 commonsourceibias.t18 commonsourceibias.t19 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 vdd.t86 vdd.t84 vdd.t85 vdd.t38 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X17 a_n3827_n3924.t32 minus.t5 a_n1996_n452.t8 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X18 a_n1986_8322.t19 a_n1996_n452.t45 a_n7636_8799.t31 vdd.t129 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X19 commonsourceibias.t15 commonsourceibias.t14 gnd.t335 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 gnd.t334 commonsourceibias.t66 CSoutput.t209 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X21 CSoutput.t188 a_n7636_8799.t36 vdd.t286 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X22 vdd.t285 a_n7636_8799.t37 CSoutput.t187 vdd.t218 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X23 a_n1996_n452.t6 minus.t6 a_n3827_n3924.t30 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X24 gnd.t127 gnd.t125 gnd.t126 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X25 gnd.t124 gnd.t121 gnd.t123 gnd.t122 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X26 vdd.t284 a_n7636_8799.t38 CSoutput.t186 vdd.t247 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X27 a_n1996_n452.t13 minus.t7 a_n3827_n3924.t38 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X28 CSoutput.t185 a_n7636_8799.t39 vdd.t283 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X29 vdd.t282 a_n7636_8799.t40 CSoutput.t184 vdd.t244 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X30 vdd.t281 a_n7636_8799.t41 CSoutput.t183 vdd.t269 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X31 commonsourceibias.t13 commonsourceibias.t12 gnd.t333 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 a_n7636_8799.t17 a_n1996_n452.t46 a_n1986_8322.t18 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X33 CSoutput.t182 a_n7636_8799.t42 vdd.t280 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X34 gnd.t332 commonsourceibias.t67 CSoutput.t210 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 CSoutput.t198 commonsourceibias.t68 gnd.t331 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 a_n3827_n3924.t42 minus.t8 a_n1996_n452.t39 gnd.t137 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X37 gnd.t330 commonsourceibias.t10 commonsourceibias.t11 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X38 CSoutput.t216 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X39 CSoutput.t199 commonsourceibias.t69 gnd.t329 gnd.t265 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 CSoutput.t181 a_n7636_8799.t43 vdd.t279 vdd.t230 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X41 vdd.t83 vdd.t81 vdd.t82 vdd.t16 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X42 CSoutput.t180 a_n7636_8799.t44 vdd.t278 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X43 a_n3827_n3924.t24 diffpairibias.t21 gnd.t10 gnd.t9 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X44 commonsourceibias.t29 commonsourceibias.t28 gnd.t312 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X45 CSoutput.t68 commonsourceibias.t70 gnd.t328 gnd.t265 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X46 CSoutput.t179 a_n7636_8799.t45 vdd.t277 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X47 a_n3827_n3924.t19 plus.t7 a_n7636_8799.t0 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X48 gnd.t327 commonsourceibias.t8 commonsourceibias.t9 gnd.t250 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 CSoutput.t69 commonsourceibias.t71 gnd.t326 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X50 a_n1808_13878.t18 a_n1996_n452.t16 a_n1996_n452.t17 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X51 vdd.t276 a_n7636_8799.t46 CSoutput.t178 vdd.t269 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X52 vdd.t80 vdd.t78 vdd.t79 vdd.t38 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X53 CSoutput.t177 a_n7636_8799.t47 vdd.t275 vdd.t222 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X54 a_n1996_n452.t35 a_n1996_n452.t34 a_n1808_13878.t17 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X55 output.t3 outputibias.t8 gnd.t179 gnd.t178 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X56 CSoutput.t217 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X57 a_n7636_8799.t10 plus.t8 a_n3827_n3924.t18 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X58 CSoutput.t176 a_n7636_8799.t48 vdd.t274 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X59 vdd.t77 vdd.t75 vdd.t76 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X60 vdd.t273 a_n7636_8799.t49 CSoutput.t175 vdd.t218 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 vdd.t108 CSoutput.t218 output.t19 gnd.t357 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X62 diffpairibias.t19 diffpairibias.t18 gnd.t363 gnd.t362 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X63 CSoutput.t52 commonsourceibias.t72 gnd.t325 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X64 a_n1996_n452.t42 minus.t9 a_n3827_n3924.t46 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X65 CSoutput.t53 commonsourceibias.t73 gnd.t324 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X66 CSoutput.t14 commonsourceibias.t74 gnd.t323 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 CSoutput.t174 a_n7636_8799.t50 vdd.t272 vdd.t226 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X68 commonsourceibias.t55 commonsourceibias.t54 gnd.t322 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X69 gnd.t120 gnd.t118 gnd.t119 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X70 vdd.t229 a_n7636_8799.t51 CSoutput.t173 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 vdd.t271 a_n7636_8799.t52 CSoutput.t172 vdd.t244 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 vdd.t270 a_n7636_8799.t53 CSoutput.t171 vdd.t269 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X73 vdd.t268 a_n7636_8799.t54 CSoutput.t170 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 plus.t3 gnd.t115 gnd.t117 gnd.t116 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X75 diffpairibias.t17 diffpairibias.t16 gnd.t361 gnd.t360 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X76 CSoutput.t169 a_n7636_8799.t55 vdd.t267 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X77 CSoutput.t168 a_n7636_8799.t56 vdd.t266 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X78 gnd.t114 gnd.t112 gnd.t113 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X79 gnd.t111 gnd.t109 gnd.t110 gnd.t30 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X80 vdd.t234 a_n7636_8799.t57 CSoutput.t167 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 CSoutput.t15 commonsourceibias.t75 gnd.t321 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 CSoutput.t166 a_n7636_8799.t58 vdd.t265 vdd.t252 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 CSoutput.t165 a_n7636_8799.t59 vdd.t264 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X84 CSoutput.t164 a_n7636_8799.t60 vdd.t263 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X85 CSoutput.t163 a_n7636_8799.t61 vdd.t262 vdd.t252 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 vdd.t261 a_n7636_8799.t62 CSoutput.t162 vdd.t249 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X87 gnd.t320 commonsourceibias.t76 CSoutput.t59 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 gnd.t108 gnd.t105 gnd.t107 gnd.t106 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X89 CSoutput.t60 commonsourceibias.t77 gnd.t319 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 gnd.t318 commonsourceibias.t78 CSoutput.t19 gnd.t205 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X91 a_n3827_n3924.t17 plus.t9 a_n7636_8799.t11 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X92 gnd.t104 gnd.t102 gnd.t103 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X93 a_n3827_n3924.t25 diffpairibias.t22 gnd.t136 gnd.t135 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X94 vdd.t260 a_n7636_8799.t63 CSoutput.t161 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X95 CSoutput.t20 commonsourceibias.t79 gnd.t317 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X96 a_n1996_n452.t31 a_n1996_n452.t30 a_n1808_13878.t16 vdd.t129 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X97 vdd.t259 a_n7636_8799.t64 CSoutput.t160 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X98 vdd.t258 a_n7636_8799.t65 CSoutput.t159 vdd.t247 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X99 a_n7636_8799.t30 a_n1996_n452.t47 a_n1986_8322.t17 vdd.t99 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X100 a_n1996_n452.t27 a_n1996_n452.t26 a_n1808_13878.t15 vdd.t124 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X101 vdd.t257 a_n7636_8799.t66 CSoutput.t158 vdd.t249 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 outputibias.t7 outputibias.t6 gnd.t147 gnd.t146 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X103 commonsourceibias.t53 commonsourceibias.t52 gnd.t316 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 gnd.t315 commonsourceibias.t80 CSoutput.t23 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X105 gnd.t101 gnd.t99 gnd.t100 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X106 CSoutput.t24 commonsourceibias.t81 gnd.t314 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X107 vdd.t256 a_n7636_8799.t67 CSoutput.t157 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X108 gnd.t313 commonsourceibias.t30 commonsourceibias.t31 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 CSoutput.t156 a_n7636_8799.t68 vdd.t239 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X110 CSoutput.t35 commonsourceibias.t82 gnd.t311 gnd.t265 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X111 diffpairibias.t15 diffpairibias.t14 gnd.t172 gnd.t171 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X112 a_n1996_n452.t40 minus.t10 a_n3827_n3924.t43 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X113 vdd.t74 vdd.t72 vdd.t73 vdd.t59 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X114 vdd.t255 a_n7636_8799.t69 CSoutput.t155 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X115 CSoutput.t154 a_n7636_8799.t70 vdd.t254 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X116 vdd.t71 vdd.t68 vdd.t70 vdd.t69 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X117 gnd.t310 commonsourceibias.t83 CSoutput.t36 gnd.t213 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X118 a_n3827_n3924.t47 minus.t11 a_n1996_n452.t43 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X119 vdd.t67 vdd.t65 vdd.t66 vdd.t12 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X120 vdd.t64 vdd.t62 vdd.t63 vdd.t55 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X121 vdd.t110 a_n1996_n452.t48 a_n1986_8322.t7 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X122 gnd.t307 commonsourceibias.t26 commonsourceibias.t27 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X123 CSoutput.t31 commonsourceibias.t84 gnd.t309 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X124 output.t18 CSoutput.t219 vdd.t104 gnd.t356 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X125 CSoutput.t32 commonsourceibias.t85 gnd.t308 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X126 a_n1986_8322.t6 a_n1996_n452.t49 vdd.t95 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X127 a_n3827_n3924.t44 diffpairibias.t23 gnd.t181 gnd.t180 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X128 CSoutput.t153 a_n7636_8799.t71 vdd.t253 vdd.t252 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X129 CSoutput.t152 a_n7636_8799.t72 vdd.t251 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X130 gnd.t306 commonsourceibias.t86 CSoutput.t27 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X131 gnd.t98 gnd.t96 gnd.t97 gnd.t41 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X132 vdd.t250 a_n7636_8799.t73 CSoutput.t151 vdd.t249 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X133 a_n3827_n3924.t33 minus.t12 a_n1996_n452.t9 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X134 commonsourceibias.t41 commonsourceibias.t40 gnd.t296 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X135 vdd.t2 a_n1996_n452.t50 a_n1808_13878.t6 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X136 gnd.t305 commonsourceibias.t87 CSoutput.t28 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X137 a_n1996_n452.t12 minus.t13 a_n3827_n3924.t37 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X138 a_n3827_n3924.t16 plus.t10 a_n7636_8799.t3 gnd.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X139 a_n3827_n3924.t15 plus.t11 a_n7636_8799.t16 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X140 vdd.t61 vdd.t58 vdd.t60 vdd.t59 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X141 gnd.t304 commonsourceibias.t46 commonsourceibias.t47 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X142 output.t17 CSoutput.t220 vdd.t105 gnd.t355 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X143 CSoutput.t205 commonsourceibias.t88 gnd.t303 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X144 gnd.t302 commonsourceibias.t89 CSoutput.t206 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X145 vdd.t57 vdd.t54 vdd.t56 vdd.t55 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X146 vdd.t248 a_n7636_8799.t74 CSoutput.t150 vdd.t247 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X147 CSoutput.t61 commonsourceibias.t90 gnd.t301 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X148 a_n7636_8799.t29 plus.t12 a_n3827_n3924.t14 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X149 a_n7636_8799.t21 plus.t13 a_n3827_n3924.t13 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X150 commonsourceibias.t45 commonsourceibias.t44 gnd.t300 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X151 vdd.t53 vdd.t50 vdd.t52 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X152 a_n1986_8322.t5 a_n1996_n452.t51 vdd.t295 vdd.t294 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X153 a_n7636_8799.t28 a_n1996_n452.t52 a_n1986_8322.t16 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X154 gnd.t299 commonsourceibias.t91 CSoutput.t62 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X155 gnd.t95 gnd.t93 gnd.t94 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X156 CSoutput.t149 a_n7636_8799.t75 vdd.t246 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X157 diffpairibias.t13 diffpairibias.t12 gnd.t160 gnd.t159 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X158 vdd.t245 a_n7636_8799.t76 CSoutput.t148 vdd.t244 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 a_n1996_n452.t38 minus.t14 a_n3827_n3924.t41 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X160 a_n1996_n452.t21 a_n1996_n452.t20 a_n1808_13878.t14 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X161 vdd.t243 a_n7636_8799.t77 CSoutput.t147 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X162 a_n7636_8799.t22 a_n1996_n452.t53 a_n1986_8322.t15 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X163 CSoutput.t146 a_n7636_8799.t78 vdd.t242 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X164 gnd.t298 commonsourceibias.t42 commonsourceibias.t43 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 a_n1808_13878.t13 a_n1996_n452.t32 a_n1996_n452.t33 vdd.t99 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X166 gnd.t92 gnd.t90 minus.t4 gnd.t91 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X167 a_n3827_n3924.t1 minus.t15 a_n1996_n452.t0 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X168 gnd.t297 commonsourceibias.t92 CSoutput.t37 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 output.t16 CSoutput.t221 vdd.t106 gnd.t354 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X170 gnd.t295 commonsourceibias.t93 CSoutput.t38 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X171 CSoutput.t145 a_n7636_8799.t79 vdd.t241 vdd.t226 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X172 vdd.t4 a_n1996_n452.t54 a_n1986_8322.t4 vdd.t3 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X173 gnd.t89 gnd.t87 gnd.t88 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X174 vdd.t240 a_n7636_8799.t80 CSoutput.t144 vdd.t224 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X175 output.t2 outputibias.t9 gnd.t365 gnd.t364 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X176 gnd.t86 gnd.t83 gnd.t85 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X177 gnd.t82 gnd.t80 gnd.t81 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X178 CSoutput.t143 a_n7636_8799.t81 vdd.t238 vdd.t222 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X179 outputibias.t5 outputibias.t4 gnd.t134 gnd.t133 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X180 vdd.t107 CSoutput.t222 output.t15 gnd.t353 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X181 vdd.t237 a_n7636_8799.t82 CSoutput.t142 vdd.t137 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X182 CSoutput.t44 commonsourceibias.t94 gnd.t294 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 gnd.t293 commonsourceibias.t95 CSoutput.t45 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X184 a_n3827_n3924.t12 plus.t14 a_n7636_8799.t2 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X185 gnd.t292 commonsourceibias.t96 CSoutput.t200 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X186 gnd.t79 gnd.t77 minus.t3 gnd.t78 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X187 vdd.t236 a_n7636_8799.t83 CSoutput.t141 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X188 a_n3827_n3924.t40 diffpairibias.t24 gnd.t177 gnd.t176 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X189 a_n3827_n3924.t39 diffpairibias.t25 gnd.t175 gnd.t174 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X190 outputibias.t3 outputibias.t2 gnd.t158 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X191 vdd.t235 a_n7636_8799.t84 CSoutput.t140 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X192 vdd.t233 a_n7636_8799.t85 CSoutput.t139 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X193 a_n7636_8799.t23 plus.t15 a_n3827_n3924.t11 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X194 gnd.t76 gnd.t74 gnd.t75 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X195 gnd.t73 gnd.t71 gnd.t72 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X196 CSoutput.t138 a_n7636_8799.t86 vdd.t232 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X197 CSoutput.t137 a_n7636_8799.t87 vdd.t231 vdd.t230 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X198 vdd.t100 CSoutput.t223 output.t14 gnd.t352 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X199 CSoutput.t136 a_n7636_8799.t88 vdd.t228 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X200 CSoutput.t1 commonsourceibias.t97 gnd.t291 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 output.t13 CSoutput.t224 vdd.t101 gnd.t351 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X202 gnd.t70 gnd.t68 gnd.t69 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X203 gnd.t290 commonsourceibias.t98 CSoutput.t67 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X204 diffpairibias.t11 diffpairibias.t10 gnd.t166 gnd.t165 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X205 a_n1808_13878.t5 a_n1996_n452.t55 vdd.t120 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X206 vdd.t49 vdd.t47 vdd.t48 vdd.t23 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X207 vdd.t6 a_n1996_n452.t56 a_n1808_13878.t4 vdd.t5 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X208 vdd.t46 vdd.t44 vdd.t45 vdd.t31 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X209 CSoutput.t135 a_n7636_8799.t89 vdd.t227 vdd.t226 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X210 gnd.t289 commonsourceibias.t99 CSoutput.t46 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X211 CSoutput.t2 commonsourceibias.t100 gnd.t288 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X212 vdd.t225 a_n7636_8799.t90 CSoutput.t134 vdd.t224 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X213 output.t12 CSoutput.t225 vdd.t102 gnd.t350 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X214 vdd.t43 vdd.t41 vdd.t42 vdd.t31 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X215 diffpairibias.t9 diffpairibias.t8 gnd.t359 gnd.t358 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X216 gnd.t287 commonsourceibias.t101 CSoutput.t47 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X217 a_n3827_n3924.t26 minus.t16 a_n1996_n452.t3 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X218 CSoutput.t133 a_n7636_8799.t91 vdd.t223 vdd.t222 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X219 vdd.t216 a_n7636_8799.t92 CSoutput.t132 vdd.t137 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X220 vdd.t221 a_n7636_8799.t93 CSoutput.t131 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X221 commonsourceibias.t33 commonsourceibias.t32 gnd.t286 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X222 a_n1986_8322.t14 a_n1996_n452.t57 a_n7636_8799.t27 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X223 CSoutput.t130 a_n7636_8799.t94 vdd.t220 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X224 outputibias.t1 outputibias.t0 gnd.t153 gnd.t152 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X225 diffpairibias.t7 diffpairibias.t6 gnd.t150 gnd.t149 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X226 vdd.t219 a_n7636_8799.t95 CSoutput.t129 vdd.t218 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X227 a_n1996_n452.t1 minus.t17 a_n3827_n3924.t22 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X228 CSoutput.t128 a_n7636_8799.t96 vdd.t217 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 a_n1996_n452.t41 minus.t18 a_n3827_n3924.t45 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X230 vdd.t215 a_n7636_8799.t97 CSoutput.t127 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X231 plus.t2 gnd.t65 gnd.t67 gnd.t66 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X232 vdd.t88 a_n1996_n452.t58 a_n1986_8322.t3 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X233 vdd.t213 a_n7636_8799.t98 CSoutput.t126 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X234 vdd.t212 a_n7636_8799.t99 CSoutput.t125 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X235 output.t1 outputibias.t10 gnd.t156 gnd.t155 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X236 CSoutput.t211 commonsourceibias.t102 gnd.t285 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X237 CSoutput.t226 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X238 a_n7636_8799.t1 plus.t16 a_n3827_n3924.t10 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X239 gnd.t64 gnd.t62 minus.t2 gnd.t63 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X240 commonsourceibias.t17 commonsourceibias.t16 gnd.t284 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X241 a_n3827_n3924.t34 minus.t19 a_n1996_n452.t10 gnd.t161 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X242 gnd.t61 gnd.t58 gnd.t60 gnd.t59 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X243 a_n1808_13878.t3 a_n1996_n452.t59 vdd.t90 vdd.t89 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X244 vdd.t291 CSoutput.t227 output.t11 gnd.t349 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X245 CSoutput.t201 commonsourceibias.t103 gnd.t283 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 vdd.t210 a_n7636_8799.t100 CSoutput.t124 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X247 gnd.t282 commonsourceibias.t104 CSoutput.t70 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X248 CSoutput.t228 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X249 CSoutput.t123 a_n7636_8799.t101 vdd.t209 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X250 CSoutput.t122 a_n7636_8799.t102 vdd.t208 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X251 gnd.t271 commonsourceibias.t58 commonsourceibias.t59 gnd.t205 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X252 gnd.t281 commonsourceibias.t105 CSoutput.t54 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 CSoutput.t16 commonsourceibias.t106 gnd.t280 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 gnd.t57 gnd.t54 gnd.t56 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X255 CSoutput.t63 commonsourceibias.t107 gnd.t279 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X256 vdd.t40 vdd.t37 vdd.t39 vdd.t38 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X257 gnd.t278 commonsourceibias.t108 CSoutput.t21 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X258 CSoutput.t25 commonsourceibias.t109 gnd.t277 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X259 minus.t1 gnd.t51 gnd.t53 gnd.t52 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X260 vdd.t36 vdd.t34 vdd.t35 vdd.t23 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X261 a_n3827_n3924.t36 diffpairibias.t26 gnd.t168 gnd.t167 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X262 gnd.t275 commonsourceibias.t110 CSoutput.t39 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X263 a_n1986_8322.t13 a_n1996_n452.t60 a_n7636_8799.t5 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X264 commonsourceibias.t61 commonsourceibias.t60 gnd.t274 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X265 vdd.t33 vdd.t30 vdd.t32 vdd.t31 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X266 vdd.t93 a_n1996_n452.t61 a_n1986_8322.t2 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X267 CSoutput.t121 a_n7636_8799.t103 vdd.t207 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X268 vdd.t205 a_n7636_8799.t104 CSoutput.t120 vdd.t131 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X269 CSoutput.t33 commonsourceibias.t111 gnd.t273 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X270 CSoutput.t119 a_n7636_8799.t105 vdd.t204 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X271 gnd.t272 commonsourceibias.t112 CSoutput.t29 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X272 vdd.t203 a_n7636_8799.t106 CSoutput.t118 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 vdd.t202 a_n7636_8799.t107 CSoutput.t117 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X274 a_n7636_8799.t9 plus.t17 a_n3827_n3924.t9 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X275 CSoutput.t207 commonsourceibias.t113 gnd.t270 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X276 gnd.t269 commonsourceibias.t114 CSoutput.t64 gnd.t250 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X277 gnd.t268 commonsourceibias.t115 CSoutput.t3 gnd.t205 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X278 CSoutput.t12 commonsourceibias.t116 gnd.t267 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X279 commonsourceibias.t57 commonsourceibias.t56 gnd.t266 gnd.t265 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X280 vdd.t29 vdd.t26 vdd.t28 vdd.t27 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X281 a_n3827_n3924.t8 plus.t18 a_n7636_8799.t6 gnd.t137 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X282 vdd.t201 a_n7636_8799.t108 CSoutput.t116 vdd.t145 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X283 CSoutput.t115 a_n7636_8799.t109 vdd.t200 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X284 CSoutput.t114 a_n7636_8799.t110 vdd.t198 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 a_n1808_13878.t12 a_n1996_n452.t28 a_n1996_n452.t29 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X286 CSoutput.t48 commonsourceibias.t117 gnd.t264 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 gnd.t50 gnd.t47 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X288 a_n1986_8322.t12 a_n1996_n452.t62 a_n7636_8799.t25 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X289 diffpairibias.t5 diffpairibias.t4 gnd.t170 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X290 gnd.t263 commonsourceibias.t118 CSoutput.t4 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X291 CSoutput.t202 commonsourceibias.t119 gnd.t261 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 gnd.t259 commonsourceibias.t50 commonsourceibias.t51 gnd.t213 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X293 gnd.t46 gnd.t44 gnd.t45 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X294 output.t10 CSoutput.t229 vdd.t292 gnd.t348 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X295 commonsourceibias.t49 commonsourceibias.t48 gnd.t258 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X296 CSoutput.t113 a_n7636_8799.t111 vdd.t197 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X297 gnd.t257 commonsourceibias.t120 CSoutput.t40 gnd.t250 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X298 CSoutput.t112 a_n7636_8799.t112 vdd.t195 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X299 a_n3827_n3924.t48 diffpairibias.t27 gnd.t369 gnd.t368 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X300 vdd.t194 a_n7636_8799.t113 CSoutput.t111 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 gnd.t256 commonsourceibias.t121 CSoutput.t49 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X302 vdd.t193 a_n7636_8799.t114 CSoutput.t110 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X303 a_n1986_8322.t1 a_n1996_n452.t63 vdd.t128 vdd.t127 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X304 gnd.t254 commonsourceibias.t122 CSoutput.t212 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X305 CSoutput.t203 commonsourceibias.t123 gnd.t253 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X306 CSoutput.t109 a_n7636_8799.t115 vdd.t191 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X307 output.t9 CSoutput.t230 vdd.t293 gnd.t347 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X308 gnd.t252 commonsourceibias.t38 commonsourceibias.t39 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X309 commonsourceibias.t37 commonsourceibias.t36 gnd.t245 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X310 vdd.t114 a_n1996_n452.t64 a_n1808_13878.t2 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X311 CSoutput.t108 a_n7636_8799.t116 vdd.t189 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X312 gnd.t251 commonsourceibias.t124 CSoutput.t50 gnd.t250 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X313 CSoutput.t213 commonsourceibias.t125 gnd.t249 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 CSoutput.t107 a_n7636_8799.t117 vdd.t187 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X315 gnd.t43 gnd.t40 gnd.t42 gnd.t41 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X316 CSoutput.t204 commonsourceibias.t126 gnd.t248 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X317 gnd.t246 commonsourceibias.t127 CSoutput.t10 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X318 commonsourceibias.t35 commonsourceibias.t34 gnd.t244 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X319 gnd.t242 commonsourceibias.t128 CSoutput.t214 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 vdd.t186 a_n7636_8799.t118 CSoutput.t106 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X321 vdd.t150 a_n7636_8799.t119 CSoutput.t105 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 vdd.t25 vdd.t22 vdd.t24 vdd.t23 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X323 gnd.t241 commonsourceibias.t62 commonsourceibias.t63 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X324 gnd.t39 gnd.t36 gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X325 minus.t0 gnd.t33 gnd.t35 gnd.t34 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X326 a_n3827_n3924.t31 minus.t20 a_n1996_n452.t7 gnd.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X327 a_n1986_8322.t11 a_n1996_n452.t65 a_n7636_8799.t19 vdd.t111 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X328 vdd.t21 vdd.t19 vdd.t20 vdd.t16 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X329 CSoutput.t104 a_n7636_8799.t120 vdd.t184 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X330 a_n7636_8799.t20 a_n1996_n452.t66 a_n1986_8322.t10 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X331 gnd.t240 commonsourceibias.t129 CSoutput.t65 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X332 vdd.t182 a_n7636_8799.t121 CSoutput.t103 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X333 a_n1808_13878.t1 a_n1996_n452.t67 vdd.t116 vdd.t115 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X334 CSoutput.t5 commonsourceibias.t130 gnd.t238 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X335 gnd.t32 gnd.t29 gnd.t31 gnd.t30 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X336 vdd.t180 a_n7636_8799.t122 CSoutput.t102 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X337 gnd.t237 commonsourceibias.t131 CSoutput.t196 gnd.t213 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X338 a_n1996_n452.t4 minus.t21 a_n3827_n3924.t28 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X339 CSoutput.t101 a_n7636_8799.t123 vdd.t179 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 vdd.t7 CSoutput.t231 output.t8 gnd.t346 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X341 vdd.t8 CSoutput.t232 output.t7 gnd.t345 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X342 gnd.t233 commonsourceibias.t2 commonsourceibias.t3 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X343 CSoutput.t41 commonsourceibias.t132 gnd.t236 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X344 CSoutput.t34 commonsourceibias.t133 gnd.t235 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X345 CSoutput.t13 commonsourceibias.t134 gnd.t234 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X346 gnd.t232 commonsourceibias.t135 CSoutput.t6 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X347 a_n7636_8799.t15 plus.t19 a_n3827_n3924.t7 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X348 CSoutput.t7 commonsourceibias.t136 gnd.t231 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X349 CSoutput.t233 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X350 a_n3827_n3924.t35 minus.t22 a_n1996_n452.t11 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X351 vdd.t177 a_n7636_8799.t124 CSoutput.t100 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X352 CSoutput.t99 a_n7636_8799.t125 vdd.t175 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X353 CSoutput.t98 a_n7636_8799.t126 vdd.t173 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X354 CSoutput.t22 commonsourceibias.t137 gnd.t229 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X355 CSoutput.t215 commonsourceibias.t138 gnd.t227 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X356 gnd.t226 commonsourceibias.t139 CSoutput.t26 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X357 CSoutput.t97 a_n7636_8799.t127 vdd.t172 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X358 CSoutput.t96 a_n7636_8799.t128 vdd.t171 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X359 a_n1808_13878.t11 a_n1996_n452.t18 a_n1996_n452.t19 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X360 a_n3827_n3924.t6 plus.t20 a_n7636_8799.t4 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X361 vdd.t170 a_n7636_8799.t129 CSoutput.t95 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X362 gnd.t225 commonsourceibias.t0 commonsourceibias.t1 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X363 gnd.t223 commonsourceibias.t4 commonsourceibias.t5 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X364 CSoutput.t94 a_n7636_8799.t130 vdd.t169 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X365 a_n3827_n3924.t49 diffpairibias.t28 gnd.t371 gnd.t370 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X366 vdd.t168 a_n7636_8799.t131 CSoutput.t93 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X367 vdd.t167 a_n7636_8799.t132 CSoutput.t92 vdd.t145 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X368 CSoutput.t66 commonsourceibias.t140 gnd.t221 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X369 gnd.t219 commonsourceibias.t141 CSoutput.t197 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X370 CSoutput.t91 a_n7636_8799.t133 vdd.t166 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X371 a_n1996_n452.t25 a_n1996_n452.t24 a_n1808_13878.t10 vdd.t111 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X372 a_n7636_8799.t12 a_n1996_n452.t68 a_n1986_8322.t9 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X373 vdd.t165 a_n7636_8799.t134 CSoutput.t90 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X374 CSoutput.t89 a_n7636_8799.t135 vdd.t164 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X375 CSoutput.t30 commonsourceibias.t142 gnd.t217 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X376 a_n7636_8799.t8 plus.t21 a_n3827_n3924.t5 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X377 vdd.t162 a_n7636_8799.t136 CSoutput.t88 vdd.t131 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X378 gnd.t28 gnd.t25 gnd.t27 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X379 gnd.t215 commonsourceibias.t143 CSoutput.t208 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X380 gnd.t17 gnd.t15 plus.t1 gnd.t16 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X381 gnd.t214 commonsourceibias.t144 CSoutput.t11 gnd.t213 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X382 gnd.t212 commonsourceibias.t145 CSoutput.t71 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X383 diffpairibias.t3 diffpairibias.t2 gnd.t367 gnd.t366 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X384 vdd.t161 a_n7636_8799.t137 CSoutput.t87 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X385 vdd.t18 vdd.t15 vdd.t17 vdd.t16 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X386 CSoutput.t55 commonsourceibias.t146 gnd.t210 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X387 CSoutput.t86 a_n7636_8799.t138 vdd.t159 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X388 output.t6 CSoutput.t234 vdd.t9 gnd.t344 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X389 gnd.t24 gnd.t21 gnd.t23 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X390 vdd.t117 CSoutput.t235 output.t5 gnd.t343 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X391 a_n3827_n3924.t4 plus.t22 a_n7636_8799.t13 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X392 gnd.t20 gnd.t18 plus.t0 gnd.t19 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X393 gnd.t208 commonsourceibias.t147 CSoutput.t17 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X394 gnd.t206 commonsourceibias.t148 CSoutput.t193 gnd.t205 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X395 vdd.t136 a_n7636_8799.t139 CSoutput.t85 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X396 gnd.t14 gnd.t11 gnd.t13 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X397 diffpairibias.t1 diffpairibias.t0 gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X398 CSoutput.t194 commonsourceibias.t149 gnd.t204 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X399 a_n3827_n3924.t3 plus.t23 a_n7636_8799.t14 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X400 CSoutput.t236 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X401 gnd.t202 commonsourceibias.t150 CSoutput.t8 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X402 vdd.t98 a_n1996_n452.t69 a_n1808_13878.t0 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X403 a_n7636_8799.t7 plus.t24 a_n3827_n3924.t2 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X404 CSoutput.t84 a_n7636_8799.t140 vdd.t157 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X405 a_n3827_n3924.t23 minus.t23 a_n1996_n452.t2 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X406 CSoutput.t83 a_n7636_8799.t141 vdd.t134 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X407 vdd.t155 a_n7636_8799.t142 CSoutput.t82 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X408 gnd.t201 commonsourceibias.t151 CSoutput.t56 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X409 vdd.t154 a_n7636_8799.t143 CSoutput.t81 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X410 CSoutput.t80 a_n7636_8799.t144 vdd.t152 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X411 gnd.t199 commonsourceibias.t152 CSoutput.t72 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X412 a_n1996_n452.t5 minus.t24 a_n3827_n3924.t29 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X413 CSoutput.t79 a_n7636_8799.t145 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X414 a_n1986_8322.t8 a_n1996_n452.t70 a_n7636_8799.t24 vdd.t124 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X415 CSoutput.t51 commonsourceibias.t153 gnd.t197 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X416 vdd.t146 a_n7636_8799.t146 CSoutput.t78 vdd.t145 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X417 vdd.t144 a_n7636_8799.t147 CSoutput.t77 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X418 output.t0 outputibias.t11 gnd.t164 gnd.t163 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X419 CSoutput.t76 a_n7636_8799.t148 vdd.t142 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X420 CSoutput.t75 a_n7636_8799.t149 vdd.t140 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X421 vdd.t138 a_n7636_8799.t150 CSoutput.t74 vdd.t137 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X422 gnd.t195 commonsourceibias.t154 CSoutput.t18 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X423 commonsourceibias.t7 commonsourceibias.t6 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X424 gnd.t191 commonsourceibias.t155 CSoutput.t195 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X425 CSoutput.t57 commonsourceibias.t156 gnd.t189 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X426 a_n1986_8322.t0 a_n1996_n452.t71 vdd.t126 vdd.t125 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X427 a_n1808_13878.t9 a_n1996_n452.t22 a_n1996_n452.t23 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X428 vdd.t118 CSoutput.t237 output.t4 gnd.t342 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X429 vdd.t132 a_n7636_8799.t151 CSoutput.t73 vdd.t131 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X430 a_n3827_n3924.t27 diffpairibias.t29 gnd.t143 gnd.t142 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X431 CSoutput.t0 commonsourceibias.t157 gnd.t187 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X432 CSoutput.t9 commonsourceibias.t158 gnd.t185 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X433 a_n1996_n452.t15 a_n1996_n452.t14 a_n1808_13878.t8 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X434 gnd.t183 commonsourceibias.t159 CSoutput.t58 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X435 vdd.t14 vdd.t11 vdd.t13 vdd.t12 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
R0 a_n7636_8799.n222 a_n7636_8799.t60 485.149
R1 a_n7636_8799.n241 a_n7636_8799.t72 485.149
R2 a_n7636_8799.n261 a_n7636_8799.t109 485.149
R3 a_n7636_8799.n161 a_n7636_8799.t132 485.149
R4 a_n7636_8799.n180 a_n7636_8799.t146 485.149
R5 a_n7636_8799.n200 a_n7636_8799.t108 485.149
R6 a_n7636_8799.n54 a_n7636_8799.t82 485.135
R7 a_n7636_8799.n234 a_n7636_8799.t81 464.166
R8 a_n7636_8799.n216 a_n7636_8799.t54 464.166
R9 a_n7636_8799.n233 a_n7636_8799.t130 464.166
R10 a_n7636_8799.n232 a_n7636_8799.t85 464.166
R11 a_n7636_8799.n217 a_n7636_8799.t61 464.166
R12 a_n7636_8799.n231 a_n7636_8799.t136 464.166
R13 a_n7636_8799.n230 a_n7636_8799.t102 464.166
R14 a_n7636_8799.n218 a_n7636_8799.t100 464.166
R15 a_n7636_8799.n229 a_n7636_8799.t35 464.166
R16 a_n7636_8799.n228 a_n7636_8799.t106 464.166
R17 a_n7636_8799.n219 a_n7636_8799.t105 464.166
R18 a_n7636_8799.n227 a_n7636_8799.t37 464.166
R19 a_n7636_8799.n226 a_n7636_8799.t36 464.166
R20 a_n7636_8799.n220 a_n7636_8799.t122 464.166
R21 a_n7636_8799.n225 a_n7636_8799.t56 464.166
R22 a_n7636_8799.n224 a_n7636_8799.t40 464.166
R23 a_n7636_8799.n221 a_n7636_8799.t126 464.166
R24 a_n7636_8799.n223 a_n7636_8799.t84 464.166
R25 a_n7636_8799.n69 a_n7636_8799.t92 485.135
R26 a_n7636_8799.n253 a_n7636_8799.t91 464.166
R27 a_n7636_8799.n235 a_n7636_8799.t69 464.166
R28 a_n7636_8799.n252 a_n7636_8799.t145 464.166
R29 a_n7636_8799.n251 a_n7636_8799.t98 464.166
R30 a_n7636_8799.n236 a_n7636_8799.t71 464.166
R31 a_n7636_8799.n250 a_n7636_8799.t151 464.166
R32 a_n7636_8799.n249 a_n7636_8799.t115 464.166
R33 a_n7636_8799.n237 a_n7636_8799.t114 464.166
R34 a_n7636_8799.n248 a_n7636_8799.t45 464.166
R35 a_n7636_8799.n247 a_n7636_8799.t118 464.166
R36 a_n7636_8799.n238 a_n7636_8799.t117 464.166
R37 a_n7636_8799.n246 a_n7636_8799.t49 464.166
R38 a_n7636_8799.n245 a_n7636_8799.t48 464.166
R39 a_n7636_8799.n239 a_n7636_8799.t139 464.166
R40 a_n7636_8799.n244 a_n7636_8799.t70 464.166
R41 a_n7636_8799.n243 a_n7636_8799.t52 464.166
R42 a_n7636_8799.n240 a_n7636_8799.t140 464.166
R43 a_n7636_8799.n242 a_n7636_8799.t99 464.166
R44 a_n7636_8799.n84 a_n7636_8799.t150 485.135
R45 a_n7636_8799.n273 a_n7636_8799.t47 464.166
R46 a_n7636_8799.n255 a_n7636_8799.t97 464.166
R47 a_n7636_8799.n272 a_n7636_8799.t34 464.166
R48 a_n7636_8799.n271 a_n7636_8799.t121 464.166
R49 a_n7636_8799.n256 a_n7636_8799.t58 464.166
R50 a_n7636_8799.n270 a_n7636_8799.t104 464.166
R51 a_n7636_8799.n269 a_n7636_8799.t39 464.166
R52 a_n7636_8799.n257 a_n7636_8799.t64 464.166
R53 a_n7636_8799.n268 a_n7636_8799.t144 464.166
R54 a_n7636_8799.n267 a_n7636_8799.t113 464.166
R55 a_n7636_8799.n258 a_n7636_8799.t138 464.166
R56 a_n7636_8799.n266 a_n7636_8799.t95 464.166
R57 a_n7636_8799.n265 a_n7636_8799.t116 464.166
R58 a_n7636_8799.n259 a_n7636_8799.t51 464.166
R59 a_n7636_8799.n264 a_n7636_8799.t135 464.166
R60 a_n7636_8799.n263 a_n7636_8799.t76 464.166
R61 a_n7636_8799.n260 a_n7636_8799.t127 464.166
R62 a_n7636_8799.n262 a_n7636_8799.t63 464.166
R63 a_n7636_8799.n162 a_n7636_8799.t133 464.166
R64 a_n7636_8799.n163 a_n7636_8799.t83 464.166
R65 a_n7636_8799.n164 a_n7636_8799.t112 464.166
R66 a_n7636_8799.n165 a_n7636_8799.t129 464.166
R67 a_n7636_8799.n160 a_n7636_8799.t79 464.166
R68 a_n7636_8799.n166 a_n7636_8799.t80 464.166
R69 a_n7636_8799.n167 a_n7636_8799.t110 464.166
R70 a_n7636_8799.n168 a_n7636_8799.t67 464.166
R71 a_n7636_8799.n169 a_n7636_8799.t68 464.166
R72 a_n7636_8799.n159 a_n7636_8799.t107 464.166
R73 a_n7636_8799.n170 a_n7636_8799.t32 464.166
R74 a_n7636_8799.n158 a_n7636_8799.t65 464.166
R75 a_n7636_8799.n171 a_n7636_8799.t88 464.166
R76 a_n7636_8799.n172 a_n7636_8799.t131 464.166
R77 a_n7636_8799.n173 a_n7636_8799.t44 464.166
R78 a_n7636_8799.n174 a_n7636_8799.t62 464.166
R79 a_n7636_8799.n157 a_n7636_8799.t128 464.166
R80 a_n7636_8799.n175 a_n7636_8799.t41 464.166
R81 a_n7636_8799.n181 a_n7636_8799.t149 464.166
R82 a_n7636_8799.n182 a_n7636_8799.t93 464.166
R83 a_n7636_8799.n183 a_n7636_8799.t125 464.166
R84 a_n7636_8799.n184 a_n7636_8799.t143 464.166
R85 a_n7636_8799.n179 a_n7636_8799.t89 464.166
R86 a_n7636_8799.n185 a_n7636_8799.t90 464.166
R87 a_n7636_8799.n186 a_n7636_8799.t123 464.166
R88 a_n7636_8799.n187 a_n7636_8799.t77 464.166
R89 a_n7636_8799.n188 a_n7636_8799.t78 464.166
R90 a_n7636_8799.n178 a_n7636_8799.t119 464.166
R91 a_n7636_8799.n189 a_n7636_8799.t43 464.166
R92 a_n7636_8799.n177 a_n7636_8799.t74 464.166
R93 a_n7636_8799.n190 a_n7636_8799.t101 464.166
R94 a_n7636_8799.n191 a_n7636_8799.t147 464.166
R95 a_n7636_8799.n192 a_n7636_8799.t59 464.166
R96 a_n7636_8799.n193 a_n7636_8799.t73 464.166
R97 a_n7636_8799.n176 a_n7636_8799.t141 464.166
R98 a_n7636_8799.n194 a_n7636_8799.t53 464.166
R99 a_n7636_8799.n201 a_n7636_8799.t86 464.166
R100 a_n7636_8799.n202 a_n7636_8799.t124 464.166
R101 a_n7636_8799.n203 a_n7636_8799.t75 464.166
R102 a_n7636_8799.n204 a_n7636_8799.t134 464.166
R103 a_n7636_8799.n199 a_n7636_8799.t50 464.166
R104 a_n7636_8799.n205 a_n7636_8799.t33 464.166
R105 a_n7636_8799.n206 a_n7636_8799.t94 464.166
R106 a_n7636_8799.n207 a_n7636_8799.t137 464.166
R107 a_n7636_8799.n208 a_n7636_8799.t111 464.166
R108 a_n7636_8799.n198 a_n7636_8799.t142 464.166
R109 a_n7636_8799.n209 a_n7636_8799.t87 464.166
R110 a_n7636_8799.n197 a_n7636_8799.t38 464.166
R111 a_n7636_8799.n210 a_n7636_8799.t103 464.166
R112 a_n7636_8799.n211 a_n7636_8799.t57 464.166
R113 a_n7636_8799.n212 a_n7636_8799.t120 464.166
R114 a_n7636_8799.n213 a_n7636_8799.t66 464.166
R115 a_n7636_8799.n196 a_n7636_8799.t96 464.166
R116 a_n7636_8799.n214 a_n7636_8799.t46 464.166
R117 a_n7636_8799.n45 a_n7636_8799.n68 71.7212
R118 a_n7636_8799.n68 a_n7636_8799.n221 17.8606
R119 a_n7636_8799.n67 a_n7636_8799.n45 76.9909
R120 a_n7636_8799.n224 a_n7636_8799.n67 7.32118
R121 a_n7636_8799.n66 a_n7636_8799.n44 78.3454
R122 a_n7636_8799.n44 a_n7636_8799.n65 72.8951
R123 a_n7636_8799.n64 a_n7636_8799.n46 70.1674
R124 a_n7636_8799.n227 a_n7636_8799.n64 20.9683
R125 a_n7636_8799.n46 a_n7636_8799.n63 72.3034
R126 a_n7636_8799.n63 a_n7636_8799.n219 16.6962
R127 a_n7636_8799.n62 a_n7636_8799.n47 77.6622
R128 a_n7636_8799.n228 a_n7636_8799.n62 5.97853
R129 a_n7636_8799.n61 a_n7636_8799.n47 77.6622
R130 a_n7636_8799.n48 a_n7636_8799.n60 72.3034
R131 a_n7636_8799.n59 a_n7636_8799.n48 70.1674
R132 a_n7636_8799.n231 a_n7636_8799.n59 20.9683
R133 a_n7636_8799.n50 a_n7636_8799.n58 72.8951
R134 a_n7636_8799.n58 a_n7636_8799.n217 15.5127
R135 a_n7636_8799.n57 a_n7636_8799.n50 78.3454
R136 a_n7636_8799.n232 a_n7636_8799.n57 4.61226
R137 a_n7636_8799.n56 a_n7636_8799.n49 76.9909
R138 a_n7636_8799.n49 a_n7636_8799.n55 71.7212
R139 a_n7636_8799.n234 a_n7636_8799.n54 20.9683
R140 a_n7636_8799.n51 a_n7636_8799.n54 70.1674
R141 a_n7636_8799.n37 a_n7636_8799.n83 71.7212
R142 a_n7636_8799.n83 a_n7636_8799.n240 17.8606
R143 a_n7636_8799.n82 a_n7636_8799.n37 76.9909
R144 a_n7636_8799.n243 a_n7636_8799.n82 7.32118
R145 a_n7636_8799.n81 a_n7636_8799.n36 78.3454
R146 a_n7636_8799.n36 a_n7636_8799.n80 72.8951
R147 a_n7636_8799.n79 a_n7636_8799.n38 70.1674
R148 a_n7636_8799.n246 a_n7636_8799.n79 20.9683
R149 a_n7636_8799.n38 a_n7636_8799.n78 72.3034
R150 a_n7636_8799.n78 a_n7636_8799.n238 16.6962
R151 a_n7636_8799.n77 a_n7636_8799.n39 77.6622
R152 a_n7636_8799.n247 a_n7636_8799.n77 5.97853
R153 a_n7636_8799.n76 a_n7636_8799.n39 77.6622
R154 a_n7636_8799.n40 a_n7636_8799.n75 72.3034
R155 a_n7636_8799.n74 a_n7636_8799.n40 70.1674
R156 a_n7636_8799.n250 a_n7636_8799.n74 20.9683
R157 a_n7636_8799.n42 a_n7636_8799.n73 72.8951
R158 a_n7636_8799.n73 a_n7636_8799.n236 15.5127
R159 a_n7636_8799.n72 a_n7636_8799.n42 78.3454
R160 a_n7636_8799.n251 a_n7636_8799.n72 4.61226
R161 a_n7636_8799.n71 a_n7636_8799.n41 76.9909
R162 a_n7636_8799.n41 a_n7636_8799.n70 71.7212
R163 a_n7636_8799.n253 a_n7636_8799.n69 20.9683
R164 a_n7636_8799.n43 a_n7636_8799.n69 70.1674
R165 a_n7636_8799.n29 a_n7636_8799.n98 71.7212
R166 a_n7636_8799.n98 a_n7636_8799.n260 17.8606
R167 a_n7636_8799.n97 a_n7636_8799.n29 76.9909
R168 a_n7636_8799.n263 a_n7636_8799.n97 7.32118
R169 a_n7636_8799.n96 a_n7636_8799.n28 78.3454
R170 a_n7636_8799.n28 a_n7636_8799.n95 72.8951
R171 a_n7636_8799.n94 a_n7636_8799.n30 70.1674
R172 a_n7636_8799.n266 a_n7636_8799.n94 20.9683
R173 a_n7636_8799.n30 a_n7636_8799.n93 72.3034
R174 a_n7636_8799.n93 a_n7636_8799.n258 16.6962
R175 a_n7636_8799.n92 a_n7636_8799.n31 77.6622
R176 a_n7636_8799.n267 a_n7636_8799.n92 5.97853
R177 a_n7636_8799.n91 a_n7636_8799.n31 77.6622
R178 a_n7636_8799.n32 a_n7636_8799.n90 72.3034
R179 a_n7636_8799.n89 a_n7636_8799.n32 70.1674
R180 a_n7636_8799.n270 a_n7636_8799.n89 20.9683
R181 a_n7636_8799.n34 a_n7636_8799.n88 72.8951
R182 a_n7636_8799.n88 a_n7636_8799.n256 15.5127
R183 a_n7636_8799.n87 a_n7636_8799.n34 78.3454
R184 a_n7636_8799.n271 a_n7636_8799.n87 4.61226
R185 a_n7636_8799.n86 a_n7636_8799.n33 76.9909
R186 a_n7636_8799.n33 a_n7636_8799.n85 71.7212
R187 a_n7636_8799.n273 a_n7636_8799.n84 20.9683
R188 a_n7636_8799.n35 a_n7636_8799.n84 70.1674
R189 a_n7636_8799.n21 a_n7636_8799.n113 70.1674
R190 a_n7636_8799.n175 a_n7636_8799.n113 20.9683
R191 a_n7636_8799.n112 a_n7636_8799.n21 71.7212
R192 a_n7636_8799.n112 a_n7636_8799.n157 17.8606
R193 a_n7636_8799.n20 a_n7636_8799.n111 76.9909
R194 a_n7636_8799.n174 a_n7636_8799.n111 7.32118
R195 a_n7636_8799.n110 a_n7636_8799.n20 78.3454
R196 a_n7636_8799.n22 a_n7636_8799.n109 72.8951
R197 a_n7636_8799.n108 a_n7636_8799.n22 70.1674
R198 a_n7636_8799.n108 a_n7636_8799.n158 20.9683
R199 a_n7636_8799.n23 a_n7636_8799.n107 72.3034
R200 a_n7636_8799.n170 a_n7636_8799.n107 16.6962
R201 a_n7636_8799.n106 a_n7636_8799.n23 77.6622
R202 a_n7636_8799.n106 a_n7636_8799.n159 5.97853
R203 a_n7636_8799.n24 a_n7636_8799.n105 77.6622
R204 a_n7636_8799.n104 a_n7636_8799.n24 72.3034
R205 a_n7636_8799.n25 a_n7636_8799.n103 70.1674
R206 a_n7636_8799.n166 a_n7636_8799.n103 20.9683
R207 a_n7636_8799.n102 a_n7636_8799.n25 72.8951
R208 a_n7636_8799.n102 a_n7636_8799.n160 15.5127
R209 a_n7636_8799.n26 a_n7636_8799.n101 78.3454
R210 a_n7636_8799.n165 a_n7636_8799.n101 4.61226
R211 a_n7636_8799.n100 a_n7636_8799.n26 76.9909
R212 a_n7636_8799.n99 a_n7636_8799.n163 17.8606
R213 a_n7636_8799.n99 a_n7636_8799.n27 71.7212
R214 a_n7636_8799.n13 a_n7636_8799.n128 70.1674
R215 a_n7636_8799.n194 a_n7636_8799.n128 20.9683
R216 a_n7636_8799.n127 a_n7636_8799.n13 71.7212
R217 a_n7636_8799.n127 a_n7636_8799.n176 17.8606
R218 a_n7636_8799.n12 a_n7636_8799.n126 76.9909
R219 a_n7636_8799.n193 a_n7636_8799.n126 7.32118
R220 a_n7636_8799.n125 a_n7636_8799.n12 78.3454
R221 a_n7636_8799.n14 a_n7636_8799.n124 72.8951
R222 a_n7636_8799.n123 a_n7636_8799.n14 70.1674
R223 a_n7636_8799.n123 a_n7636_8799.n177 20.9683
R224 a_n7636_8799.n15 a_n7636_8799.n122 72.3034
R225 a_n7636_8799.n189 a_n7636_8799.n122 16.6962
R226 a_n7636_8799.n121 a_n7636_8799.n15 77.6622
R227 a_n7636_8799.n121 a_n7636_8799.n178 5.97853
R228 a_n7636_8799.n16 a_n7636_8799.n120 77.6622
R229 a_n7636_8799.n119 a_n7636_8799.n16 72.3034
R230 a_n7636_8799.n17 a_n7636_8799.n118 70.1674
R231 a_n7636_8799.n185 a_n7636_8799.n118 20.9683
R232 a_n7636_8799.n117 a_n7636_8799.n17 72.8951
R233 a_n7636_8799.n117 a_n7636_8799.n179 15.5127
R234 a_n7636_8799.n18 a_n7636_8799.n116 78.3454
R235 a_n7636_8799.n184 a_n7636_8799.n116 4.61226
R236 a_n7636_8799.n115 a_n7636_8799.n18 76.9909
R237 a_n7636_8799.n114 a_n7636_8799.n182 17.8606
R238 a_n7636_8799.n114 a_n7636_8799.n19 71.7212
R239 a_n7636_8799.n5 a_n7636_8799.n143 70.1674
R240 a_n7636_8799.n214 a_n7636_8799.n143 20.9683
R241 a_n7636_8799.n142 a_n7636_8799.n5 71.7212
R242 a_n7636_8799.n142 a_n7636_8799.n196 17.8606
R243 a_n7636_8799.n4 a_n7636_8799.n141 76.9909
R244 a_n7636_8799.n213 a_n7636_8799.n141 7.32118
R245 a_n7636_8799.n140 a_n7636_8799.n4 78.3454
R246 a_n7636_8799.n6 a_n7636_8799.n139 72.8951
R247 a_n7636_8799.n138 a_n7636_8799.n6 70.1674
R248 a_n7636_8799.n138 a_n7636_8799.n197 20.9683
R249 a_n7636_8799.n7 a_n7636_8799.n137 72.3034
R250 a_n7636_8799.n209 a_n7636_8799.n137 16.6962
R251 a_n7636_8799.n136 a_n7636_8799.n7 77.6622
R252 a_n7636_8799.n136 a_n7636_8799.n198 5.97853
R253 a_n7636_8799.n8 a_n7636_8799.n135 77.6622
R254 a_n7636_8799.n134 a_n7636_8799.n8 72.3034
R255 a_n7636_8799.n9 a_n7636_8799.n133 70.1674
R256 a_n7636_8799.n205 a_n7636_8799.n133 20.9683
R257 a_n7636_8799.n132 a_n7636_8799.n9 72.8951
R258 a_n7636_8799.n132 a_n7636_8799.n199 15.5127
R259 a_n7636_8799.n10 a_n7636_8799.n131 78.3454
R260 a_n7636_8799.n204 a_n7636_8799.n131 4.61226
R261 a_n7636_8799.n130 a_n7636_8799.n10 76.9909
R262 a_n7636_8799.n129 a_n7636_8799.n202 17.8606
R263 a_n7636_8799.n129 a_n7636_8799.n11 71.7212
R264 a_n7636_8799.n52 a_n7636_8799.n144 98.9633
R265 a_n7636_8799.n280 a_n7636_8799.n53 98.9632
R266 a_n7636_8799.n53 a_n7636_8799.n279 98.6055
R267 a_n7636_8799.n53 a_n7636_8799.n278 98.6055
R268 a_n7636_8799.n52 a_n7636_8799.n146 98.6055
R269 a_n7636_8799.n52 a_n7636_8799.n145 98.6055
R270 a_n7636_8799.n3 a_n7636_8799.n147 81.3764
R271 a_n7636_8799.n1 a_n7636_8799.n153 81.3764
R272 a_n7636_8799.n0 a_n7636_8799.n150 81.3764
R273 a_n7636_8799.n2 a_n7636_8799.n155 80.9324
R274 a_n7636_8799.n2 a_n7636_8799.n156 80.9324
R275 a_n7636_8799.n3 a_n7636_8799.n149 80.9324
R276 a_n7636_8799.n3 a_n7636_8799.n148 80.9324
R277 a_n7636_8799.n1 a_n7636_8799.n154 80.9324
R278 a_n7636_8799.n1 a_n7636_8799.n152 80.9324
R279 a_n7636_8799.n0 a_n7636_8799.n151 80.9324
R280 a_n7636_8799.n45 a_n7636_8799.n222 70.4033
R281 a_n7636_8799.n37 a_n7636_8799.n241 70.4033
R282 a_n7636_8799.n29 a_n7636_8799.n261 70.4033
R283 a_n7636_8799.n161 a_n7636_8799.n27 70.4033
R284 a_n7636_8799.n180 a_n7636_8799.n19 70.4033
R285 a_n7636_8799.n200 a_n7636_8799.n11 70.4033
R286 a_n7636_8799.n233 a_n7636_8799.n232 48.2005
R287 a_n7636_8799.n59 a_n7636_8799.n230 20.9683
R288 a_n7636_8799.n229 a_n7636_8799.n228 48.2005
R289 a_n7636_8799.n64 a_n7636_8799.n226 20.9683
R290 a_n7636_8799.n225 a_n7636_8799.n224 48.2005
R291 a_n7636_8799.n252 a_n7636_8799.n251 48.2005
R292 a_n7636_8799.n74 a_n7636_8799.n249 20.9683
R293 a_n7636_8799.n248 a_n7636_8799.n247 48.2005
R294 a_n7636_8799.n79 a_n7636_8799.n245 20.9683
R295 a_n7636_8799.n244 a_n7636_8799.n243 48.2005
R296 a_n7636_8799.n272 a_n7636_8799.n271 48.2005
R297 a_n7636_8799.n89 a_n7636_8799.n269 20.9683
R298 a_n7636_8799.n268 a_n7636_8799.n267 48.2005
R299 a_n7636_8799.n94 a_n7636_8799.n265 20.9683
R300 a_n7636_8799.n264 a_n7636_8799.n263 48.2005
R301 a_n7636_8799.n165 a_n7636_8799.n164 48.2005
R302 a_n7636_8799.n167 a_n7636_8799.n103 20.9683
R303 a_n7636_8799.n169 a_n7636_8799.n159 48.2005
R304 a_n7636_8799.n171 a_n7636_8799.n108 20.9683
R305 a_n7636_8799.n174 a_n7636_8799.n173 48.2005
R306 a_n7636_8799.t42 a_n7636_8799.n113 485.135
R307 a_n7636_8799.n184 a_n7636_8799.n183 48.2005
R308 a_n7636_8799.n186 a_n7636_8799.n118 20.9683
R309 a_n7636_8799.n188 a_n7636_8799.n178 48.2005
R310 a_n7636_8799.n190 a_n7636_8799.n123 20.9683
R311 a_n7636_8799.n193 a_n7636_8799.n192 48.2005
R312 a_n7636_8799.t55 a_n7636_8799.n128 485.135
R313 a_n7636_8799.n204 a_n7636_8799.n203 48.2005
R314 a_n7636_8799.n206 a_n7636_8799.n133 20.9683
R315 a_n7636_8799.n208 a_n7636_8799.n198 48.2005
R316 a_n7636_8799.n210 a_n7636_8799.n138 20.9683
R317 a_n7636_8799.n213 a_n7636_8799.n212 48.2005
R318 a_n7636_8799.t148 a_n7636_8799.n143 485.135
R319 a_n7636_8799.n55 a_n7636_8799.n216 17.8606
R320 a_n7636_8799.n223 a_n7636_8799.n68 25.894
R321 a_n7636_8799.n70 a_n7636_8799.n235 17.8606
R322 a_n7636_8799.n242 a_n7636_8799.n83 25.894
R323 a_n7636_8799.n85 a_n7636_8799.n255 17.8606
R324 a_n7636_8799.n262 a_n7636_8799.n98 25.894
R325 a_n7636_8799.n175 a_n7636_8799.n112 25.894
R326 a_n7636_8799.n194 a_n7636_8799.n127 25.894
R327 a_n7636_8799.n214 a_n7636_8799.n142 25.894
R328 a_n7636_8799.n66 a_n7636_8799.n220 43.3183
R329 a_n7636_8799.n81 a_n7636_8799.n239 43.3183
R330 a_n7636_8799.n96 a_n7636_8799.n259 43.3183
R331 a_n7636_8799.n172 a_n7636_8799.n110 43.3183
R332 a_n7636_8799.n191 a_n7636_8799.n125 43.3183
R333 a_n7636_8799.n211 a_n7636_8799.n140 43.3183
R334 a_n7636_8799.n60 a_n7636_8799.n218 16.6962
R335 a_n7636_8799.n227 a_n7636_8799.n63 27.6507
R336 a_n7636_8799.n75 a_n7636_8799.n237 16.6962
R337 a_n7636_8799.n246 a_n7636_8799.n78 27.6507
R338 a_n7636_8799.n90 a_n7636_8799.n257 16.6962
R339 a_n7636_8799.n266 a_n7636_8799.n93 27.6507
R340 a_n7636_8799.n168 a_n7636_8799.n104 16.6962
R341 a_n7636_8799.n158 a_n7636_8799.n107 27.6507
R342 a_n7636_8799.n187 a_n7636_8799.n119 16.6962
R343 a_n7636_8799.n177 a_n7636_8799.n122 27.6507
R344 a_n7636_8799.n207 a_n7636_8799.n134 16.6962
R345 a_n7636_8799.n197 a_n7636_8799.n137 27.6507
R346 a_n7636_8799.n61 a_n7636_8799.n218 41.7634
R347 a_n7636_8799.n76 a_n7636_8799.n237 41.7634
R348 a_n7636_8799.n91 a_n7636_8799.n257 41.7634
R349 a_n7636_8799.n105 a_n7636_8799.n168 41.7634
R350 a_n7636_8799.n120 a_n7636_8799.n187 41.7634
R351 a_n7636_8799.n135 a_n7636_8799.n207 41.7634
R352 a_n7636_8799.n231 a_n7636_8799.n58 29.3885
R353 a_n7636_8799.n65 a_n7636_8799.n220 15.5127
R354 a_n7636_8799.n250 a_n7636_8799.n73 29.3885
R355 a_n7636_8799.n80 a_n7636_8799.n239 15.5127
R356 a_n7636_8799.n270 a_n7636_8799.n88 29.3885
R357 a_n7636_8799.n95 a_n7636_8799.n259 15.5127
R358 a_n7636_8799.n166 a_n7636_8799.n102 29.3885
R359 a_n7636_8799.n172 a_n7636_8799.n109 15.5127
R360 a_n7636_8799.n185 a_n7636_8799.n117 29.3885
R361 a_n7636_8799.n191 a_n7636_8799.n124 15.5127
R362 a_n7636_8799.n205 a_n7636_8799.n132 29.3885
R363 a_n7636_8799.n211 a_n7636_8799.n139 15.5127
R364 a_n7636_8799.n56 a_n7636_8799.n216 40.1848
R365 a_n7636_8799.n71 a_n7636_8799.n235 40.1848
R366 a_n7636_8799.n86 a_n7636_8799.n255 40.1848
R367 a_n7636_8799.n163 a_n7636_8799.n100 40.1848
R368 a_n7636_8799.n182 a_n7636_8799.n115 40.1848
R369 a_n7636_8799.n202 a_n7636_8799.n130 40.1848
R370 a_n7636_8799.n2 a_n7636_8799.n1 32.7526
R371 a_n7636_8799.n223 a_n7636_8799.n222 20.9576
R372 a_n7636_8799.n242 a_n7636_8799.n241 20.9576
R373 a_n7636_8799.n262 a_n7636_8799.n261 20.9576
R374 a_n7636_8799.n162 a_n7636_8799.n161 20.9576
R375 a_n7636_8799.n181 a_n7636_8799.n180 20.9576
R376 a_n7636_8799.n201 a_n7636_8799.n200 20.9576
R377 a_n7636_8799.n56 a_n7636_8799.n233 7.32118
R378 a_n7636_8799.n67 a_n7636_8799.n221 40.1848
R379 a_n7636_8799.n71 a_n7636_8799.n252 7.32118
R380 a_n7636_8799.n82 a_n7636_8799.n240 40.1848
R381 a_n7636_8799.n86 a_n7636_8799.n272 7.32118
R382 a_n7636_8799.n97 a_n7636_8799.n260 40.1848
R383 a_n7636_8799.n164 a_n7636_8799.n100 7.32118
R384 a_n7636_8799.n157 a_n7636_8799.n111 40.1848
R385 a_n7636_8799.n183 a_n7636_8799.n115 7.32118
R386 a_n7636_8799.n176 a_n7636_8799.n126 40.1848
R387 a_n7636_8799.n203 a_n7636_8799.n130 7.32118
R388 a_n7636_8799.n196 a_n7636_8799.n141 40.1848
R389 a_n7636_8799.n226 a_n7636_8799.n65 29.3885
R390 a_n7636_8799.n245 a_n7636_8799.n80 29.3885
R391 a_n7636_8799.n265 a_n7636_8799.n95 29.3885
R392 a_n7636_8799.n109 a_n7636_8799.n171 29.3885
R393 a_n7636_8799.n124 a_n7636_8799.n190 29.3885
R394 a_n7636_8799.n139 a_n7636_8799.n210 29.3885
R395 a_n7636_8799.n61 a_n7636_8799.n229 5.97853
R396 a_n7636_8799.n62 a_n7636_8799.n219 41.7634
R397 a_n7636_8799.n76 a_n7636_8799.n248 5.97853
R398 a_n7636_8799.n77 a_n7636_8799.n238 41.7634
R399 a_n7636_8799.n91 a_n7636_8799.n268 5.97853
R400 a_n7636_8799.n92 a_n7636_8799.n258 41.7634
R401 a_n7636_8799.n169 a_n7636_8799.n105 5.97853
R402 a_n7636_8799.n170 a_n7636_8799.n106 41.7634
R403 a_n7636_8799.n188 a_n7636_8799.n120 5.97853
R404 a_n7636_8799.n189 a_n7636_8799.n121 41.7634
R405 a_n7636_8799.n208 a_n7636_8799.n135 5.97853
R406 a_n7636_8799.n209 a_n7636_8799.n136 41.7634
R407 a_n7636_8799.n276 a_n7636_8799.n3 12.3339
R408 a_n7636_8799.n277 a_n7636_8799.n276 11.4887
R409 a_n7636_8799.n230 a_n7636_8799.n60 27.6507
R410 a_n7636_8799.n249 a_n7636_8799.n75 27.6507
R411 a_n7636_8799.n269 a_n7636_8799.n90 27.6507
R412 a_n7636_8799.n167 a_n7636_8799.n104 27.6507
R413 a_n7636_8799.n186 a_n7636_8799.n119 27.6507
R414 a_n7636_8799.n206 a_n7636_8799.n134 27.6507
R415 a_n7636_8799.n57 a_n7636_8799.n217 43.3183
R416 a_n7636_8799.n66 a_n7636_8799.n225 4.61226
R417 a_n7636_8799.n72 a_n7636_8799.n236 43.3183
R418 a_n7636_8799.n81 a_n7636_8799.n244 4.61226
R419 a_n7636_8799.n87 a_n7636_8799.n256 43.3183
R420 a_n7636_8799.n96 a_n7636_8799.n264 4.61226
R421 a_n7636_8799.n160 a_n7636_8799.n101 43.3183
R422 a_n7636_8799.n173 a_n7636_8799.n110 4.61226
R423 a_n7636_8799.n179 a_n7636_8799.n116 43.3183
R424 a_n7636_8799.n192 a_n7636_8799.n125 4.61226
R425 a_n7636_8799.n199 a_n7636_8799.n131 43.3183
R426 a_n7636_8799.n53 a_n7636_8799.n277 31.0713
R427 a_n7636_8799.n212 a_n7636_8799.n140 4.61226
R428 a_n7636_8799.n254 a_n7636_8799.n51 9.04406
R429 a_n7636_8799.n195 a_n7636_8799.n21 9.04406
R430 a_n7636_8799.n234 a_n7636_8799.n55 25.894
R431 a_n7636_8799.n253 a_n7636_8799.n70 25.894
R432 a_n7636_8799.n273 a_n7636_8799.n85 25.894
R433 a_n7636_8799.n99 a_n7636_8799.n162 25.894
R434 a_n7636_8799.n114 a_n7636_8799.n181 25.894
R435 a_n7636_8799.n129 a_n7636_8799.n201 25.894
R436 a_n7636_8799.n277 a_n7636_8799.n52 18.0938
R437 a_n7636_8799.n275 a_n7636_8799.n215 6.86985
R438 a_n7636_8799.n275 a_n7636_8799.n274 6.51296
R439 a_n7636_8799.n254 a_n7636_8799.n43 4.93611
R440 a_n7636_8799.n274 a_n7636_8799.n35 4.93611
R441 a_n7636_8799.n195 a_n7636_8799.n13 4.93611
R442 a_n7636_8799.n215 a_n7636_8799.n5 4.93611
R443 a_n7636_8799.n274 a_n7636_8799.n254 4.10845
R444 a_n7636_8799.n215 a_n7636_8799.n195 4.10845
R445 a_n7636_8799.n279 a_n7636_8799.t31 3.61217
R446 a_n7636_8799.n279 a_n7636_8799.t28 3.61217
R447 a_n7636_8799.n278 a_n7636_8799.t19 3.61217
R448 a_n7636_8799.n278 a_n7636_8799.t20 3.61217
R449 a_n7636_8799.n146 a_n7636_8799.t25 3.61217
R450 a_n7636_8799.n146 a_n7636_8799.t12 3.61217
R451 a_n7636_8799.n145 a_n7636_8799.t27 3.61217
R452 a_n7636_8799.n145 a_n7636_8799.t30 3.61217
R453 a_n7636_8799.n144 a_n7636_8799.t24 3.61217
R454 a_n7636_8799.n144 a_n7636_8799.t22 3.61217
R455 a_n7636_8799.t5 a_n7636_8799.n280 3.61217
R456 a_n7636_8799.n280 a_n7636_8799.t17 3.61217
R457 a_n7636_8799.n276 a_n7636_8799.n275 3.4105
R458 a_n7636_8799.n155 a_n7636_8799.t3 2.82907
R459 a_n7636_8799.n155 a_n7636_8799.t7 2.82907
R460 a_n7636_8799.n156 a_n7636_8799.t0 2.82907
R461 a_n7636_8799.n156 a_n7636_8799.t29 2.82907
R462 a_n7636_8799.n149 a_n7636_8799.t14 2.82907
R463 a_n7636_8799.n149 a_n7636_8799.t10 2.82907
R464 a_n7636_8799.n148 a_n7636_8799.t13 2.82907
R465 a_n7636_8799.n148 a_n7636_8799.t8 2.82907
R466 a_n7636_8799.n147 a_n7636_8799.t6 2.82907
R467 a_n7636_8799.n147 a_n7636_8799.t9 2.82907
R468 a_n7636_8799.n153 a_n7636_8799.t16 2.82907
R469 a_n7636_8799.n153 a_n7636_8799.t21 2.82907
R470 a_n7636_8799.n154 a_n7636_8799.t4 2.82907
R471 a_n7636_8799.n154 a_n7636_8799.t1 2.82907
R472 a_n7636_8799.n152 a_n7636_8799.t26 2.82907
R473 a_n7636_8799.n152 a_n7636_8799.t15 2.82907
R474 a_n7636_8799.n151 a_n7636_8799.t11 2.82907
R475 a_n7636_8799.n151 a_n7636_8799.t18 2.82907
R476 a_n7636_8799.n150 a_n7636_8799.t2 2.82907
R477 a_n7636_8799.n150 a_n7636_8799.t23 2.82907
R478 a_n7636_8799.n3 a_n7636_8799.n2 1.3324
R479 a_n7636_8799.n45 a_n7636_8799.n44 1.13686
R480 a_n7636_8799.n37 a_n7636_8799.n36 1.13686
R481 a_n7636_8799.n29 a_n7636_8799.n28 1.13686
R482 a_n7636_8799.n21 a_n7636_8799.n20 1.13686
R483 a_n7636_8799.n13 a_n7636_8799.n12 1.13686
R484 a_n7636_8799.n5 a_n7636_8799.n4 1.13686
R485 a_n7636_8799.n1 a_n7636_8799.n0 0.888431
R486 a_n7636_8799.n50 a_n7636_8799.n49 0.758076
R487 a_n7636_8799.n50 a_n7636_8799.n48 0.758076
R488 a_n7636_8799.n48 a_n7636_8799.n47 0.758076
R489 a_n7636_8799.n47 a_n7636_8799.n46 0.758076
R490 a_n7636_8799.n44 a_n7636_8799.n46 0.758076
R491 a_n7636_8799.n42 a_n7636_8799.n41 0.758076
R492 a_n7636_8799.n42 a_n7636_8799.n40 0.758076
R493 a_n7636_8799.n40 a_n7636_8799.n39 0.758076
R494 a_n7636_8799.n39 a_n7636_8799.n38 0.758076
R495 a_n7636_8799.n36 a_n7636_8799.n38 0.758076
R496 a_n7636_8799.n34 a_n7636_8799.n33 0.758076
R497 a_n7636_8799.n34 a_n7636_8799.n32 0.758076
R498 a_n7636_8799.n32 a_n7636_8799.n31 0.758076
R499 a_n7636_8799.n31 a_n7636_8799.n30 0.758076
R500 a_n7636_8799.n28 a_n7636_8799.n30 0.758076
R501 a_n7636_8799.n25 a_n7636_8799.n26 0.758076
R502 a_n7636_8799.n24 a_n7636_8799.n25 0.758076
R503 a_n7636_8799.n23 a_n7636_8799.n24 0.758076
R504 a_n7636_8799.n22 a_n7636_8799.n23 0.758076
R505 a_n7636_8799.n20 a_n7636_8799.n22 0.758076
R506 a_n7636_8799.n17 a_n7636_8799.n18 0.758076
R507 a_n7636_8799.n16 a_n7636_8799.n17 0.758076
R508 a_n7636_8799.n15 a_n7636_8799.n16 0.758076
R509 a_n7636_8799.n14 a_n7636_8799.n15 0.758076
R510 a_n7636_8799.n12 a_n7636_8799.n14 0.758076
R511 a_n7636_8799.n9 a_n7636_8799.n10 0.758076
R512 a_n7636_8799.n8 a_n7636_8799.n9 0.758076
R513 a_n7636_8799.n7 a_n7636_8799.n8 0.758076
R514 a_n7636_8799.n6 a_n7636_8799.n7 0.758076
R515 a_n7636_8799.n4 a_n7636_8799.n6 0.758076
R516 a_n7636_8799.n10 a_n7636_8799.n11 0.568682
R517 a_n7636_8799.n18 a_n7636_8799.n19 0.568682
R518 a_n7636_8799.n26 a_n7636_8799.n27 0.568682
R519 a_n7636_8799.n33 a_n7636_8799.n35 0.568682
R520 a_n7636_8799.n41 a_n7636_8799.n43 0.568682
R521 a_n7636_8799.n49 a_n7636_8799.n51 0.568682
R522 vdd.n327 vdd.n291 756.745
R523 vdd.n268 vdd.n232 756.745
R524 vdd.n225 vdd.n189 756.745
R525 vdd.n166 vdd.n130 756.745
R526 vdd.n124 vdd.n88 756.745
R527 vdd.n65 vdd.n29 756.745
R528 vdd.n1746 vdd.n1710 756.745
R529 vdd.n1805 vdd.n1769 756.745
R530 vdd.n1644 vdd.n1608 756.745
R531 vdd.n1703 vdd.n1667 756.745
R532 vdd.n1543 vdd.n1507 756.745
R533 vdd.n1602 vdd.n1566 756.745
R534 vdd.n2177 vdd.t65 640.208
R535 vdd.n965 vdd.t50 640.208
R536 vdd.n2151 vdd.t11 640.208
R537 vdd.n957 vdd.t75 640.208
R538 vdd.n2922 vdd.t26 640.208
R539 vdd.n2642 vdd.t72 640.208
R540 vdd.n832 vdd.t54 640.208
R541 vdd.n2639 vdd.t58 640.208
R542 vdd.n799 vdd.t62 640.208
R543 vdd.n1027 vdd.t68 640.208
R544 vdd.n1317 vdd.t41 592.009
R545 vdd.n1355 vdd.t30 592.009
R546 vdd.n1251 vdd.t44 592.009
R547 vdd.n2333 vdd.t22 592.009
R548 vdd.n1970 vdd.t34 592.009
R549 vdd.n1930 vdd.t47 592.009
R550 vdd.n426 vdd.t37 592.009
R551 vdd.n440 vdd.t78 592.009
R552 vdd.n452 vdd.t84 592.009
R553 vdd.n768 vdd.t15 592.009
R554 vdd.n3184 vdd.t19 592.009
R555 vdd.n688 vdd.t81 592.009
R556 vdd.n328 vdd.n327 585
R557 vdd.n326 vdd.n293 585
R558 vdd.n325 vdd.n324 585
R559 vdd.n296 vdd.n294 585
R560 vdd.n319 vdd.n318 585
R561 vdd.n317 vdd.n316 585
R562 vdd.n300 vdd.n299 585
R563 vdd.n311 vdd.n310 585
R564 vdd.n309 vdd.n308 585
R565 vdd.n304 vdd.n303 585
R566 vdd.n269 vdd.n268 585
R567 vdd.n267 vdd.n234 585
R568 vdd.n266 vdd.n265 585
R569 vdd.n237 vdd.n235 585
R570 vdd.n260 vdd.n259 585
R571 vdd.n258 vdd.n257 585
R572 vdd.n241 vdd.n240 585
R573 vdd.n252 vdd.n251 585
R574 vdd.n250 vdd.n249 585
R575 vdd.n245 vdd.n244 585
R576 vdd.n226 vdd.n225 585
R577 vdd.n224 vdd.n191 585
R578 vdd.n223 vdd.n222 585
R579 vdd.n194 vdd.n192 585
R580 vdd.n217 vdd.n216 585
R581 vdd.n215 vdd.n214 585
R582 vdd.n198 vdd.n197 585
R583 vdd.n209 vdd.n208 585
R584 vdd.n207 vdd.n206 585
R585 vdd.n202 vdd.n201 585
R586 vdd.n167 vdd.n166 585
R587 vdd.n165 vdd.n132 585
R588 vdd.n164 vdd.n163 585
R589 vdd.n135 vdd.n133 585
R590 vdd.n158 vdd.n157 585
R591 vdd.n156 vdd.n155 585
R592 vdd.n139 vdd.n138 585
R593 vdd.n150 vdd.n149 585
R594 vdd.n148 vdd.n147 585
R595 vdd.n143 vdd.n142 585
R596 vdd.n125 vdd.n124 585
R597 vdd.n123 vdd.n90 585
R598 vdd.n122 vdd.n121 585
R599 vdd.n93 vdd.n91 585
R600 vdd.n116 vdd.n115 585
R601 vdd.n114 vdd.n113 585
R602 vdd.n97 vdd.n96 585
R603 vdd.n108 vdd.n107 585
R604 vdd.n106 vdd.n105 585
R605 vdd.n101 vdd.n100 585
R606 vdd.n66 vdd.n65 585
R607 vdd.n64 vdd.n31 585
R608 vdd.n63 vdd.n62 585
R609 vdd.n34 vdd.n32 585
R610 vdd.n57 vdd.n56 585
R611 vdd.n55 vdd.n54 585
R612 vdd.n38 vdd.n37 585
R613 vdd.n49 vdd.n48 585
R614 vdd.n47 vdd.n46 585
R615 vdd.n42 vdd.n41 585
R616 vdd.n1747 vdd.n1746 585
R617 vdd.n1745 vdd.n1712 585
R618 vdd.n1744 vdd.n1743 585
R619 vdd.n1715 vdd.n1713 585
R620 vdd.n1738 vdd.n1737 585
R621 vdd.n1736 vdd.n1735 585
R622 vdd.n1719 vdd.n1718 585
R623 vdd.n1730 vdd.n1729 585
R624 vdd.n1728 vdd.n1727 585
R625 vdd.n1723 vdd.n1722 585
R626 vdd.n1806 vdd.n1805 585
R627 vdd.n1804 vdd.n1771 585
R628 vdd.n1803 vdd.n1802 585
R629 vdd.n1774 vdd.n1772 585
R630 vdd.n1797 vdd.n1796 585
R631 vdd.n1795 vdd.n1794 585
R632 vdd.n1778 vdd.n1777 585
R633 vdd.n1789 vdd.n1788 585
R634 vdd.n1787 vdd.n1786 585
R635 vdd.n1782 vdd.n1781 585
R636 vdd.n1645 vdd.n1644 585
R637 vdd.n1643 vdd.n1610 585
R638 vdd.n1642 vdd.n1641 585
R639 vdd.n1613 vdd.n1611 585
R640 vdd.n1636 vdd.n1635 585
R641 vdd.n1634 vdd.n1633 585
R642 vdd.n1617 vdd.n1616 585
R643 vdd.n1628 vdd.n1627 585
R644 vdd.n1626 vdd.n1625 585
R645 vdd.n1621 vdd.n1620 585
R646 vdd.n1704 vdd.n1703 585
R647 vdd.n1702 vdd.n1669 585
R648 vdd.n1701 vdd.n1700 585
R649 vdd.n1672 vdd.n1670 585
R650 vdd.n1695 vdd.n1694 585
R651 vdd.n1693 vdd.n1692 585
R652 vdd.n1676 vdd.n1675 585
R653 vdd.n1687 vdd.n1686 585
R654 vdd.n1685 vdd.n1684 585
R655 vdd.n1680 vdd.n1679 585
R656 vdd.n1544 vdd.n1543 585
R657 vdd.n1542 vdd.n1509 585
R658 vdd.n1541 vdd.n1540 585
R659 vdd.n1512 vdd.n1510 585
R660 vdd.n1535 vdd.n1534 585
R661 vdd.n1533 vdd.n1532 585
R662 vdd.n1516 vdd.n1515 585
R663 vdd.n1527 vdd.n1526 585
R664 vdd.n1525 vdd.n1524 585
R665 vdd.n1520 vdd.n1519 585
R666 vdd.n1603 vdd.n1602 585
R667 vdd.n1601 vdd.n1568 585
R668 vdd.n1600 vdd.n1599 585
R669 vdd.n1571 vdd.n1569 585
R670 vdd.n1594 vdd.n1593 585
R671 vdd.n1592 vdd.n1591 585
R672 vdd.n1575 vdd.n1574 585
R673 vdd.n1586 vdd.n1585 585
R674 vdd.n1584 vdd.n1583 585
R675 vdd.n1579 vdd.n1578 585
R676 vdd.n3356 vdd.n392 509.269
R677 vdd.n3352 vdd.n393 509.269
R678 vdd.n3224 vdd.n685 509.269
R679 vdd.n3221 vdd.n684 509.269
R680 vdd.n2328 vdd.n1075 509.269
R681 vdd.n2331 vdd.n2330 509.269
R682 vdd.n1224 vdd.n1188 509.269
R683 vdd.n1420 vdd.n1189 509.269
R684 vdd.n305 vdd.t263 329.043
R685 vdd.n246 vdd.t237 329.043
R686 vdd.n203 vdd.t251 329.043
R687 vdd.n144 vdd.t216 329.043
R688 vdd.n102 vdd.t200 329.043
R689 vdd.n43 vdd.t138 329.043
R690 vdd.n1724 vdd.t280 329.043
R691 vdd.n1783 vdd.t167 329.043
R692 vdd.n1622 vdd.t267 329.043
R693 vdd.n1681 vdd.t146 329.043
R694 vdd.n1521 vdd.t142 329.043
R695 vdd.n1580 vdd.t201 329.043
R696 vdd.n1317 vdd.t43 319.788
R697 vdd.n1355 vdd.t33 319.788
R698 vdd.n1251 vdd.t46 319.788
R699 vdd.n2333 vdd.t24 319.788
R700 vdd.n1970 vdd.t35 319.788
R701 vdd.n1930 vdd.t48 319.788
R702 vdd.n426 vdd.t39 319.788
R703 vdd.n440 vdd.t79 319.788
R704 vdd.n452 vdd.t85 319.788
R705 vdd.n768 vdd.t18 319.788
R706 vdd.n3184 vdd.t21 319.788
R707 vdd.n688 vdd.t83 319.788
R708 vdd.n1318 vdd.t42 303.69
R709 vdd.n1356 vdd.t32 303.69
R710 vdd.n1252 vdd.t45 303.69
R711 vdd.n2334 vdd.t25 303.69
R712 vdd.n1971 vdd.t36 303.69
R713 vdd.n1931 vdd.t49 303.69
R714 vdd.n427 vdd.t40 303.69
R715 vdd.n441 vdd.t80 303.69
R716 vdd.n453 vdd.t86 303.69
R717 vdd.n769 vdd.t17 303.69
R718 vdd.n3185 vdd.t20 303.69
R719 vdd.n689 vdd.t82 303.69
R720 vdd.n2865 vdd.n913 297.074
R721 vdd.n3058 vdd.n809 297.074
R722 vdd.n2995 vdd.n806 297.074
R723 vdd.n2788 vdd.n914 297.074
R724 vdd.n2603 vdd.n954 297.074
R725 vdd.n2534 vdd.n2533 297.074
R726 vdd.n2280 vdd.n1050 297.074
R727 vdd.n2376 vdd.n1048 297.074
R728 vdd.n2974 vdd.n807 297.074
R729 vdd.n3061 vdd.n3060 297.074
R730 vdd.n2637 vdd.n915 297.074
R731 vdd.n2863 vdd.n916 297.074
R732 vdd.n2531 vdd.n963 297.074
R733 vdd.n961 vdd.n936 297.074
R734 vdd.n2217 vdd.n1051 297.074
R735 vdd.n2374 vdd.n1052 297.074
R736 vdd.n2976 vdd.n807 185
R737 vdd.n3059 vdd.n807 185
R738 vdd.n2978 vdd.n2977 185
R739 vdd.n2977 vdd.n805 185
R740 vdd.n2979 vdd.n839 185
R741 vdd.n2989 vdd.n839 185
R742 vdd.n2980 vdd.n848 185
R743 vdd.n848 vdd.n846 185
R744 vdd.n2982 vdd.n2981 185
R745 vdd.n2983 vdd.n2982 185
R746 vdd.n2935 vdd.n847 185
R747 vdd.n847 vdd.n843 185
R748 vdd.n2934 vdd.n2933 185
R749 vdd.n2933 vdd.n2932 185
R750 vdd.n850 vdd.n849 185
R751 vdd.n851 vdd.n850 185
R752 vdd.n2925 vdd.n2924 185
R753 vdd.n2926 vdd.n2925 185
R754 vdd.n2921 vdd.n860 185
R755 vdd.n860 vdd.n857 185
R756 vdd.n2920 vdd.n2919 185
R757 vdd.n2919 vdd.n2918 185
R758 vdd.n862 vdd.n861 185
R759 vdd.n870 vdd.n862 185
R760 vdd.n2911 vdd.n2910 185
R761 vdd.n2912 vdd.n2911 185
R762 vdd.n2909 vdd.n871 185
R763 vdd.n2760 vdd.n871 185
R764 vdd.n2908 vdd.n2907 185
R765 vdd.n2907 vdd.n2906 185
R766 vdd.n873 vdd.n872 185
R767 vdd.n874 vdd.n873 185
R768 vdd.n2899 vdd.n2898 185
R769 vdd.n2900 vdd.n2899 185
R770 vdd.n2897 vdd.n883 185
R771 vdd.n883 vdd.n880 185
R772 vdd.n2896 vdd.n2895 185
R773 vdd.n2895 vdd.n2894 185
R774 vdd.n885 vdd.n884 185
R775 vdd.n893 vdd.n885 185
R776 vdd.n2887 vdd.n2886 185
R777 vdd.n2888 vdd.n2887 185
R778 vdd.n2885 vdd.n894 185
R779 vdd.n900 vdd.n894 185
R780 vdd.n2884 vdd.n2883 185
R781 vdd.n2883 vdd.n2882 185
R782 vdd.n896 vdd.n895 185
R783 vdd.n897 vdd.n896 185
R784 vdd.n2875 vdd.n2874 185
R785 vdd.n2876 vdd.n2875 185
R786 vdd.n2873 vdd.n906 185
R787 vdd.n2781 vdd.n906 185
R788 vdd.n2872 vdd.n2871 185
R789 vdd.n2871 vdd.n2870 185
R790 vdd.n908 vdd.n907 185
R791 vdd.t119 vdd.n908 185
R792 vdd.n2863 vdd.n2862 185
R793 vdd.n2864 vdd.n2863 185
R794 vdd.n2861 vdd.n916 185
R795 vdd.n2860 vdd.n2859 185
R796 vdd.n918 vdd.n917 185
R797 vdd.n2646 vdd.n2645 185
R798 vdd.n2648 vdd.n2647 185
R799 vdd.n2650 vdd.n2649 185
R800 vdd.n2652 vdd.n2651 185
R801 vdd.n2654 vdd.n2653 185
R802 vdd.n2656 vdd.n2655 185
R803 vdd.n2658 vdd.n2657 185
R804 vdd.n2660 vdd.n2659 185
R805 vdd.n2662 vdd.n2661 185
R806 vdd.n2664 vdd.n2663 185
R807 vdd.n2666 vdd.n2665 185
R808 vdd.n2668 vdd.n2667 185
R809 vdd.n2670 vdd.n2669 185
R810 vdd.n2672 vdd.n2671 185
R811 vdd.n2674 vdd.n2673 185
R812 vdd.n2676 vdd.n2675 185
R813 vdd.n2678 vdd.n2677 185
R814 vdd.n2680 vdd.n2679 185
R815 vdd.n2682 vdd.n2681 185
R816 vdd.n2684 vdd.n2683 185
R817 vdd.n2686 vdd.n2685 185
R818 vdd.n2688 vdd.n2687 185
R819 vdd.n2690 vdd.n2689 185
R820 vdd.n2692 vdd.n2691 185
R821 vdd.n2694 vdd.n2693 185
R822 vdd.n2696 vdd.n2695 185
R823 vdd.n2698 vdd.n2697 185
R824 vdd.n2700 vdd.n2699 185
R825 vdd.n2702 vdd.n2701 185
R826 vdd.n2704 vdd.n2703 185
R827 vdd.n2706 vdd.n2705 185
R828 vdd.n2707 vdd.n2637 185
R829 vdd.n2857 vdd.n2637 185
R830 vdd.n3062 vdd.n3061 185
R831 vdd.n3063 vdd.n798 185
R832 vdd.n3065 vdd.n3064 185
R833 vdd.n3067 vdd.n796 185
R834 vdd.n3069 vdd.n3068 185
R835 vdd.n3070 vdd.n795 185
R836 vdd.n3072 vdd.n3071 185
R837 vdd.n3074 vdd.n793 185
R838 vdd.n3076 vdd.n3075 185
R839 vdd.n3077 vdd.n792 185
R840 vdd.n3079 vdd.n3078 185
R841 vdd.n3081 vdd.n790 185
R842 vdd.n3083 vdd.n3082 185
R843 vdd.n3084 vdd.n789 185
R844 vdd.n3086 vdd.n3085 185
R845 vdd.n3088 vdd.n788 185
R846 vdd.n3089 vdd.n786 185
R847 vdd.n3092 vdd.n3091 185
R848 vdd.n787 vdd.n785 185
R849 vdd.n2948 vdd.n2947 185
R850 vdd.n2950 vdd.n2949 185
R851 vdd.n2952 vdd.n2944 185
R852 vdd.n2954 vdd.n2953 185
R853 vdd.n2955 vdd.n2943 185
R854 vdd.n2957 vdd.n2956 185
R855 vdd.n2959 vdd.n2941 185
R856 vdd.n2961 vdd.n2960 185
R857 vdd.n2962 vdd.n2940 185
R858 vdd.n2964 vdd.n2963 185
R859 vdd.n2966 vdd.n2938 185
R860 vdd.n2968 vdd.n2967 185
R861 vdd.n2969 vdd.n2937 185
R862 vdd.n2971 vdd.n2970 185
R863 vdd.n2973 vdd.n2936 185
R864 vdd.n2975 vdd.n2974 185
R865 vdd.n2974 vdd.n692 185
R866 vdd.n3060 vdd.n802 185
R867 vdd.n3060 vdd.n3059 185
R868 vdd.n2712 vdd.n804 185
R869 vdd.n805 vdd.n804 185
R870 vdd.n2713 vdd.n838 185
R871 vdd.n2989 vdd.n838 185
R872 vdd.n2715 vdd.n2714 185
R873 vdd.n2714 vdd.n846 185
R874 vdd.n2716 vdd.n845 185
R875 vdd.n2983 vdd.n845 185
R876 vdd.n2718 vdd.n2717 185
R877 vdd.n2717 vdd.n843 185
R878 vdd.n2719 vdd.n853 185
R879 vdd.n2932 vdd.n853 185
R880 vdd.n2721 vdd.n2720 185
R881 vdd.n2720 vdd.n851 185
R882 vdd.n2722 vdd.n859 185
R883 vdd.n2926 vdd.n859 185
R884 vdd.n2724 vdd.n2723 185
R885 vdd.n2723 vdd.n857 185
R886 vdd.n2725 vdd.n864 185
R887 vdd.n2918 vdd.n864 185
R888 vdd.n2727 vdd.n2726 185
R889 vdd.n2726 vdd.n870 185
R890 vdd.n2728 vdd.n869 185
R891 vdd.n2912 vdd.n869 185
R892 vdd.n2762 vdd.n2761 185
R893 vdd.n2761 vdd.n2760 185
R894 vdd.n2763 vdd.n876 185
R895 vdd.n2906 vdd.n876 185
R896 vdd.n2765 vdd.n2764 185
R897 vdd.n2764 vdd.n874 185
R898 vdd.n2766 vdd.n882 185
R899 vdd.n2900 vdd.n882 185
R900 vdd.n2768 vdd.n2767 185
R901 vdd.n2767 vdd.n880 185
R902 vdd.n2769 vdd.n887 185
R903 vdd.n2894 vdd.n887 185
R904 vdd.n2771 vdd.n2770 185
R905 vdd.n2770 vdd.n893 185
R906 vdd.n2772 vdd.n892 185
R907 vdd.n2888 vdd.n892 185
R908 vdd.n2774 vdd.n2773 185
R909 vdd.n2773 vdd.n900 185
R910 vdd.n2775 vdd.n899 185
R911 vdd.n2882 vdd.n899 185
R912 vdd.n2777 vdd.n2776 185
R913 vdd.n2776 vdd.n897 185
R914 vdd.n2778 vdd.n905 185
R915 vdd.n2876 vdd.n905 185
R916 vdd.n2780 vdd.n2779 185
R917 vdd.n2781 vdd.n2780 185
R918 vdd.n2711 vdd.n910 185
R919 vdd.n2870 vdd.n910 185
R920 vdd.n2710 vdd.n2709 185
R921 vdd.n2709 vdd.t119 185
R922 vdd.n2708 vdd.n915 185
R923 vdd.n2864 vdd.n915 185
R924 vdd.n2328 vdd.n2327 185
R925 vdd.n2329 vdd.n2328 185
R926 vdd.n1076 vdd.n1074 185
R927 vdd.n1894 vdd.n1074 185
R928 vdd.n1897 vdd.n1896 185
R929 vdd.n1896 vdd.n1895 185
R930 vdd.n1079 vdd.n1078 185
R931 vdd.n1080 vdd.n1079 185
R932 vdd.n1883 vdd.n1882 185
R933 vdd.n1884 vdd.n1883 185
R934 vdd.n1088 vdd.n1087 185
R935 vdd.n1875 vdd.n1087 185
R936 vdd.n1878 vdd.n1877 185
R937 vdd.n1877 vdd.n1876 185
R938 vdd.n1091 vdd.n1090 185
R939 vdd.n1098 vdd.n1091 185
R940 vdd.n1866 vdd.n1865 185
R941 vdd.n1867 vdd.n1866 185
R942 vdd.n1100 vdd.n1099 185
R943 vdd.n1099 vdd.n1097 185
R944 vdd.n1861 vdd.n1860 185
R945 vdd.n1860 vdd.n1859 185
R946 vdd.n1103 vdd.n1102 185
R947 vdd.n1104 vdd.n1103 185
R948 vdd.n1850 vdd.n1849 185
R949 vdd.n1851 vdd.n1850 185
R950 vdd.n1111 vdd.n1110 185
R951 vdd.n1842 vdd.n1110 185
R952 vdd.n1845 vdd.n1844 185
R953 vdd.n1844 vdd.n1843 185
R954 vdd.n1114 vdd.n1113 185
R955 vdd.n1120 vdd.n1114 185
R956 vdd.n1833 vdd.n1832 185
R957 vdd.n1834 vdd.n1833 185
R958 vdd.n1122 vdd.n1121 185
R959 vdd.n1825 vdd.n1121 185
R960 vdd.n1828 vdd.n1827 185
R961 vdd.n1827 vdd.n1826 185
R962 vdd.n1125 vdd.n1124 185
R963 vdd.n1126 vdd.n1125 185
R964 vdd.n1816 vdd.n1815 185
R965 vdd.n1817 vdd.n1816 185
R966 vdd.n1134 vdd.n1133 185
R967 vdd.n1133 vdd.n1132 185
R968 vdd.n1504 vdd.n1503 185
R969 vdd.n1503 vdd.n1502 185
R970 vdd.n1137 vdd.n1136 185
R971 vdd.n1143 vdd.n1137 185
R972 vdd.n1493 vdd.n1492 185
R973 vdd.n1494 vdd.n1493 185
R974 vdd.n1145 vdd.n1144 185
R975 vdd.n1485 vdd.n1144 185
R976 vdd.n1488 vdd.n1487 185
R977 vdd.n1487 vdd.n1486 185
R978 vdd.n1148 vdd.n1147 185
R979 vdd.n1155 vdd.n1148 185
R980 vdd.n1476 vdd.n1475 185
R981 vdd.n1477 vdd.n1476 185
R982 vdd.n1157 vdd.n1156 185
R983 vdd.n1156 vdd.n1154 185
R984 vdd.n1471 vdd.n1470 185
R985 vdd.n1470 vdd.n1469 185
R986 vdd.n1160 vdd.n1159 185
R987 vdd.n1161 vdd.n1160 185
R988 vdd.n1460 vdd.n1459 185
R989 vdd.n1461 vdd.n1460 185
R990 vdd.n1168 vdd.n1167 185
R991 vdd.n1452 vdd.n1167 185
R992 vdd.n1455 vdd.n1454 185
R993 vdd.n1454 vdd.n1453 185
R994 vdd.n1171 vdd.n1170 185
R995 vdd.n1177 vdd.n1171 185
R996 vdd.n1443 vdd.n1442 185
R997 vdd.n1444 vdd.n1443 185
R998 vdd.n1179 vdd.n1178 185
R999 vdd.n1435 vdd.n1178 185
R1000 vdd.n1438 vdd.n1437 185
R1001 vdd.n1437 vdd.n1436 185
R1002 vdd.n1182 vdd.n1181 185
R1003 vdd.n1183 vdd.n1182 185
R1004 vdd.n1426 vdd.n1425 185
R1005 vdd.n1427 vdd.n1426 185
R1006 vdd.n1190 vdd.n1189 185
R1007 vdd.n1225 vdd.n1189 185
R1008 vdd.n1421 vdd.n1420 185
R1009 vdd.n1193 vdd.n1192 185
R1010 vdd.n1417 vdd.n1416 185
R1011 vdd.n1418 vdd.n1417 185
R1012 vdd.n1227 vdd.n1226 185
R1013 vdd.n1412 vdd.n1229 185
R1014 vdd.n1411 vdd.n1230 185
R1015 vdd.n1410 vdd.n1231 185
R1016 vdd.n1233 vdd.n1232 185
R1017 vdd.n1406 vdd.n1235 185
R1018 vdd.n1405 vdd.n1236 185
R1019 vdd.n1404 vdd.n1237 185
R1020 vdd.n1239 vdd.n1238 185
R1021 vdd.n1400 vdd.n1241 185
R1022 vdd.n1399 vdd.n1242 185
R1023 vdd.n1398 vdd.n1243 185
R1024 vdd.n1245 vdd.n1244 185
R1025 vdd.n1394 vdd.n1247 185
R1026 vdd.n1393 vdd.n1248 185
R1027 vdd.n1392 vdd.n1249 185
R1028 vdd.n1253 vdd.n1250 185
R1029 vdd.n1388 vdd.n1255 185
R1030 vdd.n1387 vdd.n1256 185
R1031 vdd.n1386 vdd.n1257 185
R1032 vdd.n1259 vdd.n1258 185
R1033 vdd.n1382 vdd.n1261 185
R1034 vdd.n1381 vdd.n1262 185
R1035 vdd.n1380 vdd.n1263 185
R1036 vdd.n1265 vdd.n1264 185
R1037 vdd.n1376 vdd.n1267 185
R1038 vdd.n1375 vdd.n1268 185
R1039 vdd.n1374 vdd.n1269 185
R1040 vdd.n1271 vdd.n1270 185
R1041 vdd.n1370 vdd.n1273 185
R1042 vdd.n1369 vdd.n1274 185
R1043 vdd.n1368 vdd.n1275 185
R1044 vdd.n1277 vdd.n1276 185
R1045 vdd.n1364 vdd.n1279 185
R1046 vdd.n1363 vdd.n1280 185
R1047 vdd.n1362 vdd.n1281 185
R1048 vdd.n1283 vdd.n1282 185
R1049 vdd.n1358 vdd.n1285 185
R1050 vdd.n1357 vdd.n1354 185
R1051 vdd.n1353 vdd.n1286 185
R1052 vdd.n1288 vdd.n1287 185
R1053 vdd.n1349 vdd.n1290 185
R1054 vdd.n1348 vdd.n1291 185
R1055 vdd.n1347 vdd.n1292 185
R1056 vdd.n1294 vdd.n1293 185
R1057 vdd.n1343 vdd.n1296 185
R1058 vdd.n1342 vdd.n1297 185
R1059 vdd.n1341 vdd.n1298 185
R1060 vdd.n1300 vdd.n1299 185
R1061 vdd.n1337 vdd.n1302 185
R1062 vdd.n1336 vdd.n1303 185
R1063 vdd.n1335 vdd.n1304 185
R1064 vdd.n1306 vdd.n1305 185
R1065 vdd.n1331 vdd.n1308 185
R1066 vdd.n1330 vdd.n1309 185
R1067 vdd.n1329 vdd.n1310 185
R1068 vdd.n1312 vdd.n1311 185
R1069 vdd.n1325 vdd.n1314 185
R1070 vdd.n1324 vdd.n1315 185
R1071 vdd.n1323 vdd.n1316 185
R1072 vdd.n1320 vdd.n1224 185
R1073 vdd.n1418 vdd.n1224 185
R1074 vdd.n2332 vdd.n2331 185
R1075 vdd.n2336 vdd.n1069 185
R1076 vdd.n1999 vdd.n1068 185
R1077 vdd.n2002 vdd.n2001 185
R1078 vdd.n2004 vdd.n2003 185
R1079 vdd.n2007 vdd.n2006 185
R1080 vdd.n2009 vdd.n2008 185
R1081 vdd.n2011 vdd.n1997 185
R1082 vdd.n2013 vdd.n2012 185
R1083 vdd.n2014 vdd.n1991 185
R1084 vdd.n2016 vdd.n2015 185
R1085 vdd.n2018 vdd.n1989 185
R1086 vdd.n2020 vdd.n2019 185
R1087 vdd.n2021 vdd.n1984 185
R1088 vdd.n2023 vdd.n2022 185
R1089 vdd.n2025 vdd.n1982 185
R1090 vdd.n2027 vdd.n2026 185
R1091 vdd.n2028 vdd.n1978 185
R1092 vdd.n2030 vdd.n2029 185
R1093 vdd.n2032 vdd.n1975 185
R1094 vdd.n2034 vdd.n2033 185
R1095 vdd.n1976 vdd.n1969 185
R1096 vdd.n2038 vdd.n1973 185
R1097 vdd.n2039 vdd.n1965 185
R1098 vdd.n2041 vdd.n2040 185
R1099 vdd.n2043 vdd.n1963 185
R1100 vdd.n2045 vdd.n2044 185
R1101 vdd.n2046 vdd.n1958 185
R1102 vdd.n2048 vdd.n2047 185
R1103 vdd.n2050 vdd.n1956 185
R1104 vdd.n2052 vdd.n2051 185
R1105 vdd.n2053 vdd.n1951 185
R1106 vdd.n2055 vdd.n2054 185
R1107 vdd.n2057 vdd.n1949 185
R1108 vdd.n2059 vdd.n2058 185
R1109 vdd.n2060 vdd.n1944 185
R1110 vdd.n2062 vdd.n2061 185
R1111 vdd.n2064 vdd.n1942 185
R1112 vdd.n2066 vdd.n2065 185
R1113 vdd.n2067 vdd.n1938 185
R1114 vdd.n2069 vdd.n2068 185
R1115 vdd.n2071 vdd.n1935 185
R1116 vdd.n2073 vdd.n2072 185
R1117 vdd.n1936 vdd.n1929 185
R1118 vdd.n2077 vdd.n1933 185
R1119 vdd.n2078 vdd.n1925 185
R1120 vdd.n2080 vdd.n2079 185
R1121 vdd.n2082 vdd.n1923 185
R1122 vdd.n2084 vdd.n2083 185
R1123 vdd.n2085 vdd.n1918 185
R1124 vdd.n2087 vdd.n2086 185
R1125 vdd.n2089 vdd.n1916 185
R1126 vdd.n2091 vdd.n2090 185
R1127 vdd.n2092 vdd.n1911 185
R1128 vdd.n2094 vdd.n2093 185
R1129 vdd.n2096 vdd.n1910 185
R1130 vdd.n2097 vdd.n1907 185
R1131 vdd.n2100 vdd.n2099 185
R1132 vdd.n1909 vdd.n1905 185
R1133 vdd.n2317 vdd.n1903 185
R1134 vdd.n2319 vdd.n2318 185
R1135 vdd.n2321 vdd.n1901 185
R1136 vdd.n2323 vdd.n2322 185
R1137 vdd.n2324 vdd.n1075 185
R1138 vdd.n2330 vdd.n1072 185
R1139 vdd.n2330 vdd.n2329 185
R1140 vdd.n1083 vdd.n1071 185
R1141 vdd.n1894 vdd.n1071 185
R1142 vdd.n1893 vdd.n1892 185
R1143 vdd.n1895 vdd.n1893 185
R1144 vdd.n1082 vdd.n1081 185
R1145 vdd.n1081 vdd.n1080 185
R1146 vdd.n1886 vdd.n1885 185
R1147 vdd.n1885 vdd.n1884 185
R1148 vdd.n1086 vdd.n1085 185
R1149 vdd.n1875 vdd.n1086 185
R1150 vdd.n1874 vdd.n1873 185
R1151 vdd.n1876 vdd.n1874 185
R1152 vdd.n1093 vdd.n1092 185
R1153 vdd.n1098 vdd.n1092 185
R1154 vdd.n1869 vdd.n1868 185
R1155 vdd.n1868 vdd.n1867 185
R1156 vdd.n1096 vdd.n1095 185
R1157 vdd.n1097 vdd.n1096 185
R1158 vdd.n1858 vdd.n1857 185
R1159 vdd.n1859 vdd.n1858 185
R1160 vdd.n1106 vdd.n1105 185
R1161 vdd.n1105 vdd.n1104 185
R1162 vdd.n1853 vdd.n1852 185
R1163 vdd.n1852 vdd.n1851 185
R1164 vdd.n1109 vdd.n1108 185
R1165 vdd.n1842 vdd.n1109 185
R1166 vdd.n1841 vdd.n1840 185
R1167 vdd.n1843 vdd.n1841 185
R1168 vdd.n1116 vdd.n1115 185
R1169 vdd.n1120 vdd.n1115 185
R1170 vdd.n1836 vdd.n1835 185
R1171 vdd.n1835 vdd.n1834 185
R1172 vdd.n1119 vdd.n1118 185
R1173 vdd.n1825 vdd.n1119 185
R1174 vdd.n1824 vdd.n1823 185
R1175 vdd.n1826 vdd.n1824 185
R1176 vdd.n1128 vdd.n1127 185
R1177 vdd.n1127 vdd.n1126 185
R1178 vdd.n1819 vdd.n1818 185
R1179 vdd.n1818 vdd.n1817 185
R1180 vdd.n1131 vdd.n1130 185
R1181 vdd.n1132 vdd.n1131 185
R1182 vdd.n1501 vdd.n1500 185
R1183 vdd.n1502 vdd.n1501 185
R1184 vdd.n1139 vdd.n1138 185
R1185 vdd.n1143 vdd.n1138 185
R1186 vdd.n1496 vdd.n1495 185
R1187 vdd.n1495 vdd.n1494 185
R1188 vdd.n1142 vdd.n1141 185
R1189 vdd.n1485 vdd.n1142 185
R1190 vdd.n1484 vdd.n1483 185
R1191 vdd.n1486 vdd.n1484 185
R1192 vdd.n1150 vdd.n1149 185
R1193 vdd.n1155 vdd.n1149 185
R1194 vdd.n1479 vdd.n1478 185
R1195 vdd.n1478 vdd.n1477 185
R1196 vdd.n1153 vdd.n1152 185
R1197 vdd.n1154 vdd.n1153 185
R1198 vdd.n1468 vdd.n1467 185
R1199 vdd.n1469 vdd.n1468 185
R1200 vdd.n1163 vdd.n1162 185
R1201 vdd.n1162 vdd.n1161 185
R1202 vdd.n1463 vdd.n1462 185
R1203 vdd.n1462 vdd.n1461 185
R1204 vdd.n1166 vdd.n1165 185
R1205 vdd.n1452 vdd.n1166 185
R1206 vdd.n1451 vdd.n1450 185
R1207 vdd.n1453 vdd.n1451 185
R1208 vdd.n1173 vdd.n1172 185
R1209 vdd.n1177 vdd.n1172 185
R1210 vdd.n1446 vdd.n1445 185
R1211 vdd.n1445 vdd.n1444 185
R1212 vdd.n1176 vdd.n1175 185
R1213 vdd.n1435 vdd.n1176 185
R1214 vdd.n1434 vdd.n1433 185
R1215 vdd.n1436 vdd.n1434 185
R1216 vdd.n1185 vdd.n1184 185
R1217 vdd.n1184 vdd.n1183 185
R1218 vdd.n1429 vdd.n1428 185
R1219 vdd.n1428 vdd.n1427 185
R1220 vdd.n1188 vdd.n1187 185
R1221 vdd.n1225 vdd.n1188 185
R1222 vdd.n956 vdd.n954 185
R1223 vdd.n2532 vdd.n954 185
R1224 vdd.n2454 vdd.n973 185
R1225 vdd.n973 vdd.t109 185
R1226 vdd.n2456 vdd.n2455 185
R1227 vdd.n2457 vdd.n2456 185
R1228 vdd.n2453 vdd.n972 185
R1229 vdd.n2156 vdd.n972 185
R1230 vdd.n2452 vdd.n2451 185
R1231 vdd.n2451 vdd.n2450 185
R1232 vdd.n975 vdd.n974 185
R1233 vdd.n976 vdd.n975 185
R1234 vdd.n2441 vdd.n2440 185
R1235 vdd.n2442 vdd.n2441 185
R1236 vdd.n2439 vdd.n986 185
R1237 vdd.n986 vdd.n983 185
R1238 vdd.n2438 vdd.n2437 185
R1239 vdd.n2437 vdd.n2436 185
R1240 vdd.n988 vdd.n987 185
R1241 vdd.n989 vdd.n988 185
R1242 vdd.n2429 vdd.n2428 185
R1243 vdd.n2430 vdd.n2429 185
R1244 vdd.n2427 vdd.n997 185
R1245 vdd.n1002 vdd.n997 185
R1246 vdd.n2426 vdd.n2425 185
R1247 vdd.n2425 vdd.n2424 185
R1248 vdd.n999 vdd.n998 185
R1249 vdd.n1008 vdd.n999 185
R1250 vdd.n2417 vdd.n2416 185
R1251 vdd.n2418 vdd.n2417 185
R1252 vdd.n2415 vdd.n1009 185
R1253 vdd.n2257 vdd.n1009 185
R1254 vdd.n2414 vdd.n2413 185
R1255 vdd.n2413 vdd.n2412 185
R1256 vdd.n1011 vdd.n1010 185
R1257 vdd.n1012 vdd.n1011 185
R1258 vdd.n2405 vdd.n2404 185
R1259 vdd.n2406 vdd.n2405 185
R1260 vdd.n2403 vdd.n1021 185
R1261 vdd.n1021 vdd.n1018 185
R1262 vdd.n2402 vdd.n2401 185
R1263 vdd.n2401 vdd.n2400 185
R1264 vdd.n1023 vdd.n1022 185
R1265 vdd.n1033 vdd.n1023 185
R1266 vdd.n2392 vdd.n2391 185
R1267 vdd.n2393 vdd.n2392 185
R1268 vdd.n2390 vdd.n1034 185
R1269 vdd.n1034 vdd.n1030 185
R1270 vdd.n2389 vdd.n2388 185
R1271 vdd.n2388 vdd.n2387 185
R1272 vdd.n1036 vdd.n1035 185
R1273 vdd.n1037 vdd.n1036 185
R1274 vdd.n2380 vdd.n2379 185
R1275 vdd.n2381 vdd.n2380 185
R1276 vdd.n2378 vdd.n1046 185
R1277 vdd.n1046 vdd.n1043 185
R1278 vdd.n2377 vdd.n2376 185
R1279 vdd.n2376 vdd.n2375 185
R1280 vdd.n1048 vdd.n1047 185
R1281 vdd.n2112 vdd.n2111 185
R1282 vdd.n2113 vdd.n2109 185
R1283 vdd.n2109 vdd.n1049 185
R1284 vdd.n2115 vdd.n2114 185
R1285 vdd.n2117 vdd.n2108 185
R1286 vdd.n2120 vdd.n2119 185
R1287 vdd.n2121 vdd.n2107 185
R1288 vdd.n2123 vdd.n2122 185
R1289 vdd.n2125 vdd.n2106 185
R1290 vdd.n2128 vdd.n2127 185
R1291 vdd.n2129 vdd.n2105 185
R1292 vdd.n2131 vdd.n2130 185
R1293 vdd.n2133 vdd.n2104 185
R1294 vdd.n2136 vdd.n2135 185
R1295 vdd.n2137 vdd.n2103 185
R1296 vdd.n2139 vdd.n2138 185
R1297 vdd.n2141 vdd.n2102 185
R1298 vdd.n2314 vdd.n2142 185
R1299 vdd.n2313 vdd.n2312 185
R1300 vdd.n2310 vdd.n2143 185
R1301 vdd.n2308 vdd.n2307 185
R1302 vdd.n2306 vdd.n2144 185
R1303 vdd.n2305 vdd.n2304 185
R1304 vdd.n2302 vdd.n2145 185
R1305 vdd.n2300 vdd.n2299 185
R1306 vdd.n2298 vdd.n2146 185
R1307 vdd.n2297 vdd.n2296 185
R1308 vdd.n2294 vdd.n2147 185
R1309 vdd.n2292 vdd.n2291 185
R1310 vdd.n2290 vdd.n2148 185
R1311 vdd.n2289 vdd.n2288 185
R1312 vdd.n2286 vdd.n2149 185
R1313 vdd.n2284 vdd.n2283 185
R1314 vdd.n2282 vdd.n2150 185
R1315 vdd.n2281 vdd.n2280 185
R1316 vdd.n2535 vdd.n2534 185
R1317 vdd.n2537 vdd.n2536 185
R1318 vdd.n2539 vdd.n2538 185
R1319 vdd.n2542 vdd.n2541 185
R1320 vdd.n2544 vdd.n2543 185
R1321 vdd.n2546 vdd.n2545 185
R1322 vdd.n2548 vdd.n2547 185
R1323 vdd.n2550 vdd.n2549 185
R1324 vdd.n2552 vdd.n2551 185
R1325 vdd.n2554 vdd.n2553 185
R1326 vdd.n2556 vdd.n2555 185
R1327 vdd.n2558 vdd.n2557 185
R1328 vdd.n2560 vdd.n2559 185
R1329 vdd.n2562 vdd.n2561 185
R1330 vdd.n2564 vdd.n2563 185
R1331 vdd.n2566 vdd.n2565 185
R1332 vdd.n2568 vdd.n2567 185
R1333 vdd.n2570 vdd.n2569 185
R1334 vdd.n2572 vdd.n2571 185
R1335 vdd.n2574 vdd.n2573 185
R1336 vdd.n2576 vdd.n2575 185
R1337 vdd.n2578 vdd.n2577 185
R1338 vdd.n2580 vdd.n2579 185
R1339 vdd.n2582 vdd.n2581 185
R1340 vdd.n2584 vdd.n2583 185
R1341 vdd.n2586 vdd.n2585 185
R1342 vdd.n2588 vdd.n2587 185
R1343 vdd.n2590 vdd.n2589 185
R1344 vdd.n2592 vdd.n2591 185
R1345 vdd.n2594 vdd.n2593 185
R1346 vdd.n2596 vdd.n2595 185
R1347 vdd.n2598 vdd.n2597 185
R1348 vdd.n2600 vdd.n2599 185
R1349 vdd.n2601 vdd.n955 185
R1350 vdd.n2603 vdd.n2602 185
R1351 vdd.n2604 vdd.n2603 185
R1352 vdd.n2533 vdd.n959 185
R1353 vdd.n2533 vdd.n2532 185
R1354 vdd.n2154 vdd.n960 185
R1355 vdd.t109 vdd.n960 185
R1356 vdd.n2155 vdd.n970 185
R1357 vdd.n2457 vdd.n970 185
R1358 vdd.n2158 vdd.n2157 185
R1359 vdd.n2157 vdd.n2156 185
R1360 vdd.n2159 vdd.n977 185
R1361 vdd.n2450 vdd.n977 185
R1362 vdd.n2161 vdd.n2160 185
R1363 vdd.n2160 vdd.n976 185
R1364 vdd.n2162 vdd.n984 185
R1365 vdd.n2442 vdd.n984 185
R1366 vdd.n2164 vdd.n2163 185
R1367 vdd.n2163 vdd.n983 185
R1368 vdd.n2165 vdd.n990 185
R1369 vdd.n2436 vdd.n990 185
R1370 vdd.n2167 vdd.n2166 185
R1371 vdd.n2166 vdd.n989 185
R1372 vdd.n2168 vdd.n995 185
R1373 vdd.n2430 vdd.n995 185
R1374 vdd.n2170 vdd.n2169 185
R1375 vdd.n2169 vdd.n1002 185
R1376 vdd.n2171 vdd.n1000 185
R1377 vdd.n2424 vdd.n1000 185
R1378 vdd.n2173 vdd.n2172 185
R1379 vdd.n2172 vdd.n1008 185
R1380 vdd.n2174 vdd.n1006 185
R1381 vdd.n2418 vdd.n1006 185
R1382 vdd.n2259 vdd.n2258 185
R1383 vdd.n2258 vdd.n2257 185
R1384 vdd.n2260 vdd.n1013 185
R1385 vdd.n2412 vdd.n1013 185
R1386 vdd.n2262 vdd.n2261 185
R1387 vdd.n2261 vdd.n1012 185
R1388 vdd.n2263 vdd.n1019 185
R1389 vdd.n2406 vdd.n1019 185
R1390 vdd.n2265 vdd.n2264 185
R1391 vdd.n2264 vdd.n1018 185
R1392 vdd.n2266 vdd.n1024 185
R1393 vdd.n2400 vdd.n1024 185
R1394 vdd.n2268 vdd.n2267 185
R1395 vdd.n2267 vdd.n1033 185
R1396 vdd.n2269 vdd.n1031 185
R1397 vdd.n2393 vdd.n1031 185
R1398 vdd.n2271 vdd.n2270 185
R1399 vdd.n2270 vdd.n1030 185
R1400 vdd.n2272 vdd.n1038 185
R1401 vdd.n2387 vdd.n1038 185
R1402 vdd.n2274 vdd.n2273 185
R1403 vdd.n2273 vdd.n1037 185
R1404 vdd.n2275 vdd.n1044 185
R1405 vdd.n2381 vdd.n1044 185
R1406 vdd.n2277 vdd.n2276 185
R1407 vdd.n2276 vdd.n1043 185
R1408 vdd.n2278 vdd.n1050 185
R1409 vdd.n2375 vdd.n1050 185
R1410 vdd.n3357 vdd.n3356 185
R1411 vdd.n3356 vdd.n3355 185
R1412 vdd.n3358 vdd.n387 185
R1413 vdd.n387 vdd.n386 185
R1414 vdd.n3360 vdd.n3359 185
R1415 vdd.n3361 vdd.n3360 185
R1416 vdd.n382 vdd.n381 185
R1417 vdd.n3362 vdd.n382 185
R1418 vdd.n3365 vdd.n3364 185
R1419 vdd.n3364 vdd.n3363 185
R1420 vdd.n3366 vdd.n376 185
R1421 vdd.n376 vdd.n375 185
R1422 vdd.n3368 vdd.n3367 185
R1423 vdd.n3369 vdd.n3368 185
R1424 vdd.n371 vdd.n370 185
R1425 vdd.n3370 vdd.n371 185
R1426 vdd.n3373 vdd.n3372 185
R1427 vdd.n3372 vdd.n3371 185
R1428 vdd.n3374 vdd.n365 185
R1429 vdd.n3331 vdd.n365 185
R1430 vdd.n3376 vdd.n3375 185
R1431 vdd.n3377 vdd.n3376 185
R1432 vdd.n360 vdd.n359 185
R1433 vdd.n3378 vdd.n360 185
R1434 vdd.n3381 vdd.n3380 185
R1435 vdd.n3380 vdd.n3379 185
R1436 vdd.n3382 vdd.n354 185
R1437 vdd.n361 vdd.n354 185
R1438 vdd.n3384 vdd.n3383 185
R1439 vdd.n3385 vdd.n3384 185
R1440 vdd.n350 vdd.n349 185
R1441 vdd.n3386 vdd.n350 185
R1442 vdd.n3389 vdd.n3388 185
R1443 vdd.n3388 vdd.n3387 185
R1444 vdd.n3390 vdd.n345 185
R1445 vdd.n345 vdd.n344 185
R1446 vdd.n3392 vdd.n3391 185
R1447 vdd.n3393 vdd.n3392 185
R1448 vdd.n339 vdd.n337 185
R1449 vdd.n3394 vdd.n339 185
R1450 vdd.n3397 vdd.n3396 185
R1451 vdd.n3396 vdd.n3395 185
R1452 vdd.n338 vdd.n336 185
R1453 vdd.n340 vdd.n338 185
R1454 vdd.n3307 vdd.n3306 185
R1455 vdd.n3308 vdd.n3307 185
R1456 vdd.n635 vdd.n634 185
R1457 vdd.n634 vdd.n633 185
R1458 vdd.n3302 vdd.n3301 185
R1459 vdd.n3301 vdd.n3300 185
R1460 vdd.n638 vdd.n637 185
R1461 vdd.n644 vdd.n638 185
R1462 vdd.n3288 vdd.n3287 185
R1463 vdd.n3289 vdd.n3288 185
R1464 vdd.n646 vdd.n645 185
R1465 vdd.n3280 vdd.n645 185
R1466 vdd.n3283 vdd.n3282 185
R1467 vdd.n3282 vdd.n3281 185
R1468 vdd.n649 vdd.n648 185
R1469 vdd.n656 vdd.n649 185
R1470 vdd.n3271 vdd.n3270 185
R1471 vdd.n3272 vdd.n3271 185
R1472 vdd.n658 vdd.n657 185
R1473 vdd.n657 vdd.n655 185
R1474 vdd.n3266 vdd.n3265 185
R1475 vdd.n3265 vdd.n3264 185
R1476 vdd.n661 vdd.n660 185
R1477 vdd.n662 vdd.n661 185
R1478 vdd.n3255 vdd.n3254 185
R1479 vdd.n3256 vdd.n3255 185
R1480 vdd.n669 vdd.n668 185
R1481 vdd.n3247 vdd.n668 185
R1482 vdd.n3250 vdd.n3249 185
R1483 vdd.n3249 vdd.n3248 185
R1484 vdd.n672 vdd.n671 185
R1485 vdd.n679 vdd.n672 185
R1486 vdd.n3238 vdd.n3237 185
R1487 vdd.n3239 vdd.n3238 185
R1488 vdd.n681 vdd.n680 185
R1489 vdd.n680 vdd.n678 185
R1490 vdd.n3233 vdd.n3232 185
R1491 vdd.n3232 vdd.n3231 185
R1492 vdd.n684 vdd.n683 185
R1493 vdd.n723 vdd.n684 185
R1494 vdd.n3221 vdd.n3220 185
R1495 vdd.n3219 vdd.n725 185
R1496 vdd.n3218 vdd.n724 185
R1497 vdd.n3223 vdd.n724 185
R1498 vdd.n729 vdd.n728 185
R1499 vdd.n733 vdd.n732 185
R1500 vdd.n3214 vdd.n734 185
R1501 vdd.n3213 vdd.n3212 185
R1502 vdd.n3211 vdd.n3210 185
R1503 vdd.n3209 vdd.n3208 185
R1504 vdd.n3207 vdd.n3206 185
R1505 vdd.n3205 vdd.n3204 185
R1506 vdd.n3203 vdd.n3202 185
R1507 vdd.n3201 vdd.n3200 185
R1508 vdd.n3199 vdd.n3198 185
R1509 vdd.n3197 vdd.n3196 185
R1510 vdd.n3195 vdd.n3194 185
R1511 vdd.n3193 vdd.n3192 185
R1512 vdd.n3191 vdd.n3190 185
R1513 vdd.n3189 vdd.n3188 185
R1514 vdd.n3187 vdd.n3186 185
R1515 vdd.n3178 vdd.n747 185
R1516 vdd.n3180 vdd.n3179 185
R1517 vdd.n3177 vdd.n3176 185
R1518 vdd.n3175 vdd.n3174 185
R1519 vdd.n3173 vdd.n3172 185
R1520 vdd.n3171 vdd.n3170 185
R1521 vdd.n3169 vdd.n3168 185
R1522 vdd.n3167 vdd.n3166 185
R1523 vdd.n3165 vdd.n3164 185
R1524 vdd.n3163 vdd.n3162 185
R1525 vdd.n3161 vdd.n3160 185
R1526 vdd.n3159 vdd.n3158 185
R1527 vdd.n3157 vdd.n3156 185
R1528 vdd.n3155 vdd.n3154 185
R1529 vdd.n3153 vdd.n3152 185
R1530 vdd.n3151 vdd.n3150 185
R1531 vdd.n3149 vdd.n3148 185
R1532 vdd.n3147 vdd.n3146 185
R1533 vdd.n3145 vdd.n3144 185
R1534 vdd.n3143 vdd.n3142 185
R1535 vdd.n3141 vdd.n3140 185
R1536 vdd.n3139 vdd.n3138 185
R1537 vdd.n3132 vdd.n767 185
R1538 vdd.n3134 vdd.n3133 185
R1539 vdd.n3131 vdd.n3130 185
R1540 vdd.n3129 vdd.n3128 185
R1541 vdd.n3127 vdd.n3126 185
R1542 vdd.n3125 vdd.n3124 185
R1543 vdd.n3123 vdd.n3122 185
R1544 vdd.n3121 vdd.n3120 185
R1545 vdd.n3119 vdd.n3118 185
R1546 vdd.n3117 vdd.n3116 185
R1547 vdd.n3115 vdd.n3114 185
R1548 vdd.n3113 vdd.n3112 185
R1549 vdd.n3111 vdd.n3110 185
R1550 vdd.n3109 vdd.n3108 185
R1551 vdd.n3107 vdd.n3106 185
R1552 vdd.n3105 vdd.n3104 185
R1553 vdd.n3103 vdd.n3102 185
R1554 vdd.n3101 vdd.n3100 185
R1555 vdd.n3099 vdd.n3098 185
R1556 vdd.n3097 vdd.n3096 185
R1557 vdd.n3095 vdd.n691 185
R1558 vdd.n3225 vdd.n3224 185
R1559 vdd.n3224 vdd.n3223 185
R1560 vdd.n3352 vdd.n3351 185
R1561 vdd.n618 vdd.n425 185
R1562 vdd.n617 vdd.n616 185
R1563 vdd.n615 vdd.n614 185
R1564 vdd.n613 vdd.n430 185
R1565 vdd.n609 vdd.n608 185
R1566 vdd.n607 vdd.n606 185
R1567 vdd.n605 vdd.n604 185
R1568 vdd.n603 vdd.n432 185
R1569 vdd.n599 vdd.n598 185
R1570 vdd.n597 vdd.n596 185
R1571 vdd.n595 vdd.n594 185
R1572 vdd.n593 vdd.n434 185
R1573 vdd.n589 vdd.n588 185
R1574 vdd.n587 vdd.n586 185
R1575 vdd.n585 vdd.n584 185
R1576 vdd.n583 vdd.n436 185
R1577 vdd.n579 vdd.n578 185
R1578 vdd.n577 vdd.n576 185
R1579 vdd.n575 vdd.n574 185
R1580 vdd.n573 vdd.n438 185
R1581 vdd.n569 vdd.n568 185
R1582 vdd.n567 vdd.n566 185
R1583 vdd.n565 vdd.n564 185
R1584 vdd.n563 vdd.n442 185
R1585 vdd.n559 vdd.n558 185
R1586 vdd.n557 vdd.n556 185
R1587 vdd.n555 vdd.n554 185
R1588 vdd.n553 vdd.n444 185
R1589 vdd.n549 vdd.n548 185
R1590 vdd.n547 vdd.n546 185
R1591 vdd.n545 vdd.n544 185
R1592 vdd.n543 vdd.n446 185
R1593 vdd.n539 vdd.n538 185
R1594 vdd.n537 vdd.n536 185
R1595 vdd.n535 vdd.n534 185
R1596 vdd.n533 vdd.n448 185
R1597 vdd.n529 vdd.n528 185
R1598 vdd.n527 vdd.n526 185
R1599 vdd.n525 vdd.n524 185
R1600 vdd.n523 vdd.n450 185
R1601 vdd.n519 vdd.n518 185
R1602 vdd.n517 vdd.n516 185
R1603 vdd.n515 vdd.n514 185
R1604 vdd.n513 vdd.n454 185
R1605 vdd.n509 vdd.n508 185
R1606 vdd.n507 vdd.n506 185
R1607 vdd.n505 vdd.n504 185
R1608 vdd.n503 vdd.n456 185
R1609 vdd.n499 vdd.n498 185
R1610 vdd.n497 vdd.n496 185
R1611 vdd.n495 vdd.n494 185
R1612 vdd.n493 vdd.n458 185
R1613 vdd.n489 vdd.n488 185
R1614 vdd.n487 vdd.n486 185
R1615 vdd.n485 vdd.n484 185
R1616 vdd.n483 vdd.n460 185
R1617 vdd.n479 vdd.n478 185
R1618 vdd.n477 vdd.n476 185
R1619 vdd.n475 vdd.n474 185
R1620 vdd.n473 vdd.n462 185
R1621 vdd.n469 vdd.n468 185
R1622 vdd.n467 vdd.n466 185
R1623 vdd.n465 vdd.n392 185
R1624 vdd.n3348 vdd.n393 185
R1625 vdd.n3355 vdd.n393 185
R1626 vdd.n3347 vdd.n3346 185
R1627 vdd.n3346 vdd.n386 185
R1628 vdd.n3345 vdd.n385 185
R1629 vdd.n3361 vdd.n385 185
R1630 vdd.n621 vdd.n384 185
R1631 vdd.n3362 vdd.n384 185
R1632 vdd.n3341 vdd.n383 185
R1633 vdd.n3363 vdd.n383 185
R1634 vdd.n3340 vdd.n3339 185
R1635 vdd.n3339 vdd.n375 185
R1636 vdd.n3338 vdd.n374 185
R1637 vdd.n3369 vdd.n374 185
R1638 vdd.n623 vdd.n373 185
R1639 vdd.n3370 vdd.n373 185
R1640 vdd.n3334 vdd.n372 185
R1641 vdd.n3371 vdd.n372 185
R1642 vdd.n3333 vdd.n3332 185
R1643 vdd.n3332 vdd.n3331 185
R1644 vdd.n3330 vdd.n364 185
R1645 vdd.n3377 vdd.n364 185
R1646 vdd.n625 vdd.n363 185
R1647 vdd.n3378 vdd.n363 185
R1648 vdd.n3326 vdd.n362 185
R1649 vdd.n3379 vdd.n362 185
R1650 vdd.n3325 vdd.n3324 185
R1651 vdd.n3324 vdd.n361 185
R1652 vdd.n3323 vdd.n353 185
R1653 vdd.n3385 vdd.n353 185
R1654 vdd.n627 vdd.n352 185
R1655 vdd.n3386 vdd.n352 185
R1656 vdd.n3319 vdd.n351 185
R1657 vdd.n3387 vdd.n351 185
R1658 vdd.n3318 vdd.n3317 185
R1659 vdd.n3317 vdd.n344 185
R1660 vdd.n3316 vdd.n343 185
R1661 vdd.n3393 vdd.n343 185
R1662 vdd.n629 vdd.n342 185
R1663 vdd.n3394 vdd.n342 185
R1664 vdd.n3312 vdd.n341 185
R1665 vdd.n3395 vdd.n341 185
R1666 vdd.n3311 vdd.n3310 185
R1667 vdd.n3310 vdd.n340 185
R1668 vdd.n3309 vdd.n631 185
R1669 vdd.n3309 vdd.n3308 185
R1670 vdd.n3297 vdd.n632 185
R1671 vdd.n633 vdd.n632 185
R1672 vdd.n3299 vdd.n3298 185
R1673 vdd.n3300 vdd.n3299 185
R1674 vdd.n640 vdd.n639 185
R1675 vdd.n644 vdd.n639 185
R1676 vdd.n3291 vdd.n3290 185
R1677 vdd.n3290 vdd.n3289 185
R1678 vdd.n643 vdd.n642 185
R1679 vdd.n3280 vdd.n643 185
R1680 vdd.n3279 vdd.n3278 185
R1681 vdd.n3281 vdd.n3279 185
R1682 vdd.n651 vdd.n650 185
R1683 vdd.n656 vdd.n650 185
R1684 vdd.n3274 vdd.n3273 185
R1685 vdd.n3273 vdd.n3272 185
R1686 vdd.n654 vdd.n653 185
R1687 vdd.n655 vdd.n654 185
R1688 vdd.n3263 vdd.n3262 185
R1689 vdd.n3264 vdd.n3263 185
R1690 vdd.n664 vdd.n663 185
R1691 vdd.n663 vdd.n662 185
R1692 vdd.n3258 vdd.n3257 185
R1693 vdd.n3257 vdd.n3256 185
R1694 vdd.n667 vdd.n666 185
R1695 vdd.n3247 vdd.n667 185
R1696 vdd.n3246 vdd.n3245 185
R1697 vdd.n3248 vdd.n3246 185
R1698 vdd.n674 vdd.n673 185
R1699 vdd.n679 vdd.n673 185
R1700 vdd.n3241 vdd.n3240 185
R1701 vdd.n3240 vdd.n3239 185
R1702 vdd.n677 vdd.n676 185
R1703 vdd.n678 vdd.n677 185
R1704 vdd.n3230 vdd.n3229 185
R1705 vdd.n3231 vdd.n3230 185
R1706 vdd.n686 vdd.n685 185
R1707 vdd.n723 vdd.n685 185
R1708 vdd.n913 vdd.n912 185
R1709 vdd.n2855 vdd.n2854 185
R1710 vdd.n2853 vdd.n2638 185
R1711 vdd.n2857 vdd.n2638 185
R1712 vdd.n2852 vdd.n2851 185
R1713 vdd.n2850 vdd.n2849 185
R1714 vdd.n2848 vdd.n2847 185
R1715 vdd.n2846 vdd.n2845 185
R1716 vdd.n2844 vdd.n2843 185
R1717 vdd.n2842 vdd.n2841 185
R1718 vdd.n2840 vdd.n2839 185
R1719 vdd.n2838 vdd.n2837 185
R1720 vdd.n2836 vdd.n2835 185
R1721 vdd.n2834 vdd.n2833 185
R1722 vdd.n2832 vdd.n2831 185
R1723 vdd.n2830 vdd.n2829 185
R1724 vdd.n2828 vdd.n2827 185
R1725 vdd.n2826 vdd.n2825 185
R1726 vdd.n2824 vdd.n2823 185
R1727 vdd.n2822 vdd.n2821 185
R1728 vdd.n2820 vdd.n2819 185
R1729 vdd.n2818 vdd.n2817 185
R1730 vdd.n2816 vdd.n2815 185
R1731 vdd.n2814 vdd.n2813 185
R1732 vdd.n2812 vdd.n2811 185
R1733 vdd.n2810 vdd.n2809 185
R1734 vdd.n2808 vdd.n2807 185
R1735 vdd.n2806 vdd.n2805 185
R1736 vdd.n2804 vdd.n2803 185
R1737 vdd.n2802 vdd.n2801 185
R1738 vdd.n2800 vdd.n2799 185
R1739 vdd.n2798 vdd.n2797 185
R1740 vdd.n2796 vdd.n2795 185
R1741 vdd.n2793 vdd.n2792 185
R1742 vdd.n2791 vdd.n2790 185
R1743 vdd.n2789 vdd.n2788 185
R1744 vdd.n2995 vdd.n2994 185
R1745 vdd.n2997 vdd.n834 185
R1746 vdd.n2999 vdd.n2998 185
R1747 vdd.n3001 vdd.n831 185
R1748 vdd.n3003 vdd.n3002 185
R1749 vdd.n3005 vdd.n829 185
R1750 vdd.n3007 vdd.n3006 185
R1751 vdd.n3008 vdd.n828 185
R1752 vdd.n3010 vdd.n3009 185
R1753 vdd.n3012 vdd.n826 185
R1754 vdd.n3014 vdd.n3013 185
R1755 vdd.n3015 vdd.n825 185
R1756 vdd.n3017 vdd.n3016 185
R1757 vdd.n3019 vdd.n823 185
R1758 vdd.n3021 vdd.n3020 185
R1759 vdd.n3022 vdd.n822 185
R1760 vdd.n3024 vdd.n3023 185
R1761 vdd.n3026 vdd.n731 185
R1762 vdd.n3028 vdd.n3027 185
R1763 vdd.n3030 vdd.n820 185
R1764 vdd.n3032 vdd.n3031 185
R1765 vdd.n3033 vdd.n819 185
R1766 vdd.n3035 vdd.n3034 185
R1767 vdd.n3037 vdd.n817 185
R1768 vdd.n3039 vdd.n3038 185
R1769 vdd.n3040 vdd.n816 185
R1770 vdd.n3042 vdd.n3041 185
R1771 vdd.n3044 vdd.n814 185
R1772 vdd.n3046 vdd.n3045 185
R1773 vdd.n3047 vdd.n813 185
R1774 vdd.n3049 vdd.n3048 185
R1775 vdd.n3051 vdd.n812 185
R1776 vdd.n3052 vdd.n811 185
R1777 vdd.n3055 vdd.n3054 185
R1778 vdd.n3056 vdd.n809 185
R1779 vdd.n809 vdd.n692 185
R1780 vdd.n2993 vdd.n806 185
R1781 vdd.n3059 vdd.n806 185
R1782 vdd.n2992 vdd.n2991 185
R1783 vdd.n2991 vdd.n805 185
R1784 vdd.n2990 vdd.n836 185
R1785 vdd.n2990 vdd.n2989 185
R1786 vdd.n2744 vdd.n837 185
R1787 vdd.n846 vdd.n837 185
R1788 vdd.n2745 vdd.n844 185
R1789 vdd.n2983 vdd.n844 185
R1790 vdd.n2747 vdd.n2746 185
R1791 vdd.n2746 vdd.n843 185
R1792 vdd.n2748 vdd.n852 185
R1793 vdd.n2932 vdd.n852 185
R1794 vdd.n2750 vdd.n2749 185
R1795 vdd.n2749 vdd.n851 185
R1796 vdd.n2751 vdd.n858 185
R1797 vdd.n2926 vdd.n858 185
R1798 vdd.n2753 vdd.n2752 185
R1799 vdd.n2752 vdd.n857 185
R1800 vdd.n2754 vdd.n863 185
R1801 vdd.n2918 vdd.n863 185
R1802 vdd.n2756 vdd.n2755 185
R1803 vdd.n2755 vdd.n870 185
R1804 vdd.n2757 vdd.n868 185
R1805 vdd.n2912 vdd.n868 185
R1806 vdd.n2759 vdd.n2758 185
R1807 vdd.n2760 vdd.n2759 185
R1808 vdd.n2743 vdd.n875 185
R1809 vdd.n2906 vdd.n875 185
R1810 vdd.n2742 vdd.n2741 185
R1811 vdd.n2741 vdd.n874 185
R1812 vdd.n2740 vdd.n881 185
R1813 vdd.n2900 vdd.n881 185
R1814 vdd.n2739 vdd.n2738 185
R1815 vdd.n2738 vdd.n880 185
R1816 vdd.n2737 vdd.n886 185
R1817 vdd.n2894 vdd.n886 185
R1818 vdd.n2736 vdd.n2735 185
R1819 vdd.n2735 vdd.n893 185
R1820 vdd.n2734 vdd.n891 185
R1821 vdd.n2888 vdd.n891 185
R1822 vdd.n2733 vdd.n2732 185
R1823 vdd.n2732 vdd.n900 185
R1824 vdd.n2731 vdd.n898 185
R1825 vdd.n2882 vdd.n898 185
R1826 vdd.n2730 vdd.n2729 185
R1827 vdd.n2729 vdd.n897 185
R1828 vdd.n2641 vdd.n904 185
R1829 vdd.n2876 vdd.n904 185
R1830 vdd.n2783 vdd.n2782 185
R1831 vdd.n2782 vdd.n2781 185
R1832 vdd.n2784 vdd.n909 185
R1833 vdd.n2870 vdd.n909 185
R1834 vdd.n2786 vdd.n2785 185
R1835 vdd.n2785 vdd.t119 185
R1836 vdd.n2787 vdd.n914 185
R1837 vdd.n2864 vdd.n914 185
R1838 vdd.n2866 vdd.n2865 185
R1839 vdd.n2865 vdd.n2864 185
R1840 vdd.n2867 vdd.n911 185
R1841 vdd.n911 vdd.t119 185
R1842 vdd.n2869 vdd.n2868 185
R1843 vdd.n2870 vdd.n2869 185
R1844 vdd.n903 vdd.n902 185
R1845 vdd.n2781 vdd.n903 185
R1846 vdd.n2878 vdd.n2877 185
R1847 vdd.n2877 vdd.n2876 185
R1848 vdd.n2879 vdd.n901 185
R1849 vdd.n901 vdd.n897 185
R1850 vdd.n2881 vdd.n2880 185
R1851 vdd.n2882 vdd.n2881 185
R1852 vdd.n890 vdd.n889 185
R1853 vdd.n900 vdd.n890 185
R1854 vdd.n2890 vdd.n2889 185
R1855 vdd.n2889 vdd.n2888 185
R1856 vdd.n2891 vdd.n888 185
R1857 vdd.n893 vdd.n888 185
R1858 vdd.n2893 vdd.n2892 185
R1859 vdd.n2894 vdd.n2893 185
R1860 vdd.n879 vdd.n878 185
R1861 vdd.n880 vdd.n879 185
R1862 vdd.n2902 vdd.n2901 185
R1863 vdd.n2901 vdd.n2900 185
R1864 vdd.n2903 vdd.n877 185
R1865 vdd.n877 vdd.n874 185
R1866 vdd.n2905 vdd.n2904 185
R1867 vdd.n2906 vdd.n2905 185
R1868 vdd.n867 vdd.n866 185
R1869 vdd.n2760 vdd.n867 185
R1870 vdd.n2914 vdd.n2913 185
R1871 vdd.n2913 vdd.n2912 185
R1872 vdd.n2915 vdd.n865 185
R1873 vdd.n870 vdd.n865 185
R1874 vdd.n2917 vdd.n2916 185
R1875 vdd.n2918 vdd.n2917 185
R1876 vdd.n856 vdd.n855 185
R1877 vdd.n857 vdd.n856 185
R1878 vdd.n2928 vdd.n2927 185
R1879 vdd.n2927 vdd.n2926 185
R1880 vdd.n2929 vdd.n854 185
R1881 vdd.n854 vdd.n851 185
R1882 vdd.n2931 vdd.n2930 185
R1883 vdd.n2932 vdd.n2931 185
R1884 vdd.n842 vdd.n841 185
R1885 vdd.n843 vdd.n842 185
R1886 vdd.n2985 vdd.n2984 185
R1887 vdd.n2984 vdd.n2983 185
R1888 vdd.n2986 vdd.n840 185
R1889 vdd.n846 vdd.n840 185
R1890 vdd.n2988 vdd.n2987 185
R1891 vdd.n2989 vdd.n2988 185
R1892 vdd.n810 vdd.n808 185
R1893 vdd.n808 vdd.n805 185
R1894 vdd.n3058 vdd.n3057 185
R1895 vdd.n3059 vdd.n3058 185
R1896 vdd.n2531 vdd.n2530 185
R1897 vdd.n2532 vdd.n2531 185
R1898 vdd.n964 vdd.n962 185
R1899 vdd.n962 vdd.t109 185
R1900 vdd.n2446 vdd.n971 185
R1901 vdd.n2457 vdd.n971 185
R1902 vdd.n2447 vdd.n980 185
R1903 vdd.n2156 vdd.n980 185
R1904 vdd.n2449 vdd.n2448 185
R1905 vdd.n2450 vdd.n2449 185
R1906 vdd.n2445 vdd.n979 185
R1907 vdd.n979 vdd.n976 185
R1908 vdd.n2444 vdd.n2443 185
R1909 vdd.n2443 vdd.n2442 185
R1910 vdd.n982 vdd.n981 185
R1911 vdd.n983 vdd.n982 185
R1912 vdd.n2435 vdd.n2434 185
R1913 vdd.n2436 vdd.n2435 185
R1914 vdd.n2433 vdd.n992 185
R1915 vdd.n992 vdd.n989 185
R1916 vdd.n2432 vdd.n2431 185
R1917 vdd.n2431 vdd.n2430 185
R1918 vdd.n994 vdd.n993 185
R1919 vdd.n1002 vdd.n994 185
R1920 vdd.n2423 vdd.n2422 185
R1921 vdd.n2424 vdd.n2423 185
R1922 vdd.n2421 vdd.n1003 185
R1923 vdd.n1008 vdd.n1003 185
R1924 vdd.n2420 vdd.n2419 185
R1925 vdd.n2419 vdd.n2418 185
R1926 vdd.n1005 vdd.n1004 185
R1927 vdd.n2257 vdd.n1005 185
R1928 vdd.n2411 vdd.n2410 185
R1929 vdd.n2412 vdd.n2411 185
R1930 vdd.n2409 vdd.n1015 185
R1931 vdd.n1015 vdd.n1012 185
R1932 vdd.n2408 vdd.n2407 185
R1933 vdd.n2407 vdd.n2406 185
R1934 vdd.n1017 vdd.n1016 185
R1935 vdd.n1018 vdd.n1017 185
R1936 vdd.n2399 vdd.n2398 185
R1937 vdd.n2400 vdd.n2399 185
R1938 vdd.n2396 vdd.n1026 185
R1939 vdd.n1033 vdd.n1026 185
R1940 vdd.n2395 vdd.n2394 185
R1941 vdd.n2394 vdd.n2393 185
R1942 vdd.n1029 vdd.n1028 185
R1943 vdd.n1030 vdd.n1029 185
R1944 vdd.n2386 vdd.n2385 185
R1945 vdd.n2387 vdd.n2386 185
R1946 vdd.n2384 vdd.n1040 185
R1947 vdd.n1040 vdd.n1037 185
R1948 vdd.n2383 vdd.n2382 185
R1949 vdd.n2382 vdd.n2381 185
R1950 vdd.n1042 vdd.n1041 185
R1951 vdd.n1043 vdd.n1042 185
R1952 vdd.n2374 vdd.n2373 185
R1953 vdd.n2375 vdd.n2374 185
R1954 vdd.n2462 vdd.n936 185
R1955 vdd.n2604 vdd.n936 185
R1956 vdd.n2464 vdd.n2463 185
R1957 vdd.n2466 vdd.n2465 185
R1958 vdd.n2468 vdd.n2467 185
R1959 vdd.n2470 vdd.n2469 185
R1960 vdd.n2472 vdd.n2471 185
R1961 vdd.n2474 vdd.n2473 185
R1962 vdd.n2476 vdd.n2475 185
R1963 vdd.n2478 vdd.n2477 185
R1964 vdd.n2480 vdd.n2479 185
R1965 vdd.n2482 vdd.n2481 185
R1966 vdd.n2484 vdd.n2483 185
R1967 vdd.n2486 vdd.n2485 185
R1968 vdd.n2488 vdd.n2487 185
R1969 vdd.n2490 vdd.n2489 185
R1970 vdd.n2492 vdd.n2491 185
R1971 vdd.n2494 vdd.n2493 185
R1972 vdd.n2496 vdd.n2495 185
R1973 vdd.n2498 vdd.n2497 185
R1974 vdd.n2500 vdd.n2499 185
R1975 vdd.n2502 vdd.n2501 185
R1976 vdd.n2504 vdd.n2503 185
R1977 vdd.n2506 vdd.n2505 185
R1978 vdd.n2508 vdd.n2507 185
R1979 vdd.n2510 vdd.n2509 185
R1980 vdd.n2512 vdd.n2511 185
R1981 vdd.n2514 vdd.n2513 185
R1982 vdd.n2516 vdd.n2515 185
R1983 vdd.n2518 vdd.n2517 185
R1984 vdd.n2520 vdd.n2519 185
R1985 vdd.n2522 vdd.n2521 185
R1986 vdd.n2524 vdd.n2523 185
R1987 vdd.n2526 vdd.n2525 185
R1988 vdd.n2528 vdd.n2527 185
R1989 vdd.n2529 vdd.n963 185
R1990 vdd.n2461 vdd.n961 185
R1991 vdd.n2532 vdd.n961 185
R1992 vdd.n2460 vdd.n2459 185
R1993 vdd.n2459 vdd.t109 185
R1994 vdd.n2458 vdd.n968 185
R1995 vdd.n2458 vdd.n2457 185
R1996 vdd.n2238 vdd.n969 185
R1997 vdd.n2156 vdd.n969 185
R1998 vdd.n2239 vdd.n978 185
R1999 vdd.n2450 vdd.n978 185
R2000 vdd.n2241 vdd.n2240 185
R2001 vdd.n2240 vdd.n976 185
R2002 vdd.n2242 vdd.n985 185
R2003 vdd.n2442 vdd.n985 185
R2004 vdd.n2244 vdd.n2243 185
R2005 vdd.n2243 vdd.n983 185
R2006 vdd.n2245 vdd.n991 185
R2007 vdd.n2436 vdd.n991 185
R2008 vdd.n2247 vdd.n2246 185
R2009 vdd.n2246 vdd.n989 185
R2010 vdd.n2248 vdd.n996 185
R2011 vdd.n2430 vdd.n996 185
R2012 vdd.n2250 vdd.n2249 185
R2013 vdd.n2249 vdd.n1002 185
R2014 vdd.n2251 vdd.n1001 185
R2015 vdd.n2424 vdd.n1001 185
R2016 vdd.n2253 vdd.n2252 185
R2017 vdd.n2252 vdd.n1008 185
R2018 vdd.n2254 vdd.n1007 185
R2019 vdd.n2418 vdd.n1007 185
R2020 vdd.n2256 vdd.n2255 185
R2021 vdd.n2257 vdd.n2256 185
R2022 vdd.n2237 vdd.n1014 185
R2023 vdd.n2412 vdd.n1014 185
R2024 vdd.n2236 vdd.n2235 185
R2025 vdd.n2235 vdd.n1012 185
R2026 vdd.n2234 vdd.n1020 185
R2027 vdd.n2406 vdd.n1020 185
R2028 vdd.n2233 vdd.n2232 185
R2029 vdd.n2232 vdd.n1018 185
R2030 vdd.n2231 vdd.n1025 185
R2031 vdd.n2400 vdd.n1025 185
R2032 vdd.n2230 vdd.n2229 185
R2033 vdd.n2229 vdd.n1033 185
R2034 vdd.n2228 vdd.n1032 185
R2035 vdd.n2393 vdd.n1032 185
R2036 vdd.n2227 vdd.n2226 185
R2037 vdd.n2226 vdd.n1030 185
R2038 vdd.n2225 vdd.n1039 185
R2039 vdd.n2387 vdd.n1039 185
R2040 vdd.n2224 vdd.n2223 185
R2041 vdd.n2223 vdd.n1037 185
R2042 vdd.n2222 vdd.n1045 185
R2043 vdd.n2381 vdd.n1045 185
R2044 vdd.n2221 vdd.n2220 185
R2045 vdd.n2220 vdd.n1043 185
R2046 vdd.n2219 vdd.n1051 185
R2047 vdd.n2375 vdd.n1051 185
R2048 vdd.n2372 vdd.n1052 185
R2049 vdd.n2371 vdd.n2370 185
R2050 vdd.n2368 vdd.n1053 185
R2051 vdd.n2366 vdd.n2365 185
R2052 vdd.n2364 vdd.n1054 185
R2053 vdd.n2363 vdd.n2362 185
R2054 vdd.n2360 vdd.n1055 185
R2055 vdd.n2358 vdd.n2357 185
R2056 vdd.n2356 vdd.n1056 185
R2057 vdd.n2355 vdd.n2354 185
R2058 vdd.n2352 vdd.n1057 185
R2059 vdd.n2350 vdd.n2349 185
R2060 vdd.n2348 vdd.n1058 185
R2061 vdd.n2347 vdd.n2346 185
R2062 vdd.n2344 vdd.n1059 185
R2063 vdd.n2342 vdd.n2341 185
R2064 vdd.n2340 vdd.n1060 185
R2065 vdd.n2339 vdd.n1062 185
R2066 vdd.n2184 vdd.n1063 185
R2067 vdd.n2187 vdd.n2186 185
R2068 vdd.n2189 vdd.n2188 185
R2069 vdd.n2191 vdd.n2183 185
R2070 vdd.n2194 vdd.n2193 185
R2071 vdd.n2195 vdd.n2182 185
R2072 vdd.n2197 vdd.n2196 185
R2073 vdd.n2199 vdd.n2181 185
R2074 vdd.n2202 vdd.n2201 185
R2075 vdd.n2203 vdd.n2180 185
R2076 vdd.n2205 vdd.n2204 185
R2077 vdd.n2207 vdd.n2179 185
R2078 vdd.n2210 vdd.n2209 185
R2079 vdd.n2211 vdd.n2176 185
R2080 vdd.n2214 vdd.n2213 185
R2081 vdd.n2216 vdd.n2175 185
R2082 vdd.n2218 vdd.n2217 185
R2083 vdd.n2217 vdd.n1049 185
R2084 vdd.n327 vdd.n326 171.744
R2085 vdd.n326 vdd.n325 171.744
R2086 vdd.n325 vdd.n294 171.744
R2087 vdd.n318 vdd.n294 171.744
R2088 vdd.n318 vdd.n317 171.744
R2089 vdd.n317 vdd.n299 171.744
R2090 vdd.n310 vdd.n299 171.744
R2091 vdd.n310 vdd.n309 171.744
R2092 vdd.n309 vdd.n303 171.744
R2093 vdd.n268 vdd.n267 171.744
R2094 vdd.n267 vdd.n266 171.744
R2095 vdd.n266 vdd.n235 171.744
R2096 vdd.n259 vdd.n235 171.744
R2097 vdd.n259 vdd.n258 171.744
R2098 vdd.n258 vdd.n240 171.744
R2099 vdd.n251 vdd.n240 171.744
R2100 vdd.n251 vdd.n250 171.744
R2101 vdd.n250 vdd.n244 171.744
R2102 vdd.n225 vdd.n224 171.744
R2103 vdd.n224 vdd.n223 171.744
R2104 vdd.n223 vdd.n192 171.744
R2105 vdd.n216 vdd.n192 171.744
R2106 vdd.n216 vdd.n215 171.744
R2107 vdd.n215 vdd.n197 171.744
R2108 vdd.n208 vdd.n197 171.744
R2109 vdd.n208 vdd.n207 171.744
R2110 vdd.n207 vdd.n201 171.744
R2111 vdd.n166 vdd.n165 171.744
R2112 vdd.n165 vdd.n164 171.744
R2113 vdd.n164 vdd.n133 171.744
R2114 vdd.n157 vdd.n133 171.744
R2115 vdd.n157 vdd.n156 171.744
R2116 vdd.n156 vdd.n138 171.744
R2117 vdd.n149 vdd.n138 171.744
R2118 vdd.n149 vdd.n148 171.744
R2119 vdd.n148 vdd.n142 171.744
R2120 vdd.n124 vdd.n123 171.744
R2121 vdd.n123 vdd.n122 171.744
R2122 vdd.n122 vdd.n91 171.744
R2123 vdd.n115 vdd.n91 171.744
R2124 vdd.n115 vdd.n114 171.744
R2125 vdd.n114 vdd.n96 171.744
R2126 vdd.n107 vdd.n96 171.744
R2127 vdd.n107 vdd.n106 171.744
R2128 vdd.n106 vdd.n100 171.744
R2129 vdd.n65 vdd.n64 171.744
R2130 vdd.n64 vdd.n63 171.744
R2131 vdd.n63 vdd.n32 171.744
R2132 vdd.n56 vdd.n32 171.744
R2133 vdd.n56 vdd.n55 171.744
R2134 vdd.n55 vdd.n37 171.744
R2135 vdd.n48 vdd.n37 171.744
R2136 vdd.n48 vdd.n47 171.744
R2137 vdd.n47 vdd.n41 171.744
R2138 vdd.n1746 vdd.n1745 171.744
R2139 vdd.n1745 vdd.n1744 171.744
R2140 vdd.n1744 vdd.n1713 171.744
R2141 vdd.n1737 vdd.n1713 171.744
R2142 vdd.n1737 vdd.n1736 171.744
R2143 vdd.n1736 vdd.n1718 171.744
R2144 vdd.n1729 vdd.n1718 171.744
R2145 vdd.n1729 vdd.n1728 171.744
R2146 vdd.n1728 vdd.n1722 171.744
R2147 vdd.n1805 vdd.n1804 171.744
R2148 vdd.n1804 vdd.n1803 171.744
R2149 vdd.n1803 vdd.n1772 171.744
R2150 vdd.n1796 vdd.n1772 171.744
R2151 vdd.n1796 vdd.n1795 171.744
R2152 vdd.n1795 vdd.n1777 171.744
R2153 vdd.n1788 vdd.n1777 171.744
R2154 vdd.n1788 vdd.n1787 171.744
R2155 vdd.n1787 vdd.n1781 171.744
R2156 vdd.n1644 vdd.n1643 171.744
R2157 vdd.n1643 vdd.n1642 171.744
R2158 vdd.n1642 vdd.n1611 171.744
R2159 vdd.n1635 vdd.n1611 171.744
R2160 vdd.n1635 vdd.n1634 171.744
R2161 vdd.n1634 vdd.n1616 171.744
R2162 vdd.n1627 vdd.n1616 171.744
R2163 vdd.n1627 vdd.n1626 171.744
R2164 vdd.n1626 vdd.n1620 171.744
R2165 vdd.n1703 vdd.n1702 171.744
R2166 vdd.n1702 vdd.n1701 171.744
R2167 vdd.n1701 vdd.n1670 171.744
R2168 vdd.n1694 vdd.n1670 171.744
R2169 vdd.n1694 vdd.n1693 171.744
R2170 vdd.n1693 vdd.n1675 171.744
R2171 vdd.n1686 vdd.n1675 171.744
R2172 vdd.n1686 vdd.n1685 171.744
R2173 vdd.n1685 vdd.n1679 171.744
R2174 vdd.n1543 vdd.n1542 171.744
R2175 vdd.n1542 vdd.n1541 171.744
R2176 vdd.n1541 vdd.n1510 171.744
R2177 vdd.n1534 vdd.n1510 171.744
R2178 vdd.n1534 vdd.n1533 171.744
R2179 vdd.n1533 vdd.n1515 171.744
R2180 vdd.n1526 vdd.n1515 171.744
R2181 vdd.n1526 vdd.n1525 171.744
R2182 vdd.n1525 vdd.n1519 171.744
R2183 vdd.n1602 vdd.n1601 171.744
R2184 vdd.n1601 vdd.n1600 171.744
R2185 vdd.n1600 vdd.n1569 171.744
R2186 vdd.n1593 vdd.n1569 171.744
R2187 vdd.n1593 vdd.n1592 171.744
R2188 vdd.n1592 vdd.n1574 171.744
R2189 vdd.n1585 vdd.n1574 171.744
R2190 vdd.n1585 vdd.n1584 171.744
R2191 vdd.n1584 vdd.n1578 171.744
R2192 vdd.n468 vdd.n467 146.341
R2193 vdd.n474 vdd.n473 146.341
R2194 vdd.n478 vdd.n477 146.341
R2195 vdd.n484 vdd.n483 146.341
R2196 vdd.n488 vdd.n487 146.341
R2197 vdd.n494 vdd.n493 146.341
R2198 vdd.n498 vdd.n497 146.341
R2199 vdd.n504 vdd.n503 146.341
R2200 vdd.n508 vdd.n507 146.341
R2201 vdd.n514 vdd.n513 146.341
R2202 vdd.n518 vdd.n517 146.341
R2203 vdd.n524 vdd.n523 146.341
R2204 vdd.n528 vdd.n527 146.341
R2205 vdd.n534 vdd.n533 146.341
R2206 vdd.n538 vdd.n537 146.341
R2207 vdd.n544 vdd.n543 146.341
R2208 vdd.n548 vdd.n547 146.341
R2209 vdd.n554 vdd.n553 146.341
R2210 vdd.n558 vdd.n557 146.341
R2211 vdd.n564 vdd.n563 146.341
R2212 vdd.n568 vdd.n567 146.341
R2213 vdd.n574 vdd.n573 146.341
R2214 vdd.n578 vdd.n577 146.341
R2215 vdd.n584 vdd.n583 146.341
R2216 vdd.n588 vdd.n587 146.341
R2217 vdd.n594 vdd.n593 146.341
R2218 vdd.n598 vdd.n597 146.341
R2219 vdd.n604 vdd.n603 146.341
R2220 vdd.n608 vdd.n607 146.341
R2221 vdd.n614 vdd.n613 146.341
R2222 vdd.n616 vdd.n425 146.341
R2223 vdd.n3230 vdd.n685 146.341
R2224 vdd.n3230 vdd.n677 146.341
R2225 vdd.n3240 vdd.n677 146.341
R2226 vdd.n3240 vdd.n673 146.341
R2227 vdd.n3246 vdd.n673 146.341
R2228 vdd.n3246 vdd.n667 146.341
R2229 vdd.n3257 vdd.n667 146.341
R2230 vdd.n3257 vdd.n663 146.341
R2231 vdd.n3263 vdd.n663 146.341
R2232 vdd.n3263 vdd.n654 146.341
R2233 vdd.n3273 vdd.n654 146.341
R2234 vdd.n3273 vdd.n650 146.341
R2235 vdd.n3279 vdd.n650 146.341
R2236 vdd.n3279 vdd.n643 146.341
R2237 vdd.n3290 vdd.n643 146.341
R2238 vdd.n3290 vdd.n639 146.341
R2239 vdd.n3299 vdd.n639 146.341
R2240 vdd.n3299 vdd.n632 146.341
R2241 vdd.n3309 vdd.n632 146.341
R2242 vdd.n3310 vdd.n3309 146.341
R2243 vdd.n3310 vdd.n341 146.341
R2244 vdd.n342 vdd.n341 146.341
R2245 vdd.n343 vdd.n342 146.341
R2246 vdd.n3317 vdd.n343 146.341
R2247 vdd.n3317 vdd.n351 146.341
R2248 vdd.n352 vdd.n351 146.341
R2249 vdd.n353 vdd.n352 146.341
R2250 vdd.n3324 vdd.n353 146.341
R2251 vdd.n3324 vdd.n362 146.341
R2252 vdd.n363 vdd.n362 146.341
R2253 vdd.n364 vdd.n363 146.341
R2254 vdd.n3332 vdd.n364 146.341
R2255 vdd.n3332 vdd.n372 146.341
R2256 vdd.n373 vdd.n372 146.341
R2257 vdd.n374 vdd.n373 146.341
R2258 vdd.n3339 vdd.n374 146.341
R2259 vdd.n3339 vdd.n383 146.341
R2260 vdd.n384 vdd.n383 146.341
R2261 vdd.n385 vdd.n384 146.341
R2262 vdd.n3346 vdd.n385 146.341
R2263 vdd.n3346 vdd.n393 146.341
R2264 vdd.n725 vdd.n724 146.341
R2265 vdd.n728 vdd.n724 146.341
R2266 vdd.n734 vdd.n733 146.341
R2267 vdd.n3212 vdd.n3211 146.341
R2268 vdd.n3208 vdd.n3207 146.341
R2269 vdd.n3204 vdd.n3203 146.341
R2270 vdd.n3200 vdd.n3199 146.341
R2271 vdd.n3196 vdd.n3195 146.341
R2272 vdd.n3192 vdd.n3191 146.341
R2273 vdd.n3188 vdd.n3187 146.341
R2274 vdd.n3179 vdd.n3178 146.341
R2275 vdd.n3176 vdd.n3175 146.341
R2276 vdd.n3172 vdd.n3171 146.341
R2277 vdd.n3168 vdd.n3167 146.341
R2278 vdd.n3164 vdd.n3163 146.341
R2279 vdd.n3160 vdd.n3159 146.341
R2280 vdd.n3156 vdd.n3155 146.341
R2281 vdd.n3152 vdd.n3151 146.341
R2282 vdd.n3148 vdd.n3147 146.341
R2283 vdd.n3144 vdd.n3143 146.341
R2284 vdd.n3140 vdd.n3139 146.341
R2285 vdd.n3133 vdd.n3132 146.341
R2286 vdd.n3130 vdd.n3129 146.341
R2287 vdd.n3126 vdd.n3125 146.341
R2288 vdd.n3122 vdd.n3121 146.341
R2289 vdd.n3118 vdd.n3117 146.341
R2290 vdd.n3114 vdd.n3113 146.341
R2291 vdd.n3110 vdd.n3109 146.341
R2292 vdd.n3106 vdd.n3105 146.341
R2293 vdd.n3102 vdd.n3101 146.341
R2294 vdd.n3098 vdd.n3097 146.341
R2295 vdd.n3224 vdd.n691 146.341
R2296 vdd.n3232 vdd.n684 146.341
R2297 vdd.n3232 vdd.n680 146.341
R2298 vdd.n3238 vdd.n680 146.341
R2299 vdd.n3238 vdd.n672 146.341
R2300 vdd.n3249 vdd.n672 146.341
R2301 vdd.n3249 vdd.n668 146.341
R2302 vdd.n3255 vdd.n668 146.341
R2303 vdd.n3255 vdd.n661 146.341
R2304 vdd.n3265 vdd.n661 146.341
R2305 vdd.n3265 vdd.n657 146.341
R2306 vdd.n3271 vdd.n657 146.341
R2307 vdd.n3271 vdd.n649 146.341
R2308 vdd.n3282 vdd.n649 146.341
R2309 vdd.n3282 vdd.n645 146.341
R2310 vdd.n3288 vdd.n645 146.341
R2311 vdd.n3288 vdd.n638 146.341
R2312 vdd.n3301 vdd.n638 146.341
R2313 vdd.n3301 vdd.n634 146.341
R2314 vdd.n3307 vdd.n634 146.341
R2315 vdd.n3307 vdd.n338 146.341
R2316 vdd.n3396 vdd.n338 146.341
R2317 vdd.n3396 vdd.n339 146.341
R2318 vdd.n3392 vdd.n339 146.341
R2319 vdd.n3392 vdd.n345 146.341
R2320 vdd.n3388 vdd.n345 146.341
R2321 vdd.n3388 vdd.n350 146.341
R2322 vdd.n3384 vdd.n350 146.341
R2323 vdd.n3384 vdd.n354 146.341
R2324 vdd.n3380 vdd.n354 146.341
R2325 vdd.n3380 vdd.n360 146.341
R2326 vdd.n3376 vdd.n360 146.341
R2327 vdd.n3376 vdd.n365 146.341
R2328 vdd.n3372 vdd.n365 146.341
R2329 vdd.n3372 vdd.n371 146.341
R2330 vdd.n3368 vdd.n371 146.341
R2331 vdd.n3368 vdd.n376 146.341
R2332 vdd.n3364 vdd.n376 146.341
R2333 vdd.n3364 vdd.n382 146.341
R2334 vdd.n3360 vdd.n382 146.341
R2335 vdd.n3360 vdd.n387 146.341
R2336 vdd.n3356 vdd.n387 146.341
R2337 vdd.n2322 vdd.n2321 146.341
R2338 vdd.n2319 vdd.n1903 146.341
R2339 vdd.n2099 vdd.n1909 146.341
R2340 vdd.n2097 vdd.n2096 146.341
R2341 vdd.n2094 vdd.n1911 146.341
R2342 vdd.n2090 vdd.n2089 146.341
R2343 vdd.n2087 vdd.n1918 146.341
R2344 vdd.n2083 vdd.n2082 146.341
R2345 vdd.n2080 vdd.n1925 146.341
R2346 vdd.n1936 vdd.n1933 146.341
R2347 vdd.n2072 vdd.n2071 146.341
R2348 vdd.n2069 vdd.n1938 146.341
R2349 vdd.n2065 vdd.n2064 146.341
R2350 vdd.n2062 vdd.n1944 146.341
R2351 vdd.n2058 vdd.n2057 146.341
R2352 vdd.n2055 vdd.n1951 146.341
R2353 vdd.n2051 vdd.n2050 146.341
R2354 vdd.n2048 vdd.n1958 146.341
R2355 vdd.n2044 vdd.n2043 146.341
R2356 vdd.n2041 vdd.n1965 146.341
R2357 vdd.n1976 vdd.n1973 146.341
R2358 vdd.n2033 vdd.n2032 146.341
R2359 vdd.n2030 vdd.n1978 146.341
R2360 vdd.n2026 vdd.n2025 146.341
R2361 vdd.n2023 vdd.n1984 146.341
R2362 vdd.n2019 vdd.n2018 146.341
R2363 vdd.n2016 vdd.n1991 146.341
R2364 vdd.n2012 vdd.n2011 146.341
R2365 vdd.n2009 vdd.n2006 146.341
R2366 vdd.n2004 vdd.n2001 146.341
R2367 vdd.n1999 vdd.n1069 146.341
R2368 vdd.n1428 vdd.n1188 146.341
R2369 vdd.n1428 vdd.n1184 146.341
R2370 vdd.n1434 vdd.n1184 146.341
R2371 vdd.n1434 vdd.n1176 146.341
R2372 vdd.n1445 vdd.n1176 146.341
R2373 vdd.n1445 vdd.n1172 146.341
R2374 vdd.n1451 vdd.n1172 146.341
R2375 vdd.n1451 vdd.n1166 146.341
R2376 vdd.n1462 vdd.n1166 146.341
R2377 vdd.n1462 vdd.n1162 146.341
R2378 vdd.n1468 vdd.n1162 146.341
R2379 vdd.n1468 vdd.n1153 146.341
R2380 vdd.n1478 vdd.n1153 146.341
R2381 vdd.n1478 vdd.n1149 146.341
R2382 vdd.n1484 vdd.n1149 146.341
R2383 vdd.n1484 vdd.n1142 146.341
R2384 vdd.n1495 vdd.n1142 146.341
R2385 vdd.n1495 vdd.n1138 146.341
R2386 vdd.n1501 vdd.n1138 146.341
R2387 vdd.n1501 vdd.n1131 146.341
R2388 vdd.n1818 vdd.n1131 146.341
R2389 vdd.n1818 vdd.n1127 146.341
R2390 vdd.n1824 vdd.n1127 146.341
R2391 vdd.n1824 vdd.n1119 146.341
R2392 vdd.n1835 vdd.n1119 146.341
R2393 vdd.n1835 vdd.n1115 146.341
R2394 vdd.n1841 vdd.n1115 146.341
R2395 vdd.n1841 vdd.n1109 146.341
R2396 vdd.n1852 vdd.n1109 146.341
R2397 vdd.n1852 vdd.n1105 146.341
R2398 vdd.n1858 vdd.n1105 146.341
R2399 vdd.n1858 vdd.n1096 146.341
R2400 vdd.n1868 vdd.n1096 146.341
R2401 vdd.n1868 vdd.n1092 146.341
R2402 vdd.n1874 vdd.n1092 146.341
R2403 vdd.n1874 vdd.n1086 146.341
R2404 vdd.n1885 vdd.n1086 146.341
R2405 vdd.n1885 vdd.n1081 146.341
R2406 vdd.n1893 vdd.n1081 146.341
R2407 vdd.n1893 vdd.n1071 146.341
R2408 vdd.n2330 vdd.n1071 146.341
R2409 vdd.n1417 vdd.n1193 146.341
R2410 vdd.n1417 vdd.n1226 146.341
R2411 vdd.n1230 vdd.n1229 146.341
R2412 vdd.n1232 vdd.n1231 146.341
R2413 vdd.n1236 vdd.n1235 146.341
R2414 vdd.n1238 vdd.n1237 146.341
R2415 vdd.n1242 vdd.n1241 146.341
R2416 vdd.n1244 vdd.n1243 146.341
R2417 vdd.n1248 vdd.n1247 146.341
R2418 vdd.n1250 vdd.n1249 146.341
R2419 vdd.n1256 vdd.n1255 146.341
R2420 vdd.n1258 vdd.n1257 146.341
R2421 vdd.n1262 vdd.n1261 146.341
R2422 vdd.n1264 vdd.n1263 146.341
R2423 vdd.n1268 vdd.n1267 146.341
R2424 vdd.n1270 vdd.n1269 146.341
R2425 vdd.n1274 vdd.n1273 146.341
R2426 vdd.n1276 vdd.n1275 146.341
R2427 vdd.n1280 vdd.n1279 146.341
R2428 vdd.n1282 vdd.n1281 146.341
R2429 vdd.n1354 vdd.n1285 146.341
R2430 vdd.n1287 vdd.n1286 146.341
R2431 vdd.n1291 vdd.n1290 146.341
R2432 vdd.n1293 vdd.n1292 146.341
R2433 vdd.n1297 vdd.n1296 146.341
R2434 vdd.n1299 vdd.n1298 146.341
R2435 vdd.n1303 vdd.n1302 146.341
R2436 vdd.n1305 vdd.n1304 146.341
R2437 vdd.n1309 vdd.n1308 146.341
R2438 vdd.n1311 vdd.n1310 146.341
R2439 vdd.n1315 vdd.n1314 146.341
R2440 vdd.n1316 vdd.n1224 146.341
R2441 vdd.n1426 vdd.n1189 146.341
R2442 vdd.n1426 vdd.n1182 146.341
R2443 vdd.n1437 vdd.n1182 146.341
R2444 vdd.n1437 vdd.n1178 146.341
R2445 vdd.n1443 vdd.n1178 146.341
R2446 vdd.n1443 vdd.n1171 146.341
R2447 vdd.n1454 vdd.n1171 146.341
R2448 vdd.n1454 vdd.n1167 146.341
R2449 vdd.n1460 vdd.n1167 146.341
R2450 vdd.n1460 vdd.n1160 146.341
R2451 vdd.n1470 vdd.n1160 146.341
R2452 vdd.n1470 vdd.n1156 146.341
R2453 vdd.n1476 vdd.n1156 146.341
R2454 vdd.n1476 vdd.n1148 146.341
R2455 vdd.n1487 vdd.n1148 146.341
R2456 vdd.n1487 vdd.n1144 146.341
R2457 vdd.n1493 vdd.n1144 146.341
R2458 vdd.n1493 vdd.n1137 146.341
R2459 vdd.n1503 vdd.n1137 146.341
R2460 vdd.n1503 vdd.n1133 146.341
R2461 vdd.n1816 vdd.n1133 146.341
R2462 vdd.n1816 vdd.n1125 146.341
R2463 vdd.n1827 vdd.n1125 146.341
R2464 vdd.n1827 vdd.n1121 146.341
R2465 vdd.n1833 vdd.n1121 146.341
R2466 vdd.n1833 vdd.n1114 146.341
R2467 vdd.n1844 vdd.n1114 146.341
R2468 vdd.n1844 vdd.n1110 146.341
R2469 vdd.n1850 vdd.n1110 146.341
R2470 vdd.n1850 vdd.n1103 146.341
R2471 vdd.n1860 vdd.n1103 146.341
R2472 vdd.n1860 vdd.n1099 146.341
R2473 vdd.n1866 vdd.n1099 146.341
R2474 vdd.n1866 vdd.n1091 146.341
R2475 vdd.n1877 vdd.n1091 146.341
R2476 vdd.n1877 vdd.n1087 146.341
R2477 vdd.n1883 vdd.n1087 146.341
R2478 vdd.n1883 vdd.n1079 146.341
R2479 vdd.n1896 vdd.n1079 146.341
R2480 vdd.n1896 vdd.n1074 146.341
R2481 vdd.n2328 vdd.n1074 146.341
R2482 vdd.n1073 vdd.n1049 141.707
R2483 vdd.n3223 vdd.n692 141.707
R2484 vdd.n2177 vdd.t67 127.284
R2485 vdd.n965 vdd.t52 127.284
R2486 vdd.n2151 vdd.t14 127.284
R2487 vdd.n957 vdd.t76 127.284
R2488 vdd.n2922 vdd.t28 127.284
R2489 vdd.n2922 vdd.t29 127.284
R2490 vdd.n2642 vdd.t74 127.284
R2491 vdd.n832 vdd.t56 127.284
R2492 vdd.n2639 vdd.t61 127.284
R2493 vdd.n799 vdd.t63 127.284
R2494 vdd.n1027 vdd.t70 127.284
R2495 vdd.n1027 vdd.t71 127.284
R2496 vdd.n22 vdd.n20 117.314
R2497 vdd.n17 vdd.n15 117.314
R2498 vdd.n27 vdd.n26 116.927
R2499 vdd.n24 vdd.n23 116.927
R2500 vdd.n22 vdd.n21 116.927
R2501 vdd.n17 vdd.n16 116.927
R2502 vdd.n19 vdd.n18 116.927
R2503 vdd.n27 vdd.n25 116.927
R2504 vdd.n2178 vdd.t66 111.188
R2505 vdd.n966 vdd.t53 111.188
R2506 vdd.n2152 vdd.t13 111.188
R2507 vdd.n958 vdd.t77 111.188
R2508 vdd.n2643 vdd.t73 111.188
R2509 vdd.n833 vdd.t57 111.188
R2510 vdd.n2640 vdd.t60 111.188
R2511 vdd.n800 vdd.t64 111.188
R2512 vdd.n2865 vdd.n911 99.5127
R2513 vdd.n2869 vdd.n911 99.5127
R2514 vdd.n2869 vdd.n903 99.5127
R2515 vdd.n2877 vdd.n903 99.5127
R2516 vdd.n2877 vdd.n901 99.5127
R2517 vdd.n2881 vdd.n901 99.5127
R2518 vdd.n2881 vdd.n890 99.5127
R2519 vdd.n2889 vdd.n890 99.5127
R2520 vdd.n2889 vdd.n888 99.5127
R2521 vdd.n2893 vdd.n888 99.5127
R2522 vdd.n2893 vdd.n879 99.5127
R2523 vdd.n2901 vdd.n879 99.5127
R2524 vdd.n2901 vdd.n877 99.5127
R2525 vdd.n2905 vdd.n877 99.5127
R2526 vdd.n2905 vdd.n867 99.5127
R2527 vdd.n2913 vdd.n867 99.5127
R2528 vdd.n2913 vdd.n865 99.5127
R2529 vdd.n2917 vdd.n865 99.5127
R2530 vdd.n2917 vdd.n856 99.5127
R2531 vdd.n2927 vdd.n856 99.5127
R2532 vdd.n2927 vdd.n854 99.5127
R2533 vdd.n2931 vdd.n854 99.5127
R2534 vdd.n2931 vdd.n842 99.5127
R2535 vdd.n2984 vdd.n842 99.5127
R2536 vdd.n2984 vdd.n840 99.5127
R2537 vdd.n2988 vdd.n840 99.5127
R2538 vdd.n2988 vdd.n808 99.5127
R2539 vdd.n3058 vdd.n808 99.5127
R2540 vdd.n3054 vdd.n809 99.5127
R2541 vdd.n3052 vdd.n3051 99.5127
R2542 vdd.n3049 vdd.n813 99.5127
R2543 vdd.n3045 vdd.n3044 99.5127
R2544 vdd.n3042 vdd.n816 99.5127
R2545 vdd.n3038 vdd.n3037 99.5127
R2546 vdd.n3035 vdd.n819 99.5127
R2547 vdd.n3031 vdd.n3030 99.5127
R2548 vdd.n3028 vdd.n3026 99.5127
R2549 vdd.n3024 vdd.n822 99.5127
R2550 vdd.n3020 vdd.n3019 99.5127
R2551 vdd.n3017 vdd.n825 99.5127
R2552 vdd.n3013 vdd.n3012 99.5127
R2553 vdd.n3010 vdd.n828 99.5127
R2554 vdd.n3006 vdd.n3005 99.5127
R2555 vdd.n3003 vdd.n831 99.5127
R2556 vdd.n2998 vdd.n2997 99.5127
R2557 vdd.n2785 vdd.n914 99.5127
R2558 vdd.n2785 vdd.n909 99.5127
R2559 vdd.n2782 vdd.n909 99.5127
R2560 vdd.n2782 vdd.n904 99.5127
R2561 vdd.n2729 vdd.n904 99.5127
R2562 vdd.n2729 vdd.n898 99.5127
R2563 vdd.n2732 vdd.n898 99.5127
R2564 vdd.n2732 vdd.n891 99.5127
R2565 vdd.n2735 vdd.n891 99.5127
R2566 vdd.n2735 vdd.n886 99.5127
R2567 vdd.n2738 vdd.n886 99.5127
R2568 vdd.n2738 vdd.n881 99.5127
R2569 vdd.n2741 vdd.n881 99.5127
R2570 vdd.n2741 vdd.n875 99.5127
R2571 vdd.n2759 vdd.n875 99.5127
R2572 vdd.n2759 vdd.n868 99.5127
R2573 vdd.n2755 vdd.n868 99.5127
R2574 vdd.n2755 vdd.n863 99.5127
R2575 vdd.n2752 vdd.n863 99.5127
R2576 vdd.n2752 vdd.n858 99.5127
R2577 vdd.n2749 vdd.n858 99.5127
R2578 vdd.n2749 vdd.n852 99.5127
R2579 vdd.n2746 vdd.n852 99.5127
R2580 vdd.n2746 vdd.n844 99.5127
R2581 vdd.n844 vdd.n837 99.5127
R2582 vdd.n2990 vdd.n837 99.5127
R2583 vdd.n2991 vdd.n2990 99.5127
R2584 vdd.n2991 vdd.n806 99.5127
R2585 vdd.n2855 vdd.n2638 99.5127
R2586 vdd.n2851 vdd.n2638 99.5127
R2587 vdd.n2849 vdd.n2848 99.5127
R2588 vdd.n2845 vdd.n2844 99.5127
R2589 vdd.n2841 vdd.n2840 99.5127
R2590 vdd.n2837 vdd.n2836 99.5127
R2591 vdd.n2833 vdd.n2832 99.5127
R2592 vdd.n2829 vdd.n2828 99.5127
R2593 vdd.n2825 vdd.n2824 99.5127
R2594 vdd.n2821 vdd.n2820 99.5127
R2595 vdd.n2817 vdd.n2816 99.5127
R2596 vdd.n2813 vdd.n2812 99.5127
R2597 vdd.n2809 vdd.n2808 99.5127
R2598 vdd.n2805 vdd.n2804 99.5127
R2599 vdd.n2801 vdd.n2800 99.5127
R2600 vdd.n2797 vdd.n2796 99.5127
R2601 vdd.n2792 vdd.n2791 99.5127
R2602 vdd.n2603 vdd.n955 99.5127
R2603 vdd.n2599 vdd.n2598 99.5127
R2604 vdd.n2595 vdd.n2594 99.5127
R2605 vdd.n2591 vdd.n2590 99.5127
R2606 vdd.n2587 vdd.n2586 99.5127
R2607 vdd.n2583 vdd.n2582 99.5127
R2608 vdd.n2579 vdd.n2578 99.5127
R2609 vdd.n2575 vdd.n2574 99.5127
R2610 vdd.n2571 vdd.n2570 99.5127
R2611 vdd.n2567 vdd.n2566 99.5127
R2612 vdd.n2563 vdd.n2562 99.5127
R2613 vdd.n2559 vdd.n2558 99.5127
R2614 vdd.n2555 vdd.n2554 99.5127
R2615 vdd.n2551 vdd.n2550 99.5127
R2616 vdd.n2547 vdd.n2546 99.5127
R2617 vdd.n2543 vdd.n2542 99.5127
R2618 vdd.n2538 vdd.n2537 99.5127
R2619 vdd.n2276 vdd.n1050 99.5127
R2620 vdd.n2276 vdd.n1044 99.5127
R2621 vdd.n2273 vdd.n1044 99.5127
R2622 vdd.n2273 vdd.n1038 99.5127
R2623 vdd.n2270 vdd.n1038 99.5127
R2624 vdd.n2270 vdd.n1031 99.5127
R2625 vdd.n2267 vdd.n1031 99.5127
R2626 vdd.n2267 vdd.n1024 99.5127
R2627 vdd.n2264 vdd.n1024 99.5127
R2628 vdd.n2264 vdd.n1019 99.5127
R2629 vdd.n2261 vdd.n1019 99.5127
R2630 vdd.n2261 vdd.n1013 99.5127
R2631 vdd.n2258 vdd.n1013 99.5127
R2632 vdd.n2258 vdd.n1006 99.5127
R2633 vdd.n2172 vdd.n1006 99.5127
R2634 vdd.n2172 vdd.n1000 99.5127
R2635 vdd.n2169 vdd.n1000 99.5127
R2636 vdd.n2169 vdd.n995 99.5127
R2637 vdd.n2166 vdd.n995 99.5127
R2638 vdd.n2166 vdd.n990 99.5127
R2639 vdd.n2163 vdd.n990 99.5127
R2640 vdd.n2163 vdd.n984 99.5127
R2641 vdd.n2160 vdd.n984 99.5127
R2642 vdd.n2160 vdd.n977 99.5127
R2643 vdd.n2157 vdd.n977 99.5127
R2644 vdd.n2157 vdd.n970 99.5127
R2645 vdd.n970 vdd.n960 99.5127
R2646 vdd.n2533 vdd.n960 99.5127
R2647 vdd.n2111 vdd.n2109 99.5127
R2648 vdd.n2115 vdd.n2109 99.5127
R2649 vdd.n2119 vdd.n2117 99.5127
R2650 vdd.n2123 vdd.n2107 99.5127
R2651 vdd.n2127 vdd.n2125 99.5127
R2652 vdd.n2131 vdd.n2105 99.5127
R2653 vdd.n2135 vdd.n2133 99.5127
R2654 vdd.n2139 vdd.n2103 99.5127
R2655 vdd.n2142 vdd.n2141 99.5127
R2656 vdd.n2312 vdd.n2310 99.5127
R2657 vdd.n2308 vdd.n2144 99.5127
R2658 vdd.n2304 vdd.n2302 99.5127
R2659 vdd.n2300 vdd.n2146 99.5127
R2660 vdd.n2296 vdd.n2294 99.5127
R2661 vdd.n2292 vdd.n2148 99.5127
R2662 vdd.n2288 vdd.n2286 99.5127
R2663 vdd.n2284 vdd.n2150 99.5127
R2664 vdd.n2376 vdd.n1046 99.5127
R2665 vdd.n2380 vdd.n1046 99.5127
R2666 vdd.n2380 vdd.n1036 99.5127
R2667 vdd.n2388 vdd.n1036 99.5127
R2668 vdd.n2388 vdd.n1034 99.5127
R2669 vdd.n2392 vdd.n1034 99.5127
R2670 vdd.n2392 vdd.n1023 99.5127
R2671 vdd.n2401 vdd.n1023 99.5127
R2672 vdd.n2401 vdd.n1021 99.5127
R2673 vdd.n2405 vdd.n1021 99.5127
R2674 vdd.n2405 vdd.n1011 99.5127
R2675 vdd.n2413 vdd.n1011 99.5127
R2676 vdd.n2413 vdd.n1009 99.5127
R2677 vdd.n2417 vdd.n1009 99.5127
R2678 vdd.n2417 vdd.n999 99.5127
R2679 vdd.n2425 vdd.n999 99.5127
R2680 vdd.n2425 vdd.n997 99.5127
R2681 vdd.n2429 vdd.n997 99.5127
R2682 vdd.n2429 vdd.n988 99.5127
R2683 vdd.n2437 vdd.n988 99.5127
R2684 vdd.n2437 vdd.n986 99.5127
R2685 vdd.n2441 vdd.n986 99.5127
R2686 vdd.n2441 vdd.n975 99.5127
R2687 vdd.n2451 vdd.n975 99.5127
R2688 vdd.n2451 vdd.n972 99.5127
R2689 vdd.n2456 vdd.n972 99.5127
R2690 vdd.n2456 vdd.n973 99.5127
R2691 vdd.n973 vdd.n954 99.5127
R2692 vdd.n2974 vdd.n2973 99.5127
R2693 vdd.n2971 vdd.n2937 99.5127
R2694 vdd.n2967 vdd.n2966 99.5127
R2695 vdd.n2964 vdd.n2940 99.5127
R2696 vdd.n2960 vdd.n2959 99.5127
R2697 vdd.n2957 vdd.n2943 99.5127
R2698 vdd.n2953 vdd.n2952 99.5127
R2699 vdd.n2950 vdd.n2947 99.5127
R2700 vdd.n3091 vdd.n787 99.5127
R2701 vdd.n3089 vdd.n3088 99.5127
R2702 vdd.n3086 vdd.n789 99.5127
R2703 vdd.n3082 vdd.n3081 99.5127
R2704 vdd.n3079 vdd.n792 99.5127
R2705 vdd.n3075 vdd.n3074 99.5127
R2706 vdd.n3072 vdd.n795 99.5127
R2707 vdd.n3068 vdd.n3067 99.5127
R2708 vdd.n3065 vdd.n798 99.5127
R2709 vdd.n2709 vdd.n915 99.5127
R2710 vdd.n2709 vdd.n910 99.5127
R2711 vdd.n2780 vdd.n910 99.5127
R2712 vdd.n2780 vdd.n905 99.5127
R2713 vdd.n2776 vdd.n905 99.5127
R2714 vdd.n2776 vdd.n899 99.5127
R2715 vdd.n2773 vdd.n899 99.5127
R2716 vdd.n2773 vdd.n892 99.5127
R2717 vdd.n2770 vdd.n892 99.5127
R2718 vdd.n2770 vdd.n887 99.5127
R2719 vdd.n2767 vdd.n887 99.5127
R2720 vdd.n2767 vdd.n882 99.5127
R2721 vdd.n2764 vdd.n882 99.5127
R2722 vdd.n2764 vdd.n876 99.5127
R2723 vdd.n2761 vdd.n876 99.5127
R2724 vdd.n2761 vdd.n869 99.5127
R2725 vdd.n2726 vdd.n869 99.5127
R2726 vdd.n2726 vdd.n864 99.5127
R2727 vdd.n2723 vdd.n864 99.5127
R2728 vdd.n2723 vdd.n859 99.5127
R2729 vdd.n2720 vdd.n859 99.5127
R2730 vdd.n2720 vdd.n853 99.5127
R2731 vdd.n2717 vdd.n853 99.5127
R2732 vdd.n2717 vdd.n845 99.5127
R2733 vdd.n2714 vdd.n845 99.5127
R2734 vdd.n2714 vdd.n838 99.5127
R2735 vdd.n838 vdd.n804 99.5127
R2736 vdd.n3060 vdd.n804 99.5127
R2737 vdd.n2859 vdd.n918 99.5127
R2738 vdd.n2647 vdd.n2646 99.5127
R2739 vdd.n2651 vdd.n2650 99.5127
R2740 vdd.n2655 vdd.n2654 99.5127
R2741 vdd.n2659 vdd.n2658 99.5127
R2742 vdd.n2663 vdd.n2662 99.5127
R2743 vdd.n2667 vdd.n2666 99.5127
R2744 vdd.n2671 vdd.n2670 99.5127
R2745 vdd.n2675 vdd.n2674 99.5127
R2746 vdd.n2679 vdd.n2678 99.5127
R2747 vdd.n2683 vdd.n2682 99.5127
R2748 vdd.n2687 vdd.n2686 99.5127
R2749 vdd.n2691 vdd.n2690 99.5127
R2750 vdd.n2695 vdd.n2694 99.5127
R2751 vdd.n2699 vdd.n2698 99.5127
R2752 vdd.n2703 vdd.n2702 99.5127
R2753 vdd.n2705 vdd.n2637 99.5127
R2754 vdd.n2863 vdd.n908 99.5127
R2755 vdd.n2871 vdd.n908 99.5127
R2756 vdd.n2871 vdd.n906 99.5127
R2757 vdd.n2875 vdd.n906 99.5127
R2758 vdd.n2875 vdd.n896 99.5127
R2759 vdd.n2883 vdd.n896 99.5127
R2760 vdd.n2883 vdd.n894 99.5127
R2761 vdd.n2887 vdd.n894 99.5127
R2762 vdd.n2887 vdd.n885 99.5127
R2763 vdd.n2895 vdd.n885 99.5127
R2764 vdd.n2895 vdd.n883 99.5127
R2765 vdd.n2899 vdd.n883 99.5127
R2766 vdd.n2899 vdd.n873 99.5127
R2767 vdd.n2907 vdd.n873 99.5127
R2768 vdd.n2907 vdd.n871 99.5127
R2769 vdd.n2911 vdd.n871 99.5127
R2770 vdd.n2911 vdd.n862 99.5127
R2771 vdd.n2919 vdd.n862 99.5127
R2772 vdd.n2919 vdd.n860 99.5127
R2773 vdd.n2925 vdd.n860 99.5127
R2774 vdd.n2925 vdd.n850 99.5127
R2775 vdd.n2933 vdd.n850 99.5127
R2776 vdd.n2933 vdd.n847 99.5127
R2777 vdd.n2982 vdd.n847 99.5127
R2778 vdd.n2982 vdd.n848 99.5127
R2779 vdd.n848 vdd.n839 99.5127
R2780 vdd.n2977 vdd.n839 99.5127
R2781 vdd.n2977 vdd.n807 99.5127
R2782 vdd.n2527 vdd.n2526 99.5127
R2783 vdd.n2523 vdd.n2522 99.5127
R2784 vdd.n2519 vdd.n2518 99.5127
R2785 vdd.n2515 vdd.n2514 99.5127
R2786 vdd.n2511 vdd.n2510 99.5127
R2787 vdd.n2507 vdd.n2506 99.5127
R2788 vdd.n2503 vdd.n2502 99.5127
R2789 vdd.n2499 vdd.n2498 99.5127
R2790 vdd.n2495 vdd.n2494 99.5127
R2791 vdd.n2491 vdd.n2490 99.5127
R2792 vdd.n2487 vdd.n2486 99.5127
R2793 vdd.n2483 vdd.n2482 99.5127
R2794 vdd.n2479 vdd.n2478 99.5127
R2795 vdd.n2475 vdd.n2474 99.5127
R2796 vdd.n2471 vdd.n2470 99.5127
R2797 vdd.n2467 vdd.n2466 99.5127
R2798 vdd.n2463 vdd.n936 99.5127
R2799 vdd.n2220 vdd.n1051 99.5127
R2800 vdd.n2220 vdd.n1045 99.5127
R2801 vdd.n2223 vdd.n1045 99.5127
R2802 vdd.n2223 vdd.n1039 99.5127
R2803 vdd.n2226 vdd.n1039 99.5127
R2804 vdd.n2226 vdd.n1032 99.5127
R2805 vdd.n2229 vdd.n1032 99.5127
R2806 vdd.n2229 vdd.n1025 99.5127
R2807 vdd.n2232 vdd.n1025 99.5127
R2808 vdd.n2232 vdd.n1020 99.5127
R2809 vdd.n2235 vdd.n1020 99.5127
R2810 vdd.n2235 vdd.n1014 99.5127
R2811 vdd.n2256 vdd.n1014 99.5127
R2812 vdd.n2256 vdd.n1007 99.5127
R2813 vdd.n2252 vdd.n1007 99.5127
R2814 vdd.n2252 vdd.n1001 99.5127
R2815 vdd.n2249 vdd.n1001 99.5127
R2816 vdd.n2249 vdd.n996 99.5127
R2817 vdd.n2246 vdd.n996 99.5127
R2818 vdd.n2246 vdd.n991 99.5127
R2819 vdd.n2243 vdd.n991 99.5127
R2820 vdd.n2243 vdd.n985 99.5127
R2821 vdd.n2240 vdd.n985 99.5127
R2822 vdd.n2240 vdd.n978 99.5127
R2823 vdd.n978 vdd.n969 99.5127
R2824 vdd.n2458 vdd.n969 99.5127
R2825 vdd.n2459 vdd.n2458 99.5127
R2826 vdd.n2459 vdd.n961 99.5127
R2827 vdd.n2370 vdd.n2368 99.5127
R2828 vdd.n2366 vdd.n1054 99.5127
R2829 vdd.n2362 vdd.n2360 99.5127
R2830 vdd.n2358 vdd.n1056 99.5127
R2831 vdd.n2354 vdd.n2352 99.5127
R2832 vdd.n2350 vdd.n1058 99.5127
R2833 vdd.n2346 vdd.n2344 99.5127
R2834 vdd.n2342 vdd.n1060 99.5127
R2835 vdd.n2184 vdd.n1062 99.5127
R2836 vdd.n2189 vdd.n2186 99.5127
R2837 vdd.n2193 vdd.n2191 99.5127
R2838 vdd.n2197 vdd.n2182 99.5127
R2839 vdd.n2201 vdd.n2199 99.5127
R2840 vdd.n2205 vdd.n2180 99.5127
R2841 vdd.n2209 vdd.n2207 99.5127
R2842 vdd.n2214 vdd.n2176 99.5127
R2843 vdd.n2217 vdd.n2216 99.5127
R2844 vdd.n2374 vdd.n1042 99.5127
R2845 vdd.n2382 vdd.n1042 99.5127
R2846 vdd.n2382 vdd.n1040 99.5127
R2847 vdd.n2386 vdd.n1040 99.5127
R2848 vdd.n2386 vdd.n1029 99.5127
R2849 vdd.n2394 vdd.n1029 99.5127
R2850 vdd.n2394 vdd.n1026 99.5127
R2851 vdd.n2399 vdd.n1026 99.5127
R2852 vdd.n2399 vdd.n1017 99.5127
R2853 vdd.n2407 vdd.n1017 99.5127
R2854 vdd.n2407 vdd.n1015 99.5127
R2855 vdd.n2411 vdd.n1015 99.5127
R2856 vdd.n2411 vdd.n1005 99.5127
R2857 vdd.n2419 vdd.n1005 99.5127
R2858 vdd.n2419 vdd.n1003 99.5127
R2859 vdd.n2423 vdd.n1003 99.5127
R2860 vdd.n2423 vdd.n994 99.5127
R2861 vdd.n2431 vdd.n994 99.5127
R2862 vdd.n2431 vdd.n992 99.5127
R2863 vdd.n2435 vdd.n992 99.5127
R2864 vdd.n2435 vdd.n982 99.5127
R2865 vdd.n2443 vdd.n982 99.5127
R2866 vdd.n2443 vdd.n979 99.5127
R2867 vdd.n2449 vdd.n979 99.5127
R2868 vdd.n2449 vdd.n980 99.5127
R2869 vdd.n980 vdd.n971 99.5127
R2870 vdd.n971 vdd.n962 99.5127
R2871 vdd.n2531 vdd.n962 99.5127
R2872 vdd.n9 vdd.n7 98.9633
R2873 vdd.n2 vdd.n0 98.9633
R2874 vdd.n9 vdd.n8 98.6055
R2875 vdd.n11 vdd.n10 98.6055
R2876 vdd.n13 vdd.n12 98.6055
R2877 vdd.n6 vdd.n5 98.6055
R2878 vdd.n4 vdd.n3 98.6055
R2879 vdd.n2 vdd.n1 98.6055
R2880 vdd.t263 vdd.n303 85.8723
R2881 vdd.t237 vdd.n244 85.8723
R2882 vdd.t251 vdd.n201 85.8723
R2883 vdd.t216 vdd.n142 85.8723
R2884 vdd.t200 vdd.n100 85.8723
R2885 vdd.t138 vdd.n41 85.8723
R2886 vdd.t280 vdd.n1722 85.8723
R2887 vdd.t167 vdd.n1781 85.8723
R2888 vdd.t267 vdd.n1620 85.8723
R2889 vdd.t146 vdd.n1679 85.8723
R2890 vdd.t142 vdd.n1519 85.8723
R2891 vdd.t201 vdd.n1578 85.8723
R2892 vdd.n2923 vdd.n2922 78.546
R2893 vdd.n2397 vdd.n1027 78.546
R2894 vdd.n290 vdd.n289 75.1835
R2895 vdd.n288 vdd.n287 75.1835
R2896 vdd.n286 vdd.n285 75.1835
R2897 vdd.n284 vdd.n283 75.1835
R2898 vdd.n282 vdd.n281 75.1835
R2899 vdd.n280 vdd.n279 75.1835
R2900 vdd.n278 vdd.n277 75.1835
R2901 vdd.n276 vdd.n275 75.1835
R2902 vdd.n274 vdd.n273 75.1835
R2903 vdd.n188 vdd.n187 75.1835
R2904 vdd.n186 vdd.n185 75.1835
R2905 vdd.n184 vdd.n183 75.1835
R2906 vdd.n182 vdd.n181 75.1835
R2907 vdd.n180 vdd.n179 75.1835
R2908 vdd.n178 vdd.n177 75.1835
R2909 vdd.n176 vdd.n175 75.1835
R2910 vdd.n174 vdd.n173 75.1835
R2911 vdd.n172 vdd.n171 75.1835
R2912 vdd.n87 vdd.n86 75.1835
R2913 vdd.n85 vdd.n84 75.1835
R2914 vdd.n83 vdd.n82 75.1835
R2915 vdd.n81 vdd.n80 75.1835
R2916 vdd.n79 vdd.n78 75.1835
R2917 vdd.n77 vdd.n76 75.1835
R2918 vdd.n75 vdd.n74 75.1835
R2919 vdd.n73 vdd.n72 75.1835
R2920 vdd.n71 vdd.n70 75.1835
R2921 vdd.n1752 vdd.n1751 75.1835
R2922 vdd.n1754 vdd.n1753 75.1835
R2923 vdd.n1756 vdd.n1755 75.1835
R2924 vdd.n1758 vdd.n1757 75.1835
R2925 vdd.n1760 vdd.n1759 75.1835
R2926 vdd.n1762 vdd.n1761 75.1835
R2927 vdd.n1764 vdd.n1763 75.1835
R2928 vdd.n1766 vdd.n1765 75.1835
R2929 vdd.n1768 vdd.n1767 75.1835
R2930 vdd.n1650 vdd.n1649 75.1835
R2931 vdd.n1652 vdd.n1651 75.1835
R2932 vdd.n1654 vdd.n1653 75.1835
R2933 vdd.n1656 vdd.n1655 75.1835
R2934 vdd.n1658 vdd.n1657 75.1835
R2935 vdd.n1660 vdd.n1659 75.1835
R2936 vdd.n1662 vdd.n1661 75.1835
R2937 vdd.n1664 vdd.n1663 75.1835
R2938 vdd.n1666 vdd.n1665 75.1835
R2939 vdd.n1549 vdd.n1548 75.1835
R2940 vdd.n1551 vdd.n1550 75.1835
R2941 vdd.n1553 vdd.n1552 75.1835
R2942 vdd.n1555 vdd.n1554 75.1835
R2943 vdd.n1557 vdd.n1556 75.1835
R2944 vdd.n1559 vdd.n1558 75.1835
R2945 vdd.n1561 vdd.n1560 75.1835
R2946 vdd.n1563 vdd.n1562 75.1835
R2947 vdd.n1565 vdd.n1564 75.1835
R2948 vdd.n2858 vdd.n2857 72.8958
R2949 vdd.n2857 vdd.n2621 72.8958
R2950 vdd.n2857 vdd.n2622 72.8958
R2951 vdd.n2857 vdd.n2623 72.8958
R2952 vdd.n2857 vdd.n2624 72.8958
R2953 vdd.n2857 vdd.n2625 72.8958
R2954 vdd.n2857 vdd.n2626 72.8958
R2955 vdd.n2857 vdd.n2627 72.8958
R2956 vdd.n2857 vdd.n2628 72.8958
R2957 vdd.n2857 vdd.n2629 72.8958
R2958 vdd.n2857 vdd.n2630 72.8958
R2959 vdd.n2857 vdd.n2631 72.8958
R2960 vdd.n2857 vdd.n2632 72.8958
R2961 vdd.n2857 vdd.n2633 72.8958
R2962 vdd.n2857 vdd.n2634 72.8958
R2963 vdd.n2857 vdd.n2635 72.8958
R2964 vdd.n2857 vdd.n2636 72.8958
R2965 vdd.n803 vdd.n692 72.8958
R2966 vdd.n3066 vdd.n692 72.8958
R2967 vdd.n797 vdd.n692 72.8958
R2968 vdd.n3073 vdd.n692 72.8958
R2969 vdd.n794 vdd.n692 72.8958
R2970 vdd.n3080 vdd.n692 72.8958
R2971 vdd.n791 vdd.n692 72.8958
R2972 vdd.n3087 vdd.n692 72.8958
R2973 vdd.n3090 vdd.n692 72.8958
R2974 vdd.n2946 vdd.n692 72.8958
R2975 vdd.n2951 vdd.n692 72.8958
R2976 vdd.n2945 vdd.n692 72.8958
R2977 vdd.n2958 vdd.n692 72.8958
R2978 vdd.n2942 vdd.n692 72.8958
R2979 vdd.n2965 vdd.n692 72.8958
R2980 vdd.n2939 vdd.n692 72.8958
R2981 vdd.n2972 vdd.n692 72.8958
R2982 vdd.n2110 vdd.n1049 72.8958
R2983 vdd.n2116 vdd.n1049 72.8958
R2984 vdd.n2118 vdd.n1049 72.8958
R2985 vdd.n2124 vdd.n1049 72.8958
R2986 vdd.n2126 vdd.n1049 72.8958
R2987 vdd.n2132 vdd.n1049 72.8958
R2988 vdd.n2134 vdd.n1049 72.8958
R2989 vdd.n2140 vdd.n1049 72.8958
R2990 vdd.n2311 vdd.n1049 72.8958
R2991 vdd.n2309 vdd.n1049 72.8958
R2992 vdd.n2303 vdd.n1049 72.8958
R2993 vdd.n2301 vdd.n1049 72.8958
R2994 vdd.n2295 vdd.n1049 72.8958
R2995 vdd.n2293 vdd.n1049 72.8958
R2996 vdd.n2287 vdd.n1049 72.8958
R2997 vdd.n2285 vdd.n1049 72.8958
R2998 vdd.n2279 vdd.n1049 72.8958
R2999 vdd.n2604 vdd.n937 72.8958
R3000 vdd.n2604 vdd.n938 72.8958
R3001 vdd.n2604 vdd.n939 72.8958
R3002 vdd.n2604 vdd.n940 72.8958
R3003 vdd.n2604 vdd.n941 72.8958
R3004 vdd.n2604 vdd.n942 72.8958
R3005 vdd.n2604 vdd.n943 72.8958
R3006 vdd.n2604 vdd.n944 72.8958
R3007 vdd.n2604 vdd.n945 72.8958
R3008 vdd.n2604 vdd.n946 72.8958
R3009 vdd.n2604 vdd.n947 72.8958
R3010 vdd.n2604 vdd.n948 72.8958
R3011 vdd.n2604 vdd.n949 72.8958
R3012 vdd.n2604 vdd.n950 72.8958
R3013 vdd.n2604 vdd.n951 72.8958
R3014 vdd.n2604 vdd.n952 72.8958
R3015 vdd.n2604 vdd.n953 72.8958
R3016 vdd.n2857 vdd.n2856 72.8958
R3017 vdd.n2857 vdd.n2605 72.8958
R3018 vdd.n2857 vdd.n2606 72.8958
R3019 vdd.n2857 vdd.n2607 72.8958
R3020 vdd.n2857 vdd.n2608 72.8958
R3021 vdd.n2857 vdd.n2609 72.8958
R3022 vdd.n2857 vdd.n2610 72.8958
R3023 vdd.n2857 vdd.n2611 72.8958
R3024 vdd.n2857 vdd.n2612 72.8958
R3025 vdd.n2857 vdd.n2613 72.8958
R3026 vdd.n2857 vdd.n2614 72.8958
R3027 vdd.n2857 vdd.n2615 72.8958
R3028 vdd.n2857 vdd.n2616 72.8958
R3029 vdd.n2857 vdd.n2617 72.8958
R3030 vdd.n2857 vdd.n2618 72.8958
R3031 vdd.n2857 vdd.n2619 72.8958
R3032 vdd.n2857 vdd.n2620 72.8958
R3033 vdd.n2996 vdd.n692 72.8958
R3034 vdd.n835 vdd.n692 72.8958
R3035 vdd.n3004 vdd.n692 72.8958
R3036 vdd.n830 vdd.n692 72.8958
R3037 vdd.n3011 vdd.n692 72.8958
R3038 vdd.n827 vdd.n692 72.8958
R3039 vdd.n3018 vdd.n692 72.8958
R3040 vdd.n824 vdd.n692 72.8958
R3041 vdd.n3025 vdd.n692 72.8958
R3042 vdd.n3029 vdd.n692 72.8958
R3043 vdd.n821 vdd.n692 72.8958
R3044 vdd.n3036 vdd.n692 72.8958
R3045 vdd.n818 vdd.n692 72.8958
R3046 vdd.n3043 vdd.n692 72.8958
R3047 vdd.n815 vdd.n692 72.8958
R3048 vdd.n3050 vdd.n692 72.8958
R3049 vdd.n3053 vdd.n692 72.8958
R3050 vdd.n2604 vdd.n935 72.8958
R3051 vdd.n2604 vdd.n934 72.8958
R3052 vdd.n2604 vdd.n933 72.8958
R3053 vdd.n2604 vdd.n932 72.8958
R3054 vdd.n2604 vdd.n931 72.8958
R3055 vdd.n2604 vdd.n930 72.8958
R3056 vdd.n2604 vdd.n929 72.8958
R3057 vdd.n2604 vdd.n928 72.8958
R3058 vdd.n2604 vdd.n927 72.8958
R3059 vdd.n2604 vdd.n926 72.8958
R3060 vdd.n2604 vdd.n925 72.8958
R3061 vdd.n2604 vdd.n924 72.8958
R3062 vdd.n2604 vdd.n923 72.8958
R3063 vdd.n2604 vdd.n922 72.8958
R3064 vdd.n2604 vdd.n921 72.8958
R3065 vdd.n2604 vdd.n920 72.8958
R3066 vdd.n2604 vdd.n919 72.8958
R3067 vdd.n2369 vdd.n1049 72.8958
R3068 vdd.n2367 vdd.n1049 72.8958
R3069 vdd.n2361 vdd.n1049 72.8958
R3070 vdd.n2359 vdd.n1049 72.8958
R3071 vdd.n2353 vdd.n1049 72.8958
R3072 vdd.n2351 vdd.n1049 72.8958
R3073 vdd.n2345 vdd.n1049 72.8958
R3074 vdd.n2343 vdd.n1049 72.8958
R3075 vdd.n1061 vdd.n1049 72.8958
R3076 vdd.n2185 vdd.n1049 72.8958
R3077 vdd.n2190 vdd.n1049 72.8958
R3078 vdd.n2192 vdd.n1049 72.8958
R3079 vdd.n2198 vdd.n1049 72.8958
R3080 vdd.n2200 vdd.n1049 72.8958
R3081 vdd.n2206 vdd.n1049 72.8958
R3082 vdd.n2208 vdd.n1049 72.8958
R3083 vdd.n2215 vdd.n1049 72.8958
R3084 vdd.n1419 vdd.n1418 66.2847
R3085 vdd.n1418 vdd.n1194 66.2847
R3086 vdd.n1418 vdd.n1195 66.2847
R3087 vdd.n1418 vdd.n1196 66.2847
R3088 vdd.n1418 vdd.n1197 66.2847
R3089 vdd.n1418 vdd.n1198 66.2847
R3090 vdd.n1418 vdd.n1199 66.2847
R3091 vdd.n1418 vdd.n1200 66.2847
R3092 vdd.n1418 vdd.n1201 66.2847
R3093 vdd.n1418 vdd.n1202 66.2847
R3094 vdd.n1418 vdd.n1203 66.2847
R3095 vdd.n1418 vdd.n1204 66.2847
R3096 vdd.n1418 vdd.n1205 66.2847
R3097 vdd.n1418 vdd.n1206 66.2847
R3098 vdd.n1418 vdd.n1207 66.2847
R3099 vdd.n1418 vdd.n1208 66.2847
R3100 vdd.n1418 vdd.n1209 66.2847
R3101 vdd.n1418 vdd.n1210 66.2847
R3102 vdd.n1418 vdd.n1211 66.2847
R3103 vdd.n1418 vdd.n1212 66.2847
R3104 vdd.n1418 vdd.n1213 66.2847
R3105 vdd.n1418 vdd.n1214 66.2847
R3106 vdd.n1418 vdd.n1215 66.2847
R3107 vdd.n1418 vdd.n1216 66.2847
R3108 vdd.n1418 vdd.n1217 66.2847
R3109 vdd.n1418 vdd.n1218 66.2847
R3110 vdd.n1418 vdd.n1219 66.2847
R3111 vdd.n1418 vdd.n1220 66.2847
R3112 vdd.n1418 vdd.n1221 66.2847
R3113 vdd.n1418 vdd.n1222 66.2847
R3114 vdd.n1418 vdd.n1223 66.2847
R3115 vdd.n1073 vdd.n1070 66.2847
R3116 vdd.n2000 vdd.n1073 66.2847
R3117 vdd.n2005 vdd.n1073 66.2847
R3118 vdd.n2010 vdd.n1073 66.2847
R3119 vdd.n1998 vdd.n1073 66.2847
R3120 vdd.n2017 vdd.n1073 66.2847
R3121 vdd.n1990 vdd.n1073 66.2847
R3122 vdd.n2024 vdd.n1073 66.2847
R3123 vdd.n1983 vdd.n1073 66.2847
R3124 vdd.n2031 vdd.n1073 66.2847
R3125 vdd.n1977 vdd.n1073 66.2847
R3126 vdd.n1972 vdd.n1073 66.2847
R3127 vdd.n2042 vdd.n1073 66.2847
R3128 vdd.n1964 vdd.n1073 66.2847
R3129 vdd.n2049 vdd.n1073 66.2847
R3130 vdd.n1957 vdd.n1073 66.2847
R3131 vdd.n2056 vdd.n1073 66.2847
R3132 vdd.n1950 vdd.n1073 66.2847
R3133 vdd.n2063 vdd.n1073 66.2847
R3134 vdd.n1943 vdd.n1073 66.2847
R3135 vdd.n2070 vdd.n1073 66.2847
R3136 vdd.n1937 vdd.n1073 66.2847
R3137 vdd.n1932 vdd.n1073 66.2847
R3138 vdd.n2081 vdd.n1073 66.2847
R3139 vdd.n1924 vdd.n1073 66.2847
R3140 vdd.n2088 vdd.n1073 66.2847
R3141 vdd.n1917 vdd.n1073 66.2847
R3142 vdd.n2095 vdd.n1073 66.2847
R3143 vdd.n2098 vdd.n1073 66.2847
R3144 vdd.n1908 vdd.n1073 66.2847
R3145 vdd.n2320 vdd.n1073 66.2847
R3146 vdd.n1902 vdd.n1073 66.2847
R3147 vdd.n3223 vdd.n3222 66.2847
R3148 vdd.n3223 vdd.n693 66.2847
R3149 vdd.n3223 vdd.n694 66.2847
R3150 vdd.n3223 vdd.n695 66.2847
R3151 vdd.n3223 vdd.n696 66.2847
R3152 vdd.n3223 vdd.n697 66.2847
R3153 vdd.n3223 vdd.n698 66.2847
R3154 vdd.n3223 vdd.n699 66.2847
R3155 vdd.n3223 vdd.n700 66.2847
R3156 vdd.n3223 vdd.n701 66.2847
R3157 vdd.n3223 vdd.n702 66.2847
R3158 vdd.n3223 vdd.n703 66.2847
R3159 vdd.n3223 vdd.n704 66.2847
R3160 vdd.n3223 vdd.n705 66.2847
R3161 vdd.n3223 vdd.n706 66.2847
R3162 vdd.n3223 vdd.n707 66.2847
R3163 vdd.n3223 vdd.n708 66.2847
R3164 vdd.n3223 vdd.n709 66.2847
R3165 vdd.n3223 vdd.n710 66.2847
R3166 vdd.n3223 vdd.n711 66.2847
R3167 vdd.n3223 vdd.n712 66.2847
R3168 vdd.n3223 vdd.n713 66.2847
R3169 vdd.n3223 vdd.n714 66.2847
R3170 vdd.n3223 vdd.n715 66.2847
R3171 vdd.n3223 vdd.n716 66.2847
R3172 vdd.n3223 vdd.n717 66.2847
R3173 vdd.n3223 vdd.n718 66.2847
R3174 vdd.n3223 vdd.n719 66.2847
R3175 vdd.n3223 vdd.n720 66.2847
R3176 vdd.n3223 vdd.n721 66.2847
R3177 vdd.n3223 vdd.n722 66.2847
R3178 vdd.n3354 vdd.n3353 66.2847
R3179 vdd.n3354 vdd.n424 66.2847
R3180 vdd.n3354 vdd.n423 66.2847
R3181 vdd.n3354 vdd.n422 66.2847
R3182 vdd.n3354 vdd.n421 66.2847
R3183 vdd.n3354 vdd.n420 66.2847
R3184 vdd.n3354 vdd.n419 66.2847
R3185 vdd.n3354 vdd.n418 66.2847
R3186 vdd.n3354 vdd.n417 66.2847
R3187 vdd.n3354 vdd.n416 66.2847
R3188 vdd.n3354 vdd.n415 66.2847
R3189 vdd.n3354 vdd.n414 66.2847
R3190 vdd.n3354 vdd.n413 66.2847
R3191 vdd.n3354 vdd.n412 66.2847
R3192 vdd.n3354 vdd.n411 66.2847
R3193 vdd.n3354 vdd.n410 66.2847
R3194 vdd.n3354 vdd.n409 66.2847
R3195 vdd.n3354 vdd.n408 66.2847
R3196 vdd.n3354 vdd.n407 66.2847
R3197 vdd.n3354 vdd.n406 66.2847
R3198 vdd.n3354 vdd.n405 66.2847
R3199 vdd.n3354 vdd.n404 66.2847
R3200 vdd.n3354 vdd.n403 66.2847
R3201 vdd.n3354 vdd.n402 66.2847
R3202 vdd.n3354 vdd.n401 66.2847
R3203 vdd.n3354 vdd.n400 66.2847
R3204 vdd.n3354 vdd.n399 66.2847
R3205 vdd.n3354 vdd.n398 66.2847
R3206 vdd.n3354 vdd.n397 66.2847
R3207 vdd.n3354 vdd.n396 66.2847
R3208 vdd.n3354 vdd.n395 66.2847
R3209 vdd.n3354 vdd.n394 66.2847
R3210 vdd.n467 vdd.n394 52.4337
R3211 vdd.n473 vdd.n395 52.4337
R3212 vdd.n477 vdd.n396 52.4337
R3213 vdd.n483 vdd.n397 52.4337
R3214 vdd.n487 vdd.n398 52.4337
R3215 vdd.n493 vdd.n399 52.4337
R3216 vdd.n497 vdd.n400 52.4337
R3217 vdd.n503 vdd.n401 52.4337
R3218 vdd.n507 vdd.n402 52.4337
R3219 vdd.n513 vdd.n403 52.4337
R3220 vdd.n517 vdd.n404 52.4337
R3221 vdd.n523 vdd.n405 52.4337
R3222 vdd.n527 vdd.n406 52.4337
R3223 vdd.n533 vdd.n407 52.4337
R3224 vdd.n537 vdd.n408 52.4337
R3225 vdd.n543 vdd.n409 52.4337
R3226 vdd.n547 vdd.n410 52.4337
R3227 vdd.n553 vdd.n411 52.4337
R3228 vdd.n557 vdd.n412 52.4337
R3229 vdd.n563 vdd.n413 52.4337
R3230 vdd.n567 vdd.n414 52.4337
R3231 vdd.n573 vdd.n415 52.4337
R3232 vdd.n577 vdd.n416 52.4337
R3233 vdd.n583 vdd.n417 52.4337
R3234 vdd.n587 vdd.n418 52.4337
R3235 vdd.n593 vdd.n419 52.4337
R3236 vdd.n597 vdd.n420 52.4337
R3237 vdd.n603 vdd.n421 52.4337
R3238 vdd.n607 vdd.n422 52.4337
R3239 vdd.n613 vdd.n423 52.4337
R3240 vdd.n616 vdd.n424 52.4337
R3241 vdd.n3353 vdd.n3352 52.4337
R3242 vdd.n3222 vdd.n3221 52.4337
R3243 vdd.n728 vdd.n693 52.4337
R3244 vdd.n734 vdd.n694 52.4337
R3245 vdd.n3211 vdd.n695 52.4337
R3246 vdd.n3207 vdd.n696 52.4337
R3247 vdd.n3203 vdd.n697 52.4337
R3248 vdd.n3199 vdd.n698 52.4337
R3249 vdd.n3195 vdd.n699 52.4337
R3250 vdd.n3191 vdd.n700 52.4337
R3251 vdd.n3187 vdd.n701 52.4337
R3252 vdd.n3179 vdd.n702 52.4337
R3253 vdd.n3175 vdd.n703 52.4337
R3254 vdd.n3171 vdd.n704 52.4337
R3255 vdd.n3167 vdd.n705 52.4337
R3256 vdd.n3163 vdd.n706 52.4337
R3257 vdd.n3159 vdd.n707 52.4337
R3258 vdd.n3155 vdd.n708 52.4337
R3259 vdd.n3151 vdd.n709 52.4337
R3260 vdd.n3147 vdd.n710 52.4337
R3261 vdd.n3143 vdd.n711 52.4337
R3262 vdd.n3139 vdd.n712 52.4337
R3263 vdd.n3133 vdd.n713 52.4337
R3264 vdd.n3129 vdd.n714 52.4337
R3265 vdd.n3125 vdd.n715 52.4337
R3266 vdd.n3121 vdd.n716 52.4337
R3267 vdd.n3117 vdd.n717 52.4337
R3268 vdd.n3113 vdd.n718 52.4337
R3269 vdd.n3109 vdd.n719 52.4337
R3270 vdd.n3105 vdd.n720 52.4337
R3271 vdd.n3101 vdd.n721 52.4337
R3272 vdd.n3097 vdd.n722 52.4337
R3273 vdd.n2322 vdd.n1902 52.4337
R3274 vdd.n2320 vdd.n2319 52.4337
R3275 vdd.n1909 vdd.n1908 52.4337
R3276 vdd.n2098 vdd.n2097 52.4337
R3277 vdd.n2095 vdd.n2094 52.4337
R3278 vdd.n2090 vdd.n1917 52.4337
R3279 vdd.n2088 vdd.n2087 52.4337
R3280 vdd.n2083 vdd.n1924 52.4337
R3281 vdd.n2081 vdd.n2080 52.4337
R3282 vdd.n1933 vdd.n1932 52.4337
R3283 vdd.n2072 vdd.n1937 52.4337
R3284 vdd.n2070 vdd.n2069 52.4337
R3285 vdd.n2065 vdd.n1943 52.4337
R3286 vdd.n2063 vdd.n2062 52.4337
R3287 vdd.n2058 vdd.n1950 52.4337
R3288 vdd.n2056 vdd.n2055 52.4337
R3289 vdd.n2051 vdd.n1957 52.4337
R3290 vdd.n2049 vdd.n2048 52.4337
R3291 vdd.n2044 vdd.n1964 52.4337
R3292 vdd.n2042 vdd.n2041 52.4337
R3293 vdd.n1973 vdd.n1972 52.4337
R3294 vdd.n2033 vdd.n1977 52.4337
R3295 vdd.n2031 vdd.n2030 52.4337
R3296 vdd.n2026 vdd.n1983 52.4337
R3297 vdd.n2024 vdd.n2023 52.4337
R3298 vdd.n2019 vdd.n1990 52.4337
R3299 vdd.n2017 vdd.n2016 52.4337
R3300 vdd.n2012 vdd.n1998 52.4337
R3301 vdd.n2010 vdd.n2009 52.4337
R3302 vdd.n2005 vdd.n2004 52.4337
R3303 vdd.n2000 vdd.n1999 52.4337
R3304 vdd.n2331 vdd.n1070 52.4337
R3305 vdd.n1420 vdd.n1419 52.4337
R3306 vdd.n1226 vdd.n1194 52.4337
R3307 vdd.n1230 vdd.n1195 52.4337
R3308 vdd.n1232 vdd.n1196 52.4337
R3309 vdd.n1236 vdd.n1197 52.4337
R3310 vdd.n1238 vdd.n1198 52.4337
R3311 vdd.n1242 vdd.n1199 52.4337
R3312 vdd.n1244 vdd.n1200 52.4337
R3313 vdd.n1248 vdd.n1201 52.4337
R3314 vdd.n1250 vdd.n1202 52.4337
R3315 vdd.n1256 vdd.n1203 52.4337
R3316 vdd.n1258 vdd.n1204 52.4337
R3317 vdd.n1262 vdd.n1205 52.4337
R3318 vdd.n1264 vdd.n1206 52.4337
R3319 vdd.n1268 vdd.n1207 52.4337
R3320 vdd.n1270 vdd.n1208 52.4337
R3321 vdd.n1274 vdd.n1209 52.4337
R3322 vdd.n1276 vdd.n1210 52.4337
R3323 vdd.n1280 vdd.n1211 52.4337
R3324 vdd.n1282 vdd.n1212 52.4337
R3325 vdd.n1354 vdd.n1213 52.4337
R3326 vdd.n1287 vdd.n1214 52.4337
R3327 vdd.n1291 vdd.n1215 52.4337
R3328 vdd.n1293 vdd.n1216 52.4337
R3329 vdd.n1297 vdd.n1217 52.4337
R3330 vdd.n1299 vdd.n1218 52.4337
R3331 vdd.n1303 vdd.n1219 52.4337
R3332 vdd.n1305 vdd.n1220 52.4337
R3333 vdd.n1309 vdd.n1221 52.4337
R3334 vdd.n1311 vdd.n1222 52.4337
R3335 vdd.n1315 vdd.n1223 52.4337
R3336 vdd.n1419 vdd.n1193 52.4337
R3337 vdd.n1229 vdd.n1194 52.4337
R3338 vdd.n1231 vdd.n1195 52.4337
R3339 vdd.n1235 vdd.n1196 52.4337
R3340 vdd.n1237 vdd.n1197 52.4337
R3341 vdd.n1241 vdd.n1198 52.4337
R3342 vdd.n1243 vdd.n1199 52.4337
R3343 vdd.n1247 vdd.n1200 52.4337
R3344 vdd.n1249 vdd.n1201 52.4337
R3345 vdd.n1255 vdd.n1202 52.4337
R3346 vdd.n1257 vdd.n1203 52.4337
R3347 vdd.n1261 vdd.n1204 52.4337
R3348 vdd.n1263 vdd.n1205 52.4337
R3349 vdd.n1267 vdd.n1206 52.4337
R3350 vdd.n1269 vdd.n1207 52.4337
R3351 vdd.n1273 vdd.n1208 52.4337
R3352 vdd.n1275 vdd.n1209 52.4337
R3353 vdd.n1279 vdd.n1210 52.4337
R3354 vdd.n1281 vdd.n1211 52.4337
R3355 vdd.n1285 vdd.n1212 52.4337
R3356 vdd.n1286 vdd.n1213 52.4337
R3357 vdd.n1290 vdd.n1214 52.4337
R3358 vdd.n1292 vdd.n1215 52.4337
R3359 vdd.n1296 vdd.n1216 52.4337
R3360 vdd.n1298 vdd.n1217 52.4337
R3361 vdd.n1302 vdd.n1218 52.4337
R3362 vdd.n1304 vdd.n1219 52.4337
R3363 vdd.n1308 vdd.n1220 52.4337
R3364 vdd.n1310 vdd.n1221 52.4337
R3365 vdd.n1314 vdd.n1222 52.4337
R3366 vdd.n1316 vdd.n1223 52.4337
R3367 vdd.n1070 vdd.n1069 52.4337
R3368 vdd.n2001 vdd.n2000 52.4337
R3369 vdd.n2006 vdd.n2005 52.4337
R3370 vdd.n2011 vdd.n2010 52.4337
R3371 vdd.n1998 vdd.n1991 52.4337
R3372 vdd.n2018 vdd.n2017 52.4337
R3373 vdd.n1990 vdd.n1984 52.4337
R3374 vdd.n2025 vdd.n2024 52.4337
R3375 vdd.n1983 vdd.n1978 52.4337
R3376 vdd.n2032 vdd.n2031 52.4337
R3377 vdd.n1977 vdd.n1976 52.4337
R3378 vdd.n1972 vdd.n1965 52.4337
R3379 vdd.n2043 vdd.n2042 52.4337
R3380 vdd.n1964 vdd.n1958 52.4337
R3381 vdd.n2050 vdd.n2049 52.4337
R3382 vdd.n1957 vdd.n1951 52.4337
R3383 vdd.n2057 vdd.n2056 52.4337
R3384 vdd.n1950 vdd.n1944 52.4337
R3385 vdd.n2064 vdd.n2063 52.4337
R3386 vdd.n1943 vdd.n1938 52.4337
R3387 vdd.n2071 vdd.n2070 52.4337
R3388 vdd.n1937 vdd.n1936 52.4337
R3389 vdd.n1932 vdd.n1925 52.4337
R3390 vdd.n2082 vdd.n2081 52.4337
R3391 vdd.n1924 vdd.n1918 52.4337
R3392 vdd.n2089 vdd.n2088 52.4337
R3393 vdd.n1917 vdd.n1911 52.4337
R3394 vdd.n2096 vdd.n2095 52.4337
R3395 vdd.n2099 vdd.n2098 52.4337
R3396 vdd.n1908 vdd.n1903 52.4337
R3397 vdd.n2321 vdd.n2320 52.4337
R3398 vdd.n1902 vdd.n1075 52.4337
R3399 vdd.n3222 vdd.n725 52.4337
R3400 vdd.n733 vdd.n693 52.4337
R3401 vdd.n3212 vdd.n694 52.4337
R3402 vdd.n3208 vdd.n695 52.4337
R3403 vdd.n3204 vdd.n696 52.4337
R3404 vdd.n3200 vdd.n697 52.4337
R3405 vdd.n3196 vdd.n698 52.4337
R3406 vdd.n3192 vdd.n699 52.4337
R3407 vdd.n3188 vdd.n700 52.4337
R3408 vdd.n3178 vdd.n701 52.4337
R3409 vdd.n3176 vdd.n702 52.4337
R3410 vdd.n3172 vdd.n703 52.4337
R3411 vdd.n3168 vdd.n704 52.4337
R3412 vdd.n3164 vdd.n705 52.4337
R3413 vdd.n3160 vdd.n706 52.4337
R3414 vdd.n3156 vdd.n707 52.4337
R3415 vdd.n3152 vdd.n708 52.4337
R3416 vdd.n3148 vdd.n709 52.4337
R3417 vdd.n3144 vdd.n710 52.4337
R3418 vdd.n3140 vdd.n711 52.4337
R3419 vdd.n3132 vdd.n712 52.4337
R3420 vdd.n3130 vdd.n713 52.4337
R3421 vdd.n3126 vdd.n714 52.4337
R3422 vdd.n3122 vdd.n715 52.4337
R3423 vdd.n3118 vdd.n716 52.4337
R3424 vdd.n3114 vdd.n717 52.4337
R3425 vdd.n3110 vdd.n718 52.4337
R3426 vdd.n3106 vdd.n719 52.4337
R3427 vdd.n3102 vdd.n720 52.4337
R3428 vdd.n3098 vdd.n721 52.4337
R3429 vdd.n722 vdd.n691 52.4337
R3430 vdd.n3353 vdd.n425 52.4337
R3431 vdd.n614 vdd.n424 52.4337
R3432 vdd.n608 vdd.n423 52.4337
R3433 vdd.n604 vdd.n422 52.4337
R3434 vdd.n598 vdd.n421 52.4337
R3435 vdd.n594 vdd.n420 52.4337
R3436 vdd.n588 vdd.n419 52.4337
R3437 vdd.n584 vdd.n418 52.4337
R3438 vdd.n578 vdd.n417 52.4337
R3439 vdd.n574 vdd.n416 52.4337
R3440 vdd.n568 vdd.n415 52.4337
R3441 vdd.n564 vdd.n414 52.4337
R3442 vdd.n558 vdd.n413 52.4337
R3443 vdd.n554 vdd.n412 52.4337
R3444 vdd.n548 vdd.n411 52.4337
R3445 vdd.n544 vdd.n410 52.4337
R3446 vdd.n538 vdd.n409 52.4337
R3447 vdd.n534 vdd.n408 52.4337
R3448 vdd.n528 vdd.n407 52.4337
R3449 vdd.n524 vdd.n406 52.4337
R3450 vdd.n518 vdd.n405 52.4337
R3451 vdd.n514 vdd.n404 52.4337
R3452 vdd.n508 vdd.n403 52.4337
R3453 vdd.n504 vdd.n402 52.4337
R3454 vdd.n498 vdd.n401 52.4337
R3455 vdd.n494 vdd.n400 52.4337
R3456 vdd.n488 vdd.n399 52.4337
R3457 vdd.n484 vdd.n398 52.4337
R3458 vdd.n478 vdd.n397 52.4337
R3459 vdd.n474 vdd.n396 52.4337
R3460 vdd.n468 vdd.n395 52.4337
R3461 vdd.n394 vdd.n392 52.4337
R3462 vdd.t115 vdd.t87 51.4683
R3463 vdd.n274 vdd.n272 42.0461
R3464 vdd.n172 vdd.n170 42.0461
R3465 vdd.n71 vdd.n69 42.0461
R3466 vdd.n1752 vdd.n1750 42.0461
R3467 vdd.n1650 vdd.n1648 42.0461
R3468 vdd.n1549 vdd.n1547 42.0461
R3469 vdd.n332 vdd.n331 41.6884
R3470 vdd.n230 vdd.n229 41.6884
R3471 vdd.n129 vdd.n128 41.6884
R3472 vdd.n1810 vdd.n1809 41.6884
R3473 vdd.n1708 vdd.n1707 41.6884
R3474 vdd.n1607 vdd.n1606 41.6884
R3475 vdd.n1319 vdd.n1318 41.1157
R3476 vdd.n1357 vdd.n1356 41.1157
R3477 vdd.n1253 vdd.n1252 41.1157
R3478 vdd.n428 vdd.n427 41.1157
R3479 vdd.n566 vdd.n441 41.1157
R3480 vdd.n454 vdd.n453 41.1157
R3481 vdd.n3053 vdd.n3052 39.2114
R3482 vdd.n3050 vdd.n3049 39.2114
R3483 vdd.n3045 vdd.n815 39.2114
R3484 vdd.n3043 vdd.n3042 39.2114
R3485 vdd.n3038 vdd.n818 39.2114
R3486 vdd.n3036 vdd.n3035 39.2114
R3487 vdd.n3031 vdd.n821 39.2114
R3488 vdd.n3029 vdd.n3028 39.2114
R3489 vdd.n3025 vdd.n3024 39.2114
R3490 vdd.n3020 vdd.n824 39.2114
R3491 vdd.n3018 vdd.n3017 39.2114
R3492 vdd.n3013 vdd.n827 39.2114
R3493 vdd.n3011 vdd.n3010 39.2114
R3494 vdd.n3006 vdd.n830 39.2114
R3495 vdd.n3004 vdd.n3003 39.2114
R3496 vdd.n2998 vdd.n835 39.2114
R3497 vdd.n2996 vdd.n2995 39.2114
R3498 vdd.n2856 vdd.n913 39.2114
R3499 vdd.n2851 vdd.n2605 39.2114
R3500 vdd.n2848 vdd.n2606 39.2114
R3501 vdd.n2844 vdd.n2607 39.2114
R3502 vdd.n2840 vdd.n2608 39.2114
R3503 vdd.n2836 vdd.n2609 39.2114
R3504 vdd.n2832 vdd.n2610 39.2114
R3505 vdd.n2828 vdd.n2611 39.2114
R3506 vdd.n2824 vdd.n2612 39.2114
R3507 vdd.n2820 vdd.n2613 39.2114
R3508 vdd.n2816 vdd.n2614 39.2114
R3509 vdd.n2812 vdd.n2615 39.2114
R3510 vdd.n2808 vdd.n2616 39.2114
R3511 vdd.n2804 vdd.n2617 39.2114
R3512 vdd.n2800 vdd.n2618 39.2114
R3513 vdd.n2796 vdd.n2619 39.2114
R3514 vdd.n2791 vdd.n2620 39.2114
R3515 vdd.n2599 vdd.n953 39.2114
R3516 vdd.n2595 vdd.n952 39.2114
R3517 vdd.n2591 vdd.n951 39.2114
R3518 vdd.n2587 vdd.n950 39.2114
R3519 vdd.n2583 vdd.n949 39.2114
R3520 vdd.n2579 vdd.n948 39.2114
R3521 vdd.n2575 vdd.n947 39.2114
R3522 vdd.n2571 vdd.n946 39.2114
R3523 vdd.n2567 vdd.n945 39.2114
R3524 vdd.n2563 vdd.n944 39.2114
R3525 vdd.n2559 vdd.n943 39.2114
R3526 vdd.n2555 vdd.n942 39.2114
R3527 vdd.n2551 vdd.n941 39.2114
R3528 vdd.n2547 vdd.n940 39.2114
R3529 vdd.n2543 vdd.n939 39.2114
R3530 vdd.n2538 vdd.n938 39.2114
R3531 vdd.n2534 vdd.n937 39.2114
R3532 vdd.n2110 vdd.n1048 39.2114
R3533 vdd.n2116 vdd.n2115 39.2114
R3534 vdd.n2119 vdd.n2118 39.2114
R3535 vdd.n2124 vdd.n2123 39.2114
R3536 vdd.n2127 vdd.n2126 39.2114
R3537 vdd.n2132 vdd.n2131 39.2114
R3538 vdd.n2135 vdd.n2134 39.2114
R3539 vdd.n2140 vdd.n2139 39.2114
R3540 vdd.n2311 vdd.n2142 39.2114
R3541 vdd.n2310 vdd.n2309 39.2114
R3542 vdd.n2303 vdd.n2144 39.2114
R3543 vdd.n2302 vdd.n2301 39.2114
R3544 vdd.n2295 vdd.n2146 39.2114
R3545 vdd.n2294 vdd.n2293 39.2114
R3546 vdd.n2287 vdd.n2148 39.2114
R3547 vdd.n2286 vdd.n2285 39.2114
R3548 vdd.n2279 vdd.n2150 39.2114
R3549 vdd.n2972 vdd.n2971 39.2114
R3550 vdd.n2967 vdd.n2939 39.2114
R3551 vdd.n2965 vdd.n2964 39.2114
R3552 vdd.n2960 vdd.n2942 39.2114
R3553 vdd.n2958 vdd.n2957 39.2114
R3554 vdd.n2953 vdd.n2945 39.2114
R3555 vdd.n2951 vdd.n2950 39.2114
R3556 vdd.n2946 vdd.n787 39.2114
R3557 vdd.n3090 vdd.n3089 39.2114
R3558 vdd.n3087 vdd.n3086 39.2114
R3559 vdd.n3082 vdd.n791 39.2114
R3560 vdd.n3080 vdd.n3079 39.2114
R3561 vdd.n3075 vdd.n794 39.2114
R3562 vdd.n3073 vdd.n3072 39.2114
R3563 vdd.n3068 vdd.n797 39.2114
R3564 vdd.n3066 vdd.n3065 39.2114
R3565 vdd.n3061 vdd.n803 39.2114
R3566 vdd.n2858 vdd.n916 39.2114
R3567 vdd.n2621 vdd.n918 39.2114
R3568 vdd.n2647 vdd.n2622 39.2114
R3569 vdd.n2651 vdd.n2623 39.2114
R3570 vdd.n2655 vdd.n2624 39.2114
R3571 vdd.n2659 vdd.n2625 39.2114
R3572 vdd.n2663 vdd.n2626 39.2114
R3573 vdd.n2667 vdd.n2627 39.2114
R3574 vdd.n2671 vdd.n2628 39.2114
R3575 vdd.n2675 vdd.n2629 39.2114
R3576 vdd.n2679 vdd.n2630 39.2114
R3577 vdd.n2683 vdd.n2631 39.2114
R3578 vdd.n2687 vdd.n2632 39.2114
R3579 vdd.n2691 vdd.n2633 39.2114
R3580 vdd.n2695 vdd.n2634 39.2114
R3581 vdd.n2699 vdd.n2635 39.2114
R3582 vdd.n2703 vdd.n2636 39.2114
R3583 vdd.n2859 vdd.n2858 39.2114
R3584 vdd.n2646 vdd.n2621 39.2114
R3585 vdd.n2650 vdd.n2622 39.2114
R3586 vdd.n2654 vdd.n2623 39.2114
R3587 vdd.n2658 vdd.n2624 39.2114
R3588 vdd.n2662 vdd.n2625 39.2114
R3589 vdd.n2666 vdd.n2626 39.2114
R3590 vdd.n2670 vdd.n2627 39.2114
R3591 vdd.n2674 vdd.n2628 39.2114
R3592 vdd.n2678 vdd.n2629 39.2114
R3593 vdd.n2682 vdd.n2630 39.2114
R3594 vdd.n2686 vdd.n2631 39.2114
R3595 vdd.n2690 vdd.n2632 39.2114
R3596 vdd.n2694 vdd.n2633 39.2114
R3597 vdd.n2698 vdd.n2634 39.2114
R3598 vdd.n2702 vdd.n2635 39.2114
R3599 vdd.n2705 vdd.n2636 39.2114
R3600 vdd.n803 vdd.n798 39.2114
R3601 vdd.n3067 vdd.n3066 39.2114
R3602 vdd.n797 vdd.n795 39.2114
R3603 vdd.n3074 vdd.n3073 39.2114
R3604 vdd.n794 vdd.n792 39.2114
R3605 vdd.n3081 vdd.n3080 39.2114
R3606 vdd.n791 vdd.n789 39.2114
R3607 vdd.n3088 vdd.n3087 39.2114
R3608 vdd.n3091 vdd.n3090 39.2114
R3609 vdd.n2947 vdd.n2946 39.2114
R3610 vdd.n2952 vdd.n2951 39.2114
R3611 vdd.n2945 vdd.n2943 39.2114
R3612 vdd.n2959 vdd.n2958 39.2114
R3613 vdd.n2942 vdd.n2940 39.2114
R3614 vdd.n2966 vdd.n2965 39.2114
R3615 vdd.n2939 vdd.n2937 39.2114
R3616 vdd.n2973 vdd.n2972 39.2114
R3617 vdd.n2111 vdd.n2110 39.2114
R3618 vdd.n2117 vdd.n2116 39.2114
R3619 vdd.n2118 vdd.n2107 39.2114
R3620 vdd.n2125 vdd.n2124 39.2114
R3621 vdd.n2126 vdd.n2105 39.2114
R3622 vdd.n2133 vdd.n2132 39.2114
R3623 vdd.n2134 vdd.n2103 39.2114
R3624 vdd.n2141 vdd.n2140 39.2114
R3625 vdd.n2312 vdd.n2311 39.2114
R3626 vdd.n2309 vdd.n2308 39.2114
R3627 vdd.n2304 vdd.n2303 39.2114
R3628 vdd.n2301 vdd.n2300 39.2114
R3629 vdd.n2296 vdd.n2295 39.2114
R3630 vdd.n2293 vdd.n2292 39.2114
R3631 vdd.n2288 vdd.n2287 39.2114
R3632 vdd.n2285 vdd.n2284 39.2114
R3633 vdd.n2280 vdd.n2279 39.2114
R3634 vdd.n2537 vdd.n937 39.2114
R3635 vdd.n2542 vdd.n938 39.2114
R3636 vdd.n2546 vdd.n939 39.2114
R3637 vdd.n2550 vdd.n940 39.2114
R3638 vdd.n2554 vdd.n941 39.2114
R3639 vdd.n2558 vdd.n942 39.2114
R3640 vdd.n2562 vdd.n943 39.2114
R3641 vdd.n2566 vdd.n944 39.2114
R3642 vdd.n2570 vdd.n945 39.2114
R3643 vdd.n2574 vdd.n946 39.2114
R3644 vdd.n2578 vdd.n947 39.2114
R3645 vdd.n2582 vdd.n948 39.2114
R3646 vdd.n2586 vdd.n949 39.2114
R3647 vdd.n2590 vdd.n950 39.2114
R3648 vdd.n2594 vdd.n951 39.2114
R3649 vdd.n2598 vdd.n952 39.2114
R3650 vdd.n955 vdd.n953 39.2114
R3651 vdd.n2856 vdd.n2855 39.2114
R3652 vdd.n2849 vdd.n2605 39.2114
R3653 vdd.n2845 vdd.n2606 39.2114
R3654 vdd.n2841 vdd.n2607 39.2114
R3655 vdd.n2837 vdd.n2608 39.2114
R3656 vdd.n2833 vdd.n2609 39.2114
R3657 vdd.n2829 vdd.n2610 39.2114
R3658 vdd.n2825 vdd.n2611 39.2114
R3659 vdd.n2821 vdd.n2612 39.2114
R3660 vdd.n2817 vdd.n2613 39.2114
R3661 vdd.n2813 vdd.n2614 39.2114
R3662 vdd.n2809 vdd.n2615 39.2114
R3663 vdd.n2805 vdd.n2616 39.2114
R3664 vdd.n2801 vdd.n2617 39.2114
R3665 vdd.n2797 vdd.n2618 39.2114
R3666 vdd.n2792 vdd.n2619 39.2114
R3667 vdd.n2788 vdd.n2620 39.2114
R3668 vdd.n2997 vdd.n2996 39.2114
R3669 vdd.n835 vdd.n831 39.2114
R3670 vdd.n3005 vdd.n3004 39.2114
R3671 vdd.n830 vdd.n828 39.2114
R3672 vdd.n3012 vdd.n3011 39.2114
R3673 vdd.n827 vdd.n825 39.2114
R3674 vdd.n3019 vdd.n3018 39.2114
R3675 vdd.n824 vdd.n822 39.2114
R3676 vdd.n3026 vdd.n3025 39.2114
R3677 vdd.n3030 vdd.n3029 39.2114
R3678 vdd.n821 vdd.n819 39.2114
R3679 vdd.n3037 vdd.n3036 39.2114
R3680 vdd.n818 vdd.n816 39.2114
R3681 vdd.n3044 vdd.n3043 39.2114
R3682 vdd.n815 vdd.n813 39.2114
R3683 vdd.n3051 vdd.n3050 39.2114
R3684 vdd.n3054 vdd.n3053 39.2114
R3685 vdd.n963 vdd.n919 39.2114
R3686 vdd.n2526 vdd.n920 39.2114
R3687 vdd.n2522 vdd.n921 39.2114
R3688 vdd.n2518 vdd.n922 39.2114
R3689 vdd.n2514 vdd.n923 39.2114
R3690 vdd.n2510 vdd.n924 39.2114
R3691 vdd.n2506 vdd.n925 39.2114
R3692 vdd.n2502 vdd.n926 39.2114
R3693 vdd.n2498 vdd.n927 39.2114
R3694 vdd.n2494 vdd.n928 39.2114
R3695 vdd.n2490 vdd.n929 39.2114
R3696 vdd.n2486 vdd.n930 39.2114
R3697 vdd.n2482 vdd.n931 39.2114
R3698 vdd.n2478 vdd.n932 39.2114
R3699 vdd.n2474 vdd.n933 39.2114
R3700 vdd.n2470 vdd.n934 39.2114
R3701 vdd.n2466 vdd.n935 39.2114
R3702 vdd.n2369 vdd.n1052 39.2114
R3703 vdd.n2368 vdd.n2367 39.2114
R3704 vdd.n2361 vdd.n1054 39.2114
R3705 vdd.n2360 vdd.n2359 39.2114
R3706 vdd.n2353 vdd.n1056 39.2114
R3707 vdd.n2352 vdd.n2351 39.2114
R3708 vdd.n2345 vdd.n1058 39.2114
R3709 vdd.n2344 vdd.n2343 39.2114
R3710 vdd.n1061 vdd.n1060 39.2114
R3711 vdd.n2185 vdd.n2184 39.2114
R3712 vdd.n2190 vdd.n2189 39.2114
R3713 vdd.n2193 vdd.n2192 39.2114
R3714 vdd.n2198 vdd.n2197 39.2114
R3715 vdd.n2201 vdd.n2200 39.2114
R3716 vdd.n2206 vdd.n2205 39.2114
R3717 vdd.n2209 vdd.n2208 39.2114
R3718 vdd.n2215 vdd.n2214 39.2114
R3719 vdd.n2463 vdd.n935 39.2114
R3720 vdd.n2467 vdd.n934 39.2114
R3721 vdd.n2471 vdd.n933 39.2114
R3722 vdd.n2475 vdd.n932 39.2114
R3723 vdd.n2479 vdd.n931 39.2114
R3724 vdd.n2483 vdd.n930 39.2114
R3725 vdd.n2487 vdd.n929 39.2114
R3726 vdd.n2491 vdd.n928 39.2114
R3727 vdd.n2495 vdd.n927 39.2114
R3728 vdd.n2499 vdd.n926 39.2114
R3729 vdd.n2503 vdd.n925 39.2114
R3730 vdd.n2507 vdd.n924 39.2114
R3731 vdd.n2511 vdd.n923 39.2114
R3732 vdd.n2515 vdd.n922 39.2114
R3733 vdd.n2519 vdd.n921 39.2114
R3734 vdd.n2523 vdd.n920 39.2114
R3735 vdd.n2527 vdd.n919 39.2114
R3736 vdd.n2370 vdd.n2369 39.2114
R3737 vdd.n2367 vdd.n2366 39.2114
R3738 vdd.n2362 vdd.n2361 39.2114
R3739 vdd.n2359 vdd.n2358 39.2114
R3740 vdd.n2354 vdd.n2353 39.2114
R3741 vdd.n2351 vdd.n2350 39.2114
R3742 vdd.n2346 vdd.n2345 39.2114
R3743 vdd.n2343 vdd.n2342 39.2114
R3744 vdd.n1062 vdd.n1061 39.2114
R3745 vdd.n2186 vdd.n2185 39.2114
R3746 vdd.n2191 vdd.n2190 39.2114
R3747 vdd.n2192 vdd.n2182 39.2114
R3748 vdd.n2199 vdd.n2198 39.2114
R3749 vdd.n2200 vdd.n2180 39.2114
R3750 vdd.n2207 vdd.n2206 39.2114
R3751 vdd.n2208 vdd.n2176 39.2114
R3752 vdd.n2216 vdd.n2215 39.2114
R3753 vdd.n2335 vdd.n2334 37.2369
R3754 vdd.n2038 vdd.n1971 37.2369
R3755 vdd.n2077 vdd.n1931 37.2369
R3756 vdd.n3138 vdd.n769 37.2369
R3757 vdd.n3186 vdd.n3185 37.2369
R3758 vdd.n690 vdd.n689 37.2369
R3759 vdd.n2377 vdd.n1047 31.6883
R3760 vdd.n2602 vdd.n956 31.6883
R3761 vdd.n2535 vdd.n959 31.6883
R3762 vdd.n2281 vdd.n2278 31.6883
R3763 vdd.n2789 vdd.n2787 31.6883
R3764 vdd.n2994 vdd.n2993 31.6883
R3765 vdd.n2866 vdd.n912 31.6883
R3766 vdd.n3057 vdd.n3056 31.6883
R3767 vdd.n2976 vdd.n2975 31.6883
R3768 vdd.n3062 vdd.n802 31.6883
R3769 vdd.n2708 vdd.n2707 31.6883
R3770 vdd.n2862 vdd.n2861 31.6883
R3771 vdd.n2373 vdd.n2372 31.6883
R3772 vdd.n2530 vdd.n2529 31.6883
R3773 vdd.n2462 vdd.n2461 31.6883
R3774 vdd.n2219 vdd.n2218 31.6883
R3775 vdd.n2212 vdd.n2178 30.449
R3776 vdd.n967 vdd.n966 30.449
R3777 vdd.n2153 vdd.n2152 30.449
R3778 vdd.n2540 vdd.n958 30.449
R3779 vdd.n2644 vdd.n2643 30.449
R3780 vdd.n3000 vdd.n833 30.449
R3781 vdd.n2794 vdd.n2640 30.449
R3782 vdd.n801 vdd.n800 30.449
R3783 vdd.n1418 vdd.n1225 22.2201
R3784 vdd.n2329 vdd.n1073 22.2201
R3785 vdd.n3223 vdd.n723 22.2201
R3786 vdd.n3355 vdd.n3354 22.2201
R3787 vdd.n1429 vdd.n1187 19.3944
R3788 vdd.n1429 vdd.n1185 19.3944
R3789 vdd.n1433 vdd.n1185 19.3944
R3790 vdd.n1433 vdd.n1175 19.3944
R3791 vdd.n1446 vdd.n1175 19.3944
R3792 vdd.n1446 vdd.n1173 19.3944
R3793 vdd.n1450 vdd.n1173 19.3944
R3794 vdd.n1450 vdd.n1165 19.3944
R3795 vdd.n1463 vdd.n1165 19.3944
R3796 vdd.n1463 vdd.n1163 19.3944
R3797 vdd.n1467 vdd.n1163 19.3944
R3798 vdd.n1467 vdd.n1152 19.3944
R3799 vdd.n1479 vdd.n1152 19.3944
R3800 vdd.n1479 vdd.n1150 19.3944
R3801 vdd.n1483 vdd.n1150 19.3944
R3802 vdd.n1483 vdd.n1141 19.3944
R3803 vdd.n1496 vdd.n1141 19.3944
R3804 vdd.n1496 vdd.n1139 19.3944
R3805 vdd.n1500 vdd.n1139 19.3944
R3806 vdd.n1500 vdd.n1130 19.3944
R3807 vdd.n1819 vdd.n1130 19.3944
R3808 vdd.n1819 vdd.n1128 19.3944
R3809 vdd.n1823 vdd.n1128 19.3944
R3810 vdd.n1823 vdd.n1118 19.3944
R3811 vdd.n1836 vdd.n1118 19.3944
R3812 vdd.n1836 vdd.n1116 19.3944
R3813 vdd.n1840 vdd.n1116 19.3944
R3814 vdd.n1840 vdd.n1108 19.3944
R3815 vdd.n1853 vdd.n1108 19.3944
R3816 vdd.n1853 vdd.n1106 19.3944
R3817 vdd.n1857 vdd.n1106 19.3944
R3818 vdd.n1857 vdd.n1095 19.3944
R3819 vdd.n1869 vdd.n1095 19.3944
R3820 vdd.n1869 vdd.n1093 19.3944
R3821 vdd.n1873 vdd.n1093 19.3944
R3822 vdd.n1873 vdd.n1085 19.3944
R3823 vdd.n1886 vdd.n1085 19.3944
R3824 vdd.n1886 vdd.n1082 19.3944
R3825 vdd.n1892 vdd.n1082 19.3944
R3826 vdd.n1892 vdd.n1083 19.3944
R3827 vdd.n1083 vdd.n1072 19.3944
R3828 vdd.n1353 vdd.n1288 19.3944
R3829 vdd.n1349 vdd.n1288 19.3944
R3830 vdd.n1349 vdd.n1348 19.3944
R3831 vdd.n1348 vdd.n1347 19.3944
R3832 vdd.n1347 vdd.n1294 19.3944
R3833 vdd.n1343 vdd.n1294 19.3944
R3834 vdd.n1343 vdd.n1342 19.3944
R3835 vdd.n1342 vdd.n1341 19.3944
R3836 vdd.n1341 vdd.n1300 19.3944
R3837 vdd.n1337 vdd.n1300 19.3944
R3838 vdd.n1337 vdd.n1336 19.3944
R3839 vdd.n1336 vdd.n1335 19.3944
R3840 vdd.n1335 vdd.n1306 19.3944
R3841 vdd.n1331 vdd.n1306 19.3944
R3842 vdd.n1331 vdd.n1330 19.3944
R3843 vdd.n1330 vdd.n1329 19.3944
R3844 vdd.n1329 vdd.n1312 19.3944
R3845 vdd.n1325 vdd.n1312 19.3944
R3846 vdd.n1325 vdd.n1324 19.3944
R3847 vdd.n1324 vdd.n1323 19.3944
R3848 vdd.n1388 vdd.n1387 19.3944
R3849 vdd.n1387 vdd.n1386 19.3944
R3850 vdd.n1386 vdd.n1259 19.3944
R3851 vdd.n1382 vdd.n1259 19.3944
R3852 vdd.n1382 vdd.n1381 19.3944
R3853 vdd.n1381 vdd.n1380 19.3944
R3854 vdd.n1380 vdd.n1265 19.3944
R3855 vdd.n1376 vdd.n1265 19.3944
R3856 vdd.n1376 vdd.n1375 19.3944
R3857 vdd.n1375 vdd.n1374 19.3944
R3858 vdd.n1374 vdd.n1271 19.3944
R3859 vdd.n1370 vdd.n1271 19.3944
R3860 vdd.n1370 vdd.n1369 19.3944
R3861 vdd.n1369 vdd.n1368 19.3944
R3862 vdd.n1368 vdd.n1277 19.3944
R3863 vdd.n1364 vdd.n1277 19.3944
R3864 vdd.n1364 vdd.n1363 19.3944
R3865 vdd.n1363 vdd.n1362 19.3944
R3866 vdd.n1362 vdd.n1283 19.3944
R3867 vdd.n1358 vdd.n1283 19.3944
R3868 vdd.n1421 vdd.n1192 19.3944
R3869 vdd.n1416 vdd.n1192 19.3944
R3870 vdd.n1416 vdd.n1227 19.3944
R3871 vdd.n1412 vdd.n1227 19.3944
R3872 vdd.n1412 vdd.n1411 19.3944
R3873 vdd.n1411 vdd.n1410 19.3944
R3874 vdd.n1410 vdd.n1233 19.3944
R3875 vdd.n1406 vdd.n1233 19.3944
R3876 vdd.n1406 vdd.n1405 19.3944
R3877 vdd.n1405 vdd.n1404 19.3944
R3878 vdd.n1404 vdd.n1239 19.3944
R3879 vdd.n1400 vdd.n1239 19.3944
R3880 vdd.n1400 vdd.n1399 19.3944
R3881 vdd.n1399 vdd.n1398 19.3944
R3882 vdd.n1398 vdd.n1245 19.3944
R3883 vdd.n1394 vdd.n1245 19.3944
R3884 vdd.n1394 vdd.n1393 19.3944
R3885 vdd.n1393 vdd.n1392 19.3944
R3886 vdd.n2034 vdd.n1969 19.3944
R3887 vdd.n2034 vdd.n1975 19.3944
R3888 vdd.n2029 vdd.n1975 19.3944
R3889 vdd.n2029 vdd.n2028 19.3944
R3890 vdd.n2028 vdd.n2027 19.3944
R3891 vdd.n2027 vdd.n1982 19.3944
R3892 vdd.n2022 vdd.n1982 19.3944
R3893 vdd.n2022 vdd.n2021 19.3944
R3894 vdd.n2021 vdd.n2020 19.3944
R3895 vdd.n2020 vdd.n1989 19.3944
R3896 vdd.n2015 vdd.n1989 19.3944
R3897 vdd.n2015 vdd.n2014 19.3944
R3898 vdd.n2014 vdd.n2013 19.3944
R3899 vdd.n2013 vdd.n1997 19.3944
R3900 vdd.n2008 vdd.n1997 19.3944
R3901 vdd.n2008 vdd.n2007 19.3944
R3902 vdd.n2003 vdd.n2002 19.3944
R3903 vdd.n2336 vdd.n1068 19.3944
R3904 vdd.n2073 vdd.n1929 19.3944
R3905 vdd.n2073 vdd.n1935 19.3944
R3906 vdd.n2068 vdd.n1935 19.3944
R3907 vdd.n2068 vdd.n2067 19.3944
R3908 vdd.n2067 vdd.n2066 19.3944
R3909 vdd.n2066 vdd.n1942 19.3944
R3910 vdd.n2061 vdd.n1942 19.3944
R3911 vdd.n2061 vdd.n2060 19.3944
R3912 vdd.n2060 vdd.n2059 19.3944
R3913 vdd.n2059 vdd.n1949 19.3944
R3914 vdd.n2054 vdd.n1949 19.3944
R3915 vdd.n2054 vdd.n2053 19.3944
R3916 vdd.n2053 vdd.n2052 19.3944
R3917 vdd.n2052 vdd.n1956 19.3944
R3918 vdd.n2047 vdd.n1956 19.3944
R3919 vdd.n2047 vdd.n2046 19.3944
R3920 vdd.n2046 vdd.n2045 19.3944
R3921 vdd.n2045 vdd.n1963 19.3944
R3922 vdd.n2040 vdd.n1963 19.3944
R3923 vdd.n2040 vdd.n2039 19.3944
R3924 vdd.n2324 vdd.n2323 19.3944
R3925 vdd.n2323 vdd.n1901 19.3944
R3926 vdd.n2318 vdd.n2317 19.3944
R3927 vdd.n2100 vdd.n1905 19.3944
R3928 vdd.n2100 vdd.n1907 19.3944
R3929 vdd.n1910 vdd.n1907 19.3944
R3930 vdd.n2093 vdd.n1910 19.3944
R3931 vdd.n2093 vdd.n2092 19.3944
R3932 vdd.n2092 vdd.n2091 19.3944
R3933 vdd.n2091 vdd.n1916 19.3944
R3934 vdd.n2086 vdd.n1916 19.3944
R3935 vdd.n2086 vdd.n2085 19.3944
R3936 vdd.n2085 vdd.n2084 19.3944
R3937 vdd.n2084 vdd.n1923 19.3944
R3938 vdd.n2079 vdd.n1923 19.3944
R3939 vdd.n2079 vdd.n2078 19.3944
R3940 vdd.n1425 vdd.n1190 19.3944
R3941 vdd.n1425 vdd.n1181 19.3944
R3942 vdd.n1438 vdd.n1181 19.3944
R3943 vdd.n1438 vdd.n1179 19.3944
R3944 vdd.n1442 vdd.n1179 19.3944
R3945 vdd.n1442 vdd.n1170 19.3944
R3946 vdd.n1455 vdd.n1170 19.3944
R3947 vdd.n1455 vdd.n1168 19.3944
R3948 vdd.n1459 vdd.n1168 19.3944
R3949 vdd.n1459 vdd.n1159 19.3944
R3950 vdd.n1471 vdd.n1159 19.3944
R3951 vdd.n1471 vdd.n1157 19.3944
R3952 vdd.n1475 vdd.n1157 19.3944
R3953 vdd.n1475 vdd.n1147 19.3944
R3954 vdd.n1488 vdd.n1147 19.3944
R3955 vdd.n1488 vdd.n1145 19.3944
R3956 vdd.n1492 vdd.n1145 19.3944
R3957 vdd.n1492 vdd.n1136 19.3944
R3958 vdd.n1504 vdd.n1136 19.3944
R3959 vdd.n1504 vdd.n1134 19.3944
R3960 vdd.n1815 vdd.n1134 19.3944
R3961 vdd.n1815 vdd.n1124 19.3944
R3962 vdd.n1828 vdd.n1124 19.3944
R3963 vdd.n1828 vdd.n1122 19.3944
R3964 vdd.n1832 vdd.n1122 19.3944
R3965 vdd.n1832 vdd.n1113 19.3944
R3966 vdd.n1845 vdd.n1113 19.3944
R3967 vdd.n1845 vdd.n1111 19.3944
R3968 vdd.n1849 vdd.n1111 19.3944
R3969 vdd.n1849 vdd.n1102 19.3944
R3970 vdd.n1861 vdd.n1102 19.3944
R3971 vdd.n1861 vdd.n1100 19.3944
R3972 vdd.n1865 vdd.n1100 19.3944
R3973 vdd.n1865 vdd.n1090 19.3944
R3974 vdd.n1878 vdd.n1090 19.3944
R3975 vdd.n1878 vdd.n1088 19.3944
R3976 vdd.n1882 vdd.n1088 19.3944
R3977 vdd.n1882 vdd.n1078 19.3944
R3978 vdd.n1897 vdd.n1078 19.3944
R3979 vdd.n1897 vdd.n1076 19.3944
R3980 vdd.n2327 vdd.n1076 19.3944
R3981 vdd.n3229 vdd.n686 19.3944
R3982 vdd.n3229 vdd.n676 19.3944
R3983 vdd.n3241 vdd.n676 19.3944
R3984 vdd.n3241 vdd.n674 19.3944
R3985 vdd.n3245 vdd.n674 19.3944
R3986 vdd.n3245 vdd.n666 19.3944
R3987 vdd.n3258 vdd.n666 19.3944
R3988 vdd.n3258 vdd.n664 19.3944
R3989 vdd.n3262 vdd.n664 19.3944
R3990 vdd.n3262 vdd.n653 19.3944
R3991 vdd.n3274 vdd.n653 19.3944
R3992 vdd.n3274 vdd.n651 19.3944
R3993 vdd.n3278 vdd.n651 19.3944
R3994 vdd.n3278 vdd.n642 19.3944
R3995 vdd.n3291 vdd.n642 19.3944
R3996 vdd.n3291 vdd.n640 19.3944
R3997 vdd.n3298 vdd.n640 19.3944
R3998 vdd.n3298 vdd.n3297 19.3944
R3999 vdd.n3297 vdd.n631 19.3944
R4000 vdd.n3311 vdd.n631 19.3944
R4001 vdd.n3312 vdd.n3311 19.3944
R4002 vdd.n3312 vdd.n629 19.3944
R4003 vdd.n3316 vdd.n629 19.3944
R4004 vdd.n3318 vdd.n3316 19.3944
R4005 vdd.n3319 vdd.n3318 19.3944
R4006 vdd.n3319 vdd.n627 19.3944
R4007 vdd.n3323 vdd.n627 19.3944
R4008 vdd.n3325 vdd.n3323 19.3944
R4009 vdd.n3326 vdd.n3325 19.3944
R4010 vdd.n3326 vdd.n625 19.3944
R4011 vdd.n3330 vdd.n625 19.3944
R4012 vdd.n3333 vdd.n3330 19.3944
R4013 vdd.n3334 vdd.n3333 19.3944
R4014 vdd.n3334 vdd.n623 19.3944
R4015 vdd.n3338 vdd.n623 19.3944
R4016 vdd.n3340 vdd.n3338 19.3944
R4017 vdd.n3341 vdd.n3340 19.3944
R4018 vdd.n3341 vdd.n621 19.3944
R4019 vdd.n3345 vdd.n621 19.3944
R4020 vdd.n3347 vdd.n3345 19.3944
R4021 vdd.n3348 vdd.n3347 19.3944
R4022 vdd.n569 vdd.n438 19.3944
R4023 vdd.n575 vdd.n438 19.3944
R4024 vdd.n576 vdd.n575 19.3944
R4025 vdd.n579 vdd.n576 19.3944
R4026 vdd.n579 vdd.n436 19.3944
R4027 vdd.n585 vdd.n436 19.3944
R4028 vdd.n586 vdd.n585 19.3944
R4029 vdd.n589 vdd.n586 19.3944
R4030 vdd.n589 vdd.n434 19.3944
R4031 vdd.n595 vdd.n434 19.3944
R4032 vdd.n596 vdd.n595 19.3944
R4033 vdd.n599 vdd.n596 19.3944
R4034 vdd.n599 vdd.n432 19.3944
R4035 vdd.n605 vdd.n432 19.3944
R4036 vdd.n606 vdd.n605 19.3944
R4037 vdd.n609 vdd.n606 19.3944
R4038 vdd.n609 vdd.n430 19.3944
R4039 vdd.n615 vdd.n430 19.3944
R4040 vdd.n617 vdd.n615 19.3944
R4041 vdd.n618 vdd.n617 19.3944
R4042 vdd.n516 vdd.n515 19.3944
R4043 vdd.n519 vdd.n516 19.3944
R4044 vdd.n519 vdd.n450 19.3944
R4045 vdd.n525 vdd.n450 19.3944
R4046 vdd.n526 vdd.n525 19.3944
R4047 vdd.n529 vdd.n526 19.3944
R4048 vdd.n529 vdd.n448 19.3944
R4049 vdd.n535 vdd.n448 19.3944
R4050 vdd.n536 vdd.n535 19.3944
R4051 vdd.n539 vdd.n536 19.3944
R4052 vdd.n539 vdd.n446 19.3944
R4053 vdd.n545 vdd.n446 19.3944
R4054 vdd.n546 vdd.n545 19.3944
R4055 vdd.n549 vdd.n546 19.3944
R4056 vdd.n549 vdd.n444 19.3944
R4057 vdd.n555 vdd.n444 19.3944
R4058 vdd.n556 vdd.n555 19.3944
R4059 vdd.n559 vdd.n556 19.3944
R4060 vdd.n559 vdd.n442 19.3944
R4061 vdd.n565 vdd.n442 19.3944
R4062 vdd.n466 vdd.n465 19.3944
R4063 vdd.n469 vdd.n466 19.3944
R4064 vdd.n469 vdd.n462 19.3944
R4065 vdd.n475 vdd.n462 19.3944
R4066 vdd.n476 vdd.n475 19.3944
R4067 vdd.n479 vdd.n476 19.3944
R4068 vdd.n479 vdd.n460 19.3944
R4069 vdd.n485 vdd.n460 19.3944
R4070 vdd.n486 vdd.n485 19.3944
R4071 vdd.n489 vdd.n486 19.3944
R4072 vdd.n489 vdd.n458 19.3944
R4073 vdd.n495 vdd.n458 19.3944
R4074 vdd.n496 vdd.n495 19.3944
R4075 vdd.n499 vdd.n496 19.3944
R4076 vdd.n499 vdd.n456 19.3944
R4077 vdd.n505 vdd.n456 19.3944
R4078 vdd.n506 vdd.n505 19.3944
R4079 vdd.n509 vdd.n506 19.3944
R4080 vdd.n3233 vdd.n683 19.3944
R4081 vdd.n3233 vdd.n681 19.3944
R4082 vdd.n3237 vdd.n681 19.3944
R4083 vdd.n3237 vdd.n671 19.3944
R4084 vdd.n3250 vdd.n671 19.3944
R4085 vdd.n3250 vdd.n669 19.3944
R4086 vdd.n3254 vdd.n669 19.3944
R4087 vdd.n3254 vdd.n660 19.3944
R4088 vdd.n3266 vdd.n660 19.3944
R4089 vdd.n3266 vdd.n658 19.3944
R4090 vdd.n3270 vdd.n658 19.3944
R4091 vdd.n3270 vdd.n648 19.3944
R4092 vdd.n3283 vdd.n648 19.3944
R4093 vdd.n3283 vdd.n646 19.3944
R4094 vdd.n3287 vdd.n646 19.3944
R4095 vdd.n3287 vdd.n637 19.3944
R4096 vdd.n3302 vdd.n637 19.3944
R4097 vdd.n3302 vdd.n635 19.3944
R4098 vdd.n3306 vdd.n635 19.3944
R4099 vdd.n3306 vdd.n336 19.3944
R4100 vdd.n3397 vdd.n336 19.3944
R4101 vdd.n3397 vdd.n337 19.3944
R4102 vdd.n3391 vdd.n337 19.3944
R4103 vdd.n3391 vdd.n3390 19.3944
R4104 vdd.n3390 vdd.n3389 19.3944
R4105 vdd.n3389 vdd.n349 19.3944
R4106 vdd.n3383 vdd.n349 19.3944
R4107 vdd.n3383 vdd.n3382 19.3944
R4108 vdd.n3382 vdd.n3381 19.3944
R4109 vdd.n3381 vdd.n359 19.3944
R4110 vdd.n3375 vdd.n359 19.3944
R4111 vdd.n3375 vdd.n3374 19.3944
R4112 vdd.n3374 vdd.n3373 19.3944
R4113 vdd.n3373 vdd.n370 19.3944
R4114 vdd.n3367 vdd.n370 19.3944
R4115 vdd.n3367 vdd.n3366 19.3944
R4116 vdd.n3366 vdd.n3365 19.3944
R4117 vdd.n3365 vdd.n381 19.3944
R4118 vdd.n3359 vdd.n381 19.3944
R4119 vdd.n3359 vdd.n3358 19.3944
R4120 vdd.n3358 vdd.n3357 19.3944
R4121 vdd.n3180 vdd.n747 19.3944
R4122 vdd.n3180 vdd.n3177 19.3944
R4123 vdd.n3177 vdd.n3174 19.3944
R4124 vdd.n3174 vdd.n3173 19.3944
R4125 vdd.n3173 vdd.n3170 19.3944
R4126 vdd.n3170 vdd.n3169 19.3944
R4127 vdd.n3169 vdd.n3166 19.3944
R4128 vdd.n3166 vdd.n3165 19.3944
R4129 vdd.n3165 vdd.n3162 19.3944
R4130 vdd.n3162 vdd.n3161 19.3944
R4131 vdd.n3161 vdd.n3158 19.3944
R4132 vdd.n3158 vdd.n3157 19.3944
R4133 vdd.n3157 vdd.n3154 19.3944
R4134 vdd.n3154 vdd.n3153 19.3944
R4135 vdd.n3153 vdd.n3150 19.3944
R4136 vdd.n3150 vdd.n3149 19.3944
R4137 vdd.n3149 vdd.n3146 19.3944
R4138 vdd.n3146 vdd.n3145 19.3944
R4139 vdd.n3145 vdd.n3142 19.3944
R4140 vdd.n3142 vdd.n3141 19.3944
R4141 vdd.n3220 vdd.n3219 19.3944
R4142 vdd.n3219 vdd.n3218 19.3944
R4143 vdd.n732 vdd.n729 19.3944
R4144 vdd.n3214 vdd.n3213 19.3944
R4145 vdd.n3213 vdd.n3210 19.3944
R4146 vdd.n3210 vdd.n3209 19.3944
R4147 vdd.n3209 vdd.n3206 19.3944
R4148 vdd.n3206 vdd.n3205 19.3944
R4149 vdd.n3205 vdd.n3202 19.3944
R4150 vdd.n3202 vdd.n3201 19.3944
R4151 vdd.n3201 vdd.n3198 19.3944
R4152 vdd.n3198 vdd.n3197 19.3944
R4153 vdd.n3197 vdd.n3194 19.3944
R4154 vdd.n3194 vdd.n3193 19.3944
R4155 vdd.n3193 vdd.n3190 19.3944
R4156 vdd.n3190 vdd.n3189 19.3944
R4157 vdd.n3134 vdd.n767 19.3944
R4158 vdd.n3134 vdd.n3131 19.3944
R4159 vdd.n3131 vdd.n3128 19.3944
R4160 vdd.n3128 vdd.n3127 19.3944
R4161 vdd.n3127 vdd.n3124 19.3944
R4162 vdd.n3124 vdd.n3123 19.3944
R4163 vdd.n3123 vdd.n3120 19.3944
R4164 vdd.n3120 vdd.n3119 19.3944
R4165 vdd.n3119 vdd.n3116 19.3944
R4166 vdd.n3116 vdd.n3115 19.3944
R4167 vdd.n3115 vdd.n3112 19.3944
R4168 vdd.n3112 vdd.n3111 19.3944
R4169 vdd.n3111 vdd.n3108 19.3944
R4170 vdd.n3108 vdd.n3107 19.3944
R4171 vdd.n3107 vdd.n3104 19.3944
R4172 vdd.n3104 vdd.n3103 19.3944
R4173 vdd.n3100 vdd.n3099 19.3944
R4174 vdd.n3096 vdd.n3095 19.3944
R4175 vdd.n1357 vdd.n1353 19.0066
R4176 vdd.n2038 vdd.n1969 19.0066
R4177 vdd.n569 vdd.n566 19.0066
R4178 vdd.n3138 vdd.n767 19.0066
R4179 vdd.n2178 vdd.n2177 16.0975
R4180 vdd.n966 vdd.n965 16.0975
R4181 vdd.n1318 vdd.n1317 16.0975
R4182 vdd.n1356 vdd.n1355 16.0975
R4183 vdd.n1252 vdd.n1251 16.0975
R4184 vdd.n2334 vdd.n2333 16.0975
R4185 vdd.n1971 vdd.n1970 16.0975
R4186 vdd.n1931 vdd.n1930 16.0975
R4187 vdd.n2152 vdd.n2151 16.0975
R4188 vdd.n958 vdd.n957 16.0975
R4189 vdd.n2643 vdd.n2642 16.0975
R4190 vdd.n427 vdd.n426 16.0975
R4191 vdd.n441 vdd.n440 16.0975
R4192 vdd.n453 vdd.n452 16.0975
R4193 vdd.n769 vdd.n768 16.0975
R4194 vdd.n3185 vdd.n3184 16.0975
R4195 vdd.n833 vdd.n832 16.0975
R4196 vdd.n2640 vdd.n2639 16.0975
R4197 vdd.n689 vdd.n688 16.0975
R4198 vdd.n800 vdd.n799 16.0975
R4199 vdd.t87 vdd.n2604 15.4182
R4200 vdd.n2857 vdd.t115 15.4182
R4201 vdd.n28 vdd.n27 14.7125
R4202 vdd.n2375 vdd.n1049 14.5112
R4203 vdd.n3059 vdd.n692 14.5112
R4204 vdd.n328 vdd.n293 13.1884
R4205 vdd.n269 vdd.n234 13.1884
R4206 vdd.n226 vdd.n191 13.1884
R4207 vdd.n167 vdd.n132 13.1884
R4208 vdd.n125 vdd.n90 13.1884
R4209 vdd.n66 vdd.n31 13.1884
R4210 vdd.n1747 vdd.n1712 13.1884
R4211 vdd.n1806 vdd.n1771 13.1884
R4212 vdd.n1645 vdd.n1610 13.1884
R4213 vdd.n1704 vdd.n1669 13.1884
R4214 vdd.n1544 vdd.n1509 13.1884
R4215 vdd.n1603 vdd.n1568 13.1884
R4216 vdd.n1388 vdd.n1253 12.9944
R4217 vdd.n1392 vdd.n1253 12.9944
R4218 vdd.n2077 vdd.n1929 12.9944
R4219 vdd.n2078 vdd.n2077 12.9944
R4220 vdd.n515 vdd.n454 12.9944
R4221 vdd.n509 vdd.n454 12.9944
R4222 vdd.n3186 vdd.n747 12.9944
R4223 vdd.n3189 vdd.n3186 12.9944
R4224 vdd.n329 vdd.n291 12.8005
R4225 vdd.n324 vdd.n295 12.8005
R4226 vdd.n270 vdd.n232 12.8005
R4227 vdd.n265 vdd.n236 12.8005
R4228 vdd.n227 vdd.n189 12.8005
R4229 vdd.n222 vdd.n193 12.8005
R4230 vdd.n168 vdd.n130 12.8005
R4231 vdd.n163 vdd.n134 12.8005
R4232 vdd.n126 vdd.n88 12.8005
R4233 vdd.n121 vdd.n92 12.8005
R4234 vdd.n67 vdd.n29 12.8005
R4235 vdd.n62 vdd.n33 12.8005
R4236 vdd.n1748 vdd.n1710 12.8005
R4237 vdd.n1743 vdd.n1714 12.8005
R4238 vdd.n1807 vdd.n1769 12.8005
R4239 vdd.n1802 vdd.n1773 12.8005
R4240 vdd.n1646 vdd.n1608 12.8005
R4241 vdd.n1641 vdd.n1612 12.8005
R4242 vdd.n1705 vdd.n1667 12.8005
R4243 vdd.n1700 vdd.n1671 12.8005
R4244 vdd.n1545 vdd.n1507 12.8005
R4245 vdd.n1540 vdd.n1511 12.8005
R4246 vdd.n1604 vdd.n1566 12.8005
R4247 vdd.n1599 vdd.n1570 12.8005
R4248 vdd.n323 vdd.n296 12.0247
R4249 vdd.n264 vdd.n237 12.0247
R4250 vdd.n221 vdd.n194 12.0247
R4251 vdd.n162 vdd.n135 12.0247
R4252 vdd.n120 vdd.n93 12.0247
R4253 vdd.n61 vdd.n34 12.0247
R4254 vdd.n1742 vdd.n1715 12.0247
R4255 vdd.n1801 vdd.n1774 12.0247
R4256 vdd.n1640 vdd.n1613 12.0247
R4257 vdd.n1699 vdd.n1672 12.0247
R4258 vdd.n1539 vdd.n1512 12.0247
R4259 vdd.n1598 vdd.n1571 12.0247
R4260 vdd.n1427 vdd.n1183 11.337
R4261 vdd.n1436 vdd.n1183 11.337
R4262 vdd.n1436 vdd.n1435 11.337
R4263 vdd.n1444 vdd.n1177 11.337
R4264 vdd.n1453 vdd.n1452 11.337
R4265 vdd.n1469 vdd.n1161 11.337
R4266 vdd.n1477 vdd.n1154 11.337
R4267 vdd.n1486 vdd.n1485 11.337
R4268 vdd.n1494 vdd.n1143 11.337
R4269 vdd.n1817 vdd.n1132 11.337
R4270 vdd.n1826 vdd.n1126 11.337
R4271 vdd.n1834 vdd.n1120 11.337
R4272 vdd.n1843 vdd.n1842 11.337
R4273 vdd.n1859 vdd.n1104 11.337
R4274 vdd.n1867 vdd.n1097 11.337
R4275 vdd.n1876 vdd.n1875 11.337
R4276 vdd.n1884 vdd.n1080 11.337
R4277 vdd.n1895 vdd.n1080 11.337
R4278 vdd.n1895 vdd.n1894 11.337
R4279 vdd.n3231 vdd.n678 11.337
R4280 vdd.n3239 vdd.n678 11.337
R4281 vdd.n3239 vdd.n679 11.337
R4282 vdd.n3248 vdd.n3247 11.337
R4283 vdd.n3264 vdd.n662 11.337
R4284 vdd.n3272 vdd.n655 11.337
R4285 vdd.n3281 vdd.n3280 11.337
R4286 vdd.n3289 vdd.n644 11.337
R4287 vdd.n3308 vdd.n633 11.337
R4288 vdd.n3395 vdd.n340 11.337
R4289 vdd.n3393 vdd.n344 11.337
R4290 vdd.n3387 vdd.n3386 11.337
R4291 vdd.n3379 vdd.n361 11.337
R4292 vdd.n3378 vdd.n3377 11.337
R4293 vdd.n3371 vdd.n3370 11.337
R4294 vdd.n3369 vdd.n375 11.337
R4295 vdd.n3363 vdd.n3362 11.337
R4296 vdd.n3362 vdd.n3361 11.337
R4297 vdd.n3361 vdd.n386 11.337
R4298 vdd.n320 vdd.n319 11.249
R4299 vdd.n261 vdd.n260 11.249
R4300 vdd.n218 vdd.n217 11.249
R4301 vdd.n159 vdd.n158 11.249
R4302 vdd.n117 vdd.n116 11.249
R4303 vdd.n58 vdd.n57 11.249
R4304 vdd.n1739 vdd.n1738 11.249
R4305 vdd.n1798 vdd.n1797 11.249
R4306 vdd.n1637 vdd.n1636 11.249
R4307 vdd.n1696 vdd.n1695 11.249
R4308 vdd.n1536 vdd.n1535 11.249
R4309 vdd.n1595 vdd.n1594 11.249
R4310 vdd.n1225 vdd.t31 11.2237
R4311 vdd.n3355 vdd.t38 11.2237
R4312 vdd.n2532 vdd.t94 11.1103
R4313 vdd.n2864 vdd.t5 11.1103
R4314 vdd.t133 vdd.n1098 10.7702
R4315 vdd.n3256 vdd.t214 10.7702
R4316 vdd.n305 vdd.n304 10.7238
R4317 vdd.n246 vdd.n245 10.7238
R4318 vdd.n203 vdd.n202 10.7238
R4319 vdd.n144 vdd.n143 10.7238
R4320 vdd.n102 vdd.n101 10.7238
R4321 vdd.n43 vdd.n42 10.7238
R4322 vdd.n1724 vdd.n1723 10.7238
R4323 vdd.n1783 vdd.n1782 10.7238
R4324 vdd.n1622 vdd.n1621 10.7238
R4325 vdd.n1681 vdd.n1680 10.7238
R4326 vdd.n1521 vdd.n1520 10.7238
R4327 vdd.n1580 vdd.n1579 10.7238
R4328 vdd.n2378 vdd.n2377 10.6151
R4329 vdd.n2379 vdd.n2378 10.6151
R4330 vdd.n2379 vdd.n1035 10.6151
R4331 vdd.n2389 vdd.n1035 10.6151
R4332 vdd.n2390 vdd.n2389 10.6151
R4333 vdd.n2391 vdd.n2390 10.6151
R4334 vdd.n2391 vdd.n1022 10.6151
R4335 vdd.n2402 vdd.n1022 10.6151
R4336 vdd.n2403 vdd.n2402 10.6151
R4337 vdd.n2404 vdd.n2403 10.6151
R4338 vdd.n2404 vdd.n1010 10.6151
R4339 vdd.n2414 vdd.n1010 10.6151
R4340 vdd.n2415 vdd.n2414 10.6151
R4341 vdd.n2416 vdd.n2415 10.6151
R4342 vdd.n2416 vdd.n998 10.6151
R4343 vdd.n2426 vdd.n998 10.6151
R4344 vdd.n2427 vdd.n2426 10.6151
R4345 vdd.n2428 vdd.n2427 10.6151
R4346 vdd.n2428 vdd.n987 10.6151
R4347 vdd.n2438 vdd.n987 10.6151
R4348 vdd.n2439 vdd.n2438 10.6151
R4349 vdd.n2440 vdd.n2439 10.6151
R4350 vdd.n2440 vdd.n974 10.6151
R4351 vdd.n2452 vdd.n974 10.6151
R4352 vdd.n2453 vdd.n2452 10.6151
R4353 vdd.n2455 vdd.n2453 10.6151
R4354 vdd.n2455 vdd.n2454 10.6151
R4355 vdd.n2454 vdd.n956 10.6151
R4356 vdd.n2602 vdd.n2601 10.6151
R4357 vdd.n2601 vdd.n2600 10.6151
R4358 vdd.n2600 vdd.n2597 10.6151
R4359 vdd.n2597 vdd.n2596 10.6151
R4360 vdd.n2596 vdd.n2593 10.6151
R4361 vdd.n2593 vdd.n2592 10.6151
R4362 vdd.n2592 vdd.n2589 10.6151
R4363 vdd.n2589 vdd.n2588 10.6151
R4364 vdd.n2588 vdd.n2585 10.6151
R4365 vdd.n2585 vdd.n2584 10.6151
R4366 vdd.n2584 vdd.n2581 10.6151
R4367 vdd.n2581 vdd.n2580 10.6151
R4368 vdd.n2580 vdd.n2577 10.6151
R4369 vdd.n2577 vdd.n2576 10.6151
R4370 vdd.n2576 vdd.n2573 10.6151
R4371 vdd.n2573 vdd.n2572 10.6151
R4372 vdd.n2572 vdd.n2569 10.6151
R4373 vdd.n2569 vdd.n2568 10.6151
R4374 vdd.n2568 vdd.n2565 10.6151
R4375 vdd.n2565 vdd.n2564 10.6151
R4376 vdd.n2564 vdd.n2561 10.6151
R4377 vdd.n2561 vdd.n2560 10.6151
R4378 vdd.n2560 vdd.n2557 10.6151
R4379 vdd.n2557 vdd.n2556 10.6151
R4380 vdd.n2556 vdd.n2553 10.6151
R4381 vdd.n2553 vdd.n2552 10.6151
R4382 vdd.n2552 vdd.n2549 10.6151
R4383 vdd.n2549 vdd.n2548 10.6151
R4384 vdd.n2548 vdd.n2545 10.6151
R4385 vdd.n2545 vdd.n2544 10.6151
R4386 vdd.n2544 vdd.n2541 10.6151
R4387 vdd.n2539 vdd.n2536 10.6151
R4388 vdd.n2536 vdd.n2535 10.6151
R4389 vdd.n2278 vdd.n2277 10.6151
R4390 vdd.n2277 vdd.n2275 10.6151
R4391 vdd.n2275 vdd.n2274 10.6151
R4392 vdd.n2274 vdd.n2272 10.6151
R4393 vdd.n2272 vdd.n2271 10.6151
R4394 vdd.n2271 vdd.n2269 10.6151
R4395 vdd.n2269 vdd.n2268 10.6151
R4396 vdd.n2268 vdd.n2266 10.6151
R4397 vdd.n2266 vdd.n2265 10.6151
R4398 vdd.n2265 vdd.n2263 10.6151
R4399 vdd.n2263 vdd.n2262 10.6151
R4400 vdd.n2262 vdd.n2260 10.6151
R4401 vdd.n2260 vdd.n2259 10.6151
R4402 vdd.n2259 vdd.n2174 10.6151
R4403 vdd.n2174 vdd.n2173 10.6151
R4404 vdd.n2173 vdd.n2171 10.6151
R4405 vdd.n2171 vdd.n2170 10.6151
R4406 vdd.n2170 vdd.n2168 10.6151
R4407 vdd.n2168 vdd.n2167 10.6151
R4408 vdd.n2167 vdd.n2165 10.6151
R4409 vdd.n2165 vdd.n2164 10.6151
R4410 vdd.n2164 vdd.n2162 10.6151
R4411 vdd.n2162 vdd.n2161 10.6151
R4412 vdd.n2161 vdd.n2159 10.6151
R4413 vdd.n2159 vdd.n2158 10.6151
R4414 vdd.n2158 vdd.n2155 10.6151
R4415 vdd.n2155 vdd.n2154 10.6151
R4416 vdd.n2154 vdd.n959 10.6151
R4417 vdd.n2112 vdd.n1047 10.6151
R4418 vdd.n2113 vdd.n2112 10.6151
R4419 vdd.n2114 vdd.n2113 10.6151
R4420 vdd.n2114 vdd.n2108 10.6151
R4421 vdd.n2120 vdd.n2108 10.6151
R4422 vdd.n2121 vdd.n2120 10.6151
R4423 vdd.n2122 vdd.n2121 10.6151
R4424 vdd.n2122 vdd.n2106 10.6151
R4425 vdd.n2128 vdd.n2106 10.6151
R4426 vdd.n2129 vdd.n2128 10.6151
R4427 vdd.n2130 vdd.n2129 10.6151
R4428 vdd.n2130 vdd.n2104 10.6151
R4429 vdd.n2136 vdd.n2104 10.6151
R4430 vdd.n2137 vdd.n2136 10.6151
R4431 vdd.n2138 vdd.n2137 10.6151
R4432 vdd.n2138 vdd.n2102 10.6151
R4433 vdd.n2314 vdd.n2102 10.6151
R4434 vdd.n2314 vdd.n2313 10.6151
R4435 vdd.n2313 vdd.n2143 10.6151
R4436 vdd.n2307 vdd.n2143 10.6151
R4437 vdd.n2307 vdd.n2306 10.6151
R4438 vdd.n2306 vdd.n2305 10.6151
R4439 vdd.n2305 vdd.n2145 10.6151
R4440 vdd.n2299 vdd.n2145 10.6151
R4441 vdd.n2299 vdd.n2298 10.6151
R4442 vdd.n2298 vdd.n2297 10.6151
R4443 vdd.n2297 vdd.n2147 10.6151
R4444 vdd.n2291 vdd.n2147 10.6151
R4445 vdd.n2291 vdd.n2290 10.6151
R4446 vdd.n2290 vdd.n2289 10.6151
R4447 vdd.n2289 vdd.n2149 10.6151
R4448 vdd.n2283 vdd.n2282 10.6151
R4449 vdd.n2282 vdd.n2281 10.6151
R4450 vdd.n2787 vdd.n2786 10.6151
R4451 vdd.n2786 vdd.n2784 10.6151
R4452 vdd.n2784 vdd.n2783 10.6151
R4453 vdd.n2783 vdd.n2641 10.6151
R4454 vdd.n2730 vdd.n2641 10.6151
R4455 vdd.n2731 vdd.n2730 10.6151
R4456 vdd.n2733 vdd.n2731 10.6151
R4457 vdd.n2734 vdd.n2733 10.6151
R4458 vdd.n2736 vdd.n2734 10.6151
R4459 vdd.n2737 vdd.n2736 10.6151
R4460 vdd.n2739 vdd.n2737 10.6151
R4461 vdd.n2740 vdd.n2739 10.6151
R4462 vdd.n2742 vdd.n2740 10.6151
R4463 vdd.n2743 vdd.n2742 10.6151
R4464 vdd.n2758 vdd.n2743 10.6151
R4465 vdd.n2758 vdd.n2757 10.6151
R4466 vdd.n2757 vdd.n2756 10.6151
R4467 vdd.n2756 vdd.n2754 10.6151
R4468 vdd.n2754 vdd.n2753 10.6151
R4469 vdd.n2753 vdd.n2751 10.6151
R4470 vdd.n2751 vdd.n2750 10.6151
R4471 vdd.n2750 vdd.n2748 10.6151
R4472 vdd.n2748 vdd.n2747 10.6151
R4473 vdd.n2747 vdd.n2745 10.6151
R4474 vdd.n2745 vdd.n2744 10.6151
R4475 vdd.n2744 vdd.n836 10.6151
R4476 vdd.n2992 vdd.n836 10.6151
R4477 vdd.n2993 vdd.n2992 10.6151
R4478 vdd.n2854 vdd.n912 10.6151
R4479 vdd.n2854 vdd.n2853 10.6151
R4480 vdd.n2853 vdd.n2852 10.6151
R4481 vdd.n2852 vdd.n2850 10.6151
R4482 vdd.n2850 vdd.n2847 10.6151
R4483 vdd.n2847 vdd.n2846 10.6151
R4484 vdd.n2846 vdd.n2843 10.6151
R4485 vdd.n2843 vdd.n2842 10.6151
R4486 vdd.n2842 vdd.n2839 10.6151
R4487 vdd.n2839 vdd.n2838 10.6151
R4488 vdd.n2838 vdd.n2835 10.6151
R4489 vdd.n2835 vdd.n2834 10.6151
R4490 vdd.n2834 vdd.n2831 10.6151
R4491 vdd.n2831 vdd.n2830 10.6151
R4492 vdd.n2830 vdd.n2827 10.6151
R4493 vdd.n2827 vdd.n2826 10.6151
R4494 vdd.n2826 vdd.n2823 10.6151
R4495 vdd.n2823 vdd.n2822 10.6151
R4496 vdd.n2822 vdd.n2819 10.6151
R4497 vdd.n2819 vdd.n2818 10.6151
R4498 vdd.n2818 vdd.n2815 10.6151
R4499 vdd.n2815 vdd.n2814 10.6151
R4500 vdd.n2814 vdd.n2811 10.6151
R4501 vdd.n2811 vdd.n2810 10.6151
R4502 vdd.n2810 vdd.n2807 10.6151
R4503 vdd.n2807 vdd.n2806 10.6151
R4504 vdd.n2806 vdd.n2803 10.6151
R4505 vdd.n2803 vdd.n2802 10.6151
R4506 vdd.n2802 vdd.n2799 10.6151
R4507 vdd.n2799 vdd.n2798 10.6151
R4508 vdd.n2798 vdd.n2795 10.6151
R4509 vdd.n2793 vdd.n2790 10.6151
R4510 vdd.n2790 vdd.n2789 10.6151
R4511 vdd.n2867 vdd.n2866 10.6151
R4512 vdd.n2868 vdd.n2867 10.6151
R4513 vdd.n2868 vdd.n902 10.6151
R4514 vdd.n2878 vdd.n902 10.6151
R4515 vdd.n2879 vdd.n2878 10.6151
R4516 vdd.n2880 vdd.n2879 10.6151
R4517 vdd.n2880 vdd.n889 10.6151
R4518 vdd.n2890 vdd.n889 10.6151
R4519 vdd.n2891 vdd.n2890 10.6151
R4520 vdd.n2892 vdd.n2891 10.6151
R4521 vdd.n2892 vdd.n878 10.6151
R4522 vdd.n2902 vdd.n878 10.6151
R4523 vdd.n2903 vdd.n2902 10.6151
R4524 vdd.n2904 vdd.n2903 10.6151
R4525 vdd.n2904 vdd.n866 10.6151
R4526 vdd.n2914 vdd.n866 10.6151
R4527 vdd.n2915 vdd.n2914 10.6151
R4528 vdd.n2916 vdd.n2915 10.6151
R4529 vdd.n2916 vdd.n855 10.6151
R4530 vdd.n2928 vdd.n855 10.6151
R4531 vdd.n2929 vdd.n2928 10.6151
R4532 vdd.n2930 vdd.n2929 10.6151
R4533 vdd.n2930 vdd.n841 10.6151
R4534 vdd.n2985 vdd.n841 10.6151
R4535 vdd.n2986 vdd.n2985 10.6151
R4536 vdd.n2987 vdd.n2986 10.6151
R4537 vdd.n2987 vdd.n810 10.6151
R4538 vdd.n3057 vdd.n810 10.6151
R4539 vdd.n3056 vdd.n3055 10.6151
R4540 vdd.n3055 vdd.n811 10.6151
R4541 vdd.n812 vdd.n811 10.6151
R4542 vdd.n3048 vdd.n812 10.6151
R4543 vdd.n3048 vdd.n3047 10.6151
R4544 vdd.n3047 vdd.n3046 10.6151
R4545 vdd.n3046 vdd.n814 10.6151
R4546 vdd.n3041 vdd.n814 10.6151
R4547 vdd.n3041 vdd.n3040 10.6151
R4548 vdd.n3040 vdd.n3039 10.6151
R4549 vdd.n3039 vdd.n817 10.6151
R4550 vdd.n3034 vdd.n817 10.6151
R4551 vdd.n3034 vdd.n3033 10.6151
R4552 vdd.n3033 vdd.n3032 10.6151
R4553 vdd.n3032 vdd.n820 10.6151
R4554 vdd.n3027 vdd.n820 10.6151
R4555 vdd.n3027 vdd.n731 10.6151
R4556 vdd.n3023 vdd.n731 10.6151
R4557 vdd.n3023 vdd.n3022 10.6151
R4558 vdd.n3022 vdd.n3021 10.6151
R4559 vdd.n3021 vdd.n823 10.6151
R4560 vdd.n3016 vdd.n823 10.6151
R4561 vdd.n3016 vdd.n3015 10.6151
R4562 vdd.n3015 vdd.n3014 10.6151
R4563 vdd.n3014 vdd.n826 10.6151
R4564 vdd.n3009 vdd.n826 10.6151
R4565 vdd.n3009 vdd.n3008 10.6151
R4566 vdd.n3008 vdd.n3007 10.6151
R4567 vdd.n3007 vdd.n829 10.6151
R4568 vdd.n3002 vdd.n829 10.6151
R4569 vdd.n3002 vdd.n3001 10.6151
R4570 vdd.n2999 vdd.n834 10.6151
R4571 vdd.n2994 vdd.n834 10.6151
R4572 vdd.n2975 vdd.n2936 10.6151
R4573 vdd.n2970 vdd.n2936 10.6151
R4574 vdd.n2970 vdd.n2969 10.6151
R4575 vdd.n2969 vdd.n2968 10.6151
R4576 vdd.n2968 vdd.n2938 10.6151
R4577 vdd.n2963 vdd.n2938 10.6151
R4578 vdd.n2963 vdd.n2962 10.6151
R4579 vdd.n2962 vdd.n2961 10.6151
R4580 vdd.n2961 vdd.n2941 10.6151
R4581 vdd.n2956 vdd.n2941 10.6151
R4582 vdd.n2956 vdd.n2955 10.6151
R4583 vdd.n2955 vdd.n2954 10.6151
R4584 vdd.n2954 vdd.n2944 10.6151
R4585 vdd.n2949 vdd.n2944 10.6151
R4586 vdd.n2949 vdd.n2948 10.6151
R4587 vdd.n2948 vdd.n785 10.6151
R4588 vdd.n3092 vdd.n785 10.6151
R4589 vdd.n3092 vdd.n786 10.6151
R4590 vdd.n788 vdd.n786 10.6151
R4591 vdd.n3085 vdd.n788 10.6151
R4592 vdd.n3085 vdd.n3084 10.6151
R4593 vdd.n3084 vdd.n3083 10.6151
R4594 vdd.n3083 vdd.n790 10.6151
R4595 vdd.n3078 vdd.n790 10.6151
R4596 vdd.n3078 vdd.n3077 10.6151
R4597 vdd.n3077 vdd.n3076 10.6151
R4598 vdd.n3076 vdd.n793 10.6151
R4599 vdd.n3071 vdd.n793 10.6151
R4600 vdd.n3071 vdd.n3070 10.6151
R4601 vdd.n3070 vdd.n3069 10.6151
R4602 vdd.n3069 vdd.n796 10.6151
R4603 vdd.n3064 vdd.n3063 10.6151
R4604 vdd.n3063 vdd.n3062 10.6151
R4605 vdd.n2710 vdd.n2708 10.6151
R4606 vdd.n2711 vdd.n2710 10.6151
R4607 vdd.n2779 vdd.n2711 10.6151
R4608 vdd.n2779 vdd.n2778 10.6151
R4609 vdd.n2778 vdd.n2777 10.6151
R4610 vdd.n2777 vdd.n2775 10.6151
R4611 vdd.n2775 vdd.n2774 10.6151
R4612 vdd.n2774 vdd.n2772 10.6151
R4613 vdd.n2772 vdd.n2771 10.6151
R4614 vdd.n2771 vdd.n2769 10.6151
R4615 vdd.n2769 vdd.n2768 10.6151
R4616 vdd.n2768 vdd.n2766 10.6151
R4617 vdd.n2766 vdd.n2765 10.6151
R4618 vdd.n2765 vdd.n2763 10.6151
R4619 vdd.n2763 vdd.n2762 10.6151
R4620 vdd.n2762 vdd.n2728 10.6151
R4621 vdd.n2728 vdd.n2727 10.6151
R4622 vdd.n2727 vdd.n2725 10.6151
R4623 vdd.n2725 vdd.n2724 10.6151
R4624 vdd.n2724 vdd.n2722 10.6151
R4625 vdd.n2722 vdd.n2721 10.6151
R4626 vdd.n2721 vdd.n2719 10.6151
R4627 vdd.n2719 vdd.n2718 10.6151
R4628 vdd.n2718 vdd.n2716 10.6151
R4629 vdd.n2716 vdd.n2715 10.6151
R4630 vdd.n2715 vdd.n2713 10.6151
R4631 vdd.n2713 vdd.n2712 10.6151
R4632 vdd.n2712 vdd.n802 10.6151
R4633 vdd.n2861 vdd.n2860 10.6151
R4634 vdd.n2860 vdd.n917 10.6151
R4635 vdd.n2645 vdd.n917 10.6151
R4636 vdd.n2648 vdd.n2645 10.6151
R4637 vdd.n2649 vdd.n2648 10.6151
R4638 vdd.n2652 vdd.n2649 10.6151
R4639 vdd.n2653 vdd.n2652 10.6151
R4640 vdd.n2656 vdd.n2653 10.6151
R4641 vdd.n2657 vdd.n2656 10.6151
R4642 vdd.n2660 vdd.n2657 10.6151
R4643 vdd.n2661 vdd.n2660 10.6151
R4644 vdd.n2664 vdd.n2661 10.6151
R4645 vdd.n2665 vdd.n2664 10.6151
R4646 vdd.n2668 vdd.n2665 10.6151
R4647 vdd.n2669 vdd.n2668 10.6151
R4648 vdd.n2672 vdd.n2669 10.6151
R4649 vdd.n2673 vdd.n2672 10.6151
R4650 vdd.n2676 vdd.n2673 10.6151
R4651 vdd.n2677 vdd.n2676 10.6151
R4652 vdd.n2680 vdd.n2677 10.6151
R4653 vdd.n2681 vdd.n2680 10.6151
R4654 vdd.n2684 vdd.n2681 10.6151
R4655 vdd.n2685 vdd.n2684 10.6151
R4656 vdd.n2688 vdd.n2685 10.6151
R4657 vdd.n2689 vdd.n2688 10.6151
R4658 vdd.n2692 vdd.n2689 10.6151
R4659 vdd.n2693 vdd.n2692 10.6151
R4660 vdd.n2696 vdd.n2693 10.6151
R4661 vdd.n2697 vdd.n2696 10.6151
R4662 vdd.n2700 vdd.n2697 10.6151
R4663 vdd.n2701 vdd.n2700 10.6151
R4664 vdd.n2706 vdd.n2704 10.6151
R4665 vdd.n2707 vdd.n2706 10.6151
R4666 vdd.n2862 vdd.n907 10.6151
R4667 vdd.n2872 vdd.n907 10.6151
R4668 vdd.n2873 vdd.n2872 10.6151
R4669 vdd.n2874 vdd.n2873 10.6151
R4670 vdd.n2874 vdd.n895 10.6151
R4671 vdd.n2884 vdd.n895 10.6151
R4672 vdd.n2885 vdd.n2884 10.6151
R4673 vdd.n2886 vdd.n2885 10.6151
R4674 vdd.n2886 vdd.n884 10.6151
R4675 vdd.n2896 vdd.n884 10.6151
R4676 vdd.n2897 vdd.n2896 10.6151
R4677 vdd.n2898 vdd.n2897 10.6151
R4678 vdd.n2898 vdd.n872 10.6151
R4679 vdd.n2908 vdd.n872 10.6151
R4680 vdd.n2909 vdd.n2908 10.6151
R4681 vdd.n2910 vdd.n2909 10.6151
R4682 vdd.n2910 vdd.n861 10.6151
R4683 vdd.n2920 vdd.n861 10.6151
R4684 vdd.n2921 vdd.n2920 10.6151
R4685 vdd.n2924 vdd.n2921 10.6151
R4686 vdd.n2934 vdd.n849 10.6151
R4687 vdd.n2935 vdd.n2934 10.6151
R4688 vdd.n2981 vdd.n2935 10.6151
R4689 vdd.n2981 vdd.n2980 10.6151
R4690 vdd.n2980 vdd.n2979 10.6151
R4691 vdd.n2979 vdd.n2978 10.6151
R4692 vdd.n2978 vdd.n2976 10.6151
R4693 vdd.n2373 vdd.n1041 10.6151
R4694 vdd.n2383 vdd.n1041 10.6151
R4695 vdd.n2384 vdd.n2383 10.6151
R4696 vdd.n2385 vdd.n2384 10.6151
R4697 vdd.n2385 vdd.n1028 10.6151
R4698 vdd.n2395 vdd.n1028 10.6151
R4699 vdd.n2396 vdd.n2395 10.6151
R4700 vdd.n2398 vdd.n1016 10.6151
R4701 vdd.n2408 vdd.n1016 10.6151
R4702 vdd.n2409 vdd.n2408 10.6151
R4703 vdd.n2410 vdd.n2409 10.6151
R4704 vdd.n2410 vdd.n1004 10.6151
R4705 vdd.n2420 vdd.n1004 10.6151
R4706 vdd.n2421 vdd.n2420 10.6151
R4707 vdd.n2422 vdd.n2421 10.6151
R4708 vdd.n2422 vdd.n993 10.6151
R4709 vdd.n2432 vdd.n993 10.6151
R4710 vdd.n2433 vdd.n2432 10.6151
R4711 vdd.n2434 vdd.n2433 10.6151
R4712 vdd.n2434 vdd.n981 10.6151
R4713 vdd.n2444 vdd.n981 10.6151
R4714 vdd.n2445 vdd.n2444 10.6151
R4715 vdd.n2448 vdd.n2445 10.6151
R4716 vdd.n2448 vdd.n2447 10.6151
R4717 vdd.n2447 vdd.n2446 10.6151
R4718 vdd.n2446 vdd.n964 10.6151
R4719 vdd.n2530 vdd.n964 10.6151
R4720 vdd.n2529 vdd.n2528 10.6151
R4721 vdd.n2528 vdd.n2525 10.6151
R4722 vdd.n2525 vdd.n2524 10.6151
R4723 vdd.n2524 vdd.n2521 10.6151
R4724 vdd.n2521 vdd.n2520 10.6151
R4725 vdd.n2520 vdd.n2517 10.6151
R4726 vdd.n2517 vdd.n2516 10.6151
R4727 vdd.n2516 vdd.n2513 10.6151
R4728 vdd.n2513 vdd.n2512 10.6151
R4729 vdd.n2512 vdd.n2509 10.6151
R4730 vdd.n2509 vdd.n2508 10.6151
R4731 vdd.n2508 vdd.n2505 10.6151
R4732 vdd.n2505 vdd.n2504 10.6151
R4733 vdd.n2504 vdd.n2501 10.6151
R4734 vdd.n2501 vdd.n2500 10.6151
R4735 vdd.n2500 vdd.n2497 10.6151
R4736 vdd.n2497 vdd.n2496 10.6151
R4737 vdd.n2496 vdd.n2493 10.6151
R4738 vdd.n2493 vdd.n2492 10.6151
R4739 vdd.n2492 vdd.n2489 10.6151
R4740 vdd.n2489 vdd.n2488 10.6151
R4741 vdd.n2488 vdd.n2485 10.6151
R4742 vdd.n2485 vdd.n2484 10.6151
R4743 vdd.n2484 vdd.n2481 10.6151
R4744 vdd.n2481 vdd.n2480 10.6151
R4745 vdd.n2480 vdd.n2477 10.6151
R4746 vdd.n2477 vdd.n2476 10.6151
R4747 vdd.n2476 vdd.n2473 10.6151
R4748 vdd.n2473 vdd.n2472 10.6151
R4749 vdd.n2472 vdd.n2469 10.6151
R4750 vdd.n2469 vdd.n2468 10.6151
R4751 vdd.n2465 vdd.n2464 10.6151
R4752 vdd.n2464 vdd.n2462 10.6151
R4753 vdd.n2221 vdd.n2219 10.6151
R4754 vdd.n2222 vdd.n2221 10.6151
R4755 vdd.n2224 vdd.n2222 10.6151
R4756 vdd.n2225 vdd.n2224 10.6151
R4757 vdd.n2227 vdd.n2225 10.6151
R4758 vdd.n2228 vdd.n2227 10.6151
R4759 vdd.n2230 vdd.n2228 10.6151
R4760 vdd.n2231 vdd.n2230 10.6151
R4761 vdd.n2233 vdd.n2231 10.6151
R4762 vdd.n2234 vdd.n2233 10.6151
R4763 vdd.n2236 vdd.n2234 10.6151
R4764 vdd.n2237 vdd.n2236 10.6151
R4765 vdd.n2255 vdd.n2237 10.6151
R4766 vdd.n2255 vdd.n2254 10.6151
R4767 vdd.n2254 vdd.n2253 10.6151
R4768 vdd.n2253 vdd.n2251 10.6151
R4769 vdd.n2251 vdd.n2250 10.6151
R4770 vdd.n2250 vdd.n2248 10.6151
R4771 vdd.n2248 vdd.n2247 10.6151
R4772 vdd.n2247 vdd.n2245 10.6151
R4773 vdd.n2245 vdd.n2244 10.6151
R4774 vdd.n2244 vdd.n2242 10.6151
R4775 vdd.n2242 vdd.n2241 10.6151
R4776 vdd.n2241 vdd.n2239 10.6151
R4777 vdd.n2239 vdd.n2238 10.6151
R4778 vdd.n2238 vdd.n968 10.6151
R4779 vdd.n2460 vdd.n968 10.6151
R4780 vdd.n2461 vdd.n2460 10.6151
R4781 vdd.n2372 vdd.n2371 10.6151
R4782 vdd.n2371 vdd.n1053 10.6151
R4783 vdd.n2365 vdd.n1053 10.6151
R4784 vdd.n2365 vdd.n2364 10.6151
R4785 vdd.n2364 vdd.n2363 10.6151
R4786 vdd.n2363 vdd.n1055 10.6151
R4787 vdd.n2357 vdd.n1055 10.6151
R4788 vdd.n2357 vdd.n2356 10.6151
R4789 vdd.n2356 vdd.n2355 10.6151
R4790 vdd.n2355 vdd.n1057 10.6151
R4791 vdd.n2349 vdd.n1057 10.6151
R4792 vdd.n2349 vdd.n2348 10.6151
R4793 vdd.n2348 vdd.n2347 10.6151
R4794 vdd.n2347 vdd.n1059 10.6151
R4795 vdd.n2341 vdd.n1059 10.6151
R4796 vdd.n2341 vdd.n2340 10.6151
R4797 vdd.n2340 vdd.n2339 10.6151
R4798 vdd.n2339 vdd.n1063 10.6151
R4799 vdd.n2187 vdd.n1063 10.6151
R4800 vdd.n2188 vdd.n2187 10.6151
R4801 vdd.n2188 vdd.n2183 10.6151
R4802 vdd.n2194 vdd.n2183 10.6151
R4803 vdd.n2195 vdd.n2194 10.6151
R4804 vdd.n2196 vdd.n2195 10.6151
R4805 vdd.n2196 vdd.n2181 10.6151
R4806 vdd.n2202 vdd.n2181 10.6151
R4807 vdd.n2203 vdd.n2202 10.6151
R4808 vdd.n2204 vdd.n2203 10.6151
R4809 vdd.n2204 vdd.n2179 10.6151
R4810 vdd.n2210 vdd.n2179 10.6151
R4811 vdd.n2211 vdd.n2210 10.6151
R4812 vdd.n2213 vdd.n2175 10.6151
R4813 vdd.n2218 vdd.n2175 10.6151
R4814 vdd.n1851 vdd.t143 10.5435
R4815 vdd.n656 vdd.t252 10.5435
R4816 vdd.n316 vdd.n298 10.4732
R4817 vdd.n257 vdd.n239 10.4732
R4818 vdd.n214 vdd.n196 10.4732
R4819 vdd.n155 vdd.n137 10.4732
R4820 vdd.n113 vdd.n95 10.4732
R4821 vdd.n54 vdd.n36 10.4732
R4822 vdd.n1735 vdd.n1717 10.4732
R4823 vdd.n1794 vdd.n1776 10.4732
R4824 vdd.n1633 vdd.n1615 10.4732
R4825 vdd.n1692 vdd.n1674 10.4732
R4826 vdd.n1532 vdd.n1514 10.4732
R4827 vdd.n1591 vdd.n1573 10.4732
R4828 vdd.t230 vdd.n1825 10.3167
R4829 vdd.n3300 vdd.t192 10.3167
R4830 vdd.n1502 vdd.t160 10.09
R4831 vdd.n3394 vdd.t158 10.09
R4832 vdd.t226 vdd.n1155 9.86327
R4833 vdd.n3385 vdd.t135 9.86327
R4834 vdd.n315 vdd.n300 9.69747
R4835 vdd.n256 vdd.n241 9.69747
R4836 vdd.n213 vdd.n198 9.69747
R4837 vdd.n154 vdd.n139 9.69747
R4838 vdd.n112 vdd.n97 9.69747
R4839 vdd.n53 vdd.n38 9.69747
R4840 vdd.n1734 vdd.n1719 9.69747
R4841 vdd.n1793 vdd.n1778 9.69747
R4842 vdd.n1632 vdd.n1617 9.69747
R4843 vdd.n1691 vdd.n1676 9.69747
R4844 vdd.n1531 vdd.n1516 9.69747
R4845 vdd.n1590 vdd.n1575 9.69747
R4846 vdd.n2315 vdd.n2314 9.67831
R4847 vdd.n3216 vdd.n731 9.67831
R4848 vdd.n3093 vdd.n3092 9.67831
R4849 vdd.n2339 vdd.n2338 9.67831
R4850 vdd.n1461 vdd.t176 9.63654
R4851 vdd.n3331 vdd.t156 9.63654
R4852 vdd.n331 vdd.n330 9.45567
R4853 vdd.n272 vdd.n271 9.45567
R4854 vdd.n229 vdd.n228 9.45567
R4855 vdd.n170 vdd.n169 9.45567
R4856 vdd.n128 vdd.n127 9.45567
R4857 vdd.n69 vdd.n68 9.45567
R4858 vdd.n1750 vdd.n1749 9.45567
R4859 vdd.n1809 vdd.n1808 9.45567
R4860 vdd.n1648 vdd.n1647 9.45567
R4861 vdd.n1707 vdd.n1706 9.45567
R4862 vdd.n1547 vdd.n1546 9.45567
R4863 vdd.n1606 vdd.n1605 9.45567
R4864 vdd.n1435 vdd.t145 9.40981
R4865 vdd.n3363 vdd.t199 9.40981
R4866 vdd.n2075 vdd.n1929 9.3005
R4867 vdd.n2074 vdd.n2073 9.3005
R4868 vdd.n1935 vdd.n1934 9.3005
R4869 vdd.n2068 vdd.n1939 9.3005
R4870 vdd.n2067 vdd.n1940 9.3005
R4871 vdd.n2066 vdd.n1941 9.3005
R4872 vdd.n1945 vdd.n1942 9.3005
R4873 vdd.n2061 vdd.n1946 9.3005
R4874 vdd.n2060 vdd.n1947 9.3005
R4875 vdd.n2059 vdd.n1948 9.3005
R4876 vdd.n1952 vdd.n1949 9.3005
R4877 vdd.n2054 vdd.n1953 9.3005
R4878 vdd.n2053 vdd.n1954 9.3005
R4879 vdd.n2052 vdd.n1955 9.3005
R4880 vdd.n1959 vdd.n1956 9.3005
R4881 vdd.n2047 vdd.n1960 9.3005
R4882 vdd.n2046 vdd.n1961 9.3005
R4883 vdd.n2045 vdd.n1962 9.3005
R4884 vdd.n1966 vdd.n1963 9.3005
R4885 vdd.n2040 vdd.n1967 9.3005
R4886 vdd.n2039 vdd.n1968 9.3005
R4887 vdd.n2038 vdd.n2037 9.3005
R4888 vdd.n2036 vdd.n1969 9.3005
R4889 vdd.n2035 vdd.n2034 9.3005
R4890 vdd.n1975 vdd.n1974 9.3005
R4891 vdd.n2029 vdd.n1979 9.3005
R4892 vdd.n2028 vdd.n1980 9.3005
R4893 vdd.n2027 vdd.n1981 9.3005
R4894 vdd.n1985 vdd.n1982 9.3005
R4895 vdd.n2022 vdd.n1986 9.3005
R4896 vdd.n2021 vdd.n1987 9.3005
R4897 vdd.n2020 vdd.n1988 9.3005
R4898 vdd.n1992 vdd.n1989 9.3005
R4899 vdd.n2015 vdd.n1993 9.3005
R4900 vdd.n2014 vdd.n1994 9.3005
R4901 vdd.n2013 vdd.n1995 9.3005
R4902 vdd.n1997 vdd.n1996 9.3005
R4903 vdd.n2008 vdd.n1064 9.3005
R4904 vdd.n2077 vdd.n2076 9.3005
R4905 vdd.n2101 vdd.n2100 9.3005
R4906 vdd.n1907 vdd.n1906 9.3005
R4907 vdd.n1912 vdd.n1910 9.3005
R4908 vdd.n2093 vdd.n1913 9.3005
R4909 vdd.n2092 vdd.n1914 9.3005
R4910 vdd.n2091 vdd.n1915 9.3005
R4911 vdd.n1919 vdd.n1916 9.3005
R4912 vdd.n2086 vdd.n1920 9.3005
R4913 vdd.n2085 vdd.n1921 9.3005
R4914 vdd.n2084 vdd.n1922 9.3005
R4915 vdd.n1926 vdd.n1923 9.3005
R4916 vdd.n2079 vdd.n1927 9.3005
R4917 vdd.n2078 vdd.n1928 9.3005
R4918 vdd.n2323 vdd.n1900 9.3005
R4919 vdd.n2325 vdd.n2324 9.3005
R4920 vdd.n1815 vdd.n1814 9.3005
R4921 vdd.n1124 vdd.n1123 9.3005
R4922 vdd.n1829 vdd.n1828 9.3005
R4923 vdd.n1830 vdd.n1122 9.3005
R4924 vdd.n1832 vdd.n1831 9.3005
R4925 vdd.n1113 vdd.n1112 9.3005
R4926 vdd.n1846 vdd.n1845 9.3005
R4927 vdd.n1847 vdd.n1111 9.3005
R4928 vdd.n1849 vdd.n1848 9.3005
R4929 vdd.n1102 vdd.n1101 9.3005
R4930 vdd.n1862 vdd.n1861 9.3005
R4931 vdd.n1863 vdd.n1100 9.3005
R4932 vdd.n1865 vdd.n1864 9.3005
R4933 vdd.n1090 vdd.n1089 9.3005
R4934 vdd.n1879 vdd.n1878 9.3005
R4935 vdd.n1880 vdd.n1088 9.3005
R4936 vdd.n1882 vdd.n1881 9.3005
R4937 vdd.n1078 vdd.n1077 9.3005
R4938 vdd.n1898 vdd.n1897 9.3005
R4939 vdd.n1899 vdd.n1076 9.3005
R4940 vdd.n2327 vdd.n2326 9.3005
R4941 vdd.n307 vdd.n306 9.3005
R4942 vdd.n302 vdd.n301 9.3005
R4943 vdd.n313 vdd.n312 9.3005
R4944 vdd.n315 vdd.n314 9.3005
R4945 vdd.n298 vdd.n297 9.3005
R4946 vdd.n321 vdd.n320 9.3005
R4947 vdd.n323 vdd.n322 9.3005
R4948 vdd.n295 vdd.n292 9.3005
R4949 vdd.n330 vdd.n329 9.3005
R4950 vdd.n248 vdd.n247 9.3005
R4951 vdd.n243 vdd.n242 9.3005
R4952 vdd.n254 vdd.n253 9.3005
R4953 vdd.n256 vdd.n255 9.3005
R4954 vdd.n239 vdd.n238 9.3005
R4955 vdd.n262 vdd.n261 9.3005
R4956 vdd.n264 vdd.n263 9.3005
R4957 vdd.n236 vdd.n233 9.3005
R4958 vdd.n271 vdd.n270 9.3005
R4959 vdd.n205 vdd.n204 9.3005
R4960 vdd.n200 vdd.n199 9.3005
R4961 vdd.n211 vdd.n210 9.3005
R4962 vdd.n213 vdd.n212 9.3005
R4963 vdd.n196 vdd.n195 9.3005
R4964 vdd.n219 vdd.n218 9.3005
R4965 vdd.n221 vdd.n220 9.3005
R4966 vdd.n193 vdd.n190 9.3005
R4967 vdd.n228 vdd.n227 9.3005
R4968 vdd.n146 vdd.n145 9.3005
R4969 vdd.n141 vdd.n140 9.3005
R4970 vdd.n152 vdd.n151 9.3005
R4971 vdd.n154 vdd.n153 9.3005
R4972 vdd.n137 vdd.n136 9.3005
R4973 vdd.n160 vdd.n159 9.3005
R4974 vdd.n162 vdd.n161 9.3005
R4975 vdd.n134 vdd.n131 9.3005
R4976 vdd.n169 vdd.n168 9.3005
R4977 vdd.n104 vdd.n103 9.3005
R4978 vdd.n99 vdd.n98 9.3005
R4979 vdd.n110 vdd.n109 9.3005
R4980 vdd.n112 vdd.n111 9.3005
R4981 vdd.n95 vdd.n94 9.3005
R4982 vdd.n118 vdd.n117 9.3005
R4983 vdd.n120 vdd.n119 9.3005
R4984 vdd.n92 vdd.n89 9.3005
R4985 vdd.n127 vdd.n126 9.3005
R4986 vdd.n45 vdd.n44 9.3005
R4987 vdd.n40 vdd.n39 9.3005
R4988 vdd.n51 vdd.n50 9.3005
R4989 vdd.n53 vdd.n52 9.3005
R4990 vdd.n36 vdd.n35 9.3005
R4991 vdd.n59 vdd.n58 9.3005
R4992 vdd.n61 vdd.n60 9.3005
R4993 vdd.n33 vdd.n30 9.3005
R4994 vdd.n68 vdd.n67 9.3005
R4995 vdd.n3138 vdd.n3137 9.3005
R4996 vdd.n3141 vdd.n766 9.3005
R4997 vdd.n3142 vdd.n765 9.3005
R4998 vdd.n3145 vdd.n764 9.3005
R4999 vdd.n3146 vdd.n763 9.3005
R5000 vdd.n3149 vdd.n762 9.3005
R5001 vdd.n3150 vdd.n761 9.3005
R5002 vdd.n3153 vdd.n760 9.3005
R5003 vdd.n3154 vdd.n759 9.3005
R5004 vdd.n3157 vdd.n758 9.3005
R5005 vdd.n3158 vdd.n757 9.3005
R5006 vdd.n3161 vdd.n756 9.3005
R5007 vdd.n3162 vdd.n755 9.3005
R5008 vdd.n3165 vdd.n754 9.3005
R5009 vdd.n3166 vdd.n753 9.3005
R5010 vdd.n3169 vdd.n752 9.3005
R5011 vdd.n3170 vdd.n751 9.3005
R5012 vdd.n3173 vdd.n750 9.3005
R5013 vdd.n3174 vdd.n749 9.3005
R5014 vdd.n3177 vdd.n748 9.3005
R5015 vdd.n3181 vdd.n3180 9.3005
R5016 vdd.n3182 vdd.n747 9.3005
R5017 vdd.n3186 vdd.n3183 9.3005
R5018 vdd.n3189 vdd.n746 9.3005
R5019 vdd.n3190 vdd.n745 9.3005
R5020 vdd.n3193 vdd.n744 9.3005
R5021 vdd.n3194 vdd.n743 9.3005
R5022 vdd.n3197 vdd.n742 9.3005
R5023 vdd.n3198 vdd.n741 9.3005
R5024 vdd.n3201 vdd.n740 9.3005
R5025 vdd.n3202 vdd.n739 9.3005
R5026 vdd.n3205 vdd.n738 9.3005
R5027 vdd.n3206 vdd.n737 9.3005
R5028 vdd.n3209 vdd.n736 9.3005
R5029 vdd.n3210 vdd.n735 9.3005
R5030 vdd.n3213 vdd.n730 9.3005
R5031 vdd.n3219 vdd.n727 9.3005
R5032 vdd.n3220 vdd.n726 9.3005
R5033 vdd.n3234 vdd.n3233 9.3005
R5034 vdd.n3235 vdd.n681 9.3005
R5035 vdd.n3237 vdd.n3236 9.3005
R5036 vdd.n671 vdd.n670 9.3005
R5037 vdd.n3251 vdd.n3250 9.3005
R5038 vdd.n3252 vdd.n669 9.3005
R5039 vdd.n3254 vdd.n3253 9.3005
R5040 vdd.n660 vdd.n659 9.3005
R5041 vdd.n3267 vdd.n3266 9.3005
R5042 vdd.n3268 vdd.n658 9.3005
R5043 vdd.n3270 vdd.n3269 9.3005
R5044 vdd.n648 vdd.n647 9.3005
R5045 vdd.n3284 vdd.n3283 9.3005
R5046 vdd.n3285 vdd.n646 9.3005
R5047 vdd.n3287 vdd.n3286 9.3005
R5048 vdd.n637 vdd.n636 9.3005
R5049 vdd.n3303 vdd.n3302 9.3005
R5050 vdd.n3304 vdd.n635 9.3005
R5051 vdd.n3306 vdd.n3305 9.3005
R5052 vdd.n336 vdd.n334 9.3005
R5053 vdd.n683 vdd.n682 9.3005
R5054 vdd.n3398 vdd.n3397 9.3005
R5055 vdd.n337 vdd.n335 9.3005
R5056 vdd.n3391 vdd.n346 9.3005
R5057 vdd.n3390 vdd.n347 9.3005
R5058 vdd.n3389 vdd.n348 9.3005
R5059 vdd.n355 vdd.n349 9.3005
R5060 vdd.n3383 vdd.n356 9.3005
R5061 vdd.n3382 vdd.n357 9.3005
R5062 vdd.n3381 vdd.n358 9.3005
R5063 vdd.n366 vdd.n359 9.3005
R5064 vdd.n3375 vdd.n367 9.3005
R5065 vdd.n3374 vdd.n368 9.3005
R5066 vdd.n3373 vdd.n369 9.3005
R5067 vdd.n377 vdd.n370 9.3005
R5068 vdd.n3367 vdd.n378 9.3005
R5069 vdd.n3366 vdd.n379 9.3005
R5070 vdd.n3365 vdd.n380 9.3005
R5071 vdd.n388 vdd.n381 9.3005
R5072 vdd.n3359 vdd.n389 9.3005
R5073 vdd.n3358 vdd.n390 9.3005
R5074 vdd.n3357 vdd.n391 9.3005
R5075 vdd.n466 vdd.n463 9.3005
R5076 vdd.n470 vdd.n469 9.3005
R5077 vdd.n471 vdd.n462 9.3005
R5078 vdd.n475 vdd.n472 9.3005
R5079 vdd.n476 vdd.n461 9.3005
R5080 vdd.n480 vdd.n479 9.3005
R5081 vdd.n481 vdd.n460 9.3005
R5082 vdd.n485 vdd.n482 9.3005
R5083 vdd.n486 vdd.n459 9.3005
R5084 vdd.n490 vdd.n489 9.3005
R5085 vdd.n491 vdd.n458 9.3005
R5086 vdd.n495 vdd.n492 9.3005
R5087 vdd.n496 vdd.n457 9.3005
R5088 vdd.n500 vdd.n499 9.3005
R5089 vdd.n501 vdd.n456 9.3005
R5090 vdd.n505 vdd.n502 9.3005
R5091 vdd.n506 vdd.n455 9.3005
R5092 vdd.n510 vdd.n509 9.3005
R5093 vdd.n511 vdd.n454 9.3005
R5094 vdd.n515 vdd.n512 9.3005
R5095 vdd.n516 vdd.n451 9.3005
R5096 vdd.n520 vdd.n519 9.3005
R5097 vdd.n521 vdd.n450 9.3005
R5098 vdd.n525 vdd.n522 9.3005
R5099 vdd.n526 vdd.n449 9.3005
R5100 vdd.n530 vdd.n529 9.3005
R5101 vdd.n531 vdd.n448 9.3005
R5102 vdd.n535 vdd.n532 9.3005
R5103 vdd.n536 vdd.n447 9.3005
R5104 vdd.n540 vdd.n539 9.3005
R5105 vdd.n541 vdd.n446 9.3005
R5106 vdd.n545 vdd.n542 9.3005
R5107 vdd.n546 vdd.n445 9.3005
R5108 vdd.n550 vdd.n549 9.3005
R5109 vdd.n551 vdd.n444 9.3005
R5110 vdd.n555 vdd.n552 9.3005
R5111 vdd.n556 vdd.n443 9.3005
R5112 vdd.n560 vdd.n559 9.3005
R5113 vdd.n561 vdd.n442 9.3005
R5114 vdd.n565 vdd.n562 9.3005
R5115 vdd.n566 vdd.n439 9.3005
R5116 vdd.n570 vdd.n569 9.3005
R5117 vdd.n571 vdd.n438 9.3005
R5118 vdd.n575 vdd.n572 9.3005
R5119 vdd.n576 vdd.n437 9.3005
R5120 vdd.n580 vdd.n579 9.3005
R5121 vdd.n581 vdd.n436 9.3005
R5122 vdd.n585 vdd.n582 9.3005
R5123 vdd.n586 vdd.n435 9.3005
R5124 vdd.n590 vdd.n589 9.3005
R5125 vdd.n591 vdd.n434 9.3005
R5126 vdd.n595 vdd.n592 9.3005
R5127 vdd.n596 vdd.n433 9.3005
R5128 vdd.n600 vdd.n599 9.3005
R5129 vdd.n601 vdd.n432 9.3005
R5130 vdd.n605 vdd.n602 9.3005
R5131 vdd.n606 vdd.n431 9.3005
R5132 vdd.n610 vdd.n609 9.3005
R5133 vdd.n611 vdd.n430 9.3005
R5134 vdd.n615 vdd.n612 9.3005
R5135 vdd.n617 vdd.n429 9.3005
R5136 vdd.n619 vdd.n618 9.3005
R5137 vdd.n3351 vdd.n3350 9.3005
R5138 vdd.n465 vdd.n464 9.3005
R5139 vdd.n3229 vdd.n3228 9.3005
R5140 vdd.n676 vdd.n675 9.3005
R5141 vdd.n3242 vdd.n3241 9.3005
R5142 vdd.n3243 vdd.n674 9.3005
R5143 vdd.n3245 vdd.n3244 9.3005
R5144 vdd.n666 vdd.n665 9.3005
R5145 vdd.n3259 vdd.n3258 9.3005
R5146 vdd.n3260 vdd.n664 9.3005
R5147 vdd.n3262 vdd.n3261 9.3005
R5148 vdd.n653 vdd.n652 9.3005
R5149 vdd.n3275 vdd.n3274 9.3005
R5150 vdd.n3276 vdd.n651 9.3005
R5151 vdd.n3278 vdd.n3277 9.3005
R5152 vdd.n642 vdd.n641 9.3005
R5153 vdd.n3292 vdd.n3291 9.3005
R5154 vdd.n3293 vdd.n640 9.3005
R5155 vdd.n3298 vdd.n3294 9.3005
R5156 vdd.n3297 vdd.n3296 9.3005
R5157 vdd.n3295 vdd.n631 9.3005
R5158 vdd.n3311 vdd.n630 9.3005
R5159 vdd.n3313 vdd.n3312 9.3005
R5160 vdd.n3314 vdd.n629 9.3005
R5161 vdd.n3316 vdd.n3315 9.3005
R5162 vdd.n3318 vdd.n628 9.3005
R5163 vdd.n3320 vdd.n3319 9.3005
R5164 vdd.n3321 vdd.n627 9.3005
R5165 vdd.n3323 vdd.n3322 9.3005
R5166 vdd.n3325 vdd.n626 9.3005
R5167 vdd.n3327 vdd.n3326 9.3005
R5168 vdd.n3328 vdd.n625 9.3005
R5169 vdd.n3330 vdd.n3329 9.3005
R5170 vdd.n3333 vdd.n624 9.3005
R5171 vdd.n3335 vdd.n3334 9.3005
R5172 vdd.n3336 vdd.n623 9.3005
R5173 vdd.n3338 vdd.n3337 9.3005
R5174 vdd.n3340 vdd.n622 9.3005
R5175 vdd.n3342 vdd.n3341 9.3005
R5176 vdd.n3343 vdd.n621 9.3005
R5177 vdd.n3345 vdd.n3344 9.3005
R5178 vdd.n3347 vdd.n620 9.3005
R5179 vdd.n3349 vdd.n3348 9.3005
R5180 vdd.n3227 vdd.n686 9.3005
R5181 vdd.n3226 vdd.n3225 9.3005
R5182 vdd.n3095 vdd.n687 9.3005
R5183 vdd.n3104 vdd.n783 9.3005
R5184 vdd.n3107 vdd.n782 9.3005
R5185 vdd.n3108 vdd.n781 9.3005
R5186 vdd.n3111 vdd.n780 9.3005
R5187 vdd.n3112 vdd.n779 9.3005
R5188 vdd.n3115 vdd.n778 9.3005
R5189 vdd.n3116 vdd.n777 9.3005
R5190 vdd.n3119 vdd.n776 9.3005
R5191 vdd.n3120 vdd.n775 9.3005
R5192 vdd.n3123 vdd.n774 9.3005
R5193 vdd.n3124 vdd.n773 9.3005
R5194 vdd.n3127 vdd.n772 9.3005
R5195 vdd.n3128 vdd.n771 9.3005
R5196 vdd.n3131 vdd.n770 9.3005
R5197 vdd.n3135 vdd.n3134 9.3005
R5198 vdd.n3136 vdd.n767 9.3005
R5199 vdd.n2337 vdd.n2336 9.3005
R5200 vdd.n2332 vdd.n1067 9.3005
R5201 vdd.n1430 vdd.n1429 9.3005
R5202 vdd.n1431 vdd.n1185 9.3005
R5203 vdd.n1433 vdd.n1432 9.3005
R5204 vdd.n1175 vdd.n1174 9.3005
R5205 vdd.n1447 vdd.n1446 9.3005
R5206 vdd.n1448 vdd.n1173 9.3005
R5207 vdd.n1450 vdd.n1449 9.3005
R5208 vdd.n1165 vdd.n1164 9.3005
R5209 vdd.n1464 vdd.n1463 9.3005
R5210 vdd.n1465 vdd.n1163 9.3005
R5211 vdd.n1467 vdd.n1466 9.3005
R5212 vdd.n1152 vdd.n1151 9.3005
R5213 vdd.n1480 vdd.n1479 9.3005
R5214 vdd.n1481 vdd.n1150 9.3005
R5215 vdd.n1483 vdd.n1482 9.3005
R5216 vdd.n1141 vdd.n1140 9.3005
R5217 vdd.n1497 vdd.n1496 9.3005
R5218 vdd.n1498 vdd.n1139 9.3005
R5219 vdd.n1500 vdd.n1499 9.3005
R5220 vdd.n1130 vdd.n1129 9.3005
R5221 vdd.n1820 vdd.n1819 9.3005
R5222 vdd.n1821 vdd.n1128 9.3005
R5223 vdd.n1823 vdd.n1822 9.3005
R5224 vdd.n1118 vdd.n1117 9.3005
R5225 vdd.n1837 vdd.n1836 9.3005
R5226 vdd.n1838 vdd.n1116 9.3005
R5227 vdd.n1840 vdd.n1839 9.3005
R5228 vdd.n1108 vdd.n1107 9.3005
R5229 vdd.n1854 vdd.n1853 9.3005
R5230 vdd.n1855 vdd.n1106 9.3005
R5231 vdd.n1857 vdd.n1856 9.3005
R5232 vdd.n1095 vdd.n1094 9.3005
R5233 vdd.n1870 vdd.n1869 9.3005
R5234 vdd.n1871 vdd.n1093 9.3005
R5235 vdd.n1873 vdd.n1872 9.3005
R5236 vdd.n1085 vdd.n1084 9.3005
R5237 vdd.n1887 vdd.n1886 9.3005
R5238 vdd.n1888 vdd.n1082 9.3005
R5239 vdd.n1892 vdd.n1891 9.3005
R5240 vdd.n1890 vdd.n1083 9.3005
R5241 vdd.n1889 vdd.n1072 9.3005
R5242 vdd.n1187 vdd.n1186 9.3005
R5243 vdd.n1323 vdd.n1322 9.3005
R5244 vdd.n1324 vdd.n1313 9.3005
R5245 vdd.n1326 vdd.n1325 9.3005
R5246 vdd.n1327 vdd.n1312 9.3005
R5247 vdd.n1329 vdd.n1328 9.3005
R5248 vdd.n1330 vdd.n1307 9.3005
R5249 vdd.n1332 vdd.n1331 9.3005
R5250 vdd.n1333 vdd.n1306 9.3005
R5251 vdd.n1335 vdd.n1334 9.3005
R5252 vdd.n1336 vdd.n1301 9.3005
R5253 vdd.n1338 vdd.n1337 9.3005
R5254 vdd.n1339 vdd.n1300 9.3005
R5255 vdd.n1341 vdd.n1340 9.3005
R5256 vdd.n1342 vdd.n1295 9.3005
R5257 vdd.n1344 vdd.n1343 9.3005
R5258 vdd.n1345 vdd.n1294 9.3005
R5259 vdd.n1347 vdd.n1346 9.3005
R5260 vdd.n1348 vdd.n1289 9.3005
R5261 vdd.n1350 vdd.n1349 9.3005
R5262 vdd.n1351 vdd.n1288 9.3005
R5263 vdd.n1353 vdd.n1352 9.3005
R5264 vdd.n1357 vdd.n1284 9.3005
R5265 vdd.n1359 vdd.n1358 9.3005
R5266 vdd.n1360 vdd.n1283 9.3005
R5267 vdd.n1362 vdd.n1361 9.3005
R5268 vdd.n1363 vdd.n1278 9.3005
R5269 vdd.n1365 vdd.n1364 9.3005
R5270 vdd.n1366 vdd.n1277 9.3005
R5271 vdd.n1368 vdd.n1367 9.3005
R5272 vdd.n1369 vdd.n1272 9.3005
R5273 vdd.n1371 vdd.n1370 9.3005
R5274 vdd.n1372 vdd.n1271 9.3005
R5275 vdd.n1374 vdd.n1373 9.3005
R5276 vdd.n1375 vdd.n1266 9.3005
R5277 vdd.n1377 vdd.n1376 9.3005
R5278 vdd.n1378 vdd.n1265 9.3005
R5279 vdd.n1380 vdd.n1379 9.3005
R5280 vdd.n1381 vdd.n1260 9.3005
R5281 vdd.n1383 vdd.n1382 9.3005
R5282 vdd.n1384 vdd.n1259 9.3005
R5283 vdd.n1386 vdd.n1385 9.3005
R5284 vdd.n1387 vdd.n1254 9.3005
R5285 vdd.n1389 vdd.n1388 9.3005
R5286 vdd.n1390 vdd.n1253 9.3005
R5287 vdd.n1392 vdd.n1391 9.3005
R5288 vdd.n1393 vdd.n1246 9.3005
R5289 vdd.n1395 vdd.n1394 9.3005
R5290 vdd.n1396 vdd.n1245 9.3005
R5291 vdd.n1398 vdd.n1397 9.3005
R5292 vdd.n1399 vdd.n1240 9.3005
R5293 vdd.n1401 vdd.n1400 9.3005
R5294 vdd.n1402 vdd.n1239 9.3005
R5295 vdd.n1404 vdd.n1403 9.3005
R5296 vdd.n1405 vdd.n1234 9.3005
R5297 vdd.n1407 vdd.n1406 9.3005
R5298 vdd.n1408 vdd.n1233 9.3005
R5299 vdd.n1410 vdd.n1409 9.3005
R5300 vdd.n1411 vdd.n1228 9.3005
R5301 vdd.n1413 vdd.n1412 9.3005
R5302 vdd.n1414 vdd.n1227 9.3005
R5303 vdd.n1416 vdd.n1415 9.3005
R5304 vdd.n1192 vdd.n1191 9.3005
R5305 vdd.n1422 vdd.n1421 9.3005
R5306 vdd.n1321 vdd.n1320 9.3005
R5307 vdd.n1425 vdd.n1424 9.3005
R5308 vdd.n1181 vdd.n1180 9.3005
R5309 vdd.n1439 vdd.n1438 9.3005
R5310 vdd.n1440 vdd.n1179 9.3005
R5311 vdd.n1442 vdd.n1441 9.3005
R5312 vdd.n1170 vdd.n1169 9.3005
R5313 vdd.n1456 vdd.n1455 9.3005
R5314 vdd.n1457 vdd.n1168 9.3005
R5315 vdd.n1459 vdd.n1458 9.3005
R5316 vdd.n1159 vdd.n1158 9.3005
R5317 vdd.n1472 vdd.n1471 9.3005
R5318 vdd.n1473 vdd.n1157 9.3005
R5319 vdd.n1475 vdd.n1474 9.3005
R5320 vdd.n1147 vdd.n1146 9.3005
R5321 vdd.n1489 vdd.n1488 9.3005
R5322 vdd.n1490 vdd.n1145 9.3005
R5323 vdd.n1492 vdd.n1491 9.3005
R5324 vdd.n1136 vdd.n1135 9.3005
R5325 vdd.n1505 vdd.n1504 9.3005
R5326 vdd.n1506 vdd.n1134 9.3005
R5327 vdd.n1423 vdd.n1190 9.3005
R5328 vdd.n1726 vdd.n1725 9.3005
R5329 vdd.n1721 vdd.n1720 9.3005
R5330 vdd.n1732 vdd.n1731 9.3005
R5331 vdd.n1734 vdd.n1733 9.3005
R5332 vdd.n1717 vdd.n1716 9.3005
R5333 vdd.n1740 vdd.n1739 9.3005
R5334 vdd.n1742 vdd.n1741 9.3005
R5335 vdd.n1714 vdd.n1711 9.3005
R5336 vdd.n1749 vdd.n1748 9.3005
R5337 vdd.n1785 vdd.n1784 9.3005
R5338 vdd.n1780 vdd.n1779 9.3005
R5339 vdd.n1791 vdd.n1790 9.3005
R5340 vdd.n1793 vdd.n1792 9.3005
R5341 vdd.n1776 vdd.n1775 9.3005
R5342 vdd.n1799 vdd.n1798 9.3005
R5343 vdd.n1801 vdd.n1800 9.3005
R5344 vdd.n1773 vdd.n1770 9.3005
R5345 vdd.n1808 vdd.n1807 9.3005
R5346 vdd.n1624 vdd.n1623 9.3005
R5347 vdd.n1619 vdd.n1618 9.3005
R5348 vdd.n1630 vdd.n1629 9.3005
R5349 vdd.n1632 vdd.n1631 9.3005
R5350 vdd.n1615 vdd.n1614 9.3005
R5351 vdd.n1638 vdd.n1637 9.3005
R5352 vdd.n1640 vdd.n1639 9.3005
R5353 vdd.n1612 vdd.n1609 9.3005
R5354 vdd.n1647 vdd.n1646 9.3005
R5355 vdd.n1683 vdd.n1682 9.3005
R5356 vdd.n1678 vdd.n1677 9.3005
R5357 vdd.n1689 vdd.n1688 9.3005
R5358 vdd.n1691 vdd.n1690 9.3005
R5359 vdd.n1674 vdd.n1673 9.3005
R5360 vdd.n1697 vdd.n1696 9.3005
R5361 vdd.n1699 vdd.n1698 9.3005
R5362 vdd.n1671 vdd.n1668 9.3005
R5363 vdd.n1706 vdd.n1705 9.3005
R5364 vdd.n1523 vdd.n1522 9.3005
R5365 vdd.n1518 vdd.n1517 9.3005
R5366 vdd.n1529 vdd.n1528 9.3005
R5367 vdd.n1531 vdd.n1530 9.3005
R5368 vdd.n1514 vdd.n1513 9.3005
R5369 vdd.n1537 vdd.n1536 9.3005
R5370 vdd.n1539 vdd.n1538 9.3005
R5371 vdd.n1511 vdd.n1508 9.3005
R5372 vdd.n1546 vdd.n1545 9.3005
R5373 vdd.n1582 vdd.n1581 9.3005
R5374 vdd.n1577 vdd.n1576 9.3005
R5375 vdd.n1588 vdd.n1587 9.3005
R5376 vdd.n1590 vdd.n1589 9.3005
R5377 vdd.n1573 vdd.n1572 9.3005
R5378 vdd.n1596 vdd.n1595 9.3005
R5379 vdd.n1598 vdd.n1597 9.3005
R5380 vdd.n1570 vdd.n1567 9.3005
R5381 vdd.n1605 vdd.n1604 9.3005
R5382 vdd.n1461 vdd.t174 9.18308
R5383 vdd.n3331 vdd.t244 9.18308
R5384 vdd.n1155 vdd.t224 8.95635
R5385 vdd.n2329 vdd.t23 8.95635
R5386 vdd.n723 vdd.t16 8.95635
R5387 vdd.t188 vdd.n3385 8.95635
R5388 vdd.n312 vdd.n311 8.92171
R5389 vdd.n253 vdd.n252 8.92171
R5390 vdd.n210 vdd.n209 8.92171
R5391 vdd.n151 vdd.n150 8.92171
R5392 vdd.n109 vdd.n108 8.92171
R5393 vdd.n50 vdd.n49 8.92171
R5394 vdd.n1731 vdd.n1730 8.92171
R5395 vdd.n1790 vdd.n1789 8.92171
R5396 vdd.n1629 vdd.n1628 8.92171
R5397 vdd.n1688 vdd.n1687 8.92171
R5398 vdd.n1528 vdd.n1527 8.92171
R5399 vdd.n1587 vdd.n1586 8.92171
R5400 vdd.n231 vdd.n129 8.81535
R5401 vdd.n1709 vdd.n1607 8.81535
R5402 vdd.n1502 vdd.t196 8.72962
R5403 vdd.t185 vdd.n3394 8.72962
R5404 vdd.n1825 vdd.t247 8.50289
R5405 vdd.n3300 vdd.t190 8.50289
R5406 vdd.n28 vdd.n14 8.42249
R5407 vdd.n1851 vdd.t183 8.27616
R5408 vdd.t181 vdd.n656 8.27616
R5409 vdd.n3400 vdd.n3399 8.16225
R5410 vdd.n1813 vdd.n1812 8.16225
R5411 vdd.n308 vdd.n302 8.14595
R5412 vdd.n249 vdd.n243 8.14595
R5413 vdd.n206 vdd.n200 8.14595
R5414 vdd.n147 vdd.n141 8.14595
R5415 vdd.n105 vdd.n99 8.14595
R5416 vdd.n46 vdd.n40 8.14595
R5417 vdd.n1727 vdd.n1721 8.14595
R5418 vdd.n1786 vdd.n1780 8.14595
R5419 vdd.n1625 vdd.n1619 8.14595
R5420 vdd.n1684 vdd.n1678 8.14595
R5421 vdd.n1524 vdd.n1518 8.14595
R5422 vdd.n1583 vdd.n1577 8.14595
R5423 vdd.n2923 vdd.n849 8.11757
R5424 vdd.n2397 vdd.n2396 8.11757
R5425 vdd.n1098 vdd.t269 8.04943
R5426 vdd.n3256 vdd.t222 8.04943
R5427 vdd.n2375 vdd.n1043 7.70933
R5428 vdd.n2381 vdd.n1043 7.70933
R5429 vdd.n2387 vdd.n1037 7.70933
R5430 vdd.n2387 vdd.n1030 7.70933
R5431 vdd.n2393 vdd.n1030 7.70933
R5432 vdd.n2393 vdd.n1033 7.70933
R5433 vdd.n2400 vdd.n1018 7.70933
R5434 vdd.n2406 vdd.n1018 7.70933
R5435 vdd.n2412 vdd.n1012 7.70933
R5436 vdd.n2418 vdd.n1008 7.70933
R5437 vdd.n2424 vdd.n1002 7.70933
R5438 vdd.n2436 vdd.n989 7.70933
R5439 vdd.n2442 vdd.n983 7.70933
R5440 vdd.n2442 vdd.n976 7.70933
R5441 vdd.n2450 vdd.n976 7.70933
R5442 vdd.n2457 vdd.t109 7.70933
R5443 vdd.n2532 vdd.t109 7.70933
R5444 vdd.n2864 vdd.t119 7.70933
R5445 vdd.n2870 vdd.t119 7.70933
R5446 vdd.n2876 vdd.n897 7.70933
R5447 vdd.n2882 vdd.n897 7.70933
R5448 vdd.n2882 vdd.n900 7.70933
R5449 vdd.n2888 vdd.n893 7.70933
R5450 vdd.n2900 vdd.n880 7.70933
R5451 vdd.n2906 vdd.n874 7.70933
R5452 vdd.n2912 vdd.n870 7.70933
R5453 vdd.n2918 vdd.n857 7.70933
R5454 vdd.n2926 vdd.n857 7.70933
R5455 vdd.n2932 vdd.n851 7.70933
R5456 vdd.n2932 vdd.n843 7.70933
R5457 vdd.n2983 vdd.n843 7.70933
R5458 vdd.n2983 vdd.n846 7.70933
R5459 vdd.n2989 vdd.n805 7.70933
R5460 vdd.n3059 vdd.n805 7.70933
R5461 vdd.n307 vdd.n304 7.3702
R5462 vdd.n248 vdd.n245 7.3702
R5463 vdd.n205 vdd.n202 7.3702
R5464 vdd.n146 vdd.n143 7.3702
R5465 vdd.n104 vdd.n101 7.3702
R5466 vdd.n45 vdd.n42 7.3702
R5467 vdd.n1726 vdd.n1723 7.3702
R5468 vdd.n1785 vdd.n1782 7.3702
R5469 vdd.n1624 vdd.n1621 7.3702
R5470 vdd.n1683 vdd.n1680 7.3702
R5471 vdd.n1523 vdd.n1520 7.3702
R5472 vdd.n1582 vdd.n1579 7.3702
R5473 vdd.n1884 vdd.t141 7.1425
R5474 vdd.n679 vdd.t137 7.1425
R5475 vdd.n1358 vdd.n1357 6.98232
R5476 vdd.n2039 vdd.n2038 6.98232
R5477 vdd.n566 vdd.n565 6.98232
R5478 vdd.n3141 vdd.n3138 6.98232
R5479 vdd.t249 vdd.n1097 6.91577
R5480 vdd.n3264 vdd.t147 6.91577
R5481 vdd.n1843 vdd.t206 6.68904
R5482 vdd.n3280 vdd.t131 6.68904
R5483 vdd.t149 vdd.n1126 6.46231
R5484 vdd.n3308 vdd.t151 6.46231
R5485 vdd.n3400 vdd.n333 6.38151
R5486 vdd.n1812 vdd.n1811 6.38151
R5487 vdd.n1494 vdd.t178 6.23558
R5488 vdd.t218 vdd.n344 6.23558
R5489 vdd.t153 vdd.n1154 6.00885
R5490 vdd.n2412 vdd.t129 6.00885
R5491 vdd.n2912 vdd.t99 6.00885
R5492 vdd.n3379 vdd.t163 6.00885
R5493 vdd.n1033 vdd.t69 5.89549
R5494 vdd.t27 vdd.n851 5.89549
R5495 vdd.n308 vdd.n307 5.81868
R5496 vdd.n249 vdd.n248 5.81868
R5497 vdd.n206 vdd.n205 5.81868
R5498 vdd.n147 vdd.n146 5.81868
R5499 vdd.n105 vdd.n104 5.81868
R5500 vdd.n46 vdd.n45 5.81868
R5501 vdd.n1727 vdd.n1726 5.81868
R5502 vdd.n1786 vdd.n1785 5.81868
R5503 vdd.n1625 vdd.n1624 5.81868
R5504 vdd.n1684 vdd.n1683 5.81868
R5505 vdd.n1524 vdd.n1523 5.81868
R5506 vdd.n1583 vdd.n1582 5.81868
R5507 vdd.n1453 vdd.t139 5.78212
R5508 vdd.t12 vdd.n1037 5.78212
R5509 vdd.n2156 vdd.t51 5.78212
R5510 vdd.n2781 vdd.t59 5.78212
R5511 vdd.n846 vdd.t55 5.78212
R5512 vdd.n3370 vdd.t211 5.78212
R5513 vdd.n2540 vdd.n2539 5.77611
R5514 vdd.n2283 vdd.n2153 5.77611
R5515 vdd.n2794 vdd.n2793 5.77611
R5516 vdd.n3000 vdd.n2999 5.77611
R5517 vdd.n3064 vdd.n801 5.77611
R5518 vdd.n2704 vdd.n2644 5.77611
R5519 vdd.n2465 vdd.n967 5.77611
R5520 vdd.n2213 vdd.n2212 5.77611
R5521 vdd.n1320 vdd.n1319 5.62474
R5522 vdd.n2335 vdd.n2332 5.62474
R5523 vdd.n3351 vdd.n428 5.62474
R5524 vdd.n3225 vdd.n690 5.62474
R5525 vdd.n1177 vdd.t139 5.55539
R5526 vdd.t211 vdd.n3369 5.55539
R5527 vdd.t125 vdd.n989 5.44203
R5528 vdd.n893 vdd.t1 5.44203
R5529 vdd.n1469 vdd.t153 5.32866
R5530 vdd.t163 vdd.n3378 5.32866
R5531 vdd.n1485 vdd.t178 5.10193
R5532 vdd.t103 vdd.n1012 5.10193
R5533 vdd.n1002 vdd.t91 5.10193
R5534 vdd.t10 vdd.n880 5.10193
R5535 vdd.n870 vdd.t121 5.10193
R5536 vdd.n3387 vdd.t218 5.10193
R5537 vdd.n311 vdd.n302 5.04292
R5538 vdd.n252 vdd.n243 5.04292
R5539 vdd.n209 vdd.n200 5.04292
R5540 vdd.n150 vdd.n141 5.04292
R5541 vdd.n108 vdd.n99 5.04292
R5542 vdd.n49 vdd.n40 5.04292
R5543 vdd.n1730 vdd.n1721 5.04292
R5544 vdd.n1789 vdd.n1780 5.04292
R5545 vdd.n1628 vdd.n1619 5.04292
R5546 vdd.n1687 vdd.n1678 5.04292
R5547 vdd.n1527 vdd.n1518 5.04292
R5548 vdd.n1586 vdd.n1577 5.04292
R5549 vdd.n1817 vdd.t149 4.8752
R5550 vdd.t0 vdd.t92 4.8752
R5551 vdd.t112 vdd.t3 4.8752
R5552 vdd.t89 vdd.t124 4.8752
R5553 vdd.t122 vdd.t130 4.8752
R5554 vdd.t151 vdd.n340 4.8752
R5555 vdd.n2541 vdd.n2540 4.83952
R5556 vdd.n2153 vdd.n2149 4.83952
R5557 vdd.n2795 vdd.n2794 4.83952
R5558 vdd.n3001 vdd.n3000 4.83952
R5559 vdd.n801 vdd.n796 4.83952
R5560 vdd.n2701 vdd.n2644 4.83952
R5561 vdd.n2468 vdd.n967 4.83952
R5562 vdd.n2212 vdd.n2211 4.83952
R5563 vdd.n2007 vdd.n1065 4.74817
R5564 vdd.n2002 vdd.n1066 4.74817
R5565 vdd.n1904 vdd.n1901 4.74817
R5566 vdd.n2316 vdd.n1905 4.74817
R5567 vdd.n2318 vdd.n1904 4.74817
R5568 vdd.n2317 vdd.n2316 4.74817
R5569 vdd.n3218 vdd.n3217 4.74817
R5570 vdd.n3215 vdd.n3214 4.74817
R5571 vdd.n3215 vdd.n732 4.74817
R5572 vdd.n3217 vdd.n729 4.74817
R5573 vdd.n3100 vdd.n784 4.74817
R5574 vdd.n3096 vdd.n3094 4.74817
R5575 vdd.n3099 vdd.n3094 4.74817
R5576 vdd.n3103 vdd.n784 4.74817
R5577 vdd.n2003 vdd.n1065 4.74817
R5578 vdd.n1068 vdd.n1066 4.74817
R5579 vdd.n333 vdd.n332 4.7074
R5580 vdd.n231 vdd.n230 4.7074
R5581 vdd.n1811 vdd.n1810 4.7074
R5582 vdd.n1709 vdd.n1708 4.7074
R5583 vdd.n1120 vdd.t206 4.64847
R5584 vdd.n3289 vdd.t131 4.64847
R5585 vdd.n2418 vdd.t294 4.53511
R5586 vdd.n2906 vdd.t113 4.53511
R5587 vdd.n1859 vdd.t249 4.42174
R5588 vdd.t147 vdd.n655 4.42174
R5589 vdd.n2450 vdd.t127 4.30838
R5590 vdd.n2876 vdd.t97 4.30838
R5591 vdd.n312 vdd.n300 4.26717
R5592 vdd.n253 vdd.n241 4.26717
R5593 vdd.n210 vdd.n198 4.26717
R5594 vdd.n151 vdd.n139 4.26717
R5595 vdd.n109 vdd.n97 4.26717
R5596 vdd.n50 vdd.n38 4.26717
R5597 vdd.n1731 vdd.n1719 4.26717
R5598 vdd.n1790 vdd.n1778 4.26717
R5599 vdd.n1629 vdd.n1617 4.26717
R5600 vdd.n1688 vdd.n1676 4.26717
R5601 vdd.n1528 vdd.n1516 4.26717
R5602 vdd.n1587 vdd.n1575 4.26717
R5603 vdd.n1875 vdd.t141 4.19501
R5604 vdd.n3248 vdd.t137 4.19501
R5605 vdd.n333 vdd.n231 4.10845
R5606 vdd.n1811 vdd.n1709 4.10845
R5607 vdd.n289 vdd.t173 4.06363
R5608 vdd.n289 vdd.t235 4.06363
R5609 vdd.n287 vdd.t266 4.06363
R5610 vdd.n287 vdd.t282 4.06363
R5611 vdd.n285 vdd.t286 4.06363
R5612 vdd.n285 vdd.t180 4.06363
R5613 vdd.n283 vdd.t204 4.06363
R5614 vdd.n283 vdd.t285 4.06363
R5615 vdd.n281 vdd.t287 4.06363
R5616 vdd.n281 vdd.t203 4.06363
R5617 vdd.n279 vdd.t208 4.06363
R5618 vdd.n279 vdd.t210 4.06363
R5619 vdd.n277 vdd.t262 4.06363
R5620 vdd.n277 vdd.t162 4.06363
R5621 vdd.n275 vdd.t169 4.06363
R5622 vdd.n275 vdd.t233 4.06363
R5623 vdd.n273 vdd.t238 4.06363
R5624 vdd.n273 vdd.t268 4.06363
R5625 vdd.n187 vdd.t157 4.06363
R5626 vdd.n187 vdd.t212 4.06363
R5627 vdd.n185 vdd.t254 4.06363
R5628 vdd.n185 vdd.t271 4.06363
R5629 vdd.n183 vdd.t274 4.06363
R5630 vdd.n183 vdd.t136 4.06363
R5631 vdd.n181 vdd.t187 4.06363
R5632 vdd.n181 vdd.t273 4.06363
R5633 vdd.n179 vdd.t277 4.06363
R5634 vdd.n179 vdd.t186 4.06363
R5635 vdd.n177 vdd.t191 4.06363
R5636 vdd.n177 vdd.t193 4.06363
R5637 vdd.n175 vdd.t253 4.06363
R5638 vdd.n175 vdd.t132 4.06363
R5639 vdd.n173 vdd.t148 4.06363
R5640 vdd.n173 vdd.t213 4.06363
R5641 vdd.n171 vdd.t223 4.06363
R5642 vdd.n171 vdd.t255 4.06363
R5643 vdd.n86 vdd.t172 4.06363
R5644 vdd.n86 vdd.t260 4.06363
R5645 vdd.n84 vdd.t164 4.06363
R5646 vdd.n84 vdd.t245 4.06363
R5647 vdd.n82 vdd.t189 4.06363
R5648 vdd.n82 vdd.t229 4.06363
R5649 vdd.n80 vdd.t159 4.06363
R5650 vdd.n80 vdd.t219 4.06363
R5651 vdd.n78 vdd.t152 4.06363
R5652 vdd.n78 vdd.t194 4.06363
R5653 vdd.n76 vdd.t283 4.06363
R5654 vdd.n76 vdd.t259 4.06363
R5655 vdd.n74 vdd.t265 4.06363
R5656 vdd.n74 vdd.t205 4.06363
R5657 vdd.n72 vdd.t288 4.06363
R5658 vdd.n72 vdd.t182 4.06363
R5659 vdd.n70 vdd.t275 4.06363
R5660 vdd.n70 vdd.t215 4.06363
R5661 vdd.n1751 vdd.t171 4.06363
R5662 vdd.n1751 vdd.t281 4.06363
R5663 vdd.n1753 vdd.t278 4.06363
R5664 vdd.n1753 vdd.t261 4.06363
R5665 vdd.n1755 vdd.t228 4.06363
R5666 vdd.n1755 vdd.t168 4.06363
R5667 vdd.n1757 vdd.t290 4.06363
R5668 vdd.n1757 vdd.t258 4.06363
R5669 vdd.n1759 vdd.t239 4.06363
R5670 vdd.n1759 vdd.t202 4.06363
R5671 vdd.n1761 vdd.t198 4.06363
R5672 vdd.n1761 vdd.t256 4.06363
R5673 vdd.n1763 vdd.t241 4.06363
R5674 vdd.n1763 vdd.t240 4.06363
R5675 vdd.n1765 vdd.t195 4.06363
R5676 vdd.n1765 vdd.t170 4.06363
R5677 vdd.n1767 vdd.t166 4.06363
R5678 vdd.n1767 vdd.t236 4.06363
R5679 vdd.n1649 vdd.t134 4.06363
R5680 vdd.n1649 vdd.t270 4.06363
R5681 vdd.n1651 vdd.t264 4.06363
R5682 vdd.n1651 vdd.t250 4.06363
R5683 vdd.n1653 vdd.t209 4.06363
R5684 vdd.n1653 vdd.t144 4.06363
R5685 vdd.n1655 vdd.t279 4.06363
R5686 vdd.n1655 vdd.t248 4.06363
R5687 vdd.n1657 vdd.t242 4.06363
R5688 vdd.n1657 vdd.t150 4.06363
R5689 vdd.n1659 vdd.t179 4.06363
R5690 vdd.n1659 vdd.t243 4.06363
R5691 vdd.n1661 vdd.t227 4.06363
R5692 vdd.n1661 vdd.t225 4.06363
R5693 vdd.n1663 vdd.t175 4.06363
R5694 vdd.n1663 vdd.t154 4.06363
R5695 vdd.n1665 vdd.t140 4.06363
R5696 vdd.n1665 vdd.t221 4.06363
R5697 vdd.n1548 vdd.t217 4.06363
R5698 vdd.n1548 vdd.t276 4.06363
R5699 vdd.n1550 vdd.t184 4.06363
R5700 vdd.n1550 vdd.t257 4.06363
R5701 vdd.n1552 vdd.t207 4.06363
R5702 vdd.n1552 vdd.t234 4.06363
R5703 vdd.n1554 vdd.t231 4.06363
R5704 vdd.n1554 vdd.t284 4.06363
R5705 vdd.n1556 vdd.t197 4.06363
R5706 vdd.n1556 vdd.t155 4.06363
R5707 vdd.n1558 vdd.t220 4.06363
R5708 vdd.n1558 vdd.t161 4.06363
R5709 vdd.n1560 vdd.t272 4.06363
R5710 vdd.n1560 vdd.t289 4.06363
R5711 vdd.n1562 vdd.t246 4.06363
R5712 vdd.n1562 vdd.t165 4.06363
R5713 vdd.n1564 vdd.t232 4.06363
R5714 vdd.n1564 vdd.t177 4.06363
R5715 vdd.n26 vdd.t102 3.9605
R5716 vdd.n26 vdd.t291 3.9605
R5717 vdd.n23 vdd.t9 3.9605
R5718 vdd.n23 vdd.t107 3.9605
R5719 vdd.n21 vdd.t105 3.9605
R5720 vdd.n21 vdd.t108 3.9605
R5721 vdd.n20 vdd.t293 3.9605
R5722 vdd.n20 vdd.t8 3.9605
R5723 vdd.n15 vdd.t104 3.9605
R5724 vdd.n15 vdd.t7 3.9605
R5725 vdd.n16 vdd.t292 3.9605
R5726 vdd.n16 vdd.t100 3.9605
R5727 vdd.n18 vdd.t106 3.9605
R5728 vdd.n18 vdd.t117 3.9605
R5729 vdd.n25 vdd.t101 3.9605
R5730 vdd.n25 vdd.t118 3.9605
R5731 vdd.n7 vdd.t123 3.61217
R5732 vdd.n7 vdd.t114 3.61217
R5733 vdd.n8 vdd.t90 3.61217
R5734 vdd.n8 vdd.t2 3.61217
R5735 vdd.n10 vdd.t120 3.61217
R5736 vdd.n10 vdd.t98 3.61217
R5737 vdd.n12 vdd.t116 3.61217
R5738 vdd.n12 vdd.t6 3.61217
R5739 vdd.n5 vdd.t95 3.61217
R5740 vdd.n5 vdd.t88 3.61217
R5741 vdd.n3 vdd.t128 3.61217
R5742 vdd.n3 vdd.t110 3.61217
R5743 vdd.n1 vdd.t126 3.61217
R5744 vdd.n1 vdd.t4 3.61217
R5745 vdd.n0 vdd.t295 3.61217
R5746 vdd.n0 vdd.t93 3.61217
R5747 vdd.n316 vdd.n315 3.49141
R5748 vdd.n257 vdd.n256 3.49141
R5749 vdd.n214 vdd.n213 3.49141
R5750 vdd.n155 vdd.n154 3.49141
R5751 vdd.n113 vdd.n112 3.49141
R5752 vdd.n54 vdd.n53 3.49141
R5753 vdd.n1735 vdd.n1734 3.49141
R5754 vdd.n1794 vdd.n1793 3.49141
R5755 vdd.n1633 vdd.n1632 3.49141
R5756 vdd.n1692 vdd.n1691 3.49141
R5757 vdd.n1532 vdd.n1531 3.49141
R5758 vdd.n1591 vdd.n1590 3.49141
R5759 vdd.n2156 vdd.t127 3.40145
R5760 vdd.n2604 vdd.t94 3.40145
R5761 vdd.n2857 vdd.t5 3.40145
R5762 vdd.n2781 vdd.t97 3.40145
R5763 vdd.n1876 vdd.t269 3.28809
R5764 vdd.n3247 vdd.t222 3.28809
R5765 vdd.n2257 vdd.t294 3.17472
R5766 vdd.n2760 vdd.t113 3.17472
R5767 vdd.t183 vdd.n1104 3.06136
R5768 vdd.n3272 vdd.t181 3.06136
R5769 vdd.n1834 vdd.t247 2.83463
R5770 vdd.n644 vdd.t190 2.83463
R5771 vdd.n319 vdd.n298 2.71565
R5772 vdd.n260 vdd.n239 2.71565
R5773 vdd.n217 vdd.n196 2.71565
R5774 vdd.n158 vdd.n137 2.71565
R5775 vdd.n116 vdd.n95 2.71565
R5776 vdd.n57 vdd.n36 2.71565
R5777 vdd.n1738 vdd.n1717 2.71565
R5778 vdd.n1797 vdd.n1776 2.71565
R5779 vdd.n1636 vdd.n1615 2.71565
R5780 vdd.n1695 vdd.n1674 2.71565
R5781 vdd.n1535 vdd.n1514 2.71565
R5782 vdd.n1594 vdd.n1573 2.71565
R5783 vdd.t196 vdd.n1132 2.6079
R5784 vdd.n2406 vdd.t103 2.6079
R5785 vdd.n2430 vdd.t91 2.6079
R5786 vdd.n2894 vdd.t10 2.6079
R5787 vdd.n2918 vdd.t121 2.6079
R5788 vdd.n3395 vdd.t185 2.6079
R5789 vdd.n2924 vdd.n2923 2.49806
R5790 vdd.n2398 vdd.n2397 2.49806
R5791 vdd.n306 vdd.n305 2.4129
R5792 vdd.n247 vdd.n246 2.4129
R5793 vdd.n204 vdd.n203 2.4129
R5794 vdd.n145 vdd.n144 2.4129
R5795 vdd.n103 vdd.n102 2.4129
R5796 vdd.n44 vdd.n43 2.4129
R5797 vdd.n1725 vdd.n1724 2.4129
R5798 vdd.n1784 vdd.n1783 2.4129
R5799 vdd.n1623 vdd.n1622 2.4129
R5800 vdd.n1682 vdd.n1681 2.4129
R5801 vdd.n1522 vdd.n1521 2.4129
R5802 vdd.n1581 vdd.n1580 2.4129
R5803 vdd.n1486 vdd.t224 2.38117
R5804 vdd.n1894 vdd.t23 2.38117
R5805 vdd.n3231 vdd.t16 2.38117
R5806 vdd.n3386 vdd.t188 2.38117
R5807 vdd.n2315 vdd.n1904 2.27742
R5808 vdd.n2316 vdd.n2315 2.27742
R5809 vdd.n3216 vdd.n3215 2.27742
R5810 vdd.n3217 vdd.n3216 2.27742
R5811 vdd.n3094 vdd.n3093 2.27742
R5812 vdd.n3093 vdd.n784 2.27742
R5813 vdd.n2338 vdd.n1065 2.27742
R5814 vdd.n2338 vdd.n1066 2.27742
R5815 vdd.n2430 vdd.t125 2.2678
R5816 vdd.n2894 vdd.t1 2.2678
R5817 vdd.t174 vdd.n1161 2.15444
R5818 vdd.n3377 vdd.t244 2.15444
R5819 vdd.t3 vdd.n983 2.04107
R5820 vdd.n900 vdd.t89 2.04107
R5821 vdd.n320 vdd.n296 1.93989
R5822 vdd.n261 vdd.n237 1.93989
R5823 vdd.n218 vdd.n194 1.93989
R5824 vdd.n159 vdd.n135 1.93989
R5825 vdd.n117 vdd.n93 1.93989
R5826 vdd.n58 vdd.n34 1.93989
R5827 vdd.n1739 vdd.n1715 1.93989
R5828 vdd.n1798 vdd.n1774 1.93989
R5829 vdd.n1637 vdd.n1613 1.93989
R5830 vdd.n1696 vdd.n1672 1.93989
R5831 vdd.n1536 vdd.n1512 1.93989
R5832 vdd.n1595 vdd.n1571 1.93989
R5833 vdd.n1444 vdd.t145 1.92771
R5834 vdd.n2381 vdd.t12 1.92771
R5835 vdd.n2457 vdd.t51 1.92771
R5836 vdd.n2870 vdd.t59 1.92771
R5837 vdd.n2989 vdd.t55 1.92771
R5838 vdd.t199 vdd.n375 1.92771
R5839 vdd.n1452 vdd.t176 1.70098
R5840 vdd.n2257 vdd.t129 1.70098
R5841 vdd.n1008 vdd.t0 1.70098
R5842 vdd.t130 vdd.n874 1.70098
R5843 vdd.n2760 vdd.t99 1.70098
R5844 vdd.n3371 vdd.t156 1.70098
R5845 vdd.n1477 vdd.t226 1.47425
R5846 vdd.n361 vdd.t135 1.47425
R5847 vdd.n1143 vdd.t160 1.24752
R5848 vdd.t158 vdd.n3393 1.24752
R5849 vdd.n331 vdd.n291 1.16414
R5850 vdd.n324 vdd.n323 1.16414
R5851 vdd.n272 vdd.n232 1.16414
R5852 vdd.n265 vdd.n264 1.16414
R5853 vdd.n229 vdd.n189 1.16414
R5854 vdd.n222 vdd.n221 1.16414
R5855 vdd.n170 vdd.n130 1.16414
R5856 vdd.n163 vdd.n162 1.16414
R5857 vdd.n128 vdd.n88 1.16414
R5858 vdd.n121 vdd.n120 1.16414
R5859 vdd.n69 vdd.n29 1.16414
R5860 vdd.n62 vdd.n61 1.16414
R5861 vdd.n1750 vdd.n1710 1.16414
R5862 vdd.n1743 vdd.n1742 1.16414
R5863 vdd.n1809 vdd.n1769 1.16414
R5864 vdd.n1802 vdd.n1801 1.16414
R5865 vdd.n1648 vdd.n1608 1.16414
R5866 vdd.n1641 vdd.n1640 1.16414
R5867 vdd.n1707 vdd.n1667 1.16414
R5868 vdd.n1700 vdd.n1699 1.16414
R5869 vdd.n1547 vdd.n1507 1.16414
R5870 vdd.n1540 vdd.n1539 1.16414
R5871 vdd.n1606 vdd.n1566 1.16414
R5872 vdd.n1599 vdd.n1598 1.16414
R5873 vdd.n2424 vdd.t92 1.13415
R5874 vdd.n2900 vdd.t122 1.13415
R5875 vdd.n1826 vdd.t230 1.02079
R5876 vdd.t69 vdd.t111 1.02079
R5877 vdd.t96 vdd.t27 1.02079
R5878 vdd.t192 vdd.n633 1.02079
R5879 vdd.n1323 vdd.n1319 0.970197
R5880 vdd.n2336 vdd.n2335 0.970197
R5881 vdd.n618 vdd.n428 0.970197
R5882 vdd.n3095 vdd.n690 0.970197
R5883 vdd.n1812 vdd.n28 0.90431
R5884 vdd vdd.n3400 0.896477
R5885 vdd.n1842 vdd.t143 0.794056
R5886 vdd.n2400 vdd.t111 0.794056
R5887 vdd.n2436 vdd.t112 0.794056
R5888 vdd.n2888 vdd.t124 0.794056
R5889 vdd.n2926 vdd.t96 0.794056
R5890 vdd.n3281 vdd.t252 0.794056
R5891 vdd.n1867 vdd.t133 0.567326
R5892 vdd.t214 vdd.n662 0.567326
R5893 vdd.n2326 vdd.n2325 0.530988
R5894 vdd.n726 vdd.n682 0.530988
R5895 vdd.n464 vdd.n391 0.530988
R5896 vdd.n3350 vdd.n3349 0.530988
R5897 vdd.n3227 vdd.n3226 0.530988
R5898 vdd.n1889 vdd.n1067 0.530988
R5899 vdd.n1321 vdd.n1186 0.530988
R5900 vdd.n1423 vdd.n1422 0.530988
R5901 vdd.n4 vdd.n2 0.459552
R5902 vdd.n11 vdd.n9 0.459552
R5903 vdd.n329 vdd.n328 0.388379
R5904 vdd.n295 vdd.n293 0.388379
R5905 vdd.n270 vdd.n269 0.388379
R5906 vdd.n236 vdd.n234 0.388379
R5907 vdd.n227 vdd.n226 0.388379
R5908 vdd.n193 vdd.n191 0.388379
R5909 vdd.n168 vdd.n167 0.388379
R5910 vdd.n134 vdd.n132 0.388379
R5911 vdd.n126 vdd.n125 0.388379
R5912 vdd.n92 vdd.n90 0.388379
R5913 vdd.n67 vdd.n66 0.388379
R5914 vdd.n33 vdd.n31 0.388379
R5915 vdd.n1748 vdd.n1747 0.388379
R5916 vdd.n1714 vdd.n1712 0.388379
R5917 vdd.n1807 vdd.n1806 0.388379
R5918 vdd.n1773 vdd.n1771 0.388379
R5919 vdd.n1646 vdd.n1645 0.388379
R5920 vdd.n1612 vdd.n1610 0.388379
R5921 vdd.n1705 vdd.n1704 0.388379
R5922 vdd.n1671 vdd.n1669 0.388379
R5923 vdd.n1545 vdd.n1544 0.388379
R5924 vdd.n1511 vdd.n1509 0.388379
R5925 vdd.n1604 vdd.n1603 0.388379
R5926 vdd.n1570 vdd.n1568 0.388379
R5927 vdd.n19 vdd.n17 0.387128
R5928 vdd.n24 vdd.n22 0.387128
R5929 vdd.n6 vdd.n4 0.358259
R5930 vdd.n13 vdd.n11 0.358259
R5931 vdd.n276 vdd.n274 0.358259
R5932 vdd.n278 vdd.n276 0.358259
R5933 vdd.n280 vdd.n278 0.358259
R5934 vdd.n282 vdd.n280 0.358259
R5935 vdd.n284 vdd.n282 0.358259
R5936 vdd.n286 vdd.n284 0.358259
R5937 vdd.n288 vdd.n286 0.358259
R5938 vdd.n290 vdd.n288 0.358259
R5939 vdd.n332 vdd.n290 0.358259
R5940 vdd.n174 vdd.n172 0.358259
R5941 vdd.n176 vdd.n174 0.358259
R5942 vdd.n178 vdd.n176 0.358259
R5943 vdd.n180 vdd.n178 0.358259
R5944 vdd.n182 vdd.n180 0.358259
R5945 vdd.n184 vdd.n182 0.358259
R5946 vdd.n186 vdd.n184 0.358259
R5947 vdd.n188 vdd.n186 0.358259
R5948 vdd.n230 vdd.n188 0.358259
R5949 vdd.n73 vdd.n71 0.358259
R5950 vdd.n75 vdd.n73 0.358259
R5951 vdd.n77 vdd.n75 0.358259
R5952 vdd.n79 vdd.n77 0.358259
R5953 vdd.n81 vdd.n79 0.358259
R5954 vdd.n83 vdd.n81 0.358259
R5955 vdd.n85 vdd.n83 0.358259
R5956 vdd.n87 vdd.n85 0.358259
R5957 vdd.n129 vdd.n87 0.358259
R5958 vdd.n1810 vdd.n1768 0.358259
R5959 vdd.n1768 vdd.n1766 0.358259
R5960 vdd.n1766 vdd.n1764 0.358259
R5961 vdd.n1764 vdd.n1762 0.358259
R5962 vdd.n1762 vdd.n1760 0.358259
R5963 vdd.n1760 vdd.n1758 0.358259
R5964 vdd.n1758 vdd.n1756 0.358259
R5965 vdd.n1756 vdd.n1754 0.358259
R5966 vdd.n1754 vdd.n1752 0.358259
R5967 vdd.n1708 vdd.n1666 0.358259
R5968 vdd.n1666 vdd.n1664 0.358259
R5969 vdd.n1664 vdd.n1662 0.358259
R5970 vdd.n1662 vdd.n1660 0.358259
R5971 vdd.n1660 vdd.n1658 0.358259
R5972 vdd.n1658 vdd.n1656 0.358259
R5973 vdd.n1656 vdd.n1654 0.358259
R5974 vdd.n1654 vdd.n1652 0.358259
R5975 vdd.n1652 vdd.n1650 0.358259
R5976 vdd.n1607 vdd.n1565 0.358259
R5977 vdd.n1565 vdd.n1563 0.358259
R5978 vdd.n1563 vdd.n1561 0.358259
R5979 vdd.n1561 vdd.n1559 0.358259
R5980 vdd.n1559 vdd.n1557 0.358259
R5981 vdd.n1557 vdd.n1555 0.358259
R5982 vdd.n1555 vdd.n1553 0.358259
R5983 vdd.n1553 vdd.n1551 0.358259
R5984 vdd.n1551 vdd.n1549 0.358259
R5985 vdd.n14 vdd.n6 0.334552
R5986 vdd.n14 vdd.n13 0.334552
R5987 vdd.n27 vdd.n19 0.21707
R5988 vdd.n27 vdd.n24 0.21707
R5989 vdd.n330 vdd.n292 0.155672
R5990 vdd.n322 vdd.n292 0.155672
R5991 vdd.n322 vdd.n321 0.155672
R5992 vdd.n321 vdd.n297 0.155672
R5993 vdd.n314 vdd.n297 0.155672
R5994 vdd.n314 vdd.n313 0.155672
R5995 vdd.n313 vdd.n301 0.155672
R5996 vdd.n306 vdd.n301 0.155672
R5997 vdd.n271 vdd.n233 0.155672
R5998 vdd.n263 vdd.n233 0.155672
R5999 vdd.n263 vdd.n262 0.155672
R6000 vdd.n262 vdd.n238 0.155672
R6001 vdd.n255 vdd.n238 0.155672
R6002 vdd.n255 vdd.n254 0.155672
R6003 vdd.n254 vdd.n242 0.155672
R6004 vdd.n247 vdd.n242 0.155672
R6005 vdd.n228 vdd.n190 0.155672
R6006 vdd.n220 vdd.n190 0.155672
R6007 vdd.n220 vdd.n219 0.155672
R6008 vdd.n219 vdd.n195 0.155672
R6009 vdd.n212 vdd.n195 0.155672
R6010 vdd.n212 vdd.n211 0.155672
R6011 vdd.n211 vdd.n199 0.155672
R6012 vdd.n204 vdd.n199 0.155672
R6013 vdd.n169 vdd.n131 0.155672
R6014 vdd.n161 vdd.n131 0.155672
R6015 vdd.n161 vdd.n160 0.155672
R6016 vdd.n160 vdd.n136 0.155672
R6017 vdd.n153 vdd.n136 0.155672
R6018 vdd.n153 vdd.n152 0.155672
R6019 vdd.n152 vdd.n140 0.155672
R6020 vdd.n145 vdd.n140 0.155672
R6021 vdd.n127 vdd.n89 0.155672
R6022 vdd.n119 vdd.n89 0.155672
R6023 vdd.n119 vdd.n118 0.155672
R6024 vdd.n118 vdd.n94 0.155672
R6025 vdd.n111 vdd.n94 0.155672
R6026 vdd.n111 vdd.n110 0.155672
R6027 vdd.n110 vdd.n98 0.155672
R6028 vdd.n103 vdd.n98 0.155672
R6029 vdd.n68 vdd.n30 0.155672
R6030 vdd.n60 vdd.n30 0.155672
R6031 vdd.n60 vdd.n59 0.155672
R6032 vdd.n59 vdd.n35 0.155672
R6033 vdd.n52 vdd.n35 0.155672
R6034 vdd.n52 vdd.n51 0.155672
R6035 vdd.n51 vdd.n39 0.155672
R6036 vdd.n44 vdd.n39 0.155672
R6037 vdd.n1749 vdd.n1711 0.155672
R6038 vdd.n1741 vdd.n1711 0.155672
R6039 vdd.n1741 vdd.n1740 0.155672
R6040 vdd.n1740 vdd.n1716 0.155672
R6041 vdd.n1733 vdd.n1716 0.155672
R6042 vdd.n1733 vdd.n1732 0.155672
R6043 vdd.n1732 vdd.n1720 0.155672
R6044 vdd.n1725 vdd.n1720 0.155672
R6045 vdd.n1808 vdd.n1770 0.155672
R6046 vdd.n1800 vdd.n1770 0.155672
R6047 vdd.n1800 vdd.n1799 0.155672
R6048 vdd.n1799 vdd.n1775 0.155672
R6049 vdd.n1792 vdd.n1775 0.155672
R6050 vdd.n1792 vdd.n1791 0.155672
R6051 vdd.n1791 vdd.n1779 0.155672
R6052 vdd.n1784 vdd.n1779 0.155672
R6053 vdd.n1647 vdd.n1609 0.155672
R6054 vdd.n1639 vdd.n1609 0.155672
R6055 vdd.n1639 vdd.n1638 0.155672
R6056 vdd.n1638 vdd.n1614 0.155672
R6057 vdd.n1631 vdd.n1614 0.155672
R6058 vdd.n1631 vdd.n1630 0.155672
R6059 vdd.n1630 vdd.n1618 0.155672
R6060 vdd.n1623 vdd.n1618 0.155672
R6061 vdd.n1706 vdd.n1668 0.155672
R6062 vdd.n1698 vdd.n1668 0.155672
R6063 vdd.n1698 vdd.n1697 0.155672
R6064 vdd.n1697 vdd.n1673 0.155672
R6065 vdd.n1690 vdd.n1673 0.155672
R6066 vdd.n1690 vdd.n1689 0.155672
R6067 vdd.n1689 vdd.n1677 0.155672
R6068 vdd.n1682 vdd.n1677 0.155672
R6069 vdd.n1546 vdd.n1508 0.155672
R6070 vdd.n1538 vdd.n1508 0.155672
R6071 vdd.n1538 vdd.n1537 0.155672
R6072 vdd.n1537 vdd.n1513 0.155672
R6073 vdd.n1530 vdd.n1513 0.155672
R6074 vdd.n1530 vdd.n1529 0.155672
R6075 vdd.n1529 vdd.n1517 0.155672
R6076 vdd.n1522 vdd.n1517 0.155672
R6077 vdd.n1605 vdd.n1567 0.155672
R6078 vdd.n1597 vdd.n1567 0.155672
R6079 vdd.n1597 vdd.n1596 0.155672
R6080 vdd.n1596 vdd.n1572 0.155672
R6081 vdd.n1589 vdd.n1572 0.155672
R6082 vdd.n1589 vdd.n1588 0.155672
R6083 vdd.n1588 vdd.n1576 0.155672
R6084 vdd.n1581 vdd.n1576 0.155672
R6085 vdd.n2101 vdd.n1906 0.152939
R6086 vdd.n1912 vdd.n1906 0.152939
R6087 vdd.n1913 vdd.n1912 0.152939
R6088 vdd.n1914 vdd.n1913 0.152939
R6089 vdd.n1915 vdd.n1914 0.152939
R6090 vdd.n1919 vdd.n1915 0.152939
R6091 vdd.n1920 vdd.n1919 0.152939
R6092 vdd.n1921 vdd.n1920 0.152939
R6093 vdd.n1922 vdd.n1921 0.152939
R6094 vdd.n1926 vdd.n1922 0.152939
R6095 vdd.n1927 vdd.n1926 0.152939
R6096 vdd.n1928 vdd.n1927 0.152939
R6097 vdd.n2076 vdd.n1928 0.152939
R6098 vdd.n2076 vdd.n2075 0.152939
R6099 vdd.n2075 vdd.n2074 0.152939
R6100 vdd.n2074 vdd.n1934 0.152939
R6101 vdd.n1939 vdd.n1934 0.152939
R6102 vdd.n1940 vdd.n1939 0.152939
R6103 vdd.n1941 vdd.n1940 0.152939
R6104 vdd.n1945 vdd.n1941 0.152939
R6105 vdd.n1946 vdd.n1945 0.152939
R6106 vdd.n1947 vdd.n1946 0.152939
R6107 vdd.n1948 vdd.n1947 0.152939
R6108 vdd.n1952 vdd.n1948 0.152939
R6109 vdd.n1953 vdd.n1952 0.152939
R6110 vdd.n1954 vdd.n1953 0.152939
R6111 vdd.n1955 vdd.n1954 0.152939
R6112 vdd.n1959 vdd.n1955 0.152939
R6113 vdd.n1960 vdd.n1959 0.152939
R6114 vdd.n1961 vdd.n1960 0.152939
R6115 vdd.n1962 vdd.n1961 0.152939
R6116 vdd.n1966 vdd.n1962 0.152939
R6117 vdd.n1967 vdd.n1966 0.152939
R6118 vdd.n1968 vdd.n1967 0.152939
R6119 vdd.n2037 vdd.n1968 0.152939
R6120 vdd.n2037 vdd.n2036 0.152939
R6121 vdd.n2036 vdd.n2035 0.152939
R6122 vdd.n2035 vdd.n1974 0.152939
R6123 vdd.n1979 vdd.n1974 0.152939
R6124 vdd.n1980 vdd.n1979 0.152939
R6125 vdd.n1981 vdd.n1980 0.152939
R6126 vdd.n1985 vdd.n1981 0.152939
R6127 vdd.n1986 vdd.n1985 0.152939
R6128 vdd.n1987 vdd.n1986 0.152939
R6129 vdd.n1988 vdd.n1987 0.152939
R6130 vdd.n1992 vdd.n1988 0.152939
R6131 vdd.n1993 vdd.n1992 0.152939
R6132 vdd.n1994 vdd.n1993 0.152939
R6133 vdd.n1995 vdd.n1994 0.152939
R6134 vdd.n1996 vdd.n1995 0.152939
R6135 vdd.n1996 vdd.n1064 0.152939
R6136 vdd.n2325 vdd.n1900 0.152939
R6137 vdd.n1814 vdd.n1123 0.152939
R6138 vdd.n1829 vdd.n1123 0.152939
R6139 vdd.n1830 vdd.n1829 0.152939
R6140 vdd.n1831 vdd.n1830 0.152939
R6141 vdd.n1831 vdd.n1112 0.152939
R6142 vdd.n1846 vdd.n1112 0.152939
R6143 vdd.n1847 vdd.n1846 0.152939
R6144 vdd.n1848 vdd.n1847 0.152939
R6145 vdd.n1848 vdd.n1101 0.152939
R6146 vdd.n1862 vdd.n1101 0.152939
R6147 vdd.n1863 vdd.n1862 0.152939
R6148 vdd.n1864 vdd.n1863 0.152939
R6149 vdd.n1864 vdd.n1089 0.152939
R6150 vdd.n1879 vdd.n1089 0.152939
R6151 vdd.n1880 vdd.n1879 0.152939
R6152 vdd.n1881 vdd.n1880 0.152939
R6153 vdd.n1881 vdd.n1077 0.152939
R6154 vdd.n1898 vdd.n1077 0.152939
R6155 vdd.n1899 vdd.n1898 0.152939
R6156 vdd.n2326 vdd.n1899 0.152939
R6157 vdd.n735 vdd.n730 0.152939
R6158 vdd.n736 vdd.n735 0.152939
R6159 vdd.n737 vdd.n736 0.152939
R6160 vdd.n738 vdd.n737 0.152939
R6161 vdd.n739 vdd.n738 0.152939
R6162 vdd.n740 vdd.n739 0.152939
R6163 vdd.n741 vdd.n740 0.152939
R6164 vdd.n742 vdd.n741 0.152939
R6165 vdd.n743 vdd.n742 0.152939
R6166 vdd.n744 vdd.n743 0.152939
R6167 vdd.n745 vdd.n744 0.152939
R6168 vdd.n746 vdd.n745 0.152939
R6169 vdd.n3183 vdd.n746 0.152939
R6170 vdd.n3183 vdd.n3182 0.152939
R6171 vdd.n3182 vdd.n3181 0.152939
R6172 vdd.n3181 vdd.n748 0.152939
R6173 vdd.n749 vdd.n748 0.152939
R6174 vdd.n750 vdd.n749 0.152939
R6175 vdd.n751 vdd.n750 0.152939
R6176 vdd.n752 vdd.n751 0.152939
R6177 vdd.n753 vdd.n752 0.152939
R6178 vdd.n754 vdd.n753 0.152939
R6179 vdd.n755 vdd.n754 0.152939
R6180 vdd.n756 vdd.n755 0.152939
R6181 vdd.n757 vdd.n756 0.152939
R6182 vdd.n758 vdd.n757 0.152939
R6183 vdd.n759 vdd.n758 0.152939
R6184 vdd.n760 vdd.n759 0.152939
R6185 vdd.n761 vdd.n760 0.152939
R6186 vdd.n762 vdd.n761 0.152939
R6187 vdd.n763 vdd.n762 0.152939
R6188 vdd.n764 vdd.n763 0.152939
R6189 vdd.n765 vdd.n764 0.152939
R6190 vdd.n766 vdd.n765 0.152939
R6191 vdd.n3137 vdd.n766 0.152939
R6192 vdd.n3137 vdd.n3136 0.152939
R6193 vdd.n3136 vdd.n3135 0.152939
R6194 vdd.n3135 vdd.n770 0.152939
R6195 vdd.n771 vdd.n770 0.152939
R6196 vdd.n772 vdd.n771 0.152939
R6197 vdd.n773 vdd.n772 0.152939
R6198 vdd.n774 vdd.n773 0.152939
R6199 vdd.n775 vdd.n774 0.152939
R6200 vdd.n776 vdd.n775 0.152939
R6201 vdd.n777 vdd.n776 0.152939
R6202 vdd.n778 vdd.n777 0.152939
R6203 vdd.n779 vdd.n778 0.152939
R6204 vdd.n780 vdd.n779 0.152939
R6205 vdd.n781 vdd.n780 0.152939
R6206 vdd.n782 vdd.n781 0.152939
R6207 vdd.n783 vdd.n782 0.152939
R6208 vdd.n727 vdd.n726 0.152939
R6209 vdd.n3234 vdd.n682 0.152939
R6210 vdd.n3235 vdd.n3234 0.152939
R6211 vdd.n3236 vdd.n3235 0.152939
R6212 vdd.n3236 vdd.n670 0.152939
R6213 vdd.n3251 vdd.n670 0.152939
R6214 vdd.n3252 vdd.n3251 0.152939
R6215 vdd.n3253 vdd.n3252 0.152939
R6216 vdd.n3253 vdd.n659 0.152939
R6217 vdd.n3267 vdd.n659 0.152939
R6218 vdd.n3268 vdd.n3267 0.152939
R6219 vdd.n3269 vdd.n3268 0.152939
R6220 vdd.n3269 vdd.n647 0.152939
R6221 vdd.n3284 vdd.n647 0.152939
R6222 vdd.n3285 vdd.n3284 0.152939
R6223 vdd.n3286 vdd.n3285 0.152939
R6224 vdd.n3286 vdd.n636 0.152939
R6225 vdd.n3303 vdd.n636 0.152939
R6226 vdd.n3304 vdd.n3303 0.152939
R6227 vdd.n3305 vdd.n3304 0.152939
R6228 vdd.n3305 vdd.n334 0.152939
R6229 vdd.n3398 vdd.n335 0.152939
R6230 vdd.n346 vdd.n335 0.152939
R6231 vdd.n347 vdd.n346 0.152939
R6232 vdd.n348 vdd.n347 0.152939
R6233 vdd.n355 vdd.n348 0.152939
R6234 vdd.n356 vdd.n355 0.152939
R6235 vdd.n357 vdd.n356 0.152939
R6236 vdd.n358 vdd.n357 0.152939
R6237 vdd.n366 vdd.n358 0.152939
R6238 vdd.n367 vdd.n366 0.152939
R6239 vdd.n368 vdd.n367 0.152939
R6240 vdd.n369 vdd.n368 0.152939
R6241 vdd.n377 vdd.n369 0.152939
R6242 vdd.n378 vdd.n377 0.152939
R6243 vdd.n379 vdd.n378 0.152939
R6244 vdd.n380 vdd.n379 0.152939
R6245 vdd.n388 vdd.n380 0.152939
R6246 vdd.n389 vdd.n388 0.152939
R6247 vdd.n390 vdd.n389 0.152939
R6248 vdd.n391 vdd.n390 0.152939
R6249 vdd.n464 vdd.n463 0.152939
R6250 vdd.n470 vdd.n463 0.152939
R6251 vdd.n471 vdd.n470 0.152939
R6252 vdd.n472 vdd.n471 0.152939
R6253 vdd.n472 vdd.n461 0.152939
R6254 vdd.n480 vdd.n461 0.152939
R6255 vdd.n481 vdd.n480 0.152939
R6256 vdd.n482 vdd.n481 0.152939
R6257 vdd.n482 vdd.n459 0.152939
R6258 vdd.n490 vdd.n459 0.152939
R6259 vdd.n491 vdd.n490 0.152939
R6260 vdd.n492 vdd.n491 0.152939
R6261 vdd.n492 vdd.n457 0.152939
R6262 vdd.n500 vdd.n457 0.152939
R6263 vdd.n501 vdd.n500 0.152939
R6264 vdd.n502 vdd.n501 0.152939
R6265 vdd.n502 vdd.n455 0.152939
R6266 vdd.n510 vdd.n455 0.152939
R6267 vdd.n511 vdd.n510 0.152939
R6268 vdd.n512 vdd.n511 0.152939
R6269 vdd.n512 vdd.n451 0.152939
R6270 vdd.n520 vdd.n451 0.152939
R6271 vdd.n521 vdd.n520 0.152939
R6272 vdd.n522 vdd.n521 0.152939
R6273 vdd.n522 vdd.n449 0.152939
R6274 vdd.n530 vdd.n449 0.152939
R6275 vdd.n531 vdd.n530 0.152939
R6276 vdd.n532 vdd.n531 0.152939
R6277 vdd.n532 vdd.n447 0.152939
R6278 vdd.n540 vdd.n447 0.152939
R6279 vdd.n541 vdd.n540 0.152939
R6280 vdd.n542 vdd.n541 0.152939
R6281 vdd.n542 vdd.n445 0.152939
R6282 vdd.n550 vdd.n445 0.152939
R6283 vdd.n551 vdd.n550 0.152939
R6284 vdd.n552 vdd.n551 0.152939
R6285 vdd.n552 vdd.n443 0.152939
R6286 vdd.n560 vdd.n443 0.152939
R6287 vdd.n561 vdd.n560 0.152939
R6288 vdd.n562 vdd.n561 0.152939
R6289 vdd.n562 vdd.n439 0.152939
R6290 vdd.n570 vdd.n439 0.152939
R6291 vdd.n571 vdd.n570 0.152939
R6292 vdd.n572 vdd.n571 0.152939
R6293 vdd.n572 vdd.n437 0.152939
R6294 vdd.n580 vdd.n437 0.152939
R6295 vdd.n581 vdd.n580 0.152939
R6296 vdd.n582 vdd.n581 0.152939
R6297 vdd.n582 vdd.n435 0.152939
R6298 vdd.n590 vdd.n435 0.152939
R6299 vdd.n591 vdd.n590 0.152939
R6300 vdd.n592 vdd.n591 0.152939
R6301 vdd.n592 vdd.n433 0.152939
R6302 vdd.n600 vdd.n433 0.152939
R6303 vdd.n601 vdd.n600 0.152939
R6304 vdd.n602 vdd.n601 0.152939
R6305 vdd.n602 vdd.n431 0.152939
R6306 vdd.n610 vdd.n431 0.152939
R6307 vdd.n611 vdd.n610 0.152939
R6308 vdd.n612 vdd.n611 0.152939
R6309 vdd.n612 vdd.n429 0.152939
R6310 vdd.n619 vdd.n429 0.152939
R6311 vdd.n3350 vdd.n619 0.152939
R6312 vdd.n3228 vdd.n3227 0.152939
R6313 vdd.n3228 vdd.n675 0.152939
R6314 vdd.n3242 vdd.n675 0.152939
R6315 vdd.n3243 vdd.n3242 0.152939
R6316 vdd.n3244 vdd.n3243 0.152939
R6317 vdd.n3244 vdd.n665 0.152939
R6318 vdd.n3259 vdd.n665 0.152939
R6319 vdd.n3260 vdd.n3259 0.152939
R6320 vdd.n3261 vdd.n3260 0.152939
R6321 vdd.n3261 vdd.n652 0.152939
R6322 vdd.n3275 vdd.n652 0.152939
R6323 vdd.n3276 vdd.n3275 0.152939
R6324 vdd.n3277 vdd.n3276 0.152939
R6325 vdd.n3277 vdd.n641 0.152939
R6326 vdd.n3292 vdd.n641 0.152939
R6327 vdd.n3293 vdd.n3292 0.152939
R6328 vdd.n3294 vdd.n3293 0.152939
R6329 vdd.n3296 vdd.n3294 0.152939
R6330 vdd.n3296 vdd.n3295 0.152939
R6331 vdd.n3295 vdd.n630 0.152939
R6332 vdd.n3313 vdd.n630 0.152939
R6333 vdd.n3314 vdd.n3313 0.152939
R6334 vdd.n3315 vdd.n3314 0.152939
R6335 vdd.n3315 vdd.n628 0.152939
R6336 vdd.n3320 vdd.n628 0.152939
R6337 vdd.n3321 vdd.n3320 0.152939
R6338 vdd.n3322 vdd.n3321 0.152939
R6339 vdd.n3322 vdd.n626 0.152939
R6340 vdd.n3327 vdd.n626 0.152939
R6341 vdd.n3328 vdd.n3327 0.152939
R6342 vdd.n3329 vdd.n3328 0.152939
R6343 vdd.n3329 vdd.n624 0.152939
R6344 vdd.n3335 vdd.n624 0.152939
R6345 vdd.n3336 vdd.n3335 0.152939
R6346 vdd.n3337 vdd.n3336 0.152939
R6347 vdd.n3337 vdd.n622 0.152939
R6348 vdd.n3342 vdd.n622 0.152939
R6349 vdd.n3343 vdd.n3342 0.152939
R6350 vdd.n3344 vdd.n3343 0.152939
R6351 vdd.n3344 vdd.n620 0.152939
R6352 vdd.n3349 vdd.n620 0.152939
R6353 vdd.n3226 vdd.n687 0.152939
R6354 vdd.n2337 vdd.n1067 0.152939
R6355 vdd.n1430 vdd.n1186 0.152939
R6356 vdd.n1431 vdd.n1430 0.152939
R6357 vdd.n1432 vdd.n1431 0.152939
R6358 vdd.n1432 vdd.n1174 0.152939
R6359 vdd.n1447 vdd.n1174 0.152939
R6360 vdd.n1448 vdd.n1447 0.152939
R6361 vdd.n1449 vdd.n1448 0.152939
R6362 vdd.n1449 vdd.n1164 0.152939
R6363 vdd.n1464 vdd.n1164 0.152939
R6364 vdd.n1465 vdd.n1464 0.152939
R6365 vdd.n1466 vdd.n1465 0.152939
R6366 vdd.n1466 vdd.n1151 0.152939
R6367 vdd.n1480 vdd.n1151 0.152939
R6368 vdd.n1481 vdd.n1480 0.152939
R6369 vdd.n1482 vdd.n1481 0.152939
R6370 vdd.n1482 vdd.n1140 0.152939
R6371 vdd.n1497 vdd.n1140 0.152939
R6372 vdd.n1498 vdd.n1497 0.152939
R6373 vdd.n1499 vdd.n1498 0.152939
R6374 vdd.n1499 vdd.n1129 0.152939
R6375 vdd.n1820 vdd.n1129 0.152939
R6376 vdd.n1821 vdd.n1820 0.152939
R6377 vdd.n1822 vdd.n1821 0.152939
R6378 vdd.n1822 vdd.n1117 0.152939
R6379 vdd.n1837 vdd.n1117 0.152939
R6380 vdd.n1838 vdd.n1837 0.152939
R6381 vdd.n1839 vdd.n1838 0.152939
R6382 vdd.n1839 vdd.n1107 0.152939
R6383 vdd.n1854 vdd.n1107 0.152939
R6384 vdd.n1855 vdd.n1854 0.152939
R6385 vdd.n1856 vdd.n1855 0.152939
R6386 vdd.n1856 vdd.n1094 0.152939
R6387 vdd.n1870 vdd.n1094 0.152939
R6388 vdd.n1871 vdd.n1870 0.152939
R6389 vdd.n1872 vdd.n1871 0.152939
R6390 vdd.n1872 vdd.n1084 0.152939
R6391 vdd.n1887 vdd.n1084 0.152939
R6392 vdd.n1888 vdd.n1887 0.152939
R6393 vdd.n1891 vdd.n1888 0.152939
R6394 vdd.n1891 vdd.n1890 0.152939
R6395 vdd.n1890 vdd.n1889 0.152939
R6396 vdd.n1422 vdd.n1191 0.152939
R6397 vdd.n1415 vdd.n1191 0.152939
R6398 vdd.n1415 vdd.n1414 0.152939
R6399 vdd.n1414 vdd.n1413 0.152939
R6400 vdd.n1413 vdd.n1228 0.152939
R6401 vdd.n1409 vdd.n1228 0.152939
R6402 vdd.n1409 vdd.n1408 0.152939
R6403 vdd.n1408 vdd.n1407 0.152939
R6404 vdd.n1407 vdd.n1234 0.152939
R6405 vdd.n1403 vdd.n1234 0.152939
R6406 vdd.n1403 vdd.n1402 0.152939
R6407 vdd.n1402 vdd.n1401 0.152939
R6408 vdd.n1401 vdd.n1240 0.152939
R6409 vdd.n1397 vdd.n1240 0.152939
R6410 vdd.n1397 vdd.n1396 0.152939
R6411 vdd.n1396 vdd.n1395 0.152939
R6412 vdd.n1395 vdd.n1246 0.152939
R6413 vdd.n1391 vdd.n1246 0.152939
R6414 vdd.n1391 vdd.n1390 0.152939
R6415 vdd.n1390 vdd.n1389 0.152939
R6416 vdd.n1389 vdd.n1254 0.152939
R6417 vdd.n1385 vdd.n1254 0.152939
R6418 vdd.n1385 vdd.n1384 0.152939
R6419 vdd.n1384 vdd.n1383 0.152939
R6420 vdd.n1383 vdd.n1260 0.152939
R6421 vdd.n1379 vdd.n1260 0.152939
R6422 vdd.n1379 vdd.n1378 0.152939
R6423 vdd.n1378 vdd.n1377 0.152939
R6424 vdd.n1377 vdd.n1266 0.152939
R6425 vdd.n1373 vdd.n1266 0.152939
R6426 vdd.n1373 vdd.n1372 0.152939
R6427 vdd.n1372 vdd.n1371 0.152939
R6428 vdd.n1371 vdd.n1272 0.152939
R6429 vdd.n1367 vdd.n1272 0.152939
R6430 vdd.n1367 vdd.n1366 0.152939
R6431 vdd.n1366 vdd.n1365 0.152939
R6432 vdd.n1365 vdd.n1278 0.152939
R6433 vdd.n1361 vdd.n1278 0.152939
R6434 vdd.n1361 vdd.n1360 0.152939
R6435 vdd.n1360 vdd.n1359 0.152939
R6436 vdd.n1359 vdd.n1284 0.152939
R6437 vdd.n1352 vdd.n1284 0.152939
R6438 vdd.n1352 vdd.n1351 0.152939
R6439 vdd.n1351 vdd.n1350 0.152939
R6440 vdd.n1350 vdd.n1289 0.152939
R6441 vdd.n1346 vdd.n1289 0.152939
R6442 vdd.n1346 vdd.n1345 0.152939
R6443 vdd.n1345 vdd.n1344 0.152939
R6444 vdd.n1344 vdd.n1295 0.152939
R6445 vdd.n1340 vdd.n1295 0.152939
R6446 vdd.n1340 vdd.n1339 0.152939
R6447 vdd.n1339 vdd.n1338 0.152939
R6448 vdd.n1338 vdd.n1301 0.152939
R6449 vdd.n1334 vdd.n1301 0.152939
R6450 vdd.n1334 vdd.n1333 0.152939
R6451 vdd.n1333 vdd.n1332 0.152939
R6452 vdd.n1332 vdd.n1307 0.152939
R6453 vdd.n1328 vdd.n1307 0.152939
R6454 vdd.n1328 vdd.n1327 0.152939
R6455 vdd.n1327 vdd.n1326 0.152939
R6456 vdd.n1326 vdd.n1313 0.152939
R6457 vdd.n1322 vdd.n1313 0.152939
R6458 vdd.n1322 vdd.n1321 0.152939
R6459 vdd.n1424 vdd.n1423 0.152939
R6460 vdd.n1424 vdd.n1180 0.152939
R6461 vdd.n1439 vdd.n1180 0.152939
R6462 vdd.n1440 vdd.n1439 0.152939
R6463 vdd.n1441 vdd.n1440 0.152939
R6464 vdd.n1441 vdd.n1169 0.152939
R6465 vdd.n1456 vdd.n1169 0.152939
R6466 vdd.n1457 vdd.n1456 0.152939
R6467 vdd.n1458 vdd.n1457 0.152939
R6468 vdd.n1458 vdd.n1158 0.152939
R6469 vdd.n1472 vdd.n1158 0.152939
R6470 vdd.n1473 vdd.n1472 0.152939
R6471 vdd.n1474 vdd.n1473 0.152939
R6472 vdd.n1474 vdd.n1146 0.152939
R6473 vdd.n1489 vdd.n1146 0.152939
R6474 vdd.n1490 vdd.n1489 0.152939
R6475 vdd.n1491 vdd.n1490 0.152939
R6476 vdd.n1491 vdd.n1135 0.152939
R6477 vdd.n1505 vdd.n1135 0.152939
R6478 vdd.n1506 vdd.n1505 0.152939
R6479 vdd.n1427 vdd.t31 0.113865
R6480 vdd.t38 vdd.n386 0.113865
R6481 vdd.n2315 vdd.n1900 0.110256
R6482 vdd.n3216 vdd.n727 0.110256
R6483 vdd.n3093 vdd.n687 0.110256
R6484 vdd.n2338 vdd.n2337 0.110256
R6485 vdd.n1814 vdd.n1813 0.0695946
R6486 vdd.n3399 vdd.n334 0.0695946
R6487 vdd.n3399 vdd.n3398 0.0695946
R6488 vdd.n1813 vdd.n1506 0.0695946
R6489 vdd.n2315 vdd.n2101 0.0431829
R6490 vdd.n2338 vdd.n1064 0.0431829
R6491 vdd.n3216 vdd.n730 0.0431829
R6492 vdd.n3093 vdd.n783 0.0431829
R6493 vdd vdd.n28 0.00833333
R6494 CSoutput.n19 CSoutput.t230 184.661
R6495 CSoutput.n78 CSoutput.n77 165.8
R6496 CSoutput.n76 CSoutput.n0 165.8
R6497 CSoutput.n75 CSoutput.n74 165.8
R6498 CSoutput.n73 CSoutput.n72 165.8
R6499 CSoutput.n71 CSoutput.n2 165.8
R6500 CSoutput.n69 CSoutput.n68 165.8
R6501 CSoutput.n67 CSoutput.n3 165.8
R6502 CSoutput.n66 CSoutput.n65 165.8
R6503 CSoutput.n63 CSoutput.n4 165.8
R6504 CSoutput.n61 CSoutput.n60 165.8
R6505 CSoutput.n59 CSoutput.n5 165.8
R6506 CSoutput.n58 CSoutput.n57 165.8
R6507 CSoutput.n55 CSoutput.n6 165.8
R6508 CSoutput.n54 CSoutput.n53 165.8
R6509 CSoutput.n52 CSoutput.n51 165.8
R6510 CSoutput.n50 CSoutput.n8 165.8
R6511 CSoutput.n48 CSoutput.n47 165.8
R6512 CSoutput.n46 CSoutput.n9 165.8
R6513 CSoutput.n45 CSoutput.n44 165.8
R6514 CSoutput.n42 CSoutput.n10 165.8
R6515 CSoutput.n41 CSoutput.n40 165.8
R6516 CSoutput.n39 CSoutput.n38 165.8
R6517 CSoutput.n37 CSoutput.n12 165.8
R6518 CSoutput.n35 CSoutput.n34 165.8
R6519 CSoutput.n33 CSoutput.n13 165.8
R6520 CSoutput.n32 CSoutput.n31 165.8
R6521 CSoutput.n29 CSoutput.n14 165.8
R6522 CSoutput.n28 CSoutput.n27 165.8
R6523 CSoutput.n26 CSoutput.n25 165.8
R6524 CSoutput.n24 CSoutput.n16 165.8
R6525 CSoutput.n22 CSoutput.n21 165.8
R6526 CSoutput.n20 CSoutput.n17 165.8
R6527 CSoutput.n77 CSoutput.t231 162.194
R6528 CSoutput.n18 CSoutput.t232 120.501
R6529 CSoutput.n23 CSoutput.t220 120.501
R6530 CSoutput.n15 CSoutput.t218 120.501
R6531 CSoutput.n30 CSoutput.t234 120.501
R6532 CSoutput.n36 CSoutput.t222 120.501
R6533 CSoutput.n11 CSoutput.t224 120.501
R6534 CSoutput.n43 CSoutput.t237 120.501
R6535 CSoutput.n49 CSoutput.t225 120.501
R6536 CSoutput.n7 CSoutput.t227 120.501
R6537 CSoutput.n56 CSoutput.t221 120.501
R6538 CSoutput.n62 CSoutput.t235 120.501
R6539 CSoutput.n64 CSoutput.t229 120.501
R6540 CSoutput.n70 CSoutput.t223 120.501
R6541 CSoutput.n1 CSoutput.t219 120.501
R6542 CSoutput.n330 CSoutput.n328 103.469
R6543 CSoutput.n310 CSoutput.n308 103.469
R6544 CSoutput.n291 CSoutput.n289 103.469
R6545 CSoutput.n120 CSoutput.n118 103.469
R6546 CSoutput.n100 CSoutput.n98 103.469
R6547 CSoutput.n81 CSoutput.n79 103.469
R6548 CSoutput.n344 CSoutput.n343 103.111
R6549 CSoutput.n342 CSoutput.n341 103.111
R6550 CSoutput.n340 CSoutput.n339 103.111
R6551 CSoutput.n338 CSoutput.n337 103.111
R6552 CSoutput.n336 CSoutput.n335 103.111
R6553 CSoutput.n334 CSoutput.n333 103.111
R6554 CSoutput.n332 CSoutput.n331 103.111
R6555 CSoutput.n330 CSoutput.n329 103.111
R6556 CSoutput.n326 CSoutput.n325 103.111
R6557 CSoutput.n324 CSoutput.n323 103.111
R6558 CSoutput.n322 CSoutput.n321 103.111
R6559 CSoutput.n320 CSoutput.n319 103.111
R6560 CSoutput.n318 CSoutput.n317 103.111
R6561 CSoutput.n316 CSoutput.n315 103.111
R6562 CSoutput.n314 CSoutput.n313 103.111
R6563 CSoutput.n312 CSoutput.n311 103.111
R6564 CSoutput.n310 CSoutput.n309 103.111
R6565 CSoutput.n307 CSoutput.n306 103.111
R6566 CSoutput.n305 CSoutput.n304 103.111
R6567 CSoutput.n303 CSoutput.n302 103.111
R6568 CSoutput.n301 CSoutput.n300 103.111
R6569 CSoutput.n299 CSoutput.n298 103.111
R6570 CSoutput.n297 CSoutput.n296 103.111
R6571 CSoutput.n295 CSoutput.n294 103.111
R6572 CSoutput.n293 CSoutput.n292 103.111
R6573 CSoutput.n291 CSoutput.n290 103.111
R6574 CSoutput.n120 CSoutput.n119 103.111
R6575 CSoutput.n122 CSoutput.n121 103.111
R6576 CSoutput.n124 CSoutput.n123 103.111
R6577 CSoutput.n126 CSoutput.n125 103.111
R6578 CSoutput.n128 CSoutput.n127 103.111
R6579 CSoutput.n130 CSoutput.n129 103.111
R6580 CSoutput.n132 CSoutput.n131 103.111
R6581 CSoutput.n134 CSoutput.n133 103.111
R6582 CSoutput.n136 CSoutput.n135 103.111
R6583 CSoutput.n100 CSoutput.n99 103.111
R6584 CSoutput.n102 CSoutput.n101 103.111
R6585 CSoutput.n104 CSoutput.n103 103.111
R6586 CSoutput.n106 CSoutput.n105 103.111
R6587 CSoutput.n108 CSoutput.n107 103.111
R6588 CSoutput.n110 CSoutput.n109 103.111
R6589 CSoutput.n112 CSoutput.n111 103.111
R6590 CSoutput.n114 CSoutput.n113 103.111
R6591 CSoutput.n116 CSoutput.n115 103.111
R6592 CSoutput.n81 CSoutput.n80 103.111
R6593 CSoutput.n83 CSoutput.n82 103.111
R6594 CSoutput.n85 CSoutput.n84 103.111
R6595 CSoutput.n87 CSoutput.n86 103.111
R6596 CSoutput.n89 CSoutput.n88 103.111
R6597 CSoutput.n91 CSoutput.n90 103.111
R6598 CSoutput.n93 CSoutput.n92 103.111
R6599 CSoutput.n95 CSoutput.n94 103.111
R6600 CSoutput.n97 CSoutput.n96 103.111
R6601 CSoutput.n346 CSoutput.n345 103.111
R6602 CSoutput.n382 CSoutput.n380 81.5057
R6603 CSoutput.n366 CSoutput.n364 81.5057
R6604 CSoutput.n351 CSoutput.n349 81.5057
R6605 CSoutput.n430 CSoutput.n428 81.5057
R6606 CSoutput.n414 CSoutput.n412 81.5057
R6607 CSoutput.n399 CSoutput.n397 81.5057
R6608 CSoutput.n394 CSoutput.n393 80.9324
R6609 CSoutput.n392 CSoutput.n391 80.9324
R6610 CSoutput.n390 CSoutput.n389 80.9324
R6611 CSoutput.n388 CSoutput.n387 80.9324
R6612 CSoutput.n386 CSoutput.n385 80.9324
R6613 CSoutput.n384 CSoutput.n383 80.9324
R6614 CSoutput.n382 CSoutput.n381 80.9324
R6615 CSoutput.n378 CSoutput.n377 80.9324
R6616 CSoutput.n376 CSoutput.n375 80.9324
R6617 CSoutput.n374 CSoutput.n373 80.9324
R6618 CSoutput.n372 CSoutput.n371 80.9324
R6619 CSoutput.n370 CSoutput.n369 80.9324
R6620 CSoutput.n368 CSoutput.n367 80.9324
R6621 CSoutput.n366 CSoutput.n365 80.9324
R6622 CSoutput.n363 CSoutput.n362 80.9324
R6623 CSoutput.n361 CSoutput.n360 80.9324
R6624 CSoutput.n359 CSoutput.n358 80.9324
R6625 CSoutput.n357 CSoutput.n356 80.9324
R6626 CSoutput.n355 CSoutput.n354 80.9324
R6627 CSoutput.n353 CSoutput.n352 80.9324
R6628 CSoutput.n351 CSoutput.n350 80.9324
R6629 CSoutput.n430 CSoutput.n429 80.9324
R6630 CSoutput.n432 CSoutput.n431 80.9324
R6631 CSoutput.n434 CSoutput.n433 80.9324
R6632 CSoutput.n436 CSoutput.n435 80.9324
R6633 CSoutput.n438 CSoutput.n437 80.9324
R6634 CSoutput.n440 CSoutput.n439 80.9324
R6635 CSoutput.n442 CSoutput.n441 80.9324
R6636 CSoutput.n414 CSoutput.n413 80.9324
R6637 CSoutput.n416 CSoutput.n415 80.9324
R6638 CSoutput.n418 CSoutput.n417 80.9324
R6639 CSoutput.n420 CSoutput.n419 80.9324
R6640 CSoutput.n422 CSoutput.n421 80.9324
R6641 CSoutput.n424 CSoutput.n423 80.9324
R6642 CSoutput.n426 CSoutput.n425 80.9324
R6643 CSoutput.n399 CSoutput.n398 80.9324
R6644 CSoutput.n401 CSoutput.n400 80.9324
R6645 CSoutput.n403 CSoutput.n402 80.9324
R6646 CSoutput.n405 CSoutput.n404 80.9324
R6647 CSoutput.n407 CSoutput.n406 80.9324
R6648 CSoutput.n409 CSoutput.n408 80.9324
R6649 CSoutput.n411 CSoutput.n410 80.9324
R6650 CSoutput.n25 CSoutput.n24 48.1486
R6651 CSoutput.n69 CSoutput.n3 48.1486
R6652 CSoutput.n38 CSoutput.n37 48.1486
R6653 CSoutput.n42 CSoutput.n41 48.1486
R6654 CSoutput.n51 CSoutput.n50 48.1486
R6655 CSoutput.n55 CSoutput.n54 48.1486
R6656 CSoutput.n22 CSoutput.n17 46.462
R6657 CSoutput.n72 CSoutput.n71 46.462
R6658 CSoutput.n20 CSoutput.n19 44.9055
R6659 CSoutput.n29 CSoutput.n28 43.7635
R6660 CSoutput.n65 CSoutput.n63 43.7635
R6661 CSoutput.n35 CSoutput.n13 41.7396
R6662 CSoutput.n57 CSoutput.n5 41.7396
R6663 CSoutput.n44 CSoutput.n9 37.0171
R6664 CSoutput.n48 CSoutput.n9 37.0171
R6665 CSoutput.n76 CSoutput.n75 34.9932
R6666 CSoutput.n31 CSoutput.n13 32.2947
R6667 CSoutput.n61 CSoutput.n5 32.2947
R6668 CSoutput.n30 CSoutput.n29 29.6014
R6669 CSoutput.n63 CSoutput.n62 29.6014
R6670 CSoutput.n19 CSoutput.n18 28.4085
R6671 CSoutput.n18 CSoutput.n17 25.1176
R6672 CSoutput.n72 CSoutput.n1 25.1176
R6673 CSoutput.n43 CSoutput.n42 22.0922
R6674 CSoutput.n50 CSoutput.n49 22.0922
R6675 CSoutput.n77 CSoutput.n76 21.8586
R6676 CSoutput.n37 CSoutput.n36 18.9681
R6677 CSoutput.n56 CSoutput.n55 18.9681
R6678 CSoutput.n25 CSoutput.n15 17.6292
R6679 CSoutput.n64 CSoutput.n3 17.6292
R6680 CSoutput.n24 CSoutput.n23 15.844
R6681 CSoutput.n70 CSoutput.n69 15.844
R6682 CSoutput.n38 CSoutput.n11 14.5051
R6683 CSoutput.n54 CSoutput.n7 14.5051
R6684 CSoutput.n445 CSoutput.n78 11.4982
R6685 CSoutput.n41 CSoutput.n11 11.3811
R6686 CSoutput.n51 CSoutput.n7 11.3811
R6687 CSoutput.n23 CSoutput.n22 10.0422
R6688 CSoutput.n71 CSoutput.n70 10.0422
R6689 CSoutput.n327 CSoutput.n307 9.25285
R6690 CSoutput.n117 CSoutput.n97 9.25285
R6691 CSoutput.n379 CSoutput.n363 8.98182
R6692 CSoutput.n427 CSoutput.n411 8.98182
R6693 CSoutput.n396 CSoutput.n348 8.92798
R6694 CSoutput.n28 CSoutput.n15 8.25698
R6695 CSoutput.n65 CSoutput.n64 8.25698
R6696 CSoutput.n348 CSoutput.n347 7.12641
R6697 CSoutput.n138 CSoutput.n137 7.12641
R6698 CSoutput.n36 CSoutput.n35 6.91809
R6699 CSoutput.n57 CSoutput.n56 6.91809
R6700 CSoutput.n396 CSoutput.n395 6.02792
R6701 CSoutput.n444 CSoutput.n443 6.02792
R6702 CSoutput.n445 CSoutput.n138 5.33554
R6703 CSoutput.n395 CSoutput.n394 5.25266
R6704 CSoutput.n379 CSoutput.n378 5.25266
R6705 CSoutput.n443 CSoutput.n442 5.25266
R6706 CSoutput.n427 CSoutput.n426 5.25266
R6707 CSoutput.n347 CSoutput.n346 5.1449
R6708 CSoutput.n327 CSoutput.n326 5.1449
R6709 CSoutput.n137 CSoutput.n136 5.1449
R6710 CSoutput.n117 CSoutput.n116 5.1449
R6711 CSoutput.n229 CSoutput.n182 4.5005
R6712 CSoutput.n198 CSoutput.n182 4.5005
R6713 CSoutput.n193 CSoutput.n177 4.5005
R6714 CSoutput.n193 CSoutput.n179 4.5005
R6715 CSoutput.n193 CSoutput.n176 4.5005
R6716 CSoutput.n193 CSoutput.n180 4.5005
R6717 CSoutput.n193 CSoutput.n175 4.5005
R6718 CSoutput.n193 CSoutput.t233 4.5005
R6719 CSoutput.n193 CSoutput.n174 4.5005
R6720 CSoutput.n193 CSoutput.n181 4.5005
R6721 CSoutput.n193 CSoutput.n182 4.5005
R6722 CSoutput.n191 CSoutput.n177 4.5005
R6723 CSoutput.n191 CSoutput.n179 4.5005
R6724 CSoutput.n191 CSoutput.n176 4.5005
R6725 CSoutput.n191 CSoutput.n180 4.5005
R6726 CSoutput.n191 CSoutput.n175 4.5005
R6727 CSoutput.n191 CSoutput.t233 4.5005
R6728 CSoutput.n191 CSoutput.n174 4.5005
R6729 CSoutput.n191 CSoutput.n181 4.5005
R6730 CSoutput.n191 CSoutput.n182 4.5005
R6731 CSoutput.n190 CSoutput.n177 4.5005
R6732 CSoutput.n190 CSoutput.n179 4.5005
R6733 CSoutput.n190 CSoutput.n176 4.5005
R6734 CSoutput.n190 CSoutput.n180 4.5005
R6735 CSoutput.n190 CSoutput.n175 4.5005
R6736 CSoutput.n190 CSoutput.t233 4.5005
R6737 CSoutput.n190 CSoutput.n174 4.5005
R6738 CSoutput.n190 CSoutput.n181 4.5005
R6739 CSoutput.n190 CSoutput.n182 4.5005
R6740 CSoutput.n275 CSoutput.n177 4.5005
R6741 CSoutput.n275 CSoutput.n179 4.5005
R6742 CSoutput.n275 CSoutput.n176 4.5005
R6743 CSoutput.n275 CSoutput.n180 4.5005
R6744 CSoutput.n275 CSoutput.n175 4.5005
R6745 CSoutput.n275 CSoutput.t233 4.5005
R6746 CSoutput.n275 CSoutput.n174 4.5005
R6747 CSoutput.n275 CSoutput.n181 4.5005
R6748 CSoutput.n275 CSoutput.n182 4.5005
R6749 CSoutput.n273 CSoutput.n177 4.5005
R6750 CSoutput.n273 CSoutput.n179 4.5005
R6751 CSoutput.n273 CSoutput.n176 4.5005
R6752 CSoutput.n273 CSoutput.n180 4.5005
R6753 CSoutput.n273 CSoutput.n175 4.5005
R6754 CSoutput.n273 CSoutput.t233 4.5005
R6755 CSoutput.n273 CSoutput.n174 4.5005
R6756 CSoutput.n273 CSoutput.n181 4.5005
R6757 CSoutput.n271 CSoutput.n177 4.5005
R6758 CSoutput.n271 CSoutput.n179 4.5005
R6759 CSoutput.n271 CSoutput.n176 4.5005
R6760 CSoutput.n271 CSoutput.n180 4.5005
R6761 CSoutput.n271 CSoutput.n175 4.5005
R6762 CSoutput.n271 CSoutput.t233 4.5005
R6763 CSoutput.n271 CSoutput.n174 4.5005
R6764 CSoutput.n271 CSoutput.n181 4.5005
R6765 CSoutput.n201 CSoutput.n177 4.5005
R6766 CSoutput.n201 CSoutput.n179 4.5005
R6767 CSoutput.n201 CSoutput.n176 4.5005
R6768 CSoutput.n201 CSoutput.n180 4.5005
R6769 CSoutput.n201 CSoutput.n175 4.5005
R6770 CSoutput.n201 CSoutput.t233 4.5005
R6771 CSoutput.n201 CSoutput.n174 4.5005
R6772 CSoutput.n201 CSoutput.n181 4.5005
R6773 CSoutput.n201 CSoutput.n182 4.5005
R6774 CSoutput.n200 CSoutput.n177 4.5005
R6775 CSoutput.n200 CSoutput.n179 4.5005
R6776 CSoutput.n200 CSoutput.n176 4.5005
R6777 CSoutput.n200 CSoutput.n180 4.5005
R6778 CSoutput.n200 CSoutput.n175 4.5005
R6779 CSoutput.n200 CSoutput.t233 4.5005
R6780 CSoutput.n200 CSoutput.n174 4.5005
R6781 CSoutput.n200 CSoutput.n181 4.5005
R6782 CSoutput.n200 CSoutput.n182 4.5005
R6783 CSoutput.n204 CSoutput.n177 4.5005
R6784 CSoutput.n204 CSoutput.n179 4.5005
R6785 CSoutput.n204 CSoutput.n176 4.5005
R6786 CSoutput.n204 CSoutput.n180 4.5005
R6787 CSoutput.n204 CSoutput.n175 4.5005
R6788 CSoutput.n204 CSoutput.t233 4.5005
R6789 CSoutput.n204 CSoutput.n174 4.5005
R6790 CSoutput.n204 CSoutput.n181 4.5005
R6791 CSoutput.n204 CSoutput.n182 4.5005
R6792 CSoutput.n203 CSoutput.n177 4.5005
R6793 CSoutput.n203 CSoutput.n179 4.5005
R6794 CSoutput.n203 CSoutput.n176 4.5005
R6795 CSoutput.n203 CSoutput.n180 4.5005
R6796 CSoutput.n203 CSoutput.n175 4.5005
R6797 CSoutput.n203 CSoutput.t233 4.5005
R6798 CSoutput.n203 CSoutput.n174 4.5005
R6799 CSoutput.n203 CSoutput.n181 4.5005
R6800 CSoutput.n203 CSoutput.n182 4.5005
R6801 CSoutput.n186 CSoutput.n177 4.5005
R6802 CSoutput.n186 CSoutput.n179 4.5005
R6803 CSoutput.n186 CSoutput.n176 4.5005
R6804 CSoutput.n186 CSoutput.n180 4.5005
R6805 CSoutput.n186 CSoutput.n175 4.5005
R6806 CSoutput.n186 CSoutput.t233 4.5005
R6807 CSoutput.n186 CSoutput.n174 4.5005
R6808 CSoutput.n186 CSoutput.n181 4.5005
R6809 CSoutput.n186 CSoutput.n182 4.5005
R6810 CSoutput.n278 CSoutput.n177 4.5005
R6811 CSoutput.n278 CSoutput.n179 4.5005
R6812 CSoutput.n278 CSoutput.n176 4.5005
R6813 CSoutput.n278 CSoutput.n180 4.5005
R6814 CSoutput.n278 CSoutput.n175 4.5005
R6815 CSoutput.n278 CSoutput.t233 4.5005
R6816 CSoutput.n278 CSoutput.n174 4.5005
R6817 CSoutput.n278 CSoutput.n181 4.5005
R6818 CSoutput.n278 CSoutput.n182 4.5005
R6819 CSoutput.n265 CSoutput.n236 4.5005
R6820 CSoutput.n265 CSoutput.n242 4.5005
R6821 CSoutput.n223 CSoutput.n212 4.5005
R6822 CSoutput.n223 CSoutput.n214 4.5005
R6823 CSoutput.n223 CSoutput.n211 4.5005
R6824 CSoutput.n223 CSoutput.n215 4.5005
R6825 CSoutput.n223 CSoutput.n210 4.5005
R6826 CSoutput.n223 CSoutput.t226 4.5005
R6827 CSoutput.n223 CSoutput.n209 4.5005
R6828 CSoutput.n223 CSoutput.n216 4.5005
R6829 CSoutput.n265 CSoutput.n223 4.5005
R6830 CSoutput.n244 CSoutput.n212 4.5005
R6831 CSoutput.n244 CSoutput.n214 4.5005
R6832 CSoutput.n244 CSoutput.n211 4.5005
R6833 CSoutput.n244 CSoutput.n215 4.5005
R6834 CSoutput.n244 CSoutput.n210 4.5005
R6835 CSoutput.n244 CSoutput.t226 4.5005
R6836 CSoutput.n244 CSoutput.n209 4.5005
R6837 CSoutput.n244 CSoutput.n216 4.5005
R6838 CSoutput.n265 CSoutput.n244 4.5005
R6839 CSoutput.n222 CSoutput.n212 4.5005
R6840 CSoutput.n222 CSoutput.n214 4.5005
R6841 CSoutput.n222 CSoutput.n211 4.5005
R6842 CSoutput.n222 CSoutput.n215 4.5005
R6843 CSoutput.n222 CSoutput.n210 4.5005
R6844 CSoutput.n222 CSoutput.t226 4.5005
R6845 CSoutput.n222 CSoutput.n209 4.5005
R6846 CSoutput.n222 CSoutput.n216 4.5005
R6847 CSoutput.n265 CSoutput.n222 4.5005
R6848 CSoutput.n246 CSoutput.n212 4.5005
R6849 CSoutput.n246 CSoutput.n214 4.5005
R6850 CSoutput.n246 CSoutput.n211 4.5005
R6851 CSoutput.n246 CSoutput.n215 4.5005
R6852 CSoutput.n246 CSoutput.n210 4.5005
R6853 CSoutput.n246 CSoutput.t226 4.5005
R6854 CSoutput.n246 CSoutput.n209 4.5005
R6855 CSoutput.n246 CSoutput.n216 4.5005
R6856 CSoutput.n265 CSoutput.n246 4.5005
R6857 CSoutput.n212 CSoutput.n207 4.5005
R6858 CSoutput.n214 CSoutput.n207 4.5005
R6859 CSoutput.n211 CSoutput.n207 4.5005
R6860 CSoutput.n215 CSoutput.n207 4.5005
R6861 CSoutput.n210 CSoutput.n207 4.5005
R6862 CSoutput.t226 CSoutput.n207 4.5005
R6863 CSoutput.n209 CSoutput.n207 4.5005
R6864 CSoutput.n216 CSoutput.n207 4.5005
R6865 CSoutput.n268 CSoutput.n212 4.5005
R6866 CSoutput.n268 CSoutput.n214 4.5005
R6867 CSoutput.n268 CSoutput.n211 4.5005
R6868 CSoutput.n268 CSoutput.n215 4.5005
R6869 CSoutput.n268 CSoutput.n210 4.5005
R6870 CSoutput.n268 CSoutput.t226 4.5005
R6871 CSoutput.n268 CSoutput.n209 4.5005
R6872 CSoutput.n268 CSoutput.n216 4.5005
R6873 CSoutput.n266 CSoutput.n212 4.5005
R6874 CSoutput.n266 CSoutput.n214 4.5005
R6875 CSoutput.n266 CSoutput.n211 4.5005
R6876 CSoutput.n266 CSoutput.n215 4.5005
R6877 CSoutput.n266 CSoutput.n210 4.5005
R6878 CSoutput.n266 CSoutput.t226 4.5005
R6879 CSoutput.n266 CSoutput.n209 4.5005
R6880 CSoutput.n266 CSoutput.n216 4.5005
R6881 CSoutput.n266 CSoutput.n265 4.5005
R6882 CSoutput.n248 CSoutput.n212 4.5005
R6883 CSoutput.n248 CSoutput.n214 4.5005
R6884 CSoutput.n248 CSoutput.n211 4.5005
R6885 CSoutput.n248 CSoutput.n215 4.5005
R6886 CSoutput.n248 CSoutput.n210 4.5005
R6887 CSoutput.n248 CSoutput.t226 4.5005
R6888 CSoutput.n248 CSoutput.n209 4.5005
R6889 CSoutput.n248 CSoutput.n216 4.5005
R6890 CSoutput.n265 CSoutput.n248 4.5005
R6891 CSoutput.n220 CSoutput.n212 4.5005
R6892 CSoutput.n220 CSoutput.n214 4.5005
R6893 CSoutput.n220 CSoutput.n211 4.5005
R6894 CSoutput.n220 CSoutput.n215 4.5005
R6895 CSoutput.n220 CSoutput.n210 4.5005
R6896 CSoutput.n220 CSoutput.t226 4.5005
R6897 CSoutput.n220 CSoutput.n209 4.5005
R6898 CSoutput.n220 CSoutput.n216 4.5005
R6899 CSoutput.n265 CSoutput.n220 4.5005
R6900 CSoutput.n250 CSoutput.n212 4.5005
R6901 CSoutput.n250 CSoutput.n214 4.5005
R6902 CSoutput.n250 CSoutput.n211 4.5005
R6903 CSoutput.n250 CSoutput.n215 4.5005
R6904 CSoutput.n250 CSoutput.n210 4.5005
R6905 CSoutput.n250 CSoutput.t226 4.5005
R6906 CSoutput.n250 CSoutput.n209 4.5005
R6907 CSoutput.n250 CSoutput.n216 4.5005
R6908 CSoutput.n265 CSoutput.n250 4.5005
R6909 CSoutput.n219 CSoutput.n212 4.5005
R6910 CSoutput.n219 CSoutput.n214 4.5005
R6911 CSoutput.n219 CSoutput.n211 4.5005
R6912 CSoutput.n219 CSoutput.n215 4.5005
R6913 CSoutput.n219 CSoutput.n210 4.5005
R6914 CSoutput.n219 CSoutput.t226 4.5005
R6915 CSoutput.n219 CSoutput.n209 4.5005
R6916 CSoutput.n219 CSoutput.n216 4.5005
R6917 CSoutput.n265 CSoutput.n219 4.5005
R6918 CSoutput.n264 CSoutput.n212 4.5005
R6919 CSoutput.n264 CSoutput.n214 4.5005
R6920 CSoutput.n264 CSoutput.n211 4.5005
R6921 CSoutput.n264 CSoutput.n215 4.5005
R6922 CSoutput.n264 CSoutput.n210 4.5005
R6923 CSoutput.n264 CSoutput.t226 4.5005
R6924 CSoutput.n264 CSoutput.n209 4.5005
R6925 CSoutput.n264 CSoutput.n216 4.5005
R6926 CSoutput.n265 CSoutput.n264 4.5005
R6927 CSoutput.n263 CSoutput.n148 4.5005
R6928 CSoutput.n164 CSoutput.n148 4.5005
R6929 CSoutput.n159 CSoutput.n143 4.5005
R6930 CSoutput.n159 CSoutput.n145 4.5005
R6931 CSoutput.n159 CSoutput.n142 4.5005
R6932 CSoutput.n159 CSoutput.n146 4.5005
R6933 CSoutput.n159 CSoutput.n141 4.5005
R6934 CSoutput.n159 CSoutput.t216 4.5005
R6935 CSoutput.n159 CSoutput.n140 4.5005
R6936 CSoutput.n159 CSoutput.n147 4.5005
R6937 CSoutput.n159 CSoutput.n148 4.5005
R6938 CSoutput.n157 CSoutput.n143 4.5005
R6939 CSoutput.n157 CSoutput.n145 4.5005
R6940 CSoutput.n157 CSoutput.n142 4.5005
R6941 CSoutput.n157 CSoutput.n146 4.5005
R6942 CSoutput.n157 CSoutput.n141 4.5005
R6943 CSoutput.n157 CSoutput.t216 4.5005
R6944 CSoutput.n157 CSoutput.n140 4.5005
R6945 CSoutput.n157 CSoutput.n147 4.5005
R6946 CSoutput.n157 CSoutput.n148 4.5005
R6947 CSoutput.n156 CSoutput.n143 4.5005
R6948 CSoutput.n156 CSoutput.n145 4.5005
R6949 CSoutput.n156 CSoutput.n142 4.5005
R6950 CSoutput.n156 CSoutput.n146 4.5005
R6951 CSoutput.n156 CSoutput.n141 4.5005
R6952 CSoutput.n156 CSoutput.t216 4.5005
R6953 CSoutput.n156 CSoutput.n140 4.5005
R6954 CSoutput.n156 CSoutput.n147 4.5005
R6955 CSoutput.n156 CSoutput.n148 4.5005
R6956 CSoutput.n285 CSoutput.n143 4.5005
R6957 CSoutput.n285 CSoutput.n145 4.5005
R6958 CSoutput.n285 CSoutput.n142 4.5005
R6959 CSoutput.n285 CSoutput.n146 4.5005
R6960 CSoutput.n285 CSoutput.n141 4.5005
R6961 CSoutput.n285 CSoutput.t216 4.5005
R6962 CSoutput.n285 CSoutput.n140 4.5005
R6963 CSoutput.n285 CSoutput.n147 4.5005
R6964 CSoutput.n285 CSoutput.n148 4.5005
R6965 CSoutput.n283 CSoutput.n143 4.5005
R6966 CSoutput.n283 CSoutput.n145 4.5005
R6967 CSoutput.n283 CSoutput.n142 4.5005
R6968 CSoutput.n283 CSoutput.n146 4.5005
R6969 CSoutput.n283 CSoutput.n141 4.5005
R6970 CSoutput.n283 CSoutput.t216 4.5005
R6971 CSoutput.n283 CSoutput.n140 4.5005
R6972 CSoutput.n283 CSoutput.n147 4.5005
R6973 CSoutput.n281 CSoutput.n143 4.5005
R6974 CSoutput.n281 CSoutput.n145 4.5005
R6975 CSoutput.n281 CSoutput.n142 4.5005
R6976 CSoutput.n281 CSoutput.n146 4.5005
R6977 CSoutput.n281 CSoutput.n141 4.5005
R6978 CSoutput.n281 CSoutput.t216 4.5005
R6979 CSoutput.n281 CSoutput.n140 4.5005
R6980 CSoutput.n281 CSoutput.n147 4.5005
R6981 CSoutput.n167 CSoutput.n143 4.5005
R6982 CSoutput.n167 CSoutput.n145 4.5005
R6983 CSoutput.n167 CSoutput.n142 4.5005
R6984 CSoutput.n167 CSoutput.n146 4.5005
R6985 CSoutput.n167 CSoutput.n141 4.5005
R6986 CSoutput.n167 CSoutput.t216 4.5005
R6987 CSoutput.n167 CSoutput.n140 4.5005
R6988 CSoutput.n167 CSoutput.n147 4.5005
R6989 CSoutput.n167 CSoutput.n148 4.5005
R6990 CSoutput.n166 CSoutput.n143 4.5005
R6991 CSoutput.n166 CSoutput.n145 4.5005
R6992 CSoutput.n166 CSoutput.n142 4.5005
R6993 CSoutput.n166 CSoutput.n146 4.5005
R6994 CSoutput.n166 CSoutput.n141 4.5005
R6995 CSoutput.n166 CSoutput.t216 4.5005
R6996 CSoutput.n166 CSoutput.n140 4.5005
R6997 CSoutput.n166 CSoutput.n147 4.5005
R6998 CSoutput.n166 CSoutput.n148 4.5005
R6999 CSoutput.n170 CSoutput.n143 4.5005
R7000 CSoutput.n170 CSoutput.n145 4.5005
R7001 CSoutput.n170 CSoutput.n142 4.5005
R7002 CSoutput.n170 CSoutput.n146 4.5005
R7003 CSoutput.n170 CSoutput.n141 4.5005
R7004 CSoutput.n170 CSoutput.t216 4.5005
R7005 CSoutput.n170 CSoutput.n140 4.5005
R7006 CSoutput.n170 CSoutput.n147 4.5005
R7007 CSoutput.n170 CSoutput.n148 4.5005
R7008 CSoutput.n169 CSoutput.n143 4.5005
R7009 CSoutput.n169 CSoutput.n145 4.5005
R7010 CSoutput.n169 CSoutput.n142 4.5005
R7011 CSoutput.n169 CSoutput.n146 4.5005
R7012 CSoutput.n169 CSoutput.n141 4.5005
R7013 CSoutput.n169 CSoutput.t216 4.5005
R7014 CSoutput.n169 CSoutput.n140 4.5005
R7015 CSoutput.n169 CSoutput.n147 4.5005
R7016 CSoutput.n169 CSoutput.n148 4.5005
R7017 CSoutput.n152 CSoutput.n143 4.5005
R7018 CSoutput.n152 CSoutput.n145 4.5005
R7019 CSoutput.n152 CSoutput.n142 4.5005
R7020 CSoutput.n152 CSoutput.n146 4.5005
R7021 CSoutput.n152 CSoutput.n141 4.5005
R7022 CSoutput.n152 CSoutput.t216 4.5005
R7023 CSoutput.n152 CSoutput.n140 4.5005
R7024 CSoutput.n152 CSoutput.n147 4.5005
R7025 CSoutput.n152 CSoutput.n148 4.5005
R7026 CSoutput.n288 CSoutput.n143 4.5005
R7027 CSoutput.n288 CSoutput.n145 4.5005
R7028 CSoutput.n288 CSoutput.n142 4.5005
R7029 CSoutput.n288 CSoutput.n146 4.5005
R7030 CSoutput.n288 CSoutput.n141 4.5005
R7031 CSoutput.n288 CSoutput.t216 4.5005
R7032 CSoutput.n288 CSoutput.n140 4.5005
R7033 CSoutput.n288 CSoutput.n147 4.5005
R7034 CSoutput.n288 CSoutput.n148 4.5005
R7035 CSoutput.n347 CSoutput.n327 4.10845
R7036 CSoutput.n137 CSoutput.n117 4.10845
R7037 CSoutput.n345 CSoutput.t140 4.06363
R7038 CSoutput.n345 CSoutput.t164 4.06363
R7039 CSoutput.n343 CSoutput.t184 4.06363
R7040 CSoutput.n343 CSoutput.t98 4.06363
R7041 CSoutput.n341 CSoutput.t102 4.06363
R7042 CSoutput.n341 CSoutput.t168 4.06363
R7043 CSoutput.n339 CSoutput.t187 4.06363
R7044 CSoutput.n339 CSoutput.t188 4.06363
R7045 CSoutput.n337 CSoutput.t118 4.06363
R7046 CSoutput.n337 CSoutput.t119 4.06363
R7047 CSoutput.n335 CSoutput.t124 4.06363
R7048 CSoutput.n335 CSoutput.t189 4.06363
R7049 CSoutput.n333 CSoutput.t88 4.06363
R7050 CSoutput.n333 CSoutput.t122 4.06363
R7051 CSoutput.n331 CSoutput.t139 4.06363
R7052 CSoutput.n331 CSoutput.t163 4.06363
R7053 CSoutput.n329 CSoutput.t170 4.06363
R7054 CSoutput.n329 CSoutput.t94 4.06363
R7055 CSoutput.n328 CSoutput.t142 4.06363
R7056 CSoutput.n328 CSoutput.t143 4.06363
R7057 CSoutput.n325 CSoutput.t125 4.06363
R7058 CSoutput.n325 CSoutput.t152 4.06363
R7059 CSoutput.n323 CSoutput.t172 4.06363
R7060 CSoutput.n323 CSoutput.t84 4.06363
R7061 CSoutput.n321 CSoutput.t85 4.06363
R7062 CSoutput.n321 CSoutput.t154 4.06363
R7063 CSoutput.n319 CSoutput.t175 4.06363
R7064 CSoutput.n319 CSoutput.t176 4.06363
R7065 CSoutput.n317 CSoutput.t106 4.06363
R7066 CSoutput.n317 CSoutput.t107 4.06363
R7067 CSoutput.n315 CSoutput.t110 4.06363
R7068 CSoutput.n315 CSoutput.t179 4.06363
R7069 CSoutput.n313 CSoutput.t73 4.06363
R7070 CSoutput.n313 CSoutput.t109 4.06363
R7071 CSoutput.n311 CSoutput.t126 4.06363
R7072 CSoutput.n311 CSoutput.t153 4.06363
R7073 CSoutput.n309 CSoutput.t155 4.06363
R7074 CSoutput.n309 CSoutput.t79 4.06363
R7075 CSoutput.n308 CSoutput.t132 4.06363
R7076 CSoutput.n308 CSoutput.t133 4.06363
R7077 CSoutput.n306 CSoutput.t161 4.06363
R7078 CSoutput.n306 CSoutput.t115 4.06363
R7079 CSoutput.n304 CSoutput.t148 4.06363
R7080 CSoutput.n304 CSoutput.t97 4.06363
R7081 CSoutput.n302 CSoutput.t173 4.06363
R7082 CSoutput.n302 CSoutput.t89 4.06363
R7083 CSoutput.n300 CSoutput.t129 4.06363
R7084 CSoutput.n300 CSoutput.t108 4.06363
R7085 CSoutput.n298 CSoutput.t111 4.06363
R7086 CSoutput.n298 CSoutput.t86 4.06363
R7087 CSoutput.n296 CSoutput.t160 4.06363
R7088 CSoutput.n296 CSoutput.t80 4.06363
R7089 CSoutput.n294 CSoutput.t120 4.06363
R7090 CSoutput.n294 CSoutput.t185 4.06363
R7091 CSoutput.n292 CSoutput.t103 4.06363
R7092 CSoutput.n292 CSoutput.t166 4.06363
R7093 CSoutput.n290 CSoutput.t127 4.06363
R7094 CSoutput.n290 CSoutput.t190 4.06363
R7095 CSoutput.n289 CSoutput.t74 4.06363
R7096 CSoutput.n289 CSoutput.t177 4.06363
R7097 CSoutput.n118 CSoutput.t183 4.06363
R7098 CSoutput.n118 CSoutput.t182 4.06363
R7099 CSoutput.n119 CSoutput.t162 4.06363
R7100 CSoutput.n119 CSoutput.t96 4.06363
R7101 CSoutput.n121 CSoutput.t93 4.06363
R7102 CSoutput.n121 CSoutput.t180 4.06363
R7103 CSoutput.n123 CSoutput.t159 4.06363
R7104 CSoutput.n123 CSoutput.t136 4.06363
R7105 CSoutput.n125 CSoutput.t117 4.06363
R7106 CSoutput.n125 CSoutput.t192 4.06363
R7107 CSoutput.n127 CSoutput.t157 4.06363
R7108 CSoutput.n127 CSoutput.t156 4.06363
R7109 CSoutput.n129 CSoutput.t144 4.06363
R7110 CSoutput.n129 CSoutput.t114 4.06363
R7111 CSoutput.n131 CSoutput.t95 4.06363
R7112 CSoutput.n131 CSoutput.t145 4.06363
R7113 CSoutput.n133 CSoutput.t141 4.06363
R7114 CSoutput.n133 CSoutput.t112 4.06363
R7115 CSoutput.n135 CSoutput.t92 4.06363
R7116 CSoutput.n135 CSoutput.t91 4.06363
R7117 CSoutput.n98 CSoutput.t171 4.06363
R7118 CSoutput.n98 CSoutput.t169 4.06363
R7119 CSoutput.n99 CSoutput.t151 4.06363
R7120 CSoutput.n99 CSoutput.t83 4.06363
R7121 CSoutput.n101 CSoutput.t77 4.06363
R7122 CSoutput.n101 CSoutput.t165 4.06363
R7123 CSoutput.n103 CSoutput.t150 4.06363
R7124 CSoutput.n103 CSoutput.t123 4.06363
R7125 CSoutput.n105 CSoutput.t105 4.06363
R7126 CSoutput.n105 CSoutput.t181 4.06363
R7127 CSoutput.n107 CSoutput.t147 4.06363
R7128 CSoutput.n107 CSoutput.t146 4.06363
R7129 CSoutput.n109 CSoutput.t134 4.06363
R7130 CSoutput.n109 CSoutput.t101 4.06363
R7131 CSoutput.n111 CSoutput.t81 4.06363
R7132 CSoutput.n111 CSoutput.t135 4.06363
R7133 CSoutput.n113 CSoutput.t131 4.06363
R7134 CSoutput.n113 CSoutput.t99 4.06363
R7135 CSoutput.n115 CSoutput.t78 4.06363
R7136 CSoutput.n115 CSoutput.t75 4.06363
R7137 CSoutput.n79 CSoutput.t178 4.06363
R7138 CSoutput.n79 CSoutput.t76 4.06363
R7139 CSoutput.n80 CSoutput.t158 4.06363
R7140 CSoutput.n80 CSoutput.t128 4.06363
R7141 CSoutput.n82 CSoutput.t167 4.06363
R7142 CSoutput.n82 CSoutput.t104 4.06363
R7143 CSoutput.n84 CSoutput.t186 4.06363
R7144 CSoutput.n84 CSoutput.t121 4.06363
R7145 CSoutput.n86 CSoutput.t82 4.06363
R7146 CSoutput.n86 CSoutput.t137 4.06363
R7147 CSoutput.n88 CSoutput.t87 4.06363
R7148 CSoutput.n88 CSoutput.t113 4.06363
R7149 CSoutput.n90 CSoutput.t191 4.06363
R7150 CSoutput.n90 CSoutput.t130 4.06363
R7151 CSoutput.n92 CSoutput.t90 4.06363
R7152 CSoutput.n92 CSoutput.t174 4.06363
R7153 CSoutput.n94 CSoutput.t100 4.06363
R7154 CSoutput.n94 CSoutput.t149 4.06363
R7155 CSoutput.n96 CSoutput.t116 4.06363
R7156 CSoutput.n96 CSoutput.t138 4.06363
R7157 CSoutput.n44 CSoutput.n43 3.79402
R7158 CSoutput.n49 CSoutput.n48 3.79402
R7159 CSoutput.n395 CSoutput.n379 3.72967
R7160 CSoutput.n443 CSoutput.n427 3.72967
R7161 CSoutput.n445 CSoutput.n444 3.57343
R7162 CSoutput.n444 CSoutput.n396 3.3798
R7163 CSoutput.n393 CSoutput.t208 2.82907
R7164 CSoutput.n393 CSoutput.t7 2.82907
R7165 CSoutput.n391 CSoutput.t8 2.82907
R7166 CSoutput.n391 CSoutput.t68 2.82907
R7167 CSoutput.n389 CSoutput.t47 2.82907
R7168 CSoutput.n389 CSoutput.t9 2.82907
R7169 CSoutput.n387 CSoutput.t210 2.82907
R7170 CSoutput.n387 CSoutput.t24 2.82907
R7171 CSoutput.n385 CSoutput.t40 2.82907
R7172 CSoutput.n385 CSoutput.t33 2.82907
R7173 CSoutput.n383 CSoutput.t58 2.82907
R7174 CSoutput.n383 CSoutput.t14 2.82907
R7175 CSoutput.n381 CSoutput.t23 2.82907
R7176 CSoutput.n381 CSoutput.t13 2.82907
R7177 CSoutput.n380 CSoutput.t193 2.82907
R7178 CSoutput.n380 CSoutput.t198 2.82907
R7179 CSoutput.n377 CSoutput.t6 2.82907
R7180 CSoutput.n377 CSoutput.t42 2.82907
R7181 CSoutput.n375 CSoutput.t72 2.82907
R7182 CSoutput.n375 CSoutput.t199 2.82907
R7183 CSoutput.n373 CSoutput.t197 2.82907
R7184 CSoutput.n373 CSoutput.t213 2.82907
R7185 CSoutput.n371 CSoutput.t10 2.82907
R7186 CSoutput.n371 CSoutput.t194 2.82907
R7187 CSoutput.n369 CSoutput.t64 2.82907
R7188 CSoutput.n369 CSoutput.t66 2.82907
R7189 CSoutput.n367 CSoutput.t26 2.82907
R7190 CSoutput.n367 CSoutput.t204 2.82907
R7191 CSoutput.n365 CSoutput.t214 2.82907
R7192 CSoutput.n365 CSoutput.t12 2.82907
R7193 CSoutput.n364 CSoutput.t3 2.82907
R7194 CSoutput.n364 CSoutput.t215 2.82907
R7195 CSoutput.n362 CSoutput.t17 2.82907
R7196 CSoutput.n362 CSoutput.t41 2.82907
R7197 CSoutput.n360 CSoutput.t39 2.82907
R7198 CSoutput.n360 CSoutput.t35 2.82907
R7199 CSoutput.n358 CSoutput.t37 2.82907
R7200 CSoutput.n358 CSoutput.t203 2.82907
R7201 CSoutput.n356 CSoutput.t18 2.82907
R7202 CSoutput.n356 CSoutput.t16 2.82907
R7203 CSoutput.n354 CSoutput.t50 2.82907
R7204 CSoutput.n354 CSoutput.t207 2.82907
R7205 CSoutput.n352 CSoutput.t29 2.82907
R7206 CSoutput.n352 CSoutput.t15 2.82907
R7207 CSoutput.n350 CSoutput.t200 2.82907
R7208 CSoutput.n350 CSoutput.t0 2.82907
R7209 CSoutput.n349 CSoutput.t19 2.82907
R7210 CSoutput.n349 CSoutput.t55 2.82907
R7211 CSoutput.n428 CSoutput.t27 2.82907
R7212 CSoutput.n428 CSoutput.t69 2.82907
R7213 CSoutput.n429 CSoutput.t209 2.82907
R7214 CSoutput.n429 CSoutput.t1 2.82907
R7215 CSoutput.n431 CSoutput.t38 2.82907
R7216 CSoutput.n431 CSoutput.t60 2.82907
R7217 CSoutput.n433 CSoutput.t71 2.82907
R7218 CSoutput.n433 CSoutput.t201 2.82907
R7219 CSoutput.n435 CSoutput.t67 2.82907
R7220 CSoutput.n435 CSoutput.t32 2.82907
R7221 CSoutput.n437 CSoutput.t59 2.82907
R7222 CSoutput.n437 CSoutput.t44 2.82907
R7223 CSoutput.n439 CSoutput.t206 2.82907
R7224 CSoutput.n439 CSoutput.t52 2.82907
R7225 CSoutput.n441 CSoutput.t11 2.82907
R7226 CSoutput.n441 CSoutput.t34 2.82907
R7227 CSoutput.n412 CSoutput.t4 2.82907
R7228 CSoutput.n412 CSoutput.t2 2.82907
R7229 CSoutput.n413 CSoutput.t46 2.82907
R7230 CSoutput.n413 CSoutput.t25 2.82907
R7231 CSoutput.n415 CSoutput.t21 2.82907
R7232 CSoutput.n415 CSoutput.t48 2.82907
R7233 CSoutput.n417 CSoutput.t212 2.82907
R7234 CSoutput.n417 CSoutput.t5 2.82907
R7235 CSoutput.n419 CSoutput.t65 2.82907
R7236 CSoutput.n419 CSoutput.t63 2.82907
R7237 CSoutput.n421 CSoutput.t54 2.82907
R7238 CSoutput.n421 CSoutput.t57 2.82907
R7239 CSoutput.n423 CSoutput.t195 2.82907
R7240 CSoutput.n423 CSoutput.t22 2.82907
R7241 CSoutput.n425 CSoutput.t196 2.82907
R7242 CSoutput.n425 CSoutput.t30 2.82907
R7243 CSoutput.n397 CSoutput.t70 2.82907
R7244 CSoutput.n397 CSoutput.t51 2.82907
R7245 CSoutput.n398 CSoutput.t49 2.82907
R7246 CSoutput.n398 CSoutput.t53 2.82907
R7247 CSoutput.n400 CSoutput.t56 2.82907
R7248 CSoutput.n400 CSoutput.t61 2.82907
R7249 CSoutput.n402 CSoutput.t62 2.82907
R7250 CSoutput.n402 CSoutput.t211 2.82907
R7251 CSoutput.n404 CSoutput.t28 2.82907
R7252 CSoutput.n404 CSoutput.t202 2.82907
R7253 CSoutput.n406 CSoutput.t45 2.82907
R7254 CSoutput.n406 CSoutput.t20 2.82907
R7255 CSoutput.n408 CSoutput.t43 2.82907
R7256 CSoutput.n408 CSoutput.t205 2.82907
R7257 CSoutput.n410 CSoutput.t36 2.82907
R7258 CSoutput.n410 CSoutput.t31 2.82907
R7259 CSoutput.n348 CSoutput.n138 2.57547
R7260 CSoutput.n75 CSoutput.n1 2.45513
R7261 CSoutput.n229 CSoutput.n227 2.251
R7262 CSoutput.n229 CSoutput.n226 2.251
R7263 CSoutput.n229 CSoutput.n225 2.251
R7264 CSoutput.n229 CSoutput.n224 2.251
R7265 CSoutput.n198 CSoutput.n197 2.251
R7266 CSoutput.n198 CSoutput.n196 2.251
R7267 CSoutput.n198 CSoutput.n195 2.251
R7268 CSoutput.n198 CSoutput.n194 2.251
R7269 CSoutput.n271 CSoutput.n270 2.251
R7270 CSoutput.n236 CSoutput.n234 2.251
R7271 CSoutput.n236 CSoutput.n233 2.251
R7272 CSoutput.n236 CSoutput.n232 2.251
R7273 CSoutput.n254 CSoutput.n236 2.251
R7274 CSoutput.n242 CSoutput.n241 2.251
R7275 CSoutput.n242 CSoutput.n240 2.251
R7276 CSoutput.n242 CSoutput.n239 2.251
R7277 CSoutput.n242 CSoutput.n238 2.251
R7278 CSoutput.n268 CSoutput.n208 2.251
R7279 CSoutput.n263 CSoutput.n261 2.251
R7280 CSoutput.n263 CSoutput.n260 2.251
R7281 CSoutput.n263 CSoutput.n259 2.251
R7282 CSoutput.n263 CSoutput.n258 2.251
R7283 CSoutput.n164 CSoutput.n163 2.251
R7284 CSoutput.n164 CSoutput.n162 2.251
R7285 CSoutput.n164 CSoutput.n161 2.251
R7286 CSoutput.n164 CSoutput.n160 2.251
R7287 CSoutput.n281 CSoutput.n280 2.251
R7288 CSoutput.n198 CSoutput.n178 2.2505
R7289 CSoutput.n193 CSoutput.n178 2.2505
R7290 CSoutput.n191 CSoutput.n178 2.2505
R7291 CSoutput.n190 CSoutput.n178 2.2505
R7292 CSoutput.n275 CSoutput.n178 2.2505
R7293 CSoutput.n273 CSoutput.n178 2.2505
R7294 CSoutput.n271 CSoutput.n178 2.2505
R7295 CSoutput.n201 CSoutput.n178 2.2505
R7296 CSoutput.n200 CSoutput.n178 2.2505
R7297 CSoutput.n204 CSoutput.n178 2.2505
R7298 CSoutput.n203 CSoutput.n178 2.2505
R7299 CSoutput.n186 CSoutput.n178 2.2505
R7300 CSoutput.n278 CSoutput.n178 2.2505
R7301 CSoutput.n278 CSoutput.n277 2.2505
R7302 CSoutput.n242 CSoutput.n213 2.2505
R7303 CSoutput.n223 CSoutput.n213 2.2505
R7304 CSoutput.n244 CSoutput.n213 2.2505
R7305 CSoutput.n222 CSoutput.n213 2.2505
R7306 CSoutput.n246 CSoutput.n213 2.2505
R7307 CSoutput.n213 CSoutput.n207 2.2505
R7308 CSoutput.n268 CSoutput.n213 2.2505
R7309 CSoutput.n266 CSoutput.n213 2.2505
R7310 CSoutput.n248 CSoutput.n213 2.2505
R7311 CSoutput.n220 CSoutput.n213 2.2505
R7312 CSoutput.n250 CSoutput.n213 2.2505
R7313 CSoutput.n219 CSoutput.n213 2.2505
R7314 CSoutput.n264 CSoutput.n213 2.2505
R7315 CSoutput.n264 CSoutput.n217 2.2505
R7316 CSoutput.n164 CSoutput.n144 2.2505
R7317 CSoutput.n159 CSoutput.n144 2.2505
R7318 CSoutput.n157 CSoutput.n144 2.2505
R7319 CSoutput.n156 CSoutput.n144 2.2505
R7320 CSoutput.n285 CSoutput.n144 2.2505
R7321 CSoutput.n283 CSoutput.n144 2.2505
R7322 CSoutput.n281 CSoutput.n144 2.2505
R7323 CSoutput.n167 CSoutput.n144 2.2505
R7324 CSoutput.n166 CSoutput.n144 2.2505
R7325 CSoutput.n170 CSoutput.n144 2.2505
R7326 CSoutput.n169 CSoutput.n144 2.2505
R7327 CSoutput.n152 CSoutput.n144 2.2505
R7328 CSoutput.n288 CSoutput.n144 2.2505
R7329 CSoutput.n288 CSoutput.n287 2.2505
R7330 CSoutput.n206 CSoutput.n199 2.25024
R7331 CSoutput.n206 CSoutput.n192 2.25024
R7332 CSoutput.n274 CSoutput.n206 2.25024
R7333 CSoutput.n206 CSoutput.n202 2.25024
R7334 CSoutput.n206 CSoutput.n205 2.25024
R7335 CSoutput.n206 CSoutput.n173 2.25024
R7336 CSoutput.n256 CSoutput.n253 2.25024
R7337 CSoutput.n256 CSoutput.n252 2.25024
R7338 CSoutput.n256 CSoutput.n251 2.25024
R7339 CSoutput.n256 CSoutput.n218 2.25024
R7340 CSoutput.n256 CSoutput.n255 2.25024
R7341 CSoutput.n257 CSoutput.n256 2.25024
R7342 CSoutput.n172 CSoutput.n165 2.25024
R7343 CSoutput.n172 CSoutput.n158 2.25024
R7344 CSoutput.n284 CSoutput.n172 2.25024
R7345 CSoutput.n172 CSoutput.n168 2.25024
R7346 CSoutput.n172 CSoutput.n171 2.25024
R7347 CSoutput.n172 CSoutput.n139 2.25024
R7348 CSoutput.n273 CSoutput.n183 1.50111
R7349 CSoutput.n221 CSoutput.n207 1.50111
R7350 CSoutput.n283 CSoutput.n149 1.50111
R7351 CSoutput.n229 CSoutput.n228 1.501
R7352 CSoutput.n236 CSoutput.n235 1.501
R7353 CSoutput.n263 CSoutput.n262 1.501
R7354 CSoutput.n277 CSoutput.n188 1.12536
R7355 CSoutput.n277 CSoutput.n189 1.12536
R7356 CSoutput.n277 CSoutput.n276 1.12536
R7357 CSoutput.n237 CSoutput.n217 1.12536
R7358 CSoutput.n243 CSoutput.n217 1.12536
R7359 CSoutput.n245 CSoutput.n217 1.12536
R7360 CSoutput.n287 CSoutput.n154 1.12536
R7361 CSoutput.n287 CSoutput.n155 1.12536
R7362 CSoutput.n287 CSoutput.n286 1.12536
R7363 CSoutput.n277 CSoutput.n184 1.12536
R7364 CSoutput.n277 CSoutput.n185 1.12536
R7365 CSoutput.n277 CSoutput.n187 1.12536
R7366 CSoutput.n267 CSoutput.n217 1.12536
R7367 CSoutput.n247 CSoutput.n217 1.12536
R7368 CSoutput.n249 CSoutput.n217 1.12536
R7369 CSoutput.n287 CSoutput.n150 1.12536
R7370 CSoutput.n287 CSoutput.n151 1.12536
R7371 CSoutput.n287 CSoutput.n153 1.12536
R7372 CSoutput.n31 CSoutput.n30 0.669944
R7373 CSoutput.n62 CSoutput.n61 0.669944
R7374 CSoutput.n384 CSoutput.n382 0.573776
R7375 CSoutput.n386 CSoutput.n384 0.573776
R7376 CSoutput.n388 CSoutput.n386 0.573776
R7377 CSoutput.n390 CSoutput.n388 0.573776
R7378 CSoutput.n392 CSoutput.n390 0.573776
R7379 CSoutput.n394 CSoutput.n392 0.573776
R7380 CSoutput.n368 CSoutput.n366 0.573776
R7381 CSoutput.n370 CSoutput.n368 0.573776
R7382 CSoutput.n372 CSoutput.n370 0.573776
R7383 CSoutput.n374 CSoutput.n372 0.573776
R7384 CSoutput.n376 CSoutput.n374 0.573776
R7385 CSoutput.n378 CSoutput.n376 0.573776
R7386 CSoutput.n353 CSoutput.n351 0.573776
R7387 CSoutput.n355 CSoutput.n353 0.573776
R7388 CSoutput.n357 CSoutput.n355 0.573776
R7389 CSoutput.n359 CSoutput.n357 0.573776
R7390 CSoutput.n361 CSoutput.n359 0.573776
R7391 CSoutput.n363 CSoutput.n361 0.573776
R7392 CSoutput.n442 CSoutput.n440 0.573776
R7393 CSoutput.n440 CSoutput.n438 0.573776
R7394 CSoutput.n438 CSoutput.n436 0.573776
R7395 CSoutput.n436 CSoutput.n434 0.573776
R7396 CSoutput.n434 CSoutput.n432 0.573776
R7397 CSoutput.n432 CSoutput.n430 0.573776
R7398 CSoutput.n426 CSoutput.n424 0.573776
R7399 CSoutput.n424 CSoutput.n422 0.573776
R7400 CSoutput.n422 CSoutput.n420 0.573776
R7401 CSoutput.n420 CSoutput.n418 0.573776
R7402 CSoutput.n418 CSoutput.n416 0.573776
R7403 CSoutput.n416 CSoutput.n414 0.573776
R7404 CSoutput.n411 CSoutput.n409 0.573776
R7405 CSoutput.n409 CSoutput.n407 0.573776
R7406 CSoutput.n407 CSoutput.n405 0.573776
R7407 CSoutput.n405 CSoutput.n403 0.573776
R7408 CSoutput.n403 CSoutput.n401 0.573776
R7409 CSoutput.n401 CSoutput.n399 0.573776
R7410 CSoutput.n445 CSoutput.n288 0.53442
R7411 CSoutput.n332 CSoutput.n330 0.358259
R7412 CSoutput.n334 CSoutput.n332 0.358259
R7413 CSoutput.n336 CSoutput.n334 0.358259
R7414 CSoutput.n338 CSoutput.n336 0.358259
R7415 CSoutput.n340 CSoutput.n338 0.358259
R7416 CSoutput.n342 CSoutput.n340 0.358259
R7417 CSoutput.n344 CSoutput.n342 0.358259
R7418 CSoutput.n346 CSoutput.n344 0.358259
R7419 CSoutput.n312 CSoutput.n310 0.358259
R7420 CSoutput.n314 CSoutput.n312 0.358259
R7421 CSoutput.n316 CSoutput.n314 0.358259
R7422 CSoutput.n318 CSoutput.n316 0.358259
R7423 CSoutput.n320 CSoutput.n318 0.358259
R7424 CSoutput.n322 CSoutput.n320 0.358259
R7425 CSoutput.n324 CSoutput.n322 0.358259
R7426 CSoutput.n326 CSoutput.n324 0.358259
R7427 CSoutput.n293 CSoutput.n291 0.358259
R7428 CSoutput.n295 CSoutput.n293 0.358259
R7429 CSoutput.n297 CSoutput.n295 0.358259
R7430 CSoutput.n299 CSoutput.n297 0.358259
R7431 CSoutput.n301 CSoutput.n299 0.358259
R7432 CSoutput.n303 CSoutput.n301 0.358259
R7433 CSoutput.n305 CSoutput.n303 0.358259
R7434 CSoutput.n307 CSoutput.n305 0.358259
R7435 CSoutput.n136 CSoutput.n134 0.358259
R7436 CSoutput.n134 CSoutput.n132 0.358259
R7437 CSoutput.n132 CSoutput.n130 0.358259
R7438 CSoutput.n130 CSoutput.n128 0.358259
R7439 CSoutput.n128 CSoutput.n126 0.358259
R7440 CSoutput.n126 CSoutput.n124 0.358259
R7441 CSoutput.n124 CSoutput.n122 0.358259
R7442 CSoutput.n122 CSoutput.n120 0.358259
R7443 CSoutput.n116 CSoutput.n114 0.358259
R7444 CSoutput.n114 CSoutput.n112 0.358259
R7445 CSoutput.n112 CSoutput.n110 0.358259
R7446 CSoutput.n110 CSoutput.n108 0.358259
R7447 CSoutput.n108 CSoutput.n106 0.358259
R7448 CSoutput.n106 CSoutput.n104 0.358259
R7449 CSoutput.n104 CSoutput.n102 0.358259
R7450 CSoutput.n102 CSoutput.n100 0.358259
R7451 CSoutput.n97 CSoutput.n95 0.358259
R7452 CSoutput.n95 CSoutput.n93 0.358259
R7453 CSoutput.n93 CSoutput.n91 0.358259
R7454 CSoutput.n91 CSoutput.n89 0.358259
R7455 CSoutput.n89 CSoutput.n87 0.358259
R7456 CSoutput.n87 CSoutput.n85 0.358259
R7457 CSoutput.n85 CSoutput.n83 0.358259
R7458 CSoutput.n83 CSoutput.n81 0.358259
R7459 CSoutput.n21 CSoutput.n20 0.169105
R7460 CSoutput.n21 CSoutput.n16 0.169105
R7461 CSoutput.n26 CSoutput.n16 0.169105
R7462 CSoutput.n27 CSoutput.n26 0.169105
R7463 CSoutput.n27 CSoutput.n14 0.169105
R7464 CSoutput.n32 CSoutput.n14 0.169105
R7465 CSoutput.n33 CSoutput.n32 0.169105
R7466 CSoutput.n34 CSoutput.n33 0.169105
R7467 CSoutput.n34 CSoutput.n12 0.169105
R7468 CSoutput.n39 CSoutput.n12 0.169105
R7469 CSoutput.n40 CSoutput.n39 0.169105
R7470 CSoutput.n40 CSoutput.n10 0.169105
R7471 CSoutput.n45 CSoutput.n10 0.169105
R7472 CSoutput.n46 CSoutput.n45 0.169105
R7473 CSoutput.n47 CSoutput.n46 0.169105
R7474 CSoutput.n47 CSoutput.n8 0.169105
R7475 CSoutput.n52 CSoutput.n8 0.169105
R7476 CSoutput.n53 CSoutput.n52 0.169105
R7477 CSoutput.n53 CSoutput.n6 0.169105
R7478 CSoutput.n58 CSoutput.n6 0.169105
R7479 CSoutput.n59 CSoutput.n58 0.169105
R7480 CSoutput.n60 CSoutput.n59 0.169105
R7481 CSoutput.n60 CSoutput.n4 0.169105
R7482 CSoutput.n66 CSoutput.n4 0.169105
R7483 CSoutput.n67 CSoutput.n66 0.169105
R7484 CSoutput.n68 CSoutput.n67 0.169105
R7485 CSoutput.n68 CSoutput.n2 0.169105
R7486 CSoutput.n73 CSoutput.n2 0.169105
R7487 CSoutput.n74 CSoutput.n73 0.169105
R7488 CSoutput.n74 CSoutput.n0 0.169105
R7489 CSoutput.n78 CSoutput.n0 0.169105
R7490 CSoutput.n231 CSoutput.n230 0.0910737
R7491 CSoutput.n282 CSoutput.n279 0.0723685
R7492 CSoutput.n236 CSoutput.n231 0.0522944
R7493 CSoutput.n279 CSoutput.n278 0.0499135
R7494 CSoutput.n230 CSoutput.n229 0.0499135
R7495 CSoutput.n264 CSoutput.n263 0.0464294
R7496 CSoutput.n272 CSoutput.n269 0.0391444
R7497 CSoutput.n231 CSoutput.t236 0.023435
R7498 CSoutput.n279 CSoutput.t228 0.02262
R7499 CSoutput.n230 CSoutput.t217 0.02262
R7500 CSoutput CSoutput.n445 0.0052
R7501 CSoutput.n201 CSoutput.n184 0.00365111
R7502 CSoutput.n204 CSoutput.n185 0.00365111
R7503 CSoutput.n187 CSoutput.n186 0.00365111
R7504 CSoutput.n229 CSoutput.n188 0.00365111
R7505 CSoutput.n193 CSoutput.n189 0.00365111
R7506 CSoutput.n276 CSoutput.n190 0.00365111
R7507 CSoutput.n267 CSoutput.n266 0.00365111
R7508 CSoutput.n247 CSoutput.n220 0.00365111
R7509 CSoutput.n249 CSoutput.n219 0.00365111
R7510 CSoutput.n237 CSoutput.n236 0.00365111
R7511 CSoutput.n243 CSoutput.n223 0.00365111
R7512 CSoutput.n245 CSoutput.n222 0.00365111
R7513 CSoutput.n167 CSoutput.n150 0.00365111
R7514 CSoutput.n170 CSoutput.n151 0.00365111
R7515 CSoutput.n153 CSoutput.n152 0.00365111
R7516 CSoutput.n263 CSoutput.n154 0.00365111
R7517 CSoutput.n159 CSoutput.n155 0.00365111
R7518 CSoutput.n286 CSoutput.n156 0.00365111
R7519 CSoutput.n198 CSoutput.n188 0.00340054
R7520 CSoutput.n191 CSoutput.n189 0.00340054
R7521 CSoutput.n276 CSoutput.n275 0.00340054
R7522 CSoutput.n271 CSoutput.n184 0.00340054
R7523 CSoutput.n200 CSoutput.n185 0.00340054
R7524 CSoutput.n203 CSoutput.n187 0.00340054
R7525 CSoutput.n242 CSoutput.n237 0.00340054
R7526 CSoutput.n244 CSoutput.n243 0.00340054
R7527 CSoutput.n246 CSoutput.n245 0.00340054
R7528 CSoutput.n268 CSoutput.n267 0.00340054
R7529 CSoutput.n248 CSoutput.n247 0.00340054
R7530 CSoutput.n250 CSoutput.n249 0.00340054
R7531 CSoutput.n164 CSoutput.n154 0.00340054
R7532 CSoutput.n157 CSoutput.n155 0.00340054
R7533 CSoutput.n286 CSoutput.n285 0.00340054
R7534 CSoutput.n281 CSoutput.n150 0.00340054
R7535 CSoutput.n166 CSoutput.n151 0.00340054
R7536 CSoutput.n169 CSoutput.n153 0.00340054
R7537 CSoutput.n199 CSoutput.n193 0.00252698
R7538 CSoutput.n192 CSoutput.n190 0.00252698
R7539 CSoutput.n274 CSoutput.n273 0.00252698
R7540 CSoutput.n202 CSoutput.n200 0.00252698
R7541 CSoutput.n205 CSoutput.n203 0.00252698
R7542 CSoutput.n278 CSoutput.n173 0.00252698
R7543 CSoutput.n199 CSoutput.n198 0.00252698
R7544 CSoutput.n192 CSoutput.n191 0.00252698
R7545 CSoutput.n275 CSoutput.n274 0.00252698
R7546 CSoutput.n202 CSoutput.n201 0.00252698
R7547 CSoutput.n205 CSoutput.n204 0.00252698
R7548 CSoutput.n186 CSoutput.n173 0.00252698
R7549 CSoutput.n253 CSoutput.n223 0.00252698
R7550 CSoutput.n252 CSoutput.n222 0.00252698
R7551 CSoutput.n251 CSoutput.n207 0.00252698
R7552 CSoutput.n248 CSoutput.n218 0.00252698
R7553 CSoutput.n255 CSoutput.n250 0.00252698
R7554 CSoutput.n264 CSoutput.n257 0.00252698
R7555 CSoutput.n253 CSoutput.n242 0.00252698
R7556 CSoutput.n252 CSoutput.n244 0.00252698
R7557 CSoutput.n251 CSoutput.n246 0.00252698
R7558 CSoutput.n266 CSoutput.n218 0.00252698
R7559 CSoutput.n255 CSoutput.n220 0.00252698
R7560 CSoutput.n257 CSoutput.n219 0.00252698
R7561 CSoutput.n165 CSoutput.n159 0.00252698
R7562 CSoutput.n158 CSoutput.n156 0.00252698
R7563 CSoutput.n284 CSoutput.n283 0.00252698
R7564 CSoutput.n168 CSoutput.n166 0.00252698
R7565 CSoutput.n171 CSoutput.n169 0.00252698
R7566 CSoutput.n288 CSoutput.n139 0.00252698
R7567 CSoutput.n165 CSoutput.n164 0.00252698
R7568 CSoutput.n158 CSoutput.n157 0.00252698
R7569 CSoutput.n285 CSoutput.n284 0.00252698
R7570 CSoutput.n168 CSoutput.n167 0.00252698
R7571 CSoutput.n171 CSoutput.n170 0.00252698
R7572 CSoutput.n152 CSoutput.n139 0.00252698
R7573 CSoutput.n273 CSoutput.n272 0.0020275
R7574 CSoutput.n272 CSoutput.n271 0.0020275
R7575 CSoutput.n269 CSoutput.n207 0.0020275
R7576 CSoutput.n269 CSoutput.n268 0.0020275
R7577 CSoutput.n283 CSoutput.n282 0.0020275
R7578 CSoutput.n282 CSoutput.n281 0.0020275
R7579 CSoutput.n183 CSoutput.n182 0.00166668
R7580 CSoutput.n265 CSoutput.n221 0.00166668
R7581 CSoutput.n149 CSoutput.n148 0.00166668
R7582 CSoutput.n287 CSoutput.n149 0.00133328
R7583 CSoutput.n221 CSoutput.n217 0.00133328
R7584 CSoutput.n277 CSoutput.n183 0.00133328
R7585 CSoutput.n280 CSoutput.n172 0.001
R7586 CSoutput.n258 CSoutput.n172 0.001
R7587 CSoutput.n160 CSoutput.n140 0.001
R7588 CSoutput.n259 CSoutput.n140 0.001
R7589 CSoutput.n161 CSoutput.n141 0.001
R7590 CSoutput.n260 CSoutput.n141 0.001
R7591 CSoutput.n162 CSoutput.n142 0.001
R7592 CSoutput.n261 CSoutput.n142 0.001
R7593 CSoutput.n163 CSoutput.n143 0.001
R7594 CSoutput.n262 CSoutput.n143 0.001
R7595 CSoutput.n256 CSoutput.n208 0.001
R7596 CSoutput.n256 CSoutput.n254 0.001
R7597 CSoutput.n238 CSoutput.n209 0.001
R7598 CSoutput.n232 CSoutput.n209 0.001
R7599 CSoutput.n239 CSoutput.n210 0.001
R7600 CSoutput.n233 CSoutput.n210 0.001
R7601 CSoutput.n240 CSoutput.n211 0.001
R7602 CSoutput.n234 CSoutput.n211 0.001
R7603 CSoutput.n241 CSoutput.n212 0.001
R7604 CSoutput.n235 CSoutput.n212 0.001
R7605 CSoutput.n270 CSoutput.n206 0.001
R7606 CSoutput.n224 CSoutput.n206 0.001
R7607 CSoutput.n194 CSoutput.n174 0.001
R7608 CSoutput.n225 CSoutput.n174 0.001
R7609 CSoutput.n195 CSoutput.n175 0.001
R7610 CSoutput.n226 CSoutput.n175 0.001
R7611 CSoutput.n196 CSoutput.n176 0.001
R7612 CSoutput.n227 CSoutput.n176 0.001
R7613 CSoutput.n197 CSoutput.n177 0.001
R7614 CSoutput.n228 CSoutput.n177 0.001
R7615 CSoutput.n228 CSoutput.n178 0.001
R7616 CSoutput.n227 CSoutput.n179 0.001
R7617 CSoutput.n226 CSoutput.n180 0.001
R7618 CSoutput.n225 CSoutput.t233 0.001
R7619 CSoutput.n224 CSoutput.n181 0.001
R7620 CSoutput.n197 CSoutput.n179 0.001
R7621 CSoutput.n196 CSoutput.n180 0.001
R7622 CSoutput.n195 CSoutput.t233 0.001
R7623 CSoutput.n194 CSoutput.n181 0.001
R7624 CSoutput.n270 CSoutput.n182 0.001
R7625 CSoutput.n235 CSoutput.n213 0.001
R7626 CSoutput.n234 CSoutput.n214 0.001
R7627 CSoutput.n233 CSoutput.n215 0.001
R7628 CSoutput.n232 CSoutput.t226 0.001
R7629 CSoutput.n254 CSoutput.n216 0.001
R7630 CSoutput.n241 CSoutput.n214 0.001
R7631 CSoutput.n240 CSoutput.n215 0.001
R7632 CSoutput.n239 CSoutput.t226 0.001
R7633 CSoutput.n238 CSoutput.n216 0.001
R7634 CSoutput.n265 CSoutput.n208 0.001
R7635 CSoutput.n262 CSoutput.n144 0.001
R7636 CSoutput.n261 CSoutput.n145 0.001
R7637 CSoutput.n260 CSoutput.n146 0.001
R7638 CSoutput.n259 CSoutput.t216 0.001
R7639 CSoutput.n258 CSoutput.n147 0.001
R7640 CSoutput.n163 CSoutput.n145 0.001
R7641 CSoutput.n162 CSoutput.n146 0.001
R7642 CSoutput.n161 CSoutput.t216 0.001
R7643 CSoutput.n160 CSoutput.n147 0.001
R7644 CSoutput.n280 CSoutput.n148 0.001
R7645 commonsourceibias.n35 commonsourceibias.t54 223.028
R7646 commonsourceibias.n128 commonsourceibias.t132 223.028
R7647 commonsourceibias.n307 commonsourceibias.t136 223.028
R7648 commonsourceibias.n217 commonsourceibias.t64 223.028
R7649 commonsourceibias.n454 commonsourceibias.t50 223.028
R7650 commonsourceibias.n395 commonsourceibias.t83 223.028
R7651 commonsourceibias.n679 commonsourceibias.t144 223.028
R7652 commonsourceibias.n589 commonsourceibias.t131 223.028
R7653 commonsourceibias.n99 commonsourceibias.t58 207.983
R7654 commonsourceibias.n192 commonsourceibias.t78 207.983
R7655 commonsourceibias.n371 commonsourceibias.t148 207.983
R7656 commonsourceibias.n281 commonsourceibias.t115 207.983
R7657 commonsourceibias.n520 commonsourceibias.t40 207.983
R7658 commonsourceibias.n566 commonsourceibias.t153 207.983
R7659 commonsourceibias.n745 commonsourceibias.t71 207.983
R7660 commonsourceibias.n655 commonsourceibias.t100 207.983
R7661 commonsourceibias.n97 commonsourceibias.t52 168.701
R7662 commonsourceibias.n91 commonsourceibias.t4 168.701
R7663 commonsourceibias.n17 commonsourceibias.t44 168.701
R7664 commonsourceibias.n83 commonsourceibias.t18 168.701
R7665 commonsourceibias.n77 commonsourceibias.t16 168.701
R7666 commonsourceibias.n22 commonsourceibias.t8 168.701
R7667 commonsourceibias.n69 commonsourceibias.t14 168.701
R7668 commonsourceibias.n63 commonsourceibias.t46 168.701
R7669 commonsourceibias.n25 commonsourceibias.t22 168.701
R7670 commonsourceibias.n27 commonsourceibias.t2 168.701
R7671 commonsourceibias.n29 commonsourceibias.t28 168.701
R7672 commonsourceibias.n46 commonsourceibias.t20 168.701
R7673 commonsourceibias.n40 commonsourceibias.t56 168.701
R7674 commonsourceibias.n34 commonsourceibias.t30 168.701
R7675 commonsourceibias.n190 commonsourceibias.t146 168.701
R7676 commonsourceibias.n184 commonsourceibias.t96 168.701
R7677 commonsourceibias.n5 commonsourceibias.t157 168.701
R7678 commonsourceibias.n176 commonsourceibias.t112 168.701
R7679 commonsourceibias.n170 commonsourceibias.t75 168.701
R7680 commonsourceibias.n10 commonsourceibias.t124 168.701
R7681 commonsourceibias.n162 commonsourceibias.t113 168.701
R7682 commonsourceibias.n156 commonsourceibias.t154 168.701
R7683 commonsourceibias.n118 commonsourceibias.t106 168.701
R7684 commonsourceibias.n120 commonsourceibias.t92 168.701
R7685 commonsourceibias.n122 commonsourceibias.t123 168.701
R7686 commonsourceibias.n139 commonsourceibias.t110 168.701
R7687 commonsourceibias.n133 commonsourceibias.t82 168.701
R7688 commonsourceibias.n127 commonsourceibias.t147 168.701
R7689 commonsourceibias.n306 commonsourceibias.t143 168.701
R7690 commonsourceibias.n312 commonsourceibias.t70 168.701
R7691 commonsourceibias.n318 commonsourceibias.t150 168.701
R7692 commonsourceibias.n301 commonsourceibias.t158 168.701
R7693 commonsourceibias.n299 commonsourceibias.t101 168.701
R7694 commonsourceibias.n297 commonsourceibias.t81 168.701
R7695 commonsourceibias.n335 commonsourceibias.t67 168.701
R7696 commonsourceibias.n341 commonsourceibias.t111 168.701
R7697 commonsourceibias.n294 commonsourceibias.t120 168.701
R7698 commonsourceibias.n349 commonsourceibias.t74 168.701
R7699 commonsourceibias.n355 commonsourceibias.t159 168.701
R7700 commonsourceibias.n289 commonsourceibias.t134 168.701
R7701 commonsourceibias.n363 commonsourceibias.t80 168.701
R7702 commonsourceibias.n369 commonsourceibias.t68 168.701
R7703 commonsourceibias.n279 commonsourceibias.t138 168.701
R7704 commonsourceibias.n273 commonsourceibias.t128 168.701
R7705 commonsourceibias.n199 commonsourceibias.t116 168.701
R7706 commonsourceibias.n265 commonsourceibias.t139 168.701
R7707 commonsourceibias.n259 commonsourceibias.t126 168.701
R7708 commonsourceibias.n204 commonsourceibias.t114 168.701
R7709 commonsourceibias.n251 commonsourceibias.t140 168.701
R7710 commonsourceibias.n245 commonsourceibias.t127 168.701
R7711 commonsourceibias.n207 commonsourceibias.t149 168.701
R7712 commonsourceibias.n209 commonsourceibias.t141 168.701
R7713 commonsourceibias.n211 commonsourceibias.t125 168.701
R7714 commonsourceibias.n228 commonsourceibias.t152 168.701
R7715 commonsourceibias.n222 commonsourceibias.t69 168.701
R7716 commonsourceibias.n216 commonsourceibias.t135 168.701
R7717 commonsourceibias.n453 commonsourceibias.t48 168.701
R7718 commonsourceibias.n459 commonsourceibias.t42 168.701
R7719 commonsourceibias.n465 commonsourceibias.t36 168.701
R7720 commonsourceibias.n448 commonsourceibias.t0 168.701
R7721 commonsourceibias.n446 commonsourceibias.t60 168.701
R7722 commonsourceibias.n444 commonsourceibias.t38 168.701
R7723 commonsourceibias.n482 commonsourceibias.t12 168.701
R7724 commonsourceibias.n488 commonsourceibias.t62 168.701
R7725 commonsourceibias.n490 commonsourceibias.t6 168.701
R7726 commonsourceibias.n497 commonsourceibias.t26 168.701
R7727 commonsourceibias.n503 commonsourceibias.t34 168.701
R7728 commonsourceibias.n505 commonsourceibias.t10 168.701
R7729 commonsourceibias.n512 commonsourceibias.t32 168.701
R7730 commonsourceibias.n518 commonsourceibias.t24 168.701
R7731 commonsourceibias.n564 commonsourceibias.t104 168.701
R7732 commonsourceibias.n558 commonsourceibias.t73 168.701
R7733 commonsourceibias.n551 commonsourceibias.t121 168.701
R7734 commonsourceibias.n549 commonsourceibias.t90 168.701
R7735 commonsourceibias.n543 commonsourceibias.t151 168.701
R7736 commonsourceibias.n536 commonsourceibias.t102 168.701
R7737 commonsourceibias.n534 commonsourceibias.t91 168.701
R7738 commonsourceibias.n394 commonsourceibias.t84 168.701
R7739 commonsourceibias.n400 commonsourceibias.t65 168.701
R7740 commonsourceibias.n406 commonsourceibias.t88 168.701
R7741 commonsourceibias.n389 commonsourceibias.t95 168.701
R7742 commonsourceibias.n387 commonsourceibias.t79 168.701
R7743 commonsourceibias.n385 commonsourceibias.t87 168.701
R7744 commonsourceibias.n423 commonsourceibias.t119 168.701
R7745 commonsourceibias.n678 commonsourceibias.t133 168.701
R7746 commonsourceibias.n684 commonsourceibias.t89 168.701
R7747 commonsourceibias.n690 commonsourceibias.t72 168.701
R7748 commonsourceibias.n673 commonsourceibias.t76 168.701
R7749 commonsourceibias.n671 commonsourceibias.t94 168.701
R7750 commonsourceibias.n669 commonsourceibias.t98 168.701
R7751 commonsourceibias.n707 commonsourceibias.t85 168.701
R7752 commonsourceibias.n713 commonsourceibias.t145 168.701
R7753 commonsourceibias.n715 commonsourceibias.t103 168.701
R7754 commonsourceibias.n722 commonsourceibias.t93 168.701
R7755 commonsourceibias.n728 commonsourceibias.t77 168.701
R7756 commonsourceibias.n730 commonsourceibias.t66 168.701
R7757 commonsourceibias.n737 commonsourceibias.t97 168.701
R7758 commonsourceibias.n743 commonsourceibias.t86 168.701
R7759 commonsourceibias.n588 commonsourceibias.t142 168.701
R7760 commonsourceibias.n594 commonsourceibias.t155 168.701
R7761 commonsourceibias.n600 commonsourceibias.t137 168.701
R7762 commonsourceibias.n583 commonsourceibias.t105 168.701
R7763 commonsourceibias.n581 commonsourceibias.t156 168.701
R7764 commonsourceibias.n579 commonsourceibias.t129 168.701
R7765 commonsourceibias.n617 commonsourceibias.t107 168.701
R7766 commonsourceibias.n623 commonsourceibias.t122 168.701
R7767 commonsourceibias.n625 commonsourceibias.t130 168.701
R7768 commonsourceibias.n632 commonsourceibias.t108 168.701
R7769 commonsourceibias.n638 commonsourceibias.t117 168.701
R7770 commonsourceibias.n640 commonsourceibias.t99 168.701
R7771 commonsourceibias.n647 commonsourceibias.t109 168.701
R7772 commonsourceibias.n653 commonsourceibias.t118 168.701
R7773 commonsourceibias.n36 commonsourceibias.n33 161.3
R7774 commonsourceibias.n38 commonsourceibias.n37 161.3
R7775 commonsourceibias.n39 commonsourceibias.n32 161.3
R7776 commonsourceibias.n42 commonsourceibias.n41 161.3
R7777 commonsourceibias.n43 commonsourceibias.n31 161.3
R7778 commonsourceibias.n45 commonsourceibias.n44 161.3
R7779 commonsourceibias.n47 commonsourceibias.n30 161.3
R7780 commonsourceibias.n49 commonsourceibias.n48 161.3
R7781 commonsourceibias.n51 commonsourceibias.n50 161.3
R7782 commonsourceibias.n52 commonsourceibias.n28 161.3
R7783 commonsourceibias.n54 commonsourceibias.n53 161.3
R7784 commonsourceibias.n56 commonsourceibias.n55 161.3
R7785 commonsourceibias.n57 commonsourceibias.n26 161.3
R7786 commonsourceibias.n59 commonsourceibias.n58 161.3
R7787 commonsourceibias.n61 commonsourceibias.n60 161.3
R7788 commonsourceibias.n62 commonsourceibias.n24 161.3
R7789 commonsourceibias.n65 commonsourceibias.n64 161.3
R7790 commonsourceibias.n66 commonsourceibias.n23 161.3
R7791 commonsourceibias.n68 commonsourceibias.n67 161.3
R7792 commonsourceibias.n70 commonsourceibias.n21 161.3
R7793 commonsourceibias.n72 commonsourceibias.n71 161.3
R7794 commonsourceibias.n73 commonsourceibias.n20 161.3
R7795 commonsourceibias.n75 commonsourceibias.n74 161.3
R7796 commonsourceibias.n76 commonsourceibias.n19 161.3
R7797 commonsourceibias.n79 commonsourceibias.n78 161.3
R7798 commonsourceibias.n80 commonsourceibias.n18 161.3
R7799 commonsourceibias.n82 commonsourceibias.n81 161.3
R7800 commonsourceibias.n84 commonsourceibias.n16 161.3
R7801 commonsourceibias.n86 commonsourceibias.n85 161.3
R7802 commonsourceibias.n87 commonsourceibias.n15 161.3
R7803 commonsourceibias.n89 commonsourceibias.n88 161.3
R7804 commonsourceibias.n90 commonsourceibias.n14 161.3
R7805 commonsourceibias.n93 commonsourceibias.n92 161.3
R7806 commonsourceibias.n94 commonsourceibias.n13 161.3
R7807 commonsourceibias.n96 commonsourceibias.n95 161.3
R7808 commonsourceibias.n98 commonsourceibias.n12 161.3
R7809 commonsourceibias.n129 commonsourceibias.n126 161.3
R7810 commonsourceibias.n131 commonsourceibias.n130 161.3
R7811 commonsourceibias.n132 commonsourceibias.n125 161.3
R7812 commonsourceibias.n135 commonsourceibias.n134 161.3
R7813 commonsourceibias.n136 commonsourceibias.n124 161.3
R7814 commonsourceibias.n138 commonsourceibias.n137 161.3
R7815 commonsourceibias.n140 commonsourceibias.n123 161.3
R7816 commonsourceibias.n142 commonsourceibias.n141 161.3
R7817 commonsourceibias.n144 commonsourceibias.n143 161.3
R7818 commonsourceibias.n145 commonsourceibias.n121 161.3
R7819 commonsourceibias.n147 commonsourceibias.n146 161.3
R7820 commonsourceibias.n149 commonsourceibias.n148 161.3
R7821 commonsourceibias.n150 commonsourceibias.n119 161.3
R7822 commonsourceibias.n152 commonsourceibias.n151 161.3
R7823 commonsourceibias.n154 commonsourceibias.n153 161.3
R7824 commonsourceibias.n155 commonsourceibias.n117 161.3
R7825 commonsourceibias.n158 commonsourceibias.n157 161.3
R7826 commonsourceibias.n159 commonsourceibias.n11 161.3
R7827 commonsourceibias.n161 commonsourceibias.n160 161.3
R7828 commonsourceibias.n163 commonsourceibias.n9 161.3
R7829 commonsourceibias.n165 commonsourceibias.n164 161.3
R7830 commonsourceibias.n166 commonsourceibias.n8 161.3
R7831 commonsourceibias.n168 commonsourceibias.n167 161.3
R7832 commonsourceibias.n169 commonsourceibias.n7 161.3
R7833 commonsourceibias.n172 commonsourceibias.n171 161.3
R7834 commonsourceibias.n173 commonsourceibias.n6 161.3
R7835 commonsourceibias.n175 commonsourceibias.n174 161.3
R7836 commonsourceibias.n177 commonsourceibias.n4 161.3
R7837 commonsourceibias.n179 commonsourceibias.n178 161.3
R7838 commonsourceibias.n180 commonsourceibias.n3 161.3
R7839 commonsourceibias.n182 commonsourceibias.n181 161.3
R7840 commonsourceibias.n183 commonsourceibias.n2 161.3
R7841 commonsourceibias.n186 commonsourceibias.n185 161.3
R7842 commonsourceibias.n187 commonsourceibias.n1 161.3
R7843 commonsourceibias.n189 commonsourceibias.n188 161.3
R7844 commonsourceibias.n191 commonsourceibias.n0 161.3
R7845 commonsourceibias.n370 commonsourceibias.n284 161.3
R7846 commonsourceibias.n368 commonsourceibias.n367 161.3
R7847 commonsourceibias.n366 commonsourceibias.n285 161.3
R7848 commonsourceibias.n365 commonsourceibias.n364 161.3
R7849 commonsourceibias.n362 commonsourceibias.n286 161.3
R7850 commonsourceibias.n361 commonsourceibias.n360 161.3
R7851 commonsourceibias.n359 commonsourceibias.n287 161.3
R7852 commonsourceibias.n358 commonsourceibias.n357 161.3
R7853 commonsourceibias.n356 commonsourceibias.n288 161.3
R7854 commonsourceibias.n354 commonsourceibias.n353 161.3
R7855 commonsourceibias.n352 commonsourceibias.n290 161.3
R7856 commonsourceibias.n351 commonsourceibias.n350 161.3
R7857 commonsourceibias.n348 commonsourceibias.n291 161.3
R7858 commonsourceibias.n347 commonsourceibias.n346 161.3
R7859 commonsourceibias.n345 commonsourceibias.n292 161.3
R7860 commonsourceibias.n344 commonsourceibias.n343 161.3
R7861 commonsourceibias.n342 commonsourceibias.n293 161.3
R7862 commonsourceibias.n340 commonsourceibias.n339 161.3
R7863 commonsourceibias.n338 commonsourceibias.n295 161.3
R7864 commonsourceibias.n337 commonsourceibias.n336 161.3
R7865 commonsourceibias.n334 commonsourceibias.n296 161.3
R7866 commonsourceibias.n333 commonsourceibias.n332 161.3
R7867 commonsourceibias.n331 commonsourceibias.n330 161.3
R7868 commonsourceibias.n329 commonsourceibias.n298 161.3
R7869 commonsourceibias.n328 commonsourceibias.n327 161.3
R7870 commonsourceibias.n326 commonsourceibias.n325 161.3
R7871 commonsourceibias.n324 commonsourceibias.n300 161.3
R7872 commonsourceibias.n323 commonsourceibias.n322 161.3
R7873 commonsourceibias.n321 commonsourceibias.n320 161.3
R7874 commonsourceibias.n319 commonsourceibias.n302 161.3
R7875 commonsourceibias.n317 commonsourceibias.n316 161.3
R7876 commonsourceibias.n315 commonsourceibias.n303 161.3
R7877 commonsourceibias.n314 commonsourceibias.n313 161.3
R7878 commonsourceibias.n311 commonsourceibias.n304 161.3
R7879 commonsourceibias.n310 commonsourceibias.n309 161.3
R7880 commonsourceibias.n308 commonsourceibias.n305 161.3
R7881 commonsourceibias.n218 commonsourceibias.n215 161.3
R7882 commonsourceibias.n220 commonsourceibias.n219 161.3
R7883 commonsourceibias.n221 commonsourceibias.n214 161.3
R7884 commonsourceibias.n224 commonsourceibias.n223 161.3
R7885 commonsourceibias.n225 commonsourceibias.n213 161.3
R7886 commonsourceibias.n227 commonsourceibias.n226 161.3
R7887 commonsourceibias.n229 commonsourceibias.n212 161.3
R7888 commonsourceibias.n231 commonsourceibias.n230 161.3
R7889 commonsourceibias.n233 commonsourceibias.n232 161.3
R7890 commonsourceibias.n234 commonsourceibias.n210 161.3
R7891 commonsourceibias.n236 commonsourceibias.n235 161.3
R7892 commonsourceibias.n238 commonsourceibias.n237 161.3
R7893 commonsourceibias.n239 commonsourceibias.n208 161.3
R7894 commonsourceibias.n241 commonsourceibias.n240 161.3
R7895 commonsourceibias.n243 commonsourceibias.n242 161.3
R7896 commonsourceibias.n244 commonsourceibias.n206 161.3
R7897 commonsourceibias.n247 commonsourceibias.n246 161.3
R7898 commonsourceibias.n248 commonsourceibias.n205 161.3
R7899 commonsourceibias.n250 commonsourceibias.n249 161.3
R7900 commonsourceibias.n252 commonsourceibias.n203 161.3
R7901 commonsourceibias.n254 commonsourceibias.n253 161.3
R7902 commonsourceibias.n255 commonsourceibias.n202 161.3
R7903 commonsourceibias.n257 commonsourceibias.n256 161.3
R7904 commonsourceibias.n258 commonsourceibias.n201 161.3
R7905 commonsourceibias.n261 commonsourceibias.n260 161.3
R7906 commonsourceibias.n262 commonsourceibias.n200 161.3
R7907 commonsourceibias.n264 commonsourceibias.n263 161.3
R7908 commonsourceibias.n266 commonsourceibias.n198 161.3
R7909 commonsourceibias.n268 commonsourceibias.n267 161.3
R7910 commonsourceibias.n269 commonsourceibias.n197 161.3
R7911 commonsourceibias.n271 commonsourceibias.n270 161.3
R7912 commonsourceibias.n272 commonsourceibias.n196 161.3
R7913 commonsourceibias.n275 commonsourceibias.n274 161.3
R7914 commonsourceibias.n276 commonsourceibias.n195 161.3
R7915 commonsourceibias.n278 commonsourceibias.n277 161.3
R7916 commonsourceibias.n280 commonsourceibias.n194 161.3
R7917 commonsourceibias.n519 commonsourceibias.n433 161.3
R7918 commonsourceibias.n517 commonsourceibias.n516 161.3
R7919 commonsourceibias.n515 commonsourceibias.n434 161.3
R7920 commonsourceibias.n514 commonsourceibias.n513 161.3
R7921 commonsourceibias.n511 commonsourceibias.n435 161.3
R7922 commonsourceibias.n510 commonsourceibias.n509 161.3
R7923 commonsourceibias.n508 commonsourceibias.n436 161.3
R7924 commonsourceibias.n507 commonsourceibias.n506 161.3
R7925 commonsourceibias.n504 commonsourceibias.n437 161.3
R7926 commonsourceibias.n502 commonsourceibias.n501 161.3
R7927 commonsourceibias.n500 commonsourceibias.n438 161.3
R7928 commonsourceibias.n499 commonsourceibias.n498 161.3
R7929 commonsourceibias.n496 commonsourceibias.n439 161.3
R7930 commonsourceibias.n495 commonsourceibias.n494 161.3
R7931 commonsourceibias.n493 commonsourceibias.n440 161.3
R7932 commonsourceibias.n492 commonsourceibias.n491 161.3
R7933 commonsourceibias.n489 commonsourceibias.n441 161.3
R7934 commonsourceibias.n487 commonsourceibias.n486 161.3
R7935 commonsourceibias.n485 commonsourceibias.n442 161.3
R7936 commonsourceibias.n484 commonsourceibias.n483 161.3
R7937 commonsourceibias.n481 commonsourceibias.n443 161.3
R7938 commonsourceibias.n480 commonsourceibias.n479 161.3
R7939 commonsourceibias.n478 commonsourceibias.n477 161.3
R7940 commonsourceibias.n476 commonsourceibias.n445 161.3
R7941 commonsourceibias.n475 commonsourceibias.n474 161.3
R7942 commonsourceibias.n473 commonsourceibias.n472 161.3
R7943 commonsourceibias.n471 commonsourceibias.n447 161.3
R7944 commonsourceibias.n470 commonsourceibias.n469 161.3
R7945 commonsourceibias.n468 commonsourceibias.n467 161.3
R7946 commonsourceibias.n466 commonsourceibias.n449 161.3
R7947 commonsourceibias.n464 commonsourceibias.n463 161.3
R7948 commonsourceibias.n462 commonsourceibias.n450 161.3
R7949 commonsourceibias.n461 commonsourceibias.n460 161.3
R7950 commonsourceibias.n458 commonsourceibias.n451 161.3
R7951 commonsourceibias.n457 commonsourceibias.n456 161.3
R7952 commonsourceibias.n455 commonsourceibias.n452 161.3
R7953 commonsourceibias.n425 commonsourceibias.n424 161.3
R7954 commonsourceibias.n422 commonsourceibias.n384 161.3
R7955 commonsourceibias.n421 commonsourceibias.n420 161.3
R7956 commonsourceibias.n419 commonsourceibias.n418 161.3
R7957 commonsourceibias.n417 commonsourceibias.n386 161.3
R7958 commonsourceibias.n416 commonsourceibias.n415 161.3
R7959 commonsourceibias.n414 commonsourceibias.n413 161.3
R7960 commonsourceibias.n412 commonsourceibias.n388 161.3
R7961 commonsourceibias.n411 commonsourceibias.n410 161.3
R7962 commonsourceibias.n409 commonsourceibias.n408 161.3
R7963 commonsourceibias.n407 commonsourceibias.n390 161.3
R7964 commonsourceibias.n405 commonsourceibias.n404 161.3
R7965 commonsourceibias.n403 commonsourceibias.n391 161.3
R7966 commonsourceibias.n402 commonsourceibias.n401 161.3
R7967 commonsourceibias.n399 commonsourceibias.n392 161.3
R7968 commonsourceibias.n398 commonsourceibias.n397 161.3
R7969 commonsourceibias.n396 commonsourceibias.n393 161.3
R7970 commonsourceibias.n531 commonsourceibias.n383 161.3
R7971 commonsourceibias.n565 commonsourceibias.n374 161.3
R7972 commonsourceibias.n563 commonsourceibias.n562 161.3
R7973 commonsourceibias.n561 commonsourceibias.n375 161.3
R7974 commonsourceibias.n560 commonsourceibias.n559 161.3
R7975 commonsourceibias.n557 commonsourceibias.n376 161.3
R7976 commonsourceibias.n556 commonsourceibias.n555 161.3
R7977 commonsourceibias.n554 commonsourceibias.n377 161.3
R7978 commonsourceibias.n553 commonsourceibias.n552 161.3
R7979 commonsourceibias.n550 commonsourceibias.n378 161.3
R7980 commonsourceibias.n548 commonsourceibias.n547 161.3
R7981 commonsourceibias.n546 commonsourceibias.n379 161.3
R7982 commonsourceibias.n545 commonsourceibias.n544 161.3
R7983 commonsourceibias.n542 commonsourceibias.n380 161.3
R7984 commonsourceibias.n541 commonsourceibias.n540 161.3
R7985 commonsourceibias.n539 commonsourceibias.n381 161.3
R7986 commonsourceibias.n538 commonsourceibias.n537 161.3
R7987 commonsourceibias.n535 commonsourceibias.n382 161.3
R7988 commonsourceibias.n533 commonsourceibias.n532 161.3
R7989 commonsourceibias.n744 commonsourceibias.n658 161.3
R7990 commonsourceibias.n742 commonsourceibias.n741 161.3
R7991 commonsourceibias.n740 commonsourceibias.n659 161.3
R7992 commonsourceibias.n739 commonsourceibias.n738 161.3
R7993 commonsourceibias.n736 commonsourceibias.n660 161.3
R7994 commonsourceibias.n735 commonsourceibias.n734 161.3
R7995 commonsourceibias.n733 commonsourceibias.n661 161.3
R7996 commonsourceibias.n732 commonsourceibias.n731 161.3
R7997 commonsourceibias.n729 commonsourceibias.n662 161.3
R7998 commonsourceibias.n727 commonsourceibias.n726 161.3
R7999 commonsourceibias.n725 commonsourceibias.n663 161.3
R8000 commonsourceibias.n724 commonsourceibias.n723 161.3
R8001 commonsourceibias.n721 commonsourceibias.n664 161.3
R8002 commonsourceibias.n720 commonsourceibias.n719 161.3
R8003 commonsourceibias.n718 commonsourceibias.n665 161.3
R8004 commonsourceibias.n717 commonsourceibias.n716 161.3
R8005 commonsourceibias.n714 commonsourceibias.n666 161.3
R8006 commonsourceibias.n712 commonsourceibias.n711 161.3
R8007 commonsourceibias.n710 commonsourceibias.n667 161.3
R8008 commonsourceibias.n709 commonsourceibias.n708 161.3
R8009 commonsourceibias.n706 commonsourceibias.n668 161.3
R8010 commonsourceibias.n705 commonsourceibias.n704 161.3
R8011 commonsourceibias.n703 commonsourceibias.n702 161.3
R8012 commonsourceibias.n701 commonsourceibias.n670 161.3
R8013 commonsourceibias.n700 commonsourceibias.n699 161.3
R8014 commonsourceibias.n698 commonsourceibias.n697 161.3
R8015 commonsourceibias.n696 commonsourceibias.n672 161.3
R8016 commonsourceibias.n695 commonsourceibias.n694 161.3
R8017 commonsourceibias.n693 commonsourceibias.n692 161.3
R8018 commonsourceibias.n691 commonsourceibias.n674 161.3
R8019 commonsourceibias.n689 commonsourceibias.n688 161.3
R8020 commonsourceibias.n687 commonsourceibias.n675 161.3
R8021 commonsourceibias.n686 commonsourceibias.n685 161.3
R8022 commonsourceibias.n683 commonsourceibias.n676 161.3
R8023 commonsourceibias.n682 commonsourceibias.n681 161.3
R8024 commonsourceibias.n680 commonsourceibias.n677 161.3
R8025 commonsourceibias.n654 commonsourceibias.n568 161.3
R8026 commonsourceibias.n652 commonsourceibias.n651 161.3
R8027 commonsourceibias.n650 commonsourceibias.n569 161.3
R8028 commonsourceibias.n649 commonsourceibias.n648 161.3
R8029 commonsourceibias.n646 commonsourceibias.n570 161.3
R8030 commonsourceibias.n645 commonsourceibias.n644 161.3
R8031 commonsourceibias.n643 commonsourceibias.n571 161.3
R8032 commonsourceibias.n642 commonsourceibias.n641 161.3
R8033 commonsourceibias.n639 commonsourceibias.n572 161.3
R8034 commonsourceibias.n637 commonsourceibias.n636 161.3
R8035 commonsourceibias.n635 commonsourceibias.n573 161.3
R8036 commonsourceibias.n634 commonsourceibias.n633 161.3
R8037 commonsourceibias.n631 commonsourceibias.n574 161.3
R8038 commonsourceibias.n630 commonsourceibias.n629 161.3
R8039 commonsourceibias.n628 commonsourceibias.n575 161.3
R8040 commonsourceibias.n627 commonsourceibias.n626 161.3
R8041 commonsourceibias.n624 commonsourceibias.n576 161.3
R8042 commonsourceibias.n622 commonsourceibias.n621 161.3
R8043 commonsourceibias.n620 commonsourceibias.n577 161.3
R8044 commonsourceibias.n619 commonsourceibias.n618 161.3
R8045 commonsourceibias.n616 commonsourceibias.n578 161.3
R8046 commonsourceibias.n615 commonsourceibias.n614 161.3
R8047 commonsourceibias.n613 commonsourceibias.n612 161.3
R8048 commonsourceibias.n611 commonsourceibias.n580 161.3
R8049 commonsourceibias.n610 commonsourceibias.n609 161.3
R8050 commonsourceibias.n608 commonsourceibias.n607 161.3
R8051 commonsourceibias.n606 commonsourceibias.n582 161.3
R8052 commonsourceibias.n605 commonsourceibias.n604 161.3
R8053 commonsourceibias.n603 commonsourceibias.n602 161.3
R8054 commonsourceibias.n601 commonsourceibias.n584 161.3
R8055 commonsourceibias.n599 commonsourceibias.n598 161.3
R8056 commonsourceibias.n597 commonsourceibias.n585 161.3
R8057 commonsourceibias.n596 commonsourceibias.n595 161.3
R8058 commonsourceibias.n593 commonsourceibias.n586 161.3
R8059 commonsourceibias.n592 commonsourceibias.n591 161.3
R8060 commonsourceibias.n590 commonsourceibias.n587 161.3
R8061 commonsourceibias.n111 commonsourceibias.n109 81.5057
R8062 commonsourceibias.n428 commonsourceibias.n426 81.5057
R8063 commonsourceibias.n111 commonsourceibias.n110 80.9324
R8064 commonsourceibias.n113 commonsourceibias.n112 80.9324
R8065 commonsourceibias.n115 commonsourceibias.n114 80.9324
R8066 commonsourceibias.n108 commonsourceibias.n107 80.9324
R8067 commonsourceibias.n106 commonsourceibias.n105 80.9324
R8068 commonsourceibias.n104 commonsourceibias.n103 80.9324
R8069 commonsourceibias.n102 commonsourceibias.n101 80.9324
R8070 commonsourceibias.n523 commonsourceibias.n522 80.9324
R8071 commonsourceibias.n525 commonsourceibias.n524 80.9324
R8072 commonsourceibias.n527 commonsourceibias.n526 80.9324
R8073 commonsourceibias.n529 commonsourceibias.n528 80.9324
R8074 commonsourceibias.n432 commonsourceibias.n431 80.9324
R8075 commonsourceibias.n430 commonsourceibias.n429 80.9324
R8076 commonsourceibias.n428 commonsourceibias.n427 80.9324
R8077 commonsourceibias.n100 commonsourceibias.n99 80.6037
R8078 commonsourceibias.n193 commonsourceibias.n192 80.6037
R8079 commonsourceibias.n372 commonsourceibias.n371 80.6037
R8080 commonsourceibias.n282 commonsourceibias.n281 80.6037
R8081 commonsourceibias.n521 commonsourceibias.n520 80.6037
R8082 commonsourceibias.n567 commonsourceibias.n566 80.6037
R8083 commonsourceibias.n746 commonsourceibias.n745 80.6037
R8084 commonsourceibias.n656 commonsourceibias.n655 80.6037
R8085 commonsourceibias.n85 commonsourceibias.n84 56.5617
R8086 commonsourceibias.n71 commonsourceibias.n70 56.5617
R8087 commonsourceibias.n62 commonsourceibias.n61 56.5617
R8088 commonsourceibias.n48 commonsourceibias.n47 56.5617
R8089 commonsourceibias.n178 commonsourceibias.n177 56.5617
R8090 commonsourceibias.n164 commonsourceibias.n163 56.5617
R8091 commonsourceibias.n155 commonsourceibias.n154 56.5617
R8092 commonsourceibias.n141 commonsourceibias.n140 56.5617
R8093 commonsourceibias.n320 commonsourceibias.n319 56.5617
R8094 commonsourceibias.n334 commonsourceibias.n333 56.5617
R8095 commonsourceibias.n343 commonsourceibias.n342 56.5617
R8096 commonsourceibias.n357 commonsourceibias.n356 56.5617
R8097 commonsourceibias.n267 commonsourceibias.n266 56.5617
R8098 commonsourceibias.n253 commonsourceibias.n252 56.5617
R8099 commonsourceibias.n244 commonsourceibias.n243 56.5617
R8100 commonsourceibias.n230 commonsourceibias.n229 56.5617
R8101 commonsourceibias.n467 commonsourceibias.n466 56.5617
R8102 commonsourceibias.n481 commonsourceibias.n480 56.5617
R8103 commonsourceibias.n491 commonsourceibias.n489 56.5617
R8104 commonsourceibias.n506 commonsourceibias.n504 56.5617
R8105 commonsourceibias.n552 commonsourceibias.n550 56.5617
R8106 commonsourceibias.n537 commonsourceibias.n535 56.5617
R8107 commonsourceibias.n408 commonsourceibias.n407 56.5617
R8108 commonsourceibias.n422 commonsourceibias.n421 56.5617
R8109 commonsourceibias.n692 commonsourceibias.n691 56.5617
R8110 commonsourceibias.n706 commonsourceibias.n705 56.5617
R8111 commonsourceibias.n716 commonsourceibias.n714 56.5617
R8112 commonsourceibias.n731 commonsourceibias.n729 56.5617
R8113 commonsourceibias.n602 commonsourceibias.n601 56.5617
R8114 commonsourceibias.n616 commonsourceibias.n615 56.5617
R8115 commonsourceibias.n626 commonsourceibias.n624 56.5617
R8116 commonsourceibias.n641 commonsourceibias.n639 56.5617
R8117 commonsourceibias.n76 commonsourceibias.n75 56.0773
R8118 commonsourceibias.n57 commonsourceibias.n56 56.0773
R8119 commonsourceibias.n169 commonsourceibias.n168 56.0773
R8120 commonsourceibias.n150 commonsourceibias.n149 56.0773
R8121 commonsourceibias.n329 commonsourceibias.n328 56.0773
R8122 commonsourceibias.n348 commonsourceibias.n347 56.0773
R8123 commonsourceibias.n258 commonsourceibias.n257 56.0773
R8124 commonsourceibias.n239 commonsourceibias.n238 56.0773
R8125 commonsourceibias.n476 commonsourceibias.n475 56.0773
R8126 commonsourceibias.n496 commonsourceibias.n495 56.0773
R8127 commonsourceibias.n542 commonsourceibias.n541 56.0773
R8128 commonsourceibias.n417 commonsourceibias.n416 56.0773
R8129 commonsourceibias.n701 commonsourceibias.n700 56.0773
R8130 commonsourceibias.n721 commonsourceibias.n720 56.0773
R8131 commonsourceibias.n611 commonsourceibias.n610 56.0773
R8132 commonsourceibias.n631 commonsourceibias.n630 56.0773
R8133 commonsourceibias.n99 commonsourceibias.n98 55.3321
R8134 commonsourceibias.n192 commonsourceibias.n191 55.3321
R8135 commonsourceibias.n371 commonsourceibias.n370 55.3321
R8136 commonsourceibias.n281 commonsourceibias.n280 55.3321
R8137 commonsourceibias.n520 commonsourceibias.n519 55.3321
R8138 commonsourceibias.n566 commonsourceibias.n565 55.3321
R8139 commonsourceibias.n745 commonsourceibias.n744 55.3321
R8140 commonsourceibias.n655 commonsourceibias.n654 55.3321
R8141 commonsourceibias.n90 commonsourceibias.n89 55.1086
R8142 commonsourceibias.n41 commonsourceibias.n31 55.1086
R8143 commonsourceibias.n183 commonsourceibias.n182 55.1086
R8144 commonsourceibias.n134 commonsourceibias.n124 55.1086
R8145 commonsourceibias.n313 commonsourceibias.n303 55.1086
R8146 commonsourceibias.n362 commonsourceibias.n361 55.1086
R8147 commonsourceibias.n272 commonsourceibias.n271 55.1086
R8148 commonsourceibias.n223 commonsourceibias.n213 55.1086
R8149 commonsourceibias.n460 commonsourceibias.n450 55.1086
R8150 commonsourceibias.n511 commonsourceibias.n510 55.1086
R8151 commonsourceibias.n557 commonsourceibias.n556 55.1086
R8152 commonsourceibias.n401 commonsourceibias.n391 55.1086
R8153 commonsourceibias.n685 commonsourceibias.n675 55.1086
R8154 commonsourceibias.n736 commonsourceibias.n735 55.1086
R8155 commonsourceibias.n595 commonsourceibias.n585 55.1086
R8156 commonsourceibias.n646 commonsourceibias.n645 55.1086
R8157 commonsourceibias.n35 commonsourceibias.n34 47.4592
R8158 commonsourceibias.n128 commonsourceibias.n127 47.4592
R8159 commonsourceibias.n307 commonsourceibias.n306 47.4592
R8160 commonsourceibias.n217 commonsourceibias.n216 47.4592
R8161 commonsourceibias.n454 commonsourceibias.n453 47.4592
R8162 commonsourceibias.n395 commonsourceibias.n394 47.4592
R8163 commonsourceibias.n679 commonsourceibias.n678 47.4592
R8164 commonsourceibias.n589 commonsourceibias.n588 47.4592
R8165 commonsourceibias.n308 commonsourceibias.n307 44.0436
R8166 commonsourceibias.n455 commonsourceibias.n454 44.0436
R8167 commonsourceibias.n396 commonsourceibias.n395 44.0436
R8168 commonsourceibias.n680 commonsourceibias.n679 44.0436
R8169 commonsourceibias.n590 commonsourceibias.n589 44.0436
R8170 commonsourceibias.n36 commonsourceibias.n35 44.0436
R8171 commonsourceibias.n129 commonsourceibias.n128 44.0436
R8172 commonsourceibias.n218 commonsourceibias.n217 44.0436
R8173 commonsourceibias.n92 commonsourceibias.n13 42.5146
R8174 commonsourceibias.n39 commonsourceibias.n38 42.5146
R8175 commonsourceibias.n185 commonsourceibias.n1 42.5146
R8176 commonsourceibias.n132 commonsourceibias.n131 42.5146
R8177 commonsourceibias.n311 commonsourceibias.n310 42.5146
R8178 commonsourceibias.n364 commonsourceibias.n285 42.5146
R8179 commonsourceibias.n274 commonsourceibias.n195 42.5146
R8180 commonsourceibias.n221 commonsourceibias.n220 42.5146
R8181 commonsourceibias.n458 commonsourceibias.n457 42.5146
R8182 commonsourceibias.n513 commonsourceibias.n434 42.5146
R8183 commonsourceibias.n559 commonsourceibias.n375 42.5146
R8184 commonsourceibias.n399 commonsourceibias.n398 42.5146
R8185 commonsourceibias.n683 commonsourceibias.n682 42.5146
R8186 commonsourceibias.n738 commonsourceibias.n659 42.5146
R8187 commonsourceibias.n593 commonsourceibias.n592 42.5146
R8188 commonsourceibias.n648 commonsourceibias.n569 42.5146
R8189 commonsourceibias.n78 commonsourceibias.n18 41.5458
R8190 commonsourceibias.n53 commonsourceibias.n52 41.5458
R8191 commonsourceibias.n171 commonsourceibias.n6 41.5458
R8192 commonsourceibias.n146 commonsourceibias.n145 41.5458
R8193 commonsourceibias.n325 commonsourceibias.n324 41.5458
R8194 commonsourceibias.n350 commonsourceibias.n290 41.5458
R8195 commonsourceibias.n260 commonsourceibias.n200 41.5458
R8196 commonsourceibias.n235 commonsourceibias.n234 41.5458
R8197 commonsourceibias.n472 commonsourceibias.n471 41.5458
R8198 commonsourceibias.n498 commonsourceibias.n438 41.5458
R8199 commonsourceibias.n544 commonsourceibias.n379 41.5458
R8200 commonsourceibias.n413 commonsourceibias.n412 41.5458
R8201 commonsourceibias.n697 commonsourceibias.n696 41.5458
R8202 commonsourceibias.n723 commonsourceibias.n663 41.5458
R8203 commonsourceibias.n607 commonsourceibias.n606 41.5458
R8204 commonsourceibias.n633 commonsourceibias.n573 41.5458
R8205 commonsourceibias.n68 commonsourceibias.n23 40.577
R8206 commonsourceibias.n64 commonsourceibias.n23 40.577
R8207 commonsourceibias.n161 commonsourceibias.n11 40.577
R8208 commonsourceibias.n157 commonsourceibias.n11 40.577
R8209 commonsourceibias.n336 commonsourceibias.n295 40.577
R8210 commonsourceibias.n340 commonsourceibias.n295 40.577
R8211 commonsourceibias.n250 commonsourceibias.n205 40.577
R8212 commonsourceibias.n246 commonsourceibias.n205 40.577
R8213 commonsourceibias.n483 commonsourceibias.n442 40.577
R8214 commonsourceibias.n487 commonsourceibias.n442 40.577
R8215 commonsourceibias.n533 commonsourceibias.n383 40.577
R8216 commonsourceibias.n424 commonsourceibias.n383 40.577
R8217 commonsourceibias.n708 commonsourceibias.n667 40.577
R8218 commonsourceibias.n712 commonsourceibias.n667 40.577
R8219 commonsourceibias.n618 commonsourceibias.n577 40.577
R8220 commonsourceibias.n622 commonsourceibias.n577 40.577
R8221 commonsourceibias.n82 commonsourceibias.n18 39.6083
R8222 commonsourceibias.n52 commonsourceibias.n51 39.6083
R8223 commonsourceibias.n175 commonsourceibias.n6 39.6083
R8224 commonsourceibias.n145 commonsourceibias.n144 39.6083
R8225 commonsourceibias.n324 commonsourceibias.n323 39.6083
R8226 commonsourceibias.n354 commonsourceibias.n290 39.6083
R8227 commonsourceibias.n264 commonsourceibias.n200 39.6083
R8228 commonsourceibias.n234 commonsourceibias.n233 39.6083
R8229 commonsourceibias.n471 commonsourceibias.n470 39.6083
R8230 commonsourceibias.n502 commonsourceibias.n438 39.6083
R8231 commonsourceibias.n548 commonsourceibias.n379 39.6083
R8232 commonsourceibias.n412 commonsourceibias.n411 39.6083
R8233 commonsourceibias.n696 commonsourceibias.n695 39.6083
R8234 commonsourceibias.n727 commonsourceibias.n663 39.6083
R8235 commonsourceibias.n606 commonsourceibias.n605 39.6083
R8236 commonsourceibias.n637 commonsourceibias.n573 39.6083
R8237 commonsourceibias.n96 commonsourceibias.n13 38.6395
R8238 commonsourceibias.n38 commonsourceibias.n33 38.6395
R8239 commonsourceibias.n189 commonsourceibias.n1 38.6395
R8240 commonsourceibias.n131 commonsourceibias.n126 38.6395
R8241 commonsourceibias.n310 commonsourceibias.n305 38.6395
R8242 commonsourceibias.n368 commonsourceibias.n285 38.6395
R8243 commonsourceibias.n278 commonsourceibias.n195 38.6395
R8244 commonsourceibias.n220 commonsourceibias.n215 38.6395
R8245 commonsourceibias.n457 commonsourceibias.n452 38.6395
R8246 commonsourceibias.n517 commonsourceibias.n434 38.6395
R8247 commonsourceibias.n563 commonsourceibias.n375 38.6395
R8248 commonsourceibias.n398 commonsourceibias.n393 38.6395
R8249 commonsourceibias.n682 commonsourceibias.n677 38.6395
R8250 commonsourceibias.n742 commonsourceibias.n659 38.6395
R8251 commonsourceibias.n592 commonsourceibias.n587 38.6395
R8252 commonsourceibias.n652 commonsourceibias.n569 38.6395
R8253 commonsourceibias.n89 commonsourceibias.n15 26.0455
R8254 commonsourceibias.n45 commonsourceibias.n31 26.0455
R8255 commonsourceibias.n182 commonsourceibias.n3 26.0455
R8256 commonsourceibias.n138 commonsourceibias.n124 26.0455
R8257 commonsourceibias.n317 commonsourceibias.n303 26.0455
R8258 commonsourceibias.n361 commonsourceibias.n287 26.0455
R8259 commonsourceibias.n271 commonsourceibias.n197 26.0455
R8260 commonsourceibias.n227 commonsourceibias.n213 26.0455
R8261 commonsourceibias.n464 commonsourceibias.n450 26.0455
R8262 commonsourceibias.n510 commonsourceibias.n436 26.0455
R8263 commonsourceibias.n556 commonsourceibias.n377 26.0455
R8264 commonsourceibias.n405 commonsourceibias.n391 26.0455
R8265 commonsourceibias.n689 commonsourceibias.n675 26.0455
R8266 commonsourceibias.n735 commonsourceibias.n661 26.0455
R8267 commonsourceibias.n599 commonsourceibias.n585 26.0455
R8268 commonsourceibias.n645 commonsourceibias.n571 26.0455
R8269 commonsourceibias.n75 commonsourceibias.n20 25.0767
R8270 commonsourceibias.n58 commonsourceibias.n57 25.0767
R8271 commonsourceibias.n168 commonsourceibias.n8 25.0767
R8272 commonsourceibias.n151 commonsourceibias.n150 25.0767
R8273 commonsourceibias.n330 commonsourceibias.n329 25.0767
R8274 commonsourceibias.n347 commonsourceibias.n292 25.0767
R8275 commonsourceibias.n257 commonsourceibias.n202 25.0767
R8276 commonsourceibias.n240 commonsourceibias.n239 25.0767
R8277 commonsourceibias.n477 commonsourceibias.n476 25.0767
R8278 commonsourceibias.n495 commonsourceibias.n440 25.0767
R8279 commonsourceibias.n541 commonsourceibias.n381 25.0767
R8280 commonsourceibias.n418 commonsourceibias.n417 25.0767
R8281 commonsourceibias.n702 commonsourceibias.n701 25.0767
R8282 commonsourceibias.n720 commonsourceibias.n665 25.0767
R8283 commonsourceibias.n612 commonsourceibias.n611 25.0767
R8284 commonsourceibias.n630 commonsourceibias.n575 25.0767
R8285 commonsourceibias.n71 commonsourceibias.n22 24.3464
R8286 commonsourceibias.n61 commonsourceibias.n25 24.3464
R8287 commonsourceibias.n164 commonsourceibias.n10 24.3464
R8288 commonsourceibias.n154 commonsourceibias.n118 24.3464
R8289 commonsourceibias.n333 commonsourceibias.n297 24.3464
R8290 commonsourceibias.n343 commonsourceibias.n294 24.3464
R8291 commonsourceibias.n253 commonsourceibias.n204 24.3464
R8292 commonsourceibias.n243 commonsourceibias.n207 24.3464
R8293 commonsourceibias.n480 commonsourceibias.n444 24.3464
R8294 commonsourceibias.n491 commonsourceibias.n490 24.3464
R8295 commonsourceibias.n537 commonsourceibias.n536 24.3464
R8296 commonsourceibias.n421 commonsourceibias.n385 24.3464
R8297 commonsourceibias.n705 commonsourceibias.n669 24.3464
R8298 commonsourceibias.n716 commonsourceibias.n715 24.3464
R8299 commonsourceibias.n615 commonsourceibias.n579 24.3464
R8300 commonsourceibias.n626 commonsourceibias.n625 24.3464
R8301 commonsourceibias.n85 commonsourceibias.n17 23.8546
R8302 commonsourceibias.n47 commonsourceibias.n46 23.8546
R8303 commonsourceibias.n178 commonsourceibias.n5 23.8546
R8304 commonsourceibias.n140 commonsourceibias.n139 23.8546
R8305 commonsourceibias.n319 commonsourceibias.n318 23.8546
R8306 commonsourceibias.n357 commonsourceibias.n289 23.8546
R8307 commonsourceibias.n267 commonsourceibias.n199 23.8546
R8308 commonsourceibias.n229 commonsourceibias.n228 23.8546
R8309 commonsourceibias.n466 commonsourceibias.n465 23.8546
R8310 commonsourceibias.n506 commonsourceibias.n505 23.8546
R8311 commonsourceibias.n552 commonsourceibias.n551 23.8546
R8312 commonsourceibias.n407 commonsourceibias.n406 23.8546
R8313 commonsourceibias.n691 commonsourceibias.n690 23.8546
R8314 commonsourceibias.n731 commonsourceibias.n730 23.8546
R8315 commonsourceibias.n601 commonsourceibias.n600 23.8546
R8316 commonsourceibias.n641 commonsourceibias.n640 23.8546
R8317 commonsourceibias.n98 commonsourceibias.n97 17.4607
R8318 commonsourceibias.n191 commonsourceibias.n190 17.4607
R8319 commonsourceibias.n370 commonsourceibias.n369 17.4607
R8320 commonsourceibias.n280 commonsourceibias.n279 17.4607
R8321 commonsourceibias.n519 commonsourceibias.n518 17.4607
R8322 commonsourceibias.n565 commonsourceibias.n564 17.4607
R8323 commonsourceibias.n744 commonsourceibias.n743 17.4607
R8324 commonsourceibias.n654 commonsourceibias.n653 17.4607
R8325 commonsourceibias.n84 commonsourceibias.n83 16.9689
R8326 commonsourceibias.n48 commonsourceibias.n29 16.9689
R8327 commonsourceibias.n177 commonsourceibias.n176 16.9689
R8328 commonsourceibias.n141 commonsourceibias.n122 16.9689
R8329 commonsourceibias.n320 commonsourceibias.n301 16.9689
R8330 commonsourceibias.n356 commonsourceibias.n355 16.9689
R8331 commonsourceibias.n266 commonsourceibias.n265 16.9689
R8332 commonsourceibias.n230 commonsourceibias.n211 16.9689
R8333 commonsourceibias.n467 commonsourceibias.n448 16.9689
R8334 commonsourceibias.n504 commonsourceibias.n503 16.9689
R8335 commonsourceibias.n550 commonsourceibias.n549 16.9689
R8336 commonsourceibias.n408 commonsourceibias.n389 16.9689
R8337 commonsourceibias.n692 commonsourceibias.n673 16.9689
R8338 commonsourceibias.n729 commonsourceibias.n728 16.9689
R8339 commonsourceibias.n602 commonsourceibias.n583 16.9689
R8340 commonsourceibias.n639 commonsourceibias.n638 16.9689
R8341 commonsourceibias.n70 commonsourceibias.n69 16.477
R8342 commonsourceibias.n63 commonsourceibias.n62 16.477
R8343 commonsourceibias.n163 commonsourceibias.n162 16.477
R8344 commonsourceibias.n156 commonsourceibias.n155 16.477
R8345 commonsourceibias.n335 commonsourceibias.n334 16.477
R8346 commonsourceibias.n342 commonsourceibias.n341 16.477
R8347 commonsourceibias.n252 commonsourceibias.n251 16.477
R8348 commonsourceibias.n245 commonsourceibias.n244 16.477
R8349 commonsourceibias.n482 commonsourceibias.n481 16.477
R8350 commonsourceibias.n489 commonsourceibias.n488 16.477
R8351 commonsourceibias.n535 commonsourceibias.n534 16.477
R8352 commonsourceibias.n423 commonsourceibias.n422 16.477
R8353 commonsourceibias.n707 commonsourceibias.n706 16.477
R8354 commonsourceibias.n714 commonsourceibias.n713 16.477
R8355 commonsourceibias.n617 commonsourceibias.n616 16.477
R8356 commonsourceibias.n624 commonsourceibias.n623 16.477
R8357 commonsourceibias.n77 commonsourceibias.n76 15.9852
R8358 commonsourceibias.n56 commonsourceibias.n27 15.9852
R8359 commonsourceibias.n170 commonsourceibias.n169 15.9852
R8360 commonsourceibias.n149 commonsourceibias.n120 15.9852
R8361 commonsourceibias.n328 commonsourceibias.n299 15.9852
R8362 commonsourceibias.n349 commonsourceibias.n348 15.9852
R8363 commonsourceibias.n259 commonsourceibias.n258 15.9852
R8364 commonsourceibias.n238 commonsourceibias.n209 15.9852
R8365 commonsourceibias.n475 commonsourceibias.n446 15.9852
R8366 commonsourceibias.n497 commonsourceibias.n496 15.9852
R8367 commonsourceibias.n543 commonsourceibias.n542 15.9852
R8368 commonsourceibias.n416 commonsourceibias.n387 15.9852
R8369 commonsourceibias.n700 commonsourceibias.n671 15.9852
R8370 commonsourceibias.n722 commonsourceibias.n721 15.9852
R8371 commonsourceibias.n610 commonsourceibias.n581 15.9852
R8372 commonsourceibias.n632 commonsourceibias.n631 15.9852
R8373 commonsourceibias.n91 commonsourceibias.n90 15.4934
R8374 commonsourceibias.n41 commonsourceibias.n40 15.4934
R8375 commonsourceibias.n184 commonsourceibias.n183 15.4934
R8376 commonsourceibias.n134 commonsourceibias.n133 15.4934
R8377 commonsourceibias.n313 commonsourceibias.n312 15.4934
R8378 commonsourceibias.n363 commonsourceibias.n362 15.4934
R8379 commonsourceibias.n273 commonsourceibias.n272 15.4934
R8380 commonsourceibias.n223 commonsourceibias.n222 15.4934
R8381 commonsourceibias.n460 commonsourceibias.n459 15.4934
R8382 commonsourceibias.n512 commonsourceibias.n511 15.4934
R8383 commonsourceibias.n558 commonsourceibias.n557 15.4934
R8384 commonsourceibias.n401 commonsourceibias.n400 15.4934
R8385 commonsourceibias.n685 commonsourceibias.n684 15.4934
R8386 commonsourceibias.n737 commonsourceibias.n736 15.4934
R8387 commonsourceibias.n595 commonsourceibias.n594 15.4934
R8388 commonsourceibias.n647 commonsourceibias.n646 15.4934
R8389 commonsourceibias.n102 commonsourceibias.n100 13.2663
R8390 commonsourceibias.n523 commonsourceibias.n521 13.2663
R8391 commonsourceibias.n748 commonsourceibias.n373 10.4122
R8392 commonsourceibias.n159 commonsourceibias.n116 9.50363
R8393 commonsourceibias.n531 commonsourceibias.n530 9.50363
R8394 commonsourceibias.n92 commonsourceibias.n91 9.09948
R8395 commonsourceibias.n40 commonsourceibias.n39 9.09948
R8396 commonsourceibias.n185 commonsourceibias.n184 9.09948
R8397 commonsourceibias.n133 commonsourceibias.n132 9.09948
R8398 commonsourceibias.n312 commonsourceibias.n311 9.09948
R8399 commonsourceibias.n364 commonsourceibias.n363 9.09948
R8400 commonsourceibias.n274 commonsourceibias.n273 9.09948
R8401 commonsourceibias.n222 commonsourceibias.n221 9.09948
R8402 commonsourceibias.n459 commonsourceibias.n458 9.09948
R8403 commonsourceibias.n513 commonsourceibias.n512 9.09948
R8404 commonsourceibias.n559 commonsourceibias.n558 9.09948
R8405 commonsourceibias.n400 commonsourceibias.n399 9.09948
R8406 commonsourceibias.n684 commonsourceibias.n683 9.09948
R8407 commonsourceibias.n738 commonsourceibias.n737 9.09948
R8408 commonsourceibias.n594 commonsourceibias.n593 9.09948
R8409 commonsourceibias.n648 commonsourceibias.n647 9.09948
R8410 commonsourceibias.n283 commonsourceibias.n193 8.79451
R8411 commonsourceibias.n657 commonsourceibias.n567 8.79451
R8412 commonsourceibias.n78 commonsourceibias.n77 8.60764
R8413 commonsourceibias.n53 commonsourceibias.n27 8.60764
R8414 commonsourceibias.n171 commonsourceibias.n170 8.60764
R8415 commonsourceibias.n146 commonsourceibias.n120 8.60764
R8416 commonsourceibias.n325 commonsourceibias.n299 8.60764
R8417 commonsourceibias.n350 commonsourceibias.n349 8.60764
R8418 commonsourceibias.n260 commonsourceibias.n259 8.60764
R8419 commonsourceibias.n235 commonsourceibias.n209 8.60764
R8420 commonsourceibias.n472 commonsourceibias.n446 8.60764
R8421 commonsourceibias.n498 commonsourceibias.n497 8.60764
R8422 commonsourceibias.n544 commonsourceibias.n543 8.60764
R8423 commonsourceibias.n413 commonsourceibias.n387 8.60764
R8424 commonsourceibias.n697 commonsourceibias.n671 8.60764
R8425 commonsourceibias.n723 commonsourceibias.n722 8.60764
R8426 commonsourceibias.n607 commonsourceibias.n581 8.60764
R8427 commonsourceibias.n633 commonsourceibias.n632 8.60764
R8428 commonsourceibias.n748 commonsourceibias.n747 8.46921
R8429 commonsourceibias.n69 commonsourceibias.n68 8.11581
R8430 commonsourceibias.n64 commonsourceibias.n63 8.11581
R8431 commonsourceibias.n162 commonsourceibias.n161 8.11581
R8432 commonsourceibias.n157 commonsourceibias.n156 8.11581
R8433 commonsourceibias.n336 commonsourceibias.n335 8.11581
R8434 commonsourceibias.n341 commonsourceibias.n340 8.11581
R8435 commonsourceibias.n251 commonsourceibias.n250 8.11581
R8436 commonsourceibias.n246 commonsourceibias.n245 8.11581
R8437 commonsourceibias.n483 commonsourceibias.n482 8.11581
R8438 commonsourceibias.n488 commonsourceibias.n487 8.11581
R8439 commonsourceibias.n534 commonsourceibias.n533 8.11581
R8440 commonsourceibias.n424 commonsourceibias.n423 8.11581
R8441 commonsourceibias.n708 commonsourceibias.n707 8.11581
R8442 commonsourceibias.n713 commonsourceibias.n712 8.11581
R8443 commonsourceibias.n618 commonsourceibias.n617 8.11581
R8444 commonsourceibias.n623 commonsourceibias.n622 8.11581
R8445 commonsourceibias.n83 commonsourceibias.n82 7.62397
R8446 commonsourceibias.n51 commonsourceibias.n29 7.62397
R8447 commonsourceibias.n176 commonsourceibias.n175 7.62397
R8448 commonsourceibias.n144 commonsourceibias.n122 7.62397
R8449 commonsourceibias.n323 commonsourceibias.n301 7.62397
R8450 commonsourceibias.n355 commonsourceibias.n354 7.62397
R8451 commonsourceibias.n265 commonsourceibias.n264 7.62397
R8452 commonsourceibias.n233 commonsourceibias.n211 7.62397
R8453 commonsourceibias.n470 commonsourceibias.n448 7.62397
R8454 commonsourceibias.n503 commonsourceibias.n502 7.62397
R8455 commonsourceibias.n549 commonsourceibias.n548 7.62397
R8456 commonsourceibias.n411 commonsourceibias.n389 7.62397
R8457 commonsourceibias.n695 commonsourceibias.n673 7.62397
R8458 commonsourceibias.n728 commonsourceibias.n727 7.62397
R8459 commonsourceibias.n605 commonsourceibias.n583 7.62397
R8460 commonsourceibias.n638 commonsourceibias.n637 7.62397
R8461 commonsourceibias.n97 commonsourceibias.n96 7.13213
R8462 commonsourceibias.n34 commonsourceibias.n33 7.13213
R8463 commonsourceibias.n190 commonsourceibias.n189 7.13213
R8464 commonsourceibias.n127 commonsourceibias.n126 7.13213
R8465 commonsourceibias.n306 commonsourceibias.n305 7.13213
R8466 commonsourceibias.n369 commonsourceibias.n368 7.13213
R8467 commonsourceibias.n279 commonsourceibias.n278 7.13213
R8468 commonsourceibias.n216 commonsourceibias.n215 7.13213
R8469 commonsourceibias.n453 commonsourceibias.n452 7.13213
R8470 commonsourceibias.n518 commonsourceibias.n517 7.13213
R8471 commonsourceibias.n564 commonsourceibias.n563 7.13213
R8472 commonsourceibias.n394 commonsourceibias.n393 7.13213
R8473 commonsourceibias.n678 commonsourceibias.n677 7.13213
R8474 commonsourceibias.n743 commonsourceibias.n742 7.13213
R8475 commonsourceibias.n588 commonsourceibias.n587 7.13213
R8476 commonsourceibias.n653 commonsourceibias.n652 7.13213
R8477 commonsourceibias.n373 commonsourceibias.n372 5.06534
R8478 commonsourceibias.n283 commonsourceibias.n282 5.06534
R8479 commonsourceibias.n747 commonsourceibias.n746 5.06534
R8480 commonsourceibias.n657 commonsourceibias.n656 5.06534
R8481 commonsourceibias commonsourceibias.n748 4.04308
R8482 commonsourceibias.n373 commonsourceibias.n283 3.72967
R8483 commonsourceibias.n747 commonsourceibias.n657 3.72967
R8484 commonsourceibias.n109 commonsourceibias.t31 2.82907
R8485 commonsourceibias.n109 commonsourceibias.t55 2.82907
R8486 commonsourceibias.n110 commonsourceibias.t21 2.82907
R8487 commonsourceibias.n110 commonsourceibias.t57 2.82907
R8488 commonsourceibias.n112 commonsourceibias.t3 2.82907
R8489 commonsourceibias.n112 commonsourceibias.t29 2.82907
R8490 commonsourceibias.n114 commonsourceibias.t47 2.82907
R8491 commonsourceibias.n114 commonsourceibias.t23 2.82907
R8492 commonsourceibias.n107 commonsourceibias.t9 2.82907
R8493 commonsourceibias.n107 commonsourceibias.t15 2.82907
R8494 commonsourceibias.n105 commonsourceibias.t19 2.82907
R8495 commonsourceibias.n105 commonsourceibias.t17 2.82907
R8496 commonsourceibias.n103 commonsourceibias.t5 2.82907
R8497 commonsourceibias.n103 commonsourceibias.t45 2.82907
R8498 commonsourceibias.n101 commonsourceibias.t59 2.82907
R8499 commonsourceibias.n101 commonsourceibias.t53 2.82907
R8500 commonsourceibias.n522 commonsourceibias.t25 2.82907
R8501 commonsourceibias.n522 commonsourceibias.t41 2.82907
R8502 commonsourceibias.n524 commonsourceibias.t11 2.82907
R8503 commonsourceibias.n524 commonsourceibias.t33 2.82907
R8504 commonsourceibias.n526 commonsourceibias.t27 2.82907
R8505 commonsourceibias.n526 commonsourceibias.t35 2.82907
R8506 commonsourceibias.n528 commonsourceibias.t63 2.82907
R8507 commonsourceibias.n528 commonsourceibias.t7 2.82907
R8508 commonsourceibias.n431 commonsourceibias.t39 2.82907
R8509 commonsourceibias.n431 commonsourceibias.t13 2.82907
R8510 commonsourceibias.n429 commonsourceibias.t1 2.82907
R8511 commonsourceibias.n429 commonsourceibias.t61 2.82907
R8512 commonsourceibias.n427 commonsourceibias.t43 2.82907
R8513 commonsourceibias.n427 commonsourceibias.t37 2.82907
R8514 commonsourceibias.n426 commonsourceibias.t51 2.82907
R8515 commonsourceibias.n426 commonsourceibias.t49 2.82907
R8516 commonsourceibias.n17 commonsourceibias.n15 0.738255
R8517 commonsourceibias.n46 commonsourceibias.n45 0.738255
R8518 commonsourceibias.n5 commonsourceibias.n3 0.738255
R8519 commonsourceibias.n139 commonsourceibias.n138 0.738255
R8520 commonsourceibias.n318 commonsourceibias.n317 0.738255
R8521 commonsourceibias.n289 commonsourceibias.n287 0.738255
R8522 commonsourceibias.n199 commonsourceibias.n197 0.738255
R8523 commonsourceibias.n228 commonsourceibias.n227 0.738255
R8524 commonsourceibias.n465 commonsourceibias.n464 0.738255
R8525 commonsourceibias.n505 commonsourceibias.n436 0.738255
R8526 commonsourceibias.n551 commonsourceibias.n377 0.738255
R8527 commonsourceibias.n406 commonsourceibias.n405 0.738255
R8528 commonsourceibias.n690 commonsourceibias.n689 0.738255
R8529 commonsourceibias.n730 commonsourceibias.n661 0.738255
R8530 commonsourceibias.n600 commonsourceibias.n599 0.738255
R8531 commonsourceibias.n640 commonsourceibias.n571 0.738255
R8532 commonsourceibias.n104 commonsourceibias.n102 0.573776
R8533 commonsourceibias.n106 commonsourceibias.n104 0.573776
R8534 commonsourceibias.n108 commonsourceibias.n106 0.573776
R8535 commonsourceibias.n115 commonsourceibias.n113 0.573776
R8536 commonsourceibias.n113 commonsourceibias.n111 0.573776
R8537 commonsourceibias.n430 commonsourceibias.n428 0.573776
R8538 commonsourceibias.n432 commonsourceibias.n430 0.573776
R8539 commonsourceibias.n529 commonsourceibias.n527 0.573776
R8540 commonsourceibias.n527 commonsourceibias.n525 0.573776
R8541 commonsourceibias.n525 commonsourceibias.n523 0.573776
R8542 commonsourceibias.n116 commonsourceibias.n108 0.287138
R8543 commonsourceibias.n116 commonsourceibias.n115 0.287138
R8544 commonsourceibias.n530 commonsourceibias.n432 0.287138
R8545 commonsourceibias.n530 commonsourceibias.n529 0.287138
R8546 commonsourceibias.n100 commonsourceibias.n12 0.285035
R8547 commonsourceibias.n193 commonsourceibias.n0 0.285035
R8548 commonsourceibias.n372 commonsourceibias.n284 0.285035
R8549 commonsourceibias.n282 commonsourceibias.n194 0.285035
R8550 commonsourceibias.n521 commonsourceibias.n433 0.285035
R8551 commonsourceibias.n567 commonsourceibias.n374 0.285035
R8552 commonsourceibias.n746 commonsourceibias.n658 0.285035
R8553 commonsourceibias.n656 commonsourceibias.n568 0.285035
R8554 commonsourceibias.n22 commonsourceibias.n20 0.246418
R8555 commonsourceibias.n58 commonsourceibias.n25 0.246418
R8556 commonsourceibias.n10 commonsourceibias.n8 0.246418
R8557 commonsourceibias.n151 commonsourceibias.n118 0.246418
R8558 commonsourceibias.n330 commonsourceibias.n297 0.246418
R8559 commonsourceibias.n294 commonsourceibias.n292 0.246418
R8560 commonsourceibias.n204 commonsourceibias.n202 0.246418
R8561 commonsourceibias.n240 commonsourceibias.n207 0.246418
R8562 commonsourceibias.n477 commonsourceibias.n444 0.246418
R8563 commonsourceibias.n490 commonsourceibias.n440 0.246418
R8564 commonsourceibias.n536 commonsourceibias.n381 0.246418
R8565 commonsourceibias.n418 commonsourceibias.n385 0.246418
R8566 commonsourceibias.n702 commonsourceibias.n669 0.246418
R8567 commonsourceibias.n715 commonsourceibias.n665 0.246418
R8568 commonsourceibias.n612 commonsourceibias.n579 0.246418
R8569 commonsourceibias.n625 commonsourceibias.n575 0.246418
R8570 commonsourceibias.n95 commonsourceibias.n12 0.189894
R8571 commonsourceibias.n95 commonsourceibias.n94 0.189894
R8572 commonsourceibias.n94 commonsourceibias.n93 0.189894
R8573 commonsourceibias.n93 commonsourceibias.n14 0.189894
R8574 commonsourceibias.n88 commonsourceibias.n14 0.189894
R8575 commonsourceibias.n88 commonsourceibias.n87 0.189894
R8576 commonsourceibias.n87 commonsourceibias.n86 0.189894
R8577 commonsourceibias.n86 commonsourceibias.n16 0.189894
R8578 commonsourceibias.n81 commonsourceibias.n16 0.189894
R8579 commonsourceibias.n81 commonsourceibias.n80 0.189894
R8580 commonsourceibias.n80 commonsourceibias.n79 0.189894
R8581 commonsourceibias.n79 commonsourceibias.n19 0.189894
R8582 commonsourceibias.n74 commonsourceibias.n19 0.189894
R8583 commonsourceibias.n74 commonsourceibias.n73 0.189894
R8584 commonsourceibias.n73 commonsourceibias.n72 0.189894
R8585 commonsourceibias.n72 commonsourceibias.n21 0.189894
R8586 commonsourceibias.n67 commonsourceibias.n21 0.189894
R8587 commonsourceibias.n67 commonsourceibias.n66 0.189894
R8588 commonsourceibias.n66 commonsourceibias.n65 0.189894
R8589 commonsourceibias.n65 commonsourceibias.n24 0.189894
R8590 commonsourceibias.n60 commonsourceibias.n24 0.189894
R8591 commonsourceibias.n60 commonsourceibias.n59 0.189894
R8592 commonsourceibias.n59 commonsourceibias.n26 0.189894
R8593 commonsourceibias.n55 commonsourceibias.n26 0.189894
R8594 commonsourceibias.n55 commonsourceibias.n54 0.189894
R8595 commonsourceibias.n54 commonsourceibias.n28 0.189894
R8596 commonsourceibias.n50 commonsourceibias.n28 0.189894
R8597 commonsourceibias.n50 commonsourceibias.n49 0.189894
R8598 commonsourceibias.n49 commonsourceibias.n30 0.189894
R8599 commonsourceibias.n44 commonsourceibias.n30 0.189894
R8600 commonsourceibias.n44 commonsourceibias.n43 0.189894
R8601 commonsourceibias.n43 commonsourceibias.n42 0.189894
R8602 commonsourceibias.n42 commonsourceibias.n32 0.189894
R8603 commonsourceibias.n37 commonsourceibias.n32 0.189894
R8604 commonsourceibias.n37 commonsourceibias.n36 0.189894
R8605 commonsourceibias.n158 commonsourceibias.n117 0.189894
R8606 commonsourceibias.n153 commonsourceibias.n117 0.189894
R8607 commonsourceibias.n153 commonsourceibias.n152 0.189894
R8608 commonsourceibias.n152 commonsourceibias.n119 0.189894
R8609 commonsourceibias.n148 commonsourceibias.n119 0.189894
R8610 commonsourceibias.n148 commonsourceibias.n147 0.189894
R8611 commonsourceibias.n147 commonsourceibias.n121 0.189894
R8612 commonsourceibias.n143 commonsourceibias.n121 0.189894
R8613 commonsourceibias.n143 commonsourceibias.n142 0.189894
R8614 commonsourceibias.n142 commonsourceibias.n123 0.189894
R8615 commonsourceibias.n137 commonsourceibias.n123 0.189894
R8616 commonsourceibias.n137 commonsourceibias.n136 0.189894
R8617 commonsourceibias.n136 commonsourceibias.n135 0.189894
R8618 commonsourceibias.n135 commonsourceibias.n125 0.189894
R8619 commonsourceibias.n130 commonsourceibias.n125 0.189894
R8620 commonsourceibias.n130 commonsourceibias.n129 0.189894
R8621 commonsourceibias.n188 commonsourceibias.n0 0.189894
R8622 commonsourceibias.n188 commonsourceibias.n187 0.189894
R8623 commonsourceibias.n187 commonsourceibias.n186 0.189894
R8624 commonsourceibias.n186 commonsourceibias.n2 0.189894
R8625 commonsourceibias.n181 commonsourceibias.n2 0.189894
R8626 commonsourceibias.n181 commonsourceibias.n180 0.189894
R8627 commonsourceibias.n180 commonsourceibias.n179 0.189894
R8628 commonsourceibias.n179 commonsourceibias.n4 0.189894
R8629 commonsourceibias.n174 commonsourceibias.n4 0.189894
R8630 commonsourceibias.n174 commonsourceibias.n173 0.189894
R8631 commonsourceibias.n173 commonsourceibias.n172 0.189894
R8632 commonsourceibias.n172 commonsourceibias.n7 0.189894
R8633 commonsourceibias.n167 commonsourceibias.n7 0.189894
R8634 commonsourceibias.n167 commonsourceibias.n166 0.189894
R8635 commonsourceibias.n166 commonsourceibias.n165 0.189894
R8636 commonsourceibias.n165 commonsourceibias.n9 0.189894
R8637 commonsourceibias.n160 commonsourceibias.n9 0.189894
R8638 commonsourceibias.n367 commonsourceibias.n284 0.189894
R8639 commonsourceibias.n367 commonsourceibias.n366 0.189894
R8640 commonsourceibias.n366 commonsourceibias.n365 0.189894
R8641 commonsourceibias.n365 commonsourceibias.n286 0.189894
R8642 commonsourceibias.n360 commonsourceibias.n286 0.189894
R8643 commonsourceibias.n360 commonsourceibias.n359 0.189894
R8644 commonsourceibias.n359 commonsourceibias.n358 0.189894
R8645 commonsourceibias.n358 commonsourceibias.n288 0.189894
R8646 commonsourceibias.n353 commonsourceibias.n288 0.189894
R8647 commonsourceibias.n353 commonsourceibias.n352 0.189894
R8648 commonsourceibias.n352 commonsourceibias.n351 0.189894
R8649 commonsourceibias.n351 commonsourceibias.n291 0.189894
R8650 commonsourceibias.n346 commonsourceibias.n291 0.189894
R8651 commonsourceibias.n346 commonsourceibias.n345 0.189894
R8652 commonsourceibias.n345 commonsourceibias.n344 0.189894
R8653 commonsourceibias.n344 commonsourceibias.n293 0.189894
R8654 commonsourceibias.n339 commonsourceibias.n293 0.189894
R8655 commonsourceibias.n339 commonsourceibias.n338 0.189894
R8656 commonsourceibias.n338 commonsourceibias.n337 0.189894
R8657 commonsourceibias.n337 commonsourceibias.n296 0.189894
R8658 commonsourceibias.n332 commonsourceibias.n296 0.189894
R8659 commonsourceibias.n332 commonsourceibias.n331 0.189894
R8660 commonsourceibias.n331 commonsourceibias.n298 0.189894
R8661 commonsourceibias.n327 commonsourceibias.n298 0.189894
R8662 commonsourceibias.n327 commonsourceibias.n326 0.189894
R8663 commonsourceibias.n326 commonsourceibias.n300 0.189894
R8664 commonsourceibias.n322 commonsourceibias.n300 0.189894
R8665 commonsourceibias.n322 commonsourceibias.n321 0.189894
R8666 commonsourceibias.n321 commonsourceibias.n302 0.189894
R8667 commonsourceibias.n316 commonsourceibias.n302 0.189894
R8668 commonsourceibias.n316 commonsourceibias.n315 0.189894
R8669 commonsourceibias.n315 commonsourceibias.n314 0.189894
R8670 commonsourceibias.n314 commonsourceibias.n304 0.189894
R8671 commonsourceibias.n309 commonsourceibias.n304 0.189894
R8672 commonsourceibias.n309 commonsourceibias.n308 0.189894
R8673 commonsourceibias.n277 commonsourceibias.n194 0.189894
R8674 commonsourceibias.n277 commonsourceibias.n276 0.189894
R8675 commonsourceibias.n276 commonsourceibias.n275 0.189894
R8676 commonsourceibias.n275 commonsourceibias.n196 0.189894
R8677 commonsourceibias.n270 commonsourceibias.n196 0.189894
R8678 commonsourceibias.n270 commonsourceibias.n269 0.189894
R8679 commonsourceibias.n269 commonsourceibias.n268 0.189894
R8680 commonsourceibias.n268 commonsourceibias.n198 0.189894
R8681 commonsourceibias.n263 commonsourceibias.n198 0.189894
R8682 commonsourceibias.n263 commonsourceibias.n262 0.189894
R8683 commonsourceibias.n262 commonsourceibias.n261 0.189894
R8684 commonsourceibias.n261 commonsourceibias.n201 0.189894
R8685 commonsourceibias.n256 commonsourceibias.n201 0.189894
R8686 commonsourceibias.n256 commonsourceibias.n255 0.189894
R8687 commonsourceibias.n255 commonsourceibias.n254 0.189894
R8688 commonsourceibias.n254 commonsourceibias.n203 0.189894
R8689 commonsourceibias.n249 commonsourceibias.n203 0.189894
R8690 commonsourceibias.n249 commonsourceibias.n248 0.189894
R8691 commonsourceibias.n248 commonsourceibias.n247 0.189894
R8692 commonsourceibias.n247 commonsourceibias.n206 0.189894
R8693 commonsourceibias.n242 commonsourceibias.n206 0.189894
R8694 commonsourceibias.n242 commonsourceibias.n241 0.189894
R8695 commonsourceibias.n241 commonsourceibias.n208 0.189894
R8696 commonsourceibias.n237 commonsourceibias.n208 0.189894
R8697 commonsourceibias.n237 commonsourceibias.n236 0.189894
R8698 commonsourceibias.n236 commonsourceibias.n210 0.189894
R8699 commonsourceibias.n232 commonsourceibias.n210 0.189894
R8700 commonsourceibias.n232 commonsourceibias.n231 0.189894
R8701 commonsourceibias.n231 commonsourceibias.n212 0.189894
R8702 commonsourceibias.n226 commonsourceibias.n212 0.189894
R8703 commonsourceibias.n226 commonsourceibias.n225 0.189894
R8704 commonsourceibias.n225 commonsourceibias.n224 0.189894
R8705 commonsourceibias.n224 commonsourceibias.n214 0.189894
R8706 commonsourceibias.n219 commonsourceibias.n214 0.189894
R8707 commonsourceibias.n219 commonsourceibias.n218 0.189894
R8708 commonsourceibias.n456 commonsourceibias.n455 0.189894
R8709 commonsourceibias.n456 commonsourceibias.n451 0.189894
R8710 commonsourceibias.n461 commonsourceibias.n451 0.189894
R8711 commonsourceibias.n462 commonsourceibias.n461 0.189894
R8712 commonsourceibias.n463 commonsourceibias.n462 0.189894
R8713 commonsourceibias.n463 commonsourceibias.n449 0.189894
R8714 commonsourceibias.n468 commonsourceibias.n449 0.189894
R8715 commonsourceibias.n469 commonsourceibias.n468 0.189894
R8716 commonsourceibias.n469 commonsourceibias.n447 0.189894
R8717 commonsourceibias.n473 commonsourceibias.n447 0.189894
R8718 commonsourceibias.n474 commonsourceibias.n473 0.189894
R8719 commonsourceibias.n474 commonsourceibias.n445 0.189894
R8720 commonsourceibias.n478 commonsourceibias.n445 0.189894
R8721 commonsourceibias.n479 commonsourceibias.n478 0.189894
R8722 commonsourceibias.n479 commonsourceibias.n443 0.189894
R8723 commonsourceibias.n484 commonsourceibias.n443 0.189894
R8724 commonsourceibias.n485 commonsourceibias.n484 0.189894
R8725 commonsourceibias.n486 commonsourceibias.n485 0.189894
R8726 commonsourceibias.n486 commonsourceibias.n441 0.189894
R8727 commonsourceibias.n492 commonsourceibias.n441 0.189894
R8728 commonsourceibias.n493 commonsourceibias.n492 0.189894
R8729 commonsourceibias.n494 commonsourceibias.n493 0.189894
R8730 commonsourceibias.n494 commonsourceibias.n439 0.189894
R8731 commonsourceibias.n499 commonsourceibias.n439 0.189894
R8732 commonsourceibias.n500 commonsourceibias.n499 0.189894
R8733 commonsourceibias.n501 commonsourceibias.n500 0.189894
R8734 commonsourceibias.n501 commonsourceibias.n437 0.189894
R8735 commonsourceibias.n507 commonsourceibias.n437 0.189894
R8736 commonsourceibias.n508 commonsourceibias.n507 0.189894
R8737 commonsourceibias.n509 commonsourceibias.n508 0.189894
R8738 commonsourceibias.n509 commonsourceibias.n435 0.189894
R8739 commonsourceibias.n514 commonsourceibias.n435 0.189894
R8740 commonsourceibias.n515 commonsourceibias.n514 0.189894
R8741 commonsourceibias.n516 commonsourceibias.n515 0.189894
R8742 commonsourceibias.n516 commonsourceibias.n433 0.189894
R8743 commonsourceibias.n397 commonsourceibias.n396 0.189894
R8744 commonsourceibias.n397 commonsourceibias.n392 0.189894
R8745 commonsourceibias.n402 commonsourceibias.n392 0.189894
R8746 commonsourceibias.n403 commonsourceibias.n402 0.189894
R8747 commonsourceibias.n404 commonsourceibias.n403 0.189894
R8748 commonsourceibias.n404 commonsourceibias.n390 0.189894
R8749 commonsourceibias.n409 commonsourceibias.n390 0.189894
R8750 commonsourceibias.n410 commonsourceibias.n409 0.189894
R8751 commonsourceibias.n410 commonsourceibias.n388 0.189894
R8752 commonsourceibias.n414 commonsourceibias.n388 0.189894
R8753 commonsourceibias.n415 commonsourceibias.n414 0.189894
R8754 commonsourceibias.n415 commonsourceibias.n386 0.189894
R8755 commonsourceibias.n419 commonsourceibias.n386 0.189894
R8756 commonsourceibias.n420 commonsourceibias.n419 0.189894
R8757 commonsourceibias.n420 commonsourceibias.n384 0.189894
R8758 commonsourceibias.n425 commonsourceibias.n384 0.189894
R8759 commonsourceibias.n532 commonsourceibias.n382 0.189894
R8760 commonsourceibias.n538 commonsourceibias.n382 0.189894
R8761 commonsourceibias.n539 commonsourceibias.n538 0.189894
R8762 commonsourceibias.n540 commonsourceibias.n539 0.189894
R8763 commonsourceibias.n540 commonsourceibias.n380 0.189894
R8764 commonsourceibias.n545 commonsourceibias.n380 0.189894
R8765 commonsourceibias.n546 commonsourceibias.n545 0.189894
R8766 commonsourceibias.n547 commonsourceibias.n546 0.189894
R8767 commonsourceibias.n547 commonsourceibias.n378 0.189894
R8768 commonsourceibias.n553 commonsourceibias.n378 0.189894
R8769 commonsourceibias.n554 commonsourceibias.n553 0.189894
R8770 commonsourceibias.n555 commonsourceibias.n554 0.189894
R8771 commonsourceibias.n555 commonsourceibias.n376 0.189894
R8772 commonsourceibias.n560 commonsourceibias.n376 0.189894
R8773 commonsourceibias.n561 commonsourceibias.n560 0.189894
R8774 commonsourceibias.n562 commonsourceibias.n561 0.189894
R8775 commonsourceibias.n562 commonsourceibias.n374 0.189894
R8776 commonsourceibias.n681 commonsourceibias.n680 0.189894
R8777 commonsourceibias.n681 commonsourceibias.n676 0.189894
R8778 commonsourceibias.n686 commonsourceibias.n676 0.189894
R8779 commonsourceibias.n687 commonsourceibias.n686 0.189894
R8780 commonsourceibias.n688 commonsourceibias.n687 0.189894
R8781 commonsourceibias.n688 commonsourceibias.n674 0.189894
R8782 commonsourceibias.n693 commonsourceibias.n674 0.189894
R8783 commonsourceibias.n694 commonsourceibias.n693 0.189894
R8784 commonsourceibias.n694 commonsourceibias.n672 0.189894
R8785 commonsourceibias.n698 commonsourceibias.n672 0.189894
R8786 commonsourceibias.n699 commonsourceibias.n698 0.189894
R8787 commonsourceibias.n699 commonsourceibias.n670 0.189894
R8788 commonsourceibias.n703 commonsourceibias.n670 0.189894
R8789 commonsourceibias.n704 commonsourceibias.n703 0.189894
R8790 commonsourceibias.n704 commonsourceibias.n668 0.189894
R8791 commonsourceibias.n709 commonsourceibias.n668 0.189894
R8792 commonsourceibias.n710 commonsourceibias.n709 0.189894
R8793 commonsourceibias.n711 commonsourceibias.n710 0.189894
R8794 commonsourceibias.n711 commonsourceibias.n666 0.189894
R8795 commonsourceibias.n717 commonsourceibias.n666 0.189894
R8796 commonsourceibias.n718 commonsourceibias.n717 0.189894
R8797 commonsourceibias.n719 commonsourceibias.n718 0.189894
R8798 commonsourceibias.n719 commonsourceibias.n664 0.189894
R8799 commonsourceibias.n724 commonsourceibias.n664 0.189894
R8800 commonsourceibias.n725 commonsourceibias.n724 0.189894
R8801 commonsourceibias.n726 commonsourceibias.n725 0.189894
R8802 commonsourceibias.n726 commonsourceibias.n662 0.189894
R8803 commonsourceibias.n732 commonsourceibias.n662 0.189894
R8804 commonsourceibias.n733 commonsourceibias.n732 0.189894
R8805 commonsourceibias.n734 commonsourceibias.n733 0.189894
R8806 commonsourceibias.n734 commonsourceibias.n660 0.189894
R8807 commonsourceibias.n739 commonsourceibias.n660 0.189894
R8808 commonsourceibias.n740 commonsourceibias.n739 0.189894
R8809 commonsourceibias.n741 commonsourceibias.n740 0.189894
R8810 commonsourceibias.n741 commonsourceibias.n658 0.189894
R8811 commonsourceibias.n591 commonsourceibias.n590 0.189894
R8812 commonsourceibias.n591 commonsourceibias.n586 0.189894
R8813 commonsourceibias.n596 commonsourceibias.n586 0.189894
R8814 commonsourceibias.n597 commonsourceibias.n596 0.189894
R8815 commonsourceibias.n598 commonsourceibias.n597 0.189894
R8816 commonsourceibias.n598 commonsourceibias.n584 0.189894
R8817 commonsourceibias.n603 commonsourceibias.n584 0.189894
R8818 commonsourceibias.n604 commonsourceibias.n603 0.189894
R8819 commonsourceibias.n604 commonsourceibias.n582 0.189894
R8820 commonsourceibias.n608 commonsourceibias.n582 0.189894
R8821 commonsourceibias.n609 commonsourceibias.n608 0.189894
R8822 commonsourceibias.n609 commonsourceibias.n580 0.189894
R8823 commonsourceibias.n613 commonsourceibias.n580 0.189894
R8824 commonsourceibias.n614 commonsourceibias.n613 0.189894
R8825 commonsourceibias.n614 commonsourceibias.n578 0.189894
R8826 commonsourceibias.n619 commonsourceibias.n578 0.189894
R8827 commonsourceibias.n620 commonsourceibias.n619 0.189894
R8828 commonsourceibias.n621 commonsourceibias.n620 0.189894
R8829 commonsourceibias.n621 commonsourceibias.n576 0.189894
R8830 commonsourceibias.n627 commonsourceibias.n576 0.189894
R8831 commonsourceibias.n628 commonsourceibias.n627 0.189894
R8832 commonsourceibias.n629 commonsourceibias.n628 0.189894
R8833 commonsourceibias.n629 commonsourceibias.n574 0.189894
R8834 commonsourceibias.n634 commonsourceibias.n574 0.189894
R8835 commonsourceibias.n635 commonsourceibias.n634 0.189894
R8836 commonsourceibias.n636 commonsourceibias.n635 0.189894
R8837 commonsourceibias.n636 commonsourceibias.n572 0.189894
R8838 commonsourceibias.n642 commonsourceibias.n572 0.189894
R8839 commonsourceibias.n643 commonsourceibias.n642 0.189894
R8840 commonsourceibias.n644 commonsourceibias.n643 0.189894
R8841 commonsourceibias.n644 commonsourceibias.n570 0.189894
R8842 commonsourceibias.n649 commonsourceibias.n570 0.189894
R8843 commonsourceibias.n650 commonsourceibias.n649 0.189894
R8844 commonsourceibias.n651 commonsourceibias.n650 0.189894
R8845 commonsourceibias.n651 commonsourceibias.n568 0.189894
R8846 commonsourceibias.n159 commonsourceibias.n158 0.170955
R8847 commonsourceibias.n160 commonsourceibias.n159 0.170955
R8848 commonsourceibias.n531 commonsourceibias.n425 0.170955
R8849 commonsourceibias.n532 commonsourceibias.n531 0.170955
R8850 gnd.n7072 gnd.n514 1183.27
R8851 gnd.n4441 gnd.n4127 939.716
R8852 gnd.n7550 gnd.n208 795.207
R8853 gnd.n348 gnd.n211 795.207
R8854 gnd.n1576 gnd.n1464 795.207
R8855 gnd.n5958 gnd.n1578 795.207
R8856 gnd.n6411 gnd.n1064 795.207
R8857 gnd.n4794 gnd.n1067 795.207
R8858 gnd.n4281 gnd.n4164 795.207
R8859 gnd.n4320 gnd.n2639 795.207
R8860 gnd.n4035 gnd.n2650 766.379
R8861 gnd.n4038 gnd.n4037 766.379
R8862 gnd.n3276 gnd.n3179 766.379
R8863 gnd.n3272 gnd.n3177 766.379
R8864 gnd.n4126 gnd.n2672 756.769
R8865 gnd.n4029 gnd.n4028 756.769
R8866 gnd.n3369 gnd.n3086 756.769
R8867 gnd.n3367 gnd.n3089 756.769
R8868 gnd.n6653 gnd.n767 756.769
R8869 gnd.n7073 gnd.n515 756.769
R8870 gnd.n7286 gnd.n388 756.769
R8871 gnd.n6485 gnd.n937 756.769
R8872 gnd.n7548 gnd.n213 739.952
R8873 gnd.n7439 gnd.n210 739.952
R8874 gnd.n5961 gnd.n5960 739.952
R8875 gnd.n6078 gnd.n1510 739.952
R8876 gnd.n6409 gnd.n1069 739.952
R8877 gnd.n2386 gnd.n1066 739.952
R8878 gnd.n4444 gnd.n4443 739.952
R8879 gnd.n4439 gnd.n2635 739.952
R8880 gnd.n4855 gnd.n2196 711.122
R8881 gnd.n6147 gnd.n1400 711.122
R8882 gnd.n4867 gnd.n2194 711.122
R8883 gnd.n6149 gnd.n1395 711.122
R8884 gnd.n6654 gnd.n6653 585
R8885 gnd.n6653 gnd.n6652 585
R8886 gnd.n771 gnd.n770 585
R8887 gnd.n6651 gnd.n771 585
R8888 gnd.n6649 gnd.n6648 585
R8889 gnd.n6650 gnd.n6649 585
R8890 gnd.n6647 gnd.n773 585
R8891 gnd.n773 gnd.n772 585
R8892 gnd.n6646 gnd.n6645 585
R8893 gnd.n6645 gnd.n6644 585
R8894 gnd.n778 gnd.n777 585
R8895 gnd.n6643 gnd.n778 585
R8896 gnd.n6641 gnd.n6640 585
R8897 gnd.n6642 gnd.n6641 585
R8898 gnd.n6639 gnd.n780 585
R8899 gnd.n780 gnd.n779 585
R8900 gnd.n6638 gnd.n6637 585
R8901 gnd.n6637 gnd.n6636 585
R8902 gnd.n786 gnd.n785 585
R8903 gnd.n6635 gnd.n786 585
R8904 gnd.n6633 gnd.n6632 585
R8905 gnd.n6634 gnd.n6633 585
R8906 gnd.n6631 gnd.n788 585
R8907 gnd.n788 gnd.n787 585
R8908 gnd.n6630 gnd.n6629 585
R8909 gnd.n6629 gnd.n6628 585
R8910 gnd.n794 gnd.n793 585
R8911 gnd.n6627 gnd.n794 585
R8912 gnd.n6625 gnd.n6624 585
R8913 gnd.n6626 gnd.n6625 585
R8914 gnd.n6623 gnd.n796 585
R8915 gnd.n796 gnd.n795 585
R8916 gnd.n6622 gnd.n6621 585
R8917 gnd.n6621 gnd.n6620 585
R8918 gnd.n802 gnd.n801 585
R8919 gnd.n6619 gnd.n802 585
R8920 gnd.n6617 gnd.n6616 585
R8921 gnd.n6618 gnd.n6617 585
R8922 gnd.n6615 gnd.n804 585
R8923 gnd.n804 gnd.n803 585
R8924 gnd.n6614 gnd.n6613 585
R8925 gnd.n6613 gnd.n6612 585
R8926 gnd.n810 gnd.n809 585
R8927 gnd.n6611 gnd.n810 585
R8928 gnd.n6609 gnd.n6608 585
R8929 gnd.n6610 gnd.n6609 585
R8930 gnd.n6607 gnd.n812 585
R8931 gnd.n812 gnd.n811 585
R8932 gnd.n6606 gnd.n6605 585
R8933 gnd.n6605 gnd.n6604 585
R8934 gnd.n818 gnd.n817 585
R8935 gnd.n6603 gnd.n818 585
R8936 gnd.n6601 gnd.n6600 585
R8937 gnd.n6602 gnd.n6601 585
R8938 gnd.n6599 gnd.n820 585
R8939 gnd.n820 gnd.n819 585
R8940 gnd.n6598 gnd.n6597 585
R8941 gnd.n6597 gnd.n6596 585
R8942 gnd.n826 gnd.n825 585
R8943 gnd.n6595 gnd.n826 585
R8944 gnd.n6593 gnd.n6592 585
R8945 gnd.n6594 gnd.n6593 585
R8946 gnd.n6591 gnd.n828 585
R8947 gnd.n828 gnd.n827 585
R8948 gnd.n6590 gnd.n6589 585
R8949 gnd.n6589 gnd.n6588 585
R8950 gnd.n834 gnd.n833 585
R8951 gnd.n6587 gnd.n834 585
R8952 gnd.n6585 gnd.n6584 585
R8953 gnd.n6586 gnd.n6585 585
R8954 gnd.n6583 gnd.n836 585
R8955 gnd.n836 gnd.n835 585
R8956 gnd.n6582 gnd.n6581 585
R8957 gnd.n6581 gnd.n6580 585
R8958 gnd.n842 gnd.n841 585
R8959 gnd.n6579 gnd.n842 585
R8960 gnd.n6577 gnd.n6576 585
R8961 gnd.n6578 gnd.n6577 585
R8962 gnd.n6575 gnd.n844 585
R8963 gnd.n844 gnd.n843 585
R8964 gnd.n6574 gnd.n6573 585
R8965 gnd.n6573 gnd.n6572 585
R8966 gnd.n850 gnd.n849 585
R8967 gnd.n6571 gnd.n850 585
R8968 gnd.n6569 gnd.n6568 585
R8969 gnd.n6570 gnd.n6569 585
R8970 gnd.n6567 gnd.n852 585
R8971 gnd.n852 gnd.n851 585
R8972 gnd.n6566 gnd.n6565 585
R8973 gnd.n6565 gnd.n6564 585
R8974 gnd.n858 gnd.n857 585
R8975 gnd.n6563 gnd.n858 585
R8976 gnd.n6561 gnd.n6560 585
R8977 gnd.n6562 gnd.n6561 585
R8978 gnd.n6559 gnd.n860 585
R8979 gnd.n860 gnd.n859 585
R8980 gnd.n6558 gnd.n6557 585
R8981 gnd.n6557 gnd.n6556 585
R8982 gnd.n866 gnd.n865 585
R8983 gnd.n6555 gnd.n866 585
R8984 gnd.n6553 gnd.n6552 585
R8985 gnd.n6554 gnd.n6553 585
R8986 gnd.n6551 gnd.n868 585
R8987 gnd.n868 gnd.n867 585
R8988 gnd.n6550 gnd.n6549 585
R8989 gnd.n6549 gnd.n6548 585
R8990 gnd.n874 gnd.n873 585
R8991 gnd.n6547 gnd.n874 585
R8992 gnd.n6545 gnd.n6544 585
R8993 gnd.n6546 gnd.n6545 585
R8994 gnd.n6543 gnd.n876 585
R8995 gnd.n876 gnd.n875 585
R8996 gnd.n6542 gnd.n6541 585
R8997 gnd.n6541 gnd.n6540 585
R8998 gnd.n882 gnd.n881 585
R8999 gnd.n6539 gnd.n882 585
R9000 gnd.n6537 gnd.n6536 585
R9001 gnd.n6538 gnd.n6537 585
R9002 gnd.n6535 gnd.n884 585
R9003 gnd.n884 gnd.n883 585
R9004 gnd.n6534 gnd.n6533 585
R9005 gnd.n6533 gnd.n6532 585
R9006 gnd.n890 gnd.n889 585
R9007 gnd.n6531 gnd.n890 585
R9008 gnd.n6529 gnd.n6528 585
R9009 gnd.n6530 gnd.n6529 585
R9010 gnd.n6527 gnd.n892 585
R9011 gnd.n892 gnd.n891 585
R9012 gnd.n6526 gnd.n6525 585
R9013 gnd.n6525 gnd.n6524 585
R9014 gnd.n898 gnd.n897 585
R9015 gnd.n6523 gnd.n898 585
R9016 gnd.n6521 gnd.n6520 585
R9017 gnd.n6522 gnd.n6521 585
R9018 gnd.n6519 gnd.n900 585
R9019 gnd.n900 gnd.n899 585
R9020 gnd.n6518 gnd.n6517 585
R9021 gnd.n6517 gnd.n6516 585
R9022 gnd.n906 gnd.n905 585
R9023 gnd.n6515 gnd.n906 585
R9024 gnd.n6513 gnd.n6512 585
R9025 gnd.n6514 gnd.n6513 585
R9026 gnd.n6511 gnd.n908 585
R9027 gnd.n908 gnd.n907 585
R9028 gnd.n6510 gnd.n6509 585
R9029 gnd.n6509 gnd.n6508 585
R9030 gnd.n914 gnd.n913 585
R9031 gnd.n6507 gnd.n914 585
R9032 gnd.n6505 gnd.n6504 585
R9033 gnd.n6506 gnd.n6505 585
R9034 gnd.n6503 gnd.n916 585
R9035 gnd.n916 gnd.n915 585
R9036 gnd.n6502 gnd.n6501 585
R9037 gnd.n6501 gnd.n6500 585
R9038 gnd.n922 gnd.n921 585
R9039 gnd.n6499 gnd.n922 585
R9040 gnd.n6497 gnd.n6496 585
R9041 gnd.n6498 gnd.n6497 585
R9042 gnd.n6495 gnd.n924 585
R9043 gnd.n924 gnd.n923 585
R9044 gnd.n6494 gnd.n6493 585
R9045 gnd.n6493 gnd.n6492 585
R9046 gnd.n930 gnd.n929 585
R9047 gnd.n6491 gnd.n930 585
R9048 gnd.n6489 gnd.n6488 585
R9049 gnd.n6490 gnd.n6489 585
R9050 gnd.n6487 gnd.n932 585
R9051 gnd.n932 gnd.n931 585
R9052 gnd.n768 gnd.n767 585
R9053 gnd.n767 gnd.n766 585
R9054 gnd.n6659 gnd.n6658 585
R9055 gnd.n6660 gnd.n6659 585
R9056 gnd.n765 gnd.n764 585
R9057 gnd.n6661 gnd.n765 585
R9058 gnd.n6664 gnd.n6663 585
R9059 gnd.n6663 gnd.n6662 585
R9060 gnd.n762 gnd.n761 585
R9061 gnd.n761 gnd.n760 585
R9062 gnd.n6669 gnd.n6668 585
R9063 gnd.n6670 gnd.n6669 585
R9064 gnd.n759 gnd.n758 585
R9065 gnd.n6671 gnd.n759 585
R9066 gnd.n6674 gnd.n6673 585
R9067 gnd.n6673 gnd.n6672 585
R9068 gnd.n756 gnd.n755 585
R9069 gnd.n755 gnd.n754 585
R9070 gnd.n6679 gnd.n6678 585
R9071 gnd.n6680 gnd.n6679 585
R9072 gnd.n753 gnd.n752 585
R9073 gnd.n6681 gnd.n753 585
R9074 gnd.n6684 gnd.n6683 585
R9075 gnd.n6683 gnd.n6682 585
R9076 gnd.n750 gnd.n749 585
R9077 gnd.n749 gnd.n748 585
R9078 gnd.n6689 gnd.n6688 585
R9079 gnd.n6690 gnd.n6689 585
R9080 gnd.n747 gnd.n746 585
R9081 gnd.n6691 gnd.n747 585
R9082 gnd.n6694 gnd.n6693 585
R9083 gnd.n6693 gnd.n6692 585
R9084 gnd.n744 gnd.n743 585
R9085 gnd.n743 gnd.n742 585
R9086 gnd.n6699 gnd.n6698 585
R9087 gnd.n6700 gnd.n6699 585
R9088 gnd.n741 gnd.n740 585
R9089 gnd.n6701 gnd.n741 585
R9090 gnd.n6704 gnd.n6703 585
R9091 gnd.n6703 gnd.n6702 585
R9092 gnd.n738 gnd.n737 585
R9093 gnd.n737 gnd.n736 585
R9094 gnd.n6709 gnd.n6708 585
R9095 gnd.n6710 gnd.n6709 585
R9096 gnd.n735 gnd.n734 585
R9097 gnd.n6711 gnd.n735 585
R9098 gnd.n6714 gnd.n6713 585
R9099 gnd.n6713 gnd.n6712 585
R9100 gnd.n732 gnd.n731 585
R9101 gnd.n731 gnd.n730 585
R9102 gnd.n6719 gnd.n6718 585
R9103 gnd.n6720 gnd.n6719 585
R9104 gnd.n729 gnd.n728 585
R9105 gnd.n6721 gnd.n729 585
R9106 gnd.n6724 gnd.n6723 585
R9107 gnd.n6723 gnd.n6722 585
R9108 gnd.n726 gnd.n725 585
R9109 gnd.n725 gnd.n724 585
R9110 gnd.n6729 gnd.n6728 585
R9111 gnd.n6730 gnd.n6729 585
R9112 gnd.n723 gnd.n722 585
R9113 gnd.n6731 gnd.n723 585
R9114 gnd.n6734 gnd.n6733 585
R9115 gnd.n6733 gnd.n6732 585
R9116 gnd.n720 gnd.n719 585
R9117 gnd.n719 gnd.n718 585
R9118 gnd.n6739 gnd.n6738 585
R9119 gnd.n6740 gnd.n6739 585
R9120 gnd.n717 gnd.n716 585
R9121 gnd.n6741 gnd.n717 585
R9122 gnd.n6744 gnd.n6743 585
R9123 gnd.n6743 gnd.n6742 585
R9124 gnd.n714 gnd.n713 585
R9125 gnd.n713 gnd.n712 585
R9126 gnd.n6749 gnd.n6748 585
R9127 gnd.n6750 gnd.n6749 585
R9128 gnd.n711 gnd.n710 585
R9129 gnd.n6751 gnd.n711 585
R9130 gnd.n6754 gnd.n6753 585
R9131 gnd.n6753 gnd.n6752 585
R9132 gnd.n708 gnd.n707 585
R9133 gnd.n707 gnd.n706 585
R9134 gnd.n6759 gnd.n6758 585
R9135 gnd.n6760 gnd.n6759 585
R9136 gnd.n705 gnd.n704 585
R9137 gnd.n6761 gnd.n705 585
R9138 gnd.n6764 gnd.n6763 585
R9139 gnd.n6763 gnd.n6762 585
R9140 gnd.n702 gnd.n701 585
R9141 gnd.n701 gnd.n700 585
R9142 gnd.n6769 gnd.n6768 585
R9143 gnd.n6770 gnd.n6769 585
R9144 gnd.n699 gnd.n698 585
R9145 gnd.n6771 gnd.n699 585
R9146 gnd.n6774 gnd.n6773 585
R9147 gnd.n6773 gnd.n6772 585
R9148 gnd.n696 gnd.n695 585
R9149 gnd.n695 gnd.n694 585
R9150 gnd.n6779 gnd.n6778 585
R9151 gnd.n6780 gnd.n6779 585
R9152 gnd.n693 gnd.n692 585
R9153 gnd.n6781 gnd.n693 585
R9154 gnd.n6784 gnd.n6783 585
R9155 gnd.n6783 gnd.n6782 585
R9156 gnd.n690 gnd.n689 585
R9157 gnd.n689 gnd.n688 585
R9158 gnd.n6789 gnd.n6788 585
R9159 gnd.n6790 gnd.n6789 585
R9160 gnd.n687 gnd.n686 585
R9161 gnd.n6791 gnd.n687 585
R9162 gnd.n6794 gnd.n6793 585
R9163 gnd.n6793 gnd.n6792 585
R9164 gnd.n684 gnd.n683 585
R9165 gnd.n683 gnd.n682 585
R9166 gnd.n6799 gnd.n6798 585
R9167 gnd.n6800 gnd.n6799 585
R9168 gnd.n681 gnd.n680 585
R9169 gnd.n6801 gnd.n681 585
R9170 gnd.n6804 gnd.n6803 585
R9171 gnd.n6803 gnd.n6802 585
R9172 gnd.n678 gnd.n677 585
R9173 gnd.n677 gnd.n676 585
R9174 gnd.n6809 gnd.n6808 585
R9175 gnd.n6810 gnd.n6809 585
R9176 gnd.n675 gnd.n674 585
R9177 gnd.n6811 gnd.n675 585
R9178 gnd.n6814 gnd.n6813 585
R9179 gnd.n6813 gnd.n6812 585
R9180 gnd.n672 gnd.n671 585
R9181 gnd.n671 gnd.n670 585
R9182 gnd.n6819 gnd.n6818 585
R9183 gnd.n6820 gnd.n6819 585
R9184 gnd.n669 gnd.n668 585
R9185 gnd.n6821 gnd.n669 585
R9186 gnd.n6824 gnd.n6823 585
R9187 gnd.n6823 gnd.n6822 585
R9188 gnd.n666 gnd.n665 585
R9189 gnd.n665 gnd.n664 585
R9190 gnd.n6829 gnd.n6828 585
R9191 gnd.n6830 gnd.n6829 585
R9192 gnd.n663 gnd.n662 585
R9193 gnd.n6831 gnd.n663 585
R9194 gnd.n6834 gnd.n6833 585
R9195 gnd.n6833 gnd.n6832 585
R9196 gnd.n660 gnd.n659 585
R9197 gnd.n659 gnd.n658 585
R9198 gnd.n6839 gnd.n6838 585
R9199 gnd.n6840 gnd.n6839 585
R9200 gnd.n657 gnd.n656 585
R9201 gnd.n6841 gnd.n657 585
R9202 gnd.n6844 gnd.n6843 585
R9203 gnd.n6843 gnd.n6842 585
R9204 gnd.n654 gnd.n653 585
R9205 gnd.n653 gnd.n652 585
R9206 gnd.n6849 gnd.n6848 585
R9207 gnd.n6850 gnd.n6849 585
R9208 gnd.n651 gnd.n650 585
R9209 gnd.n6851 gnd.n651 585
R9210 gnd.n6854 gnd.n6853 585
R9211 gnd.n6853 gnd.n6852 585
R9212 gnd.n648 gnd.n647 585
R9213 gnd.n647 gnd.n646 585
R9214 gnd.n6859 gnd.n6858 585
R9215 gnd.n6860 gnd.n6859 585
R9216 gnd.n645 gnd.n644 585
R9217 gnd.n6861 gnd.n645 585
R9218 gnd.n6864 gnd.n6863 585
R9219 gnd.n6863 gnd.n6862 585
R9220 gnd.n642 gnd.n641 585
R9221 gnd.n641 gnd.n640 585
R9222 gnd.n6869 gnd.n6868 585
R9223 gnd.n6870 gnd.n6869 585
R9224 gnd.n639 gnd.n638 585
R9225 gnd.n6871 gnd.n639 585
R9226 gnd.n6874 gnd.n6873 585
R9227 gnd.n6873 gnd.n6872 585
R9228 gnd.n636 gnd.n635 585
R9229 gnd.n635 gnd.n634 585
R9230 gnd.n6879 gnd.n6878 585
R9231 gnd.n6880 gnd.n6879 585
R9232 gnd.n633 gnd.n632 585
R9233 gnd.n6881 gnd.n633 585
R9234 gnd.n6884 gnd.n6883 585
R9235 gnd.n6883 gnd.n6882 585
R9236 gnd.n630 gnd.n629 585
R9237 gnd.n629 gnd.n628 585
R9238 gnd.n6889 gnd.n6888 585
R9239 gnd.n6890 gnd.n6889 585
R9240 gnd.n627 gnd.n626 585
R9241 gnd.n6891 gnd.n627 585
R9242 gnd.n6894 gnd.n6893 585
R9243 gnd.n6893 gnd.n6892 585
R9244 gnd.n624 gnd.n623 585
R9245 gnd.n623 gnd.n622 585
R9246 gnd.n6899 gnd.n6898 585
R9247 gnd.n6900 gnd.n6899 585
R9248 gnd.n621 gnd.n620 585
R9249 gnd.n6901 gnd.n621 585
R9250 gnd.n6904 gnd.n6903 585
R9251 gnd.n6903 gnd.n6902 585
R9252 gnd.n618 gnd.n617 585
R9253 gnd.n617 gnd.n616 585
R9254 gnd.n6909 gnd.n6908 585
R9255 gnd.n6910 gnd.n6909 585
R9256 gnd.n615 gnd.n614 585
R9257 gnd.n6911 gnd.n615 585
R9258 gnd.n6914 gnd.n6913 585
R9259 gnd.n6913 gnd.n6912 585
R9260 gnd.n612 gnd.n611 585
R9261 gnd.n611 gnd.n610 585
R9262 gnd.n6919 gnd.n6918 585
R9263 gnd.n6920 gnd.n6919 585
R9264 gnd.n609 gnd.n608 585
R9265 gnd.n6921 gnd.n609 585
R9266 gnd.n6924 gnd.n6923 585
R9267 gnd.n6923 gnd.n6922 585
R9268 gnd.n606 gnd.n605 585
R9269 gnd.n605 gnd.n604 585
R9270 gnd.n6929 gnd.n6928 585
R9271 gnd.n6930 gnd.n6929 585
R9272 gnd.n603 gnd.n602 585
R9273 gnd.n6931 gnd.n603 585
R9274 gnd.n6934 gnd.n6933 585
R9275 gnd.n6933 gnd.n6932 585
R9276 gnd.n600 gnd.n599 585
R9277 gnd.n599 gnd.n598 585
R9278 gnd.n6939 gnd.n6938 585
R9279 gnd.n6940 gnd.n6939 585
R9280 gnd.n597 gnd.n596 585
R9281 gnd.n6941 gnd.n597 585
R9282 gnd.n6944 gnd.n6943 585
R9283 gnd.n6943 gnd.n6942 585
R9284 gnd.n594 gnd.n593 585
R9285 gnd.n593 gnd.n592 585
R9286 gnd.n6949 gnd.n6948 585
R9287 gnd.n6950 gnd.n6949 585
R9288 gnd.n591 gnd.n590 585
R9289 gnd.n6951 gnd.n591 585
R9290 gnd.n6954 gnd.n6953 585
R9291 gnd.n6953 gnd.n6952 585
R9292 gnd.n588 gnd.n587 585
R9293 gnd.n587 gnd.n586 585
R9294 gnd.n6959 gnd.n6958 585
R9295 gnd.n6960 gnd.n6959 585
R9296 gnd.n585 gnd.n584 585
R9297 gnd.n6961 gnd.n585 585
R9298 gnd.n6964 gnd.n6963 585
R9299 gnd.n6963 gnd.n6962 585
R9300 gnd.n582 gnd.n581 585
R9301 gnd.n581 gnd.n580 585
R9302 gnd.n6969 gnd.n6968 585
R9303 gnd.n6970 gnd.n6969 585
R9304 gnd.n579 gnd.n578 585
R9305 gnd.n6971 gnd.n579 585
R9306 gnd.n6974 gnd.n6973 585
R9307 gnd.n6973 gnd.n6972 585
R9308 gnd.n576 gnd.n575 585
R9309 gnd.n575 gnd.n574 585
R9310 gnd.n6979 gnd.n6978 585
R9311 gnd.n6980 gnd.n6979 585
R9312 gnd.n573 gnd.n572 585
R9313 gnd.n6981 gnd.n573 585
R9314 gnd.n6984 gnd.n6983 585
R9315 gnd.n6983 gnd.n6982 585
R9316 gnd.n570 gnd.n569 585
R9317 gnd.n569 gnd.n568 585
R9318 gnd.n6989 gnd.n6988 585
R9319 gnd.n6990 gnd.n6989 585
R9320 gnd.n567 gnd.n566 585
R9321 gnd.n6991 gnd.n567 585
R9322 gnd.n6994 gnd.n6993 585
R9323 gnd.n6993 gnd.n6992 585
R9324 gnd.n564 gnd.n563 585
R9325 gnd.n563 gnd.n562 585
R9326 gnd.n6999 gnd.n6998 585
R9327 gnd.n7000 gnd.n6999 585
R9328 gnd.n561 gnd.n560 585
R9329 gnd.n7001 gnd.n561 585
R9330 gnd.n7004 gnd.n7003 585
R9331 gnd.n7003 gnd.n7002 585
R9332 gnd.n558 gnd.n557 585
R9333 gnd.n557 gnd.n556 585
R9334 gnd.n7009 gnd.n7008 585
R9335 gnd.n7010 gnd.n7009 585
R9336 gnd.n555 gnd.n554 585
R9337 gnd.n7011 gnd.n555 585
R9338 gnd.n7014 gnd.n7013 585
R9339 gnd.n7013 gnd.n7012 585
R9340 gnd.n552 gnd.n551 585
R9341 gnd.n551 gnd.n550 585
R9342 gnd.n7019 gnd.n7018 585
R9343 gnd.n7020 gnd.n7019 585
R9344 gnd.n549 gnd.n548 585
R9345 gnd.n7021 gnd.n549 585
R9346 gnd.n7024 gnd.n7023 585
R9347 gnd.n7023 gnd.n7022 585
R9348 gnd.n546 gnd.n545 585
R9349 gnd.n545 gnd.n544 585
R9350 gnd.n7029 gnd.n7028 585
R9351 gnd.n7030 gnd.n7029 585
R9352 gnd.n543 gnd.n542 585
R9353 gnd.n7031 gnd.n543 585
R9354 gnd.n7034 gnd.n7033 585
R9355 gnd.n7033 gnd.n7032 585
R9356 gnd.n540 gnd.n539 585
R9357 gnd.n539 gnd.n538 585
R9358 gnd.n7039 gnd.n7038 585
R9359 gnd.n7040 gnd.n7039 585
R9360 gnd.n537 gnd.n536 585
R9361 gnd.n7041 gnd.n537 585
R9362 gnd.n7044 gnd.n7043 585
R9363 gnd.n7043 gnd.n7042 585
R9364 gnd.n534 gnd.n533 585
R9365 gnd.n533 gnd.n532 585
R9366 gnd.n7049 gnd.n7048 585
R9367 gnd.n7050 gnd.n7049 585
R9368 gnd.n531 gnd.n530 585
R9369 gnd.n7051 gnd.n531 585
R9370 gnd.n7054 gnd.n7053 585
R9371 gnd.n7053 gnd.n7052 585
R9372 gnd.n528 gnd.n527 585
R9373 gnd.n527 gnd.n526 585
R9374 gnd.n7059 gnd.n7058 585
R9375 gnd.n7060 gnd.n7059 585
R9376 gnd.n525 gnd.n524 585
R9377 gnd.n7061 gnd.n525 585
R9378 gnd.n7064 gnd.n7063 585
R9379 gnd.n7063 gnd.n7062 585
R9380 gnd.n522 gnd.n521 585
R9381 gnd.n521 gnd.n520 585
R9382 gnd.n7069 gnd.n7068 585
R9383 gnd.n7070 gnd.n7069 585
R9384 gnd.n519 gnd.n518 585
R9385 gnd.n7071 gnd.n519 585
R9386 gnd.n7074 gnd.n7073 585
R9387 gnd.n7073 gnd.n7072 585
R9388 gnd.n7285 gnd.n392 585
R9389 gnd.n7285 gnd.n7284 585
R9390 gnd.n7279 gnd.n393 585
R9391 gnd.n7283 gnd.n393 585
R9392 gnd.n7281 gnd.n7280 585
R9393 gnd.n7282 gnd.n7281 585
R9394 gnd.n396 gnd.n395 585
R9395 gnd.n395 gnd.n394 585
R9396 gnd.n7274 gnd.n7273 585
R9397 gnd.n7273 gnd.n7272 585
R9398 gnd.n399 gnd.n398 585
R9399 gnd.n7271 gnd.n399 585
R9400 gnd.n7269 gnd.n7268 585
R9401 gnd.n7270 gnd.n7269 585
R9402 gnd.n402 gnd.n401 585
R9403 gnd.n401 gnd.n400 585
R9404 gnd.n7264 gnd.n7263 585
R9405 gnd.n7263 gnd.n7262 585
R9406 gnd.n405 gnd.n404 585
R9407 gnd.n7261 gnd.n405 585
R9408 gnd.n7259 gnd.n7258 585
R9409 gnd.n7260 gnd.n7259 585
R9410 gnd.n408 gnd.n407 585
R9411 gnd.n407 gnd.n406 585
R9412 gnd.n7254 gnd.n7253 585
R9413 gnd.n7253 gnd.n7252 585
R9414 gnd.n411 gnd.n410 585
R9415 gnd.n7251 gnd.n411 585
R9416 gnd.n7249 gnd.n7248 585
R9417 gnd.n7250 gnd.n7249 585
R9418 gnd.n414 gnd.n413 585
R9419 gnd.n413 gnd.n412 585
R9420 gnd.n7244 gnd.n7243 585
R9421 gnd.n7243 gnd.n7242 585
R9422 gnd.n417 gnd.n416 585
R9423 gnd.n7241 gnd.n417 585
R9424 gnd.n7239 gnd.n7238 585
R9425 gnd.n7240 gnd.n7239 585
R9426 gnd.n420 gnd.n419 585
R9427 gnd.n419 gnd.n418 585
R9428 gnd.n7234 gnd.n7233 585
R9429 gnd.n7233 gnd.n7232 585
R9430 gnd.n423 gnd.n422 585
R9431 gnd.n7231 gnd.n423 585
R9432 gnd.n7229 gnd.n7228 585
R9433 gnd.n7230 gnd.n7229 585
R9434 gnd.n426 gnd.n425 585
R9435 gnd.n425 gnd.n424 585
R9436 gnd.n7224 gnd.n7223 585
R9437 gnd.n7223 gnd.n7222 585
R9438 gnd.n429 gnd.n428 585
R9439 gnd.n7221 gnd.n429 585
R9440 gnd.n7219 gnd.n7218 585
R9441 gnd.n7220 gnd.n7219 585
R9442 gnd.n432 gnd.n431 585
R9443 gnd.n431 gnd.n430 585
R9444 gnd.n7214 gnd.n7213 585
R9445 gnd.n7213 gnd.n7212 585
R9446 gnd.n435 gnd.n434 585
R9447 gnd.n7211 gnd.n435 585
R9448 gnd.n7209 gnd.n7208 585
R9449 gnd.n7210 gnd.n7209 585
R9450 gnd.n438 gnd.n437 585
R9451 gnd.n437 gnd.n436 585
R9452 gnd.n7204 gnd.n7203 585
R9453 gnd.n7203 gnd.n7202 585
R9454 gnd.n441 gnd.n440 585
R9455 gnd.n7201 gnd.n441 585
R9456 gnd.n7199 gnd.n7198 585
R9457 gnd.n7200 gnd.n7199 585
R9458 gnd.n444 gnd.n443 585
R9459 gnd.n443 gnd.n442 585
R9460 gnd.n7194 gnd.n7193 585
R9461 gnd.n7193 gnd.n7192 585
R9462 gnd.n447 gnd.n446 585
R9463 gnd.n7191 gnd.n447 585
R9464 gnd.n7189 gnd.n7188 585
R9465 gnd.n7190 gnd.n7189 585
R9466 gnd.n450 gnd.n449 585
R9467 gnd.n449 gnd.n448 585
R9468 gnd.n7184 gnd.n7183 585
R9469 gnd.n7183 gnd.n7182 585
R9470 gnd.n453 gnd.n452 585
R9471 gnd.n7181 gnd.n453 585
R9472 gnd.n7179 gnd.n7178 585
R9473 gnd.n7180 gnd.n7179 585
R9474 gnd.n456 gnd.n455 585
R9475 gnd.n455 gnd.n454 585
R9476 gnd.n7174 gnd.n7173 585
R9477 gnd.n7173 gnd.n7172 585
R9478 gnd.n459 gnd.n458 585
R9479 gnd.n7171 gnd.n459 585
R9480 gnd.n7169 gnd.n7168 585
R9481 gnd.n7170 gnd.n7169 585
R9482 gnd.n462 gnd.n461 585
R9483 gnd.n461 gnd.n460 585
R9484 gnd.n7164 gnd.n7163 585
R9485 gnd.n7163 gnd.n7162 585
R9486 gnd.n465 gnd.n464 585
R9487 gnd.n7161 gnd.n465 585
R9488 gnd.n7159 gnd.n7158 585
R9489 gnd.n7160 gnd.n7159 585
R9490 gnd.n468 gnd.n467 585
R9491 gnd.n467 gnd.n466 585
R9492 gnd.n7154 gnd.n7153 585
R9493 gnd.n7153 gnd.n7152 585
R9494 gnd.n471 gnd.n470 585
R9495 gnd.n7151 gnd.n471 585
R9496 gnd.n7149 gnd.n7148 585
R9497 gnd.n7150 gnd.n7149 585
R9498 gnd.n474 gnd.n473 585
R9499 gnd.n473 gnd.n472 585
R9500 gnd.n7144 gnd.n7143 585
R9501 gnd.n7143 gnd.n7142 585
R9502 gnd.n477 gnd.n476 585
R9503 gnd.n7141 gnd.n477 585
R9504 gnd.n7139 gnd.n7138 585
R9505 gnd.n7140 gnd.n7139 585
R9506 gnd.n480 gnd.n479 585
R9507 gnd.n479 gnd.n478 585
R9508 gnd.n7134 gnd.n7133 585
R9509 gnd.n7133 gnd.n7132 585
R9510 gnd.n483 gnd.n482 585
R9511 gnd.n7131 gnd.n483 585
R9512 gnd.n7129 gnd.n7128 585
R9513 gnd.n7130 gnd.n7129 585
R9514 gnd.n486 gnd.n485 585
R9515 gnd.n485 gnd.n484 585
R9516 gnd.n7124 gnd.n7123 585
R9517 gnd.n7123 gnd.n7122 585
R9518 gnd.n489 gnd.n488 585
R9519 gnd.n7121 gnd.n489 585
R9520 gnd.n7119 gnd.n7118 585
R9521 gnd.n7120 gnd.n7119 585
R9522 gnd.n492 gnd.n491 585
R9523 gnd.n491 gnd.n490 585
R9524 gnd.n7114 gnd.n7113 585
R9525 gnd.n7113 gnd.n7112 585
R9526 gnd.n495 gnd.n494 585
R9527 gnd.n7111 gnd.n495 585
R9528 gnd.n7109 gnd.n7108 585
R9529 gnd.n7110 gnd.n7109 585
R9530 gnd.n498 gnd.n497 585
R9531 gnd.n497 gnd.n496 585
R9532 gnd.n7104 gnd.n7103 585
R9533 gnd.n7103 gnd.n7102 585
R9534 gnd.n501 gnd.n500 585
R9535 gnd.n7101 gnd.n501 585
R9536 gnd.n7099 gnd.n7098 585
R9537 gnd.n7100 gnd.n7099 585
R9538 gnd.n504 gnd.n503 585
R9539 gnd.n503 gnd.n502 585
R9540 gnd.n7094 gnd.n7093 585
R9541 gnd.n7093 gnd.n7092 585
R9542 gnd.n507 gnd.n506 585
R9543 gnd.n7091 gnd.n507 585
R9544 gnd.n7089 gnd.n7088 585
R9545 gnd.n7090 gnd.n7089 585
R9546 gnd.n510 gnd.n509 585
R9547 gnd.n509 gnd.n508 585
R9548 gnd.n7084 gnd.n7083 585
R9549 gnd.n7083 gnd.n7082 585
R9550 gnd.n513 gnd.n512 585
R9551 gnd.n7081 gnd.n513 585
R9552 gnd.n7079 gnd.n7078 585
R9553 gnd.n7080 gnd.n7079 585
R9554 gnd.n516 gnd.n515 585
R9555 gnd.n515 gnd.n514 585
R9556 gnd.n6412 gnd.n6411 585
R9557 gnd.n6411 gnd.n6410 585
R9558 gnd.n6413 gnd.n1060 585
R9559 gnd.n4778 gnd.n1060 585
R9560 gnd.n6415 gnd.n6414 585
R9561 gnd.n6416 gnd.n6415 585
R9562 gnd.n1045 gnd.n1044 585
R9563 gnd.n4771 gnd.n1045 585
R9564 gnd.n6424 gnd.n6423 585
R9565 gnd.n6423 gnd.n6422 585
R9566 gnd.n6425 gnd.n1040 585
R9567 gnd.n4762 gnd.n1040 585
R9568 gnd.n6427 gnd.n6426 585
R9569 gnd.n6428 gnd.n6427 585
R9570 gnd.n1025 gnd.n1024 585
R9571 gnd.n4756 gnd.n1025 585
R9572 gnd.n6436 gnd.n6435 585
R9573 gnd.n6435 gnd.n6434 585
R9574 gnd.n6437 gnd.n1020 585
R9575 gnd.n4691 gnd.n1020 585
R9576 gnd.n6439 gnd.n6438 585
R9577 gnd.n6440 gnd.n6439 585
R9578 gnd.n1005 gnd.n1004 585
R9579 gnd.n4685 gnd.n1005 585
R9580 gnd.n6448 gnd.n6447 585
R9581 gnd.n6447 gnd.n6446 585
R9582 gnd.n6449 gnd.n1000 585
R9583 gnd.n4679 gnd.n1000 585
R9584 gnd.n6451 gnd.n6450 585
R9585 gnd.n6452 gnd.n6451 585
R9586 gnd.n985 gnd.n984 585
R9587 gnd.n4708 gnd.n985 585
R9588 gnd.n6460 gnd.n6459 585
R9589 gnd.n6459 gnd.n6458 585
R9590 gnd.n6461 gnd.n980 585
R9591 gnd.n4672 gnd.n980 585
R9592 gnd.n6463 gnd.n6462 585
R9593 gnd.n6464 gnd.n6463 585
R9594 gnd.n966 gnd.n965 585
R9595 gnd.n4664 gnd.n966 585
R9596 gnd.n6472 gnd.n6471 585
R9597 gnd.n6471 gnd.n6470 585
R9598 gnd.n6473 gnd.n960 585
R9599 gnd.n4657 gnd.n960 585
R9600 gnd.n6475 gnd.n6474 585
R9601 gnd.n6476 gnd.n6475 585
R9602 gnd.n961 gnd.n959 585
R9603 gnd.n4649 gnd.n959 585
R9604 gnd.n4609 gnd.n2518 585
R9605 gnd.n4619 gnd.n2518 585
R9606 gnd.n4610 gnd.n2525 585
R9607 gnd.n2525 gnd.n2516 585
R9608 gnd.n4612 gnd.n4611 585
R9609 gnd.n4613 gnd.n4612 585
R9610 gnd.n2526 gnd.n2524 585
R9611 gnd.n4600 gnd.n2524 585
R9612 gnd.n4575 gnd.n941 585
R9613 gnd.n6483 gnd.n941 585
R9614 gnd.n4577 gnd.n4576 585
R9615 gnd.n4576 gnd.n938 585
R9616 gnd.n4578 gnd.n2537 585
R9617 gnd.n4585 gnd.n2537 585
R9618 gnd.n4580 gnd.n4579 585
R9619 gnd.n4581 gnd.n4580 585
R9620 gnd.n2543 gnd.n2542 585
R9621 gnd.n2542 gnd.n2540 585
R9622 gnd.n4552 gnd.n2550 585
R9623 gnd.n4565 gnd.n2550 585
R9624 gnd.n4553 gnd.n2560 585
R9625 gnd.n2560 gnd.n2558 585
R9626 gnd.n4555 gnd.n4554 585
R9627 gnd.n4556 gnd.n4555 585
R9628 gnd.n2561 gnd.n2559 585
R9629 gnd.n4545 gnd.n2559 585
R9630 gnd.n4510 gnd.n4509 585
R9631 gnd.n4509 gnd.n2566 585
R9632 gnd.n4511 gnd.n2573 585
R9633 gnd.n4525 gnd.n2573 585
R9634 gnd.n4512 gnd.n2585 585
R9635 gnd.n2585 gnd.n2583 585
R9636 gnd.n4514 gnd.n4513 585
R9637 gnd.n4515 gnd.n4514 585
R9638 gnd.n2586 gnd.n2584 585
R9639 gnd.n2584 gnd.n2580 585
R9640 gnd.n4487 gnd.n2594 585
R9641 gnd.n4499 gnd.n2594 585
R9642 gnd.n4488 gnd.n2604 585
R9643 gnd.n2604 gnd.n2592 585
R9644 gnd.n4490 gnd.n4489 585
R9645 gnd.n4491 gnd.n4490 585
R9646 gnd.n2605 gnd.n2603 585
R9647 gnd.n2603 gnd.n2600 585
R9648 gnd.n4467 gnd.n2611 585
R9649 gnd.n4479 gnd.n2611 585
R9650 gnd.n4468 gnd.n2622 585
R9651 gnd.n2622 gnd.n2620 585
R9652 gnd.n4470 gnd.n4469 585
R9653 gnd.n4471 gnd.n4470 585
R9654 gnd.n2623 gnd.n2621 585
R9655 gnd.n2621 gnd.n2617 585
R9656 gnd.n2644 gnd.n2630 585
R9657 gnd.n4459 gnd.n2630 585
R9658 gnd.n2642 gnd.n2640 585
R9659 gnd.n2640 gnd.n2628 585
R9660 gnd.n4450 gnd.n4449 585
R9661 gnd.n4451 gnd.n4450 585
R9662 gnd.n2641 gnd.n2639 585
R9663 gnd.n2639 gnd.n2636 585
R9664 gnd.n4321 gnd.n4320 585
R9665 gnd.n4319 gnd.n4318 585
R9666 gnd.n4317 gnd.n4316 585
R9667 gnd.n4315 gnd.n4314 585
R9668 gnd.n4313 gnd.n4312 585
R9669 gnd.n4311 gnd.n4310 585
R9670 gnd.n4309 gnd.n4308 585
R9671 gnd.n4307 gnd.n4306 585
R9672 gnd.n4305 gnd.n4304 585
R9673 gnd.n4303 gnd.n4302 585
R9674 gnd.n4301 gnd.n4300 585
R9675 gnd.n4299 gnd.n4298 585
R9676 gnd.n4297 gnd.n4296 585
R9677 gnd.n4295 gnd.n4294 585
R9678 gnd.n4293 gnd.n4292 585
R9679 gnd.n4291 gnd.n4290 585
R9680 gnd.n4289 gnd.n4288 585
R9681 gnd.n4248 gnd.n4245 585
R9682 gnd.n4284 gnd.n4164 585
R9683 gnd.n4441 gnd.n4164 585
R9684 gnd.n4795 gnd.n4794 585
R9685 gnd.n4796 gnd.n2463 585
R9686 gnd.n4797 gnd.n2459 585
R9687 gnd.n2457 gnd.n2448 585
R9688 gnd.n4804 gnd.n2447 585
R9689 gnd.n4805 gnd.n2445 585
R9690 gnd.n2444 gnd.n2437 585
R9691 gnd.n4812 gnd.n2436 585
R9692 gnd.n4813 gnd.n2435 585
R9693 gnd.n2433 gnd.n2425 585
R9694 gnd.n4820 gnd.n2424 585
R9695 gnd.n4821 gnd.n2422 585
R9696 gnd.n2421 gnd.n2414 585
R9697 gnd.n4828 gnd.n2413 585
R9698 gnd.n4829 gnd.n2412 585
R9699 gnd.n2410 gnd.n2402 585
R9700 gnd.n4836 gnd.n2401 585
R9701 gnd.n4837 gnd.n2399 585
R9702 gnd.n2398 gnd.n1064 585
R9703 gnd.n1073 gnd.n1064 585
R9704 gnd.n4781 gnd.n1067 585
R9705 gnd.n6410 gnd.n1067 585
R9706 gnd.n4780 gnd.n4779 585
R9707 gnd.n4779 gnd.n4778 585
R9708 gnd.n2466 gnd.n1059 585
R9709 gnd.n6416 gnd.n1059 585
R9710 gnd.n4770 gnd.n4769 585
R9711 gnd.n4771 gnd.n4770 585
R9712 gnd.n2470 gnd.n1048 585
R9713 gnd.n6422 gnd.n1048 585
R9714 gnd.n4764 gnd.n4763 585
R9715 gnd.n4763 gnd.n4762 585
R9716 gnd.n2472 gnd.n1038 585
R9717 gnd.n6428 gnd.n1038 585
R9718 gnd.n4694 gnd.n2475 585
R9719 gnd.n4756 gnd.n2475 585
R9720 gnd.n4695 gnd.n1028 585
R9721 gnd.n6434 gnd.n1028 585
R9722 gnd.n4696 gnd.n4692 585
R9723 gnd.n4692 gnd.n4691 585
R9724 gnd.n2494 gnd.n1018 585
R9725 gnd.n6440 gnd.n1018 585
R9726 gnd.n4700 gnd.n2493 585
R9727 gnd.n4685 gnd.n2493 585
R9728 gnd.n4701 gnd.n1008 585
R9729 gnd.n6446 gnd.n1008 585
R9730 gnd.n4702 gnd.n2492 585
R9731 gnd.n4679 gnd.n2492 585
R9732 gnd.n2489 gnd.n998 585
R9733 gnd.n6452 gnd.n998 585
R9734 gnd.n4707 gnd.n4706 585
R9735 gnd.n4708 gnd.n4707 585
R9736 gnd.n2488 gnd.n988 585
R9737 gnd.n6458 gnd.n988 585
R9738 gnd.n4671 gnd.n4670 585
R9739 gnd.n4672 gnd.n4671 585
R9740 gnd.n2497 gnd.n978 585
R9741 gnd.n6464 gnd.n978 585
R9742 gnd.n4666 gnd.n4665 585
R9743 gnd.n4665 gnd.n4664 585
R9744 gnd.n2499 gnd.n969 585
R9745 gnd.n6470 gnd.n969 585
R9746 gnd.n4656 gnd.n4655 585
R9747 gnd.n4657 gnd.n4656 585
R9748 gnd.n2502 gnd.n957 585
R9749 gnd.n6476 gnd.n957 585
R9750 gnd.n4651 gnd.n4650 585
R9751 gnd.n4650 gnd.n4649 585
R9752 gnd.n2505 gnd.n2504 585
R9753 gnd.n4619 gnd.n2505 585
R9754 gnd.n4593 gnd.n4592 585
R9755 gnd.n4592 gnd.n2516 585
R9756 gnd.n4597 gnd.n2522 585
R9757 gnd.n4613 gnd.n2522 585
R9758 gnd.n4599 gnd.n4598 585
R9759 gnd.n4600 gnd.n4599 585
R9760 gnd.n2532 gnd.n940 585
R9761 gnd.n6483 gnd.n940 585
R9762 gnd.n4588 gnd.n4587 585
R9763 gnd.n4587 gnd.n938 585
R9764 gnd.n4586 gnd.n2534 585
R9765 gnd.n4586 gnd.n4585 585
R9766 gnd.n4536 gnd.n2535 585
R9767 gnd.n4581 gnd.n2535 585
R9768 gnd.n4538 gnd.n4537 585
R9769 gnd.n4537 gnd.n2540 585
R9770 gnd.n4539 gnd.n2549 585
R9771 gnd.n4565 gnd.n2549 585
R9772 gnd.n4541 gnd.n4540 585
R9773 gnd.n4540 gnd.n2558 585
R9774 gnd.n4542 gnd.n2557 585
R9775 gnd.n4556 gnd.n2557 585
R9776 gnd.n4544 gnd.n4543 585
R9777 gnd.n4545 gnd.n4544 585
R9778 gnd.n2568 gnd.n2567 585
R9779 gnd.n2567 gnd.n2566 585
R9780 gnd.n4527 gnd.n4526 585
R9781 gnd.n4526 gnd.n4525 585
R9782 gnd.n2571 gnd.n2570 585
R9783 gnd.n2583 gnd.n2571 585
R9784 gnd.n4262 gnd.n2582 585
R9785 gnd.n4515 gnd.n2582 585
R9786 gnd.n4264 gnd.n4263 585
R9787 gnd.n4263 gnd.n2580 585
R9788 gnd.n4265 gnd.n2593 585
R9789 gnd.n4499 gnd.n2593 585
R9790 gnd.n4267 gnd.n4266 585
R9791 gnd.n4266 gnd.n2592 585
R9792 gnd.n4268 gnd.n2602 585
R9793 gnd.n4491 gnd.n2602 585
R9794 gnd.n4270 gnd.n4269 585
R9795 gnd.n4269 gnd.n2600 585
R9796 gnd.n4271 gnd.n2610 585
R9797 gnd.n4479 gnd.n2610 585
R9798 gnd.n4273 gnd.n4272 585
R9799 gnd.n4272 gnd.n2620 585
R9800 gnd.n4274 gnd.n2619 585
R9801 gnd.n4471 gnd.n2619 585
R9802 gnd.n4276 gnd.n4275 585
R9803 gnd.n4275 gnd.n2617 585
R9804 gnd.n4277 gnd.n2629 585
R9805 gnd.n4459 gnd.n2629 585
R9806 gnd.n4279 gnd.n4278 585
R9807 gnd.n4278 gnd.n2628 585
R9808 gnd.n4280 gnd.n2638 585
R9809 gnd.n4451 gnd.n2638 585
R9810 gnd.n4282 gnd.n4281 585
R9811 gnd.n4281 gnd.n2636 585
R9812 gnd.n4035 gnd.n4034 585
R9813 gnd.n4036 gnd.n4035 585
R9814 gnd.n2725 gnd.n2724 585
R9815 gnd.n2731 gnd.n2724 585
R9816 gnd.n4010 gnd.n2743 585
R9817 gnd.n2743 gnd.n2730 585
R9818 gnd.n4012 gnd.n4011 585
R9819 gnd.n4013 gnd.n4012 585
R9820 gnd.n2744 gnd.n2742 585
R9821 gnd.n2742 gnd.n2738 585
R9822 gnd.n3744 gnd.n3743 585
R9823 gnd.n3743 gnd.n3742 585
R9824 gnd.n2749 gnd.n2748 585
R9825 gnd.n3712 gnd.n2749 585
R9826 gnd.n3732 gnd.n3731 585
R9827 gnd.n3731 gnd.n3730 585
R9828 gnd.n2756 gnd.n2755 585
R9829 gnd.n3718 gnd.n2756 585
R9830 gnd.n3688 gnd.n2776 585
R9831 gnd.n2776 gnd.n2775 585
R9832 gnd.n3690 gnd.n3689 585
R9833 gnd.n3691 gnd.n3690 585
R9834 gnd.n2777 gnd.n2774 585
R9835 gnd.n2785 gnd.n2774 585
R9836 gnd.n3666 gnd.n2797 585
R9837 gnd.n2797 gnd.n2784 585
R9838 gnd.n3668 gnd.n3667 585
R9839 gnd.n3669 gnd.n3668 585
R9840 gnd.n2798 gnd.n2796 585
R9841 gnd.n2796 gnd.n2792 585
R9842 gnd.n3654 gnd.n3653 585
R9843 gnd.n3653 gnd.n3652 585
R9844 gnd.n2803 gnd.n2802 585
R9845 gnd.n2813 gnd.n2803 585
R9846 gnd.n3643 gnd.n3642 585
R9847 gnd.n3642 gnd.n3641 585
R9848 gnd.n2810 gnd.n2809 585
R9849 gnd.n3629 gnd.n2810 585
R9850 gnd.n3603 gnd.n2831 585
R9851 gnd.n2831 gnd.n2820 585
R9852 gnd.n3605 gnd.n3604 585
R9853 gnd.n3606 gnd.n3605 585
R9854 gnd.n2832 gnd.n2830 585
R9855 gnd.n2840 gnd.n2830 585
R9856 gnd.n3581 gnd.n2852 585
R9857 gnd.n2852 gnd.n2839 585
R9858 gnd.n3583 gnd.n3582 585
R9859 gnd.n3584 gnd.n3583 585
R9860 gnd.n2853 gnd.n2851 585
R9861 gnd.n2851 gnd.n2847 585
R9862 gnd.n3569 gnd.n3568 585
R9863 gnd.n3568 gnd.n3567 585
R9864 gnd.n2858 gnd.n2857 585
R9865 gnd.n2867 gnd.n2858 585
R9866 gnd.n3558 gnd.n3557 585
R9867 gnd.n3557 gnd.n3556 585
R9868 gnd.n2865 gnd.n2864 585
R9869 gnd.n3544 gnd.n2865 585
R9870 gnd.n2982 gnd.n2981 585
R9871 gnd.n2982 gnd.n2874 585
R9872 gnd.n3501 gnd.n3500 585
R9873 gnd.n3500 gnd.n3499 585
R9874 gnd.n3502 gnd.n2976 585
R9875 gnd.n2987 gnd.n2976 585
R9876 gnd.n3504 gnd.n3503 585
R9877 gnd.n3505 gnd.n3504 585
R9878 gnd.n2977 gnd.n2975 585
R9879 gnd.n3000 gnd.n2975 585
R9880 gnd.n2960 gnd.n2959 585
R9881 gnd.n2963 gnd.n2960 585
R9882 gnd.n3515 gnd.n3514 585
R9883 gnd.n3514 gnd.n3513 585
R9884 gnd.n3516 gnd.n2954 585
R9885 gnd.n3475 gnd.n2954 585
R9886 gnd.n3518 gnd.n3517 585
R9887 gnd.n3519 gnd.n3518 585
R9888 gnd.n2955 gnd.n2953 585
R9889 gnd.n3014 gnd.n2953 585
R9890 gnd.n3467 gnd.n3466 585
R9891 gnd.n3466 gnd.n3465 585
R9892 gnd.n3011 gnd.n3010 585
R9893 gnd.n3449 gnd.n3011 585
R9894 gnd.n3436 gnd.n3030 585
R9895 gnd.n3030 gnd.n3029 585
R9896 gnd.n3438 gnd.n3437 585
R9897 gnd.n3439 gnd.n3438 585
R9898 gnd.n3031 gnd.n3028 585
R9899 gnd.n3037 gnd.n3028 585
R9900 gnd.n3417 gnd.n3416 585
R9901 gnd.n3418 gnd.n3417 585
R9902 gnd.n3048 gnd.n3047 585
R9903 gnd.n3047 gnd.n3043 585
R9904 gnd.n3407 gnd.n3406 585
R9905 gnd.n3408 gnd.n3407 585
R9906 gnd.n3058 gnd.n3057 585
R9907 gnd.n3063 gnd.n3057 585
R9908 gnd.n3385 gnd.n3076 585
R9909 gnd.n3076 gnd.n3062 585
R9910 gnd.n3387 gnd.n3386 585
R9911 gnd.n3388 gnd.n3387 585
R9912 gnd.n3077 gnd.n3075 585
R9913 gnd.n3075 gnd.n3071 585
R9914 gnd.n3376 gnd.n3375 585
R9915 gnd.n3377 gnd.n3376 585
R9916 gnd.n3084 gnd.n3083 585
R9917 gnd.n3088 gnd.n3083 585
R9918 gnd.n3353 gnd.n3105 585
R9919 gnd.n3105 gnd.n3087 585
R9920 gnd.n3355 gnd.n3354 585
R9921 gnd.n3356 gnd.n3355 585
R9922 gnd.n3106 gnd.n3104 585
R9923 gnd.n3104 gnd.n3095 585
R9924 gnd.n3348 gnd.n3347 585
R9925 gnd.n3347 gnd.n3346 585
R9926 gnd.n3153 gnd.n3152 585
R9927 gnd.n3154 gnd.n3153 585
R9928 gnd.n3307 gnd.n3306 585
R9929 gnd.n3308 gnd.n3307 585
R9930 gnd.n3163 gnd.n3162 585
R9931 gnd.n3162 gnd.n3161 585
R9932 gnd.n3302 gnd.n3301 585
R9933 gnd.n3301 gnd.n3300 585
R9934 gnd.n3166 gnd.n3165 585
R9935 gnd.n3167 gnd.n3166 585
R9936 gnd.n3291 gnd.n3290 585
R9937 gnd.n3292 gnd.n3291 585
R9938 gnd.n3174 gnd.n3173 585
R9939 gnd.n3283 gnd.n3173 585
R9940 gnd.n3286 gnd.n3285 585
R9941 gnd.n3285 gnd.n3284 585
R9942 gnd.n3177 gnd.n3176 585
R9943 gnd.n3178 gnd.n3177 585
R9944 gnd.n3272 gnd.n3271 585
R9945 gnd.n3270 gnd.n3196 585
R9946 gnd.n3269 gnd.n3195 585
R9947 gnd.n3274 gnd.n3195 585
R9948 gnd.n3268 gnd.n3267 585
R9949 gnd.n3266 gnd.n3265 585
R9950 gnd.n3264 gnd.n3263 585
R9951 gnd.n3262 gnd.n3261 585
R9952 gnd.n3260 gnd.n3259 585
R9953 gnd.n3258 gnd.n3257 585
R9954 gnd.n3256 gnd.n3255 585
R9955 gnd.n3254 gnd.n3253 585
R9956 gnd.n3252 gnd.n3251 585
R9957 gnd.n3250 gnd.n3249 585
R9958 gnd.n3248 gnd.n3247 585
R9959 gnd.n3246 gnd.n3245 585
R9960 gnd.n3244 gnd.n3243 585
R9961 gnd.n3242 gnd.n3241 585
R9962 gnd.n3240 gnd.n3239 585
R9963 gnd.n3238 gnd.n3237 585
R9964 gnd.n3236 gnd.n3235 585
R9965 gnd.n3234 gnd.n3233 585
R9966 gnd.n3232 gnd.n3231 585
R9967 gnd.n3230 gnd.n3229 585
R9968 gnd.n3228 gnd.n3227 585
R9969 gnd.n3226 gnd.n3225 585
R9970 gnd.n3183 gnd.n3182 585
R9971 gnd.n3277 gnd.n3276 585
R9972 gnd.n4039 gnd.n4038 585
R9973 gnd.n4041 gnd.n4040 585
R9974 gnd.n4043 gnd.n4042 585
R9975 gnd.n4045 gnd.n4044 585
R9976 gnd.n4047 gnd.n4046 585
R9977 gnd.n4049 gnd.n4048 585
R9978 gnd.n4051 gnd.n4050 585
R9979 gnd.n4053 gnd.n4052 585
R9980 gnd.n4055 gnd.n4054 585
R9981 gnd.n4057 gnd.n4056 585
R9982 gnd.n4059 gnd.n4058 585
R9983 gnd.n4061 gnd.n4060 585
R9984 gnd.n4063 gnd.n4062 585
R9985 gnd.n4065 gnd.n4064 585
R9986 gnd.n4067 gnd.n4066 585
R9987 gnd.n4069 gnd.n4068 585
R9988 gnd.n4071 gnd.n4070 585
R9989 gnd.n4073 gnd.n4072 585
R9990 gnd.n4075 gnd.n4074 585
R9991 gnd.n4077 gnd.n4076 585
R9992 gnd.n4079 gnd.n4078 585
R9993 gnd.n4081 gnd.n4080 585
R9994 gnd.n4083 gnd.n4082 585
R9995 gnd.n4085 gnd.n4084 585
R9996 gnd.n4087 gnd.n4086 585
R9997 gnd.n4088 gnd.n2692 585
R9998 gnd.n4089 gnd.n2650 585
R9999 gnd.n4127 gnd.n2650 585
R10000 gnd.n4037 gnd.n2722 585
R10001 gnd.n4037 gnd.n4036 585
R10002 gnd.n3705 gnd.n2721 585
R10003 gnd.n2731 gnd.n2721 585
R10004 gnd.n3707 gnd.n3706 585
R10005 gnd.n3706 gnd.n2730 585
R10006 gnd.n3708 gnd.n2740 585
R10007 gnd.n4013 gnd.n2740 585
R10008 gnd.n3710 gnd.n3709 585
R10009 gnd.n3709 gnd.n2738 585
R10010 gnd.n3711 gnd.n2751 585
R10011 gnd.n3742 gnd.n2751 585
R10012 gnd.n3714 gnd.n3713 585
R10013 gnd.n3713 gnd.n3712 585
R10014 gnd.n3715 gnd.n2758 585
R10015 gnd.n3730 gnd.n2758 585
R10016 gnd.n3717 gnd.n3716 585
R10017 gnd.n3718 gnd.n3717 585
R10018 gnd.n2768 gnd.n2767 585
R10019 gnd.n2775 gnd.n2767 585
R10020 gnd.n3693 gnd.n3692 585
R10021 gnd.n3692 gnd.n3691 585
R10022 gnd.n2771 gnd.n2770 585
R10023 gnd.n2785 gnd.n2771 585
R10024 gnd.n3619 gnd.n3618 585
R10025 gnd.n3618 gnd.n2784 585
R10026 gnd.n3620 gnd.n2794 585
R10027 gnd.n3669 gnd.n2794 585
R10028 gnd.n3622 gnd.n3621 585
R10029 gnd.n3621 gnd.n2792 585
R10030 gnd.n3623 gnd.n2805 585
R10031 gnd.n3652 gnd.n2805 585
R10032 gnd.n3625 gnd.n3624 585
R10033 gnd.n3624 gnd.n2813 585
R10034 gnd.n3626 gnd.n2812 585
R10035 gnd.n3641 gnd.n2812 585
R10036 gnd.n3628 gnd.n3627 585
R10037 gnd.n3629 gnd.n3628 585
R10038 gnd.n2824 gnd.n2823 585
R10039 gnd.n2823 gnd.n2820 585
R10040 gnd.n3608 gnd.n3607 585
R10041 gnd.n3607 gnd.n3606 585
R10042 gnd.n2827 gnd.n2826 585
R10043 gnd.n2840 gnd.n2827 585
R10044 gnd.n3532 gnd.n3531 585
R10045 gnd.n3531 gnd.n2839 585
R10046 gnd.n3533 gnd.n2849 585
R10047 gnd.n3584 gnd.n2849 585
R10048 gnd.n3535 gnd.n3534 585
R10049 gnd.n3534 gnd.n2847 585
R10050 gnd.n3536 gnd.n2860 585
R10051 gnd.n3567 gnd.n2860 585
R10052 gnd.n3538 gnd.n3537 585
R10053 gnd.n3537 gnd.n2867 585
R10054 gnd.n3539 gnd.n2866 585
R10055 gnd.n3556 gnd.n2866 585
R10056 gnd.n3541 gnd.n3540 585
R10057 gnd.n3544 gnd.n3541 585
R10058 gnd.n2877 gnd.n2876 585
R10059 gnd.n2876 gnd.n2874 585
R10060 gnd.n2984 gnd.n2983 585
R10061 gnd.n3499 gnd.n2983 585
R10062 gnd.n2986 gnd.n2985 585
R10063 gnd.n2987 gnd.n2986 585
R10064 gnd.n2997 gnd.n2973 585
R10065 gnd.n3505 gnd.n2973 585
R10066 gnd.n2999 gnd.n2998 585
R10067 gnd.n3000 gnd.n2999 585
R10068 gnd.n2996 gnd.n2995 585
R10069 gnd.n2996 gnd.n2963 585
R10070 gnd.n2994 gnd.n2961 585
R10071 gnd.n3513 gnd.n2961 585
R10072 gnd.n2950 gnd.n2948 585
R10073 gnd.n3475 gnd.n2950 585
R10074 gnd.n3521 gnd.n3520 585
R10075 gnd.n3520 gnd.n3519 585
R10076 gnd.n2949 gnd.n2947 585
R10077 gnd.n3014 gnd.n2949 585
R10078 gnd.n3446 gnd.n3013 585
R10079 gnd.n3465 gnd.n3013 585
R10080 gnd.n3448 gnd.n3447 585
R10081 gnd.n3449 gnd.n3448 585
R10082 gnd.n3023 gnd.n3022 585
R10083 gnd.n3029 gnd.n3022 585
R10084 gnd.n3441 gnd.n3440 585
R10085 gnd.n3440 gnd.n3439 585
R10086 gnd.n3026 gnd.n3025 585
R10087 gnd.n3037 gnd.n3026 585
R10088 gnd.n3326 gnd.n3045 585
R10089 gnd.n3418 gnd.n3045 585
R10090 gnd.n3328 gnd.n3327 585
R10091 gnd.n3327 gnd.n3043 585
R10092 gnd.n3329 gnd.n3056 585
R10093 gnd.n3408 gnd.n3056 585
R10094 gnd.n3331 gnd.n3330 585
R10095 gnd.n3331 gnd.n3063 585
R10096 gnd.n3333 gnd.n3332 585
R10097 gnd.n3332 gnd.n3062 585
R10098 gnd.n3334 gnd.n3073 585
R10099 gnd.n3388 gnd.n3073 585
R10100 gnd.n3336 gnd.n3335 585
R10101 gnd.n3335 gnd.n3071 585
R10102 gnd.n3337 gnd.n3082 585
R10103 gnd.n3377 gnd.n3082 585
R10104 gnd.n3339 gnd.n3338 585
R10105 gnd.n3339 gnd.n3088 585
R10106 gnd.n3341 gnd.n3340 585
R10107 gnd.n3340 gnd.n3087 585
R10108 gnd.n3342 gnd.n3103 585
R10109 gnd.n3356 gnd.n3103 585
R10110 gnd.n3343 gnd.n3156 585
R10111 gnd.n3156 gnd.n3095 585
R10112 gnd.n3345 gnd.n3344 585
R10113 gnd.n3346 gnd.n3345 585
R10114 gnd.n3157 gnd.n3155 585
R10115 gnd.n3155 gnd.n3154 585
R10116 gnd.n3310 gnd.n3309 585
R10117 gnd.n3309 gnd.n3308 585
R10118 gnd.n3160 gnd.n3159 585
R10119 gnd.n3161 gnd.n3160 585
R10120 gnd.n3299 gnd.n3298 585
R10121 gnd.n3300 gnd.n3299 585
R10122 gnd.n3169 gnd.n3168 585
R10123 gnd.n3168 gnd.n3167 585
R10124 gnd.n3294 gnd.n3293 585
R10125 gnd.n3293 gnd.n3292 585
R10126 gnd.n3172 gnd.n3171 585
R10127 gnd.n3283 gnd.n3172 585
R10128 gnd.n3282 gnd.n3281 585
R10129 gnd.n3284 gnd.n3282 585
R10130 gnd.n3180 gnd.n3179 585
R10131 gnd.n3179 gnd.n3178 585
R10132 gnd.n7551 gnd.n7550 585
R10133 gnd.n7550 gnd.n7549 585
R10134 gnd.n7552 gnd.n204 585
R10135 gnd.n209 gnd.n204 585
R10136 gnd.n7554 gnd.n7553 585
R10137 gnd.n7555 gnd.n7554 585
R10138 gnd.n190 gnd.n189 585
R10139 gnd.n194 gnd.n190 585
R10140 gnd.n7563 gnd.n7562 585
R10141 gnd.n7562 gnd.n7561 585
R10142 gnd.n7564 gnd.n185 585
R10143 gnd.n191 gnd.n185 585
R10144 gnd.n7566 gnd.n7565 585
R10145 gnd.n7567 gnd.n7566 585
R10146 gnd.n170 gnd.n169 585
R10147 gnd.n174 gnd.n170 585
R10148 gnd.n7575 gnd.n7574 585
R10149 gnd.n7574 gnd.n7573 585
R10150 gnd.n7576 gnd.n165 585
R10151 gnd.n171 gnd.n165 585
R10152 gnd.n7578 gnd.n7577 585
R10153 gnd.n7579 gnd.n7578 585
R10154 gnd.n152 gnd.n151 585
R10155 gnd.n162 gnd.n152 585
R10156 gnd.n7587 gnd.n7586 585
R10157 gnd.n7586 gnd.n7585 585
R10158 gnd.n7588 gnd.n147 585
R10159 gnd.n147 gnd.n146 585
R10160 gnd.n7590 gnd.n7589 585
R10161 gnd.n7591 gnd.n7590 585
R10162 gnd.n132 gnd.n131 585
R10163 gnd.n136 gnd.n132 585
R10164 gnd.n7599 gnd.n7598 585
R10165 gnd.n7598 gnd.n7597 585
R10166 gnd.n7600 gnd.n127 585
R10167 gnd.n133 gnd.n127 585
R10168 gnd.n7602 gnd.n7601 585
R10169 gnd.n7603 gnd.n7602 585
R10170 gnd.n115 gnd.n114 585
R10171 gnd.n124 gnd.n115 585
R10172 gnd.n7611 gnd.n7610 585
R10173 gnd.n7610 gnd.n7609 585
R10174 gnd.n7612 gnd.n109 585
R10175 gnd.n109 gnd.n107 585
R10176 gnd.n7614 gnd.n7613 585
R10177 gnd.n7615 gnd.n7614 585
R10178 gnd.n110 gnd.n108 585
R10179 gnd.n7357 gnd.n108 585
R10180 gnd.n7313 gnd.n7312 585
R10181 gnd.n7312 gnd.n368 585
R10182 gnd.n7311 gnd.n91 585
R10183 gnd.n7623 gnd.n91 585
R10184 gnd.n7310 gnd.n7309 585
R10185 gnd.n7309 gnd.n7308 585
R10186 gnd.n374 gnd.n372 585
R10187 gnd.n7295 gnd.n374 585
R10188 gnd.n7301 gnd.n7300 585
R10189 gnd.n7300 gnd.n7299 585
R10190 gnd.n380 gnd.n379 585
R10191 gnd.n1699 gnd.n380 585
R10192 gnd.n1691 gnd.n1690 585
R10193 gnd.n5887 gnd.n1691 585
R10194 gnd.n5893 gnd.n5892 585
R10195 gnd.n5892 gnd.n5891 585
R10196 gnd.n5894 gnd.n1686 585
R10197 gnd.n5858 gnd.n1686 585
R10198 gnd.n5896 gnd.n5895 585
R10199 gnd.n5897 gnd.n5896 585
R10200 gnd.n1671 gnd.n1670 585
R10201 gnd.n5874 gnd.n1671 585
R10202 gnd.n5905 gnd.n5904 585
R10203 gnd.n5904 gnd.n5903 585
R10204 gnd.n5906 gnd.n1666 585
R10205 gnd.n5844 gnd.n1666 585
R10206 gnd.n5908 gnd.n5907 585
R10207 gnd.n5909 gnd.n5908 585
R10208 gnd.n1651 gnd.n1650 585
R10209 gnd.n5836 gnd.n1651 585
R10210 gnd.n5917 gnd.n5916 585
R10211 gnd.n5916 gnd.n5915 585
R10212 gnd.n5918 gnd.n1646 585
R10213 gnd.n5829 gnd.n1646 585
R10214 gnd.n5920 gnd.n5919 585
R10215 gnd.n5921 gnd.n5920 585
R10216 gnd.n1631 gnd.n1630 585
R10217 gnd.n5821 gnd.n1631 585
R10218 gnd.n5929 gnd.n5928 585
R10219 gnd.n5928 gnd.n5927 585
R10220 gnd.n5930 gnd.n1626 585
R10221 gnd.n5758 gnd.n1626 585
R10222 gnd.n5932 gnd.n5931 585
R10223 gnd.n5933 gnd.n5932 585
R10224 gnd.n1611 gnd.n1610 585
R10225 gnd.n5749 gnd.n1611 585
R10226 gnd.n5941 gnd.n5940 585
R10227 gnd.n5940 gnd.n5939 585
R10228 gnd.n5942 gnd.n1604 585
R10229 gnd.n5743 gnd.n1604 585
R10230 gnd.n5944 gnd.n5943 585
R10231 gnd.n5945 gnd.n5944 585
R10232 gnd.n1605 gnd.n1603 585
R10233 gnd.n5736 gnd.n1603 585
R10234 gnd.n1587 gnd.n1581 585
R10235 gnd.n5951 gnd.n1587 585
R10236 gnd.n5956 gnd.n1579 585
R10237 gnd.n5775 gnd.n1579 585
R10238 gnd.n5958 gnd.n5957 585
R10239 gnd.n5959 gnd.n5958 585
R10240 gnd.n1578 gnd.n1418 585
R10241 gnd.n6126 gnd.n1419 585
R10242 gnd.n6125 gnd.n1420 585
R10243 gnd.n1495 gnd.n1421 585
R10244 gnd.n6118 gnd.n1427 585
R10245 gnd.n6117 gnd.n1428 585
R10246 gnd.n1498 gnd.n1429 585
R10247 gnd.n6110 gnd.n1435 585
R10248 gnd.n6109 gnd.n1436 585
R10249 gnd.n1500 gnd.n1437 585
R10250 gnd.n6102 gnd.n1443 585
R10251 gnd.n6101 gnd.n1444 585
R10252 gnd.n1503 gnd.n1445 585
R10253 gnd.n6094 gnd.n1451 585
R10254 gnd.n6093 gnd.n1452 585
R10255 gnd.n1505 gnd.n1453 585
R10256 gnd.n6086 gnd.n1461 585
R10257 gnd.n6085 gnd.n6082 585
R10258 gnd.n1464 gnd.n1462 585
R10259 gnd.n6080 gnd.n1464 585
R10260 gnd.n349 gnd.n348 585
R10261 gnd.n7405 gnd.n344 585
R10262 gnd.n7407 gnd.n7406 585
R10263 gnd.n7409 gnd.n342 585
R10264 gnd.n7411 gnd.n7410 585
R10265 gnd.n7412 gnd.n337 585
R10266 gnd.n7414 gnd.n7413 585
R10267 gnd.n7416 gnd.n335 585
R10268 gnd.n7418 gnd.n7417 585
R10269 gnd.n7419 gnd.n330 585
R10270 gnd.n7421 gnd.n7420 585
R10271 gnd.n7423 gnd.n328 585
R10272 gnd.n7425 gnd.n7424 585
R10273 gnd.n7426 gnd.n323 585
R10274 gnd.n7428 gnd.n7427 585
R10275 gnd.n7430 gnd.n321 585
R10276 gnd.n7432 gnd.n7431 585
R10277 gnd.n7433 gnd.n319 585
R10278 gnd.n7434 gnd.n208 585
R10279 gnd.n212 gnd.n208 585
R10280 gnd.n7401 gnd.n211 585
R10281 gnd.n7549 gnd.n211 585
R10282 gnd.n7400 gnd.n7399 585
R10283 gnd.n7399 gnd.n209 585
R10284 gnd.n7398 gnd.n203 585
R10285 gnd.n7555 gnd.n203 585
R10286 gnd.n354 gnd.n353 585
R10287 gnd.n353 gnd.n194 585
R10288 gnd.n7394 gnd.n193 585
R10289 gnd.n7561 gnd.n193 585
R10290 gnd.n7393 gnd.n7392 585
R10291 gnd.n7392 gnd.n191 585
R10292 gnd.n7391 gnd.n183 585
R10293 gnd.n7567 gnd.n183 585
R10294 gnd.n357 gnd.n356 585
R10295 gnd.n356 gnd.n174 585
R10296 gnd.n7387 gnd.n173 585
R10297 gnd.n7573 gnd.n173 585
R10298 gnd.n7386 gnd.n7385 585
R10299 gnd.n7385 gnd.n171 585
R10300 gnd.n7384 gnd.n164 585
R10301 gnd.n7579 gnd.n164 585
R10302 gnd.n360 gnd.n359 585
R10303 gnd.n359 gnd.n162 585
R10304 gnd.n7380 gnd.n154 585
R10305 gnd.n7585 gnd.n154 585
R10306 gnd.n7379 gnd.n7378 585
R10307 gnd.n7378 gnd.n146 585
R10308 gnd.n7377 gnd.n145 585
R10309 gnd.n7591 gnd.n145 585
R10310 gnd.n363 gnd.n362 585
R10311 gnd.n362 gnd.n136 585
R10312 gnd.n7373 gnd.n135 585
R10313 gnd.n7597 gnd.n135 585
R10314 gnd.n7372 gnd.n7371 585
R10315 gnd.n7371 gnd.n133 585
R10316 gnd.n7370 gnd.n126 585
R10317 gnd.n7603 gnd.n126 585
R10318 gnd.n366 gnd.n365 585
R10319 gnd.n365 gnd.n124 585
R10320 gnd.n7366 gnd.n117 585
R10321 gnd.n7609 gnd.n117 585
R10322 gnd.n7365 gnd.n7364 585
R10323 gnd.n7364 gnd.n107 585
R10324 gnd.n7363 gnd.n106 585
R10325 gnd.n7615 gnd.n106 585
R10326 gnd.n7359 gnd.n7358 585
R10327 gnd.n7358 gnd.n7357 585
R10328 gnd.n88 gnd.n87 585
R10329 gnd.n368 gnd.n88 585
R10330 gnd.n7625 gnd.n7624 585
R10331 gnd.n7624 gnd.n7623 585
R10332 gnd.n7626 gnd.n86 585
R10333 gnd.n7308 gnd.n86 585
R10334 gnd.n7294 gnd.n85 585
R10335 gnd.n7295 gnd.n7294 585
R10336 gnd.n5862 gnd.n383 585
R10337 gnd.n7299 gnd.n383 585
R10338 gnd.n5861 gnd.n5860 585
R10339 gnd.n5860 gnd.n1699 585
R10340 gnd.n5866 gnd.n1698 585
R10341 gnd.n5887 gnd.n1698 585
R10342 gnd.n5867 gnd.n1694 585
R10343 gnd.n5891 gnd.n1694 585
R10344 gnd.n5868 gnd.n5859 585
R10345 gnd.n5859 gnd.n5858 585
R10346 gnd.n1708 gnd.n1684 585
R10347 gnd.n5897 gnd.n1684 585
R10348 gnd.n5873 gnd.n5872 585
R10349 gnd.n5874 gnd.n5873 585
R10350 gnd.n1707 gnd.n1674 585
R10351 gnd.n5903 gnd.n1674 585
R10352 gnd.n5843 gnd.n5842 585
R10353 gnd.n5844 gnd.n5843 585
R10354 gnd.n1712 gnd.n1664 585
R10355 gnd.n5909 gnd.n1664 585
R10356 gnd.n5838 gnd.n5837 585
R10357 gnd.n5837 gnd.n5836 585
R10358 gnd.n1714 gnd.n1654 585
R10359 gnd.n5915 gnd.n1654 585
R10360 gnd.n5828 gnd.n5827 585
R10361 gnd.n5829 gnd.n5828 585
R10362 gnd.n1717 gnd.n1644 585
R10363 gnd.n5921 gnd.n1644 585
R10364 gnd.n5823 gnd.n5822 585
R10365 gnd.n5822 gnd.n5821 585
R10366 gnd.n1719 gnd.n1634 585
R10367 gnd.n5927 gnd.n1634 585
R10368 gnd.n5761 gnd.n5759 585
R10369 gnd.n5759 gnd.n5758 585
R10370 gnd.n5762 gnd.n1624 585
R10371 gnd.n5933 gnd.n1624 585
R10372 gnd.n5763 gnd.n5741 585
R10373 gnd.n5749 gnd.n5741 585
R10374 gnd.n5739 gnd.n1614 585
R10375 gnd.n5939 gnd.n1614 585
R10376 gnd.n5767 gnd.n5738 585
R10377 gnd.n5743 gnd.n5738 585
R10378 gnd.n5768 gnd.n1601 585
R10379 gnd.n5945 gnd.n1601 585
R10380 gnd.n5769 gnd.n5737 585
R10381 gnd.n5737 gnd.n5736 585
R10382 gnd.n1736 gnd.n1585 585
R10383 gnd.n5951 gnd.n1585 585
R10384 gnd.n5774 gnd.n5773 585
R10385 gnd.n5775 gnd.n5774 585
R10386 gnd.n1735 gnd.n1576 585
R10387 gnd.n5959 gnd.n1576 585
R10388 gnd.n4022 gnd.n2672 585
R10389 gnd.n2672 gnd.n2649 585
R10390 gnd.n4023 gnd.n2733 585
R10391 gnd.n2733 gnd.n2723 585
R10392 gnd.n4025 gnd.n4024 585
R10393 gnd.n4026 gnd.n4025 585
R10394 gnd.n2734 gnd.n2732 585
R10395 gnd.n2741 gnd.n2732 585
R10396 gnd.n4016 gnd.n4015 585
R10397 gnd.n4015 gnd.n4014 585
R10398 gnd.n2737 gnd.n2736 585
R10399 gnd.n3741 gnd.n2737 585
R10400 gnd.n3726 gnd.n2760 585
R10401 gnd.n2760 gnd.n2750 585
R10402 gnd.n3728 gnd.n3727 585
R10403 gnd.n3729 gnd.n3728 585
R10404 gnd.n2761 gnd.n2759 585
R10405 gnd.n2759 gnd.n2757 585
R10406 gnd.n3721 gnd.n3720 585
R10407 gnd.n3720 gnd.n3719 585
R10408 gnd.n2764 gnd.n2763 585
R10409 gnd.n2773 gnd.n2764 585
R10410 gnd.n3677 gnd.n2787 585
R10411 gnd.n2787 gnd.n2772 585
R10412 gnd.n3679 gnd.n3678 585
R10413 gnd.n3680 gnd.n3679 585
R10414 gnd.n2788 gnd.n2786 585
R10415 gnd.n2795 gnd.n2786 585
R10416 gnd.n3672 gnd.n3671 585
R10417 gnd.n3671 gnd.n3670 585
R10418 gnd.n2791 gnd.n2790 585
R10419 gnd.n3651 gnd.n2791 585
R10420 gnd.n3637 gnd.n2815 585
R10421 gnd.n2815 gnd.n2804 585
R10422 gnd.n3639 gnd.n3638 585
R10423 gnd.n3640 gnd.n3639 585
R10424 gnd.n2816 gnd.n2814 585
R10425 gnd.n2814 gnd.n2811 585
R10426 gnd.n3632 gnd.n3631 585
R10427 gnd.n3631 gnd.n3630 585
R10428 gnd.n2819 gnd.n2818 585
R10429 gnd.n2829 gnd.n2819 585
R10430 gnd.n3592 gnd.n2842 585
R10431 gnd.n2842 gnd.n2828 585
R10432 gnd.n3594 gnd.n3593 585
R10433 gnd.n3595 gnd.n3594 585
R10434 gnd.n2843 gnd.n2841 585
R10435 gnd.n2850 gnd.n2841 585
R10436 gnd.n3587 gnd.n3586 585
R10437 gnd.n3586 gnd.n3585 585
R10438 gnd.n2846 gnd.n2845 585
R10439 gnd.n3566 gnd.n2846 585
R10440 gnd.n3552 gnd.n2869 585
R10441 gnd.n2869 gnd.n2859 585
R10442 gnd.n3554 gnd.n3553 585
R10443 gnd.n3555 gnd.n3554 585
R10444 gnd.n2870 gnd.n2868 585
R10445 gnd.n3543 gnd.n2868 585
R10446 gnd.n3547 gnd.n3546 585
R10447 gnd.n3546 gnd.n3545 585
R10448 gnd.n2873 gnd.n2872 585
R10449 gnd.n3498 gnd.n2873 585
R10450 gnd.n2991 gnd.n2990 585
R10451 gnd.n2992 gnd.n2991 585
R10452 gnd.n2971 gnd.n2970 585
R10453 gnd.n2974 gnd.n2971 585
R10454 gnd.n3508 gnd.n3507 585
R10455 gnd.n3507 gnd.n3506 585
R10456 gnd.n3509 gnd.n2965 585
R10457 gnd.n3001 gnd.n2965 585
R10458 gnd.n3511 gnd.n3510 585
R10459 gnd.n3512 gnd.n3511 585
R10460 gnd.n2966 gnd.n2964 585
R10461 gnd.n3476 gnd.n2964 585
R10462 gnd.n3460 gnd.n3459 585
R10463 gnd.n3459 gnd.n2952 585
R10464 gnd.n3461 gnd.n3016 585
R10465 gnd.n3016 gnd.n2951 585
R10466 gnd.n3463 gnd.n3462 585
R10467 gnd.n3464 gnd.n3463 585
R10468 gnd.n3017 gnd.n3015 585
R10469 gnd.n3015 gnd.n3012 585
R10470 gnd.n3452 gnd.n3451 585
R10471 gnd.n3451 gnd.n3450 585
R10472 gnd.n3020 gnd.n3019 585
R10473 gnd.n3027 gnd.n3020 585
R10474 gnd.n3426 gnd.n3425 585
R10475 gnd.n3427 gnd.n3426 585
R10476 gnd.n3039 gnd.n3038 585
R10477 gnd.n3046 gnd.n3038 585
R10478 gnd.n3421 gnd.n3420 585
R10479 gnd.n3420 gnd.n3419 585
R10480 gnd.n3042 gnd.n3041 585
R10481 gnd.n3409 gnd.n3042 585
R10482 gnd.n3396 gnd.n3066 585
R10483 gnd.n3066 gnd.n3065 585
R10484 gnd.n3398 gnd.n3397 585
R10485 gnd.n3399 gnd.n3398 585
R10486 gnd.n3067 gnd.n3064 585
R10487 gnd.n3074 gnd.n3064 585
R10488 gnd.n3391 gnd.n3390 585
R10489 gnd.n3390 gnd.n3389 585
R10490 gnd.n3070 gnd.n3069 585
R10491 gnd.n3378 gnd.n3070 585
R10492 gnd.n3365 gnd.n3091 585
R10493 gnd.n3091 gnd.n3090 585
R10494 gnd.n3367 gnd.n3366 585
R10495 gnd.n3368 gnd.n3367 585
R10496 gnd.n3361 gnd.n3089 585
R10497 gnd.n3360 gnd.n3359 585
R10498 gnd.n3094 gnd.n3093 585
R10499 gnd.n3357 gnd.n3094 585
R10500 gnd.n3116 gnd.n3115 585
R10501 gnd.n3119 gnd.n3118 585
R10502 gnd.n3117 gnd.n3112 585
R10503 gnd.n3124 gnd.n3123 585
R10504 gnd.n3126 gnd.n3125 585
R10505 gnd.n3129 gnd.n3128 585
R10506 gnd.n3127 gnd.n3110 585
R10507 gnd.n3134 gnd.n3133 585
R10508 gnd.n3136 gnd.n3135 585
R10509 gnd.n3139 gnd.n3138 585
R10510 gnd.n3137 gnd.n3108 585
R10511 gnd.n3144 gnd.n3143 585
R10512 gnd.n3148 gnd.n3145 585
R10513 gnd.n3149 gnd.n3086 585
R10514 gnd.n4028 gnd.n2687 585
R10515 gnd.n4095 gnd.n4094 585
R10516 gnd.n4097 gnd.n4096 585
R10517 gnd.n4099 gnd.n4098 585
R10518 gnd.n4101 gnd.n4100 585
R10519 gnd.n4103 gnd.n4102 585
R10520 gnd.n4105 gnd.n4104 585
R10521 gnd.n4107 gnd.n4106 585
R10522 gnd.n4109 gnd.n4108 585
R10523 gnd.n4111 gnd.n4110 585
R10524 gnd.n4113 gnd.n4112 585
R10525 gnd.n4115 gnd.n4114 585
R10526 gnd.n4117 gnd.n4116 585
R10527 gnd.n4120 gnd.n4119 585
R10528 gnd.n4118 gnd.n2675 585
R10529 gnd.n4124 gnd.n2673 585
R10530 gnd.n4126 gnd.n4125 585
R10531 gnd.n4127 gnd.n4126 585
R10532 gnd.n4029 gnd.n2728 585
R10533 gnd.n4029 gnd.n2649 585
R10534 gnd.n4031 gnd.n4030 585
R10535 gnd.n4030 gnd.n2723 585
R10536 gnd.n4027 gnd.n2727 585
R10537 gnd.n4027 gnd.n4026 585
R10538 gnd.n4006 gnd.n2729 585
R10539 gnd.n2741 gnd.n2729 585
R10540 gnd.n4005 gnd.n2739 585
R10541 gnd.n4014 gnd.n2739 585
R10542 gnd.n3739 gnd.n2746 585
R10543 gnd.n3741 gnd.n3739 585
R10544 gnd.n3738 gnd.n3737 585
R10545 gnd.n3738 gnd.n2750 585
R10546 gnd.n3736 gnd.n2752 585
R10547 gnd.n3729 gnd.n2752 585
R10548 gnd.n2765 gnd.n2753 585
R10549 gnd.n2765 gnd.n2757 585
R10550 gnd.n3685 gnd.n2766 585
R10551 gnd.n3719 gnd.n2766 585
R10552 gnd.n3684 gnd.n3683 585
R10553 gnd.n3683 gnd.n2773 585
R10554 gnd.n3682 gnd.n2781 585
R10555 gnd.n3682 gnd.n2772 585
R10556 gnd.n3681 gnd.n2783 585
R10557 gnd.n3681 gnd.n3680 585
R10558 gnd.n3660 gnd.n2782 585
R10559 gnd.n2795 gnd.n2782 585
R10560 gnd.n3659 gnd.n2793 585
R10561 gnd.n3670 gnd.n2793 585
R10562 gnd.n3650 gnd.n2800 585
R10563 gnd.n3651 gnd.n3650 585
R10564 gnd.n3649 gnd.n3648 585
R10565 gnd.n3649 gnd.n2804 585
R10566 gnd.n3647 gnd.n2806 585
R10567 gnd.n3640 gnd.n2806 585
R10568 gnd.n2821 gnd.n2807 585
R10569 gnd.n2821 gnd.n2811 585
R10570 gnd.n3600 gnd.n2822 585
R10571 gnd.n3630 gnd.n2822 585
R10572 gnd.n3599 gnd.n3598 585
R10573 gnd.n3598 gnd.n2829 585
R10574 gnd.n3597 gnd.n2836 585
R10575 gnd.n3597 gnd.n2828 585
R10576 gnd.n3596 gnd.n2838 585
R10577 gnd.n3596 gnd.n3595 585
R10578 gnd.n3575 gnd.n2837 585
R10579 gnd.n2850 gnd.n2837 585
R10580 gnd.n3574 gnd.n2848 585
R10581 gnd.n3585 gnd.n2848 585
R10582 gnd.n3565 gnd.n2855 585
R10583 gnd.n3566 gnd.n3565 585
R10584 gnd.n3564 gnd.n3563 585
R10585 gnd.n3564 gnd.n2859 585
R10586 gnd.n3562 gnd.n2861 585
R10587 gnd.n3555 gnd.n2861 585
R10588 gnd.n3542 gnd.n2862 585
R10589 gnd.n3543 gnd.n3542 585
R10590 gnd.n3495 gnd.n2875 585
R10591 gnd.n3545 gnd.n2875 585
R10592 gnd.n3497 gnd.n3496 585
R10593 gnd.n3498 gnd.n3497 585
R10594 gnd.n3490 gnd.n2993 585
R10595 gnd.n2993 gnd.n2992 585
R10596 gnd.n3488 gnd.n3487 585
R10597 gnd.n3487 gnd.n2974 585
R10598 gnd.n3485 gnd.n2972 585
R10599 gnd.n3506 gnd.n2972 585
R10600 gnd.n3003 gnd.n3002 585
R10601 gnd.n3002 gnd.n3001 585
R10602 gnd.n3479 gnd.n2962 585
R10603 gnd.n3512 gnd.n2962 585
R10604 gnd.n3478 gnd.n3477 585
R10605 gnd.n3477 gnd.n3476 585
R10606 gnd.n3474 gnd.n3005 585
R10607 gnd.n3474 gnd.n2952 585
R10608 gnd.n3473 gnd.n3472 585
R10609 gnd.n3473 gnd.n2951 585
R10610 gnd.n3008 gnd.n3007 585
R10611 gnd.n3464 gnd.n3007 585
R10612 gnd.n3432 gnd.n3431 585
R10613 gnd.n3431 gnd.n3012 585
R10614 gnd.n3433 gnd.n3021 585
R10615 gnd.n3450 gnd.n3021 585
R10616 gnd.n3430 gnd.n3429 585
R10617 gnd.n3429 gnd.n3027 585
R10618 gnd.n3428 gnd.n3035 585
R10619 gnd.n3428 gnd.n3427 585
R10620 gnd.n3413 gnd.n3036 585
R10621 gnd.n3046 gnd.n3036 585
R10622 gnd.n3412 gnd.n3044 585
R10623 gnd.n3419 gnd.n3044 585
R10624 gnd.n3411 gnd.n3410 585
R10625 gnd.n3410 gnd.n3409 585
R10626 gnd.n3055 gnd.n3052 585
R10627 gnd.n3065 gnd.n3055 585
R10628 gnd.n3401 gnd.n3400 585
R10629 gnd.n3400 gnd.n3399 585
R10630 gnd.n3061 gnd.n3060 585
R10631 gnd.n3074 gnd.n3061 585
R10632 gnd.n3381 gnd.n3072 585
R10633 gnd.n3389 gnd.n3072 585
R10634 gnd.n3380 gnd.n3379 585
R10635 gnd.n3379 gnd.n3378 585
R10636 gnd.n3081 gnd.n3079 585
R10637 gnd.n3090 gnd.n3081 585
R10638 gnd.n3370 gnd.n3369 585
R10639 gnd.n3369 gnd.n3368 585
R10640 gnd.n5543 gnd.n1874 585
R10641 gnd.n1874 gnd.n1830 585
R10642 gnd.n5545 gnd.n5544 585
R10643 gnd.n5546 gnd.n5545 585
R10644 gnd.n5454 gnd.n1873 585
R10645 gnd.n1880 gnd.n1873 585
R10646 gnd.n5453 gnd.n5452 585
R10647 gnd.n5452 gnd.n5451 585
R10648 gnd.n1876 gnd.n1875 585
R10649 gnd.n1877 gnd.n1876 585
R10650 gnd.n5439 gnd.n5438 585
R10651 gnd.n5440 gnd.n5439 585
R10652 gnd.n5437 gnd.n1889 585
R10653 gnd.n1889 gnd.n1886 585
R10654 gnd.n5436 gnd.n5435 585
R10655 gnd.n5435 gnd.n5434 585
R10656 gnd.n1891 gnd.n1890 585
R10657 gnd.n5371 gnd.n1891 585
R10658 gnd.n5397 gnd.n5396 585
R10659 gnd.n5397 gnd.n1900 585
R10660 gnd.n5399 gnd.n5398 585
R10661 gnd.n5398 gnd.n1899 585
R10662 gnd.n5400 gnd.n1913 585
R10663 gnd.n5385 gnd.n1913 585
R10664 gnd.n5402 gnd.n5401 585
R10665 gnd.n5403 gnd.n5402 585
R10666 gnd.n5395 gnd.n1912 585
R10667 gnd.n1912 gnd.n1907 585
R10668 gnd.n5394 gnd.n5393 585
R10669 gnd.n5393 gnd.n5392 585
R10670 gnd.n1915 gnd.n1914 585
R10671 gnd.n5278 gnd.n1915 585
R10672 gnd.n5364 gnd.n5363 585
R10673 gnd.n5365 gnd.n5364 585
R10674 gnd.n5362 gnd.n1922 585
R10675 gnd.n1922 gnd.n1920 585
R10676 gnd.n5361 gnd.n5360 585
R10677 gnd.n5360 gnd.n5359 585
R10678 gnd.n1924 gnd.n1923 585
R10679 gnd.n1937 gnd.n1924 585
R10680 gnd.n5346 gnd.n5345 585
R10681 gnd.n5347 gnd.n5346 585
R10682 gnd.n5344 gnd.n1938 585
R10683 gnd.n5339 gnd.n1938 585
R10684 gnd.n5343 gnd.n5342 585
R10685 gnd.n5342 gnd.n5341 585
R10686 gnd.n1940 gnd.n1939 585
R10687 gnd.n1941 gnd.n1940 585
R10688 gnd.n5327 gnd.n5326 585
R10689 gnd.n5328 gnd.n5327 585
R10690 gnd.n5325 gnd.n1946 585
R10691 gnd.n5321 gnd.n1946 585
R10692 gnd.n5324 gnd.n5323 585
R10693 gnd.n5323 gnd.n5322 585
R10694 gnd.n1948 gnd.n1947 585
R10695 gnd.n5309 gnd.n1948 585
R10696 gnd.n1986 gnd.n1985 585
R10697 gnd.n1985 gnd.n1958 585
R10698 gnd.n1987 gnd.n1963 585
R10699 gnd.n5301 gnd.n1963 585
R10700 gnd.n1989 gnd.n1988 585
R10701 gnd.n5241 gnd.n1989 585
R10702 gnd.n5244 gnd.n1984 585
R10703 gnd.n5244 gnd.n5243 585
R10704 gnd.n5246 gnd.n5245 585
R10705 gnd.n5245 gnd.n1970 585
R10706 gnd.n5247 gnd.n1982 585
R10707 gnd.n5235 gnd.n1982 585
R10708 gnd.n5249 gnd.n5248 585
R10709 gnd.n5250 gnd.n5249 585
R10710 gnd.n1983 gnd.n1981 585
R10711 gnd.n1981 gnd.n1977 585
R10712 gnd.n5229 gnd.n5228 585
R10713 gnd.n5230 gnd.n5229 585
R10714 gnd.n5227 gnd.n1994 585
R10715 gnd.n1999 gnd.n1994 585
R10716 gnd.n5226 gnd.n5225 585
R10717 gnd.n5225 gnd.n5224 585
R10718 gnd.n1996 gnd.n1995 585
R10719 gnd.n5200 gnd.n1996 585
R10720 gnd.n5212 gnd.n5211 585
R10721 gnd.n5213 gnd.n5212 585
R10722 gnd.n5210 gnd.n2009 585
R10723 gnd.n2009 gnd.n2005 585
R10724 gnd.n5209 gnd.n5208 585
R10725 gnd.n5208 gnd.n5207 585
R10726 gnd.n2011 gnd.n2010 585
R10727 gnd.n2017 gnd.n2011 585
R10728 gnd.n5193 gnd.n5192 585
R10729 gnd.n5194 gnd.n5193 585
R10730 gnd.n5191 gnd.n2019 585
R10731 gnd.n2026 gnd.n2019 585
R10732 gnd.n5190 gnd.n5189 585
R10733 gnd.n5189 gnd.n5188 585
R10734 gnd.n2021 gnd.n2020 585
R10735 gnd.n5065 gnd.n2021 585
R10736 gnd.n5175 gnd.n5174 585
R10737 gnd.n5176 gnd.n5175 585
R10738 gnd.n5173 gnd.n2036 585
R10739 gnd.n2036 gnd.n2033 585
R10740 gnd.n5172 gnd.n5171 585
R10741 gnd.n5171 gnd.n5170 585
R10742 gnd.n2038 gnd.n2037 585
R10743 gnd.n5062 gnd.n2038 585
R10744 gnd.n5120 gnd.n5119 585
R10745 gnd.n5120 gnd.n2047 585
R10746 gnd.n5122 gnd.n5121 585
R10747 gnd.n5121 gnd.n2046 585
R10748 gnd.n5123 gnd.n2060 585
R10749 gnd.n2060 gnd.n2058 585
R10750 gnd.n5125 gnd.n5124 585
R10751 gnd.n5126 gnd.n5125 585
R10752 gnd.n5118 gnd.n2059 585
R10753 gnd.n2059 gnd.n2055 585
R10754 gnd.n5117 gnd.n5116 585
R10755 gnd.n5116 gnd.n5115 585
R10756 gnd.n2062 gnd.n2061 585
R10757 gnd.n2063 gnd.n2062 585
R10758 gnd.n5088 gnd.n2085 585
R10759 gnd.n5088 gnd.n5087 585
R10760 gnd.n5090 gnd.n5089 585
R10761 gnd.n5089 gnd.n2071 585
R10762 gnd.n5091 gnd.n2083 585
R10763 gnd.n5056 gnd.n2083 585
R10764 gnd.n5093 gnd.n5092 585
R10765 gnd.n5094 gnd.n5093 585
R10766 gnd.n2084 gnd.n2082 585
R10767 gnd.n2082 gnd.n2078 585
R10768 gnd.n5050 gnd.n5049 585
R10769 gnd.n5051 gnd.n5050 585
R10770 gnd.n5048 gnd.n2092 585
R10771 gnd.n2098 gnd.n2092 585
R10772 gnd.n5047 gnd.n5046 585
R10773 gnd.n5046 gnd.n5045 585
R10774 gnd.n2094 gnd.n2093 585
R10775 gnd.n2095 gnd.n2094 585
R10776 gnd.n5034 gnd.n5033 585
R10777 gnd.n5035 gnd.n5034 585
R10778 gnd.n5032 gnd.n2105 585
R10779 gnd.n5028 gnd.n2105 585
R10780 gnd.n5031 gnd.n5030 585
R10781 gnd.n5030 gnd.n5029 585
R10782 gnd.n2107 gnd.n2106 585
R10783 gnd.n2107 gnd.n1302 585
R10784 gnd.n5015 gnd.n5014 585
R10785 gnd.n5016 gnd.n5015 585
R10786 gnd.n5013 gnd.n5012 585
R10787 gnd.n5012 gnd.n5011 585
R10788 gnd.n1285 gnd.n1284 585
R10789 gnd.n1289 gnd.n1285 585
R10790 gnd.n6268 gnd.n6267 585
R10791 gnd.n6267 gnd.n6266 585
R10792 gnd.n6269 gnd.n1279 585
R10793 gnd.n1286 gnd.n1279 585
R10794 gnd.n6271 gnd.n6270 585
R10795 gnd.n6272 gnd.n6271 585
R10796 gnd.n1283 gnd.n1278 585
R10797 gnd.n1278 gnd.n1277 585
R10798 gnd.n1282 gnd.n1197 585
R10799 gnd.n6278 gnd.n1197 585
R10800 gnd.n1281 gnd.n1280 585
R10801 gnd.n1280 gnd.n1196 585
R10802 gnd.n1182 gnd.n1181 585
R10803 gnd.n1186 gnd.n1182 585
R10804 gnd.n6287 gnd.n6286 585
R10805 gnd.n6286 gnd.n6285 585
R10806 gnd.n6288 gnd.n1160 585
R10807 gnd.n1183 gnd.n1160 585
R10808 gnd.n6353 gnd.n6352 585
R10809 gnd.n6351 gnd.n1159 585
R10810 gnd.n6350 gnd.n1158 585
R10811 gnd.n6355 gnd.n1158 585
R10812 gnd.n6349 gnd.n6348 585
R10813 gnd.n6347 gnd.n6346 585
R10814 gnd.n6345 gnd.n6344 585
R10815 gnd.n6343 gnd.n6342 585
R10816 gnd.n6341 gnd.n6340 585
R10817 gnd.n6339 gnd.n6338 585
R10818 gnd.n6337 gnd.n6336 585
R10819 gnd.n6335 gnd.n6334 585
R10820 gnd.n6333 gnd.n6332 585
R10821 gnd.n6331 gnd.n6330 585
R10822 gnd.n6329 gnd.n6328 585
R10823 gnd.n6327 gnd.n6326 585
R10824 gnd.n6325 gnd.n6324 585
R10825 gnd.n6323 gnd.n6322 585
R10826 gnd.n6321 gnd.n6320 585
R10827 gnd.n6319 gnd.n6318 585
R10828 gnd.n6317 gnd.n6316 585
R10829 gnd.n6315 gnd.n6314 585
R10830 gnd.n6313 gnd.n6312 585
R10831 gnd.n6311 gnd.n6310 585
R10832 gnd.n6309 gnd.n6308 585
R10833 gnd.n6307 gnd.n6306 585
R10834 gnd.n6305 gnd.n6304 585
R10835 gnd.n6303 gnd.n6302 585
R10836 gnd.n6301 gnd.n6300 585
R10837 gnd.n6299 gnd.n6298 585
R10838 gnd.n6297 gnd.n6296 585
R10839 gnd.n6295 gnd.n6294 585
R10840 gnd.n6293 gnd.n1122 585
R10841 gnd.n6358 gnd.n6357 585
R10842 gnd.n1124 gnd.n1121 585
R10843 gnd.n1205 gnd.n1204 585
R10844 gnd.n1207 gnd.n1206 585
R10845 gnd.n1210 gnd.n1209 585
R10846 gnd.n1212 gnd.n1211 585
R10847 gnd.n1214 gnd.n1213 585
R10848 gnd.n1216 gnd.n1215 585
R10849 gnd.n1218 gnd.n1217 585
R10850 gnd.n1220 gnd.n1219 585
R10851 gnd.n1222 gnd.n1221 585
R10852 gnd.n1224 gnd.n1223 585
R10853 gnd.n1226 gnd.n1225 585
R10854 gnd.n1228 gnd.n1227 585
R10855 gnd.n1230 gnd.n1229 585
R10856 gnd.n1232 gnd.n1231 585
R10857 gnd.n1234 gnd.n1233 585
R10858 gnd.n1236 gnd.n1235 585
R10859 gnd.n1238 gnd.n1237 585
R10860 gnd.n1240 gnd.n1239 585
R10861 gnd.n1242 gnd.n1241 585
R10862 gnd.n1244 gnd.n1243 585
R10863 gnd.n1246 gnd.n1245 585
R10864 gnd.n1248 gnd.n1247 585
R10865 gnd.n1250 gnd.n1249 585
R10866 gnd.n1252 gnd.n1251 585
R10867 gnd.n1254 gnd.n1253 585
R10868 gnd.n1256 gnd.n1255 585
R10869 gnd.n1258 gnd.n1257 585
R10870 gnd.n1260 gnd.n1259 585
R10871 gnd.n1262 gnd.n1261 585
R10872 gnd.n1264 gnd.n1263 585
R10873 gnd.n1266 gnd.n1265 585
R10874 gnd.n5550 gnd.n5549 585
R10875 gnd.n5552 gnd.n5551 585
R10876 gnd.n5554 gnd.n5553 585
R10877 gnd.n5556 gnd.n5555 585
R10878 gnd.n5558 gnd.n5557 585
R10879 gnd.n5560 gnd.n5559 585
R10880 gnd.n5562 gnd.n5561 585
R10881 gnd.n5564 gnd.n5563 585
R10882 gnd.n5566 gnd.n5565 585
R10883 gnd.n5568 gnd.n5567 585
R10884 gnd.n5570 gnd.n5569 585
R10885 gnd.n5572 gnd.n5571 585
R10886 gnd.n5574 gnd.n5573 585
R10887 gnd.n5576 gnd.n5575 585
R10888 gnd.n5578 gnd.n5577 585
R10889 gnd.n5580 gnd.n5579 585
R10890 gnd.n5582 gnd.n5581 585
R10891 gnd.n5584 gnd.n5583 585
R10892 gnd.n5586 gnd.n5585 585
R10893 gnd.n5588 gnd.n5587 585
R10894 gnd.n5590 gnd.n5589 585
R10895 gnd.n5592 gnd.n5591 585
R10896 gnd.n5594 gnd.n5593 585
R10897 gnd.n5596 gnd.n5595 585
R10898 gnd.n5598 gnd.n5597 585
R10899 gnd.n5600 gnd.n5599 585
R10900 gnd.n5602 gnd.n5601 585
R10901 gnd.n5604 gnd.n5603 585
R10902 gnd.n5606 gnd.n5605 585
R10903 gnd.n5609 gnd.n5608 585
R10904 gnd.n5611 gnd.n5610 585
R10905 gnd.n5613 gnd.n5612 585
R10906 gnd.n5615 gnd.n5614 585
R10907 gnd.n5476 gnd.n1539 585
R10908 gnd.n5478 gnd.n5477 585
R10909 gnd.n5480 gnd.n5479 585
R10910 gnd.n5482 gnd.n5481 585
R10911 gnd.n5485 gnd.n5484 585
R10912 gnd.n5487 gnd.n5486 585
R10913 gnd.n5489 gnd.n5488 585
R10914 gnd.n5491 gnd.n5490 585
R10915 gnd.n5493 gnd.n5492 585
R10916 gnd.n5495 gnd.n5494 585
R10917 gnd.n5497 gnd.n5496 585
R10918 gnd.n5499 gnd.n5498 585
R10919 gnd.n5501 gnd.n5500 585
R10920 gnd.n5503 gnd.n5502 585
R10921 gnd.n5505 gnd.n5504 585
R10922 gnd.n5507 gnd.n5506 585
R10923 gnd.n5509 gnd.n5508 585
R10924 gnd.n5511 gnd.n5510 585
R10925 gnd.n5513 gnd.n5512 585
R10926 gnd.n5515 gnd.n5514 585
R10927 gnd.n5517 gnd.n5516 585
R10928 gnd.n5519 gnd.n5518 585
R10929 gnd.n5521 gnd.n5520 585
R10930 gnd.n5523 gnd.n5522 585
R10931 gnd.n5525 gnd.n5524 585
R10932 gnd.n5527 gnd.n5526 585
R10933 gnd.n5529 gnd.n5528 585
R10934 gnd.n5531 gnd.n5530 585
R10935 gnd.n5533 gnd.n5532 585
R10936 gnd.n5535 gnd.n5534 585
R10937 gnd.n5537 gnd.n5536 585
R10938 gnd.n5539 gnd.n5538 585
R10939 gnd.n5541 gnd.n5540 585
R10940 gnd.n5548 gnd.n1869 585
R10941 gnd.n5548 gnd.n1830 585
R10942 gnd.n5547 gnd.n1871 585
R10943 gnd.n5547 gnd.n5546 585
R10944 gnd.n5373 gnd.n1870 585
R10945 gnd.n1880 gnd.n1870 585
R10946 gnd.n5374 gnd.n1878 585
R10947 gnd.n5451 gnd.n1878 585
R10948 gnd.n5376 gnd.n5375 585
R10949 gnd.n5375 gnd.n1877 585
R10950 gnd.n5377 gnd.n1888 585
R10951 gnd.n5440 gnd.n1888 585
R10952 gnd.n5379 gnd.n5378 585
R10953 gnd.n5378 gnd.n1886 585
R10954 gnd.n5380 gnd.n1892 585
R10955 gnd.n5434 gnd.n1892 585
R10956 gnd.n5381 gnd.n5372 585
R10957 gnd.n5372 gnd.n5371 585
R10958 gnd.n5383 gnd.n5382 585
R10959 gnd.n5383 gnd.n1900 585
R10960 gnd.n5384 gnd.n5369 585
R10961 gnd.n5384 gnd.n1899 585
R10962 gnd.n5387 gnd.n5386 585
R10963 gnd.n5386 gnd.n5385 585
R10964 gnd.n5388 gnd.n1909 585
R10965 gnd.n5403 gnd.n1909 585
R10966 gnd.n5389 gnd.n1917 585
R10967 gnd.n1917 gnd.n1907 585
R10968 gnd.n5391 gnd.n5390 585
R10969 gnd.n5392 gnd.n5391 585
R10970 gnd.n5368 gnd.n1916 585
R10971 gnd.n5278 gnd.n1916 585
R10972 gnd.n5367 gnd.n5366 585
R10973 gnd.n5366 gnd.n5365 585
R10974 gnd.n1919 gnd.n1918 585
R10975 gnd.n1920 gnd.n1919 585
R10976 gnd.n5333 gnd.n1926 585
R10977 gnd.n5359 gnd.n1926 585
R10978 gnd.n5335 gnd.n5334 585
R10979 gnd.n5334 gnd.n1937 585
R10980 gnd.n5336 gnd.n1936 585
R10981 gnd.n5347 gnd.n1936 585
R10982 gnd.n5338 gnd.n5337 585
R10983 gnd.n5339 gnd.n5338 585
R10984 gnd.n5332 gnd.n1942 585
R10985 gnd.n5341 gnd.n1942 585
R10986 gnd.n5331 gnd.n5330 585
R10987 gnd.n5330 gnd.n1941 585
R10988 gnd.n5329 gnd.n1944 585
R10989 gnd.n5329 gnd.n5328 585
R10990 gnd.n5305 gnd.n1945 585
R10991 gnd.n5321 gnd.n1945 585
R10992 gnd.n5306 gnd.n1950 585
R10993 gnd.n5322 gnd.n1950 585
R10994 gnd.n5308 gnd.n5307 585
R10995 gnd.n5309 gnd.n5308 585
R10996 gnd.n5304 gnd.n1960 585
R10997 gnd.n1960 gnd.n1958 585
R10998 gnd.n5303 gnd.n5302 585
R10999 gnd.n5302 gnd.n5301 585
R11000 gnd.n1962 gnd.n1961 585
R11001 gnd.n5241 gnd.n1962 585
R11002 gnd.n5240 gnd.n5239 585
R11003 gnd.n5243 gnd.n5240 585
R11004 gnd.n5238 gnd.n1990 585
R11005 gnd.n1990 gnd.n1970 585
R11006 gnd.n5237 gnd.n5236 585
R11007 gnd.n5236 gnd.n5235 585
R11008 gnd.n5234 gnd.n1979 585
R11009 gnd.n5250 gnd.n1979 585
R11010 gnd.n5233 gnd.n5232 585
R11011 gnd.n5232 gnd.n1977 585
R11012 gnd.n5231 gnd.n1991 585
R11013 gnd.n5231 gnd.n5230 585
R11014 gnd.n5198 gnd.n1992 585
R11015 gnd.n1999 gnd.n1992 585
R11016 gnd.n5199 gnd.n1997 585
R11017 gnd.n5224 gnd.n1997 585
R11018 gnd.n5202 gnd.n5201 585
R11019 gnd.n5201 gnd.n5200 585
R11020 gnd.n5203 gnd.n2007 585
R11021 gnd.n5213 gnd.n2007 585
R11022 gnd.n5204 gnd.n2014 585
R11023 gnd.n2014 gnd.n2005 585
R11024 gnd.n5206 gnd.n5205 585
R11025 gnd.n5207 gnd.n5206 585
R11026 gnd.n5197 gnd.n2013 585
R11027 gnd.n2017 gnd.n2013 585
R11028 gnd.n5196 gnd.n5195 585
R11029 gnd.n5195 gnd.n5194 585
R11030 gnd.n2016 gnd.n2015 585
R11031 gnd.n2026 gnd.n2016 585
R11032 gnd.n5064 gnd.n2024 585
R11033 gnd.n5188 gnd.n2024 585
R11034 gnd.n5067 gnd.n5066 585
R11035 gnd.n5066 gnd.n5065 585
R11036 gnd.n5068 gnd.n2035 585
R11037 gnd.n5176 gnd.n2035 585
R11038 gnd.n5070 gnd.n5069 585
R11039 gnd.n5069 gnd.n2033 585
R11040 gnd.n5071 gnd.n2039 585
R11041 gnd.n5170 gnd.n2039 585
R11042 gnd.n5072 gnd.n5063 585
R11043 gnd.n5063 gnd.n5062 585
R11044 gnd.n5074 gnd.n5073 585
R11045 gnd.n5074 gnd.n2047 585
R11046 gnd.n5075 gnd.n5060 585
R11047 gnd.n5075 gnd.n2046 585
R11048 gnd.n5077 gnd.n5076 585
R11049 gnd.n5076 gnd.n2058 585
R11050 gnd.n5078 gnd.n2057 585
R11051 gnd.n5126 gnd.n2057 585
R11052 gnd.n5080 gnd.n5079 585
R11053 gnd.n5079 gnd.n2055 585
R11054 gnd.n5081 gnd.n2064 585
R11055 gnd.n5115 gnd.n2064 585
R11056 gnd.n5082 gnd.n2087 585
R11057 gnd.n2087 gnd.n2063 585
R11058 gnd.n5084 gnd.n5083 585
R11059 gnd.n5087 gnd.n5084 585
R11060 gnd.n5059 gnd.n2086 585
R11061 gnd.n2086 gnd.n2071 585
R11062 gnd.n5058 gnd.n5057 585
R11063 gnd.n5057 gnd.n5056 585
R11064 gnd.n5055 gnd.n2080 585
R11065 gnd.n5094 gnd.n2080 585
R11066 gnd.n5054 gnd.n5053 585
R11067 gnd.n5053 gnd.n2078 585
R11068 gnd.n5052 gnd.n2088 585
R11069 gnd.n5052 gnd.n5051 585
R11070 gnd.n5021 gnd.n2089 585
R11071 gnd.n2098 gnd.n2089 585
R11072 gnd.n5022 gnd.n2096 585
R11073 gnd.n5045 gnd.n2096 585
R11074 gnd.n5024 gnd.n5023 585
R11075 gnd.n5023 gnd.n2095 585
R11076 gnd.n5025 gnd.n2103 585
R11077 gnd.n5035 gnd.n2103 585
R11078 gnd.n5027 gnd.n5026 585
R11079 gnd.n5028 gnd.n5027 585
R11080 gnd.n5020 gnd.n2109 585
R11081 gnd.n5029 gnd.n2109 585
R11082 gnd.n5019 gnd.n5018 585
R11083 gnd.n5018 gnd.n1302 585
R11084 gnd.n5017 gnd.n2110 585
R11085 gnd.n5017 gnd.n5016 585
R11086 gnd.n2115 gnd.n2114 585
R11087 gnd.n5011 gnd.n2115 585
R11088 gnd.n2113 gnd.n2111 585
R11089 gnd.n2111 gnd.n1289 585
R11090 gnd.n2112 gnd.n1287 585
R11091 gnd.n6266 gnd.n1287 585
R11092 gnd.n1274 gnd.n1273 585
R11093 gnd.n1286 gnd.n1274 585
R11094 gnd.n6274 gnd.n6273 585
R11095 gnd.n6273 gnd.n6272 585
R11096 gnd.n6275 gnd.n1201 585
R11097 gnd.n1277 gnd.n1201 585
R11098 gnd.n6277 gnd.n6276 585
R11099 gnd.n6278 gnd.n6277 585
R11100 gnd.n1272 gnd.n1200 585
R11101 gnd.n1200 gnd.n1196 585
R11102 gnd.n1271 gnd.n1270 585
R11103 gnd.n1270 gnd.n1186 585
R11104 gnd.n1269 gnd.n1184 585
R11105 gnd.n6285 gnd.n1184 585
R11106 gnd.n1268 gnd.n1267 585
R11107 gnd.n1267 gnd.n1183 585
R11108 gnd.n6409 gnd.n6408 585
R11109 gnd.n6410 gnd.n6409 585
R11110 gnd.n1056 gnd.n1055 585
R11111 gnd.n4778 gnd.n1056 585
R11112 gnd.n6418 gnd.n6417 585
R11113 gnd.n6417 gnd.n6416 585
R11114 gnd.n6419 gnd.n1050 585
R11115 gnd.n4771 gnd.n1050 585
R11116 gnd.n6421 gnd.n6420 585
R11117 gnd.n6422 gnd.n6421 585
R11118 gnd.n1036 gnd.n1035 585
R11119 gnd.n4762 gnd.n1036 585
R11120 gnd.n6430 gnd.n6429 585
R11121 gnd.n6429 gnd.n6428 585
R11122 gnd.n6431 gnd.n1030 585
R11123 gnd.n4756 gnd.n1030 585
R11124 gnd.n6433 gnd.n6432 585
R11125 gnd.n6434 gnd.n6433 585
R11126 gnd.n1015 gnd.n1014 585
R11127 gnd.n4691 gnd.n1015 585
R11128 gnd.n6442 gnd.n6441 585
R11129 gnd.n6441 gnd.n6440 585
R11130 gnd.n6443 gnd.n1009 585
R11131 gnd.n4685 gnd.n1009 585
R11132 gnd.n6445 gnd.n6444 585
R11133 gnd.n6446 gnd.n6445 585
R11134 gnd.n996 gnd.n995 585
R11135 gnd.n4679 gnd.n996 585
R11136 gnd.n6454 gnd.n6453 585
R11137 gnd.n6453 gnd.n6452 585
R11138 gnd.n6455 gnd.n990 585
R11139 gnd.n4708 gnd.n990 585
R11140 gnd.n6457 gnd.n6456 585
R11141 gnd.n6458 gnd.n6457 585
R11142 gnd.n975 gnd.n974 585
R11143 gnd.n4672 gnd.n975 585
R11144 gnd.n6466 gnd.n6465 585
R11145 gnd.n6465 gnd.n6464 585
R11146 gnd.n6467 gnd.n970 585
R11147 gnd.n4664 gnd.n970 585
R11148 gnd.n6469 gnd.n6468 585
R11149 gnd.n6470 gnd.n6469 585
R11150 gnd.n955 gnd.n953 585
R11151 gnd.n4657 gnd.n955 585
R11152 gnd.n6478 gnd.n6477 585
R11153 gnd.n6477 gnd.n6476 585
R11154 gnd.n954 gnd.n952 585
R11155 gnd.n4649 gnd.n954 585
R11156 gnd.n4618 gnd.n4617 585
R11157 gnd.n4619 gnd.n4618 585
R11158 gnd.n4616 gnd.n4615 585
R11159 gnd.n4615 gnd.n2516 585
R11160 gnd.n4614 gnd.n2519 585
R11161 gnd.n4614 gnd.n4613 585
R11162 gnd.n945 gnd.n943 585
R11163 gnd.n4600 gnd.n943 585
R11164 gnd.n6482 gnd.n6481 585
R11165 gnd.n6483 gnd.n6482 585
R11166 gnd.n944 gnd.n942 585
R11167 gnd.n942 gnd.n938 585
R11168 gnd.n4584 gnd.n4583 585
R11169 gnd.n4585 gnd.n4584 585
R11170 gnd.n4582 gnd.n2539 585
R11171 gnd.n4582 gnd.n4581 585
R11172 gnd.n4562 gnd.n2538 585
R11173 gnd.n2540 gnd.n2538 585
R11174 gnd.n4564 gnd.n4563 585
R11175 gnd.n4565 gnd.n4564 585
R11176 gnd.n2552 gnd.n2551 585
R11177 gnd.n2558 gnd.n2551 585
R11178 gnd.n4558 gnd.n4557 585
R11179 gnd.n4557 gnd.n4556 585
R11180 gnd.n2555 gnd.n2554 585
R11181 gnd.n4545 gnd.n2555 585
R11182 gnd.n4522 gnd.n2575 585
R11183 gnd.n2575 gnd.n2566 585
R11184 gnd.n4524 gnd.n4523 585
R11185 gnd.n4525 gnd.n4524 585
R11186 gnd.n2576 gnd.n2574 585
R11187 gnd.n2583 gnd.n2574 585
R11188 gnd.n4517 gnd.n4516 585
R11189 gnd.n4516 gnd.n4515 585
R11190 gnd.n2579 gnd.n2578 585
R11191 gnd.n2580 gnd.n2579 585
R11192 gnd.n4498 gnd.n4497 585
R11193 gnd.n4499 gnd.n4498 585
R11194 gnd.n2596 gnd.n2595 585
R11195 gnd.n2595 gnd.n2592 585
R11196 gnd.n4493 gnd.n4492 585
R11197 gnd.n4492 gnd.n4491 585
R11198 gnd.n2599 gnd.n2598 585
R11199 gnd.n2600 gnd.n2599 585
R11200 gnd.n4478 gnd.n4477 585
R11201 gnd.n4479 gnd.n4478 585
R11202 gnd.n2613 gnd.n2612 585
R11203 gnd.n2620 gnd.n2612 585
R11204 gnd.n4473 gnd.n4472 585
R11205 gnd.n4472 gnd.n4471 585
R11206 gnd.n2616 gnd.n2615 585
R11207 gnd.n2617 gnd.n2616 585
R11208 gnd.n4458 gnd.n4457 585
R11209 gnd.n4459 gnd.n4458 585
R11210 gnd.n2632 gnd.n2631 585
R11211 gnd.n2631 gnd.n2628 585
R11212 gnd.n4453 gnd.n4452 585
R11213 gnd.n4452 gnd.n4451 585
R11214 gnd.n2635 gnd.n2634 585
R11215 gnd.n2636 gnd.n2635 585
R11216 gnd.n4439 gnd.n4438 585
R11217 gnd.n4437 gnd.n4166 585
R11218 gnd.n4436 gnd.n4165 585
R11219 gnd.n4441 gnd.n4165 585
R11220 gnd.n4435 gnd.n4434 585
R11221 gnd.n4433 gnd.n4432 585
R11222 gnd.n4431 gnd.n4430 585
R11223 gnd.n4429 gnd.n4428 585
R11224 gnd.n4427 gnd.n4426 585
R11225 gnd.n4425 gnd.n4424 585
R11226 gnd.n4423 gnd.n4422 585
R11227 gnd.n4421 gnd.n4420 585
R11228 gnd.n4419 gnd.n4418 585
R11229 gnd.n4417 gnd.n4416 585
R11230 gnd.n4415 gnd.n4414 585
R11231 gnd.n4413 gnd.n4412 585
R11232 gnd.n4411 gnd.n4410 585
R11233 gnd.n4409 gnd.n4408 585
R11234 gnd.n4407 gnd.n4406 585
R11235 gnd.n4404 gnd.n4403 585
R11236 gnd.n4402 gnd.n4401 585
R11237 gnd.n4400 gnd.n4399 585
R11238 gnd.n4398 gnd.n4397 585
R11239 gnd.n4396 gnd.n4395 585
R11240 gnd.n4394 gnd.n4393 585
R11241 gnd.n4392 gnd.n4391 585
R11242 gnd.n4390 gnd.n4389 585
R11243 gnd.n4388 gnd.n4387 585
R11244 gnd.n4386 gnd.n4385 585
R11245 gnd.n4384 gnd.n4383 585
R11246 gnd.n4382 gnd.n4381 585
R11247 gnd.n4380 gnd.n4379 585
R11248 gnd.n4378 gnd.n4377 585
R11249 gnd.n4376 gnd.n4375 585
R11250 gnd.n4374 gnd.n4373 585
R11251 gnd.n4372 gnd.n4371 585
R11252 gnd.n4370 gnd.n4369 585
R11253 gnd.n4368 gnd.n4367 585
R11254 gnd.n4366 gnd.n4365 585
R11255 gnd.n4364 gnd.n4363 585
R11256 gnd.n4362 gnd.n4361 585
R11257 gnd.n4360 gnd.n4359 585
R11258 gnd.n4358 gnd.n4357 585
R11259 gnd.n4356 gnd.n4355 585
R11260 gnd.n4354 gnd.n4353 585
R11261 gnd.n4352 gnd.n4351 585
R11262 gnd.n4350 gnd.n4349 585
R11263 gnd.n4348 gnd.n4347 585
R11264 gnd.n4346 gnd.n4345 585
R11265 gnd.n4344 gnd.n4343 585
R11266 gnd.n4342 gnd.n4341 585
R11267 gnd.n4340 gnd.n4339 585
R11268 gnd.n4338 gnd.n4337 585
R11269 gnd.n4336 gnd.n4335 585
R11270 gnd.n4334 gnd.n4333 585
R11271 gnd.n4332 gnd.n4331 585
R11272 gnd.n4330 gnd.n4329 585
R11273 gnd.n4328 gnd.n4327 585
R11274 gnd.n4326 gnd.n2648 585
R11275 gnd.n4443 gnd.n2647 585
R11276 gnd.n2387 gnd.n2386 585
R11277 gnd.n2384 gnd.n2280 585
R11278 gnd.n2383 gnd.n2382 585
R11279 gnd.n2376 gnd.n2282 585
R11280 gnd.n2378 gnd.n2377 585
R11281 gnd.n2374 gnd.n2284 585
R11282 gnd.n2373 gnd.n2372 585
R11283 gnd.n2366 gnd.n2286 585
R11284 gnd.n2368 gnd.n2367 585
R11285 gnd.n2364 gnd.n2288 585
R11286 gnd.n2363 gnd.n2362 585
R11287 gnd.n2356 gnd.n2290 585
R11288 gnd.n2358 gnd.n2357 585
R11289 gnd.n2354 gnd.n2292 585
R11290 gnd.n2353 gnd.n2352 585
R11291 gnd.n2346 gnd.n2294 585
R11292 gnd.n2348 gnd.n2347 585
R11293 gnd.n2344 gnd.n2296 585
R11294 gnd.n2343 gnd.n2342 585
R11295 gnd.n2336 gnd.n2298 585
R11296 gnd.n2338 gnd.n2337 585
R11297 gnd.n2334 gnd.n2302 585
R11298 gnd.n2333 gnd.n2332 585
R11299 gnd.n2326 gnd.n2304 585
R11300 gnd.n2328 gnd.n2327 585
R11301 gnd.n2324 gnd.n2306 585
R11302 gnd.n2323 gnd.n2322 585
R11303 gnd.n2316 gnd.n2308 585
R11304 gnd.n2318 gnd.n2317 585
R11305 gnd.n2314 gnd.n2311 585
R11306 gnd.n2313 gnd.n1117 585
R11307 gnd.n6360 gnd.n1113 585
R11308 gnd.n6362 gnd.n6361 585
R11309 gnd.n6364 gnd.n1111 585
R11310 gnd.n6366 gnd.n6365 585
R11311 gnd.n6367 gnd.n1106 585
R11312 gnd.n6369 gnd.n6368 585
R11313 gnd.n6371 gnd.n1104 585
R11314 gnd.n6373 gnd.n6372 585
R11315 gnd.n6375 gnd.n1097 585
R11316 gnd.n6377 gnd.n6376 585
R11317 gnd.n6379 gnd.n1095 585
R11318 gnd.n6381 gnd.n6380 585
R11319 gnd.n6382 gnd.n1090 585
R11320 gnd.n6384 gnd.n6383 585
R11321 gnd.n6386 gnd.n1088 585
R11322 gnd.n6388 gnd.n6387 585
R11323 gnd.n6389 gnd.n1083 585
R11324 gnd.n6391 gnd.n6390 585
R11325 gnd.n6393 gnd.n1081 585
R11326 gnd.n6395 gnd.n6394 585
R11327 gnd.n6396 gnd.n1075 585
R11328 gnd.n6398 gnd.n6397 585
R11329 gnd.n6400 gnd.n1074 585
R11330 gnd.n6401 gnd.n1072 585
R11331 gnd.n6404 gnd.n6403 585
R11332 gnd.n6405 gnd.n1069 585
R11333 gnd.n1073 gnd.n1069 585
R11334 gnd.n4775 gnd.n1066 585
R11335 gnd.n6410 gnd.n1066 585
R11336 gnd.n4777 gnd.n4776 585
R11337 gnd.n4778 gnd.n4777 585
R11338 gnd.n4774 gnd.n1058 585
R11339 gnd.n6416 gnd.n1058 585
R11340 gnd.n4773 gnd.n4772 585
R11341 gnd.n4772 gnd.n4771 585
R11342 gnd.n2468 gnd.n1047 585
R11343 gnd.n6422 gnd.n1047 585
R11344 gnd.n4761 gnd.n4760 585
R11345 gnd.n4762 gnd.n4761 585
R11346 gnd.n4759 gnd.n1037 585
R11347 gnd.n6428 gnd.n1037 585
R11348 gnd.n4758 gnd.n4757 585
R11349 gnd.n4757 gnd.n4756 585
R11350 gnd.n2473 gnd.n1027 585
R11351 gnd.n6434 gnd.n1027 585
R11352 gnd.n4690 gnd.n4689 585
R11353 gnd.n4691 gnd.n4690 585
R11354 gnd.n4688 gnd.n1017 585
R11355 gnd.n6440 gnd.n1017 585
R11356 gnd.n4687 gnd.n4686 585
R11357 gnd.n4686 gnd.n4685 585
R11358 gnd.n4682 gnd.n1007 585
R11359 gnd.n6446 gnd.n1007 585
R11360 gnd.n4681 gnd.n4680 585
R11361 gnd.n4680 gnd.n4679 585
R11362 gnd.n4678 gnd.n997 585
R11363 gnd.n6452 gnd.n997 585
R11364 gnd.n4677 gnd.n2487 585
R11365 gnd.n4708 gnd.n2487 585
R11366 gnd.n4675 gnd.n987 585
R11367 gnd.n6458 gnd.n987 585
R11368 gnd.n4674 gnd.n4673 585
R11369 gnd.n4673 gnd.n4672 585
R11370 gnd.n2496 gnd.n977 585
R11371 gnd.n6464 gnd.n977 585
R11372 gnd.n4663 gnd.n4662 585
R11373 gnd.n4664 gnd.n4663 585
R11374 gnd.n4660 gnd.n968 585
R11375 gnd.n6470 gnd.n968 585
R11376 gnd.n4659 gnd.n4658 585
R11377 gnd.n4658 gnd.n4657 585
R11378 gnd.n2501 gnd.n956 585
R11379 gnd.n6476 gnd.n956 585
R11380 gnd.n4606 gnd.n2507 585
R11381 gnd.n4649 gnd.n2507 585
R11382 gnd.n4607 gnd.n2517 585
R11383 gnd.n4619 gnd.n2517 585
R11384 gnd.n4605 gnd.n4604 585
R11385 gnd.n4604 gnd.n2516 585
R11386 gnd.n4603 gnd.n2521 585
R11387 gnd.n4613 gnd.n2521 585
R11388 gnd.n4602 gnd.n4601 585
R11389 gnd.n4601 gnd.n4600 585
R11390 gnd.n2530 gnd.n939 585
R11391 gnd.n6483 gnd.n939 585
R11392 gnd.n4572 gnd.n4571 585
R11393 gnd.n4571 gnd.n938 585
R11394 gnd.n4570 gnd.n2536 585
R11395 gnd.n4585 gnd.n2536 585
R11396 gnd.n4569 gnd.n2541 585
R11397 gnd.n4581 gnd.n2541 585
R11398 gnd.n4568 gnd.n4567 585
R11399 gnd.n4567 gnd.n2540 585
R11400 gnd.n4566 gnd.n2546 585
R11401 gnd.n4566 gnd.n4565 585
R11402 gnd.n4549 gnd.n2548 585
R11403 gnd.n2558 gnd.n2548 585
R11404 gnd.n4548 gnd.n2556 585
R11405 gnd.n4556 gnd.n2556 585
R11406 gnd.n4547 gnd.n4546 585
R11407 gnd.n4546 gnd.n4545 585
R11408 gnd.n2565 gnd.n2563 585
R11409 gnd.n2566 gnd.n2565 585
R11410 gnd.n4506 gnd.n2572 585
R11411 gnd.n4525 gnd.n2572 585
R11412 gnd.n4505 gnd.n4504 585
R11413 gnd.n4504 gnd.n2583 585
R11414 gnd.n4503 gnd.n2581 585
R11415 gnd.n4515 gnd.n2581 585
R11416 gnd.n4502 gnd.n4501 585
R11417 gnd.n4501 gnd.n2580 585
R11418 gnd.n4500 gnd.n2589 585
R11419 gnd.n4500 gnd.n4499 585
R11420 gnd.n4484 gnd.n2591 585
R11421 gnd.n2592 gnd.n2591 585
R11422 gnd.n4483 gnd.n2601 585
R11423 gnd.n4491 gnd.n2601 585
R11424 gnd.n4482 gnd.n4481 585
R11425 gnd.n4481 gnd.n2600 585
R11426 gnd.n4480 gnd.n2607 585
R11427 gnd.n4480 gnd.n4479 585
R11428 gnd.n4464 gnd.n2609 585
R11429 gnd.n2620 gnd.n2609 585
R11430 gnd.n4463 gnd.n2618 585
R11431 gnd.n4471 gnd.n2618 585
R11432 gnd.n4462 gnd.n4461 585
R11433 gnd.n4461 gnd.n2617 585
R11434 gnd.n4460 gnd.n2625 585
R11435 gnd.n4460 gnd.n4459 585
R11436 gnd.n4446 gnd.n2627 585
R11437 gnd.n2628 gnd.n2627 585
R11438 gnd.n4447 gnd.n2637 585
R11439 gnd.n4451 gnd.n2637 585
R11440 gnd.n4445 gnd.n4444 585
R11441 gnd.n4444 gnd.n2636 585
R11442 gnd.n7548 gnd.n7547 585
R11443 gnd.n7549 gnd.n7548 585
R11444 gnd.n201 gnd.n200 585
R11445 gnd.n209 gnd.n201 585
R11446 gnd.n7557 gnd.n7556 585
R11447 gnd.n7556 gnd.n7555 585
R11448 gnd.n7558 gnd.n195 585
R11449 gnd.n195 gnd.n194 585
R11450 gnd.n7560 gnd.n7559 585
R11451 gnd.n7561 gnd.n7560 585
R11452 gnd.n181 gnd.n180 585
R11453 gnd.n191 gnd.n181 585
R11454 gnd.n7569 gnd.n7568 585
R11455 gnd.n7568 gnd.n7567 585
R11456 gnd.n7570 gnd.n175 585
R11457 gnd.n175 gnd.n174 585
R11458 gnd.n7572 gnd.n7571 585
R11459 gnd.n7573 gnd.n7572 585
R11460 gnd.n161 gnd.n160 585
R11461 gnd.n171 gnd.n161 585
R11462 gnd.n7581 gnd.n7580 585
R11463 gnd.n7580 gnd.n7579 585
R11464 gnd.n7582 gnd.n155 585
R11465 gnd.n162 gnd.n155 585
R11466 gnd.n7584 gnd.n7583 585
R11467 gnd.n7585 gnd.n7584 585
R11468 gnd.n143 gnd.n142 585
R11469 gnd.n146 gnd.n143 585
R11470 gnd.n7593 gnd.n7592 585
R11471 gnd.n7592 gnd.n7591 585
R11472 gnd.n7594 gnd.n137 585
R11473 gnd.n137 gnd.n136 585
R11474 gnd.n7596 gnd.n7595 585
R11475 gnd.n7597 gnd.n7596 585
R11476 gnd.n123 gnd.n122 585
R11477 gnd.n133 gnd.n123 585
R11478 gnd.n7605 gnd.n7604 585
R11479 gnd.n7604 gnd.n7603 585
R11480 gnd.n7606 gnd.n118 585
R11481 gnd.n124 gnd.n118 585
R11482 gnd.n7608 gnd.n7607 585
R11483 gnd.n7609 gnd.n7608 585
R11484 gnd.n104 gnd.n102 585
R11485 gnd.n107 gnd.n104 585
R11486 gnd.n7617 gnd.n7616 585
R11487 gnd.n7616 gnd.n7615 585
R11488 gnd.n103 gnd.n95 585
R11489 gnd.n7357 gnd.n103 585
R11490 gnd.n7620 gnd.n93 585
R11491 gnd.n368 gnd.n93 585
R11492 gnd.n7622 gnd.n7621 585
R11493 gnd.n7623 gnd.n7622 585
R11494 gnd.n385 gnd.n92 585
R11495 gnd.n7308 gnd.n92 585
R11496 gnd.n7296 gnd.n386 585
R11497 gnd.n7296 gnd.n7295 585
R11498 gnd.n7298 gnd.n7297 585
R11499 gnd.n7299 gnd.n7298 585
R11500 gnd.n384 gnd.n100 585
R11501 gnd.n1699 gnd.n384 585
R11502 gnd.n5888 gnd.n1695 585
R11503 gnd.n5888 gnd.n5887 585
R11504 gnd.n5890 gnd.n5889 585
R11505 gnd.n5891 gnd.n5890 585
R11506 gnd.n1682 gnd.n1681 585
R11507 gnd.n5858 gnd.n1682 585
R11508 gnd.n5899 gnd.n5898 585
R11509 gnd.n5898 gnd.n5897 585
R11510 gnd.n5900 gnd.n1676 585
R11511 gnd.n5874 gnd.n1676 585
R11512 gnd.n5902 gnd.n5901 585
R11513 gnd.n5903 gnd.n5902 585
R11514 gnd.n1661 gnd.n1660 585
R11515 gnd.n5844 gnd.n1661 585
R11516 gnd.n5911 gnd.n5910 585
R11517 gnd.n5910 gnd.n5909 585
R11518 gnd.n5912 gnd.n1655 585
R11519 gnd.n5836 gnd.n1655 585
R11520 gnd.n5914 gnd.n5913 585
R11521 gnd.n5915 gnd.n5914 585
R11522 gnd.n1642 gnd.n1641 585
R11523 gnd.n5829 gnd.n1642 585
R11524 gnd.n5923 gnd.n5922 585
R11525 gnd.n5922 gnd.n5921 585
R11526 gnd.n5924 gnd.n1636 585
R11527 gnd.n5821 gnd.n1636 585
R11528 gnd.n5926 gnd.n5925 585
R11529 gnd.n5927 gnd.n5926 585
R11530 gnd.n1621 gnd.n1620 585
R11531 gnd.n5758 gnd.n1621 585
R11532 gnd.n5935 gnd.n5934 585
R11533 gnd.n5934 gnd.n5933 585
R11534 gnd.n5936 gnd.n1615 585
R11535 gnd.n5749 gnd.n1615 585
R11536 gnd.n5938 gnd.n5937 585
R11537 gnd.n5939 gnd.n5938 585
R11538 gnd.n1598 gnd.n1597 585
R11539 gnd.n5743 gnd.n1598 585
R11540 gnd.n5947 gnd.n5946 585
R11541 gnd.n5946 gnd.n5945 585
R11542 gnd.n5948 gnd.n1589 585
R11543 gnd.n5736 gnd.n1589 585
R11544 gnd.n5950 gnd.n5949 585
R11545 gnd.n5951 gnd.n5950 585
R11546 gnd.n1590 gnd.n1588 585
R11547 gnd.n5775 gnd.n1588 585
R11548 gnd.n1591 gnd.n1510 585
R11549 gnd.n5959 gnd.n1510 585
R11550 gnd.n6078 gnd.n6077 585
R11551 gnd.n6076 gnd.n1509 585
R11552 gnd.n6075 gnd.n1508 585
R11553 gnd.n6080 gnd.n1508 585
R11554 gnd.n6074 gnd.n6073 585
R11555 gnd.n6072 gnd.n6071 585
R11556 gnd.n6070 gnd.n6069 585
R11557 gnd.n6068 gnd.n6067 585
R11558 gnd.n6066 gnd.n6065 585
R11559 gnd.n6064 gnd.n6063 585
R11560 gnd.n6062 gnd.n6061 585
R11561 gnd.n6060 gnd.n6059 585
R11562 gnd.n6058 gnd.n6057 585
R11563 gnd.n6056 gnd.n6055 585
R11564 gnd.n6054 gnd.n6053 585
R11565 gnd.n6052 gnd.n6051 585
R11566 gnd.n6050 gnd.n6049 585
R11567 gnd.n6048 gnd.n6047 585
R11568 gnd.n6046 gnd.n6045 585
R11569 gnd.n6043 gnd.n6042 585
R11570 gnd.n6041 gnd.n6040 585
R11571 gnd.n6039 gnd.n6038 585
R11572 gnd.n6037 gnd.n6036 585
R11573 gnd.n6035 gnd.n6034 585
R11574 gnd.n6033 gnd.n6032 585
R11575 gnd.n6031 gnd.n6030 585
R11576 gnd.n6029 gnd.n6028 585
R11577 gnd.n6026 gnd.n6025 585
R11578 gnd.n6024 gnd.n6023 585
R11579 gnd.n6022 gnd.n6021 585
R11580 gnd.n6020 gnd.n6019 585
R11581 gnd.n6018 gnd.n6017 585
R11582 gnd.n6016 gnd.n6015 585
R11583 gnd.n6014 gnd.n6013 585
R11584 gnd.n6012 gnd.n6011 585
R11585 gnd.n6010 gnd.n6009 585
R11586 gnd.n6008 gnd.n6007 585
R11587 gnd.n6006 gnd.n6005 585
R11588 gnd.n6004 gnd.n6003 585
R11589 gnd.n6002 gnd.n6001 585
R11590 gnd.n6000 gnd.n5999 585
R11591 gnd.n5998 gnd.n5997 585
R11592 gnd.n5996 gnd.n5995 585
R11593 gnd.n5994 gnd.n5993 585
R11594 gnd.n5992 gnd.n5991 585
R11595 gnd.n5990 gnd.n5989 585
R11596 gnd.n5988 gnd.n5987 585
R11597 gnd.n5986 gnd.n5985 585
R11598 gnd.n5984 gnd.n5983 585
R11599 gnd.n5982 gnd.n5981 585
R11600 gnd.n5980 gnd.n5979 585
R11601 gnd.n5978 gnd.n5977 585
R11602 gnd.n5976 gnd.n5975 585
R11603 gnd.n5974 gnd.n5973 585
R11604 gnd.n5972 gnd.n5971 585
R11605 gnd.n5970 gnd.n5969 585
R11606 gnd.n5968 gnd.n5967 585
R11607 gnd.n5962 gnd.n5961 585
R11608 gnd.n7439 gnd.n7438 585
R11609 gnd.n7441 gnd.n315 585
R11610 gnd.n7443 gnd.n7442 585
R11611 gnd.n7444 gnd.n308 585
R11612 gnd.n7446 gnd.n7445 585
R11613 gnd.n7448 gnd.n306 585
R11614 gnd.n7450 gnd.n7449 585
R11615 gnd.n7451 gnd.n301 585
R11616 gnd.n7453 gnd.n7452 585
R11617 gnd.n7455 gnd.n299 585
R11618 gnd.n7457 gnd.n7456 585
R11619 gnd.n7458 gnd.n294 585
R11620 gnd.n7460 gnd.n7459 585
R11621 gnd.n7462 gnd.n292 585
R11622 gnd.n7464 gnd.n7463 585
R11623 gnd.n7465 gnd.n287 585
R11624 gnd.n7467 gnd.n7466 585
R11625 gnd.n7469 gnd.n286 585
R11626 gnd.n7470 gnd.n283 585
R11627 gnd.n7473 gnd.n7472 585
R11628 gnd.n285 gnd.n279 585
R11629 gnd.n7477 gnd.n276 585
R11630 gnd.n7479 gnd.n7478 585
R11631 gnd.n7481 gnd.n274 585
R11632 gnd.n7483 gnd.n7482 585
R11633 gnd.n7484 gnd.n269 585
R11634 gnd.n7486 gnd.n7485 585
R11635 gnd.n7488 gnd.n267 585
R11636 gnd.n7490 gnd.n7489 585
R11637 gnd.n7491 gnd.n262 585
R11638 gnd.n7493 gnd.n7492 585
R11639 gnd.n7495 gnd.n260 585
R11640 gnd.n7497 gnd.n7496 585
R11641 gnd.n7498 gnd.n255 585
R11642 gnd.n7500 gnd.n7499 585
R11643 gnd.n7502 gnd.n253 585
R11644 gnd.n7504 gnd.n7503 585
R11645 gnd.n7505 gnd.n248 585
R11646 gnd.n7507 gnd.n7506 585
R11647 gnd.n7509 gnd.n246 585
R11648 gnd.n7511 gnd.n7510 585
R11649 gnd.n7515 gnd.n241 585
R11650 gnd.n7517 gnd.n7516 585
R11651 gnd.n7519 gnd.n239 585
R11652 gnd.n7521 gnd.n7520 585
R11653 gnd.n7522 gnd.n234 585
R11654 gnd.n7524 gnd.n7523 585
R11655 gnd.n7526 gnd.n232 585
R11656 gnd.n7528 gnd.n7527 585
R11657 gnd.n7529 gnd.n227 585
R11658 gnd.n7531 gnd.n7530 585
R11659 gnd.n7533 gnd.n225 585
R11660 gnd.n7535 gnd.n7534 585
R11661 gnd.n7536 gnd.n220 585
R11662 gnd.n7538 gnd.n7537 585
R11663 gnd.n7540 gnd.n218 585
R11664 gnd.n7542 gnd.n7541 585
R11665 gnd.n7543 gnd.n216 585
R11666 gnd.n7544 gnd.n213 585
R11667 gnd.n213 gnd.n212 585
R11668 gnd.n7321 gnd.n210 585
R11669 gnd.n7549 gnd.n210 585
R11670 gnd.n7323 gnd.n7322 585
R11671 gnd.n7322 gnd.n209 585
R11672 gnd.n7324 gnd.n202 585
R11673 gnd.n7555 gnd.n202 585
R11674 gnd.n7326 gnd.n7325 585
R11675 gnd.n7325 gnd.n194 585
R11676 gnd.n7327 gnd.n192 585
R11677 gnd.n7561 gnd.n192 585
R11678 gnd.n7329 gnd.n7328 585
R11679 gnd.n7328 gnd.n191 585
R11680 gnd.n7330 gnd.n182 585
R11681 gnd.n7567 gnd.n182 585
R11682 gnd.n7332 gnd.n7331 585
R11683 gnd.n7331 gnd.n174 585
R11684 gnd.n7333 gnd.n172 585
R11685 gnd.n7573 gnd.n172 585
R11686 gnd.n7335 gnd.n7334 585
R11687 gnd.n7334 gnd.n171 585
R11688 gnd.n7336 gnd.n163 585
R11689 gnd.n7579 gnd.n163 585
R11690 gnd.n7338 gnd.n7337 585
R11691 gnd.n7337 gnd.n162 585
R11692 gnd.n7339 gnd.n153 585
R11693 gnd.n7585 gnd.n153 585
R11694 gnd.n7341 gnd.n7340 585
R11695 gnd.n7340 gnd.n146 585
R11696 gnd.n7342 gnd.n144 585
R11697 gnd.n7591 gnd.n144 585
R11698 gnd.n7344 gnd.n7343 585
R11699 gnd.n7343 gnd.n136 585
R11700 gnd.n7345 gnd.n134 585
R11701 gnd.n7597 gnd.n134 585
R11702 gnd.n7347 gnd.n7346 585
R11703 gnd.n7346 gnd.n133 585
R11704 gnd.n7348 gnd.n125 585
R11705 gnd.n7603 gnd.n125 585
R11706 gnd.n7350 gnd.n7349 585
R11707 gnd.n7349 gnd.n124 585
R11708 gnd.n7351 gnd.n116 585
R11709 gnd.n7609 gnd.n116 585
R11710 gnd.n7353 gnd.n7352 585
R11711 gnd.n7352 gnd.n107 585
R11712 gnd.n7354 gnd.n105 585
R11713 gnd.n7615 gnd.n105 585
R11714 gnd.n7356 gnd.n7355 585
R11715 gnd.n7357 gnd.n7356 585
R11716 gnd.n370 gnd.n369 585
R11717 gnd.n369 gnd.n368 585
R11718 gnd.n7305 gnd.n89 585
R11719 gnd.n7623 gnd.n89 585
R11720 gnd.n7307 gnd.n7306 585
R11721 gnd.n7308 gnd.n7307 585
R11722 gnd.n7304 gnd.n376 585
R11723 gnd.n7295 gnd.n376 585
R11724 gnd.n382 gnd.n377 585
R11725 gnd.n7299 gnd.n382 585
R11726 gnd.n5853 gnd.n5852 585
R11727 gnd.n5852 gnd.n1699 585
R11728 gnd.n5854 gnd.n1697 585
R11729 gnd.n5887 gnd.n1697 585
R11730 gnd.n5855 gnd.n1693 585
R11731 gnd.n5891 gnd.n1693 585
R11732 gnd.n5857 gnd.n5856 585
R11733 gnd.n5858 gnd.n5857 585
R11734 gnd.n5850 gnd.n1683 585
R11735 gnd.n5897 gnd.n1683 585
R11736 gnd.n5849 gnd.n1706 585
R11737 gnd.n5874 gnd.n1706 585
R11738 gnd.n5847 gnd.n1673 585
R11739 gnd.n5903 gnd.n1673 585
R11740 gnd.n5846 gnd.n5845 585
R11741 gnd.n5845 gnd.n5844 585
R11742 gnd.n1711 gnd.n1663 585
R11743 gnd.n5909 gnd.n1663 585
R11744 gnd.n5835 gnd.n5834 585
R11745 gnd.n5836 gnd.n5835 585
R11746 gnd.n5832 gnd.n1653 585
R11747 gnd.n5915 gnd.n1653 585
R11748 gnd.n5831 gnd.n5830 585
R11749 gnd.n5830 gnd.n5829 585
R11750 gnd.n1716 gnd.n1643 585
R11751 gnd.n5921 gnd.n1643 585
R11752 gnd.n5754 gnd.n1720 585
R11753 gnd.n5821 gnd.n1720 585
R11754 gnd.n5755 gnd.n1633 585
R11755 gnd.n5927 gnd.n1633 585
R11756 gnd.n5757 gnd.n5756 585
R11757 gnd.n5758 gnd.n5757 585
R11758 gnd.n5752 gnd.n1623 585
R11759 gnd.n5933 gnd.n1623 585
R11760 gnd.n5751 gnd.n5750 585
R11761 gnd.n5750 gnd.n5749 585
R11762 gnd.n5746 gnd.n1613 585
R11763 gnd.n5939 gnd.n1613 585
R11764 gnd.n5745 gnd.n5744 585
R11765 gnd.n5744 gnd.n5743 585
R11766 gnd.n5742 gnd.n1600 585
R11767 gnd.n5945 gnd.n1600 585
R11768 gnd.n1584 gnd.n1583 585
R11769 gnd.n5736 gnd.n1584 585
R11770 gnd.n5953 gnd.n5952 585
R11771 gnd.n5952 gnd.n5951 585
R11772 gnd.n5954 gnd.n1573 585
R11773 gnd.n5775 gnd.n1573 585
R11774 gnd.n5960 gnd.n1574 585
R11775 gnd.n5960 gnd.n5959 585
R11776 gnd.n6486 gnd.n6485 585
R11777 gnd.n6485 gnd.n6484 585
R11778 gnd.n7287 gnd.n7286 585
R11779 gnd.n7286 gnd.n90 585
R11780 gnd.n7290 gnd.n388 585
R11781 gnd.n388 gnd.n375 585
R11782 gnd.n7292 gnd.n7291 585
R11783 gnd.n7293 gnd.n7292 585
R11784 gnd.n389 gnd.n387 585
R11785 gnd.n387 gnd.n381 585
R11786 gnd.n5885 gnd.n5884 585
R11787 gnd.n5886 gnd.n5885 585
R11788 gnd.n1701 gnd.n1700 585
R11789 gnd.n1700 gnd.n1696 585
R11790 gnd.n5879 gnd.n5878 585
R11791 gnd.n5878 gnd.n1692 585
R11792 gnd.n5877 gnd.n1703 585
R11793 gnd.n5877 gnd.n1685 585
R11794 gnd.n5876 gnd.n1705 585
R11795 gnd.n5876 gnd.n5875 585
R11796 gnd.n5808 gnd.n1704 585
R11797 gnd.n1704 gnd.n1675 585
R11798 gnd.n5810 gnd.n5809 585
R11799 gnd.n5809 gnd.n1672 585
R11800 gnd.n5811 gnd.n5801 585
R11801 gnd.n5801 gnd.n1665 585
R11802 gnd.n5813 gnd.n5812 585
R11803 gnd.n5813 gnd.n1662 585
R11804 gnd.n5814 gnd.n5800 585
R11805 gnd.n5814 gnd.n1715 585
R11806 gnd.n5816 gnd.n5815 585
R11807 gnd.n5815 gnd.n1652 585
R11808 gnd.n5817 gnd.n1722 585
R11809 gnd.n1722 gnd.n1645 585
R11810 gnd.n5819 gnd.n5818 585
R11811 gnd.n5820 gnd.n5819 585
R11812 gnd.n1723 gnd.n1721 585
R11813 gnd.n1721 gnd.n1635 585
R11814 gnd.n5794 gnd.n5793 585
R11815 gnd.n5793 gnd.n1632 585
R11816 gnd.n5792 gnd.n1725 585
R11817 gnd.n5792 gnd.n1625 585
R11818 gnd.n5791 gnd.n5790 585
R11819 gnd.n5791 gnd.n1622 585
R11820 gnd.n1727 gnd.n1726 585
R11821 gnd.n5748 gnd.n1726 585
R11822 gnd.n5786 gnd.n5785 585
R11823 gnd.n5785 gnd.n1612 585
R11824 gnd.n5784 gnd.n1729 585
R11825 gnd.n5784 gnd.n1602 585
R11826 gnd.n5783 gnd.n5782 585
R11827 gnd.n5783 gnd.n1599 585
R11828 gnd.n1731 gnd.n1730 585
R11829 gnd.n1730 gnd.n1586 585
R11830 gnd.n5778 gnd.n5777 585
R11831 gnd.n5777 gnd.n5776 585
R11832 gnd.n1734 gnd.n1733 585
R11833 gnd.n1734 gnd.n1577 585
R11834 gnd.n5719 gnd.n5718 585
R11835 gnd.n5719 gnd.n1575 585
R11836 gnd.n5720 gnd.n5715 585
R11837 gnd.n5720 gnd.n1507 585
R11838 gnd.n5722 gnd.n5721 585
R11839 gnd.n5721 gnd.n1465 585
R11840 gnd.n5723 gnd.n1766 585
R11841 gnd.n1766 gnd.n1764 585
R11842 gnd.n5725 gnd.n5724 585
R11843 gnd.n5726 gnd.n5725 585
R11844 gnd.n1767 gnd.n1765 585
R11845 gnd.n1765 gnd.n1398 585
R11846 gnd.n5709 gnd.n1397 585
R11847 gnd.n6148 gnd.n1397 585
R11848 gnd.n5708 gnd.n5707 585
R11849 gnd.n5707 gnd.n1396 585
R11850 gnd.n5706 gnd.n1769 585
R11851 gnd.n5706 gnd.n5705 585
R11852 gnd.n5693 gnd.n1770 585
R11853 gnd.n1771 gnd.n1770 585
R11854 gnd.n5695 gnd.n5694 585
R11855 gnd.n5696 gnd.n5695 585
R11856 gnd.n1779 gnd.n1778 585
R11857 gnd.n1778 gnd.n1777 585
R11858 gnd.n5687 gnd.n5686 585
R11859 gnd.n5686 gnd.n5685 585
R11860 gnd.n1782 gnd.n1781 585
R11861 gnd.n1789 gnd.n1782 585
R11862 gnd.n5675 gnd.n5674 585
R11863 gnd.n5676 gnd.n5675 585
R11864 gnd.n1791 gnd.n1790 585
R11865 gnd.n1790 gnd.n1788 585
R11866 gnd.n5670 gnd.n5669 585
R11867 gnd.n5669 gnd.n5668 585
R11868 gnd.n1794 gnd.n1793 585
R11869 gnd.n1795 gnd.n1794 585
R11870 gnd.n5658 gnd.n5657 585
R11871 gnd.n5659 gnd.n5658 585
R11872 gnd.n1803 gnd.n1802 585
R11873 gnd.n1802 gnd.n1801 585
R11874 gnd.n5653 gnd.n5652 585
R11875 gnd.n5652 gnd.n5651 585
R11876 gnd.n1806 gnd.n1805 585
R11877 gnd.n1807 gnd.n1806 585
R11878 gnd.n5641 gnd.n5640 585
R11879 gnd.n5642 gnd.n5641 585
R11880 gnd.n1815 gnd.n1814 585
R11881 gnd.n1814 gnd.n1813 585
R11882 gnd.n5636 gnd.n5635 585
R11883 gnd.n5635 gnd.n5634 585
R11884 gnd.n1818 gnd.n1817 585
R11885 gnd.n1819 gnd.n1818 585
R11886 gnd.n5624 gnd.n5623 585
R11887 gnd.n5625 gnd.n5624 585
R11888 gnd.n1826 gnd.n1825 585
R11889 gnd.n1849 gnd.n1825 585
R11890 gnd.n5619 gnd.n5618 585
R11891 gnd.n5618 gnd.n5617 585
R11892 gnd.n1829 gnd.n1828 585
R11893 gnd.n1872 gnd.n1829 585
R11894 gnd.n5449 gnd.n5448 585
R11895 gnd.n5450 gnd.n5449 585
R11896 gnd.n1882 gnd.n1881 585
R11897 gnd.n1881 gnd.n1877 585
R11898 gnd.n5444 gnd.n5443 585
R11899 gnd.n5443 gnd.n5442 585
R11900 gnd.n1885 gnd.n1884 585
R11901 gnd.n5433 gnd.n1885 585
R11902 gnd.n5411 gnd.n1902 585
R11903 gnd.n5370 gnd.n1902 585
R11904 gnd.n5413 gnd.n5412 585
R11905 gnd.n5414 gnd.n5413 585
R11906 gnd.n1903 gnd.n1901 585
R11907 gnd.n1911 gnd.n1901 585
R11908 gnd.n5406 gnd.n5405 585
R11909 gnd.n5405 gnd.n5404 585
R11910 gnd.n1906 gnd.n1905 585
R11911 gnd.n5279 gnd.n1906 585
R11912 gnd.n5355 gnd.n1930 585
R11913 gnd.n1930 gnd.n1921 585
R11914 gnd.n5357 gnd.n5356 585
R11915 gnd.n5358 gnd.n5357 585
R11916 gnd.n1931 gnd.n1929 585
R11917 gnd.n1929 gnd.n1925 585
R11918 gnd.n5350 gnd.n5349 585
R11919 gnd.n5349 gnd.n5348 585
R11920 gnd.n1934 gnd.n1933 585
R11921 gnd.n5340 gnd.n1934 585
R11922 gnd.n5317 gnd.n1953 585
R11923 gnd.n5270 gnd.n1953 585
R11924 gnd.n5319 gnd.n5318 585
R11925 gnd.n5320 gnd.n5319 585
R11926 gnd.n1954 gnd.n1952 585
R11927 gnd.n1952 gnd.n1949 585
R11928 gnd.n5312 gnd.n5311 585
R11929 gnd.n5311 gnd.n5310 585
R11930 gnd.n1957 gnd.n1956 585
R11931 gnd.n5301 gnd.n1957 585
R11932 gnd.n5259 gnd.n1972 585
R11933 gnd.n5242 gnd.n1972 585
R11934 gnd.n5261 gnd.n5260 585
R11935 gnd.n5262 gnd.n5261 585
R11936 gnd.n1973 gnd.n1971 585
R11937 gnd.n1980 gnd.n1971 585
R11938 gnd.n5254 gnd.n5253 585
R11939 gnd.n5253 gnd.n5252 585
R11940 gnd.n1976 gnd.n1975 585
R11941 gnd.n1993 gnd.n1976 585
R11942 gnd.n5222 gnd.n5221 585
R11943 gnd.n5223 gnd.n5222 585
R11944 gnd.n2001 gnd.n2000 585
R11945 gnd.n2008 gnd.n2000 585
R11946 gnd.n5217 gnd.n5216 585
R11947 gnd.n5216 gnd.n5215 585
R11948 gnd.n2004 gnd.n2003 585
R11949 gnd.n2012 gnd.n2004 585
R11950 gnd.n5184 gnd.n2028 585
R11951 gnd.n2028 gnd.n2018 585
R11952 gnd.n5186 gnd.n5185 585
R11953 gnd.n5187 gnd.n5186 585
R11954 gnd.n2029 gnd.n2027 585
R11955 gnd.n2027 gnd.n2023 585
R11956 gnd.n5179 gnd.n5178 585
R11957 gnd.n5178 gnd.n5177 585
R11958 gnd.n2032 gnd.n2031 585
R11959 gnd.n5169 gnd.n2032 585
R11960 gnd.n5134 gnd.n2050 585
R11961 gnd.n5061 gnd.n2050 585
R11962 gnd.n5136 gnd.n5135 585
R11963 gnd.n5137 gnd.n5136 585
R11964 gnd.n2051 gnd.n2049 585
R11965 gnd.n2058 gnd.n2049 585
R11966 gnd.n5129 gnd.n5128 585
R11967 gnd.n5128 gnd.n5127 585
R11968 gnd.n2054 gnd.n2053 585
R11969 gnd.n5114 gnd.n2054 585
R11970 gnd.n5102 gnd.n2073 585
R11971 gnd.n5086 gnd.n2073 585
R11972 gnd.n5104 gnd.n5103 585
R11973 gnd.n5105 gnd.n5104 585
R11974 gnd.n2074 gnd.n2072 585
R11975 gnd.n2081 gnd.n2072 585
R11976 gnd.n5097 gnd.n5096 585
R11977 gnd.n5096 gnd.n5095 585
R11978 gnd.n2077 gnd.n2076 585
R11979 gnd.n2091 gnd.n2077 585
R11980 gnd.n5043 gnd.n5042 585
R11981 gnd.n5044 gnd.n5043 585
R11982 gnd.n2100 gnd.n2099 585
R11983 gnd.n2104 gnd.n2099 585
R11984 gnd.n5038 gnd.n5037 585
R11985 gnd.n5037 gnd.n5036 585
R11986 gnd.n1300 gnd.n1299 585
R11987 gnd.n2108 gnd.n1300 585
R11988 gnd.n6261 gnd.n6260 585
R11989 gnd.n6260 gnd.n6259 585
R11990 gnd.n6262 gnd.n1292 585
R11991 gnd.n5010 gnd.n1292 585
R11992 gnd.n6264 gnd.n6263 585
R11993 gnd.n6265 gnd.n6264 585
R11994 gnd.n1293 gnd.n1291 585
R11995 gnd.n1291 gnd.n1276 585
R11996 gnd.n1195 gnd.n1194 585
R11997 gnd.n1275 gnd.n1195 585
R11998 gnd.n6280 gnd.n6279 585
R11999 gnd.n6279 gnd.n6278 585
R12000 gnd.n6281 gnd.n1189 585
R12001 gnd.n4941 gnd.n1189 585
R12002 gnd.n6283 gnd.n6282 585
R12003 gnd.n6284 gnd.n6283 585
R12004 gnd.n1190 gnd.n1188 585
R12005 gnd.n1188 gnd.n1157 585
R12006 gnd.n4972 gnd.n2127 585
R12007 gnd.n2127 gnd.n1125 585
R12008 gnd.n4974 gnd.n4973 585
R12009 gnd.n4975 gnd.n4974 585
R12010 gnd.n2128 gnd.n2126 585
R12011 gnd.n2126 gnd.n2124 585
R12012 gnd.n4966 gnd.n4965 585
R12013 gnd.n4965 gnd.n4964 585
R12014 gnd.n2131 gnd.n2130 585
R12015 gnd.n2132 gnd.n2131 585
R12016 gnd.n4929 gnd.n4928 585
R12017 gnd.n4930 gnd.n4929 585
R12018 gnd.n2143 gnd.n2142 585
R12019 gnd.n2149 gnd.n2142 585
R12020 gnd.n4924 gnd.n4923 585
R12021 gnd.n4923 gnd.n4922 585
R12022 gnd.n2146 gnd.n2145 585
R12023 gnd.n2147 gnd.n2146 585
R12024 gnd.n4913 gnd.n4912 585
R12025 gnd.n4914 gnd.n4913 585
R12026 gnd.n2157 gnd.n2156 585
R12027 gnd.n2163 gnd.n2156 585
R12028 gnd.n4908 gnd.n4907 585
R12029 gnd.n4907 gnd.n4906 585
R12030 gnd.n2160 gnd.n2159 585
R12031 gnd.n2161 gnd.n2160 585
R12032 gnd.n4897 gnd.n4896 585
R12033 gnd.n4898 gnd.n4897 585
R12034 gnd.n2172 gnd.n2171 585
R12035 gnd.n2171 gnd.n2169 585
R12036 gnd.n4892 gnd.n4891 585
R12037 gnd.n4891 gnd.n4890 585
R12038 gnd.n2175 gnd.n2174 585
R12039 gnd.n2176 gnd.n2175 585
R12040 gnd.n4881 gnd.n4880 585
R12041 gnd.n4882 gnd.n4881 585
R12042 gnd.n2186 gnd.n2185 585
R12043 gnd.n2185 gnd.n2183 585
R12044 gnd.n4876 gnd.n4875 585
R12045 gnd.n4875 gnd.n4874 585
R12046 gnd.n2189 gnd.n2188 585
R12047 gnd.n2197 gnd.n2189 585
R12048 gnd.n4865 gnd.n4864 585
R12049 gnd.n4866 gnd.n4865 585
R12050 gnd.n2199 gnd.n2198 585
R12051 gnd.n2198 gnd.n2195 585
R12052 gnd.n4860 gnd.n4859 585
R12053 gnd.n4859 gnd.n4858 585
R12054 gnd.n2202 gnd.n2201 585
R12055 gnd.n2203 gnd.n2202 585
R12056 gnd.n4739 gnd.n4735 585
R12057 gnd.n4735 gnd.n4734 585
R12058 gnd.n4742 gnd.n4740 585
R12059 gnd.n4742 gnd.n4741 585
R12060 gnd.n4743 gnd.n4733 585
R12061 gnd.n4743 gnd.n1068 585
R12062 gnd.n4745 gnd.n4744 585
R12063 gnd.n4744 gnd.n1065 585
R12064 gnd.n4746 gnd.n4728 585
R12065 gnd.n4728 gnd.n2467 585
R12066 gnd.n4748 gnd.n4747 585
R12067 gnd.n4748 gnd.n1057 585
R12068 gnd.n4749 gnd.n4727 585
R12069 gnd.n4749 gnd.n1049 585
R12070 gnd.n4751 gnd.n4750 585
R12071 gnd.n4750 gnd.n1046 585
R12072 gnd.n4752 gnd.n2477 585
R12073 gnd.n2477 gnd.n1039 585
R12074 gnd.n4754 gnd.n4753 585
R12075 gnd.n4755 gnd.n4754 585
R12076 gnd.n2478 gnd.n2476 585
R12077 gnd.n2476 gnd.n1029 585
R12078 gnd.n4721 gnd.n4720 585
R12079 gnd.n4720 gnd.n1026 585
R12080 gnd.n4719 gnd.n2480 585
R12081 gnd.n4719 gnd.n1019 585
R12082 gnd.n4718 gnd.n4717 585
R12083 gnd.n4718 gnd.n1016 585
R12084 gnd.n2482 gnd.n2481 585
R12085 gnd.n4684 gnd.n2481 585
R12086 gnd.n4713 gnd.n4712 585
R12087 gnd.n4712 gnd.n1006 585
R12088 gnd.n4711 gnd.n2484 585
R12089 gnd.n4711 gnd.n999 585
R12090 gnd.n4710 gnd.n2486 585
R12091 gnd.n4710 gnd.n4709 585
R12092 gnd.n4636 gnd.n2485 585
R12093 gnd.n2485 gnd.n989 585
R12094 gnd.n4638 gnd.n4637 585
R12095 gnd.n4637 gnd.n986 585
R12096 gnd.n4639 gnd.n4629 585
R12097 gnd.n4629 gnd.n979 585
R12098 gnd.n4641 gnd.n4640 585
R12099 gnd.n4641 gnd.n976 585
R12100 gnd.n4642 gnd.n4628 585
R12101 gnd.n4642 gnd.n2500 585
R12102 gnd.n4644 gnd.n4643 585
R12103 gnd.n4643 gnd.n967 585
R12104 gnd.n4645 gnd.n2509 585
R12105 gnd.n2509 gnd.n958 585
R12106 gnd.n4647 gnd.n4646 585
R12107 gnd.n4648 gnd.n4647 585
R12108 gnd.n2510 gnd.n2508 585
R12109 gnd.n2508 gnd.n2506 585
R12110 gnd.n4622 gnd.n4621 585
R12111 gnd.n4621 gnd.n4620 585
R12112 gnd.n2515 gnd.n2514 585
R12113 gnd.n2523 gnd.n2515 585
R12114 gnd.n2511 gnd.n937 585
R12115 gnd.n2520 gnd.n937 585
R12116 gnd.n6147 gnd.n6146 585
R12117 gnd.n6148 gnd.n6147 585
R12118 gnd.n1401 gnd.n1399 585
R12119 gnd.n1399 gnd.n1396 585
R12120 gnd.n5703 gnd.n5702 585
R12121 gnd.n5705 gnd.n5703 585
R12122 gnd.n1773 gnd.n1772 585
R12123 gnd.n1772 gnd.n1771 585
R12124 gnd.n5698 gnd.n5697 585
R12125 gnd.n5697 gnd.n5696 585
R12126 gnd.n1776 gnd.n1775 585
R12127 gnd.n1777 gnd.n1776 585
R12128 gnd.n5683 gnd.n5682 585
R12129 gnd.n5685 gnd.n5683 585
R12130 gnd.n1784 gnd.n1783 585
R12131 gnd.n1789 gnd.n1783 585
R12132 gnd.n5678 gnd.n5677 585
R12133 gnd.n5677 gnd.n5676 585
R12134 gnd.n1787 gnd.n1786 585
R12135 gnd.n1788 gnd.n1787 585
R12136 gnd.n5666 gnd.n5665 585
R12137 gnd.n5668 gnd.n5666 585
R12138 gnd.n1797 gnd.n1796 585
R12139 gnd.n1796 gnd.n1795 585
R12140 gnd.n5661 gnd.n5660 585
R12141 gnd.n5660 gnd.n5659 585
R12142 gnd.n1800 gnd.n1799 585
R12143 gnd.n1801 gnd.n1800 585
R12144 gnd.n5649 gnd.n5648 585
R12145 gnd.n5651 gnd.n5649 585
R12146 gnd.n1809 gnd.n1808 585
R12147 gnd.n1808 gnd.n1807 585
R12148 gnd.n5644 gnd.n5643 585
R12149 gnd.n5643 gnd.n5642 585
R12150 gnd.n1812 gnd.n1811 585
R12151 gnd.n1813 gnd.n1812 585
R12152 gnd.n5632 gnd.n5631 585
R12153 gnd.n5634 gnd.n5632 585
R12154 gnd.n1821 gnd.n1820 585
R12155 gnd.n1820 gnd.n1819 585
R12156 gnd.n5627 gnd.n5626 585
R12157 gnd.n5626 gnd.n5625 585
R12158 gnd.n1824 gnd.n1823 585
R12159 gnd.n1849 gnd.n1824 585
R12160 gnd.n5422 gnd.n1831 585
R12161 gnd.n5617 gnd.n1831 585
R12162 gnd.n5425 gnd.n5421 585
R12163 gnd.n5421 gnd.n1872 585
R12164 gnd.n5426 gnd.n1879 585
R12165 gnd.n5450 gnd.n1879 585
R12166 gnd.n5427 gnd.n5420 585
R12167 gnd.n5420 gnd.n1877 585
R12168 gnd.n1895 gnd.n1887 585
R12169 gnd.n5442 gnd.n1887 585
R12170 gnd.n5432 gnd.n5431 585
R12171 gnd.n5433 gnd.n5432 585
R12172 gnd.n1894 gnd.n1893 585
R12173 gnd.n5370 gnd.n1893 585
R12174 gnd.n5416 gnd.n5415 585
R12175 gnd.n5415 gnd.n5414 585
R12176 gnd.n1898 gnd.n1897 585
R12177 gnd.n1911 gnd.n1898 585
R12178 gnd.n5281 gnd.n1908 585
R12179 gnd.n5404 gnd.n1908 585
R12180 gnd.n5282 gnd.n5280 585
R12181 gnd.n5280 gnd.n5279 585
R12182 gnd.n5277 gnd.n5275 585
R12183 gnd.n5277 gnd.n1921 585
R12184 gnd.n5286 gnd.n1927 585
R12185 gnd.n5358 gnd.n1927 585
R12186 gnd.n5287 gnd.n5274 585
R12187 gnd.n5274 gnd.n1925 585
R12188 gnd.n5288 gnd.n1935 585
R12189 gnd.n5348 gnd.n1935 585
R12190 gnd.n5272 gnd.n1943 585
R12191 gnd.n5340 gnd.n1943 585
R12192 gnd.n5292 gnd.n5271 585
R12193 gnd.n5271 gnd.n5270 585
R12194 gnd.n5293 gnd.n1951 585
R12195 gnd.n5320 gnd.n1951 585
R12196 gnd.n5294 gnd.n5268 585
R12197 gnd.n5268 gnd.n1949 585
R12198 gnd.n1966 gnd.n1959 585
R12199 gnd.n5310 gnd.n1959 585
R12200 gnd.n5299 gnd.n5298 585
R12201 gnd.n5301 gnd.n5299 585
R12202 gnd.n1965 gnd.n1964 585
R12203 gnd.n5242 gnd.n1964 585
R12204 gnd.n5264 gnd.n5263 585
R12205 gnd.n5263 gnd.n5262 585
R12206 gnd.n1969 gnd.n1968 585
R12207 gnd.n1980 gnd.n1969 585
R12208 gnd.n5151 gnd.n1978 585
R12209 gnd.n5252 gnd.n1978 585
R12210 gnd.n5150 gnd.n5149 585
R12211 gnd.n5149 gnd.n1993 585
R12212 gnd.n5155 gnd.n1998 585
R12213 gnd.n5223 gnd.n1998 585
R12214 gnd.n5156 gnd.n5148 585
R12215 gnd.n5148 gnd.n2008 585
R12216 gnd.n5157 gnd.n2006 585
R12217 gnd.n5215 gnd.n2006 585
R12218 gnd.n5146 gnd.n5145 585
R12219 gnd.n5145 gnd.n2012 585
R12220 gnd.n5161 gnd.n5144 585
R12221 gnd.n5144 gnd.n2018 585
R12222 gnd.n5162 gnd.n2025 585
R12223 gnd.n5187 gnd.n2025 585
R12224 gnd.n5163 gnd.n5143 585
R12225 gnd.n5143 gnd.n2023 585
R12226 gnd.n2042 gnd.n2034 585
R12227 gnd.n5177 gnd.n2034 585
R12228 gnd.n5168 gnd.n5167 585
R12229 gnd.n5169 gnd.n5168 585
R12230 gnd.n2041 gnd.n2040 585
R12231 gnd.n5061 gnd.n2040 585
R12232 gnd.n5139 gnd.n5138 585
R12233 gnd.n5138 gnd.n5137 585
R12234 gnd.n2045 gnd.n2044 585
R12235 gnd.n2058 gnd.n2045 585
R12236 gnd.n2067 gnd.n2056 585
R12237 gnd.n5127 gnd.n2056 585
R12238 gnd.n5113 gnd.n5112 585
R12239 gnd.n5114 gnd.n5113 585
R12240 gnd.n2066 gnd.n2065 585
R12241 gnd.n5086 gnd.n2065 585
R12242 gnd.n5107 gnd.n5106 585
R12243 gnd.n5106 gnd.n5105 585
R12244 gnd.n2070 gnd.n2069 585
R12245 gnd.n2081 gnd.n2070 585
R12246 gnd.n4997 gnd.n2079 585
R12247 gnd.n5095 gnd.n2079 585
R12248 gnd.n4998 gnd.n4996 585
R12249 gnd.n4996 gnd.n2091 585
R12250 gnd.n4994 gnd.n2097 585
R12251 gnd.n5044 gnd.n2097 585
R12252 gnd.n5002 gnd.n4993 585
R12253 gnd.n4993 gnd.n2104 585
R12254 gnd.n5003 gnd.n2102 585
R12255 gnd.n5036 gnd.n2102 585
R12256 gnd.n5004 gnd.n4992 585
R12257 gnd.n4992 gnd.n2108 585
R12258 gnd.n2117 gnd.n1301 585
R12259 gnd.n6259 gnd.n1301 585
R12260 gnd.n5009 gnd.n5008 585
R12261 gnd.n5010 gnd.n5009 585
R12262 gnd.n2116 gnd.n1288 585
R12263 gnd.n6265 gnd.n1288 585
R12264 gnd.n4988 gnd.n4987 585
R12265 gnd.n4987 gnd.n1276 585
R12266 gnd.n4986 gnd.n4985 585
R12267 gnd.n4986 gnd.n1275 585
R12268 gnd.n4984 gnd.n1198 585
R12269 gnd.n6278 gnd.n1198 585
R12270 gnd.n4940 gnd.n2119 585
R12271 gnd.n4941 gnd.n4940 585
R12272 gnd.n4980 gnd.n1185 585
R12273 gnd.n6284 gnd.n1185 585
R12274 gnd.n4979 gnd.n4978 585
R12275 gnd.n4978 gnd.n1157 585
R12276 gnd.n4977 gnd.n2121 585
R12277 gnd.n4977 gnd.n1125 585
R12278 gnd.n4976 gnd.n2123 585
R12279 gnd.n4976 gnd.n4975 585
R12280 gnd.n2237 gnd.n2122 585
R12281 gnd.n2124 gnd.n2122 585
R12282 gnd.n2242 gnd.n2133 585
R12283 gnd.n4964 gnd.n2133 585
R12284 gnd.n2243 gnd.n2236 585
R12285 gnd.n2236 gnd.n2132 585
R12286 gnd.n2244 gnd.n2141 585
R12287 gnd.n4930 gnd.n2141 585
R12288 gnd.n2234 gnd.n2233 585
R12289 gnd.n2233 gnd.n2149 585
R12290 gnd.n2248 gnd.n2148 585
R12291 gnd.n4922 gnd.n2148 585
R12292 gnd.n2249 gnd.n2232 585
R12293 gnd.n2232 gnd.n2147 585
R12294 gnd.n2250 gnd.n2155 585
R12295 gnd.n4914 gnd.n2155 585
R12296 gnd.n2230 gnd.n2229 585
R12297 gnd.n2229 gnd.n2163 585
R12298 gnd.n2254 gnd.n2162 585
R12299 gnd.n4906 gnd.n2162 585
R12300 gnd.n2255 gnd.n2228 585
R12301 gnd.n2228 gnd.n2161 585
R12302 gnd.n2256 gnd.n2170 585
R12303 gnd.n4898 gnd.n2170 585
R12304 gnd.n2226 gnd.n2225 585
R12305 gnd.n2225 gnd.n2169 585
R12306 gnd.n2260 gnd.n2177 585
R12307 gnd.n4890 gnd.n2177 585
R12308 gnd.n2261 gnd.n2224 585
R12309 gnd.n2224 gnd.n2176 585
R12310 gnd.n2262 gnd.n2184 585
R12311 gnd.n4882 gnd.n2184 585
R12312 gnd.n2222 gnd.n2221 585
R12313 gnd.n2221 gnd.n2183 585
R12314 gnd.n2266 gnd.n2190 585
R12315 gnd.n4874 gnd.n2190 585
R12316 gnd.n2267 gnd.n2220 585
R12317 gnd.n2220 gnd.n2197 585
R12318 gnd.n2268 gnd.n2196 585
R12319 gnd.n4866 gnd.n2196 585
R12320 gnd.n4855 gnd.n4854 585
R12321 gnd.n4853 gnd.n2218 585
R12322 gnd.n2271 gnd.n2217 585
R12323 gnd.n4857 gnd.n2217 585
R12324 gnd.n4849 gnd.n2273 585
R12325 gnd.n4848 gnd.n2274 585
R12326 gnd.n4847 gnd.n2275 585
R12327 gnd.n2391 gnd.n2276 585
R12328 gnd.n4842 gnd.n2392 585
R12329 gnd.n4841 gnd.n2393 585
R12330 gnd.n4840 gnd.n2394 585
R12331 gnd.n2404 gnd.n2395 585
R12332 gnd.n4833 gnd.n2405 585
R12333 gnd.n4832 gnd.n2406 585
R12334 gnd.n2408 gnd.n2407 585
R12335 gnd.n4825 gnd.n2416 585
R12336 gnd.n4824 gnd.n2417 585
R12337 gnd.n2427 gnd.n2418 585
R12338 gnd.n4817 gnd.n2428 585
R12339 gnd.n4816 gnd.n2429 585
R12340 gnd.n2431 gnd.n2430 585
R12341 gnd.n4809 gnd.n2439 585
R12342 gnd.n4808 gnd.n2440 585
R12343 gnd.n2450 gnd.n2441 585
R12344 gnd.n4801 gnd.n2451 585
R12345 gnd.n4800 gnd.n2452 585
R12346 gnd.n4785 gnd.n4784 585
R12347 gnd.n4787 gnd.n4786 585
R12348 gnd.n4790 gnd.n4788 585
R12349 gnd.n4789 gnd.n2194 585
R12350 gnd.n6150 gnd.n6149 585
R12351 gnd.n6149 gnd.n6148 585
R12352 gnd.n6151 gnd.n1394 585
R12353 gnd.n1396 gnd.n1394 585
R12354 gnd.n5704 gnd.n1392 585
R12355 gnd.n5705 gnd.n5704 585
R12356 gnd.n6155 gnd.n1391 585
R12357 gnd.n1771 gnd.n1391 585
R12358 gnd.n6156 gnd.n1390 585
R12359 gnd.n5696 gnd.n1390 585
R12360 gnd.n6157 gnd.n1389 585
R12361 gnd.n1777 gnd.n1389 585
R12362 gnd.n5684 gnd.n1387 585
R12363 gnd.n5685 gnd.n5684 585
R12364 gnd.n6161 gnd.n1386 585
R12365 gnd.n1789 gnd.n1386 585
R12366 gnd.n6162 gnd.n1385 585
R12367 gnd.n5676 gnd.n1385 585
R12368 gnd.n6163 gnd.n1384 585
R12369 gnd.n1788 gnd.n1384 585
R12370 gnd.n5667 gnd.n1382 585
R12371 gnd.n5668 gnd.n5667 585
R12372 gnd.n6167 gnd.n1381 585
R12373 gnd.n1795 gnd.n1381 585
R12374 gnd.n6168 gnd.n1380 585
R12375 gnd.n5659 gnd.n1380 585
R12376 gnd.n6169 gnd.n1379 585
R12377 gnd.n1801 gnd.n1379 585
R12378 gnd.n5650 gnd.n1377 585
R12379 gnd.n5651 gnd.n5650 585
R12380 gnd.n6173 gnd.n1376 585
R12381 gnd.n1807 gnd.n1376 585
R12382 gnd.n6174 gnd.n1375 585
R12383 gnd.n5642 gnd.n1375 585
R12384 gnd.n6175 gnd.n1374 585
R12385 gnd.n1813 gnd.n1374 585
R12386 gnd.n5633 gnd.n1372 585
R12387 gnd.n5634 gnd.n5633 585
R12388 gnd.n6179 gnd.n1371 585
R12389 gnd.n1819 gnd.n1371 585
R12390 gnd.n6180 gnd.n1370 585
R12391 gnd.n5625 gnd.n1370 585
R12392 gnd.n6181 gnd.n1369 585
R12393 gnd.n1849 gnd.n1369 585
R12394 gnd.n5616 gnd.n1367 585
R12395 gnd.n5617 gnd.n5616 585
R12396 gnd.n6185 gnd.n1366 585
R12397 gnd.n1872 gnd.n1366 585
R12398 gnd.n6186 gnd.n1365 585
R12399 gnd.n5450 gnd.n1365 585
R12400 gnd.n6187 gnd.n1364 585
R12401 gnd.n1877 gnd.n1364 585
R12402 gnd.n5441 gnd.n1362 585
R12403 gnd.n5442 gnd.n5441 585
R12404 gnd.n6191 gnd.n1361 585
R12405 gnd.n5433 gnd.n1361 585
R12406 gnd.n6192 gnd.n1360 585
R12407 gnd.n5370 gnd.n1360 585
R12408 gnd.n6193 gnd.n1359 585
R12409 gnd.n5414 gnd.n1359 585
R12410 gnd.n1910 gnd.n1357 585
R12411 gnd.n1911 gnd.n1910 585
R12412 gnd.n6197 gnd.n1356 585
R12413 gnd.n5404 gnd.n1356 585
R12414 gnd.n6198 gnd.n1355 585
R12415 gnd.n5279 gnd.n1355 585
R12416 gnd.n6199 gnd.n1354 585
R12417 gnd.n1921 gnd.n1354 585
R12418 gnd.n1928 gnd.n1352 585
R12419 gnd.n5358 gnd.n1928 585
R12420 gnd.n6203 gnd.n1351 585
R12421 gnd.n1925 gnd.n1351 585
R12422 gnd.n6204 gnd.n1350 585
R12423 gnd.n5348 gnd.n1350 585
R12424 gnd.n6205 gnd.n1349 585
R12425 gnd.n5340 gnd.n1349 585
R12426 gnd.n5269 gnd.n1347 585
R12427 gnd.n5270 gnd.n5269 585
R12428 gnd.n6209 gnd.n1346 585
R12429 gnd.n5320 gnd.n1346 585
R12430 gnd.n6210 gnd.n1345 585
R12431 gnd.n1949 gnd.n1345 585
R12432 gnd.n6211 gnd.n1344 585
R12433 gnd.n5310 gnd.n1344 585
R12434 gnd.n5300 gnd.n1342 585
R12435 gnd.n5301 gnd.n5300 585
R12436 gnd.n6215 gnd.n1341 585
R12437 gnd.n5242 gnd.n1341 585
R12438 gnd.n6216 gnd.n1340 585
R12439 gnd.n5262 gnd.n1340 585
R12440 gnd.n6217 gnd.n1339 585
R12441 gnd.n1980 gnd.n1339 585
R12442 gnd.n5251 gnd.n1337 585
R12443 gnd.n5252 gnd.n5251 585
R12444 gnd.n6221 gnd.n1336 585
R12445 gnd.n1993 gnd.n1336 585
R12446 gnd.n6222 gnd.n1335 585
R12447 gnd.n5223 gnd.n1335 585
R12448 gnd.n6223 gnd.n1334 585
R12449 gnd.n2008 gnd.n1334 585
R12450 gnd.n5214 gnd.n1332 585
R12451 gnd.n5215 gnd.n5214 585
R12452 gnd.n6227 gnd.n1331 585
R12453 gnd.n2012 gnd.n1331 585
R12454 gnd.n6228 gnd.n1330 585
R12455 gnd.n2018 gnd.n1330 585
R12456 gnd.n6229 gnd.n1329 585
R12457 gnd.n5187 gnd.n1329 585
R12458 gnd.n2022 gnd.n1327 585
R12459 gnd.n2023 gnd.n2022 585
R12460 gnd.n6233 gnd.n1326 585
R12461 gnd.n5177 gnd.n1326 585
R12462 gnd.n6234 gnd.n1325 585
R12463 gnd.n5169 gnd.n1325 585
R12464 gnd.n6235 gnd.n1324 585
R12465 gnd.n5061 gnd.n1324 585
R12466 gnd.n2048 gnd.n1322 585
R12467 gnd.n5137 gnd.n2048 585
R12468 gnd.n6239 gnd.n1321 585
R12469 gnd.n2058 gnd.n1321 585
R12470 gnd.n6240 gnd.n1320 585
R12471 gnd.n5127 gnd.n1320 585
R12472 gnd.n6241 gnd.n1319 585
R12473 gnd.n5114 gnd.n1319 585
R12474 gnd.n5085 gnd.n1317 585
R12475 gnd.n5086 gnd.n5085 585
R12476 gnd.n6245 gnd.n1316 585
R12477 gnd.n5105 gnd.n1316 585
R12478 gnd.n6246 gnd.n1315 585
R12479 gnd.n2081 gnd.n1315 585
R12480 gnd.n6247 gnd.n1314 585
R12481 gnd.n5095 gnd.n1314 585
R12482 gnd.n2090 gnd.n1312 585
R12483 gnd.n2091 gnd.n2090 585
R12484 gnd.n6251 gnd.n1311 585
R12485 gnd.n5044 gnd.n1311 585
R12486 gnd.n6252 gnd.n1310 585
R12487 gnd.n2104 gnd.n1310 585
R12488 gnd.n6253 gnd.n1309 585
R12489 gnd.n5036 gnd.n1309 585
R12490 gnd.n1306 gnd.n1304 585
R12491 gnd.n2108 gnd.n1304 585
R12492 gnd.n6258 gnd.n6257 585
R12493 gnd.n6259 gnd.n6258 585
R12494 gnd.n1305 gnd.n1303 585
R12495 gnd.n5010 gnd.n1303 585
R12496 gnd.n4946 gnd.n1290 585
R12497 gnd.n6265 gnd.n1290 585
R12498 gnd.n4945 gnd.n4944 585
R12499 gnd.n4944 gnd.n1276 585
R12500 gnd.n4950 gnd.n4943 585
R12501 gnd.n4943 gnd.n1275 585
R12502 gnd.n4951 gnd.n1199 585
R12503 gnd.n6278 gnd.n1199 585
R12504 gnd.n4952 gnd.n4942 585
R12505 gnd.n4942 gnd.n4941 585
R12506 gnd.n4938 gnd.n1187 585
R12507 gnd.n6284 gnd.n1187 585
R12508 gnd.n4956 gnd.n4937 585
R12509 gnd.n4937 gnd.n1157 585
R12510 gnd.n4957 gnd.n4936 585
R12511 gnd.n4936 gnd.n1125 585
R12512 gnd.n4958 gnd.n2125 585
R12513 gnd.n4975 gnd.n2125 585
R12514 gnd.n2137 gnd.n2135 585
R12515 gnd.n2135 gnd.n2124 585
R12516 gnd.n4963 gnd.n4962 585
R12517 gnd.n4964 gnd.n4963 585
R12518 gnd.n2136 gnd.n2134 585
R12519 gnd.n2134 gnd.n2132 585
R12520 gnd.n4932 gnd.n4931 585
R12521 gnd.n4931 gnd.n4930 585
R12522 gnd.n2140 gnd.n2139 585
R12523 gnd.n2149 gnd.n2140 585
R12524 gnd.n4921 gnd.n4920 585
R12525 gnd.n4922 gnd.n4921 585
R12526 gnd.n2151 gnd.n2150 585
R12527 gnd.n2150 gnd.n2147 585
R12528 gnd.n4916 gnd.n4915 585
R12529 gnd.n4915 gnd.n4914 585
R12530 gnd.n2154 gnd.n2153 585
R12531 gnd.n2163 gnd.n2154 585
R12532 gnd.n4905 gnd.n4904 585
R12533 gnd.n4906 gnd.n4905 585
R12534 gnd.n2165 gnd.n2164 585
R12535 gnd.n2164 gnd.n2161 585
R12536 gnd.n4900 gnd.n4899 585
R12537 gnd.n4899 gnd.n4898 585
R12538 gnd.n2168 gnd.n2167 585
R12539 gnd.n2169 gnd.n2168 585
R12540 gnd.n4889 gnd.n4888 585
R12541 gnd.n4890 gnd.n4889 585
R12542 gnd.n2179 gnd.n2178 585
R12543 gnd.n2178 gnd.n2176 585
R12544 gnd.n4884 gnd.n4883 585
R12545 gnd.n4883 gnd.n4882 585
R12546 gnd.n2182 gnd.n2181 585
R12547 gnd.n2183 gnd.n2182 585
R12548 gnd.n4873 gnd.n4872 585
R12549 gnd.n4874 gnd.n4873 585
R12550 gnd.n2192 gnd.n2191 585
R12551 gnd.n2197 gnd.n2191 585
R12552 gnd.n4868 gnd.n4867 585
R12553 gnd.n4867 gnd.n4866 585
R12554 gnd.n6089 gnd.n1456 585
R12555 gnd.n5727 gnd.n1456 585
R12556 gnd.n6090 gnd.n1455 585
R12557 gnd.n1759 gnd.n1449 585
R12558 gnd.n6097 gnd.n1448 585
R12559 gnd.n6098 gnd.n1447 585
R12560 gnd.n1756 gnd.n1441 585
R12561 gnd.n6105 gnd.n1440 585
R12562 gnd.n6106 gnd.n1439 585
R12563 gnd.n1754 gnd.n1433 585
R12564 gnd.n6113 gnd.n1432 585
R12565 gnd.n6114 gnd.n1431 585
R12566 gnd.n1751 gnd.n1425 585
R12567 gnd.n6121 gnd.n1424 585
R12568 gnd.n6122 gnd.n1423 585
R12569 gnd.n1749 gnd.n1416 585
R12570 gnd.n6129 gnd.n1415 585
R12571 gnd.n6130 gnd.n1414 585
R12572 gnd.n1746 gnd.n1411 585
R12573 gnd.n6135 gnd.n1410 585
R12574 gnd.n6136 gnd.n1409 585
R12575 gnd.n6137 gnd.n1408 585
R12576 gnd.n1743 gnd.n1406 585
R12577 gnd.n6141 gnd.n1405 585
R12578 gnd.n6142 gnd.n1404 585
R12579 gnd.n6143 gnd.n1400 585
R12580 gnd.n5730 gnd.n1395 585
R12581 gnd.n5731 gnd.n5729 585
R12582 gnd.n1741 gnd.n1740 585
R12583 gnd.n1762 gnd.n1761 585
R12584 gnd.n5540 gnd.n1874 473.281
R12585 gnd.n5549 gnd.n5548 473.281
R12586 gnd.n1267 gnd.n1266 473.281
R12587 gnd.n6353 gnd.n1160 473.281
R12588 gnd.n6652 gnd.n766 466.675
R12589 gnd.n1202 gnd.t109 443.966
R12590 gnd.n1867 gnd.t40 443.966
R12591 gnd.n6290 gnd.t29 443.966
R12592 gnd.n5474 gnd.t96 443.966
R12593 gnd.n2453 gnd.t58 371.625
R12594 gnd.n6083 gnd.t11 371.625
R12595 gnd.n2460 gnd.t54 371.625
R12596 gnd.n1529 gnd.t112 371.625
R12597 gnd.n1552 gnd.t118 371.625
R12598 gnd.n5963 gnd.t68 371.625
R12599 gnd.n313 gnd.t93 371.625
R12600 gnd.n280 gnd.t44 371.625
R12601 gnd.n7512 gnd.t87 371.625
R12602 gnd.n350 gnd.t36 371.625
R12603 gnd.n4185 gnd.t71 371.625
R12604 gnd.n4207 gnd.t74 371.625
R12605 gnd.n4228 gnd.t21 371.625
R12606 gnd.n4246 gnd.t99 371.625
R12607 gnd.n1101 gnd.t80 371.625
R12608 gnd.n2278 gnd.t102 371.625
R12609 gnd.n2300 gnd.t125 371.625
R12610 gnd.n1457 gnd.t25 371.625
R12611 gnd.n3146 gnd.t47 323.425
R12612 gnd.n2688 gnd.t83 323.425
R12613 gnd.n3995 gnd.n3969 289.615
R12614 gnd.n3963 gnd.n3937 289.615
R12615 gnd.n3931 gnd.n3905 289.615
R12616 gnd.n3900 gnd.n3874 289.615
R12617 gnd.n3868 gnd.n3842 289.615
R12618 gnd.n3836 gnd.n3810 289.615
R12619 gnd.n3804 gnd.n3778 289.615
R12620 gnd.n3773 gnd.n3747 289.615
R12621 gnd.n3220 gnd.t121 279.217
R12622 gnd.n2714 gnd.t105 279.217
R12623 gnd.n1167 gnd.t17 260.649
R12624 gnd.n5466 gnd.t64 260.649
R12625 gnd.n6355 gnd.n6354 256.663
R12626 gnd.n6355 gnd.n1126 256.663
R12627 gnd.n6355 gnd.n1127 256.663
R12628 gnd.n6355 gnd.n1128 256.663
R12629 gnd.n6355 gnd.n1129 256.663
R12630 gnd.n6355 gnd.n1130 256.663
R12631 gnd.n6355 gnd.n1131 256.663
R12632 gnd.n6355 gnd.n1132 256.663
R12633 gnd.n6355 gnd.n1133 256.663
R12634 gnd.n6355 gnd.n1134 256.663
R12635 gnd.n6355 gnd.n1135 256.663
R12636 gnd.n6355 gnd.n1136 256.663
R12637 gnd.n6355 gnd.n1137 256.663
R12638 gnd.n6355 gnd.n1138 256.663
R12639 gnd.n6355 gnd.n1139 256.663
R12640 gnd.n6355 gnd.n1140 256.663
R12641 gnd.n6358 gnd.n1123 256.663
R12642 gnd.n6356 gnd.n6355 256.663
R12643 gnd.n6355 gnd.n1141 256.663
R12644 gnd.n6355 gnd.n1142 256.663
R12645 gnd.n6355 gnd.n1143 256.663
R12646 gnd.n6355 gnd.n1144 256.663
R12647 gnd.n6355 gnd.n1145 256.663
R12648 gnd.n6355 gnd.n1146 256.663
R12649 gnd.n6355 gnd.n1147 256.663
R12650 gnd.n6355 gnd.n1148 256.663
R12651 gnd.n6355 gnd.n1149 256.663
R12652 gnd.n6355 gnd.n1150 256.663
R12653 gnd.n6355 gnd.n1151 256.663
R12654 gnd.n6355 gnd.n1152 256.663
R12655 gnd.n6355 gnd.n1153 256.663
R12656 gnd.n6355 gnd.n1154 256.663
R12657 gnd.n6355 gnd.n1155 256.663
R12658 gnd.n6355 gnd.n1156 256.663
R12659 gnd.n5615 gnd.n1850 256.663
R12660 gnd.n5615 gnd.n1851 256.663
R12661 gnd.n5615 gnd.n1852 256.663
R12662 gnd.n5615 gnd.n1853 256.663
R12663 gnd.n5615 gnd.n1854 256.663
R12664 gnd.n5615 gnd.n1855 256.663
R12665 gnd.n5615 gnd.n1856 256.663
R12666 gnd.n5615 gnd.n1857 256.663
R12667 gnd.n5615 gnd.n1858 256.663
R12668 gnd.n5615 gnd.n1859 256.663
R12669 gnd.n5615 gnd.n1860 256.663
R12670 gnd.n5615 gnd.n1861 256.663
R12671 gnd.n5615 gnd.n1862 256.663
R12672 gnd.n5615 gnd.n1863 256.663
R12673 gnd.n5615 gnd.n1864 256.663
R12674 gnd.n5615 gnd.n1865 256.663
R12675 gnd.n1866 gnd.n1539 256.663
R12676 gnd.n5615 gnd.n1848 256.663
R12677 gnd.n5615 gnd.n1847 256.663
R12678 gnd.n5615 gnd.n1846 256.663
R12679 gnd.n5615 gnd.n1845 256.663
R12680 gnd.n5615 gnd.n1844 256.663
R12681 gnd.n5615 gnd.n1843 256.663
R12682 gnd.n5615 gnd.n1842 256.663
R12683 gnd.n5615 gnd.n1841 256.663
R12684 gnd.n5615 gnd.n1840 256.663
R12685 gnd.n5615 gnd.n1839 256.663
R12686 gnd.n5615 gnd.n1838 256.663
R12687 gnd.n5615 gnd.n1837 256.663
R12688 gnd.n5615 gnd.n1836 256.663
R12689 gnd.n5615 gnd.n1835 256.663
R12690 gnd.n5615 gnd.n1834 256.663
R12691 gnd.n5615 gnd.n1833 256.663
R12692 gnd.n5615 gnd.n1832 256.663
R12693 gnd.n4441 gnd.n4155 242.672
R12694 gnd.n4441 gnd.n4156 242.672
R12695 gnd.n4441 gnd.n4157 242.672
R12696 gnd.n4441 gnd.n4158 242.672
R12697 gnd.n4441 gnd.n4159 242.672
R12698 gnd.n4441 gnd.n4160 242.672
R12699 gnd.n4441 gnd.n4161 242.672
R12700 gnd.n4441 gnd.n4162 242.672
R12701 gnd.n4441 gnd.n4163 242.672
R12702 gnd.n4793 gnd.n1073 242.672
R12703 gnd.n2458 gnd.n1073 242.672
R12704 gnd.n2446 gnd.n1073 242.672
R12705 gnd.n2443 gnd.n1073 242.672
R12706 gnd.n2434 gnd.n1073 242.672
R12707 gnd.n2423 gnd.n1073 242.672
R12708 gnd.n2420 gnd.n1073 242.672
R12709 gnd.n2411 gnd.n1073 242.672
R12710 gnd.n2400 gnd.n1073 242.672
R12711 gnd.n3274 gnd.n3273 242.672
R12712 gnd.n3274 gnd.n3184 242.672
R12713 gnd.n3274 gnd.n3185 242.672
R12714 gnd.n3274 gnd.n3186 242.672
R12715 gnd.n3274 gnd.n3187 242.672
R12716 gnd.n3274 gnd.n3188 242.672
R12717 gnd.n3274 gnd.n3189 242.672
R12718 gnd.n3274 gnd.n3190 242.672
R12719 gnd.n3274 gnd.n3191 242.672
R12720 gnd.n3274 gnd.n3192 242.672
R12721 gnd.n3274 gnd.n3193 242.672
R12722 gnd.n3274 gnd.n3194 242.672
R12723 gnd.n3275 gnd.n3274 242.672
R12724 gnd.n4127 gnd.n2663 242.672
R12725 gnd.n4127 gnd.n2662 242.672
R12726 gnd.n4127 gnd.n2661 242.672
R12727 gnd.n4127 gnd.n2660 242.672
R12728 gnd.n4127 gnd.n2659 242.672
R12729 gnd.n4127 gnd.n2658 242.672
R12730 gnd.n4127 gnd.n2657 242.672
R12731 gnd.n4127 gnd.n2656 242.672
R12732 gnd.n4127 gnd.n2655 242.672
R12733 gnd.n4127 gnd.n2654 242.672
R12734 gnd.n4127 gnd.n2653 242.672
R12735 gnd.n4127 gnd.n2652 242.672
R12736 gnd.n4127 gnd.n2651 242.672
R12737 gnd.n6080 gnd.n1494 242.672
R12738 gnd.n6080 gnd.n1496 242.672
R12739 gnd.n6080 gnd.n1497 242.672
R12740 gnd.n6080 gnd.n1499 242.672
R12741 gnd.n6080 gnd.n1501 242.672
R12742 gnd.n6080 gnd.n1502 242.672
R12743 gnd.n6080 gnd.n1504 242.672
R12744 gnd.n6080 gnd.n1506 242.672
R12745 gnd.n6081 gnd.n6080 242.672
R12746 gnd.n347 gnd.n212 242.672
R12747 gnd.n7408 gnd.n212 242.672
R12748 gnd.n343 gnd.n212 242.672
R12749 gnd.n7415 gnd.n212 242.672
R12750 gnd.n336 gnd.n212 242.672
R12751 gnd.n7422 gnd.n212 242.672
R12752 gnd.n329 gnd.n212 242.672
R12753 gnd.n7429 gnd.n212 242.672
R12754 gnd.n322 gnd.n212 242.672
R12755 gnd.n3358 gnd.n3357 242.672
R12756 gnd.n3357 gnd.n3096 242.672
R12757 gnd.n3357 gnd.n3097 242.672
R12758 gnd.n3357 gnd.n3098 242.672
R12759 gnd.n3357 gnd.n3099 242.672
R12760 gnd.n3357 gnd.n3100 242.672
R12761 gnd.n3357 gnd.n3101 242.672
R12762 gnd.n3357 gnd.n3102 242.672
R12763 gnd.n4127 gnd.n2664 242.672
R12764 gnd.n4127 gnd.n2665 242.672
R12765 gnd.n4127 gnd.n2666 242.672
R12766 gnd.n4127 gnd.n2667 242.672
R12767 gnd.n4127 gnd.n2668 242.672
R12768 gnd.n4127 gnd.n2669 242.672
R12769 gnd.n4127 gnd.n2670 242.672
R12770 gnd.n4127 gnd.n2671 242.672
R12771 gnd.n4441 gnd.n4440 242.672
R12772 gnd.n4441 gnd.n4128 242.672
R12773 gnd.n4441 gnd.n4129 242.672
R12774 gnd.n4441 gnd.n4130 242.672
R12775 gnd.n4441 gnd.n4131 242.672
R12776 gnd.n4441 gnd.n4132 242.672
R12777 gnd.n4441 gnd.n4133 242.672
R12778 gnd.n4441 gnd.n4134 242.672
R12779 gnd.n4441 gnd.n4135 242.672
R12780 gnd.n4441 gnd.n4136 242.672
R12781 gnd.n4441 gnd.n4137 242.672
R12782 gnd.n4441 gnd.n4138 242.672
R12783 gnd.n4441 gnd.n4139 242.672
R12784 gnd.n4441 gnd.n4140 242.672
R12785 gnd.n4441 gnd.n4141 242.672
R12786 gnd.n4441 gnd.n4142 242.672
R12787 gnd.n4441 gnd.n4143 242.672
R12788 gnd.n4441 gnd.n4144 242.672
R12789 gnd.n4441 gnd.n4145 242.672
R12790 gnd.n4441 gnd.n4146 242.672
R12791 gnd.n4441 gnd.n4147 242.672
R12792 gnd.n4441 gnd.n4148 242.672
R12793 gnd.n4441 gnd.n4149 242.672
R12794 gnd.n4441 gnd.n4150 242.672
R12795 gnd.n4441 gnd.n4151 242.672
R12796 gnd.n4441 gnd.n4152 242.672
R12797 gnd.n4441 gnd.n4153 242.672
R12798 gnd.n4441 gnd.n4154 242.672
R12799 gnd.n4442 gnd.n4441 242.672
R12800 gnd.n2385 gnd.n1073 242.672
R12801 gnd.n2281 gnd.n1073 242.672
R12802 gnd.n2375 gnd.n1073 242.672
R12803 gnd.n2285 gnd.n1073 242.672
R12804 gnd.n2365 gnd.n1073 242.672
R12805 gnd.n2289 gnd.n1073 242.672
R12806 gnd.n2355 gnd.n1073 242.672
R12807 gnd.n2293 gnd.n1073 242.672
R12808 gnd.n2345 gnd.n1073 242.672
R12809 gnd.n2297 gnd.n1073 242.672
R12810 gnd.n2335 gnd.n1073 242.672
R12811 gnd.n2303 gnd.n1073 242.672
R12812 gnd.n2325 gnd.n1073 242.672
R12813 gnd.n2307 gnd.n1073 242.672
R12814 gnd.n2315 gnd.n1073 242.672
R12815 gnd.n2312 gnd.n1073 242.672
R12816 gnd.n6359 gnd.n1119 242.672
R12817 gnd.n1118 gnd.n1073 242.672
R12818 gnd.n6363 gnd.n1073 242.672
R12819 gnd.n1112 gnd.n1073 242.672
R12820 gnd.n6370 gnd.n1073 242.672
R12821 gnd.n1105 gnd.n1073 242.672
R12822 gnd.n6378 gnd.n1073 242.672
R12823 gnd.n1096 gnd.n1073 242.672
R12824 gnd.n6385 gnd.n1073 242.672
R12825 gnd.n1089 gnd.n1073 242.672
R12826 gnd.n6392 gnd.n1073 242.672
R12827 gnd.n1082 gnd.n1073 242.672
R12828 gnd.n6399 gnd.n1073 242.672
R12829 gnd.n6402 gnd.n1073 242.672
R12830 gnd.n6080 gnd.n6079 242.672
R12831 gnd.n6080 gnd.n1466 242.672
R12832 gnd.n6080 gnd.n1467 242.672
R12833 gnd.n6080 gnd.n1468 242.672
R12834 gnd.n6080 gnd.n1469 242.672
R12835 gnd.n6080 gnd.n1470 242.672
R12836 gnd.n6080 gnd.n1471 242.672
R12837 gnd.n6080 gnd.n1472 242.672
R12838 gnd.n6080 gnd.n1473 242.672
R12839 gnd.n6080 gnd.n1474 242.672
R12840 gnd.n6080 gnd.n1475 242.672
R12841 gnd.n6080 gnd.n1476 242.672
R12842 gnd.n6080 gnd.n1477 242.672
R12843 gnd.n6027 gnd.n1540 242.672
R12844 gnd.n6080 gnd.n1478 242.672
R12845 gnd.n6080 gnd.n1479 242.672
R12846 gnd.n6080 gnd.n1480 242.672
R12847 gnd.n6080 gnd.n1481 242.672
R12848 gnd.n6080 gnd.n1482 242.672
R12849 gnd.n6080 gnd.n1483 242.672
R12850 gnd.n6080 gnd.n1484 242.672
R12851 gnd.n6080 gnd.n1485 242.672
R12852 gnd.n6080 gnd.n1486 242.672
R12853 gnd.n6080 gnd.n1487 242.672
R12854 gnd.n6080 gnd.n1488 242.672
R12855 gnd.n6080 gnd.n1489 242.672
R12856 gnd.n6080 gnd.n1490 242.672
R12857 gnd.n6080 gnd.n1491 242.672
R12858 gnd.n6080 gnd.n1492 242.672
R12859 gnd.n6080 gnd.n1493 242.672
R12860 gnd.n7440 gnd.n212 242.672
R12861 gnd.n316 gnd.n212 242.672
R12862 gnd.n7447 gnd.n212 242.672
R12863 gnd.n307 gnd.n212 242.672
R12864 gnd.n7454 gnd.n212 242.672
R12865 gnd.n300 gnd.n212 242.672
R12866 gnd.n7461 gnd.n212 242.672
R12867 gnd.n293 gnd.n212 242.672
R12868 gnd.n7468 gnd.n212 242.672
R12869 gnd.n7471 gnd.n212 242.672
R12870 gnd.n284 gnd.n212 242.672
R12871 gnd.n7480 gnd.n212 242.672
R12872 gnd.n275 gnd.n212 242.672
R12873 gnd.n7487 gnd.n212 242.672
R12874 gnd.n268 gnd.n212 242.672
R12875 gnd.n7494 gnd.n212 242.672
R12876 gnd.n261 gnd.n212 242.672
R12877 gnd.n7501 gnd.n212 242.672
R12878 gnd.n254 gnd.n212 242.672
R12879 gnd.n7508 gnd.n212 242.672
R12880 gnd.n247 gnd.n212 242.672
R12881 gnd.n7518 gnd.n212 242.672
R12882 gnd.n240 gnd.n212 242.672
R12883 gnd.n7525 gnd.n212 242.672
R12884 gnd.n233 gnd.n212 242.672
R12885 gnd.n7532 gnd.n212 242.672
R12886 gnd.n226 gnd.n212 242.672
R12887 gnd.n7539 gnd.n212 242.672
R12888 gnd.n219 gnd.n212 242.672
R12889 gnd.n4857 gnd.n4856 242.672
R12890 gnd.n4857 gnd.n2204 242.672
R12891 gnd.n4857 gnd.n2205 242.672
R12892 gnd.n4857 gnd.n2206 242.672
R12893 gnd.n4857 gnd.n2207 242.672
R12894 gnd.n4857 gnd.n2208 242.672
R12895 gnd.n4857 gnd.n2209 242.672
R12896 gnd.n4857 gnd.n2210 242.672
R12897 gnd.n4857 gnd.n2211 242.672
R12898 gnd.n4857 gnd.n2212 242.672
R12899 gnd.n4857 gnd.n2213 242.672
R12900 gnd.n4857 gnd.n2214 242.672
R12901 gnd.n4857 gnd.n2215 242.672
R12902 gnd.n4857 gnd.n2216 242.672
R12903 gnd.n5727 gnd.n1760 242.672
R12904 gnd.n5727 gnd.n1758 242.672
R12905 gnd.n5727 gnd.n1757 242.672
R12906 gnd.n5727 gnd.n1755 242.672
R12907 gnd.n5727 gnd.n1753 242.672
R12908 gnd.n5727 gnd.n1752 242.672
R12909 gnd.n5727 gnd.n1750 242.672
R12910 gnd.n5727 gnd.n1748 242.672
R12911 gnd.n5727 gnd.n1747 242.672
R12912 gnd.n5727 gnd.n1745 242.672
R12913 gnd.n5727 gnd.n1744 242.672
R12914 gnd.n5727 gnd.n1742 242.672
R12915 gnd.n5728 gnd.n5727 242.672
R12916 gnd.n5727 gnd.n1763 242.672
R12917 gnd.n216 gnd.n213 240.244
R12918 gnd.n7541 gnd.n7540 240.244
R12919 gnd.n7538 gnd.n220 240.244
R12920 gnd.n7534 gnd.n7533 240.244
R12921 gnd.n7531 gnd.n227 240.244
R12922 gnd.n7527 gnd.n7526 240.244
R12923 gnd.n7524 gnd.n234 240.244
R12924 gnd.n7520 gnd.n7519 240.244
R12925 gnd.n7517 gnd.n241 240.244
R12926 gnd.n7510 gnd.n7509 240.244
R12927 gnd.n7507 gnd.n248 240.244
R12928 gnd.n7503 gnd.n7502 240.244
R12929 gnd.n7500 gnd.n255 240.244
R12930 gnd.n7496 gnd.n7495 240.244
R12931 gnd.n7493 gnd.n262 240.244
R12932 gnd.n7489 gnd.n7488 240.244
R12933 gnd.n7486 gnd.n269 240.244
R12934 gnd.n7482 gnd.n7481 240.244
R12935 gnd.n7479 gnd.n276 240.244
R12936 gnd.n7472 gnd.n285 240.244
R12937 gnd.n7470 gnd.n7469 240.244
R12938 gnd.n7467 gnd.n287 240.244
R12939 gnd.n7463 gnd.n7462 240.244
R12940 gnd.n7460 gnd.n294 240.244
R12941 gnd.n7456 gnd.n7455 240.244
R12942 gnd.n7453 gnd.n301 240.244
R12943 gnd.n7449 gnd.n7448 240.244
R12944 gnd.n7446 gnd.n308 240.244
R12945 gnd.n7442 gnd.n7441 240.244
R12946 gnd.n5960 gnd.n1573 240.244
R12947 gnd.n5952 gnd.n1573 240.244
R12948 gnd.n5952 gnd.n1584 240.244
R12949 gnd.n1600 gnd.n1584 240.244
R12950 gnd.n5744 gnd.n1600 240.244
R12951 gnd.n5744 gnd.n1613 240.244
R12952 gnd.n5750 gnd.n1613 240.244
R12953 gnd.n5750 gnd.n1623 240.244
R12954 gnd.n5757 gnd.n1623 240.244
R12955 gnd.n5757 gnd.n1633 240.244
R12956 gnd.n1720 gnd.n1633 240.244
R12957 gnd.n1720 gnd.n1643 240.244
R12958 gnd.n5830 gnd.n1643 240.244
R12959 gnd.n5830 gnd.n1653 240.244
R12960 gnd.n5835 gnd.n1653 240.244
R12961 gnd.n5835 gnd.n1663 240.244
R12962 gnd.n5845 gnd.n1663 240.244
R12963 gnd.n5845 gnd.n1673 240.244
R12964 gnd.n1706 gnd.n1673 240.244
R12965 gnd.n1706 gnd.n1683 240.244
R12966 gnd.n5857 gnd.n1683 240.244
R12967 gnd.n5857 gnd.n1693 240.244
R12968 gnd.n1697 gnd.n1693 240.244
R12969 gnd.n5852 gnd.n1697 240.244
R12970 gnd.n5852 gnd.n382 240.244
R12971 gnd.n382 gnd.n376 240.244
R12972 gnd.n7307 gnd.n376 240.244
R12973 gnd.n7307 gnd.n89 240.244
R12974 gnd.n369 gnd.n89 240.244
R12975 gnd.n7356 gnd.n369 240.244
R12976 gnd.n7356 gnd.n105 240.244
R12977 gnd.n7352 gnd.n105 240.244
R12978 gnd.n7352 gnd.n116 240.244
R12979 gnd.n7349 gnd.n116 240.244
R12980 gnd.n7349 gnd.n125 240.244
R12981 gnd.n7346 gnd.n125 240.244
R12982 gnd.n7346 gnd.n134 240.244
R12983 gnd.n7343 gnd.n134 240.244
R12984 gnd.n7343 gnd.n144 240.244
R12985 gnd.n7340 gnd.n144 240.244
R12986 gnd.n7340 gnd.n153 240.244
R12987 gnd.n7337 gnd.n153 240.244
R12988 gnd.n7337 gnd.n163 240.244
R12989 gnd.n7334 gnd.n163 240.244
R12990 gnd.n7334 gnd.n172 240.244
R12991 gnd.n7331 gnd.n172 240.244
R12992 gnd.n7331 gnd.n182 240.244
R12993 gnd.n7328 gnd.n182 240.244
R12994 gnd.n7328 gnd.n192 240.244
R12995 gnd.n7325 gnd.n192 240.244
R12996 gnd.n7325 gnd.n202 240.244
R12997 gnd.n7322 gnd.n202 240.244
R12998 gnd.n7322 gnd.n210 240.244
R12999 gnd.n1509 gnd.n1508 240.244
R13000 gnd.n6073 gnd.n1508 240.244
R13001 gnd.n6071 gnd.n6070 240.244
R13002 gnd.n6067 gnd.n6066 240.244
R13003 gnd.n6063 gnd.n6062 240.244
R13004 gnd.n6059 gnd.n6058 240.244
R13005 gnd.n6055 gnd.n6054 240.244
R13006 gnd.n6051 gnd.n6050 240.244
R13007 gnd.n6047 gnd.n6046 240.244
R13008 gnd.n6042 gnd.n6041 240.244
R13009 gnd.n6038 gnd.n6037 240.244
R13010 gnd.n6034 gnd.n6033 240.244
R13011 gnd.n6030 gnd.n6029 240.244
R13012 gnd.n6025 gnd.n6024 240.244
R13013 gnd.n6021 gnd.n6020 240.244
R13014 gnd.n6017 gnd.n6016 240.244
R13015 gnd.n6013 gnd.n6012 240.244
R13016 gnd.n6009 gnd.n6008 240.244
R13017 gnd.n6005 gnd.n6004 240.244
R13018 gnd.n6001 gnd.n6000 240.244
R13019 gnd.n5997 gnd.n5996 240.244
R13020 gnd.n5993 gnd.n5992 240.244
R13021 gnd.n5989 gnd.n5988 240.244
R13022 gnd.n5985 gnd.n5984 240.244
R13023 gnd.n5981 gnd.n5980 240.244
R13024 gnd.n5977 gnd.n5976 240.244
R13025 gnd.n5973 gnd.n5972 240.244
R13026 gnd.n5969 gnd.n5968 240.244
R13027 gnd.n1588 gnd.n1510 240.244
R13028 gnd.n5950 gnd.n1588 240.244
R13029 gnd.n5950 gnd.n1589 240.244
R13030 gnd.n5946 gnd.n1589 240.244
R13031 gnd.n5946 gnd.n1598 240.244
R13032 gnd.n5938 gnd.n1598 240.244
R13033 gnd.n5938 gnd.n1615 240.244
R13034 gnd.n5934 gnd.n1615 240.244
R13035 gnd.n5934 gnd.n1621 240.244
R13036 gnd.n5926 gnd.n1621 240.244
R13037 gnd.n5926 gnd.n1636 240.244
R13038 gnd.n5922 gnd.n1636 240.244
R13039 gnd.n5922 gnd.n1642 240.244
R13040 gnd.n5914 gnd.n1642 240.244
R13041 gnd.n5914 gnd.n1655 240.244
R13042 gnd.n5910 gnd.n1655 240.244
R13043 gnd.n5910 gnd.n1661 240.244
R13044 gnd.n5902 gnd.n1661 240.244
R13045 gnd.n5902 gnd.n1676 240.244
R13046 gnd.n5898 gnd.n1676 240.244
R13047 gnd.n5898 gnd.n1682 240.244
R13048 gnd.n5890 gnd.n1682 240.244
R13049 gnd.n5890 gnd.n5888 240.244
R13050 gnd.n5888 gnd.n384 240.244
R13051 gnd.n7298 gnd.n384 240.244
R13052 gnd.n7298 gnd.n7296 240.244
R13053 gnd.n7296 gnd.n92 240.244
R13054 gnd.n7622 gnd.n92 240.244
R13055 gnd.n7622 gnd.n93 240.244
R13056 gnd.n103 gnd.n93 240.244
R13057 gnd.n7616 gnd.n103 240.244
R13058 gnd.n7616 gnd.n104 240.244
R13059 gnd.n7608 gnd.n104 240.244
R13060 gnd.n7608 gnd.n118 240.244
R13061 gnd.n7604 gnd.n118 240.244
R13062 gnd.n7604 gnd.n123 240.244
R13063 gnd.n7596 gnd.n123 240.244
R13064 gnd.n7596 gnd.n137 240.244
R13065 gnd.n7592 gnd.n137 240.244
R13066 gnd.n7592 gnd.n143 240.244
R13067 gnd.n7584 gnd.n143 240.244
R13068 gnd.n7584 gnd.n155 240.244
R13069 gnd.n7580 gnd.n155 240.244
R13070 gnd.n7580 gnd.n161 240.244
R13071 gnd.n7572 gnd.n161 240.244
R13072 gnd.n7572 gnd.n175 240.244
R13073 gnd.n7568 gnd.n175 240.244
R13074 gnd.n7568 gnd.n181 240.244
R13075 gnd.n7560 gnd.n181 240.244
R13076 gnd.n7560 gnd.n195 240.244
R13077 gnd.n7556 gnd.n195 240.244
R13078 gnd.n7556 gnd.n201 240.244
R13079 gnd.n7548 gnd.n201 240.244
R13080 gnd.n6403 gnd.n1069 240.244
R13081 gnd.n6401 gnd.n6400 240.244
R13082 gnd.n6398 gnd.n1075 240.244
R13083 gnd.n6394 gnd.n6393 240.244
R13084 gnd.n6391 gnd.n1083 240.244
R13085 gnd.n6387 gnd.n6386 240.244
R13086 gnd.n6384 gnd.n1090 240.244
R13087 gnd.n6380 gnd.n6379 240.244
R13088 gnd.n6377 gnd.n1097 240.244
R13089 gnd.n6372 gnd.n6371 240.244
R13090 gnd.n6369 gnd.n1106 240.244
R13091 gnd.n6365 gnd.n6364 240.244
R13092 gnd.n6362 gnd.n1113 240.244
R13093 gnd.n2314 gnd.n2313 240.244
R13094 gnd.n2317 gnd.n2316 240.244
R13095 gnd.n2324 gnd.n2323 240.244
R13096 gnd.n2327 gnd.n2326 240.244
R13097 gnd.n2334 gnd.n2333 240.244
R13098 gnd.n2337 gnd.n2336 240.244
R13099 gnd.n2344 gnd.n2343 240.244
R13100 gnd.n2347 gnd.n2346 240.244
R13101 gnd.n2354 gnd.n2353 240.244
R13102 gnd.n2357 gnd.n2356 240.244
R13103 gnd.n2364 gnd.n2363 240.244
R13104 gnd.n2367 gnd.n2366 240.244
R13105 gnd.n2374 gnd.n2373 240.244
R13106 gnd.n2377 gnd.n2376 240.244
R13107 gnd.n2384 gnd.n2383 240.244
R13108 gnd.n4444 gnd.n2637 240.244
R13109 gnd.n2637 gnd.n2627 240.244
R13110 gnd.n4460 gnd.n2627 240.244
R13111 gnd.n4461 gnd.n4460 240.244
R13112 gnd.n4461 gnd.n2618 240.244
R13113 gnd.n2618 gnd.n2609 240.244
R13114 gnd.n4480 gnd.n2609 240.244
R13115 gnd.n4481 gnd.n4480 240.244
R13116 gnd.n4481 gnd.n2601 240.244
R13117 gnd.n2601 gnd.n2591 240.244
R13118 gnd.n4500 gnd.n2591 240.244
R13119 gnd.n4501 gnd.n4500 240.244
R13120 gnd.n4501 gnd.n2581 240.244
R13121 gnd.n4504 gnd.n2581 240.244
R13122 gnd.n4504 gnd.n2572 240.244
R13123 gnd.n2572 gnd.n2565 240.244
R13124 gnd.n4546 gnd.n2565 240.244
R13125 gnd.n4546 gnd.n2556 240.244
R13126 gnd.n2556 gnd.n2548 240.244
R13127 gnd.n4566 gnd.n2548 240.244
R13128 gnd.n4567 gnd.n4566 240.244
R13129 gnd.n4567 gnd.n2541 240.244
R13130 gnd.n2541 gnd.n2536 240.244
R13131 gnd.n4571 gnd.n2536 240.244
R13132 gnd.n4571 gnd.n939 240.244
R13133 gnd.n4601 gnd.n939 240.244
R13134 gnd.n4601 gnd.n2521 240.244
R13135 gnd.n4604 gnd.n2521 240.244
R13136 gnd.n4604 gnd.n2517 240.244
R13137 gnd.n2517 gnd.n2507 240.244
R13138 gnd.n2507 gnd.n956 240.244
R13139 gnd.n4658 gnd.n956 240.244
R13140 gnd.n4658 gnd.n968 240.244
R13141 gnd.n4663 gnd.n968 240.244
R13142 gnd.n4663 gnd.n977 240.244
R13143 gnd.n4673 gnd.n977 240.244
R13144 gnd.n4673 gnd.n987 240.244
R13145 gnd.n2487 gnd.n987 240.244
R13146 gnd.n2487 gnd.n997 240.244
R13147 gnd.n4680 gnd.n997 240.244
R13148 gnd.n4680 gnd.n1007 240.244
R13149 gnd.n4686 gnd.n1007 240.244
R13150 gnd.n4686 gnd.n1017 240.244
R13151 gnd.n4690 gnd.n1017 240.244
R13152 gnd.n4690 gnd.n1027 240.244
R13153 gnd.n4757 gnd.n1027 240.244
R13154 gnd.n4757 gnd.n1037 240.244
R13155 gnd.n4761 gnd.n1037 240.244
R13156 gnd.n4761 gnd.n1047 240.244
R13157 gnd.n4772 gnd.n1047 240.244
R13158 gnd.n4772 gnd.n1058 240.244
R13159 gnd.n4777 gnd.n1058 240.244
R13160 gnd.n4777 gnd.n1066 240.244
R13161 gnd.n4166 gnd.n4165 240.244
R13162 gnd.n4434 gnd.n4165 240.244
R13163 gnd.n4432 gnd.n4431 240.244
R13164 gnd.n4428 gnd.n4427 240.244
R13165 gnd.n4424 gnd.n4423 240.244
R13166 gnd.n4420 gnd.n4419 240.244
R13167 gnd.n4416 gnd.n4415 240.244
R13168 gnd.n4412 gnd.n4411 240.244
R13169 gnd.n4408 gnd.n4407 240.244
R13170 gnd.n4403 gnd.n4402 240.244
R13171 gnd.n4399 gnd.n4398 240.244
R13172 gnd.n4395 gnd.n4394 240.244
R13173 gnd.n4391 gnd.n4390 240.244
R13174 gnd.n4387 gnd.n4386 240.244
R13175 gnd.n4383 gnd.n4382 240.244
R13176 gnd.n4379 gnd.n4378 240.244
R13177 gnd.n4375 gnd.n4374 240.244
R13178 gnd.n4371 gnd.n4370 240.244
R13179 gnd.n4367 gnd.n4366 240.244
R13180 gnd.n4363 gnd.n4362 240.244
R13181 gnd.n4359 gnd.n4358 240.244
R13182 gnd.n4355 gnd.n4354 240.244
R13183 gnd.n4351 gnd.n4350 240.244
R13184 gnd.n4347 gnd.n4346 240.244
R13185 gnd.n4343 gnd.n4342 240.244
R13186 gnd.n4339 gnd.n4338 240.244
R13187 gnd.n4335 gnd.n4334 240.244
R13188 gnd.n4331 gnd.n4330 240.244
R13189 gnd.n4327 gnd.n2648 240.244
R13190 gnd.n4452 gnd.n2635 240.244
R13191 gnd.n4452 gnd.n2631 240.244
R13192 gnd.n4458 gnd.n2631 240.244
R13193 gnd.n4458 gnd.n2616 240.244
R13194 gnd.n4472 gnd.n2616 240.244
R13195 gnd.n4472 gnd.n2612 240.244
R13196 gnd.n4478 gnd.n2612 240.244
R13197 gnd.n4478 gnd.n2599 240.244
R13198 gnd.n4492 gnd.n2599 240.244
R13199 gnd.n4492 gnd.n2595 240.244
R13200 gnd.n4498 gnd.n2595 240.244
R13201 gnd.n4498 gnd.n2579 240.244
R13202 gnd.n4516 gnd.n2579 240.244
R13203 gnd.n4516 gnd.n2574 240.244
R13204 gnd.n4524 gnd.n2574 240.244
R13205 gnd.n4524 gnd.n2575 240.244
R13206 gnd.n2575 gnd.n2555 240.244
R13207 gnd.n4557 gnd.n2555 240.244
R13208 gnd.n4557 gnd.n2551 240.244
R13209 gnd.n4564 gnd.n2551 240.244
R13210 gnd.n4564 gnd.n2538 240.244
R13211 gnd.n4582 gnd.n2538 240.244
R13212 gnd.n4584 gnd.n4582 240.244
R13213 gnd.n4584 gnd.n942 240.244
R13214 gnd.n6482 gnd.n942 240.244
R13215 gnd.n6482 gnd.n943 240.244
R13216 gnd.n4614 gnd.n943 240.244
R13217 gnd.n4615 gnd.n4614 240.244
R13218 gnd.n4618 gnd.n4615 240.244
R13219 gnd.n4618 gnd.n954 240.244
R13220 gnd.n6477 gnd.n954 240.244
R13221 gnd.n6477 gnd.n955 240.244
R13222 gnd.n6469 gnd.n955 240.244
R13223 gnd.n6469 gnd.n970 240.244
R13224 gnd.n6465 gnd.n970 240.244
R13225 gnd.n6465 gnd.n975 240.244
R13226 gnd.n6457 gnd.n975 240.244
R13227 gnd.n6457 gnd.n990 240.244
R13228 gnd.n6453 gnd.n990 240.244
R13229 gnd.n6453 gnd.n996 240.244
R13230 gnd.n6445 gnd.n996 240.244
R13231 gnd.n6445 gnd.n1009 240.244
R13232 gnd.n6441 gnd.n1009 240.244
R13233 gnd.n6441 gnd.n1015 240.244
R13234 gnd.n6433 gnd.n1015 240.244
R13235 gnd.n6433 gnd.n1030 240.244
R13236 gnd.n6429 gnd.n1030 240.244
R13237 gnd.n6429 gnd.n1036 240.244
R13238 gnd.n6421 gnd.n1036 240.244
R13239 gnd.n6421 gnd.n1050 240.244
R13240 gnd.n6417 gnd.n1050 240.244
R13241 gnd.n6417 gnd.n1056 240.244
R13242 gnd.n6409 gnd.n1056 240.244
R13243 gnd.n4126 gnd.n2673 240.244
R13244 gnd.n4119 gnd.n4118 240.244
R13245 gnd.n4116 gnd.n4115 240.244
R13246 gnd.n4112 gnd.n4111 240.244
R13247 gnd.n4108 gnd.n4107 240.244
R13248 gnd.n4104 gnd.n4103 240.244
R13249 gnd.n4100 gnd.n4099 240.244
R13250 gnd.n4096 gnd.n4095 240.244
R13251 gnd.n3369 gnd.n3081 240.244
R13252 gnd.n3379 gnd.n3081 240.244
R13253 gnd.n3379 gnd.n3072 240.244
R13254 gnd.n3072 gnd.n3061 240.244
R13255 gnd.n3400 gnd.n3061 240.244
R13256 gnd.n3400 gnd.n3055 240.244
R13257 gnd.n3410 gnd.n3055 240.244
R13258 gnd.n3410 gnd.n3044 240.244
R13259 gnd.n3044 gnd.n3036 240.244
R13260 gnd.n3428 gnd.n3036 240.244
R13261 gnd.n3429 gnd.n3428 240.244
R13262 gnd.n3429 gnd.n3021 240.244
R13263 gnd.n3431 gnd.n3021 240.244
R13264 gnd.n3431 gnd.n3007 240.244
R13265 gnd.n3473 gnd.n3007 240.244
R13266 gnd.n3474 gnd.n3473 240.244
R13267 gnd.n3477 gnd.n3474 240.244
R13268 gnd.n3477 gnd.n2962 240.244
R13269 gnd.n3002 gnd.n2962 240.244
R13270 gnd.n3002 gnd.n2972 240.244
R13271 gnd.n3487 gnd.n2972 240.244
R13272 gnd.n3487 gnd.n2993 240.244
R13273 gnd.n3497 gnd.n2993 240.244
R13274 gnd.n3497 gnd.n2875 240.244
R13275 gnd.n3542 gnd.n2875 240.244
R13276 gnd.n3542 gnd.n2861 240.244
R13277 gnd.n3564 gnd.n2861 240.244
R13278 gnd.n3565 gnd.n3564 240.244
R13279 gnd.n3565 gnd.n2848 240.244
R13280 gnd.n2848 gnd.n2837 240.244
R13281 gnd.n3596 gnd.n2837 240.244
R13282 gnd.n3597 gnd.n3596 240.244
R13283 gnd.n3598 gnd.n3597 240.244
R13284 gnd.n3598 gnd.n2822 240.244
R13285 gnd.n2822 gnd.n2821 240.244
R13286 gnd.n2821 gnd.n2806 240.244
R13287 gnd.n3649 gnd.n2806 240.244
R13288 gnd.n3650 gnd.n3649 240.244
R13289 gnd.n3650 gnd.n2793 240.244
R13290 gnd.n2793 gnd.n2782 240.244
R13291 gnd.n3681 gnd.n2782 240.244
R13292 gnd.n3682 gnd.n3681 240.244
R13293 gnd.n3683 gnd.n3682 240.244
R13294 gnd.n3683 gnd.n2766 240.244
R13295 gnd.n2766 gnd.n2765 240.244
R13296 gnd.n2765 gnd.n2752 240.244
R13297 gnd.n3738 gnd.n2752 240.244
R13298 gnd.n3739 gnd.n3738 240.244
R13299 gnd.n3739 gnd.n2739 240.244
R13300 gnd.n2739 gnd.n2729 240.244
R13301 gnd.n4027 gnd.n2729 240.244
R13302 gnd.n4030 gnd.n4027 240.244
R13303 gnd.n4030 gnd.n4029 240.244
R13304 gnd.n3359 gnd.n3094 240.244
R13305 gnd.n3115 gnd.n3094 240.244
R13306 gnd.n3118 gnd.n3117 240.244
R13307 gnd.n3125 gnd.n3124 240.244
R13308 gnd.n3128 gnd.n3127 240.244
R13309 gnd.n3135 gnd.n3134 240.244
R13310 gnd.n3138 gnd.n3137 240.244
R13311 gnd.n3145 gnd.n3144 240.244
R13312 gnd.n3367 gnd.n3091 240.244
R13313 gnd.n3091 gnd.n3070 240.244
R13314 gnd.n3390 gnd.n3070 240.244
R13315 gnd.n3390 gnd.n3064 240.244
R13316 gnd.n3398 gnd.n3064 240.244
R13317 gnd.n3398 gnd.n3066 240.244
R13318 gnd.n3066 gnd.n3042 240.244
R13319 gnd.n3420 gnd.n3042 240.244
R13320 gnd.n3420 gnd.n3038 240.244
R13321 gnd.n3426 gnd.n3038 240.244
R13322 gnd.n3426 gnd.n3020 240.244
R13323 gnd.n3451 gnd.n3020 240.244
R13324 gnd.n3451 gnd.n3015 240.244
R13325 gnd.n3463 gnd.n3015 240.244
R13326 gnd.n3463 gnd.n3016 240.244
R13327 gnd.n3459 gnd.n3016 240.244
R13328 gnd.n3459 gnd.n2964 240.244
R13329 gnd.n3511 gnd.n2964 240.244
R13330 gnd.n3511 gnd.n2965 240.244
R13331 gnd.n3507 gnd.n2965 240.244
R13332 gnd.n3507 gnd.n2971 240.244
R13333 gnd.n2991 gnd.n2971 240.244
R13334 gnd.n2991 gnd.n2873 240.244
R13335 gnd.n3546 gnd.n2873 240.244
R13336 gnd.n3546 gnd.n2868 240.244
R13337 gnd.n3554 gnd.n2868 240.244
R13338 gnd.n3554 gnd.n2869 240.244
R13339 gnd.n2869 gnd.n2846 240.244
R13340 gnd.n3586 gnd.n2846 240.244
R13341 gnd.n3586 gnd.n2841 240.244
R13342 gnd.n3594 gnd.n2841 240.244
R13343 gnd.n3594 gnd.n2842 240.244
R13344 gnd.n2842 gnd.n2819 240.244
R13345 gnd.n3631 gnd.n2819 240.244
R13346 gnd.n3631 gnd.n2814 240.244
R13347 gnd.n3639 gnd.n2814 240.244
R13348 gnd.n3639 gnd.n2815 240.244
R13349 gnd.n2815 gnd.n2791 240.244
R13350 gnd.n3671 gnd.n2791 240.244
R13351 gnd.n3671 gnd.n2786 240.244
R13352 gnd.n3679 gnd.n2786 240.244
R13353 gnd.n3679 gnd.n2787 240.244
R13354 gnd.n2787 gnd.n2764 240.244
R13355 gnd.n3720 gnd.n2764 240.244
R13356 gnd.n3720 gnd.n2759 240.244
R13357 gnd.n3728 gnd.n2759 240.244
R13358 gnd.n3728 gnd.n2760 240.244
R13359 gnd.n2760 gnd.n2737 240.244
R13360 gnd.n4015 gnd.n2737 240.244
R13361 gnd.n4015 gnd.n2732 240.244
R13362 gnd.n4025 gnd.n2732 240.244
R13363 gnd.n4025 gnd.n2733 240.244
R13364 gnd.n2733 gnd.n2672 240.244
R13365 gnd.n319 gnd.n208 240.244
R13366 gnd.n7431 gnd.n7430 240.244
R13367 gnd.n7428 gnd.n323 240.244
R13368 gnd.n7424 gnd.n7423 240.244
R13369 gnd.n7421 gnd.n330 240.244
R13370 gnd.n7417 gnd.n7416 240.244
R13371 gnd.n7414 gnd.n337 240.244
R13372 gnd.n7410 gnd.n7409 240.244
R13373 gnd.n7407 gnd.n344 240.244
R13374 gnd.n5774 gnd.n1576 240.244
R13375 gnd.n5774 gnd.n1585 240.244
R13376 gnd.n5737 gnd.n1585 240.244
R13377 gnd.n5737 gnd.n1601 240.244
R13378 gnd.n5738 gnd.n1601 240.244
R13379 gnd.n5738 gnd.n1614 240.244
R13380 gnd.n5741 gnd.n1614 240.244
R13381 gnd.n5741 gnd.n1624 240.244
R13382 gnd.n5759 gnd.n1624 240.244
R13383 gnd.n5759 gnd.n1634 240.244
R13384 gnd.n5822 gnd.n1634 240.244
R13385 gnd.n5822 gnd.n1644 240.244
R13386 gnd.n5828 gnd.n1644 240.244
R13387 gnd.n5828 gnd.n1654 240.244
R13388 gnd.n5837 gnd.n1654 240.244
R13389 gnd.n5837 gnd.n1664 240.244
R13390 gnd.n5843 gnd.n1664 240.244
R13391 gnd.n5843 gnd.n1674 240.244
R13392 gnd.n5873 gnd.n1674 240.244
R13393 gnd.n5873 gnd.n1684 240.244
R13394 gnd.n5859 gnd.n1684 240.244
R13395 gnd.n5859 gnd.n1694 240.244
R13396 gnd.n1698 gnd.n1694 240.244
R13397 gnd.n5860 gnd.n1698 240.244
R13398 gnd.n5860 gnd.n383 240.244
R13399 gnd.n7294 gnd.n383 240.244
R13400 gnd.n7294 gnd.n86 240.244
R13401 gnd.n7624 gnd.n86 240.244
R13402 gnd.n7624 gnd.n88 240.244
R13403 gnd.n7358 gnd.n88 240.244
R13404 gnd.n7358 gnd.n106 240.244
R13405 gnd.n7364 gnd.n106 240.244
R13406 gnd.n7364 gnd.n117 240.244
R13407 gnd.n365 gnd.n117 240.244
R13408 gnd.n365 gnd.n126 240.244
R13409 gnd.n7371 gnd.n126 240.244
R13410 gnd.n7371 gnd.n135 240.244
R13411 gnd.n362 gnd.n135 240.244
R13412 gnd.n362 gnd.n145 240.244
R13413 gnd.n7378 gnd.n145 240.244
R13414 gnd.n7378 gnd.n154 240.244
R13415 gnd.n359 gnd.n154 240.244
R13416 gnd.n359 gnd.n164 240.244
R13417 gnd.n7385 gnd.n164 240.244
R13418 gnd.n7385 gnd.n173 240.244
R13419 gnd.n356 gnd.n173 240.244
R13420 gnd.n356 gnd.n183 240.244
R13421 gnd.n7392 gnd.n183 240.244
R13422 gnd.n7392 gnd.n193 240.244
R13423 gnd.n353 gnd.n193 240.244
R13424 gnd.n353 gnd.n203 240.244
R13425 gnd.n7399 gnd.n203 240.244
R13426 gnd.n7399 gnd.n211 240.244
R13427 gnd.n1420 gnd.n1419 240.244
R13428 gnd.n1495 gnd.n1427 240.244
R13429 gnd.n1498 gnd.n1428 240.244
R13430 gnd.n1436 gnd.n1435 240.244
R13431 gnd.n1500 gnd.n1443 240.244
R13432 gnd.n1503 gnd.n1444 240.244
R13433 gnd.n1452 gnd.n1451 240.244
R13434 gnd.n1505 gnd.n1461 240.244
R13435 gnd.n6082 gnd.n1464 240.244
R13436 gnd.n5958 gnd.n1579 240.244
R13437 gnd.n1587 gnd.n1579 240.244
R13438 gnd.n1603 gnd.n1587 240.244
R13439 gnd.n5944 gnd.n1603 240.244
R13440 gnd.n5944 gnd.n1604 240.244
R13441 gnd.n5940 gnd.n1604 240.244
R13442 gnd.n5940 gnd.n1611 240.244
R13443 gnd.n5932 gnd.n1611 240.244
R13444 gnd.n5932 gnd.n1626 240.244
R13445 gnd.n5928 gnd.n1626 240.244
R13446 gnd.n5928 gnd.n1631 240.244
R13447 gnd.n5920 gnd.n1631 240.244
R13448 gnd.n5920 gnd.n1646 240.244
R13449 gnd.n5916 gnd.n1646 240.244
R13450 gnd.n5916 gnd.n1651 240.244
R13451 gnd.n5908 gnd.n1651 240.244
R13452 gnd.n5908 gnd.n1666 240.244
R13453 gnd.n5904 gnd.n1666 240.244
R13454 gnd.n5904 gnd.n1671 240.244
R13455 gnd.n5896 gnd.n1671 240.244
R13456 gnd.n5896 gnd.n1686 240.244
R13457 gnd.n5892 gnd.n1686 240.244
R13458 gnd.n5892 gnd.n1691 240.244
R13459 gnd.n1691 gnd.n380 240.244
R13460 gnd.n7300 gnd.n380 240.244
R13461 gnd.n7300 gnd.n374 240.244
R13462 gnd.n7309 gnd.n374 240.244
R13463 gnd.n7309 gnd.n91 240.244
R13464 gnd.n7312 gnd.n91 240.244
R13465 gnd.n7312 gnd.n108 240.244
R13466 gnd.n7614 gnd.n108 240.244
R13467 gnd.n7614 gnd.n109 240.244
R13468 gnd.n7610 gnd.n109 240.244
R13469 gnd.n7610 gnd.n115 240.244
R13470 gnd.n7602 gnd.n115 240.244
R13471 gnd.n7602 gnd.n127 240.244
R13472 gnd.n7598 gnd.n127 240.244
R13473 gnd.n7598 gnd.n132 240.244
R13474 gnd.n7590 gnd.n132 240.244
R13475 gnd.n7590 gnd.n147 240.244
R13476 gnd.n7586 gnd.n147 240.244
R13477 gnd.n7586 gnd.n152 240.244
R13478 gnd.n7578 gnd.n152 240.244
R13479 gnd.n7578 gnd.n165 240.244
R13480 gnd.n7574 gnd.n165 240.244
R13481 gnd.n7574 gnd.n170 240.244
R13482 gnd.n7566 gnd.n170 240.244
R13483 gnd.n7566 gnd.n185 240.244
R13484 gnd.n7562 gnd.n185 240.244
R13485 gnd.n7562 gnd.n190 240.244
R13486 gnd.n7554 gnd.n190 240.244
R13487 gnd.n7554 gnd.n204 240.244
R13488 gnd.n7550 gnd.n204 240.244
R13489 gnd.n2692 gnd.n2650 240.244
R13490 gnd.n4086 gnd.n4085 240.244
R13491 gnd.n4082 gnd.n4081 240.244
R13492 gnd.n4078 gnd.n4077 240.244
R13493 gnd.n4074 gnd.n4073 240.244
R13494 gnd.n4070 gnd.n4069 240.244
R13495 gnd.n4066 gnd.n4065 240.244
R13496 gnd.n4062 gnd.n4061 240.244
R13497 gnd.n4058 gnd.n4057 240.244
R13498 gnd.n4054 gnd.n4053 240.244
R13499 gnd.n4050 gnd.n4049 240.244
R13500 gnd.n4046 gnd.n4045 240.244
R13501 gnd.n4042 gnd.n4041 240.244
R13502 gnd.n3282 gnd.n3179 240.244
R13503 gnd.n3282 gnd.n3172 240.244
R13504 gnd.n3293 gnd.n3172 240.244
R13505 gnd.n3293 gnd.n3168 240.244
R13506 gnd.n3299 gnd.n3168 240.244
R13507 gnd.n3299 gnd.n3160 240.244
R13508 gnd.n3309 gnd.n3160 240.244
R13509 gnd.n3309 gnd.n3155 240.244
R13510 gnd.n3345 gnd.n3155 240.244
R13511 gnd.n3345 gnd.n3156 240.244
R13512 gnd.n3156 gnd.n3103 240.244
R13513 gnd.n3340 gnd.n3103 240.244
R13514 gnd.n3340 gnd.n3339 240.244
R13515 gnd.n3339 gnd.n3082 240.244
R13516 gnd.n3335 gnd.n3082 240.244
R13517 gnd.n3335 gnd.n3073 240.244
R13518 gnd.n3332 gnd.n3073 240.244
R13519 gnd.n3332 gnd.n3331 240.244
R13520 gnd.n3331 gnd.n3056 240.244
R13521 gnd.n3327 gnd.n3056 240.244
R13522 gnd.n3327 gnd.n3045 240.244
R13523 gnd.n3045 gnd.n3026 240.244
R13524 gnd.n3440 gnd.n3026 240.244
R13525 gnd.n3440 gnd.n3022 240.244
R13526 gnd.n3448 gnd.n3022 240.244
R13527 gnd.n3448 gnd.n3013 240.244
R13528 gnd.n3013 gnd.n2949 240.244
R13529 gnd.n3520 gnd.n2949 240.244
R13530 gnd.n3520 gnd.n2950 240.244
R13531 gnd.n2961 gnd.n2950 240.244
R13532 gnd.n2996 gnd.n2961 240.244
R13533 gnd.n2999 gnd.n2996 240.244
R13534 gnd.n2999 gnd.n2973 240.244
R13535 gnd.n2986 gnd.n2973 240.244
R13536 gnd.n2986 gnd.n2983 240.244
R13537 gnd.n2983 gnd.n2876 240.244
R13538 gnd.n3541 gnd.n2876 240.244
R13539 gnd.n3541 gnd.n2866 240.244
R13540 gnd.n3537 gnd.n2866 240.244
R13541 gnd.n3537 gnd.n2860 240.244
R13542 gnd.n3534 gnd.n2860 240.244
R13543 gnd.n3534 gnd.n2849 240.244
R13544 gnd.n3531 gnd.n2849 240.244
R13545 gnd.n3531 gnd.n2827 240.244
R13546 gnd.n3607 gnd.n2827 240.244
R13547 gnd.n3607 gnd.n2823 240.244
R13548 gnd.n3628 gnd.n2823 240.244
R13549 gnd.n3628 gnd.n2812 240.244
R13550 gnd.n3624 gnd.n2812 240.244
R13551 gnd.n3624 gnd.n2805 240.244
R13552 gnd.n3621 gnd.n2805 240.244
R13553 gnd.n3621 gnd.n2794 240.244
R13554 gnd.n3618 gnd.n2794 240.244
R13555 gnd.n3618 gnd.n2771 240.244
R13556 gnd.n3692 gnd.n2771 240.244
R13557 gnd.n3692 gnd.n2767 240.244
R13558 gnd.n3717 gnd.n2767 240.244
R13559 gnd.n3717 gnd.n2758 240.244
R13560 gnd.n3713 gnd.n2758 240.244
R13561 gnd.n3713 gnd.n2751 240.244
R13562 gnd.n3709 gnd.n2751 240.244
R13563 gnd.n3709 gnd.n2740 240.244
R13564 gnd.n3706 gnd.n2740 240.244
R13565 gnd.n3706 gnd.n2721 240.244
R13566 gnd.n4037 gnd.n2721 240.244
R13567 gnd.n3196 gnd.n3195 240.244
R13568 gnd.n3267 gnd.n3195 240.244
R13569 gnd.n3265 gnd.n3264 240.244
R13570 gnd.n3261 gnd.n3260 240.244
R13571 gnd.n3257 gnd.n3256 240.244
R13572 gnd.n3253 gnd.n3252 240.244
R13573 gnd.n3249 gnd.n3248 240.244
R13574 gnd.n3245 gnd.n3244 240.244
R13575 gnd.n3241 gnd.n3240 240.244
R13576 gnd.n3237 gnd.n3236 240.244
R13577 gnd.n3233 gnd.n3232 240.244
R13578 gnd.n3229 gnd.n3228 240.244
R13579 gnd.n3225 gnd.n3183 240.244
R13580 gnd.n3285 gnd.n3177 240.244
R13581 gnd.n3285 gnd.n3173 240.244
R13582 gnd.n3291 gnd.n3173 240.244
R13583 gnd.n3291 gnd.n3166 240.244
R13584 gnd.n3301 gnd.n3166 240.244
R13585 gnd.n3301 gnd.n3162 240.244
R13586 gnd.n3307 gnd.n3162 240.244
R13587 gnd.n3307 gnd.n3153 240.244
R13588 gnd.n3347 gnd.n3153 240.244
R13589 gnd.n3347 gnd.n3104 240.244
R13590 gnd.n3355 gnd.n3104 240.244
R13591 gnd.n3355 gnd.n3105 240.244
R13592 gnd.n3105 gnd.n3083 240.244
R13593 gnd.n3376 gnd.n3083 240.244
R13594 gnd.n3376 gnd.n3075 240.244
R13595 gnd.n3387 gnd.n3075 240.244
R13596 gnd.n3387 gnd.n3076 240.244
R13597 gnd.n3076 gnd.n3057 240.244
R13598 gnd.n3407 gnd.n3057 240.244
R13599 gnd.n3407 gnd.n3047 240.244
R13600 gnd.n3417 gnd.n3047 240.244
R13601 gnd.n3417 gnd.n3028 240.244
R13602 gnd.n3438 gnd.n3028 240.244
R13603 gnd.n3438 gnd.n3030 240.244
R13604 gnd.n3030 gnd.n3011 240.244
R13605 gnd.n3466 gnd.n3011 240.244
R13606 gnd.n3466 gnd.n2953 240.244
R13607 gnd.n3518 gnd.n2953 240.244
R13608 gnd.n3518 gnd.n2954 240.244
R13609 gnd.n3514 gnd.n2954 240.244
R13610 gnd.n3514 gnd.n2960 240.244
R13611 gnd.n2975 gnd.n2960 240.244
R13612 gnd.n3504 gnd.n2975 240.244
R13613 gnd.n3504 gnd.n2976 240.244
R13614 gnd.n3500 gnd.n2976 240.244
R13615 gnd.n3500 gnd.n2982 240.244
R13616 gnd.n2982 gnd.n2865 240.244
R13617 gnd.n3557 gnd.n2865 240.244
R13618 gnd.n3557 gnd.n2858 240.244
R13619 gnd.n3568 gnd.n2858 240.244
R13620 gnd.n3568 gnd.n2851 240.244
R13621 gnd.n3583 gnd.n2851 240.244
R13622 gnd.n3583 gnd.n2852 240.244
R13623 gnd.n2852 gnd.n2830 240.244
R13624 gnd.n3605 gnd.n2830 240.244
R13625 gnd.n3605 gnd.n2831 240.244
R13626 gnd.n2831 gnd.n2810 240.244
R13627 gnd.n3642 gnd.n2810 240.244
R13628 gnd.n3642 gnd.n2803 240.244
R13629 gnd.n3653 gnd.n2803 240.244
R13630 gnd.n3653 gnd.n2796 240.244
R13631 gnd.n3668 gnd.n2796 240.244
R13632 gnd.n3668 gnd.n2797 240.244
R13633 gnd.n2797 gnd.n2774 240.244
R13634 gnd.n3690 gnd.n2774 240.244
R13635 gnd.n3690 gnd.n2776 240.244
R13636 gnd.n2776 gnd.n2756 240.244
R13637 gnd.n3731 gnd.n2756 240.244
R13638 gnd.n3731 gnd.n2749 240.244
R13639 gnd.n3743 gnd.n2749 240.244
R13640 gnd.n3743 gnd.n2742 240.244
R13641 gnd.n4012 gnd.n2742 240.244
R13642 gnd.n4012 gnd.n2743 240.244
R13643 gnd.n2743 gnd.n2724 240.244
R13644 gnd.n4035 gnd.n2724 240.244
R13645 gnd.n2399 gnd.n1064 240.244
R13646 gnd.n2410 gnd.n2401 240.244
R13647 gnd.n2413 gnd.n2412 240.244
R13648 gnd.n2422 gnd.n2421 240.244
R13649 gnd.n2433 gnd.n2424 240.244
R13650 gnd.n2436 gnd.n2435 240.244
R13651 gnd.n2445 gnd.n2444 240.244
R13652 gnd.n2457 gnd.n2447 240.244
R13653 gnd.n2463 gnd.n2459 240.244
R13654 gnd.n4281 gnd.n2638 240.244
R13655 gnd.n4278 gnd.n2638 240.244
R13656 gnd.n4278 gnd.n2629 240.244
R13657 gnd.n4275 gnd.n2629 240.244
R13658 gnd.n4275 gnd.n2619 240.244
R13659 gnd.n4272 gnd.n2619 240.244
R13660 gnd.n4272 gnd.n2610 240.244
R13661 gnd.n4269 gnd.n2610 240.244
R13662 gnd.n4269 gnd.n2602 240.244
R13663 gnd.n4266 gnd.n2602 240.244
R13664 gnd.n4266 gnd.n2593 240.244
R13665 gnd.n4263 gnd.n2593 240.244
R13666 gnd.n4263 gnd.n2582 240.244
R13667 gnd.n2582 gnd.n2571 240.244
R13668 gnd.n4526 gnd.n2571 240.244
R13669 gnd.n4526 gnd.n2567 240.244
R13670 gnd.n4544 gnd.n2567 240.244
R13671 gnd.n4544 gnd.n2557 240.244
R13672 gnd.n4540 gnd.n2557 240.244
R13673 gnd.n4540 gnd.n2549 240.244
R13674 gnd.n4537 gnd.n2549 240.244
R13675 gnd.n4537 gnd.n2535 240.244
R13676 gnd.n4586 gnd.n2535 240.244
R13677 gnd.n4587 gnd.n4586 240.244
R13678 gnd.n4587 gnd.n940 240.244
R13679 gnd.n4599 gnd.n940 240.244
R13680 gnd.n4599 gnd.n2522 240.244
R13681 gnd.n4592 gnd.n2522 240.244
R13682 gnd.n4592 gnd.n2505 240.244
R13683 gnd.n4650 gnd.n2505 240.244
R13684 gnd.n4650 gnd.n957 240.244
R13685 gnd.n4656 gnd.n957 240.244
R13686 gnd.n4656 gnd.n969 240.244
R13687 gnd.n4665 gnd.n969 240.244
R13688 gnd.n4665 gnd.n978 240.244
R13689 gnd.n4671 gnd.n978 240.244
R13690 gnd.n4671 gnd.n988 240.244
R13691 gnd.n4707 gnd.n988 240.244
R13692 gnd.n4707 gnd.n998 240.244
R13693 gnd.n2492 gnd.n998 240.244
R13694 gnd.n2492 gnd.n1008 240.244
R13695 gnd.n2493 gnd.n1008 240.244
R13696 gnd.n2493 gnd.n1018 240.244
R13697 gnd.n4692 gnd.n1018 240.244
R13698 gnd.n4692 gnd.n1028 240.244
R13699 gnd.n2475 gnd.n1028 240.244
R13700 gnd.n2475 gnd.n1038 240.244
R13701 gnd.n4763 gnd.n1038 240.244
R13702 gnd.n4763 gnd.n1048 240.244
R13703 gnd.n4770 gnd.n1048 240.244
R13704 gnd.n4770 gnd.n1059 240.244
R13705 gnd.n4779 gnd.n1059 240.244
R13706 gnd.n4779 gnd.n1067 240.244
R13707 gnd.n4318 gnd.n4317 240.244
R13708 gnd.n4314 gnd.n4313 240.244
R13709 gnd.n4310 gnd.n4309 240.244
R13710 gnd.n4306 gnd.n4305 240.244
R13711 gnd.n4302 gnd.n4301 240.244
R13712 gnd.n4298 gnd.n4297 240.244
R13713 gnd.n4294 gnd.n4293 240.244
R13714 gnd.n4290 gnd.n4289 240.244
R13715 gnd.n4245 gnd.n4164 240.244
R13716 gnd.n4450 gnd.n2639 240.244
R13717 gnd.n4450 gnd.n2640 240.244
R13718 gnd.n2640 gnd.n2630 240.244
R13719 gnd.n2630 gnd.n2621 240.244
R13720 gnd.n4470 gnd.n2621 240.244
R13721 gnd.n4470 gnd.n2622 240.244
R13722 gnd.n2622 gnd.n2611 240.244
R13723 gnd.n2611 gnd.n2603 240.244
R13724 gnd.n4490 gnd.n2603 240.244
R13725 gnd.n4490 gnd.n2604 240.244
R13726 gnd.n2604 gnd.n2594 240.244
R13727 gnd.n2594 gnd.n2584 240.244
R13728 gnd.n4514 gnd.n2584 240.244
R13729 gnd.n4514 gnd.n2585 240.244
R13730 gnd.n2585 gnd.n2573 240.244
R13731 gnd.n4509 gnd.n2573 240.244
R13732 gnd.n4509 gnd.n2559 240.244
R13733 gnd.n4555 gnd.n2559 240.244
R13734 gnd.n4555 gnd.n2560 240.244
R13735 gnd.n2560 gnd.n2550 240.244
R13736 gnd.n2550 gnd.n2542 240.244
R13737 gnd.n4580 gnd.n2542 240.244
R13738 gnd.n4580 gnd.n2537 240.244
R13739 gnd.n4576 gnd.n2537 240.244
R13740 gnd.n4576 gnd.n941 240.244
R13741 gnd.n2524 gnd.n941 240.244
R13742 gnd.n4612 gnd.n2524 240.244
R13743 gnd.n4612 gnd.n2525 240.244
R13744 gnd.n2525 gnd.n2518 240.244
R13745 gnd.n2518 gnd.n959 240.244
R13746 gnd.n6475 gnd.n959 240.244
R13747 gnd.n6475 gnd.n960 240.244
R13748 gnd.n6471 gnd.n960 240.244
R13749 gnd.n6471 gnd.n966 240.244
R13750 gnd.n6463 gnd.n966 240.244
R13751 gnd.n6463 gnd.n980 240.244
R13752 gnd.n6459 gnd.n980 240.244
R13753 gnd.n6459 gnd.n985 240.244
R13754 gnd.n6451 gnd.n985 240.244
R13755 gnd.n6451 gnd.n1000 240.244
R13756 gnd.n6447 gnd.n1000 240.244
R13757 gnd.n6447 gnd.n1005 240.244
R13758 gnd.n6439 gnd.n1005 240.244
R13759 gnd.n6439 gnd.n1020 240.244
R13760 gnd.n6435 gnd.n1020 240.244
R13761 gnd.n6435 gnd.n1025 240.244
R13762 gnd.n6427 gnd.n1025 240.244
R13763 gnd.n6427 gnd.n1040 240.244
R13764 gnd.n6423 gnd.n1040 240.244
R13765 gnd.n6423 gnd.n1045 240.244
R13766 gnd.n6415 gnd.n1045 240.244
R13767 gnd.n6415 gnd.n1060 240.244
R13768 gnd.n6411 gnd.n1060 240.244
R13769 gnd.n6659 gnd.n767 240.244
R13770 gnd.n6659 gnd.n765 240.244
R13771 gnd.n6663 gnd.n765 240.244
R13772 gnd.n6663 gnd.n761 240.244
R13773 gnd.n6669 gnd.n761 240.244
R13774 gnd.n6669 gnd.n759 240.244
R13775 gnd.n6673 gnd.n759 240.244
R13776 gnd.n6673 gnd.n755 240.244
R13777 gnd.n6679 gnd.n755 240.244
R13778 gnd.n6679 gnd.n753 240.244
R13779 gnd.n6683 gnd.n753 240.244
R13780 gnd.n6683 gnd.n749 240.244
R13781 gnd.n6689 gnd.n749 240.244
R13782 gnd.n6689 gnd.n747 240.244
R13783 gnd.n6693 gnd.n747 240.244
R13784 gnd.n6693 gnd.n743 240.244
R13785 gnd.n6699 gnd.n743 240.244
R13786 gnd.n6699 gnd.n741 240.244
R13787 gnd.n6703 gnd.n741 240.244
R13788 gnd.n6703 gnd.n737 240.244
R13789 gnd.n6709 gnd.n737 240.244
R13790 gnd.n6709 gnd.n735 240.244
R13791 gnd.n6713 gnd.n735 240.244
R13792 gnd.n6713 gnd.n731 240.244
R13793 gnd.n6719 gnd.n731 240.244
R13794 gnd.n6719 gnd.n729 240.244
R13795 gnd.n6723 gnd.n729 240.244
R13796 gnd.n6723 gnd.n725 240.244
R13797 gnd.n6729 gnd.n725 240.244
R13798 gnd.n6729 gnd.n723 240.244
R13799 gnd.n6733 gnd.n723 240.244
R13800 gnd.n6733 gnd.n719 240.244
R13801 gnd.n6739 gnd.n719 240.244
R13802 gnd.n6739 gnd.n717 240.244
R13803 gnd.n6743 gnd.n717 240.244
R13804 gnd.n6743 gnd.n713 240.244
R13805 gnd.n6749 gnd.n713 240.244
R13806 gnd.n6749 gnd.n711 240.244
R13807 gnd.n6753 gnd.n711 240.244
R13808 gnd.n6753 gnd.n707 240.244
R13809 gnd.n6759 gnd.n707 240.244
R13810 gnd.n6759 gnd.n705 240.244
R13811 gnd.n6763 gnd.n705 240.244
R13812 gnd.n6763 gnd.n701 240.244
R13813 gnd.n6769 gnd.n701 240.244
R13814 gnd.n6769 gnd.n699 240.244
R13815 gnd.n6773 gnd.n699 240.244
R13816 gnd.n6773 gnd.n695 240.244
R13817 gnd.n6779 gnd.n695 240.244
R13818 gnd.n6779 gnd.n693 240.244
R13819 gnd.n6783 gnd.n693 240.244
R13820 gnd.n6783 gnd.n689 240.244
R13821 gnd.n6789 gnd.n689 240.244
R13822 gnd.n6789 gnd.n687 240.244
R13823 gnd.n6793 gnd.n687 240.244
R13824 gnd.n6793 gnd.n683 240.244
R13825 gnd.n6799 gnd.n683 240.244
R13826 gnd.n6799 gnd.n681 240.244
R13827 gnd.n6803 gnd.n681 240.244
R13828 gnd.n6803 gnd.n677 240.244
R13829 gnd.n6809 gnd.n677 240.244
R13830 gnd.n6809 gnd.n675 240.244
R13831 gnd.n6813 gnd.n675 240.244
R13832 gnd.n6813 gnd.n671 240.244
R13833 gnd.n6819 gnd.n671 240.244
R13834 gnd.n6819 gnd.n669 240.244
R13835 gnd.n6823 gnd.n669 240.244
R13836 gnd.n6823 gnd.n665 240.244
R13837 gnd.n6829 gnd.n665 240.244
R13838 gnd.n6829 gnd.n663 240.244
R13839 gnd.n6833 gnd.n663 240.244
R13840 gnd.n6833 gnd.n659 240.244
R13841 gnd.n6839 gnd.n659 240.244
R13842 gnd.n6839 gnd.n657 240.244
R13843 gnd.n6843 gnd.n657 240.244
R13844 gnd.n6843 gnd.n653 240.244
R13845 gnd.n6849 gnd.n653 240.244
R13846 gnd.n6849 gnd.n651 240.244
R13847 gnd.n6853 gnd.n651 240.244
R13848 gnd.n6853 gnd.n647 240.244
R13849 gnd.n6859 gnd.n647 240.244
R13850 gnd.n6859 gnd.n645 240.244
R13851 gnd.n6863 gnd.n645 240.244
R13852 gnd.n6863 gnd.n641 240.244
R13853 gnd.n6869 gnd.n641 240.244
R13854 gnd.n6869 gnd.n639 240.244
R13855 gnd.n6873 gnd.n639 240.244
R13856 gnd.n6873 gnd.n635 240.244
R13857 gnd.n6879 gnd.n635 240.244
R13858 gnd.n6879 gnd.n633 240.244
R13859 gnd.n6883 gnd.n633 240.244
R13860 gnd.n6883 gnd.n629 240.244
R13861 gnd.n6889 gnd.n629 240.244
R13862 gnd.n6889 gnd.n627 240.244
R13863 gnd.n6893 gnd.n627 240.244
R13864 gnd.n6893 gnd.n623 240.244
R13865 gnd.n6899 gnd.n623 240.244
R13866 gnd.n6899 gnd.n621 240.244
R13867 gnd.n6903 gnd.n621 240.244
R13868 gnd.n6903 gnd.n617 240.244
R13869 gnd.n6909 gnd.n617 240.244
R13870 gnd.n6909 gnd.n615 240.244
R13871 gnd.n6913 gnd.n615 240.244
R13872 gnd.n6913 gnd.n611 240.244
R13873 gnd.n6919 gnd.n611 240.244
R13874 gnd.n6919 gnd.n609 240.244
R13875 gnd.n6923 gnd.n609 240.244
R13876 gnd.n6923 gnd.n605 240.244
R13877 gnd.n6929 gnd.n605 240.244
R13878 gnd.n6929 gnd.n603 240.244
R13879 gnd.n6933 gnd.n603 240.244
R13880 gnd.n6933 gnd.n599 240.244
R13881 gnd.n6939 gnd.n599 240.244
R13882 gnd.n6939 gnd.n597 240.244
R13883 gnd.n6943 gnd.n597 240.244
R13884 gnd.n6943 gnd.n593 240.244
R13885 gnd.n6949 gnd.n593 240.244
R13886 gnd.n6949 gnd.n591 240.244
R13887 gnd.n6953 gnd.n591 240.244
R13888 gnd.n6953 gnd.n587 240.244
R13889 gnd.n6959 gnd.n587 240.244
R13890 gnd.n6959 gnd.n585 240.244
R13891 gnd.n6963 gnd.n585 240.244
R13892 gnd.n6963 gnd.n581 240.244
R13893 gnd.n6969 gnd.n581 240.244
R13894 gnd.n6969 gnd.n579 240.244
R13895 gnd.n6973 gnd.n579 240.244
R13896 gnd.n6973 gnd.n575 240.244
R13897 gnd.n6979 gnd.n575 240.244
R13898 gnd.n6979 gnd.n573 240.244
R13899 gnd.n6983 gnd.n573 240.244
R13900 gnd.n6983 gnd.n569 240.244
R13901 gnd.n6989 gnd.n569 240.244
R13902 gnd.n6989 gnd.n567 240.244
R13903 gnd.n6993 gnd.n567 240.244
R13904 gnd.n6993 gnd.n563 240.244
R13905 gnd.n6999 gnd.n563 240.244
R13906 gnd.n6999 gnd.n561 240.244
R13907 gnd.n7003 gnd.n561 240.244
R13908 gnd.n7003 gnd.n557 240.244
R13909 gnd.n7009 gnd.n557 240.244
R13910 gnd.n7009 gnd.n555 240.244
R13911 gnd.n7013 gnd.n555 240.244
R13912 gnd.n7013 gnd.n551 240.244
R13913 gnd.n7019 gnd.n551 240.244
R13914 gnd.n7019 gnd.n549 240.244
R13915 gnd.n7023 gnd.n549 240.244
R13916 gnd.n7023 gnd.n545 240.244
R13917 gnd.n7029 gnd.n545 240.244
R13918 gnd.n7029 gnd.n543 240.244
R13919 gnd.n7033 gnd.n543 240.244
R13920 gnd.n7033 gnd.n539 240.244
R13921 gnd.n7039 gnd.n539 240.244
R13922 gnd.n7039 gnd.n537 240.244
R13923 gnd.n7043 gnd.n537 240.244
R13924 gnd.n7043 gnd.n533 240.244
R13925 gnd.n7049 gnd.n533 240.244
R13926 gnd.n7049 gnd.n531 240.244
R13927 gnd.n7053 gnd.n531 240.244
R13928 gnd.n7053 gnd.n527 240.244
R13929 gnd.n7059 gnd.n527 240.244
R13930 gnd.n7059 gnd.n525 240.244
R13931 gnd.n7063 gnd.n525 240.244
R13932 gnd.n7063 gnd.n521 240.244
R13933 gnd.n7069 gnd.n521 240.244
R13934 gnd.n7069 gnd.n519 240.244
R13935 gnd.n7073 gnd.n519 240.244
R13936 gnd.n7079 gnd.n515 240.244
R13937 gnd.n7079 gnd.n513 240.244
R13938 gnd.n7083 gnd.n513 240.244
R13939 gnd.n7083 gnd.n509 240.244
R13940 gnd.n7089 gnd.n509 240.244
R13941 gnd.n7089 gnd.n507 240.244
R13942 gnd.n7093 gnd.n507 240.244
R13943 gnd.n7093 gnd.n503 240.244
R13944 gnd.n7099 gnd.n503 240.244
R13945 gnd.n7099 gnd.n501 240.244
R13946 gnd.n7103 gnd.n501 240.244
R13947 gnd.n7103 gnd.n497 240.244
R13948 gnd.n7109 gnd.n497 240.244
R13949 gnd.n7109 gnd.n495 240.244
R13950 gnd.n7113 gnd.n495 240.244
R13951 gnd.n7113 gnd.n491 240.244
R13952 gnd.n7119 gnd.n491 240.244
R13953 gnd.n7119 gnd.n489 240.244
R13954 gnd.n7123 gnd.n489 240.244
R13955 gnd.n7123 gnd.n485 240.244
R13956 gnd.n7129 gnd.n485 240.244
R13957 gnd.n7129 gnd.n483 240.244
R13958 gnd.n7133 gnd.n483 240.244
R13959 gnd.n7133 gnd.n479 240.244
R13960 gnd.n7139 gnd.n479 240.244
R13961 gnd.n7139 gnd.n477 240.244
R13962 gnd.n7143 gnd.n477 240.244
R13963 gnd.n7143 gnd.n473 240.244
R13964 gnd.n7149 gnd.n473 240.244
R13965 gnd.n7149 gnd.n471 240.244
R13966 gnd.n7153 gnd.n471 240.244
R13967 gnd.n7153 gnd.n467 240.244
R13968 gnd.n7159 gnd.n467 240.244
R13969 gnd.n7159 gnd.n465 240.244
R13970 gnd.n7163 gnd.n465 240.244
R13971 gnd.n7163 gnd.n461 240.244
R13972 gnd.n7169 gnd.n461 240.244
R13973 gnd.n7169 gnd.n459 240.244
R13974 gnd.n7173 gnd.n459 240.244
R13975 gnd.n7173 gnd.n455 240.244
R13976 gnd.n7179 gnd.n455 240.244
R13977 gnd.n7179 gnd.n453 240.244
R13978 gnd.n7183 gnd.n453 240.244
R13979 gnd.n7183 gnd.n449 240.244
R13980 gnd.n7189 gnd.n449 240.244
R13981 gnd.n7189 gnd.n447 240.244
R13982 gnd.n7193 gnd.n447 240.244
R13983 gnd.n7193 gnd.n443 240.244
R13984 gnd.n7199 gnd.n443 240.244
R13985 gnd.n7199 gnd.n441 240.244
R13986 gnd.n7203 gnd.n441 240.244
R13987 gnd.n7203 gnd.n437 240.244
R13988 gnd.n7209 gnd.n437 240.244
R13989 gnd.n7209 gnd.n435 240.244
R13990 gnd.n7213 gnd.n435 240.244
R13991 gnd.n7213 gnd.n431 240.244
R13992 gnd.n7219 gnd.n431 240.244
R13993 gnd.n7219 gnd.n429 240.244
R13994 gnd.n7223 gnd.n429 240.244
R13995 gnd.n7223 gnd.n425 240.244
R13996 gnd.n7229 gnd.n425 240.244
R13997 gnd.n7229 gnd.n423 240.244
R13998 gnd.n7233 gnd.n423 240.244
R13999 gnd.n7233 gnd.n419 240.244
R14000 gnd.n7239 gnd.n419 240.244
R14001 gnd.n7239 gnd.n417 240.244
R14002 gnd.n7243 gnd.n417 240.244
R14003 gnd.n7243 gnd.n413 240.244
R14004 gnd.n7249 gnd.n413 240.244
R14005 gnd.n7249 gnd.n411 240.244
R14006 gnd.n7253 gnd.n411 240.244
R14007 gnd.n7253 gnd.n407 240.244
R14008 gnd.n7259 gnd.n407 240.244
R14009 gnd.n7259 gnd.n405 240.244
R14010 gnd.n7263 gnd.n405 240.244
R14011 gnd.n7263 gnd.n401 240.244
R14012 gnd.n7269 gnd.n401 240.244
R14013 gnd.n7269 gnd.n399 240.244
R14014 gnd.n7273 gnd.n399 240.244
R14015 gnd.n7273 gnd.n395 240.244
R14016 gnd.n7281 gnd.n395 240.244
R14017 gnd.n7281 gnd.n393 240.244
R14018 gnd.n7285 gnd.n393 240.244
R14019 gnd.n7286 gnd.n7285 240.244
R14020 gnd.n2515 gnd.n937 240.244
R14021 gnd.n4621 gnd.n2515 240.244
R14022 gnd.n4621 gnd.n2508 240.244
R14023 gnd.n4647 gnd.n2508 240.244
R14024 gnd.n4647 gnd.n2509 240.244
R14025 gnd.n4643 gnd.n2509 240.244
R14026 gnd.n4643 gnd.n4642 240.244
R14027 gnd.n4642 gnd.n4641 240.244
R14028 gnd.n4641 gnd.n4629 240.244
R14029 gnd.n4637 gnd.n4629 240.244
R14030 gnd.n4637 gnd.n2485 240.244
R14031 gnd.n4710 gnd.n2485 240.244
R14032 gnd.n4711 gnd.n4710 240.244
R14033 gnd.n4712 gnd.n4711 240.244
R14034 gnd.n4712 gnd.n2481 240.244
R14035 gnd.n4718 gnd.n2481 240.244
R14036 gnd.n4719 gnd.n4718 240.244
R14037 gnd.n4720 gnd.n4719 240.244
R14038 gnd.n4720 gnd.n2476 240.244
R14039 gnd.n4754 gnd.n2476 240.244
R14040 gnd.n4754 gnd.n2477 240.244
R14041 gnd.n4750 gnd.n2477 240.244
R14042 gnd.n4750 gnd.n4749 240.244
R14043 gnd.n4749 gnd.n4748 240.244
R14044 gnd.n4748 gnd.n4728 240.244
R14045 gnd.n4744 gnd.n4728 240.244
R14046 gnd.n4744 gnd.n4743 240.244
R14047 gnd.n4743 gnd.n4742 240.244
R14048 gnd.n4742 gnd.n4735 240.244
R14049 gnd.n4735 gnd.n2202 240.244
R14050 gnd.n4859 gnd.n2202 240.244
R14051 gnd.n4859 gnd.n2198 240.244
R14052 gnd.n4865 gnd.n2198 240.244
R14053 gnd.n4865 gnd.n2189 240.244
R14054 gnd.n4875 gnd.n2189 240.244
R14055 gnd.n4875 gnd.n2185 240.244
R14056 gnd.n4881 gnd.n2185 240.244
R14057 gnd.n4881 gnd.n2175 240.244
R14058 gnd.n4891 gnd.n2175 240.244
R14059 gnd.n4891 gnd.n2171 240.244
R14060 gnd.n4897 gnd.n2171 240.244
R14061 gnd.n4897 gnd.n2160 240.244
R14062 gnd.n4907 gnd.n2160 240.244
R14063 gnd.n4907 gnd.n2156 240.244
R14064 gnd.n4913 gnd.n2156 240.244
R14065 gnd.n4913 gnd.n2146 240.244
R14066 gnd.n4923 gnd.n2146 240.244
R14067 gnd.n4923 gnd.n2142 240.244
R14068 gnd.n4929 gnd.n2142 240.244
R14069 gnd.n4929 gnd.n2131 240.244
R14070 gnd.n4965 gnd.n2131 240.244
R14071 gnd.n4965 gnd.n2126 240.244
R14072 gnd.n4974 gnd.n2126 240.244
R14073 gnd.n4974 gnd.n2127 240.244
R14074 gnd.n2127 gnd.n1188 240.244
R14075 gnd.n6283 gnd.n1188 240.244
R14076 gnd.n6283 gnd.n1189 240.244
R14077 gnd.n6279 gnd.n1189 240.244
R14078 gnd.n6279 gnd.n1195 240.244
R14079 gnd.n1291 gnd.n1195 240.244
R14080 gnd.n6264 gnd.n1291 240.244
R14081 gnd.n6264 gnd.n1292 240.244
R14082 gnd.n6260 gnd.n1292 240.244
R14083 gnd.n6260 gnd.n1300 240.244
R14084 gnd.n5037 gnd.n1300 240.244
R14085 gnd.n5037 gnd.n2099 240.244
R14086 gnd.n5043 gnd.n2099 240.244
R14087 gnd.n5043 gnd.n2077 240.244
R14088 gnd.n5096 gnd.n2077 240.244
R14089 gnd.n5096 gnd.n2072 240.244
R14090 gnd.n5104 gnd.n2072 240.244
R14091 gnd.n5104 gnd.n2073 240.244
R14092 gnd.n2073 gnd.n2054 240.244
R14093 gnd.n5128 gnd.n2054 240.244
R14094 gnd.n5128 gnd.n2049 240.244
R14095 gnd.n5136 gnd.n2049 240.244
R14096 gnd.n5136 gnd.n2050 240.244
R14097 gnd.n2050 gnd.n2032 240.244
R14098 gnd.n5178 gnd.n2032 240.244
R14099 gnd.n5178 gnd.n2027 240.244
R14100 gnd.n5186 gnd.n2027 240.244
R14101 gnd.n5186 gnd.n2028 240.244
R14102 gnd.n2028 gnd.n2004 240.244
R14103 gnd.n5216 gnd.n2004 240.244
R14104 gnd.n5216 gnd.n2000 240.244
R14105 gnd.n5222 gnd.n2000 240.244
R14106 gnd.n5222 gnd.n1976 240.244
R14107 gnd.n5253 gnd.n1976 240.244
R14108 gnd.n5253 gnd.n1971 240.244
R14109 gnd.n5261 gnd.n1971 240.244
R14110 gnd.n5261 gnd.n1972 240.244
R14111 gnd.n1972 gnd.n1957 240.244
R14112 gnd.n5311 gnd.n1957 240.244
R14113 gnd.n5311 gnd.n1952 240.244
R14114 gnd.n5319 gnd.n1952 240.244
R14115 gnd.n5319 gnd.n1953 240.244
R14116 gnd.n1953 gnd.n1934 240.244
R14117 gnd.n5349 gnd.n1934 240.244
R14118 gnd.n5349 gnd.n1929 240.244
R14119 gnd.n5357 gnd.n1929 240.244
R14120 gnd.n5357 gnd.n1930 240.244
R14121 gnd.n1930 gnd.n1906 240.244
R14122 gnd.n5405 gnd.n1906 240.244
R14123 gnd.n5405 gnd.n1901 240.244
R14124 gnd.n5413 gnd.n1901 240.244
R14125 gnd.n5413 gnd.n1902 240.244
R14126 gnd.n1902 gnd.n1885 240.244
R14127 gnd.n5443 gnd.n1885 240.244
R14128 gnd.n5443 gnd.n1881 240.244
R14129 gnd.n5449 gnd.n1881 240.244
R14130 gnd.n5449 gnd.n1829 240.244
R14131 gnd.n5618 gnd.n1829 240.244
R14132 gnd.n5618 gnd.n1825 240.244
R14133 gnd.n5624 gnd.n1825 240.244
R14134 gnd.n5624 gnd.n1818 240.244
R14135 gnd.n5635 gnd.n1818 240.244
R14136 gnd.n5635 gnd.n1814 240.244
R14137 gnd.n5641 gnd.n1814 240.244
R14138 gnd.n5641 gnd.n1806 240.244
R14139 gnd.n5652 gnd.n1806 240.244
R14140 gnd.n5652 gnd.n1802 240.244
R14141 gnd.n5658 gnd.n1802 240.244
R14142 gnd.n5658 gnd.n1794 240.244
R14143 gnd.n5669 gnd.n1794 240.244
R14144 gnd.n5669 gnd.n1790 240.244
R14145 gnd.n5675 gnd.n1790 240.244
R14146 gnd.n5675 gnd.n1782 240.244
R14147 gnd.n5686 gnd.n1782 240.244
R14148 gnd.n5686 gnd.n1778 240.244
R14149 gnd.n5695 gnd.n1778 240.244
R14150 gnd.n5695 gnd.n1770 240.244
R14151 gnd.n5706 gnd.n1770 240.244
R14152 gnd.n5707 gnd.n5706 240.244
R14153 gnd.n5707 gnd.n1397 240.244
R14154 gnd.n1765 gnd.n1397 240.244
R14155 gnd.n5725 gnd.n1765 240.244
R14156 gnd.n5725 gnd.n1766 240.244
R14157 gnd.n5721 gnd.n1766 240.244
R14158 gnd.n5721 gnd.n5720 240.244
R14159 gnd.n5720 gnd.n5719 240.244
R14160 gnd.n5719 gnd.n1734 240.244
R14161 gnd.n5777 gnd.n1734 240.244
R14162 gnd.n5777 gnd.n1730 240.244
R14163 gnd.n5783 gnd.n1730 240.244
R14164 gnd.n5784 gnd.n5783 240.244
R14165 gnd.n5785 gnd.n5784 240.244
R14166 gnd.n5785 gnd.n1726 240.244
R14167 gnd.n5791 gnd.n1726 240.244
R14168 gnd.n5792 gnd.n5791 240.244
R14169 gnd.n5793 gnd.n5792 240.244
R14170 gnd.n5793 gnd.n1721 240.244
R14171 gnd.n5819 gnd.n1721 240.244
R14172 gnd.n5819 gnd.n1722 240.244
R14173 gnd.n5815 gnd.n1722 240.244
R14174 gnd.n5815 gnd.n5814 240.244
R14175 gnd.n5814 gnd.n5813 240.244
R14176 gnd.n5813 gnd.n5801 240.244
R14177 gnd.n5809 gnd.n5801 240.244
R14178 gnd.n5809 gnd.n1704 240.244
R14179 gnd.n5876 gnd.n1704 240.244
R14180 gnd.n5877 gnd.n5876 240.244
R14181 gnd.n5878 gnd.n5877 240.244
R14182 gnd.n5878 gnd.n1700 240.244
R14183 gnd.n5885 gnd.n1700 240.244
R14184 gnd.n5885 gnd.n387 240.244
R14185 gnd.n7292 gnd.n387 240.244
R14186 gnd.n7292 gnd.n388 240.244
R14187 gnd.n6653 gnd.n771 240.244
R14188 gnd.n6649 gnd.n771 240.244
R14189 gnd.n6649 gnd.n773 240.244
R14190 gnd.n6645 gnd.n773 240.244
R14191 gnd.n6645 gnd.n778 240.244
R14192 gnd.n6641 gnd.n778 240.244
R14193 gnd.n6641 gnd.n780 240.244
R14194 gnd.n6637 gnd.n780 240.244
R14195 gnd.n6637 gnd.n786 240.244
R14196 gnd.n6633 gnd.n786 240.244
R14197 gnd.n6633 gnd.n788 240.244
R14198 gnd.n6629 gnd.n788 240.244
R14199 gnd.n6629 gnd.n794 240.244
R14200 gnd.n6625 gnd.n794 240.244
R14201 gnd.n6625 gnd.n796 240.244
R14202 gnd.n6621 gnd.n796 240.244
R14203 gnd.n6621 gnd.n802 240.244
R14204 gnd.n6617 gnd.n802 240.244
R14205 gnd.n6617 gnd.n804 240.244
R14206 gnd.n6613 gnd.n804 240.244
R14207 gnd.n6613 gnd.n810 240.244
R14208 gnd.n6609 gnd.n810 240.244
R14209 gnd.n6609 gnd.n812 240.244
R14210 gnd.n6605 gnd.n812 240.244
R14211 gnd.n6605 gnd.n818 240.244
R14212 gnd.n6601 gnd.n818 240.244
R14213 gnd.n6601 gnd.n820 240.244
R14214 gnd.n6597 gnd.n820 240.244
R14215 gnd.n6597 gnd.n826 240.244
R14216 gnd.n6593 gnd.n826 240.244
R14217 gnd.n6593 gnd.n828 240.244
R14218 gnd.n6589 gnd.n828 240.244
R14219 gnd.n6589 gnd.n834 240.244
R14220 gnd.n6585 gnd.n834 240.244
R14221 gnd.n6585 gnd.n836 240.244
R14222 gnd.n6581 gnd.n836 240.244
R14223 gnd.n6581 gnd.n842 240.244
R14224 gnd.n6577 gnd.n842 240.244
R14225 gnd.n6577 gnd.n844 240.244
R14226 gnd.n6573 gnd.n844 240.244
R14227 gnd.n6573 gnd.n850 240.244
R14228 gnd.n6569 gnd.n850 240.244
R14229 gnd.n6569 gnd.n852 240.244
R14230 gnd.n6565 gnd.n852 240.244
R14231 gnd.n6565 gnd.n858 240.244
R14232 gnd.n6561 gnd.n858 240.244
R14233 gnd.n6561 gnd.n860 240.244
R14234 gnd.n6557 gnd.n860 240.244
R14235 gnd.n6557 gnd.n866 240.244
R14236 gnd.n6553 gnd.n866 240.244
R14237 gnd.n6553 gnd.n868 240.244
R14238 gnd.n6549 gnd.n868 240.244
R14239 gnd.n6549 gnd.n874 240.244
R14240 gnd.n6545 gnd.n874 240.244
R14241 gnd.n6545 gnd.n876 240.244
R14242 gnd.n6541 gnd.n876 240.244
R14243 gnd.n6541 gnd.n882 240.244
R14244 gnd.n6537 gnd.n882 240.244
R14245 gnd.n6537 gnd.n884 240.244
R14246 gnd.n6533 gnd.n884 240.244
R14247 gnd.n6533 gnd.n890 240.244
R14248 gnd.n6529 gnd.n890 240.244
R14249 gnd.n6529 gnd.n892 240.244
R14250 gnd.n6525 gnd.n892 240.244
R14251 gnd.n6525 gnd.n898 240.244
R14252 gnd.n6521 gnd.n898 240.244
R14253 gnd.n6521 gnd.n900 240.244
R14254 gnd.n6517 gnd.n900 240.244
R14255 gnd.n6517 gnd.n906 240.244
R14256 gnd.n6513 gnd.n906 240.244
R14257 gnd.n6513 gnd.n908 240.244
R14258 gnd.n6509 gnd.n908 240.244
R14259 gnd.n6509 gnd.n914 240.244
R14260 gnd.n6505 gnd.n914 240.244
R14261 gnd.n6505 gnd.n916 240.244
R14262 gnd.n6501 gnd.n916 240.244
R14263 gnd.n6501 gnd.n922 240.244
R14264 gnd.n6497 gnd.n922 240.244
R14265 gnd.n6497 gnd.n924 240.244
R14266 gnd.n6493 gnd.n924 240.244
R14267 gnd.n6493 gnd.n930 240.244
R14268 gnd.n6489 gnd.n930 240.244
R14269 gnd.n6489 gnd.n932 240.244
R14270 gnd.n6485 gnd.n932 240.244
R14271 gnd.n2220 gnd.n2196 240.244
R14272 gnd.n2220 gnd.n2190 240.244
R14273 gnd.n2221 gnd.n2190 240.244
R14274 gnd.n2221 gnd.n2184 240.244
R14275 gnd.n2224 gnd.n2184 240.244
R14276 gnd.n2224 gnd.n2177 240.244
R14277 gnd.n2225 gnd.n2177 240.244
R14278 gnd.n2225 gnd.n2170 240.244
R14279 gnd.n2228 gnd.n2170 240.244
R14280 gnd.n2228 gnd.n2162 240.244
R14281 gnd.n2229 gnd.n2162 240.244
R14282 gnd.n2229 gnd.n2155 240.244
R14283 gnd.n2232 gnd.n2155 240.244
R14284 gnd.n2232 gnd.n2148 240.244
R14285 gnd.n2233 gnd.n2148 240.244
R14286 gnd.n2233 gnd.n2141 240.244
R14287 gnd.n2236 gnd.n2141 240.244
R14288 gnd.n2236 gnd.n2133 240.244
R14289 gnd.n2133 gnd.n2122 240.244
R14290 gnd.n4976 gnd.n2122 240.244
R14291 gnd.n4977 gnd.n4976 240.244
R14292 gnd.n4978 gnd.n4977 240.244
R14293 gnd.n4978 gnd.n1185 240.244
R14294 gnd.n4940 gnd.n1185 240.244
R14295 gnd.n4940 gnd.n1198 240.244
R14296 gnd.n4986 gnd.n1198 240.244
R14297 gnd.n4987 gnd.n4986 240.244
R14298 gnd.n4987 gnd.n1288 240.244
R14299 gnd.n5009 gnd.n1288 240.244
R14300 gnd.n5009 gnd.n1301 240.244
R14301 gnd.n4992 gnd.n1301 240.244
R14302 gnd.n4992 gnd.n2102 240.244
R14303 gnd.n4993 gnd.n2102 240.244
R14304 gnd.n4993 gnd.n2097 240.244
R14305 gnd.n4996 gnd.n2097 240.244
R14306 gnd.n4996 gnd.n2079 240.244
R14307 gnd.n2079 gnd.n2070 240.244
R14308 gnd.n5106 gnd.n2070 240.244
R14309 gnd.n5106 gnd.n2065 240.244
R14310 gnd.n5113 gnd.n2065 240.244
R14311 gnd.n5113 gnd.n2056 240.244
R14312 gnd.n2056 gnd.n2045 240.244
R14313 gnd.n5138 gnd.n2045 240.244
R14314 gnd.n5138 gnd.n2040 240.244
R14315 gnd.n5168 gnd.n2040 240.244
R14316 gnd.n5168 gnd.n2034 240.244
R14317 gnd.n5143 gnd.n2034 240.244
R14318 gnd.n5143 gnd.n2025 240.244
R14319 gnd.n5144 gnd.n2025 240.244
R14320 gnd.n5145 gnd.n5144 240.244
R14321 gnd.n5145 gnd.n2006 240.244
R14322 gnd.n5148 gnd.n2006 240.244
R14323 gnd.n5148 gnd.n1998 240.244
R14324 gnd.n5149 gnd.n1998 240.244
R14325 gnd.n5149 gnd.n1978 240.244
R14326 gnd.n1978 gnd.n1969 240.244
R14327 gnd.n5263 gnd.n1969 240.244
R14328 gnd.n5263 gnd.n1964 240.244
R14329 gnd.n5299 gnd.n1964 240.244
R14330 gnd.n5299 gnd.n1959 240.244
R14331 gnd.n5268 gnd.n1959 240.244
R14332 gnd.n5268 gnd.n1951 240.244
R14333 gnd.n5271 gnd.n1951 240.244
R14334 gnd.n5271 gnd.n1943 240.244
R14335 gnd.n1943 gnd.n1935 240.244
R14336 gnd.n5274 gnd.n1935 240.244
R14337 gnd.n5274 gnd.n1927 240.244
R14338 gnd.n5277 gnd.n1927 240.244
R14339 gnd.n5280 gnd.n5277 240.244
R14340 gnd.n5280 gnd.n1908 240.244
R14341 gnd.n1908 gnd.n1898 240.244
R14342 gnd.n5415 gnd.n1898 240.244
R14343 gnd.n5415 gnd.n1893 240.244
R14344 gnd.n5432 gnd.n1893 240.244
R14345 gnd.n5432 gnd.n1887 240.244
R14346 gnd.n5420 gnd.n1887 240.244
R14347 gnd.n5420 gnd.n1879 240.244
R14348 gnd.n5421 gnd.n1879 240.244
R14349 gnd.n5421 gnd.n1831 240.244
R14350 gnd.n1831 gnd.n1824 240.244
R14351 gnd.n5626 gnd.n1824 240.244
R14352 gnd.n5626 gnd.n1820 240.244
R14353 gnd.n5632 gnd.n1820 240.244
R14354 gnd.n5632 gnd.n1812 240.244
R14355 gnd.n5643 gnd.n1812 240.244
R14356 gnd.n5643 gnd.n1808 240.244
R14357 gnd.n5649 gnd.n1808 240.244
R14358 gnd.n5649 gnd.n1800 240.244
R14359 gnd.n5660 gnd.n1800 240.244
R14360 gnd.n5660 gnd.n1796 240.244
R14361 gnd.n5666 gnd.n1796 240.244
R14362 gnd.n5666 gnd.n1787 240.244
R14363 gnd.n5677 gnd.n1787 240.244
R14364 gnd.n5677 gnd.n1783 240.244
R14365 gnd.n5683 gnd.n1783 240.244
R14366 gnd.n5683 gnd.n1776 240.244
R14367 gnd.n5697 gnd.n1776 240.244
R14368 gnd.n5697 gnd.n1772 240.244
R14369 gnd.n5703 gnd.n1772 240.244
R14370 gnd.n5703 gnd.n1399 240.244
R14371 gnd.n6147 gnd.n1399 240.244
R14372 gnd.n2218 gnd.n2217 240.244
R14373 gnd.n2273 gnd.n2217 240.244
R14374 gnd.n2275 gnd.n2274 240.244
R14375 gnd.n2392 gnd.n2391 240.244
R14376 gnd.n2394 gnd.n2393 240.244
R14377 gnd.n2405 gnd.n2404 240.244
R14378 gnd.n2407 gnd.n2406 240.244
R14379 gnd.n2417 gnd.n2416 240.244
R14380 gnd.n2428 gnd.n2427 240.244
R14381 gnd.n2430 gnd.n2429 240.244
R14382 gnd.n2440 gnd.n2439 240.244
R14383 gnd.n2451 gnd.n2450 240.244
R14384 gnd.n4784 gnd.n2452 240.244
R14385 gnd.n4788 gnd.n4787 240.244
R14386 gnd.n4867 gnd.n2191 240.244
R14387 gnd.n4873 gnd.n2191 240.244
R14388 gnd.n4873 gnd.n2182 240.244
R14389 gnd.n4883 gnd.n2182 240.244
R14390 gnd.n4883 gnd.n2178 240.244
R14391 gnd.n4889 gnd.n2178 240.244
R14392 gnd.n4889 gnd.n2168 240.244
R14393 gnd.n4899 gnd.n2168 240.244
R14394 gnd.n4899 gnd.n2164 240.244
R14395 gnd.n4905 gnd.n2164 240.244
R14396 gnd.n4905 gnd.n2154 240.244
R14397 gnd.n4915 gnd.n2154 240.244
R14398 gnd.n4915 gnd.n2150 240.244
R14399 gnd.n4921 gnd.n2150 240.244
R14400 gnd.n4921 gnd.n2140 240.244
R14401 gnd.n4931 gnd.n2140 240.244
R14402 gnd.n4931 gnd.n2134 240.244
R14403 gnd.n4963 gnd.n2134 240.244
R14404 gnd.n4963 gnd.n2135 240.244
R14405 gnd.n2135 gnd.n2125 240.244
R14406 gnd.n4936 gnd.n2125 240.244
R14407 gnd.n4937 gnd.n4936 240.244
R14408 gnd.n4937 gnd.n1187 240.244
R14409 gnd.n4942 gnd.n1187 240.244
R14410 gnd.n4942 gnd.n1199 240.244
R14411 gnd.n4943 gnd.n1199 240.244
R14412 gnd.n4944 gnd.n4943 240.244
R14413 gnd.n4944 gnd.n1290 240.244
R14414 gnd.n1303 gnd.n1290 240.244
R14415 gnd.n6258 gnd.n1303 240.244
R14416 gnd.n6258 gnd.n1304 240.244
R14417 gnd.n1309 gnd.n1304 240.244
R14418 gnd.n1310 gnd.n1309 240.244
R14419 gnd.n1311 gnd.n1310 240.244
R14420 gnd.n2090 gnd.n1311 240.244
R14421 gnd.n2090 gnd.n1314 240.244
R14422 gnd.n1315 gnd.n1314 240.244
R14423 gnd.n1316 gnd.n1315 240.244
R14424 gnd.n5085 gnd.n1316 240.244
R14425 gnd.n5085 gnd.n1319 240.244
R14426 gnd.n1320 gnd.n1319 240.244
R14427 gnd.n1321 gnd.n1320 240.244
R14428 gnd.n2048 gnd.n1321 240.244
R14429 gnd.n2048 gnd.n1324 240.244
R14430 gnd.n1325 gnd.n1324 240.244
R14431 gnd.n1326 gnd.n1325 240.244
R14432 gnd.n2022 gnd.n1326 240.244
R14433 gnd.n2022 gnd.n1329 240.244
R14434 gnd.n1330 gnd.n1329 240.244
R14435 gnd.n1331 gnd.n1330 240.244
R14436 gnd.n5214 gnd.n1331 240.244
R14437 gnd.n5214 gnd.n1334 240.244
R14438 gnd.n1335 gnd.n1334 240.244
R14439 gnd.n1336 gnd.n1335 240.244
R14440 gnd.n5251 gnd.n1336 240.244
R14441 gnd.n5251 gnd.n1339 240.244
R14442 gnd.n1340 gnd.n1339 240.244
R14443 gnd.n1341 gnd.n1340 240.244
R14444 gnd.n5300 gnd.n1341 240.244
R14445 gnd.n5300 gnd.n1344 240.244
R14446 gnd.n1345 gnd.n1344 240.244
R14447 gnd.n1346 gnd.n1345 240.244
R14448 gnd.n5269 gnd.n1346 240.244
R14449 gnd.n5269 gnd.n1349 240.244
R14450 gnd.n1350 gnd.n1349 240.244
R14451 gnd.n1351 gnd.n1350 240.244
R14452 gnd.n1928 gnd.n1351 240.244
R14453 gnd.n1928 gnd.n1354 240.244
R14454 gnd.n1355 gnd.n1354 240.244
R14455 gnd.n1356 gnd.n1355 240.244
R14456 gnd.n1910 gnd.n1356 240.244
R14457 gnd.n1910 gnd.n1359 240.244
R14458 gnd.n1360 gnd.n1359 240.244
R14459 gnd.n1361 gnd.n1360 240.244
R14460 gnd.n5441 gnd.n1361 240.244
R14461 gnd.n5441 gnd.n1364 240.244
R14462 gnd.n1365 gnd.n1364 240.244
R14463 gnd.n1366 gnd.n1365 240.244
R14464 gnd.n5616 gnd.n1366 240.244
R14465 gnd.n5616 gnd.n1369 240.244
R14466 gnd.n1370 gnd.n1369 240.244
R14467 gnd.n1371 gnd.n1370 240.244
R14468 gnd.n5633 gnd.n1371 240.244
R14469 gnd.n5633 gnd.n1374 240.244
R14470 gnd.n1375 gnd.n1374 240.244
R14471 gnd.n1376 gnd.n1375 240.244
R14472 gnd.n5650 gnd.n1376 240.244
R14473 gnd.n5650 gnd.n1379 240.244
R14474 gnd.n1380 gnd.n1379 240.244
R14475 gnd.n1381 gnd.n1380 240.244
R14476 gnd.n5667 gnd.n1381 240.244
R14477 gnd.n5667 gnd.n1384 240.244
R14478 gnd.n1385 gnd.n1384 240.244
R14479 gnd.n1386 gnd.n1385 240.244
R14480 gnd.n5684 gnd.n1386 240.244
R14481 gnd.n5684 gnd.n1389 240.244
R14482 gnd.n1390 gnd.n1389 240.244
R14483 gnd.n1391 gnd.n1390 240.244
R14484 gnd.n5704 gnd.n1391 240.244
R14485 gnd.n5704 gnd.n1394 240.244
R14486 gnd.n6149 gnd.n1394 240.244
R14487 gnd.n1405 gnd.n1404 240.244
R14488 gnd.n1743 gnd.n1408 240.244
R14489 gnd.n1410 gnd.n1409 240.244
R14490 gnd.n1746 gnd.n1414 240.244
R14491 gnd.n1749 gnd.n1415 240.244
R14492 gnd.n1424 gnd.n1423 240.244
R14493 gnd.n1751 gnd.n1431 240.244
R14494 gnd.n1754 gnd.n1432 240.244
R14495 gnd.n1440 gnd.n1439 240.244
R14496 gnd.n1756 gnd.n1447 240.244
R14497 gnd.n1759 gnd.n1448 240.244
R14498 gnd.n1456 gnd.n1455 240.244
R14499 gnd.n1762 gnd.n1456 240.244
R14500 gnd.n5729 gnd.n1741 240.244
R14501 gnd.n1167 gnd.n1166 240.132
R14502 gnd.n5466 gnd.n5465 240.132
R14503 gnd.n6660 gnd.n766 225.874
R14504 gnd.n6661 gnd.n6660 225.874
R14505 gnd.n6662 gnd.n6661 225.874
R14506 gnd.n6662 gnd.n760 225.874
R14507 gnd.n6670 gnd.n760 225.874
R14508 gnd.n6671 gnd.n6670 225.874
R14509 gnd.n6672 gnd.n6671 225.874
R14510 gnd.n6672 gnd.n754 225.874
R14511 gnd.n6680 gnd.n754 225.874
R14512 gnd.n6681 gnd.n6680 225.874
R14513 gnd.n6682 gnd.n6681 225.874
R14514 gnd.n6682 gnd.n748 225.874
R14515 gnd.n6690 gnd.n748 225.874
R14516 gnd.n6691 gnd.n6690 225.874
R14517 gnd.n6692 gnd.n6691 225.874
R14518 gnd.n6692 gnd.n742 225.874
R14519 gnd.n6700 gnd.n742 225.874
R14520 gnd.n6701 gnd.n6700 225.874
R14521 gnd.n6702 gnd.n6701 225.874
R14522 gnd.n6702 gnd.n736 225.874
R14523 gnd.n6710 gnd.n736 225.874
R14524 gnd.n6711 gnd.n6710 225.874
R14525 gnd.n6712 gnd.n6711 225.874
R14526 gnd.n6712 gnd.n730 225.874
R14527 gnd.n6720 gnd.n730 225.874
R14528 gnd.n6721 gnd.n6720 225.874
R14529 gnd.n6722 gnd.n6721 225.874
R14530 gnd.n6722 gnd.n724 225.874
R14531 gnd.n6730 gnd.n724 225.874
R14532 gnd.n6731 gnd.n6730 225.874
R14533 gnd.n6732 gnd.n6731 225.874
R14534 gnd.n6732 gnd.n718 225.874
R14535 gnd.n6740 gnd.n718 225.874
R14536 gnd.n6741 gnd.n6740 225.874
R14537 gnd.n6742 gnd.n6741 225.874
R14538 gnd.n6742 gnd.n712 225.874
R14539 gnd.n6750 gnd.n712 225.874
R14540 gnd.n6751 gnd.n6750 225.874
R14541 gnd.n6752 gnd.n6751 225.874
R14542 gnd.n6752 gnd.n706 225.874
R14543 gnd.n6760 gnd.n706 225.874
R14544 gnd.n6761 gnd.n6760 225.874
R14545 gnd.n6762 gnd.n6761 225.874
R14546 gnd.n6762 gnd.n700 225.874
R14547 gnd.n6770 gnd.n700 225.874
R14548 gnd.n6771 gnd.n6770 225.874
R14549 gnd.n6772 gnd.n6771 225.874
R14550 gnd.n6772 gnd.n694 225.874
R14551 gnd.n6780 gnd.n694 225.874
R14552 gnd.n6781 gnd.n6780 225.874
R14553 gnd.n6782 gnd.n6781 225.874
R14554 gnd.n6782 gnd.n688 225.874
R14555 gnd.n6790 gnd.n688 225.874
R14556 gnd.n6791 gnd.n6790 225.874
R14557 gnd.n6792 gnd.n6791 225.874
R14558 gnd.n6792 gnd.n682 225.874
R14559 gnd.n6800 gnd.n682 225.874
R14560 gnd.n6801 gnd.n6800 225.874
R14561 gnd.n6802 gnd.n6801 225.874
R14562 gnd.n6802 gnd.n676 225.874
R14563 gnd.n6810 gnd.n676 225.874
R14564 gnd.n6811 gnd.n6810 225.874
R14565 gnd.n6812 gnd.n6811 225.874
R14566 gnd.n6812 gnd.n670 225.874
R14567 gnd.n6820 gnd.n670 225.874
R14568 gnd.n6821 gnd.n6820 225.874
R14569 gnd.n6822 gnd.n6821 225.874
R14570 gnd.n6822 gnd.n664 225.874
R14571 gnd.n6830 gnd.n664 225.874
R14572 gnd.n6831 gnd.n6830 225.874
R14573 gnd.n6832 gnd.n6831 225.874
R14574 gnd.n6832 gnd.n658 225.874
R14575 gnd.n6840 gnd.n658 225.874
R14576 gnd.n6841 gnd.n6840 225.874
R14577 gnd.n6842 gnd.n6841 225.874
R14578 gnd.n6842 gnd.n652 225.874
R14579 gnd.n6850 gnd.n652 225.874
R14580 gnd.n6851 gnd.n6850 225.874
R14581 gnd.n6852 gnd.n6851 225.874
R14582 gnd.n6852 gnd.n646 225.874
R14583 gnd.n6860 gnd.n646 225.874
R14584 gnd.n6861 gnd.n6860 225.874
R14585 gnd.n6862 gnd.n6861 225.874
R14586 gnd.n6862 gnd.n640 225.874
R14587 gnd.n6870 gnd.n640 225.874
R14588 gnd.n6871 gnd.n6870 225.874
R14589 gnd.n6872 gnd.n6871 225.874
R14590 gnd.n6872 gnd.n634 225.874
R14591 gnd.n6880 gnd.n634 225.874
R14592 gnd.n6881 gnd.n6880 225.874
R14593 gnd.n6882 gnd.n6881 225.874
R14594 gnd.n6882 gnd.n628 225.874
R14595 gnd.n6890 gnd.n628 225.874
R14596 gnd.n6891 gnd.n6890 225.874
R14597 gnd.n6892 gnd.n6891 225.874
R14598 gnd.n6892 gnd.n622 225.874
R14599 gnd.n6900 gnd.n622 225.874
R14600 gnd.n6901 gnd.n6900 225.874
R14601 gnd.n6902 gnd.n6901 225.874
R14602 gnd.n6902 gnd.n616 225.874
R14603 gnd.n6910 gnd.n616 225.874
R14604 gnd.n6911 gnd.n6910 225.874
R14605 gnd.n6912 gnd.n6911 225.874
R14606 gnd.n6912 gnd.n610 225.874
R14607 gnd.n6920 gnd.n610 225.874
R14608 gnd.n6921 gnd.n6920 225.874
R14609 gnd.n6922 gnd.n6921 225.874
R14610 gnd.n6922 gnd.n604 225.874
R14611 gnd.n6930 gnd.n604 225.874
R14612 gnd.n6931 gnd.n6930 225.874
R14613 gnd.n6932 gnd.n6931 225.874
R14614 gnd.n6932 gnd.n598 225.874
R14615 gnd.n6940 gnd.n598 225.874
R14616 gnd.n6941 gnd.n6940 225.874
R14617 gnd.n6942 gnd.n6941 225.874
R14618 gnd.n6942 gnd.n592 225.874
R14619 gnd.n6950 gnd.n592 225.874
R14620 gnd.n6951 gnd.n6950 225.874
R14621 gnd.n6952 gnd.n6951 225.874
R14622 gnd.n6952 gnd.n586 225.874
R14623 gnd.n6960 gnd.n586 225.874
R14624 gnd.n6961 gnd.n6960 225.874
R14625 gnd.n6962 gnd.n6961 225.874
R14626 gnd.n6962 gnd.n580 225.874
R14627 gnd.n6970 gnd.n580 225.874
R14628 gnd.n6971 gnd.n6970 225.874
R14629 gnd.n6972 gnd.n6971 225.874
R14630 gnd.n6972 gnd.n574 225.874
R14631 gnd.n6980 gnd.n574 225.874
R14632 gnd.n6981 gnd.n6980 225.874
R14633 gnd.n6982 gnd.n6981 225.874
R14634 gnd.n6982 gnd.n568 225.874
R14635 gnd.n6990 gnd.n568 225.874
R14636 gnd.n6991 gnd.n6990 225.874
R14637 gnd.n6992 gnd.n6991 225.874
R14638 gnd.n6992 gnd.n562 225.874
R14639 gnd.n7000 gnd.n562 225.874
R14640 gnd.n7001 gnd.n7000 225.874
R14641 gnd.n7002 gnd.n7001 225.874
R14642 gnd.n7002 gnd.n556 225.874
R14643 gnd.n7010 gnd.n556 225.874
R14644 gnd.n7011 gnd.n7010 225.874
R14645 gnd.n7012 gnd.n7011 225.874
R14646 gnd.n7012 gnd.n550 225.874
R14647 gnd.n7020 gnd.n550 225.874
R14648 gnd.n7021 gnd.n7020 225.874
R14649 gnd.n7022 gnd.n7021 225.874
R14650 gnd.n7022 gnd.n544 225.874
R14651 gnd.n7030 gnd.n544 225.874
R14652 gnd.n7031 gnd.n7030 225.874
R14653 gnd.n7032 gnd.n7031 225.874
R14654 gnd.n7032 gnd.n538 225.874
R14655 gnd.n7040 gnd.n538 225.874
R14656 gnd.n7041 gnd.n7040 225.874
R14657 gnd.n7042 gnd.n7041 225.874
R14658 gnd.n7042 gnd.n532 225.874
R14659 gnd.n7050 gnd.n532 225.874
R14660 gnd.n7051 gnd.n7050 225.874
R14661 gnd.n7052 gnd.n7051 225.874
R14662 gnd.n7052 gnd.n526 225.874
R14663 gnd.n7060 gnd.n526 225.874
R14664 gnd.n7061 gnd.n7060 225.874
R14665 gnd.n7062 gnd.n7061 225.874
R14666 gnd.n7062 gnd.n520 225.874
R14667 gnd.n7070 gnd.n520 225.874
R14668 gnd.n7071 gnd.n7070 225.874
R14669 gnd.n7072 gnd.n7071 225.874
R14670 gnd.n3220 gnd.t124 224.174
R14671 gnd.n2714 gnd.t107 224.174
R14672 gnd.n1540 gnd.n1477 199.319
R14673 gnd.n1540 gnd.n1478 199.319
R14674 gnd.n1119 gnd.n1118 199.319
R14675 gnd.n2312 gnd.n1119 199.319
R14676 gnd.n1168 gnd.n1165 186.49
R14677 gnd.n5467 gnd.n5464 186.49
R14678 gnd.n3996 gnd.n3995 185
R14679 gnd.n3994 gnd.n3993 185
R14680 gnd.n3973 gnd.n3972 185
R14681 gnd.n3988 gnd.n3987 185
R14682 gnd.n3986 gnd.n3985 185
R14683 gnd.n3977 gnd.n3976 185
R14684 gnd.n3980 gnd.n3979 185
R14685 gnd.n3964 gnd.n3963 185
R14686 gnd.n3962 gnd.n3961 185
R14687 gnd.n3941 gnd.n3940 185
R14688 gnd.n3956 gnd.n3955 185
R14689 gnd.n3954 gnd.n3953 185
R14690 gnd.n3945 gnd.n3944 185
R14691 gnd.n3948 gnd.n3947 185
R14692 gnd.n3932 gnd.n3931 185
R14693 gnd.n3930 gnd.n3929 185
R14694 gnd.n3909 gnd.n3908 185
R14695 gnd.n3924 gnd.n3923 185
R14696 gnd.n3922 gnd.n3921 185
R14697 gnd.n3913 gnd.n3912 185
R14698 gnd.n3916 gnd.n3915 185
R14699 gnd.n3901 gnd.n3900 185
R14700 gnd.n3899 gnd.n3898 185
R14701 gnd.n3878 gnd.n3877 185
R14702 gnd.n3893 gnd.n3892 185
R14703 gnd.n3891 gnd.n3890 185
R14704 gnd.n3882 gnd.n3881 185
R14705 gnd.n3885 gnd.n3884 185
R14706 gnd.n3869 gnd.n3868 185
R14707 gnd.n3867 gnd.n3866 185
R14708 gnd.n3846 gnd.n3845 185
R14709 gnd.n3861 gnd.n3860 185
R14710 gnd.n3859 gnd.n3858 185
R14711 gnd.n3850 gnd.n3849 185
R14712 gnd.n3853 gnd.n3852 185
R14713 gnd.n3837 gnd.n3836 185
R14714 gnd.n3835 gnd.n3834 185
R14715 gnd.n3814 gnd.n3813 185
R14716 gnd.n3829 gnd.n3828 185
R14717 gnd.n3827 gnd.n3826 185
R14718 gnd.n3818 gnd.n3817 185
R14719 gnd.n3821 gnd.n3820 185
R14720 gnd.n3805 gnd.n3804 185
R14721 gnd.n3803 gnd.n3802 185
R14722 gnd.n3782 gnd.n3781 185
R14723 gnd.n3797 gnd.n3796 185
R14724 gnd.n3795 gnd.n3794 185
R14725 gnd.n3786 gnd.n3785 185
R14726 gnd.n3789 gnd.n3788 185
R14727 gnd.n3774 gnd.n3773 185
R14728 gnd.n3772 gnd.n3771 185
R14729 gnd.n3751 gnd.n3750 185
R14730 gnd.n3766 gnd.n3765 185
R14731 gnd.n3764 gnd.n3763 185
R14732 gnd.n3755 gnd.n3754 185
R14733 gnd.n3758 gnd.n3757 185
R14734 gnd.n3221 gnd.t123 178.987
R14735 gnd.n2715 gnd.t108 178.987
R14736 gnd.n1 gnd.t1 170.774
R14737 gnd.n9 gnd.t369 170.103
R14738 gnd.n8 gnd.t181 170.103
R14739 gnd.n7 gnd.t371 170.103
R14740 gnd.n6 gnd.t175 170.103
R14741 gnd.n5 gnd.t143 170.103
R14742 gnd.n4 gnd.t177 170.103
R14743 gnd.n3 gnd.t10 170.103
R14744 gnd.n2 gnd.t136 170.103
R14745 gnd.n1 gnd.t168 170.103
R14746 gnd.n6027 gnd.n1539 164.544
R14747 gnd.n6359 gnd.n6358 164.544
R14748 gnd.n5538 gnd.n5537 163.367
R14749 gnd.n5534 gnd.n5533 163.367
R14750 gnd.n5530 gnd.n5529 163.367
R14751 gnd.n5526 gnd.n5525 163.367
R14752 gnd.n5522 gnd.n5521 163.367
R14753 gnd.n5518 gnd.n5517 163.367
R14754 gnd.n5514 gnd.n5513 163.367
R14755 gnd.n5510 gnd.n5509 163.367
R14756 gnd.n5506 gnd.n5505 163.367
R14757 gnd.n5502 gnd.n5501 163.367
R14758 gnd.n5498 gnd.n5497 163.367
R14759 gnd.n5494 gnd.n5493 163.367
R14760 gnd.n5490 gnd.n5489 163.367
R14761 gnd.n5486 gnd.n5485 163.367
R14762 gnd.n5481 gnd.n5480 163.367
R14763 gnd.n5477 gnd.n5476 163.367
R14764 gnd.n5614 gnd.n5613 163.367
R14765 gnd.n5610 gnd.n5609 163.367
R14766 gnd.n5605 gnd.n5604 163.367
R14767 gnd.n5601 gnd.n5600 163.367
R14768 gnd.n5597 gnd.n5596 163.367
R14769 gnd.n5593 gnd.n5592 163.367
R14770 gnd.n5589 gnd.n5588 163.367
R14771 gnd.n5585 gnd.n5584 163.367
R14772 gnd.n5581 gnd.n5580 163.367
R14773 gnd.n5577 gnd.n5576 163.367
R14774 gnd.n5573 gnd.n5572 163.367
R14775 gnd.n5569 gnd.n5568 163.367
R14776 gnd.n5565 gnd.n5564 163.367
R14777 gnd.n5561 gnd.n5560 163.367
R14778 gnd.n5557 gnd.n5556 163.367
R14779 gnd.n5553 gnd.n5552 163.367
R14780 gnd.n1267 gnd.n1184 163.367
R14781 gnd.n1270 gnd.n1184 163.367
R14782 gnd.n1270 gnd.n1200 163.367
R14783 gnd.n6277 gnd.n1200 163.367
R14784 gnd.n6277 gnd.n1201 163.367
R14785 gnd.n6273 gnd.n1201 163.367
R14786 gnd.n6273 gnd.n1274 163.367
R14787 gnd.n1287 gnd.n1274 163.367
R14788 gnd.n2111 gnd.n1287 163.367
R14789 gnd.n2115 gnd.n2111 163.367
R14790 gnd.n5017 gnd.n2115 163.367
R14791 gnd.n5018 gnd.n5017 163.367
R14792 gnd.n5018 gnd.n2109 163.367
R14793 gnd.n5027 gnd.n2109 163.367
R14794 gnd.n5027 gnd.n2103 163.367
R14795 gnd.n5023 gnd.n2103 163.367
R14796 gnd.n5023 gnd.n2096 163.367
R14797 gnd.n2096 gnd.n2089 163.367
R14798 gnd.n5052 gnd.n2089 163.367
R14799 gnd.n5053 gnd.n5052 163.367
R14800 gnd.n5053 gnd.n2080 163.367
R14801 gnd.n5057 gnd.n2080 163.367
R14802 gnd.n5057 gnd.n2086 163.367
R14803 gnd.n5084 gnd.n2086 163.367
R14804 gnd.n5084 gnd.n2087 163.367
R14805 gnd.n2087 gnd.n2064 163.367
R14806 gnd.n5079 gnd.n2064 163.367
R14807 gnd.n5079 gnd.n2057 163.367
R14808 gnd.n5076 gnd.n2057 163.367
R14809 gnd.n5076 gnd.n5075 163.367
R14810 gnd.n5075 gnd.n5074 163.367
R14811 gnd.n5074 gnd.n5063 163.367
R14812 gnd.n5063 gnd.n2039 163.367
R14813 gnd.n5069 gnd.n2039 163.367
R14814 gnd.n5069 gnd.n2035 163.367
R14815 gnd.n5066 gnd.n2035 163.367
R14816 gnd.n5066 gnd.n2024 163.367
R14817 gnd.n2024 gnd.n2016 163.367
R14818 gnd.n5195 gnd.n2016 163.367
R14819 gnd.n5195 gnd.n2013 163.367
R14820 gnd.n5206 gnd.n2013 163.367
R14821 gnd.n5206 gnd.n2014 163.367
R14822 gnd.n2014 gnd.n2007 163.367
R14823 gnd.n5201 gnd.n2007 163.367
R14824 gnd.n5201 gnd.n1997 163.367
R14825 gnd.n1997 gnd.n1992 163.367
R14826 gnd.n5231 gnd.n1992 163.367
R14827 gnd.n5232 gnd.n5231 163.367
R14828 gnd.n5232 gnd.n1979 163.367
R14829 gnd.n5236 gnd.n1979 163.367
R14830 gnd.n5236 gnd.n1990 163.367
R14831 gnd.n5240 gnd.n1990 163.367
R14832 gnd.n5240 gnd.n1962 163.367
R14833 gnd.n5302 gnd.n1962 163.367
R14834 gnd.n5302 gnd.n1960 163.367
R14835 gnd.n5308 gnd.n1960 163.367
R14836 gnd.n5308 gnd.n1950 163.367
R14837 gnd.n1950 gnd.n1945 163.367
R14838 gnd.n5329 gnd.n1945 163.367
R14839 gnd.n5330 gnd.n5329 163.367
R14840 gnd.n5330 gnd.n1942 163.367
R14841 gnd.n5338 gnd.n1942 163.367
R14842 gnd.n5338 gnd.n1936 163.367
R14843 gnd.n5334 gnd.n1936 163.367
R14844 gnd.n5334 gnd.n1926 163.367
R14845 gnd.n1926 gnd.n1919 163.367
R14846 gnd.n5366 gnd.n1919 163.367
R14847 gnd.n5366 gnd.n1916 163.367
R14848 gnd.n5391 gnd.n1916 163.367
R14849 gnd.n5391 gnd.n1917 163.367
R14850 gnd.n1917 gnd.n1909 163.367
R14851 gnd.n5386 gnd.n1909 163.367
R14852 gnd.n5386 gnd.n5384 163.367
R14853 gnd.n5384 gnd.n5383 163.367
R14854 gnd.n5383 gnd.n5372 163.367
R14855 gnd.n5372 gnd.n1892 163.367
R14856 gnd.n5378 gnd.n1892 163.367
R14857 gnd.n5378 gnd.n1888 163.367
R14858 gnd.n5375 gnd.n1888 163.367
R14859 gnd.n5375 gnd.n1878 163.367
R14860 gnd.n1878 gnd.n1870 163.367
R14861 gnd.n5547 gnd.n1870 163.367
R14862 gnd.n5548 gnd.n5547 163.367
R14863 gnd.n1159 gnd.n1158 163.367
R14864 gnd.n6348 gnd.n1158 163.367
R14865 gnd.n6346 gnd.n6345 163.367
R14866 gnd.n6342 gnd.n6341 163.367
R14867 gnd.n6338 gnd.n6337 163.367
R14868 gnd.n6334 gnd.n6333 163.367
R14869 gnd.n6330 gnd.n6329 163.367
R14870 gnd.n6326 gnd.n6325 163.367
R14871 gnd.n6322 gnd.n6321 163.367
R14872 gnd.n6318 gnd.n6317 163.367
R14873 gnd.n6314 gnd.n6313 163.367
R14874 gnd.n6310 gnd.n6309 163.367
R14875 gnd.n6306 gnd.n6305 163.367
R14876 gnd.n6302 gnd.n6301 163.367
R14877 gnd.n6298 gnd.n6297 163.367
R14878 gnd.n6294 gnd.n6293 163.367
R14879 gnd.n6357 gnd.n1124 163.367
R14880 gnd.n1206 gnd.n1205 163.367
R14881 gnd.n1211 gnd.n1210 163.367
R14882 gnd.n1215 gnd.n1214 163.367
R14883 gnd.n1219 gnd.n1218 163.367
R14884 gnd.n1223 gnd.n1222 163.367
R14885 gnd.n1227 gnd.n1226 163.367
R14886 gnd.n1231 gnd.n1230 163.367
R14887 gnd.n1235 gnd.n1234 163.367
R14888 gnd.n1239 gnd.n1238 163.367
R14889 gnd.n1243 gnd.n1242 163.367
R14890 gnd.n1247 gnd.n1246 163.367
R14891 gnd.n1251 gnd.n1250 163.367
R14892 gnd.n1255 gnd.n1254 163.367
R14893 gnd.n1259 gnd.n1258 163.367
R14894 gnd.n1263 gnd.n1262 163.367
R14895 gnd.n6286 gnd.n1160 163.367
R14896 gnd.n6286 gnd.n1182 163.367
R14897 gnd.n1280 gnd.n1182 163.367
R14898 gnd.n1280 gnd.n1197 163.367
R14899 gnd.n1278 gnd.n1197 163.367
R14900 gnd.n6271 gnd.n1278 163.367
R14901 gnd.n6271 gnd.n1279 163.367
R14902 gnd.n6267 gnd.n1279 163.367
R14903 gnd.n6267 gnd.n1285 163.367
R14904 gnd.n5012 gnd.n1285 163.367
R14905 gnd.n5015 gnd.n5012 163.367
R14906 gnd.n5015 gnd.n2107 163.367
R14907 gnd.n5030 gnd.n2107 163.367
R14908 gnd.n5030 gnd.n2105 163.367
R14909 gnd.n5034 gnd.n2105 163.367
R14910 gnd.n5034 gnd.n2094 163.367
R14911 gnd.n5046 gnd.n2094 163.367
R14912 gnd.n5046 gnd.n2092 163.367
R14913 gnd.n5050 gnd.n2092 163.367
R14914 gnd.n5050 gnd.n2082 163.367
R14915 gnd.n5093 gnd.n2082 163.367
R14916 gnd.n5093 gnd.n2083 163.367
R14917 gnd.n5089 gnd.n2083 163.367
R14918 gnd.n5089 gnd.n5088 163.367
R14919 gnd.n5088 gnd.n2062 163.367
R14920 gnd.n5116 gnd.n2062 163.367
R14921 gnd.n5116 gnd.n2059 163.367
R14922 gnd.n5125 gnd.n2059 163.367
R14923 gnd.n5125 gnd.n2060 163.367
R14924 gnd.n5121 gnd.n2060 163.367
R14925 gnd.n5121 gnd.n5120 163.367
R14926 gnd.n5120 gnd.n2038 163.367
R14927 gnd.n5171 gnd.n2038 163.367
R14928 gnd.n5171 gnd.n2036 163.367
R14929 gnd.n5175 gnd.n2036 163.367
R14930 gnd.n5175 gnd.n2021 163.367
R14931 gnd.n5189 gnd.n2021 163.367
R14932 gnd.n5189 gnd.n2019 163.367
R14933 gnd.n5193 gnd.n2019 163.367
R14934 gnd.n5193 gnd.n2011 163.367
R14935 gnd.n5208 gnd.n2011 163.367
R14936 gnd.n5208 gnd.n2009 163.367
R14937 gnd.n5212 gnd.n2009 163.367
R14938 gnd.n5212 gnd.n1996 163.367
R14939 gnd.n5225 gnd.n1996 163.367
R14940 gnd.n5225 gnd.n1994 163.367
R14941 gnd.n5229 gnd.n1994 163.367
R14942 gnd.n5229 gnd.n1981 163.367
R14943 gnd.n5249 gnd.n1981 163.367
R14944 gnd.n5249 gnd.n1982 163.367
R14945 gnd.n5245 gnd.n1982 163.367
R14946 gnd.n5245 gnd.n5244 163.367
R14947 gnd.n5244 gnd.n1989 163.367
R14948 gnd.n1989 gnd.n1963 163.367
R14949 gnd.n1985 gnd.n1963 163.367
R14950 gnd.n1985 gnd.n1948 163.367
R14951 gnd.n5323 gnd.n1948 163.367
R14952 gnd.n5323 gnd.n1946 163.367
R14953 gnd.n5327 gnd.n1946 163.367
R14954 gnd.n5327 gnd.n1940 163.367
R14955 gnd.n5342 gnd.n1940 163.367
R14956 gnd.n5342 gnd.n1938 163.367
R14957 gnd.n5346 gnd.n1938 163.367
R14958 gnd.n5346 gnd.n1924 163.367
R14959 gnd.n5360 gnd.n1924 163.367
R14960 gnd.n5360 gnd.n1922 163.367
R14961 gnd.n5364 gnd.n1922 163.367
R14962 gnd.n5364 gnd.n1915 163.367
R14963 gnd.n5393 gnd.n1915 163.367
R14964 gnd.n5393 gnd.n1912 163.367
R14965 gnd.n5402 gnd.n1912 163.367
R14966 gnd.n5402 gnd.n1913 163.367
R14967 gnd.n5398 gnd.n1913 163.367
R14968 gnd.n5398 gnd.n5397 163.367
R14969 gnd.n5397 gnd.n1891 163.367
R14970 gnd.n5435 gnd.n1891 163.367
R14971 gnd.n5435 gnd.n1889 163.367
R14972 gnd.n5439 gnd.n1889 163.367
R14973 gnd.n5439 gnd.n1876 163.367
R14974 gnd.n5452 gnd.n1876 163.367
R14975 gnd.n5452 gnd.n1873 163.367
R14976 gnd.n5545 gnd.n1873 163.367
R14977 gnd.n5545 gnd.n1874 163.367
R14978 gnd.n5473 gnd.n5472 156.462
R14979 gnd.n3936 gnd.n3904 153.042
R14980 gnd.n4000 gnd.n3999 152.079
R14981 gnd.n3968 gnd.n3967 152.079
R14982 gnd.n3936 gnd.n3935 152.079
R14983 gnd.n1173 gnd.n1172 152
R14984 gnd.n1174 gnd.n1163 152
R14985 gnd.n1176 gnd.n1175 152
R14986 gnd.n1178 gnd.n1161 152
R14987 gnd.n1180 gnd.n1179 152
R14988 gnd.n5471 gnd.n5455 152
R14989 gnd.n5463 gnd.n5456 152
R14990 gnd.n5462 gnd.n5461 152
R14991 gnd.n5460 gnd.n5457 152
R14992 gnd.n5458 gnd.t62 150.546
R14993 gnd.t365 gnd.n3978 147.661
R14994 gnd.t156 gnd.n3946 147.661
R14995 gnd.t179 gnd.n3914 147.661
R14996 gnd.t164 gnd.n3883 147.661
R14997 gnd.t134 gnd.n3851 147.661
R14998 gnd.t147 gnd.n3819 147.661
R14999 gnd.t153 gnd.n3787 147.661
R15000 gnd.t158 gnd.n3756 147.661
R15001 gnd.n1866 gnd.n1848 143.351
R15002 gnd.n1140 gnd.n1123 143.351
R15003 gnd.n6356 gnd.n1123 143.351
R15004 gnd.n1170 gnd.t18 130.484
R15005 gnd.n1179 gnd.t15 126.766
R15006 gnd.n1177 gnd.t115 126.766
R15007 gnd.n1163 gnd.t128 126.766
R15008 gnd.n1171 gnd.t65 126.766
R15009 gnd.n5459 gnd.t33 126.766
R15010 gnd.n5461 gnd.t77 126.766
R15011 gnd.n5470 gnd.t51 126.766
R15012 gnd.n5472 gnd.t90 126.766
R15013 gnd.n7080 gnd.n514 106.77
R15014 gnd.n7081 gnd.n7080 106.77
R15015 gnd.n7082 gnd.n7081 106.77
R15016 gnd.n7082 gnd.n508 106.77
R15017 gnd.n7090 gnd.n508 106.77
R15018 gnd.n7091 gnd.n7090 106.77
R15019 gnd.n7092 gnd.n7091 106.77
R15020 gnd.n7092 gnd.n502 106.77
R15021 gnd.n7100 gnd.n502 106.77
R15022 gnd.n7101 gnd.n7100 106.77
R15023 gnd.n7102 gnd.n7101 106.77
R15024 gnd.n7102 gnd.n496 106.77
R15025 gnd.n7110 gnd.n496 106.77
R15026 gnd.n7111 gnd.n7110 106.77
R15027 gnd.n7112 gnd.n7111 106.77
R15028 gnd.n7112 gnd.n490 106.77
R15029 gnd.n7120 gnd.n490 106.77
R15030 gnd.n7121 gnd.n7120 106.77
R15031 gnd.n7122 gnd.n7121 106.77
R15032 gnd.n7122 gnd.n484 106.77
R15033 gnd.n7130 gnd.n484 106.77
R15034 gnd.n7131 gnd.n7130 106.77
R15035 gnd.n7132 gnd.n7131 106.77
R15036 gnd.n7132 gnd.n478 106.77
R15037 gnd.n7140 gnd.n478 106.77
R15038 gnd.n7141 gnd.n7140 106.77
R15039 gnd.n7142 gnd.n7141 106.77
R15040 gnd.n7142 gnd.n472 106.77
R15041 gnd.n7150 gnd.n472 106.77
R15042 gnd.n7151 gnd.n7150 106.77
R15043 gnd.n7152 gnd.n7151 106.77
R15044 gnd.n7152 gnd.n466 106.77
R15045 gnd.n7160 gnd.n466 106.77
R15046 gnd.n7161 gnd.n7160 106.77
R15047 gnd.n7162 gnd.n7161 106.77
R15048 gnd.n7162 gnd.n460 106.77
R15049 gnd.n7170 gnd.n460 106.77
R15050 gnd.n7171 gnd.n7170 106.77
R15051 gnd.n7172 gnd.n7171 106.77
R15052 gnd.n7172 gnd.n454 106.77
R15053 gnd.n7180 gnd.n454 106.77
R15054 gnd.n7181 gnd.n7180 106.77
R15055 gnd.n7182 gnd.n7181 106.77
R15056 gnd.n7182 gnd.n448 106.77
R15057 gnd.n7190 gnd.n448 106.77
R15058 gnd.n7191 gnd.n7190 106.77
R15059 gnd.n7192 gnd.n7191 106.77
R15060 gnd.n7192 gnd.n442 106.77
R15061 gnd.n7200 gnd.n442 106.77
R15062 gnd.n7201 gnd.n7200 106.77
R15063 gnd.n7202 gnd.n7201 106.77
R15064 gnd.n7202 gnd.n436 106.77
R15065 gnd.n7210 gnd.n436 106.77
R15066 gnd.n7211 gnd.n7210 106.77
R15067 gnd.n7212 gnd.n7211 106.77
R15068 gnd.n7212 gnd.n430 106.77
R15069 gnd.n7220 gnd.n430 106.77
R15070 gnd.n7221 gnd.n7220 106.77
R15071 gnd.n7222 gnd.n7221 106.77
R15072 gnd.n7222 gnd.n424 106.77
R15073 gnd.n7230 gnd.n424 106.77
R15074 gnd.n7231 gnd.n7230 106.77
R15075 gnd.n7232 gnd.n7231 106.77
R15076 gnd.n7232 gnd.n418 106.77
R15077 gnd.n7240 gnd.n418 106.77
R15078 gnd.n7241 gnd.n7240 106.77
R15079 gnd.n7242 gnd.n7241 106.77
R15080 gnd.n7242 gnd.n412 106.77
R15081 gnd.n7250 gnd.n412 106.77
R15082 gnd.n7251 gnd.n7250 106.77
R15083 gnd.n7252 gnd.n7251 106.77
R15084 gnd.n7252 gnd.n406 106.77
R15085 gnd.n7260 gnd.n406 106.77
R15086 gnd.n7261 gnd.n7260 106.77
R15087 gnd.n7262 gnd.n7261 106.77
R15088 gnd.n7262 gnd.n400 106.77
R15089 gnd.n7270 gnd.n400 106.77
R15090 gnd.n7271 gnd.n7270 106.77
R15091 gnd.n7272 gnd.n7271 106.77
R15092 gnd.n7272 gnd.n394 106.77
R15093 gnd.n7282 gnd.n394 106.77
R15094 gnd.n7283 gnd.n7282 106.77
R15095 gnd.n7284 gnd.n7283 106.77
R15096 gnd.n3995 gnd.n3994 104.615
R15097 gnd.n3994 gnd.n3972 104.615
R15098 gnd.n3987 gnd.n3972 104.615
R15099 gnd.n3987 gnd.n3986 104.615
R15100 gnd.n3986 gnd.n3976 104.615
R15101 gnd.n3979 gnd.n3976 104.615
R15102 gnd.n3963 gnd.n3962 104.615
R15103 gnd.n3962 gnd.n3940 104.615
R15104 gnd.n3955 gnd.n3940 104.615
R15105 gnd.n3955 gnd.n3954 104.615
R15106 gnd.n3954 gnd.n3944 104.615
R15107 gnd.n3947 gnd.n3944 104.615
R15108 gnd.n3931 gnd.n3930 104.615
R15109 gnd.n3930 gnd.n3908 104.615
R15110 gnd.n3923 gnd.n3908 104.615
R15111 gnd.n3923 gnd.n3922 104.615
R15112 gnd.n3922 gnd.n3912 104.615
R15113 gnd.n3915 gnd.n3912 104.615
R15114 gnd.n3900 gnd.n3899 104.615
R15115 gnd.n3899 gnd.n3877 104.615
R15116 gnd.n3892 gnd.n3877 104.615
R15117 gnd.n3892 gnd.n3891 104.615
R15118 gnd.n3891 gnd.n3881 104.615
R15119 gnd.n3884 gnd.n3881 104.615
R15120 gnd.n3868 gnd.n3867 104.615
R15121 gnd.n3867 gnd.n3845 104.615
R15122 gnd.n3860 gnd.n3845 104.615
R15123 gnd.n3860 gnd.n3859 104.615
R15124 gnd.n3859 gnd.n3849 104.615
R15125 gnd.n3852 gnd.n3849 104.615
R15126 gnd.n3836 gnd.n3835 104.615
R15127 gnd.n3835 gnd.n3813 104.615
R15128 gnd.n3828 gnd.n3813 104.615
R15129 gnd.n3828 gnd.n3827 104.615
R15130 gnd.n3827 gnd.n3817 104.615
R15131 gnd.n3820 gnd.n3817 104.615
R15132 gnd.n3804 gnd.n3803 104.615
R15133 gnd.n3803 gnd.n3781 104.615
R15134 gnd.n3796 gnd.n3781 104.615
R15135 gnd.n3796 gnd.n3795 104.615
R15136 gnd.n3795 gnd.n3785 104.615
R15137 gnd.n3788 gnd.n3785 104.615
R15138 gnd.n3773 gnd.n3772 104.615
R15139 gnd.n3772 gnd.n3750 104.615
R15140 gnd.n3765 gnd.n3750 104.615
R15141 gnd.n3765 gnd.n3764 104.615
R15142 gnd.n3764 gnd.n3754 104.615
R15143 gnd.n3757 gnd.n3754 104.615
R15144 gnd.n3146 gnd.t50 100.632
R15145 gnd.n2688 gnd.t85 100.632
R15146 gnd.n7541 gnd.n219 99.6594
R15147 gnd.n7539 gnd.n7538 99.6594
R15148 gnd.n7534 gnd.n226 99.6594
R15149 gnd.n7532 gnd.n7531 99.6594
R15150 gnd.n7527 gnd.n233 99.6594
R15151 gnd.n7525 gnd.n7524 99.6594
R15152 gnd.n7520 gnd.n240 99.6594
R15153 gnd.n7518 gnd.n7517 99.6594
R15154 gnd.n7510 gnd.n247 99.6594
R15155 gnd.n7508 gnd.n7507 99.6594
R15156 gnd.n7503 gnd.n254 99.6594
R15157 gnd.n7501 gnd.n7500 99.6594
R15158 gnd.n7496 gnd.n261 99.6594
R15159 gnd.n7494 gnd.n7493 99.6594
R15160 gnd.n7489 gnd.n268 99.6594
R15161 gnd.n7487 gnd.n7486 99.6594
R15162 gnd.n7482 gnd.n275 99.6594
R15163 gnd.n7480 gnd.n7479 99.6594
R15164 gnd.n285 gnd.n284 99.6594
R15165 gnd.n7471 gnd.n7470 99.6594
R15166 gnd.n7468 gnd.n7467 99.6594
R15167 gnd.n7463 gnd.n293 99.6594
R15168 gnd.n7461 gnd.n7460 99.6594
R15169 gnd.n7456 gnd.n300 99.6594
R15170 gnd.n7454 gnd.n7453 99.6594
R15171 gnd.n7449 gnd.n307 99.6594
R15172 gnd.n7447 gnd.n7446 99.6594
R15173 gnd.n7442 gnd.n316 99.6594
R15174 gnd.n7440 gnd.n7439 99.6594
R15175 gnd.n6079 gnd.n6078 99.6594
R15176 gnd.n6073 gnd.n1466 99.6594
R15177 gnd.n6070 gnd.n1467 99.6594
R15178 gnd.n6066 gnd.n1468 99.6594
R15179 gnd.n6062 gnd.n1469 99.6594
R15180 gnd.n6058 gnd.n1470 99.6594
R15181 gnd.n6054 gnd.n1471 99.6594
R15182 gnd.n6050 gnd.n1472 99.6594
R15183 gnd.n6046 gnd.n1473 99.6594
R15184 gnd.n6041 gnd.n1474 99.6594
R15185 gnd.n6037 gnd.n1475 99.6594
R15186 gnd.n6033 gnd.n1476 99.6594
R15187 gnd.n6029 gnd.n1477 99.6594
R15188 gnd.n6024 gnd.n1479 99.6594
R15189 gnd.n6020 gnd.n1480 99.6594
R15190 gnd.n6016 gnd.n1481 99.6594
R15191 gnd.n6012 gnd.n1482 99.6594
R15192 gnd.n6008 gnd.n1483 99.6594
R15193 gnd.n6004 gnd.n1484 99.6594
R15194 gnd.n6000 gnd.n1485 99.6594
R15195 gnd.n5996 gnd.n1486 99.6594
R15196 gnd.n5992 gnd.n1487 99.6594
R15197 gnd.n5988 gnd.n1488 99.6594
R15198 gnd.n5984 gnd.n1489 99.6594
R15199 gnd.n5980 gnd.n1490 99.6594
R15200 gnd.n5976 gnd.n1491 99.6594
R15201 gnd.n5972 gnd.n1492 99.6594
R15202 gnd.n5968 gnd.n1493 99.6594
R15203 gnd.n6402 gnd.n6401 99.6594
R15204 gnd.n6399 gnd.n6398 99.6594
R15205 gnd.n6394 gnd.n1082 99.6594
R15206 gnd.n6392 gnd.n6391 99.6594
R15207 gnd.n6387 gnd.n1089 99.6594
R15208 gnd.n6385 gnd.n6384 99.6594
R15209 gnd.n6380 gnd.n1096 99.6594
R15210 gnd.n6378 gnd.n6377 99.6594
R15211 gnd.n6372 gnd.n1105 99.6594
R15212 gnd.n6370 gnd.n6369 99.6594
R15213 gnd.n6365 gnd.n1112 99.6594
R15214 gnd.n6363 gnd.n6362 99.6594
R15215 gnd.n2313 gnd.n2312 99.6594
R15216 gnd.n2317 gnd.n2315 99.6594
R15217 gnd.n2323 gnd.n2307 99.6594
R15218 gnd.n2327 gnd.n2325 99.6594
R15219 gnd.n2333 gnd.n2303 99.6594
R15220 gnd.n2337 gnd.n2335 99.6594
R15221 gnd.n2343 gnd.n2297 99.6594
R15222 gnd.n2347 gnd.n2345 99.6594
R15223 gnd.n2353 gnd.n2293 99.6594
R15224 gnd.n2357 gnd.n2355 99.6594
R15225 gnd.n2363 gnd.n2289 99.6594
R15226 gnd.n2367 gnd.n2365 99.6594
R15227 gnd.n2373 gnd.n2285 99.6594
R15228 gnd.n2377 gnd.n2375 99.6594
R15229 gnd.n2383 gnd.n2281 99.6594
R15230 gnd.n2386 gnd.n2385 99.6594
R15231 gnd.n4440 gnd.n4439 99.6594
R15232 gnd.n4434 gnd.n4128 99.6594
R15233 gnd.n4431 gnd.n4129 99.6594
R15234 gnd.n4427 gnd.n4130 99.6594
R15235 gnd.n4423 gnd.n4131 99.6594
R15236 gnd.n4419 gnd.n4132 99.6594
R15237 gnd.n4415 gnd.n4133 99.6594
R15238 gnd.n4411 gnd.n4134 99.6594
R15239 gnd.n4407 gnd.n4135 99.6594
R15240 gnd.n4402 gnd.n4136 99.6594
R15241 gnd.n4398 gnd.n4137 99.6594
R15242 gnd.n4394 gnd.n4138 99.6594
R15243 gnd.n4390 gnd.n4139 99.6594
R15244 gnd.n4386 gnd.n4140 99.6594
R15245 gnd.n4382 gnd.n4141 99.6594
R15246 gnd.n4378 gnd.n4142 99.6594
R15247 gnd.n4374 gnd.n4143 99.6594
R15248 gnd.n4370 gnd.n4144 99.6594
R15249 gnd.n4366 gnd.n4145 99.6594
R15250 gnd.n4362 gnd.n4146 99.6594
R15251 gnd.n4358 gnd.n4147 99.6594
R15252 gnd.n4354 gnd.n4148 99.6594
R15253 gnd.n4350 gnd.n4149 99.6594
R15254 gnd.n4346 gnd.n4150 99.6594
R15255 gnd.n4342 gnd.n4151 99.6594
R15256 gnd.n4338 gnd.n4152 99.6594
R15257 gnd.n4334 gnd.n4153 99.6594
R15258 gnd.n4330 gnd.n4154 99.6594
R15259 gnd.n4442 gnd.n2648 99.6594
R15260 gnd.n4118 gnd.n2671 99.6594
R15261 gnd.n4116 gnd.n2670 99.6594
R15262 gnd.n4112 gnd.n2669 99.6594
R15263 gnd.n4108 gnd.n2668 99.6594
R15264 gnd.n4104 gnd.n2667 99.6594
R15265 gnd.n4100 gnd.n2666 99.6594
R15266 gnd.n4096 gnd.n2665 99.6594
R15267 gnd.n4028 gnd.n2664 99.6594
R15268 gnd.n3358 gnd.n3089 99.6594
R15269 gnd.n3115 gnd.n3096 99.6594
R15270 gnd.n3117 gnd.n3097 99.6594
R15271 gnd.n3125 gnd.n3098 99.6594
R15272 gnd.n3127 gnd.n3099 99.6594
R15273 gnd.n3135 gnd.n3100 99.6594
R15274 gnd.n3137 gnd.n3101 99.6594
R15275 gnd.n3145 gnd.n3102 99.6594
R15276 gnd.n7431 gnd.n322 99.6594
R15277 gnd.n7429 gnd.n7428 99.6594
R15278 gnd.n7424 gnd.n329 99.6594
R15279 gnd.n7422 gnd.n7421 99.6594
R15280 gnd.n7417 gnd.n336 99.6594
R15281 gnd.n7415 gnd.n7414 99.6594
R15282 gnd.n7410 gnd.n343 99.6594
R15283 gnd.n7408 gnd.n7407 99.6594
R15284 gnd.n348 gnd.n347 99.6594
R15285 gnd.n1578 gnd.n1494 99.6594
R15286 gnd.n1496 gnd.n1420 99.6594
R15287 gnd.n1497 gnd.n1427 99.6594
R15288 gnd.n1499 gnd.n1498 99.6594
R15289 gnd.n1501 gnd.n1436 99.6594
R15290 gnd.n1502 gnd.n1443 99.6594
R15291 gnd.n1504 gnd.n1503 99.6594
R15292 gnd.n1506 gnd.n1452 99.6594
R15293 gnd.n6081 gnd.n1461 99.6594
R15294 gnd.n4086 gnd.n2651 99.6594
R15295 gnd.n4082 gnd.n2652 99.6594
R15296 gnd.n4078 gnd.n2653 99.6594
R15297 gnd.n4074 gnd.n2654 99.6594
R15298 gnd.n4070 gnd.n2655 99.6594
R15299 gnd.n4066 gnd.n2656 99.6594
R15300 gnd.n4062 gnd.n2657 99.6594
R15301 gnd.n4058 gnd.n2658 99.6594
R15302 gnd.n4054 gnd.n2659 99.6594
R15303 gnd.n4050 gnd.n2660 99.6594
R15304 gnd.n4046 gnd.n2661 99.6594
R15305 gnd.n4042 gnd.n2662 99.6594
R15306 gnd.n4038 gnd.n2663 99.6594
R15307 gnd.n3273 gnd.n3272 99.6594
R15308 gnd.n3267 gnd.n3184 99.6594
R15309 gnd.n3264 gnd.n3185 99.6594
R15310 gnd.n3260 gnd.n3186 99.6594
R15311 gnd.n3256 gnd.n3187 99.6594
R15312 gnd.n3252 gnd.n3188 99.6594
R15313 gnd.n3248 gnd.n3189 99.6594
R15314 gnd.n3244 gnd.n3190 99.6594
R15315 gnd.n3240 gnd.n3191 99.6594
R15316 gnd.n3236 gnd.n3192 99.6594
R15317 gnd.n3232 gnd.n3193 99.6594
R15318 gnd.n3228 gnd.n3194 99.6594
R15319 gnd.n3275 gnd.n3183 99.6594
R15320 gnd.n2401 gnd.n2400 99.6594
R15321 gnd.n2412 gnd.n2411 99.6594
R15322 gnd.n2421 gnd.n2420 99.6594
R15323 gnd.n2424 gnd.n2423 99.6594
R15324 gnd.n2435 gnd.n2434 99.6594
R15325 gnd.n2444 gnd.n2443 99.6594
R15326 gnd.n2447 gnd.n2446 99.6594
R15327 gnd.n2459 gnd.n2458 99.6594
R15328 gnd.n4794 gnd.n4793 99.6594
R15329 gnd.n4320 gnd.n4155 99.6594
R15330 gnd.n4317 gnd.n4156 99.6594
R15331 gnd.n4313 gnd.n4157 99.6594
R15332 gnd.n4309 gnd.n4158 99.6594
R15333 gnd.n4305 gnd.n4159 99.6594
R15334 gnd.n4301 gnd.n4160 99.6594
R15335 gnd.n4297 gnd.n4161 99.6594
R15336 gnd.n4293 gnd.n4162 99.6594
R15337 gnd.n4289 gnd.n4163 99.6594
R15338 gnd.n4318 gnd.n4155 99.6594
R15339 gnd.n4314 gnd.n4156 99.6594
R15340 gnd.n4310 gnd.n4157 99.6594
R15341 gnd.n4306 gnd.n4158 99.6594
R15342 gnd.n4302 gnd.n4159 99.6594
R15343 gnd.n4298 gnd.n4160 99.6594
R15344 gnd.n4294 gnd.n4161 99.6594
R15345 gnd.n4290 gnd.n4162 99.6594
R15346 gnd.n4245 gnd.n4163 99.6594
R15347 gnd.n4793 gnd.n2463 99.6594
R15348 gnd.n2458 gnd.n2457 99.6594
R15349 gnd.n2446 gnd.n2445 99.6594
R15350 gnd.n2443 gnd.n2436 99.6594
R15351 gnd.n2434 gnd.n2433 99.6594
R15352 gnd.n2423 gnd.n2422 99.6594
R15353 gnd.n2420 gnd.n2413 99.6594
R15354 gnd.n2411 gnd.n2410 99.6594
R15355 gnd.n2400 gnd.n2399 99.6594
R15356 gnd.n3273 gnd.n3196 99.6594
R15357 gnd.n3265 gnd.n3184 99.6594
R15358 gnd.n3261 gnd.n3185 99.6594
R15359 gnd.n3257 gnd.n3186 99.6594
R15360 gnd.n3253 gnd.n3187 99.6594
R15361 gnd.n3249 gnd.n3188 99.6594
R15362 gnd.n3245 gnd.n3189 99.6594
R15363 gnd.n3241 gnd.n3190 99.6594
R15364 gnd.n3237 gnd.n3191 99.6594
R15365 gnd.n3233 gnd.n3192 99.6594
R15366 gnd.n3229 gnd.n3193 99.6594
R15367 gnd.n3225 gnd.n3194 99.6594
R15368 gnd.n3276 gnd.n3275 99.6594
R15369 gnd.n4041 gnd.n2663 99.6594
R15370 gnd.n4045 gnd.n2662 99.6594
R15371 gnd.n4049 gnd.n2661 99.6594
R15372 gnd.n4053 gnd.n2660 99.6594
R15373 gnd.n4057 gnd.n2659 99.6594
R15374 gnd.n4061 gnd.n2658 99.6594
R15375 gnd.n4065 gnd.n2657 99.6594
R15376 gnd.n4069 gnd.n2656 99.6594
R15377 gnd.n4073 gnd.n2655 99.6594
R15378 gnd.n4077 gnd.n2654 99.6594
R15379 gnd.n4081 gnd.n2653 99.6594
R15380 gnd.n4085 gnd.n2652 99.6594
R15381 gnd.n2692 gnd.n2651 99.6594
R15382 gnd.n1494 gnd.n1419 99.6594
R15383 gnd.n1496 gnd.n1495 99.6594
R15384 gnd.n1497 gnd.n1428 99.6594
R15385 gnd.n1499 gnd.n1435 99.6594
R15386 gnd.n1501 gnd.n1500 99.6594
R15387 gnd.n1502 gnd.n1444 99.6594
R15388 gnd.n1504 gnd.n1451 99.6594
R15389 gnd.n1506 gnd.n1505 99.6594
R15390 gnd.n6082 gnd.n6081 99.6594
R15391 gnd.n347 gnd.n344 99.6594
R15392 gnd.n7409 gnd.n7408 99.6594
R15393 gnd.n343 gnd.n337 99.6594
R15394 gnd.n7416 gnd.n7415 99.6594
R15395 gnd.n336 gnd.n330 99.6594
R15396 gnd.n7423 gnd.n7422 99.6594
R15397 gnd.n329 gnd.n323 99.6594
R15398 gnd.n7430 gnd.n7429 99.6594
R15399 gnd.n322 gnd.n319 99.6594
R15400 gnd.n3359 gnd.n3358 99.6594
R15401 gnd.n3118 gnd.n3096 99.6594
R15402 gnd.n3124 gnd.n3097 99.6594
R15403 gnd.n3128 gnd.n3098 99.6594
R15404 gnd.n3134 gnd.n3099 99.6594
R15405 gnd.n3138 gnd.n3100 99.6594
R15406 gnd.n3144 gnd.n3101 99.6594
R15407 gnd.n3102 gnd.n3086 99.6594
R15408 gnd.n4095 gnd.n2664 99.6594
R15409 gnd.n4099 gnd.n2665 99.6594
R15410 gnd.n4103 gnd.n2666 99.6594
R15411 gnd.n4107 gnd.n2667 99.6594
R15412 gnd.n4111 gnd.n2668 99.6594
R15413 gnd.n4115 gnd.n2669 99.6594
R15414 gnd.n4119 gnd.n2670 99.6594
R15415 gnd.n2673 gnd.n2671 99.6594
R15416 gnd.n4440 gnd.n4166 99.6594
R15417 gnd.n4432 gnd.n4128 99.6594
R15418 gnd.n4428 gnd.n4129 99.6594
R15419 gnd.n4424 gnd.n4130 99.6594
R15420 gnd.n4420 gnd.n4131 99.6594
R15421 gnd.n4416 gnd.n4132 99.6594
R15422 gnd.n4412 gnd.n4133 99.6594
R15423 gnd.n4408 gnd.n4134 99.6594
R15424 gnd.n4403 gnd.n4135 99.6594
R15425 gnd.n4399 gnd.n4136 99.6594
R15426 gnd.n4395 gnd.n4137 99.6594
R15427 gnd.n4391 gnd.n4138 99.6594
R15428 gnd.n4387 gnd.n4139 99.6594
R15429 gnd.n4383 gnd.n4140 99.6594
R15430 gnd.n4379 gnd.n4141 99.6594
R15431 gnd.n4375 gnd.n4142 99.6594
R15432 gnd.n4371 gnd.n4143 99.6594
R15433 gnd.n4367 gnd.n4144 99.6594
R15434 gnd.n4363 gnd.n4145 99.6594
R15435 gnd.n4359 gnd.n4146 99.6594
R15436 gnd.n4355 gnd.n4147 99.6594
R15437 gnd.n4351 gnd.n4148 99.6594
R15438 gnd.n4347 gnd.n4149 99.6594
R15439 gnd.n4343 gnd.n4150 99.6594
R15440 gnd.n4339 gnd.n4151 99.6594
R15441 gnd.n4335 gnd.n4152 99.6594
R15442 gnd.n4331 gnd.n4153 99.6594
R15443 gnd.n4327 gnd.n4154 99.6594
R15444 gnd.n4443 gnd.n4442 99.6594
R15445 gnd.n2385 gnd.n2384 99.6594
R15446 gnd.n2376 gnd.n2281 99.6594
R15447 gnd.n2375 gnd.n2374 99.6594
R15448 gnd.n2366 gnd.n2285 99.6594
R15449 gnd.n2365 gnd.n2364 99.6594
R15450 gnd.n2356 gnd.n2289 99.6594
R15451 gnd.n2355 gnd.n2354 99.6594
R15452 gnd.n2346 gnd.n2293 99.6594
R15453 gnd.n2345 gnd.n2344 99.6594
R15454 gnd.n2336 gnd.n2297 99.6594
R15455 gnd.n2335 gnd.n2334 99.6594
R15456 gnd.n2326 gnd.n2303 99.6594
R15457 gnd.n2325 gnd.n2324 99.6594
R15458 gnd.n2316 gnd.n2307 99.6594
R15459 gnd.n2315 gnd.n2314 99.6594
R15460 gnd.n1118 gnd.n1113 99.6594
R15461 gnd.n6364 gnd.n6363 99.6594
R15462 gnd.n1112 gnd.n1106 99.6594
R15463 gnd.n6371 gnd.n6370 99.6594
R15464 gnd.n1105 gnd.n1097 99.6594
R15465 gnd.n6379 gnd.n6378 99.6594
R15466 gnd.n1096 gnd.n1090 99.6594
R15467 gnd.n6386 gnd.n6385 99.6594
R15468 gnd.n1089 gnd.n1083 99.6594
R15469 gnd.n6393 gnd.n6392 99.6594
R15470 gnd.n1082 gnd.n1075 99.6594
R15471 gnd.n6400 gnd.n6399 99.6594
R15472 gnd.n6403 gnd.n6402 99.6594
R15473 gnd.n6079 gnd.n1509 99.6594
R15474 gnd.n6071 gnd.n1466 99.6594
R15475 gnd.n6067 gnd.n1467 99.6594
R15476 gnd.n6063 gnd.n1468 99.6594
R15477 gnd.n6059 gnd.n1469 99.6594
R15478 gnd.n6055 gnd.n1470 99.6594
R15479 gnd.n6051 gnd.n1471 99.6594
R15480 gnd.n6047 gnd.n1472 99.6594
R15481 gnd.n6042 gnd.n1473 99.6594
R15482 gnd.n6038 gnd.n1474 99.6594
R15483 gnd.n6034 gnd.n1475 99.6594
R15484 gnd.n6030 gnd.n1476 99.6594
R15485 gnd.n6025 gnd.n1478 99.6594
R15486 gnd.n6021 gnd.n1479 99.6594
R15487 gnd.n6017 gnd.n1480 99.6594
R15488 gnd.n6013 gnd.n1481 99.6594
R15489 gnd.n6009 gnd.n1482 99.6594
R15490 gnd.n6005 gnd.n1483 99.6594
R15491 gnd.n6001 gnd.n1484 99.6594
R15492 gnd.n5997 gnd.n1485 99.6594
R15493 gnd.n5993 gnd.n1486 99.6594
R15494 gnd.n5989 gnd.n1487 99.6594
R15495 gnd.n5985 gnd.n1488 99.6594
R15496 gnd.n5981 gnd.n1489 99.6594
R15497 gnd.n5977 gnd.n1490 99.6594
R15498 gnd.n5973 gnd.n1491 99.6594
R15499 gnd.n5969 gnd.n1492 99.6594
R15500 gnd.n5961 gnd.n1493 99.6594
R15501 gnd.n7441 gnd.n7440 99.6594
R15502 gnd.n316 gnd.n308 99.6594
R15503 gnd.n7448 gnd.n7447 99.6594
R15504 gnd.n307 gnd.n301 99.6594
R15505 gnd.n7455 gnd.n7454 99.6594
R15506 gnd.n300 gnd.n294 99.6594
R15507 gnd.n7462 gnd.n7461 99.6594
R15508 gnd.n293 gnd.n287 99.6594
R15509 gnd.n7469 gnd.n7468 99.6594
R15510 gnd.n7472 gnd.n7471 99.6594
R15511 gnd.n284 gnd.n276 99.6594
R15512 gnd.n7481 gnd.n7480 99.6594
R15513 gnd.n275 gnd.n269 99.6594
R15514 gnd.n7488 gnd.n7487 99.6594
R15515 gnd.n268 gnd.n262 99.6594
R15516 gnd.n7495 gnd.n7494 99.6594
R15517 gnd.n261 gnd.n255 99.6594
R15518 gnd.n7502 gnd.n7501 99.6594
R15519 gnd.n254 gnd.n248 99.6594
R15520 gnd.n7509 gnd.n7508 99.6594
R15521 gnd.n247 gnd.n241 99.6594
R15522 gnd.n7519 gnd.n7518 99.6594
R15523 gnd.n240 gnd.n234 99.6594
R15524 gnd.n7526 gnd.n7525 99.6594
R15525 gnd.n233 gnd.n227 99.6594
R15526 gnd.n7533 gnd.n7532 99.6594
R15527 gnd.n226 gnd.n220 99.6594
R15528 gnd.n7540 gnd.n7539 99.6594
R15529 gnd.n219 gnd.n216 99.6594
R15530 gnd.n4856 gnd.n4855 99.6594
R15531 gnd.n2273 gnd.n2204 99.6594
R15532 gnd.n2275 gnd.n2205 99.6594
R15533 gnd.n2392 gnd.n2206 99.6594
R15534 gnd.n2394 gnd.n2207 99.6594
R15535 gnd.n2405 gnd.n2208 99.6594
R15536 gnd.n2407 gnd.n2209 99.6594
R15537 gnd.n2417 gnd.n2210 99.6594
R15538 gnd.n2428 gnd.n2211 99.6594
R15539 gnd.n2430 gnd.n2212 99.6594
R15540 gnd.n2440 gnd.n2213 99.6594
R15541 gnd.n2451 gnd.n2214 99.6594
R15542 gnd.n4784 gnd.n2215 99.6594
R15543 gnd.n4788 gnd.n2216 99.6594
R15544 gnd.n4856 gnd.n2218 99.6594
R15545 gnd.n2274 gnd.n2204 99.6594
R15546 gnd.n2391 gnd.n2205 99.6594
R15547 gnd.n2393 gnd.n2206 99.6594
R15548 gnd.n2404 gnd.n2207 99.6594
R15549 gnd.n2406 gnd.n2208 99.6594
R15550 gnd.n2416 gnd.n2209 99.6594
R15551 gnd.n2427 gnd.n2210 99.6594
R15552 gnd.n2429 gnd.n2211 99.6594
R15553 gnd.n2439 gnd.n2212 99.6594
R15554 gnd.n2450 gnd.n2213 99.6594
R15555 gnd.n2452 gnd.n2214 99.6594
R15556 gnd.n4787 gnd.n2215 99.6594
R15557 gnd.n2216 gnd.n2194 99.6594
R15558 gnd.n1742 gnd.n1404 99.6594
R15559 gnd.n1744 gnd.n1743 99.6594
R15560 gnd.n1745 gnd.n1409 99.6594
R15561 gnd.n1747 gnd.n1746 99.6594
R15562 gnd.n1748 gnd.n1415 99.6594
R15563 gnd.n1750 gnd.n1423 99.6594
R15564 gnd.n1752 gnd.n1751 99.6594
R15565 gnd.n1753 gnd.n1432 99.6594
R15566 gnd.n1755 gnd.n1439 99.6594
R15567 gnd.n1757 gnd.n1756 99.6594
R15568 gnd.n1758 gnd.n1448 99.6594
R15569 gnd.n1760 gnd.n1455 99.6594
R15570 gnd.n1763 gnd.n1762 99.6594
R15571 gnd.n5729 gnd.n5728 99.6594
R15572 gnd.n1760 gnd.n1759 99.6594
R15573 gnd.n1758 gnd.n1447 99.6594
R15574 gnd.n1757 gnd.n1440 99.6594
R15575 gnd.n1755 gnd.n1754 99.6594
R15576 gnd.n1753 gnd.n1431 99.6594
R15577 gnd.n1752 gnd.n1424 99.6594
R15578 gnd.n1750 gnd.n1749 99.6594
R15579 gnd.n1748 gnd.n1414 99.6594
R15580 gnd.n1747 gnd.n1410 99.6594
R15581 gnd.n1745 gnd.n1408 99.6594
R15582 gnd.n1744 gnd.n1405 99.6594
R15583 gnd.n1742 gnd.n1400 99.6594
R15584 gnd.n5728 gnd.n1395 99.6594
R15585 gnd.n1763 gnd.n1741 99.6594
R15586 gnd.n2453 gnd.t61 98.63
R15587 gnd.n6083 gnd.t14 98.63
R15588 gnd.n2460 gnd.t56 98.63
R15589 gnd.n1529 gnd.t114 98.63
R15590 gnd.n1552 gnd.t120 98.63
R15591 gnd.n5963 gnd.t70 98.63
R15592 gnd.n313 gnd.t94 98.63
R15593 gnd.n280 gnd.t45 98.63
R15594 gnd.n7512 gnd.t88 98.63
R15595 gnd.n350 gnd.t38 98.63
R15596 gnd.n4185 gnd.t73 98.63
R15597 gnd.n4207 gnd.t76 98.63
R15598 gnd.n4228 gnd.t24 98.63
R15599 gnd.n4246 gnd.t101 98.63
R15600 gnd.n1101 gnd.t81 98.63
R15601 gnd.n2278 gnd.t103 98.63
R15602 gnd.n2300 gnd.t126 98.63
R15603 gnd.n1457 gnd.t27 98.63
R15604 gnd.n1202 gnd.t111 92.8196
R15605 gnd.n1867 gnd.t42 92.8196
R15606 gnd.n6290 gnd.t32 92.8118
R15607 gnd.n5474 gnd.t97 92.8118
R15608 gnd.n1170 gnd.n1169 81.8399
R15609 gnd.n3147 gnd.t49 74.8376
R15610 gnd.n2689 gnd.t86 74.8376
R15611 gnd.n1203 gnd.t110 72.8438
R15612 gnd.n1868 gnd.t43 72.8438
R15613 gnd.n1171 gnd.n1164 72.8411
R15614 gnd.n1177 gnd.n1162 72.8411
R15615 gnd.n5470 gnd.n5469 72.8411
R15616 gnd.n2454 gnd.t60 72.836
R15617 gnd.n6291 gnd.t31 72.836
R15618 gnd.n5475 gnd.t98 72.836
R15619 gnd.n6084 gnd.t13 72.836
R15620 gnd.n2461 gnd.t57 72.836
R15621 gnd.n1530 gnd.t113 72.836
R15622 gnd.n1553 gnd.t119 72.836
R15623 gnd.n5964 gnd.t69 72.836
R15624 gnd.n314 gnd.t95 72.836
R15625 gnd.n281 gnd.t46 72.836
R15626 gnd.n7513 gnd.t89 72.836
R15627 gnd.n351 gnd.t39 72.836
R15628 gnd.n4186 gnd.t72 72.836
R15629 gnd.n4208 gnd.t75 72.836
R15630 gnd.n4229 gnd.t23 72.836
R15631 gnd.n4247 gnd.t100 72.836
R15632 gnd.n1102 gnd.t82 72.836
R15633 gnd.n2279 gnd.t104 72.836
R15634 gnd.n2301 gnd.t127 72.836
R15635 gnd.n1458 gnd.t28 72.836
R15636 gnd.n5538 gnd.n1832 71.676
R15637 gnd.n5534 gnd.n1833 71.676
R15638 gnd.n5530 gnd.n1834 71.676
R15639 gnd.n5526 gnd.n1835 71.676
R15640 gnd.n5522 gnd.n1836 71.676
R15641 gnd.n5518 gnd.n1837 71.676
R15642 gnd.n5514 gnd.n1838 71.676
R15643 gnd.n5510 gnd.n1839 71.676
R15644 gnd.n5506 gnd.n1840 71.676
R15645 gnd.n5502 gnd.n1841 71.676
R15646 gnd.n5498 gnd.n1842 71.676
R15647 gnd.n5494 gnd.n1843 71.676
R15648 gnd.n5490 gnd.n1844 71.676
R15649 gnd.n5486 gnd.n1845 71.676
R15650 gnd.n5481 gnd.n1846 71.676
R15651 gnd.n5477 gnd.n1847 71.676
R15652 gnd.n5614 gnd.n1866 71.676
R15653 gnd.n5610 gnd.n1865 71.676
R15654 gnd.n5605 gnd.n1864 71.676
R15655 gnd.n5601 gnd.n1863 71.676
R15656 gnd.n5597 gnd.n1862 71.676
R15657 gnd.n5593 gnd.n1861 71.676
R15658 gnd.n5589 gnd.n1860 71.676
R15659 gnd.n5585 gnd.n1859 71.676
R15660 gnd.n5581 gnd.n1858 71.676
R15661 gnd.n5577 gnd.n1857 71.676
R15662 gnd.n5573 gnd.n1856 71.676
R15663 gnd.n5569 gnd.n1855 71.676
R15664 gnd.n5565 gnd.n1854 71.676
R15665 gnd.n5561 gnd.n1853 71.676
R15666 gnd.n5557 gnd.n1852 71.676
R15667 gnd.n5553 gnd.n1851 71.676
R15668 gnd.n5549 gnd.n1850 71.676
R15669 gnd.n6354 gnd.n6353 71.676
R15670 gnd.n6348 gnd.n1126 71.676
R15671 gnd.n6345 gnd.n1127 71.676
R15672 gnd.n6341 gnd.n1128 71.676
R15673 gnd.n6337 gnd.n1129 71.676
R15674 gnd.n6333 gnd.n1130 71.676
R15675 gnd.n6329 gnd.n1131 71.676
R15676 gnd.n6325 gnd.n1132 71.676
R15677 gnd.n6321 gnd.n1133 71.676
R15678 gnd.n6317 gnd.n1134 71.676
R15679 gnd.n6313 gnd.n1135 71.676
R15680 gnd.n6309 gnd.n1136 71.676
R15681 gnd.n6305 gnd.n1137 71.676
R15682 gnd.n6301 gnd.n1138 71.676
R15683 gnd.n6297 gnd.n1139 71.676
R15684 gnd.n6293 gnd.n1140 71.676
R15685 gnd.n1141 gnd.n1124 71.676
R15686 gnd.n1206 gnd.n1142 71.676
R15687 gnd.n1211 gnd.n1143 71.676
R15688 gnd.n1215 gnd.n1144 71.676
R15689 gnd.n1219 gnd.n1145 71.676
R15690 gnd.n1223 gnd.n1146 71.676
R15691 gnd.n1227 gnd.n1147 71.676
R15692 gnd.n1231 gnd.n1148 71.676
R15693 gnd.n1235 gnd.n1149 71.676
R15694 gnd.n1239 gnd.n1150 71.676
R15695 gnd.n1243 gnd.n1151 71.676
R15696 gnd.n1247 gnd.n1152 71.676
R15697 gnd.n1251 gnd.n1153 71.676
R15698 gnd.n1255 gnd.n1154 71.676
R15699 gnd.n1259 gnd.n1155 71.676
R15700 gnd.n1263 gnd.n1156 71.676
R15701 gnd.n6354 gnd.n1159 71.676
R15702 gnd.n6346 gnd.n1126 71.676
R15703 gnd.n6342 gnd.n1127 71.676
R15704 gnd.n6338 gnd.n1128 71.676
R15705 gnd.n6334 gnd.n1129 71.676
R15706 gnd.n6330 gnd.n1130 71.676
R15707 gnd.n6326 gnd.n1131 71.676
R15708 gnd.n6322 gnd.n1132 71.676
R15709 gnd.n6318 gnd.n1133 71.676
R15710 gnd.n6314 gnd.n1134 71.676
R15711 gnd.n6310 gnd.n1135 71.676
R15712 gnd.n6306 gnd.n1136 71.676
R15713 gnd.n6302 gnd.n1137 71.676
R15714 gnd.n6298 gnd.n1138 71.676
R15715 gnd.n6294 gnd.n1139 71.676
R15716 gnd.n6357 gnd.n6356 71.676
R15717 gnd.n1205 gnd.n1141 71.676
R15718 gnd.n1210 gnd.n1142 71.676
R15719 gnd.n1214 gnd.n1143 71.676
R15720 gnd.n1218 gnd.n1144 71.676
R15721 gnd.n1222 gnd.n1145 71.676
R15722 gnd.n1226 gnd.n1146 71.676
R15723 gnd.n1230 gnd.n1147 71.676
R15724 gnd.n1234 gnd.n1148 71.676
R15725 gnd.n1238 gnd.n1149 71.676
R15726 gnd.n1242 gnd.n1150 71.676
R15727 gnd.n1246 gnd.n1151 71.676
R15728 gnd.n1250 gnd.n1152 71.676
R15729 gnd.n1254 gnd.n1153 71.676
R15730 gnd.n1258 gnd.n1154 71.676
R15731 gnd.n1262 gnd.n1155 71.676
R15732 gnd.n1266 gnd.n1156 71.676
R15733 gnd.n5552 gnd.n1850 71.676
R15734 gnd.n5556 gnd.n1851 71.676
R15735 gnd.n5560 gnd.n1852 71.676
R15736 gnd.n5564 gnd.n1853 71.676
R15737 gnd.n5568 gnd.n1854 71.676
R15738 gnd.n5572 gnd.n1855 71.676
R15739 gnd.n5576 gnd.n1856 71.676
R15740 gnd.n5580 gnd.n1857 71.676
R15741 gnd.n5584 gnd.n1858 71.676
R15742 gnd.n5588 gnd.n1859 71.676
R15743 gnd.n5592 gnd.n1860 71.676
R15744 gnd.n5596 gnd.n1861 71.676
R15745 gnd.n5600 gnd.n1862 71.676
R15746 gnd.n5604 gnd.n1863 71.676
R15747 gnd.n5609 gnd.n1864 71.676
R15748 gnd.n5613 gnd.n1865 71.676
R15749 gnd.n5476 gnd.n1848 71.676
R15750 gnd.n5480 gnd.n1847 71.676
R15751 gnd.n5485 gnd.n1846 71.676
R15752 gnd.n5489 gnd.n1845 71.676
R15753 gnd.n5493 gnd.n1844 71.676
R15754 gnd.n5497 gnd.n1843 71.676
R15755 gnd.n5501 gnd.n1842 71.676
R15756 gnd.n5505 gnd.n1841 71.676
R15757 gnd.n5509 gnd.n1840 71.676
R15758 gnd.n5513 gnd.n1839 71.676
R15759 gnd.n5517 gnd.n1838 71.676
R15760 gnd.n5521 gnd.n1837 71.676
R15761 gnd.n5525 gnd.n1836 71.676
R15762 gnd.n5529 gnd.n1835 71.676
R15763 gnd.n5533 gnd.n1834 71.676
R15764 gnd.n5537 gnd.n1833 71.676
R15765 gnd.n5540 gnd.n1832 71.676
R15766 gnd.n10 gnd.t359 69.1507
R15767 gnd.n18 gnd.t172 68.4792
R15768 gnd.n17 gnd.t7 68.4792
R15769 gnd.n16 gnd.t166 68.4792
R15770 gnd.n15 gnd.t160 68.4792
R15771 gnd.n14 gnd.t150 68.4792
R15772 gnd.n13 gnd.t367 68.4792
R15773 gnd.n12 gnd.t361 68.4792
R15774 gnd.n11 gnd.t170 68.4792
R15775 gnd.n10 gnd.t363 68.4792
R15776 gnd.n3274 gnd.n3178 64.369
R15777 gnd.n7284 gnd.n184 64.0626
R15778 gnd.n1208 gnd.n1203 59.5399
R15779 gnd.n5607 gnd.n1868 59.5399
R15780 gnd.n6292 gnd.n6291 59.5399
R15781 gnd.n5483 gnd.n5475 59.5399
R15782 gnd.n6289 gnd.n1180 59.1804
R15783 gnd.n4127 gnd.n2649 57.3586
R15784 gnd.n4441 gnd.n2636 57.3586
R15785 gnd.n7549 gnd.n212 57.3586
R15786 gnd.n2929 gnd.t296 56.407
R15787 gnd.n2882 gnd.t326 56.407
R15788 gnd.n2897 gnd.t288 56.407
R15789 gnd.n2913 gnd.t197 56.407
R15790 gnd.n68 gnd.t271 56.407
R15791 gnd.n21 gnd.t206 56.407
R15792 gnd.n36 gnd.t268 56.407
R15793 gnd.n52 gnd.t318 56.407
R15794 gnd.n2942 gnd.t259 55.8337
R15795 gnd.n2895 gnd.t214 55.8337
R15796 gnd.n2910 gnd.t237 55.8337
R15797 gnd.n2926 gnd.t310 55.8337
R15798 gnd.n81 gnd.t322 55.8337
R15799 gnd.n34 gnd.t231 55.8337
R15800 gnd.n49 gnd.t340 55.8337
R15801 gnd.n65 gnd.t236 55.8337
R15802 gnd.n1168 gnd.n1167 54.358
R15803 gnd.n5467 gnd.n5466 54.358
R15804 gnd.n2929 gnd.n2928 53.0052
R15805 gnd.n2931 gnd.n2930 53.0052
R15806 gnd.n2933 gnd.n2932 53.0052
R15807 gnd.n2935 gnd.n2934 53.0052
R15808 gnd.n2937 gnd.n2936 53.0052
R15809 gnd.n2939 gnd.n2938 53.0052
R15810 gnd.n2941 gnd.n2940 53.0052
R15811 gnd.n2882 gnd.n2881 53.0052
R15812 gnd.n2884 gnd.n2883 53.0052
R15813 gnd.n2886 gnd.n2885 53.0052
R15814 gnd.n2888 gnd.n2887 53.0052
R15815 gnd.n2890 gnd.n2889 53.0052
R15816 gnd.n2892 gnd.n2891 53.0052
R15817 gnd.n2894 gnd.n2893 53.0052
R15818 gnd.n2897 gnd.n2896 53.0052
R15819 gnd.n2899 gnd.n2898 53.0052
R15820 gnd.n2901 gnd.n2900 53.0052
R15821 gnd.n2903 gnd.n2902 53.0052
R15822 gnd.n2905 gnd.n2904 53.0052
R15823 gnd.n2907 gnd.n2906 53.0052
R15824 gnd.n2909 gnd.n2908 53.0052
R15825 gnd.n2913 gnd.n2912 53.0052
R15826 gnd.n2915 gnd.n2914 53.0052
R15827 gnd.n2917 gnd.n2916 53.0052
R15828 gnd.n2919 gnd.n2918 53.0052
R15829 gnd.n2921 gnd.n2920 53.0052
R15830 gnd.n2923 gnd.n2922 53.0052
R15831 gnd.n2925 gnd.n2924 53.0052
R15832 gnd.n80 gnd.n79 53.0052
R15833 gnd.n78 gnd.n77 53.0052
R15834 gnd.n76 gnd.n75 53.0052
R15835 gnd.n74 gnd.n73 53.0052
R15836 gnd.n72 gnd.n71 53.0052
R15837 gnd.n70 gnd.n69 53.0052
R15838 gnd.n68 gnd.n67 53.0052
R15839 gnd.n33 gnd.n32 53.0052
R15840 gnd.n31 gnd.n30 53.0052
R15841 gnd.n29 gnd.n28 53.0052
R15842 gnd.n27 gnd.n26 53.0052
R15843 gnd.n25 gnd.n24 53.0052
R15844 gnd.n23 gnd.n22 53.0052
R15845 gnd.n21 gnd.n20 53.0052
R15846 gnd.n48 gnd.n47 53.0052
R15847 gnd.n46 gnd.n45 53.0052
R15848 gnd.n44 gnd.n43 53.0052
R15849 gnd.n42 gnd.n41 53.0052
R15850 gnd.n40 gnd.n39 53.0052
R15851 gnd.n38 gnd.n37 53.0052
R15852 gnd.n36 gnd.n35 53.0052
R15853 gnd.n64 gnd.n63 53.0052
R15854 gnd.n62 gnd.n61 53.0052
R15855 gnd.n60 gnd.n59 53.0052
R15856 gnd.n58 gnd.n57 53.0052
R15857 gnd.n56 gnd.n55 53.0052
R15858 gnd.n54 gnd.n53 53.0052
R15859 gnd.n52 gnd.n51 53.0052
R15860 gnd.n5458 gnd.n5457 52.4801
R15861 gnd.n3979 gnd.t365 52.3082
R15862 gnd.n3947 gnd.t156 52.3082
R15863 gnd.n3915 gnd.t179 52.3082
R15864 gnd.n3884 gnd.t164 52.3082
R15865 gnd.n3852 gnd.t134 52.3082
R15866 gnd.n3820 gnd.t147 52.3082
R15867 gnd.n3788 gnd.t153 52.3082
R15868 gnd.n3757 gnd.t158 52.3082
R15869 gnd.n3809 gnd.n3777 51.4173
R15870 gnd.n3873 gnd.n3872 50.455
R15871 gnd.n3841 gnd.n3840 50.455
R15872 gnd.n3809 gnd.n3808 50.455
R15873 gnd.n3221 gnd.n3220 45.1884
R15874 gnd.n2715 gnd.n2714 45.1884
R15875 gnd.n5542 gnd.n5473 44.3322
R15876 gnd.n1171 gnd.n1170 44.3189
R15877 gnd.n2455 gnd.n2454 42.4732
R15878 gnd.n1459 gnd.n1458 42.4732
R15879 gnd.n6085 gnd.n6084 42.2793
R15880 gnd.n3222 gnd.n3221 42.2793
R15881 gnd.n2716 gnd.n2715 42.2793
R15882 gnd.n3148 gnd.n3147 42.2793
R15883 gnd.n4094 gnd.n2689 42.2793
R15884 gnd.n4796 gnd.n2461 42.2793
R15885 gnd.n6044 gnd.n1530 42.2793
R15886 gnd.n6007 gnd.n1553 42.2793
R15887 gnd.n5967 gnd.n5964 42.2793
R15888 gnd.n315 gnd.n314 42.2793
R15889 gnd.n7477 gnd.n281 42.2793
R15890 gnd.n7514 gnd.n7513 42.2793
R15891 gnd.n7405 gnd.n351 42.2793
R15892 gnd.n4405 gnd.n4186 42.2793
R15893 gnd.n4365 gnd.n4208 42.2793
R15894 gnd.n4326 gnd.n4229 42.2793
R15895 gnd.n4248 gnd.n4247 42.2793
R15896 gnd.n6374 gnd.n1102 42.2793
R15897 gnd.n2280 gnd.n2279 42.2793
R15898 gnd.n2302 gnd.n2301 42.2793
R15899 gnd.n1169 gnd.n1168 41.6274
R15900 gnd.n5468 gnd.n5467 41.6274
R15901 gnd.n1178 gnd.n1177 40.8975
R15902 gnd.n5471 gnd.n5470 40.8975
R15903 gnd.n1177 gnd.n1176 35.055
R15904 gnd.n1172 gnd.n1171 35.055
R15905 gnd.n5460 gnd.n5459 35.055
R15906 gnd.n5470 gnd.n5456 35.055
R15907 gnd.n6652 gnd.n6651 34.6789
R15908 gnd.n6651 gnd.n6650 34.6789
R15909 gnd.n6650 gnd.n772 34.6789
R15910 gnd.n6644 gnd.n772 34.6789
R15911 gnd.n6644 gnd.n6643 34.6789
R15912 gnd.n6643 gnd.n6642 34.6789
R15913 gnd.n6642 gnd.n779 34.6789
R15914 gnd.n6636 gnd.n779 34.6789
R15915 gnd.n6636 gnd.n6635 34.6789
R15916 gnd.n6635 gnd.n6634 34.6789
R15917 gnd.n6634 gnd.n787 34.6789
R15918 gnd.n6628 gnd.n787 34.6789
R15919 gnd.n6628 gnd.n6627 34.6789
R15920 gnd.n6627 gnd.n6626 34.6789
R15921 gnd.n6626 gnd.n795 34.6789
R15922 gnd.n6620 gnd.n795 34.6789
R15923 gnd.n6620 gnd.n6619 34.6789
R15924 gnd.n6619 gnd.n6618 34.6789
R15925 gnd.n6618 gnd.n803 34.6789
R15926 gnd.n6612 gnd.n803 34.6789
R15927 gnd.n6612 gnd.n6611 34.6789
R15928 gnd.n6611 gnd.n6610 34.6789
R15929 gnd.n6610 gnd.n811 34.6789
R15930 gnd.n6604 gnd.n811 34.6789
R15931 gnd.n6604 gnd.n6603 34.6789
R15932 gnd.n6603 gnd.n6602 34.6789
R15933 gnd.n6602 gnd.n819 34.6789
R15934 gnd.n6596 gnd.n819 34.6789
R15935 gnd.n6596 gnd.n6595 34.6789
R15936 gnd.n6595 gnd.n6594 34.6789
R15937 gnd.n6594 gnd.n827 34.6789
R15938 gnd.n6588 gnd.n827 34.6789
R15939 gnd.n6588 gnd.n6587 34.6789
R15940 gnd.n6587 gnd.n6586 34.6789
R15941 gnd.n6586 gnd.n835 34.6789
R15942 gnd.n6580 gnd.n835 34.6789
R15943 gnd.n6580 gnd.n6579 34.6789
R15944 gnd.n6579 gnd.n6578 34.6789
R15945 gnd.n6578 gnd.n843 34.6789
R15946 gnd.n6572 gnd.n843 34.6789
R15947 gnd.n6572 gnd.n6571 34.6789
R15948 gnd.n6571 gnd.n6570 34.6789
R15949 gnd.n6570 gnd.n851 34.6789
R15950 gnd.n6564 gnd.n851 34.6789
R15951 gnd.n6564 gnd.n6563 34.6789
R15952 gnd.n6563 gnd.n6562 34.6789
R15953 gnd.n6562 gnd.n859 34.6789
R15954 gnd.n6556 gnd.n859 34.6789
R15955 gnd.n6556 gnd.n6555 34.6789
R15956 gnd.n6555 gnd.n6554 34.6789
R15957 gnd.n6554 gnd.n867 34.6789
R15958 gnd.n6548 gnd.n867 34.6789
R15959 gnd.n6548 gnd.n6547 34.6789
R15960 gnd.n6547 gnd.n6546 34.6789
R15961 gnd.n6546 gnd.n875 34.6789
R15962 gnd.n6540 gnd.n875 34.6789
R15963 gnd.n6540 gnd.n6539 34.6789
R15964 gnd.n6539 gnd.n6538 34.6789
R15965 gnd.n6538 gnd.n883 34.6789
R15966 gnd.n6532 gnd.n883 34.6789
R15967 gnd.n6532 gnd.n6531 34.6789
R15968 gnd.n6531 gnd.n6530 34.6789
R15969 gnd.n6530 gnd.n891 34.6789
R15970 gnd.n6524 gnd.n891 34.6789
R15971 gnd.n6524 gnd.n6523 34.6789
R15972 gnd.n6523 gnd.n6522 34.6789
R15973 gnd.n6522 gnd.n899 34.6789
R15974 gnd.n6516 gnd.n899 34.6789
R15975 gnd.n6516 gnd.n6515 34.6789
R15976 gnd.n6515 gnd.n6514 34.6789
R15977 gnd.n6514 gnd.n907 34.6789
R15978 gnd.n6508 gnd.n907 34.6789
R15979 gnd.n6508 gnd.n6507 34.6789
R15980 gnd.n6507 gnd.n6506 34.6789
R15981 gnd.n6506 gnd.n915 34.6789
R15982 gnd.n6500 gnd.n915 34.6789
R15983 gnd.n6500 gnd.n6499 34.6789
R15984 gnd.n6499 gnd.n6498 34.6789
R15985 gnd.n6498 gnd.n923 34.6789
R15986 gnd.n6492 gnd.n923 34.6789
R15987 gnd.n6492 gnd.n6491 34.6789
R15988 gnd.n6491 gnd.n6490 34.6789
R15989 gnd.n6490 gnd.n931 34.6789
R15990 gnd.n3284 gnd.n3178 31.8661
R15991 gnd.n3284 gnd.n3283 31.8661
R15992 gnd.n3292 gnd.n3167 31.8661
R15993 gnd.n3300 gnd.n3167 31.8661
R15994 gnd.n3300 gnd.n3161 31.8661
R15995 gnd.n3308 gnd.n3161 31.8661
R15996 gnd.n3308 gnd.n3154 31.8661
R15997 gnd.n3346 gnd.n3154 31.8661
R15998 gnd.n3356 gnd.n3087 31.8661
R15999 gnd.n4451 gnd.n2636 31.8661
R16000 gnd.n4459 gnd.n2628 31.8661
R16001 gnd.n4459 gnd.n2617 31.8661
R16002 gnd.n4471 gnd.n2617 31.8661
R16003 gnd.n4471 gnd.n2620 31.8661
R16004 gnd.n4479 gnd.n2600 31.8661
R16005 gnd.n4491 gnd.n2600 31.8661
R16006 gnd.n4499 gnd.n2592 31.8661
R16007 gnd.n4515 gnd.n2580 31.8661
R16008 gnd.n4515 gnd.n2583 31.8661
R16009 gnd.n4525 gnd.n2566 31.8661
R16010 gnd.n4545 gnd.n2566 31.8661
R16011 gnd.n4556 gnd.n2558 31.8661
R16012 gnd.n4565 gnd.n2540 31.8661
R16013 gnd.n4581 gnd.n2540 31.8661
R16014 gnd.n4585 gnd.n938 31.8661
R16015 gnd.n4741 gnd.n1068 31.8661
R16016 gnd.n4734 gnd.n2203 31.8661
R16017 gnd.n4858 gnd.n2203 31.8661
R16018 gnd.n4866 gnd.n2195 31.8661
R16019 gnd.n4866 gnd.n2197 31.8661
R16020 gnd.n4874 gnd.n2183 31.8661
R16021 gnd.n4882 gnd.n2183 31.8661
R16022 gnd.n4882 gnd.n2176 31.8661
R16023 gnd.n4890 gnd.n2176 31.8661
R16024 gnd.n4898 gnd.n2169 31.8661
R16025 gnd.n4898 gnd.n2161 31.8661
R16026 gnd.n4906 gnd.n2161 31.8661
R16027 gnd.n4906 gnd.n2163 31.8661
R16028 gnd.n4914 gnd.n2147 31.8661
R16029 gnd.n4922 gnd.n2147 31.8661
R16030 gnd.n4922 gnd.n2149 31.8661
R16031 gnd.n4930 gnd.n2132 31.8661
R16032 gnd.n4964 gnd.n2132 31.8661
R16033 gnd.n4964 gnd.n2124 31.8661
R16034 gnd.n4975 gnd.n2124 31.8661
R16035 gnd.n5625 gnd.n1819 31.8661
R16036 gnd.n5634 gnd.n1819 31.8661
R16037 gnd.n5634 gnd.n1813 31.8661
R16038 gnd.n5642 gnd.n1813 31.8661
R16039 gnd.n5651 gnd.n1807 31.8661
R16040 gnd.n5651 gnd.n1801 31.8661
R16041 gnd.n5659 gnd.n1801 31.8661
R16042 gnd.n5668 gnd.n1795 31.8661
R16043 gnd.n5668 gnd.n1788 31.8661
R16044 gnd.n5676 gnd.n1788 31.8661
R16045 gnd.n5676 gnd.n1789 31.8661
R16046 gnd.n5685 gnd.n1777 31.8661
R16047 gnd.n5696 gnd.n1777 31.8661
R16048 gnd.n5696 gnd.n1771 31.8661
R16049 gnd.n5705 gnd.n1771 31.8661
R16050 gnd.n6148 gnd.n1396 31.8661
R16051 gnd.n6148 gnd.n1398 31.8661
R16052 gnd.n5726 gnd.n1764 31.8661
R16053 gnd.n1764 gnd.n1465 31.8661
R16054 gnd.n1575 gnd.n1507 31.8661
R16055 gnd.n7357 gnd.n368 31.8661
R16056 gnd.n7615 gnd.n107 31.8661
R16057 gnd.n7609 gnd.n107 31.8661
R16058 gnd.n7603 gnd.n124 31.8661
R16059 gnd.n7597 gnd.n133 31.8661
R16060 gnd.n7597 gnd.n136 31.8661
R16061 gnd.n7591 gnd.n146 31.8661
R16062 gnd.n7585 gnd.n146 31.8661
R16063 gnd.n7579 gnd.n162 31.8661
R16064 gnd.n7573 gnd.n171 31.8661
R16065 gnd.n7573 gnd.n174 31.8661
R16066 gnd.n7561 gnd.n191 31.8661
R16067 gnd.n7561 gnd.n194 31.8661
R16068 gnd.n7555 gnd.n194 31.8661
R16069 gnd.n7549 gnd.n209 31.8661
R16070 gnd.n5550 gnd.n1869 30.7517
R16071 gnd.n1268 gnd.n1265 30.7517
R16072 gnd.n6355 gnd.n1157 28.9982
R16073 gnd.n5617 gnd.n5615 28.9982
R16074 gnd.n4499 gnd.t190 27.7236
R16075 gnd.n162 gnd.t265 27.7236
R16076 gnd.n2558 gnd.t188 27.0862
R16077 gnd.n2149 gnd.t167 27.0862
R16078 gnd.t6 gnd.n1807 27.0862
R16079 gnd.n124 gnd.t218 27.0862
R16080 gnd.n4600 gnd.t260 26.4489
R16081 gnd.n7308 gnd.t194 26.4489
R16082 gnd.n4556 gnd.t224 25.8116
R16083 gnd.n7603 gnd.t184 25.8116
R16084 gnd.n2454 gnd.n2453 25.7944
R16085 gnd.n6084 gnd.n6083 25.7944
R16086 gnd.n3147 gnd.n3146 25.7944
R16087 gnd.n2689 gnd.n2688 25.7944
R16088 gnd.n2461 gnd.n2460 25.7944
R16089 gnd.n1530 gnd.n1529 25.7944
R16090 gnd.n1553 gnd.n1552 25.7944
R16091 gnd.n5964 gnd.n5963 25.7944
R16092 gnd.n314 gnd.n313 25.7944
R16093 gnd.n281 gnd.n280 25.7944
R16094 gnd.n7513 gnd.n7512 25.7944
R16095 gnd.n351 gnd.n350 25.7944
R16096 gnd.n4186 gnd.n4185 25.7944
R16097 gnd.n4208 gnd.n4207 25.7944
R16098 gnd.n4229 gnd.n4228 25.7944
R16099 gnd.n4247 gnd.n4246 25.7944
R16100 gnd.n1102 gnd.n1101 25.7944
R16101 gnd.n2279 gnd.n2278 25.7944
R16102 gnd.n2301 gnd.n2300 25.7944
R16103 gnd.n1458 gnd.n1457 25.7944
R16104 gnd.t216 gnd.n2592 25.1743
R16105 gnd.n7579 gnd.t207 25.1743
R16106 gnd.n3368 gnd.n3088 24.8557
R16107 gnd.n3378 gnd.n3071 24.8557
R16108 gnd.n3074 gnd.n3062 24.8557
R16109 gnd.n3399 gnd.n3063 24.8557
R16110 gnd.n3409 gnd.n3043 24.8557
R16111 gnd.n3419 gnd.n3418 24.8557
R16112 gnd.n3029 gnd.n3027 24.8557
R16113 gnd.n3450 gnd.n3449 24.8557
R16114 gnd.n3465 gnd.n3012 24.8557
R16115 gnd.n3519 gnd.n2951 24.8557
R16116 gnd.n3475 gnd.n2952 24.8557
R16117 gnd.n3512 gnd.n2963 24.8557
R16118 gnd.n3001 gnd.n3000 24.8557
R16119 gnd.n3506 gnd.n3505 24.8557
R16120 gnd.n2987 gnd.n2974 24.8557
R16121 gnd.n3545 gnd.n3544 24.8557
R16122 gnd.n3555 gnd.n2867 24.8557
R16123 gnd.n3567 gnd.n2859 24.8557
R16124 gnd.n3566 gnd.n2847 24.8557
R16125 gnd.n3585 gnd.n3584 24.8557
R16126 gnd.n3595 gnd.n2840 24.8557
R16127 gnd.n3606 gnd.n2828 24.8557
R16128 gnd.n3630 gnd.n3629 24.8557
R16129 gnd.n3641 gnd.n2811 24.8557
R16130 gnd.n3640 gnd.n2813 24.8557
R16131 gnd.n3652 gnd.n2804 24.8557
R16132 gnd.n3670 gnd.n3669 24.8557
R16133 gnd.n2795 gnd.n2784 24.8557
R16134 gnd.n3691 gnd.n2772 24.8557
R16135 gnd.n3719 gnd.n3718 24.8557
R16136 gnd.n3730 gnd.n2757 24.8557
R16137 gnd.n3742 gnd.n2750 24.8557
R16138 gnd.n4014 gnd.n4013 24.8557
R16139 gnd.n4036 gnd.n2723 24.8557
R16140 gnd.n2197 gnd.t59 24.537
R16141 gnd.n4914 gnd.t358 24.537
R16142 gnd.n5659 gnd.t368 24.537
R16143 gnd.t26 gnd.n1396 24.537
R16144 gnd.n4857 gnd.n2195 23.8997
R16145 gnd.n5727 gnd.n1398 23.8997
R16146 gnd.n3389 gnd.t157 23.2624
R16147 gnd.n7567 gnd.n184 23.2624
R16148 gnd.n3090 gnd.t48 22.6251
R16149 gnd.n4451 gnd.t22 22.6251
R16150 gnd.n209 gnd.t37 22.6251
R16151 gnd.n6285 gnd.n1183 21.6691
R16152 gnd.n6278 gnd.n1196 21.6691
R16153 gnd.n5029 gnd.n5028 21.6691
R16154 gnd.n5045 gnd.n2095 21.6691
R16155 gnd.n5051 gnd.n2078 21.6691
R16156 gnd.n5056 gnd.n2071 21.6691
R16157 gnd.n5115 gnd.n2063 21.6691
R16158 gnd.n5126 gnd.n2058 21.6691
R16159 gnd.n5207 gnd.n2005 21.6691
R16160 gnd.n5301 gnd.n1958 21.6691
R16161 gnd.n5322 gnd.n5321 21.6691
R16162 gnd.n5341 gnd.n1941 21.6691
R16163 gnd.n5347 gnd.n1937 21.6691
R16164 gnd.n5365 gnd.n1920 21.6691
R16165 gnd.n5392 gnd.n1907 21.6691
R16166 gnd.n5451 gnd.n1877 21.6691
R16167 gnd.t163 gnd.n3095 21.3504
R16168 gnd.n6266 gnd.t66 21.0318
R16169 gnd.n3740 gnd.n931 20.8076
R16170 gnd.t352 gnd.n2785 20.7131
R16171 gnd.n6284 gnd.n1186 20.3945
R16172 gnd.n6272 gnd.n1276 20.3945
R16173 gnd.n5433 gnd.n1886 20.3945
R16174 gnd.n1880 gnd.n1872 20.3945
R16175 gnd.t354 gnd.n2820 20.0758
R16176 gnd.n5011 gnd.t169 20.0758
R16177 gnd.t370 gnd.n1899 20.0758
R16178 gnd.n1203 gnd.n1202 19.9763
R16179 gnd.n1868 gnd.n1867 19.9763
R16180 gnd.n6291 gnd.n6290 19.9763
R16181 gnd.n5475 gnd.n5474 19.9763
R16182 gnd.n1166 gnd.t117 19.8005
R16183 gnd.n1166 gnd.t130 19.8005
R16184 gnd.n1165 gnd.t67 19.8005
R16185 gnd.n1165 gnd.t20 19.8005
R16186 gnd.n5465 gnd.t35 19.8005
R16187 gnd.n5465 gnd.t79 19.8005
R16188 gnd.n5464 gnd.t53 19.8005
R16189 gnd.n5464 gnd.t92 19.8005
R16190 gnd.n4734 gnd.n1073 19.7572
R16191 gnd.n6080 gnd.n1465 19.7572
R16192 gnd.n1162 gnd.n1161 19.5087
R16193 gnd.n1175 gnd.n1162 19.5087
R16194 gnd.n1173 gnd.n1164 19.5087
R16195 gnd.n5469 gnd.n5463 19.5087
R16196 gnd.n3556 gnd.t342 19.4385
R16197 gnd.n4890 gnd.t0 19.4385
R16198 gnd.n5685 gnd.t171 19.4385
R16199 gnd.n4868 gnd.n2192 19.3944
R16200 gnd.n4872 gnd.n2192 19.3944
R16201 gnd.n4872 gnd.n2181 19.3944
R16202 gnd.n4884 gnd.n2181 19.3944
R16203 gnd.n4884 gnd.n2179 19.3944
R16204 gnd.n4888 gnd.n2179 19.3944
R16205 gnd.n4888 gnd.n2167 19.3944
R16206 gnd.n4900 gnd.n2167 19.3944
R16207 gnd.n4900 gnd.n2165 19.3944
R16208 gnd.n4904 gnd.n2165 19.3944
R16209 gnd.n4904 gnd.n2153 19.3944
R16210 gnd.n4916 gnd.n2153 19.3944
R16211 gnd.n4916 gnd.n2151 19.3944
R16212 gnd.n4920 gnd.n2151 19.3944
R16213 gnd.n4920 gnd.n2139 19.3944
R16214 gnd.n4932 gnd.n2139 19.3944
R16215 gnd.n4932 gnd.n2136 19.3944
R16216 gnd.n4962 gnd.n2136 19.3944
R16217 gnd.n4962 gnd.n2137 19.3944
R16218 gnd.n4958 gnd.n2137 19.3944
R16219 gnd.n4958 gnd.n4957 19.3944
R16220 gnd.n4957 gnd.n4956 19.3944
R16221 gnd.n4956 gnd.n4938 19.3944
R16222 gnd.n4952 gnd.n4938 19.3944
R16223 gnd.n4952 gnd.n4951 19.3944
R16224 gnd.n4951 gnd.n4950 19.3944
R16225 gnd.n4950 gnd.n4945 19.3944
R16226 gnd.n4946 gnd.n4945 19.3944
R16227 gnd.n4946 gnd.n1305 19.3944
R16228 gnd.n6257 gnd.n1305 19.3944
R16229 gnd.n6257 gnd.n1306 19.3944
R16230 gnd.n6253 gnd.n1306 19.3944
R16231 gnd.n6253 gnd.n6252 19.3944
R16232 gnd.n6252 gnd.n6251 19.3944
R16233 gnd.n6251 gnd.n1312 19.3944
R16234 gnd.n6247 gnd.n1312 19.3944
R16235 gnd.n6247 gnd.n6246 19.3944
R16236 gnd.n6246 gnd.n6245 19.3944
R16237 gnd.n6245 gnd.n1317 19.3944
R16238 gnd.n6241 gnd.n1317 19.3944
R16239 gnd.n6241 gnd.n6240 19.3944
R16240 gnd.n6240 gnd.n6239 19.3944
R16241 gnd.n6239 gnd.n1322 19.3944
R16242 gnd.n6235 gnd.n1322 19.3944
R16243 gnd.n6235 gnd.n6234 19.3944
R16244 gnd.n6234 gnd.n6233 19.3944
R16245 gnd.n6233 gnd.n1327 19.3944
R16246 gnd.n6229 gnd.n1327 19.3944
R16247 gnd.n6229 gnd.n6228 19.3944
R16248 gnd.n6228 gnd.n6227 19.3944
R16249 gnd.n6227 gnd.n1332 19.3944
R16250 gnd.n6223 gnd.n1332 19.3944
R16251 gnd.n6223 gnd.n6222 19.3944
R16252 gnd.n6222 gnd.n6221 19.3944
R16253 gnd.n6221 gnd.n1337 19.3944
R16254 gnd.n6217 gnd.n1337 19.3944
R16255 gnd.n6217 gnd.n6216 19.3944
R16256 gnd.n6216 gnd.n6215 19.3944
R16257 gnd.n6215 gnd.n1342 19.3944
R16258 gnd.n6211 gnd.n1342 19.3944
R16259 gnd.n6211 gnd.n6210 19.3944
R16260 gnd.n6210 gnd.n6209 19.3944
R16261 gnd.n6209 gnd.n1347 19.3944
R16262 gnd.n6205 gnd.n1347 19.3944
R16263 gnd.n6205 gnd.n6204 19.3944
R16264 gnd.n6204 gnd.n6203 19.3944
R16265 gnd.n6203 gnd.n1352 19.3944
R16266 gnd.n6199 gnd.n1352 19.3944
R16267 gnd.n6199 gnd.n6198 19.3944
R16268 gnd.n6198 gnd.n6197 19.3944
R16269 gnd.n6197 gnd.n1357 19.3944
R16270 gnd.n6193 gnd.n1357 19.3944
R16271 gnd.n6193 gnd.n6192 19.3944
R16272 gnd.n6192 gnd.n6191 19.3944
R16273 gnd.n6191 gnd.n1362 19.3944
R16274 gnd.n6187 gnd.n1362 19.3944
R16275 gnd.n6187 gnd.n6186 19.3944
R16276 gnd.n6186 gnd.n6185 19.3944
R16277 gnd.n6185 gnd.n1367 19.3944
R16278 gnd.n6181 gnd.n1367 19.3944
R16279 gnd.n6181 gnd.n6180 19.3944
R16280 gnd.n6180 gnd.n6179 19.3944
R16281 gnd.n6179 gnd.n1372 19.3944
R16282 gnd.n6175 gnd.n1372 19.3944
R16283 gnd.n6175 gnd.n6174 19.3944
R16284 gnd.n6174 gnd.n6173 19.3944
R16285 gnd.n6173 gnd.n1377 19.3944
R16286 gnd.n6169 gnd.n1377 19.3944
R16287 gnd.n6169 gnd.n6168 19.3944
R16288 gnd.n6168 gnd.n6167 19.3944
R16289 gnd.n6167 gnd.n1382 19.3944
R16290 gnd.n6163 gnd.n1382 19.3944
R16291 gnd.n6163 gnd.n6162 19.3944
R16292 gnd.n6162 gnd.n6161 19.3944
R16293 gnd.n6161 gnd.n1387 19.3944
R16294 gnd.n6157 gnd.n1387 19.3944
R16295 gnd.n6157 gnd.n6156 19.3944
R16296 gnd.n6156 gnd.n6155 19.3944
R16297 gnd.n6155 gnd.n1392 19.3944
R16298 gnd.n6151 gnd.n1392 19.3944
R16299 gnd.n6151 gnd.n6150 19.3944
R16300 gnd.n4786 gnd.n4785 19.3944
R16301 gnd.n4790 gnd.n4786 19.3944
R16302 gnd.n4790 gnd.n4789 19.3944
R16303 gnd.n4854 gnd.n4853 19.3944
R16304 gnd.n4853 gnd.n2271 19.3944
R16305 gnd.n4849 gnd.n2271 19.3944
R16306 gnd.n4849 gnd.n4848 19.3944
R16307 gnd.n4848 gnd.n4847 19.3944
R16308 gnd.n4847 gnd.n2276 19.3944
R16309 gnd.n4842 gnd.n2276 19.3944
R16310 gnd.n4842 gnd.n4841 19.3944
R16311 gnd.n4841 gnd.n4840 19.3944
R16312 gnd.n4840 gnd.n2395 19.3944
R16313 gnd.n4833 gnd.n2395 19.3944
R16314 gnd.n4833 gnd.n4832 19.3944
R16315 gnd.n4832 gnd.n2408 19.3944
R16316 gnd.n4825 gnd.n2408 19.3944
R16317 gnd.n4825 gnd.n4824 19.3944
R16318 gnd.n4824 gnd.n2418 19.3944
R16319 gnd.n4817 gnd.n2418 19.3944
R16320 gnd.n4817 gnd.n4816 19.3944
R16321 gnd.n4816 gnd.n2431 19.3944
R16322 gnd.n4809 gnd.n2431 19.3944
R16323 gnd.n4809 gnd.n4808 19.3944
R16324 gnd.n4808 gnd.n2441 19.3944
R16325 gnd.n4801 gnd.n2441 19.3944
R16326 gnd.n4801 gnd.n4800 19.3944
R16327 gnd.n6126 gnd.n1418 19.3944
R16328 gnd.n6126 gnd.n6125 19.3944
R16329 gnd.n6125 gnd.n1421 19.3944
R16330 gnd.n6118 gnd.n1421 19.3944
R16331 gnd.n6118 gnd.n6117 19.3944
R16332 gnd.n6117 gnd.n1429 19.3944
R16333 gnd.n6110 gnd.n1429 19.3944
R16334 gnd.n6110 gnd.n6109 19.3944
R16335 gnd.n6109 gnd.n1437 19.3944
R16336 gnd.n6102 gnd.n1437 19.3944
R16337 gnd.n6102 gnd.n6101 19.3944
R16338 gnd.n6101 gnd.n1445 19.3944
R16339 gnd.n6094 gnd.n1445 19.3944
R16340 gnd.n6094 gnd.n6093 19.3944
R16341 gnd.n6093 gnd.n1453 19.3944
R16342 gnd.n6086 gnd.n1453 19.3944
R16343 gnd.n3271 gnd.n3270 19.3944
R16344 gnd.n3270 gnd.n3269 19.3944
R16345 gnd.n3269 gnd.n3268 19.3944
R16346 gnd.n3268 gnd.n3266 19.3944
R16347 gnd.n3266 gnd.n3263 19.3944
R16348 gnd.n3263 gnd.n3262 19.3944
R16349 gnd.n3262 gnd.n3259 19.3944
R16350 gnd.n3259 gnd.n3258 19.3944
R16351 gnd.n3258 gnd.n3255 19.3944
R16352 gnd.n3255 gnd.n3254 19.3944
R16353 gnd.n3254 gnd.n3251 19.3944
R16354 gnd.n3251 gnd.n3250 19.3944
R16355 gnd.n3250 gnd.n3247 19.3944
R16356 gnd.n3247 gnd.n3246 19.3944
R16357 gnd.n3246 gnd.n3243 19.3944
R16358 gnd.n3243 gnd.n3242 19.3944
R16359 gnd.n3242 gnd.n3239 19.3944
R16360 gnd.n3239 gnd.n3238 19.3944
R16361 gnd.n3238 gnd.n3235 19.3944
R16362 gnd.n3235 gnd.n3234 19.3944
R16363 gnd.n3234 gnd.n3231 19.3944
R16364 gnd.n3231 gnd.n3230 19.3944
R16365 gnd.n3227 gnd.n3226 19.3944
R16366 gnd.n3226 gnd.n3182 19.3944
R16367 gnd.n3277 gnd.n3182 19.3944
R16368 gnd.n4044 gnd.n4043 19.3944
R16369 gnd.n4043 gnd.n4040 19.3944
R16370 gnd.n4040 gnd.n4039 19.3944
R16371 gnd.n4089 gnd.n4088 19.3944
R16372 gnd.n4088 gnd.n4087 19.3944
R16373 gnd.n4087 gnd.n4084 19.3944
R16374 gnd.n4084 gnd.n4083 19.3944
R16375 gnd.n4083 gnd.n4080 19.3944
R16376 gnd.n4080 gnd.n4079 19.3944
R16377 gnd.n4079 gnd.n4076 19.3944
R16378 gnd.n4076 gnd.n4075 19.3944
R16379 gnd.n4075 gnd.n4072 19.3944
R16380 gnd.n4072 gnd.n4071 19.3944
R16381 gnd.n4071 gnd.n4068 19.3944
R16382 gnd.n4068 gnd.n4067 19.3944
R16383 gnd.n4067 gnd.n4064 19.3944
R16384 gnd.n4064 gnd.n4063 19.3944
R16385 gnd.n4063 gnd.n4060 19.3944
R16386 gnd.n4060 gnd.n4059 19.3944
R16387 gnd.n4059 gnd.n4056 19.3944
R16388 gnd.n4056 gnd.n4055 19.3944
R16389 gnd.n4055 gnd.n4052 19.3944
R16390 gnd.n4052 gnd.n4051 19.3944
R16391 gnd.n4051 gnd.n4048 19.3944
R16392 gnd.n4048 gnd.n4047 19.3944
R16393 gnd.n3370 gnd.n3079 19.3944
R16394 gnd.n3380 gnd.n3079 19.3944
R16395 gnd.n3381 gnd.n3380 19.3944
R16396 gnd.n3381 gnd.n3060 19.3944
R16397 gnd.n3401 gnd.n3060 19.3944
R16398 gnd.n3401 gnd.n3052 19.3944
R16399 gnd.n3411 gnd.n3052 19.3944
R16400 gnd.n3412 gnd.n3411 19.3944
R16401 gnd.n3413 gnd.n3412 19.3944
R16402 gnd.n3413 gnd.n3035 19.3944
R16403 gnd.n3430 gnd.n3035 19.3944
R16404 gnd.n3433 gnd.n3430 19.3944
R16405 gnd.n3433 gnd.n3432 19.3944
R16406 gnd.n3432 gnd.n3008 19.3944
R16407 gnd.n3472 gnd.n3008 19.3944
R16408 gnd.n3472 gnd.n3005 19.3944
R16409 gnd.n3478 gnd.n3005 19.3944
R16410 gnd.n3479 gnd.n3478 19.3944
R16411 gnd.n3479 gnd.n3003 19.3944
R16412 gnd.n3485 gnd.n3003 19.3944
R16413 gnd.n3488 gnd.n3485 19.3944
R16414 gnd.n3490 gnd.n3488 19.3944
R16415 gnd.n3496 gnd.n3490 19.3944
R16416 gnd.n3496 gnd.n3495 19.3944
R16417 gnd.n3495 gnd.n2862 19.3944
R16418 gnd.n3562 gnd.n2862 19.3944
R16419 gnd.n3563 gnd.n3562 19.3944
R16420 gnd.n3563 gnd.n2855 19.3944
R16421 gnd.n3574 gnd.n2855 19.3944
R16422 gnd.n3575 gnd.n3574 19.3944
R16423 gnd.n3575 gnd.n2838 19.3944
R16424 gnd.n2838 gnd.n2836 19.3944
R16425 gnd.n3599 gnd.n2836 19.3944
R16426 gnd.n3600 gnd.n3599 19.3944
R16427 gnd.n3600 gnd.n2807 19.3944
R16428 gnd.n3647 gnd.n2807 19.3944
R16429 gnd.n3648 gnd.n3647 19.3944
R16430 gnd.n3648 gnd.n2800 19.3944
R16431 gnd.n3659 gnd.n2800 19.3944
R16432 gnd.n3660 gnd.n3659 19.3944
R16433 gnd.n3660 gnd.n2783 19.3944
R16434 gnd.n2783 gnd.n2781 19.3944
R16435 gnd.n3684 gnd.n2781 19.3944
R16436 gnd.n3685 gnd.n3684 19.3944
R16437 gnd.n3685 gnd.n2753 19.3944
R16438 gnd.n3736 gnd.n2753 19.3944
R16439 gnd.n3737 gnd.n3736 19.3944
R16440 gnd.n3737 gnd.n2746 19.3944
R16441 gnd.n4005 gnd.n2746 19.3944
R16442 gnd.n4006 gnd.n4005 19.3944
R16443 gnd.n4006 gnd.n2727 19.3944
R16444 gnd.n4031 gnd.n2727 19.3944
R16445 gnd.n4031 gnd.n2728 19.3944
R16446 gnd.n3361 gnd.n3360 19.3944
R16447 gnd.n3360 gnd.n3093 19.3944
R16448 gnd.n3116 gnd.n3093 19.3944
R16449 gnd.n3119 gnd.n3116 19.3944
R16450 gnd.n3119 gnd.n3112 19.3944
R16451 gnd.n3123 gnd.n3112 19.3944
R16452 gnd.n3126 gnd.n3123 19.3944
R16453 gnd.n3129 gnd.n3126 19.3944
R16454 gnd.n3129 gnd.n3110 19.3944
R16455 gnd.n3133 gnd.n3110 19.3944
R16456 gnd.n3136 gnd.n3133 19.3944
R16457 gnd.n3139 gnd.n3136 19.3944
R16458 gnd.n3139 gnd.n3108 19.3944
R16459 gnd.n3143 gnd.n3108 19.3944
R16460 gnd.n3366 gnd.n3365 19.3944
R16461 gnd.n3365 gnd.n3069 19.3944
R16462 gnd.n3391 gnd.n3069 19.3944
R16463 gnd.n3391 gnd.n3067 19.3944
R16464 gnd.n3397 gnd.n3067 19.3944
R16465 gnd.n3397 gnd.n3396 19.3944
R16466 gnd.n3396 gnd.n3041 19.3944
R16467 gnd.n3421 gnd.n3041 19.3944
R16468 gnd.n3421 gnd.n3039 19.3944
R16469 gnd.n3425 gnd.n3039 19.3944
R16470 gnd.n3425 gnd.n3019 19.3944
R16471 gnd.n3452 gnd.n3019 19.3944
R16472 gnd.n3452 gnd.n3017 19.3944
R16473 gnd.n3462 gnd.n3017 19.3944
R16474 gnd.n3462 gnd.n3461 19.3944
R16475 gnd.n3461 gnd.n3460 19.3944
R16476 gnd.n3460 gnd.n2966 19.3944
R16477 gnd.n3510 gnd.n2966 19.3944
R16478 gnd.n3510 gnd.n3509 19.3944
R16479 gnd.n3509 gnd.n3508 19.3944
R16480 gnd.n3508 gnd.n2970 19.3944
R16481 gnd.n2990 gnd.n2970 19.3944
R16482 gnd.n2990 gnd.n2872 19.3944
R16483 gnd.n3547 gnd.n2872 19.3944
R16484 gnd.n3547 gnd.n2870 19.3944
R16485 gnd.n3553 gnd.n2870 19.3944
R16486 gnd.n3553 gnd.n3552 19.3944
R16487 gnd.n3552 gnd.n2845 19.3944
R16488 gnd.n3587 gnd.n2845 19.3944
R16489 gnd.n3587 gnd.n2843 19.3944
R16490 gnd.n3593 gnd.n2843 19.3944
R16491 gnd.n3593 gnd.n3592 19.3944
R16492 gnd.n3592 gnd.n2818 19.3944
R16493 gnd.n3632 gnd.n2818 19.3944
R16494 gnd.n3632 gnd.n2816 19.3944
R16495 gnd.n3638 gnd.n2816 19.3944
R16496 gnd.n3638 gnd.n3637 19.3944
R16497 gnd.n3637 gnd.n2790 19.3944
R16498 gnd.n3672 gnd.n2790 19.3944
R16499 gnd.n3672 gnd.n2788 19.3944
R16500 gnd.n3678 gnd.n2788 19.3944
R16501 gnd.n3678 gnd.n3677 19.3944
R16502 gnd.n3677 gnd.n2763 19.3944
R16503 gnd.n3721 gnd.n2763 19.3944
R16504 gnd.n3721 gnd.n2761 19.3944
R16505 gnd.n3727 gnd.n2761 19.3944
R16506 gnd.n3727 gnd.n3726 19.3944
R16507 gnd.n3726 gnd.n2736 19.3944
R16508 gnd.n4016 gnd.n2736 19.3944
R16509 gnd.n4016 gnd.n2734 19.3944
R16510 gnd.n4024 gnd.n2734 19.3944
R16511 gnd.n4024 gnd.n4023 19.3944
R16512 gnd.n4023 gnd.n4022 19.3944
R16513 gnd.n4125 gnd.n4124 19.3944
R16514 gnd.n4124 gnd.n2675 19.3944
R16515 gnd.n4120 gnd.n2675 19.3944
R16516 gnd.n4120 gnd.n4117 19.3944
R16517 gnd.n4117 gnd.n4114 19.3944
R16518 gnd.n4114 gnd.n4113 19.3944
R16519 gnd.n4113 gnd.n4110 19.3944
R16520 gnd.n4110 gnd.n4109 19.3944
R16521 gnd.n4109 gnd.n4106 19.3944
R16522 gnd.n4106 gnd.n4105 19.3944
R16523 gnd.n4105 gnd.n4102 19.3944
R16524 gnd.n4102 gnd.n4101 19.3944
R16525 gnd.n4101 gnd.n4098 19.3944
R16526 gnd.n4098 gnd.n4097 19.3944
R16527 gnd.n3281 gnd.n3180 19.3944
R16528 gnd.n3281 gnd.n3171 19.3944
R16529 gnd.n3294 gnd.n3171 19.3944
R16530 gnd.n3294 gnd.n3169 19.3944
R16531 gnd.n3298 gnd.n3169 19.3944
R16532 gnd.n3298 gnd.n3159 19.3944
R16533 gnd.n3310 gnd.n3159 19.3944
R16534 gnd.n3310 gnd.n3157 19.3944
R16535 gnd.n3344 gnd.n3157 19.3944
R16536 gnd.n3344 gnd.n3343 19.3944
R16537 gnd.n3343 gnd.n3342 19.3944
R16538 gnd.n3342 gnd.n3341 19.3944
R16539 gnd.n3341 gnd.n3338 19.3944
R16540 gnd.n3338 gnd.n3337 19.3944
R16541 gnd.n3337 gnd.n3336 19.3944
R16542 gnd.n3336 gnd.n3334 19.3944
R16543 gnd.n3334 gnd.n3333 19.3944
R16544 gnd.n3333 gnd.n3330 19.3944
R16545 gnd.n3330 gnd.n3329 19.3944
R16546 gnd.n3329 gnd.n3328 19.3944
R16547 gnd.n3328 gnd.n3326 19.3944
R16548 gnd.n3326 gnd.n3025 19.3944
R16549 gnd.n3441 gnd.n3025 19.3944
R16550 gnd.n3441 gnd.n3023 19.3944
R16551 gnd.n3447 gnd.n3023 19.3944
R16552 gnd.n3447 gnd.n3446 19.3944
R16553 gnd.n3446 gnd.n2947 19.3944
R16554 gnd.n3521 gnd.n2947 19.3944
R16555 gnd.n3521 gnd.n2948 19.3944
R16556 gnd.n2995 gnd.n2994 19.3944
R16557 gnd.n2998 gnd.n2997 19.3944
R16558 gnd.n2985 gnd.n2984 19.3944
R16559 gnd.n3540 gnd.n2877 19.3944
R16560 gnd.n3540 gnd.n3539 19.3944
R16561 gnd.n3539 gnd.n3538 19.3944
R16562 gnd.n3538 gnd.n3536 19.3944
R16563 gnd.n3536 gnd.n3535 19.3944
R16564 gnd.n3535 gnd.n3533 19.3944
R16565 gnd.n3533 gnd.n3532 19.3944
R16566 gnd.n3532 gnd.n2826 19.3944
R16567 gnd.n3608 gnd.n2826 19.3944
R16568 gnd.n3608 gnd.n2824 19.3944
R16569 gnd.n3627 gnd.n2824 19.3944
R16570 gnd.n3627 gnd.n3626 19.3944
R16571 gnd.n3626 gnd.n3625 19.3944
R16572 gnd.n3625 gnd.n3623 19.3944
R16573 gnd.n3623 gnd.n3622 19.3944
R16574 gnd.n3622 gnd.n3620 19.3944
R16575 gnd.n3620 gnd.n3619 19.3944
R16576 gnd.n3619 gnd.n2770 19.3944
R16577 gnd.n3693 gnd.n2770 19.3944
R16578 gnd.n3693 gnd.n2768 19.3944
R16579 gnd.n3716 gnd.n2768 19.3944
R16580 gnd.n3716 gnd.n3715 19.3944
R16581 gnd.n3715 gnd.n3714 19.3944
R16582 gnd.n3714 gnd.n3711 19.3944
R16583 gnd.n3711 gnd.n3710 19.3944
R16584 gnd.n3710 gnd.n3708 19.3944
R16585 gnd.n3708 gnd.n3707 19.3944
R16586 gnd.n3707 gnd.n3705 19.3944
R16587 gnd.n3705 gnd.n2722 19.3944
R16588 gnd.n3286 gnd.n3176 19.3944
R16589 gnd.n3286 gnd.n3174 19.3944
R16590 gnd.n3290 gnd.n3174 19.3944
R16591 gnd.n3290 gnd.n3165 19.3944
R16592 gnd.n3302 gnd.n3165 19.3944
R16593 gnd.n3302 gnd.n3163 19.3944
R16594 gnd.n3306 gnd.n3163 19.3944
R16595 gnd.n3306 gnd.n3152 19.3944
R16596 gnd.n3348 gnd.n3152 19.3944
R16597 gnd.n3348 gnd.n3106 19.3944
R16598 gnd.n3354 gnd.n3106 19.3944
R16599 gnd.n3354 gnd.n3353 19.3944
R16600 gnd.n3353 gnd.n3084 19.3944
R16601 gnd.n3375 gnd.n3084 19.3944
R16602 gnd.n3375 gnd.n3077 19.3944
R16603 gnd.n3386 gnd.n3077 19.3944
R16604 gnd.n3386 gnd.n3385 19.3944
R16605 gnd.n3385 gnd.n3058 19.3944
R16606 gnd.n3406 gnd.n3058 19.3944
R16607 gnd.n3406 gnd.n3048 19.3944
R16608 gnd.n3416 gnd.n3048 19.3944
R16609 gnd.n3416 gnd.n3031 19.3944
R16610 gnd.n3437 gnd.n3031 19.3944
R16611 gnd.n3437 gnd.n3436 19.3944
R16612 gnd.n3436 gnd.n3010 19.3944
R16613 gnd.n3467 gnd.n3010 19.3944
R16614 gnd.n3467 gnd.n2955 19.3944
R16615 gnd.n3517 gnd.n2955 19.3944
R16616 gnd.n3517 gnd.n3516 19.3944
R16617 gnd.n3516 gnd.n3515 19.3944
R16618 gnd.n3515 gnd.n2959 19.3944
R16619 gnd.n2977 gnd.n2959 19.3944
R16620 gnd.n3503 gnd.n2977 19.3944
R16621 gnd.n3503 gnd.n3502 19.3944
R16622 gnd.n3502 gnd.n3501 19.3944
R16623 gnd.n3501 gnd.n2981 19.3944
R16624 gnd.n2981 gnd.n2864 19.3944
R16625 gnd.n3558 gnd.n2864 19.3944
R16626 gnd.n3558 gnd.n2857 19.3944
R16627 gnd.n3569 gnd.n2857 19.3944
R16628 gnd.n3569 gnd.n2853 19.3944
R16629 gnd.n3582 gnd.n2853 19.3944
R16630 gnd.n3582 gnd.n3581 19.3944
R16631 gnd.n3581 gnd.n2832 19.3944
R16632 gnd.n3604 gnd.n2832 19.3944
R16633 gnd.n3604 gnd.n3603 19.3944
R16634 gnd.n3603 gnd.n2809 19.3944
R16635 gnd.n3643 gnd.n2809 19.3944
R16636 gnd.n3643 gnd.n2802 19.3944
R16637 gnd.n3654 gnd.n2802 19.3944
R16638 gnd.n3654 gnd.n2798 19.3944
R16639 gnd.n3667 gnd.n2798 19.3944
R16640 gnd.n3667 gnd.n3666 19.3944
R16641 gnd.n3666 gnd.n2777 19.3944
R16642 gnd.n3689 gnd.n2777 19.3944
R16643 gnd.n3689 gnd.n3688 19.3944
R16644 gnd.n3688 gnd.n2755 19.3944
R16645 gnd.n3732 gnd.n2755 19.3944
R16646 gnd.n3732 gnd.n2748 19.3944
R16647 gnd.n3744 gnd.n2748 19.3944
R16648 gnd.n3744 gnd.n2744 19.3944
R16649 gnd.n4011 gnd.n2744 19.3944
R16650 gnd.n4011 gnd.n4010 19.3944
R16651 gnd.n4010 gnd.n2725 19.3944
R16652 gnd.n4034 gnd.n2725 19.3944
R16653 gnd.n4837 gnd.n2398 19.3944
R16654 gnd.n4837 gnd.n4836 19.3944
R16655 gnd.n4836 gnd.n2402 19.3944
R16656 gnd.n4829 gnd.n2402 19.3944
R16657 gnd.n4829 gnd.n4828 19.3944
R16658 gnd.n4828 gnd.n2414 19.3944
R16659 gnd.n4821 gnd.n2414 19.3944
R16660 gnd.n4821 gnd.n4820 19.3944
R16661 gnd.n4820 gnd.n2425 19.3944
R16662 gnd.n4813 gnd.n2425 19.3944
R16663 gnd.n4813 gnd.n4812 19.3944
R16664 gnd.n4812 gnd.n2437 19.3944
R16665 gnd.n4805 gnd.n2437 19.3944
R16666 gnd.n4805 gnd.n4804 19.3944
R16667 gnd.n4804 gnd.n2448 19.3944
R16668 gnd.n4797 gnd.n2448 19.3944
R16669 gnd.n2514 gnd.n2511 19.3944
R16670 gnd.n4622 gnd.n2514 19.3944
R16671 gnd.n4622 gnd.n2510 19.3944
R16672 gnd.n4646 gnd.n2510 19.3944
R16673 gnd.n4646 gnd.n4645 19.3944
R16674 gnd.n4645 gnd.n4644 19.3944
R16675 gnd.n4644 gnd.n4628 19.3944
R16676 gnd.n4640 gnd.n4628 19.3944
R16677 gnd.n4640 gnd.n4639 19.3944
R16678 gnd.n4639 gnd.n4638 19.3944
R16679 gnd.n4638 gnd.n4636 19.3944
R16680 gnd.n4636 gnd.n2486 19.3944
R16681 gnd.n2486 gnd.n2484 19.3944
R16682 gnd.n4713 gnd.n2484 19.3944
R16683 gnd.n4713 gnd.n2482 19.3944
R16684 gnd.n4717 gnd.n2482 19.3944
R16685 gnd.n4717 gnd.n2480 19.3944
R16686 gnd.n4721 gnd.n2480 19.3944
R16687 gnd.n4721 gnd.n2478 19.3944
R16688 gnd.n4753 gnd.n2478 19.3944
R16689 gnd.n4753 gnd.n4752 19.3944
R16690 gnd.n4752 gnd.n4751 19.3944
R16691 gnd.n4751 gnd.n4727 19.3944
R16692 gnd.n4747 gnd.n4727 19.3944
R16693 gnd.n4747 gnd.n4746 19.3944
R16694 gnd.n4746 gnd.n4745 19.3944
R16695 gnd.n4745 gnd.n4733 19.3944
R16696 gnd.n4740 gnd.n4733 19.3944
R16697 gnd.n4740 gnd.n4739 19.3944
R16698 gnd.n4739 gnd.n2201 19.3944
R16699 gnd.n4860 gnd.n2201 19.3944
R16700 gnd.n4860 gnd.n2199 19.3944
R16701 gnd.n4864 gnd.n2199 19.3944
R16702 gnd.n4864 gnd.n2188 19.3944
R16703 gnd.n4876 gnd.n2188 19.3944
R16704 gnd.n4876 gnd.n2186 19.3944
R16705 gnd.n4880 gnd.n2186 19.3944
R16706 gnd.n4880 gnd.n2174 19.3944
R16707 gnd.n4892 gnd.n2174 19.3944
R16708 gnd.n4892 gnd.n2172 19.3944
R16709 gnd.n4896 gnd.n2172 19.3944
R16710 gnd.n4896 gnd.n2159 19.3944
R16711 gnd.n4908 gnd.n2159 19.3944
R16712 gnd.n4908 gnd.n2157 19.3944
R16713 gnd.n4912 gnd.n2157 19.3944
R16714 gnd.n4912 gnd.n2145 19.3944
R16715 gnd.n4924 gnd.n2145 19.3944
R16716 gnd.n4924 gnd.n2143 19.3944
R16717 gnd.n4928 gnd.n2143 19.3944
R16718 gnd.n4928 gnd.n2130 19.3944
R16719 gnd.n4966 gnd.n2130 19.3944
R16720 gnd.n4966 gnd.n2128 19.3944
R16721 gnd.n4973 gnd.n2128 19.3944
R16722 gnd.n4973 gnd.n4972 19.3944
R16723 gnd.n4972 gnd.n1190 19.3944
R16724 gnd.n6282 gnd.n1190 19.3944
R16725 gnd.n6282 gnd.n6281 19.3944
R16726 gnd.n6281 gnd.n6280 19.3944
R16727 gnd.n6280 gnd.n1194 19.3944
R16728 gnd.n1293 gnd.n1194 19.3944
R16729 gnd.n6263 gnd.n1293 19.3944
R16730 gnd.n6263 gnd.n6262 19.3944
R16731 gnd.n6262 gnd.n6261 19.3944
R16732 gnd.n6261 gnd.n1299 19.3944
R16733 gnd.n5038 gnd.n1299 19.3944
R16734 gnd.n5038 gnd.n2100 19.3944
R16735 gnd.n5042 gnd.n2100 19.3944
R16736 gnd.n5042 gnd.n2076 19.3944
R16737 gnd.n5097 gnd.n2076 19.3944
R16738 gnd.n5097 gnd.n2074 19.3944
R16739 gnd.n5103 gnd.n2074 19.3944
R16740 gnd.n5103 gnd.n5102 19.3944
R16741 gnd.n5102 gnd.n2053 19.3944
R16742 gnd.n5129 gnd.n2053 19.3944
R16743 gnd.n5129 gnd.n2051 19.3944
R16744 gnd.n5135 gnd.n2051 19.3944
R16745 gnd.n5135 gnd.n5134 19.3944
R16746 gnd.n5134 gnd.n2031 19.3944
R16747 gnd.n5179 gnd.n2031 19.3944
R16748 gnd.n5179 gnd.n2029 19.3944
R16749 gnd.n5185 gnd.n2029 19.3944
R16750 gnd.n5185 gnd.n5184 19.3944
R16751 gnd.n5184 gnd.n2003 19.3944
R16752 gnd.n5217 gnd.n2003 19.3944
R16753 gnd.n5217 gnd.n2001 19.3944
R16754 gnd.n5221 gnd.n2001 19.3944
R16755 gnd.n5221 gnd.n1975 19.3944
R16756 gnd.n5254 gnd.n1975 19.3944
R16757 gnd.n5254 gnd.n1973 19.3944
R16758 gnd.n5260 gnd.n1973 19.3944
R16759 gnd.n5260 gnd.n5259 19.3944
R16760 gnd.n5259 gnd.n1956 19.3944
R16761 gnd.n5312 gnd.n1956 19.3944
R16762 gnd.n5312 gnd.n1954 19.3944
R16763 gnd.n5318 gnd.n1954 19.3944
R16764 gnd.n5318 gnd.n5317 19.3944
R16765 gnd.n5317 gnd.n1933 19.3944
R16766 gnd.n5350 gnd.n1933 19.3944
R16767 gnd.n5350 gnd.n1931 19.3944
R16768 gnd.n5356 gnd.n1931 19.3944
R16769 gnd.n5356 gnd.n5355 19.3944
R16770 gnd.n5355 gnd.n1905 19.3944
R16771 gnd.n5406 gnd.n1905 19.3944
R16772 gnd.n5406 gnd.n1903 19.3944
R16773 gnd.n5412 gnd.n1903 19.3944
R16774 gnd.n5412 gnd.n5411 19.3944
R16775 gnd.n5411 gnd.n1884 19.3944
R16776 gnd.n5444 gnd.n1884 19.3944
R16777 gnd.n5444 gnd.n1882 19.3944
R16778 gnd.n5448 gnd.n1882 19.3944
R16779 gnd.n5448 gnd.n1828 19.3944
R16780 gnd.n5619 gnd.n1828 19.3944
R16781 gnd.n5619 gnd.n1826 19.3944
R16782 gnd.n5623 gnd.n1826 19.3944
R16783 gnd.n5623 gnd.n1817 19.3944
R16784 gnd.n5636 gnd.n1817 19.3944
R16785 gnd.n5636 gnd.n1815 19.3944
R16786 gnd.n5640 gnd.n1815 19.3944
R16787 gnd.n5640 gnd.n1805 19.3944
R16788 gnd.n5653 gnd.n1805 19.3944
R16789 gnd.n5653 gnd.n1803 19.3944
R16790 gnd.n5657 gnd.n1803 19.3944
R16791 gnd.n5657 gnd.n1793 19.3944
R16792 gnd.n5670 gnd.n1793 19.3944
R16793 gnd.n5670 gnd.n1791 19.3944
R16794 gnd.n5674 gnd.n1791 19.3944
R16795 gnd.n5674 gnd.n1781 19.3944
R16796 gnd.n5687 gnd.n1781 19.3944
R16797 gnd.n5687 gnd.n1779 19.3944
R16798 gnd.n5694 gnd.n1779 19.3944
R16799 gnd.n5694 gnd.n5693 19.3944
R16800 gnd.n5693 gnd.n1769 19.3944
R16801 gnd.n5708 gnd.n1769 19.3944
R16802 gnd.n5709 gnd.n5708 19.3944
R16803 gnd.n5709 gnd.n1767 19.3944
R16804 gnd.n5724 gnd.n1767 19.3944
R16805 gnd.n5724 gnd.n5723 19.3944
R16806 gnd.n5723 gnd.n5722 19.3944
R16807 gnd.n5722 gnd.n5715 19.3944
R16808 gnd.n5718 gnd.n5715 19.3944
R16809 gnd.n5718 gnd.n1733 19.3944
R16810 gnd.n5778 gnd.n1733 19.3944
R16811 gnd.n5778 gnd.n1731 19.3944
R16812 gnd.n5782 gnd.n1731 19.3944
R16813 gnd.n5782 gnd.n1729 19.3944
R16814 gnd.n5786 gnd.n1729 19.3944
R16815 gnd.n5786 gnd.n1727 19.3944
R16816 gnd.n5790 gnd.n1727 19.3944
R16817 gnd.n5790 gnd.n1725 19.3944
R16818 gnd.n5794 gnd.n1725 19.3944
R16819 gnd.n5794 gnd.n1723 19.3944
R16820 gnd.n5818 gnd.n1723 19.3944
R16821 gnd.n5818 gnd.n5817 19.3944
R16822 gnd.n5817 gnd.n5816 19.3944
R16823 gnd.n5816 gnd.n5800 19.3944
R16824 gnd.n5812 gnd.n5800 19.3944
R16825 gnd.n5812 gnd.n5811 19.3944
R16826 gnd.n5811 gnd.n5810 19.3944
R16827 gnd.n5810 gnd.n5808 19.3944
R16828 gnd.n5808 gnd.n1705 19.3944
R16829 gnd.n1705 gnd.n1703 19.3944
R16830 gnd.n5879 gnd.n1703 19.3944
R16831 gnd.n5879 gnd.n1701 19.3944
R16832 gnd.n5884 gnd.n1701 19.3944
R16833 gnd.n5884 gnd.n389 19.3944
R16834 gnd.n7291 gnd.n389 19.3944
R16835 gnd.n7291 gnd.n7290 19.3944
R16836 gnd.n7078 gnd.n516 19.3944
R16837 gnd.n7078 gnd.n512 19.3944
R16838 gnd.n7084 gnd.n512 19.3944
R16839 gnd.n7084 gnd.n510 19.3944
R16840 gnd.n7088 gnd.n510 19.3944
R16841 gnd.n7088 gnd.n506 19.3944
R16842 gnd.n7094 gnd.n506 19.3944
R16843 gnd.n7094 gnd.n504 19.3944
R16844 gnd.n7098 gnd.n504 19.3944
R16845 gnd.n7098 gnd.n500 19.3944
R16846 gnd.n7104 gnd.n500 19.3944
R16847 gnd.n7104 gnd.n498 19.3944
R16848 gnd.n7108 gnd.n498 19.3944
R16849 gnd.n7108 gnd.n494 19.3944
R16850 gnd.n7114 gnd.n494 19.3944
R16851 gnd.n7114 gnd.n492 19.3944
R16852 gnd.n7118 gnd.n492 19.3944
R16853 gnd.n7118 gnd.n488 19.3944
R16854 gnd.n7124 gnd.n488 19.3944
R16855 gnd.n7124 gnd.n486 19.3944
R16856 gnd.n7128 gnd.n486 19.3944
R16857 gnd.n7128 gnd.n482 19.3944
R16858 gnd.n7134 gnd.n482 19.3944
R16859 gnd.n7134 gnd.n480 19.3944
R16860 gnd.n7138 gnd.n480 19.3944
R16861 gnd.n7138 gnd.n476 19.3944
R16862 gnd.n7144 gnd.n476 19.3944
R16863 gnd.n7144 gnd.n474 19.3944
R16864 gnd.n7148 gnd.n474 19.3944
R16865 gnd.n7148 gnd.n470 19.3944
R16866 gnd.n7154 gnd.n470 19.3944
R16867 gnd.n7154 gnd.n468 19.3944
R16868 gnd.n7158 gnd.n468 19.3944
R16869 gnd.n7158 gnd.n464 19.3944
R16870 gnd.n7164 gnd.n464 19.3944
R16871 gnd.n7164 gnd.n462 19.3944
R16872 gnd.n7168 gnd.n462 19.3944
R16873 gnd.n7168 gnd.n458 19.3944
R16874 gnd.n7174 gnd.n458 19.3944
R16875 gnd.n7174 gnd.n456 19.3944
R16876 gnd.n7178 gnd.n456 19.3944
R16877 gnd.n7178 gnd.n452 19.3944
R16878 gnd.n7184 gnd.n452 19.3944
R16879 gnd.n7184 gnd.n450 19.3944
R16880 gnd.n7188 gnd.n450 19.3944
R16881 gnd.n7188 gnd.n446 19.3944
R16882 gnd.n7194 gnd.n446 19.3944
R16883 gnd.n7194 gnd.n444 19.3944
R16884 gnd.n7198 gnd.n444 19.3944
R16885 gnd.n7198 gnd.n440 19.3944
R16886 gnd.n7204 gnd.n440 19.3944
R16887 gnd.n7204 gnd.n438 19.3944
R16888 gnd.n7208 gnd.n438 19.3944
R16889 gnd.n7208 gnd.n434 19.3944
R16890 gnd.n7214 gnd.n434 19.3944
R16891 gnd.n7214 gnd.n432 19.3944
R16892 gnd.n7218 gnd.n432 19.3944
R16893 gnd.n7218 gnd.n428 19.3944
R16894 gnd.n7224 gnd.n428 19.3944
R16895 gnd.n7224 gnd.n426 19.3944
R16896 gnd.n7228 gnd.n426 19.3944
R16897 gnd.n7228 gnd.n422 19.3944
R16898 gnd.n7234 gnd.n422 19.3944
R16899 gnd.n7234 gnd.n420 19.3944
R16900 gnd.n7238 gnd.n420 19.3944
R16901 gnd.n7238 gnd.n416 19.3944
R16902 gnd.n7244 gnd.n416 19.3944
R16903 gnd.n7244 gnd.n414 19.3944
R16904 gnd.n7248 gnd.n414 19.3944
R16905 gnd.n7248 gnd.n410 19.3944
R16906 gnd.n7254 gnd.n410 19.3944
R16907 gnd.n7254 gnd.n408 19.3944
R16908 gnd.n7258 gnd.n408 19.3944
R16909 gnd.n7258 gnd.n404 19.3944
R16910 gnd.n7264 gnd.n404 19.3944
R16911 gnd.n7264 gnd.n402 19.3944
R16912 gnd.n7268 gnd.n402 19.3944
R16913 gnd.n7268 gnd.n398 19.3944
R16914 gnd.n7274 gnd.n398 19.3944
R16915 gnd.n7274 gnd.n396 19.3944
R16916 gnd.n7280 gnd.n396 19.3944
R16917 gnd.n7280 gnd.n7279 19.3944
R16918 gnd.n7279 gnd.n392 19.3944
R16919 gnd.n7287 gnd.n392 19.3944
R16920 gnd.n6658 gnd.n768 19.3944
R16921 gnd.n6658 gnd.n764 19.3944
R16922 gnd.n6664 gnd.n764 19.3944
R16923 gnd.n6664 gnd.n762 19.3944
R16924 gnd.n6668 gnd.n762 19.3944
R16925 gnd.n6668 gnd.n758 19.3944
R16926 gnd.n6674 gnd.n758 19.3944
R16927 gnd.n6674 gnd.n756 19.3944
R16928 gnd.n6678 gnd.n756 19.3944
R16929 gnd.n6678 gnd.n752 19.3944
R16930 gnd.n6684 gnd.n752 19.3944
R16931 gnd.n6684 gnd.n750 19.3944
R16932 gnd.n6688 gnd.n750 19.3944
R16933 gnd.n6688 gnd.n746 19.3944
R16934 gnd.n6694 gnd.n746 19.3944
R16935 gnd.n6694 gnd.n744 19.3944
R16936 gnd.n6698 gnd.n744 19.3944
R16937 gnd.n6698 gnd.n740 19.3944
R16938 gnd.n6704 gnd.n740 19.3944
R16939 gnd.n6704 gnd.n738 19.3944
R16940 gnd.n6708 gnd.n738 19.3944
R16941 gnd.n6708 gnd.n734 19.3944
R16942 gnd.n6714 gnd.n734 19.3944
R16943 gnd.n6714 gnd.n732 19.3944
R16944 gnd.n6718 gnd.n732 19.3944
R16945 gnd.n6718 gnd.n728 19.3944
R16946 gnd.n6724 gnd.n728 19.3944
R16947 gnd.n6724 gnd.n726 19.3944
R16948 gnd.n6728 gnd.n726 19.3944
R16949 gnd.n6728 gnd.n722 19.3944
R16950 gnd.n6734 gnd.n722 19.3944
R16951 gnd.n6734 gnd.n720 19.3944
R16952 gnd.n6738 gnd.n720 19.3944
R16953 gnd.n6738 gnd.n716 19.3944
R16954 gnd.n6744 gnd.n716 19.3944
R16955 gnd.n6744 gnd.n714 19.3944
R16956 gnd.n6748 gnd.n714 19.3944
R16957 gnd.n6748 gnd.n710 19.3944
R16958 gnd.n6754 gnd.n710 19.3944
R16959 gnd.n6754 gnd.n708 19.3944
R16960 gnd.n6758 gnd.n708 19.3944
R16961 gnd.n6758 gnd.n704 19.3944
R16962 gnd.n6764 gnd.n704 19.3944
R16963 gnd.n6764 gnd.n702 19.3944
R16964 gnd.n6768 gnd.n702 19.3944
R16965 gnd.n6768 gnd.n698 19.3944
R16966 gnd.n6774 gnd.n698 19.3944
R16967 gnd.n6774 gnd.n696 19.3944
R16968 gnd.n6778 gnd.n696 19.3944
R16969 gnd.n6778 gnd.n692 19.3944
R16970 gnd.n6784 gnd.n692 19.3944
R16971 gnd.n6784 gnd.n690 19.3944
R16972 gnd.n6788 gnd.n690 19.3944
R16973 gnd.n6788 gnd.n686 19.3944
R16974 gnd.n6794 gnd.n686 19.3944
R16975 gnd.n6794 gnd.n684 19.3944
R16976 gnd.n6798 gnd.n684 19.3944
R16977 gnd.n6798 gnd.n680 19.3944
R16978 gnd.n6804 gnd.n680 19.3944
R16979 gnd.n6804 gnd.n678 19.3944
R16980 gnd.n6808 gnd.n678 19.3944
R16981 gnd.n6808 gnd.n674 19.3944
R16982 gnd.n6814 gnd.n674 19.3944
R16983 gnd.n6814 gnd.n672 19.3944
R16984 gnd.n6818 gnd.n672 19.3944
R16985 gnd.n6818 gnd.n668 19.3944
R16986 gnd.n6824 gnd.n668 19.3944
R16987 gnd.n6824 gnd.n666 19.3944
R16988 gnd.n6828 gnd.n666 19.3944
R16989 gnd.n6828 gnd.n662 19.3944
R16990 gnd.n6834 gnd.n662 19.3944
R16991 gnd.n6834 gnd.n660 19.3944
R16992 gnd.n6838 gnd.n660 19.3944
R16993 gnd.n6838 gnd.n656 19.3944
R16994 gnd.n6844 gnd.n656 19.3944
R16995 gnd.n6844 gnd.n654 19.3944
R16996 gnd.n6848 gnd.n654 19.3944
R16997 gnd.n6848 gnd.n650 19.3944
R16998 gnd.n6854 gnd.n650 19.3944
R16999 gnd.n6854 gnd.n648 19.3944
R17000 gnd.n6858 gnd.n648 19.3944
R17001 gnd.n6858 gnd.n644 19.3944
R17002 gnd.n6864 gnd.n644 19.3944
R17003 gnd.n6864 gnd.n642 19.3944
R17004 gnd.n6868 gnd.n642 19.3944
R17005 gnd.n6868 gnd.n638 19.3944
R17006 gnd.n6874 gnd.n638 19.3944
R17007 gnd.n6874 gnd.n636 19.3944
R17008 gnd.n6878 gnd.n636 19.3944
R17009 gnd.n6878 gnd.n632 19.3944
R17010 gnd.n6884 gnd.n632 19.3944
R17011 gnd.n6884 gnd.n630 19.3944
R17012 gnd.n6888 gnd.n630 19.3944
R17013 gnd.n6888 gnd.n626 19.3944
R17014 gnd.n6894 gnd.n626 19.3944
R17015 gnd.n6894 gnd.n624 19.3944
R17016 gnd.n6898 gnd.n624 19.3944
R17017 gnd.n6898 gnd.n620 19.3944
R17018 gnd.n6904 gnd.n620 19.3944
R17019 gnd.n6904 gnd.n618 19.3944
R17020 gnd.n6908 gnd.n618 19.3944
R17021 gnd.n6908 gnd.n614 19.3944
R17022 gnd.n6914 gnd.n614 19.3944
R17023 gnd.n6914 gnd.n612 19.3944
R17024 gnd.n6918 gnd.n612 19.3944
R17025 gnd.n6918 gnd.n608 19.3944
R17026 gnd.n6924 gnd.n608 19.3944
R17027 gnd.n6924 gnd.n606 19.3944
R17028 gnd.n6928 gnd.n606 19.3944
R17029 gnd.n6928 gnd.n602 19.3944
R17030 gnd.n6934 gnd.n602 19.3944
R17031 gnd.n6934 gnd.n600 19.3944
R17032 gnd.n6938 gnd.n600 19.3944
R17033 gnd.n6938 gnd.n596 19.3944
R17034 gnd.n6944 gnd.n596 19.3944
R17035 gnd.n6944 gnd.n594 19.3944
R17036 gnd.n6948 gnd.n594 19.3944
R17037 gnd.n6948 gnd.n590 19.3944
R17038 gnd.n6954 gnd.n590 19.3944
R17039 gnd.n6954 gnd.n588 19.3944
R17040 gnd.n6958 gnd.n588 19.3944
R17041 gnd.n6958 gnd.n584 19.3944
R17042 gnd.n6964 gnd.n584 19.3944
R17043 gnd.n6964 gnd.n582 19.3944
R17044 gnd.n6968 gnd.n582 19.3944
R17045 gnd.n6968 gnd.n578 19.3944
R17046 gnd.n6974 gnd.n578 19.3944
R17047 gnd.n6974 gnd.n576 19.3944
R17048 gnd.n6978 gnd.n576 19.3944
R17049 gnd.n6978 gnd.n572 19.3944
R17050 gnd.n6984 gnd.n572 19.3944
R17051 gnd.n6984 gnd.n570 19.3944
R17052 gnd.n6988 gnd.n570 19.3944
R17053 gnd.n6988 gnd.n566 19.3944
R17054 gnd.n6994 gnd.n566 19.3944
R17055 gnd.n6994 gnd.n564 19.3944
R17056 gnd.n6998 gnd.n564 19.3944
R17057 gnd.n6998 gnd.n560 19.3944
R17058 gnd.n7004 gnd.n560 19.3944
R17059 gnd.n7004 gnd.n558 19.3944
R17060 gnd.n7008 gnd.n558 19.3944
R17061 gnd.n7008 gnd.n554 19.3944
R17062 gnd.n7014 gnd.n554 19.3944
R17063 gnd.n7014 gnd.n552 19.3944
R17064 gnd.n7018 gnd.n552 19.3944
R17065 gnd.n7018 gnd.n548 19.3944
R17066 gnd.n7024 gnd.n548 19.3944
R17067 gnd.n7024 gnd.n546 19.3944
R17068 gnd.n7028 gnd.n546 19.3944
R17069 gnd.n7028 gnd.n542 19.3944
R17070 gnd.n7034 gnd.n542 19.3944
R17071 gnd.n7034 gnd.n540 19.3944
R17072 gnd.n7038 gnd.n540 19.3944
R17073 gnd.n7038 gnd.n536 19.3944
R17074 gnd.n7044 gnd.n536 19.3944
R17075 gnd.n7044 gnd.n534 19.3944
R17076 gnd.n7048 gnd.n534 19.3944
R17077 gnd.n7048 gnd.n530 19.3944
R17078 gnd.n7054 gnd.n530 19.3944
R17079 gnd.n7054 gnd.n528 19.3944
R17080 gnd.n7058 gnd.n528 19.3944
R17081 gnd.n7058 gnd.n524 19.3944
R17082 gnd.n7064 gnd.n524 19.3944
R17083 gnd.n7064 gnd.n522 19.3944
R17084 gnd.n7068 gnd.n522 19.3944
R17085 gnd.n7068 gnd.n518 19.3944
R17086 gnd.n7074 gnd.n518 19.3944
R17087 gnd.n6077 gnd.n6076 19.3944
R17088 gnd.n6076 gnd.n6075 19.3944
R17089 gnd.n6075 gnd.n6074 19.3944
R17090 gnd.n6074 gnd.n6072 19.3944
R17091 gnd.n6072 gnd.n6069 19.3944
R17092 gnd.n6069 gnd.n6068 19.3944
R17093 gnd.n6068 gnd.n6065 19.3944
R17094 gnd.n6065 gnd.n6064 19.3944
R17095 gnd.n6064 gnd.n6061 19.3944
R17096 gnd.n6061 gnd.n6060 19.3944
R17097 gnd.n6060 gnd.n6057 19.3944
R17098 gnd.n6057 gnd.n6056 19.3944
R17099 gnd.n6056 gnd.n6053 19.3944
R17100 gnd.n6053 gnd.n6052 19.3944
R17101 gnd.n6052 gnd.n6049 19.3944
R17102 gnd.n6049 gnd.n6048 19.3944
R17103 gnd.n6048 gnd.n6045 19.3944
R17104 gnd.n6043 gnd.n6040 19.3944
R17105 gnd.n6040 gnd.n6039 19.3944
R17106 gnd.n6039 gnd.n6036 19.3944
R17107 gnd.n6036 gnd.n6035 19.3944
R17108 gnd.n6035 gnd.n6032 19.3944
R17109 gnd.n6032 gnd.n6031 19.3944
R17110 gnd.n6031 gnd.n6028 19.3944
R17111 gnd.n6026 gnd.n6023 19.3944
R17112 gnd.n6023 gnd.n6022 19.3944
R17113 gnd.n6022 gnd.n6019 19.3944
R17114 gnd.n6019 gnd.n6018 19.3944
R17115 gnd.n6018 gnd.n6015 19.3944
R17116 gnd.n6015 gnd.n6014 19.3944
R17117 gnd.n6014 gnd.n6011 19.3944
R17118 gnd.n6011 gnd.n6010 19.3944
R17119 gnd.n6006 gnd.n6003 19.3944
R17120 gnd.n6003 gnd.n6002 19.3944
R17121 gnd.n6002 gnd.n5999 19.3944
R17122 gnd.n5999 gnd.n5998 19.3944
R17123 gnd.n5998 gnd.n5995 19.3944
R17124 gnd.n5995 gnd.n5994 19.3944
R17125 gnd.n5994 gnd.n5991 19.3944
R17126 gnd.n5991 gnd.n5990 19.3944
R17127 gnd.n5990 gnd.n5987 19.3944
R17128 gnd.n5987 gnd.n5986 19.3944
R17129 gnd.n5986 gnd.n5983 19.3944
R17130 gnd.n5983 gnd.n5982 19.3944
R17131 gnd.n5982 gnd.n5979 19.3944
R17132 gnd.n5979 gnd.n5978 19.3944
R17133 gnd.n5978 gnd.n5975 19.3944
R17134 gnd.n5975 gnd.n5974 19.3944
R17135 gnd.n5974 gnd.n5971 19.3944
R17136 gnd.n5971 gnd.n5970 19.3944
R17137 gnd.n5954 gnd.n1574 19.3944
R17138 gnd.n5954 gnd.n5953 19.3944
R17139 gnd.n5953 gnd.n1583 19.3944
R17140 gnd.n5742 gnd.n1583 19.3944
R17141 gnd.n5745 gnd.n5742 19.3944
R17142 gnd.n5746 gnd.n5745 19.3944
R17143 gnd.n5751 gnd.n5746 19.3944
R17144 gnd.n5752 gnd.n5751 19.3944
R17145 gnd.n5756 gnd.n5752 19.3944
R17146 gnd.n5756 gnd.n5755 19.3944
R17147 gnd.n5755 gnd.n5754 19.3944
R17148 gnd.n5754 gnd.n1716 19.3944
R17149 gnd.n5831 gnd.n1716 19.3944
R17150 gnd.n5832 gnd.n5831 19.3944
R17151 gnd.n5834 gnd.n5832 19.3944
R17152 gnd.n5834 gnd.n1711 19.3944
R17153 gnd.n5846 gnd.n1711 19.3944
R17154 gnd.n5847 gnd.n5846 19.3944
R17155 gnd.n5849 gnd.n5847 19.3944
R17156 gnd.n5850 gnd.n5849 19.3944
R17157 gnd.n5856 gnd.n5850 19.3944
R17158 gnd.n5856 gnd.n5855 19.3944
R17159 gnd.n5855 gnd.n5854 19.3944
R17160 gnd.n5854 gnd.n5853 19.3944
R17161 gnd.n5853 gnd.n377 19.3944
R17162 gnd.n7304 gnd.n377 19.3944
R17163 gnd.n7306 gnd.n7304 19.3944
R17164 gnd.n7306 gnd.n7305 19.3944
R17165 gnd.n7305 gnd.n370 19.3944
R17166 gnd.n7355 gnd.n370 19.3944
R17167 gnd.n7355 gnd.n7354 19.3944
R17168 gnd.n7354 gnd.n7353 19.3944
R17169 gnd.n7353 gnd.n7351 19.3944
R17170 gnd.n7351 gnd.n7350 19.3944
R17171 gnd.n7350 gnd.n7348 19.3944
R17172 gnd.n7348 gnd.n7347 19.3944
R17173 gnd.n7347 gnd.n7345 19.3944
R17174 gnd.n7345 gnd.n7344 19.3944
R17175 gnd.n7344 gnd.n7342 19.3944
R17176 gnd.n7342 gnd.n7341 19.3944
R17177 gnd.n7341 gnd.n7339 19.3944
R17178 gnd.n7339 gnd.n7338 19.3944
R17179 gnd.n7338 gnd.n7336 19.3944
R17180 gnd.n7336 gnd.n7335 19.3944
R17181 gnd.n7335 gnd.n7333 19.3944
R17182 gnd.n7333 gnd.n7332 19.3944
R17183 gnd.n7332 gnd.n7330 19.3944
R17184 gnd.n7330 gnd.n7329 19.3944
R17185 gnd.n7329 gnd.n7327 19.3944
R17186 gnd.n7327 gnd.n7326 19.3944
R17187 gnd.n7326 gnd.n7324 19.3944
R17188 gnd.n7324 gnd.n7323 19.3944
R17189 gnd.n7323 gnd.n7321 19.3944
R17190 gnd.n5957 gnd.n5956 19.3944
R17191 gnd.n5956 gnd.n1581 19.3944
R17192 gnd.n1605 gnd.n1581 19.3944
R17193 gnd.n5943 gnd.n1605 19.3944
R17194 gnd.n5943 gnd.n5942 19.3944
R17195 gnd.n5942 gnd.n5941 19.3944
R17196 gnd.n5941 gnd.n1610 19.3944
R17197 gnd.n5931 gnd.n1610 19.3944
R17198 gnd.n5931 gnd.n5930 19.3944
R17199 gnd.n5930 gnd.n5929 19.3944
R17200 gnd.n5929 gnd.n1630 19.3944
R17201 gnd.n5919 gnd.n1630 19.3944
R17202 gnd.n5919 gnd.n5918 19.3944
R17203 gnd.n5918 gnd.n5917 19.3944
R17204 gnd.n5917 gnd.n1650 19.3944
R17205 gnd.n5907 gnd.n1650 19.3944
R17206 gnd.n5907 gnd.n5906 19.3944
R17207 gnd.n5906 gnd.n5905 19.3944
R17208 gnd.n5905 gnd.n1670 19.3944
R17209 gnd.n5895 gnd.n1670 19.3944
R17210 gnd.n5895 gnd.n5894 19.3944
R17211 gnd.n5894 gnd.n5893 19.3944
R17212 gnd.n5893 gnd.n1690 19.3944
R17213 gnd.n1690 gnd.n379 19.3944
R17214 gnd.n7301 gnd.n379 19.3944
R17215 gnd.n7301 gnd.n372 19.3944
R17216 gnd.n7310 gnd.n372 19.3944
R17217 gnd.n7311 gnd.n7310 19.3944
R17218 gnd.n7313 gnd.n7311 19.3944
R17219 gnd.n7313 gnd.n110 19.3944
R17220 gnd.n7613 gnd.n110 19.3944
R17221 gnd.n7613 gnd.n7612 19.3944
R17222 gnd.n7612 gnd.n7611 19.3944
R17223 gnd.n7611 gnd.n114 19.3944
R17224 gnd.n7601 gnd.n114 19.3944
R17225 gnd.n7601 gnd.n7600 19.3944
R17226 gnd.n7600 gnd.n7599 19.3944
R17227 gnd.n7599 gnd.n131 19.3944
R17228 gnd.n7589 gnd.n131 19.3944
R17229 gnd.n7589 gnd.n7588 19.3944
R17230 gnd.n7588 gnd.n7587 19.3944
R17231 gnd.n7587 gnd.n151 19.3944
R17232 gnd.n7577 gnd.n151 19.3944
R17233 gnd.n7577 gnd.n7576 19.3944
R17234 gnd.n7576 gnd.n7575 19.3944
R17235 gnd.n7575 gnd.n169 19.3944
R17236 gnd.n7565 gnd.n169 19.3944
R17237 gnd.n7565 gnd.n7564 19.3944
R17238 gnd.n7564 gnd.n7563 19.3944
R17239 gnd.n7563 gnd.n189 19.3944
R17240 gnd.n7553 gnd.n189 19.3944
R17241 gnd.n7553 gnd.n7552 19.3944
R17242 gnd.n7552 gnd.n7551 19.3944
R17243 gnd.n7473 gnd.n279 19.3944
R17244 gnd.n7473 gnd.n283 19.3944
R17245 gnd.n286 gnd.n283 19.3944
R17246 gnd.n7466 gnd.n286 19.3944
R17247 gnd.n7466 gnd.n7465 19.3944
R17248 gnd.n7465 gnd.n7464 19.3944
R17249 gnd.n7464 gnd.n292 19.3944
R17250 gnd.n7459 gnd.n292 19.3944
R17251 gnd.n7459 gnd.n7458 19.3944
R17252 gnd.n7458 gnd.n7457 19.3944
R17253 gnd.n7457 gnd.n299 19.3944
R17254 gnd.n7452 gnd.n299 19.3944
R17255 gnd.n7452 gnd.n7451 19.3944
R17256 gnd.n7451 gnd.n7450 19.3944
R17257 gnd.n7450 gnd.n306 19.3944
R17258 gnd.n7445 gnd.n306 19.3944
R17259 gnd.n7445 gnd.n7444 19.3944
R17260 gnd.n7444 gnd.n7443 19.3944
R17261 gnd.n7511 gnd.n246 19.3944
R17262 gnd.n7506 gnd.n246 19.3944
R17263 gnd.n7506 gnd.n7505 19.3944
R17264 gnd.n7505 gnd.n7504 19.3944
R17265 gnd.n7504 gnd.n253 19.3944
R17266 gnd.n7499 gnd.n253 19.3944
R17267 gnd.n7499 gnd.n7498 19.3944
R17268 gnd.n7498 gnd.n7497 19.3944
R17269 gnd.n7497 gnd.n260 19.3944
R17270 gnd.n7492 gnd.n260 19.3944
R17271 gnd.n7492 gnd.n7491 19.3944
R17272 gnd.n7491 gnd.n7490 19.3944
R17273 gnd.n7490 gnd.n267 19.3944
R17274 gnd.n7485 gnd.n267 19.3944
R17275 gnd.n7485 gnd.n7484 19.3944
R17276 gnd.n7484 gnd.n7483 19.3944
R17277 gnd.n7483 gnd.n274 19.3944
R17278 gnd.n7478 gnd.n274 19.3944
R17279 gnd.n7544 gnd.n7543 19.3944
R17280 gnd.n7543 gnd.n7542 19.3944
R17281 gnd.n7542 gnd.n218 19.3944
R17282 gnd.n7537 gnd.n218 19.3944
R17283 gnd.n7537 gnd.n7536 19.3944
R17284 gnd.n7536 gnd.n7535 19.3944
R17285 gnd.n7535 gnd.n225 19.3944
R17286 gnd.n7530 gnd.n225 19.3944
R17287 gnd.n7530 gnd.n7529 19.3944
R17288 gnd.n7529 gnd.n7528 19.3944
R17289 gnd.n7528 gnd.n232 19.3944
R17290 gnd.n7523 gnd.n232 19.3944
R17291 gnd.n7523 gnd.n7522 19.3944
R17292 gnd.n7522 gnd.n7521 19.3944
R17293 gnd.n7521 gnd.n239 19.3944
R17294 gnd.n7516 gnd.n239 19.3944
R17295 gnd.n7516 gnd.n7515 19.3944
R17296 gnd.n7434 gnd.n7433 19.3944
R17297 gnd.n7433 gnd.n7432 19.3944
R17298 gnd.n7432 gnd.n321 19.3944
R17299 gnd.n7427 gnd.n321 19.3944
R17300 gnd.n7427 gnd.n7426 19.3944
R17301 gnd.n7426 gnd.n7425 19.3944
R17302 gnd.n7425 gnd.n328 19.3944
R17303 gnd.n7420 gnd.n328 19.3944
R17304 gnd.n7420 gnd.n7419 19.3944
R17305 gnd.n7419 gnd.n7418 19.3944
R17306 gnd.n7418 gnd.n335 19.3944
R17307 gnd.n7413 gnd.n335 19.3944
R17308 gnd.n7413 gnd.n7412 19.3944
R17309 gnd.n7412 gnd.n7411 19.3944
R17310 gnd.n7411 gnd.n342 19.3944
R17311 gnd.n7406 gnd.n342 19.3944
R17312 gnd.n5773 gnd.n1735 19.3944
R17313 gnd.n5773 gnd.n1736 19.3944
R17314 gnd.n5769 gnd.n1736 19.3944
R17315 gnd.n5769 gnd.n5768 19.3944
R17316 gnd.n5768 gnd.n5767 19.3944
R17317 gnd.n5767 gnd.n5739 19.3944
R17318 gnd.n5763 gnd.n5739 19.3944
R17319 gnd.n5763 gnd.n5762 19.3944
R17320 gnd.n5762 gnd.n5761 19.3944
R17321 gnd.n5761 gnd.n1719 19.3944
R17322 gnd.n5823 gnd.n1719 19.3944
R17323 gnd.n5823 gnd.n1717 19.3944
R17324 gnd.n5827 gnd.n1717 19.3944
R17325 gnd.n5827 gnd.n1714 19.3944
R17326 gnd.n5838 gnd.n1714 19.3944
R17327 gnd.n5838 gnd.n1712 19.3944
R17328 gnd.n5842 gnd.n1712 19.3944
R17329 gnd.n5842 gnd.n1707 19.3944
R17330 gnd.n5872 gnd.n1707 19.3944
R17331 gnd.n5872 gnd.n1708 19.3944
R17332 gnd.n5868 gnd.n1708 19.3944
R17333 gnd.n5868 gnd.n5867 19.3944
R17334 gnd.n5867 gnd.n5866 19.3944
R17335 gnd.n5866 gnd.n5861 19.3944
R17336 gnd.n5862 gnd.n5861 19.3944
R17337 gnd.n5862 gnd.n85 19.3944
R17338 gnd.n7626 gnd.n85 19.3944
R17339 gnd.n7626 gnd.n7625 19.3944
R17340 gnd.n7625 gnd.n87 19.3944
R17341 gnd.n7359 gnd.n87 19.3944
R17342 gnd.n7363 gnd.n7359 19.3944
R17343 gnd.n7365 gnd.n7363 19.3944
R17344 gnd.n7366 gnd.n7365 19.3944
R17345 gnd.n7366 gnd.n366 19.3944
R17346 gnd.n7370 gnd.n366 19.3944
R17347 gnd.n7372 gnd.n7370 19.3944
R17348 gnd.n7373 gnd.n7372 19.3944
R17349 gnd.n7373 gnd.n363 19.3944
R17350 gnd.n7377 gnd.n363 19.3944
R17351 gnd.n7379 gnd.n7377 19.3944
R17352 gnd.n7380 gnd.n7379 19.3944
R17353 gnd.n7380 gnd.n360 19.3944
R17354 gnd.n7384 gnd.n360 19.3944
R17355 gnd.n7386 gnd.n7384 19.3944
R17356 gnd.n7387 gnd.n7386 19.3944
R17357 gnd.n7387 gnd.n357 19.3944
R17358 gnd.n7391 gnd.n357 19.3944
R17359 gnd.n7393 gnd.n7391 19.3944
R17360 gnd.n7394 gnd.n7393 19.3944
R17361 gnd.n7394 gnd.n354 19.3944
R17362 gnd.n7398 gnd.n354 19.3944
R17363 gnd.n7400 gnd.n7398 19.3944
R17364 gnd.n7401 gnd.n7400 19.3944
R17365 gnd.n1591 gnd.n1590 19.3944
R17366 gnd.n5949 gnd.n1590 19.3944
R17367 gnd.n5949 gnd.n5948 19.3944
R17368 gnd.n5948 gnd.n5947 19.3944
R17369 gnd.n5947 gnd.n1597 19.3944
R17370 gnd.n5937 gnd.n1597 19.3944
R17371 gnd.n5937 gnd.n5936 19.3944
R17372 gnd.n5936 gnd.n5935 19.3944
R17373 gnd.n5935 gnd.n1620 19.3944
R17374 gnd.n5925 gnd.n1620 19.3944
R17375 gnd.n5925 gnd.n5924 19.3944
R17376 gnd.n5924 gnd.n5923 19.3944
R17377 gnd.n5923 gnd.n1641 19.3944
R17378 gnd.n5913 gnd.n1641 19.3944
R17379 gnd.n5913 gnd.n5912 19.3944
R17380 gnd.n5912 gnd.n5911 19.3944
R17381 gnd.n5911 gnd.n1660 19.3944
R17382 gnd.n5901 gnd.n1660 19.3944
R17383 gnd.n5901 gnd.n5900 19.3944
R17384 gnd.n5900 gnd.n5899 19.3944
R17385 gnd.n5899 gnd.n1681 19.3944
R17386 gnd.n5889 gnd.n1681 19.3944
R17387 gnd.n1695 gnd.n100 19.3944
R17388 gnd.n7297 gnd.n100 19.3944
R17389 gnd.n386 gnd.n385 19.3944
R17390 gnd.n7621 gnd.n7620 19.3944
R17391 gnd.n7617 gnd.n95 19.3944
R17392 gnd.n7617 gnd.n102 19.3944
R17393 gnd.n7607 gnd.n102 19.3944
R17394 gnd.n7607 gnd.n7606 19.3944
R17395 gnd.n7606 gnd.n7605 19.3944
R17396 gnd.n7605 gnd.n122 19.3944
R17397 gnd.n7595 gnd.n122 19.3944
R17398 gnd.n7595 gnd.n7594 19.3944
R17399 gnd.n7594 gnd.n7593 19.3944
R17400 gnd.n7593 gnd.n142 19.3944
R17401 gnd.n7583 gnd.n142 19.3944
R17402 gnd.n7583 gnd.n7582 19.3944
R17403 gnd.n7582 gnd.n7581 19.3944
R17404 gnd.n7581 gnd.n160 19.3944
R17405 gnd.n7571 gnd.n160 19.3944
R17406 gnd.n7571 gnd.n7570 19.3944
R17407 gnd.n7570 gnd.n7569 19.3944
R17408 gnd.n7569 gnd.n180 19.3944
R17409 gnd.n7559 gnd.n180 19.3944
R17410 gnd.n7559 gnd.n7558 19.3944
R17411 gnd.n7558 gnd.n7557 19.3944
R17412 gnd.n7557 gnd.n200 19.3944
R17413 gnd.n7547 gnd.n200 19.3944
R17414 gnd.n4438 gnd.n4437 19.3944
R17415 gnd.n4437 gnd.n4436 19.3944
R17416 gnd.n4436 gnd.n4435 19.3944
R17417 gnd.n4435 gnd.n4433 19.3944
R17418 gnd.n4433 gnd.n4430 19.3944
R17419 gnd.n4430 gnd.n4429 19.3944
R17420 gnd.n4429 gnd.n4426 19.3944
R17421 gnd.n4426 gnd.n4425 19.3944
R17422 gnd.n4425 gnd.n4422 19.3944
R17423 gnd.n4422 gnd.n4421 19.3944
R17424 gnd.n4421 gnd.n4418 19.3944
R17425 gnd.n4418 gnd.n4417 19.3944
R17426 gnd.n4417 gnd.n4414 19.3944
R17427 gnd.n4414 gnd.n4413 19.3944
R17428 gnd.n4413 gnd.n4410 19.3944
R17429 gnd.n4410 gnd.n4409 19.3944
R17430 gnd.n4409 gnd.n4406 19.3944
R17431 gnd.n4404 gnd.n4401 19.3944
R17432 gnd.n4401 gnd.n4400 19.3944
R17433 gnd.n4400 gnd.n4397 19.3944
R17434 gnd.n4397 gnd.n4396 19.3944
R17435 gnd.n4396 gnd.n4393 19.3944
R17436 gnd.n4393 gnd.n4392 19.3944
R17437 gnd.n4392 gnd.n4389 19.3944
R17438 gnd.n4389 gnd.n4388 19.3944
R17439 gnd.n4388 gnd.n4385 19.3944
R17440 gnd.n4385 gnd.n4384 19.3944
R17441 gnd.n4384 gnd.n4381 19.3944
R17442 gnd.n4381 gnd.n4380 19.3944
R17443 gnd.n4380 gnd.n4377 19.3944
R17444 gnd.n4377 gnd.n4376 19.3944
R17445 gnd.n4376 gnd.n4373 19.3944
R17446 gnd.n4373 gnd.n4372 19.3944
R17447 gnd.n4372 gnd.n4369 19.3944
R17448 gnd.n4369 gnd.n4368 19.3944
R17449 gnd.n4364 gnd.n4361 19.3944
R17450 gnd.n4361 gnd.n4360 19.3944
R17451 gnd.n4360 gnd.n4357 19.3944
R17452 gnd.n4357 gnd.n4356 19.3944
R17453 gnd.n4356 gnd.n4353 19.3944
R17454 gnd.n4353 gnd.n4352 19.3944
R17455 gnd.n4352 gnd.n4349 19.3944
R17456 gnd.n4349 gnd.n4348 19.3944
R17457 gnd.n4348 gnd.n4345 19.3944
R17458 gnd.n4345 gnd.n4344 19.3944
R17459 gnd.n4344 gnd.n4341 19.3944
R17460 gnd.n4341 gnd.n4340 19.3944
R17461 gnd.n4340 gnd.n4337 19.3944
R17462 gnd.n4337 gnd.n4336 19.3944
R17463 gnd.n4336 gnd.n4333 19.3944
R17464 gnd.n4333 gnd.n4332 19.3944
R17465 gnd.n4332 gnd.n4329 19.3944
R17466 gnd.n4329 gnd.n4328 19.3944
R17467 gnd.n4321 gnd.n4319 19.3944
R17468 gnd.n4319 gnd.n4316 19.3944
R17469 gnd.n4316 gnd.n4315 19.3944
R17470 gnd.n4315 gnd.n4312 19.3944
R17471 gnd.n4312 gnd.n4311 19.3944
R17472 gnd.n4311 gnd.n4308 19.3944
R17473 gnd.n4308 gnd.n4307 19.3944
R17474 gnd.n4307 gnd.n4304 19.3944
R17475 gnd.n4304 gnd.n4303 19.3944
R17476 gnd.n4303 gnd.n4300 19.3944
R17477 gnd.n4300 gnd.n4299 19.3944
R17478 gnd.n4299 gnd.n4296 19.3944
R17479 gnd.n4296 gnd.n4295 19.3944
R17480 gnd.n4295 gnd.n4292 19.3944
R17481 gnd.n4292 gnd.n4291 19.3944
R17482 gnd.n4291 gnd.n4288 19.3944
R17483 gnd.n4282 gnd.n4280 19.3944
R17484 gnd.n4280 gnd.n4279 19.3944
R17485 gnd.n4279 gnd.n4277 19.3944
R17486 gnd.n4277 gnd.n4276 19.3944
R17487 gnd.n4276 gnd.n4274 19.3944
R17488 gnd.n4274 gnd.n4273 19.3944
R17489 gnd.n4273 gnd.n4271 19.3944
R17490 gnd.n4271 gnd.n4270 19.3944
R17491 gnd.n4270 gnd.n4268 19.3944
R17492 gnd.n4268 gnd.n4267 19.3944
R17493 gnd.n4267 gnd.n4265 19.3944
R17494 gnd.n4265 gnd.n4264 19.3944
R17495 gnd.n4264 gnd.n4262 19.3944
R17496 gnd.n4262 gnd.n2570 19.3944
R17497 gnd.n4527 gnd.n2570 19.3944
R17498 gnd.n4527 gnd.n2568 19.3944
R17499 gnd.n4543 gnd.n2568 19.3944
R17500 gnd.n4543 gnd.n4542 19.3944
R17501 gnd.n4542 gnd.n4541 19.3944
R17502 gnd.n4541 gnd.n4539 19.3944
R17503 gnd.n4539 gnd.n4538 19.3944
R17504 gnd.n4538 gnd.n4536 19.3944
R17505 gnd.n4536 gnd.n2534 19.3944
R17506 gnd.n4588 gnd.n2534 19.3944
R17507 gnd.n4588 gnd.n2532 19.3944
R17508 gnd.n4598 gnd.n2532 19.3944
R17509 gnd.n4598 gnd.n4597 19.3944
R17510 gnd.n4597 gnd.n4593 19.3944
R17511 gnd.n4593 gnd.n2504 19.3944
R17512 gnd.n4651 gnd.n2504 19.3944
R17513 gnd.n4651 gnd.n2502 19.3944
R17514 gnd.n4655 gnd.n2502 19.3944
R17515 gnd.n4655 gnd.n2499 19.3944
R17516 gnd.n4666 gnd.n2499 19.3944
R17517 gnd.n4666 gnd.n2497 19.3944
R17518 gnd.n4670 gnd.n2497 19.3944
R17519 gnd.n4670 gnd.n2488 19.3944
R17520 gnd.n4706 gnd.n2488 19.3944
R17521 gnd.n4706 gnd.n2489 19.3944
R17522 gnd.n4702 gnd.n2489 19.3944
R17523 gnd.n4702 gnd.n4701 19.3944
R17524 gnd.n4701 gnd.n4700 19.3944
R17525 gnd.n4700 gnd.n2494 19.3944
R17526 gnd.n4696 gnd.n2494 19.3944
R17527 gnd.n4696 gnd.n4695 19.3944
R17528 gnd.n4695 gnd.n4694 19.3944
R17529 gnd.n4694 gnd.n2472 19.3944
R17530 gnd.n4764 gnd.n2472 19.3944
R17531 gnd.n4764 gnd.n2470 19.3944
R17532 gnd.n4769 gnd.n2470 19.3944
R17533 gnd.n4769 gnd.n2466 19.3944
R17534 gnd.n4780 gnd.n2466 19.3944
R17535 gnd.n4781 gnd.n4780 19.3944
R17536 gnd.n4447 gnd.n4445 19.3944
R17537 gnd.n4447 gnd.n4446 19.3944
R17538 gnd.n4446 gnd.n2625 19.3944
R17539 gnd.n4462 gnd.n2625 19.3944
R17540 gnd.n4463 gnd.n4462 19.3944
R17541 gnd.n4464 gnd.n4463 19.3944
R17542 gnd.n4464 gnd.n2607 19.3944
R17543 gnd.n4482 gnd.n2607 19.3944
R17544 gnd.n4483 gnd.n4482 19.3944
R17545 gnd.n4484 gnd.n4483 19.3944
R17546 gnd.n4484 gnd.n2589 19.3944
R17547 gnd.n4502 gnd.n2589 19.3944
R17548 gnd.n4503 gnd.n4502 19.3944
R17549 gnd.n4505 gnd.n4503 19.3944
R17550 gnd.n4506 gnd.n4505 19.3944
R17551 gnd.n4506 gnd.n2563 19.3944
R17552 gnd.n4547 gnd.n2563 19.3944
R17553 gnd.n4548 gnd.n4547 19.3944
R17554 gnd.n4549 gnd.n4548 19.3944
R17555 gnd.n4549 gnd.n2546 19.3944
R17556 gnd.n4568 gnd.n2546 19.3944
R17557 gnd.n4569 gnd.n4568 19.3944
R17558 gnd.n4570 gnd.n4569 19.3944
R17559 gnd.n4572 gnd.n4570 19.3944
R17560 gnd.n4572 gnd.n2530 19.3944
R17561 gnd.n4602 gnd.n2530 19.3944
R17562 gnd.n4603 gnd.n4602 19.3944
R17563 gnd.n4605 gnd.n4603 19.3944
R17564 gnd.n4607 gnd.n4605 19.3944
R17565 gnd.n4607 gnd.n4606 19.3944
R17566 gnd.n4606 gnd.n2501 19.3944
R17567 gnd.n4659 gnd.n2501 19.3944
R17568 gnd.n4660 gnd.n4659 19.3944
R17569 gnd.n4662 gnd.n4660 19.3944
R17570 gnd.n4662 gnd.n2496 19.3944
R17571 gnd.n4674 gnd.n2496 19.3944
R17572 gnd.n4675 gnd.n4674 19.3944
R17573 gnd.n4677 gnd.n4675 19.3944
R17574 gnd.n4678 gnd.n4677 19.3944
R17575 gnd.n4681 gnd.n4678 19.3944
R17576 gnd.n4682 gnd.n4681 19.3944
R17577 gnd.n4687 gnd.n4682 19.3944
R17578 gnd.n4688 gnd.n4687 19.3944
R17579 gnd.n4689 gnd.n4688 19.3944
R17580 gnd.n4689 gnd.n2473 19.3944
R17581 gnd.n4758 gnd.n2473 19.3944
R17582 gnd.n4759 gnd.n4758 19.3944
R17583 gnd.n4760 gnd.n4759 19.3944
R17584 gnd.n4760 gnd.n2468 19.3944
R17585 gnd.n4773 gnd.n2468 19.3944
R17586 gnd.n4774 gnd.n4773 19.3944
R17587 gnd.n4776 gnd.n4774 19.3944
R17588 gnd.n4776 gnd.n4775 19.3944
R17589 gnd.n4449 gnd.n2641 19.3944
R17590 gnd.n4449 gnd.n2642 19.3944
R17591 gnd.n2644 gnd.n2642 19.3944
R17592 gnd.n2644 gnd.n2623 19.3944
R17593 gnd.n4469 gnd.n2623 19.3944
R17594 gnd.n4469 gnd.n4468 19.3944
R17595 gnd.n4468 gnd.n4467 19.3944
R17596 gnd.n4467 gnd.n2605 19.3944
R17597 gnd.n4489 gnd.n2605 19.3944
R17598 gnd.n4489 gnd.n4488 19.3944
R17599 gnd.n4488 gnd.n4487 19.3944
R17600 gnd.n4487 gnd.n2586 19.3944
R17601 gnd.n4513 gnd.n2586 19.3944
R17602 gnd.n4513 gnd.n4512 19.3944
R17603 gnd.n4512 gnd.n4511 19.3944
R17604 gnd.n4511 gnd.n4510 19.3944
R17605 gnd.n4510 gnd.n2561 19.3944
R17606 gnd.n4554 gnd.n2561 19.3944
R17607 gnd.n4554 gnd.n4553 19.3944
R17608 gnd.n4553 gnd.n4552 19.3944
R17609 gnd.n4552 gnd.n2543 19.3944
R17610 gnd.n4579 gnd.n2543 19.3944
R17611 gnd.n4579 gnd.n4578 19.3944
R17612 gnd.n4578 gnd.n4577 19.3944
R17613 gnd.n4577 gnd.n4575 19.3944
R17614 gnd.n4575 gnd.n2526 19.3944
R17615 gnd.n4611 gnd.n2526 19.3944
R17616 gnd.n4611 gnd.n4610 19.3944
R17617 gnd.n4610 gnd.n4609 19.3944
R17618 gnd.n4609 gnd.n961 19.3944
R17619 gnd.n6474 gnd.n961 19.3944
R17620 gnd.n6474 gnd.n6473 19.3944
R17621 gnd.n6473 gnd.n6472 19.3944
R17622 gnd.n6472 gnd.n965 19.3944
R17623 gnd.n6462 gnd.n965 19.3944
R17624 gnd.n6462 gnd.n6461 19.3944
R17625 gnd.n6461 gnd.n6460 19.3944
R17626 gnd.n6460 gnd.n984 19.3944
R17627 gnd.n6450 gnd.n984 19.3944
R17628 gnd.n6450 gnd.n6449 19.3944
R17629 gnd.n6449 gnd.n6448 19.3944
R17630 gnd.n6448 gnd.n1004 19.3944
R17631 gnd.n6438 gnd.n1004 19.3944
R17632 gnd.n6438 gnd.n6437 19.3944
R17633 gnd.n6437 gnd.n6436 19.3944
R17634 gnd.n6436 gnd.n1024 19.3944
R17635 gnd.n6426 gnd.n1024 19.3944
R17636 gnd.n6426 gnd.n6425 19.3944
R17637 gnd.n6425 gnd.n6424 19.3944
R17638 gnd.n6424 gnd.n1044 19.3944
R17639 gnd.n6414 gnd.n1044 19.3944
R17640 gnd.n6414 gnd.n6413 19.3944
R17641 gnd.n6413 gnd.n6412 19.3944
R17642 gnd.n6405 gnd.n6404 19.3944
R17643 gnd.n6404 gnd.n1072 19.3944
R17644 gnd.n1074 gnd.n1072 19.3944
R17645 gnd.n6397 gnd.n1074 19.3944
R17646 gnd.n6397 gnd.n6396 19.3944
R17647 gnd.n6396 gnd.n6395 19.3944
R17648 gnd.n6395 gnd.n1081 19.3944
R17649 gnd.n6390 gnd.n1081 19.3944
R17650 gnd.n6390 gnd.n6389 19.3944
R17651 gnd.n6389 gnd.n6388 19.3944
R17652 gnd.n6388 gnd.n1088 19.3944
R17653 gnd.n6383 gnd.n1088 19.3944
R17654 gnd.n6383 gnd.n6382 19.3944
R17655 gnd.n6382 gnd.n6381 19.3944
R17656 gnd.n6381 gnd.n1095 19.3944
R17657 gnd.n6376 gnd.n1095 19.3944
R17658 gnd.n6376 gnd.n6375 19.3944
R17659 gnd.n2338 gnd.n2298 19.3944
R17660 gnd.n2342 gnd.n2298 19.3944
R17661 gnd.n2342 gnd.n2296 19.3944
R17662 gnd.n2348 gnd.n2296 19.3944
R17663 gnd.n2348 gnd.n2294 19.3944
R17664 gnd.n2352 gnd.n2294 19.3944
R17665 gnd.n2352 gnd.n2292 19.3944
R17666 gnd.n2358 gnd.n2292 19.3944
R17667 gnd.n2358 gnd.n2290 19.3944
R17668 gnd.n2362 gnd.n2290 19.3944
R17669 gnd.n2362 gnd.n2288 19.3944
R17670 gnd.n2368 gnd.n2288 19.3944
R17671 gnd.n2368 gnd.n2286 19.3944
R17672 gnd.n2372 gnd.n2286 19.3944
R17673 gnd.n2372 gnd.n2284 19.3944
R17674 gnd.n2378 gnd.n2284 19.3944
R17675 gnd.n2378 gnd.n2282 19.3944
R17676 gnd.n2382 gnd.n2282 19.3944
R17677 gnd.n2311 gnd.n1117 19.3944
R17678 gnd.n2318 gnd.n2311 19.3944
R17679 gnd.n2318 gnd.n2308 19.3944
R17680 gnd.n2322 gnd.n2308 19.3944
R17681 gnd.n2322 gnd.n2306 19.3944
R17682 gnd.n2328 gnd.n2306 19.3944
R17683 gnd.n2328 gnd.n2304 19.3944
R17684 gnd.n2332 gnd.n2304 19.3944
R17685 gnd.n6373 gnd.n1104 19.3944
R17686 gnd.n6368 gnd.n1104 19.3944
R17687 gnd.n6368 gnd.n6367 19.3944
R17688 gnd.n6367 gnd.n6366 19.3944
R17689 gnd.n6366 gnd.n1111 19.3944
R17690 gnd.n6361 gnd.n1111 19.3944
R17691 gnd.n6361 gnd.n6360 19.3944
R17692 gnd.n4453 gnd.n2634 19.3944
R17693 gnd.n4453 gnd.n2632 19.3944
R17694 gnd.n4457 gnd.n2632 19.3944
R17695 gnd.n4457 gnd.n2615 19.3944
R17696 gnd.n4473 gnd.n2615 19.3944
R17697 gnd.n4473 gnd.n2613 19.3944
R17698 gnd.n4477 gnd.n2613 19.3944
R17699 gnd.n4477 gnd.n2598 19.3944
R17700 gnd.n4493 gnd.n2598 19.3944
R17701 gnd.n4493 gnd.n2596 19.3944
R17702 gnd.n4497 gnd.n2596 19.3944
R17703 gnd.n4497 gnd.n2578 19.3944
R17704 gnd.n4517 gnd.n2578 19.3944
R17705 gnd.n4517 gnd.n2576 19.3944
R17706 gnd.n4523 gnd.n2576 19.3944
R17707 gnd.n4523 gnd.n4522 19.3944
R17708 gnd.n4522 gnd.n2554 19.3944
R17709 gnd.n4558 gnd.n2554 19.3944
R17710 gnd.n4558 gnd.n2552 19.3944
R17711 gnd.n4563 gnd.n2552 19.3944
R17712 gnd.n4563 gnd.n4562 19.3944
R17713 gnd.n4562 gnd.n2539 19.3944
R17714 gnd.n4583 gnd.n944 19.3944
R17715 gnd.n6481 gnd.n944 19.3944
R17716 gnd.n2519 gnd.n945 19.3944
R17717 gnd.n4617 gnd.n4616 19.3944
R17718 gnd.n6478 gnd.n952 19.3944
R17719 gnd.n6478 gnd.n953 19.3944
R17720 gnd.n6468 gnd.n953 19.3944
R17721 gnd.n6468 gnd.n6467 19.3944
R17722 gnd.n6467 gnd.n6466 19.3944
R17723 gnd.n6466 gnd.n974 19.3944
R17724 gnd.n6456 gnd.n974 19.3944
R17725 gnd.n6456 gnd.n6455 19.3944
R17726 gnd.n6455 gnd.n6454 19.3944
R17727 gnd.n6454 gnd.n995 19.3944
R17728 gnd.n6444 gnd.n995 19.3944
R17729 gnd.n6444 gnd.n6443 19.3944
R17730 gnd.n6443 gnd.n6442 19.3944
R17731 gnd.n6442 gnd.n1014 19.3944
R17732 gnd.n6432 gnd.n1014 19.3944
R17733 gnd.n6432 gnd.n6431 19.3944
R17734 gnd.n6431 gnd.n6430 19.3944
R17735 gnd.n6430 gnd.n1035 19.3944
R17736 gnd.n6420 gnd.n1035 19.3944
R17737 gnd.n6420 gnd.n6419 19.3944
R17738 gnd.n6419 gnd.n6418 19.3944
R17739 gnd.n6418 gnd.n1055 19.3944
R17740 gnd.n6408 gnd.n1055 19.3944
R17741 gnd.n6654 gnd.n770 19.3944
R17742 gnd.n6648 gnd.n770 19.3944
R17743 gnd.n6648 gnd.n6647 19.3944
R17744 gnd.n6647 gnd.n6646 19.3944
R17745 gnd.n6646 gnd.n777 19.3944
R17746 gnd.n6640 gnd.n777 19.3944
R17747 gnd.n6640 gnd.n6639 19.3944
R17748 gnd.n6639 gnd.n6638 19.3944
R17749 gnd.n6638 gnd.n785 19.3944
R17750 gnd.n6632 gnd.n785 19.3944
R17751 gnd.n6632 gnd.n6631 19.3944
R17752 gnd.n6631 gnd.n6630 19.3944
R17753 gnd.n6630 gnd.n793 19.3944
R17754 gnd.n6624 gnd.n793 19.3944
R17755 gnd.n6624 gnd.n6623 19.3944
R17756 gnd.n6623 gnd.n6622 19.3944
R17757 gnd.n6622 gnd.n801 19.3944
R17758 gnd.n6616 gnd.n801 19.3944
R17759 gnd.n6616 gnd.n6615 19.3944
R17760 gnd.n6615 gnd.n6614 19.3944
R17761 gnd.n6614 gnd.n809 19.3944
R17762 gnd.n6608 gnd.n809 19.3944
R17763 gnd.n6608 gnd.n6607 19.3944
R17764 gnd.n6607 gnd.n6606 19.3944
R17765 gnd.n6606 gnd.n817 19.3944
R17766 gnd.n6600 gnd.n817 19.3944
R17767 gnd.n6600 gnd.n6599 19.3944
R17768 gnd.n6599 gnd.n6598 19.3944
R17769 gnd.n6598 gnd.n825 19.3944
R17770 gnd.n6592 gnd.n825 19.3944
R17771 gnd.n6592 gnd.n6591 19.3944
R17772 gnd.n6591 gnd.n6590 19.3944
R17773 gnd.n6590 gnd.n833 19.3944
R17774 gnd.n6584 gnd.n833 19.3944
R17775 gnd.n6584 gnd.n6583 19.3944
R17776 gnd.n6583 gnd.n6582 19.3944
R17777 gnd.n6582 gnd.n841 19.3944
R17778 gnd.n6576 gnd.n841 19.3944
R17779 gnd.n6576 gnd.n6575 19.3944
R17780 gnd.n6575 gnd.n6574 19.3944
R17781 gnd.n6574 gnd.n849 19.3944
R17782 gnd.n6568 gnd.n849 19.3944
R17783 gnd.n6568 gnd.n6567 19.3944
R17784 gnd.n6567 gnd.n6566 19.3944
R17785 gnd.n6566 gnd.n857 19.3944
R17786 gnd.n6560 gnd.n857 19.3944
R17787 gnd.n6560 gnd.n6559 19.3944
R17788 gnd.n6559 gnd.n6558 19.3944
R17789 gnd.n6558 gnd.n865 19.3944
R17790 gnd.n6552 gnd.n865 19.3944
R17791 gnd.n6552 gnd.n6551 19.3944
R17792 gnd.n6551 gnd.n6550 19.3944
R17793 gnd.n6550 gnd.n873 19.3944
R17794 gnd.n6544 gnd.n873 19.3944
R17795 gnd.n6544 gnd.n6543 19.3944
R17796 gnd.n6543 gnd.n6542 19.3944
R17797 gnd.n6542 gnd.n881 19.3944
R17798 gnd.n6536 gnd.n881 19.3944
R17799 gnd.n6536 gnd.n6535 19.3944
R17800 gnd.n6535 gnd.n6534 19.3944
R17801 gnd.n6534 gnd.n889 19.3944
R17802 gnd.n6528 gnd.n889 19.3944
R17803 gnd.n6528 gnd.n6527 19.3944
R17804 gnd.n6527 gnd.n6526 19.3944
R17805 gnd.n6526 gnd.n897 19.3944
R17806 gnd.n6520 gnd.n897 19.3944
R17807 gnd.n6520 gnd.n6519 19.3944
R17808 gnd.n6519 gnd.n6518 19.3944
R17809 gnd.n6518 gnd.n905 19.3944
R17810 gnd.n6512 gnd.n905 19.3944
R17811 gnd.n6512 gnd.n6511 19.3944
R17812 gnd.n6511 gnd.n6510 19.3944
R17813 gnd.n6510 gnd.n913 19.3944
R17814 gnd.n6504 gnd.n913 19.3944
R17815 gnd.n6504 gnd.n6503 19.3944
R17816 gnd.n6503 gnd.n6502 19.3944
R17817 gnd.n6502 gnd.n921 19.3944
R17818 gnd.n6496 gnd.n921 19.3944
R17819 gnd.n6496 gnd.n6495 19.3944
R17820 gnd.n6495 gnd.n6494 19.3944
R17821 gnd.n6494 gnd.n929 19.3944
R17822 gnd.n6488 gnd.n929 19.3944
R17823 gnd.n6488 gnd.n6487 19.3944
R17824 gnd.n6487 gnd.n6486 19.3944
R17825 gnd.n2268 gnd.n2267 19.3944
R17826 gnd.n2267 gnd.n2266 19.3944
R17827 gnd.n2266 gnd.n2222 19.3944
R17828 gnd.n2262 gnd.n2222 19.3944
R17829 gnd.n2262 gnd.n2261 19.3944
R17830 gnd.n2261 gnd.n2260 19.3944
R17831 gnd.n2260 gnd.n2226 19.3944
R17832 gnd.n2256 gnd.n2226 19.3944
R17833 gnd.n2256 gnd.n2255 19.3944
R17834 gnd.n2255 gnd.n2254 19.3944
R17835 gnd.n2254 gnd.n2230 19.3944
R17836 gnd.n2250 gnd.n2230 19.3944
R17837 gnd.n2250 gnd.n2249 19.3944
R17838 gnd.n2249 gnd.n2248 19.3944
R17839 gnd.n2248 gnd.n2234 19.3944
R17840 gnd.n2244 gnd.n2234 19.3944
R17841 gnd.n2244 gnd.n2243 19.3944
R17842 gnd.n2243 gnd.n2242 19.3944
R17843 gnd.n2242 gnd.n2237 19.3944
R17844 gnd.n2237 gnd.n2123 19.3944
R17845 gnd.n2123 gnd.n2121 19.3944
R17846 gnd.n4979 gnd.n2121 19.3944
R17847 gnd.n4980 gnd.n4979 19.3944
R17848 gnd.n4980 gnd.n2119 19.3944
R17849 gnd.n4984 gnd.n2119 19.3944
R17850 gnd.n4985 gnd.n4984 19.3944
R17851 gnd.n4988 gnd.n4985 19.3944
R17852 gnd.n4988 gnd.n2116 19.3944
R17853 gnd.n5008 gnd.n2116 19.3944
R17854 gnd.n5008 gnd.n2117 19.3944
R17855 gnd.n5004 gnd.n2117 19.3944
R17856 gnd.n5004 gnd.n5003 19.3944
R17857 gnd.n5003 gnd.n5002 19.3944
R17858 gnd.n5002 gnd.n4994 19.3944
R17859 gnd.n4998 gnd.n4994 19.3944
R17860 gnd.n4998 gnd.n4997 19.3944
R17861 gnd.n4997 gnd.n2069 19.3944
R17862 gnd.n5107 gnd.n2069 19.3944
R17863 gnd.n5107 gnd.n2066 19.3944
R17864 gnd.n5112 gnd.n2066 19.3944
R17865 gnd.n5112 gnd.n2067 19.3944
R17866 gnd.n2067 gnd.n2044 19.3944
R17867 gnd.n5139 gnd.n2044 19.3944
R17868 gnd.n5139 gnd.n2041 19.3944
R17869 gnd.n5167 gnd.n2041 19.3944
R17870 gnd.n5167 gnd.n2042 19.3944
R17871 gnd.n5163 gnd.n2042 19.3944
R17872 gnd.n5163 gnd.n5162 19.3944
R17873 gnd.n5162 gnd.n5161 19.3944
R17874 gnd.n5161 gnd.n5146 19.3944
R17875 gnd.n5157 gnd.n5146 19.3944
R17876 gnd.n5157 gnd.n5156 19.3944
R17877 gnd.n5156 gnd.n5155 19.3944
R17878 gnd.n5155 gnd.n5150 19.3944
R17879 gnd.n5151 gnd.n5150 19.3944
R17880 gnd.n5151 gnd.n1968 19.3944
R17881 gnd.n5264 gnd.n1968 19.3944
R17882 gnd.n5264 gnd.n1965 19.3944
R17883 gnd.n5298 gnd.n1965 19.3944
R17884 gnd.n5298 gnd.n1966 19.3944
R17885 gnd.n5294 gnd.n1966 19.3944
R17886 gnd.n5294 gnd.n5293 19.3944
R17887 gnd.n5293 gnd.n5292 19.3944
R17888 gnd.n5292 gnd.n5272 19.3944
R17889 gnd.n5288 gnd.n5272 19.3944
R17890 gnd.n5288 gnd.n5287 19.3944
R17891 gnd.n5287 gnd.n5286 19.3944
R17892 gnd.n5286 gnd.n5275 19.3944
R17893 gnd.n5282 gnd.n5275 19.3944
R17894 gnd.n5282 gnd.n5281 19.3944
R17895 gnd.n5281 gnd.n1897 19.3944
R17896 gnd.n5416 gnd.n1897 19.3944
R17897 gnd.n5416 gnd.n1894 19.3944
R17898 gnd.n5431 gnd.n1894 19.3944
R17899 gnd.n5431 gnd.n1895 19.3944
R17900 gnd.n5427 gnd.n1895 19.3944
R17901 gnd.n5427 gnd.n5426 19.3944
R17902 gnd.n5426 gnd.n5425 19.3944
R17903 gnd.n5425 gnd.n5422 19.3944
R17904 gnd.n5422 gnd.n1823 19.3944
R17905 gnd.n5627 gnd.n1823 19.3944
R17906 gnd.n5627 gnd.n1821 19.3944
R17907 gnd.n5631 gnd.n1821 19.3944
R17908 gnd.n5631 gnd.n1811 19.3944
R17909 gnd.n5644 gnd.n1811 19.3944
R17910 gnd.n5644 gnd.n1809 19.3944
R17911 gnd.n5648 gnd.n1809 19.3944
R17912 gnd.n5648 gnd.n1799 19.3944
R17913 gnd.n5661 gnd.n1799 19.3944
R17914 gnd.n5661 gnd.n1797 19.3944
R17915 gnd.n5665 gnd.n1797 19.3944
R17916 gnd.n5665 gnd.n1786 19.3944
R17917 gnd.n5678 gnd.n1786 19.3944
R17918 gnd.n5678 gnd.n1784 19.3944
R17919 gnd.n5682 gnd.n1784 19.3944
R17920 gnd.n5682 gnd.n1775 19.3944
R17921 gnd.n5698 gnd.n1775 19.3944
R17922 gnd.n5698 gnd.n1773 19.3944
R17923 gnd.n5702 gnd.n1773 19.3944
R17924 gnd.n5702 gnd.n1401 19.3944
R17925 gnd.n6146 gnd.n1401 19.3944
R17926 gnd.n6143 gnd.n6142 19.3944
R17927 gnd.n6142 gnd.n6141 19.3944
R17928 gnd.n6141 gnd.n1406 19.3944
R17929 gnd.n6137 gnd.n1406 19.3944
R17930 gnd.n6137 gnd.n6136 19.3944
R17931 gnd.n6136 gnd.n6135 19.3944
R17932 gnd.n6135 gnd.n1411 19.3944
R17933 gnd.n6130 gnd.n1411 19.3944
R17934 gnd.n6130 gnd.n6129 19.3944
R17935 gnd.n6129 gnd.n1416 19.3944
R17936 gnd.n6122 gnd.n1416 19.3944
R17937 gnd.n6122 gnd.n6121 19.3944
R17938 gnd.n6121 gnd.n1425 19.3944
R17939 gnd.n6114 gnd.n1425 19.3944
R17940 gnd.n6114 gnd.n6113 19.3944
R17941 gnd.n6113 gnd.n1433 19.3944
R17942 gnd.n6106 gnd.n1433 19.3944
R17943 gnd.n6106 gnd.n6105 19.3944
R17944 gnd.n6105 gnd.n1441 19.3944
R17945 gnd.n6098 gnd.n1441 19.3944
R17946 gnd.n6098 gnd.n6097 19.3944
R17947 gnd.n6097 gnd.n1449 19.3944
R17948 gnd.n6090 gnd.n1449 19.3944
R17949 gnd.n6090 gnd.n6089 19.3944
R17950 gnd.n1761 gnd.n1740 19.3944
R17951 gnd.n5731 gnd.n1740 19.3944
R17952 gnd.n5731 gnd.n5730 19.3944
R17953 gnd.n5177 gnd.n2033 19.1199
R17954 gnd.n5252 gnd.n5250 19.1199
R17955 gnd.n5414 gnd.n1900 19.1199
R17956 gnd.n3513 gnd.t344 18.8012
R17957 gnd.n3498 gnd.t155 18.8012
R17958 gnd.n6289 gnd.n6288 18.5761
R17959 gnd.n5543 gnd.n5542 18.5761
R17960 gnd.n3357 gnd.n3356 18.4825
R17961 gnd.n4613 gnd.n2520 18.4825
R17962 gnd.n4620 gnd.n4619 18.4825
R17963 gnd.n4649 gnd.n2506 18.4825
R17964 gnd.n4657 gnd.n958 18.4825
R17965 gnd.n6470 gnd.n967 18.4825
R17966 gnd.n4664 gnd.n2500 18.4825
R17967 gnd.n6464 gnd.n976 18.4825
R17968 gnd.n6458 gnd.n986 18.4825
R17969 gnd.n4708 gnd.n989 18.4825
R17970 gnd.n4679 gnd.n999 18.4825
R17971 gnd.n6446 gnd.n1006 18.4825
R17972 gnd.n4685 gnd.n4684 18.4825
R17973 gnd.n6440 gnd.n1016 18.4825
R17974 gnd.n6434 gnd.n1026 18.4825
R17975 gnd.n4756 gnd.n1029 18.4825
R17976 gnd.n4762 gnd.n1039 18.4825
R17977 gnd.n6422 gnd.n1046 18.4825
R17978 gnd.n4771 gnd.n1049 18.4825
R17979 gnd.n6416 gnd.n1057 18.4825
R17980 gnd.n4778 gnd.n2467 18.4825
R17981 gnd.n6410 gnd.n1065 18.4825
R17982 gnd.n5959 gnd.n1577 18.4825
R17983 gnd.n5776 gnd.n5775 18.4825
R17984 gnd.n5951 gnd.n1586 18.4825
R17985 gnd.n5736 gnd.n1599 18.4825
R17986 gnd.n5945 gnd.n1602 18.4825
R17987 gnd.n5743 gnd.n1612 18.4825
R17988 gnd.n5749 gnd.n1622 18.4825
R17989 gnd.n5933 gnd.n1625 18.4825
R17990 gnd.n5927 gnd.n1635 18.4825
R17991 gnd.n5821 gnd.n5820 18.4825
R17992 gnd.n5921 gnd.n1645 18.4825
R17993 gnd.n5829 gnd.n1652 18.4825
R17994 gnd.n5836 gnd.n1662 18.4825
R17995 gnd.n5909 gnd.n1665 18.4825
R17996 gnd.n5903 gnd.n1675 18.4825
R17997 gnd.n5875 gnd.n5874 18.4825
R17998 gnd.n5897 gnd.n1685 18.4825
R17999 gnd.n5858 gnd.n1692 18.4825
R18000 gnd.n5887 gnd.n5886 18.4825
R18001 gnd.n1699 gnd.n381 18.4825
R18002 gnd.n7295 gnd.n375 18.4825
R18003 gnd.n6028 gnd.n6027 18.4247
R18004 gnd.n6360 gnd.n6359 18.4247
R18005 gnd.n6086 gnd.n6085 18.2308
R18006 gnd.n4797 gnd.n4796 18.2308
R18007 gnd.n7406 gnd.n7405 18.2308
R18008 gnd.n4288 gnd.n4248 18.2308
R18009 gnd.t345 gnd.n3037 18.1639
R18010 gnd.n2108 gnd.n1302 17.8452
R18011 gnd.n5188 gnd.n5187 17.8452
R18012 gnd.n5223 gnd.n1999 17.8452
R18013 gnd.n5404 gnd.n5403 17.8452
R18014 gnd.n3065 gnd.t347 17.5266
R18015 gnd.n2620 gnd.t213 17.5266
R18016 gnd.n6428 gnd.t196 17.5266
R18017 gnd.n5939 gnd.t205 17.5266
R18018 gnd.n7567 gnd.t230 17.5266
R18019 gnd.t173 gnd.n5094 17.2079
R18020 gnd.n5339 gnd.t3 17.2079
R18021 gnd.n5434 gnd.t63 17.2079
R18022 gnd.n3464 gnd.t357 16.8893
R18023 gnd.n3741 gnd.n3740 16.8893
R18024 gnd.n2583 gnd.t228 16.8893
R18025 gnd.n6484 gnd.n6483 16.8893
R18026 gnd.n6452 gnd.t255 16.8893
R18027 gnd.t362 gnd.n1125 16.8893
R18028 gnd.n5915 gnd.t186 16.8893
R18029 gnd.n7623 gnd.n90 16.8893
R18030 gnd.n7591 gnd.t198 16.8893
R18031 gnd.n6010 gnd.n6007 16.6793
R18032 gnd.n7478 gnd.n7477 16.6793
R18033 gnd.n4368 gnd.n4365 16.6793
R18034 gnd.n2332 gnd.n2302 16.6793
R18035 gnd.n5035 gnd.n2104 16.5706
R18036 gnd.n5087 gnd.t161 16.5706
R18037 gnd.n2017 gnd.n2012 16.5706
R18038 gnd.n5215 gnd.n5213 16.5706
R18039 gnd.n5328 gnd.t4 16.5706
R18040 gnd.n5278 gnd.n1921 16.5706
R18041 gnd.n3292 gnd.t122 16.2519
R18042 gnd.n2992 gnd.t351 16.2519
R18043 gnd.n4581 gnd.t239 16.2519
R18044 gnd.n6476 gnd.t192 16.2519
R18045 gnd.t41 gnd.t165 16.2519
R18046 gnd.n5891 gnd.t250 16.2519
R18047 gnd.n7615 gnd.t203 16.2519
R18048 gnd.t162 gnd.n2055 15.9333
R18049 gnd.n5309 gnd.t154 15.9333
R18050 gnd.n3980 gnd.n3978 15.6674
R18051 gnd.n3948 gnd.n3946 15.6674
R18052 gnd.n3916 gnd.n3914 15.6674
R18053 gnd.n3885 gnd.n3883 15.6674
R18054 gnd.n3853 gnd.n3851 15.6674
R18055 gnd.n3821 gnd.n3819 15.6674
R18056 gnd.n3789 gnd.n3787 15.6674
R18057 gnd.n3758 gnd.n3756 15.6674
R18058 gnd.n3283 gnd.t122 15.6146
R18059 gnd.t106 gnd.n2730 15.6146
R18060 gnd.t84 gnd.n2731 15.6146
R18061 gnd.n4585 gnd.t239 15.6146
R18062 gnd.n7357 gnd.t203 15.6146
R18063 gnd.n5967 gnd.n5962 15.3217
R18064 gnd.n7438 gnd.n315 15.3217
R18065 gnd.n4326 gnd.n2647 15.3217
R18066 gnd.n2387 gnd.n2280 15.3217
R18067 gnd.n5036 gnd.n5035 15.296
R18068 gnd.n2098 gnd.n2091 15.296
R18069 gnd.t2 gnd.n2046 15.296
R18070 gnd.n2018 gnd.n2017 15.296
R18071 gnd.n5213 gnd.n2008 15.296
R18072 gnd.n5241 gnd.t139 15.296
R18073 gnd.n5359 gnd.n1925 15.296
R18074 gnd.n5279 gnd.n5278 15.296
R18075 gnd.n5459 gnd.n5458 15.0827
R18076 gnd.n1169 gnd.n1164 15.0481
R18077 gnd.n5469 gnd.n5468 15.0481
R18078 gnd.n3651 gnd.t348 14.9773
R18079 gnd.n4525 gnd.t228 14.9773
R18080 gnd.n6484 gnd.n938 14.9773
R18081 gnd.n4975 gnd.t362 14.9773
R18082 gnd.t91 gnd.t180 14.9773
R18083 gnd.n5625 gnd.t180 14.9773
R18084 gnd.n368 gnd.n90 14.9773
R18085 gnd.t198 gnd.n136 14.9773
R18086 gnd.n5170 gnd.t8 14.6587
R18087 gnd.n5235 gnd.t148 14.6587
R18088 gnd.t133 gnd.n2773 14.34
R18089 gnd.n3729 gnd.t346 14.34
R18090 gnd.n4479 gnd.t213 14.34
R18091 gnd.t230 gnd.n174 14.34
R18092 gnd.n6259 gnd.n1302 14.0214
R18093 gnd.n5094 gnd.n2081 14.0214
R18094 gnd.n5065 gnd.t5 14.0214
R18095 gnd.n5188 gnd.n2023 14.0214
R18096 gnd.n1999 gnd.n1993 14.0214
R18097 gnd.n5230 gnd.t140 14.0214
R18098 gnd.n5340 gnd.n5339 14.0214
R18099 gnd.n5403 gnd.n1911 14.0214
R18100 gnd.n3439 gnd.t178 13.7027
R18101 gnd.n5061 gnd.t176 13.7027
R18102 gnd.n5262 gnd.t149 13.7027
R18103 gnd.n3149 gnd.n3148 13.5763
R18104 gnd.n4094 gnd.n2687 13.5763
R18105 gnd.n3357 gnd.n3095 13.384
R18106 gnd.n4600 gnd.n2520 13.384
R18107 gnd.n4613 gnd.n2523 13.384
R18108 gnd.n4620 gnd.n2516 13.384
R18109 gnd.n4619 gnd.n2506 13.384
R18110 gnd.n4649 gnd.n4648 13.384
R18111 gnd.n6476 gnd.n958 13.384
R18112 gnd.n4657 gnd.n967 13.384
R18113 gnd.n4664 gnd.n976 13.384
R18114 gnd.n6464 gnd.n979 13.384
R18115 gnd.n4672 gnd.n986 13.384
R18116 gnd.n6458 gnd.n989 13.384
R18117 gnd.n4709 gnd.n4708 13.384
R18118 gnd.n6452 gnd.n999 13.384
R18119 gnd.n4679 gnd.n1006 13.384
R18120 gnd.n4685 gnd.n1016 13.384
R18121 gnd.n6440 gnd.n1019 13.384
R18122 gnd.n4691 gnd.n1026 13.384
R18123 gnd.n6434 gnd.n1029 13.384
R18124 gnd.n4756 gnd.n4755 13.384
R18125 gnd.n6428 gnd.n1039 13.384
R18126 gnd.n4762 gnd.n1046 13.384
R18127 gnd.n6422 gnd.n1049 13.384
R18128 gnd.n4771 gnd.n1057 13.384
R18129 gnd.n4778 gnd.n1065 13.384
R18130 gnd.n6410 gnd.n1068 13.384
R18131 gnd.n5194 gnd.t145 13.384
R18132 gnd.n5200 gnd.t137 13.384
R18133 gnd.n5959 gnd.n1575 13.384
R18134 gnd.n5775 gnd.n1577 13.384
R18135 gnd.n5736 gnd.n1586 13.384
R18136 gnd.n5945 gnd.n1599 13.384
R18137 gnd.n5743 gnd.n1602 13.384
R18138 gnd.n5939 gnd.n1612 13.384
R18139 gnd.n5749 gnd.n5748 13.384
R18140 gnd.n5933 gnd.n1622 13.384
R18141 gnd.n5758 gnd.n1625 13.384
R18142 gnd.n5927 gnd.n1632 13.384
R18143 gnd.n5821 gnd.n1635 13.384
R18144 gnd.n5829 gnd.n1645 13.384
R18145 gnd.n5915 gnd.n1652 13.384
R18146 gnd.n5836 gnd.n1715 13.384
R18147 gnd.n5909 gnd.n1662 13.384
R18148 gnd.n5844 gnd.n1665 13.384
R18149 gnd.n5903 gnd.n1672 13.384
R18150 gnd.n5874 gnd.n1675 13.384
R18151 gnd.n5858 gnd.n1685 13.384
R18152 gnd.n5891 gnd.n1692 13.384
R18153 gnd.n5887 gnd.n1696 13.384
R18154 gnd.n5886 gnd.n1699 13.384
R18155 gnd.n7299 gnd.n381 13.384
R18156 gnd.n7295 gnd.n7293 13.384
R18157 gnd.n7308 gnd.n375 13.384
R18158 gnd.n1180 gnd.n1161 13.1884
R18159 gnd.n1175 gnd.n1174 13.1884
R18160 gnd.n1174 gnd.n1173 13.1884
R18161 gnd.n5462 gnd.n5457 13.1884
R18162 gnd.n5463 gnd.n5462 13.1884
R18163 gnd.n1176 gnd.n1163 13.146
R18164 gnd.n1172 gnd.n1163 13.146
R18165 gnd.n5461 gnd.n5460 13.146
R18166 gnd.n5461 gnd.n5456 13.146
R18167 gnd.n2523 gnd.t211 13.0654
R18168 gnd.n7293 gnd.t220 13.0654
R18169 gnd.n3981 gnd.n3977 12.8005
R18170 gnd.n3949 gnd.n3945 12.8005
R18171 gnd.n3917 gnd.n3913 12.8005
R18172 gnd.n3886 gnd.n3882 12.8005
R18173 gnd.n3854 gnd.n3850 12.8005
R18174 gnd.n3822 gnd.n3818 12.8005
R18175 gnd.n3790 gnd.n3786 12.8005
R18176 gnd.n3759 gnd.n3755 12.8005
R18177 gnd.n6265 gnd.n1289 12.7467
R18178 gnd.n5169 gnd.n2033 12.7467
R18179 gnd.n5250 gnd.n1980 12.7467
R18180 gnd.n5370 gnd.n1900 12.7467
R18181 gnd.t243 gnd.n979 12.4281
R18182 gnd.t0 gnd.n2169 12.4281
R18183 gnd.n1789 gnd.t171 12.4281
R18184 gnd.t182 gnd.n1672 12.4281
R18185 gnd.n3148 gnd.n3143 12.4126
R18186 gnd.n4097 gnd.n4094 12.4126
R18187 gnd.n6352 gnd.n6289 12.1761
R18188 gnd.n5542 gnd.n5541 12.1761
R18189 gnd.n4741 gnd.n1073 12.1094
R18190 gnd.n6080 gnd.n1507 12.1094
R18191 gnd.n3985 gnd.n3984 12.0247
R18192 gnd.n3953 gnd.n3952 12.0247
R18193 gnd.n3921 gnd.n3920 12.0247
R18194 gnd.n3890 gnd.n3889 12.0247
R18195 gnd.n3858 gnd.n3857 12.0247
R18196 gnd.n3826 gnd.n3825 12.0247
R18197 gnd.n3794 gnd.n3793 12.0247
R18198 gnd.n3763 gnd.n3762 12.0247
R18199 gnd.t262 gnd.n1019 11.7908
R18200 gnd.t209 gnd.n1632 11.7908
R18201 gnd.n6272 gnd.n1275 11.4721
R18202 gnd.n5127 gnd.n2055 11.4721
R18203 gnd.n5137 gnd.n2047 11.4721
R18204 gnd.n5243 gnd.n5242 11.4721
R18205 gnd.n5310 gnd.n5309 11.4721
R18206 gnd.n5442 gnd.n1886 11.4721
R18207 gnd.n5450 gnd.n1880 11.4721
R18208 gnd.n5546 gnd.t52 11.4721
R18209 gnd.n3988 gnd.n3975 11.249
R18210 gnd.n3956 gnd.n3943 11.249
R18211 gnd.n3924 gnd.n3911 11.249
R18212 gnd.n3893 gnd.n3880 11.249
R18213 gnd.n3861 gnd.n3848 11.249
R18214 gnd.n3829 gnd.n3816 11.249
R18215 gnd.n3797 gnd.n3784 11.249
R18216 gnd.n3766 gnd.n3753 11.249
R18217 gnd.n3427 gnd.t178 11.1535
R18218 gnd.n5087 gnd.t360 11.1535
R18219 gnd.n5328 gnd.t174 11.1535
R18220 gnd.n5970 gnd.n5967 10.6672
R18221 gnd.n7443 gnd.n315 10.6672
R18222 gnd.n4328 gnd.n4326 10.6672
R18223 gnd.n2382 gnd.n2280 10.6672
R18224 gnd.n5612 gnd.n5611 10.6151
R18225 gnd.n5611 gnd.n5608 10.6151
R18226 gnd.n5606 gnd.n5603 10.6151
R18227 gnd.n5603 gnd.n5602 10.6151
R18228 gnd.n5602 gnd.n5599 10.6151
R18229 gnd.n5599 gnd.n5598 10.6151
R18230 gnd.n5598 gnd.n5595 10.6151
R18231 gnd.n5595 gnd.n5594 10.6151
R18232 gnd.n5594 gnd.n5591 10.6151
R18233 gnd.n5591 gnd.n5590 10.6151
R18234 gnd.n5590 gnd.n5587 10.6151
R18235 gnd.n5587 gnd.n5586 10.6151
R18236 gnd.n5586 gnd.n5583 10.6151
R18237 gnd.n5583 gnd.n5582 10.6151
R18238 gnd.n5582 gnd.n5579 10.6151
R18239 gnd.n5579 gnd.n5578 10.6151
R18240 gnd.n5578 gnd.n5575 10.6151
R18241 gnd.n5575 gnd.n5574 10.6151
R18242 gnd.n5574 gnd.n5571 10.6151
R18243 gnd.n5571 gnd.n5570 10.6151
R18244 gnd.n5570 gnd.n5567 10.6151
R18245 gnd.n5567 gnd.n5566 10.6151
R18246 gnd.n5566 gnd.n5563 10.6151
R18247 gnd.n5563 gnd.n5562 10.6151
R18248 gnd.n5562 gnd.n5559 10.6151
R18249 gnd.n5559 gnd.n5558 10.6151
R18250 gnd.n5558 gnd.n5555 10.6151
R18251 gnd.n5555 gnd.n5554 10.6151
R18252 gnd.n5554 gnd.n5551 10.6151
R18253 gnd.n5551 gnd.n5550 10.6151
R18254 gnd.n1269 gnd.n1268 10.6151
R18255 gnd.n1271 gnd.n1269 10.6151
R18256 gnd.n1272 gnd.n1271 10.6151
R18257 gnd.n6276 gnd.n1272 10.6151
R18258 gnd.n6276 gnd.n6275 10.6151
R18259 gnd.n6275 gnd.n6274 10.6151
R18260 gnd.n6274 gnd.n1273 10.6151
R18261 gnd.n2112 gnd.n1273 10.6151
R18262 gnd.n2113 gnd.n2112 10.6151
R18263 gnd.n2114 gnd.n2113 10.6151
R18264 gnd.n2114 gnd.n2110 10.6151
R18265 gnd.n5019 gnd.n2110 10.6151
R18266 gnd.n5020 gnd.n5019 10.6151
R18267 gnd.n5026 gnd.n5020 10.6151
R18268 gnd.n5026 gnd.n5025 10.6151
R18269 gnd.n5025 gnd.n5024 10.6151
R18270 gnd.n5024 gnd.n5022 10.6151
R18271 gnd.n5022 gnd.n5021 10.6151
R18272 gnd.n5021 gnd.n2088 10.6151
R18273 gnd.n5054 gnd.n2088 10.6151
R18274 gnd.n5055 gnd.n5054 10.6151
R18275 gnd.n5058 gnd.n5055 10.6151
R18276 gnd.n5059 gnd.n5058 10.6151
R18277 gnd.n5083 gnd.n5059 10.6151
R18278 gnd.n5083 gnd.n5082 10.6151
R18279 gnd.n5082 gnd.n5081 10.6151
R18280 gnd.n5081 gnd.n5080 10.6151
R18281 gnd.n5080 gnd.n5078 10.6151
R18282 gnd.n5078 gnd.n5077 10.6151
R18283 gnd.n5077 gnd.n5060 10.6151
R18284 gnd.n5073 gnd.n5060 10.6151
R18285 gnd.n5073 gnd.n5072 10.6151
R18286 gnd.n5072 gnd.n5071 10.6151
R18287 gnd.n5071 gnd.n5070 10.6151
R18288 gnd.n5070 gnd.n5068 10.6151
R18289 gnd.n5068 gnd.n5067 10.6151
R18290 gnd.n5067 gnd.n5064 10.6151
R18291 gnd.n5064 gnd.n2015 10.6151
R18292 gnd.n5196 gnd.n2015 10.6151
R18293 gnd.n5197 gnd.n5196 10.6151
R18294 gnd.n5205 gnd.n5197 10.6151
R18295 gnd.n5205 gnd.n5204 10.6151
R18296 gnd.n5204 gnd.n5203 10.6151
R18297 gnd.n5203 gnd.n5202 10.6151
R18298 gnd.n5202 gnd.n5199 10.6151
R18299 gnd.n5199 gnd.n5198 10.6151
R18300 gnd.n5198 gnd.n1991 10.6151
R18301 gnd.n5233 gnd.n1991 10.6151
R18302 gnd.n5234 gnd.n5233 10.6151
R18303 gnd.n5237 gnd.n5234 10.6151
R18304 gnd.n5238 gnd.n5237 10.6151
R18305 gnd.n5239 gnd.n5238 10.6151
R18306 gnd.n5239 gnd.n1961 10.6151
R18307 gnd.n5303 gnd.n1961 10.6151
R18308 gnd.n5304 gnd.n5303 10.6151
R18309 gnd.n5307 gnd.n5304 10.6151
R18310 gnd.n5307 gnd.n5306 10.6151
R18311 gnd.n5306 gnd.n5305 10.6151
R18312 gnd.n5305 gnd.n1944 10.6151
R18313 gnd.n5331 gnd.n1944 10.6151
R18314 gnd.n5332 gnd.n5331 10.6151
R18315 gnd.n5337 gnd.n5332 10.6151
R18316 gnd.n5337 gnd.n5336 10.6151
R18317 gnd.n5336 gnd.n5335 10.6151
R18318 gnd.n5335 gnd.n5333 10.6151
R18319 gnd.n5333 gnd.n1918 10.6151
R18320 gnd.n5367 gnd.n1918 10.6151
R18321 gnd.n5368 gnd.n5367 10.6151
R18322 gnd.n5390 gnd.n5368 10.6151
R18323 gnd.n5390 gnd.n5389 10.6151
R18324 gnd.n5389 gnd.n5388 10.6151
R18325 gnd.n5388 gnd.n5387 10.6151
R18326 gnd.n5387 gnd.n5369 10.6151
R18327 gnd.n5382 gnd.n5369 10.6151
R18328 gnd.n5382 gnd.n5381 10.6151
R18329 gnd.n5381 gnd.n5380 10.6151
R18330 gnd.n5380 gnd.n5379 10.6151
R18331 gnd.n5379 gnd.n5377 10.6151
R18332 gnd.n5377 gnd.n5376 10.6151
R18333 gnd.n5376 gnd.n5374 10.6151
R18334 gnd.n5374 gnd.n5373 10.6151
R18335 gnd.n5373 gnd.n1871 10.6151
R18336 gnd.n1871 gnd.n1869 10.6151
R18337 gnd.n1204 gnd.n1121 10.6151
R18338 gnd.n1207 gnd.n1204 10.6151
R18339 gnd.n1212 gnd.n1209 10.6151
R18340 gnd.n1213 gnd.n1212 10.6151
R18341 gnd.n1216 gnd.n1213 10.6151
R18342 gnd.n1217 gnd.n1216 10.6151
R18343 gnd.n1220 gnd.n1217 10.6151
R18344 gnd.n1221 gnd.n1220 10.6151
R18345 gnd.n1224 gnd.n1221 10.6151
R18346 gnd.n1225 gnd.n1224 10.6151
R18347 gnd.n1228 gnd.n1225 10.6151
R18348 gnd.n1229 gnd.n1228 10.6151
R18349 gnd.n1232 gnd.n1229 10.6151
R18350 gnd.n1233 gnd.n1232 10.6151
R18351 gnd.n1236 gnd.n1233 10.6151
R18352 gnd.n1237 gnd.n1236 10.6151
R18353 gnd.n1240 gnd.n1237 10.6151
R18354 gnd.n1241 gnd.n1240 10.6151
R18355 gnd.n1244 gnd.n1241 10.6151
R18356 gnd.n1245 gnd.n1244 10.6151
R18357 gnd.n1248 gnd.n1245 10.6151
R18358 gnd.n1249 gnd.n1248 10.6151
R18359 gnd.n1252 gnd.n1249 10.6151
R18360 gnd.n1253 gnd.n1252 10.6151
R18361 gnd.n1256 gnd.n1253 10.6151
R18362 gnd.n1257 gnd.n1256 10.6151
R18363 gnd.n1260 gnd.n1257 10.6151
R18364 gnd.n1261 gnd.n1260 10.6151
R18365 gnd.n1264 gnd.n1261 10.6151
R18366 gnd.n1265 gnd.n1264 10.6151
R18367 gnd.n6352 gnd.n6351 10.6151
R18368 gnd.n6351 gnd.n6350 10.6151
R18369 gnd.n6350 gnd.n6349 10.6151
R18370 gnd.n6349 gnd.n6347 10.6151
R18371 gnd.n6347 gnd.n6344 10.6151
R18372 gnd.n6344 gnd.n6343 10.6151
R18373 gnd.n6343 gnd.n6340 10.6151
R18374 gnd.n6340 gnd.n6339 10.6151
R18375 gnd.n6339 gnd.n6336 10.6151
R18376 gnd.n6336 gnd.n6335 10.6151
R18377 gnd.n6335 gnd.n6332 10.6151
R18378 gnd.n6332 gnd.n6331 10.6151
R18379 gnd.n6331 gnd.n6328 10.6151
R18380 gnd.n6328 gnd.n6327 10.6151
R18381 gnd.n6327 gnd.n6324 10.6151
R18382 gnd.n6324 gnd.n6323 10.6151
R18383 gnd.n6323 gnd.n6320 10.6151
R18384 gnd.n6320 gnd.n6319 10.6151
R18385 gnd.n6319 gnd.n6316 10.6151
R18386 gnd.n6316 gnd.n6315 10.6151
R18387 gnd.n6315 gnd.n6312 10.6151
R18388 gnd.n6312 gnd.n6311 10.6151
R18389 gnd.n6311 gnd.n6308 10.6151
R18390 gnd.n6308 gnd.n6307 10.6151
R18391 gnd.n6307 gnd.n6304 10.6151
R18392 gnd.n6304 gnd.n6303 10.6151
R18393 gnd.n6303 gnd.n6300 10.6151
R18394 gnd.n6300 gnd.n6299 10.6151
R18395 gnd.n6296 gnd.n6295 10.6151
R18396 gnd.n6295 gnd.n1122 10.6151
R18397 gnd.n5541 gnd.n5539 10.6151
R18398 gnd.n5539 gnd.n5536 10.6151
R18399 gnd.n5536 gnd.n5535 10.6151
R18400 gnd.n5535 gnd.n5532 10.6151
R18401 gnd.n5532 gnd.n5531 10.6151
R18402 gnd.n5531 gnd.n5528 10.6151
R18403 gnd.n5528 gnd.n5527 10.6151
R18404 gnd.n5527 gnd.n5524 10.6151
R18405 gnd.n5524 gnd.n5523 10.6151
R18406 gnd.n5523 gnd.n5520 10.6151
R18407 gnd.n5520 gnd.n5519 10.6151
R18408 gnd.n5519 gnd.n5516 10.6151
R18409 gnd.n5516 gnd.n5515 10.6151
R18410 gnd.n5515 gnd.n5512 10.6151
R18411 gnd.n5512 gnd.n5511 10.6151
R18412 gnd.n5511 gnd.n5508 10.6151
R18413 gnd.n5508 gnd.n5507 10.6151
R18414 gnd.n5507 gnd.n5504 10.6151
R18415 gnd.n5504 gnd.n5503 10.6151
R18416 gnd.n5503 gnd.n5500 10.6151
R18417 gnd.n5500 gnd.n5499 10.6151
R18418 gnd.n5499 gnd.n5496 10.6151
R18419 gnd.n5496 gnd.n5495 10.6151
R18420 gnd.n5495 gnd.n5492 10.6151
R18421 gnd.n5492 gnd.n5491 10.6151
R18422 gnd.n5491 gnd.n5488 10.6151
R18423 gnd.n5488 gnd.n5487 10.6151
R18424 gnd.n5487 gnd.n5484 10.6151
R18425 gnd.n5482 gnd.n5479 10.6151
R18426 gnd.n5479 gnd.n5478 10.6151
R18427 gnd.n6288 gnd.n6287 10.6151
R18428 gnd.n6287 gnd.n1181 10.6151
R18429 gnd.n1281 gnd.n1181 10.6151
R18430 gnd.n1282 gnd.n1281 10.6151
R18431 gnd.n1283 gnd.n1282 10.6151
R18432 gnd.n6270 gnd.n1283 10.6151
R18433 gnd.n6270 gnd.n6269 10.6151
R18434 gnd.n6269 gnd.n6268 10.6151
R18435 gnd.n6268 gnd.n1284 10.6151
R18436 gnd.n5013 gnd.n1284 10.6151
R18437 gnd.n5014 gnd.n5013 10.6151
R18438 gnd.n5014 gnd.n2106 10.6151
R18439 gnd.n5031 gnd.n2106 10.6151
R18440 gnd.n5032 gnd.n5031 10.6151
R18441 gnd.n5033 gnd.n5032 10.6151
R18442 gnd.n5033 gnd.n2093 10.6151
R18443 gnd.n5047 gnd.n2093 10.6151
R18444 gnd.n5048 gnd.n5047 10.6151
R18445 gnd.n5049 gnd.n5048 10.6151
R18446 gnd.n5049 gnd.n2084 10.6151
R18447 gnd.n5092 gnd.n2084 10.6151
R18448 gnd.n5092 gnd.n5091 10.6151
R18449 gnd.n5091 gnd.n5090 10.6151
R18450 gnd.n5090 gnd.n2085 10.6151
R18451 gnd.n2085 gnd.n2061 10.6151
R18452 gnd.n5117 gnd.n2061 10.6151
R18453 gnd.n5118 gnd.n5117 10.6151
R18454 gnd.n5124 gnd.n5118 10.6151
R18455 gnd.n5124 gnd.n5123 10.6151
R18456 gnd.n5123 gnd.n5122 10.6151
R18457 gnd.n5122 gnd.n5119 10.6151
R18458 gnd.n5119 gnd.n2037 10.6151
R18459 gnd.n5172 gnd.n2037 10.6151
R18460 gnd.n5173 gnd.n5172 10.6151
R18461 gnd.n5174 gnd.n5173 10.6151
R18462 gnd.n5174 gnd.n2020 10.6151
R18463 gnd.n5190 gnd.n2020 10.6151
R18464 gnd.n5191 gnd.n5190 10.6151
R18465 gnd.n5192 gnd.n5191 10.6151
R18466 gnd.n5192 gnd.n2010 10.6151
R18467 gnd.n5209 gnd.n2010 10.6151
R18468 gnd.n5210 gnd.n5209 10.6151
R18469 gnd.n5211 gnd.n5210 10.6151
R18470 gnd.n5211 gnd.n1995 10.6151
R18471 gnd.n5226 gnd.n1995 10.6151
R18472 gnd.n5227 gnd.n5226 10.6151
R18473 gnd.n5228 gnd.n5227 10.6151
R18474 gnd.n5228 gnd.n1983 10.6151
R18475 gnd.n5248 gnd.n1983 10.6151
R18476 gnd.n5248 gnd.n5247 10.6151
R18477 gnd.n5247 gnd.n5246 10.6151
R18478 gnd.n5246 gnd.n1984 10.6151
R18479 gnd.n1988 gnd.n1984 10.6151
R18480 gnd.n1988 gnd.n1987 10.6151
R18481 gnd.n1987 gnd.n1986 10.6151
R18482 gnd.n1986 gnd.n1947 10.6151
R18483 gnd.n5324 gnd.n1947 10.6151
R18484 gnd.n5325 gnd.n5324 10.6151
R18485 gnd.n5326 gnd.n5325 10.6151
R18486 gnd.n5326 gnd.n1939 10.6151
R18487 gnd.n5343 gnd.n1939 10.6151
R18488 gnd.n5344 gnd.n5343 10.6151
R18489 gnd.n5345 gnd.n5344 10.6151
R18490 gnd.n5345 gnd.n1923 10.6151
R18491 gnd.n5361 gnd.n1923 10.6151
R18492 gnd.n5362 gnd.n5361 10.6151
R18493 gnd.n5363 gnd.n5362 10.6151
R18494 gnd.n5363 gnd.n1914 10.6151
R18495 gnd.n5394 gnd.n1914 10.6151
R18496 gnd.n5395 gnd.n5394 10.6151
R18497 gnd.n5401 gnd.n5395 10.6151
R18498 gnd.n5401 gnd.n5400 10.6151
R18499 gnd.n5400 gnd.n5399 10.6151
R18500 gnd.n5399 gnd.n5396 10.6151
R18501 gnd.n5396 gnd.n1890 10.6151
R18502 gnd.n5436 gnd.n1890 10.6151
R18503 gnd.n5437 gnd.n5436 10.6151
R18504 gnd.n5438 gnd.n5437 10.6151
R18505 gnd.n5438 gnd.n1875 10.6151
R18506 gnd.n5453 gnd.n1875 10.6151
R18507 gnd.n5454 gnd.n5453 10.6151
R18508 gnd.n5544 gnd.n5454 10.6151
R18509 gnd.n5544 gnd.n5543 10.6151
R18510 gnd.n3346 gnd.t163 10.5161
R18511 gnd.n2775 gnd.t133 10.5161
R18512 gnd.n3712 gnd.t346 10.5161
R18513 gnd.n5044 gnd.t9 10.5161
R18514 gnd.t159 gnd.n5358 10.5161
R18515 gnd.n3989 gnd.n3973 10.4732
R18516 gnd.n3957 gnd.n3941 10.4732
R18517 gnd.n3925 gnd.n3909 10.4732
R18518 gnd.n3894 gnd.n3878 10.4732
R18519 gnd.n3862 gnd.n3846 10.4732
R18520 gnd.n3830 gnd.n3814 10.4732
R18521 gnd.n3798 gnd.n3782 10.4732
R18522 gnd.n3767 gnd.n3751 10.4732
R18523 gnd.n4941 gnd.n1196 10.1975
R18524 gnd.n1277 gnd.n1275 10.1975
R18525 gnd.t19 gnd.n1289 10.1975
R18526 gnd.n5127 gnd.n5126 10.1975
R18527 gnd.n5137 gnd.n2046 10.1975
R18528 gnd.n5242 gnd.n5241 10.1975
R18529 gnd.n5310 gnd.n1958 10.1975
R18530 gnd.t52 gnd.n1830 10.1975
R18531 gnd.t348 gnd.n2792 9.87883
R18532 gnd.t129 gnd.t135 9.87883
R18533 gnd.n3993 gnd.n3992 9.69747
R18534 gnd.n3961 gnd.n3960 9.69747
R18535 gnd.n3929 gnd.n3928 9.69747
R18536 gnd.n3898 gnd.n3897 9.69747
R18537 gnd.n3866 gnd.n3865 9.69747
R18538 gnd.n3834 gnd.n3833 9.69747
R18539 gnd.n3802 gnd.n3801 9.69747
R18540 gnd.n3771 gnd.n3770 9.69747
R18541 gnd.n3999 gnd.n3998 9.45567
R18542 gnd.n3967 gnd.n3966 9.45567
R18543 gnd.n3935 gnd.n3934 9.45567
R18544 gnd.n3904 gnd.n3903 9.45567
R18545 gnd.n3872 gnd.n3871 9.45567
R18546 gnd.n3840 gnd.n3839 9.45567
R18547 gnd.n3808 gnd.n3807 9.45567
R18548 gnd.n3777 gnd.n3776 9.45567
R18549 gnd.n6007 gnd.n6006 9.30959
R18550 gnd.n7477 gnd.n279 9.30959
R18551 gnd.n4365 gnd.n4364 9.30959
R18552 gnd.n2338 gnd.n2302 9.30959
R18553 gnd.n3998 gnd.n3997 9.3005
R18554 gnd.n3971 gnd.n3970 9.3005
R18555 gnd.n3992 gnd.n3991 9.3005
R18556 gnd.n3990 gnd.n3989 9.3005
R18557 gnd.n3975 gnd.n3974 9.3005
R18558 gnd.n3984 gnd.n3983 9.3005
R18559 gnd.n3982 gnd.n3981 9.3005
R18560 gnd.n3966 gnd.n3965 9.3005
R18561 gnd.n3939 gnd.n3938 9.3005
R18562 gnd.n3960 gnd.n3959 9.3005
R18563 gnd.n3958 gnd.n3957 9.3005
R18564 gnd.n3943 gnd.n3942 9.3005
R18565 gnd.n3952 gnd.n3951 9.3005
R18566 gnd.n3950 gnd.n3949 9.3005
R18567 gnd.n3934 gnd.n3933 9.3005
R18568 gnd.n3907 gnd.n3906 9.3005
R18569 gnd.n3928 gnd.n3927 9.3005
R18570 gnd.n3926 gnd.n3925 9.3005
R18571 gnd.n3911 gnd.n3910 9.3005
R18572 gnd.n3920 gnd.n3919 9.3005
R18573 gnd.n3918 gnd.n3917 9.3005
R18574 gnd.n3903 gnd.n3902 9.3005
R18575 gnd.n3876 gnd.n3875 9.3005
R18576 gnd.n3897 gnd.n3896 9.3005
R18577 gnd.n3895 gnd.n3894 9.3005
R18578 gnd.n3880 gnd.n3879 9.3005
R18579 gnd.n3889 gnd.n3888 9.3005
R18580 gnd.n3887 gnd.n3886 9.3005
R18581 gnd.n3871 gnd.n3870 9.3005
R18582 gnd.n3844 gnd.n3843 9.3005
R18583 gnd.n3865 gnd.n3864 9.3005
R18584 gnd.n3863 gnd.n3862 9.3005
R18585 gnd.n3848 gnd.n3847 9.3005
R18586 gnd.n3857 gnd.n3856 9.3005
R18587 gnd.n3855 gnd.n3854 9.3005
R18588 gnd.n3839 gnd.n3838 9.3005
R18589 gnd.n3812 gnd.n3811 9.3005
R18590 gnd.n3833 gnd.n3832 9.3005
R18591 gnd.n3831 gnd.n3830 9.3005
R18592 gnd.n3816 gnd.n3815 9.3005
R18593 gnd.n3825 gnd.n3824 9.3005
R18594 gnd.n3823 gnd.n3822 9.3005
R18595 gnd.n3807 gnd.n3806 9.3005
R18596 gnd.n3780 gnd.n3779 9.3005
R18597 gnd.n3801 gnd.n3800 9.3005
R18598 gnd.n3799 gnd.n3798 9.3005
R18599 gnd.n3784 gnd.n3783 9.3005
R18600 gnd.n3793 gnd.n3792 9.3005
R18601 gnd.n3791 gnd.n3790 9.3005
R18602 gnd.n3776 gnd.n3775 9.3005
R18603 gnd.n3749 gnd.n3748 9.3005
R18604 gnd.n3770 gnd.n3769 9.3005
R18605 gnd.n3768 gnd.n3767 9.3005
R18606 gnd.n3753 gnd.n3752 9.3005
R18607 gnd.n3762 gnd.n3761 9.3005
R18608 gnd.n3760 gnd.n3759 9.3005
R18609 gnd.n4124 gnd.n4123 9.3005
R18610 gnd.n4122 gnd.n2675 9.3005
R18611 gnd.n4121 gnd.n4120 9.3005
R18612 gnd.n4117 gnd.n2676 9.3005
R18613 gnd.n4114 gnd.n2677 9.3005
R18614 gnd.n4113 gnd.n2678 9.3005
R18615 gnd.n4110 gnd.n2679 9.3005
R18616 gnd.n4109 gnd.n2680 9.3005
R18617 gnd.n4106 gnd.n2681 9.3005
R18618 gnd.n4105 gnd.n2682 9.3005
R18619 gnd.n4102 gnd.n2683 9.3005
R18620 gnd.n4101 gnd.n2684 9.3005
R18621 gnd.n4098 gnd.n2685 9.3005
R18622 gnd.n4097 gnd.n2686 9.3005
R18623 gnd.n4094 gnd.n4093 9.3005
R18624 gnd.n4092 gnd.n2687 9.3005
R18625 gnd.n4125 gnd.n2674 9.3005
R18626 gnd.n3365 gnd.n3364 9.3005
R18627 gnd.n3069 gnd.n3068 9.3005
R18628 gnd.n3392 gnd.n3391 9.3005
R18629 gnd.n3393 gnd.n3067 9.3005
R18630 gnd.n3397 gnd.n3394 9.3005
R18631 gnd.n3396 gnd.n3395 9.3005
R18632 gnd.n3041 gnd.n3040 9.3005
R18633 gnd.n3422 gnd.n3421 9.3005
R18634 gnd.n3423 gnd.n3039 9.3005
R18635 gnd.n3425 gnd.n3424 9.3005
R18636 gnd.n3019 gnd.n3018 9.3005
R18637 gnd.n3453 gnd.n3452 9.3005
R18638 gnd.n3454 gnd.n3017 9.3005
R18639 gnd.n3462 gnd.n3455 9.3005
R18640 gnd.n3461 gnd.n3456 9.3005
R18641 gnd.n3460 gnd.n3458 9.3005
R18642 gnd.n3457 gnd.n2966 9.3005
R18643 gnd.n3510 gnd.n2967 9.3005
R18644 gnd.n3509 gnd.n2968 9.3005
R18645 gnd.n3508 gnd.n2969 9.3005
R18646 gnd.n2988 gnd.n2970 9.3005
R18647 gnd.n2990 gnd.n2989 9.3005
R18648 gnd.n2872 gnd.n2871 9.3005
R18649 gnd.n3548 gnd.n3547 9.3005
R18650 gnd.n3549 gnd.n2870 9.3005
R18651 gnd.n3553 gnd.n3550 9.3005
R18652 gnd.n3552 gnd.n3551 9.3005
R18653 gnd.n2845 gnd.n2844 9.3005
R18654 gnd.n3588 gnd.n3587 9.3005
R18655 gnd.n3589 gnd.n2843 9.3005
R18656 gnd.n3593 gnd.n3590 9.3005
R18657 gnd.n3592 gnd.n3591 9.3005
R18658 gnd.n2818 gnd.n2817 9.3005
R18659 gnd.n3633 gnd.n3632 9.3005
R18660 gnd.n3634 gnd.n2816 9.3005
R18661 gnd.n3638 gnd.n3635 9.3005
R18662 gnd.n3637 gnd.n3636 9.3005
R18663 gnd.n2790 gnd.n2789 9.3005
R18664 gnd.n3673 gnd.n3672 9.3005
R18665 gnd.n3674 gnd.n2788 9.3005
R18666 gnd.n3678 gnd.n3675 9.3005
R18667 gnd.n3677 gnd.n3676 9.3005
R18668 gnd.n2763 gnd.n2762 9.3005
R18669 gnd.n3722 gnd.n3721 9.3005
R18670 gnd.n3723 gnd.n2761 9.3005
R18671 gnd.n3727 gnd.n3724 9.3005
R18672 gnd.n3726 gnd.n3725 9.3005
R18673 gnd.n2736 gnd.n2735 9.3005
R18674 gnd.n4017 gnd.n4016 9.3005
R18675 gnd.n4018 gnd.n2734 9.3005
R18676 gnd.n4024 gnd.n4019 9.3005
R18677 gnd.n4023 gnd.n4020 9.3005
R18678 gnd.n4022 gnd.n4021 9.3005
R18679 gnd.n3366 gnd.n3363 9.3005
R18680 gnd.n3148 gnd.n3107 9.3005
R18681 gnd.n3143 gnd.n3142 9.3005
R18682 gnd.n3141 gnd.n3108 9.3005
R18683 gnd.n3140 gnd.n3139 9.3005
R18684 gnd.n3136 gnd.n3109 9.3005
R18685 gnd.n3133 gnd.n3132 9.3005
R18686 gnd.n3131 gnd.n3110 9.3005
R18687 gnd.n3130 gnd.n3129 9.3005
R18688 gnd.n3126 gnd.n3111 9.3005
R18689 gnd.n3123 gnd.n3122 9.3005
R18690 gnd.n3121 gnd.n3112 9.3005
R18691 gnd.n3120 gnd.n3119 9.3005
R18692 gnd.n3116 gnd.n3114 9.3005
R18693 gnd.n3113 gnd.n3093 9.3005
R18694 gnd.n3360 gnd.n3092 9.3005
R18695 gnd.n3362 gnd.n3361 9.3005
R18696 gnd.n3150 gnd.n3149 9.3005
R18697 gnd.n3373 gnd.n3079 9.3005
R18698 gnd.n3380 gnd.n3080 9.3005
R18699 gnd.n3382 gnd.n3381 9.3005
R18700 gnd.n3383 gnd.n3060 9.3005
R18701 gnd.n3402 gnd.n3401 9.3005
R18702 gnd.n3404 gnd.n3052 9.3005
R18703 gnd.n3411 gnd.n3054 9.3005
R18704 gnd.n3412 gnd.n3049 9.3005
R18705 gnd.n3414 gnd.n3413 9.3005
R18706 gnd.n3050 gnd.n3035 9.3005
R18707 gnd.n3430 gnd.n3033 9.3005
R18708 gnd.n3434 gnd.n3433 9.3005
R18709 gnd.n3432 gnd.n3009 9.3005
R18710 gnd.n3469 gnd.n3008 9.3005
R18711 gnd.n3472 gnd.n3471 9.3005
R18712 gnd.n3005 gnd.n3004 9.3005
R18713 gnd.n3478 gnd.n3006 9.3005
R18714 gnd.n3480 gnd.n3479 9.3005
R18715 gnd.n3482 gnd.n3003 9.3005
R18716 gnd.n3485 gnd.n3484 9.3005
R18717 gnd.n3488 gnd.n3486 9.3005
R18718 gnd.n3490 gnd.n3489 9.3005
R18719 gnd.n3496 gnd.n3491 9.3005
R18720 gnd.n3495 gnd.n3494 9.3005
R18721 gnd.n2863 gnd.n2862 9.3005
R18722 gnd.n3562 gnd.n3561 9.3005
R18723 gnd.n3563 gnd.n2856 9.3005
R18724 gnd.n3571 gnd.n2855 9.3005
R18725 gnd.n3574 gnd.n3573 9.3005
R18726 gnd.n3576 gnd.n3575 9.3005
R18727 gnd.n3579 gnd.n2838 9.3005
R18728 gnd.n3577 gnd.n2836 9.3005
R18729 gnd.n3599 gnd.n2834 9.3005
R18730 gnd.n3601 gnd.n3600 9.3005
R18731 gnd.n2808 gnd.n2807 9.3005
R18732 gnd.n3647 gnd.n3646 9.3005
R18733 gnd.n3648 gnd.n2801 9.3005
R18734 gnd.n3656 gnd.n2800 9.3005
R18735 gnd.n3659 gnd.n3658 9.3005
R18736 gnd.n3661 gnd.n3660 9.3005
R18737 gnd.n3664 gnd.n2783 9.3005
R18738 gnd.n3662 gnd.n2781 9.3005
R18739 gnd.n3684 gnd.n2779 9.3005
R18740 gnd.n3686 gnd.n3685 9.3005
R18741 gnd.n2754 gnd.n2753 9.3005
R18742 gnd.n3736 gnd.n3735 9.3005
R18743 gnd.n3737 gnd.n2747 9.3005
R18744 gnd.n3746 gnd.n2746 9.3005
R18745 gnd.n4005 gnd.n4004 9.3005
R18746 gnd.n4007 gnd.n4006 9.3005
R18747 gnd.n4008 gnd.n2727 9.3005
R18748 gnd.n4032 gnd.n4031 9.3005
R18749 gnd.n2728 gnd.n2690 9.3005
R18750 gnd.n3371 gnd.n3370 9.3005
R18751 gnd.n4088 gnd.n2691 9.3005
R18752 gnd.n4087 gnd.n2693 9.3005
R18753 gnd.n4084 gnd.n2694 9.3005
R18754 gnd.n4083 gnd.n2695 9.3005
R18755 gnd.n4080 gnd.n2696 9.3005
R18756 gnd.n4079 gnd.n2697 9.3005
R18757 gnd.n4076 gnd.n2698 9.3005
R18758 gnd.n4075 gnd.n2699 9.3005
R18759 gnd.n4072 gnd.n2700 9.3005
R18760 gnd.n4071 gnd.n2701 9.3005
R18761 gnd.n4068 gnd.n2702 9.3005
R18762 gnd.n4067 gnd.n2703 9.3005
R18763 gnd.n4064 gnd.n2704 9.3005
R18764 gnd.n4063 gnd.n2705 9.3005
R18765 gnd.n4060 gnd.n2706 9.3005
R18766 gnd.n4059 gnd.n2707 9.3005
R18767 gnd.n4056 gnd.n2708 9.3005
R18768 gnd.n4055 gnd.n2709 9.3005
R18769 gnd.n4052 gnd.n2710 9.3005
R18770 gnd.n4051 gnd.n2711 9.3005
R18771 gnd.n4048 gnd.n2712 9.3005
R18772 gnd.n4047 gnd.n2713 9.3005
R18773 gnd.n4044 gnd.n2717 9.3005
R18774 gnd.n4043 gnd.n2718 9.3005
R18775 gnd.n4040 gnd.n2719 9.3005
R18776 gnd.n4039 gnd.n2720 9.3005
R18777 gnd.n4090 gnd.n4089 9.3005
R18778 gnd.n3540 gnd.n3524 9.3005
R18779 gnd.n3539 gnd.n3525 9.3005
R18780 gnd.n3538 gnd.n3526 9.3005
R18781 gnd.n3536 gnd.n3527 9.3005
R18782 gnd.n3535 gnd.n3528 9.3005
R18783 gnd.n3533 gnd.n3529 9.3005
R18784 gnd.n3532 gnd.n3530 9.3005
R18785 gnd.n2826 gnd.n2825 9.3005
R18786 gnd.n3609 gnd.n3608 9.3005
R18787 gnd.n3610 gnd.n2824 9.3005
R18788 gnd.n3627 gnd.n3611 9.3005
R18789 gnd.n3626 gnd.n3612 9.3005
R18790 gnd.n3625 gnd.n3613 9.3005
R18791 gnd.n3623 gnd.n3614 9.3005
R18792 gnd.n3622 gnd.n3615 9.3005
R18793 gnd.n3620 gnd.n3616 9.3005
R18794 gnd.n3619 gnd.n3617 9.3005
R18795 gnd.n2770 gnd.n2769 9.3005
R18796 gnd.n3694 gnd.n3693 9.3005
R18797 gnd.n3695 gnd.n2768 9.3005
R18798 gnd.n3716 gnd.n3696 9.3005
R18799 gnd.n3715 gnd.n3697 9.3005
R18800 gnd.n3714 gnd.n3698 9.3005
R18801 gnd.n3711 gnd.n3699 9.3005
R18802 gnd.n3710 gnd.n3700 9.3005
R18803 gnd.n3708 gnd.n3701 9.3005
R18804 gnd.n3707 gnd.n3702 9.3005
R18805 gnd.n3705 gnd.n3704 9.3005
R18806 gnd.n3703 gnd.n2722 9.3005
R18807 gnd.n3281 gnd.n3280 9.3005
R18808 gnd.n3171 gnd.n3170 9.3005
R18809 gnd.n3295 gnd.n3294 9.3005
R18810 gnd.n3296 gnd.n3169 9.3005
R18811 gnd.n3298 gnd.n3297 9.3005
R18812 gnd.n3159 gnd.n3158 9.3005
R18813 gnd.n3311 gnd.n3310 9.3005
R18814 gnd.n3312 gnd.n3157 9.3005
R18815 gnd.n3344 gnd.n3313 9.3005
R18816 gnd.n3343 gnd.n3314 9.3005
R18817 gnd.n3342 gnd.n3315 9.3005
R18818 gnd.n3341 gnd.n3316 9.3005
R18819 gnd.n3338 gnd.n3317 9.3005
R18820 gnd.n3337 gnd.n3318 9.3005
R18821 gnd.n3336 gnd.n3319 9.3005
R18822 gnd.n3334 gnd.n3320 9.3005
R18823 gnd.n3333 gnd.n3321 9.3005
R18824 gnd.n3330 gnd.n3322 9.3005
R18825 gnd.n3329 gnd.n3323 9.3005
R18826 gnd.n3328 gnd.n3324 9.3005
R18827 gnd.n3326 gnd.n3325 9.3005
R18828 gnd.n3025 gnd.n3024 9.3005
R18829 gnd.n3442 gnd.n3441 9.3005
R18830 gnd.n3443 gnd.n3023 9.3005
R18831 gnd.n3447 gnd.n3444 9.3005
R18832 gnd.n3446 gnd.n3445 9.3005
R18833 gnd.n2947 gnd.n2946 9.3005
R18834 gnd.n3522 gnd.n3521 9.3005
R18835 gnd.n3279 gnd.n3180 9.3005
R18836 gnd.n3182 gnd.n3181 9.3005
R18837 gnd.n3226 gnd.n3224 9.3005
R18838 gnd.n3227 gnd.n3223 9.3005
R18839 gnd.n3230 gnd.n3219 9.3005
R18840 gnd.n3231 gnd.n3218 9.3005
R18841 gnd.n3234 gnd.n3217 9.3005
R18842 gnd.n3235 gnd.n3216 9.3005
R18843 gnd.n3238 gnd.n3215 9.3005
R18844 gnd.n3239 gnd.n3214 9.3005
R18845 gnd.n3242 gnd.n3213 9.3005
R18846 gnd.n3243 gnd.n3212 9.3005
R18847 gnd.n3246 gnd.n3211 9.3005
R18848 gnd.n3247 gnd.n3210 9.3005
R18849 gnd.n3250 gnd.n3209 9.3005
R18850 gnd.n3251 gnd.n3208 9.3005
R18851 gnd.n3254 gnd.n3207 9.3005
R18852 gnd.n3255 gnd.n3206 9.3005
R18853 gnd.n3258 gnd.n3205 9.3005
R18854 gnd.n3259 gnd.n3204 9.3005
R18855 gnd.n3262 gnd.n3203 9.3005
R18856 gnd.n3263 gnd.n3202 9.3005
R18857 gnd.n3266 gnd.n3201 9.3005
R18858 gnd.n3268 gnd.n3200 9.3005
R18859 gnd.n3269 gnd.n3199 9.3005
R18860 gnd.n3270 gnd.n3198 9.3005
R18861 gnd.n3271 gnd.n3197 9.3005
R18862 gnd.n3278 gnd.n3277 9.3005
R18863 gnd.n3287 gnd.n3286 9.3005
R18864 gnd.n3288 gnd.n3174 9.3005
R18865 gnd.n3290 gnd.n3289 9.3005
R18866 gnd.n3165 gnd.n3164 9.3005
R18867 gnd.n3303 gnd.n3302 9.3005
R18868 gnd.n3304 gnd.n3163 9.3005
R18869 gnd.n3306 gnd.n3305 9.3005
R18870 gnd.n3152 gnd.n3151 9.3005
R18871 gnd.n3349 gnd.n3348 9.3005
R18872 gnd.n3350 gnd.n3106 9.3005
R18873 gnd.n3354 gnd.n3352 9.3005
R18874 gnd.n3353 gnd.n3085 9.3005
R18875 gnd.n3372 gnd.n3084 9.3005
R18876 gnd.n3375 gnd.n3374 9.3005
R18877 gnd.n3078 gnd.n3077 9.3005
R18878 gnd.n3386 gnd.n3384 9.3005
R18879 gnd.n3385 gnd.n3059 9.3005
R18880 gnd.n3403 gnd.n3058 9.3005
R18881 gnd.n3406 gnd.n3405 9.3005
R18882 gnd.n3053 gnd.n3048 9.3005
R18883 gnd.n3416 gnd.n3415 9.3005
R18884 gnd.n3051 gnd.n3031 9.3005
R18885 gnd.n3437 gnd.n3032 9.3005
R18886 gnd.n3436 gnd.n3435 9.3005
R18887 gnd.n3034 gnd.n3010 9.3005
R18888 gnd.n3468 gnd.n3467 9.3005
R18889 gnd.n3470 gnd.n2955 9.3005
R18890 gnd.n3517 gnd.n2956 9.3005
R18891 gnd.n3516 gnd.n2957 9.3005
R18892 gnd.n3515 gnd.n2958 9.3005
R18893 gnd.n3481 gnd.n2959 9.3005
R18894 gnd.n3483 gnd.n2977 9.3005
R18895 gnd.n3503 gnd.n2978 9.3005
R18896 gnd.n3502 gnd.n2979 9.3005
R18897 gnd.n3501 gnd.n2980 9.3005
R18898 gnd.n3492 gnd.n2981 9.3005
R18899 gnd.n3493 gnd.n2864 9.3005
R18900 gnd.n3559 gnd.n3558 9.3005
R18901 gnd.n3560 gnd.n2857 9.3005
R18902 gnd.n3570 gnd.n3569 9.3005
R18903 gnd.n3572 gnd.n2853 9.3005
R18904 gnd.n3582 gnd.n2854 9.3005
R18905 gnd.n3581 gnd.n3580 9.3005
R18906 gnd.n3578 gnd.n2832 9.3005
R18907 gnd.n3604 gnd.n2833 9.3005
R18908 gnd.n3603 gnd.n3602 9.3005
R18909 gnd.n2835 gnd.n2809 9.3005
R18910 gnd.n3644 gnd.n3643 9.3005
R18911 gnd.n3645 gnd.n2802 9.3005
R18912 gnd.n3655 gnd.n3654 9.3005
R18913 gnd.n3657 gnd.n2798 9.3005
R18914 gnd.n3667 gnd.n2799 9.3005
R18915 gnd.n3666 gnd.n3665 9.3005
R18916 gnd.n3663 gnd.n2777 9.3005
R18917 gnd.n3689 gnd.n2778 9.3005
R18918 gnd.n3688 gnd.n3687 9.3005
R18919 gnd.n2780 gnd.n2755 9.3005
R18920 gnd.n3733 gnd.n3732 9.3005
R18921 gnd.n3734 gnd.n2748 9.3005
R18922 gnd.n3745 gnd.n3744 9.3005
R18923 gnd.n4003 gnd.n2744 9.3005
R18924 gnd.n4011 gnd.n2745 9.3005
R18925 gnd.n4010 gnd.n4009 9.3005
R18926 gnd.n2726 gnd.n2725 9.3005
R18927 gnd.n4034 gnd.n4033 9.3005
R18928 gnd.n3176 gnd.n3175 9.3005
R18929 gnd.n6656 gnd.n768 9.3005
R18930 gnd.n6658 gnd.n6657 9.3005
R18931 gnd.n764 gnd.n763 9.3005
R18932 gnd.n6665 gnd.n6664 9.3005
R18933 gnd.n6666 gnd.n762 9.3005
R18934 gnd.n6668 gnd.n6667 9.3005
R18935 gnd.n758 gnd.n757 9.3005
R18936 gnd.n6675 gnd.n6674 9.3005
R18937 gnd.n6676 gnd.n756 9.3005
R18938 gnd.n6678 gnd.n6677 9.3005
R18939 gnd.n752 gnd.n751 9.3005
R18940 gnd.n6685 gnd.n6684 9.3005
R18941 gnd.n6686 gnd.n750 9.3005
R18942 gnd.n6688 gnd.n6687 9.3005
R18943 gnd.n746 gnd.n745 9.3005
R18944 gnd.n6695 gnd.n6694 9.3005
R18945 gnd.n6696 gnd.n744 9.3005
R18946 gnd.n6698 gnd.n6697 9.3005
R18947 gnd.n740 gnd.n739 9.3005
R18948 gnd.n6705 gnd.n6704 9.3005
R18949 gnd.n6706 gnd.n738 9.3005
R18950 gnd.n6708 gnd.n6707 9.3005
R18951 gnd.n734 gnd.n733 9.3005
R18952 gnd.n6715 gnd.n6714 9.3005
R18953 gnd.n6716 gnd.n732 9.3005
R18954 gnd.n6718 gnd.n6717 9.3005
R18955 gnd.n728 gnd.n727 9.3005
R18956 gnd.n6725 gnd.n6724 9.3005
R18957 gnd.n6726 gnd.n726 9.3005
R18958 gnd.n6728 gnd.n6727 9.3005
R18959 gnd.n722 gnd.n721 9.3005
R18960 gnd.n6735 gnd.n6734 9.3005
R18961 gnd.n6736 gnd.n720 9.3005
R18962 gnd.n6738 gnd.n6737 9.3005
R18963 gnd.n716 gnd.n715 9.3005
R18964 gnd.n6745 gnd.n6744 9.3005
R18965 gnd.n6746 gnd.n714 9.3005
R18966 gnd.n6748 gnd.n6747 9.3005
R18967 gnd.n710 gnd.n709 9.3005
R18968 gnd.n6755 gnd.n6754 9.3005
R18969 gnd.n6756 gnd.n708 9.3005
R18970 gnd.n6758 gnd.n6757 9.3005
R18971 gnd.n704 gnd.n703 9.3005
R18972 gnd.n6765 gnd.n6764 9.3005
R18973 gnd.n6766 gnd.n702 9.3005
R18974 gnd.n6768 gnd.n6767 9.3005
R18975 gnd.n698 gnd.n697 9.3005
R18976 gnd.n6775 gnd.n6774 9.3005
R18977 gnd.n6776 gnd.n696 9.3005
R18978 gnd.n6778 gnd.n6777 9.3005
R18979 gnd.n692 gnd.n691 9.3005
R18980 gnd.n6785 gnd.n6784 9.3005
R18981 gnd.n6786 gnd.n690 9.3005
R18982 gnd.n6788 gnd.n6787 9.3005
R18983 gnd.n686 gnd.n685 9.3005
R18984 gnd.n6795 gnd.n6794 9.3005
R18985 gnd.n6796 gnd.n684 9.3005
R18986 gnd.n6798 gnd.n6797 9.3005
R18987 gnd.n680 gnd.n679 9.3005
R18988 gnd.n6805 gnd.n6804 9.3005
R18989 gnd.n6806 gnd.n678 9.3005
R18990 gnd.n6808 gnd.n6807 9.3005
R18991 gnd.n674 gnd.n673 9.3005
R18992 gnd.n6815 gnd.n6814 9.3005
R18993 gnd.n6816 gnd.n672 9.3005
R18994 gnd.n6818 gnd.n6817 9.3005
R18995 gnd.n668 gnd.n667 9.3005
R18996 gnd.n6825 gnd.n6824 9.3005
R18997 gnd.n6826 gnd.n666 9.3005
R18998 gnd.n6828 gnd.n6827 9.3005
R18999 gnd.n662 gnd.n661 9.3005
R19000 gnd.n6835 gnd.n6834 9.3005
R19001 gnd.n6836 gnd.n660 9.3005
R19002 gnd.n6838 gnd.n6837 9.3005
R19003 gnd.n656 gnd.n655 9.3005
R19004 gnd.n6845 gnd.n6844 9.3005
R19005 gnd.n6846 gnd.n654 9.3005
R19006 gnd.n6848 gnd.n6847 9.3005
R19007 gnd.n650 gnd.n649 9.3005
R19008 gnd.n6855 gnd.n6854 9.3005
R19009 gnd.n6856 gnd.n648 9.3005
R19010 gnd.n6858 gnd.n6857 9.3005
R19011 gnd.n644 gnd.n643 9.3005
R19012 gnd.n6865 gnd.n6864 9.3005
R19013 gnd.n6866 gnd.n642 9.3005
R19014 gnd.n6868 gnd.n6867 9.3005
R19015 gnd.n638 gnd.n637 9.3005
R19016 gnd.n6875 gnd.n6874 9.3005
R19017 gnd.n6876 gnd.n636 9.3005
R19018 gnd.n6878 gnd.n6877 9.3005
R19019 gnd.n632 gnd.n631 9.3005
R19020 gnd.n6885 gnd.n6884 9.3005
R19021 gnd.n6886 gnd.n630 9.3005
R19022 gnd.n6888 gnd.n6887 9.3005
R19023 gnd.n626 gnd.n625 9.3005
R19024 gnd.n6895 gnd.n6894 9.3005
R19025 gnd.n6896 gnd.n624 9.3005
R19026 gnd.n6898 gnd.n6897 9.3005
R19027 gnd.n620 gnd.n619 9.3005
R19028 gnd.n6905 gnd.n6904 9.3005
R19029 gnd.n6906 gnd.n618 9.3005
R19030 gnd.n6908 gnd.n6907 9.3005
R19031 gnd.n614 gnd.n613 9.3005
R19032 gnd.n6915 gnd.n6914 9.3005
R19033 gnd.n6916 gnd.n612 9.3005
R19034 gnd.n6918 gnd.n6917 9.3005
R19035 gnd.n608 gnd.n607 9.3005
R19036 gnd.n6925 gnd.n6924 9.3005
R19037 gnd.n6926 gnd.n606 9.3005
R19038 gnd.n6928 gnd.n6927 9.3005
R19039 gnd.n602 gnd.n601 9.3005
R19040 gnd.n6935 gnd.n6934 9.3005
R19041 gnd.n6936 gnd.n600 9.3005
R19042 gnd.n6938 gnd.n6937 9.3005
R19043 gnd.n596 gnd.n595 9.3005
R19044 gnd.n6945 gnd.n6944 9.3005
R19045 gnd.n6946 gnd.n594 9.3005
R19046 gnd.n6948 gnd.n6947 9.3005
R19047 gnd.n590 gnd.n589 9.3005
R19048 gnd.n6955 gnd.n6954 9.3005
R19049 gnd.n6956 gnd.n588 9.3005
R19050 gnd.n6958 gnd.n6957 9.3005
R19051 gnd.n584 gnd.n583 9.3005
R19052 gnd.n6965 gnd.n6964 9.3005
R19053 gnd.n6966 gnd.n582 9.3005
R19054 gnd.n6968 gnd.n6967 9.3005
R19055 gnd.n578 gnd.n577 9.3005
R19056 gnd.n6975 gnd.n6974 9.3005
R19057 gnd.n6976 gnd.n576 9.3005
R19058 gnd.n6978 gnd.n6977 9.3005
R19059 gnd.n572 gnd.n571 9.3005
R19060 gnd.n6985 gnd.n6984 9.3005
R19061 gnd.n6986 gnd.n570 9.3005
R19062 gnd.n6988 gnd.n6987 9.3005
R19063 gnd.n566 gnd.n565 9.3005
R19064 gnd.n6995 gnd.n6994 9.3005
R19065 gnd.n6996 gnd.n564 9.3005
R19066 gnd.n6998 gnd.n6997 9.3005
R19067 gnd.n560 gnd.n559 9.3005
R19068 gnd.n7005 gnd.n7004 9.3005
R19069 gnd.n7006 gnd.n558 9.3005
R19070 gnd.n7008 gnd.n7007 9.3005
R19071 gnd.n554 gnd.n553 9.3005
R19072 gnd.n7015 gnd.n7014 9.3005
R19073 gnd.n7016 gnd.n552 9.3005
R19074 gnd.n7018 gnd.n7017 9.3005
R19075 gnd.n548 gnd.n547 9.3005
R19076 gnd.n7025 gnd.n7024 9.3005
R19077 gnd.n7026 gnd.n546 9.3005
R19078 gnd.n7028 gnd.n7027 9.3005
R19079 gnd.n542 gnd.n541 9.3005
R19080 gnd.n7035 gnd.n7034 9.3005
R19081 gnd.n7036 gnd.n540 9.3005
R19082 gnd.n7038 gnd.n7037 9.3005
R19083 gnd.n536 gnd.n535 9.3005
R19084 gnd.n7045 gnd.n7044 9.3005
R19085 gnd.n7046 gnd.n534 9.3005
R19086 gnd.n7048 gnd.n7047 9.3005
R19087 gnd.n530 gnd.n529 9.3005
R19088 gnd.n7055 gnd.n7054 9.3005
R19089 gnd.n7056 gnd.n528 9.3005
R19090 gnd.n7058 gnd.n7057 9.3005
R19091 gnd.n524 gnd.n523 9.3005
R19092 gnd.n7065 gnd.n7064 9.3005
R19093 gnd.n7066 gnd.n522 9.3005
R19094 gnd.n7068 gnd.n7067 9.3005
R19095 gnd.n518 gnd.n517 9.3005
R19096 gnd.n7075 gnd.n7074 9.3005
R19097 gnd.n7078 gnd.n7077 9.3005
R19098 gnd.n512 gnd.n511 9.3005
R19099 gnd.n7085 gnd.n7084 9.3005
R19100 gnd.n7086 gnd.n510 9.3005
R19101 gnd.n7088 gnd.n7087 9.3005
R19102 gnd.n506 gnd.n505 9.3005
R19103 gnd.n7095 gnd.n7094 9.3005
R19104 gnd.n7096 gnd.n504 9.3005
R19105 gnd.n7098 gnd.n7097 9.3005
R19106 gnd.n500 gnd.n499 9.3005
R19107 gnd.n7105 gnd.n7104 9.3005
R19108 gnd.n7106 gnd.n498 9.3005
R19109 gnd.n7108 gnd.n7107 9.3005
R19110 gnd.n494 gnd.n493 9.3005
R19111 gnd.n7115 gnd.n7114 9.3005
R19112 gnd.n7116 gnd.n492 9.3005
R19113 gnd.n7118 gnd.n7117 9.3005
R19114 gnd.n488 gnd.n487 9.3005
R19115 gnd.n7125 gnd.n7124 9.3005
R19116 gnd.n7126 gnd.n486 9.3005
R19117 gnd.n7128 gnd.n7127 9.3005
R19118 gnd.n482 gnd.n481 9.3005
R19119 gnd.n7135 gnd.n7134 9.3005
R19120 gnd.n7136 gnd.n480 9.3005
R19121 gnd.n7138 gnd.n7137 9.3005
R19122 gnd.n476 gnd.n475 9.3005
R19123 gnd.n7145 gnd.n7144 9.3005
R19124 gnd.n7146 gnd.n474 9.3005
R19125 gnd.n7148 gnd.n7147 9.3005
R19126 gnd.n470 gnd.n469 9.3005
R19127 gnd.n7155 gnd.n7154 9.3005
R19128 gnd.n7156 gnd.n468 9.3005
R19129 gnd.n7158 gnd.n7157 9.3005
R19130 gnd.n464 gnd.n463 9.3005
R19131 gnd.n7165 gnd.n7164 9.3005
R19132 gnd.n7166 gnd.n462 9.3005
R19133 gnd.n7168 gnd.n7167 9.3005
R19134 gnd.n458 gnd.n457 9.3005
R19135 gnd.n7175 gnd.n7174 9.3005
R19136 gnd.n7176 gnd.n456 9.3005
R19137 gnd.n7178 gnd.n7177 9.3005
R19138 gnd.n452 gnd.n451 9.3005
R19139 gnd.n7185 gnd.n7184 9.3005
R19140 gnd.n7186 gnd.n450 9.3005
R19141 gnd.n7188 gnd.n7187 9.3005
R19142 gnd.n446 gnd.n445 9.3005
R19143 gnd.n7195 gnd.n7194 9.3005
R19144 gnd.n7196 gnd.n444 9.3005
R19145 gnd.n7198 gnd.n7197 9.3005
R19146 gnd.n440 gnd.n439 9.3005
R19147 gnd.n7205 gnd.n7204 9.3005
R19148 gnd.n7206 gnd.n438 9.3005
R19149 gnd.n7208 gnd.n7207 9.3005
R19150 gnd.n434 gnd.n433 9.3005
R19151 gnd.n7215 gnd.n7214 9.3005
R19152 gnd.n7216 gnd.n432 9.3005
R19153 gnd.n7218 gnd.n7217 9.3005
R19154 gnd.n428 gnd.n427 9.3005
R19155 gnd.n7225 gnd.n7224 9.3005
R19156 gnd.n7226 gnd.n426 9.3005
R19157 gnd.n7228 gnd.n7227 9.3005
R19158 gnd.n422 gnd.n421 9.3005
R19159 gnd.n7235 gnd.n7234 9.3005
R19160 gnd.n7236 gnd.n420 9.3005
R19161 gnd.n7238 gnd.n7237 9.3005
R19162 gnd.n416 gnd.n415 9.3005
R19163 gnd.n7245 gnd.n7244 9.3005
R19164 gnd.n7246 gnd.n414 9.3005
R19165 gnd.n7248 gnd.n7247 9.3005
R19166 gnd.n410 gnd.n409 9.3005
R19167 gnd.n7255 gnd.n7254 9.3005
R19168 gnd.n7256 gnd.n408 9.3005
R19169 gnd.n7258 gnd.n7257 9.3005
R19170 gnd.n404 gnd.n403 9.3005
R19171 gnd.n7265 gnd.n7264 9.3005
R19172 gnd.n7266 gnd.n402 9.3005
R19173 gnd.n7268 gnd.n7267 9.3005
R19174 gnd.n398 gnd.n397 9.3005
R19175 gnd.n7275 gnd.n7274 9.3005
R19176 gnd.n7276 gnd.n396 9.3005
R19177 gnd.n7280 gnd.n7277 9.3005
R19178 gnd.n7279 gnd.n7278 9.3005
R19179 gnd.n392 gnd.n391 9.3005
R19180 gnd.n7288 gnd.n7287 9.3005
R19181 gnd.n7076 gnd.n516 9.3005
R19182 gnd.n7627 gnd.n7626 9.3005
R19183 gnd.n7625 gnd.n84 9.3005
R19184 gnd.n7360 gnd.n87 9.3005
R19185 gnd.n7361 gnd.n7359 9.3005
R19186 gnd.n7363 gnd.n7362 9.3005
R19187 gnd.n7365 gnd.n367 9.3005
R19188 gnd.n7367 gnd.n7366 9.3005
R19189 gnd.n7368 gnd.n366 9.3005
R19190 gnd.n7370 gnd.n7369 9.3005
R19191 gnd.n7372 gnd.n364 9.3005
R19192 gnd.n7374 gnd.n7373 9.3005
R19193 gnd.n7375 gnd.n363 9.3005
R19194 gnd.n7377 gnd.n7376 9.3005
R19195 gnd.n7379 gnd.n361 9.3005
R19196 gnd.n7381 gnd.n7380 9.3005
R19197 gnd.n7382 gnd.n360 9.3005
R19198 gnd.n7384 gnd.n7383 9.3005
R19199 gnd.n7386 gnd.n358 9.3005
R19200 gnd.n7388 gnd.n7387 9.3005
R19201 gnd.n7389 gnd.n357 9.3005
R19202 gnd.n7391 gnd.n7390 9.3005
R19203 gnd.n7393 gnd.n355 9.3005
R19204 gnd.n7395 gnd.n7394 9.3005
R19205 gnd.n7396 gnd.n354 9.3005
R19206 gnd.n7398 gnd.n7397 9.3005
R19207 gnd.n7400 gnd.n352 9.3005
R19208 gnd.n7402 gnd.n7401 9.3005
R19209 gnd.n7433 gnd.n318 9.3005
R19210 gnd.n7432 gnd.n320 9.3005
R19211 gnd.n324 gnd.n321 9.3005
R19212 gnd.n7427 gnd.n325 9.3005
R19213 gnd.n7426 gnd.n326 9.3005
R19214 gnd.n7425 gnd.n327 9.3005
R19215 gnd.n331 gnd.n328 9.3005
R19216 gnd.n7420 gnd.n332 9.3005
R19217 gnd.n7419 gnd.n333 9.3005
R19218 gnd.n7418 gnd.n334 9.3005
R19219 gnd.n338 gnd.n335 9.3005
R19220 gnd.n7413 gnd.n339 9.3005
R19221 gnd.n7412 gnd.n340 9.3005
R19222 gnd.n7411 gnd.n341 9.3005
R19223 gnd.n345 gnd.n342 9.3005
R19224 gnd.n7406 gnd.n346 9.3005
R19225 gnd.n7405 gnd.n7404 9.3005
R19226 gnd.n7403 gnd.n349 9.3005
R19227 gnd.n7435 gnd.n7434 9.3005
R19228 gnd.n7543 gnd.n215 9.3005
R19229 gnd.n7542 gnd.n217 9.3005
R19230 gnd.n221 gnd.n218 9.3005
R19231 gnd.n7537 gnd.n222 9.3005
R19232 gnd.n7536 gnd.n223 9.3005
R19233 gnd.n7535 gnd.n224 9.3005
R19234 gnd.n228 gnd.n225 9.3005
R19235 gnd.n7530 gnd.n229 9.3005
R19236 gnd.n7529 gnd.n230 9.3005
R19237 gnd.n7528 gnd.n231 9.3005
R19238 gnd.n235 gnd.n232 9.3005
R19239 gnd.n7523 gnd.n236 9.3005
R19240 gnd.n7522 gnd.n237 9.3005
R19241 gnd.n7521 gnd.n238 9.3005
R19242 gnd.n242 gnd.n239 9.3005
R19243 gnd.n7516 gnd.n243 9.3005
R19244 gnd.n7515 gnd.n244 9.3005
R19245 gnd.n7511 gnd.n245 9.3005
R19246 gnd.n249 gnd.n246 9.3005
R19247 gnd.n7506 gnd.n250 9.3005
R19248 gnd.n7505 gnd.n251 9.3005
R19249 gnd.n7504 gnd.n252 9.3005
R19250 gnd.n256 gnd.n253 9.3005
R19251 gnd.n7499 gnd.n257 9.3005
R19252 gnd.n7498 gnd.n258 9.3005
R19253 gnd.n7497 gnd.n259 9.3005
R19254 gnd.n263 gnd.n260 9.3005
R19255 gnd.n7492 gnd.n264 9.3005
R19256 gnd.n7491 gnd.n265 9.3005
R19257 gnd.n7490 gnd.n266 9.3005
R19258 gnd.n270 gnd.n267 9.3005
R19259 gnd.n7485 gnd.n271 9.3005
R19260 gnd.n7484 gnd.n272 9.3005
R19261 gnd.n7483 gnd.n273 9.3005
R19262 gnd.n277 gnd.n274 9.3005
R19263 gnd.n7478 gnd.n278 9.3005
R19264 gnd.n7477 gnd.n7476 9.3005
R19265 gnd.n7475 gnd.n279 9.3005
R19266 gnd.n7474 gnd.n7473 9.3005
R19267 gnd.n283 gnd.n282 9.3005
R19268 gnd.n288 gnd.n286 9.3005
R19269 gnd.n7466 gnd.n289 9.3005
R19270 gnd.n7465 gnd.n290 9.3005
R19271 gnd.n7464 gnd.n291 9.3005
R19272 gnd.n295 gnd.n292 9.3005
R19273 gnd.n7459 gnd.n296 9.3005
R19274 gnd.n7458 gnd.n297 9.3005
R19275 gnd.n7457 gnd.n298 9.3005
R19276 gnd.n302 gnd.n299 9.3005
R19277 gnd.n7452 gnd.n303 9.3005
R19278 gnd.n7451 gnd.n304 9.3005
R19279 gnd.n7450 gnd.n305 9.3005
R19280 gnd.n309 gnd.n306 9.3005
R19281 gnd.n7445 gnd.n310 9.3005
R19282 gnd.n7444 gnd.n311 9.3005
R19283 gnd.n7443 gnd.n312 9.3005
R19284 gnd.n317 gnd.n315 9.3005
R19285 gnd.n7438 gnd.n7437 9.3005
R19286 gnd.n7545 gnd.n7544 9.3005
R19287 gnd.n5956 gnd.n5955 9.3005
R19288 gnd.n1582 gnd.n1581 9.3005
R19289 gnd.n1606 gnd.n1605 9.3005
R19290 gnd.n5943 gnd.n1607 9.3005
R19291 gnd.n5942 gnd.n1608 9.3005
R19292 gnd.n5941 gnd.n1609 9.3005
R19293 gnd.n5747 gnd.n1610 9.3005
R19294 gnd.n5931 gnd.n1627 9.3005
R19295 gnd.n5930 gnd.n1628 9.3005
R19296 gnd.n5929 gnd.n1629 9.3005
R19297 gnd.n5753 gnd.n1630 9.3005
R19298 gnd.n5919 gnd.n1647 9.3005
R19299 gnd.n5918 gnd.n1648 9.3005
R19300 gnd.n5917 gnd.n1649 9.3005
R19301 gnd.n5833 gnd.n1650 9.3005
R19302 gnd.n5907 gnd.n1667 9.3005
R19303 gnd.n5906 gnd.n1668 9.3005
R19304 gnd.n5905 gnd.n1669 9.3005
R19305 gnd.n5848 gnd.n1670 9.3005
R19306 gnd.n5895 gnd.n1687 9.3005
R19307 gnd.n5894 gnd.n1688 9.3005
R19308 gnd.n5893 gnd.n1689 9.3005
R19309 gnd.n5851 gnd.n1690 9.3005
R19310 gnd.n379 gnd.n378 9.3005
R19311 gnd.n7302 gnd.n7301 9.3005
R19312 gnd.n7303 gnd.n372 9.3005
R19313 gnd.n7310 gnd.n373 9.3005
R19314 gnd.n7311 gnd.n371 9.3005
R19315 gnd.n7314 gnd.n7313 9.3005
R19316 gnd.n7315 gnd.n110 9.3005
R19317 gnd.n7613 gnd.n111 9.3005
R19318 gnd.n7612 gnd.n112 9.3005
R19319 gnd.n7611 gnd.n113 9.3005
R19320 gnd.n7316 gnd.n114 9.3005
R19321 gnd.n7601 gnd.n128 9.3005
R19322 gnd.n7600 gnd.n129 9.3005
R19323 gnd.n7599 gnd.n130 9.3005
R19324 gnd.n7317 gnd.n131 9.3005
R19325 gnd.n7589 gnd.n148 9.3005
R19326 gnd.n7588 gnd.n149 9.3005
R19327 gnd.n7587 gnd.n150 9.3005
R19328 gnd.n7318 gnd.n151 9.3005
R19329 gnd.n7577 gnd.n166 9.3005
R19330 gnd.n7576 gnd.n167 9.3005
R19331 gnd.n7575 gnd.n168 9.3005
R19332 gnd.n7319 gnd.n169 9.3005
R19333 gnd.n7565 gnd.n186 9.3005
R19334 gnd.n7564 gnd.n187 9.3005
R19335 gnd.n7563 gnd.n188 9.3005
R19336 gnd.n7320 gnd.n189 9.3005
R19337 gnd.n7553 gnd.n205 9.3005
R19338 gnd.n7552 gnd.n206 9.3005
R19339 gnd.n7551 gnd.n207 9.3005
R19340 gnd.n5957 gnd.n1580 9.3005
R19341 gnd.n5955 gnd.n5954 9.3005
R19342 gnd.n5953 gnd.n1582 9.3005
R19343 gnd.n1606 gnd.n1583 9.3005
R19344 gnd.n5742 gnd.n1607 9.3005
R19345 gnd.n5745 gnd.n1608 9.3005
R19346 gnd.n5746 gnd.n1609 9.3005
R19347 gnd.n5751 gnd.n5747 9.3005
R19348 gnd.n5752 gnd.n1627 9.3005
R19349 gnd.n5756 gnd.n1628 9.3005
R19350 gnd.n5755 gnd.n1629 9.3005
R19351 gnd.n5754 gnd.n5753 9.3005
R19352 gnd.n1716 gnd.n1647 9.3005
R19353 gnd.n5831 gnd.n1648 9.3005
R19354 gnd.n5832 gnd.n1649 9.3005
R19355 gnd.n5834 gnd.n5833 9.3005
R19356 gnd.n1711 gnd.n1667 9.3005
R19357 gnd.n5846 gnd.n1668 9.3005
R19358 gnd.n5847 gnd.n1669 9.3005
R19359 gnd.n5849 gnd.n5848 9.3005
R19360 gnd.n5850 gnd.n1687 9.3005
R19361 gnd.n5856 gnd.n1688 9.3005
R19362 gnd.n5855 gnd.n1689 9.3005
R19363 gnd.n5854 gnd.n5851 9.3005
R19364 gnd.n5853 gnd.n378 9.3005
R19365 gnd.n7302 gnd.n377 9.3005
R19366 gnd.n7304 gnd.n7303 9.3005
R19367 gnd.n7306 gnd.n373 9.3005
R19368 gnd.n7305 gnd.n371 9.3005
R19369 gnd.n7314 gnd.n370 9.3005
R19370 gnd.n7355 gnd.n7315 9.3005
R19371 gnd.n7354 gnd.n111 9.3005
R19372 gnd.n7353 gnd.n112 9.3005
R19373 gnd.n7351 gnd.n113 9.3005
R19374 gnd.n7350 gnd.n7316 9.3005
R19375 gnd.n7348 gnd.n128 9.3005
R19376 gnd.n7347 gnd.n129 9.3005
R19377 gnd.n7345 gnd.n130 9.3005
R19378 gnd.n7344 gnd.n7317 9.3005
R19379 gnd.n7342 gnd.n148 9.3005
R19380 gnd.n7341 gnd.n149 9.3005
R19381 gnd.n7339 gnd.n150 9.3005
R19382 gnd.n7338 gnd.n7318 9.3005
R19383 gnd.n7336 gnd.n166 9.3005
R19384 gnd.n7335 gnd.n167 9.3005
R19385 gnd.n7333 gnd.n168 9.3005
R19386 gnd.n7332 gnd.n7319 9.3005
R19387 gnd.n7330 gnd.n186 9.3005
R19388 gnd.n7329 gnd.n187 9.3005
R19389 gnd.n7327 gnd.n188 9.3005
R19390 gnd.n7326 gnd.n7320 9.3005
R19391 gnd.n7324 gnd.n205 9.3005
R19392 gnd.n7323 gnd.n206 9.3005
R19393 gnd.n7321 gnd.n207 9.3005
R19394 gnd.n1580 gnd.n1574 9.3005
R19395 gnd.n5967 gnd.n5966 9.3005
R19396 gnd.n5970 gnd.n1572 9.3005
R19397 gnd.n5971 gnd.n1571 9.3005
R19398 gnd.n5974 gnd.n1570 9.3005
R19399 gnd.n5975 gnd.n1569 9.3005
R19400 gnd.n5978 gnd.n1568 9.3005
R19401 gnd.n5979 gnd.n1567 9.3005
R19402 gnd.n5982 gnd.n1566 9.3005
R19403 gnd.n5983 gnd.n1565 9.3005
R19404 gnd.n5986 gnd.n1564 9.3005
R19405 gnd.n5987 gnd.n1563 9.3005
R19406 gnd.n5990 gnd.n1562 9.3005
R19407 gnd.n5991 gnd.n1561 9.3005
R19408 gnd.n5994 gnd.n1560 9.3005
R19409 gnd.n5995 gnd.n1559 9.3005
R19410 gnd.n5998 gnd.n1558 9.3005
R19411 gnd.n5999 gnd.n1557 9.3005
R19412 gnd.n6002 gnd.n1556 9.3005
R19413 gnd.n6003 gnd.n1555 9.3005
R19414 gnd.n6006 gnd.n1554 9.3005
R19415 gnd.n6010 gnd.n1550 9.3005
R19416 gnd.n6011 gnd.n1549 9.3005
R19417 gnd.n6014 gnd.n1548 9.3005
R19418 gnd.n6015 gnd.n1547 9.3005
R19419 gnd.n6018 gnd.n1546 9.3005
R19420 gnd.n6019 gnd.n1545 9.3005
R19421 gnd.n6022 gnd.n1544 9.3005
R19422 gnd.n6023 gnd.n1543 9.3005
R19423 gnd.n6026 gnd.n1542 9.3005
R19424 gnd.n6028 gnd.n1538 9.3005
R19425 gnd.n6031 gnd.n1537 9.3005
R19426 gnd.n6032 gnd.n1536 9.3005
R19427 gnd.n6035 gnd.n1535 9.3005
R19428 gnd.n6036 gnd.n1534 9.3005
R19429 gnd.n6039 gnd.n1533 9.3005
R19430 gnd.n6040 gnd.n1532 9.3005
R19431 gnd.n6043 gnd.n1531 9.3005
R19432 gnd.n6045 gnd.n1528 9.3005
R19433 gnd.n6048 gnd.n1527 9.3005
R19434 gnd.n6049 gnd.n1526 9.3005
R19435 gnd.n6052 gnd.n1525 9.3005
R19436 gnd.n6053 gnd.n1524 9.3005
R19437 gnd.n6056 gnd.n1523 9.3005
R19438 gnd.n6057 gnd.n1522 9.3005
R19439 gnd.n6060 gnd.n1521 9.3005
R19440 gnd.n6061 gnd.n1520 9.3005
R19441 gnd.n6064 gnd.n1519 9.3005
R19442 gnd.n6065 gnd.n1518 9.3005
R19443 gnd.n6068 gnd.n1517 9.3005
R19444 gnd.n6069 gnd.n1516 9.3005
R19445 gnd.n6072 gnd.n1515 9.3005
R19446 gnd.n6074 gnd.n1514 9.3005
R19447 gnd.n6075 gnd.n1513 9.3005
R19448 gnd.n6076 gnd.n1512 9.3005
R19449 gnd.n6077 gnd.n1511 9.3005
R19450 gnd.n6007 gnd.n1551 9.3005
R19451 gnd.n5965 gnd.n5962 9.3005
R19452 gnd.n1593 gnd.n1590 9.3005
R19453 gnd.n5949 gnd.n1594 9.3005
R19454 gnd.n5948 gnd.n1595 9.3005
R19455 gnd.n5947 gnd.n1596 9.3005
R19456 gnd.n1616 gnd.n1597 9.3005
R19457 gnd.n5937 gnd.n1617 9.3005
R19458 gnd.n5936 gnd.n1618 9.3005
R19459 gnd.n5935 gnd.n1619 9.3005
R19460 gnd.n1637 gnd.n1620 9.3005
R19461 gnd.n5925 gnd.n1638 9.3005
R19462 gnd.n5924 gnd.n1639 9.3005
R19463 gnd.n5923 gnd.n1640 9.3005
R19464 gnd.n1656 gnd.n1641 9.3005
R19465 gnd.n5913 gnd.n1657 9.3005
R19466 gnd.n5912 gnd.n1658 9.3005
R19467 gnd.n5911 gnd.n1659 9.3005
R19468 gnd.n1677 gnd.n1660 9.3005
R19469 gnd.n5901 gnd.n1678 9.3005
R19470 gnd.n5900 gnd.n1679 9.3005
R19471 gnd.n5899 gnd.n1680 9.3005
R19472 gnd.n1681 gnd.n97 9.3005
R19473 gnd.n102 gnd.n96 9.3005
R19474 gnd.n7607 gnd.n119 9.3005
R19475 gnd.n7606 gnd.n120 9.3005
R19476 gnd.n7605 gnd.n121 9.3005
R19477 gnd.n138 gnd.n122 9.3005
R19478 gnd.n7595 gnd.n139 9.3005
R19479 gnd.n7594 gnd.n140 9.3005
R19480 gnd.n7593 gnd.n141 9.3005
R19481 gnd.n156 gnd.n142 9.3005
R19482 gnd.n7583 gnd.n157 9.3005
R19483 gnd.n7582 gnd.n158 9.3005
R19484 gnd.n7581 gnd.n159 9.3005
R19485 gnd.n176 gnd.n160 9.3005
R19486 gnd.n7571 gnd.n177 9.3005
R19487 gnd.n7570 gnd.n178 9.3005
R19488 gnd.n7569 gnd.n179 9.3005
R19489 gnd.n196 gnd.n180 9.3005
R19490 gnd.n7559 gnd.n197 9.3005
R19491 gnd.n7558 gnd.n198 9.3005
R19492 gnd.n7557 gnd.n199 9.3005
R19493 gnd.n214 gnd.n200 9.3005
R19494 gnd.n7547 gnd.n7546 9.3005
R19495 gnd.n1592 gnd.n1591 9.3005
R19496 gnd.n7618 gnd.n100 9.3005
R19497 gnd.n7618 gnd.n7617 9.3005
R19498 gnd.n5880 gnd.n5879 9.3005
R19499 gnd.n5881 gnd.n1701 9.3005
R19500 gnd.n5884 gnd.n5883 9.3005
R19501 gnd.n5882 gnd.n389 9.3005
R19502 gnd.n7291 gnd.n390 9.3005
R19503 gnd.n7290 gnd.n7289 9.3005
R19504 gnd.n4644 gnd.n4627 9.3005
R19505 gnd.n4630 gnd.n4628 9.3005
R19506 gnd.n4640 gnd.n4631 9.3005
R19507 gnd.n4639 gnd.n4632 9.3005
R19508 gnd.n4638 gnd.n4633 9.3005
R19509 gnd.n4636 gnd.n4635 9.3005
R19510 gnd.n4634 gnd.n2486 9.3005
R19511 gnd.n2484 gnd.n2483 9.3005
R19512 gnd.n4714 gnd.n4713 9.3005
R19513 gnd.n4715 gnd.n2482 9.3005
R19514 gnd.n4717 gnd.n4716 9.3005
R19515 gnd.n2480 gnd.n2479 9.3005
R19516 gnd.n4722 gnd.n4721 9.3005
R19517 gnd.n4723 gnd.n2478 9.3005
R19518 gnd.n4753 gnd.n4724 9.3005
R19519 gnd.n4752 gnd.n4725 9.3005
R19520 gnd.n4751 gnd.n4726 9.3005
R19521 gnd.n4729 gnd.n4727 9.3005
R19522 gnd.n4747 gnd.n4730 9.3005
R19523 gnd.n4746 gnd.n4731 9.3005
R19524 gnd.n4745 gnd.n4732 9.3005
R19525 gnd.n4736 gnd.n4733 9.3005
R19526 gnd.n4740 gnd.n4737 9.3005
R19527 gnd.n4739 gnd.n4738 9.3005
R19528 gnd.n2201 gnd.n2200 9.3005
R19529 gnd.n4861 gnd.n4860 9.3005
R19530 gnd.n4862 gnd.n2199 9.3005
R19531 gnd.n4864 gnd.n4863 9.3005
R19532 gnd.n2188 gnd.n2187 9.3005
R19533 gnd.n4877 gnd.n4876 9.3005
R19534 gnd.n4878 gnd.n2186 9.3005
R19535 gnd.n4880 gnd.n4879 9.3005
R19536 gnd.n2174 gnd.n2173 9.3005
R19537 gnd.n4893 gnd.n4892 9.3005
R19538 gnd.n4894 gnd.n2172 9.3005
R19539 gnd.n4896 gnd.n4895 9.3005
R19540 gnd.n2159 gnd.n2158 9.3005
R19541 gnd.n4909 gnd.n4908 9.3005
R19542 gnd.n4910 gnd.n2157 9.3005
R19543 gnd.n4912 gnd.n4911 9.3005
R19544 gnd.n2145 gnd.n2144 9.3005
R19545 gnd.n4925 gnd.n4924 9.3005
R19546 gnd.n4926 gnd.n2143 9.3005
R19547 gnd.n4928 gnd.n4927 9.3005
R19548 gnd.n2130 gnd.n2129 9.3005
R19549 gnd.n4967 gnd.n4966 9.3005
R19550 gnd.n4968 gnd.n2128 9.3005
R19551 gnd.n4973 gnd.n4969 9.3005
R19552 gnd.n4972 gnd.n4971 9.3005
R19553 gnd.n4970 gnd.n1190 9.3005
R19554 gnd.n6282 gnd.n1191 9.3005
R19555 gnd.n6281 gnd.n1192 9.3005
R19556 gnd.n6280 gnd.n1193 9.3005
R19557 gnd.n1294 gnd.n1194 9.3005
R19558 gnd.n1295 gnd.n1293 9.3005
R19559 gnd.n6263 gnd.n1296 9.3005
R19560 gnd.n6262 gnd.n1297 9.3005
R19561 gnd.n6261 gnd.n1298 9.3005
R19562 gnd.n2101 gnd.n1299 9.3005
R19563 gnd.n5039 gnd.n5038 9.3005
R19564 gnd.n5040 gnd.n2100 9.3005
R19565 gnd.n5042 gnd.n5041 9.3005
R19566 gnd.n2076 gnd.n2075 9.3005
R19567 gnd.n5098 gnd.n5097 9.3005
R19568 gnd.n5099 gnd.n2074 9.3005
R19569 gnd.n5103 gnd.n5100 9.3005
R19570 gnd.n5102 gnd.n5101 9.3005
R19571 gnd.n2053 gnd.n2052 9.3005
R19572 gnd.n5130 gnd.n5129 9.3005
R19573 gnd.n5131 gnd.n2051 9.3005
R19574 gnd.n5135 gnd.n5132 9.3005
R19575 gnd.n5134 gnd.n5133 9.3005
R19576 gnd.n2031 gnd.n2030 9.3005
R19577 gnd.n5180 gnd.n5179 9.3005
R19578 gnd.n5181 gnd.n2029 9.3005
R19579 gnd.n5185 gnd.n5182 9.3005
R19580 gnd.n5184 gnd.n5183 9.3005
R19581 gnd.n2003 gnd.n2002 9.3005
R19582 gnd.n5218 gnd.n5217 9.3005
R19583 gnd.n5219 gnd.n2001 9.3005
R19584 gnd.n5221 gnd.n5220 9.3005
R19585 gnd.n1975 gnd.n1974 9.3005
R19586 gnd.n5255 gnd.n5254 9.3005
R19587 gnd.n5256 gnd.n1973 9.3005
R19588 gnd.n5260 gnd.n5257 9.3005
R19589 gnd.n5259 gnd.n5258 9.3005
R19590 gnd.n1956 gnd.n1955 9.3005
R19591 gnd.n5313 gnd.n5312 9.3005
R19592 gnd.n5314 gnd.n1954 9.3005
R19593 gnd.n5318 gnd.n5315 9.3005
R19594 gnd.n5317 gnd.n5316 9.3005
R19595 gnd.n1933 gnd.n1932 9.3005
R19596 gnd.n5351 gnd.n5350 9.3005
R19597 gnd.n5352 gnd.n1931 9.3005
R19598 gnd.n5356 gnd.n5353 9.3005
R19599 gnd.n5355 gnd.n5354 9.3005
R19600 gnd.n1905 gnd.n1904 9.3005
R19601 gnd.n5407 gnd.n5406 9.3005
R19602 gnd.n5408 gnd.n1903 9.3005
R19603 gnd.n5412 gnd.n5409 9.3005
R19604 gnd.n5411 gnd.n5410 9.3005
R19605 gnd.n1884 gnd.n1883 9.3005
R19606 gnd.n5445 gnd.n5444 9.3005
R19607 gnd.n5446 gnd.n1882 9.3005
R19608 gnd.n5448 gnd.n5447 9.3005
R19609 gnd.n1828 gnd.n1827 9.3005
R19610 gnd.n5620 gnd.n5619 9.3005
R19611 gnd.n5621 gnd.n1826 9.3005
R19612 gnd.n5623 gnd.n5622 9.3005
R19613 gnd.n1817 gnd.n1816 9.3005
R19614 gnd.n5637 gnd.n5636 9.3005
R19615 gnd.n5638 gnd.n1815 9.3005
R19616 gnd.n5640 gnd.n5639 9.3005
R19617 gnd.n1805 gnd.n1804 9.3005
R19618 gnd.n5654 gnd.n5653 9.3005
R19619 gnd.n5655 gnd.n1803 9.3005
R19620 gnd.n5657 gnd.n5656 9.3005
R19621 gnd.n1793 gnd.n1792 9.3005
R19622 gnd.n5671 gnd.n5670 9.3005
R19623 gnd.n5672 gnd.n1791 9.3005
R19624 gnd.n5674 gnd.n5673 9.3005
R19625 gnd.n1781 gnd.n1780 9.3005
R19626 gnd.n5688 gnd.n5687 9.3005
R19627 gnd.n5689 gnd.n1779 9.3005
R19628 gnd.n5694 gnd.n5690 9.3005
R19629 gnd.n5693 gnd.n5692 9.3005
R19630 gnd.n5691 gnd.n1769 9.3005
R19631 gnd.n5708 gnd.n1768 9.3005
R19632 gnd.n5710 gnd.n5709 9.3005
R19633 gnd.n5711 gnd.n1767 9.3005
R19634 gnd.n5724 gnd.n5712 9.3005
R19635 gnd.n5723 gnd.n5713 9.3005
R19636 gnd.n5722 gnd.n5714 9.3005
R19637 gnd.n5716 gnd.n5715 9.3005
R19638 gnd.n5718 gnd.n5717 9.3005
R19639 gnd.n1733 gnd.n1732 9.3005
R19640 gnd.n5779 gnd.n5778 9.3005
R19641 gnd.n5780 gnd.n1731 9.3005
R19642 gnd.n5782 gnd.n5781 9.3005
R19643 gnd.n1729 gnd.n1728 9.3005
R19644 gnd.n5787 gnd.n5786 9.3005
R19645 gnd.n5788 gnd.n1727 9.3005
R19646 gnd.n5790 gnd.n5789 9.3005
R19647 gnd.n1725 gnd.n1724 9.3005
R19648 gnd.n5795 gnd.n5794 9.3005
R19649 gnd.n5796 gnd.n1723 9.3005
R19650 gnd.n5818 gnd.n5797 9.3005
R19651 gnd.n5817 gnd.n5798 9.3005
R19652 gnd.n5816 gnd.n5799 9.3005
R19653 gnd.n5802 gnd.n5800 9.3005
R19654 gnd.n5812 gnd.n5803 9.3005
R19655 gnd.n5811 gnd.n5804 9.3005
R19656 gnd.n5810 gnd.n5805 9.3005
R19657 gnd.n5808 gnd.n5807 9.3005
R19658 gnd.n5806 gnd.n1705 9.3005
R19659 gnd.n1703 gnd.n1702 9.3005
R19660 gnd.n4280 gnd.n4249 9.3005
R19661 gnd.n4279 gnd.n4250 9.3005
R19662 gnd.n4277 gnd.n4251 9.3005
R19663 gnd.n4276 gnd.n4252 9.3005
R19664 gnd.n4274 gnd.n4253 9.3005
R19665 gnd.n4273 gnd.n4254 9.3005
R19666 gnd.n4271 gnd.n4255 9.3005
R19667 gnd.n4270 gnd.n4256 9.3005
R19668 gnd.n4268 gnd.n4257 9.3005
R19669 gnd.n4267 gnd.n4258 9.3005
R19670 gnd.n4265 gnd.n4259 9.3005
R19671 gnd.n4264 gnd.n4260 9.3005
R19672 gnd.n4262 gnd.n4261 9.3005
R19673 gnd.n2570 gnd.n2569 9.3005
R19674 gnd.n4528 gnd.n4527 9.3005
R19675 gnd.n4529 gnd.n2568 9.3005
R19676 gnd.n4543 gnd.n4530 9.3005
R19677 gnd.n4542 gnd.n4531 9.3005
R19678 gnd.n4541 gnd.n4532 9.3005
R19679 gnd.n4539 gnd.n4533 9.3005
R19680 gnd.n4538 gnd.n4534 9.3005
R19681 gnd.n4536 gnd.n4535 9.3005
R19682 gnd.n2534 gnd.n2533 9.3005
R19683 gnd.n4589 gnd.n4588 9.3005
R19684 gnd.n4590 gnd.n2532 9.3005
R19685 gnd.n4598 gnd.n4591 9.3005
R19686 gnd.n4283 gnd.n4282 9.3005
R19687 gnd.n4288 gnd.n4287 9.3005
R19688 gnd.n4291 gnd.n4244 9.3005
R19689 gnd.n4292 gnd.n4243 9.3005
R19690 gnd.n4295 gnd.n4242 9.3005
R19691 gnd.n4296 gnd.n4241 9.3005
R19692 gnd.n4299 gnd.n4240 9.3005
R19693 gnd.n4300 gnd.n4239 9.3005
R19694 gnd.n4303 gnd.n4238 9.3005
R19695 gnd.n4304 gnd.n4237 9.3005
R19696 gnd.n4307 gnd.n4236 9.3005
R19697 gnd.n4308 gnd.n4235 9.3005
R19698 gnd.n4311 gnd.n4234 9.3005
R19699 gnd.n4312 gnd.n4233 9.3005
R19700 gnd.n4315 gnd.n4232 9.3005
R19701 gnd.n4316 gnd.n4231 9.3005
R19702 gnd.n4319 gnd.n4230 9.3005
R19703 gnd.n4322 gnd.n4321 9.3005
R19704 gnd.n4286 gnd.n4248 9.3005
R19705 gnd.n4285 gnd.n4284 9.3005
R19706 gnd.n6360 gnd.n1116 9.3005
R19707 gnd.n6361 gnd.n1115 9.3005
R19708 gnd.n1114 gnd.n1111 9.3005
R19709 gnd.n6366 gnd.n1110 9.3005
R19710 gnd.n6367 gnd.n1109 9.3005
R19711 gnd.n6368 gnd.n1108 9.3005
R19712 gnd.n1107 gnd.n1104 9.3005
R19713 gnd.n6373 gnd.n1103 9.3005
R19714 gnd.n6375 gnd.n1100 9.3005
R19715 gnd.n6376 gnd.n1099 9.3005
R19716 gnd.n1098 gnd.n1095 9.3005
R19717 gnd.n6381 gnd.n1094 9.3005
R19718 gnd.n6382 gnd.n1093 9.3005
R19719 gnd.n6383 gnd.n1092 9.3005
R19720 gnd.n1091 gnd.n1088 9.3005
R19721 gnd.n6388 gnd.n1087 9.3005
R19722 gnd.n6389 gnd.n1086 9.3005
R19723 gnd.n6390 gnd.n1085 9.3005
R19724 gnd.n1084 gnd.n1081 9.3005
R19725 gnd.n6395 gnd.n1080 9.3005
R19726 gnd.n6396 gnd.n1079 9.3005
R19727 gnd.n6397 gnd.n1078 9.3005
R19728 gnd.n1077 gnd.n1074 9.3005
R19729 gnd.n1076 gnd.n1072 9.3005
R19730 gnd.n6404 gnd.n1071 9.3005
R19731 gnd.n6406 gnd.n6405 9.3005
R19732 gnd.n2311 gnd.n2310 9.3005
R19733 gnd.n2319 gnd.n2318 9.3005
R19734 gnd.n2320 gnd.n2308 9.3005
R19735 gnd.n2322 gnd.n2321 9.3005
R19736 gnd.n2306 gnd.n2305 9.3005
R19737 gnd.n2329 gnd.n2328 9.3005
R19738 gnd.n2330 gnd.n2304 9.3005
R19739 gnd.n2332 gnd.n2331 9.3005
R19740 gnd.n2302 gnd.n2299 9.3005
R19741 gnd.n2339 gnd.n2338 9.3005
R19742 gnd.n2340 gnd.n2298 9.3005
R19743 gnd.n2342 gnd.n2341 9.3005
R19744 gnd.n2296 gnd.n2295 9.3005
R19745 gnd.n2349 gnd.n2348 9.3005
R19746 gnd.n2350 gnd.n2294 9.3005
R19747 gnd.n2352 gnd.n2351 9.3005
R19748 gnd.n2292 gnd.n2291 9.3005
R19749 gnd.n2359 gnd.n2358 9.3005
R19750 gnd.n2360 gnd.n2290 9.3005
R19751 gnd.n2362 gnd.n2361 9.3005
R19752 gnd.n2288 gnd.n2287 9.3005
R19753 gnd.n2369 gnd.n2368 9.3005
R19754 gnd.n2370 gnd.n2286 9.3005
R19755 gnd.n2372 gnd.n2371 9.3005
R19756 gnd.n2284 gnd.n2283 9.3005
R19757 gnd.n2379 gnd.n2378 9.3005
R19758 gnd.n2380 gnd.n2282 9.3005
R19759 gnd.n2382 gnd.n2381 9.3005
R19760 gnd.n2280 gnd.n2277 9.3005
R19761 gnd.n2388 gnd.n2387 9.3005
R19762 gnd.n2309 gnd.n1117 9.3005
R19763 gnd.n4449 gnd.n4448 9.3005
R19764 gnd.n2646 gnd.n2642 9.3005
R19765 gnd.n2645 gnd.n2644 9.3005
R19766 gnd.n2626 gnd.n2623 9.3005
R19767 gnd.n4469 gnd.n2624 9.3005
R19768 gnd.n4468 gnd.n4465 9.3005
R19769 gnd.n4467 gnd.n4466 9.3005
R19770 gnd.n2608 gnd.n2605 9.3005
R19771 gnd.n4489 gnd.n2606 9.3005
R19772 gnd.n4488 gnd.n4485 9.3005
R19773 gnd.n4487 gnd.n4486 9.3005
R19774 gnd.n2590 gnd.n2586 9.3005
R19775 gnd.n4513 gnd.n2587 9.3005
R19776 gnd.n4512 gnd.n2588 9.3005
R19777 gnd.n4511 gnd.n4507 9.3005
R19778 gnd.n4510 gnd.n4508 9.3005
R19779 gnd.n2564 gnd.n2561 9.3005
R19780 gnd.n4554 gnd.n2562 9.3005
R19781 gnd.n4553 gnd.n4550 9.3005
R19782 gnd.n4552 gnd.n4551 9.3005
R19783 gnd.n2547 gnd.n2543 9.3005
R19784 gnd.n4579 gnd.n2544 9.3005
R19785 gnd.n4578 gnd.n2545 9.3005
R19786 gnd.n4577 gnd.n4573 9.3005
R19787 gnd.n4575 gnd.n4574 9.3005
R19788 gnd.n2531 gnd.n2526 9.3005
R19789 gnd.n4611 gnd.n2527 9.3005
R19790 gnd.n4610 gnd.n2528 9.3005
R19791 gnd.n4609 gnd.n4608 9.3005
R19792 gnd.n2529 gnd.n961 9.3005
R19793 gnd.n6474 gnd.n962 9.3005
R19794 gnd.n6473 gnd.n963 9.3005
R19795 gnd.n6472 gnd.n964 9.3005
R19796 gnd.n4661 gnd.n965 9.3005
R19797 gnd.n6462 gnd.n981 9.3005
R19798 gnd.n6461 gnd.n982 9.3005
R19799 gnd.n6460 gnd.n983 9.3005
R19800 gnd.n4676 gnd.n984 9.3005
R19801 gnd.n6450 gnd.n1001 9.3005
R19802 gnd.n6449 gnd.n1002 9.3005
R19803 gnd.n6448 gnd.n1003 9.3005
R19804 gnd.n4683 gnd.n1004 9.3005
R19805 gnd.n6438 gnd.n1021 9.3005
R19806 gnd.n6437 gnd.n1022 9.3005
R19807 gnd.n6436 gnd.n1023 9.3005
R19808 gnd.n2474 gnd.n1024 9.3005
R19809 gnd.n6426 gnd.n1041 9.3005
R19810 gnd.n6425 gnd.n1042 9.3005
R19811 gnd.n6424 gnd.n1043 9.3005
R19812 gnd.n2469 gnd.n1044 9.3005
R19813 gnd.n6414 gnd.n1061 9.3005
R19814 gnd.n6413 gnd.n1062 9.3005
R19815 gnd.n6412 gnd.n1063 9.3005
R19816 gnd.n2643 gnd.n2641 9.3005
R19817 gnd.n4448 gnd.n4447 9.3005
R19818 gnd.n4446 gnd.n2646 9.3005
R19819 gnd.n2645 gnd.n2625 9.3005
R19820 gnd.n4462 gnd.n2626 9.3005
R19821 gnd.n4463 gnd.n2624 9.3005
R19822 gnd.n4465 gnd.n4464 9.3005
R19823 gnd.n4466 gnd.n2607 9.3005
R19824 gnd.n4482 gnd.n2608 9.3005
R19825 gnd.n4483 gnd.n2606 9.3005
R19826 gnd.n4485 gnd.n4484 9.3005
R19827 gnd.n4486 gnd.n2589 9.3005
R19828 gnd.n4502 gnd.n2590 9.3005
R19829 gnd.n4503 gnd.n2587 9.3005
R19830 gnd.n4505 gnd.n2588 9.3005
R19831 gnd.n4507 gnd.n4506 9.3005
R19832 gnd.n4508 gnd.n2563 9.3005
R19833 gnd.n4547 gnd.n2564 9.3005
R19834 gnd.n4548 gnd.n2562 9.3005
R19835 gnd.n4550 gnd.n4549 9.3005
R19836 gnd.n4551 gnd.n2546 9.3005
R19837 gnd.n4568 gnd.n2547 9.3005
R19838 gnd.n4569 gnd.n2544 9.3005
R19839 gnd.n4570 gnd.n2545 9.3005
R19840 gnd.n4573 gnd.n4572 9.3005
R19841 gnd.n4574 gnd.n2530 9.3005
R19842 gnd.n4602 gnd.n2531 9.3005
R19843 gnd.n4603 gnd.n2527 9.3005
R19844 gnd.n4605 gnd.n2528 9.3005
R19845 gnd.n4608 gnd.n4607 9.3005
R19846 gnd.n4606 gnd.n2529 9.3005
R19847 gnd.n2501 gnd.n962 9.3005
R19848 gnd.n4659 gnd.n963 9.3005
R19849 gnd.n4660 gnd.n964 9.3005
R19850 gnd.n4662 gnd.n4661 9.3005
R19851 gnd.n2496 gnd.n981 9.3005
R19852 gnd.n4674 gnd.n982 9.3005
R19853 gnd.n4675 gnd.n983 9.3005
R19854 gnd.n4677 gnd.n4676 9.3005
R19855 gnd.n4678 gnd.n1001 9.3005
R19856 gnd.n4681 gnd.n1002 9.3005
R19857 gnd.n4682 gnd.n1003 9.3005
R19858 gnd.n4687 gnd.n4683 9.3005
R19859 gnd.n4688 gnd.n1021 9.3005
R19860 gnd.n4689 gnd.n1022 9.3005
R19861 gnd.n2473 gnd.n1023 9.3005
R19862 gnd.n4758 gnd.n2474 9.3005
R19863 gnd.n4759 gnd.n1041 9.3005
R19864 gnd.n4760 gnd.n1042 9.3005
R19865 gnd.n2468 gnd.n1043 9.3005
R19866 gnd.n4773 gnd.n2469 9.3005
R19867 gnd.n4774 gnd.n1061 9.3005
R19868 gnd.n4776 gnd.n1062 9.3005
R19869 gnd.n4775 gnd.n1063 9.3005
R19870 gnd.n4445 gnd.n2643 9.3005
R19871 gnd.n4326 gnd.n4325 9.3005
R19872 gnd.n4328 gnd.n4227 9.3005
R19873 gnd.n4329 gnd.n4226 9.3005
R19874 gnd.n4332 gnd.n4225 9.3005
R19875 gnd.n4333 gnd.n4224 9.3005
R19876 gnd.n4336 gnd.n4223 9.3005
R19877 gnd.n4337 gnd.n4222 9.3005
R19878 gnd.n4340 gnd.n4221 9.3005
R19879 gnd.n4341 gnd.n4220 9.3005
R19880 gnd.n4344 gnd.n4219 9.3005
R19881 gnd.n4345 gnd.n4218 9.3005
R19882 gnd.n4348 gnd.n4217 9.3005
R19883 gnd.n4349 gnd.n4216 9.3005
R19884 gnd.n4352 gnd.n4215 9.3005
R19885 gnd.n4353 gnd.n4214 9.3005
R19886 gnd.n4356 gnd.n4213 9.3005
R19887 gnd.n4357 gnd.n4212 9.3005
R19888 gnd.n4360 gnd.n4211 9.3005
R19889 gnd.n4361 gnd.n4210 9.3005
R19890 gnd.n4364 gnd.n4209 9.3005
R19891 gnd.n4368 gnd.n4205 9.3005
R19892 gnd.n4369 gnd.n4204 9.3005
R19893 gnd.n4372 gnd.n4203 9.3005
R19894 gnd.n4373 gnd.n4202 9.3005
R19895 gnd.n4376 gnd.n4201 9.3005
R19896 gnd.n4377 gnd.n4200 9.3005
R19897 gnd.n4380 gnd.n4199 9.3005
R19898 gnd.n4381 gnd.n4198 9.3005
R19899 gnd.n4384 gnd.n4197 9.3005
R19900 gnd.n4385 gnd.n4196 9.3005
R19901 gnd.n4388 gnd.n4195 9.3005
R19902 gnd.n4389 gnd.n4194 9.3005
R19903 gnd.n4392 gnd.n4193 9.3005
R19904 gnd.n4393 gnd.n4192 9.3005
R19905 gnd.n4396 gnd.n4191 9.3005
R19906 gnd.n4397 gnd.n4190 9.3005
R19907 gnd.n4400 gnd.n4189 9.3005
R19908 gnd.n4401 gnd.n4188 9.3005
R19909 gnd.n4404 gnd.n4187 9.3005
R19910 gnd.n4406 gnd.n4184 9.3005
R19911 gnd.n4409 gnd.n4183 9.3005
R19912 gnd.n4410 gnd.n4182 9.3005
R19913 gnd.n4413 gnd.n4181 9.3005
R19914 gnd.n4414 gnd.n4180 9.3005
R19915 gnd.n4417 gnd.n4179 9.3005
R19916 gnd.n4418 gnd.n4178 9.3005
R19917 gnd.n4421 gnd.n4177 9.3005
R19918 gnd.n4422 gnd.n4176 9.3005
R19919 gnd.n4425 gnd.n4175 9.3005
R19920 gnd.n4426 gnd.n4174 9.3005
R19921 gnd.n4429 gnd.n4173 9.3005
R19922 gnd.n4430 gnd.n4172 9.3005
R19923 gnd.n4433 gnd.n4171 9.3005
R19924 gnd.n4435 gnd.n4170 9.3005
R19925 gnd.n4436 gnd.n4169 9.3005
R19926 gnd.n4437 gnd.n4168 9.3005
R19927 gnd.n4438 gnd.n4167 9.3005
R19928 gnd.n4365 gnd.n4206 9.3005
R19929 gnd.n4324 gnd.n2647 9.3005
R19930 gnd.n4454 gnd.n4453 9.3005
R19931 gnd.n4455 gnd.n2632 9.3005
R19932 gnd.n4457 gnd.n4456 9.3005
R19933 gnd.n2615 gnd.n2614 9.3005
R19934 gnd.n4474 gnd.n4473 9.3005
R19935 gnd.n4475 gnd.n2613 9.3005
R19936 gnd.n4477 gnd.n4476 9.3005
R19937 gnd.n2598 gnd.n2597 9.3005
R19938 gnd.n4494 gnd.n4493 9.3005
R19939 gnd.n4495 gnd.n2596 9.3005
R19940 gnd.n4497 gnd.n4496 9.3005
R19941 gnd.n2578 gnd.n2577 9.3005
R19942 gnd.n4518 gnd.n4517 9.3005
R19943 gnd.n4519 gnd.n2576 9.3005
R19944 gnd.n4523 gnd.n4520 9.3005
R19945 gnd.n4522 gnd.n4521 9.3005
R19946 gnd.n2554 gnd.n2553 9.3005
R19947 gnd.n4559 gnd.n4558 9.3005
R19948 gnd.n4560 gnd.n2552 9.3005
R19949 gnd.n4563 gnd.n4561 9.3005
R19950 gnd.n4562 gnd.n947 9.3005
R19951 gnd.n953 gnd.n946 9.3005
R19952 gnd.n6468 gnd.n971 9.3005
R19953 gnd.n6467 gnd.n972 9.3005
R19954 gnd.n6466 gnd.n973 9.3005
R19955 gnd.n991 gnd.n974 9.3005
R19956 gnd.n6456 gnd.n992 9.3005
R19957 gnd.n6455 gnd.n993 9.3005
R19958 gnd.n6454 gnd.n994 9.3005
R19959 gnd.n1010 gnd.n995 9.3005
R19960 gnd.n6444 gnd.n1011 9.3005
R19961 gnd.n6443 gnd.n1012 9.3005
R19962 gnd.n6442 gnd.n1013 9.3005
R19963 gnd.n1031 gnd.n1014 9.3005
R19964 gnd.n6432 gnd.n1032 9.3005
R19965 gnd.n6431 gnd.n1033 9.3005
R19966 gnd.n6430 gnd.n1034 9.3005
R19967 gnd.n1051 gnd.n1035 9.3005
R19968 gnd.n6420 gnd.n1052 9.3005
R19969 gnd.n6419 gnd.n1053 9.3005
R19970 gnd.n6418 gnd.n1054 9.3005
R19971 gnd.n1070 gnd.n1055 9.3005
R19972 gnd.n6408 gnd.n6407 9.3005
R19973 gnd.n2634 gnd.n2633 9.3005
R19974 gnd.n6479 gnd.n944 9.3005
R19975 gnd.n6479 gnd.n6478 9.3005
R19976 gnd.n2514 gnd.n2513 9.3005
R19977 gnd.n4623 gnd.n4622 9.3005
R19978 gnd.n4624 gnd.n2510 9.3005
R19979 gnd.n4646 gnd.n4625 9.3005
R19980 gnd.n4645 gnd.n4626 9.3005
R19981 gnd.n2512 gnd.n2511 9.3005
R19982 gnd.n6487 gnd.n935 9.3005
R19983 gnd.n6488 gnd.n934 9.3005
R19984 gnd.n933 gnd.n929 9.3005
R19985 gnd.n6494 gnd.n928 9.3005
R19986 gnd.n6495 gnd.n927 9.3005
R19987 gnd.n6496 gnd.n926 9.3005
R19988 gnd.n925 gnd.n921 9.3005
R19989 gnd.n6502 gnd.n920 9.3005
R19990 gnd.n6503 gnd.n919 9.3005
R19991 gnd.n6504 gnd.n918 9.3005
R19992 gnd.n917 gnd.n913 9.3005
R19993 gnd.n6510 gnd.n912 9.3005
R19994 gnd.n6511 gnd.n911 9.3005
R19995 gnd.n6512 gnd.n910 9.3005
R19996 gnd.n909 gnd.n905 9.3005
R19997 gnd.n6518 gnd.n904 9.3005
R19998 gnd.n6519 gnd.n903 9.3005
R19999 gnd.n6520 gnd.n902 9.3005
R20000 gnd.n901 gnd.n897 9.3005
R20001 gnd.n6526 gnd.n896 9.3005
R20002 gnd.n6527 gnd.n895 9.3005
R20003 gnd.n6528 gnd.n894 9.3005
R20004 gnd.n893 gnd.n889 9.3005
R20005 gnd.n6534 gnd.n888 9.3005
R20006 gnd.n6535 gnd.n887 9.3005
R20007 gnd.n6536 gnd.n886 9.3005
R20008 gnd.n885 gnd.n881 9.3005
R20009 gnd.n6542 gnd.n880 9.3005
R20010 gnd.n6543 gnd.n879 9.3005
R20011 gnd.n6544 gnd.n878 9.3005
R20012 gnd.n877 gnd.n873 9.3005
R20013 gnd.n6550 gnd.n872 9.3005
R20014 gnd.n6551 gnd.n871 9.3005
R20015 gnd.n6552 gnd.n870 9.3005
R20016 gnd.n869 gnd.n865 9.3005
R20017 gnd.n6558 gnd.n864 9.3005
R20018 gnd.n6559 gnd.n863 9.3005
R20019 gnd.n6560 gnd.n862 9.3005
R20020 gnd.n861 gnd.n857 9.3005
R20021 gnd.n6566 gnd.n856 9.3005
R20022 gnd.n6567 gnd.n855 9.3005
R20023 gnd.n6568 gnd.n854 9.3005
R20024 gnd.n853 gnd.n849 9.3005
R20025 gnd.n6574 gnd.n848 9.3005
R20026 gnd.n6575 gnd.n847 9.3005
R20027 gnd.n6576 gnd.n846 9.3005
R20028 gnd.n845 gnd.n841 9.3005
R20029 gnd.n6582 gnd.n840 9.3005
R20030 gnd.n6583 gnd.n839 9.3005
R20031 gnd.n6584 gnd.n838 9.3005
R20032 gnd.n837 gnd.n833 9.3005
R20033 gnd.n6590 gnd.n832 9.3005
R20034 gnd.n6591 gnd.n831 9.3005
R20035 gnd.n6592 gnd.n830 9.3005
R20036 gnd.n829 gnd.n825 9.3005
R20037 gnd.n6598 gnd.n824 9.3005
R20038 gnd.n6599 gnd.n823 9.3005
R20039 gnd.n6600 gnd.n822 9.3005
R20040 gnd.n821 gnd.n817 9.3005
R20041 gnd.n6606 gnd.n816 9.3005
R20042 gnd.n6607 gnd.n815 9.3005
R20043 gnd.n6608 gnd.n814 9.3005
R20044 gnd.n813 gnd.n809 9.3005
R20045 gnd.n6614 gnd.n808 9.3005
R20046 gnd.n6615 gnd.n807 9.3005
R20047 gnd.n6616 gnd.n806 9.3005
R20048 gnd.n805 gnd.n801 9.3005
R20049 gnd.n6622 gnd.n800 9.3005
R20050 gnd.n6623 gnd.n799 9.3005
R20051 gnd.n6624 gnd.n798 9.3005
R20052 gnd.n797 gnd.n793 9.3005
R20053 gnd.n6630 gnd.n792 9.3005
R20054 gnd.n6631 gnd.n791 9.3005
R20055 gnd.n6632 gnd.n790 9.3005
R20056 gnd.n789 gnd.n785 9.3005
R20057 gnd.n6638 gnd.n784 9.3005
R20058 gnd.n6639 gnd.n783 9.3005
R20059 gnd.n6640 gnd.n782 9.3005
R20060 gnd.n781 gnd.n777 9.3005
R20061 gnd.n6646 gnd.n776 9.3005
R20062 gnd.n6647 gnd.n775 9.3005
R20063 gnd.n6648 gnd.n774 9.3005
R20064 gnd.n770 gnd.n769 9.3005
R20065 gnd.n6655 gnd.n6654 9.3005
R20066 gnd.n6486 gnd.n936 9.3005
R20067 gnd.n5730 gnd.n1737 9.3005
R20068 gnd.n4870 gnd.n2192 9.3005
R20069 gnd.n4872 gnd.n4871 9.3005
R20070 gnd.n2181 gnd.n2180 9.3005
R20071 gnd.n4885 gnd.n4884 9.3005
R20072 gnd.n4886 gnd.n2179 9.3005
R20073 gnd.n4888 gnd.n4887 9.3005
R20074 gnd.n2167 gnd.n2166 9.3005
R20075 gnd.n4901 gnd.n4900 9.3005
R20076 gnd.n4902 gnd.n2165 9.3005
R20077 gnd.n4904 gnd.n4903 9.3005
R20078 gnd.n2153 gnd.n2152 9.3005
R20079 gnd.n4917 gnd.n4916 9.3005
R20080 gnd.n4918 gnd.n2151 9.3005
R20081 gnd.n4920 gnd.n4919 9.3005
R20082 gnd.n2139 gnd.n2138 9.3005
R20083 gnd.n4933 gnd.n4932 9.3005
R20084 gnd.n4934 gnd.n2136 9.3005
R20085 gnd.n4962 gnd.n4961 9.3005
R20086 gnd.n4960 gnd.n2137 9.3005
R20087 gnd.n4959 gnd.n4958 9.3005
R20088 gnd.n4957 gnd.n4935 9.3005
R20089 gnd.n4956 gnd.n4955 9.3005
R20090 gnd.n4954 gnd.n4938 9.3005
R20091 gnd.n4953 gnd.n4952 9.3005
R20092 gnd.n4951 gnd.n4939 9.3005
R20093 gnd.n4950 gnd.n4949 9.3005
R20094 gnd.n4948 gnd.n4945 9.3005
R20095 gnd.n4947 gnd.n4946 9.3005
R20096 gnd.n1307 gnd.n1305 9.3005
R20097 gnd.n6257 gnd.n6256 9.3005
R20098 gnd.n6255 gnd.n1306 9.3005
R20099 gnd.n6254 gnd.n6253 9.3005
R20100 gnd.n6252 gnd.n1308 9.3005
R20101 gnd.n6251 gnd.n6250 9.3005
R20102 gnd.n6249 gnd.n1312 9.3005
R20103 gnd.n6248 gnd.n6247 9.3005
R20104 gnd.n6246 gnd.n1313 9.3005
R20105 gnd.n6245 gnd.n6244 9.3005
R20106 gnd.n6243 gnd.n1317 9.3005
R20107 gnd.n6242 gnd.n6241 9.3005
R20108 gnd.n6240 gnd.n1318 9.3005
R20109 gnd.n6239 gnd.n6238 9.3005
R20110 gnd.n6237 gnd.n1322 9.3005
R20111 gnd.n6236 gnd.n6235 9.3005
R20112 gnd.n6234 gnd.n1323 9.3005
R20113 gnd.n6233 gnd.n6232 9.3005
R20114 gnd.n6231 gnd.n1327 9.3005
R20115 gnd.n6230 gnd.n6229 9.3005
R20116 gnd.n6228 gnd.n1328 9.3005
R20117 gnd.n6227 gnd.n6226 9.3005
R20118 gnd.n6225 gnd.n1332 9.3005
R20119 gnd.n6224 gnd.n6223 9.3005
R20120 gnd.n6222 gnd.n1333 9.3005
R20121 gnd.n6221 gnd.n6220 9.3005
R20122 gnd.n6219 gnd.n1337 9.3005
R20123 gnd.n6218 gnd.n6217 9.3005
R20124 gnd.n6216 gnd.n1338 9.3005
R20125 gnd.n6215 gnd.n6214 9.3005
R20126 gnd.n6213 gnd.n1342 9.3005
R20127 gnd.n6212 gnd.n6211 9.3005
R20128 gnd.n6210 gnd.n1343 9.3005
R20129 gnd.n6209 gnd.n6208 9.3005
R20130 gnd.n6207 gnd.n1347 9.3005
R20131 gnd.n6206 gnd.n6205 9.3005
R20132 gnd.n6204 gnd.n1348 9.3005
R20133 gnd.n6203 gnd.n6202 9.3005
R20134 gnd.n6201 gnd.n1352 9.3005
R20135 gnd.n6200 gnd.n6199 9.3005
R20136 gnd.n6198 gnd.n1353 9.3005
R20137 gnd.n6197 gnd.n6196 9.3005
R20138 gnd.n6195 gnd.n1357 9.3005
R20139 gnd.n6194 gnd.n6193 9.3005
R20140 gnd.n6192 gnd.n1358 9.3005
R20141 gnd.n6191 gnd.n6190 9.3005
R20142 gnd.n6189 gnd.n1362 9.3005
R20143 gnd.n6188 gnd.n6187 9.3005
R20144 gnd.n6186 gnd.n1363 9.3005
R20145 gnd.n6185 gnd.n6184 9.3005
R20146 gnd.n6183 gnd.n1367 9.3005
R20147 gnd.n6182 gnd.n6181 9.3005
R20148 gnd.n6180 gnd.n1368 9.3005
R20149 gnd.n6179 gnd.n6178 9.3005
R20150 gnd.n6177 gnd.n1372 9.3005
R20151 gnd.n6176 gnd.n6175 9.3005
R20152 gnd.n6174 gnd.n1373 9.3005
R20153 gnd.n6173 gnd.n6172 9.3005
R20154 gnd.n6171 gnd.n1377 9.3005
R20155 gnd.n6170 gnd.n6169 9.3005
R20156 gnd.n6168 gnd.n1378 9.3005
R20157 gnd.n6167 gnd.n6166 9.3005
R20158 gnd.n6165 gnd.n1382 9.3005
R20159 gnd.n6164 gnd.n6163 9.3005
R20160 gnd.n6162 gnd.n1383 9.3005
R20161 gnd.n6161 gnd.n6160 9.3005
R20162 gnd.n6159 gnd.n1387 9.3005
R20163 gnd.n6158 gnd.n6157 9.3005
R20164 gnd.n6156 gnd.n1388 9.3005
R20165 gnd.n6155 gnd.n6154 9.3005
R20166 gnd.n6153 gnd.n1392 9.3005
R20167 gnd.n6152 gnd.n6151 9.3005
R20168 gnd.n6150 gnd.n1393 9.3005
R20169 gnd.n4869 gnd.n4868 9.3005
R20170 gnd.n4789 gnd.n2193 9.3005
R20171 gnd.n4597 gnd.n4596 9.3005
R20172 gnd.n4595 gnd.n4593 9.3005
R20173 gnd.n2504 gnd.n2503 9.3005
R20174 gnd.n4652 gnd.n4651 9.3005
R20175 gnd.n4653 gnd.n2502 9.3005
R20176 gnd.n4655 gnd.n4654 9.3005
R20177 gnd.n2499 gnd.n2498 9.3005
R20178 gnd.n4667 gnd.n4666 9.3005
R20179 gnd.n4668 gnd.n2497 9.3005
R20180 gnd.n4670 gnd.n4669 9.3005
R20181 gnd.n2490 gnd.n2488 9.3005
R20182 gnd.n4706 gnd.n4705 9.3005
R20183 gnd.n4704 gnd.n2489 9.3005
R20184 gnd.n4703 gnd.n4702 9.3005
R20185 gnd.n4701 gnd.n2491 9.3005
R20186 gnd.n4700 gnd.n4699 9.3005
R20187 gnd.n4698 gnd.n2494 9.3005
R20188 gnd.n4697 gnd.n4696 9.3005
R20189 gnd.n4695 gnd.n2495 9.3005
R20190 gnd.n4694 gnd.n4693 9.3005
R20191 gnd.n2472 gnd.n2471 9.3005
R20192 gnd.n4765 gnd.n4764 9.3005
R20193 gnd.n4766 gnd.n2470 9.3005
R20194 gnd.n4769 gnd.n4768 9.3005
R20195 gnd.n4767 gnd.n2466 9.3005
R20196 gnd.n4780 gnd.n2465 9.3005
R20197 gnd.n4782 gnd.n4781 9.3005
R20198 gnd.n4838 gnd.n4837 9.3005
R20199 gnd.n4836 gnd.n4835 9.3005
R20200 gnd.n2403 gnd.n2402 9.3005
R20201 gnd.n4830 gnd.n4829 9.3005
R20202 gnd.n4828 gnd.n4827 9.3005
R20203 gnd.n2415 gnd.n2414 9.3005
R20204 gnd.n4822 gnd.n4821 9.3005
R20205 gnd.n4820 gnd.n4819 9.3005
R20206 gnd.n2426 gnd.n2425 9.3005
R20207 gnd.n4814 gnd.n4813 9.3005
R20208 gnd.n4812 gnd.n4811 9.3005
R20209 gnd.n2438 gnd.n2437 9.3005
R20210 gnd.n4806 gnd.n4805 9.3005
R20211 gnd.n4804 gnd.n4803 9.3005
R20212 gnd.n2449 gnd.n2448 9.3005
R20213 gnd.n4798 gnd.n4797 9.3005
R20214 gnd.n4796 gnd.n2462 9.3005
R20215 gnd.n4795 gnd.n4792 9.3005
R20216 gnd.n2398 gnd.n2396 9.3005
R20217 gnd.n4791 gnd.n4790 9.3005
R20218 gnd.n4786 gnd.n2464 9.3005
R20219 gnd.n4785 gnd.n2456 9.3005
R20220 gnd.n4800 gnd.n4799 9.3005
R20221 gnd.n4802 gnd.n4801 9.3005
R20222 gnd.n2442 gnd.n2441 9.3005
R20223 gnd.n4808 gnd.n4807 9.3005
R20224 gnd.n4810 gnd.n4809 9.3005
R20225 gnd.n2432 gnd.n2431 9.3005
R20226 gnd.n4816 gnd.n4815 9.3005
R20227 gnd.n4818 gnd.n4817 9.3005
R20228 gnd.n2419 gnd.n2418 9.3005
R20229 gnd.n4824 gnd.n4823 9.3005
R20230 gnd.n4826 gnd.n4825 9.3005
R20231 gnd.n2409 gnd.n2408 9.3005
R20232 gnd.n4832 gnd.n4831 9.3005
R20233 gnd.n4834 gnd.n4833 9.3005
R20234 gnd.n2397 gnd.n2395 9.3005
R20235 gnd.n4840 gnd.n4839 9.3005
R20236 gnd.n4841 gnd.n2390 9.3005
R20237 gnd.n4843 gnd.n4842 9.3005
R20238 gnd.n4845 gnd.n2276 9.3005
R20239 gnd.n4847 gnd.n4846 9.3005
R20240 gnd.n4848 gnd.n2272 9.3005
R20241 gnd.n4850 gnd.n4849 9.3005
R20242 gnd.n4851 gnd.n2271 9.3005
R20243 gnd.n4853 gnd.n4852 9.3005
R20244 gnd.n4854 gnd.n2270 9.3005
R20245 gnd.n2267 gnd.n2219 9.3005
R20246 gnd.n2266 gnd.n2265 9.3005
R20247 gnd.n2264 gnd.n2222 9.3005
R20248 gnd.n2263 gnd.n2262 9.3005
R20249 gnd.n2261 gnd.n2223 9.3005
R20250 gnd.n2260 gnd.n2259 9.3005
R20251 gnd.n2258 gnd.n2226 9.3005
R20252 gnd.n2257 gnd.n2256 9.3005
R20253 gnd.n2255 gnd.n2227 9.3005
R20254 gnd.n2254 gnd.n2253 9.3005
R20255 gnd.n2252 gnd.n2230 9.3005
R20256 gnd.n2251 gnd.n2250 9.3005
R20257 gnd.n2249 gnd.n2231 9.3005
R20258 gnd.n2248 gnd.n2247 9.3005
R20259 gnd.n2246 gnd.n2234 9.3005
R20260 gnd.n2245 gnd.n2244 9.3005
R20261 gnd.n2243 gnd.n2235 9.3005
R20262 gnd.n2242 gnd.n2241 9.3005
R20263 gnd.n2240 gnd.n2237 9.3005
R20264 gnd.n2239 gnd.n2123 9.3005
R20265 gnd.n2238 gnd.n2121 9.3005
R20266 gnd.n4979 gnd.n2120 9.3005
R20267 gnd.n4981 gnd.n4980 9.3005
R20268 gnd.n4982 gnd.n2119 9.3005
R20269 gnd.n4984 gnd.n4983 9.3005
R20270 gnd.n4985 gnd.n2118 9.3005
R20271 gnd.n4989 gnd.n4988 9.3005
R20272 gnd.n4990 gnd.n2116 9.3005
R20273 gnd.n5008 gnd.n5007 9.3005
R20274 gnd.n5006 gnd.n2117 9.3005
R20275 gnd.n5005 gnd.n5004 9.3005
R20276 gnd.n5003 gnd.n4991 9.3005
R20277 gnd.n5002 gnd.n5001 9.3005
R20278 gnd.n5000 gnd.n4994 9.3005
R20279 gnd.n4999 gnd.n4998 9.3005
R20280 gnd.n4997 gnd.n4995 9.3005
R20281 gnd.n2069 gnd.n2068 9.3005
R20282 gnd.n5108 gnd.n5107 9.3005
R20283 gnd.n5109 gnd.n2066 9.3005
R20284 gnd.n5112 gnd.n5111 9.3005
R20285 gnd.n5110 gnd.n2067 9.3005
R20286 gnd.n2044 gnd.n2043 9.3005
R20287 gnd.n5140 gnd.n5139 9.3005
R20288 gnd.n5141 gnd.n2041 9.3005
R20289 gnd.n5167 gnd.n5166 9.3005
R20290 gnd.n5165 gnd.n2042 9.3005
R20291 gnd.n5164 gnd.n5163 9.3005
R20292 gnd.n5162 gnd.n5142 9.3005
R20293 gnd.n5161 gnd.n5160 9.3005
R20294 gnd.n5159 gnd.n5146 9.3005
R20295 gnd.n5158 gnd.n5157 9.3005
R20296 gnd.n5156 gnd.n5147 9.3005
R20297 gnd.n5155 gnd.n5154 9.3005
R20298 gnd.n5153 gnd.n5150 9.3005
R20299 gnd.n5152 gnd.n5151 9.3005
R20300 gnd.n1968 gnd.n1967 9.3005
R20301 gnd.n5265 gnd.n5264 9.3005
R20302 gnd.n5266 gnd.n1965 9.3005
R20303 gnd.n5298 gnd.n5297 9.3005
R20304 gnd.n5296 gnd.n1966 9.3005
R20305 gnd.n5295 gnd.n5294 9.3005
R20306 gnd.n5293 gnd.n5267 9.3005
R20307 gnd.n5292 gnd.n5291 9.3005
R20308 gnd.n5290 gnd.n5272 9.3005
R20309 gnd.n5289 gnd.n5288 9.3005
R20310 gnd.n5287 gnd.n5273 9.3005
R20311 gnd.n5286 gnd.n5285 9.3005
R20312 gnd.n5284 gnd.n5275 9.3005
R20313 gnd.n5283 gnd.n5282 9.3005
R20314 gnd.n5281 gnd.n5276 9.3005
R20315 gnd.n1897 gnd.n1896 9.3005
R20316 gnd.n5417 gnd.n5416 9.3005
R20317 gnd.n5418 gnd.n1894 9.3005
R20318 gnd.n5431 gnd.n5430 9.3005
R20319 gnd.n5429 gnd.n1895 9.3005
R20320 gnd.n5428 gnd.n5427 9.3005
R20321 gnd.n5426 gnd.n5419 9.3005
R20322 gnd.n5425 gnd.n5424 9.3005
R20323 gnd.n5423 gnd.n5422 9.3005
R20324 gnd.n1823 gnd.n1822 9.3005
R20325 gnd.n5628 gnd.n5627 9.3005
R20326 gnd.n5629 gnd.n1821 9.3005
R20327 gnd.n5631 gnd.n5630 9.3005
R20328 gnd.n1811 gnd.n1810 9.3005
R20329 gnd.n5645 gnd.n5644 9.3005
R20330 gnd.n5646 gnd.n1809 9.3005
R20331 gnd.n5648 gnd.n5647 9.3005
R20332 gnd.n1799 gnd.n1798 9.3005
R20333 gnd.n5662 gnd.n5661 9.3005
R20334 gnd.n5663 gnd.n1797 9.3005
R20335 gnd.n5665 gnd.n5664 9.3005
R20336 gnd.n1786 gnd.n1785 9.3005
R20337 gnd.n5679 gnd.n5678 9.3005
R20338 gnd.n5680 gnd.n1784 9.3005
R20339 gnd.n5682 gnd.n5681 9.3005
R20340 gnd.n1775 gnd.n1774 9.3005
R20341 gnd.n5699 gnd.n5698 9.3005
R20342 gnd.n5700 gnd.n1773 9.3005
R20343 gnd.n5702 gnd.n5701 9.3005
R20344 gnd.n1402 gnd.n1401 9.3005
R20345 gnd.n6146 gnd.n6145 9.3005
R20346 gnd.n2269 gnd.n2268 9.3005
R20347 gnd.n6142 gnd.n1403 9.3005
R20348 gnd.n6141 gnd.n6140 9.3005
R20349 gnd.n6139 gnd.n1406 9.3005
R20350 gnd.n6138 gnd.n6137 9.3005
R20351 gnd.n6136 gnd.n1407 9.3005
R20352 gnd.n6135 gnd.n6134 9.3005
R20353 gnd.n6144 gnd.n6143 9.3005
R20354 gnd.n6087 gnd.n6086 9.3005
R20355 gnd.n1454 gnd.n1453 9.3005
R20356 gnd.n6093 gnd.n6092 9.3005
R20357 gnd.n6095 gnd.n6094 9.3005
R20358 gnd.n1446 gnd.n1445 9.3005
R20359 gnd.n6101 gnd.n6100 9.3005
R20360 gnd.n6103 gnd.n6102 9.3005
R20361 gnd.n1438 gnd.n1437 9.3005
R20362 gnd.n6109 gnd.n6108 9.3005
R20363 gnd.n6111 gnd.n6110 9.3005
R20364 gnd.n1430 gnd.n1429 9.3005
R20365 gnd.n6117 gnd.n6116 9.3005
R20366 gnd.n6119 gnd.n6118 9.3005
R20367 gnd.n1422 gnd.n1421 9.3005
R20368 gnd.n6125 gnd.n6124 9.3005
R20369 gnd.n6127 gnd.n6126 9.3005
R20370 gnd.n1418 gnd.n1413 9.3005
R20371 gnd.n6085 gnd.n1463 9.3005
R20372 gnd.n1738 gnd.n1462 9.3005
R20373 gnd.n6132 gnd.n1411 9.3005
R20374 gnd.n6131 gnd.n6130 9.3005
R20375 gnd.n6129 gnd.n6128 9.3005
R20376 gnd.n1417 gnd.n1416 9.3005
R20377 gnd.n6123 gnd.n6122 9.3005
R20378 gnd.n6121 gnd.n6120 9.3005
R20379 gnd.n1426 gnd.n1425 9.3005
R20380 gnd.n6115 gnd.n6114 9.3005
R20381 gnd.n6113 gnd.n6112 9.3005
R20382 gnd.n1434 gnd.n1433 9.3005
R20383 gnd.n6107 gnd.n6106 9.3005
R20384 gnd.n6105 gnd.n6104 9.3005
R20385 gnd.n1442 gnd.n1441 9.3005
R20386 gnd.n6099 gnd.n6098 9.3005
R20387 gnd.n6097 gnd.n6096 9.3005
R20388 gnd.n1450 gnd.n1449 9.3005
R20389 gnd.n6091 gnd.n6090 9.3005
R20390 gnd.n6089 gnd.n6088 9.3005
R20391 gnd.n1761 gnd.n1460 9.3005
R20392 gnd.n1740 gnd.n1739 9.3005
R20393 gnd.n5732 gnd.n5731 9.3005
R20394 gnd.n5773 gnd.n5772 9.3005
R20395 gnd.n5771 gnd.n1736 9.3005
R20396 gnd.n5770 gnd.n5769 9.3005
R20397 gnd.n5768 gnd.n5735 9.3005
R20398 gnd.n5767 gnd.n5766 9.3005
R20399 gnd.n5765 gnd.n5739 9.3005
R20400 gnd.n5764 gnd.n5763 9.3005
R20401 gnd.n5762 gnd.n5740 9.3005
R20402 gnd.n5761 gnd.n5760 9.3005
R20403 gnd.n1719 gnd.n1718 9.3005
R20404 gnd.n5824 gnd.n5823 9.3005
R20405 gnd.n5825 gnd.n1717 9.3005
R20406 gnd.n5827 gnd.n5826 9.3005
R20407 gnd.n1714 gnd.n1713 9.3005
R20408 gnd.n5839 gnd.n5838 9.3005
R20409 gnd.n5840 gnd.n1712 9.3005
R20410 gnd.n5842 gnd.n5841 9.3005
R20411 gnd.n1709 gnd.n1707 9.3005
R20412 gnd.n5872 gnd.n5871 9.3005
R20413 gnd.n5870 gnd.n1708 9.3005
R20414 gnd.n5869 gnd.n5868 9.3005
R20415 gnd.n5867 gnd.n1710 9.3005
R20416 gnd.n5866 gnd.n5865 9.3005
R20417 gnd.n5864 gnd.n5861 9.3005
R20418 gnd.n5863 gnd.n5862 9.3005
R20419 gnd.n85 gnd.n83 9.3005
R20420 gnd.n5734 gnd.n1735 9.3005
R20421 gnd.t349 gnd.n2839 9.24152
R20422 gnd.n2741 gnd.t106 9.24152
R20423 gnd.n4026 gnd.t84 9.24152
R20424 gnd.t22 gnd.n2628 9.24152
R20425 gnd.n4684 gnd.t276 9.24152
R20426 gnd.n6416 gnd.t55 9.24152
R20427 gnd.n5951 gnd.t12 9.24152
R20428 gnd.n5820 gnd.t222 9.24152
R20429 gnd.n7555 gnd.t37 9.24152
R20430 gnd.t146 gnd.t349 8.92286
R20431 gnd.n6266 gnd.n6265 8.92286
R20432 gnd.n5010 gnd.t19 8.92286
R20433 gnd.n5086 gnd.n2063 8.92286
R20434 gnd.n5170 gnd.n5169 8.92286
R20435 gnd.n5235 gnd.n1980 8.92286
R20436 gnd.n5321 gnd.n5320 8.92286
R20437 gnd.n5371 gnd.n5370 8.92286
R20438 gnd.n5617 gnd.n1830 8.92286
R20439 gnd.n3996 gnd.n3971 8.92171
R20440 gnd.n3964 gnd.n3939 8.92171
R20441 gnd.n3932 gnd.n3907 8.92171
R20442 gnd.n3901 gnd.n3876 8.92171
R20443 gnd.n3869 gnd.n3844 8.92171
R20444 gnd.n3837 gnd.n3812 8.92171
R20445 gnd.n3805 gnd.n3780 8.92171
R20446 gnd.n3774 gnd.n3749 8.92171
R20447 gnd.n5473 gnd.n5455 8.72777
R20448 gnd.n3499 gnd.t351 8.60421
R20449 gnd.n2500 gnd.t200 8.60421
R20450 gnd.n5875 gnd.t247 8.60421
R20451 gnd.n191 gnd.n184 8.60421
R20452 gnd.n2911 gnd.n2895 8.43656
R20453 gnd.n50 gnd.n34 8.43656
R20454 gnd.n4941 gnd.t116 8.28555
R20455 gnd.t78 gnd.n5450 8.28555
R20456 gnd.n3997 gnd.n3969 8.14595
R20457 gnd.n3965 gnd.n3937 8.14595
R20458 gnd.n3933 gnd.n3905 8.14595
R20459 gnd.n3902 gnd.n3874 8.14595
R20460 gnd.n3870 gnd.n3842 8.14595
R20461 gnd.n3838 gnd.n3810 8.14595
R20462 gnd.n3806 gnd.n3778 8.14595
R20463 gnd.n3775 gnd.n3747 8.14595
R20464 gnd.n4594 gnd.n0 8.10675
R20465 gnd.n7629 gnd.n7628 8.10675
R20466 gnd.n4002 gnd.n4001 7.97301
R20467 gnd.t357 gnd.n3014 7.9669
R20468 gnd.n3740 gnd.n2738 7.9669
R20469 gnd.n4858 gnd.n4857 7.9669
R20470 gnd.n5727 gnd.n5726 7.9669
R20471 gnd.n7629 gnd.n82 7.86902
R20472 gnd.n6085 gnd.n1462 7.75808
R20473 gnd.n4796 gnd.n4795 7.75808
R20474 gnd.n7405 gnd.n349 7.75808
R20475 gnd.n4284 gnd.n4248 7.75808
R20476 gnd.n5056 gnd.n2081 7.64824
R20477 gnd.n5176 gnd.t5 7.64824
R20478 gnd.n5065 gnd.n2023 7.64824
R20479 gnd.n5230 gnd.n1993 7.64824
R20480 gnd.t140 gnd.n1977 7.64824
R20481 gnd.n5341 gnd.n5340 7.64824
R20482 gnd.t34 gnd.n5440 7.64824
R20483 gnd.n2944 gnd.n2943 7.53171
R20484 gnd.n3408 gnd.t347 7.32958
R20485 gnd.n4874 gnd.t59 7.32958
R20486 gnd.n2163 gnd.t358 7.32958
R20487 gnd.t368 gnd.n1795 7.32958
R20488 gnd.n5705 gnd.t26 7.32958
R20489 gnd.n1179 gnd.n1178 7.30353
R20490 gnd.n5472 gnd.n5471 7.30353
R20491 gnd.n3368 gnd.n3087 7.01093
R20492 gnd.n3090 gnd.n3088 7.01093
R20493 gnd.n3378 gnd.n3377 7.01093
R20494 gnd.n3389 gnd.n3071 7.01093
R20495 gnd.n3388 gnd.n3074 7.01093
R20496 gnd.n3399 gnd.n3062 7.01093
R20497 gnd.n3065 gnd.n3063 7.01093
R20498 gnd.n3409 gnd.n3408 7.01093
R20499 gnd.n3419 gnd.n3043 7.01093
R20500 gnd.n3418 gnd.n3046 7.01093
R20501 gnd.n3427 gnd.n3037 7.01093
R20502 gnd.n3439 gnd.n3027 7.01093
R20503 gnd.n3449 gnd.n3012 7.01093
R20504 gnd.n3465 gnd.n3464 7.01093
R20505 gnd.n3014 gnd.n2951 7.01093
R20506 gnd.n3519 gnd.n2952 7.01093
R20507 gnd.n3513 gnd.n3512 7.01093
R20508 gnd.n3001 gnd.n2963 7.01093
R20509 gnd.n3505 gnd.n2974 7.01093
R20510 gnd.n2992 gnd.n2987 7.01093
R20511 gnd.n3499 gnd.n3498 7.01093
R20512 gnd.n3545 gnd.n2874 7.01093
R20513 gnd.n3544 gnd.n3543 7.01093
R20514 gnd.n3556 gnd.n3555 7.01093
R20515 gnd.n2867 gnd.n2859 7.01093
R20516 gnd.n3585 gnd.n2847 7.01093
R20517 gnd.n3584 gnd.n2850 7.01093
R20518 gnd.n3595 gnd.n2839 7.01093
R20519 gnd.n2840 gnd.n2828 7.01093
R20520 gnd.n3606 gnd.n2829 7.01093
R20521 gnd.n3630 gnd.n2820 7.01093
R20522 gnd.n3629 gnd.n2811 7.01093
R20523 gnd.n3652 gnd.n3651 7.01093
R20524 gnd.n3670 gnd.n2792 7.01093
R20525 gnd.n3669 gnd.n2795 7.01093
R20526 gnd.n3680 gnd.n2784 7.01093
R20527 gnd.n2785 gnd.n2772 7.01093
R20528 gnd.n3691 gnd.n2773 7.01093
R20529 gnd.n3718 gnd.n2757 7.01093
R20530 gnd.n3730 gnd.n3729 7.01093
R20531 gnd.n3712 gnd.n2750 7.01093
R20532 gnd.n3742 gnd.n3741 7.01093
R20533 gnd.n4014 gnd.n2738 7.01093
R20534 gnd.n4013 gnd.n2741 7.01093
R20535 gnd.n4026 gnd.n2730 7.01093
R20536 gnd.n2731 gnd.n2723 7.01093
R20537 gnd.n4036 gnd.n2649 7.01093
R20538 gnd.n5062 gnd.t8 7.01093
R20539 gnd.t148 gnd.n1970 7.01093
R20540 gnd.n3046 gnd.t345 6.69227
R20541 gnd.n2850 gnd.t146 6.69227
R20542 gnd.n3719 gnd.t356 6.69227
R20543 gnd.n4491 gnd.t216 6.69227
R20544 gnd.n4691 gnd.t262 6.69227
R20545 gnd.t176 gnd.n2047 6.69227
R20546 gnd.n5243 gnd.t149 6.69227
R20547 gnd.n5758 gnd.t209 6.69227
R20548 gnd.n171 gnd.t207 6.69227
R20549 gnd.n5608 gnd.n5607 6.5566
R20550 gnd.n1208 gnd.n1207 6.5566
R20551 gnd.n6296 gnd.n6292 6.5566
R20552 gnd.n5483 gnd.n5482 6.5566
R20553 gnd.n1183 gnd.t16 6.37362
R20554 gnd.t30 gnd.t129 6.37362
R20555 gnd.n5051 gnd.n2091 6.37362
R20556 gnd.n2058 gnd.t2 6.37362
R20557 gnd.n5194 gnd.n2018 6.37362
R20558 gnd.n5200 gnd.n2008 6.37362
R20559 gnd.n5301 gnd.t139 6.37362
R20560 gnd.n1937 gnd.n1925 6.37362
R20561 gnd.n4785 gnd.n2455 6.20656
R20562 gnd.n1761 gnd.n1459 6.20656
R20563 gnd.t152 gnd.n3475 6.05496
R20564 gnd.n3476 gnd.t344 6.05496
R20565 gnd.t155 gnd.n2874 6.05496
R20566 gnd.t343 gnd.n3640 6.05496
R20567 gnd.n4545 gnd.t224 6.05496
R20568 gnd.n4672 gnd.t243 6.05496
R20569 gnd.t9 gnd.n2098 6.05496
R20570 gnd.t366 gnd.t145 6.05496
R20571 gnd.t137 gnd.t142 6.05496
R20572 gnd.n5359 gnd.t159 6.05496
R20573 gnd.n5844 gnd.t182 6.05496
R20574 gnd.n133 gnd.t184 6.05496
R20575 gnd.n3999 gnd.n3969 5.81868
R20576 gnd.n3967 gnd.n3937 5.81868
R20577 gnd.n3935 gnd.n3905 5.81868
R20578 gnd.n3904 gnd.n3874 5.81868
R20579 gnd.n3872 gnd.n3842 5.81868
R20580 gnd.n3840 gnd.n3810 5.81868
R20581 gnd.n3808 gnd.n3778 5.81868
R20582 gnd.n3777 gnd.n3747 5.81868
R20583 gnd.n5612 gnd.n1539 5.62001
R20584 gnd.n6358 gnd.n1121 5.62001
R20585 gnd.n6358 gnd.n1122 5.62001
R20586 gnd.n5478 gnd.n1539 5.62001
R20587 gnd.n3227 gnd.n3222 5.4308
R20588 gnd.n4044 gnd.n2716 5.4308
R20589 gnd.n3543 gnd.t342 5.41765
R20590 gnd.t350 gnd.n3566 5.41765
R20591 gnd.t364 gnd.n2804 5.41765
R20592 gnd.n6483 gnd.t260 5.41765
R20593 gnd.t211 gnd.n2516 5.41765
R20594 gnd.n7299 gnd.t220 5.41765
R20595 gnd.n7623 gnd.t194 5.41765
R20596 gnd.n6259 gnd.t131 5.09899
R20597 gnd.n2104 gnd.n2095 5.09899
R20598 gnd.n5207 gnd.n2012 5.09899
R20599 gnd.n5215 gnd.n2005 5.09899
R20600 gnd.n5365 gnd.n1921 5.09899
R20601 gnd.t138 gnd.n1911 5.09899
R20602 gnd.n3997 gnd.n3996 5.04292
R20603 gnd.n3965 gnd.n3964 5.04292
R20604 gnd.n3933 gnd.n3932 5.04292
R20605 gnd.n3902 gnd.n3901 5.04292
R20606 gnd.n3870 gnd.n3869 5.04292
R20607 gnd.n3838 gnd.n3837 5.04292
R20608 gnd.n3806 gnd.n3805 5.04292
R20609 gnd.n3775 gnd.n3774 5.04292
R20610 gnd.n3506 gnd.t353 4.78034
R20611 gnd.n2829 gnd.t354 4.78034
R20612 gnd.n4565 gnd.t188 4.78034
R20613 gnd.n6470 gnd.t200 4.78034
R20614 gnd.n4930 gnd.t167 4.78034
R20615 gnd.n5642 gnd.t6 4.78034
R20616 gnd.n5897 gnd.t247 4.78034
R20617 gnd.n7609 gnd.t218 4.78034
R20618 gnd.n2948 gnd.n2945 4.74817
R20619 gnd.n2998 gnd.n2880 4.74817
R20620 gnd.n2985 gnd.n2879 4.74817
R20621 gnd.n2878 gnd.n2877 4.74817
R20622 gnd.n2994 gnd.n2945 4.74817
R20623 gnd.n2995 gnd.n2880 4.74817
R20624 gnd.n2997 gnd.n2879 4.74817
R20625 gnd.n2984 gnd.n2878 4.74817
R20626 gnd.n5889 gnd.n101 4.74817
R20627 gnd.n386 gnd.n99 4.74817
R20628 gnd.n7621 gnd.n94 4.74817
R20629 gnd.n7619 gnd.n95 4.74817
R20630 gnd.n1695 gnd.n101 4.74817
R20631 gnd.n7297 gnd.n99 4.74817
R20632 gnd.n385 gnd.n94 4.74817
R20633 gnd.n7620 gnd.n7619 4.74817
R20634 gnd.n2539 gnd.n951 4.74817
R20635 gnd.n6480 gnd.n945 4.74817
R20636 gnd.n4616 gnd.n950 4.74817
R20637 gnd.n952 gnd.n949 4.74817
R20638 gnd.n4583 gnd.n951 4.74817
R20639 gnd.n6481 gnd.n6480 4.74817
R20640 gnd.n2519 gnd.n950 4.74817
R20641 gnd.n4617 gnd.n949 4.74817
R20642 gnd.n2943 gnd.n2942 4.74296
R20643 gnd.n82 gnd.n81 4.74296
R20644 gnd.n2911 gnd.n2910 4.7074
R20645 gnd.n2927 gnd.n2926 4.7074
R20646 gnd.n50 gnd.n49 4.7074
R20647 gnd.n66 gnd.n65 4.7074
R20648 gnd.n2943 gnd.n2927 4.65959
R20649 gnd.n82 gnd.n66 4.65959
R20650 gnd.n6027 gnd.n1541 4.6132
R20651 gnd.n6359 gnd.n1120 4.6132
R20652 gnd.n5114 gnd.t162 4.46168
R20653 gnd.t154 gnd.n1949 4.46168
R20654 gnd.n5371 gnd.t63 4.46168
R20655 gnd.n5468 gnd.n5455 4.46111
R20656 gnd.n3982 gnd.n3978 4.38594
R20657 gnd.n3950 gnd.n3946 4.38594
R20658 gnd.n3918 gnd.n3914 4.38594
R20659 gnd.n3887 gnd.n3883 4.38594
R20660 gnd.n3855 gnd.n3851 4.38594
R20661 gnd.n3823 gnd.n3819 4.38594
R20662 gnd.n3791 gnd.n3787 4.38594
R20663 gnd.n3760 gnd.n3756 4.38594
R20664 gnd.n3993 gnd.n3971 4.26717
R20665 gnd.n3961 gnd.n3939 4.26717
R20666 gnd.n3929 gnd.n3907 4.26717
R20667 gnd.n3898 gnd.n3876 4.26717
R20668 gnd.n3866 gnd.n3844 4.26717
R20669 gnd.n3834 gnd.n3812 4.26717
R20670 gnd.n3802 gnd.n3780 4.26717
R20671 gnd.n3771 gnd.n3749 4.26717
R20672 gnd.n3450 gnd.t355 4.14303
R20673 gnd.n3680 gnd.t352 4.14303
R20674 gnd.t190 gnd.n2580 4.14303
R20675 gnd.n6446 gnd.t276 4.14303
R20676 gnd.n2467 gnd.t55 4.14303
R20677 gnd.n5776 gnd.t12 4.14303
R20678 gnd.n5921 gnd.t222 4.14303
R20679 gnd.n7585 gnd.t265 4.14303
R20680 gnd.n4001 gnd.n4000 4.08274
R20681 gnd.n5607 gnd.n5606 4.05904
R20682 gnd.n1209 gnd.n1208 4.05904
R20683 gnd.n6299 gnd.n6292 4.05904
R20684 gnd.n5484 gnd.n5483 4.05904
R20685 gnd.n19 gnd.n9 3.99943
R20686 gnd.n5029 gnd.n2108 3.82437
R20687 gnd.n5045 gnd.t141 3.82437
R20688 gnd.n5095 gnd.n2078 3.82437
R20689 gnd.n5187 gnd.n2026 3.82437
R20690 gnd.n5224 gnd.n5223 3.82437
R20691 gnd.n5348 gnd.n5347 3.82437
R20692 gnd.t144 gnd.n1920 3.82437
R20693 gnd.n5404 gnd.n1907 3.82437
R20694 gnd.n3523 gnd.n2944 3.81325
R20695 gnd.n2927 gnd.n2911 3.72967
R20696 gnd.n66 gnd.n50 3.72967
R20697 gnd.n4001 gnd.n3873 3.70378
R20698 gnd.n19 gnd.n18 3.60163
R20699 gnd.n3992 gnd.n3973 3.49141
R20700 gnd.n3960 gnd.n3941 3.49141
R20701 gnd.n3928 gnd.n3909 3.49141
R20702 gnd.n3897 gnd.n3878 3.49141
R20703 gnd.n3865 gnd.n3846 3.49141
R20704 gnd.n3833 gnd.n3814 3.49141
R20705 gnd.n3801 gnd.n3782 3.49141
R20706 gnd.n3770 gnd.n3751 3.49141
R20707 gnd.n6045 gnd.n6044 3.29747
R20708 gnd.n6044 gnd.n6043 3.29747
R20709 gnd.n7514 gnd.n7511 3.29747
R20710 gnd.n7515 gnd.n7514 3.29747
R20711 gnd.n4406 gnd.n4405 3.29747
R20712 gnd.n4405 gnd.n4404 3.29747
R20713 gnd.n6375 gnd.n6374 3.29747
R20714 gnd.n6374 gnd.n6373 3.29747
R20715 gnd.t116 gnd.n1186 3.18706
R20716 gnd.n5028 gnd.t151 3.18706
R20717 gnd.n5036 gnd.t151 3.18706
R20718 gnd.n5279 gnd.t132 3.18706
R20719 gnd.n5392 gnd.t132 3.18706
R20720 gnd.n3029 gnd.t355 2.8684
R20721 gnd.n6355 gnd.n1125 2.8684
R20722 gnd.n6278 gnd.t135 2.8684
R20723 gnd.t165 gnd.n1877 2.8684
R20724 gnd.n5615 gnd.n1849 2.8684
R20725 gnd.n2928 gnd.t286 2.82907
R20726 gnd.n2928 gnd.t341 2.82907
R20727 gnd.n2930 gnd.t244 2.82907
R20728 gnd.n2930 gnd.t330 2.82907
R20729 gnd.n2932 gnd.t193 2.82907
R20730 gnd.n2932 gnd.t307 2.82907
R20731 gnd.n2934 gnd.t333 2.82907
R20732 gnd.n2934 gnd.t241 2.82907
R20733 gnd.n2936 gnd.t274 2.82907
R20734 gnd.n2936 gnd.t252 2.82907
R20735 gnd.n2938 gnd.t245 2.82907
R20736 gnd.n2938 gnd.t225 2.82907
R20737 gnd.n2940 gnd.t258 2.82907
R20738 gnd.n2940 gnd.t298 2.82907
R20739 gnd.n2881 gnd.t291 2.82907
R20740 gnd.n2881 gnd.t306 2.82907
R20741 gnd.n2883 gnd.t319 2.82907
R20742 gnd.n2883 gnd.t334 2.82907
R20743 gnd.n2885 gnd.t283 2.82907
R20744 gnd.n2885 gnd.t295 2.82907
R20745 gnd.n2887 gnd.t308 2.82907
R20746 gnd.n2887 gnd.t212 2.82907
R20747 gnd.n2889 gnd.t294 2.82907
R20748 gnd.n2889 gnd.t290 2.82907
R20749 gnd.n2891 gnd.t325 2.82907
R20750 gnd.n2891 gnd.t320 2.82907
R20751 gnd.n2893 gnd.t235 2.82907
R20752 gnd.n2893 gnd.t302 2.82907
R20753 gnd.n2896 gnd.t277 2.82907
R20754 gnd.n2896 gnd.t263 2.82907
R20755 gnd.n2898 gnd.t264 2.82907
R20756 gnd.n2898 gnd.t289 2.82907
R20757 gnd.n2900 gnd.t238 2.82907
R20758 gnd.n2900 gnd.t278 2.82907
R20759 gnd.n2902 gnd.t279 2.82907
R20760 gnd.n2902 gnd.t254 2.82907
R20761 gnd.n2904 gnd.t189 2.82907
R20762 gnd.n2904 gnd.t240 2.82907
R20763 gnd.n2906 gnd.t229 2.82907
R20764 gnd.n2906 gnd.t281 2.82907
R20765 gnd.n2908 gnd.t217 2.82907
R20766 gnd.n2908 gnd.t191 2.82907
R20767 gnd.n2912 gnd.t324 2.82907
R20768 gnd.n2912 gnd.t282 2.82907
R20769 gnd.n2914 gnd.t301 2.82907
R20770 gnd.n2914 gnd.t256 2.82907
R20771 gnd.n2916 gnd.t285 2.82907
R20772 gnd.n2916 gnd.t201 2.82907
R20773 gnd.n2918 gnd.t261 2.82907
R20774 gnd.n2918 gnd.t299 2.82907
R20775 gnd.n2920 gnd.t317 2.82907
R20776 gnd.n2920 gnd.t305 2.82907
R20777 gnd.n2922 gnd.t303 2.82907
R20778 gnd.n2922 gnd.t293 2.82907
R20779 gnd.n2924 gnd.t309 2.82907
R20780 gnd.n2924 gnd.t338 2.82907
R20781 gnd.n79 gnd.t266 2.82907
R20782 gnd.n79 gnd.t313 2.82907
R20783 gnd.n77 gnd.t312 2.82907
R20784 gnd.n77 gnd.t337 2.82907
R20785 gnd.n75 gnd.t339 2.82907
R20786 gnd.n75 gnd.t233 2.82907
R20787 gnd.n73 gnd.t335 2.82907
R20788 gnd.n73 gnd.t304 2.82907
R20789 gnd.n71 gnd.t284 2.82907
R20790 gnd.n71 gnd.t327 2.82907
R20791 gnd.n69 gnd.t300 2.82907
R20792 gnd.n69 gnd.t336 2.82907
R20793 gnd.n67 gnd.t316 2.82907
R20794 gnd.n67 gnd.t223 2.82907
R20795 gnd.n32 gnd.t328 2.82907
R20796 gnd.n32 gnd.t215 2.82907
R20797 gnd.n30 gnd.t185 2.82907
R20798 gnd.n30 gnd.t202 2.82907
R20799 gnd.n28 gnd.t314 2.82907
R20800 gnd.n28 gnd.t287 2.82907
R20801 gnd.n26 gnd.t273 2.82907
R20802 gnd.n26 gnd.t332 2.82907
R20803 gnd.n24 gnd.t323 2.82907
R20804 gnd.n24 gnd.t257 2.82907
R20805 gnd.n22 gnd.t234 2.82907
R20806 gnd.n22 gnd.t183 2.82907
R20807 gnd.n20 gnd.t331 2.82907
R20808 gnd.n20 gnd.t315 2.82907
R20809 gnd.n47 gnd.t329 2.82907
R20810 gnd.n47 gnd.t232 2.82907
R20811 gnd.n45 gnd.t249 2.82907
R20812 gnd.n45 gnd.t199 2.82907
R20813 gnd.n43 gnd.t204 2.82907
R20814 gnd.n43 gnd.t219 2.82907
R20815 gnd.n41 gnd.t221 2.82907
R20816 gnd.n41 gnd.t246 2.82907
R20817 gnd.n39 gnd.t248 2.82907
R20818 gnd.n39 gnd.t269 2.82907
R20819 gnd.n37 gnd.t267 2.82907
R20820 gnd.n37 gnd.t226 2.82907
R20821 gnd.n35 gnd.t227 2.82907
R20822 gnd.n35 gnd.t242 2.82907
R20823 gnd.n63 gnd.t311 2.82907
R20824 gnd.n63 gnd.t208 2.82907
R20825 gnd.n61 gnd.t253 2.82907
R20826 gnd.n61 gnd.t275 2.82907
R20827 gnd.n59 gnd.t280 2.82907
R20828 gnd.n59 gnd.t297 2.82907
R20829 gnd.n57 gnd.t270 2.82907
R20830 gnd.n57 gnd.t195 2.82907
R20831 gnd.n55 gnd.t321 2.82907
R20832 gnd.n55 gnd.t251 2.82907
R20833 gnd.n53 gnd.t187 2.82907
R20834 gnd.n53 gnd.t272 2.82907
R20835 gnd.n51 gnd.t210 2.82907
R20836 gnd.n51 gnd.t292 2.82907
R20837 gnd.n3989 gnd.n3988 2.71565
R20838 gnd.n3957 gnd.n3956 2.71565
R20839 gnd.n3925 gnd.n3924 2.71565
R20840 gnd.n3894 gnd.n3893 2.71565
R20841 gnd.n3862 gnd.n3861 2.71565
R20842 gnd.n3830 gnd.n3829 2.71565
R20843 gnd.n3798 gnd.n3797 2.71565
R20844 gnd.n3767 gnd.n3766 2.71565
R20845 gnd.t16 gnd.n1157 2.54975
R20846 gnd.n1277 gnd.t30 2.54975
R20847 gnd.n5011 gnd.n5010 2.54975
R20848 gnd.n5016 gnd.t131 2.54975
R20849 gnd.n5105 gnd.n2071 2.54975
R20850 gnd.n5105 gnd.t161 2.54975
R20851 gnd.n5177 gnd.n5176 2.54975
R20852 gnd.n5252 gnd.n1977 2.54975
R20853 gnd.n5270 gnd.t4 2.54975
R20854 gnd.n5270 gnd.n1941 2.54975
R20855 gnd.n5385 gnd.t138 2.54975
R20856 gnd.n5414 gnd.n1899 2.54975
R20857 gnd.n5442 gnd.t34 2.54975
R20858 gnd.n5440 gnd.t41 2.54975
R20859 gnd.n3523 gnd.n2945 2.27742
R20860 gnd.n3523 gnd.n2880 2.27742
R20861 gnd.n3523 gnd.n2879 2.27742
R20862 gnd.n3523 gnd.n2878 2.27742
R20863 gnd.n7618 gnd.n101 2.27742
R20864 gnd.n7618 gnd.n99 2.27742
R20865 gnd.n7618 gnd.n94 2.27742
R20866 gnd.n7619 gnd.n7618 2.27742
R20867 gnd.n6479 gnd.n951 2.27742
R20868 gnd.n6480 gnd.n6479 2.27742
R20869 gnd.n6479 gnd.n950 2.27742
R20870 gnd.n6479 gnd.n949 2.27742
R20871 gnd.n3377 gnd.t48 2.23109
R20872 gnd.n3000 gnd.t353 2.23109
R20873 gnd.n4648 gnd.t192 2.23109
R20874 gnd.n2026 gnd.t366 2.23109
R20875 gnd.n5224 gnd.t142 2.23109
R20876 gnd.n1696 gnd.t250 2.23109
R20877 gnd.n3985 gnd.n3975 1.93989
R20878 gnd.n3953 gnd.n3943 1.93989
R20879 gnd.n3921 gnd.n3911 1.93989
R20880 gnd.n3890 gnd.n3880 1.93989
R20881 gnd.n3858 gnd.n3848 1.93989
R20882 gnd.n3826 gnd.n3816 1.93989
R20883 gnd.n3794 gnd.n3784 1.93989
R20884 gnd.n3763 gnd.n3753 1.93989
R20885 gnd.n5451 gnd.t78 1.91244
R20886 gnd.n1849 gnd.t91 1.91244
R20887 gnd.t157 gnd.n3388 1.59378
R20888 gnd.n3567 gnd.t350 1.59378
R20889 gnd.n2813 gnd.t364 1.59378
R20890 gnd.n4709 gnd.t255 1.59378
R20891 gnd.n5016 gnd.t169 1.59378
R20892 gnd.t360 gnd.n5086 1.59378
R20893 gnd.n5320 gnd.t174 1.59378
R20894 gnd.n5385 gnd.t370 1.59378
R20895 gnd.n1715 gnd.t186 1.59378
R20896 gnd.n6285 gnd.n6284 1.27512
R20897 gnd.n1286 gnd.n1276 1.27512
R20898 gnd.t141 gnd.n5044 1.27512
R20899 gnd.n5115 gnd.n5114 1.27512
R20900 gnd.n5062 gnd.n5061 1.27512
R20901 gnd.n5262 gnd.n1970 1.27512
R20902 gnd.n5322 gnd.n1949 1.27512
R20903 gnd.n5358 gnd.t144 1.27512
R20904 gnd.n5434 gnd.n5433 1.27512
R20905 gnd.n5546 gnd.n1872 1.27512
R20906 gnd.n3230 gnd.n3222 1.16414
R20907 gnd.n4047 gnd.n2716 1.16414
R20908 gnd.n3984 gnd.n3977 1.16414
R20909 gnd.n3952 gnd.n3945 1.16414
R20910 gnd.n3920 gnd.n3913 1.16414
R20911 gnd.n3889 gnd.n3882 1.16414
R20912 gnd.n3857 gnd.n3850 1.16414
R20913 gnd.n3825 gnd.n3818 1.16414
R20914 gnd.n3793 gnd.n3786 1.16414
R20915 gnd.n3762 gnd.n3755 1.16414
R20916 gnd.n6027 gnd.n6026 0.970197
R20917 gnd.n6359 gnd.n1117 0.970197
R20918 gnd.n3968 gnd.n3936 0.962709
R20919 gnd.n4000 gnd.n3968 0.962709
R20920 gnd.n3841 gnd.n3809 0.962709
R20921 gnd.n3873 gnd.n3841 0.962709
R20922 gnd.n3476 gnd.t152 0.956468
R20923 gnd.n3641 gnd.t343 0.956468
R20924 gnd.n4755 gnd.t196 0.956468
R20925 gnd.n5748 gnd.t205 0.956468
R20926 gnd.n2 gnd.n1 0.672012
R20927 gnd.n3 gnd.n2 0.672012
R20928 gnd.n4 gnd.n3 0.672012
R20929 gnd.n5 gnd.n4 0.672012
R20930 gnd.n6 gnd.n5 0.672012
R20931 gnd.n7 gnd.n6 0.672012
R20932 gnd.n8 gnd.n7 0.672012
R20933 gnd.n9 gnd.n8 0.672012
R20934 gnd.n11 gnd.n10 0.672012
R20935 gnd.n12 gnd.n11 0.672012
R20936 gnd.n13 gnd.n12 0.672012
R20937 gnd.n14 gnd.n13 0.672012
R20938 gnd.n15 gnd.n14 0.672012
R20939 gnd.n16 gnd.n15 0.672012
R20940 gnd.n17 gnd.n16 0.672012
R20941 gnd.n18 gnd.n17 0.672012
R20942 gnd gnd.n0 0.665707
R20943 gnd.t66 gnd.n1286 0.637812
R20944 gnd.n5095 gnd.t173 0.637812
R20945 gnd.n5348 gnd.t3 0.637812
R20946 gnd.n2942 gnd.n2941 0.573776
R20947 gnd.n2941 gnd.n2939 0.573776
R20948 gnd.n2939 gnd.n2937 0.573776
R20949 gnd.n2937 gnd.n2935 0.573776
R20950 gnd.n2935 gnd.n2933 0.573776
R20951 gnd.n2933 gnd.n2931 0.573776
R20952 gnd.n2931 gnd.n2929 0.573776
R20953 gnd.n2895 gnd.n2894 0.573776
R20954 gnd.n2894 gnd.n2892 0.573776
R20955 gnd.n2892 gnd.n2890 0.573776
R20956 gnd.n2890 gnd.n2888 0.573776
R20957 gnd.n2888 gnd.n2886 0.573776
R20958 gnd.n2886 gnd.n2884 0.573776
R20959 gnd.n2884 gnd.n2882 0.573776
R20960 gnd.n2910 gnd.n2909 0.573776
R20961 gnd.n2909 gnd.n2907 0.573776
R20962 gnd.n2907 gnd.n2905 0.573776
R20963 gnd.n2905 gnd.n2903 0.573776
R20964 gnd.n2903 gnd.n2901 0.573776
R20965 gnd.n2901 gnd.n2899 0.573776
R20966 gnd.n2899 gnd.n2897 0.573776
R20967 gnd.n2926 gnd.n2925 0.573776
R20968 gnd.n2925 gnd.n2923 0.573776
R20969 gnd.n2923 gnd.n2921 0.573776
R20970 gnd.n2921 gnd.n2919 0.573776
R20971 gnd.n2919 gnd.n2917 0.573776
R20972 gnd.n2917 gnd.n2915 0.573776
R20973 gnd.n2915 gnd.n2913 0.573776
R20974 gnd.n70 gnd.n68 0.573776
R20975 gnd.n72 gnd.n70 0.573776
R20976 gnd.n74 gnd.n72 0.573776
R20977 gnd.n76 gnd.n74 0.573776
R20978 gnd.n78 gnd.n76 0.573776
R20979 gnd.n80 gnd.n78 0.573776
R20980 gnd.n81 gnd.n80 0.573776
R20981 gnd.n23 gnd.n21 0.573776
R20982 gnd.n25 gnd.n23 0.573776
R20983 gnd.n27 gnd.n25 0.573776
R20984 gnd.n29 gnd.n27 0.573776
R20985 gnd.n31 gnd.n29 0.573776
R20986 gnd.n33 gnd.n31 0.573776
R20987 gnd.n34 gnd.n33 0.573776
R20988 gnd.n38 gnd.n36 0.573776
R20989 gnd.n40 gnd.n38 0.573776
R20990 gnd.n42 gnd.n40 0.573776
R20991 gnd.n44 gnd.n42 0.573776
R20992 gnd.n46 gnd.n44 0.573776
R20993 gnd.n48 gnd.n46 0.573776
R20994 gnd.n49 gnd.n48 0.573776
R20995 gnd.n54 gnd.n52 0.573776
R20996 gnd.n56 gnd.n54 0.573776
R20997 gnd.n58 gnd.n56 0.573776
R20998 gnd.n60 gnd.n58 0.573776
R20999 gnd.n62 gnd.n60 0.573776
R21000 gnd.n64 gnd.n62 0.573776
R21001 gnd.n65 gnd.n64 0.573776
R21002 gnd.n7630 gnd.n7629 0.553847
R21003 gnd.n7403 gnd.n7402 0.505073
R21004 gnd.n4285 gnd.n4283 0.505073
R21005 gnd.n3703 gnd.n2720 0.486781
R21006 gnd.n3279 gnd.n3278 0.48678
R21007 gnd.n4021 gnd.n2674 0.480683
R21008 gnd.n3363 gnd.n3362 0.480683
R21009 gnd.n6656 gnd.n6655 0.480683
R21010 gnd.n7076 gnd.n7075 0.480683
R21011 gnd.n7289 gnd.n7288 0.480683
R21012 gnd.n2512 gnd.n936 0.480683
R21013 gnd.n7546 gnd.n7545 0.470012
R21014 gnd.n1592 gnd.n1511 0.470012
R21015 gnd.n6407 gnd.n6406 0.470012
R21016 gnd.n4167 gnd.n2633 0.470012
R21017 gnd.n1737 gnd.n1393 0.451719
R21018 gnd.n4869 gnd.n2193 0.451719
R21019 gnd.n2270 gnd.n2269 0.451719
R21020 gnd.n6145 gnd.n6144 0.451719
R21021 gnd.n7618 gnd.n98 0.420375
R21022 gnd.n6479 gnd.n948 0.420375
R21023 gnd.n4800 gnd.n2455 0.388379
R21024 gnd.n3981 gnd.n3980 0.388379
R21025 gnd.n3949 gnd.n3948 0.388379
R21026 gnd.n3917 gnd.n3916 0.388379
R21027 gnd.n3886 gnd.n3885 0.388379
R21028 gnd.n3854 gnd.n3853 0.388379
R21029 gnd.n3822 gnd.n3821 0.388379
R21030 gnd.n3790 gnd.n3789 0.388379
R21031 gnd.n3759 gnd.n3758 0.388379
R21032 gnd.n6089 gnd.n1459 0.388379
R21033 gnd.n7630 gnd.n19 0.374463
R21034 gnd gnd.n7630 0.367492
R21035 gnd.n2775 gnd.t356 0.319156
R21036 gnd.n3197 gnd.n3175 0.311721
R21037 gnd.n7436 gnd.n7435 0.293183
R21038 gnd.n4323 gnd.n4322 0.293183
R21039 gnd.n4783 gnd.n4782 0.27489
R21040 gnd.n5734 gnd.n5733 0.27489
R21041 gnd.n4092 gnd.n4091 0.268793
R21042 gnd.n7437 gnd.n7436 0.258122
R21043 gnd.n5965 gnd.n1412 0.258122
R21044 gnd.n2389 gnd.n2388 0.258122
R21045 gnd.n4324 gnd.n4323 0.258122
R21046 gnd.n4091 gnd.n4090 0.241354
R21047 gnd.n1541 gnd.n1538 0.229039
R21048 gnd.n1542 gnd.n1541 0.229039
R21049 gnd.n1120 gnd.n1116 0.229039
R21050 gnd.n2309 gnd.n1120 0.229039
R21051 gnd.n3351 gnd.n3150 0.206293
R21052 gnd.n2944 gnd.n0 0.169152
R21053 gnd.n3998 gnd.n3970 0.155672
R21054 gnd.n3991 gnd.n3970 0.155672
R21055 gnd.n3991 gnd.n3990 0.155672
R21056 gnd.n3990 gnd.n3974 0.155672
R21057 gnd.n3983 gnd.n3974 0.155672
R21058 gnd.n3983 gnd.n3982 0.155672
R21059 gnd.n3966 gnd.n3938 0.155672
R21060 gnd.n3959 gnd.n3938 0.155672
R21061 gnd.n3959 gnd.n3958 0.155672
R21062 gnd.n3958 gnd.n3942 0.155672
R21063 gnd.n3951 gnd.n3942 0.155672
R21064 gnd.n3951 gnd.n3950 0.155672
R21065 gnd.n3934 gnd.n3906 0.155672
R21066 gnd.n3927 gnd.n3906 0.155672
R21067 gnd.n3927 gnd.n3926 0.155672
R21068 gnd.n3926 gnd.n3910 0.155672
R21069 gnd.n3919 gnd.n3910 0.155672
R21070 gnd.n3919 gnd.n3918 0.155672
R21071 gnd.n3903 gnd.n3875 0.155672
R21072 gnd.n3896 gnd.n3875 0.155672
R21073 gnd.n3896 gnd.n3895 0.155672
R21074 gnd.n3895 gnd.n3879 0.155672
R21075 gnd.n3888 gnd.n3879 0.155672
R21076 gnd.n3888 gnd.n3887 0.155672
R21077 gnd.n3871 gnd.n3843 0.155672
R21078 gnd.n3864 gnd.n3843 0.155672
R21079 gnd.n3864 gnd.n3863 0.155672
R21080 gnd.n3863 gnd.n3847 0.155672
R21081 gnd.n3856 gnd.n3847 0.155672
R21082 gnd.n3856 gnd.n3855 0.155672
R21083 gnd.n3839 gnd.n3811 0.155672
R21084 gnd.n3832 gnd.n3811 0.155672
R21085 gnd.n3832 gnd.n3831 0.155672
R21086 gnd.n3831 gnd.n3815 0.155672
R21087 gnd.n3824 gnd.n3815 0.155672
R21088 gnd.n3824 gnd.n3823 0.155672
R21089 gnd.n3807 gnd.n3779 0.155672
R21090 gnd.n3800 gnd.n3779 0.155672
R21091 gnd.n3800 gnd.n3799 0.155672
R21092 gnd.n3799 gnd.n3783 0.155672
R21093 gnd.n3792 gnd.n3783 0.155672
R21094 gnd.n3792 gnd.n3791 0.155672
R21095 gnd.n3776 gnd.n3748 0.155672
R21096 gnd.n3769 gnd.n3748 0.155672
R21097 gnd.n3769 gnd.n3768 0.155672
R21098 gnd.n3768 gnd.n3752 0.155672
R21099 gnd.n3761 gnd.n3752 0.155672
R21100 gnd.n3761 gnd.n3760 0.155672
R21101 gnd.n4123 gnd.n2674 0.152939
R21102 gnd.n4123 gnd.n4122 0.152939
R21103 gnd.n4122 gnd.n4121 0.152939
R21104 gnd.n4121 gnd.n2676 0.152939
R21105 gnd.n2677 gnd.n2676 0.152939
R21106 gnd.n2678 gnd.n2677 0.152939
R21107 gnd.n2679 gnd.n2678 0.152939
R21108 gnd.n2680 gnd.n2679 0.152939
R21109 gnd.n2681 gnd.n2680 0.152939
R21110 gnd.n2682 gnd.n2681 0.152939
R21111 gnd.n2683 gnd.n2682 0.152939
R21112 gnd.n2684 gnd.n2683 0.152939
R21113 gnd.n2685 gnd.n2684 0.152939
R21114 gnd.n2686 gnd.n2685 0.152939
R21115 gnd.n4093 gnd.n2686 0.152939
R21116 gnd.n4093 gnd.n4092 0.152939
R21117 gnd.n3364 gnd.n3363 0.152939
R21118 gnd.n3364 gnd.n3068 0.152939
R21119 gnd.n3392 gnd.n3068 0.152939
R21120 gnd.n3393 gnd.n3392 0.152939
R21121 gnd.n3394 gnd.n3393 0.152939
R21122 gnd.n3395 gnd.n3394 0.152939
R21123 gnd.n3395 gnd.n3040 0.152939
R21124 gnd.n3422 gnd.n3040 0.152939
R21125 gnd.n3423 gnd.n3422 0.152939
R21126 gnd.n3424 gnd.n3423 0.152939
R21127 gnd.n3424 gnd.n3018 0.152939
R21128 gnd.n3453 gnd.n3018 0.152939
R21129 gnd.n3454 gnd.n3453 0.152939
R21130 gnd.n3455 gnd.n3454 0.152939
R21131 gnd.n3456 gnd.n3455 0.152939
R21132 gnd.n3458 gnd.n3456 0.152939
R21133 gnd.n3458 gnd.n3457 0.152939
R21134 gnd.n3457 gnd.n2967 0.152939
R21135 gnd.n2968 gnd.n2967 0.152939
R21136 gnd.n2969 gnd.n2968 0.152939
R21137 gnd.n2988 gnd.n2969 0.152939
R21138 gnd.n2989 gnd.n2988 0.152939
R21139 gnd.n2989 gnd.n2871 0.152939
R21140 gnd.n3548 gnd.n2871 0.152939
R21141 gnd.n3549 gnd.n3548 0.152939
R21142 gnd.n3550 gnd.n3549 0.152939
R21143 gnd.n3551 gnd.n3550 0.152939
R21144 gnd.n3551 gnd.n2844 0.152939
R21145 gnd.n3588 gnd.n2844 0.152939
R21146 gnd.n3589 gnd.n3588 0.152939
R21147 gnd.n3590 gnd.n3589 0.152939
R21148 gnd.n3591 gnd.n3590 0.152939
R21149 gnd.n3591 gnd.n2817 0.152939
R21150 gnd.n3633 gnd.n2817 0.152939
R21151 gnd.n3634 gnd.n3633 0.152939
R21152 gnd.n3635 gnd.n3634 0.152939
R21153 gnd.n3636 gnd.n3635 0.152939
R21154 gnd.n3636 gnd.n2789 0.152939
R21155 gnd.n3673 gnd.n2789 0.152939
R21156 gnd.n3674 gnd.n3673 0.152939
R21157 gnd.n3675 gnd.n3674 0.152939
R21158 gnd.n3676 gnd.n3675 0.152939
R21159 gnd.n3676 gnd.n2762 0.152939
R21160 gnd.n3722 gnd.n2762 0.152939
R21161 gnd.n3723 gnd.n3722 0.152939
R21162 gnd.n3724 gnd.n3723 0.152939
R21163 gnd.n3725 gnd.n3724 0.152939
R21164 gnd.n3725 gnd.n2735 0.152939
R21165 gnd.n4017 gnd.n2735 0.152939
R21166 gnd.n4018 gnd.n4017 0.152939
R21167 gnd.n4019 gnd.n4018 0.152939
R21168 gnd.n4020 gnd.n4019 0.152939
R21169 gnd.n4021 gnd.n4020 0.152939
R21170 gnd.n3362 gnd.n3092 0.152939
R21171 gnd.n3113 gnd.n3092 0.152939
R21172 gnd.n3114 gnd.n3113 0.152939
R21173 gnd.n3120 gnd.n3114 0.152939
R21174 gnd.n3121 gnd.n3120 0.152939
R21175 gnd.n3122 gnd.n3121 0.152939
R21176 gnd.n3122 gnd.n3111 0.152939
R21177 gnd.n3130 gnd.n3111 0.152939
R21178 gnd.n3131 gnd.n3130 0.152939
R21179 gnd.n3132 gnd.n3131 0.152939
R21180 gnd.n3132 gnd.n3109 0.152939
R21181 gnd.n3140 gnd.n3109 0.152939
R21182 gnd.n3141 gnd.n3140 0.152939
R21183 gnd.n3142 gnd.n3141 0.152939
R21184 gnd.n3142 gnd.n3107 0.152939
R21185 gnd.n3150 gnd.n3107 0.152939
R21186 gnd.n4090 gnd.n2691 0.152939
R21187 gnd.n2693 gnd.n2691 0.152939
R21188 gnd.n2694 gnd.n2693 0.152939
R21189 gnd.n2695 gnd.n2694 0.152939
R21190 gnd.n2696 gnd.n2695 0.152939
R21191 gnd.n2697 gnd.n2696 0.152939
R21192 gnd.n2698 gnd.n2697 0.152939
R21193 gnd.n2699 gnd.n2698 0.152939
R21194 gnd.n2700 gnd.n2699 0.152939
R21195 gnd.n2701 gnd.n2700 0.152939
R21196 gnd.n2702 gnd.n2701 0.152939
R21197 gnd.n2703 gnd.n2702 0.152939
R21198 gnd.n2704 gnd.n2703 0.152939
R21199 gnd.n2705 gnd.n2704 0.152939
R21200 gnd.n2706 gnd.n2705 0.152939
R21201 gnd.n2707 gnd.n2706 0.152939
R21202 gnd.n2708 gnd.n2707 0.152939
R21203 gnd.n2709 gnd.n2708 0.152939
R21204 gnd.n2710 gnd.n2709 0.152939
R21205 gnd.n2711 gnd.n2710 0.152939
R21206 gnd.n2712 gnd.n2711 0.152939
R21207 gnd.n2713 gnd.n2712 0.152939
R21208 gnd.n2717 gnd.n2713 0.152939
R21209 gnd.n2718 gnd.n2717 0.152939
R21210 gnd.n2719 gnd.n2718 0.152939
R21211 gnd.n2720 gnd.n2719 0.152939
R21212 gnd.n3525 gnd.n3524 0.152939
R21213 gnd.n3526 gnd.n3525 0.152939
R21214 gnd.n3527 gnd.n3526 0.152939
R21215 gnd.n3528 gnd.n3527 0.152939
R21216 gnd.n3529 gnd.n3528 0.152939
R21217 gnd.n3530 gnd.n3529 0.152939
R21218 gnd.n3530 gnd.n2825 0.152939
R21219 gnd.n3609 gnd.n2825 0.152939
R21220 gnd.n3610 gnd.n3609 0.152939
R21221 gnd.n3611 gnd.n3610 0.152939
R21222 gnd.n3612 gnd.n3611 0.152939
R21223 gnd.n3613 gnd.n3612 0.152939
R21224 gnd.n3614 gnd.n3613 0.152939
R21225 gnd.n3615 gnd.n3614 0.152939
R21226 gnd.n3616 gnd.n3615 0.152939
R21227 gnd.n3617 gnd.n3616 0.152939
R21228 gnd.n3617 gnd.n2769 0.152939
R21229 gnd.n3694 gnd.n2769 0.152939
R21230 gnd.n3695 gnd.n3694 0.152939
R21231 gnd.n3696 gnd.n3695 0.152939
R21232 gnd.n3697 gnd.n3696 0.152939
R21233 gnd.n3698 gnd.n3697 0.152939
R21234 gnd.n3699 gnd.n3698 0.152939
R21235 gnd.n3700 gnd.n3699 0.152939
R21236 gnd.n3701 gnd.n3700 0.152939
R21237 gnd.n3702 gnd.n3701 0.152939
R21238 gnd.n3704 gnd.n3702 0.152939
R21239 gnd.n3704 gnd.n3703 0.152939
R21240 gnd.n3280 gnd.n3279 0.152939
R21241 gnd.n3280 gnd.n3170 0.152939
R21242 gnd.n3295 gnd.n3170 0.152939
R21243 gnd.n3296 gnd.n3295 0.152939
R21244 gnd.n3297 gnd.n3296 0.152939
R21245 gnd.n3297 gnd.n3158 0.152939
R21246 gnd.n3311 gnd.n3158 0.152939
R21247 gnd.n3312 gnd.n3311 0.152939
R21248 gnd.n3313 gnd.n3312 0.152939
R21249 gnd.n3314 gnd.n3313 0.152939
R21250 gnd.n3315 gnd.n3314 0.152939
R21251 gnd.n3316 gnd.n3315 0.152939
R21252 gnd.n3317 gnd.n3316 0.152939
R21253 gnd.n3318 gnd.n3317 0.152939
R21254 gnd.n3319 gnd.n3318 0.152939
R21255 gnd.n3320 gnd.n3319 0.152939
R21256 gnd.n3321 gnd.n3320 0.152939
R21257 gnd.n3322 gnd.n3321 0.152939
R21258 gnd.n3323 gnd.n3322 0.152939
R21259 gnd.n3324 gnd.n3323 0.152939
R21260 gnd.n3325 gnd.n3324 0.152939
R21261 gnd.n3325 gnd.n3024 0.152939
R21262 gnd.n3442 gnd.n3024 0.152939
R21263 gnd.n3443 gnd.n3442 0.152939
R21264 gnd.n3444 gnd.n3443 0.152939
R21265 gnd.n3445 gnd.n3444 0.152939
R21266 gnd.n3445 gnd.n2946 0.152939
R21267 gnd.n3522 gnd.n2946 0.152939
R21268 gnd.n3198 gnd.n3197 0.152939
R21269 gnd.n3199 gnd.n3198 0.152939
R21270 gnd.n3200 gnd.n3199 0.152939
R21271 gnd.n3201 gnd.n3200 0.152939
R21272 gnd.n3202 gnd.n3201 0.152939
R21273 gnd.n3203 gnd.n3202 0.152939
R21274 gnd.n3204 gnd.n3203 0.152939
R21275 gnd.n3205 gnd.n3204 0.152939
R21276 gnd.n3206 gnd.n3205 0.152939
R21277 gnd.n3207 gnd.n3206 0.152939
R21278 gnd.n3208 gnd.n3207 0.152939
R21279 gnd.n3209 gnd.n3208 0.152939
R21280 gnd.n3210 gnd.n3209 0.152939
R21281 gnd.n3211 gnd.n3210 0.152939
R21282 gnd.n3212 gnd.n3211 0.152939
R21283 gnd.n3213 gnd.n3212 0.152939
R21284 gnd.n3214 gnd.n3213 0.152939
R21285 gnd.n3215 gnd.n3214 0.152939
R21286 gnd.n3216 gnd.n3215 0.152939
R21287 gnd.n3217 gnd.n3216 0.152939
R21288 gnd.n3218 gnd.n3217 0.152939
R21289 gnd.n3219 gnd.n3218 0.152939
R21290 gnd.n3223 gnd.n3219 0.152939
R21291 gnd.n3224 gnd.n3223 0.152939
R21292 gnd.n3224 gnd.n3181 0.152939
R21293 gnd.n3278 gnd.n3181 0.152939
R21294 gnd.n6657 gnd.n6656 0.152939
R21295 gnd.n6657 gnd.n763 0.152939
R21296 gnd.n6665 gnd.n763 0.152939
R21297 gnd.n6666 gnd.n6665 0.152939
R21298 gnd.n6667 gnd.n6666 0.152939
R21299 gnd.n6667 gnd.n757 0.152939
R21300 gnd.n6675 gnd.n757 0.152939
R21301 gnd.n6676 gnd.n6675 0.152939
R21302 gnd.n6677 gnd.n6676 0.152939
R21303 gnd.n6677 gnd.n751 0.152939
R21304 gnd.n6685 gnd.n751 0.152939
R21305 gnd.n6686 gnd.n6685 0.152939
R21306 gnd.n6687 gnd.n6686 0.152939
R21307 gnd.n6687 gnd.n745 0.152939
R21308 gnd.n6695 gnd.n745 0.152939
R21309 gnd.n6696 gnd.n6695 0.152939
R21310 gnd.n6697 gnd.n6696 0.152939
R21311 gnd.n6697 gnd.n739 0.152939
R21312 gnd.n6705 gnd.n739 0.152939
R21313 gnd.n6706 gnd.n6705 0.152939
R21314 gnd.n6707 gnd.n6706 0.152939
R21315 gnd.n6707 gnd.n733 0.152939
R21316 gnd.n6715 gnd.n733 0.152939
R21317 gnd.n6716 gnd.n6715 0.152939
R21318 gnd.n6717 gnd.n6716 0.152939
R21319 gnd.n6717 gnd.n727 0.152939
R21320 gnd.n6725 gnd.n727 0.152939
R21321 gnd.n6726 gnd.n6725 0.152939
R21322 gnd.n6727 gnd.n6726 0.152939
R21323 gnd.n6727 gnd.n721 0.152939
R21324 gnd.n6735 gnd.n721 0.152939
R21325 gnd.n6736 gnd.n6735 0.152939
R21326 gnd.n6737 gnd.n6736 0.152939
R21327 gnd.n6737 gnd.n715 0.152939
R21328 gnd.n6745 gnd.n715 0.152939
R21329 gnd.n6746 gnd.n6745 0.152939
R21330 gnd.n6747 gnd.n6746 0.152939
R21331 gnd.n6747 gnd.n709 0.152939
R21332 gnd.n6755 gnd.n709 0.152939
R21333 gnd.n6756 gnd.n6755 0.152939
R21334 gnd.n6757 gnd.n6756 0.152939
R21335 gnd.n6757 gnd.n703 0.152939
R21336 gnd.n6765 gnd.n703 0.152939
R21337 gnd.n6766 gnd.n6765 0.152939
R21338 gnd.n6767 gnd.n6766 0.152939
R21339 gnd.n6767 gnd.n697 0.152939
R21340 gnd.n6775 gnd.n697 0.152939
R21341 gnd.n6776 gnd.n6775 0.152939
R21342 gnd.n6777 gnd.n6776 0.152939
R21343 gnd.n6777 gnd.n691 0.152939
R21344 gnd.n6785 gnd.n691 0.152939
R21345 gnd.n6786 gnd.n6785 0.152939
R21346 gnd.n6787 gnd.n6786 0.152939
R21347 gnd.n6787 gnd.n685 0.152939
R21348 gnd.n6795 gnd.n685 0.152939
R21349 gnd.n6796 gnd.n6795 0.152939
R21350 gnd.n6797 gnd.n6796 0.152939
R21351 gnd.n6797 gnd.n679 0.152939
R21352 gnd.n6805 gnd.n679 0.152939
R21353 gnd.n6806 gnd.n6805 0.152939
R21354 gnd.n6807 gnd.n6806 0.152939
R21355 gnd.n6807 gnd.n673 0.152939
R21356 gnd.n6815 gnd.n673 0.152939
R21357 gnd.n6816 gnd.n6815 0.152939
R21358 gnd.n6817 gnd.n6816 0.152939
R21359 gnd.n6817 gnd.n667 0.152939
R21360 gnd.n6825 gnd.n667 0.152939
R21361 gnd.n6826 gnd.n6825 0.152939
R21362 gnd.n6827 gnd.n6826 0.152939
R21363 gnd.n6827 gnd.n661 0.152939
R21364 gnd.n6835 gnd.n661 0.152939
R21365 gnd.n6836 gnd.n6835 0.152939
R21366 gnd.n6837 gnd.n6836 0.152939
R21367 gnd.n6837 gnd.n655 0.152939
R21368 gnd.n6845 gnd.n655 0.152939
R21369 gnd.n6846 gnd.n6845 0.152939
R21370 gnd.n6847 gnd.n6846 0.152939
R21371 gnd.n6847 gnd.n649 0.152939
R21372 gnd.n6855 gnd.n649 0.152939
R21373 gnd.n6856 gnd.n6855 0.152939
R21374 gnd.n6857 gnd.n6856 0.152939
R21375 gnd.n6857 gnd.n643 0.152939
R21376 gnd.n6865 gnd.n643 0.152939
R21377 gnd.n6866 gnd.n6865 0.152939
R21378 gnd.n6867 gnd.n6866 0.152939
R21379 gnd.n6867 gnd.n637 0.152939
R21380 gnd.n6875 gnd.n637 0.152939
R21381 gnd.n6876 gnd.n6875 0.152939
R21382 gnd.n6877 gnd.n6876 0.152939
R21383 gnd.n6877 gnd.n631 0.152939
R21384 gnd.n6885 gnd.n631 0.152939
R21385 gnd.n6886 gnd.n6885 0.152939
R21386 gnd.n6887 gnd.n6886 0.152939
R21387 gnd.n6887 gnd.n625 0.152939
R21388 gnd.n6895 gnd.n625 0.152939
R21389 gnd.n6896 gnd.n6895 0.152939
R21390 gnd.n6897 gnd.n6896 0.152939
R21391 gnd.n6897 gnd.n619 0.152939
R21392 gnd.n6905 gnd.n619 0.152939
R21393 gnd.n6906 gnd.n6905 0.152939
R21394 gnd.n6907 gnd.n6906 0.152939
R21395 gnd.n6907 gnd.n613 0.152939
R21396 gnd.n6915 gnd.n613 0.152939
R21397 gnd.n6916 gnd.n6915 0.152939
R21398 gnd.n6917 gnd.n6916 0.152939
R21399 gnd.n6917 gnd.n607 0.152939
R21400 gnd.n6925 gnd.n607 0.152939
R21401 gnd.n6926 gnd.n6925 0.152939
R21402 gnd.n6927 gnd.n6926 0.152939
R21403 gnd.n6927 gnd.n601 0.152939
R21404 gnd.n6935 gnd.n601 0.152939
R21405 gnd.n6936 gnd.n6935 0.152939
R21406 gnd.n6937 gnd.n6936 0.152939
R21407 gnd.n6937 gnd.n595 0.152939
R21408 gnd.n6945 gnd.n595 0.152939
R21409 gnd.n6946 gnd.n6945 0.152939
R21410 gnd.n6947 gnd.n6946 0.152939
R21411 gnd.n6947 gnd.n589 0.152939
R21412 gnd.n6955 gnd.n589 0.152939
R21413 gnd.n6956 gnd.n6955 0.152939
R21414 gnd.n6957 gnd.n6956 0.152939
R21415 gnd.n6957 gnd.n583 0.152939
R21416 gnd.n6965 gnd.n583 0.152939
R21417 gnd.n6966 gnd.n6965 0.152939
R21418 gnd.n6967 gnd.n6966 0.152939
R21419 gnd.n6967 gnd.n577 0.152939
R21420 gnd.n6975 gnd.n577 0.152939
R21421 gnd.n6976 gnd.n6975 0.152939
R21422 gnd.n6977 gnd.n6976 0.152939
R21423 gnd.n6977 gnd.n571 0.152939
R21424 gnd.n6985 gnd.n571 0.152939
R21425 gnd.n6986 gnd.n6985 0.152939
R21426 gnd.n6987 gnd.n6986 0.152939
R21427 gnd.n6987 gnd.n565 0.152939
R21428 gnd.n6995 gnd.n565 0.152939
R21429 gnd.n6996 gnd.n6995 0.152939
R21430 gnd.n6997 gnd.n6996 0.152939
R21431 gnd.n6997 gnd.n559 0.152939
R21432 gnd.n7005 gnd.n559 0.152939
R21433 gnd.n7006 gnd.n7005 0.152939
R21434 gnd.n7007 gnd.n7006 0.152939
R21435 gnd.n7007 gnd.n553 0.152939
R21436 gnd.n7015 gnd.n553 0.152939
R21437 gnd.n7016 gnd.n7015 0.152939
R21438 gnd.n7017 gnd.n7016 0.152939
R21439 gnd.n7017 gnd.n547 0.152939
R21440 gnd.n7025 gnd.n547 0.152939
R21441 gnd.n7026 gnd.n7025 0.152939
R21442 gnd.n7027 gnd.n7026 0.152939
R21443 gnd.n7027 gnd.n541 0.152939
R21444 gnd.n7035 gnd.n541 0.152939
R21445 gnd.n7036 gnd.n7035 0.152939
R21446 gnd.n7037 gnd.n7036 0.152939
R21447 gnd.n7037 gnd.n535 0.152939
R21448 gnd.n7045 gnd.n535 0.152939
R21449 gnd.n7046 gnd.n7045 0.152939
R21450 gnd.n7047 gnd.n7046 0.152939
R21451 gnd.n7047 gnd.n529 0.152939
R21452 gnd.n7055 gnd.n529 0.152939
R21453 gnd.n7056 gnd.n7055 0.152939
R21454 gnd.n7057 gnd.n7056 0.152939
R21455 gnd.n7057 gnd.n523 0.152939
R21456 gnd.n7065 gnd.n523 0.152939
R21457 gnd.n7066 gnd.n7065 0.152939
R21458 gnd.n7067 gnd.n7066 0.152939
R21459 gnd.n7067 gnd.n517 0.152939
R21460 gnd.n7075 gnd.n517 0.152939
R21461 gnd.n7077 gnd.n7076 0.152939
R21462 gnd.n7077 gnd.n511 0.152939
R21463 gnd.n7085 gnd.n511 0.152939
R21464 gnd.n7086 gnd.n7085 0.152939
R21465 gnd.n7087 gnd.n7086 0.152939
R21466 gnd.n7087 gnd.n505 0.152939
R21467 gnd.n7095 gnd.n505 0.152939
R21468 gnd.n7096 gnd.n7095 0.152939
R21469 gnd.n7097 gnd.n7096 0.152939
R21470 gnd.n7097 gnd.n499 0.152939
R21471 gnd.n7105 gnd.n499 0.152939
R21472 gnd.n7106 gnd.n7105 0.152939
R21473 gnd.n7107 gnd.n7106 0.152939
R21474 gnd.n7107 gnd.n493 0.152939
R21475 gnd.n7115 gnd.n493 0.152939
R21476 gnd.n7116 gnd.n7115 0.152939
R21477 gnd.n7117 gnd.n7116 0.152939
R21478 gnd.n7117 gnd.n487 0.152939
R21479 gnd.n7125 gnd.n487 0.152939
R21480 gnd.n7126 gnd.n7125 0.152939
R21481 gnd.n7127 gnd.n7126 0.152939
R21482 gnd.n7127 gnd.n481 0.152939
R21483 gnd.n7135 gnd.n481 0.152939
R21484 gnd.n7136 gnd.n7135 0.152939
R21485 gnd.n7137 gnd.n7136 0.152939
R21486 gnd.n7137 gnd.n475 0.152939
R21487 gnd.n7145 gnd.n475 0.152939
R21488 gnd.n7146 gnd.n7145 0.152939
R21489 gnd.n7147 gnd.n7146 0.152939
R21490 gnd.n7147 gnd.n469 0.152939
R21491 gnd.n7155 gnd.n469 0.152939
R21492 gnd.n7156 gnd.n7155 0.152939
R21493 gnd.n7157 gnd.n7156 0.152939
R21494 gnd.n7157 gnd.n463 0.152939
R21495 gnd.n7165 gnd.n463 0.152939
R21496 gnd.n7166 gnd.n7165 0.152939
R21497 gnd.n7167 gnd.n7166 0.152939
R21498 gnd.n7167 gnd.n457 0.152939
R21499 gnd.n7175 gnd.n457 0.152939
R21500 gnd.n7176 gnd.n7175 0.152939
R21501 gnd.n7177 gnd.n7176 0.152939
R21502 gnd.n7177 gnd.n451 0.152939
R21503 gnd.n7185 gnd.n451 0.152939
R21504 gnd.n7186 gnd.n7185 0.152939
R21505 gnd.n7187 gnd.n7186 0.152939
R21506 gnd.n7187 gnd.n445 0.152939
R21507 gnd.n7195 gnd.n445 0.152939
R21508 gnd.n7196 gnd.n7195 0.152939
R21509 gnd.n7197 gnd.n7196 0.152939
R21510 gnd.n7197 gnd.n439 0.152939
R21511 gnd.n7205 gnd.n439 0.152939
R21512 gnd.n7206 gnd.n7205 0.152939
R21513 gnd.n7207 gnd.n7206 0.152939
R21514 gnd.n7207 gnd.n433 0.152939
R21515 gnd.n7215 gnd.n433 0.152939
R21516 gnd.n7216 gnd.n7215 0.152939
R21517 gnd.n7217 gnd.n7216 0.152939
R21518 gnd.n7217 gnd.n427 0.152939
R21519 gnd.n7225 gnd.n427 0.152939
R21520 gnd.n7226 gnd.n7225 0.152939
R21521 gnd.n7227 gnd.n7226 0.152939
R21522 gnd.n7227 gnd.n421 0.152939
R21523 gnd.n7235 gnd.n421 0.152939
R21524 gnd.n7236 gnd.n7235 0.152939
R21525 gnd.n7237 gnd.n7236 0.152939
R21526 gnd.n7237 gnd.n415 0.152939
R21527 gnd.n7245 gnd.n415 0.152939
R21528 gnd.n7246 gnd.n7245 0.152939
R21529 gnd.n7247 gnd.n7246 0.152939
R21530 gnd.n7247 gnd.n409 0.152939
R21531 gnd.n7255 gnd.n409 0.152939
R21532 gnd.n7256 gnd.n7255 0.152939
R21533 gnd.n7257 gnd.n7256 0.152939
R21534 gnd.n7257 gnd.n403 0.152939
R21535 gnd.n7265 gnd.n403 0.152939
R21536 gnd.n7266 gnd.n7265 0.152939
R21537 gnd.n7267 gnd.n7266 0.152939
R21538 gnd.n7267 gnd.n397 0.152939
R21539 gnd.n7275 gnd.n397 0.152939
R21540 gnd.n7276 gnd.n7275 0.152939
R21541 gnd.n7277 gnd.n7276 0.152939
R21542 gnd.n7278 gnd.n7277 0.152939
R21543 gnd.n7278 gnd.n391 0.152939
R21544 gnd.n7288 gnd.n391 0.152939
R21545 gnd.n119 gnd.n96 0.152939
R21546 gnd.n120 gnd.n119 0.152939
R21547 gnd.n121 gnd.n120 0.152939
R21548 gnd.n138 gnd.n121 0.152939
R21549 gnd.n139 gnd.n138 0.152939
R21550 gnd.n140 gnd.n139 0.152939
R21551 gnd.n141 gnd.n140 0.152939
R21552 gnd.n156 gnd.n141 0.152939
R21553 gnd.n157 gnd.n156 0.152939
R21554 gnd.n158 gnd.n157 0.152939
R21555 gnd.n159 gnd.n158 0.152939
R21556 gnd.n176 gnd.n159 0.152939
R21557 gnd.n177 gnd.n176 0.152939
R21558 gnd.n178 gnd.n177 0.152939
R21559 gnd.n179 gnd.n178 0.152939
R21560 gnd.n196 gnd.n179 0.152939
R21561 gnd.n197 gnd.n196 0.152939
R21562 gnd.n198 gnd.n197 0.152939
R21563 gnd.n199 gnd.n198 0.152939
R21564 gnd.n214 gnd.n199 0.152939
R21565 gnd.n7546 gnd.n214 0.152939
R21566 gnd.n7627 gnd.n84 0.152939
R21567 gnd.n7360 gnd.n84 0.152939
R21568 gnd.n7361 gnd.n7360 0.152939
R21569 gnd.n7362 gnd.n7361 0.152939
R21570 gnd.n7362 gnd.n367 0.152939
R21571 gnd.n7367 gnd.n367 0.152939
R21572 gnd.n7368 gnd.n7367 0.152939
R21573 gnd.n7369 gnd.n7368 0.152939
R21574 gnd.n7369 gnd.n364 0.152939
R21575 gnd.n7374 gnd.n364 0.152939
R21576 gnd.n7375 gnd.n7374 0.152939
R21577 gnd.n7376 gnd.n7375 0.152939
R21578 gnd.n7376 gnd.n361 0.152939
R21579 gnd.n7381 gnd.n361 0.152939
R21580 gnd.n7382 gnd.n7381 0.152939
R21581 gnd.n7383 gnd.n7382 0.152939
R21582 gnd.n7383 gnd.n358 0.152939
R21583 gnd.n7388 gnd.n358 0.152939
R21584 gnd.n7389 gnd.n7388 0.152939
R21585 gnd.n7390 gnd.n7389 0.152939
R21586 gnd.n7390 gnd.n355 0.152939
R21587 gnd.n7395 gnd.n355 0.152939
R21588 gnd.n7396 gnd.n7395 0.152939
R21589 gnd.n7397 gnd.n7396 0.152939
R21590 gnd.n7397 gnd.n352 0.152939
R21591 gnd.n7402 gnd.n352 0.152939
R21592 gnd.n7435 gnd.n318 0.152939
R21593 gnd.n320 gnd.n318 0.152939
R21594 gnd.n324 gnd.n320 0.152939
R21595 gnd.n325 gnd.n324 0.152939
R21596 gnd.n326 gnd.n325 0.152939
R21597 gnd.n327 gnd.n326 0.152939
R21598 gnd.n331 gnd.n327 0.152939
R21599 gnd.n332 gnd.n331 0.152939
R21600 gnd.n333 gnd.n332 0.152939
R21601 gnd.n334 gnd.n333 0.152939
R21602 gnd.n338 gnd.n334 0.152939
R21603 gnd.n339 gnd.n338 0.152939
R21604 gnd.n340 gnd.n339 0.152939
R21605 gnd.n341 gnd.n340 0.152939
R21606 gnd.n345 gnd.n341 0.152939
R21607 gnd.n346 gnd.n345 0.152939
R21608 gnd.n7404 gnd.n346 0.152939
R21609 gnd.n7404 gnd.n7403 0.152939
R21610 gnd.n7545 gnd.n215 0.152939
R21611 gnd.n217 gnd.n215 0.152939
R21612 gnd.n221 gnd.n217 0.152939
R21613 gnd.n222 gnd.n221 0.152939
R21614 gnd.n223 gnd.n222 0.152939
R21615 gnd.n224 gnd.n223 0.152939
R21616 gnd.n228 gnd.n224 0.152939
R21617 gnd.n229 gnd.n228 0.152939
R21618 gnd.n230 gnd.n229 0.152939
R21619 gnd.n231 gnd.n230 0.152939
R21620 gnd.n235 gnd.n231 0.152939
R21621 gnd.n236 gnd.n235 0.152939
R21622 gnd.n237 gnd.n236 0.152939
R21623 gnd.n238 gnd.n237 0.152939
R21624 gnd.n242 gnd.n238 0.152939
R21625 gnd.n243 gnd.n242 0.152939
R21626 gnd.n244 gnd.n243 0.152939
R21627 gnd.n245 gnd.n244 0.152939
R21628 gnd.n249 gnd.n245 0.152939
R21629 gnd.n250 gnd.n249 0.152939
R21630 gnd.n251 gnd.n250 0.152939
R21631 gnd.n252 gnd.n251 0.152939
R21632 gnd.n256 gnd.n252 0.152939
R21633 gnd.n257 gnd.n256 0.152939
R21634 gnd.n258 gnd.n257 0.152939
R21635 gnd.n259 gnd.n258 0.152939
R21636 gnd.n263 gnd.n259 0.152939
R21637 gnd.n264 gnd.n263 0.152939
R21638 gnd.n265 gnd.n264 0.152939
R21639 gnd.n266 gnd.n265 0.152939
R21640 gnd.n270 gnd.n266 0.152939
R21641 gnd.n271 gnd.n270 0.152939
R21642 gnd.n272 gnd.n271 0.152939
R21643 gnd.n273 gnd.n272 0.152939
R21644 gnd.n277 gnd.n273 0.152939
R21645 gnd.n278 gnd.n277 0.152939
R21646 gnd.n7476 gnd.n278 0.152939
R21647 gnd.n7476 gnd.n7475 0.152939
R21648 gnd.n7475 gnd.n7474 0.152939
R21649 gnd.n7474 gnd.n282 0.152939
R21650 gnd.n288 gnd.n282 0.152939
R21651 gnd.n289 gnd.n288 0.152939
R21652 gnd.n290 gnd.n289 0.152939
R21653 gnd.n291 gnd.n290 0.152939
R21654 gnd.n295 gnd.n291 0.152939
R21655 gnd.n296 gnd.n295 0.152939
R21656 gnd.n297 gnd.n296 0.152939
R21657 gnd.n298 gnd.n297 0.152939
R21658 gnd.n302 gnd.n298 0.152939
R21659 gnd.n303 gnd.n302 0.152939
R21660 gnd.n304 gnd.n303 0.152939
R21661 gnd.n305 gnd.n304 0.152939
R21662 gnd.n309 gnd.n305 0.152939
R21663 gnd.n310 gnd.n309 0.152939
R21664 gnd.n311 gnd.n310 0.152939
R21665 gnd.n312 gnd.n311 0.152939
R21666 gnd.n317 gnd.n312 0.152939
R21667 gnd.n7437 gnd.n317 0.152939
R21668 gnd.n1512 gnd.n1511 0.152939
R21669 gnd.n1513 gnd.n1512 0.152939
R21670 gnd.n1514 gnd.n1513 0.152939
R21671 gnd.n1515 gnd.n1514 0.152939
R21672 gnd.n1516 gnd.n1515 0.152939
R21673 gnd.n1517 gnd.n1516 0.152939
R21674 gnd.n1518 gnd.n1517 0.152939
R21675 gnd.n1519 gnd.n1518 0.152939
R21676 gnd.n1520 gnd.n1519 0.152939
R21677 gnd.n1521 gnd.n1520 0.152939
R21678 gnd.n1522 gnd.n1521 0.152939
R21679 gnd.n1523 gnd.n1522 0.152939
R21680 gnd.n1524 gnd.n1523 0.152939
R21681 gnd.n1525 gnd.n1524 0.152939
R21682 gnd.n1526 gnd.n1525 0.152939
R21683 gnd.n1527 gnd.n1526 0.152939
R21684 gnd.n1528 gnd.n1527 0.152939
R21685 gnd.n1531 gnd.n1528 0.152939
R21686 gnd.n1532 gnd.n1531 0.152939
R21687 gnd.n1533 gnd.n1532 0.152939
R21688 gnd.n1534 gnd.n1533 0.152939
R21689 gnd.n1535 gnd.n1534 0.152939
R21690 gnd.n1536 gnd.n1535 0.152939
R21691 gnd.n1537 gnd.n1536 0.152939
R21692 gnd.n1538 gnd.n1537 0.152939
R21693 gnd.n1543 gnd.n1542 0.152939
R21694 gnd.n1544 gnd.n1543 0.152939
R21695 gnd.n1545 gnd.n1544 0.152939
R21696 gnd.n1546 gnd.n1545 0.152939
R21697 gnd.n1547 gnd.n1546 0.152939
R21698 gnd.n1548 gnd.n1547 0.152939
R21699 gnd.n1549 gnd.n1548 0.152939
R21700 gnd.n1550 gnd.n1549 0.152939
R21701 gnd.n1551 gnd.n1550 0.152939
R21702 gnd.n1554 gnd.n1551 0.152939
R21703 gnd.n1555 gnd.n1554 0.152939
R21704 gnd.n1556 gnd.n1555 0.152939
R21705 gnd.n1557 gnd.n1556 0.152939
R21706 gnd.n1558 gnd.n1557 0.152939
R21707 gnd.n1559 gnd.n1558 0.152939
R21708 gnd.n1560 gnd.n1559 0.152939
R21709 gnd.n1561 gnd.n1560 0.152939
R21710 gnd.n1562 gnd.n1561 0.152939
R21711 gnd.n1563 gnd.n1562 0.152939
R21712 gnd.n1564 gnd.n1563 0.152939
R21713 gnd.n1565 gnd.n1564 0.152939
R21714 gnd.n1566 gnd.n1565 0.152939
R21715 gnd.n1567 gnd.n1566 0.152939
R21716 gnd.n1568 gnd.n1567 0.152939
R21717 gnd.n1569 gnd.n1568 0.152939
R21718 gnd.n1570 gnd.n1569 0.152939
R21719 gnd.n1571 gnd.n1570 0.152939
R21720 gnd.n1572 gnd.n1571 0.152939
R21721 gnd.n5966 gnd.n1572 0.152939
R21722 gnd.n5966 gnd.n5965 0.152939
R21723 gnd.n1593 gnd.n1592 0.152939
R21724 gnd.n1594 gnd.n1593 0.152939
R21725 gnd.n1595 gnd.n1594 0.152939
R21726 gnd.n1596 gnd.n1595 0.152939
R21727 gnd.n1616 gnd.n1596 0.152939
R21728 gnd.n1617 gnd.n1616 0.152939
R21729 gnd.n1618 gnd.n1617 0.152939
R21730 gnd.n1619 gnd.n1618 0.152939
R21731 gnd.n1637 gnd.n1619 0.152939
R21732 gnd.n1638 gnd.n1637 0.152939
R21733 gnd.n1639 gnd.n1638 0.152939
R21734 gnd.n1640 gnd.n1639 0.152939
R21735 gnd.n1656 gnd.n1640 0.152939
R21736 gnd.n1657 gnd.n1656 0.152939
R21737 gnd.n1658 gnd.n1657 0.152939
R21738 gnd.n1659 gnd.n1658 0.152939
R21739 gnd.n1677 gnd.n1659 0.152939
R21740 gnd.n1678 gnd.n1677 0.152939
R21741 gnd.n1679 gnd.n1678 0.152939
R21742 gnd.n1680 gnd.n1679 0.152939
R21743 gnd.n1680 gnd.n97 0.152939
R21744 gnd.n5880 gnd.n1702 0.152939
R21745 gnd.n5881 gnd.n5880 0.152939
R21746 gnd.n5883 gnd.n5881 0.152939
R21747 gnd.n5883 gnd.n5882 0.152939
R21748 gnd.n7289 gnd.n390 0.152939
R21749 gnd.n4627 gnd.n4626 0.152939
R21750 gnd.n4630 gnd.n4627 0.152939
R21751 gnd.n4631 gnd.n4630 0.152939
R21752 gnd.n4632 gnd.n4631 0.152939
R21753 gnd.n4633 gnd.n4632 0.152939
R21754 gnd.n4635 gnd.n4633 0.152939
R21755 gnd.n4635 gnd.n4634 0.152939
R21756 gnd.n4634 gnd.n2483 0.152939
R21757 gnd.n4714 gnd.n2483 0.152939
R21758 gnd.n4715 gnd.n4714 0.152939
R21759 gnd.n4716 gnd.n4715 0.152939
R21760 gnd.n4716 gnd.n2479 0.152939
R21761 gnd.n4722 gnd.n2479 0.152939
R21762 gnd.n4723 gnd.n4722 0.152939
R21763 gnd.n4724 gnd.n4723 0.152939
R21764 gnd.n4725 gnd.n4724 0.152939
R21765 gnd.n4726 gnd.n4725 0.152939
R21766 gnd.n4729 gnd.n4726 0.152939
R21767 gnd.n4730 gnd.n4729 0.152939
R21768 gnd.n4731 gnd.n4730 0.152939
R21769 gnd.n4732 gnd.n4731 0.152939
R21770 gnd.n4736 gnd.n4732 0.152939
R21771 gnd.n4737 gnd.n4736 0.152939
R21772 gnd.n4738 gnd.n4737 0.152939
R21773 gnd.n4738 gnd.n2200 0.152939
R21774 gnd.n4861 gnd.n2200 0.152939
R21775 gnd.n4862 gnd.n4861 0.152939
R21776 gnd.n4863 gnd.n4862 0.152939
R21777 gnd.n4863 gnd.n2187 0.152939
R21778 gnd.n4877 gnd.n2187 0.152939
R21779 gnd.n4878 gnd.n4877 0.152939
R21780 gnd.n4879 gnd.n4878 0.152939
R21781 gnd.n4879 gnd.n2173 0.152939
R21782 gnd.n4893 gnd.n2173 0.152939
R21783 gnd.n4894 gnd.n4893 0.152939
R21784 gnd.n4895 gnd.n4894 0.152939
R21785 gnd.n4895 gnd.n2158 0.152939
R21786 gnd.n4909 gnd.n2158 0.152939
R21787 gnd.n4910 gnd.n4909 0.152939
R21788 gnd.n4911 gnd.n4910 0.152939
R21789 gnd.n4911 gnd.n2144 0.152939
R21790 gnd.n4925 gnd.n2144 0.152939
R21791 gnd.n4926 gnd.n4925 0.152939
R21792 gnd.n4927 gnd.n4926 0.152939
R21793 gnd.n4927 gnd.n2129 0.152939
R21794 gnd.n4967 gnd.n2129 0.152939
R21795 gnd.n4968 gnd.n4967 0.152939
R21796 gnd.n4969 gnd.n4968 0.152939
R21797 gnd.n4971 gnd.n4969 0.152939
R21798 gnd.n4971 gnd.n4970 0.152939
R21799 gnd.n4970 gnd.n1191 0.152939
R21800 gnd.n1192 gnd.n1191 0.152939
R21801 gnd.n1193 gnd.n1192 0.152939
R21802 gnd.n1294 gnd.n1193 0.152939
R21803 gnd.n1295 gnd.n1294 0.152939
R21804 gnd.n1296 gnd.n1295 0.152939
R21805 gnd.n1297 gnd.n1296 0.152939
R21806 gnd.n1298 gnd.n1297 0.152939
R21807 gnd.n2101 gnd.n1298 0.152939
R21808 gnd.n5039 gnd.n2101 0.152939
R21809 gnd.n5040 gnd.n5039 0.152939
R21810 gnd.n5041 gnd.n5040 0.152939
R21811 gnd.n5041 gnd.n2075 0.152939
R21812 gnd.n5098 gnd.n2075 0.152939
R21813 gnd.n5099 gnd.n5098 0.152939
R21814 gnd.n5100 gnd.n5099 0.152939
R21815 gnd.n5101 gnd.n5100 0.152939
R21816 gnd.n5101 gnd.n2052 0.152939
R21817 gnd.n5130 gnd.n2052 0.152939
R21818 gnd.n5131 gnd.n5130 0.152939
R21819 gnd.n5132 gnd.n5131 0.152939
R21820 gnd.n5133 gnd.n5132 0.152939
R21821 gnd.n5133 gnd.n2030 0.152939
R21822 gnd.n5180 gnd.n2030 0.152939
R21823 gnd.n5181 gnd.n5180 0.152939
R21824 gnd.n5182 gnd.n5181 0.152939
R21825 gnd.n5183 gnd.n5182 0.152939
R21826 gnd.n5183 gnd.n2002 0.152939
R21827 gnd.n5218 gnd.n2002 0.152939
R21828 gnd.n5219 gnd.n5218 0.152939
R21829 gnd.n5220 gnd.n5219 0.152939
R21830 gnd.n5220 gnd.n1974 0.152939
R21831 gnd.n5255 gnd.n1974 0.152939
R21832 gnd.n5256 gnd.n5255 0.152939
R21833 gnd.n5257 gnd.n5256 0.152939
R21834 gnd.n5258 gnd.n5257 0.152939
R21835 gnd.n5258 gnd.n1955 0.152939
R21836 gnd.n5313 gnd.n1955 0.152939
R21837 gnd.n5314 gnd.n5313 0.152939
R21838 gnd.n5315 gnd.n5314 0.152939
R21839 gnd.n5316 gnd.n5315 0.152939
R21840 gnd.n5316 gnd.n1932 0.152939
R21841 gnd.n5351 gnd.n1932 0.152939
R21842 gnd.n5352 gnd.n5351 0.152939
R21843 gnd.n5353 gnd.n5352 0.152939
R21844 gnd.n5354 gnd.n5353 0.152939
R21845 gnd.n5354 gnd.n1904 0.152939
R21846 gnd.n5407 gnd.n1904 0.152939
R21847 gnd.n5408 gnd.n5407 0.152939
R21848 gnd.n5409 gnd.n5408 0.152939
R21849 gnd.n5410 gnd.n5409 0.152939
R21850 gnd.n5410 gnd.n1883 0.152939
R21851 gnd.n5445 gnd.n1883 0.152939
R21852 gnd.n5446 gnd.n5445 0.152939
R21853 gnd.n5447 gnd.n5446 0.152939
R21854 gnd.n5447 gnd.n1827 0.152939
R21855 gnd.n5620 gnd.n1827 0.152939
R21856 gnd.n5621 gnd.n5620 0.152939
R21857 gnd.n5622 gnd.n5621 0.152939
R21858 gnd.n5622 gnd.n1816 0.152939
R21859 gnd.n5637 gnd.n1816 0.152939
R21860 gnd.n5638 gnd.n5637 0.152939
R21861 gnd.n5639 gnd.n5638 0.152939
R21862 gnd.n5639 gnd.n1804 0.152939
R21863 gnd.n5654 gnd.n1804 0.152939
R21864 gnd.n5655 gnd.n5654 0.152939
R21865 gnd.n5656 gnd.n5655 0.152939
R21866 gnd.n5656 gnd.n1792 0.152939
R21867 gnd.n5671 gnd.n1792 0.152939
R21868 gnd.n5672 gnd.n5671 0.152939
R21869 gnd.n5673 gnd.n5672 0.152939
R21870 gnd.n5673 gnd.n1780 0.152939
R21871 gnd.n5688 gnd.n1780 0.152939
R21872 gnd.n5689 gnd.n5688 0.152939
R21873 gnd.n5690 gnd.n5689 0.152939
R21874 gnd.n5692 gnd.n5690 0.152939
R21875 gnd.n5692 gnd.n5691 0.152939
R21876 gnd.n5691 gnd.n1768 0.152939
R21877 gnd.n5710 gnd.n1768 0.152939
R21878 gnd.n5711 gnd.n5710 0.152939
R21879 gnd.n5712 gnd.n5711 0.152939
R21880 gnd.n5713 gnd.n5712 0.152939
R21881 gnd.n5714 gnd.n5713 0.152939
R21882 gnd.n5716 gnd.n5714 0.152939
R21883 gnd.n5717 gnd.n5716 0.152939
R21884 gnd.n5717 gnd.n1732 0.152939
R21885 gnd.n5779 gnd.n1732 0.152939
R21886 gnd.n5780 gnd.n5779 0.152939
R21887 gnd.n5781 gnd.n5780 0.152939
R21888 gnd.n5781 gnd.n1728 0.152939
R21889 gnd.n5787 gnd.n1728 0.152939
R21890 gnd.n5788 gnd.n5787 0.152939
R21891 gnd.n5789 gnd.n5788 0.152939
R21892 gnd.n5789 gnd.n1724 0.152939
R21893 gnd.n5795 gnd.n1724 0.152939
R21894 gnd.n5796 gnd.n5795 0.152939
R21895 gnd.n5797 gnd.n5796 0.152939
R21896 gnd.n5798 gnd.n5797 0.152939
R21897 gnd.n5799 gnd.n5798 0.152939
R21898 gnd.n5802 gnd.n5799 0.152939
R21899 gnd.n5803 gnd.n5802 0.152939
R21900 gnd.n5804 gnd.n5803 0.152939
R21901 gnd.n5805 gnd.n5804 0.152939
R21902 gnd.n5807 gnd.n5805 0.152939
R21903 gnd.n5807 gnd.n5806 0.152939
R21904 gnd.n5806 gnd.n1702 0.152939
R21905 gnd.n4283 gnd.n4249 0.152939
R21906 gnd.n4250 gnd.n4249 0.152939
R21907 gnd.n4251 gnd.n4250 0.152939
R21908 gnd.n4252 gnd.n4251 0.152939
R21909 gnd.n4253 gnd.n4252 0.152939
R21910 gnd.n4254 gnd.n4253 0.152939
R21911 gnd.n4255 gnd.n4254 0.152939
R21912 gnd.n4256 gnd.n4255 0.152939
R21913 gnd.n4257 gnd.n4256 0.152939
R21914 gnd.n4258 gnd.n4257 0.152939
R21915 gnd.n4259 gnd.n4258 0.152939
R21916 gnd.n4260 gnd.n4259 0.152939
R21917 gnd.n4261 gnd.n4260 0.152939
R21918 gnd.n4261 gnd.n2569 0.152939
R21919 gnd.n4528 gnd.n2569 0.152939
R21920 gnd.n4529 gnd.n4528 0.152939
R21921 gnd.n4530 gnd.n4529 0.152939
R21922 gnd.n4531 gnd.n4530 0.152939
R21923 gnd.n4532 gnd.n4531 0.152939
R21924 gnd.n4533 gnd.n4532 0.152939
R21925 gnd.n4534 gnd.n4533 0.152939
R21926 gnd.n4535 gnd.n4534 0.152939
R21927 gnd.n4535 gnd.n2533 0.152939
R21928 gnd.n4589 gnd.n2533 0.152939
R21929 gnd.n4590 gnd.n4589 0.152939
R21930 gnd.n4591 gnd.n4590 0.152939
R21931 gnd.n4322 gnd.n4230 0.152939
R21932 gnd.n4231 gnd.n4230 0.152939
R21933 gnd.n4232 gnd.n4231 0.152939
R21934 gnd.n4233 gnd.n4232 0.152939
R21935 gnd.n4234 gnd.n4233 0.152939
R21936 gnd.n4235 gnd.n4234 0.152939
R21937 gnd.n4236 gnd.n4235 0.152939
R21938 gnd.n4237 gnd.n4236 0.152939
R21939 gnd.n4238 gnd.n4237 0.152939
R21940 gnd.n4239 gnd.n4238 0.152939
R21941 gnd.n4240 gnd.n4239 0.152939
R21942 gnd.n4241 gnd.n4240 0.152939
R21943 gnd.n4242 gnd.n4241 0.152939
R21944 gnd.n4243 gnd.n4242 0.152939
R21945 gnd.n4244 gnd.n4243 0.152939
R21946 gnd.n4287 gnd.n4244 0.152939
R21947 gnd.n4287 gnd.n4286 0.152939
R21948 gnd.n4286 gnd.n4285 0.152939
R21949 gnd.n971 gnd.n946 0.152939
R21950 gnd.n972 gnd.n971 0.152939
R21951 gnd.n973 gnd.n972 0.152939
R21952 gnd.n991 gnd.n973 0.152939
R21953 gnd.n992 gnd.n991 0.152939
R21954 gnd.n993 gnd.n992 0.152939
R21955 gnd.n994 gnd.n993 0.152939
R21956 gnd.n1010 gnd.n994 0.152939
R21957 gnd.n1011 gnd.n1010 0.152939
R21958 gnd.n1012 gnd.n1011 0.152939
R21959 gnd.n1013 gnd.n1012 0.152939
R21960 gnd.n1031 gnd.n1013 0.152939
R21961 gnd.n1032 gnd.n1031 0.152939
R21962 gnd.n1033 gnd.n1032 0.152939
R21963 gnd.n1034 gnd.n1033 0.152939
R21964 gnd.n1051 gnd.n1034 0.152939
R21965 gnd.n1052 gnd.n1051 0.152939
R21966 gnd.n1053 gnd.n1052 0.152939
R21967 gnd.n1054 gnd.n1053 0.152939
R21968 gnd.n1070 gnd.n1054 0.152939
R21969 gnd.n6407 gnd.n1070 0.152939
R21970 gnd.n6406 gnd.n1071 0.152939
R21971 gnd.n1076 gnd.n1071 0.152939
R21972 gnd.n1077 gnd.n1076 0.152939
R21973 gnd.n1078 gnd.n1077 0.152939
R21974 gnd.n1079 gnd.n1078 0.152939
R21975 gnd.n1080 gnd.n1079 0.152939
R21976 gnd.n1084 gnd.n1080 0.152939
R21977 gnd.n1085 gnd.n1084 0.152939
R21978 gnd.n1086 gnd.n1085 0.152939
R21979 gnd.n1087 gnd.n1086 0.152939
R21980 gnd.n1091 gnd.n1087 0.152939
R21981 gnd.n1092 gnd.n1091 0.152939
R21982 gnd.n1093 gnd.n1092 0.152939
R21983 gnd.n1094 gnd.n1093 0.152939
R21984 gnd.n1098 gnd.n1094 0.152939
R21985 gnd.n1099 gnd.n1098 0.152939
R21986 gnd.n1100 gnd.n1099 0.152939
R21987 gnd.n1103 gnd.n1100 0.152939
R21988 gnd.n1107 gnd.n1103 0.152939
R21989 gnd.n1108 gnd.n1107 0.152939
R21990 gnd.n1109 gnd.n1108 0.152939
R21991 gnd.n1110 gnd.n1109 0.152939
R21992 gnd.n1114 gnd.n1110 0.152939
R21993 gnd.n1115 gnd.n1114 0.152939
R21994 gnd.n1116 gnd.n1115 0.152939
R21995 gnd.n2310 gnd.n2309 0.152939
R21996 gnd.n2319 gnd.n2310 0.152939
R21997 gnd.n2320 gnd.n2319 0.152939
R21998 gnd.n2321 gnd.n2320 0.152939
R21999 gnd.n2321 gnd.n2305 0.152939
R22000 gnd.n2329 gnd.n2305 0.152939
R22001 gnd.n2330 gnd.n2329 0.152939
R22002 gnd.n2331 gnd.n2330 0.152939
R22003 gnd.n2331 gnd.n2299 0.152939
R22004 gnd.n2339 gnd.n2299 0.152939
R22005 gnd.n2340 gnd.n2339 0.152939
R22006 gnd.n2341 gnd.n2340 0.152939
R22007 gnd.n2341 gnd.n2295 0.152939
R22008 gnd.n2349 gnd.n2295 0.152939
R22009 gnd.n2350 gnd.n2349 0.152939
R22010 gnd.n2351 gnd.n2350 0.152939
R22011 gnd.n2351 gnd.n2291 0.152939
R22012 gnd.n2359 gnd.n2291 0.152939
R22013 gnd.n2360 gnd.n2359 0.152939
R22014 gnd.n2361 gnd.n2360 0.152939
R22015 gnd.n2361 gnd.n2287 0.152939
R22016 gnd.n2369 gnd.n2287 0.152939
R22017 gnd.n2370 gnd.n2369 0.152939
R22018 gnd.n2371 gnd.n2370 0.152939
R22019 gnd.n2371 gnd.n2283 0.152939
R22020 gnd.n2379 gnd.n2283 0.152939
R22021 gnd.n2380 gnd.n2379 0.152939
R22022 gnd.n2381 gnd.n2380 0.152939
R22023 gnd.n2381 gnd.n2277 0.152939
R22024 gnd.n2388 gnd.n2277 0.152939
R22025 gnd.n4168 gnd.n4167 0.152939
R22026 gnd.n4169 gnd.n4168 0.152939
R22027 gnd.n4170 gnd.n4169 0.152939
R22028 gnd.n4171 gnd.n4170 0.152939
R22029 gnd.n4172 gnd.n4171 0.152939
R22030 gnd.n4173 gnd.n4172 0.152939
R22031 gnd.n4174 gnd.n4173 0.152939
R22032 gnd.n4175 gnd.n4174 0.152939
R22033 gnd.n4176 gnd.n4175 0.152939
R22034 gnd.n4177 gnd.n4176 0.152939
R22035 gnd.n4178 gnd.n4177 0.152939
R22036 gnd.n4179 gnd.n4178 0.152939
R22037 gnd.n4180 gnd.n4179 0.152939
R22038 gnd.n4181 gnd.n4180 0.152939
R22039 gnd.n4182 gnd.n4181 0.152939
R22040 gnd.n4183 gnd.n4182 0.152939
R22041 gnd.n4184 gnd.n4183 0.152939
R22042 gnd.n4187 gnd.n4184 0.152939
R22043 gnd.n4188 gnd.n4187 0.152939
R22044 gnd.n4189 gnd.n4188 0.152939
R22045 gnd.n4190 gnd.n4189 0.152939
R22046 gnd.n4191 gnd.n4190 0.152939
R22047 gnd.n4192 gnd.n4191 0.152939
R22048 gnd.n4193 gnd.n4192 0.152939
R22049 gnd.n4194 gnd.n4193 0.152939
R22050 gnd.n4195 gnd.n4194 0.152939
R22051 gnd.n4196 gnd.n4195 0.152939
R22052 gnd.n4197 gnd.n4196 0.152939
R22053 gnd.n4198 gnd.n4197 0.152939
R22054 gnd.n4199 gnd.n4198 0.152939
R22055 gnd.n4200 gnd.n4199 0.152939
R22056 gnd.n4201 gnd.n4200 0.152939
R22057 gnd.n4202 gnd.n4201 0.152939
R22058 gnd.n4203 gnd.n4202 0.152939
R22059 gnd.n4204 gnd.n4203 0.152939
R22060 gnd.n4205 gnd.n4204 0.152939
R22061 gnd.n4206 gnd.n4205 0.152939
R22062 gnd.n4209 gnd.n4206 0.152939
R22063 gnd.n4210 gnd.n4209 0.152939
R22064 gnd.n4211 gnd.n4210 0.152939
R22065 gnd.n4212 gnd.n4211 0.152939
R22066 gnd.n4213 gnd.n4212 0.152939
R22067 gnd.n4214 gnd.n4213 0.152939
R22068 gnd.n4215 gnd.n4214 0.152939
R22069 gnd.n4216 gnd.n4215 0.152939
R22070 gnd.n4217 gnd.n4216 0.152939
R22071 gnd.n4218 gnd.n4217 0.152939
R22072 gnd.n4219 gnd.n4218 0.152939
R22073 gnd.n4220 gnd.n4219 0.152939
R22074 gnd.n4221 gnd.n4220 0.152939
R22075 gnd.n4222 gnd.n4221 0.152939
R22076 gnd.n4223 gnd.n4222 0.152939
R22077 gnd.n4224 gnd.n4223 0.152939
R22078 gnd.n4225 gnd.n4224 0.152939
R22079 gnd.n4226 gnd.n4225 0.152939
R22080 gnd.n4227 gnd.n4226 0.152939
R22081 gnd.n4325 gnd.n4227 0.152939
R22082 gnd.n4325 gnd.n4324 0.152939
R22083 gnd.n4454 gnd.n2633 0.152939
R22084 gnd.n4455 gnd.n4454 0.152939
R22085 gnd.n4456 gnd.n4455 0.152939
R22086 gnd.n4456 gnd.n2614 0.152939
R22087 gnd.n4474 gnd.n2614 0.152939
R22088 gnd.n4475 gnd.n4474 0.152939
R22089 gnd.n4476 gnd.n4475 0.152939
R22090 gnd.n4476 gnd.n2597 0.152939
R22091 gnd.n4494 gnd.n2597 0.152939
R22092 gnd.n4495 gnd.n4494 0.152939
R22093 gnd.n4496 gnd.n4495 0.152939
R22094 gnd.n4496 gnd.n2577 0.152939
R22095 gnd.n4518 gnd.n2577 0.152939
R22096 gnd.n4519 gnd.n4518 0.152939
R22097 gnd.n4520 gnd.n4519 0.152939
R22098 gnd.n4521 gnd.n4520 0.152939
R22099 gnd.n4521 gnd.n2553 0.152939
R22100 gnd.n4559 gnd.n2553 0.152939
R22101 gnd.n4560 gnd.n4559 0.152939
R22102 gnd.n4561 gnd.n4560 0.152939
R22103 gnd.n4561 gnd.n947 0.152939
R22104 gnd.n2513 gnd.n2512 0.152939
R22105 gnd.n4624 gnd.n4623 0.152939
R22106 gnd.n4625 gnd.n4624 0.152939
R22107 gnd.n4626 gnd.n4625 0.152939
R22108 gnd.n6655 gnd.n769 0.152939
R22109 gnd.n774 gnd.n769 0.152939
R22110 gnd.n775 gnd.n774 0.152939
R22111 gnd.n776 gnd.n775 0.152939
R22112 gnd.n781 gnd.n776 0.152939
R22113 gnd.n782 gnd.n781 0.152939
R22114 gnd.n783 gnd.n782 0.152939
R22115 gnd.n784 gnd.n783 0.152939
R22116 gnd.n789 gnd.n784 0.152939
R22117 gnd.n790 gnd.n789 0.152939
R22118 gnd.n791 gnd.n790 0.152939
R22119 gnd.n792 gnd.n791 0.152939
R22120 gnd.n797 gnd.n792 0.152939
R22121 gnd.n798 gnd.n797 0.152939
R22122 gnd.n799 gnd.n798 0.152939
R22123 gnd.n800 gnd.n799 0.152939
R22124 gnd.n805 gnd.n800 0.152939
R22125 gnd.n806 gnd.n805 0.152939
R22126 gnd.n807 gnd.n806 0.152939
R22127 gnd.n808 gnd.n807 0.152939
R22128 gnd.n813 gnd.n808 0.152939
R22129 gnd.n814 gnd.n813 0.152939
R22130 gnd.n815 gnd.n814 0.152939
R22131 gnd.n816 gnd.n815 0.152939
R22132 gnd.n821 gnd.n816 0.152939
R22133 gnd.n822 gnd.n821 0.152939
R22134 gnd.n823 gnd.n822 0.152939
R22135 gnd.n824 gnd.n823 0.152939
R22136 gnd.n829 gnd.n824 0.152939
R22137 gnd.n830 gnd.n829 0.152939
R22138 gnd.n831 gnd.n830 0.152939
R22139 gnd.n832 gnd.n831 0.152939
R22140 gnd.n837 gnd.n832 0.152939
R22141 gnd.n838 gnd.n837 0.152939
R22142 gnd.n839 gnd.n838 0.152939
R22143 gnd.n840 gnd.n839 0.152939
R22144 gnd.n845 gnd.n840 0.152939
R22145 gnd.n846 gnd.n845 0.152939
R22146 gnd.n847 gnd.n846 0.152939
R22147 gnd.n848 gnd.n847 0.152939
R22148 gnd.n853 gnd.n848 0.152939
R22149 gnd.n854 gnd.n853 0.152939
R22150 gnd.n855 gnd.n854 0.152939
R22151 gnd.n856 gnd.n855 0.152939
R22152 gnd.n861 gnd.n856 0.152939
R22153 gnd.n862 gnd.n861 0.152939
R22154 gnd.n863 gnd.n862 0.152939
R22155 gnd.n864 gnd.n863 0.152939
R22156 gnd.n869 gnd.n864 0.152939
R22157 gnd.n870 gnd.n869 0.152939
R22158 gnd.n871 gnd.n870 0.152939
R22159 gnd.n872 gnd.n871 0.152939
R22160 gnd.n877 gnd.n872 0.152939
R22161 gnd.n878 gnd.n877 0.152939
R22162 gnd.n879 gnd.n878 0.152939
R22163 gnd.n880 gnd.n879 0.152939
R22164 gnd.n885 gnd.n880 0.152939
R22165 gnd.n886 gnd.n885 0.152939
R22166 gnd.n887 gnd.n886 0.152939
R22167 gnd.n888 gnd.n887 0.152939
R22168 gnd.n893 gnd.n888 0.152939
R22169 gnd.n894 gnd.n893 0.152939
R22170 gnd.n895 gnd.n894 0.152939
R22171 gnd.n896 gnd.n895 0.152939
R22172 gnd.n901 gnd.n896 0.152939
R22173 gnd.n902 gnd.n901 0.152939
R22174 gnd.n903 gnd.n902 0.152939
R22175 gnd.n904 gnd.n903 0.152939
R22176 gnd.n909 gnd.n904 0.152939
R22177 gnd.n910 gnd.n909 0.152939
R22178 gnd.n911 gnd.n910 0.152939
R22179 gnd.n912 gnd.n911 0.152939
R22180 gnd.n917 gnd.n912 0.152939
R22181 gnd.n918 gnd.n917 0.152939
R22182 gnd.n919 gnd.n918 0.152939
R22183 gnd.n920 gnd.n919 0.152939
R22184 gnd.n925 gnd.n920 0.152939
R22185 gnd.n926 gnd.n925 0.152939
R22186 gnd.n927 gnd.n926 0.152939
R22187 gnd.n928 gnd.n927 0.152939
R22188 gnd.n933 gnd.n928 0.152939
R22189 gnd.n934 gnd.n933 0.152939
R22190 gnd.n935 gnd.n934 0.152939
R22191 gnd.n936 gnd.n935 0.152939
R22192 gnd.n4870 gnd.n4869 0.152939
R22193 gnd.n4871 gnd.n4870 0.152939
R22194 gnd.n4871 gnd.n2180 0.152939
R22195 gnd.n4885 gnd.n2180 0.152939
R22196 gnd.n4886 gnd.n4885 0.152939
R22197 gnd.n4887 gnd.n4886 0.152939
R22198 gnd.n4887 gnd.n2166 0.152939
R22199 gnd.n4901 gnd.n2166 0.152939
R22200 gnd.n4902 gnd.n4901 0.152939
R22201 gnd.n4903 gnd.n4902 0.152939
R22202 gnd.n4903 gnd.n2152 0.152939
R22203 gnd.n4917 gnd.n2152 0.152939
R22204 gnd.n4918 gnd.n4917 0.152939
R22205 gnd.n4919 gnd.n4918 0.152939
R22206 gnd.n4919 gnd.n2138 0.152939
R22207 gnd.n4933 gnd.n2138 0.152939
R22208 gnd.n4934 gnd.n4933 0.152939
R22209 gnd.n4961 gnd.n4934 0.152939
R22210 gnd.n4961 gnd.n4960 0.152939
R22211 gnd.n4960 gnd.n4959 0.152939
R22212 gnd.n4959 gnd.n4935 0.152939
R22213 gnd.n4955 gnd.n4935 0.152939
R22214 gnd.n4955 gnd.n4954 0.152939
R22215 gnd.n4954 gnd.n4953 0.152939
R22216 gnd.n4953 gnd.n4939 0.152939
R22217 gnd.n4949 gnd.n4939 0.152939
R22218 gnd.n4949 gnd.n4948 0.152939
R22219 gnd.n4948 gnd.n4947 0.152939
R22220 gnd.n4947 gnd.n1307 0.152939
R22221 gnd.n6256 gnd.n1307 0.152939
R22222 gnd.n6256 gnd.n6255 0.152939
R22223 gnd.n6255 gnd.n6254 0.152939
R22224 gnd.n6254 gnd.n1308 0.152939
R22225 gnd.n6250 gnd.n1308 0.152939
R22226 gnd.n6250 gnd.n6249 0.152939
R22227 gnd.n6249 gnd.n6248 0.152939
R22228 gnd.n6248 gnd.n1313 0.152939
R22229 gnd.n6244 gnd.n1313 0.152939
R22230 gnd.n6244 gnd.n6243 0.152939
R22231 gnd.n6243 gnd.n6242 0.152939
R22232 gnd.n6242 gnd.n1318 0.152939
R22233 gnd.n6238 gnd.n1318 0.152939
R22234 gnd.n6238 gnd.n6237 0.152939
R22235 gnd.n6237 gnd.n6236 0.152939
R22236 gnd.n6236 gnd.n1323 0.152939
R22237 gnd.n6232 gnd.n1323 0.152939
R22238 gnd.n6232 gnd.n6231 0.152939
R22239 gnd.n6231 gnd.n6230 0.152939
R22240 gnd.n6230 gnd.n1328 0.152939
R22241 gnd.n6226 gnd.n1328 0.152939
R22242 gnd.n6226 gnd.n6225 0.152939
R22243 gnd.n6225 gnd.n6224 0.152939
R22244 gnd.n6224 gnd.n1333 0.152939
R22245 gnd.n6220 gnd.n1333 0.152939
R22246 gnd.n6220 gnd.n6219 0.152939
R22247 gnd.n6219 gnd.n6218 0.152939
R22248 gnd.n6218 gnd.n1338 0.152939
R22249 gnd.n6214 gnd.n1338 0.152939
R22250 gnd.n6214 gnd.n6213 0.152939
R22251 gnd.n6213 gnd.n6212 0.152939
R22252 gnd.n6212 gnd.n1343 0.152939
R22253 gnd.n6208 gnd.n1343 0.152939
R22254 gnd.n6208 gnd.n6207 0.152939
R22255 gnd.n6207 gnd.n6206 0.152939
R22256 gnd.n6206 gnd.n1348 0.152939
R22257 gnd.n6202 gnd.n1348 0.152939
R22258 gnd.n6202 gnd.n6201 0.152939
R22259 gnd.n6201 gnd.n6200 0.152939
R22260 gnd.n6200 gnd.n1353 0.152939
R22261 gnd.n6196 gnd.n1353 0.152939
R22262 gnd.n6196 gnd.n6195 0.152939
R22263 gnd.n6195 gnd.n6194 0.152939
R22264 gnd.n6194 gnd.n1358 0.152939
R22265 gnd.n6190 gnd.n1358 0.152939
R22266 gnd.n6190 gnd.n6189 0.152939
R22267 gnd.n6189 gnd.n6188 0.152939
R22268 gnd.n6188 gnd.n1363 0.152939
R22269 gnd.n6184 gnd.n1363 0.152939
R22270 gnd.n6184 gnd.n6183 0.152939
R22271 gnd.n6183 gnd.n6182 0.152939
R22272 gnd.n6182 gnd.n1368 0.152939
R22273 gnd.n6178 gnd.n1368 0.152939
R22274 gnd.n6178 gnd.n6177 0.152939
R22275 gnd.n6177 gnd.n6176 0.152939
R22276 gnd.n6176 gnd.n1373 0.152939
R22277 gnd.n6172 gnd.n1373 0.152939
R22278 gnd.n6172 gnd.n6171 0.152939
R22279 gnd.n6171 gnd.n6170 0.152939
R22280 gnd.n6170 gnd.n1378 0.152939
R22281 gnd.n6166 gnd.n1378 0.152939
R22282 gnd.n6166 gnd.n6165 0.152939
R22283 gnd.n6165 gnd.n6164 0.152939
R22284 gnd.n6164 gnd.n1383 0.152939
R22285 gnd.n6160 gnd.n1383 0.152939
R22286 gnd.n6160 gnd.n6159 0.152939
R22287 gnd.n6159 gnd.n6158 0.152939
R22288 gnd.n6158 gnd.n1388 0.152939
R22289 gnd.n6154 gnd.n1388 0.152939
R22290 gnd.n6154 gnd.n6153 0.152939
R22291 gnd.n6153 gnd.n6152 0.152939
R22292 gnd.n6152 gnd.n1393 0.152939
R22293 gnd.n4596 gnd.n4595 0.152939
R22294 gnd.n4595 gnd.n2503 0.152939
R22295 gnd.n4652 gnd.n2503 0.152939
R22296 gnd.n4653 gnd.n4652 0.152939
R22297 gnd.n4654 gnd.n4653 0.152939
R22298 gnd.n4654 gnd.n2498 0.152939
R22299 gnd.n4667 gnd.n2498 0.152939
R22300 gnd.n4668 gnd.n4667 0.152939
R22301 gnd.n4669 gnd.n4668 0.152939
R22302 gnd.n4669 gnd.n2490 0.152939
R22303 gnd.n4705 gnd.n2490 0.152939
R22304 gnd.n4705 gnd.n4704 0.152939
R22305 gnd.n4704 gnd.n4703 0.152939
R22306 gnd.n4703 gnd.n2491 0.152939
R22307 gnd.n4699 gnd.n2491 0.152939
R22308 gnd.n4699 gnd.n4698 0.152939
R22309 gnd.n4698 gnd.n4697 0.152939
R22310 gnd.n4697 gnd.n2495 0.152939
R22311 gnd.n4693 gnd.n2495 0.152939
R22312 gnd.n4693 gnd.n2471 0.152939
R22313 gnd.n4765 gnd.n2471 0.152939
R22314 gnd.n4766 gnd.n4765 0.152939
R22315 gnd.n4768 gnd.n4766 0.152939
R22316 gnd.n4768 gnd.n4767 0.152939
R22317 gnd.n4767 gnd.n2465 0.152939
R22318 gnd.n4782 gnd.n2465 0.152939
R22319 gnd.n4852 gnd.n2270 0.152939
R22320 gnd.n4852 gnd.n4851 0.152939
R22321 gnd.n4851 gnd.n4850 0.152939
R22322 gnd.n4850 gnd.n2272 0.152939
R22323 gnd.n4846 gnd.n2272 0.152939
R22324 gnd.n4846 gnd.n4845 0.152939
R22325 gnd.n2269 gnd.n2219 0.152939
R22326 gnd.n2265 gnd.n2219 0.152939
R22327 gnd.n2265 gnd.n2264 0.152939
R22328 gnd.n2264 gnd.n2263 0.152939
R22329 gnd.n2263 gnd.n2223 0.152939
R22330 gnd.n2259 gnd.n2223 0.152939
R22331 gnd.n2259 gnd.n2258 0.152939
R22332 gnd.n2258 gnd.n2257 0.152939
R22333 gnd.n2257 gnd.n2227 0.152939
R22334 gnd.n2253 gnd.n2227 0.152939
R22335 gnd.n2253 gnd.n2252 0.152939
R22336 gnd.n2252 gnd.n2251 0.152939
R22337 gnd.n2251 gnd.n2231 0.152939
R22338 gnd.n2247 gnd.n2231 0.152939
R22339 gnd.n2247 gnd.n2246 0.152939
R22340 gnd.n2246 gnd.n2245 0.152939
R22341 gnd.n2245 gnd.n2235 0.152939
R22342 gnd.n2241 gnd.n2235 0.152939
R22343 gnd.n2241 gnd.n2240 0.152939
R22344 gnd.n2240 gnd.n2239 0.152939
R22345 gnd.n2239 gnd.n2238 0.152939
R22346 gnd.n2238 gnd.n2120 0.152939
R22347 gnd.n4981 gnd.n2120 0.152939
R22348 gnd.n4982 gnd.n4981 0.152939
R22349 gnd.n4983 gnd.n4982 0.152939
R22350 gnd.n4983 gnd.n2118 0.152939
R22351 gnd.n4989 gnd.n2118 0.152939
R22352 gnd.n4990 gnd.n4989 0.152939
R22353 gnd.n5007 gnd.n4990 0.152939
R22354 gnd.n5007 gnd.n5006 0.152939
R22355 gnd.n5006 gnd.n5005 0.152939
R22356 gnd.n5005 gnd.n4991 0.152939
R22357 gnd.n5001 gnd.n4991 0.152939
R22358 gnd.n5001 gnd.n5000 0.152939
R22359 gnd.n5000 gnd.n4999 0.152939
R22360 gnd.n4999 gnd.n4995 0.152939
R22361 gnd.n4995 gnd.n2068 0.152939
R22362 gnd.n5108 gnd.n2068 0.152939
R22363 gnd.n5109 gnd.n5108 0.152939
R22364 gnd.n5111 gnd.n5109 0.152939
R22365 gnd.n5111 gnd.n5110 0.152939
R22366 gnd.n5110 gnd.n2043 0.152939
R22367 gnd.n5140 gnd.n2043 0.152939
R22368 gnd.n5141 gnd.n5140 0.152939
R22369 gnd.n5166 gnd.n5141 0.152939
R22370 gnd.n5166 gnd.n5165 0.152939
R22371 gnd.n5165 gnd.n5164 0.152939
R22372 gnd.n5164 gnd.n5142 0.152939
R22373 gnd.n5160 gnd.n5142 0.152939
R22374 gnd.n5160 gnd.n5159 0.152939
R22375 gnd.n5159 gnd.n5158 0.152939
R22376 gnd.n5158 gnd.n5147 0.152939
R22377 gnd.n5154 gnd.n5147 0.152939
R22378 gnd.n5154 gnd.n5153 0.152939
R22379 gnd.n5153 gnd.n5152 0.152939
R22380 gnd.n5152 gnd.n1967 0.152939
R22381 gnd.n5265 gnd.n1967 0.152939
R22382 gnd.n5266 gnd.n5265 0.152939
R22383 gnd.n5297 gnd.n5266 0.152939
R22384 gnd.n5297 gnd.n5296 0.152939
R22385 gnd.n5296 gnd.n5295 0.152939
R22386 gnd.n5295 gnd.n5267 0.152939
R22387 gnd.n5291 gnd.n5267 0.152939
R22388 gnd.n5291 gnd.n5290 0.152939
R22389 gnd.n5290 gnd.n5289 0.152939
R22390 gnd.n5289 gnd.n5273 0.152939
R22391 gnd.n5285 gnd.n5273 0.152939
R22392 gnd.n5285 gnd.n5284 0.152939
R22393 gnd.n5284 gnd.n5283 0.152939
R22394 gnd.n5283 gnd.n5276 0.152939
R22395 gnd.n5276 gnd.n1896 0.152939
R22396 gnd.n5417 gnd.n1896 0.152939
R22397 gnd.n5418 gnd.n5417 0.152939
R22398 gnd.n5430 gnd.n5418 0.152939
R22399 gnd.n5430 gnd.n5429 0.152939
R22400 gnd.n5429 gnd.n5428 0.152939
R22401 gnd.n5428 gnd.n5419 0.152939
R22402 gnd.n5424 gnd.n5419 0.152939
R22403 gnd.n5424 gnd.n5423 0.152939
R22404 gnd.n5423 gnd.n1822 0.152939
R22405 gnd.n5628 gnd.n1822 0.152939
R22406 gnd.n5629 gnd.n5628 0.152939
R22407 gnd.n5630 gnd.n5629 0.152939
R22408 gnd.n5630 gnd.n1810 0.152939
R22409 gnd.n5645 gnd.n1810 0.152939
R22410 gnd.n5646 gnd.n5645 0.152939
R22411 gnd.n5647 gnd.n5646 0.152939
R22412 gnd.n5647 gnd.n1798 0.152939
R22413 gnd.n5662 gnd.n1798 0.152939
R22414 gnd.n5663 gnd.n5662 0.152939
R22415 gnd.n5664 gnd.n5663 0.152939
R22416 gnd.n5664 gnd.n1785 0.152939
R22417 gnd.n5679 gnd.n1785 0.152939
R22418 gnd.n5680 gnd.n5679 0.152939
R22419 gnd.n5681 gnd.n5680 0.152939
R22420 gnd.n5681 gnd.n1774 0.152939
R22421 gnd.n5699 gnd.n1774 0.152939
R22422 gnd.n5700 gnd.n5699 0.152939
R22423 gnd.n5701 gnd.n5700 0.152939
R22424 gnd.n5701 gnd.n1402 0.152939
R22425 gnd.n6145 gnd.n1402 0.152939
R22426 gnd.n6144 gnd.n1403 0.152939
R22427 gnd.n6140 gnd.n1403 0.152939
R22428 gnd.n6140 gnd.n6139 0.152939
R22429 gnd.n6139 gnd.n6138 0.152939
R22430 gnd.n6138 gnd.n1407 0.152939
R22431 gnd.n6134 gnd.n1407 0.152939
R22432 gnd.n5772 gnd.n5734 0.152939
R22433 gnd.n5772 gnd.n5771 0.152939
R22434 gnd.n5771 gnd.n5770 0.152939
R22435 gnd.n5770 gnd.n5735 0.152939
R22436 gnd.n5766 gnd.n5735 0.152939
R22437 gnd.n5766 gnd.n5765 0.152939
R22438 gnd.n5765 gnd.n5764 0.152939
R22439 gnd.n5764 gnd.n5740 0.152939
R22440 gnd.n5760 gnd.n5740 0.152939
R22441 gnd.n5760 gnd.n1718 0.152939
R22442 gnd.n5824 gnd.n1718 0.152939
R22443 gnd.n5825 gnd.n5824 0.152939
R22444 gnd.n5826 gnd.n5825 0.152939
R22445 gnd.n5826 gnd.n1713 0.152939
R22446 gnd.n5839 gnd.n1713 0.152939
R22447 gnd.n5840 gnd.n5839 0.152939
R22448 gnd.n5841 gnd.n5840 0.152939
R22449 gnd.n5841 gnd.n1709 0.152939
R22450 gnd.n5871 gnd.n1709 0.152939
R22451 gnd.n5871 gnd.n5870 0.152939
R22452 gnd.n5870 gnd.n5869 0.152939
R22453 gnd.n5869 gnd.n1710 0.152939
R22454 gnd.n5865 gnd.n1710 0.152939
R22455 gnd.n5865 gnd.n5864 0.152939
R22456 gnd.n5864 gnd.n5863 0.152939
R22457 gnd.n5863 gnd.n83 0.152939
R22458 gnd.n4845 gnd.n4844 0.128549
R22459 gnd.n6134 gnd.n6133 0.128549
R22460 gnd.n5882 gnd.n98 0.098061
R22461 gnd.n4623 gnd.n948 0.098061
R22462 gnd.n3524 gnd.n3523 0.0767195
R22463 gnd.n3523 gnd.n3522 0.0767195
R22464 gnd.n7618 gnd.n96 0.0767195
R22465 gnd.n7618 gnd.n97 0.0767195
R22466 gnd.n6479 gnd.n946 0.0767195
R22467 gnd.n6479 gnd.n947 0.0767195
R22468 gnd.n7628 gnd.n7627 0.0695946
R22469 gnd.n4594 gnd.n4591 0.0695946
R22470 gnd.n4596 gnd.n4594 0.0695946
R22471 gnd.n7628 gnd.n83 0.0695946
R22472 gnd.n4844 gnd.n2389 0.063
R22473 gnd.n6133 gnd.n1412 0.063
R22474 gnd.n390 gnd.n98 0.055378
R22475 gnd.n2513 gnd.n948 0.055378
R22476 gnd.n4091 gnd.n2690 0.0477147
R22477 gnd.n1580 gnd.n1412 0.0477147
R22478 gnd.n7436 gnd.n207 0.0477147
R22479 gnd.n4323 gnd.n2643 0.0477147
R22480 gnd.n2389 gnd.n1063 0.0477147
R22481 gnd.n3287 gnd.n3175 0.0442063
R22482 gnd.n3288 gnd.n3287 0.0442063
R22483 gnd.n3289 gnd.n3288 0.0442063
R22484 gnd.n3289 gnd.n3164 0.0442063
R22485 gnd.n3303 gnd.n3164 0.0442063
R22486 gnd.n3304 gnd.n3303 0.0442063
R22487 gnd.n3305 gnd.n3304 0.0442063
R22488 gnd.n3305 gnd.n3151 0.0442063
R22489 gnd.n3349 gnd.n3151 0.0442063
R22490 gnd.n3350 gnd.n3349 0.0442063
R22491 gnd.n3352 gnd.n3085 0.0344674
R22492 gnd.n5955 gnd.n1580 0.0344674
R22493 gnd.n5955 gnd.n1582 0.0344674
R22494 gnd.n1606 gnd.n1582 0.0344674
R22495 gnd.n1607 gnd.n1606 0.0344674
R22496 gnd.n1608 gnd.n1607 0.0344674
R22497 gnd.n1609 gnd.n1608 0.0344674
R22498 gnd.n5747 gnd.n1609 0.0344674
R22499 gnd.n5747 gnd.n1627 0.0344674
R22500 gnd.n1628 gnd.n1627 0.0344674
R22501 gnd.n1629 gnd.n1628 0.0344674
R22502 gnd.n5753 gnd.n1629 0.0344674
R22503 gnd.n5753 gnd.n1647 0.0344674
R22504 gnd.n1648 gnd.n1647 0.0344674
R22505 gnd.n1649 gnd.n1648 0.0344674
R22506 gnd.n5833 gnd.n1649 0.0344674
R22507 gnd.n5833 gnd.n1667 0.0344674
R22508 gnd.n1668 gnd.n1667 0.0344674
R22509 gnd.n1669 gnd.n1668 0.0344674
R22510 gnd.n5848 gnd.n1669 0.0344674
R22511 gnd.n5848 gnd.n1687 0.0344674
R22512 gnd.n1688 gnd.n1687 0.0344674
R22513 gnd.n1689 gnd.n1688 0.0344674
R22514 gnd.n5851 gnd.n1689 0.0344674
R22515 gnd.n5851 gnd.n378 0.0344674
R22516 gnd.n7302 gnd.n378 0.0344674
R22517 gnd.n7303 gnd.n7302 0.0344674
R22518 gnd.n7303 gnd.n373 0.0344674
R22519 gnd.n373 gnd.n371 0.0344674
R22520 gnd.n7314 gnd.n371 0.0344674
R22521 gnd.n7315 gnd.n7314 0.0344674
R22522 gnd.n7315 gnd.n111 0.0344674
R22523 gnd.n112 gnd.n111 0.0344674
R22524 gnd.n113 gnd.n112 0.0344674
R22525 gnd.n7316 gnd.n113 0.0344674
R22526 gnd.n7316 gnd.n128 0.0344674
R22527 gnd.n129 gnd.n128 0.0344674
R22528 gnd.n130 gnd.n129 0.0344674
R22529 gnd.n7317 gnd.n130 0.0344674
R22530 gnd.n7317 gnd.n148 0.0344674
R22531 gnd.n149 gnd.n148 0.0344674
R22532 gnd.n150 gnd.n149 0.0344674
R22533 gnd.n7318 gnd.n150 0.0344674
R22534 gnd.n7318 gnd.n166 0.0344674
R22535 gnd.n167 gnd.n166 0.0344674
R22536 gnd.n168 gnd.n167 0.0344674
R22537 gnd.n7319 gnd.n168 0.0344674
R22538 gnd.n7319 gnd.n186 0.0344674
R22539 gnd.n187 gnd.n186 0.0344674
R22540 gnd.n188 gnd.n187 0.0344674
R22541 gnd.n7320 gnd.n188 0.0344674
R22542 gnd.n7320 gnd.n205 0.0344674
R22543 gnd.n206 gnd.n205 0.0344674
R22544 gnd.n207 gnd.n206 0.0344674
R22545 gnd.n4448 gnd.n2643 0.0344674
R22546 gnd.n4448 gnd.n2646 0.0344674
R22547 gnd.n2646 gnd.n2645 0.0344674
R22548 gnd.n2645 gnd.n2626 0.0344674
R22549 gnd.n2626 gnd.n2624 0.0344674
R22550 gnd.n4465 gnd.n2624 0.0344674
R22551 gnd.n4466 gnd.n4465 0.0344674
R22552 gnd.n4466 gnd.n2608 0.0344674
R22553 gnd.n2608 gnd.n2606 0.0344674
R22554 gnd.n4485 gnd.n2606 0.0344674
R22555 gnd.n4486 gnd.n4485 0.0344674
R22556 gnd.n4486 gnd.n2590 0.0344674
R22557 gnd.n2590 gnd.n2587 0.0344674
R22558 gnd.n2588 gnd.n2587 0.0344674
R22559 gnd.n4507 gnd.n2588 0.0344674
R22560 gnd.n4508 gnd.n4507 0.0344674
R22561 gnd.n4508 gnd.n2564 0.0344674
R22562 gnd.n2564 gnd.n2562 0.0344674
R22563 gnd.n4550 gnd.n2562 0.0344674
R22564 gnd.n4551 gnd.n4550 0.0344674
R22565 gnd.n4551 gnd.n2547 0.0344674
R22566 gnd.n2547 gnd.n2544 0.0344674
R22567 gnd.n2545 gnd.n2544 0.0344674
R22568 gnd.n4573 gnd.n2545 0.0344674
R22569 gnd.n4574 gnd.n4573 0.0344674
R22570 gnd.n4574 gnd.n2531 0.0344674
R22571 gnd.n2531 gnd.n2527 0.0344674
R22572 gnd.n2528 gnd.n2527 0.0344674
R22573 gnd.n4608 gnd.n2528 0.0344674
R22574 gnd.n4608 gnd.n2529 0.0344674
R22575 gnd.n2529 gnd.n962 0.0344674
R22576 gnd.n963 gnd.n962 0.0344674
R22577 gnd.n964 gnd.n963 0.0344674
R22578 gnd.n4661 gnd.n964 0.0344674
R22579 gnd.n4661 gnd.n981 0.0344674
R22580 gnd.n982 gnd.n981 0.0344674
R22581 gnd.n983 gnd.n982 0.0344674
R22582 gnd.n4676 gnd.n983 0.0344674
R22583 gnd.n4676 gnd.n1001 0.0344674
R22584 gnd.n1002 gnd.n1001 0.0344674
R22585 gnd.n1003 gnd.n1002 0.0344674
R22586 gnd.n4683 gnd.n1003 0.0344674
R22587 gnd.n4683 gnd.n1021 0.0344674
R22588 gnd.n1022 gnd.n1021 0.0344674
R22589 gnd.n1023 gnd.n1022 0.0344674
R22590 gnd.n2474 gnd.n1023 0.0344674
R22591 gnd.n2474 gnd.n1041 0.0344674
R22592 gnd.n1042 gnd.n1041 0.0344674
R22593 gnd.n1043 gnd.n1042 0.0344674
R22594 gnd.n2469 gnd.n1043 0.0344674
R22595 gnd.n2469 gnd.n1061 0.0344674
R22596 gnd.n1062 gnd.n1061 0.0344674
R22597 gnd.n1063 gnd.n1062 0.0344674
R22598 gnd.n4843 gnd.n2390 0.0343753
R22599 gnd.n6132 gnd.n6131 0.0343753
R22600 gnd.n4791 gnd.n4783 0.0296328
R22601 gnd.n5733 gnd.n5732 0.0296328
R22602 gnd.n3372 gnd.n3371 0.0269946
R22603 gnd.n3374 gnd.n3373 0.0269946
R22604 gnd.n3080 gnd.n3078 0.0269946
R22605 gnd.n3384 gnd.n3382 0.0269946
R22606 gnd.n3383 gnd.n3059 0.0269946
R22607 gnd.n3403 gnd.n3402 0.0269946
R22608 gnd.n3405 gnd.n3404 0.0269946
R22609 gnd.n3054 gnd.n3053 0.0269946
R22610 gnd.n3415 gnd.n3049 0.0269946
R22611 gnd.n3414 gnd.n3051 0.0269946
R22612 gnd.n3050 gnd.n3032 0.0269946
R22613 gnd.n3435 gnd.n3033 0.0269946
R22614 gnd.n3434 gnd.n3034 0.0269946
R22615 gnd.n3468 gnd.n3009 0.0269946
R22616 gnd.n3470 gnd.n3469 0.0269946
R22617 gnd.n3471 gnd.n2956 0.0269946
R22618 gnd.n3004 gnd.n2957 0.0269946
R22619 gnd.n3006 gnd.n2958 0.0269946
R22620 gnd.n3481 gnd.n3480 0.0269946
R22621 gnd.n3483 gnd.n3482 0.0269946
R22622 gnd.n3484 gnd.n2978 0.0269946
R22623 gnd.n3486 gnd.n2979 0.0269946
R22624 gnd.n3489 gnd.n2980 0.0269946
R22625 gnd.n3492 gnd.n3491 0.0269946
R22626 gnd.n3494 gnd.n3493 0.0269946
R22627 gnd.n3559 gnd.n2863 0.0269946
R22628 gnd.n3561 gnd.n3560 0.0269946
R22629 gnd.n3570 gnd.n2856 0.0269946
R22630 gnd.n3572 gnd.n3571 0.0269946
R22631 gnd.n3573 gnd.n2854 0.0269946
R22632 gnd.n3580 gnd.n3576 0.0269946
R22633 gnd.n3579 gnd.n3578 0.0269946
R22634 gnd.n3577 gnd.n2833 0.0269946
R22635 gnd.n3602 gnd.n2834 0.0269946
R22636 gnd.n3601 gnd.n2835 0.0269946
R22637 gnd.n3644 gnd.n2808 0.0269946
R22638 gnd.n3646 gnd.n3645 0.0269946
R22639 gnd.n3655 gnd.n2801 0.0269946
R22640 gnd.n3657 gnd.n3656 0.0269946
R22641 gnd.n3658 gnd.n2799 0.0269946
R22642 gnd.n3665 gnd.n3661 0.0269946
R22643 gnd.n3664 gnd.n3663 0.0269946
R22644 gnd.n3662 gnd.n2778 0.0269946
R22645 gnd.n3687 gnd.n2779 0.0269946
R22646 gnd.n3686 gnd.n2780 0.0269946
R22647 gnd.n3733 gnd.n2754 0.0269946
R22648 gnd.n3735 gnd.n3734 0.0269946
R22649 gnd.n3745 gnd.n2747 0.0269946
R22650 gnd.n4004 gnd.n2745 0.0269946
R22651 gnd.n4009 gnd.n4007 0.0269946
R22652 gnd.n4008 gnd.n2726 0.0269946
R22653 gnd.n4033 gnd.n4032 0.0269946
R22654 gnd.n4839 gnd.n2396 0.022519
R22655 gnd.n4838 gnd.n2397 0.022519
R22656 gnd.n4835 gnd.n4834 0.022519
R22657 gnd.n4831 gnd.n2403 0.022519
R22658 gnd.n4830 gnd.n2409 0.022519
R22659 gnd.n4827 gnd.n4826 0.022519
R22660 gnd.n4823 gnd.n2415 0.022519
R22661 gnd.n4822 gnd.n2419 0.022519
R22662 gnd.n4819 gnd.n4818 0.022519
R22663 gnd.n4815 gnd.n2426 0.022519
R22664 gnd.n4814 gnd.n2432 0.022519
R22665 gnd.n4811 gnd.n4810 0.022519
R22666 gnd.n4807 gnd.n2438 0.022519
R22667 gnd.n4806 gnd.n2442 0.022519
R22668 gnd.n4803 gnd.n4802 0.022519
R22669 gnd.n4799 gnd.n2449 0.022519
R22670 gnd.n4798 gnd.n2456 0.022519
R22671 gnd.n2464 gnd.n2462 0.022519
R22672 gnd.n4792 gnd.n4791 0.022519
R22673 gnd.n6128 gnd.n1413 0.022519
R22674 gnd.n6127 gnd.n1417 0.022519
R22675 gnd.n6124 gnd.n6123 0.022519
R22676 gnd.n6120 gnd.n1422 0.022519
R22677 gnd.n6119 gnd.n1426 0.022519
R22678 gnd.n6116 gnd.n6115 0.022519
R22679 gnd.n6112 gnd.n1430 0.022519
R22680 gnd.n6111 gnd.n1434 0.022519
R22681 gnd.n6108 gnd.n6107 0.022519
R22682 gnd.n6104 gnd.n1438 0.022519
R22683 gnd.n6103 gnd.n1442 0.022519
R22684 gnd.n6100 gnd.n6099 0.022519
R22685 gnd.n6096 gnd.n1446 0.022519
R22686 gnd.n6095 gnd.n1450 0.022519
R22687 gnd.n6092 gnd.n6091 0.022519
R22688 gnd.n6088 gnd.n1454 0.022519
R22689 gnd.n6087 gnd.n1460 0.022519
R22690 gnd.n1739 gnd.n1463 0.022519
R22691 gnd.n5732 gnd.n1738 0.022519
R22692 gnd.n5733 gnd.n1737 0.0218415
R22693 gnd.n4783 gnd.n2193 0.0218415
R22694 gnd.n3352 gnd.n3351 0.0202011
R22695 gnd.n3351 gnd.n3350 0.0148637
R22696 gnd.n4002 gnd.n3746 0.0144266
R22697 gnd.n4003 gnd.n4002 0.0130679
R22698 gnd.n2396 gnd.n2390 0.0123564
R22699 gnd.n4839 gnd.n4838 0.0123564
R22700 gnd.n4835 gnd.n2397 0.0123564
R22701 gnd.n4834 gnd.n2403 0.0123564
R22702 gnd.n4831 gnd.n4830 0.0123564
R22703 gnd.n4827 gnd.n2409 0.0123564
R22704 gnd.n4826 gnd.n2415 0.0123564
R22705 gnd.n4823 gnd.n4822 0.0123564
R22706 gnd.n4819 gnd.n2419 0.0123564
R22707 gnd.n4818 gnd.n2426 0.0123564
R22708 gnd.n4815 gnd.n4814 0.0123564
R22709 gnd.n4811 gnd.n2432 0.0123564
R22710 gnd.n4810 gnd.n2438 0.0123564
R22711 gnd.n4807 gnd.n4806 0.0123564
R22712 gnd.n4803 gnd.n2442 0.0123564
R22713 gnd.n4802 gnd.n2449 0.0123564
R22714 gnd.n4799 gnd.n4798 0.0123564
R22715 gnd.n2462 gnd.n2456 0.0123564
R22716 gnd.n4792 gnd.n2464 0.0123564
R22717 gnd.n6131 gnd.n1413 0.0123564
R22718 gnd.n6128 gnd.n6127 0.0123564
R22719 gnd.n6124 gnd.n1417 0.0123564
R22720 gnd.n6123 gnd.n1422 0.0123564
R22721 gnd.n6120 gnd.n6119 0.0123564
R22722 gnd.n6116 gnd.n1426 0.0123564
R22723 gnd.n6115 gnd.n1430 0.0123564
R22724 gnd.n6112 gnd.n6111 0.0123564
R22725 gnd.n6108 gnd.n1434 0.0123564
R22726 gnd.n6107 gnd.n1438 0.0123564
R22727 gnd.n6104 gnd.n6103 0.0123564
R22728 gnd.n6100 gnd.n1442 0.0123564
R22729 gnd.n6099 gnd.n1446 0.0123564
R22730 gnd.n6096 gnd.n6095 0.0123564
R22731 gnd.n6092 gnd.n1450 0.0123564
R22732 gnd.n6091 gnd.n1454 0.0123564
R22733 gnd.n6088 gnd.n6087 0.0123564
R22734 gnd.n1463 gnd.n1460 0.0123564
R22735 gnd.n1739 gnd.n1738 0.0123564
R22736 gnd.n3371 gnd.n3085 0.00797283
R22737 gnd.n3373 gnd.n3372 0.00797283
R22738 gnd.n3374 gnd.n3080 0.00797283
R22739 gnd.n3382 gnd.n3078 0.00797283
R22740 gnd.n3384 gnd.n3383 0.00797283
R22741 gnd.n3402 gnd.n3059 0.00797283
R22742 gnd.n3404 gnd.n3403 0.00797283
R22743 gnd.n3405 gnd.n3054 0.00797283
R22744 gnd.n3053 gnd.n3049 0.00797283
R22745 gnd.n3415 gnd.n3414 0.00797283
R22746 gnd.n3051 gnd.n3050 0.00797283
R22747 gnd.n3033 gnd.n3032 0.00797283
R22748 gnd.n3435 gnd.n3434 0.00797283
R22749 gnd.n3034 gnd.n3009 0.00797283
R22750 gnd.n3469 gnd.n3468 0.00797283
R22751 gnd.n3471 gnd.n3470 0.00797283
R22752 gnd.n3004 gnd.n2956 0.00797283
R22753 gnd.n3006 gnd.n2957 0.00797283
R22754 gnd.n3480 gnd.n2958 0.00797283
R22755 gnd.n3482 gnd.n3481 0.00797283
R22756 gnd.n3484 gnd.n3483 0.00797283
R22757 gnd.n3486 gnd.n2978 0.00797283
R22758 gnd.n3489 gnd.n2979 0.00797283
R22759 gnd.n3491 gnd.n2980 0.00797283
R22760 gnd.n3494 gnd.n3492 0.00797283
R22761 gnd.n3493 gnd.n2863 0.00797283
R22762 gnd.n3561 gnd.n3559 0.00797283
R22763 gnd.n3560 gnd.n2856 0.00797283
R22764 gnd.n3571 gnd.n3570 0.00797283
R22765 gnd.n3573 gnd.n3572 0.00797283
R22766 gnd.n3576 gnd.n2854 0.00797283
R22767 gnd.n3580 gnd.n3579 0.00797283
R22768 gnd.n3578 gnd.n3577 0.00797283
R22769 gnd.n2834 gnd.n2833 0.00797283
R22770 gnd.n3602 gnd.n3601 0.00797283
R22771 gnd.n2835 gnd.n2808 0.00797283
R22772 gnd.n3646 gnd.n3644 0.00797283
R22773 gnd.n3645 gnd.n2801 0.00797283
R22774 gnd.n3656 gnd.n3655 0.00797283
R22775 gnd.n3658 gnd.n3657 0.00797283
R22776 gnd.n3661 gnd.n2799 0.00797283
R22777 gnd.n3665 gnd.n3664 0.00797283
R22778 gnd.n3663 gnd.n3662 0.00797283
R22779 gnd.n2779 gnd.n2778 0.00797283
R22780 gnd.n3687 gnd.n3686 0.00797283
R22781 gnd.n2780 gnd.n2754 0.00797283
R22782 gnd.n3735 gnd.n3733 0.00797283
R22783 gnd.n3734 gnd.n2747 0.00797283
R22784 gnd.n3746 gnd.n3745 0.00797283
R22785 gnd.n4004 gnd.n4003 0.00797283
R22786 gnd.n4007 gnd.n2745 0.00797283
R22787 gnd.n4009 gnd.n4008 0.00797283
R22788 gnd.n4032 gnd.n2726 0.00797283
R22789 gnd.n4033 gnd.n2690 0.00797283
R22790 gnd.n4844 gnd.n4843 0.00592005
R22791 gnd.n6133 gnd.n6132 0.00592005
R22792 plus.n43 plus.t18 322.512
R22793 plus.n9 plus.t13 322.512
R22794 plus.n42 plus.t17 297.12
R22795 plus.n46 plus.t22 297.12
R22796 plus.n48 plus.t21 297.12
R22797 plus.n52 plus.t23 297.12
R22798 plus.n54 plus.t8 297.12
R22799 plus.n58 plus.t7 297.12
R22800 plus.n60 plus.t12 297.12
R22801 plus.n64 plus.t10 297.12
R22802 plus.n66 plus.t24 297.12
R22803 plus.n32 plus.t14 297.12
R22804 plus.n30 plus.t15 297.12
R22805 plus.n2 plus.t9 297.12
R22806 plus.n24 plus.t5 297.12
R22807 plus.n4 plus.t6 297.12
R22808 plus.n18 plus.t19 297.12
R22809 plus.n6 plus.t20 297.12
R22810 plus.n12 plus.t16 297.12
R22811 plus.n8 plus.t11 297.12
R22812 plus.n70 plus.t0 243.97
R22813 plus.n70 plus.n69 223.454
R22814 plus.n72 plus.n71 223.454
R22815 plus.n67 plus.n66 161.3
R22816 plus.n65 plus.n34 161.3
R22817 plus.n64 plus.n63 161.3
R22818 plus.n62 plus.n35 161.3
R22819 plus.n61 plus.n60 161.3
R22820 plus.n59 plus.n36 161.3
R22821 plus.n58 plus.n57 161.3
R22822 plus.n56 plus.n37 161.3
R22823 plus.n55 plus.n54 161.3
R22824 plus.n53 plus.n38 161.3
R22825 plus.n52 plus.n51 161.3
R22826 plus.n50 plus.n39 161.3
R22827 plus.n49 plus.n48 161.3
R22828 plus.n47 plus.n40 161.3
R22829 plus.n46 plus.n45 161.3
R22830 plus.n44 plus.n41 161.3
R22831 plus.n11 plus.n10 161.3
R22832 plus.n12 plus.n7 161.3
R22833 plus.n14 plus.n13 161.3
R22834 plus.n15 plus.n6 161.3
R22835 plus.n17 plus.n16 161.3
R22836 plus.n18 plus.n5 161.3
R22837 plus.n20 plus.n19 161.3
R22838 plus.n21 plus.n4 161.3
R22839 plus.n23 plus.n22 161.3
R22840 plus.n24 plus.n3 161.3
R22841 plus.n26 plus.n25 161.3
R22842 plus.n27 plus.n2 161.3
R22843 plus.n29 plus.n28 161.3
R22844 plus.n30 plus.n1 161.3
R22845 plus.n31 plus.n0 161.3
R22846 plus.n33 plus.n32 161.3
R22847 plus.n44 plus.n43 45.0031
R22848 plus.n10 plus.n9 45.0031
R22849 plus.n66 plus.n65 41.6278
R22850 plus.n32 plus.n31 41.6278
R22851 plus.n42 plus.n41 37.246
R22852 plus.n64 plus.n35 37.246
R22853 plus.n30 plus.n29 37.246
R22854 plus.n11 plus.n8 37.246
R22855 plus.n47 plus.n46 32.8641
R22856 plus.n60 plus.n59 32.8641
R22857 plus.n25 plus.n2 32.8641
R22858 plus.n13 plus.n12 32.8641
R22859 plus.n68 plus.n67 31.6047
R22860 plus.n48 plus.n39 28.4823
R22861 plus.n58 plus.n37 28.4823
R22862 plus.n24 plus.n23 28.4823
R22863 plus.n17 plus.n6 28.4823
R22864 plus.n53 plus.n52 24.1005
R22865 plus.n54 plus.n53 24.1005
R22866 plus.n19 plus.n4 24.1005
R22867 plus.n19 plus.n18 24.1005
R22868 plus.n69 plus.t4 19.8005
R22869 plus.n69 plus.t2 19.8005
R22870 plus.n71 plus.t1 19.8005
R22871 plus.n71 plus.t3 19.8005
R22872 plus.n52 plus.n39 19.7187
R22873 plus.n54 plus.n37 19.7187
R22874 plus.n23 plus.n4 19.7187
R22875 plus.n18 plus.n17 19.7187
R22876 plus.n43 plus.n42 15.6319
R22877 plus.n9 plus.n8 15.6319
R22878 plus.n48 plus.n47 15.3369
R22879 plus.n59 plus.n58 15.3369
R22880 plus.n25 plus.n24 15.3369
R22881 plus.n13 plus.n6 15.3369
R22882 plus plus.n73 14.734
R22883 plus.n68 plus.n33 11.866
R22884 plus.n46 plus.n41 10.955
R22885 plus.n60 plus.n35 10.955
R22886 plus.n29 plus.n2 10.955
R22887 plus.n12 plus.n11 10.955
R22888 plus.n65 plus.n64 6.57323
R22889 plus.n31 plus.n30 6.57323
R22890 plus.n73 plus.n72 5.40567
R22891 plus.n73 plus.n68 1.188
R22892 plus.n72 plus.n70 0.716017
R22893 plus.n45 plus.n44 0.189894
R22894 plus.n45 plus.n40 0.189894
R22895 plus.n49 plus.n40 0.189894
R22896 plus.n50 plus.n49 0.189894
R22897 plus.n51 plus.n50 0.189894
R22898 plus.n51 plus.n38 0.189894
R22899 plus.n55 plus.n38 0.189894
R22900 plus.n56 plus.n55 0.189894
R22901 plus.n57 plus.n56 0.189894
R22902 plus.n57 plus.n36 0.189894
R22903 plus.n61 plus.n36 0.189894
R22904 plus.n62 plus.n61 0.189894
R22905 plus.n63 plus.n62 0.189894
R22906 plus.n63 plus.n34 0.189894
R22907 plus.n67 plus.n34 0.189894
R22908 plus.n33 plus.n0 0.189894
R22909 plus.n1 plus.n0 0.189894
R22910 plus.n28 plus.n1 0.189894
R22911 plus.n28 plus.n27 0.189894
R22912 plus.n27 plus.n26 0.189894
R22913 plus.n26 plus.n3 0.189894
R22914 plus.n22 plus.n3 0.189894
R22915 plus.n22 plus.n21 0.189894
R22916 plus.n21 plus.n20 0.189894
R22917 plus.n20 plus.n5 0.189894
R22918 plus.n16 plus.n5 0.189894
R22919 plus.n16 plus.n15 0.189894
R22920 plus.n15 plus.n14 0.189894
R22921 plus.n14 plus.n7 0.189894
R22922 plus.n10 plus.n7 0.189894
R22923 a_n3827_n3924.n32 a_n3827_n3924.t48 214.994
R22924 a_n3827_n3924.n24 a_n3827_n3924.t0 214.994
R22925 a_n3827_n3924.n32 a_n3827_n3924.t44 214.321
R22926 a_n3827_n3924.n31 a_n3827_n3924.t49 214.321
R22927 a_n3827_n3924.n30 a_n3827_n3924.t39 214.321
R22928 a_n3827_n3924.n29 a_n3827_n3924.t27 214.321
R22929 a_n3827_n3924.n28 a_n3827_n3924.t40 214.321
R22930 a_n3827_n3924.n27 a_n3827_n3924.t24 214.321
R22931 a_n3827_n3924.n26 a_n3827_n3924.t25 214.321
R22932 a_n3827_n3924.n24 a_n3827_n3924.t36 214.321
R22933 a_n3827_n3924.n11 a_n3827_n3924.t8 55.8337
R22934 a_n3827_n3924.n12 a_n3827_n3924.t29 55.8337
R22935 a_n3827_n3924.n21 a_n3827_n3924.t32 55.8337
R22936 a_n3827_n3924.n2 a_n3827_n3924.t2 55.8335
R22937 a_n3827_n3924.n35 a_n3827_n3924.t37 55.8335
R22938 a_n3827_n3924.n44 a_n3827_n3924.t42 55.8335
R22939 a_n3827_n3924.n45 a_n3827_n3924.t13 55.8335
R22940 a_n3827_n3924.n22 a_n3827_n3924.t12 55.8335
R22941 a_n3827_n3924.n51 a_n3827_n3924.n50 53.0054
R22942 a_n3827_n3924.n4 a_n3827_n3924.n3 53.0052
R22943 a_n3827_n3924.n6 a_n3827_n3924.n5 53.0052
R22944 a_n3827_n3924.n8 a_n3827_n3924.n7 53.0052
R22945 a_n3827_n3924.n10 a_n3827_n3924.n9 53.0052
R22946 a_n3827_n3924.n14 a_n3827_n3924.n13 53.0052
R22947 a_n3827_n3924.n16 a_n3827_n3924.n15 53.0052
R22948 a_n3827_n3924.n18 a_n3827_n3924.n17 53.0052
R22949 a_n3827_n3924.n20 a_n3827_n3924.n19 53.0052
R22950 a_n3827_n3924.n37 a_n3827_n3924.n36 53.0051
R22951 a_n3827_n3924.n39 a_n3827_n3924.n38 53.0051
R22952 a_n3827_n3924.n41 a_n3827_n3924.n40 53.0051
R22953 a_n3827_n3924.n43 a_n3827_n3924.n42 53.0051
R22954 a_n3827_n3924.n47 a_n3827_n3924.n46 53.0051
R22955 a_n3827_n3924.n49 a_n3827_n3924.n48 53.0051
R22956 a_n3827_n3924.n1 a_n3827_n3924.n0 53.0051
R22957 a_n3827_n3924.n23 a_n3827_n3924.n21 12.1986
R22958 a_n3827_n3924.n34 a_n3827_n3924.n2 12.1986
R22959 a_n3827_n3924.n23 a_n3827_n3924.n22 5.11903
R22960 a_n3827_n3924.n35 a_n3827_n3924.n34 5.11903
R22961 a_n3827_n3924.n36 a_n3827_n3924.t28 2.82907
R22962 a_n3827_n3924.n36 a_n3827_n3924.t31 2.82907
R22963 a_n3827_n3924.n38 a_n3827_n3924.t22 2.82907
R22964 a_n3827_n3924.n38 a_n3827_n3924.t26 2.82907
R22965 a_n3827_n3924.n40 a_n3827_n3924.t43 2.82907
R22966 a_n3827_n3924.n40 a_n3827_n3924.t33 2.82907
R22967 a_n3827_n3924.n42 a_n3827_n3924.t38 2.82907
R22968 a_n3827_n3924.n42 a_n3827_n3924.t47 2.82907
R22969 a_n3827_n3924.n46 a_n3827_n3924.t10 2.82907
R22970 a_n3827_n3924.n46 a_n3827_n3924.t15 2.82907
R22971 a_n3827_n3924.n48 a_n3827_n3924.t7 2.82907
R22972 a_n3827_n3924.n48 a_n3827_n3924.t6 2.82907
R22973 a_n3827_n3924.n0 a_n3827_n3924.t11 2.82907
R22974 a_n3827_n3924.n0 a_n3827_n3924.t17 2.82907
R22975 a_n3827_n3924.n3 a_n3827_n3924.t14 2.82907
R22976 a_n3827_n3924.n3 a_n3827_n3924.t16 2.82907
R22977 a_n3827_n3924.n5 a_n3827_n3924.t18 2.82907
R22978 a_n3827_n3924.n5 a_n3827_n3924.t19 2.82907
R22979 a_n3827_n3924.n7 a_n3827_n3924.t5 2.82907
R22980 a_n3827_n3924.n7 a_n3827_n3924.t3 2.82907
R22981 a_n3827_n3924.n9 a_n3827_n3924.t9 2.82907
R22982 a_n3827_n3924.n9 a_n3827_n3924.t4 2.82907
R22983 a_n3827_n3924.n13 a_n3827_n3924.t46 2.82907
R22984 a_n3827_n3924.n13 a_n3827_n3924.t23 2.82907
R22985 a_n3827_n3924.n15 a_n3827_n3924.t41 2.82907
R22986 a_n3827_n3924.n15 a_n3827_n3924.t1 2.82907
R22987 a_n3827_n3924.n17 a_n3827_n3924.t45 2.82907
R22988 a_n3827_n3924.n17 a_n3827_n3924.t34 2.82907
R22989 a_n3827_n3924.n19 a_n3827_n3924.t30 2.82907
R22990 a_n3827_n3924.n19 a_n3827_n3924.t35 2.82907
R22991 a_n3827_n3924.t21 a_n3827_n3924.n51 2.82907
R22992 a_n3827_n3924.n51 a_n3827_n3924.t20 2.82907
R22993 a_n3827_n3924.n25 a_n3827_n3924.n23 1.95694
R22994 a_n3827_n3924.n34 a_n3827_n3924.n33 1.95694
R22995 a_n3827_n3924.n27 a_n3827_n3924.n26 0.672012
R22996 a_n3827_n3924.n28 a_n3827_n3924.n27 0.672012
R22997 a_n3827_n3924.n29 a_n3827_n3924.n28 0.672012
R22998 a_n3827_n3924.n30 a_n3827_n3924.n29 0.672012
R22999 a_n3827_n3924.n31 a_n3827_n3924.n30 0.672012
R23000 a_n3827_n3924.n25 a_n3827_n3924.n24 0.621866
R23001 a_n3827_n3924.n33 a_n3827_n3924.n31 0.579715
R23002 a_n3827_n3924.n21 a_n3827_n3924.n20 0.444466
R23003 a_n3827_n3924.n20 a_n3827_n3924.n18 0.444466
R23004 a_n3827_n3924.n18 a_n3827_n3924.n16 0.444466
R23005 a_n3827_n3924.n16 a_n3827_n3924.n14 0.444466
R23006 a_n3827_n3924.n14 a_n3827_n3924.n12 0.444466
R23007 a_n3827_n3924.n11 a_n3827_n3924.n10 0.444466
R23008 a_n3827_n3924.n10 a_n3827_n3924.n8 0.444466
R23009 a_n3827_n3924.n8 a_n3827_n3924.n6 0.444466
R23010 a_n3827_n3924.n6 a_n3827_n3924.n4 0.444466
R23011 a_n3827_n3924.n4 a_n3827_n3924.n2 0.444466
R23012 a_n3827_n3924.n22 a_n3827_n3924.n1 0.444466
R23013 a_n3827_n3924.n50 a_n3827_n3924.n1 0.444466
R23014 a_n3827_n3924.n50 a_n3827_n3924.n49 0.444466
R23015 a_n3827_n3924.n49 a_n3827_n3924.n47 0.444466
R23016 a_n3827_n3924.n47 a_n3827_n3924.n45 0.444466
R23017 a_n3827_n3924.n44 a_n3827_n3924.n43 0.444466
R23018 a_n3827_n3924.n43 a_n3827_n3924.n41 0.444466
R23019 a_n3827_n3924.n41 a_n3827_n3924.n39 0.444466
R23020 a_n3827_n3924.n39 a_n3827_n3924.n37 0.444466
R23021 a_n3827_n3924.n37 a_n3827_n3924.n35 0.444466
R23022 a_n3827_n3924.n12 a_n3827_n3924.n11 0.235414
R23023 a_n3827_n3924.n45 a_n3827_n3924.n44 0.235414
R23024 a_n3827_n3924.n33 a_n3827_n3924.n32 0.0927965
R23025 a_n3827_n3924.n26 a_n3827_n3924.n25 0.0506453
R23026 a_n1996_n452.n80 a_n1996_n452.t59 512.366
R23027 a_n1996_n452.n79 a_n1996_n452.t50 512.366
R23028 a_n1996_n452.n78 a_n1996_n452.t44 512.366
R23029 a_n1996_n452.n82 a_n1996_n452.t67 512.366
R23030 a_n1996_n452.n81 a_n1996_n452.t56 512.366
R23031 a_n1996_n452.n77 a_n1996_n452.t55 512.366
R23032 a_n1996_n452.n84 a_n1996_n452.t63 512.366
R23033 a_n1996_n452.n83 a_n1996_n452.t48 512.366
R23034 a_n1996_n452.n76 a_n1996_n452.t49 512.366
R23035 a_n1996_n452.n86 a_n1996_n452.t51 512.366
R23036 a_n1996_n452.n85 a_n1996_n452.t61 512.366
R23037 a_n1996_n452.n75 a_n1996_n452.t71 512.366
R23038 a_n1996_n452.n25 a_n1996_n452.t70 539.01
R23039 a_n1996_n452.n67 a_n1996_n452.t53 512.366
R23040 a_n1996_n452.n66 a_n1996_n452.t57 512.366
R23041 a_n1996_n452.n64 a_n1996_n452.t47 512.366
R23042 a_n1996_n452.n65 a_n1996_n452.t62 512.366
R23043 a_n1996_n452.n21 a_n1996_n452.t24 539.01
R23044 a_n1996_n452.n70 a_n1996_n452.t28 512.366
R23045 a_n1996_n452.n69 a_n1996_n452.t30 512.366
R23046 a_n1996_n452.n53 a_n1996_n452.t18 512.366
R23047 a_n1996_n452.n68 a_n1996_n452.t20 512.366
R23048 a_n1996_n452.n15 a_n1996_n452.t26 539.01
R23049 a_n1996_n452.n91 a_n1996_n452.t36 512.366
R23050 a_n1996_n452.n92 a_n1996_n452.t14 512.366
R23051 a_n1996_n452.n51 a_n1996_n452.t32 512.366
R23052 a_n1996_n452.n93 a_n1996_n452.t34 512.366
R23053 a_n1996_n452.n19 a_n1996_n452.t65 539.01
R23054 a_n1996_n452.n88 a_n1996_n452.t66 512.366
R23055 a_n1996_n452.n89 a_n1996_n452.t45 512.366
R23056 a_n1996_n452.n52 a_n1996_n452.t52 512.366
R23057 a_n1996_n452.n90 a_n1996_n452.t60 512.366
R23058 a_n1996_n452.n4 a_n1996_n452.n49 70.1674
R23059 a_n1996_n452.n6 a_n1996_n452.n47 70.1674
R23060 a_n1996_n452.n8 a_n1996_n452.n45 70.1674
R23061 a_n1996_n452.n10 a_n1996_n452.n43 70.1674
R23062 a_n1996_n452.n32 a_n1996_n452.n23 70.3058
R23063 a_n1996_n452.n50 a_n1996_n452.n28 70.3058
R23064 a_n1996_n452.n24 a_n1996_n452.n30 70.1674
R23065 a_n1996_n452.n30 a_n1996_n452.n64 20.9683
R23066 a_n1996_n452.n29 a_n1996_n452.n24 75.0448
R23067 a_n1996_n452.n66 a_n1996_n452.n29 11.2134
R23068 a_n1996_n452.n22 a_n1996_n452.n25 44.8194
R23069 a_n1996_n452.n28 a_n1996_n452.n35 70.1674
R23070 a_n1996_n452.n35 a_n1996_n452.n53 20.9683
R23071 a_n1996_n452.n34 a_n1996_n452.n33 75.0448
R23072 a_n1996_n452.n69 a_n1996_n452.n34 11.2134
R23073 a_n1996_n452.n20 a_n1996_n452.n21 44.8194
R23074 a_n1996_n452.n12 a_n1996_n452.n41 70.3058
R23075 a_n1996_n452.n16 a_n1996_n452.n38 70.3058
R23076 a_n1996_n452.n37 a_n1996_n452.n17 70.1674
R23077 a_n1996_n452.n37 a_n1996_n452.n52 20.9683
R23078 a_n1996_n452.n17 a_n1996_n452.n36 75.0448
R23079 a_n1996_n452.n89 a_n1996_n452.n36 11.2134
R23080 a_n1996_n452.n18 a_n1996_n452.n19 44.8194
R23081 a_n1996_n452.n40 a_n1996_n452.n13 70.1674
R23082 a_n1996_n452.n40 a_n1996_n452.n51 20.9683
R23083 a_n1996_n452.n13 a_n1996_n452.n39 75.0448
R23084 a_n1996_n452.n92 a_n1996_n452.n39 11.2134
R23085 a_n1996_n452.n14 a_n1996_n452.n15 44.8194
R23086 a_n1996_n452.n43 a_n1996_n452.n75 20.9683
R23087 a_n1996_n452.n42 a_n1996_n452.n11 75.0448
R23088 a_n1996_n452.n85 a_n1996_n452.n42 11.2134
R23089 a_n1996_n452.n11 a_n1996_n452.n86 161.3
R23090 a_n1996_n452.n45 a_n1996_n452.n76 20.9683
R23091 a_n1996_n452.n44 a_n1996_n452.n9 75.0448
R23092 a_n1996_n452.n83 a_n1996_n452.n44 11.2134
R23093 a_n1996_n452.n9 a_n1996_n452.n84 161.3
R23094 a_n1996_n452.n47 a_n1996_n452.n77 20.9683
R23095 a_n1996_n452.n46 a_n1996_n452.n7 75.0448
R23096 a_n1996_n452.n81 a_n1996_n452.n46 11.2134
R23097 a_n1996_n452.n7 a_n1996_n452.n82 161.3
R23098 a_n1996_n452.n49 a_n1996_n452.n78 20.9683
R23099 a_n1996_n452.n48 a_n1996_n452.n5 75.0448
R23100 a_n1996_n452.n79 a_n1996_n452.n48 11.2134
R23101 a_n1996_n452.n5 a_n1996_n452.n80 161.3
R23102 a_n1996_n452.n3 a_n1996_n452.n62 81.3764
R23103 a_n1996_n452.n1 a_n1996_n452.n57 81.3764
R23104 a_n1996_n452.n0 a_n1996_n452.n54 81.3764
R23105 a_n1996_n452.n3 a_n1996_n452.n63 80.9324
R23106 a_n1996_n452.n3 a_n1996_n452.n61 80.9324
R23107 a_n1996_n452.n2 a_n1996_n452.n60 80.9324
R23108 a_n1996_n452.n2 a_n1996_n452.n59 80.9324
R23109 a_n1996_n452.n1 a_n1996_n452.n58 80.9324
R23110 a_n1996_n452.n1 a_n1996_n452.n56 80.9324
R23111 a_n1996_n452.n0 a_n1996_n452.n55 80.9324
R23112 a_n1996_n452.n96 a_n1996_n452.t27 74.6477
R23113 a_n1996_n452.n26 a_n1996_n452.t23 74.6477
R23114 a_n1996_n452.n73 a_n1996_n452.t25 74.2899
R23115 a_n1996_n452.n27 a_n1996_n452.t17 74.2897
R23116 a_n1996_n452.n27 a_n1996_n452.n95 70.6783
R23117 a_n1996_n452.n26 a_n1996_n452.n71 70.6783
R23118 a_n1996_n452.n26 a_n1996_n452.n72 70.6783
R23119 a_n1996_n452.n97 a_n1996_n452.n96 70.6782
R23120 a_n1996_n452.n80 a_n1996_n452.n79 48.2005
R23121 a_n1996_n452.t64 a_n1996_n452.n49 533.335
R23122 a_n1996_n452.n82 a_n1996_n452.n81 48.2005
R23123 a_n1996_n452.t69 a_n1996_n452.n47 533.335
R23124 a_n1996_n452.n84 a_n1996_n452.n83 48.2005
R23125 a_n1996_n452.t58 a_n1996_n452.n45 533.335
R23126 a_n1996_n452.n86 a_n1996_n452.n85 48.2005
R23127 a_n1996_n452.t54 a_n1996_n452.n43 533.335
R23128 a_n1996_n452.n67 a_n1996_n452.n66 48.2005
R23129 a_n1996_n452.n65 a_n1996_n452.n30 20.9683
R23130 a_n1996_n452.n70 a_n1996_n452.n69 48.2005
R23131 a_n1996_n452.n68 a_n1996_n452.n35 20.9683
R23132 a_n1996_n452.n92 a_n1996_n452.n91 48.2005
R23133 a_n1996_n452.n93 a_n1996_n452.n40 20.9683
R23134 a_n1996_n452.n89 a_n1996_n452.n88 48.2005
R23135 a_n1996_n452.n90 a_n1996_n452.n37 20.9683
R23136 a_n1996_n452.n32 a_n1996_n452.t68 533.058
R23137 a_n1996_n452.n50 a_n1996_n452.t22 533.058
R23138 a_n1996_n452.t16 a_n1996_n452.n41 533.058
R23139 a_n1996_n452.t46 a_n1996_n452.n38 533.058
R23140 a_n1996_n452.n2 a_n1996_n452.n1 32.0139
R23141 a_n1996_n452.n48 a_n1996_n452.n78 35.3134
R23142 a_n1996_n452.n46 a_n1996_n452.n77 35.3134
R23143 a_n1996_n452.n44 a_n1996_n452.n76 35.3134
R23144 a_n1996_n452.n42 a_n1996_n452.n75 35.3134
R23145 a_n1996_n452.n29 a_n1996_n452.n64 35.3134
R23146 a_n1996_n452.n34 a_n1996_n452.n53 35.3134
R23147 a_n1996_n452.n51 a_n1996_n452.n39 35.3134
R23148 a_n1996_n452.n52 a_n1996_n452.n36 35.3134
R23149 a_n1996_n452.n28 a_n1996_n452.n3 23.891
R23150 a_n1996_n452.n18 a_n1996_n452.n87 12.046
R23151 a_n1996_n452.n23 a_n1996_n452.n31 11.8414
R23152 a_n1996_n452.n74 a_n1996_n452.n20 10.5365
R23153 a_n1996_n452.n27 a_n1996_n452.n94 9.50122
R23154 a_n1996_n452.n87 a_n1996_n452.n11 7.47588
R23155 a_n1996_n452.n4 a_n1996_n452.n31 7.47588
R23156 a_n1996_n452.n94 a_n1996_n452.n12 6.70126
R23157 a_n1996_n452.n74 a_n1996_n452.n73 5.65783
R23158 a_n1996_n452.n94 a_n1996_n452.n31 5.3452
R23159 a_n1996_n452.n28 a_n1996_n452.n22 3.95126
R23160 a_n1996_n452.n14 a_n1996_n452.n16 3.95126
R23161 a_n1996_n452.n95 a_n1996_n452.t33 3.61217
R23162 a_n1996_n452.n95 a_n1996_n452.t35 3.61217
R23163 a_n1996_n452.n71 a_n1996_n452.t19 3.61217
R23164 a_n1996_n452.n71 a_n1996_n452.t21 3.61217
R23165 a_n1996_n452.n72 a_n1996_n452.t29 3.61217
R23166 a_n1996_n452.n72 a_n1996_n452.t31 3.61217
R23167 a_n1996_n452.n97 a_n1996_n452.t37 3.61217
R23168 a_n1996_n452.t15 a_n1996_n452.n97 3.61217
R23169 a_n1996_n452.n62 a_n1996_n452.t2 2.82907
R23170 a_n1996_n452.n62 a_n1996_n452.t5 2.82907
R23171 a_n1996_n452.n63 a_n1996_n452.t0 2.82907
R23172 a_n1996_n452.n63 a_n1996_n452.t42 2.82907
R23173 a_n1996_n452.n61 a_n1996_n452.t10 2.82907
R23174 a_n1996_n452.n61 a_n1996_n452.t38 2.82907
R23175 a_n1996_n452.n60 a_n1996_n452.t11 2.82907
R23176 a_n1996_n452.n60 a_n1996_n452.t41 2.82907
R23177 a_n1996_n452.n59 a_n1996_n452.t8 2.82907
R23178 a_n1996_n452.n59 a_n1996_n452.t6 2.82907
R23179 a_n1996_n452.n57 a_n1996_n452.t7 2.82907
R23180 a_n1996_n452.n57 a_n1996_n452.t12 2.82907
R23181 a_n1996_n452.n58 a_n1996_n452.t3 2.82907
R23182 a_n1996_n452.n58 a_n1996_n452.t4 2.82907
R23183 a_n1996_n452.n56 a_n1996_n452.t9 2.82907
R23184 a_n1996_n452.n56 a_n1996_n452.t1 2.82907
R23185 a_n1996_n452.n55 a_n1996_n452.t43 2.82907
R23186 a_n1996_n452.n55 a_n1996_n452.t40 2.82907
R23187 a_n1996_n452.n54 a_n1996_n452.t39 2.82907
R23188 a_n1996_n452.n54 a_n1996_n452.t13 2.82907
R23189 a_n1996_n452.n87 a_n1996_n452.n74 1.30542
R23190 a_n1996_n452.n8 a_n1996_n452.n7 1.04595
R23191 a_n1996_n452.n25 a_n1996_n452.n67 13.657
R23192 a_n1996_n452.n65 a_n1996_n452.n32 21.4216
R23193 a_n1996_n452.n21 a_n1996_n452.n70 13.657
R23194 a_n1996_n452.n68 a_n1996_n452.n50 21.4216
R23195 a_n1996_n452.n91 a_n1996_n452.n15 13.657
R23196 a_n1996_n452.n41 a_n1996_n452.n93 21.4216
R23197 a_n1996_n452.n88 a_n1996_n452.n19 13.657
R23198 a_n1996_n452.n38 a_n1996_n452.n90 21.4216
R23199 a_n1996_n452.n3 a_n1996_n452.n2 1.3324
R23200 a_n1996_n452.n1 a_n1996_n452.n0 0.888431
R23201 a_n1996_n452.n24 a_n1996_n452.n22 0.758076
R23202 a_n1996_n452.n24 a_n1996_n452.n23 0.758076
R23203 a_n1996_n452.n33 a_n1996_n452.n20 0.758076
R23204 a_n1996_n452.n18 a_n1996_n452.n17 0.758076
R23205 a_n1996_n452.n17 a_n1996_n452.n16 0.758076
R23206 a_n1996_n452.n14 a_n1996_n452.n13 0.758076
R23207 a_n1996_n452.n13 a_n1996_n452.n12 0.758076
R23208 a_n1996_n452.n11 a_n1996_n452.n10 0.758076
R23209 a_n1996_n452.n9 a_n1996_n452.n8 0.758076
R23210 a_n1996_n452.n7 a_n1996_n452.n6 0.758076
R23211 a_n1996_n452.n5 a_n1996_n452.n4 0.758076
R23212 a_n1996_n452.n33 a_n1996_n452.n28 0.720197
R23213 a_n1996_n452.n96 a_n1996_n452.n27 0.716017
R23214 a_n1996_n452.n73 a_n1996_n452.n26 0.716017
R23215 a_n1996_n452.n10 a_n1996_n452.n9 0.67853
R23216 a_n1996_n452.n6 a_n1996_n452.n5 0.67853
R23217 a_n1808_13878.n2 a_n1808_13878.n0 98.9633
R23218 a_n1808_13878.n5 a_n1808_13878.n3 98.7517
R23219 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R23220 a_n1808_13878.n7 a_n1808_13878.n6 98.6055
R23221 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R23222 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R23223 a_n1808_13878.n9 a_n1808_13878.t1 74.6477
R23224 a_n1808_13878.n14 a_n1808_13878.t2 74.2899
R23225 a_n1808_13878.n11 a_n1808_13878.t3 74.2899
R23226 a_n1808_13878.n10 a_n1808_13878.t0 74.2899
R23227 a_n1808_13878.n13 a_n1808_13878.n12 70.6783
R23228 a_n1808_13878.n9 a_n1808_13878.n8 70.6783
R23229 a_n1808_13878.n15 a_n1808_13878.n7 13.5694
R23230 a_n1808_13878.n16 a_n1808_13878.n15 11.5762
R23231 a_n1808_13878.n15 a_n1808_13878.n14 6.2408
R23232 a_n1808_13878.n1 a_n1808_13878.t8 3.61217
R23233 a_n1808_13878.n1 a_n1808_13878.t13 3.61217
R23234 a_n1808_13878.n0 a_n1808_13878.t15 3.61217
R23235 a_n1808_13878.n0 a_n1808_13878.t19 3.61217
R23236 a_n1808_13878.n12 a_n1808_13878.t6 3.61217
R23237 a_n1808_13878.n12 a_n1808_13878.t7 3.61217
R23238 a_n1808_13878.n8 a_n1808_13878.t4 3.61217
R23239 a_n1808_13878.n8 a_n1808_13878.t5 3.61217
R23240 a_n1808_13878.n6 a_n1808_13878.t14 3.61217
R23241 a_n1808_13878.n6 a_n1808_13878.t9 3.61217
R23242 a_n1808_13878.n4 a_n1808_13878.t16 3.61217
R23243 a_n1808_13878.n4 a_n1808_13878.t11 3.61217
R23244 a_n1808_13878.n3 a_n1808_13878.t10 3.61217
R23245 a_n1808_13878.n3 a_n1808_13878.t12 3.61217
R23246 a_n1808_13878.n17 a_n1808_13878.t17 3.61217
R23247 a_n1808_13878.t18 a_n1808_13878.n17 3.61217
R23248 a_n1808_13878.n10 a_n1808_13878.n9 0.358259
R23249 a_n1808_13878.n13 a_n1808_13878.n11 0.358259
R23250 a_n1808_13878.n14 a_n1808_13878.n13 0.358259
R23251 a_n1808_13878.n16 a_n1808_13878.n2 0.358259
R23252 a_n1808_13878.n7 a_n1808_13878.n5 0.146627
R23253 a_n1808_13878.n11 a_n1808_13878.n10 0.101793
R23254 diffpairibias.n0 diffpairibias.t27 436.822
R23255 diffpairibias.n27 diffpairibias.t24 435.479
R23256 diffpairibias.n26 diffpairibias.t21 435.479
R23257 diffpairibias.n25 diffpairibias.t22 435.479
R23258 diffpairibias.n24 diffpairibias.t26 435.479
R23259 diffpairibias.n23 diffpairibias.t20 435.479
R23260 diffpairibias.n0 diffpairibias.t23 435.479
R23261 diffpairibias.n1 diffpairibias.t28 435.479
R23262 diffpairibias.n2 diffpairibias.t25 435.479
R23263 diffpairibias.n3 diffpairibias.t29 435.479
R23264 diffpairibias.n13 diffpairibias.t14 377.536
R23265 diffpairibias.n13 diffpairibias.t0 376.193
R23266 diffpairibias.n14 diffpairibias.t10 376.193
R23267 diffpairibias.n15 diffpairibias.t12 376.193
R23268 diffpairibias.n16 diffpairibias.t6 376.193
R23269 diffpairibias.n17 diffpairibias.t2 376.193
R23270 diffpairibias.n18 diffpairibias.t16 376.193
R23271 diffpairibias.n19 diffpairibias.t4 376.193
R23272 diffpairibias.n20 diffpairibias.t18 376.193
R23273 diffpairibias.n21 diffpairibias.t8 376.193
R23274 diffpairibias.n4 diffpairibias.t15 113.368
R23275 diffpairibias.n4 diffpairibias.t1 112.698
R23276 diffpairibias.n5 diffpairibias.t11 112.698
R23277 diffpairibias.n6 diffpairibias.t13 112.698
R23278 diffpairibias.n7 diffpairibias.t7 112.698
R23279 diffpairibias.n8 diffpairibias.t3 112.698
R23280 diffpairibias.n9 diffpairibias.t17 112.698
R23281 diffpairibias.n10 diffpairibias.t5 112.698
R23282 diffpairibias.n11 diffpairibias.t19 112.698
R23283 diffpairibias.n12 diffpairibias.t9 112.698
R23284 diffpairibias.n22 diffpairibias.n21 4.77242
R23285 diffpairibias.n22 diffpairibias.n12 4.30807
R23286 diffpairibias.n23 diffpairibias.n22 4.13945
R23287 diffpairibias.n21 diffpairibias.n20 1.34352
R23288 diffpairibias.n20 diffpairibias.n19 1.34352
R23289 diffpairibias.n19 diffpairibias.n18 1.34352
R23290 diffpairibias.n18 diffpairibias.n17 1.34352
R23291 diffpairibias.n17 diffpairibias.n16 1.34352
R23292 diffpairibias.n16 diffpairibias.n15 1.34352
R23293 diffpairibias.n15 diffpairibias.n14 1.34352
R23294 diffpairibias.n14 diffpairibias.n13 1.34352
R23295 diffpairibias.n3 diffpairibias.n2 1.34352
R23296 diffpairibias.n2 diffpairibias.n1 1.34352
R23297 diffpairibias.n1 diffpairibias.n0 1.34352
R23298 diffpairibias.n24 diffpairibias.n23 1.34352
R23299 diffpairibias.n25 diffpairibias.n24 1.34352
R23300 diffpairibias.n26 diffpairibias.n25 1.34352
R23301 diffpairibias.n27 diffpairibias.n26 1.34352
R23302 diffpairibias.n28 diffpairibias.n27 0.862419
R23303 diffpairibias diffpairibias.n28 0.684875
R23304 diffpairibias.n12 diffpairibias.n11 0.672012
R23305 diffpairibias.n11 diffpairibias.n10 0.672012
R23306 diffpairibias.n10 diffpairibias.n9 0.672012
R23307 diffpairibias.n9 diffpairibias.n8 0.672012
R23308 diffpairibias.n8 diffpairibias.n7 0.672012
R23309 diffpairibias.n7 diffpairibias.n6 0.672012
R23310 diffpairibias.n6 diffpairibias.n5 0.672012
R23311 diffpairibias.n5 diffpairibias.n4 0.672012
R23312 diffpairibias.n28 diffpairibias.n3 0.190907
R23313 minus.n43 minus.t24 322.512
R23314 minus.n9 minus.t8 322.512
R23315 minus.n66 minus.t5 297.12
R23316 minus.n64 minus.t6 297.12
R23317 minus.n36 minus.t22 297.12
R23318 minus.n58 minus.t18 297.12
R23319 minus.n38 minus.t19 297.12
R23320 minus.n52 minus.t14 297.12
R23321 minus.n40 minus.t15 297.12
R23322 minus.n46 minus.t9 297.12
R23323 minus.n42 minus.t23 297.12
R23324 minus.n8 minus.t7 297.12
R23325 minus.n12 minus.t11 297.12
R23326 minus.n14 minus.t10 297.12
R23327 minus.n18 minus.t12 297.12
R23328 minus.n20 minus.t17 297.12
R23329 minus.n24 minus.t16 297.12
R23330 minus.n26 minus.t21 297.12
R23331 minus.n30 minus.t20 297.12
R23332 minus.n32 minus.t13 297.12
R23333 minus.n72 minus.t4 243.255
R23334 minus.n71 minus.n69 224.169
R23335 minus.n71 minus.n70 223.454
R23336 minus.n45 minus.n44 161.3
R23337 minus.n46 minus.n41 161.3
R23338 minus.n48 minus.n47 161.3
R23339 minus.n49 minus.n40 161.3
R23340 minus.n51 minus.n50 161.3
R23341 minus.n52 minus.n39 161.3
R23342 minus.n54 minus.n53 161.3
R23343 minus.n55 minus.n38 161.3
R23344 minus.n57 minus.n56 161.3
R23345 minus.n58 minus.n37 161.3
R23346 minus.n60 minus.n59 161.3
R23347 minus.n61 minus.n36 161.3
R23348 minus.n63 minus.n62 161.3
R23349 minus.n64 minus.n35 161.3
R23350 minus.n65 minus.n34 161.3
R23351 minus.n67 minus.n66 161.3
R23352 minus.n33 minus.n32 161.3
R23353 minus.n31 minus.n0 161.3
R23354 minus.n30 minus.n29 161.3
R23355 minus.n28 minus.n1 161.3
R23356 minus.n27 minus.n26 161.3
R23357 minus.n25 minus.n2 161.3
R23358 minus.n24 minus.n23 161.3
R23359 minus.n22 minus.n3 161.3
R23360 minus.n21 minus.n20 161.3
R23361 minus.n19 minus.n4 161.3
R23362 minus.n18 minus.n17 161.3
R23363 minus.n16 minus.n5 161.3
R23364 minus.n15 minus.n14 161.3
R23365 minus.n13 minus.n6 161.3
R23366 minus.n12 minus.n11 161.3
R23367 minus.n10 minus.n7 161.3
R23368 minus.n44 minus.n43 45.0031
R23369 minus.n10 minus.n9 45.0031
R23370 minus.n66 minus.n65 41.6278
R23371 minus.n32 minus.n31 41.6278
R23372 minus.n64 minus.n63 37.246
R23373 minus.n45 minus.n42 37.246
R23374 minus.n8 minus.n7 37.246
R23375 minus.n30 minus.n1 37.246
R23376 minus.n59 minus.n36 32.8641
R23377 minus.n47 minus.n46 32.8641
R23378 minus.n13 minus.n12 32.8641
R23379 minus.n26 minus.n25 32.8641
R23380 minus.n68 minus.n67 31.8206
R23381 minus.n58 minus.n57 28.4823
R23382 minus.n51 minus.n40 28.4823
R23383 minus.n14 minus.n5 28.4823
R23384 minus.n24 minus.n3 28.4823
R23385 minus.n53 minus.n38 24.1005
R23386 minus.n53 minus.n52 24.1005
R23387 minus.n19 minus.n18 24.1005
R23388 minus.n20 minus.n19 24.1005
R23389 minus.n70 minus.t3 19.8005
R23390 minus.n70 minus.t1 19.8005
R23391 minus.n69 minus.t2 19.8005
R23392 minus.n69 minus.t0 19.8005
R23393 minus.n57 minus.n38 19.7187
R23394 minus.n52 minus.n51 19.7187
R23395 minus.n18 minus.n5 19.7187
R23396 minus.n20 minus.n3 19.7187
R23397 minus.n43 minus.n42 15.6319
R23398 minus.n9 minus.n8 15.6319
R23399 minus.n59 minus.n58 15.3369
R23400 minus.n47 minus.n40 15.3369
R23401 minus.n14 minus.n13 15.3369
R23402 minus.n25 minus.n24 15.3369
R23403 minus.n68 minus.n33 12.0819
R23404 minus minus.n73 11.8293
R23405 minus.n63 minus.n36 10.955
R23406 minus.n46 minus.n45 10.955
R23407 minus.n12 minus.n7 10.955
R23408 minus.n26 minus.n1 10.955
R23409 minus.n65 minus.n64 6.57323
R23410 minus.n31 minus.n30 6.57323
R23411 minus.n73 minus.n72 4.80222
R23412 minus.n73 minus.n68 0.972091
R23413 minus.n72 minus.n71 0.716017
R23414 minus.n67 minus.n34 0.189894
R23415 minus.n35 minus.n34 0.189894
R23416 minus.n62 minus.n35 0.189894
R23417 minus.n62 minus.n61 0.189894
R23418 minus.n61 minus.n60 0.189894
R23419 minus.n60 minus.n37 0.189894
R23420 minus.n56 minus.n37 0.189894
R23421 minus.n56 minus.n55 0.189894
R23422 minus.n55 minus.n54 0.189894
R23423 minus.n54 minus.n39 0.189894
R23424 minus.n50 minus.n39 0.189894
R23425 minus.n50 minus.n49 0.189894
R23426 minus.n49 minus.n48 0.189894
R23427 minus.n48 minus.n41 0.189894
R23428 minus.n44 minus.n41 0.189894
R23429 minus.n11 minus.n10 0.189894
R23430 minus.n11 minus.n6 0.189894
R23431 minus.n15 minus.n6 0.189894
R23432 minus.n16 minus.n15 0.189894
R23433 minus.n17 minus.n16 0.189894
R23434 minus.n17 minus.n4 0.189894
R23435 minus.n21 minus.n4 0.189894
R23436 minus.n22 minus.n21 0.189894
R23437 minus.n23 minus.n22 0.189894
R23438 minus.n23 minus.n2 0.189894
R23439 minus.n27 minus.n2 0.189894
R23440 minus.n28 minus.n27 0.189894
R23441 minus.n29 minus.n28 0.189894
R23442 minus.n29 minus.n0 0.189894
R23443 minus.n33 minus.n0 0.189894
R23444 a_n1986_8322.n6 a_n1986_8322.t3 74.6477
R23445 a_n1986_8322.n1 a_n1986_8322.t9 74.6477
R23446 a_n1986_8322.n16 a_n1986_8322.t18 74.6474
R23447 a_n1986_8322.n14 a_n1986_8322.t11 74.2899
R23448 a_n1986_8322.n7 a_n1986_8322.t1 74.2899
R23449 a_n1986_8322.n8 a_n1986_8322.t4 74.2899
R23450 a_n1986_8322.n11 a_n1986_8322.t5 74.2899
R23451 a_n1986_8322.n4 a_n1986_8322.t8 74.2899
R23452 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R23453 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R23454 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R23455 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R23456 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R23457 a_n1986_8322.n18 a_n1986_8322.n17 70.6782
R23458 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R23459 a_n1986_8322.n13 a_n1986_8322.t20 10.109
R23460 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R23461 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R23462 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R23463 a_n1986_8322.n15 a_n1986_8322.t16 3.61217
R23464 a_n1986_8322.n15 a_n1986_8322.t13 3.61217
R23465 a_n1986_8322.n5 a_n1986_8322.t7 3.61217
R23466 a_n1986_8322.n5 a_n1986_8322.t6 3.61217
R23467 a_n1986_8322.n9 a_n1986_8322.t2 3.61217
R23468 a_n1986_8322.n9 a_n1986_8322.t0 3.61217
R23469 a_n1986_8322.n0 a_n1986_8322.t17 3.61217
R23470 a_n1986_8322.n0 a_n1986_8322.t12 3.61217
R23471 a_n1986_8322.n2 a_n1986_8322.t15 3.61217
R23472 a_n1986_8322.n2 a_n1986_8322.t14 3.61217
R23473 a_n1986_8322.n18 a_n1986_8322.t10 3.61217
R23474 a_n1986_8322.t19 a_n1986_8322.n18 3.61217
R23475 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R23476 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R23477 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R23478 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R23479 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R23480 a_n1986_8322.n17 a_n1986_8322.n14 0.358259
R23481 a_n1986_8322.n17 a_n1986_8322.n16 0.358259
R23482 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R23483 a_n1986_8322.t20 a_n1986_8322.t21 0.057021
R23484 outputibias.n27 outputibias.n1 289.615
R23485 outputibias.n58 outputibias.n32 289.615
R23486 outputibias.n90 outputibias.n64 289.615
R23487 outputibias.n122 outputibias.n96 289.615
R23488 outputibias.n28 outputibias.n27 185
R23489 outputibias.n26 outputibias.n25 185
R23490 outputibias.n5 outputibias.n4 185
R23491 outputibias.n20 outputibias.n19 185
R23492 outputibias.n18 outputibias.n17 185
R23493 outputibias.n9 outputibias.n8 185
R23494 outputibias.n12 outputibias.n11 185
R23495 outputibias.n59 outputibias.n58 185
R23496 outputibias.n57 outputibias.n56 185
R23497 outputibias.n36 outputibias.n35 185
R23498 outputibias.n51 outputibias.n50 185
R23499 outputibias.n49 outputibias.n48 185
R23500 outputibias.n40 outputibias.n39 185
R23501 outputibias.n43 outputibias.n42 185
R23502 outputibias.n91 outputibias.n90 185
R23503 outputibias.n89 outputibias.n88 185
R23504 outputibias.n68 outputibias.n67 185
R23505 outputibias.n83 outputibias.n82 185
R23506 outputibias.n81 outputibias.n80 185
R23507 outputibias.n72 outputibias.n71 185
R23508 outputibias.n75 outputibias.n74 185
R23509 outputibias.n123 outputibias.n122 185
R23510 outputibias.n121 outputibias.n120 185
R23511 outputibias.n100 outputibias.n99 185
R23512 outputibias.n115 outputibias.n114 185
R23513 outputibias.n113 outputibias.n112 185
R23514 outputibias.n104 outputibias.n103 185
R23515 outputibias.n107 outputibias.n106 185
R23516 outputibias.n0 outputibias.t9 178.945
R23517 outputibias.n133 outputibias.t8 177.018
R23518 outputibias.n132 outputibias.t11 177.018
R23519 outputibias.n0 outputibias.t10 177.018
R23520 outputibias.t5 outputibias.n10 147.661
R23521 outputibias.t7 outputibias.n41 147.661
R23522 outputibias.t1 outputibias.n73 147.661
R23523 outputibias.t3 outputibias.n105 147.661
R23524 outputibias.n128 outputibias.t4 132.363
R23525 outputibias.n128 outputibias.t6 130.436
R23526 outputibias.n129 outputibias.t0 130.436
R23527 outputibias.n130 outputibias.t2 130.436
R23528 outputibias.n27 outputibias.n26 104.615
R23529 outputibias.n26 outputibias.n4 104.615
R23530 outputibias.n19 outputibias.n4 104.615
R23531 outputibias.n19 outputibias.n18 104.615
R23532 outputibias.n18 outputibias.n8 104.615
R23533 outputibias.n11 outputibias.n8 104.615
R23534 outputibias.n58 outputibias.n57 104.615
R23535 outputibias.n57 outputibias.n35 104.615
R23536 outputibias.n50 outputibias.n35 104.615
R23537 outputibias.n50 outputibias.n49 104.615
R23538 outputibias.n49 outputibias.n39 104.615
R23539 outputibias.n42 outputibias.n39 104.615
R23540 outputibias.n90 outputibias.n89 104.615
R23541 outputibias.n89 outputibias.n67 104.615
R23542 outputibias.n82 outputibias.n67 104.615
R23543 outputibias.n82 outputibias.n81 104.615
R23544 outputibias.n81 outputibias.n71 104.615
R23545 outputibias.n74 outputibias.n71 104.615
R23546 outputibias.n122 outputibias.n121 104.615
R23547 outputibias.n121 outputibias.n99 104.615
R23548 outputibias.n114 outputibias.n99 104.615
R23549 outputibias.n114 outputibias.n113 104.615
R23550 outputibias.n113 outputibias.n103 104.615
R23551 outputibias.n106 outputibias.n103 104.615
R23552 outputibias.n63 outputibias.n31 95.6354
R23553 outputibias.n63 outputibias.n62 94.6732
R23554 outputibias.n95 outputibias.n94 94.6732
R23555 outputibias.n127 outputibias.n126 94.6732
R23556 outputibias.n11 outputibias.t5 52.3082
R23557 outputibias.n42 outputibias.t7 52.3082
R23558 outputibias.n74 outputibias.t1 52.3082
R23559 outputibias.n106 outputibias.t3 52.3082
R23560 outputibias.n12 outputibias.n10 15.6674
R23561 outputibias.n43 outputibias.n41 15.6674
R23562 outputibias.n75 outputibias.n73 15.6674
R23563 outputibias.n107 outputibias.n105 15.6674
R23564 outputibias.n13 outputibias.n9 12.8005
R23565 outputibias.n44 outputibias.n40 12.8005
R23566 outputibias.n76 outputibias.n72 12.8005
R23567 outputibias.n108 outputibias.n104 12.8005
R23568 outputibias.n17 outputibias.n16 12.0247
R23569 outputibias.n48 outputibias.n47 12.0247
R23570 outputibias.n80 outputibias.n79 12.0247
R23571 outputibias.n112 outputibias.n111 12.0247
R23572 outputibias.n20 outputibias.n7 11.249
R23573 outputibias.n51 outputibias.n38 11.249
R23574 outputibias.n83 outputibias.n70 11.249
R23575 outputibias.n115 outputibias.n102 11.249
R23576 outputibias.n21 outputibias.n5 10.4732
R23577 outputibias.n52 outputibias.n36 10.4732
R23578 outputibias.n84 outputibias.n68 10.4732
R23579 outputibias.n116 outputibias.n100 10.4732
R23580 outputibias.n25 outputibias.n24 9.69747
R23581 outputibias.n56 outputibias.n55 9.69747
R23582 outputibias.n88 outputibias.n87 9.69747
R23583 outputibias.n120 outputibias.n119 9.69747
R23584 outputibias.n31 outputibias.n30 9.45567
R23585 outputibias.n62 outputibias.n61 9.45567
R23586 outputibias.n94 outputibias.n93 9.45567
R23587 outputibias.n126 outputibias.n125 9.45567
R23588 outputibias.n30 outputibias.n29 9.3005
R23589 outputibias.n3 outputibias.n2 9.3005
R23590 outputibias.n24 outputibias.n23 9.3005
R23591 outputibias.n22 outputibias.n21 9.3005
R23592 outputibias.n7 outputibias.n6 9.3005
R23593 outputibias.n16 outputibias.n15 9.3005
R23594 outputibias.n14 outputibias.n13 9.3005
R23595 outputibias.n61 outputibias.n60 9.3005
R23596 outputibias.n34 outputibias.n33 9.3005
R23597 outputibias.n55 outputibias.n54 9.3005
R23598 outputibias.n53 outputibias.n52 9.3005
R23599 outputibias.n38 outputibias.n37 9.3005
R23600 outputibias.n47 outputibias.n46 9.3005
R23601 outputibias.n45 outputibias.n44 9.3005
R23602 outputibias.n93 outputibias.n92 9.3005
R23603 outputibias.n66 outputibias.n65 9.3005
R23604 outputibias.n87 outputibias.n86 9.3005
R23605 outputibias.n85 outputibias.n84 9.3005
R23606 outputibias.n70 outputibias.n69 9.3005
R23607 outputibias.n79 outputibias.n78 9.3005
R23608 outputibias.n77 outputibias.n76 9.3005
R23609 outputibias.n125 outputibias.n124 9.3005
R23610 outputibias.n98 outputibias.n97 9.3005
R23611 outputibias.n119 outputibias.n118 9.3005
R23612 outputibias.n117 outputibias.n116 9.3005
R23613 outputibias.n102 outputibias.n101 9.3005
R23614 outputibias.n111 outputibias.n110 9.3005
R23615 outputibias.n109 outputibias.n108 9.3005
R23616 outputibias.n28 outputibias.n3 8.92171
R23617 outputibias.n59 outputibias.n34 8.92171
R23618 outputibias.n91 outputibias.n66 8.92171
R23619 outputibias.n123 outputibias.n98 8.92171
R23620 outputibias.n29 outputibias.n1 8.14595
R23621 outputibias.n60 outputibias.n32 8.14595
R23622 outputibias.n92 outputibias.n64 8.14595
R23623 outputibias.n124 outputibias.n96 8.14595
R23624 outputibias.n31 outputibias.n1 5.81868
R23625 outputibias.n62 outputibias.n32 5.81868
R23626 outputibias.n94 outputibias.n64 5.81868
R23627 outputibias.n126 outputibias.n96 5.81868
R23628 outputibias.n131 outputibias.n130 5.20947
R23629 outputibias.n29 outputibias.n28 5.04292
R23630 outputibias.n60 outputibias.n59 5.04292
R23631 outputibias.n92 outputibias.n91 5.04292
R23632 outputibias.n124 outputibias.n123 5.04292
R23633 outputibias.n131 outputibias.n127 4.42209
R23634 outputibias.n14 outputibias.n10 4.38594
R23635 outputibias.n45 outputibias.n41 4.38594
R23636 outputibias.n77 outputibias.n73 4.38594
R23637 outputibias.n109 outputibias.n105 4.38594
R23638 outputibias.n132 outputibias.n131 4.28454
R23639 outputibias.n25 outputibias.n3 4.26717
R23640 outputibias.n56 outputibias.n34 4.26717
R23641 outputibias.n88 outputibias.n66 4.26717
R23642 outputibias.n120 outputibias.n98 4.26717
R23643 outputibias.n24 outputibias.n5 3.49141
R23644 outputibias.n55 outputibias.n36 3.49141
R23645 outputibias.n87 outputibias.n68 3.49141
R23646 outputibias.n119 outputibias.n100 3.49141
R23647 outputibias.n21 outputibias.n20 2.71565
R23648 outputibias.n52 outputibias.n51 2.71565
R23649 outputibias.n84 outputibias.n83 2.71565
R23650 outputibias.n116 outputibias.n115 2.71565
R23651 outputibias.n17 outputibias.n7 1.93989
R23652 outputibias.n48 outputibias.n38 1.93989
R23653 outputibias.n80 outputibias.n70 1.93989
R23654 outputibias.n112 outputibias.n102 1.93989
R23655 outputibias.n130 outputibias.n129 1.9266
R23656 outputibias.n129 outputibias.n128 1.9266
R23657 outputibias.n133 outputibias.n132 1.92658
R23658 outputibias.n134 outputibias.n133 1.29913
R23659 outputibias.n16 outputibias.n9 1.16414
R23660 outputibias.n47 outputibias.n40 1.16414
R23661 outputibias.n79 outputibias.n72 1.16414
R23662 outputibias.n111 outputibias.n104 1.16414
R23663 outputibias.n127 outputibias.n95 0.962709
R23664 outputibias.n95 outputibias.n63 0.962709
R23665 outputibias.n13 outputibias.n12 0.388379
R23666 outputibias.n44 outputibias.n43 0.388379
R23667 outputibias.n76 outputibias.n75 0.388379
R23668 outputibias.n108 outputibias.n107 0.388379
R23669 outputibias.n134 outputibias.n0 0.337251
R23670 outputibias outputibias.n134 0.302375
R23671 outputibias.n30 outputibias.n2 0.155672
R23672 outputibias.n23 outputibias.n2 0.155672
R23673 outputibias.n23 outputibias.n22 0.155672
R23674 outputibias.n22 outputibias.n6 0.155672
R23675 outputibias.n15 outputibias.n6 0.155672
R23676 outputibias.n15 outputibias.n14 0.155672
R23677 outputibias.n61 outputibias.n33 0.155672
R23678 outputibias.n54 outputibias.n33 0.155672
R23679 outputibias.n54 outputibias.n53 0.155672
R23680 outputibias.n53 outputibias.n37 0.155672
R23681 outputibias.n46 outputibias.n37 0.155672
R23682 outputibias.n46 outputibias.n45 0.155672
R23683 outputibias.n93 outputibias.n65 0.155672
R23684 outputibias.n86 outputibias.n65 0.155672
R23685 outputibias.n86 outputibias.n85 0.155672
R23686 outputibias.n85 outputibias.n69 0.155672
R23687 outputibias.n78 outputibias.n69 0.155672
R23688 outputibias.n78 outputibias.n77 0.155672
R23689 outputibias.n125 outputibias.n97 0.155672
R23690 outputibias.n118 outputibias.n97 0.155672
R23691 outputibias.n118 outputibias.n117 0.155672
R23692 outputibias.n117 outputibias.n101 0.155672
R23693 outputibias.n110 outputibias.n101 0.155672
R23694 outputibias.n110 outputibias.n109 0.155672
R23695 output.n41 output.n15 289.615
R23696 output.n72 output.n46 289.615
R23697 output.n104 output.n78 289.615
R23698 output.n136 output.n110 289.615
R23699 output.n77 output.n45 197.26
R23700 output.n77 output.n76 196.298
R23701 output.n109 output.n108 196.298
R23702 output.n141 output.n140 196.298
R23703 output.n42 output.n41 185
R23704 output.n40 output.n39 185
R23705 output.n19 output.n18 185
R23706 output.n34 output.n33 185
R23707 output.n32 output.n31 185
R23708 output.n23 output.n22 185
R23709 output.n26 output.n25 185
R23710 output.n73 output.n72 185
R23711 output.n71 output.n70 185
R23712 output.n50 output.n49 185
R23713 output.n65 output.n64 185
R23714 output.n63 output.n62 185
R23715 output.n54 output.n53 185
R23716 output.n57 output.n56 185
R23717 output.n105 output.n104 185
R23718 output.n103 output.n102 185
R23719 output.n82 output.n81 185
R23720 output.n97 output.n96 185
R23721 output.n95 output.n94 185
R23722 output.n86 output.n85 185
R23723 output.n89 output.n88 185
R23724 output.n137 output.n136 185
R23725 output.n135 output.n134 185
R23726 output.n114 output.n113 185
R23727 output.n129 output.n128 185
R23728 output.n127 output.n126 185
R23729 output.n118 output.n117 185
R23730 output.n121 output.n120 185
R23731 output.t2 output.n24 147.661
R23732 output.t1 output.n55 147.661
R23733 output.t3 output.n87 147.661
R23734 output.t0 output.n119 147.661
R23735 output.n41 output.n40 104.615
R23736 output.n40 output.n18 104.615
R23737 output.n33 output.n18 104.615
R23738 output.n33 output.n32 104.615
R23739 output.n32 output.n22 104.615
R23740 output.n25 output.n22 104.615
R23741 output.n72 output.n71 104.615
R23742 output.n71 output.n49 104.615
R23743 output.n64 output.n49 104.615
R23744 output.n64 output.n63 104.615
R23745 output.n63 output.n53 104.615
R23746 output.n56 output.n53 104.615
R23747 output.n104 output.n103 104.615
R23748 output.n103 output.n81 104.615
R23749 output.n96 output.n81 104.615
R23750 output.n96 output.n95 104.615
R23751 output.n95 output.n85 104.615
R23752 output.n88 output.n85 104.615
R23753 output.n136 output.n135 104.615
R23754 output.n135 output.n113 104.615
R23755 output.n128 output.n113 104.615
R23756 output.n128 output.n127 104.615
R23757 output.n127 output.n117 104.615
R23758 output.n120 output.n117 104.615
R23759 output.n1 output.t8 77.056
R23760 output.n14 output.t9 76.6694
R23761 output.n1 output.n0 72.7095
R23762 output.n3 output.n2 72.7095
R23763 output.n5 output.n4 72.7095
R23764 output.n7 output.n6 72.7095
R23765 output.n9 output.n8 72.7095
R23766 output.n11 output.n10 72.7095
R23767 output.n13 output.n12 72.7095
R23768 output.n25 output.t2 52.3082
R23769 output.n56 output.t1 52.3082
R23770 output.n88 output.t3 52.3082
R23771 output.n120 output.t0 52.3082
R23772 output.n26 output.n24 15.6674
R23773 output.n57 output.n55 15.6674
R23774 output.n89 output.n87 15.6674
R23775 output.n121 output.n119 15.6674
R23776 output.n27 output.n23 12.8005
R23777 output.n58 output.n54 12.8005
R23778 output.n90 output.n86 12.8005
R23779 output.n122 output.n118 12.8005
R23780 output.n31 output.n30 12.0247
R23781 output.n62 output.n61 12.0247
R23782 output.n94 output.n93 12.0247
R23783 output.n126 output.n125 12.0247
R23784 output.n34 output.n21 11.249
R23785 output.n65 output.n52 11.249
R23786 output.n97 output.n84 11.249
R23787 output.n129 output.n116 11.249
R23788 output.n35 output.n19 10.4732
R23789 output.n66 output.n50 10.4732
R23790 output.n98 output.n82 10.4732
R23791 output.n130 output.n114 10.4732
R23792 output.n39 output.n38 9.69747
R23793 output.n70 output.n69 9.69747
R23794 output.n102 output.n101 9.69747
R23795 output.n134 output.n133 9.69747
R23796 output.n45 output.n44 9.45567
R23797 output.n76 output.n75 9.45567
R23798 output.n108 output.n107 9.45567
R23799 output.n140 output.n139 9.45567
R23800 output.n44 output.n43 9.3005
R23801 output.n17 output.n16 9.3005
R23802 output.n38 output.n37 9.3005
R23803 output.n36 output.n35 9.3005
R23804 output.n21 output.n20 9.3005
R23805 output.n30 output.n29 9.3005
R23806 output.n28 output.n27 9.3005
R23807 output.n75 output.n74 9.3005
R23808 output.n48 output.n47 9.3005
R23809 output.n69 output.n68 9.3005
R23810 output.n67 output.n66 9.3005
R23811 output.n52 output.n51 9.3005
R23812 output.n61 output.n60 9.3005
R23813 output.n59 output.n58 9.3005
R23814 output.n107 output.n106 9.3005
R23815 output.n80 output.n79 9.3005
R23816 output.n101 output.n100 9.3005
R23817 output.n99 output.n98 9.3005
R23818 output.n84 output.n83 9.3005
R23819 output.n93 output.n92 9.3005
R23820 output.n91 output.n90 9.3005
R23821 output.n139 output.n138 9.3005
R23822 output.n112 output.n111 9.3005
R23823 output.n133 output.n132 9.3005
R23824 output.n131 output.n130 9.3005
R23825 output.n116 output.n115 9.3005
R23826 output.n125 output.n124 9.3005
R23827 output.n123 output.n122 9.3005
R23828 output.n42 output.n17 8.92171
R23829 output.n73 output.n48 8.92171
R23830 output.n105 output.n80 8.92171
R23831 output.n137 output.n112 8.92171
R23832 output output.n141 8.15037
R23833 output.n43 output.n15 8.14595
R23834 output.n74 output.n46 8.14595
R23835 output.n106 output.n78 8.14595
R23836 output.n138 output.n110 8.14595
R23837 output.n45 output.n15 5.81868
R23838 output.n76 output.n46 5.81868
R23839 output.n108 output.n78 5.81868
R23840 output.n140 output.n110 5.81868
R23841 output.n43 output.n42 5.04292
R23842 output.n74 output.n73 5.04292
R23843 output.n106 output.n105 5.04292
R23844 output.n138 output.n137 5.04292
R23845 output.n28 output.n24 4.38594
R23846 output.n59 output.n55 4.38594
R23847 output.n91 output.n87 4.38594
R23848 output.n123 output.n119 4.38594
R23849 output.n39 output.n17 4.26717
R23850 output.n70 output.n48 4.26717
R23851 output.n102 output.n80 4.26717
R23852 output.n134 output.n112 4.26717
R23853 output.n0 output.t14 3.9605
R23854 output.n0 output.t18 3.9605
R23855 output.n2 output.t5 3.9605
R23856 output.n2 output.t10 3.9605
R23857 output.n4 output.t11 3.9605
R23858 output.n4 output.t16 3.9605
R23859 output.n6 output.t4 3.9605
R23860 output.n6 output.t12 3.9605
R23861 output.n8 output.t15 3.9605
R23862 output.n8 output.t13 3.9605
R23863 output.n10 output.t19 3.9605
R23864 output.n10 output.t6 3.9605
R23865 output.n12 output.t7 3.9605
R23866 output.n12 output.t17 3.9605
R23867 output.n38 output.n19 3.49141
R23868 output.n69 output.n50 3.49141
R23869 output.n101 output.n82 3.49141
R23870 output.n133 output.n114 3.49141
R23871 output.n35 output.n34 2.71565
R23872 output.n66 output.n65 2.71565
R23873 output.n98 output.n97 2.71565
R23874 output.n130 output.n129 2.71565
R23875 output.n31 output.n21 1.93989
R23876 output.n62 output.n52 1.93989
R23877 output.n94 output.n84 1.93989
R23878 output.n126 output.n116 1.93989
R23879 output.n30 output.n23 1.16414
R23880 output.n61 output.n54 1.16414
R23881 output.n93 output.n86 1.16414
R23882 output.n125 output.n118 1.16414
R23883 output.n141 output.n109 0.962709
R23884 output.n109 output.n77 0.962709
R23885 output.n27 output.n26 0.388379
R23886 output.n58 output.n57 0.388379
R23887 output.n90 output.n89 0.388379
R23888 output.n122 output.n121 0.388379
R23889 output.n14 output.n13 0.387128
R23890 output.n13 output.n11 0.387128
R23891 output.n11 output.n9 0.387128
R23892 output.n9 output.n7 0.387128
R23893 output.n7 output.n5 0.387128
R23894 output.n5 output.n3 0.387128
R23895 output.n3 output.n1 0.387128
R23896 output.n44 output.n16 0.155672
R23897 output.n37 output.n16 0.155672
R23898 output.n37 output.n36 0.155672
R23899 output.n36 output.n20 0.155672
R23900 output.n29 output.n20 0.155672
R23901 output.n29 output.n28 0.155672
R23902 output.n75 output.n47 0.155672
R23903 output.n68 output.n47 0.155672
R23904 output.n68 output.n67 0.155672
R23905 output.n67 output.n51 0.155672
R23906 output.n60 output.n51 0.155672
R23907 output.n60 output.n59 0.155672
R23908 output.n107 output.n79 0.155672
R23909 output.n100 output.n79 0.155672
R23910 output.n100 output.n99 0.155672
R23911 output.n99 output.n83 0.155672
R23912 output.n92 output.n83 0.155672
R23913 output.n92 output.n91 0.155672
R23914 output.n139 output.n111 0.155672
R23915 output.n132 output.n111 0.155672
R23916 output.n132 output.n131 0.155672
R23917 output.n131 output.n115 0.155672
R23918 output.n124 output.n115 0.155672
R23919 output.n124 output.n123 0.155672
R23920 output output.n14 0.126227
C0 minus commonsourceibias 0.332601f
C1 plus commonsourceibias 0.278362f
C2 output outputibias 2.34152f
C3 vdd output 7.23429f
C4 CSoutput output 6.13881f
C5 CSoutput outputibias 0.032386f
C6 vdd CSoutput 0.140616p
C7 commonsourceibias output 0.006808f
C8 minus diffpairibias 3.4e-19
C9 CSoutput minus 3.00028f
C10 vdd plus 0.089709f
C11 plus diffpairibias 3.42e-19
C12 commonsourceibias outputibias 0.003832f
C13 vdd commonsourceibias 0.004218f
C14 CSoutput plus 0.876209f
C15 commonsourceibias diffpairibias 0.064336f
C16 CSoutput commonsourceibias 54.554f
C17 minus plus 9.55573f
C18 diffpairibias gnd 60.00273f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.18415p
C22 plus gnd 34.301804f
C23 minus gnd 28.74923f
C24 CSoutput gnd 0.12625p
C25 vdd gnd 0.439015p
C26 output.t8 gnd 0.464308f
C27 output.t14 gnd 0.044422f
C28 output.t18 gnd 0.044422f
C29 output.n0 gnd 0.364624f
C30 output.n1 gnd 0.614102f
C31 output.t5 gnd 0.044422f
C32 output.t10 gnd 0.044422f
C33 output.n2 gnd 0.364624f
C34 output.n3 gnd 0.350265f
C35 output.t11 gnd 0.044422f
C36 output.t16 gnd 0.044422f
C37 output.n4 gnd 0.364624f
C38 output.n5 gnd 0.350265f
C39 output.t4 gnd 0.044422f
C40 output.t12 gnd 0.044422f
C41 output.n6 gnd 0.364624f
C42 output.n7 gnd 0.350265f
C43 output.t15 gnd 0.044422f
C44 output.t13 gnd 0.044422f
C45 output.n8 gnd 0.364624f
C46 output.n9 gnd 0.350265f
C47 output.t19 gnd 0.044422f
C48 output.t6 gnd 0.044422f
C49 output.n10 gnd 0.364624f
C50 output.n11 gnd 0.350265f
C51 output.t7 gnd 0.044422f
C52 output.t17 gnd 0.044422f
C53 output.n12 gnd 0.364624f
C54 output.n13 gnd 0.350265f
C55 output.t9 gnd 0.462979f
C56 output.n14 gnd 0.28994f
C57 output.n15 gnd 0.015803f
C58 output.n16 gnd 0.011243f
C59 output.n17 gnd 0.006041f
C60 output.n18 gnd 0.01428f
C61 output.n19 gnd 0.006397f
C62 output.n20 gnd 0.011243f
C63 output.n21 gnd 0.006041f
C64 output.n22 gnd 0.01428f
C65 output.n23 gnd 0.006397f
C66 output.n24 gnd 0.048111f
C67 output.t2 gnd 0.023274f
C68 output.n25 gnd 0.01071f
C69 output.n26 gnd 0.008435f
C70 output.n27 gnd 0.006041f
C71 output.n28 gnd 0.267512f
C72 output.n29 gnd 0.011243f
C73 output.n30 gnd 0.006041f
C74 output.n31 gnd 0.006397f
C75 output.n32 gnd 0.01428f
C76 output.n33 gnd 0.01428f
C77 output.n34 gnd 0.006397f
C78 output.n35 gnd 0.006041f
C79 output.n36 gnd 0.011243f
C80 output.n37 gnd 0.011243f
C81 output.n38 gnd 0.006041f
C82 output.n39 gnd 0.006397f
C83 output.n40 gnd 0.01428f
C84 output.n41 gnd 0.030913f
C85 output.n42 gnd 0.006397f
C86 output.n43 gnd 0.006041f
C87 output.n44 gnd 0.025987f
C88 output.n45 gnd 0.097665f
C89 output.n46 gnd 0.015803f
C90 output.n47 gnd 0.011243f
C91 output.n48 gnd 0.006041f
C92 output.n49 gnd 0.01428f
C93 output.n50 gnd 0.006397f
C94 output.n51 gnd 0.011243f
C95 output.n52 gnd 0.006041f
C96 output.n53 gnd 0.01428f
C97 output.n54 gnd 0.006397f
C98 output.n55 gnd 0.048111f
C99 output.t1 gnd 0.023274f
C100 output.n56 gnd 0.01071f
C101 output.n57 gnd 0.008435f
C102 output.n58 gnd 0.006041f
C103 output.n59 gnd 0.267512f
C104 output.n60 gnd 0.011243f
C105 output.n61 gnd 0.006041f
C106 output.n62 gnd 0.006397f
C107 output.n63 gnd 0.01428f
C108 output.n64 gnd 0.01428f
C109 output.n65 gnd 0.006397f
C110 output.n66 gnd 0.006041f
C111 output.n67 gnd 0.011243f
C112 output.n68 gnd 0.011243f
C113 output.n69 gnd 0.006041f
C114 output.n70 gnd 0.006397f
C115 output.n71 gnd 0.01428f
C116 output.n72 gnd 0.030913f
C117 output.n73 gnd 0.006397f
C118 output.n74 gnd 0.006041f
C119 output.n75 gnd 0.025987f
C120 output.n76 gnd 0.09306f
C121 output.n77 gnd 1.65264f
C122 output.n78 gnd 0.015803f
C123 output.n79 gnd 0.011243f
C124 output.n80 gnd 0.006041f
C125 output.n81 gnd 0.01428f
C126 output.n82 gnd 0.006397f
C127 output.n83 gnd 0.011243f
C128 output.n84 gnd 0.006041f
C129 output.n85 gnd 0.01428f
C130 output.n86 gnd 0.006397f
C131 output.n87 gnd 0.048111f
C132 output.t3 gnd 0.023274f
C133 output.n88 gnd 0.01071f
C134 output.n89 gnd 0.008435f
C135 output.n90 gnd 0.006041f
C136 output.n91 gnd 0.267512f
C137 output.n92 gnd 0.011243f
C138 output.n93 gnd 0.006041f
C139 output.n94 gnd 0.006397f
C140 output.n95 gnd 0.01428f
C141 output.n96 gnd 0.01428f
C142 output.n97 gnd 0.006397f
C143 output.n98 gnd 0.006041f
C144 output.n99 gnd 0.011243f
C145 output.n100 gnd 0.011243f
C146 output.n101 gnd 0.006041f
C147 output.n102 gnd 0.006397f
C148 output.n103 gnd 0.01428f
C149 output.n104 gnd 0.030913f
C150 output.n105 gnd 0.006397f
C151 output.n106 gnd 0.006041f
C152 output.n107 gnd 0.025987f
C153 output.n108 gnd 0.09306f
C154 output.n109 gnd 0.713089f
C155 output.n110 gnd 0.015803f
C156 output.n111 gnd 0.011243f
C157 output.n112 gnd 0.006041f
C158 output.n113 gnd 0.01428f
C159 output.n114 gnd 0.006397f
C160 output.n115 gnd 0.011243f
C161 output.n116 gnd 0.006041f
C162 output.n117 gnd 0.01428f
C163 output.n118 gnd 0.006397f
C164 output.n119 gnd 0.048111f
C165 output.t0 gnd 0.023274f
C166 output.n120 gnd 0.01071f
C167 output.n121 gnd 0.008435f
C168 output.n122 gnd 0.006041f
C169 output.n123 gnd 0.267512f
C170 output.n124 gnd 0.011243f
C171 output.n125 gnd 0.006041f
C172 output.n126 gnd 0.006397f
C173 output.n127 gnd 0.01428f
C174 output.n128 gnd 0.01428f
C175 output.n129 gnd 0.006397f
C176 output.n130 gnd 0.006041f
C177 output.n131 gnd 0.011243f
C178 output.n132 gnd 0.011243f
C179 output.n133 gnd 0.006041f
C180 output.n134 gnd 0.006397f
C181 output.n135 gnd 0.01428f
C182 output.n136 gnd 0.030913f
C183 output.n137 gnd 0.006397f
C184 output.n138 gnd 0.006041f
C185 output.n139 gnd 0.025987f
C186 output.n140 gnd 0.09306f
C187 output.n141 gnd 1.67353f
C188 outputibias.t10 gnd 0.11477f
C189 outputibias.t9 gnd 0.115567f
C190 outputibias.n0 gnd 0.130108f
C191 outputibias.n1 gnd 0.001372f
C192 outputibias.n2 gnd 9.76e-19
C193 outputibias.n3 gnd 5.24e-19
C194 outputibias.n4 gnd 0.001239f
C195 outputibias.n5 gnd 5.55e-19
C196 outputibias.n6 gnd 9.76e-19
C197 outputibias.n7 gnd 5.24e-19
C198 outputibias.n8 gnd 0.001239f
C199 outputibias.n9 gnd 5.55e-19
C200 outputibias.n10 gnd 0.004176f
C201 outputibias.t5 gnd 0.00202f
C202 outputibias.n11 gnd 9.3e-19
C203 outputibias.n12 gnd 7.32e-19
C204 outputibias.n13 gnd 5.24e-19
C205 outputibias.n14 gnd 0.02322f
C206 outputibias.n15 gnd 9.76e-19
C207 outputibias.n16 gnd 5.24e-19
C208 outputibias.n17 gnd 5.55e-19
C209 outputibias.n18 gnd 0.001239f
C210 outputibias.n19 gnd 0.001239f
C211 outputibias.n20 gnd 5.55e-19
C212 outputibias.n21 gnd 5.24e-19
C213 outputibias.n22 gnd 9.76e-19
C214 outputibias.n23 gnd 9.76e-19
C215 outputibias.n24 gnd 5.24e-19
C216 outputibias.n25 gnd 5.55e-19
C217 outputibias.n26 gnd 0.001239f
C218 outputibias.n27 gnd 0.002683f
C219 outputibias.n28 gnd 5.55e-19
C220 outputibias.n29 gnd 5.24e-19
C221 outputibias.n30 gnd 0.002256f
C222 outputibias.n31 gnd 0.005781f
C223 outputibias.n32 gnd 0.001372f
C224 outputibias.n33 gnd 9.76e-19
C225 outputibias.n34 gnd 5.24e-19
C226 outputibias.n35 gnd 0.001239f
C227 outputibias.n36 gnd 5.55e-19
C228 outputibias.n37 gnd 9.76e-19
C229 outputibias.n38 gnd 5.24e-19
C230 outputibias.n39 gnd 0.001239f
C231 outputibias.n40 gnd 5.55e-19
C232 outputibias.n41 gnd 0.004176f
C233 outputibias.t7 gnd 0.00202f
C234 outputibias.n42 gnd 9.3e-19
C235 outputibias.n43 gnd 7.32e-19
C236 outputibias.n44 gnd 5.24e-19
C237 outputibias.n45 gnd 0.02322f
C238 outputibias.n46 gnd 9.76e-19
C239 outputibias.n47 gnd 5.24e-19
C240 outputibias.n48 gnd 5.55e-19
C241 outputibias.n49 gnd 0.001239f
C242 outputibias.n50 gnd 0.001239f
C243 outputibias.n51 gnd 5.55e-19
C244 outputibias.n52 gnd 5.24e-19
C245 outputibias.n53 gnd 9.76e-19
C246 outputibias.n54 gnd 9.76e-19
C247 outputibias.n55 gnd 5.24e-19
C248 outputibias.n56 gnd 5.55e-19
C249 outputibias.n57 gnd 0.001239f
C250 outputibias.n58 gnd 0.002683f
C251 outputibias.n59 gnd 5.55e-19
C252 outputibias.n60 gnd 5.24e-19
C253 outputibias.n61 gnd 0.002256f
C254 outputibias.n62 gnd 0.005197f
C255 outputibias.n63 gnd 0.121892f
C256 outputibias.n64 gnd 0.001372f
C257 outputibias.n65 gnd 9.76e-19
C258 outputibias.n66 gnd 5.24e-19
C259 outputibias.n67 gnd 0.001239f
C260 outputibias.n68 gnd 5.55e-19
C261 outputibias.n69 gnd 9.76e-19
C262 outputibias.n70 gnd 5.24e-19
C263 outputibias.n71 gnd 0.001239f
C264 outputibias.n72 gnd 5.55e-19
C265 outputibias.n73 gnd 0.004176f
C266 outputibias.t1 gnd 0.00202f
C267 outputibias.n74 gnd 9.3e-19
C268 outputibias.n75 gnd 7.32e-19
C269 outputibias.n76 gnd 5.24e-19
C270 outputibias.n77 gnd 0.02322f
C271 outputibias.n78 gnd 9.76e-19
C272 outputibias.n79 gnd 5.24e-19
C273 outputibias.n80 gnd 5.55e-19
C274 outputibias.n81 gnd 0.001239f
C275 outputibias.n82 gnd 0.001239f
C276 outputibias.n83 gnd 5.55e-19
C277 outputibias.n84 gnd 5.24e-19
C278 outputibias.n85 gnd 9.76e-19
C279 outputibias.n86 gnd 9.76e-19
C280 outputibias.n87 gnd 5.24e-19
C281 outputibias.n88 gnd 5.55e-19
C282 outputibias.n89 gnd 0.001239f
C283 outputibias.n90 gnd 0.002683f
C284 outputibias.n91 gnd 5.55e-19
C285 outputibias.n92 gnd 5.24e-19
C286 outputibias.n93 gnd 0.002256f
C287 outputibias.n94 gnd 0.005197f
C288 outputibias.n95 gnd 0.064513f
C289 outputibias.n96 gnd 0.001372f
C290 outputibias.n97 gnd 9.76e-19
C291 outputibias.n98 gnd 5.24e-19
C292 outputibias.n99 gnd 0.001239f
C293 outputibias.n100 gnd 5.55e-19
C294 outputibias.n101 gnd 9.76e-19
C295 outputibias.n102 gnd 5.24e-19
C296 outputibias.n103 gnd 0.001239f
C297 outputibias.n104 gnd 5.55e-19
C298 outputibias.n105 gnd 0.004176f
C299 outputibias.t3 gnd 0.00202f
C300 outputibias.n106 gnd 9.3e-19
C301 outputibias.n107 gnd 7.32e-19
C302 outputibias.n108 gnd 5.24e-19
C303 outputibias.n109 gnd 0.02322f
C304 outputibias.n110 gnd 9.76e-19
C305 outputibias.n111 gnd 5.24e-19
C306 outputibias.n112 gnd 5.55e-19
C307 outputibias.n113 gnd 0.001239f
C308 outputibias.n114 gnd 0.001239f
C309 outputibias.n115 gnd 5.55e-19
C310 outputibias.n116 gnd 5.24e-19
C311 outputibias.n117 gnd 9.76e-19
C312 outputibias.n118 gnd 9.76e-19
C313 outputibias.n119 gnd 5.24e-19
C314 outputibias.n120 gnd 5.55e-19
C315 outputibias.n121 gnd 0.001239f
C316 outputibias.n122 gnd 0.002683f
C317 outputibias.n123 gnd 5.55e-19
C318 outputibias.n124 gnd 5.24e-19
C319 outputibias.n125 gnd 0.002256f
C320 outputibias.n126 gnd 0.005197f
C321 outputibias.n127 gnd 0.084814f
C322 outputibias.t2 gnd 0.108319f
C323 outputibias.t0 gnd 0.108319f
C324 outputibias.t6 gnd 0.108319f
C325 outputibias.t4 gnd 0.109238f
C326 outputibias.n128 gnd 0.134674f
C327 outputibias.n129 gnd 0.07244f
C328 outputibias.n130 gnd 0.079818f
C329 outputibias.n131 gnd 0.164901f
C330 outputibias.t11 gnd 0.11477f
C331 outputibias.n132 gnd 0.067481f
C332 outputibias.t8 gnd 0.11477f
C333 outputibias.n133 gnd 0.065115f
C334 outputibias.n134 gnd 0.029159f
C335 a_n1986_8322.t21 gnd 49.3316f
C336 a_n1986_8322.t20 gnd 76.0671f
C337 a_n1986_8322.t10 gnd 0.093483f
C338 a_n1986_8322.t9 gnd 0.875324f
C339 a_n1986_8322.t17 gnd 0.093483f
C340 a_n1986_8322.t12 gnd 0.093483f
C341 a_n1986_8322.n0 gnd 0.658492f
C342 a_n1986_8322.n1 gnd 0.735768f
C343 a_n1986_8322.t15 gnd 0.093483f
C344 a_n1986_8322.t14 gnd 0.093483f
C345 a_n1986_8322.n2 gnd 0.658492f
C346 a_n1986_8322.n3 gnd 0.373834f
C347 a_n1986_8322.t8 gnd 0.873581f
C348 a_n1986_8322.n4 gnd 1.39821f
C349 a_n1986_8322.t3 gnd 0.875324f
C350 a_n1986_8322.t7 gnd 0.093483f
C351 a_n1986_8322.t6 gnd 0.093483f
C352 a_n1986_8322.n5 gnd 0.658492f
C353 a_n1986_8322.n6 gnd 0.735768f
C354 a_n1986_8322.t1 gnd 0.873581f
C355 a_n1986_8322.n7 gnd 0.370248f
C356 a_n1986_8322.t4 gnd 0.873581f
C357 a_n1986_8322.n8 gnd 0.370248f
C358 a_n1986_8322.t2 gnd 0.093483f
C359 a_n1986_8322.t0 gnd 0.093483f
C360 a_n1986_8322.n9 gnd 0.658492f
C361 a_n1986_8322.n10 gnd 0.373834f
C362 a_n1986_8322.t5 gnd 0.873581f
C363 a_n1986_8322.n11 gnd 0.871851f
C364 a_n1986_8322.n12 gnd 1.58986f
C365 a_n1986_8322.n13 gnd 3.73938f
C366 a_n1986_8322.t11 gnd 0.873581f
C367 a_n1986_8322.n14 gnd 0.766111f
C368 a_n1986_8322.t18 gnd 0.875322f
C369 a_n1986_8322.t16 gnd 0.093483f
C370 a_n1986_8322.t13 gnd 0.093483f
C371 a_n1986_8322.n15 gnd 0.658492f
C372 a_n1986_8322.n16 gnd 0.73577f
C373 a_n1986_8322.n17 gnd 0.373832f
C374 a_n1986_8322.n18 gnd 0.658494f
C375 a_n1986_8322.t19 gnd 0.093483f
C376 minus.n0 gnd 0.031208f
C377 minus.n1 gnd 0.007082f
C378 minus.n2 gnd 0.031208f
C379 minus.n3 gnd 0.007082f
C380 minus.n4 gnd 0.031208f
C381 minus.n5 gnd 0.007082f
C382 minus.n6 gnd 0.031208f
C383 minus.n7 gnd 0.007082f
C384 minus.t8 gnd 0.45688f
C385 minus.t7 gnd 0.441415f
C386 minus.n8 gnd 0.201311f
C387 minus.n9 gnd 0.182867f
C388 minus.n10 gnd 0.133211f
C389 minus.n11 gnd 0.031208f
C390 minus.t11 gnd 0.441415f
C391 minus.n12 gnd 0.196091f
C392 minus.n13 gnd 0.007082f
C393 minus.t10 gnd 0.441415f
C394 minus.n14 gnd 0.196091f
C395 minus.n15 gnd 0.031208f
C396 minus.n16 gnd 0.031208f
C397 minus.n17 gnd 0.031208f
C398 minus.t12 gnd 0.441415f
C399 minus.n18 gnd 0.196091f
C400 minus.n19 gnd 0.007082f
C401 minus.t17 gnd 0.441415f
C402 minus.n20 gnd 0.196091f
C403 minus.n21 gnd 0.031208f
C404 minus.n22 gnd 0.031208f
C405 minus.n23 gnd 0.031208f
C406 minus.t16 gnd 0.441415f
C407 minus.n24 gnd 0.196091f
C408 minus.n25 gnd 0.007082f
C409 minus.t21 gnd 0.441415f
C410 minus.n26 gnd 0.196091f
C411 minus.n27 gnd 0.031208f
C412 minus.n28 gnd 0.031208f
C413 minus.n29 gnd 0.031208f
C414 minus.t20 gnd 0.441415f
C415 minus.n30 gnd 0.196091f
C416 minus.n31 gnd 0.007082f
C417 minus.t13 gnd 0.441415f
C418 minus.n32 gnd 0.195802f
C419 minus.n33 gnd 0.36059f
C420 minus.n34 gnd 0.031208f
C421 minus.t5 gnd 0.441415f
C422 minus.t6 gnd 0.441415f
C423 minus.n35 gnd 0.031208f
C424 minus.t22 gnd 0.441415f
C425 minus.n36 gnd 0.196091f
C426 minus.n37 gnd 0.031208f
C427 minus.t18 gnd 0.441415f
C428 minus.t19 gnd 0.441415f
C429 minus.n38 gnd 0.196091f
C430 minus.n39 gnd 0.031208f
C431 minus.t14 gnd 0.441415f
C432 minus.t15 gnd 0.441415f
C433 minus.n40 gnd 0.196091f
C434 minus.n41 gnd 0.031208f
C435 minus.t9 gnd 0.441415f
C436 minus.t23 gnd 0.441415f
C437 minus.n42 gnd 0.201311f
C438 minus.t24 gnd 0.45688f
C439 minus.n43 gnd 0.182867f
C440 minus.n44 gnd 0.133211f
C441 minus.n45 gnd 0.007082f
C442 minus.n46 gnd 0.196091f
C443 minus.n47 gnd 0.007082f
C444 minus.n48 gnd 0.031208f
C445 minus.n49 gnd 0.031208f
C446 minus.n50 gnd 0.031208f
C447 minus.n51 gnd 0.007082f
C448 minus.n52 gnd 0.196091f
C449 minus.n53 gnd 0.007082f
C450 minus.n54 gnd 0.031208f
C451 minus.n55 gnd 0.031208f
C452 minus.n56 gnd 0.031208f
C453 minus.n57 gnd 0.007082f
C454 minus.n58 gnd 0.196091f
C455 minus.n59 gnd 0.007082f
C456 minus.n60 gnd 0.031208f
C457 minus.n61 gnd 0.031208f
C458 minus.n62 gnd 0.031208f
C459 minus.n63 gnd 0.007082f
C460 minus.n64 gnd 0.196091f
C461 minus.n65 gnd 0.007082f
C462 minus.n66 gnd 0.195802f
C463 minus.n67 gnd 0.975177f
C464 minus.n68 gnd 1.46812f
C465 minus.t2 gnd 0.009621f
C466 minus.t0 gnd 0.009621f
C467 minus.n69 gnd 0.031635f
C468 minus.t3 gnd 0.009621f
C469 minus.t1 gnd 0.009621f
C470 minus.n70 gnd 0.031202f
C471 minus.n71 gnd 0.266291f
C472 minus.t4 gnd 0.053548f
C473 minus.n72 gnd 0.145312f
C474 minus.n73 gnd 2.16209f
C475 diffpairibias.t27 gnd 0.090128f
C476 diffpairibias.t23 gnd 0.08996f
C477 diffpairibias.n0 gnd 0.105991f
C478 diffpairibias.t28 gnd 0.08996f
C479 diffpairibias.n1 gnd 0.051736f
C480 diffpairibias.t25 gnd 0.08996f
C481 diffpairibias.n2 gnd 0.051736f
C482 diffpairibias.t29 gnd 0.08996f
C483 diffpairibias.n3 gnd 0.041084f
C484 diffpairibias.t15 gnd 0.086371f
C485 diffpairibias.t1 gnd 0.085993f
C486 diffpairibias.n4 gnd 0.13579f
C487 diffpairibias.t11 gnd 0.085993f
C488 diffpairibias.n5 gnd 0.072463f
C489 diffpairibias.t13 gnd 0.085993f
C490 diffpairibias.n6 gnd 0.072463f
C491 diffpairibias.t7 gnd 0.085993f
C492 diffpairibias.n7 gnd 0.072463f
C493 diffpairibias.t3 gnd 0.085993f
C494 diffpairibias.n8 gnd 0.072463f
C495 diffpairibias.t17 gnd 0.085993f
C496 diffpairibias.n9 gnd 0.072463f
C497 diffpairibias.t5 gnd 0.085993f
C498 diffpairibias.n10 gnd 0.072463f
C499 diffpairibias.t19 gnd 0.085993f
C500 diffpairibias.n11 gnd 0.072463f
C501 diffpairibias.t9 gnd 0.085993f
C502 diffpairibias.n12 gnd 0.102883f
C503 diffpairibias.t14 gnd 0.086899f
C504 diffpairibias.t0 gnd 0.086748f
C505 diffpairibias.n13 gnd 0.094648f
C506 diffpairibias.t10 gnd 0.086748f
C507 diffpairibias.n14 gnd 0.052262f
C508 diffpairibias.t12 gnd 0.086748f
C509 diffpairibias.n15 gnd 0.052262f
C510 diffpairibias.t6 gnd 0.086748f
C511 diffpairibias.n16 gnd 0.052262f
C512 diffpairibias.t2 gnd 0.086748f
C513 diffpairibias.n17 gnd 0.052262f
C514 diffpairibias.t16 gnd 0.086748f
C515 diffpairibias.n18 gnd 0.052262f
C516 diffpairibias.t4 gnd 0.086748f
C517 diffpairibias.n19 gnd 0.052262f
C518 diffpairibias.t18 gnd 0.086748f
C519 diffpairibias.n20 gnd 0.052262f
C520 diffpairibias.t8 gnd 0.086748f
C521 diffpairibias.n21 gnd 0.061849f
C522 diffpairibias.n22 gnd 0.233513f
C523 diffpairibias.t20 gnd 0.08996f
C524 diffpairibias.n23 gnd 0.051747f
C525 diffpairibias.t26 gnd 0.08996f
C526 diffpairibias.n24 gnd 0.051736f
C527 diffpairibias.t22 gnd 0.08996f
C528 diffpairibias.n25 gnd 0.051736f
C529 diffpairibias.t21 gnd 0.08996f
C530 diffpairibias.n26 gnd 0.051736f
C531 diffpairibias.t24 gnd 0.08996f
C532 diffpairibias.n27 gnd 0.04729f
C533 diffpairibias.n28 gnd 0.047711f
C534 a_n1808_13878.t17 gnd 0.185195f
C535 a_n1808_13878.t15 gnd 0.185195f
C536 a_n1808_13878.t19 gnd 0.185195f
C537 a_n1808_13878.n0 gnd 1.46067f
C538 a_n1808_13878.t8 gnd 0.185195f
C539 a_n1808_13878.t13 gnd 0.185195f
C540 a_n1808_13878.n1 gnd 1.45825f
C541 a_n1808_13878.n2 gnd 1.31079f
C542 a_n1808_13878.t10 gnd 0.185195f
C543 a_n1808_13878.t12 gnd 0.185195f
C544 a_n1808_13878.n3 gnd 1.4598f
C545 a_n1808_13878.t16 gnd 0.185195f
C546 a_n1808_13878.t11 gnd 0.185195f
C547 a_n1808_13878.n4 gnd 1.45825f
C548 a_n1808_13878.n5 gnd 2.03762f
C549 a_n1808_13878.t14 gnd 0.185195f
C550 a_n1808_13878.t9 gnd 0.185195f
C551 a_n1808_13878.n6 gnd 1.45825f
C552 a_n1808_13878.n7 gnd 3.69301f
C553 a_n1808_13878.t1 gnd 1.73408f
C554 a_n1808_13878.t4 gnd 0.185195f
C555 a_n1808_13878.t5 gnd 0.185195f
C556 a_n1808_13878.n8 gnd 1.30452f
C557 a_n1808_13878.n9 gnd 1.4576f
C558 a_n1808_13878.t0 gnd 1.73062f
C559 a_n1808_13878.n10 gnd 0.733487f
C560 a_n1808_13878.t3 gnd 1.73062f
C561 a_n1808_13878.n11 gnd 0.733487f
C562 a_n1808_13878.t6 gnd 0.185195f
C563 a_n1808_13878.t7 gnd 0.185195f
C564 a_n1808_13878.n12 gnd 1.30452f
C565 a_n1808_13878.n13 gnd 0.74059f
C566 a_n1808_13878.t2 gnd 1.73062f
C567 a_n1808_13878.n14 gnd 1.7272f
C568 a_n1808_13878.n15 gnd 2.51438f
C569 a_n1808_13878.n16 gnd 1.80025f
C570 a_n1808_13878.n17 gnd 1.45826f
C571 a_n1808_13878.t18 gnd 0.185195f
C572 a_n1996_n452.n0 gnd 0.822727f
C573 a_n1996_n452.n1 gnd 3.34433f
C574 a_n1996_n452.n2 gnd 3.17111f
C575 a_n1996_n452.n3 gnd 3.91594f
C576 a_n1996_n452.n4 gnd 0.527811f
C577 a_n1996_n452.n5 gnd 0.205584f
C578 a_n1996_n452.n6 gnd 0.151417f
C579 a_n1996_n452.n7 gnd 0.237979f
C580 a_n1996_n452.n8 gnd 0.183812f
C581 a_n1996_n452.n9 gnd 0.205584f
C582 a_n1996_n452.n10 gnd 0.151417f
C583 a_n1996_n452.n11 gnd 0.581979f
C584 a_n1996_n452.n12 gnd 0.433746f
C585 a_n1996_n452.n13 gnd 0.21667f
C586 a_n1996_n452.n14 gnd 0.494132f
C587 a_n1996_n452.n15 gnd 0.283464f
C588 a_n1996_n452.n16 gnd 0.439964f
C589 a_n1996_n452.n17 gnd 0.21667f
C590 a_n1996_n452.n18 gnd 0.734001f
C591 a_n1996_n452.n19 gnd 0.283464f
C592 a_n1996_n452.n20 gnd 0.641354f
C593 a_n1996_n452.n21 gnd 0.283464f
C594 a_n1996_n452.n22 gnd 0.494132f
C595 a_n1996_n452.n23 gnd 0.666675f
C596 a_n1996_n452.n24 gnd 0.21667f
C597 a_n1996_n452.n25 gnd 0.283464f
C598 a_n1996_n452.n26 gnd 1.78382f
C599 a_n1996_n452.n27 gnd 1.92214f
C600 a_n1996_n452.n28 gnd 3.22512f
C601 a_n1996_n452.n29 gnd 0.008389f
C602 a_n1996_n452.n31 gnd 1.34296f
C603 a_n1996_n452.n32 gnd 0.286629f
C604 a_n1996_n452.n33 gnd 0.108335f
C605 a_n1996_n452.n34 gnd 0.008389f
C606 a_n1996_n452.n36 gnd 0.008389f
C607 a_n1996_n452.n38 gnd 0.286629f
C608 a_n1996_n452.n39 gnd 0.008389f
C609 a_n1996_n452.n41 gnd 0.286629f
C610 a_n1996_n452.n42 gnd 0.008389f
C611 a_n1996_n452.n43 gnd 0.286221f
C612 a_n1996_n452.n44 gnd 0.008389f
C613 a_n1996_n452.n45 gnd 0.286221f
C614 a_n1996_n452.n46 gnd 0.008389f
C615 a_n1996_n452.n47 gnd 0.286221f
C616 a_n1996_n452.n48 gnd 0.008389f
C617 a_n1996_n452.n49 gnd 0.286221f
C618 a_n1996_n452.n50 gnd 0.286629f
C619 a_n1996_n452.t37 gnd 0.150285f
C620 a_n1996_n452.t27 gnd 1.40719f
C621 a_n1996_n452.t32 gnd 0.699053f
C622 a_n1996_n452.n51 gnd 0.307348f
C623 a_n1996_n452.t34 gnd 0.699053f
C624 a_n1996_n452.t36 gnd 0.699053f
C625 a_n1996_n452.t52 gnd 0.699053f
C626 a_n1996_n452.n52 gnd 0.307348f
C627 a_n1996_n452.t60 gnd 0.699053f
C628 a_n1996_n452.t66 gnd 0.699053f
C629 a_n1996_n452.t24 gnd 0.713776f
C630 a_n1996_n452.t28 gnd 0.699053f
C631 a_n1996_n452.t30 gnd 0.699053f
C632 a_n1996_n452.t18 gnd 0.699053f
C633 a_n1996_n452.n53 gnd 0.307348f
C634 a_n1996_n452.t20 gnd 0.699053f
C635 a_n1996_n452.t22 gnd 0.710611f
C636 a_n1996_n452.t39 gnd 0.116888f
C637 a_n1996_n452.t13 gnd 0.116888f
C638 a_n1996_n452.n54 gnd 1.03516f
C639 a_n1996_n452.t43 gnd 0.116888f
C640 a_n1996_n452.t40 gnd 0.116888f
C641 a_n1996_n452.n55 gnd 1.03287f
C642 a_n1996_n452.t9 gnd 0.116888f
C643 a_n1996_n452.t1 gnd 0.116888f
C644 a_n1996_n452.n56 gnd 1.03287f
C645 a_n1996_n452.t7 gnd 0.116888f
C646 a_n1996_n452.t12 gnd 0.116888f
C647 a_n1996_n452.n57 gnd 1.03516f
C648 a_n1996_n452.t3 gnd 0.116888f
C649 a_n1996_n452.t4 gnd 0.116888f
C650 a_n1996_n452.n58 gnd 1.03287f
C651 a_n1996_n452.t8 gnd 0.116888f
C652 a_n1996_n452.t6 gnd 0.116888f
C653 a_n1996_n452.n59 gnd 1.03287f
C654 a_n1996_n452.t11 gnd 0.116888f
C655 a_n1996_n452.t41 gnd 0.116888f
C656 a_n1996_n452.n60 gnd 1.03287f
C657 a_n1996_n452.t10 gnd 0.116888f
C658 a_n1996_n452.t38 gnd 0.116888f
C659 a_n1996_n452.n61 gnd 1.03287f
C660 a_n1996_n452.t2 gnd 0.116888f
C661 a_n1996_n452.t5 gnd 0.116888f
C662 a_n1996_n452.n62 gnd 1.03516f
C663 a_n1996_n452.t0 gnd 0.116888f
C664 a_n1996_n452.t42 gnd 0.116888f
C665 a_n1996_n452.n63 gnd 1.03287f
C666 a_n1996_n452.t70 gnd 0.713776f
C667 a_n1996_n452.t53 gnd 0.699053f
C668 a_n1996_n452.t57 gnd 0.699053f
C669 a_n1996_n452.t47 gnd 0.699053f
C670 a_n1996_n452.n64 gnd 0.307348f
C671 a_n1996_n452.t62 gnd 0.699053f
C672 a_n1996_n452.t68 gnd 0.710611f
C673 a_n1996_n452.n65 gnd 0.309974f
C674 a_n1996_n452.n66 gnd 0.303445f
C675 a_n1996_n452.n67 gnd 0.309973f
C676 a_n1996_n452.n68 gnd 0.309974f
C677 a_n1996_n452.n69 gnd 0.303445f
C678 a_n1996_n452.n70 gnd 0.309973f
C679 a_n1996_n452.t23 gnd 1.40719f
C680 a_n1996_n452.t19 gnd 0.150285f
C681 a_n1996_n452.t21 gnd 0.150285f
C682 a_n1996_n452.n71 gnd 1.05861f
C683 a_n1996_n452.t29 gnd 0.150285f
C684 a_n1996_n452.t31 gnd 0.150285f
C685 a_n1996_n452.n72 gnd 1.05861f
C686 a_n1996_n452.t25 gnd 1.40439f
C687 a_n1996_n452.n73 gnd 1.14844f
C688 a_n1996_n452.n74 gnd 0.789587f
C689 a_n1996_n452.t51 gnd 0.699053f
C690 a_n1996_n452.t61 gnd 0.699053f
C691 a_n1996_n452.t71 gnd 0.699053f
C692 a_n1996_n452.n75 gnd 0.307348f
C693 a_n1996_n452.t63 gnd 0.699053f
C694 a_n1996_n452.t48 gnd 0.699053f
C695 a_n1996_n452.t49 gnd 0.699053f
C696 a_n1996_n452.n76 gnd 0.307348f
C697 a_n1996_n452.t67 gnd 0.699053f
C698 a_n1996_n452.t56 gnd 0.699053f
C699 a_n1996_n452.t55 gnd 0.699053f
C700 a_n1996_n452.n77 gnd 0.307348f
C701 a_n1996_n452.t59 gnd 0.699053f
C702 a_n1996_n452.t50 gnd 0.699053f
C703 a_n1996_n452.t44 gnd 0.699053f
C704 a_n1996_n452.n78 gnd 0.307348f
C705 a_n1996_n452.t64 gnd 0.710766f
C706 a_n1996_n452.n79 gnd 0.303445f
C707 a_n1996_n452.n80 gnd 0.297934f
C708 a_n1996_n452.t69 gnd 0.710766f
C709 a_n1996_n452.n81 gnd 0.303445f
C710 a_n1996_n452.n82 gnd 0.297934f
C711 a_n1996_n452.t58 gnd 0.710766f
C712 a_n1996_n452.n83 gnd 0.303445f
C713 a_n1996_n452.n84 gnd 0.297934f
C714 a_n1996_n452.t54 gnd 0.710766f
C715 a_n1996_n452.n85 gnd 0.303445f
C716 a_n1996_n452.n86 gnd 0.297934f
C717 a_n1996_n452.n87 gnd 1.00969f
C718 a_n1996_n452.t65 gnd 0.713776f
C719 a_n1996_n452.n88 gnd 0.309973f
C720 a_n1996_n452.t45 gnd 0.699053f
C721 a_n1996_n452.n89 gnd 0.303445f
C722 a_n1996_n452.n90 gnd 0.309974f
C723 a_n1996_n452.t46 gnd 0.710611f
C724 a_n1996_n452.t26 gnd 0.713776f
C725 a_n1996_n452.n91 gnd 0.309973f
C726 a_n1996_n452.t14 gnd 0.699053f
C727 a_n1996_n452.n92 gnd 0.303445f
C728 a_n1996_n452.n93 gnd 0.309974f
C729 a_n1996_n452.t16 gnd 0.710611f
C730 a_n1996_n452.n94 gnd 1.13585f
C731 a_n1996_n452.t17 gnd 1.40439f
C732 a_n1996_n452.t33 gnd 0.150285f
C733 a_n1996_n452.t35 gnd 0.150285f
C734 a_n1996_n452.n95 gnd 1.05861f
C735 a_n1996_n452.n96 gnd 1.18283f
C736 a_n1996_n452.n97 gnd 1.05861f
C737 a_n1996_n452.t15 gnd 0.150285f
C738 a_n3827_n3924.t11 gnd 0.091917f
C739 a_n3827_n3924.t17 gnd 0.091917f
C740 a_n3827_n3924.n0 gnd 0.750696f
C741 a_n3827_n3924.n1 gnd 0.341384f
C742 a_n3827_n3924.t2 gnd 0.955301f
C743 a_n3827_n3924.n2 gnd 0.859345f
C744 a_n3827_n3924.t14 gnd 0.091917f
C745 a_n3827_n3924.t16 gnd 0.091917f
C746 a_n3827_n3924.n3 gnd 0.750697f
C747 a_n3827_n3924.n4 gnd 0.341383f
C748 a_n3827_n3924.t18 gnd 0.091917f
C749 a_n3827_n3924.t19 gnd 0.091917f
C750 a_n3827_n3924.n5 gnd 0.750697f
C751 a_n3827_n3924.n6 gnd 0.341383f
C752 a_n3827_n3924.t5 gnd 0.091917f
C753 a_n3827_n3924.t3 gnd 0.091917f
C754 a_n3827_n3924.n7 gnd 0.750697f
C755 a_n3827_n3924.n8 gnd 0.341383f
C756 a_n3827_n3924.t9 gnd 0.091917f
C757 a_n3827_n3924.t4 gnd 0.091917f
C758 a_n3827_n3924.n9 gnd 0.750697f
C759 a_n3827_n3924.n10 gnd 0.341383f
C760 a_n3827_n3924.t8 gnd 0.955305f
C761 a_n3827_n3924.n11 gnd 0.342685f
C762 a_n3827_n3924.t29 gnd 0.955305f
C763 a_n3827_n3924.n12 gnd 0.342685f
C764 a_n3827_n3924.t46 gnd 0.091917f
C765 a_n3827_n3924.t23 gnd 0.091917f
C766 a_n3827_n3924.n13 gnd 0.750697f
C767 a_n3827_n3924.n14 gnd 0.341383f
C768 a_n3827_n3924.t41 gnd 0.091917f
C769 a_n3827_n3924.t1 gnd 0.091917f
C770 a_n3827_n3924.n15 gnd 0.750697f
C771 a_n3827_n3924.n16 gnd 0.341383f
C772 a_n3827_n3924.t45 gnd 0.091917f
C773 a_n3827_n3924.t34 gnd 0.091917f
C774 a_n3827_n3924.n17 gnd 0.750697f
C775 a_n3827_n3924.n18 gnd 0.341383f
C776 a_n3827_n3924.t30 gnd 0.091917f
C777 a_n3827_n3924.t35 gnd 0.091917f
C778 a_n3827_n3924.n19 gnd 0.750697f
C779 a_n3827_n3924.n20 gnd 0.341383f
C780 a_n3827_n3924.t32 gnd 0.955305f
C781 a_n3827_n3924.n21 gnd 0.859341f
C782 a_n3827_n3924.t12 gnd 0.955301f
C783 a_n3827_n3924.n22 gnd 0.558761f
C784 a_n3827_n3924.n23 gnd 0.862207f
C785 a_n3827_n3924.t0 gnd 1.18864f
C786 a_n3827_n3924.t36 gnd 1.18694f
C787 a_n3827_n3924.n24 gnd 1.35306f
C788 a_n3827_n3924.n25 gnd 0.451836f
C789 a_n3827_n3924.t25 gnd 1.18694f
C790 a_n3827_n3924.n26 gnd 0.543403f
C791 a_n3827_n3924.t24 gnd 1.18694f
C792 a_n3827_n3924.n27 gnd 0.835985f
C793 a_n3827_n3924.t40 gnd 1.18694f
C794 a_n3827_n3924.n28 gnd 0.835985f
C795 a_n3827_n3924.t27 gnd 1.18694f
C796 a_n3827_n3924.n29 gnd 0.835985f
C797 a_n3827_n3924.t39 gnd 1.18694f
C798 a_n3827_n3924.n30 gnd 0.835985f
C799 a_n3827_n3924.t49 gnd 1.18694f
C800 a_n3827_n3924.n31 gnd 0.792525f
C801 a_n3827_n3924.t48 gnd 1.19019f
C802 a_n3827_n3924.t44 gnd 1.18694f
C803 a_n3827_n3924.n32 gnd 1.60062f
C804 a_n3827_n3924.n33 gnd 0.451836f
C805 a_n3827_n3924.n34 gnd 0.862207f
C806 a_n3827_n3924.t37 gnd 0.955301f
C807 a_n3827_n3924.n35 gnd 0.558761f
C808 a_n3827_n3924.t28 gnd 0.091917f
C809 a_n3827_n3924.t31 gnd 0.091917f
C810 a_n3827_n3924.n36 gnd 0.750696f
C811 a_n3827_n3924.n37 gnd 0.341384f
C812 a_n3827_n3924.t22 gnd 0.091917f
C813 a_n3827_n3924.t26 gnd 0.091917f
C814 a_n3827_n3924.n38 gnd 0.750696f
C815 a_n3827_n3924.n39 gnd 0.341384f
C816 a_n3827_n3924.t43 gnd 0.091917f
C817 a_n3827_n3924.t33 gnd 0.091917f
C818 a_n3827_n3924.n40 gnd 0.750696f
C819 a_n3827_n3924.n41 gnd 0.341384f
C820 a_n3827_n3924.t38 gnd 0.091917f
C821 a_n3827_n3924.t47 gnd 0.091917f
C822 a_n3827_n3924.n42 gnd 0.750696f
C823 a_n3827_n3924.n43 gnd 0.341384f
C824 a_n3827_n3924.t42 gnd 0.955301f
C825 a_n3827_n3924.n44 gnd 0.342688f
C826 a_n3827_n3924.t13 gnd 0.955301f
C827 a_n3827_n3924.n45 gnd 0.342688f
C828 a_n3827_n3924.t10 gnd 0.091917f
C829 a_n3827_n3924.t15 gnd 0.091917f
C830 a_n3827_n3924.n46 gnd 0.750696f
C831 a_n3827_n3924.n47 gnd 0.341384f
C832 a_n3827_n3924.t7 gnd 0.091917f
C833 a_n3827_n3924.t6 gnd 0.091917f
C834 a_n3827_n3924.n48 gnd 0.750696f
C835 a_n3827_n3924.n49 gnd 0.341384f
C836 a_n3827_n3924.n50 gnd 0.341387f
C837 a_n3827_n3924.t20 gnd 0.091917f
C838 a_n3827_n3924.n51 gnd 0.750693f
C839 a_n3827_n3924.t21 gnd 0.091917f
C840 plus.n0 gnd 0.0228f
C841 plus.t14 gnd 0.32248f
C842 plus.n1 gnd 0.0228f
C843 plus.t15 gnd 0.32248f
C844 plus.t9 gnd 0.32248f
C845 plus.n2 gnd 0.143256f
C846 plus.n3 gnd 0.0228f
C847 plus.t5 gnd 0.32248f
C848 plus.t6 gnd 0.32248f
C849 plus.n4 gnd 0.143256f
C850 plus.n5 gnd 0.0228f
C851 plus.t19 gnd 0.32248f
C852 plus.t20 gnd 0.32248f
C853 plus.n6 gnd 0.143256f
C854 plus.n7 gnd 0.0228f
C855 plus.t16 gnd 0.32248f
C856 plus.t11 gnd 0.32248f
C857 plus.n8 gnd 0.147069f
C858 plus.t13 gnd 0.333778f
C859 plus.n9 gnd 0.133595f
C860 plus.n10 gnd 0.097318f
C861 plus.n11 gnd 0.005174f
C862 plus.n12 gnd 0.143256f
C863 plus.n13 gnd 0.005174f
C864 plus.n14 gnd 0.0228f
C865 plus.n15 gnd 0.0228f
C866 plus.n16 gnd 0.0228f
C867 plus.n17 gnd 0.005174f
C868 plus.n18 gnd 0.143256f
C869 plus.n19 gnd 0.005174f
C870 plus.n20 gnd 0.0228f
C871 plus.n21 gnd 0.0228f
C872 plus.n22 gnd 0.0228f
C873 plus.n23 gnd 0.005174f
C874 plus.n24 gnd 0.143256f
C875 plus.n25 gnd 0.005174f
C876 plus.n26 gnd 0.0228f
C877 plus.n27 gnd 0.0228f
C878 plus.n28 gnd 0.0228f
C879 plus.n29 gnd 0.005174f
C880 plus.n30 gnd 0.143256f
C881 plus.n31 gnd 0.005174f
C882 plus.n32 gnd 0.143045f
C883 plus.n33 gnd 0.257559f
C884 plus.n34 gnd 0.0228f
C885 plus.n35 gnd 0.005174f
C886 plus.t10 gnd 0.32248f
C887 plus.n36 gnd 0.0228f
C888 plus.n37 gnd 0.005174f
C889 plus.t7 gnd 0.32248f
C890 plus.n38 gnd 0.0228f
C891 plus.n39 gnd 0.005174f
C892 plus.t23 gnd 0.32248f
C893 plus.n40 gnd 0.0228f
C894 plus.n41 gnd 0.005174f
C895 plus.t22 gnd 0.32248f
C896 plus.t18 gnd 0.333778f
C897 plus.t17 gnd 0.32248f
C898 plus.n42 gnd 0.147069f
C899 plus.n43 gnd 0.133595f
C900 plus.n44 gnd 0.097318f
C901 plus.n45 gnd 0.0228f
C902 plus.n46 gnd 0.143256f
C903 plus.n47 gnd 0.005174f
C904 plus.t21 gnd 0.32248f
C905 plus.n48 gnd 0.143256f
C906 plus.n49 gnd 0.0228f
C907 plus.n50 gnd 0.0228f
C908 plus.n51 gnd 0.0228f
C909 plus.n52 gnd 0.143256f
C910 plus.n53 gnd 0.005174f
C911 plus.t8 gnd 0.32248f
C912 plus.n54 gnd 0.143256f
C913 plus.n55 gnd 0.0228f
C914 plus.n56 gnd 0.0228f
C915 plus.n57 gnd 0.0228f
C916 plus.n58 gnd 0.143256f
C917 plus.n59 gnd 0.005174f
C918 plus.t12 gnd 0.32248f
C919 plus.n60 gnd 0.143256f
C920 plus.n61 gnd 0.0228f
C921 plus.n62 gnd 0.0228f
C922 plus.n63 gnd 0.0228f
C923 plus.n64 gnd 0.143256f
C924 plus.n65 gnd 0.005174f
C925 plus.t24 gnd 0.32248f
C926 plus.n66 gnd 0.143045f
C927 plus.n67 gnd 0.703278f
C928 plus.n68 gnd 1.06353f
C929 plus.t0 gnd 0.039359f
C930 plus.t4 gnd 0.007028f
C931 plus.t2 gnd 0.007028f
C932 plus.n69 gnd 0.022794f
C933 plus.n70 gnd 0.176956f
C934 plus.t1 gnd 0.007028f
C935 plus.t3 gnd 0.007028f
C936 plus.n71 gnd 0.022794f
C937 plus.n72 gnd 0.132827f
C938 plus.n73 gnd 2.78062f
C939 commonsourceibias.n0 gnd 0.012626f
C940 commonsourceibias.t78 gnd 0.191194f
C941 commonsourceibias.t146 gnd 0.176786f
C942 commonsourceibias.n1 gnd 0.007691f
C943 commonsourceibias.n2 gnd 0.009462f
C944 commonsourceibias.t96 gnd 0.176786f
C945 commonsourceibias.n3 gnd 0.009599f
C946 commonsourceibias.n4 gnd 0.009462f
C947 commonsourceibias.t157 gnd 0.176786f
C948 commonsourceibias.n5 gnd 0.070538f
C949 commonsourceibias.t112 gnd 0.176786f
C950 commonsourceibias.n6 gnd 0.007654f
C951 commonsourceibias.n7 gnd 0.009462f
C952 commonsourceibias.t75 gnd 0.176786f
C953 commonsourceibias.n8 gnd 0.009135f
C954 commonsourceibias.n9 gnd 0.009462f
C955 commonsourceibias.t124 gnd 0.176786f
C956 commonsourceibias.n10 gnd 0.070538f
C957 commonsourceibias.t113 gnd 0.176786f
C958 commonsourceibias.n11 gnd 0.007642f
C959 commonsourceibias.n12 gnd 0.012626f
C960 commonsourceibias.t58 gnd 0.191194f
C961 commonsourceibias.t52 gnd 0.176786f
C962 commonsourceibias.n13 gnd 0.007691f
C963 commonsourceibias.n14 gnd 0.009462f
C964 commonsourceibias.t4 gnd 0.176786f
C965 commonsourceibias.n15 gnd 0.009599f
C966 commonsourceibias.n16 gnd 0.009462f
C967 commonsourceibias.t44 gnd 0.176786f
C968 commonsourceibias.n17 gnd 0.070538f
C969 commonsourceibias.t18 gnd 0.176786f
C970 commonsourceibias.n18 gnd 0.007654f
C971 commonsourceibias.n19 gnd 0.009462f
C972 commonsourceibias.t16 gnd 0.176786f
C973 commonsourceibias.n20 gnd 0.009135f
C974 commonsourceibias.n21 gnd 0.009462f
C975 commonsourceibias.t8 gnd 0.176786f
C976 commonsourceibias.n22 gnd 0.070538f
C977 commonsourceibias.t14 gnd 0.176786f
C978 commonsourceibias.n23 gnd 0.007642f
C979 commonsourceibias.n24 gnd 0.009462f
C980 commonsourceibias.t46 gnd 0.176786f
C981 commonsourceibias.t22 gnd 0.176786f
C982 commonsourceibias.n25 gnd 0.070538f
C983 commonsourceibias.n26 gnd 0.009462f
C984 commonsourceibias.t2 gnd 0.176786f
C985 commonsourceibias.n27 gnd 0.070538f
C986 commonsourceibias.n28 gnd 0.009462f
C987 commonsourceibias.t28 gnd 0.176786f
C988 commonsourceibias.n29 gnd 0.070538f
C989 commonsourceibias.n30 gnd 0.009462f
C990 commonsourceibias.t20 gnd 0.176786f
C991 commonsourceibias.n31 gnd 0.010756f
C992 commonsourceibias.n32 gnd 0.009462f
C993 commonsourceibias.t56 gnd 0.176786f
C994 commonsourceibias.n33 gnd 0.012719f
C995 commonsourceibias.t54 gnd 0.196936f
C996 commonsourceibias.t30 gnd 0.176786f
C997 commonsourceibias.n34 gnd 0.078597f
C998 commonsourceibias.n35 gnd 0.084205f
C999 commonsourceibias.n36 gnd 0.040277f
C1000 commonsourceibias.n37 gnd 0.009462f
C1001 commonsourceibias.n38 gnd 0.007691f
C1002 commonsourceibias.n39 gnd 0.013039f
C1003 commonsourceibias.n40 gnd 0.070538f
C1004 commonsourceibias.n41 gnd 0.013095f
C1005 commonsourceibias.n42 gnd 0.009462f
C1006 commonsourceibias.n43 gnd 0.009462f
C1007 commonsourceibias.n44 gnd 0.009462f
C1008 commonsourceibias.n45 gnd 0.009599f
C1009 commonsourceibias.n46 gnd 0.070538f
C1010 commonsourceibias.n47 gnd 0.011663f
C1011 commonsourceibias.n48 gnd 0.012902f
C1012 commonsourceibias.n49 gnd 0.009462f
C1013 commonsourceibias.n50 gnd 0.009462f
C1014 commonsourceibias.n51 gnd 0.012818f
C1015 commonsourceibias.n52 gnd 0.007654f
C1016 commonsourceibias.n53 gnd 0.012977f
C1017 commonsourceibias.n54 gnd 0.009462f
C1018 commonsourceibias.n55 gnd 0.009462f
C1019 commonsourceibias.n56 gnd 0.013056f
C1020 commonsourceibias.n57 gnd 0.011258f
C1021 commonsourceibias.n58 gnd 0.009135f
C1022 commonsourceibias.n59 gnd 0.009462f
C1023 commonsourceibias.n60 gnd 0.009462f
C1024 commonsourceibias.n61 gnd 0.011574f
C1025 commonsourceibias.n62 gnd 0.012991f
C1026 commonsourceibias.n63 gnd 0.070538f
C1027 commonsourceibias.n64 gnd 0.012903f
C1028 commonsourceibias.n65 gnd 0.009462f
C1029 commonsourceibias.n66 gnd 0.009462f
C1030 commonsourceibias.n67 gnd 0.009462f
C1031 commonsourceibias.n68 gnd 0.012903f
C1032 commonsourceibias.n69 gnd 0.070538f
C1033 commonsourceibias.n70 gnd 0.012991f
C1034 commonsourceibias.n71 gnd 0.011574f
C1035 commonsourceibias.n72 gnd 0.009462f
C1036 commonsourceibias.n73 gnd 0.009462f
C1037 commonsourceibias.n74 gnd 0.009462f
C1038 commonsourceibias.n75 gnd 0.011258f
C1039 commonsourceibias.n76 gnd 0.013056f
C1040 commonsourceibias.n77 gnd 0.070538f
C1041 commonsourceibias.n78 gnd 0.012977f
C1042 commonsourceibias.n79 gnd 0.009462f
C1043 commonsourceibias.n80 gnd 0.009462f
C1044 commonsourceibias.n81 gnd 0.009462f
C1045 commonsourceibias.n82 gnd 0.012818f
C1046 commonsourceibias.n83 gnd 0.070538f
C1047 commonsourceibias.n84 gnd 0.012902f
C1048 commonsourceibias.n85 gnd 0.011663f
C1049 commonsourceibias.n86 gnd 0.009462f
C1050 commonsourceibias.n87 gnd 0.009462f
C1051 commonsourceibias.n88 gnd 0.009462f
C1052 commonsourceibias.n89 gnd 0.010756f
C1053 commonsourceibias.n90 gnd 0.013095f
C1054 commonsourceibias.n91 gnd 0.070538f
C1055 commonsourceibias.n92 gnd 0.013039f
C1056 commonsourceibias.n93 gnd 0.009462f
C1057 commonsourceibias.n94 gnd 0.009462f
C1058 commonsourceibias.n95 gnd 0.009462f
C1059 commonsourceibias.n96 gnd 0.012719f
C1060 commonsourceibias.n97 gnd 0.070538f
C1061 commonsourceibias.n98 gnd 0.01275f
C1062 commonsourceibias.n99 gnd 0.085058f
C1063 commonsourceibias.n100 gnd 0.095108f
C1064 commonsourceibias.t59 gnd 0.020419f
C1065 commonsourceibias.t53 gnd 0.020419f
C1066 commonsourceibias.n101 gnd 0.180428f
C1067 commonsourceibias.n102 gnd 0.15629f
C1068 commonsourceibias.t5 gnd 0.020419f
C1069 commonsourceibias.t45 gnd 0.020419f
C1070 commonsourceibias.n103 gnd 0.180428f
C1071 commonsourceibias.n104 gnd 0.082878f
C1072 commonsourceibias.t19 gnd 0.020419f
C1073 commonsourceibias.t17 gnd 0.020419f
C1074 commonsourceibias.n105 gnd 0.180428f
C1075 commonsourceibias.n106 gnd 0.082878f
C1076 commonsourceibias.t9 gnd 0.020419f
C1077 commonsourceibias.t15 gnd 0.020419f
C1078 commonsourceibias.n107 gnd 0.180428f
C1079 commonsourceibias.n108 gnd 0.06924f
C1080 commonsourceibias.t31 gnd 0.020419f
C1081 commonsourceibias.t55 gnd 0.020419f
C1082 commonsourceibias.n109 gnd 0.181032f
C1083 commonsourceibias.t21 gnd 0.020419f
C1084 commonsourceibias.t57 gnd 0.020419f
C1085 commonsourceibias.n110 gnd 0.180428f
C1086 commonsourceibias.n111 gnd 0.168125f
C1087 commonsourceibias.t3 gnd 0.020419f
C1088 commonsourceibias.t29 gnd 0.020419f
C1089 commonsourceibias.n112 gnd 0.180428f
C1090 commonsourceibias.n113 gnd 0.082878f
C1091 commonsourceibias.t47 gnd 0.020419f
C1092 commonsourceibias.t23 gnd 0.020419f
C1093 commonsourceibias.n114 gnd 0.180428f
C1094 commonsourceibias.n115 gnd 0.06924f
C1095 commonsourceibias.n116 gnd 0.083843f
C1096 commonsourceibias.n117 gnd 0.009462f
C1097 commonsourceibias.t154 gnd 0.176786f
C1098 commonsourceibias.t106 gnd 0.176786f
C1099 commonsourceibias.n118 gnd 0.070538f
C1100 commonsourceibias.n119 gnd 0.009462f
C1101 commonsourceibias.t92 gnd 0.176786f
C1102 commonsourceibias.n120 gnd 0.070538f
C1103 commonsourceibias.n121 gnd 0.009462f
C1104 commonsourceibias.t123 gnd 0.176786f
C1105 commonsourceibias.n122 gnd 0.070538f
C1106 commonsourceibias.n123 gnd 0.009462f
C1107 commonsourceibias.t110 gnd 0.176786f
C1108 commonsourceibias.n124 gnd 0.010756f
C1109 commonsourceibias.n125 gnd 0.009462f
C1110 commonsourceibias.t82 gnd 0.176786f
C1111 commonsourceibias.n126 gnd 0.012719f
C1112 commonsourceibias.t132 gnd 0.196936f
C1113 commonsourceibias.t147 gnd 0.176786f
C1114 commonsourceibias.n127 gnd 0.078597f
C1115 commonsourceibias.n128 gnd 0.084205f
C1116 commonsourceibias.n129 gnd 0.040277f
C1117 commonsourceibias.n130 gnd 0.009462f
C1118 commonsourceibias.n131 gnd 0.007691f
C1119 commonsourceibias.n132 gnd 0.013039f
C1120 commonsourceibias.n133 gnd 0.070538f
C1121 commonsourceibias.n134 gnd 0.013095f
C1122 commonsourceibias.n135 gnd 0.009462f
C1123 commonsourceibias.n136 gnd 0.009462f
C1124 commonsourceibias.n137 gnd 0.009462f
C1125 commonsourceibias.n138 gnd 0.009599f
C1126 commonsourceibias.n139 gnd 0.070538f
C1127 commonsourceibias.n140 gnd 0.011663f
C1128 commonsourceibias.n141 gnd 0.012902f
C1129 commonsourceibias.n142 gnd 0.009462f
C1130 commonsourceibias.n143 gnd 0.009462f
C1131 commonsourceibias.n144 gnd 0.012818f
C1132 commonsourceibias.n145 gnd 0.007654f
C1133 commonsourceibias.n146 gnd 0.012977f
C1134 commonsourceibias.n147 gnd 0.009462f
C1135 commonsourceibias.n148 gnd 0.009462f
C1136 commonsourceibias.n149 gnd 0.013056f
C1137 commonsourceibias.n150 gnd 0.011258f
C1138 commonsourceibias.n151 gnd 0.009135f
C1139 commonsourceibias.n152 gnd 0.009462f
C1140 commonsourceibias.n153 gnd 0.009462f
C1141 commonsourceibias.n154 gnd 0.011574f
C1142 commonsourceibias.n155 gnd 0.012991f
C1143 commonsourceibias.n156 gnd 0.070538f
C1144 commonsourceibias.n157 gnd 0.012903f
C1145 commonsourceibias.n158 gnd 0.009417f
C1146 commonsourceibias.n159 gnd 0.068402f
C1147 commonsourceibias.n160 gnd 0.009417f
C1148 commonsourceibias.n161 gnd 0.012903f
C1149 commonsourceibias.n162 gnd 0.070538f
C1150 commonsourceibias.n163 gnd 0.012991f
C1151 commonsourceibias.n164 gnd 0.011574f
C1152 commonsourceibias.n165 gnd 0.009462f
C1153 commonsourceibias.n166 gnd 0.009462f
C1154 commonsourceibias.n167 gnd 0.009462f
C1155 commonsourceibias.n168 gnd 0.011258f
C1156 commonsourceibias.n169 gnd 0.013056f
C1157 commonsourceibias.n170 gnd 0.070538f
C1158 commonsourceibias.n171 gnd 0.012977f
C1159 commonsourceibias.n172 gnd 0.009462f
C1160 commonsourceibias.n173 gnd 0.009462f
C1161 commonsourceibias.n174 gnd 0.009462f
C1162 commonsourceibias.n175 gnd 0.012818f
C1163 commonsourceibias.n176 gnd 0.070538f
C1164 commonsourceibias.n177 gnd 0.012902f
C1165 commonsourceibias.n178 gnd 0.011663f
C1166 commonsourceibias.n179 gnd 0.009462f
C1167 commonsourceibias.n180 gnd 0.009462f
C1168 commonsourceibias.n181 gnd 0.009462f
C1169 commonsourceibias.n182 gnd 0.010756f
C1170 commonsourceibias.n183 gnd 0.013095f
C1171 commonsourceibias.n184 gnd 0.070538f
C1172 commonsourceibias.n185 gnd 0.013039f
C1173 commonsourceibias.n186 gnd 0.009462f
C1174 commonsourceibias.n187 gnd 0.009462f
C1175 commonsourceibias.n188 gnd 0.009462f
C1176 commonsourceibias.n189 gnd 0.012719f
C1177 commonsourceibias.n190 gnd 0.070538f
C1178 commonsourceibias.n191 gnd 0.01275f
C1179 commonsourceibias.n192 gnd 0.085058f
C1180 commonsourceibias.n193 gnd 0.056191f
C1181 commonsourceibias.n194 gnd 0.012626f
C1182 commonsourceibias.t115 gnd 0.191194f
C1183 commonsourceibias.t138 gnd 0.176786f
C1184 commonsourceibias.n195 gnd 0.007691f
C1185 commonsourceibias.n196 gnd 0.009462f
C1186 commonsourceibias.t128 gnd 0.176786f
C1187 commonsourceibias.n197 gnd 0.009599f
C1188 commonsourceibias.n198 gnd 0.009462f
C1189 commonsourceibias.t116 gnd 0.176786f
C1190 commonsourceibias.n199 gnd 0.070538f
C1191 commonsourceibias.t139 gnd 0.176786f
C1192 commonsourceibias.n200 gnd 0.007654f
C1193 commonsourceibias.n201 gnd 0.009462f
C1194 commonsourceibias.t126 gnd 0.176786f
C1195 commonsourceibias.n202 gnd 0.009135f
C1196 commonsourceibias.n203 gnd 0.009462f
C1197 commonsourceibias.t114 gnd 0.176786f
C1198 commonsourceibias.n204 gnd 0.070538f
C1199 commonsourceibias.t140 gnd 0.176786f
C1200 commonsourceibias.n205 gnd 0.007642f
C1201 commonsourceibias.n206 gnd 0.009462f
C1202 commonsourceibias.t127 gnd 0.176786f
C1203 commonsourceibias.t149 gnd 0.176786f
C1204 commonsourceibias.n207 gnd 0.070538f
C1205 commonsourceibias.n208 gnd 0.009462f
C1206 commonsourceibias.t141 gnd 0.176786f
C1207 commonsourceibias.n209 gnd 0.070538f
C1208 commonsourceibias.n210 gnd 0.009462f
C1209 commonsourceibias.t125 gnd 0.176786f
C1210 commonsourceibias.n211 gnd 0.070538f
C1211 commonsourceibias.n212 gnd 0.009462f
C1212 commonsourceibias.t152 gnd 0.176786f
C1213 commonsourceibias.n213 gnd 0.010756f
C1214 commonsourceibias.n214 gnd 0.009462f
C1215 commonsourceibias.t69 gnd 0.176786f
C1216 commonsourceibias.n215 gnd 0.012719f
C1217 commonsourceibias.t64 gnd 0.196936f
C1218 commonsourceibias.t135 gnd 0.176786f
C1219 commonsourceibias.n216 gnd 0.078597f
C1220 commonsourceibias.n217 gnd 0.084205f
C1221 commonsourceibias.n218 gnd 0.040277f
C1222 commonsourceibias.n219 gnd 0.009462f
C1223 commonsourceibias.n220 gnd 0.007691f
C1224 commonsourceibias.n221 gnd 0.013039f
C1225 commonsourceibias.n222 gnd 0.070538f
C1226 commonsourceibias.n223 gnd 0.013095f
C1227 commonsourceibias.n224 gnd 0.009462f
C1228 commonsourceibias.n225 gnd 0.009462f
C1229 commonsourceibias.n226 gnd 0.009462f
C1230 commonsourceibias.n227 gnd 0.009599f
C1231 commonsourceibias.n228 gnd 0.070538f
C1232 commonsourceibias.n229 gnd 0.011663f
C1233 commonsourceibias.n230 gnd 0.012902f
C1234 commonsourceibias.n231 gnd 0.009462f
C1235 commonsourceibias.n232 gnd 0.009462f
C1236 commonsourceibias.n233 gnd 0.012818f
C1237 commonsourceibias.n234 gnd 0.007654f
C1238 commonsourceibias.n235 gnd 0.012977f
C1239 commonsourceibias.n236 gnd 0.009462f
C1240 commonsourceibias.n237 gnd 0.009462f
C1241 commonsourceibias.n238 gnd 0.013056f
C1242 commonsourceibias.n239 gnd 0.011258f
C1243 commonsourceibias.n240 gnd 0.009135f
C1244 commonsourceibias.n241 gnd 0.009462f
C1245 commonsourceibias.n242 gnd 0.009462f
C1246 commonsourceibias.n243 gnd 0.011574f
C1247 commonsourceibias.n244 gnd 0.012991f
C1248 commonsourceibias.n245 gnd 0.070538f
C1249 commonsourceibias.n246 gnd 0.012903f
C1250 commonsourceibias.n247 gnd 0.009462f
C1251 commonsourceibias.n248 gnd 0.009462f
C1252 commonsourceibias.n249 gnd 0.009462f
C1253 commonsourceibias.n250 gnd 0.012903f
C1254 commonsourceibias.n251 gnd 0.070538f
C1255 commonsourceibias.n252 gnd 0.012991f
C1256 commonsourceibias.n253 gnd 0.011574f
C1257 commonsourceibias.n254 gnd 0.009462f
C1258 commonsourceibias.n255 gnd 0.009462f
C1259 commonsourceibias.n256 gnd 0.009462f
C1260 commonsourceibias.n257 gnd 0.011258f
C1261 commonsourceibias.n258 gnd 0.013056f
C1262 commonsourceibias.n259 gnd 0.070538f
C1263 commonsourceibias.n260 gnd 0.012977f
C1264 commonsourceibias.n261 gnd 0.009462f
C1265 commonsourceibias.n262 gnd 0.009462f
C1266 commonsourceibias.n263 gnd 0.009462f
C1267 commonsourceibias.n264 gnd 0.012818f
C1268 commonsourceibias.n265 gnd 0.070538f
C1269 commonsourceibias.n266 gnd 0.012902f
C1270 commonsourceibias.n267 gnd 0.011663f
C1271 commonsourceibias.n268 gnd 0.009462f
C1272 commonsourceibias.n269 gnd 0.009462f
C1273 commonsourceibias.n270 gnd 0.009462f
C1274 commonsourceibias.n271 gnd 0.010756f
C1275 commonsourceibias.n272 gnd 0.013095f
C1276 commonsourceibias.n273 gnd 0.070538f
C1277 commonsourceibias.n274 gnd 0.013039f
C1278 commonsourceibias.n275 gnd 0.009462f
C1279 commonsourceibias.n276 gnd 0.009462f
C1280 commonsourceibias.n277 gnd 0.009462f
C1281 commonsourceibias.n278 gnd 0.012719f
C1282 commonsourceibias.n279 gnd 0.070538f
C1283 commonsourceibias.n280 gnd 0.01275f
C1284 commonsourceibias.n281 gnd 0.085058f
C1285 commonsourceibias.n282 gnd 0.030353f
C1286 commonsourceibias.n283 gnd 0.151535f
C1287 commonsourceibias.n284 gnd 0.012626f
C1288 commonsourceibias.t68 gnd 0.176786f
C1289 commonsourceibias.n285 gnd 0.007691f
C1290 commonsourceibias.n286 gnd 0.009462f
C1291 commonsourceibias.t80 gnd 0.176786f
C1292 commonsourceibias.n287 gnd 0.009599f
C1293 commonsourceibias.n288 gnd 0.009462f
C1294 commonsourceibias.t134 gnd 0.176786f
C1295 commonsourceibias.n289 gnd 0.070538f
C1296 commonsourceibias.t159 gnd 0.176786f
C1297 commonsourceibias.n290 gnd 0.007654f
C1298 commonsourceibias.n291 gnd 0.009462f
C1299 commonsourceibias.t74 gnd 0.176786f
C1300 commonsourceibias.n292 gnd 0.009135f
C1301 commonsourceibias.n293 gnd 0.009462f
C1302 commonsourceibias.t120 gnd 0.176786f
C1303 commonsourceibias.n294 gnd 0.070538f
C1304 commonsourceibias.t111 gnd 0.176786f
C1305 commonsourceibias.n295 gnd 0.007642f
C1306 commonsourceibias.n296 gnd 0.009462f
C1307 commonsourceibias.t67 gnd 0.176786f
C1308 commonsourceibias.t81 gnd 0.176786f
C1309 commonsourceibias.n297 gnd 0.070538f
C1310 commonsourceibias.n298 gnd 0.009462f
C1311 commonsourceibias.t101 gnd 0.176786f
C1312 commonsourceibias.n299 gnd 0.070538f
C1313 commonsourceibias.n300 gnd 0.009462f
C1314 commonsourceibias.t158 gnd 0.176786f
C1315 commonsourceibias.n301 gnd 0.070538f
C1316 commonsourceibias.n302 gnd 0.009462f
C1317 commonsourceibias.t150 gnd 0.176786f
C1318 commonsourceibias.n303 gnd 0.010756f
C1319 commonsourceibias.n304 gnd 0.009462f
C1320 commonsourceibias.t70 gnd 0.176786f
C1321 commonsourceibias.n305 gnd 0.012719f
C1322 commonsourceibias.t136 gnd 0.196936f
C1323 commonsourceibias.t143 gnd 0.176786f
C1324 commonsourceibias.n306 gnd 0.078597f
C1325 commonsourceibias.n307 gnd 0.084205f
C1326 commonsourceibias.n308 gnd 0.040277f
C1327 commonsourceibias.n309 gnd 0.009462f
C1328 commonsourceibias.n310 gnd 0.007691f
C1329 commonsourceibias.n311 gnd 0.013039f
C1330 commonsourceibias.n312 gnd 0.070538f
C1331 commonsourceibias.n313 gnd 0.013095f
C1332 commonsourceibias.n314 gnd 0.009462f
C1333 commonsourceibias.n315 gnd 0.009462f
C1334 commonsourceibias.n316 gnd 0.009462f
C1335 commonsourceibias.n317 gnd 0.009599f
C1336 commonsourceibias.n318 gnd 0.070538f
C1337 commonsourceibias.n319 gnd 0.011663f
C1338 commonsourceibias.n320 gnd 0.012902f
C1339 commonsourceibias.n321 gnd 0.009462f
C1340 commonsourceibias.n322 gnd 0.009462f
C1341 commonsourceibias.n323 gnd 0.012818f
C1342 commonsourceibias.n324 gnd 0.007654f
C1343 commonsourceibias.n325 gnd 0.012977f
C1344 commonsourceibias.n326 gnd 0.009462f
C1345 commonsourceibias.n327 gnd 0.009462f
C1346 commonsourceibias.n328 gnd 0.013056f
C1347 commonsourceibias.n329 gnd 0.011258f
C1348 commonsourceibias.n330 gnd 0.009135f
C1349 commonsourceibias.n331 gnd 0.009462f
C1350 commonsourceibias.n332 gnd 0.009462f
C1351 commonsourceibias.n333 gnd 0.011574f
C1352 commonsourceibias.n334 gnd 0.012991f
C1353 commonsourceibias.n335 gnd 0.070538f
C1354 commonsourceibias.n336 gnd 0.012903f
C1355 commonsourceibias.n337 gnd 0.009462f
C1356 commonsourceibias.n338 gnd 0.009462f
C1357 commonsourceibias.n339 gnd 0.009462f
C1358 commonsourceibias.n340 gnd 0.012903f
C1359 commonsourceibias.n341 gnd 0.070538f
C1360 commonsourceibias.n342 gnd 0.012991f
C1361 commonsourceibias.n343 gnd 0.011574f
C1362 commonsourceibias.n344 gnd 0.009462f
C1363 commonsourceibias.n345 gnd 0.009462f
C1364 commonsourceibias.n346 gnd 0.009462f
C1365 commonsourceibias.n347 gnd 0.011258f
C1366 commonsourceibias.n348 gnd 0.013056f
C1367 commonsourceibias.n349 gnd 0.070538f
C1368 commonsourceibias.n350 gnd 0.012977f
C1369 commonsourceibias.n351 gnd 0.009462f
C1370 commonsourceibias.n352 gnd 0.009462f
C1371 commonsourceibias.n353 gnd 0.009462f
C1372 commonsourceibias.n354 gnd 0.012818f
C1373 commonsourceibias.n355 gnd 0.070538f
C1374 commonsourceibias.n356 gnd 0.012902f
C1375 commonsourceibias.n357 gnd 0.011663f
C1376 commonsourceibias.n358 gnd 0.009462f
C1377 commonsourceibias.n359 gnd 0.009462f
C1378 commonsourceibias.n360 gnd 0.009462f
C1379 commonsourceibias.n361 gnd 0.010756f
C1380 commonsourceibias.n362 gnd 0.013095f
C1381 commonsourceibias.n363 gnd 0.070538f
C1382 commonsourceibias.n364 gnd 0.013039f
C1383 commonsourceibias.n365 gnd 0.009462f
C1384 commonsourceibias.n366 gnd 0.009462f
C1385 commonsourceibias.n367 gnd 0.009462f
C1386 commonsourceibias.n368 gnd 0.012719f
C1387 commonsourceibias.n369 gnd 0.070538f
C1388 commonsourceibias.n370 gnd 0.01275f
C1389 commonsourceibias.t148 gnd 0.191194f
C1390 commonsourceibias.n371 gnd 0.085058f
C1391 commonsourceibias.n372 gnd 0.030353f
C1392 commonsourceibias.n373 gnd 0.53129f
C1393 commonsourceibias.n374 gnd 0.012626f
C1394 commonsourceibias.t153 gnd 0.191194f
C1395 commonsourceibias.t104 gnd 0.176786f
C1396 commonsourceibias.n375 gnd 0.007691f
C1397 commonsourceibias.n376 gnd 0.009462f
C1398 commonsourceibias.t73 gnd 0.176786f
C1399 commonsourceibias.n377 gnd 0.009599f
C1400 commonsourceibias.n378 gnd 0.009462f
C1401 commonsourceibias.t90 gnd 0.176786f
C1402 commonsourceibias.n379 gnd 0.007654f
C1403 commonsourceibias.n380 gnd 0.009462f
C1404 commonsourceibias.t151 gnd 0.176786f
C1405 commonsourceibias.n381 gnd 0.009135f
C1406 commonsourceibias.n382 gnd 0.009462f
C1407 commonsourceibias.t91 gnd 0.176786f
C1408 commonsourceibias.n383 gnd 0.007642f
C1409 commonsourceibias.n384 gnd 0.009462f
C1410 commonsourceibias.t119 gnd 0.176786f
C1411 commonsourceibias.t87 gnd 0.176786f
C1412 commonsourceibias.n385 gnd 0.070538f
C1413 commonsourceibias.n386 gnd 0.009462f
C1414 commonsourceibias.t79 gnd 0.176786f
C1415 commonsourceibias.n387 gnd 0.070538f
C1416 commonsourceibias.n388 gnd 0.009462f
C1417 commonsourceibias.t95 gnd 0.176786f
C1418 commonsourceibias.n389 gnd 0.070538f
C1419 commonsourceibias.n390 gnd 0.009462f
C1420 commonsourceibias.t88 gnd 0.176786f
C1421 commonsourceibias.n391 gnd 0.010756f
C1422 commonsourceibias.n392 gnd 0.009462f
C1423 commonsourceibias.t65 gnd 0.176786f
C1424 commonsourceibias.n393 gnd 0.012719f
C1425 commonsourceibias.t83 gnd 0.196936f
C1426 commonsourceibias.t84 gnd 0.176786f
C1427 commonsourceibias.n394 gnd 0.078597f
C1428 commonsourceibias.n395 gnd 0.084205f
C1429 commonsourceibias.n396 gnd 0.040277f
C1430 commonsourceibias.n397 gnd 0.009462f
C1431 commonsourceibias.n398 gnd 0.007691f
C1432 commonsourceibias.n399 gnd 0.013039f
C1433 commonsourceibias.n400 gnd 0.070538f
C1434 commonsourceibias.n401 gnd 0.013095f
C1435 commonsourceibias.n402 gnd 0.009462f
C1436 commonsourceibias.n403 gnd 0.009462f
C1437 commonsourceibias.n404 gnd 0.009462f
C1438 commonsourceibias.n405 gnd 0.009599f
C1439 commonsourceibias.n406 gnd 0.070538f
C1440 commonsourceibias.n407 gnd 0.011663f
C1441 commonsourceibias.n408 gnd 0.012902f
C1442 commonsourceibias.n409 gnd 0.009462f
C1443 commonsourceibias.n410 gnd 0.009462f
C1444 commonsourceibias.n411 gnd 0.012818f
C1445 commonsourceibias.n412 gnd 0.007654f
C1446 commonsourceibias.n413 gnd 0.012977f
C1447 commonsourceibias.n414 gnd 0.009462f
C1448 commonsourceibias.n415 gnd 0.009462f
C1449 commonsourceibias.n416 gnd 0.013056f
C1450 commonsourceibias.n417 gnd 0.011258f
C1451 commonsourceibias.n418 gnd 0.009135f
C1452 commonsourceibias.n419 gnd 0.009462f
C1453 commonsourceibias.n420 gnd 0.009462f
C1454 commonsourceibias.n421 gnd 0.011574f
C1455 commonsourceibias.n422 gnd 0.012991f
C1456 commonsourceibias.n423 gnd 0.070538f
C1457 commonsourceibias.n424 gnd 0.012903f
C1458 commonsourceibias.n425 gnd 0.009417f
C1459 commonsourceibias.t51 gnd 0.020419f
C1460 commonsourceibias.t49 gnd 0.020419f
C1461 commonsourceibias.n426 gnd 0.181032f
C1462 commonsourceibias.t43 gnd 0.020419f
C1463 commonsourceibias.t37 gnd 0.020419f
C1464 commonsourceibias.n427 gnd 0.180428f
C1465 commonsourceibias.n428 gnd 0.168125f
C1466 commonsourceibias.t1 gnd 0.020419f
C1467 commonsourceibias.t61 gnd 0.020419f
C1468 commonsourceibias.n429 gnd 0.180428f
C1469 commonsourceibias.n430 gnd 0.082878f
C1470 commonsourceibias.t39 gnd 0.020419f
C1471 commonsourceibias.t13 gnd 0.020419f
C1472 commonsourceibias.n431 gnd 0.180428f
C1473 commonsourceibias.n432 gnd 0.06924f
C1474 commonsourceibias.n433 gnd 0.012626f
C1475 commonsourceibias.t24 gnd 0.176786f
C1476 commonsourceibias.n434 gnd 0.007691f
C1477 commonsourceibias.n435 gnd 0.009462f
C1478 commonsourceibias.t32 gnd 0.176786f
C1479 commonsourceibias.n436 gnd 0.009599f
C1480 commonsourceibias.n437 gnd 0.009462f
C1481 commonsourceibias.t34 gnd 0.176786f
C1482 commonsourceibias.n438 gnd 0.007654f
C1483 commonsourceibias.n439 gnd 0.009462f
C1484 commonsourceibias.t26 gnd 0.176786f
C1485 commonsourceibias.n440 gnd 0.009135f
C1486 commonsourceibias.n441 gnd 0.009462f
C1487 commonsourceibias.t62 gnd 0.176786f
C1488 commonsourceibias.n442 gnd 0.007642f
C1489 commonsourceibias.n443 gnd 0.009462f
C1490 commonsourceibias.t12 gnd 0.176786f
C1491 commonsourceibias.t38 gnd 0.176786f
C1492 commonsourceibias.n444 gnd 0.070538f
C1493 commonsourceibias.n445 gnd 0.009462f
C1494 commonsourceibias.t60 gnd 0.176786f
C1495 commonsourceibias.n446 gnd 0.070538f
C1496 commonsourceibias.n447 gnd 0.009462f
C1497 commonsourceibias.t0 gnd 0.176786f
C1498 commonsourceibias.n448 gnd 0.070538f
C1499 commonsourceibias.n449 gnd 0.009462f
C1500 commonsourceibias.t36 gnd 0.176786f
C1501 commonsourceibias.n450 gnd 0.010756f
C1502 commonsourceibias.n451 gnd 0.009462f
C1503 commonsourceibias.t42 gnd 0.176786f
C1504 commonsourceibias.n452 gnd 0.012719f
C1505 commonsourceibias.t50 gnd 0.196936f
C1506 commonsourceibias.t48 gnd 0.176786f
C1507 commonsourceibias.n453 gnd 0.078597f
C1508 commonsourceibias.n454 gnd 0.084205f
C1509 commonsourceibias.n455 gnd 0.040277f
C1510 commonsourceibias.n456 gnd 0.009462f
C1511 commonsourceibias.n457 gnd 0.007691f
C1512 commonsourceibias.n458 gnd 0.013039f
C1513 commonsourceibias.n459 gnd 0.070538f
C1514 commonsourceibias.n460 gnd 0.013095f
C1515 commonsourceibias.n461 gnd 0.009462f
C1516 commonsourceibias.n462 gnd 0.009462f
C1517 commonsourceibias.n463 gnd 0.009462f
C1518 commonsourceibias.n464 gnd 0.009599f
C1519 commonsourceibias.n465 gnd 0.070538f
C1520 commonsourceibias.n466 gnd 0.011663f
C1521 commonsourceibias.n467 gnd 0.012902f
C1522 commonsourceibias.n468 gnd 0.009462f
C1523 commonsourceibias.n469 gnd 0.009462f
C1524 commonsourceibias.n470 gnd 0.012818f
C1525 commonsourceibias.n471 gnd 0.007654f
C1526 commonsourceibias.n472 gnd 0.012977f
C1527 commonsourceibias.n473 gnd 0.009462f
C1528 commonsourceibias.n474 gnd 0.009462f
C1529 commonsourceibias.n475 gnd 0.013056f
C1530 commonsourceibias.n476 gnd 0.011258f
C1531 commonsourceibias.n477 gnd 0.009135f
C1532 commonsourceibias.n478 gnd 0.009462f
C1533 commonsourceibias.n479 gnd 0.009462f
C1534 commonsourceibias.n480 gnd 0.011574f
C1535 commonsourceibias.n481 gnd 0.012991f
C1536 commonsourceibias.n482 gnd 0.070538f
C1537 commonsourceibias.n483 gnd 0.012903f
C1538 commonsourceibias.n484 gnd 0.009462f
C1539 commonsourceibias.n485 gnd 0.009462f
C1540 commonsourceibias.n486 gnd 0.009462f
C1541 commonsourceibias.n487 gnd 0.012903f
C1542 commonsourceibias.n488 gnd 0.070538f
C1543 commonsourceibias.n489 gnd 0.012991f
C1544 commonsourceibias.t6 gnd 0.176786f
C1545 commonsourceibias.n490 gnd 0.070538f
C1546 commonsourceibias.n491 gnd 0.011574f
C1547 commonsourceibias.n492 gnd 0.009462f
C1548 commonsourceibias.n493 gnd 0.009462f
C1549 commonsourceibias.n494 gnd 0.009462f
C1550 commonsourceibias.n495 gnd 0.011258f
C1551 commonsourceibias.n496 gnd 0.013056f
C1552 commonsourceibias.n497 gnd 0.070538f
C1553 commonsourceibias.n498 gnd 0.012977f
C1554 commonsourceibias.n499 gnd 0.009462f
C1555 commonsourceibias.n500 gnd 0.009462f
C1556 commonsourceibias.n501 gnd 0.009462f
C1557 commonsourceibias.n502 gnd 0.012818f
C1558 commonsourceibias.n503 gnd 0.070538f
C1559 commonsourceibias.n504 gnd 0.012902f
C1560 commonsourceibias.t10 gnd 0.176786f
C1561 commonsourceibias.n505 gnd 0.070538f
C1562 commonsourceibias.n506 gnd 0.011663f
C1563 commonsourceibias.n507 gnd 0.009462f
C1564 commonsourceibias.n508 gnd 0.009462f
C1565 commonsourceibias.n509 gnd 0.009462f
C1566 commonsourceibias.n510 gnd 0.010756f
C1567 commonsourceibias.n511 gnd 0.013095f
C1568 commonsourceibias.n512 gnd 0.070538f
C1569 commonsourceibias.n513 gnd 0.013039f
C1570 commonsourceibias.n514 gnd 0.009462f
C1571 commonsourceibias.n515 gnd 0.009462f
C1572 commonsourceibias.n516 gnd 0.009462f
C1573 commonsourceibias.n517 gnd 0.012719f
C1574 commonsourceibias.n518 gnd 0.070538f
C1575 commonsourceibias.n519 gnd 0.01275f
C1576 commonsourceibias.t40 gnd 0.191194f
C1577 commonsourceibias.n520 gnd 0.085058f
C1578 commonsourceibias.n521 gnd 0.095108f
C1579 commonsourceibias.t25 gnd 0.020419f
C1580 commonsourceibias.t41 gnd 0.020419f
C1581 commonsourceibias.n522 gnd 0.180428f
C1582 commonsourceibias.n523 gnd 0.15629f
C1583 commonsourceibias.t11 gnd 0.020419f
C1584 commonsourceibias.t33 gnd 0.020419f
C1585 commonsourceibias.n524 gnd 0.180428f
C1586 commonsourceibias.n525 gnd 0.082878f
C1587 commonsourceibias.t27 gnd 0.020419f
C1588 commonsourceibias.t35 gnd 0.020419f
C1589 commonsourceibias.n526 gnd 0.180428f
C1590 commonsourceibias.n527 gnd 0.082878f
C1591 commonsourceibias.t63 gnd 0.020419f
C1592 commonsourceibias.t7 gnd 0.020419f
C1593 commonsourceibias.n528 gnd 0.180428f
C1594 commonsourceibias.n529 gnd 0.06924f
C1595 commonsourceibias.n530 gnd 0.083843f
C1596 commonsourceibias.n531 gnd 0.068402f
C1597 commonsourceibias.n532 gnd 0.009417f
C1598 commonsourceibias.n533 gnd 0.012903f
C1599 commonsourceibias.n534 gnd 0.070538f
C1600 commonsourceibias.n535 gnd 0.012991f
C1601 commonsourceibias.t102 gnd 0.176786f
C1602 commonsourceibias.n536 gnd 0.070538f
C1603 commonsourceibias.n537 gnd 0.011574f
C1604 commonsourceibias.n538 gnd 0.009462f
C1605 commonsourceibias.n539 gnd 0.009462f
C1606 commonsourceibias.n540 gnd 0.009462f
C1607 commonsourceibias.n541 gnd 0.011258f
C1608 commonsourceibias.n542 gnd 0.013056f
C1609 commonsourceibias.n543 gnd 0.070538f
C1610 commonsourceibias.n544 gnd 0.012977f
C1611 commonsourceibias.n545 gnd 0.009462f
C1612 commonsourceibias.n546 gnd 0.009462f
C1613 commonsourceibias.n547 gnd 0.009462f
C1614 commonsourceibias.n548 gnd 0.012818f
C1615 commonsourceibias.n549 gnd 0.070538f
C1616 commonsourceibias.n550 gnd 0.012902f
C1617 commonsourceibias.t121 gnd 0.176786f
C1618 commonsourceibias.n551 gnd 0.070538f
C1619 commonsourceibias.n552 gnd 0.011663f
C1620 commonsourceibias.n553 gnd 0.009462f
C1621 commonsourceibias.n554 gnd 0.009462f
C1622 commonsourceibias.n555 gnd 0.009462f
C1623 commonsourceibias.n556 gnd 0.010756f
C1624 commonsourceibias.n557 gnd 0.013095f
C1625 commonsourceibias.n558 gnd 0.070538f
C1626 commonsourceibias.n559 gnd 0.013039f
C1627 commonsourceibias.n560 gnd 0.009462f
C1628 commonsourceibias.n561 gnd 0.009462f
C1629 commonsourceibias.n562 gnd 0.009462f
C1630 commonsourceibias.n563 gnd 0.012719f
C1631 commonsourceibias.n564 gnd 0.070538f
C1632 commonsourceibias.n565 gnd 0.01275f
C1633 commonsourceibias.n566 gnd 0.085058f
C1634 commonsourceibias.n567 gnd 0.056191f
C1635 commonsourceibias.n568 gnd 0.012626f
C1636 commonsourceibias.t118 gnd 0.176786f
C1637 commonsourceibias.n569 gnd 0.007691f
C1638 commonsourceibias.n570 gnd 0.009462f
C1639 commonsourceibias.t109 gnd 0.176786f
C1640 commonsourceibias.n571 gnd 0.009599f
C1641 commonsourceibias.n572 gnd 0.009462f
C1642 commonsourceibias.t117 gnd 0.176786f
C1643 commonsourceibias.n573 gnd 0.007654f
C1644 commonsourceibias.n574 gnd 0.009462f
C1645 commonsourceibias.t108 gnd 0.176786f
C1646 commonsourceibias.n575 gnd 0.009135f
C1647 commonsourceibias.n576 gnd 0.009462f
C1648 commonsourceibias.t122 gnd 0.176786f
C1649 commonsourceibias.n577 gnd 0.007642f
C1650 commonsourceibias.n578 gnd 0.009462f
C1651 commonsourceibias.t107 gnd 0.176786f
C1652 commonsourceibias.t129 gnd 0.176786f
C1653 commonsourceibias.n579 gnd 0.070538f
C1654 commonsourceibias.n580 gnd 0.009462f
C1655 commonsourceibias.t156 gnd 0.176786f
C1656 commonsourceibias.n581 gnd 0.070538f
C1657 commonsourceibias.n582 gnd 0.009462f
C1658 commonsourceibias.t105 gnd 0.176786f
C1659 commonsourceibias.n583 gnd 0.070538f
C1660 commonsourceibias.n584 gnd 0.009462f
C1661 commonsourceibias.t137 gnd 0.176786f
C1662 commonsourceibias.n585 gnd 0.010756f
C1663 commonsourceibias.n586 gnd 0.009462f
C1664 commonsourceibias.t155 gnd 0.176786f
C1665 commonsourceibias.n587 gnd 0.012719f
C1666 commonsourceibias.t131 gnd 0.196936f
C1667 commonsourceibias.t142 gnd 0.176786f
C1668 commonsourceibias.n588 gnd 0.078597f
C1669 commonsourceibias.n589 gnd 0.084205f
C1670 commonsourceibias.n590 gnd 0.040277f
C1671 commonsourceibias.n591 gnd 0.009462f
C1672 commonsourceibias.n592 gnd 0.007691f
C1673 commonsourceibias.n593 gnd 0.013039f
C1674 commonsourceibias.n594 gnd 0.070538f
C1675 commonsourceibias.n595 gnd 0.013095f
C1676 commonsourceibias.n596 gnd 0.009462f
C1677 commonsourceibias.n597 gnd 0.009462f
C1678 commonsourceibias.n598 gnd 0.009462f
C1679 commonsourceibias.n599 gnd 0.009599f
C1680 commonsourceibias.n600 gnd 0.070538f
C1681 commonsourceibias.n601 gnd 0.011663f
C1682 commonsourceibias.n602 gnd 0.012902f
C1683 commonsourceibias.n603 gnd 0.009462f
C1684 commonsourceibias.n604 gnd 0.009462f
C1685 commonsourceibias.n605 gnd 0.012818f
C1686 commonsourceibias.n606 gnd 0.007654f
C1687 commonsourceibias.n607 gnd 0.012977f
C1688 commonsourceibias.n608 gnd 0.009462f
C1689 commonsourceibias.n609 gnd 0.009462f
C1690 commonsourceibias.n610 gnd 0.013056f
C1691 commonsourceibias.n611 gnd 0.011258f
C1692 commonsourceibias.n612 gnd 0.009135f
C1693 commonsourceibias.n613 gnd 0.009462f
C1694 commonsourceibias.n614 gnd 0.009462f
C1695 commonsourceibias.n615 gnd 0.011574f
C1696 commonsourceibias.n616 gnd 0.012991f
C1697 commonsourceibias.n617 gnd 0.070538f
C1698 commonsourceibias.n618 gnd 0.012903f
C1699 commonsourceibias.n619 gnd 0.009462f
C1700 commonsourceibias.n620 gnd 0.009462f
C1701 commonsourceibias.n621 gnd 0.009462f
C1702 commonsourceibias.n622 gnd 0.012903f
C1703 commonsourceibias.n623 gnd 0.070538f
C1704 commonsourceibias.n624 gnd 0.012991f
C1705 commonsourceibias.t130 gnd 0.176786f
C1706 commonsourceibias.n625 gnd 0.070538f
C1707 commonsourceibias.n626 gnd 0.011574f
C1708 commonsourceibias.n627 gnd 0.009462f
C1709 commonsourceibias.n628 gnd 0.009462f
C1710 commonsourceibias.n629 gnd 0.009462f
C1711 commonsourceibias.n630 gnd 0.011258f
C1712 commonsourceibias.n631 gnd 0.013056f
C1713 commonsourceibias.n632 gnd 0.070538f
C1714 commonsourceibias.n633 gnd 0.012977f
C1715 commonsourceibias.n634 gnd 0.009462f
C1716 commonsourceibias.n635 gnd 0.009462f
C1717 commonsourceibias.n636 gnd 0.009462f
C1718 commonsourceibias.n637 gnd 0.012818f
C1719 commonsourceibias.n638 gnd 0.070538f
C1720 commonsourceibias.n639 gnd 0.012902f
C1721 commonsourceibias.t99 gnd 0.176786f
C1722 commonsourceibias.n640 gnd 0.070538f
C1723 commonsourceibias.n641 gnd 0.011663f
C1724 commonsourceibias.n642 gnd 0.009462f
C1725 commonsourceibias.n643 gnd 0.009462f
C1726 commonsourceibias.n644 gnd 0.009462f
C1727 commonsourceibias.n645 gnd 0.010756f
C1728 commonsourceibias.n646 gnd 0.013095f
C1729 commonsourceibias.n647 gnd 0.070538f
C1730 commonsourceibias.n648 gnd 0.013039f
C1731 commonsourceibias.n649 gnd 0.009462f
C1732 commonsourceibias.n650 gnd 0.009462f
C1733 commonsourceibias.n651 gnd 0.009462f
C1734 commonsourceibias.n652 gnd 0.012719f
C1735 commonsourceibias.n653 gnd 0.070538f
C1736 commonsourceibias.n654 gnd 0.01275f
C1737 commonsourceibias.t100 gnd 0.191194f
C1738 commonsourceibias.n655 gnd 0.085058f
C1739 commonsourceibias.n656 gnd 0.030353f
C1740 commonsourceibias.n657 gnd 0.151535f
C1741 commonsourceibias.n658 gnd 0.012626f
C1742 commonsourceibias.t86 gnd 0.176786f
C1743 commonsourceibias.n659 gnd 0.007691f
C1744 commonsourceibias.n660 gnd 0.009462f
C1745 commonsourceibias.t97 gnd 0.176786f
C1746 commonsourceibias.n661 gnd 0.009599f
C1747 commonsourceibias.n662 gnd 0.009462f
C1748 commonsourceibias.t77 gnd 0.176786f
C1749 commonsourceibias.n663 gnd 0.007654f
C1750 commonsourceibias.n664 gnd 0.009462f
C1751 commonsourceibias.t93 gnd 0.176786f
C1752 commonsourceibias.n665 gnd 0.009135f
C1753 commonsourceibias.n666 gnd 0.009462f
C1754 commonsourceibias.t145 gnd 0.176786f
C1755 commonsourceibias.n667 gnd 0.007642f
C1756 commonsourceibias.n668 gnd 0.009462f
C1757 commonsourceibias.t85 gnd 0.176786f
C1758 commonsourceibias.t98 gnd 0.176786f
C1759 commonsourceibias.n669 gnd 0.070538f
C1760 commonsourceibias.n670 gnd 0.009462f
C1761 commonsourceibias.t94 gnd 0.176786f
C1762 commonsourceibias.n671 gnd 0.070538f
C1763 commonsourceibias.n672 gnd 0.009462f
C1764 commonsourceibias.t76 gnd 0.176786f
C1765 commonsourceibias.n673 gnd 0.070538f
C1766 commonsourceibias.n674 gnd 0.009462f
C1767 commonsourceibias.t72 gnd 0.176786f
C1768 commonsourceibias.n675 gnd 0.010756f
C1769 commonsourceibias.n676 gnd 0.009462f
C1770 commonsourceibias.t89 gnd 0.176786f
C1771 commonsourceibias.n677 gnd 0.012719f
C1772 commonsourceibias.t144 gnd 0.196936f
C1773 commonsourceibias.t133 gnd 0.176786f
C1774 commonsourceibias.n678 gnd 0.078597f
C1775 commonsourceibias.n679 gnd 0.084205f
C1776 commonsourceibias.n680 gnd 0.040277f
C1777 commonsourceibias.n681 gnd 0.009462f
C1778 commonsourceibias.n682 gnd 0.007691f
C1779 commonsourceibias.n683 gnd 0.013039f
C1780 commonsourceibias.n684 gnd 0.070538f
C1781 commonsourceibias.n685 gnd 0.013095f
C1782 commonsourceibias.n686 gnd 0.009462f
C1783 commonsourceibias.n687 gnd 0.009462f
C1784 commonsourceibias.n688 gnd 0.009462f
C1785 commonsourceibias.n689 gnd 0.009599f
C1786 commonsourceibias.n690 gnd 0.070538f
C1787 commonsourceibias.n691 gnd 0.011663f
C1788 commonsourceibias.n692 gnd 0.012902f
C1789 commonsourceibias.n693 gnd 0.009462f
C1790 commonsourceibias.n694 gnd 0.009462f
C1791 commonsourceibias.n695 gnd 0.012818f
C1792 commonsourceibias.n696 gnd 0.007654f
C1793 commonsourceibias.n697 gnd 0.012977f
C1794 commonsourceibias.n698 gnd 0.009462f
C1795 commonsourceibias.n699 gnd 0.009462f
C1796 commonsourceibias.n700 gnd 0.013056f
C1797 commonsourceibias.n701 gnd 0.011258f
C1798 commonsourceibias.n702 gnd 0.009135f
C1799 commonsourceibias.n703 gnd 0.009462f
C1800 commonsourceibias.n704 gnd 0.009462f
C1801 commonsourceibias.n705 gnd 0.011574f
C1802 commonsourceibias.n706 gnd 0.012991f
C1803 commonsourceibias.n707 gnd 0.070538f
C1804 commonsourceibias.n708 gnd 0.012903f
C1805 commonsourceibias.n709 gnd 0.009462f
C1806 commonsourceibias.n710 gnd 0.009462f
C1807 commonsourceibias.n711 gnd 0.009462f
C1808 commonsourceibias.n712 gnd 0.012903f
C1809 commonsourceibias.n713 gnd 0.070538f
C1810 commonsourceibias.n714 gnd 0.012991f
C1811 commonsourceibias.t103 gnd 0.176786f
C1812 commonsourceibias.n715 gnd 0.070538f
C1813 commonsourceibias.n716 gnd 0.011574f
C1814 commonsourceibias.n717 gnd 0.009462f
C1815 commonsourceibias.n718 gnd 0.009462f
C1816 commonsourceibias.n719 gnd 0.009462f
C1817 commonsourceibias.n720 gnd 0.011258f
C1818 commonsourceibias.n721 gnd 0.013056f
C1819 commonsourceibias.n722 gnd 0.070538f
C1820 commonsourceibias.n723 gnd 0.012977f
C1821 commonsourceibias.n724 gnd 0.009462f
C1822 commonsourceibias.n725 gnd 0.009462f
C1823 commonsourceibias.n726 gnd 0.009462f
C1824 commonsourceibias.n727 gnd 0.012818f
C1825 commonsourceibias.n728 gnd 0.070538f
C1826 commonsourceibias.n729 gnd 0.012902f
C1827 commonsourceibias.t66 gnd 0.176786f
C1828 commonsourceibias.n730 gnd 0.070538f
C1829 commonsourceibias.n731 gnd 0.011663f
C1830 commonsourceibias.n732 gnd 0.009462f
C1831 commonsourceibias.n733 gnd 0.009462f
C1832 commonsourceibias.n734 gnd 0.009462f
C1833 commonsourceibias.n735 gnd 0.010756f
C1834 commonsourceibias.n736 gnd 0.013095f
C1835 commonsourceibias.n737 gnd 0.070538f
C1836 commonsourceibias.n738 gnd 0.013039f
C1837 commonsourceibias.n739 gnd 0.009462f
C1838 commonsourceibias.n740 gnd 0.009462f
C1839 commonsourceibias.n741 gnd 0.009462f
C1840 commonsourceibias.n742 gnd 0.012719f
C1841 commonsourceibias.n743 gnd 0.070538f
C1842 commonsourceibias.n744 gnd 0.01275f
C1843 commonsourceibias.t71 gnd 0.191194f
C1844 commonsourceibias.n745 gnd 0.085058f
C1845 commonsourceibias.n746 gnd 0.030353f
C1846 commonsourceibias.n747 gnd 0.199689f
C1847 commonsourceibias.n748 gnd 5.4246f
C1848 CSoutput.n0 gnd 0.048998f
C1849 CSoutput.t219 gnd 0.324111f
C1850 CSoutput.n1 gnd 0.146352f
C1851 CSoutput.n2 gnd 0.048998f
C1852 CSoutput.t223 gnd 0.324111f
C1853 CSoutput.n3 gnd 0.038835f
C1854 CSoutput.n4 gnd 0.048998f
C1855 CSoutput.t235 gnd 0.324111f
C1856 CSoutput.n5 gnd 0.033488f
C1857 CSoutput.n6 gnd 0.048998f
C1858 CSoutput.t221 gnd 0.324111f
C1859 CSoutput.t227 gnd 0.324111f
C1860 CSoutput.n7 gnd 0.144757f
C1861 CSoutput.n8 gnd 0.048998f
C1862 CSoutput.t225 gnd 0.324111f
C1863 CSoutput.n9 gnd 0.031929f
C1864 CSoutput.n10 gnd 0.048998f
C1865 CSoutput.t237 gnd 0.324111f
C1866 CSoutput.t224 gnd 0.324111f
C1867 CSoutput.n11 gnd 0.144757f
C1868 CSoutput.n12 gnd 0.048998f
C1869 CSoutput.t222 gnd 0.324111f
C1870 CSoutput.n13 gnd 0.033488f
C1871 CSoutput.n14 gnd 0.048998f
C1872 CSoutput.t234 gnd 0.324111f
C1873 CSoutput.t218 gnd 0.324111f
C1874 CSoutput.n15 gnd 0.144757f
C1875 CSoutput.n16 gnd 0.048998f
C1876 CSoutput.t220 gnd 0.324111f
C1877 CSoutput.n17 gnd 0.035766f
C1878 CSoutput.t230 gnd 0.387321f
C1879 CSoutput.t232 gnd 0.324111f
C1880 CSoutput.n18 gnd 0.184799f
C1881 CSoutput.n19 gnd 0.179319f
C1882 CSoutput.n20 gnd 0.208031f
C1883 CSoutput.n21 gnd 0.048998f
C1884 CSoutput.n22 gnd 0.040894f
C1885 CSoutput.n23 gnd 0.144757f
C1886 CSoutput.n24 gnd 0.039421f
C1887 CSoutput.n25 gnd 0.038835f
C1888 CSoutput.n26 gnd 0.048998f
C1889 CSoutput.n27 gnd 0.048998f
C1890 CSoutput.n28 gnd 0.04058f
C1891 CSoutput.n29 gnd 0.034453f
C1892 CSoutput.n30 gnd 0.14798f
C1893 CSoutput.n31 gnd 0.034928f
C1894 CSoutput.n32 gnd 0.048998f
C1895 CSoutput.n33 gnd 0.048998f
C1896 CSoutput.n34 gnd 0.048998f
C1897 CSoutput.n35 gnd 0.040148f
C1898 CSoutput.n36 gnd 0.144757f
C1899 CSoutput.n37 gnd 0.038395f
C1900 CSoutput.n38 gnd 0.03986f
C1901 CSoutput.n39 gnd 0.048998f
C1902 CSoutput.n40 gnd 0.048998f
C1903 CSoutput.n41 gnd 0.040886f
C1904 CSoutput.n42 gnd 0.03737f
C1905 CSoutput.n43 gnd 0.144757f
C1906 CSoutput.n44 gnd 0.038317f
C1907 CSoutput.n45 gnd 0.048998f
C1908 CSoutput.n46 gnd 0.048998f
C1909 CSoutput.n47 gnd 0.048998f
C1910 CSoutput.n48 gnd 0.038317f
C1911 CSoutput.n49 gnd 0.144757f
C1912 CSoutput.n50 gnd 0.03737f
C1913 CSoutput.n51 gnd 0.040886f
C1914 CSoutput.n52 gnd 0.048998f
C1915 CSoutput.n53 gnd 0.048998f
C1916 CSoutput.n54 gnd 0.03986f
C1917 CSoutput.n55 gnd 0.038395f
C1918 CSoutput.n56 gnd 0.144757f
C1919 CSoutput.n57 gnd 0.040148f
C1920 CSoutput.n58 gnd 0.048998f
C1921 CSoutput.n59 gnd 0.048998f
C1922 CSoutput.n60 gnd 0.048998f
C1923 CSoutput.n61 gnd 0.034928f
C1924 CSoutput.n62 gnd 0.14798f
C1925 CSoutput.n63 gnd 0.034453f
C1926 CSoutput.t229 gnd 0.324111f
C1927 CSoutput.n64 gnd 0.144757f
C1928 CSoutput.n65 gnd 0.04058f
C1929 CSoutput.n66 gnd 0.048998f
C1930 CSoutput.n67 gnd 0.048998f
C1931 CSoutput.n68 gnd 0.048998f
C1932 CSoutput.n69 gnd 0.039421f
C1933 CSoutput.n70 gnd 0.144757f
C1934 CSoutput.n71 gnd 0.040894f
C1935 CSoutput.n72 gnd 0.035766f
C1936 CSoutput.n73 gnd 0.048998f
C1937 CSoutput.n74 gnd 0.048998f
C1938 CSoutput.n75 gnd 0.037092f
C1939 CSoutput.n76 gnd 0.022029f
C1940 CSoutput.t231 gnd 0.364162f
C1941 CSoutput.n77 gnd 0.180901f
C1942 CSoutput.n78 gnd 0.740057f
C1943 CSoutput.t178 gnd 0.061118f
C1944 CSoutput.t76 gnd 0.061118f
C1945 CSoutput.n79 gnd 0.473197f
C1946 CSoutput.t158 gnd 0.061118f
C1947 CSoutput.t128 gnd 0.061118f
C1948 CSoutput.n80 gnd 0.472353f
C1949 CSoutput.n81 gnd 0.479438f
C1950 CSoutput.t167 gnd 0.061118f
C1951 CSoutput.t104 gnd 0.061118f
C1952 CSoutput.n82 gnd 0.472353f
C1953 CSoutput.n83 gnd 0.236247f
C1954 CSoutput.t186 gnd 0.061118f
C1955 CSoutput.t121 gnd 0.061118f
C1956 CSoutput.n84 gnd 0.472353f
C1957 CSoutput.n85 gnd 0.236247f
C1958 CSoutput.t82 gnd 0.061118f
C1959 CSoutput.t137 gnd 0.061118f
C1960 CSoutput.n86 gnd 0.472353f
C1961 CSoutput.n87 gnd 0.236247f
C1962 CSoutput.t87 gnd 0.061118f
C1963 CSoutput.t113 gnd 0.061118f
C1964 CSoutput.n88 gnd 0.472353f
C1965 CSoutput.n89 gnd 0.236247f
C1966 CSoutput.t191 gnd 0.061118f
C1967 CSoutput.t130 gnd 0.061118f
C1968 CSoutput.n90 gnd 0.472353f
C1969 CSoutput.n91 gnd 0.236247f
C1970 CSoutput.t90 gnd 0.061118f
C1971 CSoutput.t174 gnd 0.061118f
C1972 CSoutput.n92 gnd 0.472353f
C1973 CSoutput.n93 gnd 0.236247f
C1974 CSoutput.t100 gnd 0.061118f
C1975 CSoutput.t149 gnd 0.061118f
C1976 CSoutput.n94 gnd 0.472353f
C1977 CSoutput.n95 gnd 0.236247f
C1978 CSoutput.t116 gnd 0.061118f
C1979 CSoutput.t138 gnd 0.061118f
C1980 CSoutput.n96 gnd 0.472353f
C1981 CSoutput.n97 gnd 0.433222f
C1982 CSoutput.t171 gnd 0.061118f
C1983 CSoutput.t169 gnd 0.061118f
C1984 CSoutput.n98 gnd 0.473197f
C1985 CSoutput.t151 gnd 0.061118f
C1986 CSoutput.t83 gnd 0.061118f
C1987 CSoutput.n99 gnd 0.472353f
C1988 CSoutput.n100 gnd 0.479438f
C1989 CSoutput.t77 gnd 0.061118f
C1990 CSoutput.t165 gnd 0.061118f
C1991 CSoutput.n101 gnd 0.472353f
C1992 CSoutput.n102 gnd 0.236247f
C1993 CSoutput.t150 gnd 0.061118f
C1994 CSoutput.t123 gnd 0.061118f
C1995 CSoutput.n103 gnd 0.472353f
C1996 CSoutput.n104 gnd 0.236247f
C1997 CSoutput.t105 gnd 0.061118f
C1998 CSoutput.t181 gnd 0.061118f
C1999 CSoutput.n105 gnd 0.472353f
C2000 CSoutput.n106 gnd 0.236247f
C2001 CSoutput.t147 gnd 0.061118f
C2002 CSoutput.t146 gnd 0.061118f
C2003 CSoutput.n107 gnd 0.472353f
C2004 CSoutput.n108 gnd 0.236247f
C2005 CSoutput.t134 gnd 0.061118f
C2006 CSoutput.t101 gnd 0.061118f
C2007 CSoutput.n109 gnd 0.472353f
C2008 CSoutput.n110 gnd 0.236247f
C2009 CSoutput.t81 gnd 0.061118f
C2010 CSoutput.t135 gnd 0.061118f
C2011 CSoutput.n111 gnd 0.472353f
C2012 CSoutput.n112 gnd 0.236247f
C2013 CSoutput.t131 gnd 0.061118f
C2014 CSoutput.t99 gnd 0.061118f
C2015 CSoutput.n113 gnd 0.472353f
C2016 CSoutput.n114 gnd 0.236247f
C2017 CSoutput.t78 gnd 0.061118f
C2018 CSoutput.t75 gnd 0.061118f
C2019 CSoutput.n115 gnd 0.472353f
C2020 CSoutput.n116 gnd 0.352303f
C2021 CSoutput.n117 gnd 0.444252f
C2022 CSoutput.t183 gnd 0.061118f
C2023 CSoutput.t182 gnd 0.061118f
C2024 CSoutput.n118 gnd 0.473197f
C2025 CSoutput.t162 gnd 0.061118f
C2026 CSoutput.t96 gnd 0.061118f
C2027 CSoutput.n119 gnd 0.472353f
C2028 CSoutput.n120 gnd 0.479438f
C2029 CSoutput.t93 gnd 0.061118f
C2030 CSoutput.t180 gnd 0.061118f
C2031 CSoutput.n121 gnd 0.472353f
C2032 CSoutput.n122 gnd 0.236247f
C2033 CSoutput.t159 gnd 0.061118f
C2034 CSoutput.t136 gnd 0.061118f
C2035 CSoutput.n123 gnd 0.472353f
C2036 CSoutput.n124 gnd 0.236247f
C2037 CSoutput.t117 gnd 0.061118f
C2038 CSoutput.t192 gnd 0.061118f
C2039 CSoutput.n125 gnd 0.472353f
C2040 CSoutput.n126 gnd 0.236247f
C2041 CSoutput.t157 gnd 0.061118f
C2042 CSoutput.t156 gnd 0.061118f
C2043 CSoutput.n127 gnd 0.472353f
C2044 CSoutput.n128 gnd 0.236247f
C2045 CSoutput.t144 gnd 0.061118f
C2046 CSoutput.t114 gnd 0.061118f
C2047 CSoutput.n129 gnd 0.472353f
C2048 CSoutput.n130 gnd 0.236247f
C2049 CSoutput.t95 gnd 0.061118f
C2050 CSoutput.t145 gnd 0.061118f
C2051 CSoutput.n131 gnd 0.472353f
C2052 CSoutput.n132 gnd 0.236247f
C2053 CSoutput.t141 gnd 0.061118f
C2054 CSoutput.t112 gnd 0.061118f
C2055 CSoutput.n133 gnd 0.472353f
C2056 CSoutput.n134 gnd 0.236247f
C2057 CSoutput.t92 gnd 0.061118f
C2058 CSoutput.t91 gnd 0.061118f
C2059 CSoutput.n135 gnd 0.472353f
C2060 CSoutput.n136 gnd 0.352303f
C2061 CSoutput.n137 gnd 0.49656f
C2062 CSoutput.n138 gnd 9.73103f
C2063 CSoutput.n140 gnd 0.866766f
C2064 CSoutput.n141 gnd 0.650075f
C2065 CSoutput.n142 gnd 0.866766f
C2066 CSoutput.n143 gnd 0.866766f
C2067 CSoutput.n144 gnd 2.3336f
C2068 CSoutput.n145 gnd 0.866766f
C2069 CSoutput.n146 gnd 0.866766f
C2070 CSoutput.t216 gnd 1.08346f
C2071 CSoutput.n147 gnd 0.866766f
C2072 CSoutput.n148 gnd 0.866766f
C2073 CSoutput.n152 gnd 0.866766f
C2074 CSoutput.n156 gnd 0.866766f
C2075 CSoutput.n157 gnd 0.866766f
C2076 CSoutput.n159 gnd 0.866766f
C2077 CSoutput.n164 gnd 0.866766f
C2078 CSoutput.n166 gnd 0.866766f
C2079 CSoutput.n167 gnd 0.866766f
C2080 CSoutput.n169 gnd 0.866766f
C2081 CSoutput.n170 gnd 0.866766f
C2082 CSoutput.n172 gnd 0.866766f
C2083 CSoutput.t228 gnd 14.4836f
C2084 CSoutput.n174 gnd 0.866766f
C2085 CSoutput.n175 gnd 0.650075f
C2086 CSoutput.n176 gnd 0.866766f
C2087 CSoutput.n177 gnd 0.866766f
C2088 CSoutput.n178 gnd 2.3336f
C2089 CSoutput.n179 gnd 0.866766f
C2090 CSoutput.n180 gnd 0.866766f
C2091 CSoutput.t233 gnd 1.08346f
C2092 CSoutput.n181 gnd 0.866766f
C2093 CSoutput.n182 gnd 0.866766f
C2094 CSoutput.n186 gnd 0.866766f
C2095 CSoutput.n190 gnd 0.866766f
C2096 CSoutput.n191 gnd 0.866766f
C2097 CSoutput.n193 gnd 0.866766f
C2098 CSoutput.n198 gnd 0.866766f
C2099 CSoutput.n200 gnd 0.866766f
C2100 CSoutput.n201 gnd 0.866766f
C2101 CSoutput.n203 gnd 0.866766f
C2102 CSoutput.n204 gnd 0.866766f
C2103 CSoutput.n206 gnd 0.866766f
C2104 CSoutput.n207 gnd 0.650075f
C2105 CSoutput.n209 gnd 0.866766f
C2106 CSoutput.n210 gnd 0.650075f
C2107 CSoutput.n211 gnd 0.866766f
C2108 CSoutput.n212 gnd 0.866766f
C2109 CSoutput.n213 gnd 2.3336f
C2110 CSoutput.n214 gnd 0.866766f
C2111 CSoutput.n215 gnd 0.866766f
C2112 CSoutput.t226 gnd 1.08346f
C2113 CSoutput.n216 gnd 0.866766f
C2114 CSoutput.n217 gnd 2.3336f
C2115 CSoutput.n219 gnd 0.866766f
C2116 CSoutput.n220 gnd 0.866766f
C2117 CSoutput.n222 gnd 0.866766f
C2118 CSoutput.n223 gnd 0.866766f
C2119 CSoutput.t236 gnd 14.2475f
C2120 CSoutput.t217 gnd 14.4836f
C2121 CSoutput.n229 gnd 2.71917f
C2122 CSoutput.n230 gnd 11.0769f
C2123 CSoutput.n231 gnd 11.540401f
C2124 CSoutput.n236 gnd 2.9456f
C2125 CSoutput.n242 gnd 0.866766f
C2126 CSoutput.n244 gnd 0.866766f
C2127 CSoutput.n246 gnd 0.866766f
C2128 CSoutput.n248 gnd 0.866766f
C2129 CSoutput.n250 gnd 0.866766f
C2130 CSoutput.n256 gnd 0.866766f
C2131 CSoutput.n263 gnd 1.59018f
C2132 CSoutput.n264 gnd 1.59018f
C2133 CSoutput.n265 gnd 0.866766f
C2134 CSoutput.n266 gnd 0.866766f
C2135 CSoutput.n268 gnd 0.650075f
C2136 CSoutput.n269 gnd 0.556731f
C2137 CSoutput.n271 gnd 0.650075f
C2138 CSoutput.n272 gnd 0.556731f
C2139 CSoutput.n273 gnd 0.650075f
C2140 CSoutput.n275 gnd 0.866766f
C2141 CSoutput.n277 gnd 2.3336f
C2142 CSoutput.n278 gnd 2.71917f
C2143 CSoutput.n279 gnd 10.187901f
C2144 CSoutput.n281 gnd 0.650075f
C2145 CSoutput.n282 gnd 1.67268f
C2146 CSoutput.n283 gnd 0.650075f
C2147 CSoutput.n285 gnd 0.866766f
C2148 CSoutput.n287 gnd 2.3336f
C2149 CSoutput.n288 gnd 5.08296f
C2150 CSoutput.t74 gnd 0.061118f
C2151 CSoutput.t177 gnd 0.061118f
C2152 CSoutput.n289 gnd 0.473197f
C2153 CSoutput.t127 gnd 0.061118f
C2154 CSoutput.t190 gnd 0.061118f
C2155 CSoutput.n290 gnd 0.472353f
C2156 CSoutput.n291 gnd 0.479438f
C2157 CSoutput.t103 gnd 0.061118f
C2158 CSoutput.t166 gnd 0.061118f
C2159 CSoutput.n292 gnd 0.472353f
C2160 CSoutput.n293 gnd 0.236247f
C2161 CSoutput.t120 gnd 0.061118f
C2162 CSoutput.t185 gnd 0.061118f
C2163 CSoutput.n294 gnd 0.472353f
C2164 CSoutput.n295 gnd 0.236247f
C2165 CSoutput.t160 gnd 0.061118f
C2166 CSoutput.t80 gnd 0.061118f
C2167 CSoutput.n296 gnd 0.472353f
C2168 CSoutput.n297 gnd 0.236247f
C2169 CSoutput.t111 gnd 0.061118f
C2170 CSoutput.t86 gnd 0.061118f
C2171 CSoutput.n298 gnd 0.472353f
C2172 CSoutput.n299 gnd 0.236247f
C2173 CSoutput.t129 gnd 0.061118f
C2174 CSoutput.t108 gnd 0.061118f
C2175 CSoutput.n300 gnd 0.472353f
C2176 CSoutput.n301 gnd 0.236247f
C2177 CSoutput.t173 gnd 0.061118f
C2178 CSoutput.t89 gnd 0.061118f
C2179 CSoutput.n302 gnd 0.472353f
C2180 CSoutput.n303 gnd 0.236247f
C2181 CSoutput.t148 gnd 0.061118f
C2182 CSoutput.t97 gnd 0.061118f
C2183 CSoutput.n304 gnd 0.472353f
C2184 CSoutput.n305 gnd 0.236247f
C2185 CSoutput.t161 gnd 0.061118f
C2186 CSoutput.t115 gnd 0.061118f
C2187 CSoutput.n306 gnd 0.472353f
C2188 CSoutput.n307 gnd 0.433222f
C2189 CSoutput.t132 gnd 0.061118f
C2190 CSoutput.t133 gnd 0.061118f
C2191 CSoutput.n308 gnd 0.473197f
C2192 CSoutput.t155 gnd 0.061118f
C2193 CSoutput.t79 gnd 0.061118f
C2194 CSoutput.n309 gnd 0.472353f
C2195 CSoutput.n310 gnd 0.479438f
C2196 CSoutput.t126 gnd 0.061118f
C2197 CSoutput.t153 gnd 0.061118f
C2198 CSoutput.n311 gnd 0.472353f
C2199 CSoutput.n312 gnd 0.236247f
C2200 CSoutput.t73 gnd 0.061118f
C2201 CSoutput.t109 gnd 0.061118f
C2202 CSoutput.n313 gnd 0.472353f
C2203 CSoutput.n314 gnd 0.236247f
C2204 CSoutput.t110 gnd 0.061118f
C2205 CSoutput.t179 gnd 0.061118f
C2206 CSoutput.n315 gnd 0.472353f
C2207 CSoutput.n316 gnd 0.236247f
C2208 CSoutput.t106 gnd 0.061118f
C2209 CSoutput.t107 gnd 0.061118f
C2210 CSoutput.n317 gnd 0.472353f
C2211 CSoutput.n318 gnd 0.236247f
C2212 CSoutput.t175 gnd 0.061118f
C2213 CSoutput.t176 gnd 0.061118f
C2214 CSoutput.n319 gnd 0.472353f
C2215 CSoutput.n320 gnd 0.236247f
C2216 CSoutput.t85 gnd 0.061118f
C2217 CSoutput.t154 gnd 0.061118f
C2218 CSoutput.n321 gnd 0.472353f
C2219 CSoutput.n322 gnd 0.236247f
C2220 CSoutput.t172 gnd 0.061118f
C2221 CSoutput.t84 gnd 0.061118f
C2222 CSoutput.n323 gnd 0.472353f
C2223 CSoutput.n324 gnd 0.236247f
C2224 CSoutput.t125 gnd 0.061118f
C2225 CSoutput.t152 gnd 0.061118f
C2226 CSoutput.n325 gnd 0.472353f
C2227 CSoutput.n326 gnd 0.352303f
C2228 CSoutput.n327 gnd 0.444252f
C2229 CSoutput.t142 gnd 0.061118f
C2230 CSoutput.t143 gnd 0.061118f
C2231 CSoutput.n328 gnd 0.473197f
C2232 CSoutput.t170 gnd 0.061118f
C2233 CSoutput.t94 gnd 0.061118f
C2234 CSoutput.n329 gnd 0.472353f
C2235 CSoutput.n330 gnd 0.479438f
C2236 CSoutput.t139 gnd 0.061118f
C2237 CSoutput.t163 gnd 0.061118f
C2238 CSoutput.n331 gnd 0.472353f
C2239 CSoutput.n332 gnd 0.236247f
C2240 CSoutput.t88 gnd 0.061118f
C2241 CSoutput.t122 gnd 0.061118f
C2242 CSoutput.n333 gnd 0.472353f
C2243 CSoutput.n334 gnd 0.236247f
C2244 CSoutput.t124 gnd 0.061118f
C2245 CSoutput.t189 gnd 0.061118f
C2246 CSoutput.n335 gnd 0.472353f
C2247 CSoutput.n336 gnd 0.236247f
C2248 CSoutput.t118 gnd 0.061118f
C2249 CSoutput.t119 gnd 0.061118f
C2250 CSoutput.n337 gnd 0.472353f
C2251 CSoutput.n338 gnd 0.236247f
C2252 CSoutput.t187 gnd 0.061118f
C2253 CSoutput.t188 gnd 0.061118f
C2254 CSoutput.n339 gnd 0.472353f
C2255 CSoutput.n340 gnd 0.236247f
C2256 CSoutput.t102 gnd 0.061118f
C2257 CSoutput.t168 gnd 0.061118f
C2258 CSoutput.n341 gnd 0.472353f
C2259 CSoutput.n342 gnd 0.236247f
C2260 CSoutput.t184 gnd 0.061118f
C2261 CSoutput.t98 gnd 0.061118f
C2262 CSoutput.n343 gnd 0.472353f
C2263 CSoutput.n344 gnd 0.236247f
C2264 CSoutput.t140 gnd 0.061118f
C2265 CSoutput.t164 gnd 0.061118f
C2266 CSoutput.n345 gnd 0.472351f
C2267 CSoutput.n346 gnd 0.352305f
C2268 CSoutput.n347 gnd 0.49656f
C2269 CSoutput.n348 gnd 13.6443f
C2270 CSoutput.t19 gnd 0.053478f
C2271 CSoutput.t55 gnd 0.053478f
C2272 CSoutput.n349 gnd 0.474135f
C2273 CSoutput.t200 gnd 0.053478f
C2274 CSoutput.t0 gnd 0.053478f
C2275 CSoutput.n350 gnd 0.472553f
C2276 CSoutput.n351 gnd 0.440332f
C2277 CSoutput.t29 gnd 0.053478f
C2278 CSoutput.t15 gnd 0.053478f
C2279 CSoutput.n352 gnd 0.472553f
C2280 CSoutput.n353 gnd 0.217063f
C2281 CSoutput.t50 gnd 0.053478f
C2282 CSoutput.t207 gnd 0.053478f
C2283 CSoutput.n354 gnd 0.472553f
C2284 CSoutput.n355 gnd 0.217063f
C2285 CSoutput.t18 gnd 0.053478f
C2286 CSoutput.t16 gnd 0.053478f
C2287 CSoutput.n356 gnd 0.472553f
C2288 CSoutput.n357 gnd 0.217063f
C2289 CSoutput.t37 gnd 0.053478f
C2290 CSoutput.t203 gnd 0.053478f
C2291 CSoutput.n358 gnd 0.472553f
C2292 CSoutput.n359 gnd 0.217063f
C2293 CSoutput.t39 gnd 0.053478f
C2294 CSoutput.t35 gnd 0.053478f
C2295 CSoutput.n360 gnd 0.472553f
C2296 CSoutput.n361 gnd 0.217063f
C2297 CSoutput.t17 gnd 0.053478f
C2298 CSoutput.t41 gnd 0.053478f
C2299 CSoutput.n362 gnd 0.472553f
C2300 CSoutput.n363 gnd 0.40036f
C2301 CSoutput.t3 gnd 0.053478f
C2302 CSoutput.t215 gnd 0.053478f
C2303 CSoutput.n364 gnd 0.474135f
C2304 CSoutput.t214 gnd 0.053478f
C2305 CSoutput.t12 gnd 0.053478f
C2306 CSoutput.n365 gnd 0.472553f
C2307 CSoutput.n366 gnd 0.440332f
C2308 CSoutput.t26 gnd 0.053478f
C2309 CSoutput.t204 gnd 0.053478f
C2310 CSoutput.n367 gnd 0.472553f
C2311 CSoutput.n368 gnd 0.217063f
C2312 CSoutput.t64 gnd 0.053478f
C2313 CSoutput.t66 gnd 0.053478f
C2314 CSoutput.n369 gnd 0.472553f
C2315 CSoutput.n370 gnd 0.217063f
C2316 CSoutput.t10 gnd 0.053478f
C2317 CSoutput.t194 gnd 0.053478f
C2318 CSoutput.n371 gnd 0.472553f
C2319 CSoutput.n372 gnd 0.217063f
C2320 CSoutput.t197 gnd 0.053478f
C2321 CSoutput.t213 gnd 0.053478f
C2322 CSoutput.n373 gnd 0.472553f
C2323 CSoutput.n374 gnd 0.217063f
C2324 CSoutput.t72 gnd 0.053478f
C2325 CSoutput.t199 gnd 0.053478f
C2326 CSoutput.n375 gnd 0.472553f
C2327 CSoutput.n376 gnd 0.217063f
C2328 CSoutput.t6 gnd 0.053478f
C2329 CSoutput.t42 gnd 0.053478f
C2330 CSoutput.n377 gnd 0.472553f
C2331 CSoutput.n378 gnd 0.329548f
C2332 CSoutput.n379 gnd 0.415662f
C2333 CSoutput.t193 gnd 0.053478f
C2334 CSoutput.t198 gnd 0.053478f
C2335 CSoutput.n380 gnd 0.474135f
C2336 CSoutput.t23 gnd 0.053478f
C2337 CSoutput.t13 gnd 0.053478f
C2338 CSoutput.n381 gnd 0.472553f
C2339 CSoutput.n382 gnd 0.440332f
C2340 CSoutput.t58 gnd 0.053478f
C2341 CSoutput.t14 gnd 0.053478f
C2342 CSoutput.n383 gnd 0.472553f
C2343 CSoutput.n384 gnd 0.217063f
C2344 CSoutput.t40 gnd 0.053478f
C2345 CSoutput.t33 gnd 0.053478f
C2346 CSoutput.n385 gnd 0.472553f
C2347 CSoutput.n386 gnd 0.217063f
C2348 CSoutput.t210 gnd 0.053478f
C2349 CSoutput.t24 gnd 0.053478f
C2350 CSoutput.n387 gnd 0.472553f
C2351 CSoutput.n388 gnd 0.217063f
C2352 CSoutput.t47 gnd 0.053478f
C2353 CSoutput.t9 gnd 0.053478f
C2354 CSoutput.n389 gnd 0.472553f
C2355 CSoutput.n390 gnd 0.217063f
C2356 CSoutput.t8 gnd 0.053478f
C2357 CSoutput.t68 gnd 0.053478f
C2358 CSoutput.n391 gnd 0.472553f
C2359 CSoutput.n392 gnd 0.217063f
C2360 CSoutput.t208 gnd 0.053478f
C2361 CSoutput.t7 gnd 0.053478f
C2362 CSoutput.n393 gnd 0.472553f
C2363 CSoutput.n394 gnd 0.329548f
C2364 CSoutput.n395 gnd 0.446356f
C2365 CSoutput.n396 gnd 14.2415f
C2366 CSoutput.t70 gnd 0.053478f
C2367 CSoutput.t51 gnd 0.053478f
C2368 CSoutput.n397 gnd 0.474135f
C2369 CSoutput.t49 gnd 0.053478f
C2370 CSoutput.t53 gnd 0.053478f
C2371 CSoutput.n398 gnd 0.472553f
C2372 CSoutput.n399 gnd 0.440332f
C2373 CSoutput.t56 gnd 0.053478f
C2374 CSoutput.t61 gnd 0.053478f
C2375 CSoutput.n400 gnd 0.472553f
C2376 CSoutput.n401 gnd 0.217063f
C2377 CSoutput.t62 gnd 0.053478f
C2378 CSoutput.t211 gnd 0.053478f
C2379 CSoutput.n402 gnd 0.472553f
C2380 CSoutput.n403 gnd 0.217063f
C2381 CSoutput.t28 gnd 0.053478f
C2382 CSoutput.t202 gnd 0.053478f
C2383 CSoutput.n404 gnd 0.472553f
C2384 CSoutput.n405 gnd 0.217063f
C2385 CSoutput.t45 gnd 0.053478f
C2386 CSoutput.t20 gnd 0.053478f
C2387 CSoutput.n406 gnd 0.472553f
C2388 CSoutput.n407 gnd 0.217063f
C2389 CSoutput.t43 gnd 0.053478f
C2390 CSoutput.t205 gnd 0.053478f
C2391 CSoutput.n408 gnd 0.472553f
C2392 CSoutput.n409 gnd 0.217063f
C2393 CSoutput.t36 gnd 0.053478f
C2394 CSoutput.t31 gnd 0.053478f
C2395 CSoutput.n410 gnd 0.472553f
C2396 CSoutput.n411 gnd 0.40036f
C2397 CSoutput.t4 gnd 0.053478f
C2398 CSoutput.t2 gnd 0.053478f
C2399 CSoutput.n412 gnd 0.474135f
C2400 CSoutput.t46 gnd 0.053478f
C2401 CSoutput.t25 gnd 0.053478f
C2402 CSoutput.n413 gnd 0.472553f
C2403 CSoutput.n414 gnd 0.440332f
C2404 CSoutput.t21 gnd 0.053478f
C2405 CSoutput.t48 gnd 0.053478f
C2406 CSoutput.n415 gnd 0.472553f
C2407 CSoutput.n416 gnd 0.217063f
C2408 CSoutput.t212 gnd 0.053478f
C2409 CSoutput.t5 gnd 0.053478f
C2410 CSoutput.n417 gnd 0.472553f
C2411 CSoutput.n418 gnd 0.217063f
C2412 CSoutput.t65 gnd 0.053478f
C2413 CSoutput.t63 gnd 0.053478f
C2414 CSoutput.n419 gnd 0.472553f
C2415 CSoutput.n420 gnd 0.217063f
C2416 CSoutput.t54 gnd 0.053478f
C2417 CSoutput.t57 gnd 0.053478f
C2418 CSoutput.n421 gnd 0.472553f
C2419 CSoutput.n422 gnd 0.217063f
C2420 CSoutput.t195 gnd 0.053478f
C2421 CSoutput.t22 gnd 0.053478f
C2422 CSoutput.n423 gnd 0.472553f
C2423 CSoutput.n424 gnd 0.217063f
C2424 CSoutput.t196 gnd 0.053478f
C2425 CSoutput.t30 gnd 0.053478f
C2426 CSoutput.n425 gnd 0.472553f
C2427 CSoutput.n426 gnd 0.329548f
C2428 CSoutput.n427 gnd 0.415662f
C2429 CSoutput.t27 gnd 0.053478f
C2430 CSoutput.t69 gnd 0.053478f
C2431 CSoutput.n428 gnd 0.474135f
C2432 CSoutput.t209 gnd 0.053478f
C2433 CSoutput.t1 gnd 0.053478f
C2434 CSoutput.n429 gnd 0.472553f
C2435 CSoutput.n430 gnd 0.440332f
C2436 CSoutput.t38 gnd 0.053478f
C2437 CSoutput.t60 gnd 0.053478f
C2438 CSoutput.n431 gnd 0.472553f
C2439 CSoutput.n432 gnd 0.217063f
C2440 CSoutput.t71 gnd 0.053478f
C2441 CSoutput.t201 gnd 0.053478f
C2442 CSoutput.n433 gnd 0.472553f
C2443 CSoutput.n434 gnd 0.217063f
C2444 CSoutput.t67 gnd 0.053478f
C2445 CSoutput.t32 gnd 0.053478f
C2446 CSoutput.n435 gnd 0.472553f
C2447 CSoutput.n436 gnd 0.217063f
C2448 CSoutput.t59 gnd 0.053478f
C2449 CSoutput.t44 gnd 0.053478f
C2450 CSoutput.n437 gnd 0.472553f
C2451 CSoutput.n438 gnd 0.217063f
C2452 CSoutput.t206 gnd 0.053478f
C2453 CSoutput.t52 gnd 0.053478f
C2454 CSoutput.n439 gnd 0.472553f
C2455 CSoutput.n440 gnd 0.217063f
C2456 CSoutput.t11 gnd 0.053478f
C2457 CSoutput.t34 gnd 0.053478f
C2458 CSoutput.n441 gnd 0.472553f
C2459 CSoutput.n442 gnd 0.329548f
C2460 CSoutput.n443 gnd 0.446356f
C2461 CSoutput.n444 gnd 8.42933f
C2462 CSoutput.n445 gnd 14.9667f
C2463 vdd.t295 gnd 0.040751f
C2464 vdd.t93 gnd 0.040751f
C2465 vdd.n0 gnd 0.321411f
C2466 vdd.t126 gnd 0.040751f
C2467 vdd.t4 gnd 0.040751f
C2468 vdd.n1 gnd 0.32088f
C2469 vdd.n2 gnd 0.295913f
C2470 vdd.t128 gnd 0.040751f
C2471 vdd.t110 gnd 0.040751f
C2472 vdd.n3 gnd 0.32088f
C2473 vdd.n4 gnd 0.149654f
C2474 vdd.t95 gnd 0.040751f
C2475 vdd.t88 gnd 0.040751f
C2476 vdd.n5 gnd 0.32088f
C2477 vdd.n6 gnd 0.140423f
C2478 vdd.t123 gnd 0.040751f
C2479 vdd.t114 gnd 0.040751f
C2480 vdd.n7 gnd 0.321411f
C2481 vdd.t90 gnd 0.040751f
C2482 vdd.t2 gnd 0.040751f
C2483 vdd.n8 gnd 0.32088f
C2484 vdd.n9 gnd 0.295913f
C2485 vdd.t120 gnd 0.040751f
C2486 vdd.t98 gnd 0.040751f
C2487 vdd.n10 gnd 0.32088f
C2488 vdd.n11 gnd 0.149654f
C2489 vdd.t116 gnd 0.040751f
C2490 vdd.t6 gnd 0.040751f
C2491 vdd.n12 gnd 0.32088f
C2492 vdd.n13 gnd 0.140423f
C2493 vdd.n14 gnd 0.099276f
C2494 vdd.t104 gnd 0.022639f
C2495 vdd.t7 gnd 0.022639f
C2496 vdd.n15 gnd 0.208387f
C2497 vdd.t292 gnd 0.022639f
C2498 vdd.t100 gnd 0.022639f
C2499 vdd.n16 gnd 0.207777f
C2500 vdd.n17 gnd 0.361597f
C2501 vdd.t106 gnd 0.022639f
C2502 vdd.t117 gnd 0.022639f
C2503 vdd.n18 gnd 0.207777f
C2504 vdd.n19 gnd 0.149598f
C2505 vdd.t293 gnd 0.022639f
C2506 vdd.t8 gnd 0.022639f
C2507 vdd.n20 gnd 0.208387f
C2508 vdd.t105 gnd 0.022639f
C2509 vdd.t108 gnd 0.022639f
C2510 vdd.n21 gnd 0.207777f
C2511 vdd.n22 gnd 0.361597f
C2512 vdd.t9 gnd 0.022639f
C2513 vdd.t107 gnd 0.022639f
C2514 vdd.n23 gnd 0.207777f
C2515 vdd.n24 gnd 0.149598f
C2516 vdd.t101 gnd 0.022639f
C2517 vdd.t118 gnd 0.022639f
C2518 vdd.n25 gnd 0.207777f
C2519 vdd.t102 gnd 0.022639f
C2520 vdd.t291 gnd 0.022639f
C2521 vdd.n26 gnd 0.207777f
C2522 vdd.n27 gnd 22.996801f
C2523 vdd.n28 gnd 8.87883f
C2524 vdd.n29 gnd 0.006175f
C2525 vdd.n30 gnd 0.00573f
C2526 vdd.n31 gnd 0.00317f
C2527 vdd.n32 gnd 0.007278f
C2528 vdd.n33 gnd 0.003079f
C2529 vdd.n34 gnd 0.00326f
C2530 vdd.n35 gnd 0.00573f
C2531 vdd.n36 gnd 0.003079f
C2532 vdd.n37 gnd 0.007278f
C2533 vdd.n38 gnd 0.00326f
C2534 vdd.n39 gnd 0.00573f
C2535 vdd.n40 gnd 0.003079f
C2536 vdd.n41 gnd 0.005458f
C2537 vdd.n42 gnd 0.005474f
C2538 vdd.t138 gnd 0.015635f
C2539 vdd.n43 gnd 0.034788f
C2540 vdd.n44 gnd 0.181046f
C2541 vdd.n45 gnd 0.003079f
C2542 vdd.n46 gnd 0.00326f
C2543 vdd.n47 gnd 0.007278f
C2544 vdd.n48 gnd 0.007278f
C2545 vdd.n49 gnd 0.00326f
C2546 vdd.n50 gnd 0.003079f
C2547 vdd.n51 gnd 0.00573f
C2548 vdd.n52 gnd 0.00573f
C2549 vdd.n53 gnd 0.003079f
C2550 vdd.n54 gnd 0.00326f
C2551 vdd.n55 gnd 0.007278f
C2552 vdd.n56 gnd 0.007278f
C2553 vdd.n57 gnd 0.00326f
C2554 vdd.n58 gnd 0.003079f
C2555 vdd.n59 gnd 0.00573f
C2556 vdd.n60 gnd 0.00573f
C2557 vdd.n61 gnd 0.003079f
C2558 vdd.n62 gnd 0.00326f
C2559 vdd.n63 gnd 0.007278f
C2560 vdd.n64 gnd 0.007278f
C2561 vdd.n65 gnd 0.017206f
C2562 vdd.n66 gnd 0.00317f
C2563 vdd.n67 gnd 0.003079f
C2564 vdd.n68 gnd 0.01481f
C2565 vdd.n69 gnd 0.010339f
C2566 vdd.t275 gnd 0.036223f
C2567 vdd.t215 gnd 0.036223f
C2568 vdd.n70 gnd 0.248951f
C2569 vdd.n71 gnd 0.195762f
C2570 vdd.t288 gnd 0.036223f
C2571 vdd.t182 gnd 0.036223f
C2572 vdd.n72 gnd 0.248951f
C2573 vdd.n73 gnd 0.157979f
C2574 vdd.t265 gnd 0.036223f
C2575 vdd.t205 gnd 0.036223f
C2576 vdd.n74 gnd 0.248951f
C2577 vdd.n75 gnd 0.157979f
C2578 vdd.t283 gnd 0.036223f
C2579 vdd.t259 gnd 0.036223f
C2580 vdd.n76 gnd 0.248951f
C2581 vdd.n77 gnd 0.157979f
C2582 vdd.t152 gnd 0.036223f
C2583 vdd.t194 gnd 0.036223f
C2584 vdd.n78 gnd 0.248951f
C2585 vdd.n79 gnd 0.157979f
C2586 vdd.t159 gnd 0.036223f
C2587 vdd.t219 gnd 0.036223f
C2588 vdd.n80 gnd 0.248951f
C2589 vdd.n81 gnd 0.157979f
C2590 vdd.t189 gnd 0.036223f
C2591 vdd.t229 gnd 0.036223f
C2592 vdd.n82 gnd 0.248951f
C2593 vdd.n83 gnd 0.157979f
C2594 vdd.t164 gnd 0.036223f
C2595 vdd.t245 gnd 0.036223f
C2596 vdd.n84 gnd 0.248951f
C2597 vdd.n85 gnd 0.157979f
C2598 vdd.t172 gnd 0.036223f
C2599 vdd.t260 gnd 0.036223f
C2600 vdd.n86 gnd 0.248951f
C2601 vdd.n87 gnd 0.157979f
C2602 vdd.n88 gnd 0.006175f
C2603 vdd.n89 gnd 0.00573f
C2604 vdd.n90 gnd 0.00317f
C2605 vdd.n91 gnd 0.007278f
C2606 vdd.n92 gnd 0.003079f
C2607 vdd.n93 gnd 0.00326f
C2608 vdd.n94 gnd 0.00573f
C2609 vdd.n95 gnd 0.003079f
C2610 vdd.n96 gnd 0.007278f
C2611 vdd.n97 gnd 0.00326f
C2612 vdd.n98 gnd 0.00573f
C2613 vdd.n99 gnd 0.003079f
C2614 vdd.n100 gnd 0.005458f
C2615 vdd.n101 gnd 0.005474f
C2616 vdd.t200 gnd 0.015635f
C2617 vdd.n102 gnd 0.034788f
C2618 vdd.n103 gnd 0.181046f
C2619 vdd.n104 gnd 0.003079f
C2620 vdd.n105 gnd 0.00326f
C2621 vdd.n106 gnd 0.007278f
C2622 vdd.n107 gnd 0.007278f
C2623 vdd.n108 gnd 0.00326f
C2624 vdd.n109 gnd 0.003079f
C2625 vdd.n110 gnd 0.00573f
C2626 vdd.n111 gnd 0.00573f
C2627 vdd.n112 gnd 0.003079f
C2628 vdd.n113 gnd 0.00326f
C2629 vdd.n114 gnd 0.007278f
C2630 vdd.n115 gnd 0.007278f
C2631 vdd.n116 gnd 0.00326f
C2632 vdd.n117 gnd 0.003079f
C2633 vdd.n118 gnd 0.00573f
C2634 vdd.n119 gnd 0.00573f
C2635 vdd.n120 gnd 0.003079f
C2636 vdd.n121 gnd 0.00326f
C2637 vdd.n122 gnd 0.007278f
C2638 vdd.n123 gnd 0.007278f
C2639 vdd.n124 gnd 0.017206f
C2640 vdd.n125 gnd 0.00317f
C2641 vdd.n126 gnd 0.003079f
C2642 vdd.n127 gnd 0.01481f
C2643 vdd.n128 gnd 0.010015f
C2644 vdd.n129 gnd 0.117537f
C2645 vdd.n130 gnd 0.006175f
C2646 vdd.n131 gnd 0.00573f
C2647 vdd.n132 gnd 0.00317f
C2648 vdd.n133 gnd 0.007278f
C2649 vdd.n134 gnd 0.003079f
C2650 vdd.n135 gnd 0.00326f
C2651 vdd.n136 gnd 0.00573f
C2652 vdd.n137 gnd 0.003079f
C2653 vdd.n138 gnd 0.007278f
C2654 vdd.n139 gnd 0.00326f
C2655 vdd.n140 gnd 0.00573f
C2656 vdd.n141 gnd 0.003079f
C2657 vdd.n142 gnd 0.005458f
C2658 vdd.n143 gnd 0.005474f
C2659 vdd.t216 gnd 0.015635f
C2660 vdd.n144 gnd 0.034788f
C2661 vdd.n145 gnd 0.181046f
C2662 vdd.n146 gnd 0.003079f
C2663 vdd.n147 gnd 0.00326f
C2664 vdd.n148 gnd 0.007278f
C2665 vdd.n149 gnd 0.007278f
C2666 vdd.n150 gnd 0.00326f
C2667 vdd.n151 gnd 0.003079f
C2668 vdd.n152 gnd 0.00573f
C2669 vdd.n153 gnd 0.00573f
C2670 vdd.n154 gnd 0.003079f
C2671 vdd.n155 gnd 0.00326f
C2672 vdd.n156 gnd 0.007278f
C2673 vdd.n157 gnd 0.007278f
C2674 vdd.n158 gnd 0.00326f
C2675 vdd.n159 gnd 0.003079f
C2676 vdd.n160 gnd 0.00573f
C2677 vdd.n161 gnd 0.00573f
C2678 vdd.n162 gnd 0.003079f
C2679 vdd.n163 gnd 0.00326f
C2680 vdd.n164 gnd 0.007278f
C2681 vdd.n165 gnd 0.007278f
C2682 vdd.n166 gnd 0.017206f
C2683 vdd.n167 gnd 0.00317f
C2684 vdd.n168 gnd 0.003079f
C2685 vdd.n169 gnd 0.01481f
C2686 vdd.n170 gnd 0.010339f
C2687 vdd.t223 gnd 0.036223f
C2688 vdd.t255 gnd 0.036223f
C2689 vdd.n171 gnd 0.248951f
C2690 vdd.n172 gnd 0.195762f
C2691 vdd.t148 gnd 0.036223f
C2692 vdd.t213 gnd 0.036223f
C2693 vdd.n173 gnd 0.248951f
C2694 vdd.n174 gnd 0.157979f
C2695 vdd.t253 gnd 0.036223f
C2696 vdd.t132 gnd 0.036223f
C2697 vdd.n175 gnd 0.248951f
C2698 vdd.n176 gnd 0.157979f
C2699 vdd.t191 gnd 0.036223f
C2700 vdd.t193 gnd 0.036223f
C2701 vdd.n177 gnd 0.248951f
C2702 vdd.n178 gnd 0.157979f
C2703 vdd.t277 gnd 0.036223f
C2704 vdd.t186 gnd 0.036223f
C2705 vdd.n179 gnd 0.248951f
C2706 vdd.n180 gnd 0.157979f
C2707 vdd.t187 gnd 0.036223f
C2708 vdd.t273 gnd 0.036223f
C2709 vdd.n181 gnd 0.248951f
C2710 vdd.n182 gnd 0.157979f
C2711 vdd.t274 gnd 0.036223f
C2712 vdd.t136 gnd 0.036223f
C2713 vdd.n183 gnd 0.248951f
C2714 vdd.n184 gnd 0.157979f
C2715 vdd.t254 gnd 0.036223f
C2716 vdd.t271 gnd 0.036223f
C2717 vdd.n185 gnd 0.248951f
C2718 vdd.n186 gnd 0.157979f
C2719 vdd.t157 gnd 0.036223f
C2720 vdd.t212 gnd 0.036223f
C2721 vdd.n187 gnd 0.248951f
C2722 vdd.n188 gnd 0.157979f
C2723 vdd.n189 gnd 0.006175f
C2724 vdd.n190 gnd 0.00573f
C2725 vdd.n191 gnd 0.00317f
C2726 vdd.n192 gnd 0.007278f
C2727 vdd.n193 gnd 0.003079f
C2728 vdd.n194 gnd 0.00326f
C2729 vdd.n195 gnd 0.00573f
C2730 vdd.n196 gnd 0.003079f
C2731 vdd.n197 gnd 0.007278f
C2732 vdd.n198 gnd 0.00326f
C2733 vdd.n199 gnd 0.00573f
C2734 vdd.n200 gnd 0.003079f
C2735 vdd.n201 gnd 0.005458f
C2736 vdd.n202 gnd 0.005474f
C2737 vdd.t251 gnd 0.015635f
C2738 vdd.n203 gnd 0.034788f
C2739 vdd.n204 gnd 0.181046f
C2740 vdd.n205 gnd 0.003079f
C2741 vdd.n206 gnd 0.00326f
C2742 vdd.n207 gnd 0.007278f
C2743 vdd.n208 gnd 0.007278f
C2744 vdd.n209 gnd 0.00326f
C2745 vdd.n210 gnd 0.003079f
C2746 vdd.n211 gnd 0.00573f
C2747 vdd.n212 gnd 0.00573f
C2748 vdd.n213 gnd 0.003079f
C2749 vdd.n214 gnd 0.00326f
C2750 vdd.n215 gnd 0.007278f
C2751 vdd.n216 gnd 0.007278f
C2752 vdd.n217 gnd 0.00326f
C2753 vdd.n218 gnd 0.003079f
C2754 vdd.n219 gnd 0.00573f
C2755 vdd.n220 gnd 0.00573f
C2756 vdd.n221 gnd 0.003079f
C2757 vdd.n222 gnd 0.00326f
C2758 vdd.n223 gnd 0.007278f
C2759 vdd.n224 gnd 0.007278f
C2760 vdd.n225 gnd 0.017206f
C2761 vdd.n226 gnd 0.00317f
C2762 vdd.n227 gnd 0.003079f
C2763 vdd.n228 gnd 0.01481f
C2764 vdd.n229 gnd 0.010015f
C2765 vdd.n230 gnd 0.069923f
C2766 vdd.n231 gnd 0.25195f
C2767 vdd.n232 gnd 0.006175f
C2768 vdd.n233 gnd 0.00573f
C2769 vdd.n234 gnd 0.00317f
C2770 vdd.n235 gnd 0.007278f
C2771 vdd.n236 gnd 0.003079f
C2772 vdd.n237 gnd 0.00326f
C2773 vdd.n238 gnd 0.00573f
C2774 vdd.n239 gnd 0.003079f
C2775 vdd.n240 gnd 0.007278f
C2776 vdd.n241 gnd 0.00326f
C2777 vdd.n242 gnd 0.00573f
C2778 vdd.n243 gnd 0.003079f
C2779 vdd.n244 gnd 0.005458f
C2780 vdd.n245 gnd 0.005474f
C2781 vdd.t237 gnd 0.015635f
C2782 vdd.n246 gnd 0.034788f
C2783 vdd.n247 gnd 0.181046f
C2784 vdd.n248 gnd 0.003079f
C2785 vdd.n249 gnd 0.00326f
C2786 vdd.n250 gnd 0.007278f
C2787 vdd.n251 gnd 0.007278f
C2788 vdd.n252 gnd 0.00326f
C2789 vdd.n253 gnd 0.003079f
C2790 vdd.n254 gnd 0.00573f
C2791 vdd.n255 gnd 0.00573f
C2792 vdd.n256 gnd 0.003079f
C2793 vdd.n257 gnd 0.00326f
C2794 vdd.n258 gnd 0.007278f
C2795 vdd.n259 gnd 0.007278f
C2796 vdd.n260 gnd 0.00326f
C2797 vdd.n261 gnd 0.003079f
C2798 vdd.n262 gnd 0.00573f
C2799 vdd.n263 gnd 0.00573f
C2800 vdd.n264 gnd 0.003079f
C2801 vdd.n265 gnd 0.00326f
C2802 vdd.n266 gnd 0.007278f
C2803 vdd.n267 gnd 0.007278f
C2804 vdd.n268 gnd 0.017206f
C2805 vdd.n269 gnd 0.00317f
C2806 vdd.n270 gnd 0.003079f
C2807 vdd.n271 gnd 0.01481f
C2808 vdd.n272 gnd 0.010339f
C2809 vdd.t238 gnd 0.036223f
C2810 vdd.t268 gnd 0.036223f
C2811 vdd.n273 gnd 0.248951f
C2812 vdd.n274 gnd 0.195762f
C2813 vdd.t169 gnd 0.036223f
C2814 vdd.t233 gnd 0.036223f
C2815 vdd.n275 gnd 0.248951f
C2816 vdd.n276 gnd 0.157979f
C2817 vdd.t262 gnd 0.036223f
C2818 vdd.t162 gnd 0.036223f
C2819 vdd.n277 gnd 0.248951f
C2820 vdd.n278 gnd 0.157979f
C2821 vdd.t208 gnd 0.036223f
C2822 vdd.t210 gnd 0.036223f
C2823 vdd.n279 gnd 0.248951f
C2824 vdd.n280 gnd 0.157979f
C2825 vdd.t287 gnd 0.036223f
C2826 vdd.t203 gnd 0.036223f
C2827 vdd.n281 gnd 0.248951f
C2828 vdd.n282 gnd 0.157979f
C2829 vdd.t204 gnd 0.036223f
C2830 vdd.t285 gnd 0.036223f
C2831 vdd.n283 gnd 0.248951f
C2832 vdd.n284 gnd 0.157979f
C2833 vdd.t286 gnd 0.036223f
C2834 vdd.t180 gnd 0.036223f
C2835 vdd.n285 gnd 0.248951f
C2836 vdd.n286 gnd 0.157979f
C2837 vdd.t266 gnd 0.036223f
C2838 vdd.t282 gnd 0.036223f
C2839 vdd.n287 gnd 0.248951f
C2840 vdd.n288 gnd 0.157979f
C2841 vdd.t173 gnd 0.036223f
C2842 vdd.t235 gnd 0.036223f
C2843 vdd.n289 gnd 0.248951f
C2844 vdd.n290 gnd 0.157979f
C2845 vdd.n291 gnd 0.006175f
C2846 vdd.n292 gnd 0.00573f
C2847 vdd.n293 gnd 0.00317f
C2848 vdd.n294 gnd 0.007278f
C2849 vdd.n295 gnd 0.003079f
C2850 vdd.n296 gnd 0.00326f
C2851 vdd.n297 gnd 0.00573f
C2852 vdd.n298 gnd 0.003079f
C2853 vdd.n299 gnd 0.007278f
C2854 vdd.n300 gnd 0.00326f
C2855 vdd.n301 gnd 0.00573f
C2856 vdd.n302 gnd 0.003079f
C2857 vdd.n303 gnd 0.005458f
C2858 vdd.n304 gnd 0.005474f
C2859 vdd.t263 gnd 0.015635f
C2860 vdd.n305 gnd 0.034788f
C2861 vdd.n306 gnd 0.181046f
C2862 vdd.n307 gnd 0.003079f
C2863 vdd.n308 gnd 0.00326f
C2864 vdd.n309 gnd 0.007278f
C2865 vdd.n310 gnd 0.007278f
C2866 vdd.n311 gnd 0.00326f
C2867 vdd.n312 gnd 0.003079f
C2868 vdd.n313 gnd 0.00573f
C2869 vdd.n314 gnd 0.00573f
C2870 vdd.n315 gnd 0.003079f
C2871 vdd.n316 gnd 0.00326f
C2872 vdd.n317 gnd 0.007278f
C2873 vdd.n318 gnd 0.007278f
C2874 vdd.n319 gnd 0.00326f
C2875 vdd.n320 gnd 0.003079f
C2876 vdd.n321 gnd 0.00573f
C2877 vdd.n322 gnd 0.00573f
C2878 vdd.n323 gnd 0.003079f
C2879 vdd.n324 gnd 0.00326f
C2880 vdd.n325 gnd 0.007278f
C2881 vdd.n326 gnd 0.007278f
C2882 vdd.n327 gnd 0.017206f
C2883 vdd.n328 gnd 0.00317f
C2884 vdd.n329 gnd 0.003079f
C2885 vdd.n330 gnd 0.01481f
C2886 vdd.n331 gnd 0.010015f
C2887 vdd.n332 gnd 0.069923f
C2888 vdd.n333 gnd 0.288427f
C2889 vdd.n334 gnd 0.008647f
C2890 vdd.n335 gnd 0.011251f
C2891 vdd.n336 gnd 0.009056f
C2892 vdd.n337 gnd 0.009056f
C2893 vdd.n338 gnd 0.011251f
C2894 vdd.n339 gnd 0.011251f
C2895 vdd.n340 gnd 0.822116f
C2896 vdd.n341 gnd 0.011251f
C2897 vdd.n342 gnd 0.011251f
C2898 vdd.n343 gnd 0.011251f
C2899 vdd.n344 gnd 0.891105f
C2900 vdd.n345 gnd 0.011251f
C2901 vdd.n346 gnd 0.011251f
C2902 vdd.n347 gnd 0.011251f
C2903 vdd.n348 gnd 0.011251f
C2904 vdd.n349 gnd 0.009056f
C2905 vdd.n350 gnd 0.011251f
C2906 vdd.t218 gnd 0.574906f
C2907 vdd.n351 gnd 0.011251f
C2908 vdd.n352 gnd 0.011251f
C2909 vdd.n353 gnd 0.011251f
C2910 vdd.t135 gnd 0.574906f
C2911 vdd.n354 gnd 0.011251f
C2912 vdd.n355 gnd 0.011251f
C2913 vdd.n356 gnd 0.011251f
C2914 vdd.n357 gnd 0.011251f
C2915 vdd.n358 gnd 0.011251f
C2916 vdd.n359 gnd 0.009056f
C2917 vdd.n360 gnd 0.011251f
C2918 vdd.n361 gnd 0.649644f
C2919 vdd.n362 gnd 0.011251f
C2920 vdd.n363 gnd 0.011251f
C2921 vdd.n364 gnd 0.011251f
C2922 vdd.t244 gnd 0.574906f
C2923 vdd.n365 gnd 0.011251f
C2924 vdd.n366 gnd 0.011251f
C2925 vdd.n367 gnd 0.011251f
C2926 vdd.n368 gnd 0.011251f
C2927 vdd.n369 gnd 0.011251f
C2928 vdd.n370 gnd 0.009056f
C2929 vdd.n371 gnd 0.011251f
C2930 vdd.t156 gnd 0.574906f
C2931 vdd.n372 gnd 0.011251f
C2932 vdd.n373 gnd 0.011251f
C2933 vdd.n374 gnd 0.011251f
C2934 vdd.n375 gnd 0.67264f
C2935 vdd.n376 gnd 0.011251f
C2936 vdd.n377 gnd 0.011251f
C2937 vdd.n378 gnd 0.011251f
C2938 vdd.n379 gnd 0.011251f
C2939 vdd.n380 gnd 0.011251f
C2940 vdd.n381 gnd 0.009056f
C2941 vdd.n382 gnd 0.011251f
C2942 vdd.t199 gnd 0.574906f
C2943 vdd.n383 gnd 0.011251f
C2944 vdd.n384 gnd 0.011251f
C2945 vdd.n385 gnd 0.011251f
C2946 vdd.n386 gnd 0.580655f
C2947 vdd.n387 gnd 0.011251f
C2948 vdd.n388 gnd 0.011251f
C2949 vdd.n389 gnd 0.011251f
C2950 vdd.n390 gnd 0.011251f
C2951 vdd.n391 gnd 0.027217f
C2952 vdd.n392 gnd 0.027801f
C2953 vdd.t38 gnd 0.574906f
C2954 vdd.n393 gnd 0.027217f
C2955 vdd.n425 gnd 0.011251f
C2956 vdd.t40 gnd 0.138418f
C2957 vdd.t39 gnd 0.147931f
C2958 vdd.t37 gnd 0.180773f
C2959 vdd.n426 gnd 0.231725f
C2960 vdd.n427 gnd 0.195597f
C2961 vdd.n428 gnd 0.014852f
C2962 vdd.n429 gnd 0.011251f
C2963 vdd.n430 gnd 0.009056f
C2964 vdd.n431 gnd 0.011251f
C2965 vdd.n432 gnd 0.009056f
C2966 vdd.n433 gnd 0.011251f
C2967 vdd.n434 gnd 0.009056f
C2968 vdd.n435 gnd 0.011251f
C2969 vdd.n436 gnd 0.009056f
C2970 vdd.n437 gnd 0.011251f
C2971 vdd.n438 gnd 0.009056f
C2972 vdd.n439 gnd 0.011251f
C2973 vdd.t80 gnd 0.138418f
C2974 vdd.t79 gnd 0.147931f
C2975 vdd.t78 gnd 0.180773f
C2976 vdd.n440 gnd 0.231725f
C2977 vdd.n441 gnd 0.195597f
C2978 vdd.n442 gnd 0.009056f
C2979 vdd.n443 gnd 0.011251f
C2980 vdd.n444 gnd 0.009056f
C2981 vdd.n445 gnd 0.011251f
C2982 vdd.n446 gnd 0.009056f
C2983 vdd.n447 gnd 0.011251f
C2984 vdd.n448 gnd 0.009056f
C2985 vdd.n449 gnd 0.011251f
C2986 vdd.n450 gnd 0.009056f
C2987 vdd.n451 gnd 0.011251f
C2988 vdd.t86 gnd 0.138418f
C2989 vdd.t85 gnd 0.147931f
C2990 vdd.t84 gnd 0.180773f
C2991 vdd.n452 gnd 0.231725f
C2992 vdd.n453 gnd 0.195597f
C2993 vdd.n454 gnd 0.019379f
C2994 vdd.n455 gnd 0.011251f
C2995 vdd.n456 gnd 0.009056f
C2996 vdd.n457 gnd 0.011251f
C2997 vdd.n458 gnd 0.009056f
C2998 vdd.n459 gnd 0.011251f
C2999 vdd.n460 gnd 0.009056f
C3000 vdd.n461 gnd 0.011251f
C3001 vdd.n462 gnd 0.009056f
C3002 vdd.n463 gnd 0.011251f
C3003 vdd.n464 gnd 0.027801f
C3004 vdd.n465 gnd 0.007516f
C3005 vdd.n466 gnd 0.009056f
C3006 vdd.n467 gnd 0.011251f
C3007 vdd.n468 gnd 0.011251f
C3008 vdd.n469 gnd 0.009056f
C3009 vdd.n470 gnd 0.011251f
C3010 vdd.n471 gnd 0.011251f
C3011 vdd.n472 gnd 0.011251f
C3012 vdd.n473 gnd 0.011251f
C3013 vdd.n474 gnd 0.011251f
C3014 vdd.n475 gnd 0.009056f
C3015 vdd.n476 gnd 0.009056f
C3016 vdd.n477 gnd 0.011251f
C3017 vdd.n478 gnd 0.011251f
C3018 vdd.n479 gnd 0.009056f
C3019 vdd.n480 gnd 0.011251f
C3020 vdd.n481 gnd 0.011251f
C3021 vdd.n482 gnd 0.011251f
C3022 vdd.n483 gnd 0.011251f
C3023 vdd.n484 gnd 0.011251f
C3024 vdd.n485 gnd 0.009056f
C3025 vdd.n486 gnd 0.009056f
C3026 vdd.n487 gnd 0.011251f
C3027 vdd.n488 gnd 0.011251f
C3028 vdd.n489 gnd 0.009056f
C3029 vdd.n490 gnd 0.011251f
C3030 vdd.n491 gnd 0.011251f
C3031 vdd.n492 gnd 0.011251f
C3032 vdd.n493 gnd 0.011251f
C3033 vdd.n494 gnd 0.011251f
C3034 vdd.n495 gnd 0.009056f
C3035 vdd.n496 gnd 0.009056f
C3036 vdd.n497 gnd 0.011251f
C3037 vdd.n498 gnd 0.011251f
C3038 vdd.n499 gnd 0.009056f
C3039 vdd.n500 gnd 0.011251f
C3040 vdd.n501 gnd 0.011251f
C3041 vdd.n502 gnd 0.011251f
C3042 vdd.n503 gnd 0.011251f
C3043 vdd.n504 gnd 0.011251f
C3044 vdd.n505 gnd 0.009056f
C3045 vdd.n506 gnd 0.009056f
C3046 vdd.n507 gnd 0.011251f
C3047 vdd.n508 gnd 0.011251f
C3048 vdd.n509 gnd 0.007562f
C3049 vdd.n510 gnd 0.011251f
C3050 vdd.n511 gnd 0.011251f
C3051 vdd.n512 gnd 0.011251f
C3052 vdd.n513 gnd 0.011251f
C3053 vdd.n514 gnd 0.011251f
C3054 vdd.n515 gnd 0.007562f
C3055 vdd.n516 gnd 0.009056f
C3056 vdd.n517 gnd 0.011251f
C3057 vdd.n518 gnd 0.011251f
C3058 vdd.n519 gnd 0.009056f
C3059 vdd.n520 gnd 0.011251f
C3060 vdd.n521 gnd 0.011251f
C3061 vdd.n522 gnd 0.011251f
C3062 vdd.n523 gnd 0.011251f
C3063 vdd.n524 gnd 0.011251f
C3064 vdd.n525 gnd 0.009056f
C3065 vdd.n526 gnd 0.009056f
C3066 vdd.n527 gnd 0.011251f
C3067 vdd.n528 gnd 0.011251f
C3068 vdd.n529 gnd 0.009056f
C3069 vdd.n530 gnd 0.011251f
C3070 vdd.n531 gnd 0.011251f
C3071 vdd.n532 gnd 0.011251f
C3072 vdd.n533 gnd 0.011251f
C3073 vdd.n534 gnd 0.011251f
C3074 vdd.n535 gnd 0.009056f
C3075 vdd.n536 gnd 0.009056f
C3076 vdd.n537 gnd 0.011251f
C3077 vdd.n538 gnd 0.011251f
C3078 vdd.n539 gnd 0.009056f
C3079 vdd.n540 gnd 0.011251f
C3080 vdd.n541 gnd 0.011251f
C3081 vdd.n542 gnd 0.011251f
C3082 vdd.n543 gnd 0.011251f
C3083 vdd.n544 gnd 0.011251f
C3084 vdd.n545 gnd 0.009056f
C3085 vdd.n546 gnd 0.009056f
C3086 vdd.n547 gnd 0.011251f
C3087 vdd.n548 gnd 0.011251f
C3088 vdd.n549 gnd 0.009056f
C3089 vdd.n550 gnd 0.011251f
C3090 vdd.n551 gnd 0.011251f
C3091 vdd.n552 gnd 0.011251f
C3092 vdd.n553 gnd 0.011251f
C3093 vdd.n554 gnd 0.011251f
C3094 vdd.n555 gnd 0.009056f
C3095 vdd.n556 gnd 0.009056f
C3096 vdd.n557 gnd 0.011251f
C3097 vdd.n558 gnd 0.011251f
C3098 vdd.n559 gnd 0.009056f
C3099 vdd.n560 gnd 0.011251f
C3100 vdd.n561 gnd 0.011251f
C3101 vdd.n562 gnd 0.011251f
C3102 vdd.n563 gnd 0.011251f
C3103 vdd.n564 gnd 0.011251f
C3104 vdd.n565 gnd 0.006158f
C3105 vdd.n566 gnd 0.019379f
C3106 vdd.n567 gnd 0.011251f
C3107 vdd.n568 gnd 0.011251f
C3108 vdd.n569 gnd 0.008965f
C3109 vdd.n570 gnd 0.011251f
C3110 vdd.n571 gnd 0.011251f
C3111 vdd.n572 gnd 0.011251f
C3112 vdd.n573 gnd 0.011251f
C3113 vdd.n574 gnd 0.011251f
C3114 vdd.n575 gnd 0.009056f
C3115 vdd.n576 gnd 0.009056f
C3116 vdd.n577 gnd 0.011251f
C3117 vdd.n578 gnd 0.011251f
C3118 vdd.n579 gnd 0.009056f
C3119 vdd.n580 gnd 0.011251f
C3120 vdd.n581 gnd 0.011251f
C3121 vdd.n582 gnd 0.011251f
C3122 vdd.n583 gnd 0.011251f
C3123 vdd.n584 gnd 0.011251f
C3124 vdd.n585 gnd 0.009056f
C3125 vdd.n586 gnd 0.009056f
C3126 vdd.n587 gnd 0.011251f
C3127 vdd.n588 gnd 0.011251f
C3128 vdd.n589 gnd 0.009056f
C3129 vdd.n590 gnd 0.011251f
C3130 vdd.n591 gnd 0.011251f
C3131 vdd.n592 gnd 0.011251f
C3132 vdd.n593 gnd 0.011251f
C3133 vdd.n594 gnd 0.011251f
C3134 vdd.n595 gnd 0.009056f
C3135 vdd.n596 gnd 0.009056f
C3136 vdd.n597 gnd 0.011251f
C3137 vdd.n598 gnd 0.011251f
C3138 vdd.n599 gnd 0.009056f
C3139 vdd.n600 gnd 0.011251f
C3140 vdd.n601 gnd 0.011251f
C3141 vdd.n602 gnd 0.011251f
C3142 vdd.n603 gnd 0.011251f
C3143 vdd.n604 gnd 0.011251f
C3144 vdd.n605 gnd 0.009056f
C3145 vdd.n606 gnd 0.009056f
C3146 vdd.n607 gnd 0.011251f
C3147 vdd.n608 gnd 0.011251f
C3148 vdd.n609 gnd 0.009056f
C3149 vdd.n610 gnd 0.011251f
C3150 vdd.n611 gnd 0.011251f
C3151 vdd.n612 gnd 0.011251f
C3152 vdd.n613 gnd 0.011251f
C3153 vdd.n614 gnd 0.011251f
C3154 vdd.n615 gnd 0.009056f
C3155 vdd.n616 gnd 0.011251f
C3156 vdd.n617 gnd 0.009056f
C3157 vdd.n618 gnd 0.004754f
C3158 vdd.n619 gnd 0.011251f
C3159 vdd.n620 gnd 0.011251f
C3160 vdd.n621 gnd 0.009056f
C3161 vdd.n622 gnd 0.011251f
C3162 vdd.n623 gnd 0.009056f
C3163 vdd.n624 gnd 0.011251f
C3164 vdd.n625 gnd 0.009056f
C3165 vdd.n626 gnd 0.011251f
C3166 vdd.n627 gnd 0.009056f
C3167 vdd.n628 gnd 0.011251f
C3168 vdd.n629 gnd 0.009056f
C3169 vdd.n630 gnd 0.011251f
C3170 vdd.n631 gnd 0.009056f
C3171 vdd.n632 gnd 0.011251f
C3172 vdd.n633 gnd 0.626648f
C3173 vdd.t151 gnd 0.574906f
C3174 vdd.n634 gnd 0.011251f
C3175 vdd.n635 gnd 0.009056f
C3176 vdd.n636 gnd 0.011251f
C3177 vdd.n637 gnd 0.009056f
C3178 vdd.n638 gnd 0.011251f
C3179 vdd.t190 gnd 0.574906f
C3180 vdd.n639 gnd 0.011251f
C3181 vdd.n640 gnd 0.009056f
C3182 vdd.n641 gnd 0.011251f
C3183 vdd.n642 gnd 0.009056f
C3184 vdd.n643 gnd 0.011251f
C3185 vdd.t131 gnd 0.574906f
C3186 vdd.n644 gnd 0.718633f
C3187 vdd.n645 gnd 0.011251f
C3188 vdd.n646 gnd 0.009056f
C3189 vdd.n647 gnd 0.011251f
C3190 vdd.n648 gnd 0.009056f
C3191 vdd.n649 gnd 0.011251f
C3192 vdd.t252 gnd 0.574906f
C3193 vdd.n650 gnd 0.011251f
C3194 vdd.n651 gnd 0.009056f
C3195 vdd.n652 gnd 0.011251f
C3196 vdd.n653 gnd 0.009056f
C3197 vdd.n654 gnd 0.011251f
C3198 vdd.n655 gnd 0.79912f
C3199 vdd.n656 gnd 0.954345f
C3200 vdd.t181 gnd 0.574906f
C3201 vdd.n657 gnd 0.011251f
C3202 vdd.n658 gnd 0.009056f
C3203 vdd.n659 gnd 0.011251f
C3204 vdd.n660 gnd 0.009056f
C3205 vdd.n661 gnd 0.011251f
C3206 vdd.n662 gnd 0.603652f
C3207 vdd.n663 gnd 0.011251f
C3208 vdd.n664 gnd 0.009056f
C3209 vdd.n665 gnd 0.011251f
C3210 vdd.n666 gnd 0.009056f
C3211 vdd.n667 gnd 0.011251f
C3212 vdd.t222 gnd 0.574906f
C3213 vdd.t214 gnd 0.574906f
C3214 vdd.n668 gnd 0.011251f
C3215 vdd.n669 gnd 0.009056f
C3216 vdd.n670 gnd 0.011251f
C3217 vdd.n671 gnd 0.009056f
C3218 vdd.n672 gnd 0.011251f
C3219 vdd.t137 gnd 0.574906f
C3220 vdd.n673 gnd 0.011251f
C3221 vdd.n674 gnd 0.009056f
C3222 vdd.n675 gnd 0.011251f
C3223 vdd.n676 gnd 0.009056f
C3224 vdd.n677 gnd 0.011251f
C3225 vdd.n678 gnd 1.14981f
C3226 vdd.n679 gnd 0.937097f
C3227 vdd.n680 gnd 0.011251f
C3228 vdd.n681 gnd 0.009056f
C3229 vdd.n682 gnd 0.027217f
C3230 vdd.n683 gnd 0.007516f
C3231 vdd.n684 gnd 0.027217f
C3232 vdd.t16 gnd 0.574906f
C3233 vdd.n685 gnd 0.027217f
C3234 vdd.n686 gnd 0.007516f
C3235 vdd.n687 gnd 0.009676f
C3236 vdd.t82 gnd 0.138418f
C3237 vdd.t83 gnd 0.147931f
C3238 vdd.t81 gnd 0.180773f
C3239 vdd.n688 gnd 0.231725f
C3240 vdd.n689 gnd 0.194691f
C3241 vdd.n690 gnd 0.013946f
C3242 vdd.n691 gnd 0.011251f
C3243 vdd.n692 gnd 7.92221f
C3244 vdd.n723 gnd 1.58099f
C3245 vdd.n724 gnd 0.011251f
C3246 vdd.n725 gnd 0.011251f
C3247 vdd.n726 gnd 0.027801f
C3248 vdd.n727 gnd 0.009676f
C3249 vdd.n728 gnd 0.011251f
C3250 vdd.n729 gnd 0.009056f
C3251 vdd.n730 gnd 0.007201f
C3252 vdd.n731 gnd 0.018385f
C3253 vdd.n732 gnd 0.009056f
C3254 vdd.n733 gnd 0.011251f
C3255 vdd.n734 gnd 0.011251f
C3256 vdd.n735 gnd 0.011251f
C3257 vdd.n736 gnd 0.011251f
C3258 vdd.n737 gnd 0.011251f
C3259 vdd.n738 gnd 0.011251f
C3260 vdd.n739 gnd 0.011251f
C3261 vdd.n740 gnd 0.011251f
C3262 vdd.n741 gnd 0.011251f
C3263 vdd.n742 gnd 0.011251f
C3264 vdd.n743 gnd 0.011251f
C3265 vdd.n744 gnd 0.011251f
C3266 vdd.n745 gnd 0.011251f
C3267 vdd.n746 gnd 0.011251f
C3268 vdd.n747 gnd 0.007562f
C3269 vdd.n748 gnd 0.011251f
C3270 vdd.n749 gnd 0.011251f
C3271 vdd.n750 gnd 0.011251f
C3272 vdd.n751 gnd 0.011251f
C3273 vdd.n752 gnd 0.011251f
C3274 vdd.n753 gnd 0.011251f
C3275 vdd.n754 gnd 0.011251f
C3276 vdd.n755 gnd 0.011251f
C3277 vdd.n756 gnd 0.011251f
C3278 vdd.n757 gnd 0.011251f
C3279 vdd.n758 gnd 0.011251f
C3280 vdd.n759 gnd 0.011251f
C3281 vdd.n760 gnd 0.011251f
C3282 vdd.n761 gnd 0.011251f
C3283 vdd.n762 gnd 0.011251f
C3284 vdd.n763 gnd 0.011251f
C3285 vdd.n764 gnd 0.011251f
C3286 vdd.n765 gnd 0.011251f
C3287 vdd.n766 gnd 0.011251f
C3288 vdd.n767 gnd 0.008965f
C3289 vdd.t17 gnd 0.138418f
C3290 vdd.t18 gnd 0.147931f
C3291 vdd.t15 gnd 0.180773f
C3292 vdd.n768 gnd 0.231725f
C3293 vdd.n769 gnd 0.194691f
C3294 vdd.n770 gnd 0.011251f
C3295 vdd.n771 gnd 0.011251f
C3296 vdd.n772 gnd 0.011251f
C3297 vdd.n773 gnd 0.011251f
C3298 vdd.n774 gnd 0.011251f
C3299 vdd.n775 gnd 0.011251f
C3300 vdd.n776 gnd 0.011251f
C3301 vdd.n777 gnd 0.011251f
C3302 vdd.n778 gnd 0.011251f
C3303 vdd.n779 gnd 0.011251f
C3304 vdd.n780 gnd 0.011251f
C3305 vdd.n781 gnd 0.011251f
C3306 vdd.n782 gnd 0.011251f
C3307 vdd.n783 gnd 0.007201f
C3308 vdd.n785 gnd 0.007651f
C3309 vdd.n786 gnd 0.007651f
C3310 vdd.n787 gnd 0.007651f
C3311 vdd.n788 gnd 0.007651f
C3312 vdd.n789 gnd 0.007651f
C3313 vdd.n790 gnd 0.007651f
C3314 vdd.n792 gnd 0.007651f
C3315 vdd.n793 gnd 0.007651f
C3316 vdd.n795 gnd 0.007651f
C3317 vdd.n796 gnd 0.005569f
C3318 vdd.n798 gnd 0.007651f
C3319 vdd.t64 gnd 0.309167f
C3320 vdd.t63 gnd 0.316471f
C3321 vdd.t62 gnd 0.201836f
C3322 vdd.n799 gnd 0.109081f
C3323 vdd.n800 gnd 0.061874f
C3324 vdd.n801 gnd 0.010934f
C3325 vdd.n802 gnd 0.017881f
C3326 vdd.n804 gnd 0.007651f
C3327 vdd.n805 gnd 0.781873f
C3328 vdd.n806 gnd 0.01695f
C3329 vdd.n807 gnd 0.01695f
C3330 vdd.n808 gnd 0.007651f
C3331 vdd.n809 gnd 0.018154f
C3332 vdd.n810 gnd 0.007651f
C3333 vdd.n811 gnd 0.007651f
C3334 vdd.n812 gnd 0.007651f
C3335 vdd.n813 gnd 0.007651f
C3336 vdd.n814 gnd 0.007651f
C3337 vdd.n816 gnd 0.007651f
C3338 vdd.n817 gnd 0.007651f
C3339 vdd.n819 gnd 0.007651f
C3340 vdd.n820 gnd 0.007651f
C3341 vdd.n822 gnd 0.007651f
C3342 vdd.n823 gnd 0.007651f
C3343 vdd.n825 gnd 0.007651f
C3344 vdd.n826 gnd 0.007651f
C3345 vdd.n828 gnd 0.007651f
C3346 vdd.n829 gnd 0.007651f
C3347 vdd.n831 gnd 0.007651f
C3348 vdd.t57 gnd 0.309167f
C3349 vdd.t56 gnd 0.316471f
C3350 vdd.t54 gnd 0.201836f
C3351 vdd.n832 gnd 0.109081f
C3352 vdd.n833 gnd 0.061874f
C3353 vdd.n834 gnd 0.007651f
C3354 vdd.n836 gnd 0.007651f
C3355 vdd.n837 gnd 0.007651f
C3356 vdd.t55 gnd 0.390936f
C3357 vdd.n838 gnd 0.007651f
C3358 vdd.n839 gnd 0.007651f
C3359 vdd.n840 gnd 0.007651f
C3360 vdd.n841 gnd 0.007651f
C3361 vdd.n842 gnd 0.007651f
C3362 vdd.n843 gnd 0.781873f
C3363 vdd.n844 gnd 0.007651f
C3364 vdd.n845 gnd 0.007651f
C3365 vdd.n846 gnd 0.684139f
C3366 vdd.n847 gnd 0.007651f
C3367 vdd.n848 gnd 0.007651f
C3368 vdd.n849 gnd 0.006751f
C3369 vdd.n850 gnd 0.007651f
C3370 vdd.n851 gnd 0.689888f
C3371 vdd.n852 gnd 0.007651f
C3372 vdd.n853 gnd 0.007651f
C3373 vdd.n854 gnd 0.007651f
C3374 vdd.n855 gnd 0.007651f
C3375 vdd.n856 gnd 0.007651f
C3376 vdd.n857 gnd 0.781873f
C3377 vdd.n858 gnd 0.007651f
C3378 vdd.n859 gnd 0.007651f
C3379 vdd.t27 gnd 0.350693f
C3380 vdd.t96 gnd 0.091985f
C3381 vdd.n860 gnd 0.007651f
C3382 vdd.n861 gnd 0.007651f
C3383 vdd.n862 gnd 0.007651f
C3384 vdd.t121 gnd 0.390936f
C3385 vdd.n863 gnd 0.007651f
C3386 vdd.n864 gnd 0.007651f
C3387 vdd.n865 gnd 0.007651f
C3388 vdd.n866 gnd 0.007651f
C3389 vdd.n867 gnd 0.007651f
C3390 vdd.t99 gnd 0.390936f
C3391 vdd.n868 gnd 0.007651f
C3392 vdd.n869 gnd 0.007651f
C3393 vdd.n870 gnd 0.649644f
C3394 vdd.n871 gnd 0.007651f
C3395 vdd.n872 gnd 0.007651f
C3396 vdd.n873 gnd 0.007651f
C3397 vdd.n874 gnd 0.477172f
C3398 vdd.n875 gnd 0.007651f
C3399 vdd.n876 gnd 0.007651f
C3400 vdd.t113 gnd 0.390936f
C3401 vdd.n877 gnd 0.007651f
C3402 vdd.n878 gnd 0.007651f
C3403 vdd.n879 gnd 0.007651f
C3404 vdd.n880 gnd 0.649644f
C3405 vdd.n881 gnd 0.007651f
C3406 vdd.n882 gnd 0.007651f
C3407 vdd.t130 gnd 0.333446f
C3408 vdd.t122 gnd 0.3047f
C3409 vdd.n883 gnd 0.007651f
C3410 vdd.n884 gnd 0.007651f
C3411 vdd.n885 gnd 0.007651f
C3412 vdd.t1 gnd 0.390936f
C3413 vdd.n886 gnd 0.007651f
C3414 vdd.n887 gnd 0.007651f
C3415 vdd.t10 gnd 0.390936f
C3416 vdd.n888 gnd 0.007651f
C3417 vdd.n889 gnd 0.007651f
C3418 vdd.n890 gnd 0.007651f
C3419 vdd.t124 gnd 0.287453f
C3420 vdd.n891 gnd 0.007651f
C3421 vdd.n892 gnd 0.007651f
C3422 vdd.n893 gnd 0.666891f
C3423 vdd.n894 gnd 0.007651f
C3424 vdd.n895 gnd 0.007651f
C3425 vdd.n896 gnd 0.007651f
C3426 vdd.n897 gnd 0.781873f
C3427 vdd.n898 gnd 0.007651f
C3428 vdd.n899 gnd 0.007651f
C3429 vdd.t89 gnd 0.350693f
C3430 vdd.n900 gnd 0.494419f
C3431 vdd.n901 gnd 0.007651f
C3432 vdd.n902 gnd 0.007651f
C3433 vdd.n903 gnd 0.007651f
C3434 vdd.t97 gnd 0.390936f
C3435 vdd.n904 gnd 0.007651f
C3436 vdd.n905 gnd 0.007651f
C3437 vdd.n906 gnd 0.007651f
C3438 vdd.n907 gnd 0.007651f
C3439 vdd.n908 gnd 0.007651f
C3440 vdd.t119 gnd 0.781873f
C3441 vdd.n909 gnd 0.007651f
C3442 vdd.n910 gnd 0.007651f
C3443 vdd.t59 gnd 0.390936f
C3444 vdd.n911 gnd 0.007651f
C3445 vdd.n912 gnd 0.018154f
C3446 vdd.n913 gnd 0.018154f
C3447 vdd.t5 gnd 0.73588f
C3448 vdd.n914 gnd 0.01695f
C3449 vdd.n915 gnd 0.01695f
C3450 vdd.n916 gnd 0.018154f
C3451 vdd.n917 gnd 0.007651f
C3452 vdd.n918 gnd 0.007651f
C3453 vdd.t94 gnd 0.73588f
C3454 vdd.n936 gnd 0.018154f
C3455 vdd.n954 gnd 0.01695f
C3456 vdd.n955 gnd 0.007651f
C3457 vdd.n956 gnd 0.01695f
C3458 vdd.t77 gnd 0.309167f
C3459 vdd.t76 gnd 0.316471f
C3460 vdd.t75 gnd 0.201836f
C3461 vdd.n957 gnd 0.109081f
C3462 vdd.n958 gnd 0.061874f
C3463 vdd.n959 gnd 0.017881f
C3464 vdd.n960 gnd 0.007651f
C3465 vdd.t109 gnd 0.781873f
C3466 vdd.n961 gnd 0.01695f
C3467 vdd.n962 gnd 0.007651f
C3468 vdd.n963 gnd 0.018154f
C3469 vdd.n964 gnd 0.007651f
C3470 vdd.t53 gnd 0.309167f
C3471 vdd.t52 gnd 0.316471f
C3472 vdd.t50 gnd 0.201836f
C3473 vdd.n965 gnd 0.109081f
C3474 vdd.n966 gnd 0.061874f
C3475 vdd.n967 gnd 0.010934f
C3476 vdd.n968 gnd 0.007651f
C3477 vdd.n969 gnd 0.007651f
C3478 vdd.t51 gnd 0.390936f
C3479 vdd.n970 gnd 0.007651f
C3480 vdd.n971 gnd 0.007651f
C3481 vdd.n972 gnd 0.007651f
C3482 vdd.n973 gnd 0.007651f
C3483 vdd.n974 gnd 0.007651f
C3484 vdd.n975 gnd 0.007651f
C3485 vdd.n976 gnd 0.781873f
C3486 vdd.n977 gnd 0.007651f
C3487 vdd.n978 gnd 0.007651f
C3488 vdd.t127 gnd 0.390936f
C3489 vdd.n979 gnd 0.007651f
C3490 vdd.n980 gnd 0.007651f
C3491 vdd.n981 gnd 0.007651f
C3492 vdd.n982 gnd 0.007651f
C3493 vdd.n983 gnd 0.494419f
C3494 vdd.n984 gnd 0.007651f
C3495 vdd.n985 gnd 0.007651f
C3496 vdd.n986 gnd 0.007651f
C3497 vdd.n987 gnd 0.007651f
C3498 vdd.n988 gnd 0.007651f
C3499 vdd.n989 gnd 0.666891f
C3500 vdd.n990 gnd 0.007651f
C3501 vdd.n991 gnd 0.007651f
C3502 vdd.t3 gnd 0.350693f
C3503 vdd.t112 gnd 0.287453f
C3504 vdd.n992 gnd 0.007651f
C3505 vdd.n993 gnd 0.007651f
C3506 vdd.n994 gnd 0.007651f
C3507 vdd.t91 gnd 0.390936f
C3508 vdd.n995 gnd 0.007651f
C3509 vdd.n996 gnd 0.007651f
C3510 vdd.t125 gnd 0.390936f
C3511 vdd.n997 gnd 0.007651f
C3512 vdd.n998 gnd 0.007651f
C3513 vdd.n999 gnd 0.007651f
C3514 vdd.t92 gnd 0.3047f
C3515 vdd.n1000 gnd 0.007651f
C3516 vdd.n1001 gnd 0.007651f
C3517 vdd.n1002 gnd 0.649644f
C3518 vdd.n1003 gnd 0.007651f
C3519 vdd.n1004 gnd 0.007651f
C3520 vdd.n1005 gnd 0.007651f
C3521 vdd.t294 gnd 0.390936f
C3522 vdd.n1006 gnd 0.007651f
C3523 vdd.n1007 gnd 0.007651f
C3524 vdd.t0 gnd 0.333446f
C3525 vdd.n1008 gnd 0.477172f
C3526 vdd.n1009 gnd 0.007651f
C3527 vdd.n1010 gnd 0.007651f
C3528 vdd.n1011 gnd 0.007651f
C3529 vdd.n1012 gnd 0.649644f
C3530 vdd.n1013 gnd 0.007651f
C3531 vdd.n1014 gnd 0.007651f
C3532 vdd.t129 gnd 0.390936f
C3533 vdd.n1015 gnd 0.007651f
C3534 vdd.n1016 gnd 0.007651f
C3535 vdd.n1017 gnd 0.007651f
C3536 vdd.n1018 gnd 0.781873f
C3537 vdd.n1019 gnd 0.007651f
C3538 vdd.n1020 gnd 0.007651f
C3539 vdd.t103 gnd 0.390936f
C3540 vdd.n1021 gnd 0.007651f
C3541 vdd.n1022 gnd 0.007651f
C3542 vdd.n1023 gnd 0.007651f
C3543 vdd.t111 gnd 0.091985f
C3544 vdd.n1024 gnd 0.007651f
C3545 vdd.n1025 gnd 0.007651f
C3546 vdd.n1026 gnd 0.007651f
C3547 vdd.t70 gnd 0.316471f
C3548 vdd.t68 gnd 0.201836f
C3549 vdd.t71 gnd 0.316471f
C3550 vdd.n1027 gnd 0.177869f
C3551 vdd.n1028 gnd 0.007651f
C3552 vdd.n1029 gnd 0.007651f
C3553 vdd.n1030 gnd 0.781873f
C3554 vdd.n1031 gnd 0.007651f
C3555 vdd.n1032 gnd 0.007651f
C3556 vdd.t69 gnd 0.350693f
C3557 vdd.n1033 gnd 0.689888f
C3558 vdd.n1034 gnd 0.007651f
C3559 vdd.n1035 gnd 0.007651f
C3560 vdd.n1036 gnd 0.007651f
C3561 vdd.n1037 gnd 0.684139f
C3562 vdd.n1038 gnd 0.007651f
C3563 vdd.n1039 gnd 0.007651f
C3564 vdd.n1040 gnd 0.007651f
C3565 vdd.n1041 gnd 0.007651f
C3566 vdd.n1042 gnd 0.007651f
C3567 vdd.n1043 gnd 0.781873f
C3568 vdd.n1044 gnd 0.007651f
C3569 vdd.n1045 gnd 0.007651f
C3570 vdd.t12 gnd 0.390936f
C3571 vdd.n1046 gnd 0.007651f
C3572 vdd.n1047 gnd 0.018154f
C3573 vdd.n1048 gnd 0.018154f
C3574 vdd.n1049 gnd 7.92221f
C3575 vdd.n1050 gnd 0.01695f
C3576 vdd.n1051 gnd 0.01695f
C3577 vdd.n1052 gnd 0.018154f
C3578 vdd.n1053 gnd 0.007651f
C3579 vdd.n1054 gnd 0.007651f
C3580 vdd.n1055 gnd 0.007651f
C3581 vdd.n1056 gnd 0.007651f
C3582 vdd.n1057 gnd 0.007651f
C3583 vdd.n1058 gnd 0.007651f
C3584 vdd.n1059 gnd 0.007651f
C3585 vdd.n1060 gnd 0.007651f
C3586 vdd.n1062 gnd 0.007651f
C3587 vdd.n1063 gnd 0.007651f
C3588 vdd.n1064 gnd 0.007201f
C3589 vdd.n1067 gnd 0.027801f
C3590 vdd.n1068 gnd 0.009056f
C3591 vdd.n1069 gnd 0.011251f
C3592 vdd.n1071 gnd 0.011251f
C3593 vdd.n1072 gnd 0.007516f
C3594 vdd.t23 gnd 0.574906f
C3595 vdd.n1073 gnd 8.31315f
C3596 vdd.n1074 gnd 0.011251f
C3597 vdd.n1075 gnd 0.027801f
C3598 vdd.n1076 gnd 0.009056f
C3599 vdd.n1077 gnd 0.011251f
C3600 vdd.n1078 gnd 0.009056f
C3601 vdd.n1079 gnd 0.011251f
C3602 vdd.n1080 gnd 1.14981f
C3603 vdd.n1081 gnd 0.011251f
C3604 vdd.n1082 gnd 0.009056f
C3605 vdd.n1083 gnd 0.009056f
C3606 vdd.n1084 gnd 0.011251f
C3607 vdd.n1085 gnd 0.009056f
C3608 vdd.n1086 gnd 0.011251f
C3609 vdd.t141 gnd 0.574906f
C3610 vdd.n1087 gnd 0.011251f
C3611 vdd.n1088 gnd 0.009056f
C3612 vdd.n1089 gnd 0.011251f
C3613 vdd.n1090 gnd 0.009056f
C3614 vdd.n1091 gnd 0.011251f
C3615 vdd.t269 gnd 0.574906f
C3616 vdd.n1092 gnd 0.011251f
C3617 vdd.n1093 gnd 0.009056f
C3618 vdd.n1094 gnd 0.011251f
C3619 vdd.n1095 gnd 0.009056f
C3620 vdd.n1096 gnd 0.011251f
C3621 vdd.n1097 gnd 0.925599f
C3622 vdd.n1098 gnd 0.954345f
C3623 vdd.t133 gnd 0.574906f
C3624 vdd.n1099 gnd 0.011251f
C3625 vdd.n1100 gnd 0.009056f
C3626 vdd.n1101 gnd 0.011251f
C3627 vdd.n1102 gnd 0.009056f
C3628 vdd.n1103 gnd 0.011251f
C3629 vdd.n1104 gnd 0.730131f
C3630 vdd.n1105 gnd 0.011251f
C3631 vdd.n1106 gnd 0.009056f
C3632 vdd.n1107 gnd 0.011251f
C3633 vdd.n1108 gnd 0.009056f
C3634 vdd.n1109 gnd 0.011251f
C3635 vdd.t143 gnd 0.574906f
C3636 vdd.t183 gnd 0.574906f
C3637 vdd.n1110 gnd 0.011251f
C3638 vdd.n1111 gnd 0.009056f
C3639 vdd.n1112 gnd 0.011251f
C3640 vdd.n1113 gnd 0.009056f
C3641 vdd.n1114 gnd 0.011251f
C3642 vdd.t206 gnd 0.574906f
C3643 vdd.n1115 gnd 0.011251f
C3644 vdd.n1116 gnd 0.009056f
C3645 vdd.n1117 gnd 0.011251f
C3646 vdd.n1118 gnd 0.009056f
C3647 vdd.n1119 gnd 0.011251f
C3648 vdd.t247 gnd 0.574906f
C3649 vdd.n1120 gnd 0.810618f
C3650 vdd.n1121 gnd 0.011251f
C3651 vdd.n1122 gnd 0.009056f
C3652 vdd.n1123 gnd 0.011251f
C3653 vdd.n1124 gnd 0.009056f
C3654 vdd.n1125 gnd 0.011251f
C3655 vdd.n1126 gnd 0.902603f
C3656 vdd.n1127 gnd 0.011251f
C3657 vdd.n1128 gnd 0.009056f
C3658 vdd.n1129 gnd 0.011251f
C3659 vdd.n1130 gnd 0.009056f
C3660 vdd.n1131 gnd 0.011251f
C3661 vdd.n1132 gnd 0.707135f
C3662 vdd.t149 gnd 0.574906f
C3663 vdd.n1133 gnd 0.011251f
C3664 vdd.n1134 gnd 0.009056f
C3665 vdd.n1135 gnd 0.011251f
C3666 vdd.n1136 gnd 0.009056f
C3667 vdd.n1137 gnd 0.011251f
C3668 vdd.t160 gnd 0.574906f
C3669 vdd.n1138 gnd 0.011251f
C3670 vdd.n1139 gnd 0.009056f
C3671 vdd.n1140 gnd 0.011251f
C3672 vdd.n1141 gnd 0.009056f
C3673 vdd.n1142 gnd 0.011251f
C3674 vdd.t178 gnd 0.574906f
C3675 vdd.n1143 gnd 0.638146f
C3676 vdd.n1144 gnd 0.011251f
C3677 vdd.n1145 gnd 0.009056f
C3678 vdd.n1146 gnd 0.011251f
C3679 vdd.n1147 gnd 0.009056f
C3680 vdd.n1148 gnd 0.011251f
C3681 vdd.t224 gnd 0.574906f
C3682 vdd.n1149 gnd 0.011251f
C3683 vdd.n1150 gnd 0.009056f
C3684 vdd.n1151 gnd 0.011251f
C3685 vdd.n1152 gnd 0.009056f
C3686 vdd.n1153 gnd 0.011251f
C3687 vdd.n1154 gnd 0.879607f
C3688 vdd.n1155 gnd 0.954345f
C3689 vdd.t226 gnd 0.574906f
C3690 vdd.n1156 gnd 0.011251f
C3691 vdd.n1157 gnd 0.009056f
C3692 vdd.n1158 gnd 0.011251f
C3693 vdd.n1159 gnd 0.009056f
C3694 vdd.n1160 gnd 0.011251f
C3695 vdd.n1161 gnd 0.684139f
C3696 vdd.n1162 gnd 0.011251f
C3697 vdd.n1163 gnd 0.009056f
C3698 vdd.n1164 gnd 0.011251f
C3699 vdd.n1165 gnd 0.009056f
C3700 vdd.n1166 gnd 0.011251f
C3701 vdd.t176 gnd 0.574906f
C3702 vdd.t174 gnd 0.574906f
C3703 vdd.n1167 gnd 0.011251f
C3704 vdd.n1168 gnd 0.009056f
C3705 vdd.n1169 gnd 0.011251f
C3706 vdd.n1170 gnd 0.009056f
C3707 vdd.n1171 gnd 0.011251f
C3708 vdd.t139 gnd 0.574906f
C3709 vdd.n1172 gnd 0.011251f
C3710 vdd.n1173 gnd 0.009056f
C3711 vdd.n1174 gnd 0.011251f
C3712 vdd.n1175 gnd 0.009056f
C3713 vdd.n1176 gnd 0.011251f
C3714 vdd.t145 gnd 0.574906f
C3715 vdd.n1177 gnd 0.85661f
C3716 vdd.n1178 gnd 0.011251f
C3717 vdd.n1179 gnd 0.009056f
C3718 vdd.n1180 gnd 0.011251f
C3719 vdd.n1181 gnd 0.009056f
C3720 vdd.n1182 gnd 0.011251f
C3721 vdd.n1183 gnd 1.14981f
C3722 vdd.n1184 gnd 0.011251f
C3723 vdd.n1185 gnd 0.009056f
C3724 vdd.n1186 gnd 0.027217f
C3725 vdd.n1187 gnd 0.007516f
C3726 vdd.n1188 gnd 0.027217f
C3727 vdd.t31 gnd 0.574906f
C3728 vdd.n1189 gnd 0.027217f
C3729 vdd.n1190 gnd 0.007516f
C3730 vdd.n1191 gnd 0.011251f
C3731 vdd.n1192 gnd 0.009056f
C3732 vdd.n1193 gnd 0.011251f
C3733 vdd.n1224 gnd 0.027801f
C3734 vdd.n1225 gnd 1.69597f
C3735 vdd.n1226 gnd 0.011251f
C3736 vdd.n1227 gnd 0.009056f
C3737 vdd.n1228 gnd 0.011251f
C3738 vdd.n1229 gnd 0.011251f
C3739 vdd.n1230 gnd 0.011251f
C3740 vdd.n1231 gnd 0.011251f
C3741 vdd.n1232 gnd 0.011251f
C3742 vdd.n1233 gnd 0.009056f
C3743 vdd.n1234 gnd 0.011251f
C3744 vdd.n1235 gnd 0.011251f
C3745 vdd.n1236 gnd 0.011251f
C3746 vdd.n1237 gnd 0.011251f
C3747 vdd.n1238 gnd 0.011251f
C3748 vdd.n1239 gnd 0.009056f
C3749 vdd.n1240 gnd 0.011251f
C3750 vdd.n1241 gnd 0.011251f
C3751 vdd.n1242 gnd 0.011251f
C3752 vdd.n1243 gnd 0.011251f
C3753 vdd.n1244 gnd 0.011251f
C3754 vdd.n1245 gnd 0.009056f
C3755 vdd.n1246 gnd 0.011251f
C3756 vdd.n1247 gnd 0.011251f
C3757 vdd.n1248 gnd 0.011251f
C3758 vdd.n1249 gnd 0.011251f
C3759 vdd.n1250 gnd 0.011251f
C3760 vdd.t45 gnd 0.138418f
C3761 vdd.t46 gnd 0.147931f
C3762 vdd.t44 gnd 0.180773f
C3763 vdd.n1251 gnd 0.231725f
C3764 vdd.n1252 gnd 0.195597f
C3765 vdd.n1253 gnd 0.019379f
C3766 vdd.n1254 gnd 0.011251f
C3767 vdd.n1255 gnd 0.011251f
C3768 vdd.n1256 gnd 0.011251f
C3769 vdd.n1257 gnd 0.011251f
C3770 vdd.n1258 gnd 0.011251f
C3771 vdd.n1259 gnd 0.009056f
C3772 vdd.n1260 gnd 0.011251f
C3773 vdd.n1261 gnd 0.011251f
C3774 vdd.n1262 gnd 0.011251f
C3775 vdd.n1263 gnd 0.011251f
C3776 vdd.n1264 gnd 0.011251f
C3777 vdd.n1265 gnd 0.009056f
C3778 vdd.n1266 gnd 0.011251f
C3779 vdd.n1267 gnd 0.011251f
C3780 vdd.n1268 gnd 0.011251f
C3781 vdd.n1269 gnd 0.011251f
C3782 vdd.n1270 gnd 0.011251f
C3783 vdd.n1271 gnd 0.009056f
C3784 vdd.n1272 gnd 0.011251f
C3785 vdd.n1273 gnd 0.011251f
C3786 vdd.n1274 gnd 0.011251f
C3787 vdd.n1275 gnd 0.011251f
C3788 vdd.n1276 gnd 0.011251f
C3789 vdd.n1277 gnd 0.009056f
C3790 vdd.n1278 gnd 0.011251f
C3791 vdd.n1279 gnd 0.011251f
C3792 vdd.n1280 gnd 0.011251f
C3793 vdd.n1281 gnd 0.011251f
C3794 vdd.n1282 gnd 0.011251f
C3795 vdd.n1283 gnd 0.009056f
C3796 vdd.n1284 gnd 0.011251f
C3797 vdd.n1285 gnd 0.011251f
C3798 vdd.n1286 gnd 0.011251f
C3799 vdd.n1287 gnd 0.011251f
C3800 vdd.n1288 gnd 0.009056f
C3801 vdd.n1289 gnd 0.011251f
C3802 vdd.n1290 gnd 0.011251f
C3803 vdd.n1291 gnd 0.011251f
C3804 vdd.n1292 gnd 0.011251f
C3805 vdd.n1293 gnd 0.011251f
C3806 vdd.n1294 gnd 0.009056f
C3807 vdd.n1295 gnd 0.011251f
C3808 vdd.n1296 gnd 0.011251f
C3809 vdd.n1297 gnd 0.011251f
C3810 vdd.n1298 gnd 0.011251f
C3811 vdd.n1299 gnd 0.011251f
C3812 vdd.n1300 gnd 0.009056f
C3813 vdd.n1301 gnd 0.011251f
C3814 vdd.n1302 gnd 0.011251f
C3815 vdd.n1303 gnd 0.011251f
C3816 vdd.n1304 gnd 0.011251f
C3817 vdd.n1305 gnd 0.011251f
C3818 vdd.n1306 gnd 0.009056f
C3819 vdd.n1307 gnd 0.011251f
C3820 vdd.n1308 gnd 0.011251f
C3821 vdd.n1309 gnd 0.011251f
C3822 vdd.n1310 gnd 0.011251f
C3823 vdd.n1311 gnd 0.011251f
C3824 vdd.n1312 gnd 0.009056f
C3825 vdd.n1313 gnd 0.011251f
C3826 vdd.n1314 gnd 0.011251f
C3827 vdd.n1315 gnd 0.011251f
C3828 vdd.n1316 gnd 0.011251f
C3829 vdd.t42 gnd 0.138418f
C3830 vdd.t43 gnd 0.147931f
C3831 vdd.t41 gnd 0.180773f
C3832 vdd.n1317 gnd 0.231725f
C3833 vdd.n1318 gnd 0.195597f
C3834 vdd.n1319 gnd 0.014852f
C3835 vdd.n1320 gnd 0.004302f
C3836 vdd.n1321 gnd 0.027801f
C3837 vdd.n1322 gnd 0.011251f
C3838 vdd.n1323 gnd 0.004754f
C3839 vdd.n1324 gnd 0.009056f
C3840 vdd.n1325 gnd 0.009056f
C3841 vdd.n1326 gnd 0.011251f
C3842 vdd.n1327 gnd 0.011251f
C3843 vdd.n1328 gnd 0.011251f
C3844 vdd.n1329 gnd 0.009056f
C3845 vdd.n1330 gnd 0.009056f
C3846 vdd.n1331 gnd 0.009056f
C3847 vdd.n1332 gnd 0.011251f
C3848 vdd.n1333 gnd 0.011251f
C3849 vdd.n1334 gnd 0.011251f
C3850 vdd.n1335 gnd 0.009056f
C3851 vdd.n1336 gnd 0.009056f
C3852 vdd.n1337 gnd 0.009056f
C3853 vdd.n1338 gnd 0.011251f
C3854 vdd.n1339 gnd 0.011251f
C3855 vdd.n1340 gnd 0.011251f
C3856 vdd.n1341 gnd 0.009056f
C3857 vdd.n1342 gnd 0.009056f
C3858 vdd.n1343 gnd 0.009056f
C3859 vdd.n1344 gnd 0.011251f
C3860 vdd.n1345 gnd 0.011251f
C3861 vdd.n1346 gnd 0.011251f
C3862 vdd.n1347 gnd 0.009056f
C3863 vdd.n1348 gnd 0.009056f
C3864 vdd.n1349 gnd 0.009056f
C3865 vdd.n1350 gnd 0.011251f
C3866 vdd.n1351 gnd 0.011251f
C3867 vdd.n1352 gnd 0.011251f
C3868 vdd.n1353 gnd 0.008965f
C3869 vdd.n1354 gnd 0.011251f
C3870 vdd.t32 gnd 0.138418f
C3871 vdd.t33 gnd 0.147931f
C3872 vdd.t30 gnd 0.180773f
C3873 vdd.n1355 gnd 0.231725f
C3874 vdd.n1356 gnd 0.195597f
C3875 vdd.n1357 gnd 0.019379f
C3876 vdd.n1358 gnd 0.006158f
C3877 vdd.n1359 gnd 0.011251f
C3878 vdd.n1360 gnd 0.011251f
C3879 vdd.n1361 gnd 0.011251f
C3880 vdd.n1362 gnd 0.009056f
C3881 vdd.n1363 gnd 0.009056f
C3882 vdd.n1364 gnd 0.009056f
C3883 vdd.n1365 gnd 0.011251f
C3884 vdd.n1366 gnd 0.011251f
C3885 vdd.n1367 gnd 0.011251f
C3886 vdd.n1368 gnd 0.009056f
C3887 vdd.n1369 gnd 0.009056f
C3888 vdd.n1370 gnd 0.009056f
C3889 vdd.n1371 gnd 0.011251f
C3890 vdd.n1372 gnd 0.011251f
C3891 vdd.n1373 gnd 0.011251f
C3892 vdd.n1374 gnd 0.009056f
C3893 vdd.n1375 gnd 0.009056f
C3894 vdd.n1376 gnd 0.009056f
C3895 vdd.n1377 gnd 0.011251f
C3896 vdd.n1378 gnd 0.011251f
C3897 vdd.n1379 gnd 0.011251f
C3898 vdd.n1380 gnd 0.009056f
C3899 vdd.n1381 gnd 0.009056f
C3900 vdd.n1382 gnd 0.009056f
C3901 vdd.n1383 gnd 0.011251f
C3902 vdd.n1384 gnd 0.011251f
C3903 vdd.n1385 gnd 0.011251f
C3904 vdd.n1386 gnd 0.009056f
C3905 vdd.n1387 gnd 0.009056f
C3906 vdd.n1388 gnd 0.007562f
C3907 vdd.n1389 gnd 0.011251f
C3908 vdd.n1390 gnd 0.011251f
C3909 vdd.n1391 gnd 0.011251f
C3910 vdd.n1392 gnd 0.007562f
C3911 vdd.n1393 gnd 0.009056f
C3912 vdd.n1394 gnd 0.009056f
C3913 vdd.n1395 gnd 0.011251f
C3914 vdd.n1396 gnd 0.011251f
C3915 vdd.n1397 gnd 0.011251f
C3916 vdd.n1398 gnd 0.009056f
C3917 vdd.n1399 gnd 0.009056f
C3918 vdd.n1400 gnd 0.009056f
C3919 vdd.n1401 gnd 0.011251f
C3920 vdd.n1402 gnd 0.011251f
C3921 vdd.n1403 gnd 0.011251f
C3922 vdd.n1404 gnd 0.009056f
C3923 vdd.n1405 gnd 0.009056f
C3924 vdd.n1406 gnd 0.009056f
C3925 vdd.n1407 gnd 0.011251f
C3926 vdd.n1408 gnd 0.011251f
C3927 vdd.n1409 gnd 0.011251f
C3928 vdd.n1410 gnd 0.009056f
C3929 vdd.n1411 gnd 0.009056f
C3930 vdd.n1412 gnd 0.009056f
C3931 vdd.n1413 gnd 0.011251f
C3932 vdd.n1414 gnd 0.011251f
C3933 vdd.n1415 gnd 0.011251f
C3934 vdd.n1416 gnd 0.009056f
C3935 vdd.n1417 gnd 0.011251f
C3936 vdd.n1418 gnd 2.72506f
C3937 vdd.n1420 gnd 0.027801f
C3938 vdd.n1421 gnd 0.007516f
C3939 vdd.n1422 gnd 0.027801f
C3940 vdd.n1423 gnd 0.027217f
C3941 vdd.n1424 gnd 0.011251f
C3942 vdd.n1425 gnd 0.009056f
C3943 vdd.n1426 gnd 0.011251f
C3944 vdd.n1427 gnd 0.580655f
C3945 vdd.n1428 gnd 0.011251f
C3946 vdd.n1429 gnd 0.009056f
C3947 vdd.n1430 gnd 0.011251f
C3948 vdd.n1431 gnd 0.011251f
C3949 vdd.n1432 gnd 0.011251f
C3950 vdd.n1433 gnd 0.009056f
C3951 vdd.n1434 gnd 0.011251f
C3952 vdd.n1435 gnd 1.05208f
C3953 vdd.n1436 gnd 1.14981f
C3954 vdd.n1437 gnd 0.011251f
C3955 vdd.n1438 gnd 0.009056f
C3956 vdd.n1439 gnd 0.011251f
C3957 vdd.n1440 gnd 0.011251f
C3958 vdd.n1441 gnd 0.011251f
C3959 vdd.n1442 gnd 0.009056f
C3960 vdd.n1443 gnd 0.011251f
C3961 vdd.n1444 gnd 0.67264f
C3962 vdd.n1445 gnd 0.011251f
C3963 vdd.n1446 gnd 0.009056f
C3964 vdd.n1447 gnd 0.011251f
C3965 vdd.n1448 gnd 0.011251f
C3966 vdd.n1449 gnd 0.011251f
C3967 vdd.n1450 gnd 0.009056f
C3968 vdd.n1451 gnd 0.011251f
C3969 vdd.n1452 gnd 0.661142f
C3970 vdd.n1453 gnd 0.868109f
C3971 vdd.n1454 gnd 0.011251f
C3972 vdd.n1455 gnd 0.009056f
C3973 vdd.n1456 gnd 0.011251f
C3974 vdd.n1457 gnd 0.011251f
C3975 vdd.n1458 gnd 0.011251f
C3976 vdd.n1459 gnd 0.009056f
C3977 vdd.n1460 gnd 0.011251f
C3978 vdd.n1461 gnd 0.954345f
C3979 vdd.n1462 gnd 0.011251f
C3980 vdd.n1463 gnd 0.009056f
C3981 vdd.n1464 gnd 0.011251f
C3982 vdd.n1465 gnd 0.011251f
C3983 vdd.n1466 gnd 0.011251f
C3984 vdd.n1467 gnd 0.009056f
C3985 vdd.n1468 gnd 0.011251f
C3986 vdd.t153 gnd 0.574906f
C3987 vdd.n1469 gnd 0.845112f
C3988 vdd.n1470 gnd 0.011251f
C3989 vdd.n1471 gnd 0.009056f
C3990 vdd.n1472 gnd 0.011251f
C3991 vdd.n1473 gnd 0.011251f
C3992 vdd.n1474 gnd 0.011251f
C3993 vdd.n1475 gnd 0.009056f
C3994 vdd.n1476 gnd 0.011251f
C3995 vdd.n1477 gnd 0.649644f
C3996 vdd.n1478 gnd 0.011251f
C3997 vdd.n1479 gnd 0.009056f
C3998 vdd.n1480 gnd 0.011251f
C3999 vdd.n1481 gnd 0.011251f
C4000 vdd.n1482 gnd 0.011251f
C4001 vdd.n1483 gnd 0.009056f
C4002 vdd.n1484 gnd 0.011251f
C4003 vdd.n1485 gnd 0.833614f
C4004 vdd.n1486 gnd 0.695637f
C4005 vdd.n1487 gnd 0.011251f
C4006 vdd.n1488 gnd 0.009056f
C4007 vdd.n1489 gnd 0.011251f
C4008 vdd.n1490 gnd 0.011251f
C4009 vdd.n1491 gnd 0.011251f
C4010 vdd.n1492 gnd 0.009056f
C4011 vdd.n1493 gnd 0.011251f
C4012 vdd.n1494 gnd 0.891105f
C4013 vdd.n1495 gnd 0.011251f
C4014 vdd.n1496 gnd 0.009056f
C4015 vdd.n1497 gnd 0.011251f
C4016 vdd.n1498 gnd 0.011251f
C4017 vdd.n1499 gnd 0.011251f
C4018 vdd.n1500 gnd 0.009056f
C4019 vdd.n1501 gnd 0.011251f
C4020 vdd.t196 gnd 0.574906f
C4021 vdd.n1502 gnd 0.954345f
C4022 vdd.n1503 gnd 0.011251f
C4023 vdd.n1504 gnd 0.009056f
C4024 vdd.n1505 gnd 0.011251f
C4025 vdd.n1506 gnd 0.008647f
C4026 vdd.n1507 gnd 0.006175f
C4027 vdd.n1508 gnd 0.00573f
C4028 vdd.n1509 gnd 0.00317f
C4029 vdd.n1510 gnd 0.007278f
C4030 vdd.n1511 gnd 0.003079f
C4031 vdd.n1512 gnd 0.00326f
C4032 vdd.n1513 gnd 0.00573f
C4033 vdd.n1514 gnd 0.003079f
C4034 vdd.n1515 gnd 0.007278f
C4035 vdd.n1516 gnd 0.00326f
C4036 vdd.n1517 gnd 0.00573f
C4037 vdd.n1518 gnd 0.003079f
C4038 vdd.n1519 gnd 0.005458f
C4039 vdd.n1520 gnd 0.005474f
C4040 vdd.t142 gnd 0.015635f
C4041 vdd.n1521 gnd 0.034788f
C4042 vdd.n1522 gnd 0.181046f
C4043 vdd.n1523 gnd 0.003079f
C4044 vdd.n1524 gnd 0.00326f
C4045 vdd.n1525 gnd 0.007278f
C4046 vdd.n1526 gnd 0.007278f
C4047 vdd.n1527 gnd 0.00326f
C4048 vdd.n1528 gnd 0.003079f
C4049 vdd.n1529 gnd 0.00573f
C4050 vdd.n1530 gnd 0.00573f
C4051 vdd.n1531 gnd 0.003079f
C4052 vdd.n1532 gnd 0.00326f
C4053 vdd.n1533 gnd 0.007278f
C4054 vdd.n1534 gnd 0.007278f
C4055 vdd.n1535 gnd 0.00326f
C4056 vdd.n1536 gnd 0.003079f
C4057 vdd.n1537 gnd 0.00573f
C4058 vdd.n1538 gnd 0.00573f
C4059 vdd.n1539 gnd 0.003079f
C4060 vdd.n1540 gnd 0.00326f
C4061 vdd.n1541 gnd 0.007278f
C4062 vdd.n1542 gnd 0.007278f
C4063 vdd.n1543 gnd 0.017206f
C4064 vdd.n1544 gnd 0.00317f
C4065 vdd.n1545 gnd 0.003079f
C4066 vdd.n1546 gnd 0.01481f
C4067 vdd.n1547 gnd 0.010339f
C4068 vdd.t217 gnd 0.036223f
C4069 vdd.t276 gnd 0.036223f
C4070 vdd.n1548 gnd 0.248951f
C4071 vdd.n1549 gnd 0.195762f
C4072 vdd.t184 gnd 0.036223f
C4073 vdd.t257 gnd 0.036223f
C4074 vdd.n1550 gnd 0.248951f
C4075 vdd.n1551 gnd 0.157979f
C4076 vdd.t207 gnd 0.036223f
C4077 vdd.t234 gnd 0.036223f
C4078 vdd.n1552 gnd 0.248951f
C4079 vdd.n1553 gnd 0.157979f
C4080 vdd.t231 gnd 0.036223f
C4081 vdd.t284 gnd 0.036223f
C4082 vdd.n1554 gnd 0.248951f
C4083 vdd.n1555 gnd 0.157979f
C4084 vdd.t197 gnd 0.036223f
C4085 vdd.t155 gnd 0.036223f
C4086 vdd.n1556 gnd 0.248951f
C4087 vdd.n1557 gnd 0.157979f
C4088 vdd.t220 gnd 0.036223f
C4089 vdd.t161 gnd 0.036223f
C4090 vdd.n1558 gnd 0.248951f
C4091 vdd.n1559 gnd 0.157979f
C4092 vdd.t272 gnd 0.036223f
C4093 vdd.t289 gnd 0.036223f
C4094 vdd.n1560 gnd 0.248951f
C4095 vdd.n1561 gnd 0.157979f
C4096 vdd.t246 gnd 0.036223f
C4097 vdd.t165 gnd 0.036223f
C4098 vdd.n1562 gnd 0.248951f
C4099 vdd.n1563 gnd 0.157979f
C4100 vdd.t232 gnd 0.036223f
C4101 vdd.t177 gnd 0.036223f
C4102 vdd.n1564 gnd 0.248951f
C4103 vdd.n1565 gnd 0.157979f
C4104 vdd.n1566 gnd 0.006175f
C4105 vdd.n1567 gnd 0.00573f
C4106 vdd.n1568 gnd 0.00317f
C4107 vdd.n1569 gnd 0.007278f
C4108 vdd.n1570 gnd 0.003079f
C4109 vdd.n1571 gnd 0.00326f
C4110 vdd.n1572 gnd 0.00573f
C4111 vdd.n1573 gnd 0.003079f
C4112 vdd.n1574 gnd 0.007278f
C4113 vdd.n1575 gnd 0.00326f
C4114 vdd.n1576 gnd 0.00573f
C4115 vdd.n1577 gnd 0.003079f
C4116 vdd.n1578 gnd 0.005458f
C4117 vdd.n1579 gnd 0.005474f
C4118 vdd.t201 gnd 0.015635f
C4119 vdd.n1580 gnd 0.034788f
C4120 vdd.n1581 gnd 0.181046f
C4121 vdd.n1582 gnd 0.003079f
C4122 vdd.n1583 gnd 0.00326f
C4123 vdd.n1584 gnd 0.007278f
C4124 vdd.n1585 gnd 0.007278f
C4125 vdd.n1586 gnd 0.00326f
C4126 vdd.n1587 gnd 0.003079f
C4127 vdd.n1588 gnd 0.00573f
C4128 vdd.n1589 gnd 0.00573f
C4129 vdd.n1590 gnd 0.003079f
C4130 vdd.n1591 gnd 0.00326f
C4131 vdd.n1592 gnd 0.007278f
C4132 vdd.n1593 gnd 0.007278f
C4133 vdd.n1594 gnd 0.00326f
C4134 vdd.n1595 gnd 0.003079f
C4135 vdd.n1596 gnd 0.00573f
C4136 vdd.n1597 gnd 0.00573f
C4137 vdd.n1598 gnd 0.003079f
C4138 vdd.n1599 gnd 0.00326f
C4139 vdd.n1600 gnd 0.007278f
C4140 vdd.n1601 gnd 0.007278f
C4141 vdd.n1602 gnd 0.017206f
C4142 vdd.n1603 gnd 0.00317f
C4143 vdd.n1604 gnd 0.003079f
C4144 vdd.n1605 gnd 0.01481f
C4145 vdd.n1606 gnd 0.010015f
C4146 vdd.n1607 gnd 0.117537f
C4147 vdd.n1608 gnd 0.006175f
C4148 vdd.n1609 gnd 0.00573f
C4149 vdd.n1610 gnd 0.00317f
C4150 vdd.n1611 gnd 0.007278f
C4151 vdd.n1612 gnd 0.003079f
C4152 vdd.n1613 gnd 0.00326f
C4153 vdd.n1614 gnd 0.00573f
C4154 vdd.n1615 gnd 0.003079f
C4155 vdd.n1616 gnd 0.007278f
C4156 vdd.n1617 gnd 0.00326f
C4157 vdd.n1618 gnd 0.00573f
C4158 vdd.n1619 gnd 0.003079f
C4159 vdd.n1620 gnd 0.005458f
C4160 vdd.n1621 gnd 0.005474f
C4161 vdd.t267 gnd 0.015635f
C4162 vdd.n1622 gnd 0.034788f
C4163 vdd.n1623 gnd 0.181046f
C4164 vdd.n1624 gnd 0.003079f
C4165 vdd.n1625 gnd 0.00326f
C4166 vdd.n1626 gnd 0.007278f
C4167 vdd.n1627 gnd 0.007278f
C4168 vdd.n1628 gnd 0.00326f
C4169 vdd.n1629 gnd 0.003079f
C4170 vdd.n1630 gnd 0.00573f
C4171 vdd.n1631 gnd 0.00573f
C4172 vdd.n1632 gnd 0.003079f
C4173 vdd.n1633 gnd 0.00326f
C4174 vdd.n1634 gnd 0.007278f
C4175 vdd.n1635 gnd 0.007278f
C4176 vdd.n1636 gnd 0.00326f
C4177 vdd.n1637 gnd 0.003079f
C4178 vdd.n1638 gnd 0.00573f
C4179 vdd.n1639 gnd 0.00573f
C4180 vdd.n1640 gnd 0.003079f
C4181 vdd.n1641 gnd 0.00326f
C4182 vdd.n1642 gnd 0.007278f
C4183 vdd.n1643 gnd 0.007278f
C4184 vdd.n1644 gnd 0.017206f
C4185 vdd.n1645 gnd 0.00317f
C4186 vdd.n1646 gnd 0.003079f
C4187 vdd.n1647 gnd 0.01481f
C4188 vdd.n1648 gnd 0.010339f
C4189 vdd.t134 gnd 0.036223f
C4190 vdd.t270 gnd 0.036223f
C4191 vdd.n1649 gnd 0.248951f
C4192 vdd.n1650 gnd 0.195762f
C4193 vdd.t264 gnd 0.036223f
C4194 vdd.t250 gnd 0.036223f
C4195 vdd.n1651 gnd 0.248951f
C4196 vdd.n1652 gnd 0.157979f
C4197 vdd.t209 gnd 0.036223f
C4198 vdd.t144 gnd 0.036223f
C4199 vdd.n1653 gnd 0.248951f
C4200 vdd.n1654 gnd 0.157979f
C4201 vdd.t279 gnd 0.036223f
C4202 vdd.t248 gnd 0.036223f
C4203 vdd.n1655 gnd 0.248951f
C4204 vdd.n1656 gnd 0.157979f
C4205 vdd.t242 gnd 0.036223f
C4206 vdd.t150 gnd 0.036223f
C4207 vdd.n1657 gnd 0.248951f
C4208 vdd.n1658 gnd 0.157979f
C4209 vdd.t179 gnd 0.036223f
C4210 vdd.t243 gnd 0.036223f
C4211 vdd.n1659 gnd 0.248951f
C4212 vdd.n1660 gnd 0.157979f
C4213 vdd.t227 gnd 0.036223f
C4214 vdd.t225 gnd 0.036223f
C4215 vdd.n1661 gnd 0.248951f
C4216 vdd.n1662 gnd 0.157979f
C4217 vdd.t175 gnd 0.036223f
C4218 vdd.t154 gnd 0.036223f
C4219 vdd.n1663 gnd 0.248951f
C4220 vdd.n1664 gnd 0.157979f
C4221 vdd.t140 gnd 0.036223f
C4222 vdd.t221 gnd 0.036223f
C4223 vdd.n1665 gnd 0.248951f
C4224 vdd.n1666 gnd 0.157979f
C4225 vdd.n1667 gnd 0.006175f
C4226 vdd.n1668 gnd 0.00573f
C4227 vdd.n1669 gnd 0.00317f
C4228 vdd.n1670 gnd 0.007278f
C4229 vdd.n1671 gnd 0.003079f
C4230 vdd.n1672 gnd 0.00326f
C4231 vdd.n1673 gnd 0.00573f
C4232 vdd.n1674 gnd 0.003079f
C4233 vdd.n1675 gnd 0.007278f
C4234 vdd.n1676 gnd 0.00326f
C4235 vdd.n1677 gnd 0.00573f
C4236 vdd.n1678 gnd 0.003079f
C4237 vdd.n1679 gnd 0.005458f
C4238 vdd.n1680 gnd 0.005474f
C4239 vdd.t146 gnd 0.015635f
C4240 vdd.n1681 gnd 0.034788f
C4241 vdd.n1682 gnd 0.181046f
C4242 vdd.n1683 gnd 0.003079f
C4243 vdd.n1684 gnd 0.00326f
C4244 vdd.n1685 gnd 0.007278f
C4245 vdd.n1686 gnd 0.007278f
C4246 vdd.n1687 gnd 0.00326f
C4247 vdd.n1688 gnd 0.003079f
C4248 vdd.n1689 gnd 0.00573f
C4249 vdd.n1690 gnd 0.00573f
C4250 vdd.n1691 gnd 0.003079f
C4251 vdd.n1692 gnd 0.00326f
C4252 vdd.n1693 gnd 0.007278f
C4253 vdd.n1694 gnd 0.007278f
C4254 vdd.n1695 gnd 0.00326f
C4255 vdd.n1696 gnd 0.003079f
C4256 vdd.n1697 gnd 0.00573f
C4257 vdd.n1698 gnd 0.00573f
C4258 vdd.n1699 gnd 0.003079f
C4259 vdd.n1700 gnd 0.00326f
C4260 vdd.n1701 gnd 0.007278f
C4261 vdd.n1702 gnd 0.007278f
C4262 vdd.n1703 gnd 0.017206f
C4263 vdd.n1704 gnd 0.00317f
C4264 vdd.n1705 gnd 0.003079f
C4265 vdd.n1706 gnd 0.01481f
C4266 vdd.n1707 gnd 0.010015f
C4267 vdd.n1708 gnd 0.069923f
C4268 vdd.n1709 gnd 0.25195f
C4269 vdd.n1710 gnd 0.006175f
C4270 vdd.n1711 gnd 0.00573f
C4271 vdd.n1712 gnd 0.00317f
C4272 vdd.n1713 gnd 0.007278f
C4273 vdd.n1714 gnd 0.003079f
C4274 vdd.n1715 gnd 0.00326f
C4275 vdd.n1716 gnd 0.00573f
C4276 vdd.n1717 gnd 0.003079f
C4277 vdd.n1718 gnd 0.007278f
C4278 vdd.n1719 gnd 0.00326f
C4279 vdd.n1720 gnd 0.00573f
C4280 vdd.n1721 gnd 0.003079f
C4281 vdd.n1722 gnd 0.005458f
C4282 vdd.n1723 gnd 0.005474f
C4283 vdd.t280 gnd 0.015635f
C4284 vdd.n1724 gnd 0.034788f
C4285 vdd.n1725 gnd 0.181046f
C4286 vdd.n1726 gnd 0.003079f
C4287 vdd.n1727 gnd 0.00326f
C4288 vdd.n1728 gnd 0.007278f
C4289 vdd.n1729 gnd 0.007278f
C4290 vdd.n1730 gnd 0.00326f
C4291 vdd.n1731 gnd 0.003079f
C4292 vdd.n1732 gnd 0.00573f
C4293 vdd.n1733 gnd 0.00573f
C4294 vdd.n1734 gnd 0.003079f
C4295 vdd.n1735 gnd 0.00326f
C4296 vdd.n1736 gnd 0.007278f
C4297 vdd.n1737 gnd 0.007278f
C4298 vdd.n1738 gnd 0.00326f
C4299 vdd.n1739 gnd 0.003079f
C4300 vdd.n1740 gnd 0.00573f
C4301 vdd.n1741 gnd 0.00573f
C4302 vdd.n1742 gnd 0.003079f
C4303 vdd.n1743 gnd 0.00326f
C4304 vdd.n1744 gnd 0.007278f
C4305 vdd.n1745 gnd 0.007278f
C4306 vdd.n1746 gnd 0.017206f
C4307 vdd.n1747 gnd 0.00317f
C4308 vdd.n1748 gnd 0.003079f
C4309 vdd.n1749 gnd 0.01481f
C4310 vdd.n1750 gnd 0.010339f
C4311 vdd.t171 gnd 0.036223f
C4312 vdd.t281 gnd 0.036223f
C4313 vdd.n1751 gnd 0.248951f
C4314 vdd.n1752 gnd 0.195762f
C4315 vdd.t278 gnd 0.036223f
C4316 vdd.t261 gnd 0.036223f
C4317 vdd.n1753 gnd 0.248951f
C4318 vdd.n1754 gnd 0.157979f
C4319 vdd.t228 gnd 0.036223f
C4320 vdd.t168 gnd 0.036223f
C4321 vdd.n1755 gnd 0.248951f
C4322 vdd.n1756 gnd 0.157979f
C4323 vdd.t290 gnd 0.036223f
C4324 vdd.t258 gnd 0.036223f
C4325 vdd.n1757 gnd 0.248951f
C4326 vdd.n1758 gnd 0.157979f
C4327 vdd.t239 gnd 0.036223f
C4328 vdd.t202 gnd 0.036223f
C4329 vdd.n1759 gnd 0.248951f
C4330 vdd.n1760 gnd 0.157979f
C4331 vdd.t198 gnd 0.036223f
C4332 vdd.t256 gnd 0.036223f
C4333 vdd.n1761 gnd 0.248951f
C4334 vdd.n1762 gnd 0.157979f
C4335 vdd.t241 gnd 0.036223f
C4336 vdd.t240 gnd 0.036223f
C4337 vdd.n1763 gnd 0.248951f
C4338 vdd.n1764 gnd 0.157979f
C4339 vdd.t195 gnd 0.036223f
C4340 vdd.t170 gnd 0.036223f
C4341 vdd.n1765 gnd 0.248951f
C4342 vdd.n1766 gnd 0.157979f
C4343 vdd.t166 gnd 0.036223f
C4344 vdd.t236 gnd 0.036223f
C4345 vdd.n1767 gnd 0.248951f
C4346 vdd.n1768 gnd 0.157979f
C4347 vdd.n1769 gnd 0.006175f
C4348 vdd.n1770 gnd 0.00573f
C4349 vdd.n1771 gnd 0.00317f
C4350 vdd.n1772 gnd 0.007278f
C4351 vdd.n1773 gnd 0.003079f
C4352 vdd.n1774 gnd 0.00326f
C4353 vdd.n1775 gnd 0.00573f
C4354 vdd.n1776 gnd 0.003079f
C4355 vdd.n1777 gnd 0.007278f
C4356 vdd.n1778 gnd 0.00326f
C4357 vdd.n1779 gnd 0.00573f
C4358 vdd.n1780 gnd 0.003079f
C4359 vdd.n1781 gnd 0.005458f
C4360 vdd.n1782 gnd 0.005474f
C4361 vdd.t167 gnd 0.015635f
C4362 vdd.n1783 gnd 0.034788f
C4363 vdd.n1784 gnd 0.181046f
C4364 vdd.n1785 gnd 0.003079f
C4365 vdd.n1786 gnd 0.00326f
C4366 vdd.n1787 gnd 0.007278f
C4367 vdd.n1788 gnd 0.007278f
C4368 vdd.n1789 gnd 0.00326f
C4369 vdd.n1790 gnd 0.003079f
C4370 vdd.n1791 gnd 0.00573f
C4371 vdd.n1792 gnd 0.00573f
C4372 vdd.n1793 gnd 0.003079f
C4373 vdd.n1794 gnd 0.00326f
C4374 vdd.n1795 gnd 0.007278f
C4375 vdd.n1796 gnd 0.007278f
C4376 vdd.n1797 gnd 0.00326f
C4377 vdd.n1798 gnd 0.003079f
C4378 vdd.n1799 gnd 0.00573f
C4379 vdd.n1800 gnd 0.00573f
C4380 vdd.n1801 gnd 0.003079f
C4381 vdd.n1802 gnd 0.00326f
C4382 vdd.n1803 gnd 0.007278f
C4383 vdd.n1804 gnd 0.007278f
C4384 vdd.n1805 gnd 0.017206f
C4385 vdd.n1806 gnd 0.00317f
C4386 vdd.n1807 gnd 0.003079f
C4387 vdd.n1808 gnd 0.01481f
C4388 vdd.n1809 gnd 0.010015f
C4389 vdd.n1810 gnd 0.069923f
C4390 vdd.n1811 gnd 0.288427f
C4391 vdd.n1812 gnd 2.88974f
C4392 vdd.n1813 gnd 0.663635f
C4393 vdd.n1814 gnd 0.008647f
C4394 vdd.n1815 gnd 0.009056f
C4395 vdd.n1816 gnd 0.011251f
C4396 vdd.n1817 gnd 0.822116f
C4397 vdd.n1818 gnd 0.011251f
C4398 vdd.n1819 gnd 0.009056f
C4399 vdd.n1820 gnd 0.011251f
C4400 vdd.n1821 gnd 0.011251f
C4401 vdd.n1822 gnd 0.011251f
C4402 vdd.n1823 gnd 0.009056f
C4403 vdd.n1824 gnd 0.011251f
C4404 vdd.n1825 gnd 0.954345f
C4405 vdd.t230 gnd 0.574906f
C4406 vdd.n1826 gnd 0.626648f
C4407 vdd.n1827 gnd 0.011251f
C4408 vdd.n1828 gnd 0.009056f
C4409 vdd.n1829 gnd 0.011251f
C4410 vdd.n1830 gnd 0.011251f
C4411 vdd.n1831 gnd 0.011251f
C4412 vdd.n1832 gnd 0.009056f
C4413 vdd.n1833 gnd 0.011251f
C4414 vdd.n1834 gnd 0.718633f
C4415 vdd.n1835 gnd 0.011251f
C4416 vdd.n1836 gnd 0.009056f
C4417 vdd.n1837 gnd 0.011251f
C4418 vdd.n1838 gnd 0.011251f
C4419 vdd.n1839 gnd 0.011251f
C4420 vdd.n1840 gnd 0.009056f
C4421 vdd.n1841 gnd 0.011251f
C4422 vdd.n1842 gnd 0.61515f
C4423 vdd.n1843 gnd 0.914101f
C4424 vdd.n1844 gnd 0.011251f
C4425 vdd.n1845 gnd 0.009056f
C4426 vdd.n1846 gnd 0.011251f
C4427 vdd.n1847 gnd 0.011251f
C4428 vdd.n1848 gnd 0.011251f
C4429 vdd.n1849 gnd 0.009056f
C4430 vdd.n1850 gnd 0.011251f
C4431 vdd.n1851 gnd 0.954345f
C4432 vdd.n1852 gnd 0.011251f
C4433 vdd.n1853 gnd 0.009056f
C4434 vdd.n1854 gnd 0.011251f
C4435 vdd.n1855 gnd 0.011251f
C4436 vdd.n1856 gnd 0.011251f
C4437 vdd.n1857 gnd 0.009056f
C4438 vdd.n1858 gnd 0.011251f
C4439 vdd.t249 gnd 0.574906f
C4440 vdd.n1859 gnd 0.79912f
C4441 vdd.n1860 gnd 0.011251f
C4442 vdd.n1861 gnd 0.009056f
C4443 vdd.n1862 gnd 0.011251f
C4444 vdd.n1863 gnd 0.011251f
C4445 vdd.n1864 gnd 0.011251f
C4446 vdd.n1865 gnd 0.009056f
C4447 vdd.n1866 gnd 0.011251f
C4448 vdd.n1867 gnd 0.603652f
C4449 vdd.n1868 gnd 0.011251f
C4450 vdd.n1869 gnd 0.009056f
C4451 vdd.n1870 gnd 0.011251f
C4452 vdd.n1871 gnd 0.011251f
C4453 vdd.n1872 gnd 0.011251f
C4454 vdd.n1873 gnd 0.009056f
C4455 vdd.n1874 gnd 0.011251f
C4456 vdd.n1875 gnd 0.787622f
C4457 vdd.n1876 gnd 0.741629f
C4458 vdd.n1877 gnd 0.011251f
C4459 vdd.n1878 gnd 0.009056f
C4460 vdd.n1879 gnd 0.011251f
C4461 vdd.n1880 gnd 0.011251f
C4462 vdd.n1881 gnd 0.011251f
C4463 vdd.n1882 gnd 0.009056f
C4464 vdd.n1883 gnd 0.011251f
C4465 vdd.n1884 gnd 0.937097f
C4466 vdd.n1885 gnd 0.011251f
C4467 vdd.n1886 gnd 0.009056f
C4468 vdd.n1887 gnd 0.011251f
C4469 vdd.n1888 gnd 0.011251f
C4470 vdd.n1889 gnd 0.027217f
C4471 vdd.n1890 gnd 0.011251f
C4472 vdd.n1891 gnd 0.011251f
C4473 vdd.n1892 gnd 0.009056f
C4474 vdd.n1893 gnd 0.011251f
C4475 vdd.n1894 gnd 0.695637f
C4476 vdd.n1895 gnd 1.14981f
C4477 vdd.n1896 gnd 0.011251f
C4478 vdd.n1897 gnd 0.009056f
C4479 vdd.n1898 gnd 0.011251f
C4480 vdd.n1899 gnd 0.011251f
C4481 vdd.n1900 gnd 0.009676f
C4482 vdd.n1901 gnd 0.009056f
C4483 vdd.n1903 gnd 0.011251f
C4484 vdd.n1905 gnd 0.009056f
C4485 vdd.n1906 gnd 0.011251f
C4486 vdd.n1907 gnd 0.009056f
C4487 vdd.n1909 gnd 0.011251f
C4488 vdd.n1910 gnd 0.009056f
C4489 vdd.n1911 gnd 0.011251f
C4490 vdd.n1912 gnd 0.011251f
C4491 vdd.n1913 gnd 0.011251f
C4492 vdd.n1914 gnd 0.011251f
C4493 vdd.n1915 gnd 0.011251f
C4494 vdd.n1916 gnd 0.009056f
C4495 vdd.n1918 gnd 0.011251f
C4496 vdd.n1919 gnd 0.011251f
C4497 vdd.n1920 gnd 0.011251f
C4498 vdd.n1921 gnd 0.011251f
C4499 vdd.n1922 gnd 0.011251f
C4500 vdd.n1923 gnd 0.009056f
C4501 vdd.n1925 gnd 0.011251f
C4502 vdd.n1926 gnd 0.011251f
C4503 vdd.n1927 gnd 0.011251f
C4504 vdd.n1928 gnd 0.011251f
C4505 vdd.n1929 gnd 0.007562f
C4506 vdd.t49 gnd 0.138418f
C4507 vdd.t48 gnd 0.147931f
C4508 vdd.t47 gnd 0.180773f
C4509 vdd.n1930 gnd 0.231725f
C4510 vdd.n1931 gnd 0.194691f
C4511 vdd.n1933 gnd 0.011251f
C4512 vdd.n1934 gnd 0.011251f
C4513 vdd.n1935 gnd 0.009056f
C4514 vdd.n1936 gnd 0.011251f
C4515 vdd.n1938 gnd 0.011251f
C4516 vdd.n1939 gnd 0.011251f
C4517 vdd.n1940 gnd 0.011251f
C4518 vdd.n1941 gnd 0.011251f
C4519 vdd.n1942 gnd 0.009056f
C4520 vdd.n1944 gnd 0.011251f
C4521 vdd.n1945 gnd 0.011251f
C4522 vdd.n1946 gnd 0.011251f
C4523 vdd.n1947 gnd 0.011251f
C4524 vdd.n1948 gnd 0.011251f
C4525 vdd.n1949 gnd 0.009056f
C4526 vdd.n1951 gnd 0.011251f
C4527 vdd.n1952 gnd 0.011251f
C4528 vdd.n1953 gnd 0.011251f
C4529 vdd.n1954 gnd 0.011251f
C4530 vdd.n1955 gnd 0.011251f
C4531 vdd.n1956 gnd 0.009056f
C4532 vdd.n1958 gnd 0.011251f
C4533 vdd.n1959 gnd 0.011251f
C4534 vdd.n1960 gnd 0.011251f
C4535 vdd.n1961 gnd 0.011251f
C4536 vdd.n1962 gnd 0.011251f
C4537 vdd.n1963 gnd 0.009056f
C4538 vdd.n1965 gnd 0.011251f
C4539 vdd.n1966 gnd 0.011251f
C4540 vdd.n1967 gnd 0.011251f
C4541 vdd.n1968 gnd 0.011251f
C4542 vdd.n1969 gnd 0.008965f
C4543 vdd.t36 gnd 0.138418f
C4544 vdd.t35 gnd 0.147931f
C4545 vdd.t34 gnd 0.180773f
C4546 vdd.n1970 gnd 0.231725f
C4547 vdd.n1971 gnd 0.194691f
C4548 vdd.n1973 gnd 0.011251f
C4549 vdd.n1974 gnd 0.011251f
C4550 vdd.n1975 gnd 0.009056f
C4551 vdd.n1976 gnd 0.011251f
C4552 vdd.n1978 gnd 0.011251f
C4553 vdd.n1979 gnd 0.011251f
C4554 vdd.n1980 gnd 0.011251f
C4555 vdd.n1981 gnd 0.011251f
C4556 vdd.n1982 gnd 0.009056f
C4557 vdd.n1984 gnd 0.011251f
C4558 vdd.n1985 gnd 0.011251f
C4559 vdd.n1986 gnd 0.011251f
C4560 vdd.n1987 gnd 0.011251f
C4561 vdd.n1988 gnd 0.011251f
C4562 vdd.n1989 gnd 0.009056f
C4563 vdd.n1991 gnd 0.011251f
C4564 vdd.n1992 gnd 0.011251f
C4565 vdd.n1993 gnd 0.011251f
C4566 vdd.n1994 gnd 0.011251f
C4567 vdd.n1995 gnd 0.011251f
C4568 vdd.n1996 gnd 0.011251f
C4569 vdd.n1997 gnd 0.009056f
C4570 vdd.n1999 gnd 0.011251f
C4571 vdd.n2001 gnd 0.011251f
C4572 vdd.n2002 gnd 0.009056f
C4573 vdd.n2003 gnd 0.009056f
C4574 vdd.n2004 gnd 0.011251f
C4575 vdd.n2006 gnd 0.011251f
C4576 vdd.n2007 gnd 0.009056f
C4577 vdd.n2008 gnd 0.009056f
C4578 vdd.n2009 gnd 0.011251f
C4579 vdd.n2011 gnd 0.011251f
C4580 vdd.n2012 gnd 0.011251f
C4581 vdd.n2013 gnd 0.009056f
C4582 vdd.n2014 gnd 0.009056f
C4583 vdd.n2015 gnd 0.009056f
C4584 vdd.n2016 gnd 0.011251f
C4585 vdd.n2018 gnd 0.011251f
C4586 vdd.n2019 gnd 0.011251f
C4587 vdd.n2020 gnd 0.009056f
C4588 vdd.n2021 gnd 0.009056f
C4589 vdd.n2022 gnd 0.009056f
C4590 vdd.n2023 gnd 0.011251f
C4591 vdd.n2025 gnd 0.011251f
C4592 vdd.n2026 gnd 0.011251f
C4593 vdd.n2027 gnd 0.009056f
C4594 vdd.n2028 gnd 0.009056f
C4595 vdd.n2029 gnd 0.009056f
C4596 vdd.n2030 gnd 0.011251f
C4597 vdd.n2032 gnd 0.011251f
C4598 vdd.n2033 gnd 0.011251f
C4599 vdd.n2034 gnd 0.009056f
C4600 vdd.n2035 gnd 0.011251f
C4601 vdd.n2036 gnd 0.011251f
C4602 vdd.n2037 gnd 0.011251f
C4603 vdd.n2038 gnd 0.018474f
C4604 vdd.n2039 gnd 0.006158f
C4605 vdd.n2040 gnd 0.009056f
C4606 vdd.n2041 gnd 0.011251f
C4607 vdd.n2043 gnd 0.011251f
C4608 vdd.n2044 gnd 0.011251f
C4609 vdd.n2045 gnd 0.009056f
C4610 vdd.n2046 gnd 0.009056f
C4611 vdd.n2047 gnd 0.009056f
C4612 vdd.n2048 gnd 0.011251f
C4613 vdd.n2050 gnd 0.011251f
C4614 vdd.n2051 gnd 0.011251f
C4615 vdd.n2052 gnd 0.009056f
C4616 vdd.n2053 gnd 0.009056f
C4617 vdd.n2054 gnd 0.009056f
C4618 vdd.n2055 gnd 0.011251f
C4619 vdd.n2057 gnd 0.011251f
C4620 vdd.n2058 gnd 0.011251f
C4621 vdd.n2059 gnd 0.009056f
C4622 vdd.n2060 gnd 0.009056f
C4623 vdd.n2061 gnd 0.009056f
C4624 vdd.n2062 gnd 0.011251f
C4625 vdd.n2064 gnd 0.011251f
C4626 vdd.n2065 gnd 0.011251f
C4627 vdd.n2066 gnd 0.009056f
C4628 vdd.n2067 gnd 0.009056f
C4629 vdd.n2068 gnd 0.009056f
C4630 vdd.n2069 gnd 0.011251f
C4631 vdd.n2071 gnd 0.011251f
C4632 vdd.n2072 gnd 0.011251f
C4633 vdd.n2073 gnd 0.009056f
C4634 vdd.n2074 gnd 0.011251f
C4635 vdd.n2075 gnd 0.011251f
C4636 vdd.n2076 gnd 0.011251f
C4637 vdd.n2077 gnd 0.018474f
C4638 vdd.n2078 gnd 0.007562f
C4639 vdd.n2079 gnd 0.009056f
C4640 vdd.n2080 gnd 0.011251f
C4641 vdd.n2082 gnd 0.011251f
C4642 vdd.n2083 gnd 0.011251f
C4643 vdd.n2084 gnd 0.009056f
C4644 vdd.n2085 gnd 0.009056f
C4645 vdd.n2086 gnd 0.009056f
C4646 vdd.n2087 gnd 0.011251f
C4647 vdd.n2089 gnd 0.011251f
C4648 vdd.n2090 gnd 0.011251f
C4649 vdd.n2091 gnd 0.009056f
C4650 vdd.n2092 gnd 0.009056f
C4651 vdd.n2093 gnd 0.009056f
C4652 vdd.n2094 gnd 0.011251f
C4653 vdd.n2096 gnd 0.011251f
C4654 vdd.n2097 gnd 0.011251f
C4655 vdd.n2099 gnd 0.011251f
C4656 vdd.n2100 gnd 0.009056f
C4657 vdd.n2101 gnd 0.007201f
C4658 vdd.n2102 gnd 0.007651f
C4659 vdd.n2103 gnd 0.007651f
C4660 vdd.n2104 gnd 0.007651f
C4661 vdd.n2105 gnd 0.007651f
C4662 vdd.n2106 gnd 0.007651f
C4663 vdd.n2107 gnd 0.007651f
C4664 vdd.n2108 gnd 0.007651f
C4665 vdd.n2109 gnd 0.007651f
C4666 vdd.n2111 gnd 0.007651f
C4667 vdd.n2112 gnd 0.007651f
C4668 vdd.n2113 gnd 0.007651f
C4669 vdd.n2114 gnd 0.007651f
C4670 vdd.n2115 gnd 0.007651f
C4671 vdd.n2117 gnd 0.007651f
C4672 vdd.n2119 gnd 0.007651f
C4673 vdd.n2120 gnd 0.007651f
C4674 vdd.n2121 gnd 0.007651f
C4675 vdd.n2122 gnd 0.007651f
C4676 vdd.n2123 gnd 0.007651f
C4677 vdd.n2125 gnd 0.007651f
C4678 vdd.n2127 gnd 0.007651f
C4679 vdd.n2128 gnd 0.007651f
C4680 vdd.n2129 gnd 0.007651f
C4681 vdd.n2130 gnd 0.007651f
C4682 vdd.n2131 gnd 0.007651f
C4683 vdd.n2133 gnd 0.007651f
C4684 vdd.n2135 gnd 0.007651f
C4685 vdd.n2136 gnd 0.007651f
C4686 vdd.n2137 gnd 0.007651f
C4687 vdd.n2138 gnd 0.007651f
C4688 vdd.n2139 gnd 0.007651f
C4689 vdd.n2141 gnd 0.007651f
C4690 vdd.n2142 gnd 0.007651f
C4691 vdd.n2143 gnd 0.007651f
C4692 vdd.n2144 gnd 0.007651f
C4693 vdd.n2145 gnd 0.007651f
C4694 vdd.n2146 gnd 0.007651f
C4695 vdd.n2147 gnd 0.007651f
C4696 vdd.n2148 gnd 0.007651f
C4697 vdd.n2149 gnd 0.005569f
C4698 vdd.n2150 gnd 0.007651f
C4699 vdd.t13 gnd 0.309167f
C4700 vdd.t14 gnd 0.316471f
C4701 vdd.t11 gnd 0.201836f
C4702 vdd.n2151 gnd 0.109081f
C4703 vdd.n2152 gnd 0.061874f
C4704 vdd.n2153 gnd 0.010934f
C4705 vdd.n2154 gnd 0.007651f
C4706 vdd.n2155 gnd 0.007651f
C4707 vdd.n2156 gnd 0.465674f
C4708 vdd.n2157 gnd 0.007651f
C4709 vdd.n2158 gnd 0.007651f
C4710 vdd.n2159 gnd 0.007651f
C4711 vdd.n2160 gnd 0.007651f
C4712 vdd.n2161 gnd 0.007651f
C4713 vdd.n2162 gnd 0.007651f
C4714 vdd.n2163 gnd 0.007651f
C4715 vdd.n2164 gnd 0.007651f
C4716 vdd.n2165 gnd 0.007651f
C4717 vdd.n2166 gnd 0.007651f
C4718 vdd.n2167 gnd 0.007651f
C4719 vdd.n2168 gnd 0.007651f
C4720 vdd.n2169 gnd 0.007651f
C4721 vdd.n2170 gnd 0.007651f
C4722 vdd.n2171 gnd 0.007651f
C4723 vdd.n2172 gnd 0.007651f
C4724 vdd.n2173 gnd 0.007651f
C4725 vdd.n2174 gnd 0.007651f
C4726 vdd.n2175 gnd 0.007651f
C4727 vdd.n2176 gnd 0.007651f
C4728 vdd.t66 gnd 0.309167f
C4729 vdd.t67 gnd 0.316471f
C4730 vdd.t65 gnd 0.201836f
C4731 vdd.n2177 gnd 0.109081f
C4732 vdd.n2178 gnd 0.061874f
C4733 vdd.n2179 gnd 0.007651f
C4734 vdd.n2180 gnd 0.007651f
C4735 vdd.n2181 gnd 0.007651f
C4736 vdd.n2182 gnd 0.007651f
C4737 vdd.n2183 gnd 0.007651f
C4738 vdd.n2184 gnd 0.007651f
C4739 vdd.n2186 gnd 0.007651f
C4740 vdd.n2187 gnd 0.007651f
C4741 vdd.n2188 gnd 0.007651f
C4742 vdd.n2189 gnd 0.007651f
C4743 vdd.n2191 gnd 0.007651f
C4744 vdd.n2193 gnd 0.007651f
C4745 vdd.n2194 gnd 0.007651f
C4746 vdd.n2195 gnd 0.007651f
C4747 vdd.n2196 gnd 0.007651f
C4748 vdd.n2197 gnd 0.007651f
C4749 vdd.n2199 gnd 0.007651f
C4750 vdd.n2201 gnd 0.007651f
C4751 vdd.n2202 gnd 0.007651f
C4752 vdd.n2203 gnd 0.007651f
C4753 vdd.n2204 gnd 0.007651f
C4754 vdd.n2205 gnd 0.007651f
C4755 vdd.n2207 gnd 0.007651f
C4756 vdd.n2209 gnd 0.007651f
C4757 vdd.n2210 gnd 0.007651f
C4758 vdd.n2211 gnd 0.005569f
C4759 vdd.n2212 gnd 0.010934f
C4760 vdd.n2213 gnd 0.005907f
C4761 vdd.n2214 gnd 0.007651f
C4762 vdd.n2216 gnd 0.007651f
C4763 vdd.n2217 gnd 0.018154f
C4764 vdd.n2218 gnd 0.018154f
C4765 vdd.n2219 gnd 0.01695f
C4766 vdd.n2220 gnd 0.007651f
C4767 vdd.n2221 gnd 0.007651f
C4768 vdd.n2222 gnd 0.007651f
C4769 vdd.n2223 gnd 0.007651f
C4770 vdd.n2224 gnd 0.007651f
C4771 vdd.n2225 gnd 0.007651f
C4772 vdd.n2226 gnd 0.007651f
C4773 vdd.n2227 gnd 0.007651f
C4774 vdd.n2228 gnd 0.007651f
C4775 vdd.n2229 gnd 0.007651f
C4776 vdd.n2230 gnd 0.007651f
C4777 vdd.n2231 gnd 0.007651f
C4778 vdd.n2232 gnd 0.007651f
C4779 vdd.n2233 gnd 0.007651f
C4780 vdd.n2234 gnd 0.007651f
C4781 vdd.n2235 gnd 0.007651f
C4782 vdd.n2236 gnd 0.007651f
C4783 vdd.n2237 gnd 0.007651f
C4784 vdd.n2238 gnd 0.007651f
C4785 vdd.n2239 gnd 0.007651f
C4786 vdd.n2240 gnd 0.007651f
C4787 vdd.n2241 gnd 0.007651f
C4788 vdd.n2242 gnd 0.007651f
C4789 vdd.n2243 gnd 0.007651f
C4790 vdd.n2244 gnd 0.007651f
C4791 vdd.n2245 gnd 0.007651f
C4792 vdd.n2246 gnd 0.007651f
C4793 vdd.n2247 gnd 0.007651f
C4794 vdd.n2248 gnd 0.007651f
C4795 vdd.n2249 gnd 0.007651f
C4796 vdd.n2250 gnd 0.007651f
C4797 vdd.n2251 gnd 0.007651f
C4798 vdd.n2252 gnd 0.007651f
C4799 vdd.n2253 gnd 0.007651f
C4800 vdd.n2254 gnd 0.007651f
C4801 vdd.n2255 gnd 0.007651f
C4802 vdd.n2256 gnd 0.007651f
C4803 vdd.n2257 gnd 0.24721f
C4804 vdd.n2258 gnd 0.007651f
C4805 vdd.n2259 gnd 0.007651f
C4806 vdd.n2260 gnd 0.007651f
C4807 vdd.n2261 gnd 0.007651f
C4808 vdd.n2262 gnd 0.007651f
C4809 vdd.n2263 gnd 0.007651f
C4810 vdd.n2264 gnd 0.007651f
C4811 vdd.n2265 gnd 0.007651f
C4812 vdd.n2266 gnd 0.007651f
C4813 vdd.n2267 gnd 0.007651f
C4814 vdd.n2268 gnd 0.007651f
C4815 vdd.n2269 gnd 0.007651f
C4816 vdd.n2270 gnd 0.007651f
C4817 vdd.n2271 gnd 0.007651f
C4818 vdd.n2272 gnd 0.007651f
C4819 vdd.n2273 gnd 0.007651f
C4820 vdd.n2274 gnd 0.007651f
C4821 vdd.n2275 gnd 0.007651f
C4822 vdd.n2276 gnd 0.007651f
C4823 vdd.n2277 gnd 0.007651f
C4824 vdd.n2278 gnd 0.01695f
C4825 vdd.n2280 gnd 0.018154f
C4826 vdd.n2281 gnd 0.018154f
C4827 vdd.n2282 gnd 0.007651f
C4828 vdd.n2283 gnd 0.005907f
C4829 vdd.n2284 gnd 0.007651f
C4830 vdd.n2286 gnd 0.007651f
C4831 vdd.n2288 gnd 0.007651f
C4832 vdd.n2289 gnd 0.007651f
C4833 vdd.n2290 gnd 0.007651f
C4834 vdd.n2291 gnd 0.007651f
C4835 vdd.n2292 gnd 0.007651f
C4836 vdd.n2294 gnd 0.007651f
C4837 vdd.n2296 gnd 0.007651f
C4838 vdd.n2297 gnd 0.007651f
C4839 vdd.n2298 gnd 0.007651f
C4840 vdd.n2299 gnd 0.007651f
C4841 vdd.n2300 gnd 0.007651f
C4842 vdd.n2302 gnd 0.007651f
C4843 vdd.n2304 gnd 0.007651f
C4844 vdd.n2305 gnd 0.007651f
C4845 vdd.n2306 gnd 0.007651f
C4846 vdd.n2307 gnd 0.007651f
C4847 vdd.n2308 gnd 0.007651f
C4848 vdd.n2310 gnd 0.007651f
C4849 vdd.n2312 gnd 0.007651f
C4850 vdd.n2313 gnd 0.007651f
C4851 vdd.n2314 gnd 0.022821f
C4852 vdd.n2315 gnd 0.676502f
C4853 vdd.n2317 gnd 0.009056f
C4854 vdd.n2318 gnd 0.009056f
C4855 vdd.n2319 gnd 0.011251f
C4856 vdd.n2321 gnd 0.011251f
C4857 vdd.n2322 gnd 0.011251f
C4858 vdd.n2323 gnd 0.009056f
C4859 vdd.n2324 gnd 0.007516f
C4860 vdd.n2325 gnd 0.027801f
C4861 vdd.n2326 gnd 0.027217f
C4862 vdd.n2327 gnd 0.007516f
C4863 vdd.n2328 gnd 0.027217f
C4864 vdd.n2329 gnd 1.58099f
C4865 vdd.n2330 gnd 0.027217f
C4866 vdd.n2331 gnd 0.027801f
C4867 vdd.n2332 gnd 0.004302f
C4868 vdd.t25 gnd 0.138418f
C4869 vdd.t24 gnd 0.147931f
C4870 vdd.t22 gnd 0.180773f
C4871 vdd.n2333 gnd 0.231725f
C4872 vdd.n2334 gnd 0.194691f
C4873 vdd.n2335 gnd 0.013946f
C4874 vdd.n2336 gnd 0.004754f
C4875 vdd.n2337 gnd 0.009676f
C4876 vdd.n2338 gnd 0.676502f
C4877 vdd.n2339 gnd 0.022821f
C4878 vdd.n2340 gnd 0.007651f
C4879 vdd.n2341 gnd 0.007651f
C4880 vdd.n2342 gnd 0.007651f
C4881 vdd.n2344 gnd 0.007651f
C4882 vdd.n2346 gnd 0.007651f
C4883 vdd.n2347 gnd 0.007651f
C4884 vdd.n2348 gnd 0.007651f
C4885 vdd.n2349 gnd 0.007651f
C4886 vdd.n2350 gnd 0.007651f
C4887 vdd.n2352 gnd 0.007651f
C4888 vdd.n2354 gnd 0.007651f
C4889 vdd.n2355 gnd 0.007651f
C4890 vdd.n2356 gnd 0.007651f
C4891 vdd.n2357 gnd 0.007651f
C4892 vdd.n2358 gnd 0.007651f
C4893 vdd.n2360 gnd 0.007651f
C4894 vdd.n2362 gnd 0.007651f
C4895 vdd.n2363 gnd 0.007651f
C4896 vdd.n2364 gnd 0.007651f
C4897 vdd.n2365 gnd 0.007651f
C4898 vdd.n2366 gnd 0.007651f
C4899 vdd.n2368 gnd 0.007651f
C4900 vdd.n2370 gnd 0.007651f
C4901 vdd.n2371 gnd 0.007651f
C4902 vdd.n2372 gnd 0.018154f
C4903 vdd.n2373 gnd 0.01695f
C4904 vdd.n2374 gnd 0.01695f
C4905 vdd.n2375 gnd 1.12682f
C4906 vdd.n2376 gnd 0.01695f
C4907 vdd.n2377 gnd 0.01695f
C4908 vdd.n2378 gnd 0.007651f
C4909 vdd.n2379 gnd 0.007651f
C4910 vdd.n2380 gnd 0.007651f
C4911 vdd.n2381 gnd 0.48867f
C4912 vdd.n2382 gnd 0.007651f
C4913 vdd.n2383 gnd 0.007651f
C4914 vdd.n2384 gnd 0.007651f
C4915 vdd.n2385 gnd 0.007651f
C4916 vdd.n2386 gnd 0.007651f
C4917 vdd.n2387 gnd 0.781873f
C4918 vdd.n2388 gnd 0.007651f
C4919 vdd.n2389 gnd 0.007651f
C4920 vdd.n2390 gnd 0.007651f
C4921 vdd.n2391 gnd 0.007651f
C4922 vdd.n2392 gnd 0.007651f
C4923 vdd.n2393 gnd 0.781873f
C4924 vdd.n2394 gnd 0.007651f
C4925 vdd.n2395 gnd 0.007651f
C4926 vdd.n2396 gnd 0.006751f
C4927 vdd.n2397 gnd 0.022163f
C4928 vdd.n2398 gnd 0.004725f
C4929 vdd.n2399 gnd 0.007651f
C4930 vdd.n2400 gnd 0.43118f
C4931 vdd.n2401 gnd 0.007651f
C4932 vdd.n2402 gnd 0.007651f
C4933 vdd.n2403 gnd 0.007651f
C4934 vdd.n2404 gnd 0.007651f
C4935 vdd.n2405 gnd 0.007651f
C4936 vdd.n2406 gnd 0.523165f
C4937 vdd.n2407 gnd 0.007651f
C4938 vdd.n2408 gnd 0.007651f
C4939 vdd.n2409 gnd 0.007651f
C4940 vdd.n2410 gnd 0.007651f
C4941 vdd.n2411 gnd 0.007651f
C4942 vdd.n2412 gnd 0.695637f
C4943 vdd.n2413 gnd 0.007651f
C4944 vdd.n2414 gnd 0.007651f
C4945 vdd.n2415 gnd 0.007651f
C4946 vdd.n2416 gnd 0.007651f
C4947 vdd.n2417 gnd 0.007651f
C4948 vdd.n2418 gnd 0.620899f
C4949 vdd.n2419 gnd 0.007651f
C4950 vdd.n2420 gnd 0.007651f
C4951 vdd.n2421 gnd 0.007651f
C4952 vdd.n2422 gnd 0.007651f
C4953 vdd.n2423 gnd 0.007651f
C4954 vdd.n2424 gnd 0.448427f
C4955 vdd.n2425 gnd 0.007651f
C4956 vdd.n2426 gnd 0.007651f
C4957 vdd.n2427 gnd 0.007651f
C4958 vdd.n2428 gnd 0.007651f
C4959 vdd.n2429 gnd 0.007651f
C4960 vdd.n2430 gnd 0.24721f
C4961 vdd.n2431 gnd 0.007651f
C4962 vdd.n2432 gnd 0.007651f
C4963 vdd.n2433 gnd 0.007651f
C4964 vdd.n2434 gnd 0.007651f
C4965 vdd.n2435 gnd 0.007651f
C4966 vdd.n2436 gnd 0.43118f
C4967 vdd.n2437 gnd 0.007651f
C4968 vdd.n2438 gnd 0.007651f
C4969 vdd.n2439 gnd 0.007651f
C4970 vdd.n2440 gnd 0.007651f
C4971 vdd.n2441 gnd 0.007651f
C4972 vdd.n2442 gnd 0.781873f
C4973 vdd.n2443 gnd 0.007651f
C4974 vdd.n2444 gnd 0.007651f
C4975 vdd.n2445 gnd 0.007651f
C4976 vdd.n2446 gnd 0.007651f
C4977 vdd.n2447 gnd 0.007651f
C4978 vdd.n2448 gnd 0.007651f
C4979 vdd.n2449 gnd 0.007651f
C4980 vdd.n2450 gnd 0.609401f
C4981 vdd.n2451 gnd 0.007651f
C4982 vdd.n2452 gnd 0.007651f
C4983 vdd.n2453 gnd 0.007651f
C4984 vdd.n2454 gnd 0.007651f
C4985 vdd.n2455 gnd 0.007651f
C4986 vdd.n2456 gnd 0.007651f
C4987 vdd.n2457 gnd 0.48867f
C4988 vdd.n2458 gnd 0.007651f
C4989 vdd.n2459 gnd 0.007651f
C4990 vdd.n2460 gnd 0.007651f
C4991 vdd.n2461 gnd 0.017881f
C4992 vdd.n2462 gnd 0.017222f
C4993 vdd.n2463 gnd 0.007651f
C4994 vdd.n2464 gnd 0.007651f
C4995 vdd.n2465 gnd 0.005907f
C4996 vdd.n2466 gnd 0.007651f
C4997 vdd.n2467 gnd 0.007651f
C4998 vdd.n2468 gnd 0.005569f
C4999 vdd.n2469 gnd 0.007651f
C5000 vdd.n2470 gnd 0.007651f
C5001 vdd.n2471 gnd 0.007651f
C5002 vdd.n2472 gnd 0.007651f
C5003 vdd.n2473 gnd 0.007651f
C5004 vdd.n2474 gnd 0.007651f
C5005 vdd.n2475 gnd 0.007651f
C5006 vdd.n2476 gnd 0.007651f
C5007 vdd.n2477 gnd 0.007651f
C5008 vdd.n2478 gnd 0.007651f
C5009 vdd.n2479 gnd 0.007651f
C5010 vdd.n2480 gnd 0.007651f
C5011 vdd.n2481 gnd 0.007651f
C5012 vdd.n2482 gnd 0.007651f
C5013 vdd.n2483 gnd 0.007651f
C5014 vdd.n2484 gnd 0.007651f
C5015 vdd.n2485 gnd 0.007651f
C5016 vdd.n2486 gnd 0.007651f
C5017 vdd.n2487 gnd 0.007651f
C5018 vdd.n2488 gnd 0.007651f
C5019 vdd.n2489 gnd 0.007651f
C5020 vdd.n2490 gnd 0.007651f
C5021 vdd.n2491 gnd 0.007651f
C5022 vdd.n2492 gnd 0.007651f
C5023 vdd.n2493 gnd 0.007651f
C5024 vdd.n2494 gnd 0.007651f
C5025 vdd.n2495 gnd 0.007651f
C5026 vdd.n2496 gnd 0.007651f
C5027 vdd.n2497 gnd 0.007651f
C5028 vdd.n2498 gnd 0.007651f
C5029 vdd.n2499 gnd 0.007651f
C5030 vdd.n2500 gnd 0.007651f
C5031 vdd.n2501 gnd 0.007651f
C5032 vdd.n2502 gnd 0.007651f
C5033 vdd.n2503 gnd 0.007651f
C5034 vdd.n2504 gnd 0.007651f
C5035 vdd.n2505 gnd 0.007651f
C5036 vdd.n2506 gnd 0.007651f
C5037 vdd.n2507 gnd 0.007651f
C5038 vdd.n2508 gnd 0.007651f
C5039 vdd.n2509 gnd 0.007651f
C5040 vdd.n2510 gnd 0.007651f
C5041 vdd.n2511 gnd 0.007651f
C5042 vdd.n2512 gnd 0.007651f
C5043 vdd.n2513 gnd 0.007651f
C5044 vdd.n2514 gnd 0.007651f
C5045 vdd.n2515 gnd 0.007651f
C5046 vdd.n2516 gnd 0.007651f
C5047 vdd.n2517 gnd 0.007651f
C5048 vdd.n2518 gnd 0.007651f
C5049 vdd.n2519 gnd 0.007651f
C5050 vdd.n2520 gnd 0.007651f
C5051 vdd.n2521 gnd 0.007651f
C5052 vdd.n2522 gnd 0.007651f
C5053 vdd.n2523 gnd 0.007651f
C5054 vdd.n2524 gnd 0.007651f
C5055 vdd.n2525 gnd 0.007651f
C5056 vdd.n2526 gnd 0.007651f
C5057 vdd.n2527 gnd 0.007651f
C5058 vdd.n2528 gnd 0.007651f
C5059 vdd.n2529 gnd 0.018154f
C5060 vdd.n2530 gnd 0.01695f
C5061 vdd.n2531 gnd 0.01695f
C5062 vdd.n2532 gnd 0.954345f
C5063 vdd.n2533 gnd 0.01695f
C5064 vdd.n2534 gnd 0.018154f
C5065 vdd.n2535 gnd 0.017222f
C5066 vdd.n2536 gnd 0.007651f
C5067 vdd.n2537 gnd 0.007651f
C5068 vdd.n2538 gnd 0.007651f
C5069 vdd.n2539 gnd 0.005907f
C5070 vdd.n2540 gnd 0.010934f
C5071 vdd.n2541 gnd 0.005569f
C5072 vdd.n2542 gnd 0.007651f
C5073 vdd.n2543 gnd 0.007651f
C5074 vdd.n2544 gnd 0.007651f
C5075 vdd.n2545 gnd 0.007651f
C5076 vdd.n2546 gnd 0.007651f
C5077 vdd.n2547 gnd 0.007651f
C5078 vdd.n2548 gnd 0.007651f
C5079 vdd.n2549 gnd 0.007651f
C5080 vdd.n2550 gnd 0.007651f
C5081 vdd.n2551 gnd 0.007651f
C5082 vdd.n2552 gnd 0.007651f
C5083 vdd.n2553 gnd 0.007651f
C5084 vdd.n2554 gnd 0.007651f
C5085 vdd.n2555 gnd 0.007651f
C5086 vdd.n2556 gnd 0.007651f
C5087 vdd.n2557 gnd 0.007651f
C5088 vdd.n2558 gnd 0.007651f
C5089 vdd.n2559 gnd 0.007651f
C5090 vdd.n2560 gnd 0.007651f
C5091 vdd.n2561 gnd 0.007651f
C5092 vdd.n2562 gnd 0.007651f
C5093 vdd.n2563 gnd 0.007651f
C5094 vdd.n2564 gnd 0.007651f
C5095 vdd.n2565 gnd 0.007651f
C5096 vdd.n2566 gnd 0.007651f
C5097 vdd.n2567 gnd 0.007651f
C5098 vdd.n2568 gnd 0.007651f
C5099 vdd.n2569 gnd 0.007651f
C5100 vdd.n2570 gnd 0.007651f
C5101 vdd.n2571 gnd 0.007651f
C5102 vdd.n2572 gnd 0.007651f
C5103 vdd.n2573 gnd 0.007651f
C5104 vdd.n2574 gnd 0.007651f
C5105 vdd.n2575 gnd 0.007651f
C5106 vdd.n2576 gnd 0.007651f
C5107 vdd.n2577 gnd 0.007651f
C5108 vdd.n2578 gnd 0.007651f
C5109 vdd.n2579 gnd 0.007651f
C5110 vdd.n2580 gnd 0.007651f
C5111 vdd.n2581 gnd 0.007651f
C5112 vdd.n2582 gnd 0.007651f
C5113 vdd.n2583 gnd 0.007651f
C5114 vdd.n2584 gnd 0.007651f
C5115 vdd.n2585 gnd 0.007651f
C5116 vdd.n2586 gnd 0.007651f
C5117 vdd.n2587 gnd 0.007651f
C5118 vdd.n2588 gnd 0.007651f
C5119 vdd.n2589 gnd 0.007651f
C5120 vdd.n2590 gnd 0.007651f
C5121 vdd.n2591 gnd 0.007651f
C5122 vdd.n2592 gnd 0.007651f
C5123 vdd.n2593 gnd 0.007651f
C5124 vdd.n2594 gnd 0.007651f
C5125 vdd.n2595 gnd 0.007651f
C5126 vdd.n2596 gnd 0.007651f
C5127 vdd.n2597 gnd 0.007651f
C5128 vdd.n2598 gnd 0.007651f
C5129 vdd.n2599 gnd 0.007651f
C5130 vdd.n2600 gnd 0.007651f
C5131 vdd.n2601 gnd 0.007651f
C5132 vdd.n2602 gnd 0.018154f
C5133 vdd.n2603 gnd 0.018154f
C5134 vdd.n2604 gnd 0.954345f
C5135 vdd.t87 gnd 3.39195f
C5136 vdd.t115 gnd 3.39195f
C5137 vdd.n2637 gnd 0.018154f
C5138 vdd.n2638 gnd 0.007651f
C5139 vdd.t60 gnd 0.309167f
C5140 vdd.t61 gnd 0.316471f
C5141 vdd.t58 gnd 0.201836f
C5142 vdd.n2639 gnd 0.109081f
C5143 vdd.n2640 gnd 0.061874f
C5144 vdd.n2641 gnd 0.007651f
C5145 vdd.t73 gnd 0.309167f
C5146 vdd.t74 gnd 0.316471f
C5147 vdd.t72 gnd 0.201836f
C5148 vdd.n2642 gnd 0.109081f
C5149 vdd.n2643 gnd 0.061874f
C5150 vdd.n2644 gnd 0.010934f
C5151 vdd.n2645 gnd 0.007651f
C5152 vdd.n2646 gnd 0.007651f
C5153 vdd.n2647 gnd 0.007651f
C5154 vdd.n2648 gnd 0.007651f
C5155 vdd.n2649 gnd 0.007651f
C5156 vdd.n2650 gnd 0.007651f
C5157 vdd.n2651 gnd 0.007651f
C5158 vdd.n2652 gnd 0.007651f
C5159 vdd.n2653 gnd 0.007651f
C5160 vdd.n2654 gnd 0.007651f
C5161 vdd.n2655 gnd 0.007651f
C5162 vdd.n2656 gnd 0.007651f
C5163 vdd.n2657 gnd 0.007651f
C5164 vdd.n2658 gnd 0.007651f
C5165 vdd.n2659 gnd 0.007651f
C5166 vdd.n2660 gnd 0.007651f
C5167 vdd.n2661 gnd 0.007651f
C5168 vdd.n2662 gnd 0.007651f
C5169 vdd.n2663 gnd 0.007651f
C5170 vdd.n2664 gnd 0.007651f
C5171 vdd.n2665 gnd 0.007651f
C5172 vdd.n2666 gnd 0.007651f
C5173 vdd.n2667 gnd 0.007651f
C5174 vdd.n2668 gnd 0.007651f
C5175 vdd.n2669 gnd 0.007651f
C5176 vdd.n2670 gnd 0.007651f
C5177 vdd.n2671 gnd 0.007651f
C5178 vdd.n2672 gnd 0.007651f
C5179 vdd.n2673 gnd 0.007651f
C5180 vdd.n2674 gnd 0.007651f
C5181 vdd.n2675 gnd 0.007651f
C5182 vdd.n2676 gnd 0.007651f
C5183 vdd.n2677 gnd 0.007651f
C5184 vdd.n2678 gnd 0.007651f
C5185 vdd.n2679 gnd 0.007651f
C5186 vdd.n2680 gnd 0.007651f
C5187 vdd.n2681 gnd 0.007651f
C5188 vdd.n2682 gnd 0.007651f
C5189 vdd.n2683 gnd 0.007651f
C5190 vdd.n2684 gnd 0.007651f
C5191 vdd.n2685 gnd 0.007651f
C5192 vdd.n2686 gnd 0.007651f
C5193 vdd.n2687 gnd 0.007651f
C5194 vdd.n2688 gnd 0.007651f
C5195 vdd.n2689 gnd 0.007651f
C5196 vdd.n2690 gnd 0.007651f
C5197 vdd.n2691 gnd 0.007651f
C5198 vdd.n2692 gnd 0.007651f
C5199 vdd.n2693 gnd 0.007651f
C5200 vdd.n2694 gnd 0.007651f
C5201 vdd.n2695 gnd 0.007651f
C5202 vdd.n2696 gnd 0.007651f
C5203 vdd.n2697 gnd 0.007651f
C5204 vdd.n2698 gnd 0.007651f
C5205 vdd.n2699 gnd 0.007651f
C5206 vdd.n2700 gnd 0.007651f
C5207 vdd.n2701 gnd 0.005569f
C5208 vdd.n2702 gnd 0.007651f
C5209 vdd.n2703 gnd 0.007651f
C5210 vdd.n2704 gnd 0.005907f
C5211 vdd.n2705 gnd 0.007651f
C5212 vdd.n2706 gnd 0.007651f
C5213 vdd.n2707 gnd 0.018154f
C5214 vdd.n2708 gnd 0.01695f
C5215 vdd.n2709 gnd 0.007651f
C5216 vdd.n2710 gnd 0.007651f
C5217 vdd.n2711 gnd 0.007651f
C5218 vdd.n2712 gnd 0.007651f
C5219 vdd.n2713 gnd 0.007651f
C5220 vdd.n2714 gnd 0.007651f
C5221 vdd.n2715 gnd 0.007651f
C5222 vdd.n2716 gnd 0.007651f
C5223 vdd.n2717 gnd 0.007651f
C5224 vdd.n2718 gnd 0.007651f
C5225 vdd.n2719 gnd 0.007651f
C5226 vdd.n2720 gnd 0.007651f
C5227 vdd.n2721 gnd 0.007651f
C5228 vdd.n2722 gnd 0.007651f
C5229 vdd.n2723 gnd 0.007651f
C5230 vdd.n2724 gnd 0.007651f
C5231 vdd.n2725 gnd 0.007651f
C5232 vdd.n2726 gnd 0.007651f
C5233 vdd.n2727 gnd 0.007651f
C5234 vdd.n2728 gnd 0.007651f
C5235 vdd.n2729 gnd 0.007651f
C5236 vdd.n2730 gnd 0.007651f
C5237 vdd.n2731 gnd 0.007651f
C5238 vdd.n2732 gnd 0.007651f
C5239 vdd.n2733 gnd 0.007651f
C5240 vdd.n2734 gnd 0.007651f
C5241 vdd.n2735 gnd 0.007651f
C5242 vdd.n2736 gnd 0.007651f
C5243 vdd.n2737 gnd 0.007651f
C5244 vdd.n2738 gnd 0.007651f
C5245 vdd.n2739 gnd 0.007651f
C5246 vdd.n2740 gnd 0.007651f
C5247 vdd.n2741 gnd 0.007651f
C5248 vdd.n2742 gnd 0.007651f
C5249 vdd.n2743 gnd 0.007651f
C5250 vdd.n2744 gnd 0.007651f
C5251 vdd.n2745 gnd 0.007651f
C5252 vdd.n2746 gnd 0.007651f
C5253 vdd.n2747 gnd 0.007651f
C5254 vdd.n2748 gnd 0.007651f
C5255 vdd.n2749 gnd 0.007651f
C5256 vdd.n2750 gnd 0.007651f
C5257 vdd.n2751 gnd 0.007651f
C5258 vdd.n2752 gnd 0.007651f
C5259 vdd.n2753 gnd 0.007651f
C5260 vdd.n2754 gnd 0.007651f
C5261 vdd.n2755 gnd 0.007651f
C5262 vdd.n2756 gnd 0.007651f
C5263 vdd.n2757 gnd 0.007651f
C5264 vdd.n2758 gnd 0.007651f
C5265 vdd.n2759 gnd 0.007651f
C5266 vdd.n2760 gnd 0.24721f
C5267 vdd.n2761 gnd 0.007651f
C5268 vdd.n2762 gnd 0.007651f
C5269 vdd.n2763 gnd 0.007651f
C5270 vdd.n2764 gnd 0.007651f
C5271 vdd.n2765 gnd 0.007651f
C5272 vdd.n2766 gnd 0.007651f
C5273 vdd.n2767 gnd 0.007651f
C5274 vdd.n2768 gnd 0.007651f
C5275 vdd.n2769 gnd 0.007651f
C5276 vdd.n2770 gnd 0.007651f
C5277 vdd.n2771 gnd 0.007651f
C5278 vdd.n2772 gnd 0.007651f
C5279 vdd.n2773 gnd 0.007651f
C5280 vdd.n2774 gnd 0.007651f
C5281 vdd.n2775 gnd 0.007651f
C5282 vdd.n2776 gnd 0.007651f
C5283 vdd.n2777 gnd 0.007651f
C5284 vdd.n2778 gnd 0.007651f
C5285 vdd.n2779 gnd 0.007651f
C5286 vdd.n2780 gnd 0.007651f
C5287 vdd.n2781 gnd 0.465674f
C5288 vdd.n2782 gnd 0.007651f
C5289 vdd.n2783 gnd 0.007651f
C5290 vdd.n2784 gnd 0.007651f
C5291 vdd.n2785 gnd 0.007651f
C5292 vdd.n2786 gnd 0.007651f
C5293 vdd.n2787 gnd 0.01695f
C5294 vdd.n2788 gnd 0.018154f
C5295 vdd.n2789 gnd 0.018154f
C5296 vdd.n2790 gnd 0.007651f
C5297 vdd.n2791 gnd 0.007651f
C5298 vdd.n2792 gnd 0.007651f
C5299 vdd.n2793 gnd 0.005907f
C5300 vdd.n2794 gnd 0.010934f
C5301 vdd.n2795 gnd 0.005569f
C5302 vdd.n2796 gnd 0.007651f
C5303 vdd.n2797 gnd 0.007651f
C5304 vdd.n2798 gnd 0.007651f
C5305 vdd.n2799 gnd 0.007651f
C5306 vdd.n2800 gnd 0.007651f
C5307 vdd.n2801 gnd 0.007651f
C5308 vdd.n2802 gnd 0.007651f
C5309 vdd.n2803 gnd 0.007651f
C5310 vdd.n2804 gnd 0.007651f
C5311 vdd.n2805 gnd 0.007651f
C5312 vdd.n2806 gnd 0.007651f
C5313 vdd.n2807 gnd 0.007651f
C5314 vdd.n2808 gnd 0.007651f
C5315 vdd.n2809 gnd 0.007651f
C5316 vdd.n2810 gnd 0.007651f
C5317 vdd.n2811 gnd 0.007651f
C5318 vdd.n2812 gnd 0.007651f
C5319 vdd.n2813 gnd 0.007651f
C5320 vdd.n2814 gnd 0.007651f
C5321 vdd.n2815 gnd 0.007651f
C5322 vdd.n2816 gnd 0.007651f
C5323 vdd.n2817 gnd 0.007651f
C5324 vdd.n2818 gnd 0.007651f
C5325 vdd.n2819 gnd 0.007651f
C5326 vdd.n2820 gnd 0.007651f
C5327 vdd.n2821 gnd 0.007651f
C5328 vdd.n2822 gnd 0.007651f
C5329 vdd.n2823 gnd 0.007651f
C5330 vdd.n2824 gnd 0.007651f
C5331 vdd.n2825 gnd 0.007651f
C5332 vdd.n2826 gnd 0.007651f
C5333 vdd.n2827 gnd 0.007651f
C5334 vdd.n2828 gnd 0.007651f
C5335 vdd.n2829 gnd 0.007651f
C5336 vdd.n2830 gnd 0.007651f
C5337 vdd.n2831 gnd 0.007651f
C5338 vdd.n2832 gnd 0.007651f
C5339 vdd.n2833 gnd 0.007651f
C5340 vdd.n2834 gnd 0.007651f
C5341 vdd.n2835 gnd 0.007651f
C5342 vdd.n2836 gnd 0.007651f
C5343 vdd.n2837 gnd 0.007651f
C5344 vdd.n2838 gnd 0.007651f
C5345 vdd.n2839 gnd 0.007651f
C5346 vdd.n2840 gnd 0.007651f
C5347 vdd.n2841 gnd 0.007651f
C5348 vdd.n2842 gnd 0.007651f
C5349 vdd.n2843 gnd 0.007651f
C5350 vdd.n2844 gnd 0.007651f
C5351 vdd.n2845 gnd 0.007651f
C5352 vdd.n2846 gnd 0.007651f
C5353 vdd.n2847 gnd 0.007651f
C5354 vdd.n2848 gnd 0.007651f
C5355 vdd.n2849 gnd 0.007651f
C5356 vdd.n2850 gnd 0.007651f
C5357 vdd.n2851 gnd 0.007651f
C5358 vdd.n2852 gnd 0.007651f
C5359 vdd.n2853 gnd 0.007651f
C5360 vdd.n2854 gnd 0.007651f
C5361 vdd.n2855 gnd 0.007651f
C5362 vdd.n2857 gnd 0.954345f
C5363 vdd.n2859 gnd 0.007651f
C5364 vdd.n2860 gnd 0.007651f
C5365 vdd.n2861 gnd 0.018154f
C5366 vdd.n2862 gnd 0.01695f
C5367 vdd.n2863 gnd 0.01695f
C5368 vdd.n2864 gnd 0.954345f
C5369 vdd.n2865 gnd 0.01695f
C5370 vdd.n2866 gnd 0.01695f
C5371 vdd.n2867 gnd 0.007651f
C5372 vdd.n2868 gnd 0.007651f
C5373 vdd.n2869 gnd 0.007651f
C5374 vdd.n2870 gnd 0.48867f
C5375 vdd.n2871 gnd 0.007651f
C5376 vdd.n2872 gnd 0.007651f
C5377 vdd.n2873 gnd 0.007651f
C5378 vdd.n2874 gnd 0.007651f
C5379 vdd.n2875 gnd 0.007651f
C5380 vdd.n2876 gnd 0.609401f
C5381 vdd.n2877 gnd 0.007651f
C5382 vdd.n2878 gnd 0.007651f
C5383 vdd.n2879 gnd 0.007651f
C5384 vdd.n2880 gnd 0.007651f
C5385 vdd.n2881 gnd 0.007651f
C5386 vdd.n2882 gnd 0.781873f
C5387 vdd.n2883 gnd 0.007651f
C5388 vdd.n2884 gnd 0.007651f
C5389 vdd.n2885 gnd 0.007651f
C5390 vdd.n2886 gnd 0.007651f
C5391 vdd.n2887 gnd 0.007651f
C5392 vdd.n2888 gnd 0.43118f
C5393 vdd.n2889 gnd 0.007651f
C5394 vdd.n2890 gnd 0.007651f
C5395 vdd.n2891 gnd 0.007651f
C5396 vdd.n2892 gnd 0.007651f
C5397 vdd.n2893 gnd 0.007651f
C5398 vdd.n2894 gnd 0.24721f
C5399 vdd.n2895 gnd 0.007651f
C5400 vdd.n2896 gnd 0.007651f
C5401 vdd.n2897 gnd 0.007651f
C5402 vdd.n2898 gnd 0.007651f
C5403 vdd.n2899 gnd 0.007651f
C5404 vdd.n2900 gnd 0.448427f
C5405 vdd.n2901 gnd 0.007651f
C5406 vdd.n2902 gnd 0.007651f
C5407 vdd.n2903 gnd 0.007651f
C5408 vdd.n2904 gnd 0.007651f
C5409 vdd.n2905 gnd 0.007651f
C5410 vdd.n2906 gnd 0.620899f
C5411 vdd.n2907 gnd 0.007651f
C5412 vdd.n2908 gnd 0.007651f
C5413 vdd.n2909 gnd 0.007651f
C5414 vdd.n2910 gnd 0.007651f
C5415 vdd.n2911 gnd 0.007651f
C5416 vdd.n2912 gnd 0.695637f
C5417 vdd.n2913 gnd 0.007651f
C5418 vdd.n2914 gnd 0.007651f
C5419 vdd.n2915 gnd 0.007651f
C5420 vdd.n2916 gnd 0.007651f
C5421 vdd.n2917 gnd 0.007651f
C5422 vdd.n2918 gnd 0.523165f
C5423 vdd.n2919 gnd 0.007651f
C5424 vdd.n2920 gnd 0.007651f
C5425 vdd.n2921 gnd 0.007651f
C5426 vdd.t28 gnd 0.316471f
C5427 vdd.t26 gnd 0.201836f
C5428 vdd.t29 gnd 0.316471f
C5429 vdd.n2922 gnd 0.177869f
C5430 vdd.n2923 gnd 0.022163f
C5431 vdd.n2924 gnd 0.004725f
C5432 vdd.n2925 gnd 0.007651f
C5433 vdd.n2926 gnd 0.43118f
C5434 vdd.n2927 gnd 0.007651f
C5435 vdd.n2928 gnd 0.007651f
C5436 vdd.n2929 gnd 0.007651f
C5437 vdd.n2930 gnd 0.007651f
C5438 vdd.n2931 gnd 0.007651f
C5439 vdd.n2932 gnd 0.781873f
C5440 vdd.n2933 gnd 0.007651f
C5441 vdd.n2934 gnd 0.007651f
C5442 vdd.n2935 gnd 0.007651f
C5443 vdd.n2936 gnd 0.007651f
C5444 vdd.n2937 gnd 0.007651f
C5445 vdd.n2938 gnd 0.007651f
C5446 vdd.n2940 gnd 0.007651f
C5447 vdd.n2941 gnd 0.007651f
C5448 vdd.n2943 gnd 0.007651f
C5449 vdd.n2944 gnd 0.007651f
C5450 vdd.n2947 gnd 0.007651f
C5451 vdd.n2948 gnd 0.007651f
C5452 vdd.n2949 gnd 0.007651f
C5453 vdd.n2950 gnd 0.007651f
C5454 vdd.n2952 gnd 0.007651f
C5455 vdd.n2953 gnd 0.007651f
C5456 vdd.n2954 gnd 0.007651f
C5457 vdd.n2955 gnd 0.007651f
C5458 vdd.n2956 gnd 0.007651f
C5459 vdd.n2957 gnd 0.007651f
C5460 vdd.n2959 gnd 0.007651f
C5461 vdd.n2960 gnd 0.007651f
C5462 vdd.n2961 gnd 0.007651f
C5463 vdd.n2962 gnd 0.007651f
C5464 vdd.n2963 gnd 0.007651f
C5465 vdd.n2964 gnd 0.007651f
C5466 vdd.n2966 gnd 0.007651f
C5467 vdd.n2967 gnd 0.007651f
C5468 vdd.n2968 gnd 0.007651f
C5469 vdd.n2969 gnd 0.007651f
C5470 vdd.n2970 gnd 0.007651f
C5471 vdd.n2971 gnd 0.007651f
C5472 vdd.n2973 gnd 0.007651f
C5473 vdd.n2974 gnd 0.018154f
C5474 vdd.n2975 gnd 0.018154f
C5475 vdd.n2976 gnd 0.01695f
C5476 vdd.n2977 gnd 0.007651f
C5477 vdd.n2978 gnd 0.007651f
C5478 vdd.n2979 gnd 0.007651f
C5479 vdd.n2980 gnd 0.007651f
C5480 vdd.n2981 gnd 0.007651f
C5481 vdd.n2982 gnd 0.007651f
C5482 vdd.n2983 gnd 0.781873f
C5483 vdd.n2984 gnd 0.007651f
C5484 vdd.n2985 gnd 0.007651f
C5485 vdd.n2986 gnd 0.007651f
C5486 vdd.n2987 gnd 0.007651f
C5487 vdd.n2988 gnd 0.007651f
C5488 vdd.n2989 gnd 0.48867f
C5489 vdd.n2990 gnd 0.007651f
C5490 vdd.n2991 gnd 0.007651f
C5491 vdd.n2992 gnd 0.007651f
C5492 vdd.n2993 gnd 0.017881f
C5493 vdd.n2994 gnd 0.017222f
C5494 vdd.n2995 gnd 0.018154f
C5495 vdd.n2997 gnd 0.007651f
C5496 vdd.n2998 gnd 0.007651f
C5497 vdd.n2999 gnd 0.005907f
C5498 vdd.n3000 gnd 0.010934f
C5499 vdd.n3001 gnd 0.005569f
C5500 vdd.n3002 gnd 0.007651f
C5501 vdd.n3003 gnd 0.007651f
C5502 vdd.n3005 gnd 0.007651f
C5503 vdd.n3006 gnd 0.007651f
C5504 vdd.n3007 gnd 0.007651f
C5505 vdd.n3008 gnd 0.007651f
C5506 vdd.n3009 gnd 0.007651f
C5507 vdd.n3010 gnd 0.007651f
C5508 vdd.n3012 gnd 0.007651f
C5509 vdd.n3013 gnd 0.007651f
C5510 vdd.n3014 gnd 0.007651f
C5511 vdd.n3015 gnd 0.007651f
C5512 vdd.n3016 gnd 0.007651f
C5513 vdd.n3017 gnd 0.007651f
C5514 vdd.n3019 gnd 0.007651f
C5515 vdd.n3020 gnd 0.007651f
C5516 vdd.n3021 gnd 0.007651f
C5517 vdd.n3022 gnd 0.007651f
C5518 vdd.n3023 gnd 0.007651f
C5519 vdd.n3024 gnd 0.007651f
C5520 vdd.n3026 gnd 0.007651f
C5521 vdd.n3027 gnd 0.007651f
C5522 vdd.n3028 gnd 0.007651f
C5523 vdd.n3030 gnd 0.007651f
C5524 vdd.n3031 gnd 0.007651f
C5525 vdd.n3032 gnd 0.007651f
C5526 vdd.n3033 gnd 0.007651f
C5527 vdd.n3034 gnd 0.007651f
C5528 vdd.n3035 gnd 0.007651f
C5529 vdd.n3037 gnd 0.007651f
C5530 vdd.n3038 gnd 0.007651f
C5531 vdd.n3039 gnd 0.007651f
C5532 vdd.n3040 gnd 0.007651f
C5533 vdd.n3041 gnd 0.007651f
C5534 vdd.n3042 gnd 0.007651f
C5535 vdd.n3044 gnd 0.007651f
C5536 vdd.n3045 gnd 0.007651f
C5537 vdd.n3046 gnd 0.007651f
C5538 vdd.n3047 gnd 0.007651f
C5539 vdd.n3048 gnd 0.007651f
C5540 vdd.n3049 gnd 0.007651f
C5541 vdd.n3051 gnd 0.007651f
C5542 vdd.n3052 gnd 0.007651f
C5543 vdd.n3054 gnd 0.007651f
C5544 vdd.n3055 gnd 0.007651f
C5545 vdd.n3056 gnd 0.018154f
C5546 vdd.n3057 gnd 0.01695f
C5547 vdd.n3058 gnd 0.01695f
C5548 vdd.n3059 gnd 1.12682f
C5549 vdd.n3060 gnd 0.01695f
C5550 vdd.n3061 gnd 0.018154f
C5551 vdd.n3062 gnd 0.017222f
C5552 vdd.n3063 gnd 0.007651f
C5553 vdd.n3064 gnd 0.005907f
C5554 vdd.n3065 gnd 0.007651f
C5555 vdd.n3067 gnd 0.007651f
C5556 vdd.n3068 gnd 0.007651f
C5557 vdd.n3069 gnd 0.007651f
C5558 vdd.n3070 gnd 0.007651f
C5559 vdd.n3071 gnd 0.007651f
C5560 vdd.n3072 gnd 0.007651f
C5561 vdd.n3074 gnd 0.007651f
C5562 vdd.n3075 gnd 0.007651f
C5563 vdd.n3076 gnd 0.007651f
C5564 vdd.n3077 gnd 0.007651f
C5565 vdd.n3078 gnd 0.007651f
C5566 vdd.n3079 gnd 0.007651f
C5567 vdd.n3081 gnd 0.007651f
C5568 vdd.n3082 gnd 0.007651f
C5569 vdd.n3083 gnd 0.007651f
C5570 vdd.n3084 gnd 0.007651f
C5571 vdd.n3085 gnd 0.007651f
C5572 vdd.n3086 gnd 0.007651f
C5573 vdd.n3088 gnd 0.007651f
C5574 vdd.n3089 gnd 0.007651f
C5575 vdd.n3091 gnd 0.007651f
C5576 vdd.n3092 gnd 0.018385f
C5577 vdd.n3093 gnd 0.680937f
C5578 vdd.n3095 gnd 0.004754f
C5579 vdd.n3096 gnd 0.009056f
C5580 vdd.n3097 gnd 0.011251f
C5581 vdd.n3098 gnd 0.011251f
C5582 vdd.n3099 gnd 0.009056f
C5583 vdd.n3100 gnd 0.009056f
C5584 vdd.n3101 gnd 0.011251f
C5585 vdd.n3102 gnd 0.011251f
C5586 vdd.n3103 gnd 0.009056f
C5587 vdd.n3104 gnd 0.009056f
C5588 vdd.n3105 gnd 0.011251f
C5589 vdd.n3106 gnd 0.011251f
C5590 vdd.n3107 gnd 0.009056f
C5591 vdd.n3108 gnd 0.009056f
C5592 vdd.n3109 gnd 0.011251f
C5593 vdd.n3110 gnd 0.011251f
C5594 vdd.n3111 gnd 0.009056f
C5595 vdd.n3112 gnd 0.009056f
C5596 vdd.n3113 gnd 0.011251f
C5597 vdd.n3114 gnd 0.011251f
C5598 vdd.n3115 gnd 0.009056f
C5599 vdd.n3116 gnd 0.009056f
C5600 vdd.n3117 gnd 0.011251f
C5601 vdd.n3118 gnd 0.011251f
C5602 vdd.n3119 gnd 0.009056f
C5603 vdd.n3120 gnd 0.009056f
C5604 vdd.n3121 gnd 0.011251f
C5605 vdd.n3122 gnd 0.011251f
C5606 vdd.n3123 gnd 0.009056f
C5607 vdd.n3124 gnd 0.009056f
C5608 vdd.n3125 gnd 0.011251f
C5609 vdd.n3126 gnd 0.011251f
C5610 vdd.n3127 gnd 0.009056f
C5611 vdd.n3128 gnd 0.009056f
C5612 vdd.n3129 gnd 0.011251f
C5613 vdd.n3130 gnd 0.011251f
C5614 vdd.n3131 gnd 0.009056f
C5615 vdd.n3132 gnd 0.011251f
C5616 vdd.n3133 gnd 0.011251f
C5617 vdd.n3134 gnd 0.009056f
C5618 vdd.n3135 gnd 0.011251f
C5619 vdd.n3136 gnd 0.011251f
C5620 vdd.n3137 gnd 0.011251f
C5621 vdd.n3138 gnd 0.018474f
C5622 vdd.n3139 gnd 0.011251f
C5623 vdd.n3140 gnd 0.011251f
C5624 vdd.n3141 gnd 0.006158f
C5625 vdd.n3142 gnd 0.009056f
C5626 vdd.n3143 gnd 0.011251f
C5627 vdd.n3144 gnd 0.011251f
C5628 vdd.n3145 gnd 0.009056f
C5629 vdd.n3146 gnd 0.009056f
C5630 vdd.n3147 gnd 0.011251f
C5631 vdd.n3148 gnd 0.011251f
C5632 vdd.n3149 gnd 0.009056f
C5633 vdd.n3150 gnd 0.009056f
C5634 vdd.n3151 gnd 0.011251f
C5635 vdd.n3152 gnd 0.011251f
C5636 vdd.n3153 gnd 0.009056f
C5637 vdd.n3154 gnd 0.009056f
C5638 vdd.n3155 gnd 0.011251f
C5639 vdd.n3156 gnd 0.011251f
C5640 vdd.n3157 gnd 0.009056f
C5641 vdd.n3158 gnd 0.009056f
C5642 vdd.n3159 gnd 0.011251f
C5643 vdd.n3160 gnd 0.011251f
C5644 vdd.n3161 gnd 0.009056f
C5645 vdd.n3162 gnd 0.009056f
C5646 vdd.n3163 gnd 0.011251f
C5647 vdd.n3164 gnd 0.011251f
C5648 vdd.n3165 gnd 0.009056f
C5649 vdd.n3166 gnd 0.009056f
C5650 vdd.n3167 gnd 0.011251f
C5651 vdd.n3168 gnd 0.011251f
C5652 vdd.n3169 gnd 0.009056f
C5653 vdd.n3170 gnd 0.009056f
C5654 vdd.n3171 gnd 0.011251f
C5655 vdd.n3172 gnd 0.011251f
C5656 vdd.n3173 gnd 0.009056f
C5657 vdd.n3174 gnd 0.009056f
C5658 vdd.n3175 gnd 0.011251f
C5659 vdd.n3176 gnd 0.011251f
C5660 vdd.n3177 gnd 0.009056f
C5661 vdd.n3178 gnd 0.011251f
C5662 vdd.n3179 gnd 0.011251f
C5663 vdd.n3180 gnd 0.009056f
C5664 vdd.n3181 gnd 0.011251f
C5665 vdd.n3182 gnd 0.011251f
C5666 vdd.n3183 gnd 0.011251f
C5667 vdd.t20 gnd 0.138418f
C5668 vdd.t21 gnd 0.147931f
C5669 vdd.t19 gnd 0.180773f
C5670 vdd.n3184 gnd 0.231725f
C5671 vdd.n3185 gnd 0.194691f
C5672 vdd.n3186 gnd 0.018474f
C5673 vdd.n3187 gnd 0.011251f
C5674 vdd.n3188 gnd 0.011251f
C5675 vdd.n3189 gnd 0.007562f
C5676 vdd.n3190 gnd 0.009056f
C5677 vdd.n3191 gnd 0.011251f
C5678 vdd.n3192 gnd 0.011251f
C5679 vdd.n3193 gnd 0.009056f
C5680 vdd.n3194 gnd 0.009056f
C5681 vdd.n3195 gnd 0.011251f
C5682 vdd.n3196 gnd 0.011251f
C5683 vdd.n3197 gnd 0.009056f
C5684 vdd.n3198 gnd 0.009056f
C5685 vdd.n3199 gnd 0.011251f
C5686 vdd.n3200 gnd 0.011251f
C5687 vdd.n3201 gnd 0.009056f
C5688 vdd.n3202 gnd 0.009056f
C5689 vdd.n3203 gnd 0.011251f
C5690 vdd.n3204 gnd 0.011251f
C5691 vdd.n3205 gnd 0.009056f
C5692 vdd.n3206 gnd 0.009056f
C5693 vdd.n3207 gnd 0.011251f
C5694 vdd.n3208 gnd 0.011251f
C5695 vdd.n3209 gnd 0.009056f
C5696 vdd.n3210 gnd 0.009056f
C5697 vdd.n3211 gnd 0.011251f
C5698 vdd.n3212 gnd 0.011251f
C5699 vdd.n3213 gnd 0.009056f
C5700 vdd.n3214 gnd 0.009056f
C5701 vdd.n3216 gnd 0.680937f
C5702 vdd.n3218 gnd 0.009056f
C5703 vdd.n3219 gnd 0.009056f
C5704 vdd.n3220 gnd 0.007516f
C5705 vdd.n3221 gnd 0.027801f
C5706 vdd.n3223 gnd 8.31315f
C5707 vdd.n3224 gnd 0.027801f
C5708 vdd.n3225 gnd 0.004302f
C5709 vdd.n3226 gnd 0.027801f
C5710 vdd.n3227 gnd 0.027217f
C5711 vdd.n3228 gnd 0.011251f
C5712 vdd.n3229 gnd 0.009056f
C5713 vdd.n3230 gnd 0.011251f
C5714 vdd.n3231 gnd 0.695637f
C5715 vdd.n3232 gnd 0.011251f
C5716 vdd.n3233 gnd 0.009056f
C5717 vdd.n3234 gnd 0.011251f
C5718 vdd.n3235 gnd 0.011251f
C5719 vdd.n3236 gnd 0.011251f
C5720 vdd.n3237 gnd 0.009056f
C5721 vdd.n3238 gnd 0.011251f
C5722 vdd.n3239 gnd 1.14981f
C5723 vdd.n3240 gnd 0.011251f
C5724 vdd.n3241 gnd 0.009056f
C5725 vdd.n3242 gnd 0.011251f
C5726 vdd.n3243 gnd 0.011251f
C5727 vdd.n3244 gnd 0.011251f
C5728 vdd.n3245 gnd 0.009056f
C5729 vdd.n3246 gnd 0.011251f
C5730 vdd.n3247 gnd 0.741629f
C5731 vdd.n3248 gnd 0.787622f
C5732 vdd.n3249 gnd 0.011251f
C5733 vdd.n3250 gnd 0.009056f
C5734 vdd.n3251 gnd 0.011251f
C5735 vdd.n3252 gnd 0.011251f
C5736 vdd.n3253 gnd 0.011251f
C5737 vdd.n3254 gnd 0.009056f
C5738 vdd.n3255 gnd 0.011251f
C5739 vdd.n3256 gnd 0.954345f
C5740 vdd.n3257 gnd 0.011251f
C5741 vdd.n3258 gnd 0.009056f
C5742 vdd.n3259 gnd 0.011251f
C5743 vdd.n3260 gnd 0.011251f
C5744 vdd.n3261 gnd 0.011251f
C5745 vdd.n3262 gnd 0.009056f
C5746 vdd.n3263 gnd 0.011251f
C5747 vdd.t147 gnd 0.574906f
C5748 vdd.n3264 gnd 0.925599f
C5749 vdd.n3265 gnd 0.011251f
C5750 vdd.n3266 gnd 0.009056f
C5751 vdd.n3267 gnd 0.011251f
C5752 vdd.n3268 gnd 0.011251f
C5753 vdd.n3269 gnd 0.011251f
C5754 vdd.n3270 gnd 0.009056f
C5755 vdd.n3271 gnd 0.011251f
C5756 vdd.n3272 gnd 0.730131f
C5757 vdd.n3273 gnd 0.011251f
C5758 vdd.n3274 gnd 0.009056f
C5759 vdd.n3275 gnd 0.011251f
C5760 vdd.n3276 gnd 0.011251f
C5761 vdd.n3277 gnd 0.011251f
C5762 vdd.n3278 gnd 0.009056f
C5763 vdd.n3279 gnd 0.011251f
C5764 vdd.n3280 gnd 0.914101f
C5765 vdd.n3281 gnd 0.61515f
C5766 vdd.n3282 gnd 0.011251f
C5767 vdd.n3283 gnd 0.009056f
C5768 vdd.n3284 gnd 0.011251f
C5769 vdd.n3285 gnd 0.011251f
C5770 vdd.n3286 gnd 0.011251f
C5771 vdd.n3287 gnd 0.009056f
C5772 vdd.n3288 gnd 0.011251f
C5773 vdd.n3289 gnd 0.810618f
C5774 vdd.n3290 gnd 0.011251f
C5775 vdd.n3291 gnd 0.009056f
C5776 vdd.n3292 gnd 0.011251f
C5777 vdd.n3293 gnd 0.011251f
C5778 vdd.n3294 gnd 0.011251f
C5779 vdd.n3295 gnd 0.011251f
C5780 vdd.n3296 gnd 0.011251f
C5781 vdd.n3297 gnd 0.009056f
C5782 vdd.n3298 gnd 0.009056f
C5783 vdd.n3299 gnd 0.011251f
C5784 vdd.t192 gnd 0.574906f
C5785 vdd.n3300 gnd 0.954345f
C5786 vdd.n3301 gnd 0.011251f
C5787 vdd.n3302 gnd 0.009056f
C5788 vdd.n3303 gnd 0.011251f
C5789 vdd.n3304 gnd 0.011251f
C5790 vdd.n3305 gnd 0.011251f
C5791 vdd.n3306 gnd 0.009056f
C5792 vdd.n3307 gnd 0.011251f
C5793 vdd.n3308 gnd 0.902603f
C5794 vdd.n3309 gnd 0.011251f
C5795 vdd.n3310 gnd 0.011251f
C5796 vdd.n3311 gnd 0.009056f
C5797 vdd.n3312 gnd 0.009056f
C5798 vdd.n3313 gnd 0.011251f
C5799 vdd.n3314 gnd 0.011251f
C5800 vdd.n3315 gnd 0.011251f
C5801 vdd.n3316 gnd 0.009056f
C5802 vdd.n3317 gnd 0.011251f
C5803 vdd.n3318 gnd 0.009056f
C5804 vdd.n3319 gnd 0.009056f
C5805 vdd.n3320 gnd 0.011251f
C5806 vdd.n3321 gnd 0.011251f
C5807 vdd.n3322 gnd 0.011251f
C5808 vdd.n3323 gnd 0.009056f
C5809 vdd.n3324 gnd 0.011251f
C5810 vdd.n3325 gnd 0.009056f
C5811 vdd.n3326 gnd 0.009056f
C5812 vdd.n3327 gnd 0.011251f
C5813 vdd.n3328 gnd 0.011251f
C5814 vdd.n3329 gnd 0.011251f
C5815 vdd.n3330 gnd 0.009056f
C5816 vdd.n3331 gnd 0.954345f
C5817 vdd.n3332 gnd 0.011251f
C5818 vdd.n3333 gnd 0.009056f
C5819 vdd.n3334 gnd 0.009056f
C5820 vdd.n3335 gnd 0.011251f
C5821 vdd.n3336 gnd 0.011251f
C5822 vdd.n3337 gnd 0.011251f
C5823 vdd.n3338 gnd 0.009056f
C5824 vdd.n3339 gnd 0.011251f
C5825 vdd.n3340 gnd 0.009056f
C5826 vdd.n3341 gnd 0.009056f
C5827 vdd.n3342 gnd 0.011251f
C5828 vdd.n3343 gnd 0.011251f
C5829 vdd.n3344 gnd 0.011251f
C5830 vdd.n3345 gnd 0.009056f
C5831 vdd.n3346 gnd 0.011251f
C5832 vdd.n3347 gnd 0.009056f
C5833 vdd.n3348 gnd 0.007516f
C5834 vdd.n3349 gnd 0.027217f
C5835 vdd.n3350 gnd 0.027801f
C5836 vdd.n3351 gnd 0.004302f
C5837 vdd.n3352 gnd 0.027801f
C5838 vdd.n3354 gnd 2.72506f
C5839 vdd.n3355 gnd 1.69597f
C5840 vdd.n3356 gnd 0.027217f
C5841 vdd.n3357 gnd 0.007516f
C5842 vdd.n3358 gnd 0.009056f
C5843 vdd.n3359 gnd 0.009056f
C5844 vdd.n3360 gnd 0.011251f
C5845 vdd.n3361 gnd 1.14981f
C5846 vdd.n3362 gnd 1.14981f
C5847 vdd.n3363 gnd 1.05208f
C5848 vdd.n3364 gnd 0.011251f
C5849 vdd.n3365 gnd 0.009056f
C5850 vdd.n3366 gnd 0.009056f
C5851 vdd.n3367 gnd 0.009056f
C5852 vdd.n3368 gnd 0.011251f
C5853 vdd.n3369 gnd 0.85661f
C5854 vdd.t211 gnd 0.574906f
C5855 vdd.n3370 gnd 0.868109f
C5856 vdd.n3371 gnd 0.661142f
C5857 vdd.n3372 gnd 0.011251f
C5858 vdd.n3373 gnd 0.009056f
C5859 vdd.n3374 gnd 0.009056f
C5860 vdd.n3375 gnd 0.009056f
C5861 vdd.n3376 gnd 0.011251f
C5862 vdd.n3377 gnd 0.684139f
C5863 vdd.n3378 gnd 0.845112f
C5864 vdd.t163 gnd 0.574906f
C5865 vdd.n3379 gnd 0.879607f
C5866 vdd.n3380 gnd 0.011251f
C5867 vdd.n3381 gnd 0.009056f
C5868 vdd.n3382 gnd 0.009056f
C5869 vdd.n3383 gnd 0.009056f
C5870 vdd.n3384 gnd 0.011251f
C5871 vdd.n3385 gnd 0.954345f
C5872 vdd.t188 gnd 0.574906f
C5873 vdd.n3386 gnd 0.695637f
C5874 vdd.n3387 gnd 0.833614f
C5875 vdd.n3388 gnd 0.011251f
C5876 vdd.n3389 gnd 0.009056f
C5877 vdd.n3390 gnd 0.009056f
C5878 vdd.n3391 gnd 0.009056f
C5879 vdd.n3392 gnd 0.011251f
C5880 vdd.n3393 gnd 0.638146f
C5881 vdd.t158 gnd 0.574906f
C5882 vdd.n3394 gnd 0.954345f
C5883 vdd.t185 gnd 0.574906f
C5884 vdd.n3395 gnd 0.707135f
C5885 vdd.n3396 gnd 0.011251f
C5886 vdd.n3397 gnd 0.009056f
C5887 vdd.n3398 gnd 0.008647f
C5888 vdd.n3399 gnd 0.663635f
C5889 vdd.n3400 gnd 2.87708f
C5890 a_n7636_8799.n0 gnd 0.789434f
C5891 a_n7636_8799.n1 gnd 3.25763f
C5892 a_n7636_8799.n2 gnd 3.09896f
C5893 a_n7636_8799.n3 gnd 1.53168f
C5894 a_n7636_8799.n4 gnd 0.207903f
C5895 a_n7636_8799.n5 gnd 0.285477f
C5896 a_n7636_8799.n6 gnd 0.207903f
C5897 a_n7636_8799.n7 gnd 0.207903f
C5898 a_n7636_8799.n8 gnd 0.207903f
C5899 a_n7636_8799.n9 gnd 0.207903f
C5900 a_n7636_8799.n10 gnd 0.207903f
C5901 a_n7636_8799.n11 gnd 0.216181f
C5902 a_n7636_8799.n12 gnd 0.207903f
C5903 a_n7636_8799.n13 gnd 0.285477f
C5904 a_n7636_8799.n14 gnd 0.207903f
C5905 a_n7636_8799.n15 gnd 0.207903f
C5906 a_n7636_8799.n16 gnd 0.207903f
C5907 a_n7636_8799.n17 gnd 0.207903f
C5908 a_n7636_8799.n18 gnd 0.207903f
C5909 a_n7636_8799.n19 gnd 0.216181f
C5910 a_n7636_8799.n20 gnd 0.207903f
C5911 a_n7636_8799.n21 gnd 0.450615f
C5912 a_n7636_8799.n22 gnd 0.207903f
C5913 a_n7636_8799.n23 gnd 0.207903f
C5914 a_n7636_8799.n24 gnd 0.207903f
C5915 a_n7636_8799.n25 gnd 0.207903f
C5916 a_n7636_8799.n26 gnd 0.207903f
C5917 a_n7636_8799.n27 gnd 0.216181f
C5918 a_n7636_8799.n28 gnd 0.207903f
C5919 a_n7636_8799.n29 gnd 0.320132f
C5920 a_n7636_8799.n30 gnd 0.207903f
C5921 a_n7636_8799.n31 gnd 0.207903f
C5922 a_n7636_8799.n32 gnd 0.207903f
C5923 a_n7636_8799.n33 gnd 0.207903f
C5924 a_n7636_8799.n34 gnd 0.207903f
C5925 a_n7636_8799.n35 gnd 0.181526f
C5926 a_n7636_8799.n36 gnd 0.207903f
C5927 a_n7636_8799.n37 gnd 0.320132f
C5928 a_n7636_8799.n38 gnd 0.207903f
C5929 a_n7636_8799.n39 gnd 0.207903f
C5930 a_n7636_8799.n40 gnd 0.207903f
C5931 a_n7636_8799.n41 gnd 0.207903f
C5932 a_n7636_8799.n42 gnd 0.207903f
C5933 a_n7636_8799.n43 gnd 0.181526f
C5934 a_n7636_8799.n44 gnd 0.207903f
C5935 a_n7636_8799.n45 gnd 0.320132f
C5936 a_n7636_8799.n46 gnd 0.207903f
C5937 a_n7636_8799.n47 gnd 0.207903f
C5938 a_n7636_8799.n48 gnd 0.207903f
C5939 a_n7636_8799.n49 gnd 0.207903f
C5940 a_n7636_8799.n50 gnd 0.207903f
C5941 a_n7636_8799.n51 gnd 0.346664f
C5942 a_n7636_8799.n52 gnd 2.83385f
C5943 a_n7636_8799.n53 gnd 3.97496f
C5944 a_n7636_8799.n54 gnd 0.250295f
C5945 a_n7636_8799.n55 gnd 0.003659f
C5946 a_n7636_8799.n56 gnd 0.009646f
C5947 a_n7636_8799.n57 gnd 0.010539f
C5948 a_n7636_8799.n58 gnd 0.005569f
C5949 a_n7636_8799.n60 gnd 0.004673f
C5950 a_n7636_8799.n61 gnd 0.010106f
C5951 a_n7636_8799.n62 gnd 0.010106f
C5952 a_n7636_8799.n63 gnd 0.004673f
C5953 a_n7636_8799.n65 gnd 0.005569f
C5954 a_n7636_8799.n66 gnd 0.010539f
C5955 a_n7636_8799.n67 gnd 0.009646f
C5956 a_n7636_8799.n68 gnd 0.003659f
C5957 a_n7636_8799.n69 gnd 0.250295f
C5958 a_n7636_8799.n70 gnd 0.003659f
C5959 a_n7636_8799.n71 gnd 0.009646f
C5960 a_n7636_8799.n72 gnd 0.010539f
C5961 a_n7636_8799.n73 gnd 0.005569f
C5962 a_n7636_8799.n75 gnd 0.004673f
C5963 a_n7636_8799.n76 gnd 0.010106f
C5964 a_n7636_8799.n77 gnd 0.010106f
C5965 a_n7636_8799.n78 gnd 0.004673f
C5966 a_n7636_8799.n80 gnd 0.005569f
C5967 a_n7636_8799.n81 gnd 0.010539f
C5968 a_n7636_8799.n82 gnd 0.009646f
C5969 a_n7636_8799.n83 gnd 0.003659f
C5970 a_n7636_8799.n84 gnd 0.250295f
C5971 a_n7636_8799.n85 gnd 0.003659f
C5972 a_n7636_8799.n86 gnd 0.009646f
C5973 a_n7636_8799.n87 gnd 0.010539f
C5974 a_n7636_8799.n88 gnd 0.005569f
C5975 a_n7636_8799.n90 gnd 0.004673f
C5976 a_n7636_8799.n91 gnd 0.010106f
C5977 a_n7636_8799.n92 gnd 0.010106f
C5978 a_n7636_8799.n93 gnd 0.004673f
C5979 a_n7636_8799.n95 gnd 0.005569f
C5980 a_n7636_8799.n96 gnd 0.010539f
C5981 a_n7636_8799.n97 gnd 0.009646f
C5982 a_n7636_8799.n98 gnd 0.003659f
C5983 a_n7636_8799.n99 gnd 0.003659f
C5984 a_n7636_8799.n100 gnd 0.009646f
C5985 a_n7636_8799.n101 gnd 0.010539f
C5986 a_n7636_8799.n102 gnd 0.005569f
C5987 a_n7636_8799.n104 gnd 0.004673f
C5988 a_n7636_8799.n105 gnd 0.010106f
C5989 a_n7636_8799.n106 gnd 0.010106f
C5990 a_n7636_8799.n107 gnd 0.004673f
C5991 a_n7636_8799.n109 gnd 0.005569f
C5992 a_n7636_8799.n110 gnd 0.010539f
C5993 a_n7636_8799.n111 gnd 0.009646f
C5994 a_n7636_8799.n112 gnd 0.003659f
C5995 a_n7636_8799.n113 gnd 0.250295f
C5996 a_n7636_8799.n114 gnd 0.003659f
C5997 a_n7636_8799.n115 gnd 0.009646f
C5998 a_n7636_8799.n116 gnd 0.010539f
C5999 a_n7636_8799.n117 gnd 0.005569f
C6000 a_n7636_8799.n119 gnd 0.004673f
C6001 a_n7636_8799.n120 gnd 0.010106f
C6002 a_n7636_8799.n121 gnd 0.010106f
C6003 a_n7636_8799.n122 gnd 0.004673f
C6004 a_n7636_8799.n124 gnd 0.005569f
C6005 a_n7636_8799.n125 gnd 0.010539f
C6006 a_n7636_8799.n126 gnd 0.009646f
C6007 a_n7636_8799.n127 gnd 0.003659f
C6008 a_n7636_8799.n128 gnd 0.250295f
C6009 a_n7636_8799.n129 gnd 0.003659f
C6010 a_n7636_8799.n130 gnd 0.009646f
C6011 a_n7636_8799.n131 gnd 0.010539f
C6012 a_n7636_8799.n132 gnd 0.005569f
C6013 a_n7636_8799.n134 gnd 0.004673f
C6014 a_n7636_8799.n135 gnd 0.010106f
C6015 a_n7636_8799.n136 gnd 0.010106f
C6016 a_n7636_8799.n137 gnd 0.004673f
C6017 a_n7636_8799.n139 gnd 0.005569f
C6018 a_n7636_8799.n140 gnd 0.010539f
C6019 a_n7636_8799.n141 gnd 0.009646f
C6020 a_n7636_8799.n142 gnd 0.003659f
C6021 a_n7636_8799.n143 gnd 0.250295f
C6022 a_n7636_8799.t17 gnd 0.144203f
C6023 a_n7636_8799.t24 gnd 0.144203f
C6024 a_n7636_8799.t22 gnd 0.144203f
C6025 a_n7636_8799.n144 gnd 1.13736f
C6026 a_n7636_8799.t27 gnd 0.144203f
C6027 a_n7636_8799.t30 gnd 0.144203f
C6028 a_n7636_8799.n145 gnd 1.13548f
C6029 a_n7636_8799.t25 gnd 0.144203f
C6030 a_n7636_8799.t12 gnd 0.144203f
C6031 a_n7636_8799.n146 gnd 1.13548f
C6032 a_n7636_8799.t6 gnd 0.112158f
C6033 a_n7636_8799.t9 gnd 0.112158f
C6034 a_n7636_8799.n147 gnd 0.993274f
C6035 a_n7636_8799.t13 gnd 0.112158f
C6036 a_n7636_8799.t8 gnd 0.112158f
C6037 a_n7636_8799.n148 gnd 0.99107f
C6038 a_n7636_8799.t14 gnd 0.112158f
C6039 a_n7636_8799.t10 gnd 0.112158f
C6040 a_n7636_8799.n149 gnd 0.99107f
C6041 a_n7636_8799.t2 gnd 0.112158f
C6042 a_n7636_8799.t23 gnd 0.112158f
C6043 a_n7636_8799.n150 gnd 0.993273f
C6044 a_n7636_8799.t11 gnd 0.112158f
C6045 a_n7636_8799.t18 gnd 0.112158f
C6046 a_n7636_8799.n151 gnd 0.991069f
C6047 a_n7636_8799.t26 gnd 0.112158f
C6048 a_n7636_8799.t15 gnd 0.112158f
C6049 a_n7636_8799.n152 gnd 0.991069f
C6050 a_n7636_8799.t16 gnd 0.112158f
C6051 a_n7636_8799.t21 gnd 0.112158f
C6052 a_n7636_8799.n153 gnd 0.993273f
C6053 a_n7636_8799.t4 gnd 0.112158f
C6054 a_n7636_8799.t1 gnd 0.112158f
C6055 a_n7636_8799.n154 gnd 0.991069f
C6056 a_n7636_8799.t3 gnd 0.112158f
C6057 a_n7636_8799.t7 gnd 0.112158f
C6058 a_n7636_8799.n155 gnd 0.99107f
C6059 a_n7636_8799.t0 gnd 0.112158f
C6060 a_n7636_8799.t29 gnd 0.112158f
C6061 a_n7636_8799.n156 gnd 0.99107f
C6062 a_n7636_8799.t128 gnd 0.597935f
C6063 a_n7636_8799.n157 gnd 0.269198f
C6064 a_n7636_8799.t44 gnd 0.597935f
C6065 a_n7636_8799.t65 gnd 0.597935f
C6066 a_n7636_8799.n158 gnd 0.271126f
C6067 a_n7636_8799.t88 gnd 0.597935f
C6068 a_n7636_8799.t107 gnd 0.597935f
C6069 a_n7636_8799.n159 gnd 0.264325f
C6070 a_n7636_8799.t67 gnd 0.597935f
C6071 a_n7636_8799.t79 gnd 0.597935f
C6072 a_n7636_8799.n160 gnd 0.268305f
C6073 a_n7636_8799.t112 gnd 0.597935f
C6074 a_n7636_8799.t133 gnd 0.597935f
C6075 a_n7636_8799.t132 gnd 0.609251f
C6076 a_n7636_8799.n161 gnd 0.250658f
C6077 a_n7636_8799.n162 gnd 0.271499f
C6078 a_n7636_8799.t83 gnd 0.597935f
C6079 a_n7636_8799.n163 gnd 0.269198f
C6080 a_n7636_8799.n164 gnd 0.264966f
C6081 a_n7636_8799.t129 gnd 0.597935f
C6082 a_n7636_8799.n165 gnd 0.263684f
C6083 a_n7636_8799.t80 gnd 0.597935f
C6084 a_n7636_8799.n166 gnd 0.270871f
C6085 a_n7636_8799.t110 gnd 0.597935f
C6086 a_n7636_8799.n167 gnd 0.271126f
C6087 a_n7636_8799.n168 gnd 0.268737f
C6088 a_n7636_8799.t68 gnd 0.597935f
C6089 a_n7636_8799.n169 gnd 0.264325f
C6090 a_n7636_8799.t32 gnd 0.597935f
C6091 a_n7636_8799.n170 gnd 0.268737f
C6092 a_n7636_8799.n171 gnd 0.270871f
C6093 a_n7636_8799.t131 gnd 0.597935f
C6094 a_n7636_8799.n172 gnd 0.268305f
C6095 a_n7636_8799.n173 gnd 0.263684f
C6096 a_n7636_8799.t62 gnd 0.597935f
C6097 a_n7636_8799.n174 gnd 0.264966f
C6098 a_n7636_8799.t41 gnd 0.597935f
C6099 a_n7636_8799.n175 gnd 0.271499f
C6100 a_n7636_8799.t42 gnd 0.609241f
C6101 a_n7636_8799.t141 gnd 0.597935f
C6102 a_n7636_8799.n176 gnd 0.269198f
C6103 a_n7636_8799.t59 gnd 0.597935f
C6104 a_n7636_8799.t74 gnd 0.597935f
C6105 a_n7636_8799.n177 gnd 0.271126f
C6106 a_n7636_8799.t101 gnd 0.597935f
C6107 a_n7636_8799.t119 gnd 0.597935f
C6108 a_n7636_8799.n178 gnd 0.264325f
C6109 a_n7636_8799.t77 gnd 0.597935f
C6110 a_n7636_8799.t89 gnd 0.597935f
C6111 a_n7636_8799.n179 gnd 0.268305f
C6112 a_n7636_8799.t125 gnd 0.597935f
C6113 a_n7636_8799.t149 gnd 0.597935f
C6114 a_n7636_8799.t146 gnd 0.609251f
C6115 a_n7636_8799.n180 gnd 0.250658f
C6116 a_n7636_8799.n181 gnd 0.271499f
C6117 a_n7636_8799.t93 gnd 0.597935f
C6118 a_n7636_8799.n182 gnd 0.269198f
C6119 a_n7636_8799.n183 gnd 0.264966f
C6120 a_n7636_8799.t143 gnd 0.597935f
C6121 a_n7636_8799.n184 gnd 0.263684f
C6122 a_n7636_8799.t90 gnd 0.597935f
C6123 a_n7636_8799.n185 gnd 0.270871f
C6124 a_n7636_8799.t123 gnd 0.597935f
C6125 a_n7636_8799.n186 gnd 0.271126f
C6126 a_n7636_8799.n187 gnd 0.268737f
C6127 a_n7636_8799.t78 gnd 0.597935f
C6128 a_n7636_8799.n188 gnd 0.264325f
C6129 a_n7636_8799.t43 gnd 0.597935f
C6130 a_n7636_8799.n189 gnd 0.268737f
C6131 a_n7636_8799.n190 gnd 0.270871f
C6132 a_n7636_8799.t147 gnd 0.597935f
C6133 a_n7636_8799.n191 gnd 0.268305f
C6134 a_n7636_8799.n192 gnd 0.263684f
C6135 a_n7636_8799.t73 gnd 0.597935f
C6136 a_n7636_8799.n193 gnd 0.264966f
C6137 a_n7636_8799.t53 gnd 0.597935f
C6138 a_n7636_8799.n194 gnd 0.271499f
C6139 a_n7636_8799.t55 gnd 0.609241f
C6140 a_n7636_8799.n195 gnd 0.898912f
C6141 a_n7636_8799.t96 gnd 0.597935f
C6142 a_n7636_8799.n196 gnd 0.269198f
C6143 a_n7636_8799.t120 gnd 0.597935f
C6144 a_n7636_8799.t38 gnd 0.597935f
C6145 a_n7636_8799.n197 gnd 0.271126f
C6146 a_n7636_8799.t103 gnd 0.597935f
C6147 a_n7636_8799.t142 gnd 0.597935f
C6148 a_n7636_8799.n198 gnd 0.264325f
C6149 a_n7636_8799.t137 gnd 0.597935f
C6150 a_n7636_8799.t50 gnd 0.597935f
C6151 a_n7636_8799.n199 gnd 0.268305f
C6152 a_n7636_8799.t75 gnd 0.597935f
C6153 a_n7636_8799.t86 gnd 0.597935f
C6154 a_n7636_8799.t108 gnd 0.609251f
C6155 a_n7636_8799.n200 gnd 0.250658f
C6156 a_n7636_8799.n201 gnd 0.271499f
C6157 a_n7636_8799.t124 gnd 0.597935f
C6158 a_n7636_8799.n202 gnd 0.269198f
C6159 a_n7636_8799.n203 gnd 0.264966f
C6160 a_n7636_8799.t134 gnd 0.597935f
C6161 a_n7636_8799.n204 gnd 0.263684f
C6162 a_n7636_8799.t33 gnd 0.597935f
C6163 a_n7636_8799.n205 gnd 0.270871f
C6164 a_n7636_8799.t94 gnd 0.597935f
C6165 a_n7636_8799.n206 gnd 0.271126f
C6166 a_n7636_8799.n207 gnd 0.268737f
C6167 a_n7636_8799.t111 gnd 0.597935f
C6168 a_n7636_8799.n208 gnd 0.264325f
C6169 a_n7636_8799.t87 gnd 0.597935f
C6170 a_n7636_8799.n209 gnd 0.268737f
C6171 a_n7636_8799.n210 gnd 0.270871f
C6172 a_n7636_8799.t57 gnd 0.597935f
C6173 a_n7636_8799.n211 gnd 0.268305f
C6174 a_n7636_8799.n212 gnd 0.263684f
C6175 a_n7636_8799.t66 gnd 0.597935f
C6176 a_n7636_8799.n213 gnd 0.264966f
C6177 a_n7636_8799.t46 gnd 0.597935f
C6178 a_n7636_8799.n214 gnd 0.271499f
C6179 a_n7636_8799.t148 gnd 0.609241f
C6180 a_n7636_8799.n215 gnd 1.45959f
C6181 a_n7636_8799.t82 gnd 0.609241f
C6182 a_n7636_8799.t81 gnd 0.597935f
C6183 a_n7636_8799.t54 gnd 0.597935f
C6184 a_n7636_8799.n216 gnd 0.269198f
C6185 a_n7636_8799.t130 gnd 0.597935f
C6186 a_n7636_8799.t85 gnd 0.597935f
C6187 a_n7636_8799.t61 gnd 0.597935f
C6188 a_n7636_8799.n217 gnd 0.268305f
C6189 a_n7636_8799.t136 gnd 0.597935f
C6190 a_n7636_8799.t102 gnd 0.597935f
C6191 a_n7636_8799.t100 gnd 0.597935f
C6192 a_n7636_8799.n218 gnd 0.268737f
C6193 a_n7636_8799.t35 gnd 0.597935f
C6194 a_n7636_8799.t106 gnd 0.597935f
C6195 a_n7636_8799.t105 gnd 0.597935f
C6196 a_n7636_8799.n219 gnd 0.268737f
C6197 a_n7636_8799.t37 gnd 0.597935f
C6198 a_n7636_8799.t36 gnd 0.597935f
C6199 a_n7636_8799.t122 gnd 0.597935f
C6200 a_n7636_8799.n220 gnd 0.268305f
C6201 a_n7636_8799.t56 gnd 0.597935f
C6202 a_n7636_8799.t40 gnd 0.597935f
C6203 a_n7636_8799.t126 gnd 0.597935f
C6204 a_n7636_8799.n221 gnd 0.269198f
C6205 a_n7636_8799.t60 gnd 0.609251f
C6206 a_n7636_8799.n222 gnd 0.250658f
C6207 a_n7636_8799.t84 gnd 0.597935f
C6208 a_n7636_8799.n223 gnd 0.271499f
C6209 a_n7636_8799.n224 gnd 0.264966f
C6210 a_n7636_8799.n225 gnd 0.263684f
C6211 a_n7636_8799.n226 gnd 0.270871f
C6212 a_n7636_8799.n227 gnd 0.271126f
C6213 a_n7636_8799.n228 gnd 0.264325f
C6214 a_n7636_8799.n229 gnd 0.264325f
C6215 a_n7636_8799.n230 gnd 0.271126f
C6216 a_n7636_8799.n231 gnd 0.270871f
C6217 a_n7636_8799.n232 gnd 0.263684f
C6218 a_n7636_8799.n233 gnd 0.264966f
C6219 a_n7636_8799.n234 gnd 0.271499f
C6220 a_n7636_8799.t92 gnd 0.609241f
C6221 a_n7636_8799.t91 gnd 0.597935f
C6222 a_n7636_8799.t69 gnd 0.597935f
C6223 a_n7636_8799.n235 gnd 0.269198f
C6224 a_n7636_8799.t145 gnd 0.597935f
C6225 a_n7636_8799.t98 gnd 0.597935f
C6226 a_n7636_8799.t71 gnd 0.597935f
C6227 a_n7636_8799.n236 gnd 0.268305f
C6228 a_n7636_8799.t151 gnd 0.597935f
C6229 a_n7636_8799.t115 gnd 0.597935f
C6230 a_n7636_8799.t114 gnd 0.597935f
C6231 a_n7636_8799.n237 gnd 0.268737f
C6232 a_n7636_8799.t45 gnd 0.597935f
C6233 a_n7636_8799.t118 gnd 0.597935f
C6234 a_n7636_8799.t117 gnd 0.597935f
C6235 a_n7636_8799.n238 gnd 0.268737f
C6236 a_n7636_8799.t49 gnd 0.597935f
C6237 a_n7636_8799.t48 gnd 0.597935f
C6238 a_n7636_8799.t139 gnd 0.597935f
C6239 a_n7636_8799.n239 gnd 0.268305f
C6240 a_n7636_8799.t70 gnd 0.597935f
C6241 a_n7636_8799.t52 gnd 0.597935f
C6242 a_n7636_8799.t140 gnd 0.597935f
C6243 a_n7636_8799.n240 gnd 0.269198f
C6244 a_n7636_8799.t72 gnd 0.609251f
C6245 a_n7636_8799.n241 gnd 0.250658f
C6246 a_n7636_8799.t99 gnd 0.597935f
C6247 a_n7636_8799.n242 gnd 0.271499f
C6248 a_n7636_8799.n243 gnd 0.264966f
C6249 a_n7636_8799.n244 gnd 0.263684f
C6250 a_n7636_8799.n245 gnd 0.270871f
C6251 a_n7636_8799.n246 gnd 0.271126f
C6252 a_n7636_8799.n247 gnd 0.264325f
C6253 a_n7636_8799.n248 gnd 0.264325f
C6254 a_n7636_8799.n249 gnd 0.271126f
C6255 a_n7636_8799.n250 gnd 0.270871f
C6256 a_n7636_8799.n251 gnd 0.263684f
C6257 a_n7636_8799.n252 gnd 0.264966f
C6258 a_n7636_8799.n253 gnd 0.271499f
C6259 a_n7636_8799.n254 gnd 0.898912f
C6260 a_n7636_8799.t150 gnd 0.609241f
C6261 a_n7636_8799.t47 gnd 0.597935f
C6262 a_n7636_8799.t97 gnd 0.597935f
C6263 a_n7636_8799.n255 gnd 0.269198f
C6264 a_n7636_8799.t34 gnd 0.597935f
C6265 a_n7636_8799.t121 gnd 0.597935f
C6266 a_n7636_8799.t58 gnd 0.597935f
C6267 a_n7636_8799.n256 gnd 0.268305f
C6268 a_n7636_8799.t104 gnd 0.597935f
C6269 a_n7636_8799.t39 gnd 0.597935f
C6270 a_n7636_8799.t64 gnd 0.597935f
C6271 a_n7636_8799.n257 gnd 0.268737f
C6272 a_n7636_8799.t144 gnd 0.597935f
C6273 a_n7636_8799.t113 gnd 0.597935f
C6274 a_n7636_8799.t138 gnd 0.597935f
C6275 a_n7636_8799.n258 gnd 0.268737f
C6276 a_n7636_8799.t95 gnd 0.597935f
C6277 a_n7636_8799.t116 gnd 0.597935f
C6278 a_n7636_8799.t51 gnd 0.597935f
C6279 a_n7636_8799.n259 gnd 0.268305f
C6280 a_n7636_8799.t135 gnd 0.597935f
C6281 a_n7636_8799.t76 gnd 0.597935f
C6282 a_n7636_8799.t127 gnd 0.597935f
C6283 a_n7636_8799.n260 gnd 0.269198f
C6284 a_n7636_8799.t109 gnd 0.609251f
C6285 a_n7636_8799.n261 gnd 0.250658f
C6286 a_n7636_8799.t63 gnd 0.597935f
C6287 a_n7636_8799.n262 gnd 0.271499f
C6288 a_n7636_8799.n263 gnd 0.264966f
C6289 a_n7636_8799.n264 gnd 0.263684f
C6290 a_n7636_8799.n265 gnd 0.270871f
C6291 a_n7636_8799.n266 gnd 0.271126f
C6292 a_n7636_8799.n267 gnd 0.264325f
C6293 a_n7636_8799.n268 gnd 0.264325f
C6294 a_n7636_8799.n269 gnd 0.271126f
C6295 a_n7636_8799.n270 gnd 0.270871f
C6296 a_n7636_8799.n271 gnd 0.263684f
C6297 a_n7636_8799.n272 gnd 0.264966f
C6298 a_n7636_8799.n273 gnd 0.271499f
C6299 a_n7636_8799.n274 gnd 1.133f
C6300 a_n7636_8799.n275 gnd 12.2459f
C6301 a_n7636_8799.n276 gnd 4.37601f
C6302 a_n7636_8799.n277 gnd 5.69264f
C6303 a_n7636_8799.t19 gnd 0.144203f
C6304 a_n7636_8799.t20 gnd 0.144203f
C6305 a_n7636_8799.n278 gnd 1.13548f
C6306 a_n7636_8799.t31 gnd 0.144203f
C6307 a_n7636_8799.t28 gnd 0.144203f
C6308 a_n7636_8799.n279 gnd 1.13548f
C6309 a_n7636_8799.n280 gnd 1.13736f
C6310 a_n7636_8799.t5 gnd 0.144203f
.ends

