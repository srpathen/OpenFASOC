* NGSPICE file created from opamp619.ext - technology: sky130A

.subckt opamp619 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 gnd.t351 commonsourceibias.t6 commonsourceibias.t7 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 CSoutput.t95 a_n7636_8799.t32 vdd.t263 vdd.t218 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X2 a_n2140_13878.t15 a_n2318_13878.t7 a_n2318_13878.t8 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 a_n2140_13878.t23 a_n2318_13878.t48 vdd.t16 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 CSoutput.t191 commonsourceibias.t64 gnd.t350 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X5 vdd.t262 a_n7636_8799.t33 CSoutput.t94 vdd.t213 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 commonsourceibias.t5 commonsourceibias.t4 gnd.t349 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 gnd.t348 commonsourceibias.t65 CSoutput.t190 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 a_n7636_8799.t5 plus.t5 a_n3827_n3924.t29 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X9 gnd.t347 commonsourceibias.t2 commonsourceibias.t3 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 a_n3827_n3924.t0 diffpairibias.t20 gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X11 CSoutput.t93 a_n7636_8799.t34 vdd.t261 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X12 minus.t4 gnd.t189 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X13 gnd.t346 commonsourceibias.t0 commonsourceibias.t1 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X14 vdd.t124 vdd.t122 vdd.t123 vdd.t83 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X15 a_n2318_8322.t23 a_n2318_13878.t49 a_n7636_8799.t8 vdd.t5 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X16 commonsourceibias.t59 commonsourceibias.t58 gnd.t345 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 gnd.t344 commonsourceibias.t66 CSoutput.t189 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 CSoutput.t92 a_n7636_8799.t35 vdd.t260 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X19 vdd.t259 a_n7636_8799.t36 CSoutput.t91 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X20 gnd.t188 gnd.t186 gnd.t187 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X21 a_n2318_13878.t45 minus.t5 a_n3827_n3924.t39 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X22 gnd.t185 gnd.t182 gnd.t184 gnd.t183 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X23 a_n7636_8799.t1 plus.t6 a_n3827_n3924.t28 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X24 a_n7636_8799.t9 a_n2318_13878.t50 a_n2318_8322.t22 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X25 a_n2318_13878.t2 minus.t6 a_n3827_n3924.t4 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X26 vdd.t258 a_n7636_8799.t37 CSoutput.t90 vdd.t231 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X27 CSoutput.t89 a_n7636_8799.t38 vdd.t257 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X28 vdd.t256 a_n7636_8799.t39 CSoutput.t88 vdd.t228 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X29 commonsourceibias.t57 commonsourceibias.t56 gnd.t343 gnd.t273 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X30 a_n7636_8799.t10 a_n2318_13878.t51 a_n2318_8322.t21 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X31 gnd.t342 commonsourceibias.t67 CSoutput.t188 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 CSoutput.t187 commonsourceibias.t68 gnd.t341 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X33 vdd.t121 vdd.t119 vdd.t120 vdd.t50 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X34 gnd.t340 commonsourceibias.t54 commonsourceibias.t55 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 CSoutput.t192 a_n2318_8322.t27 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X36 CSoutput.t186 commonsourceibias.t69 gnd.t339 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 CSoutput.t87 a_n7636_8799.t40 vdd.t255 vdd.t218 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X38 a_n3827_n3924.t27 plus.t7 a_n7636_8799.t12 gnd.t39 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X39 a_n3827_n3924.t5 diffpairibias.t21 gnd.t18 gnd.t17 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X40 CSoutput.t86 a_n7636_8799.t41 vdd.t254 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X41 commonsourceibias.t53 commonsourceibias.t52 gnd.t338 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X42 a_n3827_n3924.t13 minus.t7 a_n2318_13878.t38 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X43 CSoutput.t185 commonsourceibias.t70 gnd.t337 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X44 CSoutput.t85 a_n7636_8799.t42 vdd.t253 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X45 gnd.t336 commonsourceibias.t50 commonsourceibias.t51 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X46 CSoutput.t184 commonsourceibias.t71 gnd.t335 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X47 a_n2140_13878.t14 a_n2318_13878.t29 a_n2318_13878.t30 vdd.t34 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X48 vdd.t118 vdd.t116 vdd.t117 vdd.t83 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X49 a_n2318_13878.t34 a_n2318_13878.t33 a_n2140_13878.t13 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X50 output.t3 outputibias.t8 gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X51 CSoutput.t193 a_n2318_8322.t25 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X52 gnd.t181 gnd.t179 plus.t4 gnd.t180 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X53 CSoutput.t84 a_n7636_8799.t43 vdd.t252 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X54 vdd.t115 vdd.t113 vdd.t114 vdd.t96 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X55 a_n3827_n3924.t26 plus.t8 a_n7636_8799.t4 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X56 vdd.t251 a_n7636_8799.t44 CSoutput.t83 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X57 vdd.t2 CSoutput.t194 output.t19 gnd.t2 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X58 diffpairibias.t19 diffpairibias.t18 gnd.t70 gnd.t69 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X59 CSoutput.t183 commonsourceibias.t72 gnd.t334 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X60 CSoutput.t182 commonsourceibias.t73 gnd.t333 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X61 CSoutput.t181 commonsourceibias.t74 gnd.t332 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X62 a_n7636_8799.t6 a_n2318_13878.t52 a_n2318_8322.t20 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X63 CSoutput.t82 a_n7636_8799.t45 vdd.t250 vdd.t215 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X64 commonsourceibias.t49 commonsourceibias.t48 gnd.t331 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X65 gnd.t178 gnd.t176 gnd.t177 gnd.t77 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X66 vdd.t249 a_n7636_8799.t46 CSoutput.t81 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X67 vdd.t244 a_n7636_8799.t47 CSoutput.t80 vdd.t228 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X68 diffpairibias.t17 diffpairibias.t16 gnd.t68 gnd.t67 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X69 CSoutput.t79 a_n7636_8799.t48 vdd.t248 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X70 gnd.t175 gnd.t173 gnd.t174 gnd.t77 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X71 vdd.t247 a_n7636_8799.t49 CSoutput.t78 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 CSoutput.t180 commonsourceibias.t75 gnd.t330 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X73 CSoutput.t77 a_n7636_8799.t50 vdd.t245 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 CSoutput.t76 a_n7636_8799.t51 vdd.t246 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X75 CSoutput.t75 a_n7636_8799.t52 vdd.t243 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X76 CSoutput.t74 a_n7636_8799.t53 vdd.t242 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X77 a_n3827_n3924.t40 minus.t8 a_n2318_13878.t46 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X78 a_n3827_n3924.t25 plus.t9 a_n7636_8799.t11 gnd.t14 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X79 gnd.t329 commonsourceibias.t76 CSoutput.t179 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 gnd.t172 gnd.t169 gnd.t171 gnd.t170 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X81 CSoutput.t178 commonsourceibias.t77 gnd.t299 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 gnd.t328 commonsourceibias.t78 CSoutput.t177 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X83 gnd.t168 gnd.t166 gnd.t167 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X84 a_n3827_n3924.t30 diffpairibias.t22 gnd.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X85 vdd.t241 a_n7636_8799.t54 CSoutput.t73 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 CSoutput.t176 commonsourceibias.t79 gnd.t327 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 a_n2318_13878.t4 a_n2318_13878.t3 a_n2140_13878.t12 vdd.t5 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X88 vdd.t240 a_n7636_8799.t55 CSoutput.t72 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X89 a_n3827_n3924.t24 plus.t10 a_n7636_8799.t25 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X90 a_n7636_8799.t7 a_n2318_13878.t53 a_n2318_8322.t19 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X91 vdd.t239 a_n7636_8799.t56 CSoutput.t71 vdd.t231 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X92 a_n2318_13878.t12 a_n2318_13878.t11 a_n2140_13878.t11 vdd.t8 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X93 outputibias.t7 outputibias.t6 gnd.t26 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X94 commonsourceibias.t33 commonsourceibias.t32 gnd.t326 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X95 gnd.t325 commonsourceibias.t80 CSoutput.t175 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X96 gnd.t165 gnd.t163 gnd.t164 gnd.t81 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X97 CSoutput.t174 commonsourceibias.t81 gnd.t324 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X98 gnd.t323 commonsourceibias.t30 commonsourceibias.t31 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X99 vdd.t238 a_n7636_8799.t57 CSoutput.t70 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X100 CSoutput.t173 commonsourceibias.t82 gnd.t322 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X101 CSoutput.t69 a_n7636_8799.t58 vdd.t237 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 diffpairibias.t15 diffpairibias.t14 gnd.t353 gnd.t352 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X103 vdd.t112 vdd.t110 vdd.t111 vdd.t100 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X104 vdd.t109 vdd.t107 vdd.t108 vdd.t62 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X105 CSoutput.t68 a_n7636_8799.t59 vdd.t236 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X106 vdd.t106 vdd.t103 vdd.t105 vdd.t104 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X107 gnd.t306 commonsourceibias.t83 CSoutput.t172 gnd.t225 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X108 vdd.t18 a_n2318_13878.t54 a_n2318_8322.t7 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X109 gnd.t321 commonsourceibias.t28 commonsourceibias.t29 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X110 a_n2318_13878.t32 a_n2318_13878.t31 a_n2140_13878.t10 vdd.t125 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X111 CSoutput.t171 commonsourceibias.t84 gnd.t320 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X112 gnd.t162 gnd.t160 minus.t3 gnd.t161 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X113 output.t18 CSoutput.t195 vdd.t3 gnd.t3 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X114 CSoutput.t170 commonsourceibias.t85 gnd.t319 gnd.t273 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X115 a_n2318_8322.t6 a_n2318_13878.t55 vdd.t20 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X116 a_n3827_n3924.t6 diffpairibias.t23 gnd.t20 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X117 CSoutput.t67 a_n7636_8799.t60 vdd.t235 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X118 CSoutput.t66 a_n7636_8799.t61 vdd.t233 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X119 gnd.t318 commonsourceibias.t86 CSoutput.t169 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 gnd.t159 gnd.t157 gnd.t158 gnd.t102 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X121 commonsourceibias.t27 commonsourceibias.t26 gnd.t317 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X122 vdd.t10 a_n2318_13878.t56 a_n2140_13878.t22 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X123 gnd.t308 commonsourceibias.t87 CSoutput.t168 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X124 vdd.t102 vdd.t99 vdd.t101 vdd.t100 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X125 gnd.t316 commonsourceibias.t24 commonsourceibias.t25 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X126 output.t17 CSoutput.t196 vdd.t4 gnd.t4 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X127 CSoutput.t167 commonsourceibias.t88 gnd.t315 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X128 gnd.t314 commonsourceibias.t89 CSoutput.t166 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X129 vdd.t232 a_n7636_8799.t62 CSoutput.t65 vdd.t231 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X130 CSoutput.t165 commonsourceibias.t90 gnd.t309 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X131 a_n7636_8799.t23 plus.t11 a_n3827_n3924.t23 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X132 commonsourceibias.t21 commonsourceibias.t20 gnd.t313 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 vdd.t98 vdd.t95 vdd.t97 vdd.t96 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X134 a_n2318_8322.t5 a_n2318_13878.t57 vdd.t12 vdd.t11 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X135 gnd.t312 commonsourceibias.t91 CSoutput.t164 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X136 a_n7636_8799.t18 a_n2318_13878.t58 a_n2318_8322.t18 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X137 a_n7636_8799.t3 plus.t12 a_n3827_n3924.t22 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X138 gnd.t156 gnd.t154 gnd.t155 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X139 CSoutput.t64 a_n7636_8799.t63 vdd.t230 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X140 diffpairibias.t13 diffpairibias.t12 gnd.t367 gnd.t366 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X141 vdd.t229 a_n7636_8799.t64 CSoutput.t63 vdd.t228 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X142 a_n2318_13878.t6 a_n2318_13878.t5 a_n2140_13878.t9 vdd.t131 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X143 vdd.t227 a_n7636_8799.t65 CSoutput.t62 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X144 a_n7636_8799.t19 a_n2318_13878.t59 a_n2318_8322.t17 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X145 CSoutput.t61 a_n7636_8799.t66 vdd.t226 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X146 gnd.t311 commonsourceibias.t18 commonsourceibias.t19 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X147 a_n2140_13878.t8 a_n2318_13878.t21 a_n2318_13878.t22 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X148 gnd.t153 gnd.t151 gnd.t152 gnd.t73 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X149 vdd.t94 vdd.t92 vdd.t93 vdd.t62 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X150 gnd.t310 commonsourceibias.t92 CSoutput.t163 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X151 output.t16 CSoutput.t197 vdd.t26 gnd.t31 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X152 gnd.t307 commonsourceibias.t93 CSoutput.t162 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X153 CSoutput.t60 a_n7636_8799.t67 vdd.t225 vdd.t215 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X154 vdd.t46 a_n2318_13878.t60 a_n2318_8322.t4 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X155 a_n2140_13878.t7 a_n2318_13878.t23 a_n2318_13878.t24 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X156 gnd.t150 gnd.t148 gnd.t149 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X157 vdd.t224 a_n7636_8799.t68 CSoutput.t59 vdd.t213 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X158 output.t2 outputibias.t9 gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X159 a_n2318_13878.t37 minus.t9 a_n3827_n3924.t9 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X160 a_n3827_n3924.t21 plus.t13 a_n7636_8799.t13 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X161 a_n2318_13878.t20 a_n2318_13878.t19 a_n2140_13878.t6 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X162 gnd.t147 gnd.t144 gnd.t146 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X163 gnd.t143 gnd.t141 gnd.t142 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X164 outputibias.t5 outputibias.t4 gnd.t55 gnd.t54 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X165 vdd.t27 CSoutput.t198 output.t15 gnd.t32 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X166 CSoutput.t161 commonsourceibias.t94 gnd.t305 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X167 plus.t3 gnd.t138 gnd.t140 gnd.t139 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X168 gnd.t304 commonsourceibias.t95 CSoutput.t160 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 gnd.t303 commonsourceibias.t96 CSoutput.t159 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X170 vdd.t223 a_n7636_8799.t69 CSoutput.t58 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X171 a_n3827_n3924.t1 diffpairibias.t24 gnd.t12 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X172 gnd.t137 gnd.t135 minus.t2 gnd.t136 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X173 a_n3827_n3924.t37 diffpairibias.t25 gnd.t355 gnd.t354 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X174 outputibias.t3 outputibias.t2 gnd.t359 gnd.t358 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X175 a_n7636_8799.t29 plus.t14 a_n3827_n3924.t20 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X176 vdd.t222 a_n7636_8799.t70 CSoutput.t57 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X177 vdd.t220 a_n7636_8799.t71 CSoutput.t56 vdd.t177 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X178 gnd.t134 gnd.t132 gnd.t133 gnd.t81 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X179 a_n7636_8799.t2 plus.t15 a_n3827_n3924.t19 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X180 gnd.t131 gnd.t129 gnd.t130 gnd.t81 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X181 CSoutput.t55 a_n7636_8799.t72 vdd.t221 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X182 CSoutput.t54 a_n7636_8799.t73 vdd.t219 vdd.t218 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X183 vdd.t28 CSoutput.t199 output.t14 gnd.t33 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X184 CSoutput.t53 a_n7636_8799.t74 vdd.t217 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X185 CSoutput.t158 commonsourceibias.t97 gnd.t302 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X186 output.t13 CSoutput.t200 vdd.t6 gnd.t9 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X187 gnd.t128 gnd.t126 gnd.t127 gnd.t77 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X188 gnd.t301 commonsourceibias.t98 CSoutput.t157 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 diffpairibias.t11 diffpairibias.t10 gnd.t28 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X190 a_n2140_13878.t21 a_n2318_13878.t61 vdd.t48 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X191 a_n2318_13878.t47 minus.t10 a_n3827_n3924.t41 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X192 vdd.t39 a_n2318_13878.t62 a_n2140_13878.t20 vdd.t38 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X193 vdd.t91 vdd.t89 vdd.t90 vdd.t79 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X194 CSoutput.t52 a_n7636_8799.t75 vdd.t216 vdd.t215 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X195 gnd.t300 commonsourceibias.t99 CSoutput.t156 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 CSoutput.t155 commonsourceibias.t100 gnd.t298 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X197 a_n3827_n3924.t18 plus.t16 a_n7636_8799.t20 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X198 vdd.t214 a_n7636_8799.t76 CSoutput.t51 vdd.t213 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X199 output.t12 CSoutput.t201 vdd.t7 gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X200 vdd.t88 vdd.t86 vdd.t87 vdd.t79 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X201 a_n2140_13878.t5 a_n2318_13878.t15 a_n2318_13878.t16 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X202 diffpairibias.t9 diffpairibias.t8 gnd.t361 gnd.t360 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X203 gnd.t297 commonsourceibias.t101 CSoutput.t154 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X204 vdd.t212 a_n7636_8799.t77 CSoutput.t50 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X205 commonsourceibias.t41 commonsourceibias.t40 gnd.t296 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X206 a_n3827_n3924.t35 minus.t11 a_n2318_13878.t43 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X207 a_n2318_8322.t16 a_n2318_13878.t63 a_n7636_8799.t16 vdd.t40 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X208 CSoutput.t49 a_n7636_8799.t78 vdd.t211 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X209 outputibias.t1 outputibias.t0 gnd.t41 gnd.t40 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X210 diffpairibias.t7 diffpairibias.t6 gnd.t48 gnd.t47 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X211 vdd.t205 a_n7636_8799.t79 CSoutput.t48 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X212 vdd.t133 a_n2318_13878.t64 a_n2318_8322.t3 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X213 vdd.t210 a_n7636_8799.t80 CSoutput.t47 vdd.t177 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X214 vdd.t207 a_n7636_8799.t81 CSoutput.t46 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X215 output.t1 outputibias.t10 gnd.t357 gnd.t356 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X216 CSoutput.t153 commonsourceibias.t102 gnd.t295 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X217 plus.t2 gnd.t123 gnd.t125 gnd.t124 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X218 CSoutput.t202 a_n2318_8322.t27 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X219 gnd.t122 gnd.t120 minus.t1 gnd.t121 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X220 commonsourceibias.t39 commonsourceibias.t38 gnd.t294 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X221 gnd.t119 gnd.t116 gnd.t118 gnd.t117 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X222 a_n2140_13878.t19 a_n2318_13878.t65 vdd.t135 vdd.t134 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X223 vdd.t0 CSoutput.t203 output.t11 gnd.t0 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X224 CSoutput.t152 commonsourceibias.t103 gnd.t293 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X225 vdd.t209 a_n7636_8799.t82 CSoutput.t45 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X226 gnd.t292 commonsourceibias.t104 CSoutput.t151 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X227 CSoutput.t204 a_n2318_8322.t26 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X228 CSoutput.t44 a_n7636_8799.t83 vdd.t208 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 CSoutput.t43 a_n7636_8799.t84 vdd.t203 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X230 gnd.t291 commonsourceibias.t36 commonsourceibias.t37 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X231 gnd.t290 commonsourceibias.t105 CSoutput.t150 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X232 CSoutput.t149 commonsourceibias.t106 gnd.t289 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X233 gnd.t115 gnd.t112 gnd.t114 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X234 CSoutput.t148 commonsourceibias.t107 gnd.t288 gnd.t273 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 vdd.t85 vdd.t82 vdd.t84 vdd.t83 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X236 gnd.t287 commonsourceibias.t108 CSoutput.t147 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X237 CSoutput.t146 commonsourceibias.t109 gnd.t286 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X238 a_n3827_n3924.t11 diffpairibias.t26 gnd.t53 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X239 gnd.t284 commonsourceibias.t110 CSoutput.t145 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 commonsourceibias.t35 commonsourceibias.t34 gnd.t283 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X241 vdd.t81 vdd.t78 vdd.t80 vdd.t79 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X242 vdd.t130 a_n2318_13878.t66 a_n2318_8322.t2 vdd.t129 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X243 a_n2318_8322.t15 a_n2318_13878.t67 a_n7636_8799.t27 vdd.t131 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X244 CSoutput.t42 a_n7636_8799.t85 vdd.t200 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X245 a_n7636_8799.t15 plus.t17 a_n3827_n3924.t17 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X246 vdd.t202 a_n7636_8799.t86 CSoutput.t41 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X247 a_n2318_13878.t42 minus.t12 a_n3827_n3924.t34 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X248 CSoutput.t144 commonsourceibias.t111 gnd.t282 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X249 CSoutput.t40 a_n7636_8799.t87 vdd.t201 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X250 gnd.t281 commonsourceibias.t112 CSoutput.t143 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X251 a_n3827_n3924.t3 minus.t13 a_n2318_13878.t1 gnd.t14 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X252 vdd.t198 a_n7636_8799.t88 CSoutput.t39 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X253 vdd.t197 a_n7636_8799.t89 CSoutput.t38 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X254 CSoutput.t142 commonsourceibias.t113 gnd.t280 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X255 gnd.t254 commonsourceibias.t114 CSoutput.t141 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X256 vdd.t77 vdd.t75 vdd.t76 vdd.t58 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X257 gnd.t278 commonsourceibias.t115 CSoutput.t140 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X258 CSoutput.t139 commonsourceibias.t116 gnd.t279 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X259 commonsourceibias.t17 commonsourceibias.t16 gnd.t277 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 vdd.t74 vdd.t71 vdd.t73 vdd.t72 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X261 a_n3827_n3924.t2 minus.t14 a_n2318_13878.t0 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X262 vdd.t196 a_n7636_8799.t90 CSoutput.t37 vdd.t142 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X263 CSoutput.t36 a_n7636_8799.t91 vdd.t195 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X264 a_n3827_n3924.t8 minus.t15 a_n2318_13878.t36 gnd.t39 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X265 a_n2140_13878.t4 a_n2318_13878.t27 a_n2318_13878.t28 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X266 CSoutput.t35 a_n7636_8799.t92 vdd.t193 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X267 CSoutput.t138 commonsourceibias.t117 gnd.t275 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X268 gnd.t111 gnd.t108 gnd.t110 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X269 a_n2318_8322.t14 a_n2318_13878.t68 a_n7636_8799.t26 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X270 diffpairibias.t5 diffpairibias.t4 gnd.t60 gnd.t59 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X271 gnd.t272 commonsourceibias.t118 CSoutput.t137 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X272 CSoutput.t136 commonsourceibias.t119 gnd.t274 gnd.t273 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X273 gnd.t270 commonsourceibias.t14 commonsourceibias.t15 gnd.t225 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X274 gnd.t107 gnd.t105 gnd.t106 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X275 output.t10 CSoutput.t205 vdd.t1 gnd.t1 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X276 commonsourceibias.t13 commonsourceibias.t12 gnd.t269 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X277 CSoutput.t34 a_n7636_8799.t93 vdd.t192 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X278 gnd.t259 commonsourceibias.t120 CSoutput.t135 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X279 CSoutput.t33 a_n7636_8799.t94 vdd.t190 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X280 a_n3827_n3924.t10 diffpairibias.t27 gnd.t50 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X281 vdd.t189 a_n7636_8799.t95 CSoutput.t32 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X282 gnd.t258 commonsourceibias.t121 CSoutput.t134 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X283 vdd.t188 a_n7636_8799.t96 CSoutput.t31 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X284 a_n2318_8322.t1 a_n2318_13878.t69 vdd.t128 vdd.t127 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X285 gnd.t268 commonsourceibias.t122 CSoutput.t133 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 CSoutput.t132 commonsourceibias.t123 gnd.t266 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 CSoutput.t30 a_n7636_8799.t97 vdd.t186 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 output.t9 CSoutput.t206 vdd.t29 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X289 gnd.t267 commonsourceibias.t10 commonsourceibias.t11 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X290 a_n3827_n3924.t33 minus.t16 a_n2318_13878.t41 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X291 vdd.t70 vdd.t68 vdd.t69 vdd.t54 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X292 commonsourceibias.t9 commonsourceibias.t8 gnd.t265 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X293 vdd.t265 a_n2318_13878.t70 a_n2140_13878.t18 vdd.t264 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X294 CSoutput.t29 a_n7636_8799.t98 vdd.t184 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X295 gnd.t263 commonsourceibias.t124 CSoutput.t131 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X296 CSoutput.t130 commonsourceibias.t125 gnd.t264 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X297 CSoutput.t28 a_n7636_8799.t99 vdd.t182 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X298 CSoutput.t129 commonsourceibias.t126 gnd.t262 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X299 gnd.t260 commonsourceibias.t127 CSoutput.t128 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X300 commonsourceibias.t63 commonsourceibias.t62 gnd.t256 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 gnd.t252 commonsourceibias.t128 CSoutput.t127 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X302 vdd.t181 a_n7636_8799.t100 CSoutput.t27 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X303 vdd.t179 a_n7636_8799.t101 CSoutput.t26 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X304 gnd.t104 gnd.t101 gnd.t103 gnd.t102 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X305 gnd.t251 commonsourceibias.t60 commonsourceibias.t61 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X306 gnd.t100 gnd.t98 plus.t1 gnd.t99 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X307 gnd.t97 gnd.t94 gnd.t96 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X308 vdd.t67 vdd.t65 vdd.t66 vdd.t58 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X309 a_n2318_8322.t13 a_n2318_13878.t71 a_n7636_8799.t28 vdd.t36 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X310 CSoutput.t25 a_n7636_8799.t102 vdd.t173 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X311 a_n7636_8799.t31 a_n2318_13878.t72 a_n2318_8322.t12 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X312 gnd.t250 commonsourceibias.t129 CSoutput.t126 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X313 vdd.t178 a_n7636_8799.t103 CSoutput.t24 vdd.t177 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X314 a_n2140_13878.t17 a_n2318_13878.t73 vdd.t267 vdd.t266 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X315 CSoutput.t125 commonsourceibias.t130 gnd.t248 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X316 vdd.t176 a_n7636_8799.t104 CSoutput.t23 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X317 gnd.t247 commonsourceibias.t131 CSoutput.t124 gnd.t225 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X318 CSoutput.t22 a_n7636_8799.t105 vdd.t175 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 vdd.t30 CSoutput.t207 output.t8 gnd.t35 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X320 vdd.t31 CSoutput.t208 output.t7 gnd.t36 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X321 gnd.t246 commonsourceibias.t46 commonsourceibias.t47 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X322 CSoutput.t123 commonsourceibias.t132 gnd.t245 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X323 CSoutput.t122 commonsourceibias.t133 gnd.t244 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X324 a_n3827_n3924.t16 plus.t18 a_n7636_8799.t0 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X325 a_n2318_13878.t39 minus.t17 a_n3827_n3924.t31 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X326 CSoutput.t121 commonsourceibias.t134 gnd.t243 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X327 gnd.t242 commonsourceibias.t135 CSoutput.t120 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X328 CSoutput.t119 commonsourceibias.t136 gnd.t241 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X329 a_n2318_8322.t11 a_n2318_13878.t74 a_n7636_8799.t21 vdd.t125 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X330 CSoutput.t209 a_n2318_8322.t25 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X331 vdd.t171 a_n7636_8799.t106 CSoutput.t21 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X332 CSoutput.t20 a_n7636_8799.t107 vdd.t169 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X333 CSoutput.t19 a_n7636_8799.t108 vdd.t162 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X334 CSoutput.t118 commonsourceibias.t137 gnd.t239 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X335 CSoutput.t117 commonsourceibias.t138 gnd.t237 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 gnd.t236 commonsourceibias.t139 CSoutput.t116 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X337 CSoutput.t18 a_n7636_8799.t109 vdd.t164 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X338 a_n2140_13878.t3 a_n2318_13878.t9 a_n2318_13878.t10 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X339 vdd.t167 a_n7636_8799.t110 CSoutput.t17 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 vdd.t64 vdd.t61 vdd.t63 vdd.t62 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X341 gnd.t235 commonsourceibias.t44 commonsourceibias.t45 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X342 vdd.t60 vdd.t57 vdd.t59 vdd.t58 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X343 gnd.t233 commonsourceibias.t42 commonsourceibias.t43 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X344 a_n3827_n3924.t32 minus.t18 a_n2318_13878.t40 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X345 a_n3827_n3924.t12 diffpairibias.t28 gnd.t57 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X346 vdd.t166 a_n7636_8799.t111 CSoutput.t16 vdd.t142 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X347 vdd.t165 a_n7636_8799.t112 CSoutput.t15 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X348 CSoutput.t115 commonsourceibias.t140 gnd.t231 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 gnd.t224 commonsourceibias.t141 CSoutput.t114 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X350 CSoutput.t14 a_n7636_8799.t113 vdd.t163 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X351 a_n2318_13878.t18 a_n2318_13878.t17 a_n2140_13878.t2 vdd.t36 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X352 a_n7636_8799.t22 a_n2318_13878.t75 a_n2318_8322.t10 vdd.t34 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X353 vdd.t161 a_n7636_8799.t114 CSoutput.t13 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X354 CSoutput.t12 a_n7636_8799.t115 vdd.t160 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X355 CSoutput.t113 commonsourceibias.t142 gnd.t229 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X356 vdd.t158 a_n7636_8799.t116 CSoutput.t11 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X357 gnd.t93 gnd.t90 gnd.t92 gnd.t91 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X358 gnd.t227 commonsourceibias.t143 CSoutput.t112 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X359 gnd.t226 commonsourceibias.t144 CSoutput.t111 gnd.t225 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X360 gnd.t222 commonsourceibias.t145 CSoutput.t110 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X361 diffpairibias.t3 diffpairibias.t2 gnd.t365 gnd.t364 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X362 vdd.t157 a_n7636_8799.t117 CSoutput.t10 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X363 gnd.t89 gnd.t87 plus.t0 gnd.t88 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X364 CSoutput.t109 commonsourceibias.t146 gnd.t220 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X365 minus.t0 gnd.t84 gnd.t86 gnd.t85 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X366 CSoutput.t9 a_n7636_8799.t118 vdd.t155 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X367 output.t6 CSoutput.t210 vdd.t24 gnd.t29 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X368 a_n2318_8322.t9 a_n2318_13878.t76 a_n7636_8799.t17 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X369 gnd.t83 gnd.t80 gnd.t82 gnd.t81 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X370 vdd.t25 CSoutput.t211 output.t5 gnd.t30 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X371 a_n2318_13878.t35 minus.t19 a_n3827_n3924.t7 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X372 gnd.t213 commonsourceibias.t147 CSoutput.t108 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X373 gnd.t218 commonsourceibias.t148 CSoutput.t107 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X374 vdd.t153 a_n7636_8799.t119 CSoutput.t8 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X375 gnd.t79 gnd.t76 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X376 diffpairibias.t1 diffpairibias.t0 gnd.t44 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X377 CSoutput.t106 commonsourceibias.t149 gnd.t216 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X378 CSoutput.t212 a_n2318_8322.t24 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X379 gnd.t214 commonsourceibias.t150 CSoutput.t105 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X380 vdd.t56 vdd.t53 vdd.t55 vdd.t54 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X381 vdd.t43 a_n2318_13878.t77 a_n2140_13878.t16 vdd.t42 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X382 CSoutput.t7 a_n7636_8799.t120 vdd.t151 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X383 vdd.t52 vdd.t49 vdd.t51 vdd.t50 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X384 vdd.t149 a_n7636_8799.t121 CSoutput.t6 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X385 gnd.t211 commonsourceibias.t151 CSoutput.t104 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X386 vdd.t147 a_n7636_8799.t122 CSoutput.t5 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X387 CSoutput.t4 a_n7636_8799.t123 vdd.t145 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X388 a_n7636_8799.t24 plus.t19 a_n3827_n3924.t15 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X389 gnd.t209 commonsourceibias.t152 CSoutput.t103 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X390 a_n2318_13878.t44 minus.t20 a_n3827_n3924.t36 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X391 a_n2318_8322.t8 a_n2318_13878.t78 a_n7636_8799.t14 vdd.t8 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X392 CSoutput.t102 commonsourceibias.t153 gnd.t207 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X393 vdd.t143 a_n7636_8799.t124 CSoutput.t3 vdd.t142 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X394 vdd.t141 a_n7636_8799.t125 CSoutput.t2 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X395 output.t0 outputibias.t11 gnd.t46 gnd.t45 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X396 CSoutput.t1 a_n7636_8799.t126 vdd.t139 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X397 gnd.t205 commonsourceibias.t154 CSoutput.t101 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X398 commonsourceibias.t23 commonsourceibias.t22 gnd.t203 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X399 gnd.t201 commonsourceibias.t155 CSoutput.t100 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X400 CSoutput.t99 commonsourceibias.t156 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X401 a_n2318_8322.t0 a_n2318_13878.t79 vdd.t33 vdd.t32 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X402 gnd.t75 gnd.t72 gnd.t74 gnd.t73 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X403 a_n2140_13878.t1 a_n2318_13878.t25 a_n2318_13878.t26 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X404 vdd.t23 CSoutput.t213 output.t4 gnd.t24 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X405 vdd.t137 a_n7636_8799.t127 CSoutput.t0 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X406 a_n3827_n3924.t14 plus.t20 a_n7636_8799.t30 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X407 a_n3827_n3924.t38 diffpairibias.t29 gnd.t363 gnd.t362 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X408 CSoutput.t98 commonsourceibias.t157 gnd.t197 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X409 CSoutput.t97 commonsourceibias.t158 gnd.t195 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X410 a_n2318_13878.t14 a_n2318_13878.t13 a_n2140_13878.t0 vdd.t40 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X411 gnd.t193 commonsourceibias.t159 CSoutput.t96 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
R0 commonsourceibias.n35 commonsourceibias.t48 223.028
R1 commonsourceibias.n128 commonsourceibias.t132 223.028
R2 commonsourceibias.n307 commonsourceibias.t136 223.028
R3 commonsourceibias.n217 commonsourceibias.t64 223.028
R4 commonsourceibias.n454 commonsourceibias.t14 223.028
R5 commonsourceibias.n395 commonsourceibias.t83 223.028
R6 commonsourceibias.n679 commonsourceibias.t144 223.028
R7 commonsourceibias.n589 commonsourceibias.t131 223.028
R8 commonsourceibias.n99 commonsourceibias.t36 207.983
R9 commonsourceibias.n192 commonsourceibias.t78 207.983
R10 commonsourceibias.n371 commonsourceibias.t148 207.983
R11 commonsourceibias.n281 commonsourceibias.t115 207.983
R12 commonsourceibias.n520 commonsourceibias.t26 207.983
R13 commonsourceibias.n566 commonsourceibias.t153 207.983
R14 commonsourceibias.n745 commonsourceibias.t71 207.983
R15 commonsourceibias.n655 commonsourceibias.t100 207.983
R16 commonsourceibias.n97 commonsourceibias.t32 168.701
R17 commonsourceibias.n91 commonsourceibias.t42 168.701
R18 commonsourceibias.n17 commonsourceibias.t20 168.701
R19 commonsourceibias.n83 commonsourceibias.t0 168.701
R20 commonsourceibias.n77 commonsourceibias.t38 168.701
R21 commonsourceibias.n22 commonsourceibias.t50 168.701
R22 commonsourceibias.n69 commonsourceibias.t58 168.701
R23 commonsourceibias.n63 commonsourceibias.t24 168.701
R24 commonsourceibias.n25 commonsourceibias.t4 168.701
R25 commonsourceibias.n27 commonsourceibias.t46 168.701
R26 commonsourceibias.n29 commonsourceibias.t52 168.701
R27 commonsourceibias.n46 commonsourceibias.t2 168.701
R28 commonsourceibias.n40 commonsourceibias.t16 168.701
R29 commonsourceibias.n34 commonsourceibias.t30 168.701
R30 commonsourceibias.n190 commonsourceibias.t146 168.701
R31 commonsourceibias.n184 commonsourceibias.t96 168.701
R32 commonsourceibias.n5 commonsourceibias.t157 168.701
R33 commonsourceibias.n176 commonsourceibias.t112 168.701
R34 commonsourceibias.n170 commonsourceibias.t75 168.701
R35 commonsourceibias.n10 commonsourceibias.t124 168.701
R36 commonsourceibias.n162 commonsourceibias.t113 168.701
R37 commonsourceibias.n156 commonsourceibias.t154 168.701
R38 commonsourceibias.n118 commonsourceibias.t106 168.701
R39 commonsourceibias.n120 commonsourceibias.t92 168.701
R40 commonsourceibias.n122 commonsourceibias.t123 168.701
R41 commonsourceibias.n139 commonsourceibias.t110 168.701
R42 commonsourceibias.n133 commonsourceibias.t82 168.701
R43 commonsourceibias.n127 commonsourceibias.t147 168.701
R44 commonsourceibias.n306 commonsourceibias.t143 168.701
R45 commonsourceibias.n312 commonsourceibias.t70 168.701
R46 commonsourceibias.n318 commonsourceibias.t150 168.701
R47 commonsourceibias.n301 commonsourceibias.t158 168.701
R48 commonsourceibias.n299 commonsourceibias.t101 168.701
R49 commonsourceibias.n297 commonsourceibias.t81 168.701
R50 commonsourceibias.n335 commonsourceibias.t67 168.701
R51 commonsourceibias.n341 commonsourceibias.t111 168.701
R52 commonsourceibias.n294 commonsourceibias.t120 168.701
R53 commonsourceibias.n349 commonsourceibias.t74 168.701
R54 commonsourceibias.n355 commonsourceibias.t159 168.701
R55 commonsourceibias.n289 commonsourceibias.t134 168.701
R56 commonsourceibias.n363 commonsourceibias.t80 168.701
R57 commonsourceibias.n369 commonsourceibias.t68 168.701
R58 commonsourceibias.n279 commonsourceibias.t138 168.701
R59 commonsourceibias.n273 commonsourceibias.t128 168.701
R60 commonsourceibias.n199 commonsourceibias.t116 168.701
R61 commonsourceibias.n265 commonsourceibias.t139 168.701
R62 commonsourceibias.n259 commonsourceibias.t126 168.701
R63 commonsourceibias.n204 commonsourceibias.t114 168.701
R64 commonsourceibias.n251 commonsourceibias.t140 168.701
R65 commonsourceibias.n245 commonsourceibias.t127 168.701
R66 commonsourceibias.n207 commonsourceibias.t149 168.701
R67 commonsourceibias.n209 commonsourceibias.t141 168.701
R68 commonsourceibias.n211 commonsourceibias.t125 168.701
R69 commonsourceibias.n228 commonsourceibias.t152 168.701
R70 commonsourceibias.n222 commonsourceibias.t69 168.701
R71 commonsourceibias.n216 commonsourceibias.t135 168.701
R72 commonsourceibias.n453 commonsourceibias.t12 168.701
R73 commonsourceibias.n459 commonsourceibias.t18 168.701
R74 commonsourceibias.n465 commonsourceibias.t8 168.701
R75 commonsourceibias.n448 commonsourceibias.t44 168.701
R76 commonsourceibias.n446 commonsourceibias.t34 168.701
R77 commonsourceibias.n444 commonsourceibias.t10 168.701
R78 commonsourceibias.n482 commonsourceibias.t56 168.701
R79 commonsourceibias.n488 commonsourceibias.t60 168.701
R80 commonsourceibias.n490 commonsourceibias.t22 168.701
R81 commonsourceibias.n497 commonsourceibias.t28 168.701
R82 commonsourceibias.n503 commonsourceibias.t62 168.701
R83 commonsourceibias.n505 commonsourceibias.t54 168.701
R84 commonsourceibias.n512 commonsourceibias.t40 168.701
R85 commonsourceibias.n518 commonsourceibias.t6 168.701
R86 commonsourceibias.n564 commonsourceibias.t104 168.701
R87 commonsourceibias.n558 commonsourceibias.t73 168.701
R88 commonsourceibias.n551 commonsourceibias.t121 168.701
R89 commonsourceibias.n549 commonsourceibias.t90 168.701
R90 commonsourceibias.n543 commonsourceibias.t151 168.701
R91 commonsourceibias.n536 commonsourceibias.t102 168.701
R92 commonsourceibias.n534 commonsourceibias.t91 168.701
R93 commonsourceibias.n394 commonsourceibias.t84 168.701
R94 commonsourceibias.n400 commonsourceibias.t65 168.701
R95 commonsourceibias.n406 commonsourceibias.t88 168.701
R96 commonsourceibias.n389 commonsourceibias.t95 168.701
R97 commonsourceibias.n387 commonsourceibias.t79 168.701
R98 commonsourceibias.n385 commonsourceibias.t87 168.701
R99 commonsourceibias.n423 commonsourceibias.t119 168.701
R100 commonsourceibias.n678 commonsourceibias.t133 168.701
R101 commonsourceibias.n684 commonsourceibias.t89 168.701
R102 commonsourceibias.n690 commonsourceibias.t72 168.701
R103 commonsourceibias.n673 commonsourceibias.t76 168.701
R104 commonsourceibias.n671 commonsourceibias.t94 168.701
R105 commonsourceibias.n669 commonsourceibias.t98 168.701
R106 commonsourceibias.n707 commonsourceibias.t85 168.701
R107 commonsourceibias.n713 commonsourceibias.t145 168.701
R108 commonsourceibias.n715 commonsourceibias.t103 168.701
R109 commonsourceibias.n722 commonsourceibias.t93 168.701
R110 commonsourceibias.n728 commonsourceibias.t77 168.701
R111 commonsourceibias.n730 commonsourceibias.t66 168.701
R112 commonsourceibias.n737 commonsourceibias.t97 168.701
R113 commonsourceibias.n743 commonsourceibias.t86 168.701
R114 commonsourceibias.n588 commonsourceibias.t142 168.701
R115 commonsourceibias.n594 commonsourceibias.t155 168.701
R116 commonsourceibias.n600 commonsourceibias.t137 168.701
R117 commonsourceibias.n583 commonsourceibias.t105 168.701
R118 commonsourceibias.n581 commonsourceibias.t156 168.701
R119 commonsourceibias.n579 commonsourceibias.t129 168.701
R120 commonsourceibias.n617 commonsourceibias.t107 168.701
R121 commonsourceibias.n623 commonsourceibias.t122 168.701
R122 commonsourceibias.n625 commonsourceibias.t130 168.701
R123 commonsourceibias.n632 commonsourceibias.t108 168.701
R124 commonsourceibias.n638 commonsourceibias.t117 168.701
R125 commonsourceibias.n640 commonsourceibias.t99 168.701
R126 commonsourceibias.n647 commonsourceibias.t109 168.701
R127 commonsourceibias.n653 commonsourceibias.t118 168.701
R128 commonsourceibias.n36 commonsourceibias.n33 161.3
R129 commonsourceibias.n38 commonsourceibias.n37 161.3
R130 commonsourceibias.n39 commonsourceibias.n32 161.3
R131 commonsourceibias.n42 commonsourceibias.n41 161.3
R132 commonsourceibias.n43 commonsourceibias.n31 161.3
R133 commonsourceibias.n45 commonsourceibias.n44 161.3
R134 commonsourceibias.n47 commonsourceibias.n30 161.3
R135 commonsourceibias.n49 commonsourceibias.n48 161.3
R136 commonsourceibias.n51 commonsourceibias.n50 161.3
R137 commonsourceibias.n52 commonsourceibias.n28 161.3
R138 commonsourceibias.n54 commonsourceibias.n53 161.3
R139 commonsourceibias.n56 commonsourceibias.n55 161.3
R140 commonsourceibias.n57 commonsourceibias.n26 161.3
R141 commonsourceibias.n59 commonsourceibias.n58 161.3
R142 commonsourceibias.n61 commonsourceibias.n60 161.3
R143 commonsourceibias.n62 commonsourceibias.n24 161.3
R144 commonsourceibias.n65 commonsourceibias.n64 161.3
R145 commonsourceibias.n66 commonsourceibias.n23 161.3
R146 commonsourceibias.n68 commonsourceibias.n67 161.3
R147 commonsourceibias.n70 commonsourceibias.n21 161.3
R148 commonsourceibias.n72 commonsourceibias.n71 161.3
R149 commonsourceibias.n73 commonsourceibias.n20 161.3
R150 commonsourceibias.n75 commonsourceibias.n74 161.3
R151 commonsourceibias.n76 commonsourceibias.n19 161.3
R152 commonsourceibias.n79 commonsourceibias.n78 161.3
R153 commonsourceibias.n80 commonsourceibias.n18 161.3
R154 commonsourceibias.n82 commonsourceibias.n81 161.3
R155 commonsourceibias.n84 commonsourceibias.n16 161.3
R156 commonsourceibias.n86 commonsourceibias.n85 161.3
R157 commonsourceibias.n87 commonsourceibias.n15 161.3
R158 commonsourceibias.n89 commonsourceibias.n88 161.3
R159 commonsourceibias.n90 commonsourceibias.n14 161.3
R160 commonsourceibias.n93 commonsourceibias.n92 161.3
R161 commonsourceibias.n94 commonsourceibias.n13 161.3
R162 commonsourceibias.n96 commonsourceibias.n95 161.3
R163 commonsourceibias.n98 commonsourceibias.n12 161.3
R164 commonsourceibias.n129 commonsourceibias.n126 161.3
R165 commonsourceibias.n131 commonsourceibias.n130 161.3
R166 commonsourceibias.n132 commonsourceibias.n125 161.3
R167 commonsourceibias.n135 commonsourceibias.n134 161.3
R168 commonsourceibias.n136 commonsourceibias.n124 161.3
R169 commonsourceibias.n138 commonsourceibias.n137 161.3
R170 commonsourceibias.n140 commonsourceibias.n123 161.3
R171 commonsourceibias.n142 commonsourceibias.n141 161.3
R172 commonsourceibias.n144 commonsourceibias.n143 161.3
R173 commonsourceibias.n145 commonsourceibias.n121 161.3
R174 commonsourceibias.n147 commonsourceibias.n146 161.3
R175 commonsourceibias.n149 commonsourceibias.n148 161.3
R176 commonsourceibias.n150 commonsourceibias.n119 161.3
R177 commonsourceibias.n152 commonsourceibias.n151 161.3
R178 commonsourceibias.n154 commonsourceibias.n153 161.3
R179 commonsourceibias.n155 commonsourceibias.n117 161.3
R180 commonsourceibias.n158 commonsourceibias.n157 161.3
R181 commonsourceibias.n159 commonsourceibias.n11 161.3
R182 commonsourceibias.n161 commonsourceibias.n160 161.3
R183 commonsourceibias.n163 commonsourceibias.n9 161.3
R184 commonsourceibias.n165 commonsourceibias.n164 161.3
R185 commonsourceibias.n166 commonsourceibias.n8 161.3
R186 commonsourceibias.n168 commonsourceibias.n167 161.3
R187 commonsourceibias.n169 commonsourceibias.n7 161.3
R188 commonsourceibias.n172 commonsourceibias.n171 161.3
R189 commonsourceibias.n173 commonsourceibias.n6 161.3
R190 commonsourceibias.n175 commonsourceibias.n174 161.3
R191 commonsourceibias.n177 commonsourceibias.n4 161.3
R192 commonsourceibias.n179 commonsourceibias.n178 161.3
R193 commonsourceibias.n180 commonsourceibias.n3 161.3
R194 commonsourceibias.n182 commonsourceibias.n181 161.3
R195 commonsourceibias.n183 commonsourceibias.n2 161.3
R196 commonsourceibias.n186 commonsourceibias.n185 161.3
R197 commonsourceibias.n187 commonsourceibias.n1 161.3
R198 commonsourceibias.n189 commonsourceibias.n188 161.3
R199 commonsourceibias.n191 commonsourceibias.n0 161.3
R200 commonsourceibias.n370 commonsourceibias.n284 161.3
R201 commonsourceibias.n368 commonsourceibias.n367 161.3
R202 commonsourceibias.n366 commonsourceibias.n285 161.3
R203 commonsourceibias.n365 commonsourceibias.n364 161.3
R204 commonsourceibias.n362 commonsourceibias.n286 161.3
R205 commonsourceibias.n361 commonsourceibias.n360 161.3
R206 commonsourceibias.n359 commonsourceibias.n287 161.3
R207 commonsourceibias.n358 commonsourceibias.n357 161.3
R208 commonsourceibias.n356 commonsourceibias.n288 161.3
R209 commonsourceibias.n354 commonsourceibias.n353 161.3
R210 commonsourceibias.n352 commonsourceibias.n290 161.3
R211 commonsourceibias.n351 commonsourceibias.n350 161.3
R212 commonsourceibias.n348 commonsourceibias.n291 161.3
R213 commonsourceibias.n347 commonsourceibias.n346 161.3
R214 commonsourceibias.n345 commonsourceibias.n292 161.3
R215 commonsourceibias.n344 commonsourceibias.n343 161.3
R216 commonsourceibias.n342 commonsourceibias.n293 161.3
R217 commonsourceibias.n340 commonsourceibias.n339 161.3
R218 commonsourceibias.n338 commonsourceibias.n295 161.3
R219 commonsourceibias.n337 commonsourceibias.n336 161.3
R220 commonsourceibias.n334 commonsourceibias.n296 161.3
R221 commonsourceibias.n333 commonsourceibias.n332 161.3
R222 commonsourceibias.n331 commonsourceibias.n330 161.3
R223 commonsourceibias.n329 commonsourceibias.n298 161.3
R224 commonsourceibias.n328 commonsourceibias.n327 161.3
R225 commonsourceibias.n326 commonsourceibias.n325 161.3
R226 commonsourceibias.n324 commonsourceibias.n300 161.3
R227 commonsourceibias.n323 commonsourceibias.n322 161.3
R228 commonsourceibias.n321 commonsourceibias.n320 161.3
R229 commonsourceibias.n319 commonsourceibias.n302 161.3
R230 commonsourceibias.n317 commonsourceibias.n316 161.3
R231 commonsourceibias.n315 commonsourceibias.n303 161.3
R232 commonsourceibias.n314 commonsourceibias.n313 161.3
R233 commonsourceibias.n311 commonsourceibias.n304 161.3
R234 commonsourceibias.n310 commonsourceibias.n309 161.3
R235 commonsourceibias.n308 commonsourceibias.n305 161.3
R236 commonsourceibias.n218 commonsourceibias.n215 161.3
R237 commonsourceibias.n220 commonsourceibias.n219 161.3
R238 commonsourceibias.n221 commonsourceibias.n214 161.3
R239 commonsourceibias.n224 commonsourceibias.n223 161.3
R240 commonsourceibias.n225 commonsourceibias.n213 161.3
R241 commonsourceibias.n227 commonsourceibias.n226 161.3
R242 commonsourceibias.n229 commonsourceibias.n212 161.3
R243 commonsourceibias.n231 commonsourceibias.n230 161.3
R244 commonsourceibias.n233 commonsourceibias.n232 161.3
R245 commonsourceibias.n234 commonsourceibias.n210 161.3
R246 commonsourceibias.n236 commonsourceibias.n235 161.3
R247 commonsourceibias.n238 commonsourceibias.n237 161.3
R248 commonsourceibias.n239 commonsourceibias.n208 161.3
R249 commonsourceibias.n241 commonsourceibias.n240 161.3
R250 commonsourceibias.n243 commonsourceibias.n242 161.3
R251 commonsourceibias.n244 commonsourceibias.n206 161.3
R252 commonsourceibias.n247 commonsourceibias.n246 161.3
R253 commonsourceibias.n248 commonsourceibias.n205 161.3
R254 commonsourceibias.n250 commonsourceibias.n249 161.3
R255 commonsourceibias.n252 commonsourceibias.n203 161.3
R256 commonsourceibias.n254 commonsourceibias.n253 161.3
R257 commonsourceibias.n255 commonsourceibias.n202 161.3
R258 commonsourceibias.n257 commonsourceibias.n256 161.3
R259 commonsourceibias.n258 commonsourceibias.n201 161.3
R260 commonsourceibias.n261 commonsourceibias.n260 161.3
R261 commonsourceibias.n262 commonsourceibias.n200 161.3
R262 commonsourceibias.n264 commonsourceibias.n263 161.3
R263 commonsourceibias.n266 commonsourceibias.n198 161.3
R264 commonsourceibias.n268 commonsourceibias.n267 161.3
R265 commonsourceibias.n269 commonsourceibias.n197 161.3
R266 commonsourceibias.n271 commonsourceibias.n270 161.3
R267 commonsourceibias.n272 commonsourceibias.n196 161.3
R268 commonsourceibias.n275 commonsourceibias.n274 161.3
R269 commonsourceibias.n276 commonsourceibias.n195 161.3
R270 commonsourceibias.n278 commonsourceibias.n277 161.3
R271 commonsourceibias.n280 commonsourceibias.n194 161.3
R272 commonsourceibias.n519 commonsourceibias.n433 161.3
R273 commonsourceibias.n517 commonsourceibias.n516 161.3
R274 commonsourceibias.n515 commonsourceibias.n434 161.3
R275 commonsourceibias.n514 commonsourceibias.n513 161.3
R276 commonsourceibias.n511 commonsourceibias.n435 161.3
R277 commonsourceibias.n510 commonsourceibias.n509 161.3
R278 commonsourceibias.n508 commonsourceibias.n436 161.3
R279 commonsourceibias.n507 commonsourceibias.n506 161.3
R280 commonsourceibias.n504 commonsourceibias.n437 161.3
R281 commonsourceibias.n502 commonsourceibias.n501 161.3
R282 commonsourceibias.n500 commonsourceibias.n438 161.3
R283 commonsourceibias.n499 commonsourceibias.n498 161.3
R284 commonsourceibias.n496 commonsourceibias.n439 161.3
R285 commonsourceibias.n495 commonsourceibias.n494 161.3
R286 commonsourceibias.n493 commonsourceibias.n440 161.3
R287 commonsourceibias.n492 commonsourceibias.n491 161.3
R288 commonsourceibias.n489 commonsourceibias.n441 161.3
R289 commonsourceibias.n487 commonsourceibias.n486 161.3
R290 commonsourceibias.n485 commonsourceibias.n442 161.3
R291 commonsourceibias.n484 commonsourceibias.n483 161.3
R292 commonsourceibias.n481 commonsourceibias.n443 161.3
R293 commonsourceibias.n480 commonsourceibias.n479 161.3
R294 commonsourceibias.n478 commonsourceibias.n477 161.3
R295 commonsourceibias.n476 commonsourceibias.n445 161.3
R296 commonsourceibias.n475 commonsourceibias.n474 161.3
R297 commonsourceibias.n473 commonsourceibias.n472 161.3
R298 commonsourceibias.n471 commonsourceibias.n447 161.3
R299 commonsourceibias.n470 commonsourceibias.n469 161.3
R300 commonsourceibias.n468 commonsourceibias.n467 161.3
R301 commonsourceibias.n466 commonsourceibias.n449 161.3
R302 commonsourceibias.n464 commonsourceibias.n463 161.3
R303 commonsourceibias.n462 commonsourceibias.n450 161.3
R304 commonsourceibias.n461 commonsourceibias.n460 161.3
R305 commonsourceibias.n458 commonsourceibias.n451 161.3
R306 commonsourceibias.n457 commonsourceibias.n456 161.3
R307 commonsourceibias.n455 commonsourceibias.n452 161.3
R308 commonsourceibias.n425 commonsourceibias.n424 161.3
R309 commonsourceibias.n422 commonsourceibias.n384 161.3
R310 commonsourceibias.n421 commonsourceibias.n420 161.3
R311 commonsourceibias.n419 commonsourceibias.n418 161.3
R312 commonsourceibias.n417 commonsourceibias.n386 161.3
R313 commonsourceibias.n416 commonsourceibias.n415 161.3
R314 commonsourceibias.n414 commonsourceibias.n413 161.3
R315 commonsourceibias.n412 commonsourceibias.n388 161.3
R316 commonsourceibias.n411 commonsourceibias.n410 161.3
R317 commonsourceibias.n409 commonsourceibias.n408 161.3
R318 commonsourceibias.n407 commonsourceibias.n390 161.3
R319 commonsourceibias.n405 commonsourceibias.n404 161.3
R320 commonsourceibias.n403 commonsourceibias.n391 161.3
R321 commonsourceibias.n402 commonsourceibias.n401 161.3
R322 commonsourceibias.n399 commonsourceibias.n392 161.3
R323 commonsourceibias.n398 commonsourceibias.n397 161.3
R324 commonsourceibias.n396 commonsourceibias.n393 161.3
R325 commonsourceibias.n531 commonsourceibias.n383 161.3
R326 commonsourceibias.n565 commonsourceibias.n374 161.3
R327 commonsourceibias.n563 commonsourceibias.n562 161.3
R328 commonsourceibias.n561 commonsourceibias.n375 161.3
R329 commonsourceibias.n560 commonsourceibias.n559 161.3
R330 commonsourceibias.n557 commonsourceibias.n376 161.3
R331 commonsourceibias.n556 commonsourceibias.n555 161.3
R332 commonsourceibias.n554 commonsourceibias.n377 161.3
R333 commonsourceibias.n553 commonsourceibias.n552 161.3
R334 commonsourceibias.n550 commonsourceibias.n378 161.3
R335 commonsourceibias.n548 commonsourceibias.n547 161.3
R336 commonsourceibias.n546 commonsourceibias.n379 161.3
R337 commonsourceibias.n545 commonsourceibias.n544 161.3
R338 commonsourceibias.n542 commonsourceibias.n380 161.3
R339 commonsourceibias.n541 commonsourceibias.n540 161.3
R340 commonsourceibias.n539 commonsourceibias.n381 161.3
R341 commonsourceibias.n538 commonsourceibias.n537 161.3
R342 commonsourceibias.n535 commonsourceibias.n382 161.3
R343 commonsourceibias.n533 commonsourceibias.n532 161.3
R344 commonsourceibias.n744 commonsourceibias.n658 161.3
R345 commonsourceibias.n742 commonsourceibias.n741 161.3
R346 commonsourceibias.n740 commonsourceibias.n659 161.3
R347 commonsourceibias.n739 commonsourceibias.n738 161.3
R348 commonsourceibias.n736 commonsourceibias.n660 161.3
R349 commonsourceibias.n735 commonsourceibias.n734 161.3
R350 commonsourceibias.n733 commonsourceibias.n661 161.3
R351 commonsourceibias.n732 commonsourceibias.n731 161.3
R352 commonsourceibias.n729 commonsourceibias.n662 161.3
R353 commonsourceibias.n727 commonsourceibias.n726 161.3
R354 commonsourceibias.n725 commonsourceibias.n663 161.3
R355 commonsourceibias.n724 commonsourceibias.n723 161.3
R356 commonsourceibias.n721 commonsourceibias.n664 161.3
R357 commonsourceibias.n720 commonsourceibias.n719 161.3
R358 commonsourceibias.n718 commonsourceibias.n665 161.3
R359 commonsourceibias.n717 commonsourceibias.n716 161.3
R360 commonsourceibias.n714 commonsourceibias.n666 161.3
R361 commonsourceibias.n712 commonsourceibias.n711 161.3
R362 commonsourceibias.n710 commonsourceibias.n667 161.3
R363 commonsourceibias.n709 commonsourceibias.n708 161.3
R364 commonsourceibias.n706 commonsourceibias.n668 161.3
R365 commonsourceibias.n705 commonsourceibias.n704 161.3
R366 commonsourceibias.n703 commonsourceibias.n702 161.3
R367 commonsourceibias.n701 commonsourceibias.n670 161.3
R368 commonsourceibias.n700 commonsourceibias.n699 161.3
R369 commonsourceibias.n698 commonsourceibias.n697 161.3
R370 commonsourceibias.n696 commonsourceibias.n672 161.3
R371 commonsourceibias.n695 commonsourceibias.n694 161.3
R372 commonsourceibias.n693 commonsourceibias.n692 161.3
R373 commonsourceibias.n691 commonsourceibias.n674 161.3
R374 commonsourceibias.n689 commonsourceibias.n688 161.3
R375 commonsourceibias.n687 commonsourceibias.n675 161.3
R376 commonsourceibias.n686 commonsourceibias.n685 161.3
R377 commonsourceibias.n683 commonsourceibias.n676 161.3
R378 commonsourceibias.n682 commonsourceibias.n681 161.3
R379 commonsourceibias.n680 commonsourceibias.n677 161.3
R380 commonsourceibias.n654 commonsourceibias.n568 161.3
R381 commonsourceibias.n652 commonsourceibias.n651 161.3
R382 commonsourceibias.n650 commonsourceibias.n569 161.3
R383 commonsourceibias.n649 commonsourceibias.n648 161.3
R384 commonsourceibias.n646 commonsourceibias.n570 161.3
R385 commonsourceibias.n645 commonsourceibias.n644 161.3
R386 commonsourceibias.n643 commonsourceibias.n571 161.3
R387 commonsourceibias.n642 commonsourceibias.n641 161.3
R388 commonsourceibias.n639 commonsourceibias.n572 161.3
R389 commonsourceibias.n637 commonsourceibias.n636 161.3
R390 commonsourceibias.n635 commonsourceibias.n573 161.3
R391 commonsourceibias.n634 commonsourceibias.n633 161.3
R392 commonsourceibias.n631 commonsourceibias.n574 161.3
R393 commonsourceibias.n630 commonsourceibias.n629 161.3
R394 commonsourceibias.n628 commonsourceibias.n575 161.3
R395 commonsourceibias.n627 commonsourceibias.n626 161.3
R396 commonsourceibias.n624 commonsourceibias.n576 161.3
R397 commonsourceibias.n622 commonsourceibias.n621 161.3
R398 commonsourceibias.n620 commonsourceibias.n577 161.3
R399 commonsourceibias.n619 commonsourceibias.n618 161.3
R400 commonsourceibias.n616 commonsourceibias.n578 161.3
R401 commonsourceibias.n615 commonsourceibias.n614 161.3
R402 commonsourceibias.n613 commonsourceibias.n612 161.3
R403 commonsourceibias.n611 commonsourceibias.n580 161.3
R404 commonsourceibias.n610 commonsourceibias.n609 161.3
R405 commonsourceibias.n608 commonsourceibias.n607 161.3
R406 commonsourceibias.n606 commonsourceibias.n582 161.3
R407 commonsourceibias.n605 commonsourceibias.n604 161.3
R408 commonsourceibias.n603 commonsourceibias.n602 161.3
R409 commonsourceibias.n601 commonsourceibias.n584 161.3
R410 commonsourceibias.n599 commonsourceibias.n598 161.3
R411 commonsourceibias.n597 commonsourceibias.n585 161.3
R412 commonsourceibias.n596 commonsourceibias.n595 161.3
R413 commonsourceibias.n593 commonsourceibias.n586 161.3
R414 commonsourceibias.n592 commonsourceibias.n591 161.3
R415 commonsourceibias.n590 commonsourceibias.n587 161.3
R416 commonsourceibias.n111 commonsourceibias.n109 81.5057
R417 commonsourceibias.n428 commonsourceibias.n426 81.5057
R418 commonsourceibias.n111 commonsourceibias.n110 80.9324
R419 commonsourceibias.n113 commonsourceibias.n112 80.9324
R420 commonsourceibias.n115 commonsourceibias.n114 80.9324
R421 commonsourceibias.n108 commonsourceibias.n107 80.9324
R422 commonsourceibias.n106 commonsourceibias.n105 80.9324
R423 commonsourceibias.n104 commonsourceibias.n103 80.9324
R424 commonsourceibias.n102 commonsourceibias.n101 80.9324
R425 commonsourceibias.n523 commonsourceibias.n522 80.9324
R426 commonsourceibias.n525 commonsourceibias.n524 80.9324
R427 commonsourceibias.n527 commonsourceibias.n526 80.9324
R428 commonsourceibias.n529 commonsourceibias.n528 80.9324
R429 commonsourceibias.n432 commonsourceibias.n431 80.9324
R430 commonsourceibias.n430 commonsourceibias.n429 80.9324
R431 commonsourceibias.n428 commonsourceibias.n427 80.9324
R432 commonsourceibias.n100 commonsourceibias.n99 80.6037
R433 commonsourceibias.n193 commonsourceibias.n192 80.6037
R434 commonsourceibias.n372 commonsourceibias.n371 80.6037
R435 commonsourceibias.n282 commonsourceibias.n281 80.6037
R436 commonsourceibias.n521 commonsourceibias.n520 80.6037
R437 commonsourceibias.n567 commonsourceibias.n566 80.6037
R438 commonsourceibias.n746 commonsourceibias.n745 80.6037
R439 commonsourceibias.n656 commonsourceibias.n655 80.6037
R440 commonsourceibias.n85 commonsourceibias.n84 56.5617
R441 commonsourceibias.n71 commonsourceibias.n70 56.5617
R442 commonsourceibias.n62 commonsourceibias.n61 56.5617
R443 commonsourceibias.n48 commonsourceibias.n47 56.5617
R444 commonsourceibias.n178 commonsourceibias.n177 56.5617
R445 commonsourceibias.n164 commonsourceibias.n163 56.5617
R446 commonsourceibias.n155 commonsourceibias.n154 56.5617
R447 commonsourceibias.n141 commonsourceibias.n140 56.5617
R448 commonsourceibias.n320 commonsourceibias.n319 56.5617
R449 commonsourceibias.n334 commonsourceibias.n333 56.5617
R450 commonsourceibias.n343 commonsourceibias.n342 56.5617
R451 commonsourceibias.n357 commonsourceibias.n356 56.5617
R452 commonsourceibias.n267 commonsourceibias.n266 56.5617
R453 commonsourceibias.n253 commonsourceibias.n252 56.5617
R454 commonsourceibias.n244 commonsourceibias.n243 56.5617
R455 commonsourceibias.n230 commonsourceibias.n229 56.5617
R456 commonsourceibias.n467 commonsourceibias.n466 56.5617
R457 commonsourceibias.n481 commonsourceibias.n480 56.5617
R458 commonsourceibias.n491 commonsourceibias.n489 56.5617
R459 commonsourceibias.n506 commonsourceibias.n504 56.5617
R460 commonsourceibias.n552 commonsourceibias.n550 56.5617
R461 commonsourceibias.n537 commonsourceibias.n535 56.5617
R462 commonsourceibias.n408 commonsourceibias.n407 56.5617
R463 commonsourceibias.n422 commonsourceibias.n421 56.5617
R464 commonsourceibias.n692 commonsourceibias.n691 56.5617
R465 commonsourceibias.n706 commonsourceibias.n705 56.5617
R466 commonsourceibias.n716 commonsourceibias.n714 56.5617
R467 commonsourceibias.n731 commonsourceibias.n729 56.5617
R468 commonsourceibias.n602 commonsourceibias.n601 56.5617
R469 commonsourceibias.n616 commonsourceibias.n615 56.5617
R470 commonsourceibias.n626 commonsourceibias.n624 56.5617
R471 commonsourceibias.n641 commonsourceibias.n639 56.5617
R472 commonsourceibias.n76 commonsourceibias.n75 56.0773
R473 commonsourceibias.n57 commonsourceibias.n56 56.0773
R474 commonsourceibias.n169 commonsourceibias.n168 56.0773
R475 commonsourceibias.n150 commonsourceibias.n149 56.0773
R476 commonsourceibias.n329 commonsourceibias.n328 56.0773
R477 commonsourceibias.n348 commonsourceibias.n347 56.0773
R478 commonsourceibias.n258 commonsourceibias.n257 56.0773
R479 commonsourceibias.n239 commonsourceibias.n238 56.0773
R480 commonsourceibias.n476 commonsourceibias.n475 56.0773
R481 commonsourceibias.n496 commonsourceibias.n495 56.0773
R482 commonsourceibias.n542 commonsourceibias.n541 56.0773
R483 commonsourceibias.n417 commonsourceibias.n416 56.0773
R484 commonsourceibias.n701 commonsourceibias.n700 56.0773
R485 commonsourceibias.n721 commonsourceibias.n720 56.0773
R486 commonsourceibias.n611 commonsourceibias.n610 56.0773
R487 commonsourceibias.n631 commonsourceibias.n630 56.0773
R488 commonsourceibias.n99 commonsourceibias.n98 55.3321
R489 commonsourceibias.n192 commonsourceibias.n191 55.3321
R490 commonsourceibias.n371 commonsourceibias.n370 55.3321
R491 commonsourceibias.n281 commonsourceibias.n280 55.3321
R492 commonsourceibias.n520 commonsourceibias.n519 55.3321
R493 commonsourceibias.n566 commonsourceibias.n565 55.3321
R494 commonsourceibias.n745 commonsourceibias.n744 55.3321
R495 commonsourceibias.n655 commonsourceibias.n654 55.3321
R496 commonsourceibias.n90 commonsourceibias.n89 55.1086
R497 commonsourceibias.n41 commonsourceibias.n31 55.1086
R498 commonsourceibias.n183 commonsourceibias.n182 55.1086
R499 commonsourceibias.n134 commonsourceibias.n124 55.1086
R500 commonsourceibias.n313 commonsourceibias.n303 55.1086
R501 commonsourceibias.n362 commonsourceibias.n361 55.1086
R502 commonsourceibias.n272 commonsourceibias.n271 55.1086
R503 commonsourceibias.n223 commonsourceibias.n213 55.1086
R504 commonsourceibias.n460 commonsourceibias.n450 55.1086
R505 commonsourceibias.n511 commonsourceibias.n510 55.1086
R506 commonsourceibias.n557 commonsourceibias.n556 55.1086
R507 commonsourceibias.n401 commonsourceibias.n391 55.1086
R508 commonsourceibias.n685 commonsourceibias.n675 55.1086
R509 commonsourceibias.n736 commonsourceibias.n735 55.1086
R510 commonsourceibias.n595 commonsourceibias.n585 55.1086
R511 commonsourceibias.n646 commonsourceibias.n645 55.1086
R512 commonsourceibias.n35 commonsourceibias.n34 47.4592
R513 commonsourceibias.n128 commonsourceibias.n127 47.4592
R514 commonsourceibias.n307 commonsourceibias.n306 47.4592
R515 commonsourceibias.n217 commonsourceibias.n216 47.4592
R516 commonsourceibias.n454 commonsourceibias.n453 47.4592
R517 commonsourceibias.n395 commonsourceibias.n394 47.4592
R518 commonsourceibias.n679 commonsourceibias.n678 47.4592
R519 commonsourceibias.n589 commonsourceibias.n588 47.4592
R520 commonsourceibias.n308 commonsourceibias.n307 44.0436
R521 commonsourceibias.n455 commonsourceibias.n454 44.0436
R522 commonsourceibias.n396 commonsourceibias.n395 44.0436
R523 commonsourceibias.n680 commonsourceibias.n679 44.0436
R524 commonsourceibias.n590 commonsourceibias.n589 44.0436
R525 commonsourceibias.n36 commonsourceibias.n35 44.0436
R526 commonsourceibias.n129 commonsourceibias.n128 44.0436
R527 commonsourceibias.n218 commonsourceibias.n217 44.0436
R528 commonsourceibias.n92 commonsourceibias.n13 42.5146
R529 commonsourceibias.n39 commonsourceibias.n38 42.5146
R530 commonsourceibias.n185 commonsourceibias.n1 42.5146
R531 commonsourceibias.n132 commonsourceibias.n131 42.5146
R532 commonsourceibias.n311 commonsourceibias.n310 42.5146
R533 commonsourceibias.n364 commonsourceibias.n285 42.5146
R534 commonsourceibias.n274 commonsourceibias.n195 42.5146
R535 commonsourceibias.n221 commonsourceibias.n220 42.5146
R536 commonsourceibias.n458 commonsourceibias.n457 42.5146
R537 commonsourceibias.n513 commonsourceibias.n434 42.5146
R538 commonsourceibias.n559 commonsourceibias.n375 42.5146
R539 commonsourceibias.n399 commonsourceibias.n398 42.5146
R540 commonsourceibias.n683 commonsourceibias.n682 42.5146
R541 commonsourceibias.n738 commonsourceibias.n659 42.5146
R542 commonsourceibias.n593 commonsourceibias.n592 42.5146
R543 commonsourceibias.n648 commonsourceibias.n569 42.5146
R544 commonsourceibias.n78 commonsourceibias.n18 41.5458
R545 commonsourceibias.n53 commonsourceibias.n52 41.5458
R546 commonsourceibias.n171 commonsourceibias.n6 41.5458
R547 commonsourceibias.n146 commonsourceibias.n145 41.5458
R548 commonsourceibias.n325 commonsourceibias.n324 41.5458
R549 commonsourceibias.n350 commonsourceibias.n290 41.5458
R550 commonsourceibias.n260 commonsourceibias.n200 41.5458
R551 commonsourceibias.n235 commonsourceibias.n234 41.5458
R552 commonsourceibias.n472 commonsourceibias.n471 41.5458
R553 commonsourceibias.n498 commonsourceibias.n438 41.5458
R554 commonsourceibias.n544 commonsourceibias.n379 41.5458
R555 commonsourceibias.n413 commonsourceibias.n412 41.5458
R556 commonsourceibias.n697 commonsourceibias.n696 41.5458
R557 commonsourceibias.n723 commonsourceibias.n663 41.5458
R558 commonsourceibias.n607 commonsourceibias.n606 41.5458
R559 commonsourceibias.n633 commonsourceibias.n573 41.5458
R560 commonsourceibias.n68 commonsourceibias.n23 40.577
R561 commonsourceibias.n64 commonsourceibias.n23 40.577
R562 commonsourceibias.n161 commonsourceibias.n11 40.577
R563 commonsourceibias.n157 commonsourceibias.n11 40.577
R564 commonsourceibias.n336 commonsourceibias.n295 40.577
R565 commonsourceibias.n340 commonsourceibias.n295 40.577
R566 commonsourceibias.n250 commonsourceibias.n205 40.577
R567 commonsourceibias.n246 commonsourceibias.n205 40.577
R568 commonsourceibias.n483 commonsourceibias.n442 40.577
R569 commonsourceibias.n487 commonsourceibias.n442 40.577
R570 commonsourceibias.n533 commonsourceibias.n383 40.577
R571 commonsourceibias.n424 commonsourceibias.n383 40.577
R572 commonsourceibias.n708 commonsourceibias.n667 40.577
R573 commonsourceibias.n712 commonsourceibias.n667 40.577
R574 commonsourceibias.n618 commonsourceibias.n577 40.577
R575 commonsourceibias.n622 commonsourceibias.n577 40.577
R576 commonsourceibias.n82 commonsourceibias.n18 39.6083
R577 commonsourceibias.n52 commonsourceibias.n51 39.6083
R578 commonsourceibias.n175 commonsourceibias.n6 39.6083
R579 commonsourceibias.n145 commonsourceibias.n144 39.6083
R580 commonsourceibias.n324 commonsourceibias.n323 39.6083
R581 commonsourceibias.n354 commonsourceibias.n290 39.6083
R582 commonsourceibias.n264 commonsourceibias.n200 39.6083
R583 commonsourceibias.n234 commonsourceibias.n233 39.6083
R584 commonsourceibias.n471 commonsourceibias.n470 39.6083
R585 commonsourceibias.n502 commonsourceibias.n438 39.6083
R586 commonsourceibias.n548 commonsourceibias.n379 39.6083
R587 commonsourceibias.n412 commonsourceibias.n411 39.6083
R588 commonsourceibias.n696 commonsourceibias.n695 39.6083
R589 commonsourceibias.n727 commonsourceibias.n663 39.6083
R590 commonsourceibias.n606 commonsourceibias.n605 39.6083
R591 commonsourceibias.n637 commonsourceibias.n573 39.6083
R592 commonsourceibias.n96 commonsourceibias.n13 38.6395
R593 commonsourceibias.n38 commonsourceibias.n33 38.6395
R594 commonsourceibias.n189 commonsourceibias.n1 38.6395
R595 commonsourceibias.n131 commonsourceibias.n126 38.6395
R596 commonsourceibias.n310 commonsourceibias.n305 38.6395
R597 commonsourceibias.n368 commonsourceibias.n285 38.6395
R598 commonsourceibias.n278 commonsourceibias.n195 38.6395
R599 commonsourceibias.n220 commonsourceibias.n215 38.6395
R600 commonsourceibias.n457 commonsourceibias.n452 38.6395
R601 commonsourceibias.n517 commonsourceibias.n434 38.6395
R602 commonsourceibias.n563 commonsourceibias.n375 38.6395
R603 commonsourceibias.n398 commonsourceibias.n393 38.6395
R604 commonsourceibias.n682 commonsourceibias.n677 38.6395
R605 commonsourceibias.n742 commonsourceibias.n659 38.6395
R606 commonsourceibias.n592 commonsourceibias.n587 38.6395
R607 commonsourceibias.n652 commonsourceibias.n569 38.6395
R608 commonsourceibias.n89 commonsourceibias.n15 26.0455
R609 commonsourceibias.n45 commonsourceibias.n31 26.0455
R610 commonsourceibias.n182 commonsourceibias.n3 26.0455
R611 commonsourceibias.n138 commonsourceibias.n124 26.0455
R612 commonsourceibias.n317 commonsourceibias.n303 26.0455
R613 commonsourceibias.n361 commonsourceibias.n287 26.0455
R614 commonsourceibias.n271 commonsourceibias.n197 26.0455
R615 commonsourceibias.n227 commonsourceibias.n213 26.0455
R616 commonsourceibias.n464 commonsourceibias.n450 26.0455
R617 commonsourceibias.n510 commonsourceibias.n436 26.0455
R618 commonsourceibias.n556 commonsourceibias.n377 26.0455
R619 commonsourceibias.n405 commonsourceibias.n391 26.0455
R620 commonsourceibias.n689 commonsourceibias.n675 26.0455
R621 commonsourceibias.n735 commonsourceibias.n661 26.0455
R622 commonsourceibias.n599 commonsourceibias.n585 26.0455
R623 commonsourceibias.n645 commonsourceibias.n571 26.0455
R624 commonsourceibias.n75 commonsourceibias.n20 25.0767
R625 commonsourceibias.n58 commonsourceibias.n57 25.0767
R626 commonsourceibias.n168 commonsourceibias.n8 25.0767
R627 commonsourceibias.n151 commonsourceibias.n150 25.0767
R628 commonsourceibias.n330 commonsourceibias.n329 25.0767
R629 commonsourceibias.n347 commonsourceibias.n292 25.0767
R630 commonsourceibias.n257 commonsourceibias.n202 25.0767
R631 commonsourceibias.n240 commonsourceibias.n239 25.0767
R632 commonsourceibias.n477 commonsourceibias.n476 25.0767
R633 commonsourceibias.n495 commonsourceibias.n440 25.0767
R634 commonsourceibias.n541 commonsourceibias.n381 25.0767
R635 commonsourceibias.n418 commonsourceibias.n417 25.0767
R636 commonsourceibias.n702 commonsourceibias.n701 25.0767
R637 commonsourceibias.n720 commonsourceibias.n665 25.0767
R638 commonsourceibias.n612 commonsourceibias.n611 25.0767
R639 commonsourceibias.n630 commonsourceibias.n575 25.0767
R640 commonsourceibias.n71 commonsourceibias.n22 24.3464
R641 commonsourceibias.n61 commonsourceibias.n25 24.3464
R642 commonsourceibias.n164 commonsourceibias.n10 24.3464
R643 commonsourceibias.n154 commonsourceibias.n118 24.3464
R644 commonsourceibias.n333 commonsourceibias.n297 24.3464
R645 commonsourceibias.n343 commonsourceibias.n294 24.3464
R646 commonsourceibias.n253 commonsourceibias.n204 24.3464
R647 commonsourceibias.n243 commonsourceibias.n207 24.3464
R648 commonsourceibias.n480 commonsourceibias.n444 24.3464
R649 commonsourceibias.n491 commonsourceibias.n490 24.3464
R650 commonsourceibias.n537 commonsourceibias.n536 24.3464
R651 commonsourceibias.n421 commonsourceibias.n385 24.3464
R652 commonsourceibias.n705 commonsourceibias.n669 24.3464
R653 commonsourceibias.n716 commonsourceibias.n715 24.3464
R654 commonsourceibias.n615 commonsourceibias.n579 24.3464
R655 commonsourceibias.n626 commonsourceibias.n625 24.3464
R656 commonsourceibias.n85 commonsourceibias.n17 23.8546
R657 commonsourceibias.n47 commonsourceibias.n46 23.8546
R658 commonsourceibias.n178 commonsourceibias.n5 23.8546
R659 commonsourceibias.n140 commonsourceibias.n139 23.8546
R660 commonsourceibias.n319 commonsourceibias.n318 23.8546
R661 commonsourceibias.n357 commonsourceibias.n289 23.8546
R662 commonsourceibias.n267 commonsourceibias.n199 23.8546
R663 commonsourceibias.n229 commonsourceibias.n228 23.8546
R664 commonsourceibias.n466 commonsourceibias.n465 23.8546
R665 commonsourceibias.n506 commonsourceibias.n505 23.8546
R666 commonsourceibias.n552 commonsourceibias.n551 23.8546
R667 commonsourceibias.n407 commonsourceibias.n406 23.8546
R668 commonsourceibias.n691 commonsourceibias.n690 23.8546
R669 commonsourceibias.n731 commonsourceibias.n730 23.8546
R670 commonsourceibias.n601 commonsourceibias.n600 23.8546
R671 commonsourceibias.n641 commonsourceibias.n640 23.8546
R672 commonsourceibias.n98 commonsourceibias.n97 17.4607
R673 commonsourceibias.n191 commonsourceibias.n190 17.4607
R674 commonsourceibias.n370 commonsourceibias.n369 17.4607
R675 commonsourceibias.n280 commonsourceibias.n279 17.4607
R676 commonsourceibias.n519 commonsourceibias.n518 17.4607
R677 commonsourceibias.n565 commonsourceibias.n564 17.4607
R678 commonsourceibias.n744 commonsourceibias.n743 17.4607
R679 commonsourceibias.n654 commonsourceibias.n653 17.4607
R680 commonsourceibias.n84 commonsourceibias.n83 16.9689
R681 commonsourceibias.n48 commonsourceibias.n29 16.9689
R682 commonsourceibias.n177 commonsourceibias.n176 16.9689
R683 commonsourceibias.n141 commonsourceibias.n122 16.9689
R684 commonsourceibias.n320 commonsourceibias.n301 16.9689
R685 commonsourceibias.n356 commonsourceibias.n355 16.9689
R686 commonsourceibias.n266 commonsourceibias.n265 16.9689
R687 commonsourceibias.n230 commonsourceibias.n211 16.9689
R688 commonsourceibias.n467 commonsourceibias.n448 16.9689
R689 commonsourceibias.n504 commonsourceibias.n503 16.9689
R690 commonsourceibias.n550 commonsourceibias.n549 16.9689
R691 commonsourceibias.n408 commonsourceibias.n389 16.9689
R692 commonsourceibias.n692 commonsourceibias.n673 16.9689
R693 commonsourceibias.n729 commonsourceibias.n728 16.9689
R694 commonsourceibias.n602 commonsourceibias.n583 16.9689
R695 commonsourceibias.n639 commonsourceibias.n638 16.9689
R696 commonsourceibias.n70 commonsourceibias.n69 16.477
R697 commonsourceibias.n63 commonsourceibias.n62 16.477
R698 commonsourceibias.n163 commonsourceibias.n162 16.477
R699 commonsourceibias.n156 commonsourceibias.n155 16.477
R700 commonsourceibias.n335 commonsourceibias.n334 16.477
R701 commonsourceibias.n342 commonsourceibias.n341 16.477
R702 commonsourceibias.n252 commonsourceibias.n251 16.477
R703 commonsourceibias.n245 commonsourceibias.n244 16.477
R704 commonsourceibias.n482 commonsourceibias.n481 16.477
R705 commonsourceibias.n489 commonsourceibias.n488 16.477
R706 commonsourceibias.n535 commonsourceibias.n534 16.477
R707 commonsourceibias.n423 commonsourceibias.n422 16.477
R708 commonsourceibias.n707 commonsourceibias.n706 16.477
R709 commonsourceibias.n714 commonsourceibias.n713 16.477
R710 commonsourceibias.n617 commonsourceibias.n616 16.477
R711 commonsourceibias.n624 commonsourceibias.n623 16.477
R712 commonsourceibias.n77 commonsourceibias.n76 15.9852
R713 commonsourceibias.n56 commonsourceibias.n27 15.9852
R714 commonsourceibias.n170 commonsourceibias.n169 15.9852
R715 commonsourceibias.n149 commonsourceibias.n120 15.9852
R716 commonsourceibias.n328 commonsourceibias.n299 15.9852
R717 commonsourceibias.n349 commonsourceibias.n348 15.9852
R718 commonsourceibias.n259 commonsourceibias.n258 15.9852
R719 commonsourceibias.n238 commonsourceibias.n209 15.9852
R720 commonsourceibias.n475 commonsourceibias.n446 15.9852
R721 commonsourceibias.n497 commonsourceibias.n496 15.9852
R722 commonsourceibias.n543 commonsourceibias.n542 15.9852
R723 commonsourceibias.n416 commonsourceibias.n387 15.9852
R724 commonsourceibias.n700 commonsourceibias.n671 15.9852
R725 commonsourceibias.n722 commonsourceibias.n721 15.9852
R726 commonsourceibias.n610 commonsourceibias.n581 15.9852
R727 commonsourceibias.n632 commonsourceibias.n631 15.9852
R728 commonsourceibias.n91 commonsourceibias.n90 15.4934
R729 commonsourceibias.n41 commonsourceibias.n40 15.4934
R730 commonsourceibias.n184 commonsourceibias.n183 15.4934
R731 commonsourceibias.n134 commonsourceibias.n133 15.4934
R732 commonsourceibias.n313 commonsourceibias.n312 15.4934
R733 commonsourceibias.n363 commonsourceibias.n362 15.4934
R734 commonsourceibias.n273 commonsourceibias.n272 15.4934
R735 commonsourceibias.n223 commonsourceibias.n222 15.4934
R736 commonsourceibias.n460 commonsourceibias.n459 15.4934
R737 commonsourceibias.n512 commonsourceibias.n511 15.4934
R738 commonsourceibias.n558 commonsourceibias.n557 15.4934
R739 commonsourceibias.n401 commonsourceibias.n400 15.4934
R740 commonsourceibias.n685 commonsourceibias.n684 15.4934
R741 commonsourceibias.n737 commonsourceibias.n736 15.4934
R742 commonsourceibias.n595 commonsourceibias.n594 15.4934
R743 commonsourceibias.n647 commonsourceibias.n646 15.4934
R744 commonsourceibias.n102 commonsourceibias.n100 13.2663
R745 commonsourceibias.n523 commonsourceibias.n521 13.2663
R746 commonsourceibias.n748 commonsourceibias.n373 10.4122
R747 commonsourceibias.n159 commonsourceibias.n116 9.50363
R748 commonsourceibias.n531 commonsourceibias.n530 9.50363
R749 commonsourceibias.n92 commonsourceibias.n91 9.09948
R750 commonsourceibias.n40 commonsourceibias.n39 9.09948
R751 commonsourceibias.n185 commonsourceibias.n184 9.09948
R752 commonsourceibias.n133 commonsourceibias.n132 9.09948
R753 commonsourceibias.n312 commonsourceibias.n311 9.09948
R754 commonsourceibias.n364 commonsourceibias.n363 9.09948
R755 commonsourceibias.n274 commonsourceibias.n273 9.09948
R756 commonsourceibias.n222 commonsourceibias.n221 9.09948
R757 commonsourceibias.n459 commonsourceibias.n458 9.09948
R758 commonsourceibias.n513 commonsourceibias.n512 9.09948
R759 commonsourceibias.n559 commonsourceibias.n558 9.09948
R760 commonsourceibias.n400 commonsourceibias.n399 9.09948
R761 commonsourceibias.n684 commonsourceibias.n683 9.09948
R762 commonsourceibias.n738 commonsourceibias.n737 9.09948
R763 commonsourceibias.n594 commonsourceibias.n593 9.09948
R764 commonsourceibias.n648 commonsourceibias.n647 9.09948
R765 commonsourceibias.n283 commonsourceibias.n193 8.79451
R766 commonsourceibias.n657 commonsourceibias.n567 8.79451
R767 commonsourceibias.n78 commonsourceibias.n77 8.60764
R768 commonsourceibias.n53 commonsourceibias.n27 8.60764
R769 commonsourceibias.n171 commonsourceibias.n170 8.60764
R770 commonsourceibias.n146 commonsourceibias.n120 8.60764
R771 commonsourceibias.n325 commonsourceibias.n299 8.60764
R772 commonsourceibias.n350 commonsourceibias.n349 8.60764
R773 commonsourceibias.n260 commonsourceibias.n259 8.60764
R774 commonsourceibias.n235 commonsourceibias.n209 8.60764
R775 commonsourceibias.n472 commonsourceibias.n446 8.60764
R776 commonsourceibias.n498 commonsourceibias.n497 8.60764
R777 commonsourceibias.n544 commonsourceibias.n543 8.60764
R778 commonsourceibias.n413 commonsourceibias.n387 8.60764
R779 commonsourceibias.n697 commonsourceibias.n671 8.60764
R780 commonsourceibias.n723 commonsourceibias.n722 8.60764
R781 commonsourceibias.n607 commonsourceibias.n581 8.60764
R782 commonsourceibias.n633 commonsourceibias.n632 8.60764
R783 commonsourceibias.n748 commonsourceibias.n747 8.46921
R784 commonsourceibias.n69 commonsourceibias.n68 8.11581
R785 commonsourceibias.n64 commonsourceibias.n63 8.11581
R786 commonsourceibias.n162 commonsourceibias.n161 8.11581
R787 commonsourceibias.n157 commonsourceibias.n156 8.11581
R788 commonsourceibias.n336 commonsourceibias.n335 8.11581
R789 commonsourceibias.n341 commonsourceibias.n340 8.11581
R790 commonsourceibias.n251 commonsourceibias.n250 8.11581
R791 commonsourceibias.n246 commonsourceibias.n245 8.11581
R792 commonsourceibias.n483 commonsourceibias.n482 8.11581
R793 commonsourceibias.n488 commonsourceibias.n487 8.11581
R794 commonsourceibias.n534 commonsourceibias.n533 8.11581
R795 commonsourceibias.n424 commonsourceibias.n423 8.11581
R796 commonsourceibias.n708 commonsourceibias.n707 8.11581
R797 commonsourceibias.n713 commonsourceibias.n712 8.11581
R798 commonsourceibias.n618 commonsourceibias.n617 8.11581
R799 commonsourceibias.n623 commonsourceibias.n622 8.11581
R800 commonsourceibias.n83 commonsourceibias.n82 7.62397
R801 commonsourceibias.n51 commonsourceibias.n29 7.62397
R802 commonsourceibias.n176 commonsourceibias.n175 7.62397
R803 commonsourceibias.n144 commonsourceibias.n122 7.62397
R804 commonsourceibias.n323 commonsourceibias.n301 7.62397
R805 commonsourceibias.n355 commonsourceibias.n354 7.62397
R806 commonsourceibias.n265 commonsourceibias.n264 7.62397
R807 commonsourceibias.n233 commonsourceibias.n211 7.62397
R808 commonsourceibias.n470 commonsourceibias.n448 7.62397
R809 commonsourceibias.n503 commonsourceibias.n502 7.62397
R810 commonsourceibias.n549 commonsourceibias.n548 7.62397
R811 commonsourceibias.n411 commonsourceibias.n389 7.62397
R812 commonsourceibias.n695 commonsourceibias.n673 7.62397
R813 commonsourceibias.n728 commonsourceibias.n727 7.62397
R814 commonsourceibias.n605 commonsourceibias.n583 7.62397
R815 commonsourceibias.n638 commonsourceibias.n637 7.62397
R816 commonsourceibias.n97 commonsourceibias.n96 7.13213
R817 commonsourceibias.n34 commonsourceibias.n33 7.13213
R818 commonsourceibias.n190 commonsourceibias.n189 7.13213
R819 commonsourceibias.n127 commonsourceibias.n126 7.13213
R820 commonsourceibias.n306 commonsourceibias.n305 7.13213
R821 commonsourceibias.n369 commonsourceibias.n368 7.13213
R822 commonsourceibias.n279 commonsourceibias.n278 7.13213
R823 commonsourceibias.n216 commonsourceibias.n215 7.13213
R824 commonsourceibias.n453 commonsourceibias.n452 7.13213
R825 commonsourceibias.n518 commonsourceibias.n517 7.13213
R826 commonsourceibias.n564 commonsourceibias.n563 7.13213
R827 commonsourceibias.n394 commonsourceibias.n393 7.13213
R828 commonsourceibias.n678 commonsourceibias.n677 7.13213
R829 commonsourceibias.n743 commonsourceibias.n742 7.13213
R830 commonsourceibias.n588 commonsourceibias.n587 7.13213
R831 commonsourceibias.n653 commonsourceibias.n652 7.13213
R832 commonsourceibias.n373 commonsourceibias.n372 5.06534
R833 commonsourceibias.n283 commonsourceibias.n282 5.06534
R834 commonsourceibias.n747 commonsourceibias.n746 5.06534
R835 commonsourceibias.n657 commonsourceibias.n656 5.06534
R836 commonsourceibias commonsourceibias.n748 4.04308
R837 commonsourceibias.n373 commonsourceibias.n283 3.72967
R838 commonsourceibias.n747 commonsourceibias.n657 3.72967
R839 commonsourceibias.n109 commonsourceibias.t31 2.82907
R840 commonsourceibias.n109 commonsourceibias.t49 2.82907
R841 commonsourceibias.n110 commonsourceibias.t3 2.82907
R842 commonsourceibias.n110 commonsourceibias.t17 2.82907
R843 commonsourceibias.n112 commonsourceibias.t47 2.82907
R844 commonsourceibias.n112 commonsourceibias.t53 2.82907
R845 commonsourceibias.n114 commonsourceibias.t25 2.82907
R846 commonsourceibias.n114 commonsourceibias.t5 2.82907
R847 commonsourceibias.n107 commonsourceibias.t51 2.82907
R848 commonsourceibias.n107 commonsourceibias.t59 2.82907
R849 commonsourceibias.n105 commonsourceibias.t1 2.82907
R850 commonsourceibias.n105 commonsourceibias.t39 2.82907
R851 commonsourceibias.n103 commonsourceibias.t43 2.82907
R852 commonsourceibias.n103 commonsourceibias.t21 2.82907
R853 commonsourceibias.n101 commonsourceibias.t37 2.82907
R854 commonsourceibias.n101 commonsourceibias.t33 2.82907
R855 commonsourceibias.n522 commonsourceibias.t7 2.82907
R856 commonsourceibias.n522 commonsourceibias.t27 2.82907
R857 commonsourceibias.n524 commonsourceibias.t55 2.82907
R858 commonsourceibias.n524 commonsourceibias.t41 2.82907
R859 commonsourceibias.n526 commonsourceibias.t29 2.82907
R860 commonsourceibias.n526 commonsourceibias.t63 2.82907
R861 commonsourceibias.n528 commonsourceibias.t61 2.82907
R862 commonsourceibias.n528 commonsourceibias.t23 2.82907
R863 commonsourceibias.n431 commonsourceibias.t11 2.82907
R864 commonsourceibias.n431 commonsourceibias.t57 2.82907
R865 commonsourceibias.n429 commonsourceibias.t45 2.82907
R866 commonsourceibias.n429 commonsourceibias.t35 2.82907
R867 commonsourceibias.n427 commonsourceibias.t19 2.82907
R868 commonsourceibias.n427 commonsourceibias.t9 2.82907
R869 commonsourceibias.n426 commonsourceibias.t15 2.82907
R870 commonsourceibias.n426 commonsourceibias.t13 2.82907
R871 commonsourceibias.n17 commonsourceibias.n15 0.738255
R872 commonsourceibias.n46 commonsourceibias.n45 0.738255
R873 commonsourceibias.n5 commonsourceibias.n3 0.738255
R874 commonsourceibias.n139 commonsourceibias.n138 0.738255
R875 commonsourceibias.n318 commonsourceibias.n317 0.738255
R876 commonsourceibias.n289 commonsourceibias.n287 0.738255
R877 commonsourceibias.n199 commonsourceibias.n197 0.738255
R878 commonsourceibias.n228 commonsourceibias.n227 0.738255
R879 commonsourceibias.n465 commonsourceibias.n464 0.738255
R880 commonsourceibias.n505 commonsourceibias.n436 0.738255
R881 commonsourceibias.n551 commonsourceibias.n377 0.738255
R882 commonsourceibias.n406 commonsourceibias.n405 0.738255
R883 commonsourceibias.n690 commonsourceibias.n689 0.738255
R884 commonsourceibias.n730 commonsourceibias.n661 0.738255
R885 commonsourceibias.n600 commonsourceibias.n599 0.738255
R886 commonsourceibias.n640 commonsourceibias.n571 0.738255
R887 commonsourceibias.n104 commonsourceibias.n102 0.573776
R888 commonsourceibias.n106 commonsourceibias.n104 0.573776
R889 commonsourceibias.n108 commonsourceibias.n106 0.573776
R890 commonsourceibias.n115 commonsourceibias.n113 0.573776
R891 commonsourceibias.n113 commonsourceibias.n111 0.573776
R892 commonsourceibias.n430 commonsourceibias.n428 0.573776
R893 commonsourceibias.n432 commonsourceibias.n430 0.573776
R894 commonsourceibias.n529 commonsourceibias.n527 0.573776
R895 commonsourceibias.n527 commonsourceibias.n525 0.573776
R896 commonsourceibias.n525 commonsourceibias.n523 0.573776
R897 commonsourceibias.n116 commonsourceibias.n108 0.287138
R898 commonsourceibias.n116 commonsourceibias.n115 0.287138
R899 commonsourceibias.n530 commonsourceibias.n432 0.287138
R900 commonsourceibias.n530 commonsourceibias.n529 0.287138
R901 commonsourceibias.n100 commonsourceibias.n12 0.285035
R902 commonsourceibias.n193 commonsourceibias.n0 0.285035
R903 commonsourceibias.n372 commonsourceibias.n284 0.285035
R904 commonsourceibias.n282 commonsourceibias.n194 0.285035
R905 commonsourceibias.n521 commonsourceibias.n433 0.285035
R906 commonsourceibias.n567 commonsourceibias.n374 0.285035
R907 commonsourceibias.n746 commonsourceibias.n658 0.285035
R908 commonsourceibias.n656 commonsourceibias.n568 0.285035
R909 commonsourceibias.n22 commonsourceibias.n20 0.246418
R910 commonsourceibias.n58 commonsourceibias.n25 0.246418
R911 commonsourceibias.n10 commonsourceibias.n8 0.246418
R912 commonsourceibias.n151 commonsourceibias.n118 0.246418
R913 commonsourceibias.n330 commonsourceibias.n297 0.246418
R914 commonsourceibias.n294 commonsourceibias.n292 0.246418
R915 commonsourceibias.n204 commonsourceibias.n202 0.246418
R916 commonsourceibias.n240 commonsourceibias.n207 0.246418
R917 commonsourceibias.n477 commonsourceibias.n444 0.246418
R918 commonsourceibias.n490 commonsourceibias.n440 0.246418
R919 commonsourceibias.n536 commonsourceibias.n381 0.246418
R920 commonsourceibias.n418 commonsourceibias.n385 0.246418
R921 commonsourceibias.n702 commonsourceibias.n669 0.246418
R922 commonsourceibias.n715 commonsourceibias.n665 0.246418
R923 commonsourceibias.n612 commonsourceibias.n579 0.246418
R924 commonsourceibias.n625 commonsourceibias.n575 0.246418
R925 commonsourceibias.n95 commonsourceibias.n12 0.189894
R926 commonsourceibias.n95 commonsourceibias.n94 0.189894
R927 commonsourceibias.n94 commonsourceibias.n93 0.189894
R928 commonsourceibias.n93 commonsourceibias.n14 0.189894
R929 commonsourceibias.n88 commonsourceibias.n14 0.189894
R930 commonsourceibias.n88 commonsourceibias.n87 0.189894
R931 commonsourceibias.n87 commonsourceibias.n86 0.189894
R932 commonsourceibias.n86 commonsourceibias.n16 0.189894
R933 commonsourceibias.n81 commonsourceibias.n16 0.189894
R934 commonsourceibias.n81 commonsourceibias.n80 0.189894
R935 commonsourceibias.n80 commonsourceibias.n79 0.189894
R936 commonsourceibias.n79 commonsourceibias.n19 0.189894
R937 commonsourceibias.n74 commonsourceibias.n19 0.189894
R938 commonsourceibias.n74 commonsourceibias.n73 0.189894
R939 commonsourceibias.n73 commonsourceibias.n72 0.189894
R940 commonsourceibias.n72 commonsourceibias.n21 0.189894
R941 commonsourceibias.n67 commonsourceibias.n21 0.189894
R942 commonsourceibias.n67 commonsourceibias.n66 0.189894
R943 commonsourceibias.n66 commonsourceibias.n65 0.189894
R944 commonsourceibias.n65 commonsourceibias.n24 0.189894
R945 commonsourceibias.n60 commonsourceibias.n24 0.189894
R946 commonsourceibias.n60 commonsourceibias.n59 0.189894
R947 commonsourceibias.n59 commonsourceibias.n26 0.189894
R948 commonsourceibias.n55 commonsourceibias.n26 0.189894
R949 commonsourceibias.n55 commonsourceibias.n54 0.189894
R950 commonsourceibias.n54 commonsourceibias.n28 0.189894
R951 commonsourceibias.n50 commonsourceibias.n28 0.189894
R952 commonsourceibias.n50 commonsourceibias.n49 0.189894
R953 commonsourceibias.n49 commonsourceibias.n30 0.189894
R954 commonsourceibias.n44 commonsourceibias.n30 0.189894
R955 commonsourceibias.n44 commonsourceibias.n43 0.189894
R956 commonsourceibias.n43 commonsourceibias.n42 0.189894
R957 commonsourceibias.n42 commonsourceibias.n32 0.189894
R958 commonsourceibias.n37 commonsourceibias.n32 0.189894
R959 commonsourceibias.n37 commonsourceibias.n36 0.189894
R960 commonsourceibias.n158 commonsourceibias.n117 0.189894
R961 commonsourceibias.n153 commonsourceibias.n117 0.189894
R962 commonsourceibias.n153 commonsourceibias.n152 0.189894
R963 commonsourceibias.n152 commonsourceibias.n119 0.189894
R964 commonsourceibias.n148 commonsourceibias.n119 0.189894
R965 commonsourceibias.n148 commonsourceibias.n147 0.189894
R966 commonsourceibias.n147 commonsourceibias.n121 0.189894
R967 commonsourceibias.n143 commonsourceibias.n121 0.189894
R968 commonsourceibias.n143 commonsourceibias.n142 0.189894
R969 commonsourceibias.n142 commonsourceibias.n123 0.189894
R970 commonsourceibias.n137 commonsourceibias.n123 0.189894
R971 commonsourceibias.n137 commonsourceibias.n136 0.189894
R972 commonsourceibias.n136 commonsourceibias.n135 0.189894
R973 commonsourceibias.n135 commonsourceibias.n125 0.189894
R974 commonsourceibias.n130 commonsourceibias.n125 0.189894
R975 commonsourceibias.n130 commonsourceibias.n129 0.189894
R976 commonsourceibias.n188 commonsourceibias.n0 0.189894
R977 commonsourceibias.n188 commonsourceibias.n187 0.189894
R978 commonsourceibias.n187 commonsourceibias.n186 0.189894
R979 commonsourceibias.n186 commonsourceibias.n2 0.189894
R980 commonsourceibias.n181 commonsourceibias.n2 0.189894
R981 commonsourceibias.n181 commonsourceibias.n180 0.189894
R982 commonsourceibias.n180 commonsourceibias.n179 0.189894
R983 commonsourceibias.n179 commonsourceibias.n4 0.189894
R984 commonsourceibias.n174 commonsourceibias.n4 0.189894
R985 commonsourceibias.n174 commonsourceibias.n173 0.189894
R986 commonsourceibias.n173 commonsourceibias.n172 0.189894
R987 commonsourceibias.n172 commonsourceibias.n7 0.189894
R988 commonsourceibias.n167 commonsourceibias.n7 0.189894
R989 commonsourceibias.n167 commonsourceibias.n166 0.189894
R990 commonsourceibias.n166 commonsourceibias.n165 0.189894
R991 commonsourceibias.n165 commonsourceibias.n9 0.189894
R992 commonsourceibias.n160 commonsourceibias.n9 0.189894
R993 commonsourceibias.n367 commonsourceibias.n284 0.189894
R994 commonsourceibias.n367 commonsourceibias.n366 0.189894
R995 commonsourceibias.n366 commonsourceibias.n365 0.189894
R996 commonsourceibias.n365 commonsourceibias.n286 0.189894
R997 commonsourceibias.n360 commonsourceibias.n286 0.189894
R998 commonsourceibias.n360 commonsourceibias.n359 0.189894
R999 commonsourceibias.n359 commonsourceibias.n358 0.189894
R1000 commonsourceibias.n358 commonsourceibias.n288 0.189894
R1001 commonsourceibias.n353 commonsourceibias.n288 0.189894
R1002 commonsourceibias.n353 commonsourceibias.n352 0.189894
R1003 commonsourceibias.n352 commonsourceibias.n351 0.189894
R1004 commonsourceibias.n351 commonsourceibias.n291 0.189894
R1005 commonsourceibias.n346 commonsourceibias.n291 0.189894
R1006 commonsourceibias.n346 commonsourceibias.n345 0.189894
R1007 commonsourceibias.n345 commonsourceibias.n344 0.189894
R1008 commonsourceibias.n344 commonsourceibias.n293 0.189894
R1009 commonsourceibias.n339 commonsourceibias.n293 0.189894
R1010 commonsourceibias.n339 commonsourceibias.n338 0.189894
R1011 commonsourceibias.n338 commonsourceibias.n337 0.189894
R1012 commonsourceibias.n337 commonsourceibias.n296 0.189894
R1013 commonsourceibias.n332 commonsourceibias.n296 0.189894
R1014 commonsourceibias.n332 commonsourceibias.n331 0.189894
R1015 commonsourceibias.n331 commonsourceibias.n298 0.189894
R1016 commonsourceibias.n327 commonsourceibias.n298 0.189894
R1017 commonsourceibias.n327 commonsourceibias.n326 0.189894
R1018 commonsourceibias.n326 commonsourceibias.n300 0.189894
R1019 commonsourceibias.n322 commonsourceibias.n300 0.189894
R1020 commonsourceibias.n322 commonsourceibias.n321 0.189894
R1021 commonsourceibias.n321 commonsourceibias.n302 0.189894
R1022 commonsourceibias.n316 commonsourceibias.n302 0.189894
R1023 commonsourceibias.n316 commonsourceibias.n315 0.189894
R1024 commonsourceibias.n315 commonsourceibias.n314 0.189894
R1025 commonsourceibias.n314 commonsourceibias.n304 0.189894
R1026 commonsourceibias.n309 commonsourceibias.n304 0.189894
R1027 commonsourceibias.n309 commonsourceibias.n308 0.189894
R1028 commonsourceibias.n277 commonsourceibias.n194 0.189894
R1029 commonsourceibias.n277 commonsourceibias.n276 0.189894
R1030 commonsourceibias.n276 commonsourceibias.n275 0.189894
R1031 commonsourceibias.n275 commonsourceibias.n196 0.189894
R1032 commonsourceibias.n270 commonsourceibias.n196 0.189894
R1033 commonsourceibias.n270 commonsourceibias.n269 0.189894
R1034 commonsourceibias.n269 commonsourceibias.n268 0.189894
R1035 commonsourceibias.n268 commonsourceibias.n198 0.189894
R1036 commonsourceibias.n263 commonsourceibias.n198 0.189894
R1037 commonsourceibias.n263 commonsourceibias.n262 0.189894
R1038 commonsourceibias.n262 commonsourceibias.n261 0.189894
R1039 commonsourceibias.n261 commonsourceibias.n201 0.189894
R1040 commonsourceibias.n256 commonsourceibias.n201 0.189894
R1041 commonsourceibias.n256 commonsourceibias.n255 0.189894
R1042 commonsourceibias.n255 commonsourceibias.n254 0.189894
R1043 commonsourceibias.n254 commonsourceibias.n203 0.189894
R1044 commonsourceibias.n249 commonsourceibias.n203 0.189894
R1045 commonsourceibias.n249 commonsourceibias.n248 0.189894
R1046 commonsourceibias.n248 commonsourceibias.n247 0.189894
R1047 commonsourceibias.n247 commonsourceibias.n206 0.189894
R1048 commonsourceibias.n242 commonsourceibias.n206 0.189894
R1049 commonsourceibias.n242 commonsourceibias.n241 0.189894
R1050 commonsourceibias.n241 commonsourceibias.n208 0.189894
R1051 commonsourceibias.n237 commonsourceibias.n208 0.189894
R1052 commonsourceibias.n237 commonsourceibias.n236 0.189894
R1053 commonsourceibias.n236 commonsourceibias.n210 0.189894
R1054 commonsourceibias.n232 commonsourceibias.n210 0.189894
R1055 commonsourceibias.n232 commonsourceibias.n231 0.189894
R1056 commonsourceibias.n231 commonsourceibias.n212 0.189894
R1057 commonsourceibias.n226 commonsourceibias.n212 0.189894
R1058 commonsourceibias.n226 commonsourceibias.n225 0.189894
R1059 commonsourceibias.n225 commonsourceibias.n224 0.189894
R1060 commonsourceibias.n224 commonsourceibias.n214 0.189894
R1061 commonsourceibias.n219 commonsourceibias.n214 0.189894
R1062 commonsourceibias.n219 commonsourceibias.n218 0.189894
R1063 commonsourceibias.n456 commonsourceibias.n455 0.189894
R1064 commonsourceibias.n456 commonsourceibias.n451 0.189894
R1065 commonsourceibias.n461 commonsourceibias.n451 0.189894
R1066 commonsourceibias.n462 commonsourceibias.n461 0.189894
R1067 commonsourceibias.n463 commonsourceibias.n462 0.189894
R1068 commonsourceibias.n463 commonsourceibias.n449 0.189894
R1069 commonsourceibias.n468 commonsourceibias.n449 0.189894
R1070 commonsourceibias.n469 commonsourceibias.n468 0.189894
R1071 commonsourceibias.n469 commonsourceibias.n447 0.189894
R1072 commonsourceibias.n473 commonsourceibias.n447 0.189894
R1073 commonsourceibias.n474 commonsourceibias.n473 0.189894
R1074 commonsourceibias.n474 commonsourceibias.n445 0.189894
R1075 commonsourceibias.n478 commonsourceibias.n445 0.189894
R1076 commonsourceibias.n479 commonsourceibias.n478 0.189894
R1077 commonsourceibias.n479 commonsourceibias.n443 0.189894
R1078 commonsourceibias.n484 commonsourceibias.n443 0.189894
R1079 commonsourceibias.n485 commonsourceibias.n484 0.189894
R1080 commonsourceibias.n486 commonsourceibias.n485 0.189894
R1081 commonsourceibias.n486 commonsourceibias.n441 0.189894
R1082 commonsourceibias.n492 commonsourceibias.n441 0.189894
R1083 commonsourceibias.n493 commonsourceibias.n492 0.189894
R1084 commonsourceibias.n494 commonsourceibias.n493 0.189894
R1085 commonsourceibias.n494 commonsourceibias.n439 0.189894
R1086 commonsourceibias.n499 commonsourceibias.n439 0.189894
R1087 commonsourceibias.n500 commonsourceibias.n499 0.189894
R1088 commonsourceibias.n501 commonsourceibias.n500 0.189894
R1089 commonsourceibias.n501 commonsourceibias.n437 0.189894
R1090 commonsourceibias.n507 commonsourceibias.n437 0.189894
R1091 commonsourceibias.n508 commonsourceibias.n507 0.189894
R1092 commonsourceibias.n509 commonsourceibias.n508 0.189894
R1093 commonsourceibias.n509 commonsourceibias.n435 0.189894
R1094 commonsourceibias.n514 commonsourceibias.n435 0.189894
R1095 commonsourceibias.n515 commonsourceibias.n514 0.189894
R1096 commonsourceibias.n516 commonsourceibias.n515 0.189894
R1097 commonsourceibias.n516 commonsourceibias.n433 0.189894
R1098 commonsourceibias.n397 commonsourceibias.n396 0.189894
R1099 commonsourceibias.n397 commonsourceibias.n392 0.189894
R1100 commonsourceibias.n402 commonsourceibias.n392 0.189894
R1101 commonsourceibias.n403 commonsourceibias.n402 0.189894
R1102 commonsourceibias.n404 commonsourceibias.n403 0.189894
R1103 commonsourceibias.n404 commonsourceibias.n390 0.189894
R1104 commonsourceibias.n409 commonsourceibias.n390 0.189894
R1105 commonsourceibias.n410 commonsourceibias.n409 0.189894
R1106 commonsourceibias.n410 commonsourceibias.n388 0.189894
R1107 commonsourceibias.n414 commonsourceibias.n388 0.189894
R1108 commonsourceibias.n415 commonsourceibias.n414 0.189894
R1109 commonsourceibias.n415 commonsourceibias.n386 0.189894
R1110 commonsourceibias.n419 commonsourceibias.n386 0.189894
R1111 commonsourceibias.n420 commonsourceibias.n419 0.189894
R1112 commonsourceibias.n420 commonsourceibias.n384 0.189894
R1113 commonsourceibias.n425 commonsourceibias.n384 0.189894
R1114 commonsourceibias.n532 commonsourceibias.n382 0.189894
R1115 commonsourceibias.n538 commonsourceibias.n382 0.189894
R1116 commonsourceibias.n539 commonsourceibias.n538 0.189894
R1117 commonsourceibias.n540 commonsourceibias.n539 0.189894
R1118 commonsourceibias.n540 commonsourceibias.n380 0.189894
R1119 commonsourceibias.n545 commonsourceibias.n380 0.189894
R1120 commonsourceibias.n546 commonsourceibias.n545 0.189894
R1121 commonsourceibias.n547 commonsourceibias.n546 0.189894
R1122 commonsourceibias.n547 commonsourceibias.n378 0.189894
R1123 commonsourceibias.n553 commonsourceibias.n378 0.189894
R1124 commonsourceibias.n554 commonsourceibias.n553 0.189894
R1125 commonsourceibias.n555 commonsourceibias.n554 0.189894
R1126 commonsourceibias.n555 commonsourceibias.n376 0.189894
R1127 commonsourceibias.n560 commonsourceibias.n376 0.189894
R1128 commonsourceibias.n561 commonsourceibias.n560 0.189894
R1129 commonsourceibias.n562 commonsourceibias.n561 0.189894
R1130 commonsourceibias.n562 commonsourceibias.n374 0.189894
R1131 commonsourceibias.n681 commonsourceibias.n680 0.189894
R1132 commonsourceibias.n681 commonsourceibias.n676 0.189894
R1133 commonsourceibias.n686 commonsourceibias.n676 0.189894
R1134 commonsourceibias.n687 commonsourceibias.n686 0.189894
R1135 commonsourceibias.n688 commonsourceibias.n687 0.189894
R1136 commonsourceibias.n688 commonsourceibias.n674 0.189894
R1137 commonsourceibias.n693 commonsourceibias.n674 0.189894
R1138 commonsourceibias.n694 commonsourceibias.n693 0.189894
R1139 commonsourceibias.n694 commonsourceibias.n672 0.189894
R1140 commonsourceibias.n698 commonsourceibias.n672 0.189894
R1141 commonsourceibias.n699 commonsourceibias.n698 0.189894
R1142 commonsourceibias.n699 commonsourceibias.n670 0.189894
R1143 commonsourceibias.n703 commonsourceibias.n670 0.189894
R1144 commonsourceibias.n704 commonsourceibias.n703 0.189894
R1145 commonsourceibias.n704 commonsourceibias.n668 0.189894
R1146 commonsourceibias.n709 commonsourceibias.n668 0.189894
R1147 commonsourceibias.n710 commonsourceibias.n709 0.189894
R1148 commonsourceibias.n711 commonsourceibias.n710 0.189894
R1149 commonsourceibias.n711 commonsourceibias.n666 0.189894
R1150 commonsourceibias.n717 commonsourceibias.n666 0.189894
R1151 commonsourceibias.n718 commonsourceibias.n717 0.189894
R1152 commonsourceibias.n719 commonsourceibias.n718 0.189894
R1153 commonsourceibias.n719 commonsourceibias.n664 0.189894
R1154 commonsourceibias.n724 commonsourceibias.n664 0.189894
R1155 commonsourceibias.n725 commonsourceibias.n724 0.189894
R1156 commonsourceibias.n726 commonsourceibias.n725 0.189894
R1157 commonsourceibias.n726 commonsourceibias.n662 0.189894
R1158 commonsourceibias.n732 commonsourceibias.n662 0.189894
R1159 commonsourceibias.n733 commonsourceibias.n732 0.189894
R1160 commonsourceibias.n734 commonsourceibias.n733 0.189894
R1161 commonsourceibias.n734 commonsourceibias.n660 0.189894
R1162 commonsourceibias.n739 commonsourceibias.n660 0.189894
R1163 commonsourceibias.n740 commonsourceibias.n739 0.189894
R1164 commonsourceibias.n741 commonsourceibias.n740 0.189894
R1165 commonsourceibias.n741 commonsourceibias.n658 0.189894
R1166 commonsourceibias.n591 commonsourceibias.n590 0.189894
R1167 commonsourceibias.n591 commonsourceibias.n586 0.189894
R1168 commonsourceibias.n596 commonsourceibias.n586 0.189894
R1169 commonsourceibias.n597 commonsourceibias.n596 0.189894
R1170 commonsourceibias.n598 commonsourceibias.n597 0.189894
R1171 commonsourceibias.n598 commonsourceibias.n584 0.189894
R1172 commonsourceibias.n603 commonsourceibias.n584 0.189894
R1173 commonsourceibias.n604 commonsourceibias.n603 0.189894
R1174 commonsourceibias.n604 commonsourceibias.n582 0.189894
R1175 commonsourceibias.n608 commonsourceibias.n582 0.189894
R1176 commonsourceibias.n609 commonsourceibias.n608 0.189894
R1177 commonsourceibias.n609 commonsourceibias.n580 0.189894
R1178 commonsourceibias.n613 commonsourceibias.n580 0.189894
R1179 commonsourceibias.n614 commonsourceibias.n613 0.189894
R1180 commonsourceibias.n614 commonsourceibias.n578 0.189894
R1181 commonsourceibias.n619 commonsourceibias.n578 0.189894
R1182 commonsourceibias.n620 commonsourceibias.n619 0.189894
R1183 commonsourceibias.n621 commonsourceibias.n620 0.189894
R1184 commonsourceibias.n621 commonsourceibias.n576 0.189894
R1185 commonsourceibias.n627 commonsourceibias.n576 0.189894
R1186 commonsourceibias.n628 commonsourceibias.n627 0.189894
R1187 commonsourceibias.n629 commonsourceibias.n628 0.189894
R1188 commonsourceibias.n629 commonsourceibias.n574 0.189894
R1189 commonsourceibias.n634 commonsourceibias.n574 0.189894
R1190 commonsourceibias.n635 commonsourceibias.n634 0.189894
R1191 commonsourceibias.n636 commonsourceibias.n635 0.189894
R1192 commonsourceibias.n636 commonsourceibias.n572 0.189894
R1193 commonsourceibias.n642 commonsourceibias.n572 0.189894
R1194 commonsourceibias.n643 commonsourceibias.n642 0.189894
R1195 commonsourceibias.n644 commonsourceibias.n643 0.189894
R1196 commonsourceibias.n644 commonsourceibias.n570 0.189894
R1197 commonsourceibias.n649 commonsourceibias.n570 0.189894
R1198 commonsourceibias.n650 commonsourceibias.n649 0.189894
R1199 commonsourceibias.n651 commonsourceibias.n650 0.189894
R1200 commonsourceibias.n651 commonsourceibias.n568 0.189894
R1201 commonsourceibias.n159 commonsourceibias.n158 0.170955
R1202 commonsourceibias.n160 commonsourceibias.n159 0.170955
R1203 commonsourceibias.n531 commonsourceibias.n425 0.170955
R1204 commonsourceibias.n532 commonsourceibias.n531 0.170955
R1205 gnd.n7060 gnd.n514 1183.27
R1206 gnd.n4357 gnd.n4043 939.716
R1207 gnd.n7538 gnd.n208 795.207
R1208 gnd.n348 gnd.n211 795.207
R1209 gnd.n1474 gnd.n1362 795.207
R1210 gnd.n5959 gnd.n1476 795.207
R1211 gnd.n6399 gnd.n1064 795.207
R1212 gnd.n4710 gnd.n1067 795.207
R1213 gnd.n4197 gnd.n4080 795.207
R1214 gnd.n4236 gnd.n2555 795.207
R1215 gnd.n3951 gnd.n2566 766.379
R1216 gnd.n3954 gnd.n3953 766.379
R1217 gnd.n3192 gnd.n3095 766.379
R1218 gnd.n3188 gnd.n3093 766.379
R1219 gnd.n4042 gnd.n2588 756.769
R1220 gnd.n3945 gnd.n3944 756.769
R1221 gnd.n3285 gnd.n3002 756.769
R1222 gnd.n3283 gnd.n3005 756.769
R1223 gnd.n6641 gnd.n767 756.769
R1224 gnd.n7061 gnd.n515 756.769
R1225 gnd.n7274 gnd.n388 756.769
R1226 gnd.n6473 gnd.n937 756.769
R1227 gnd.n7536 gnd.n213 739.952
R1228 gnd.n7427 gnd.n210 739.952
R1229 gnd.n5962 gnd.n5961 739.952
R1230 gnd.n6079 gnd.n1408 739.952
R1231 gnd.n6397 gnd.n1069 739.952
R1232 gnd.n2302 gnd.n1066 739.952
R1233 gnd.n4360 gnd.n4359 739.952
R1234 gnd.n4355 gnd.n2551 739.952
R1235 gnd.n4771 gnd.n2113 711.122
R1236 gnd.n6148 gnd.n1298 711.122
R1237 gnd.n4783 gnd.n2111 711.122
R1238 gnd.n6150 gnd.n1293 711.122
R1239 gnd.n6642 gnd.n6641 585
R1240 gnd.n6641 gnd.n6640 585
R1241 gnd.n771 gnd.n770 585
R1242 gnd.n6639 gnd.n771 585
R1243 gnd.n6637 gnd.n6636 585
R1244 gnd.n6638 gnd.n6637 585
R1245 gnd.n6635 gnd.n773 585
R1246 gnd.n773 gnd.n772 585
R1247 gnd.n6634 gnd.n6633 585
R1248 gnd.n6633 gnd.n6632 585
R1249 gnd.n778 gnd.n777 585
R1250 gnd.n6631 gnd.n778 585
R1251 gnd.n6629 gnd.n6628 585
R1252 gnd.n6630 gnd.n6629 585
R1253 gnd.n6627 gnd.n780 585
R1254 gnd.n780 gnd.n779 585
R1255 gnd.n6626 gnd.n6625 585
R1256 gnd.n6625 gnd.n6624 585
R1257 gnd.n786 gnd.n785 585
R1258 gnd.n6623 gnd.n786 585
R1259 gnd.n6621 gnd.n6620 585
R1260 gnd.n6622 gnd.n6621 585
R1261 gnd.n6619 gnd.n788 585
R1262 gnd.n788 gnd.n787 585
R1263 gnd.n6618 gnd.n6617 585
R1264 gnd.n6617 gnd.n6616 585
R1265 gnd.n794 gnd.n793 585
R1266 gnd.n6615 gnd.n794 585
R1267 gnd.n6613 gnd.n6612 585
R1268 gnd.n6614 gnd.n6613 585
R1269 gnd.n6611 gnd.n796 585
R1270 gnd.n796 gnd.n795 585
R1271 gnd.n6610 gnd.n6609 585
R1272 gnd.n6609 gnd.n6608 585
R1273 gnd.n802 gnd.n801 585
R1274 gnd.n6607 gnd.n802 585
R1275 gnd.n6605 gnd.n6604 585
R1276 gnd.n6606 gnd.n6605 585
R1277 gnd.n6603 gnd.n804 585
R1278 gnd.n804 gnd.n803 585
R1279 gnd.n6602 gnd.n6601 585
R1280 gnd.n6601 gnd.n6600 585
R1281 gnd.n810 gnd.n809 585
R1282 gnd.n6599 gnd.n810 585
R1283 gnd.n6597 gnd.n6596 585
R1284 gnd.n6598 gnd.n6597 585
R1285 gnd.n6595 gnd.n812 585
R1286 gnd.n812 gnd.n811 585
R1287 gnd.n6594 gnd.n6593 585
R1288 gnd.n6593 gnd.n6592 585
R1289 gnd.n818 gnd.n817 585
R1290 gnd.n6591 gnd.n818 585
R1291 gnd.n6589 gnd.n6588 585
R1292 gnd.n6590 gnd.n6589 585
R1293 gnd.n6587 gnd.n820 585
R1294 gnd.n820 gnd.n819 585
R1295 gnd.n6586 gnd.n6585 585
R1296 gnd.n6585 gnd.n6584 585
R1297 gnd.n826 gnd.n825 585
R1298 gnd.n6583 gnd.n826 585
R1299 gnd.n6581 gnd.n6580 585
R1300 gnd.n6582 gnd.n6581 585
R1301 gnd.n6579 gnd.n828 585
R1302 gnd.n828 gnd.n827 585
R1303 gnd.n6578 gnd.n6577 585
R1304 gnd.n6577 gnd.n6576 585
R1305 gnd.n834 gnd.n833 585
R1306 gnd.n6575 gnd.n834 585
R1307 gnd.n6573 gnd.n6572 585
R1308 gnd.n6574 gnd.n6573 585
R1309 gnd.n6571 gnd.n836 585
R1310 gnd.n836 gnd.n835 585
R1311 gnd.n6570 gnd.n6569 585
R1312 gnd.n6569 gnd.n6568 585
R1313 gnd.n842 gnd.n841 585
R1314 gnd.n6567 gnd.n842 585
R1315 gnd.n6565 gnd.n6564 585
R1316 gnd.n6566 gnd.n6565 585
R1317 gnd.n6563 gnd.n844 585
R1318 gnd.n844 gnd.n843 585
R1319 gnd.n6562 gnd.n6561 585
R1320 gnd.n6561 gnd.n6560 585
R1321 gnd.n850 gnd.n849 585
R1322 gnd.n6559 gnd.n850 585
R1323 gnd.n6557 gnd.n6556 585
R1324 gnd.n6558 gnd.n6557 585
R1325 gnd.n6555 gnd.n852 585
R1326 gnd.n852 gnd.n851 585
R1327 gnd.n6554 gnd.n6553 585
R1328 gnd.n6553 gnd.n6552 585
R1329 gnd.n858 gnd.n857 585
R1330 gnd.n6551 gnd.n858 585
R1331 gnd.n6549 gnd.n6548 585
R1332 gnd.n6550 gnd.n6549 585
R1333 gnd.n6547 gnd.n860 585
R1334 gnd.n860 gnd.n859 585
R1335 gnd.n6546 gnd.n6545 585
R1336 gnd.n6545 gnd.n6544 585
R1337 gnd.n866 gnd.n865 585
R1338 gnd.n6543 gnd.n866 585
R1339 gnd.n6541 gnd.n6540 585
R1340 gnd.n6542 gnd.n6541 585
R1341 gnd.n6539 gnd.n868 585
R1342 gnd.n868 gnd.n867 585
R1343 gnd.n6538 gnd.n6537 585
R1344 gnd.n6537 gnd.n6536 585
R1345 gnd.n874 gnd.n873 585
R1346 gnd.n6535 gnd.n874 585
R1347 gnd.n6533 gnd.n6532 585
R1348 gnd.n6534 gnd.n6533 585
R1349 gnd.n6531 gnd.n876 585
R1350 gnd.n876 gnd.n875 585
R1351 gnd.n6530 gnd.n6529 585
R1352 gnd.n6529 gnd.n6528 585
R1353 gnd.n882 gnd.n881 585
R1354 gnd.n6527 gnd.n882 585
R1355 gnd.n6525 gnd.n6524 585
R1356 gnd.n6526 gnd.n6525 585
R1357 gnd.n6523 gnd.n884 585
R1358 gnd.n884 gnd.n883 585
R1359 gnd.n6522 gnd.n6521 585
R1360 gnd.n6521 gnd.n6520 585
R1361 gnd.n890 gnd.n889 585
R1362 gnd.n6519 gnd.n890 585
R1363 gnd.n6517 gnd.n6516 585
R1364 gnd.n6518 gnd.n6517 585
R1365 gnd.n6515 gnd.n892 585
R1366 gnd.n892 gnd.n891 585
R1367 gnd.n6514 gnd.n6513 585
R1368 gnd.n6513 gnd.n6512 585
R1369 gnd.n898 gnd.n897 585
R1370 gnd.n6511 gnd.n898 585
R1371 gnd.n6509 gnd.n6508 585
R1372 gnd.n6510 gnd.n6509 585
R1373 gnd.n6507 gnd.n900 585
R1374 gnd.n900 gnd.n899 585
R1375 gnd.n6506 gnd.n6505 585
R1376 gnd.n6505 gnd.n6504 585
R1377 gnd.n906 gnd.n905 585
R1378 gnd.n6503 gnd.n906 585
R1379 gnd.n6501 gnd.n6500 585
R1380 gnd.n6502 gnd.n6501 585
R1381 gnd.n6499 gnd.n908 585
R1382 gnd.n908 gnd.n907 585
R1383 gnd.n6498 gnd.n6497 585
R1384 gnd.n6497 gnd.n6496 585
R1385 gnd.n914 gnd.n913 585
R1386 gnd.n6495 gnd.n914 585
R1387 gnd.n6493 gnd.n6492 585
R1388 gnd.n6494 gnd.n6493 585
R1389 gnd.n6491 gnd.n916 585
R1390 gnd.n916 gnd.n915 585
R1391 gnd.n6490 gnd.n6489 585
R1392 gnd.n6489 gnd.n6488 585
R1393 gnd.n922 gnd.n921 585
R1394 gnd.n6487 gnd.n922 585
R1395 gnd.n6485 gnd.n6484 585
R1396 gnd.n6486 gnd.n6485 585
R1397 gnd.n6483 gnd.n924 585
R1398 gnd.n924 gnd.n923 585
R1399 gnd.n6482 gnd.n6481 585
R1400 gnd.n6481 gnd.n6480 585
R1401 gnd.n930 gnd.n929 585
R1402 gnd.n6479 gnd.n930 585
R1403 gnd.n6477 gnd.n6476 585
R1404 gnd.n6478 gnd.n6477 585
R1405 gnd.n6475 gnd.n932 585
R1406 gnd.n932 gnd.n931 585
R1407 gnd.n768 gnd.n767 585
R1408 gnd.n767 gnd.n766 585
R1409 gnd.n6647 gnd.n6646 585
R1410 gnd.n6648 gnd.n6647 585
R1411 gnd.n765 gnd.n764 585
R1412 gnd.n6649 gnd.n765 585
R1413 gnd.n6652 gnd.n6651 585
R1414 gnd.n6651 gnd.n6650 585
R1415 gnd.n762 gnd.n761 585
R1416 gnd.n761 gnd.n760 585
R1417 gnd.n6657 gnd.n6656 585
R1418 gnd.n6658 gnd.n6657 585
R1419 gnd.n759 gnd.n758 585
R1420 gnd.n6659 gnd.n759 585
R1421 gnd.n6662 gnd.n6661 585
R1422 gnd.n6661 gnd.n6660 585
R1423 gnd.n756 gnd.n755 585
R1424 gnd.n755 gnd.n754 585
R1425 gnd.n6667 gnd.n6666 585
R1426 gnd.n6668 gnd.n6667 585
R1427 gnd.n753 gnd.n752 585
R1428 gnd.n6669 gnd.n753 585
R1429 gnd.n6672 gnd.n6671 585
R1430 gnd.n6671 gnd.n6670 585
R1431 gnd.n750 gnd.n749 585
R1432 gnd.n749 gnd.n748 585
R1433 gnd.n6677 gnd.n6676 585
R1434 gnd.n6678 gnd.n6677 585
R1435 gnd.n747 gnd.n746 585
R1436 gnd.n6679 gnd.n747 585
R1437 gnd.n6682 gnd.n6681 585
R1438 gnd.n6681 gnd.n6680 585
R1439 gnd.n744 gnd.n743 585
R1440 gnd.n743 gnd.n742 585
R1441 gnd.n6687 gnd.n6686 585
R1442 gnd.n6688 gnd.n6687 585
R1443 gnd.n741 gnd.n740 585
R1444 gnd.n6689 gnd.n741 585
R1445 gnd.n6692 gnd.n6691 585
R1446 gnd.n6691 gnd.n6690 585
R1447 gnd.n738 gnd.n737 585
R1448 gnd.n737 gnd.n736 585
R1449 gnd.n6697 gnd.n6696 585
R1450 gnd.n6698 gnd.n6697 585
R1451 gnd.n735 gnd.n734 585
R1452 gnd.n6699 gnd.n735 585
R1453 gnd.n6702 gnd.n6701 585
R1454 gnd.n6701 gnd.n6700 585
R1455 gnd.n732 gnd.n731 585
R1456 gnd.n731 gnd.n730 585
R1457 gnd.n6707 gnd.n6706 585
R1458 gnd.n6708 gnd.n6707 585
R1459 gnd.n729 gnd.n728 585
R1460 gnd.n6709 gnd.n729 585
R1461 gnd.n6712 gnd.n6711 585
R1462 gnd.n6711 gnd.n6710 585
R1463 gnd.n726 gnd.n725 585
R1464 gnd.n725 gnd.n724 585
R1465 gnd.n6717 gnd.n6716 585
R1466 gnd.n6718 gnd.n6717 585
R1467 gnd.n723 gnd.n722 585
R1468 gnd.n6719 gnd.n723 585
R1469 gnd.n6722 gnd.n6721 585
R1470 gnd.n6721 gnd.n6720 585
R1471 gnd.n720 gnd.n719 585
R1472 gnd.n719 gnd.n718 585
R1473 gnd.n6727 gnd.n6726 585
R1474 gnd.n6728 gnd.n6727 585
R1475 gnd.n717 gnd.n716 585
R1476 gnd.n6729 gnd.n717 585
R1477 gnd.n6732 gnd.n6731 585
R1478 gnd.n6731 gnd.n6730 585
R1479 gnd.n714 gnd.n713 585
R1480 gnd.n713 gnd.n712 585
R1481 gnd.n6737 gnd.n6736 585
R1482 gnd.n6738 gnd.n6737 585
R1483 gnd.n711 gnd.n710 585
R1484 gnd.n6739 gnd.n711 585
R1485 gnd.n6742 gnd.n6741 585
R1486 gnd.n6741 gnd.n6740 585
R1487 gnd.n708 gnd.n707 585
R1488 gnd.n707 gnd.n706 585
R1489 gnd.n6747 gnd.n6746 585
R1490 gnd.n6748 gnd.n6747 585
R1491 gnd.n705 gnd.n704 585
R1492 gnd.n6749 gnd.n705 585
R1493 gnd.n6752 gnd.n6751 585
R1494 gnd.n6751 gnd.n6750 585
R1495 gnd.n702 gnd.n701 585
R1496 gnd.n701 gnd.n700 585
R1497 gnd.n6757 gnd.n6756 585
R1498 gnd.n6758 gnd.n6757 585
R1499 gnd.n699 gnd.n698 585
R1500 gnd.n6759 gnd.n699 585
R1501 gnd.n6762 gnd.n6761 585
R1502 gnd.n6761 gnd.n6760 585
R1503 gnd.n696 gnd.n695 585
R1504 gnd.n695 gnd.n694 585
R1505 gnd.n6767 gnd.n6766 585
R1506 gnd.n6768 gnd.n6767 585
R1507 gnd.n693 gnd.n692 585
R1508 gnd.n6769 gnd.n693 585
R1509 gnd.n6772 gnd.n6771 585
R1510 gnd.n6771 gnd.n6770 585
R1511 gnd.n690 gnd.n689 585
R1512 gnd.n689 gnd.n688 585
R1513 gnd.n6777 gnd.n6776 585
R1514 gnd.n6778 gnd.n6777 585
R1515 gnd.n687 gnd.n686 585
R1516 gnd.n6779 gnd.n687 585
R1517 gnd.n6782 gnd.n6781 585
R1518 gnd.n6781 gnd.n6780 585
R1519 gnd.n684 gnd.n683 585
R1520 gnd.n683 gnd.n682 585
R1521 gnd.n6787 gnd.n6786 585
R1522 gnd.n6788 gnd.n6787 585
R1523 gnd.n681 gnd.n680 585
R1524 gnd.n6789 gnd.n681 585
R1525 gnd.n6792 gnd.n6791 585
R1526 gnd.n6791 gnd.n6790 585
R1527 gnd.n678 gnd.n677 585
R1528 gnd.n677 gnd.n676 585
R1529 gnd.n6797 gnd.n6796 585
R1530 gnd.n6798 gnd.n6797 585
R1531 gnd.n675 gnd.n674 585
R1532 gnd.n6799 gnd.n675 585
R1533 gnd.n6802 gnd.n6801 585
R1534 gnd.n6801 gnd.n6800 585
R1535 gnd.n672 gnd.n671 585
R1536 gnd.n671 gnd.n670 585
R1537 gnd.n6807 gnd.n6806 585
R1538 gnd.n6808 gnd.n6807 585
R1539 gnd.n669 gnd.n668 585
R1540 gnd.n6809 gnd.n669 585
R1541 gnd.n6812 gnd.n6811 585
R1542 gnd.n6811 gnd.n6810 585
R1543 gnd.n666 gnd.n665 585
R1544 gnd.n665 gnd.n664 585
R1545 gnd.n6817 gnd.n6816 585
R1546 gnd.n6818 gnd.n6817 585
R1547 gnd.n663 gnd.n662 585
R1548 gnd.n6819 gnd.n663 585
R1549 gnd.n6822 gnd.n6821 585
R1550 gnd.n6821 gnd.n6820 585
R1551 gnd.n660 gnd.n659 585
R1552 gnd.n659 gnd.n658 585
R1553 gnd.n6827 gnd.n6826 585
R1554 gnd.n6828 gnd.n6827 585
R1555 gnd.n657 gnd.n656 585
R1556 gnd.n6829 gnd.n657 585
R1557 gnd.n6832 gnd.n6831 585
R1558 gnd.n6831 gnd.n6830 585
R1559 gnd.n654 gnd.n653 585
R1560 gnd.n653 gnd.n652 585
R1561 gnd.n6837 gnd.n6836 585
R1562 gnd.n6838 gnd.n6837 585
R1563 gnd.n651 gnd.n650 585
R1564 gnd.n6839 gnd.n651 585
R1565 gnd.n6842 gnd.n6841 585
R1566 gnd.n6841 gnd.n6840 585
R1567 gnd.n648 gnd.n647 585
R1568 gnd.n647 gnd.n646 585
R1569 gnd.n6847 gnd.n6846 585
R1570 gnd.n6848 gnd.n6847 585
R1571 gnd.n645 gnd.n644 585
R1572 gnd.n6849 gnd.n645 585
R1573 gnd.n6852 gnd.n6851 585
R1574 gnd.n6851 gnd.n6850 585
R1575 gnd.n642 gnd.n641 585
R1576 gnd.n641 gnd.n640 585
R1577 gnd.n6857 gnd.n6856 585
R1578 gnd.n6858 gnd.n6857 585
R1579 gnd.n639 gnd.n638 585
R1580 gnd.n6859 gnd.n639 585
R1581 gnd.n6862 gnd.n6861 585
R1582 gnd.n6861 gnd.n6860 585
R1583 gnd.n636 gnd.n635 585
R1584 gnd.n635 gnd.n634 585
R1585 gnd.n6867 gnd.n6866 585
R1586 gnd.n6868 gnd.n6867 585
R1587 gnd.n633 gnd.n632 585
R1588 gnd.n6869 gnd.n633 585
R1589 gnd.n6872 gnd.n6871 585
R1590 gnd.n6871 gnd.n6870 585
R1591 gnd.n630 gnd.n629 585
R1592 gnd.n629 gnd.n628 585
R1593 gnd.n6877 gnd.n6876 585
R1594 gnd.n6878 gnd.n6877 585
R1595 gnd.n627 gnd.n626 585
R1596 gnd.n6879 gnd.n627 585
R1597 gnd.n6882 gnd.n6881 585
R1598 gnd.n6881 gnd.n6880 585
R1599 gnd.n624 gnd.n623 585
R1600 gnd.n623 gnd.n622 585
R1601 gnd.n6887 gnd.n6886 585
R1602 gnd.n6888 gnd.n6887 585
R1603 gnd.n621 gnd.n620 585
R1604 gnd.n6889 gnd.n621 585
R1605 gnd.n6892 gnd.n6891 585
R1606 gnd.n6891 gnd.n6890 585
R1607 gnd.n618 gnd.n617 585
R1608 gnd.n617 gnd.n616 585
R1609 gnd.n6897 gnd.n6896 585
R1610 gnd.n6898 gnd.n6897 585
R1611 gnd.n615 gnd.n614 585
R1612 gnd.n6899 gnd.n615 585
R1613 gnd.n6902 gnd.n6901 585
R1614 gnd.n6901 gnd.n6900 585
R1615 gnd.n612 gnd.n611 585
R1616 gnd.n611 gnd.n610 585
R1617 gnd.n6907 gnd.n6906 585
R1618 gnd.n6908 gnd.n6907 585
R1619 gnd.n609 gnd.n608 585
R1620 gnd.n6909 gnd.n609 585
R1621 gnd.n6912 gnd.n6911 585
R1622 gnd.n6911 gnd.n6910 585
R1623 gnd.n606 gnd.n605 585
R1624 gnd.n605 gnd.n604 585
R1625 gnd.n6917 gnd.n6916 585
R1626 gnd.n6918 gnd.n6917 585
R1627 gnd.n603 gnd.n602 585
R1628 gnd.n6919 gnd.n603 585
R1629 gnd.n6922 gnd.n6921 585
R1630 gnd.n6921 gnd.n6920 585
R1631 gnd.n600 gnd.n599 585
R1632 gnd.n599 gnd.n598 585
R1633 gnd.n6927 gnd.n6926 585
R1634 gnd.n6928 gnd.n6927 585
R1635 gnd.n597 gnd.n596 585
R1636 gnd.n6929 gnd.n597 585
R1637 gnd.n6932 gnd.n6931 585
R1638 gnd.n6931 gnd.n6930 585
R1639 gnd.n594 gnd.n593 585
R1640 gnd.n593 gnd.n592 585
R1641 gnd.n6937 gnd.n6936 585
R1642 gnd.n6938 gnd.n6937 585
R1643 gnd.n591 gnd.n590 585
R1644 gnd.n6939 gnd.n591 585
R1645 gnd.n6942 gnd.n6941 585
R1646 gnd.n6941 gnd.n6940 585
R1647 gnd.n588 gnd.n587 585
R1648 gnd.n587 gnd.n586 585
R1649 gnd.n6947 gnd.n6946 585
R1650 gnd.n6948 gnd.n6947 585
R1651 gnd.n585 gnd.n584 585
R1652 gnd.n6949 gnd.n585 585
R1653 gnd.n6952 gnd.n6951 585
R1654 gnd.n6951 gnd.n6950 585
R1655 gnd.n582 gnd.n581 585
R1656 gnd.n581 gnd.n580 585
R1657 gnd.n6957 gnd.n6956 585
R1658 gnd.n6958 gnd.n6957 585
R1659 gnd.n579 gnd.n578 585
R1660 gnd.n6959 gnd.n579 585
R1661 gnd.n6962 gnd.n6961 585
R1662 gnd.n6961 gnd.n6960 585
R1663 gnd.n576 gnd.n575 585
R1664 gnd.n575 gnd.n574 585
R1665 gnd.n6967 gnd.n6966 585
R1666 gnd.n6968 gnd.n6967 585
R1667 gnd.n573 gnd.n572 585
R1668 gnd.n6969 gnd.n573 585
R1669 gnd.n6972 gnd.n6971 585
R1670 gnd.n6971 gnd.n6970 585
R1671 gnd.n570 gnd.n569 585
R1672 gnd.n569 gnd.n568 585
R1673 gnd.n6977 gnd.n6976 585
R1674 gnd.n6978 gnd.n6977 585
R1675 gnd.n567 gnd.n566 585
R1676 gnd.n6979 gnd.n567 585
R1677 gnd.n6982 gnd.n6981 585
R1678 gnd.n6981 gnd.n6980 585
R1679 gnd.n564 gnd.n563 585
R1680 gnd.n563 gnd.n562 585
R1681 gnd.n6987 gnd.n6986 585
R1682 gnd.n6988 gnd.n6987 585
R1683 gnd.n561 gnd.n560 585
R1684 gnd.n6989 gnd.n561 585
R1685 gnd.n6992 gnd.n6991 585
R1686 gnd.n6991 gnd.n6990 585
R1687 gnd.n558 gnd.n557 585
R1688 gnd.n557 gnd.n556 585
R1689 gnd.n6997 gnd.n6996 585
R1690 gnd.n6998 gnd.n6997 585
R1691 gnd.n555 gnd.n554 585
R1692 gnd.n6999 gnd.n555 585
R1693 gnd.n7002 gnd.n7001 585
R1694 gnd.n7001 gnd.n7000 585
R1695 gnd.n552 gnd.n551 585
R1696 gnd.n551 gnd.n550 585
R1697 gnd.n7007 gnd.n7006 585
R1698 gnd.n7008 gnd.n7007 585
R1699 gnd.n549 gnd.n548 585
R1700 gnd.n7009 gnd.n549 585
R1701 gnd.n7012 gnd.n7011 585
R1702 gnd.n7011 gnd.n7010 585
R1703 gnd.n546 gnd.n545 585
R1704 gnd.n545 gnd.n544 585
R1705 gnd.n7017 gnd.n7016 585
R1706 gnd.n7018 gnd.n7017 585
R1707 gnd.n543 gnd.n542 585
R1708 gnd.n7019 gnd.n543 585
R1709 gnd.n7022 gnd.n7021 585
R1710 gnd.n7021 gnd.n7020 585
R1711 gnd.n540 gnd.n539 585
R1712 gnd.n539 gnd.n538 585
R1713 gnd.n7027 gnd.n7026 585
R1714 gnd.n7028 gnd.n7027 585
R1715 gnd.n537 gnd.n536 585
R1716 gnd.n7029 gnd.n537 585
R1717 gnd.n7032 gnd.n7031 585
R1718 gnd.n7031 gnd.n7030 585
R1719 gnd.n534 gnd.n533 585
R1720 gnd.n533 gnd.n532 585
R1721 gnd.n7037 gnd.n7036 585
R1722 gnd.n7038 gnd.n7037 585
R1723 gnd.n531 gnd.n530 585
R1724 gnd.n7039 gnd.n531 585
R1725 gnd.n7042 gnd.n7041 585
R1726 gnd.n7041 gnd.n7040 585
R1727 gnd.n528 gnd.n527 585
R1728 gnd.n527 gnd.n526 585
R1729 gnd.n7047 gnd.n7046 585
R1730 gnd.n7048 gnd.n7047 585
R1731 gnd.n525 gnd.n524 585
R1732 gnd.n7049 gnd.n525 585
R1733 gnd.n7052 gnd.n7051 585
R1734 gnd.n7051 gnd.n7050 585
R1735 gnd.n522 gnd.n521 585
R1736 gnd.n521 gnd.n520 585
R1737 gnd.n7057 gnd.n7056 585
R1738 gnd.n7058 gnd.n7057 585
R1739 gnd.n519 gnd.n518 585
R1740 gnd.n7059 gnd.n519 585
R1741 gnd.n7062 gnd.n7061 585
R1742 gnd.n7061 gnd.n7060 585
R1743 gnd.n7273 gnd.n392 585
R1744 gnd.n7273 gnd.n7272 585
R1745 gnd.n7267 gnd.n393 585
R1746 gnd.n7271 gnd.n393 585
R1747 gnd.n7269 gnd.n7268 585
R1748 gnd.n7270 gnd.n7269 585
R1749 gnd.n396 gnd.n395 585
R1750 gnd.n395 gnd.n394 585
R1751 gnd.n7262 gnd.n7261 585
R1752 gnd.n7261 gnd.n7260 585
R1753 gnd.n399 gnd.n398 585
R1754 gnd.n7259 gnd.n399 585
R1755 gnd.n7257 gnd.n7256 585
R1756 gnd.n7258 gnd.n7257 585
R1757 gnd.n402 gnd.n401 585
R1758 gnd.n401 gnd.n400 585
R1759 gnd.n7252 gnd.n7251 585
R1760 gnd.n7251 gnd.n7250 585
R1761 gnd.n405 gnd.n404 585
R1762 gnd.n7249 gnd.n405 585
R1763 gnd.n7247 gnd.n7246 585
R1764 gnd.n7248 gnd.n7247 585
R1765 gnd.n408 gnd.n407 585
R1766 gnd.n407 gnd.n406 585
R1767 gnd.n7242 gnd.n7241 585
R1768 gnd.n7241 gnd.n7240 585
R1769 gnd.n411 gnd.n410 585
R1770 gnd.n7239 gnd.n411 585
R1771 gnd.n7237 gnd.n7236 585
R1772 gnd.n7238 gnd.n7237 585
R1773 gnd.n414 gnd.n413 585
R1774 gnd.n413 gnd.n412 585
R1775 gnd.n7232 gnd.n7231 585
R1776 gnd.n7231 gnd.n7230 585
R1777 gnd.n417 gnd.n416 585
R1778 gnd.n7229 gnd.n417 585
R1779 gnd.n7227 gnd.n7226 585
R1780 gnd.n7228 gnd.n7227 585
R1781 gnd.n420 gnd.n419 585
R1782 gnd.n419 gnd.n418 585
R1783 gnd.n7222 gnd.n7221 585
R1784 gnd.n7221 gnd.n7220 585
R1785 gnd.n423 gnd.n422 585
R1786 gnd.n7219 gnd.n423 585
R1787 gnd.n7217 gnd.n7216 585
R1788 gnd.n7218 gnd.n7217 585
R1789 gnd.n426 gnd.n425 585
R1790 gnd.n425 gnd.n424 585
R1791 gnd.n7212 gnd.n7211 585
R1792 gnd.n7211 gnd.n7210 585
R1793 gnd.n429 gnd.n428 585
R1794 gnd.n7209 gnd.n429 585
R1795 gnd.n7207 gnd.n7206 585
R1796 gnd.n7208 gnd.n7207 585
R1797 gnd.n432 gnd.n431 585
R1798 gnd.n431 gnd.n430 585
R1799 gnd.n7202 gnd.n7201 585
R1800 gnd.n7201 gnd.n7200 585
R1801 gnd.n435 gnd.n434 585
R1802 gnd.n7199 gnd.n435 585
R1803 gnd.n7197 gnd.n7196 585
R1804 gnd.n7198 gnd.n7197 585
R1805 gnd.n438 gnd.n437 585
R1806 gnd.n437 gnd.n436 585
R1807 gnd.n7192 gnd.n7191 585
R1808 gnd.n7191 gnd.n7190 585
R1809 gnd.n441 gnd.n440 585
R1810 gnd.n7189 gnd.n441 585
R1811 gnd.n7187 gnd.n7186 585
R1812 gnd.n7188 gnd.n7187 585
R1813 gnd.n444 gnd.n443 585
R1814 gnd.n443 gnd.n442 585
R1815 gnd.n7182 gnd.n7181 585
R1816 gnd.n7181 gnd.n7180 585
R1817 gnd.n447 gnd.n446 585
R1818 gnd.n7179 gnd.n447 585
R1819 gnd.n7177 gnd.n7176 585
R1820 gnd.n7178 gnd.n7177 585
R1821 gnd.n450 gnd.n449 585
R1822 gnd.n449 gnd.n448 585
R1823 gnd.n7172 gnd.n7171 585
R1824 gnd.n7171 gnd.n7170 585
R1825 gnd.n453 gnd.n452 585
R1826 gnd.n7169 gnd.n453 585
R1827 gnd.n7167 gnd.n7166 585
R1828 gnd.n7168 gnd.n7167 585
R1829 gnd.n456 gnd.n455 585
R1830 gnd.n455 gnd.n454 585
R1831 gnd.n7162 gnd.n7161 585
R1832 gnd.n7161 gnd.n7160 585
R1833 gnd.n459 gnd.n458 585
R1834 gnd.n7159 gnd.n459 585
R1835 gnd.n7157 gnd.n7156 585
R1836 gnd.n7158 gnd.n7157 585
R1837 gnd.n462 gnd.n461 585
R1838 gnd.n461 gnd.n460 585
R1839 gnd.n7152 gnd.n7151 585
R1840 gnd.n7151 gnd.n7150 585
R1841 gnd.n465 gnd.n464 585
R1842 gnd.n7149 gnd.n465 585
R1843 gnd.n7147 gnd.n7146 585
R1844 gnd.n7148 gnd.n7147 585
R1845 gnd.n468 gnd.n467 585
R1846 gnd.n467 gnd.n466 585
R1847 gnd.n7142 gnd.n7141 585
R1848 gnd.n7141 gnd.n7140 585
R1849 gnd.n471 gnd.n470 585
R1850 gnd.n7139 gnd.n471 585
R1851 gnd.n7137 gnd.n7136 585
R1852 gnd.n7138 gnd.n7137 585
R1853 gnd.n474 gnd.n473 585
R1854 gnd.n473 gnd.n472 585
R1855 gnd.n7132 gnd.n7131 585
R1856 gnd.n7131 gnd.n7130 585
R1857 gnd.n477 gnd.n476 585
R1858 gnd.n7129 gnd.n477 585
R1859 gnd.n7127 gnd.n7126 585
R1860 gnd.n7128 gnd.n7127 585
R1861 gnd.n480 gnd.n479 585
R1862 gnd.n479 gnd.n478 585
R1863 gnd.n7122 gnd.n7121 585
R1864 gnd.n7121 gnd.n7120 585
R1865 gnd.n483 gnd.n482 585
R1866 gnd.n7119 gnd.n483 585
R1867 gnd.n7117 gnd.n7116 585
R1868 gnd.n7118 gnd.n7117 585
R1869 gnd.n486 gnd.n485 585
R1870 gnd.n485 gnd.n484 585
R1871 gnd.n7112 gnd.n7111 585
R1872 gnd.n7111 gnd.n7110 585
R1873 gnd.n489 gnd.n488 585
R1874 gnd.n7109 gnd.n489 585
R1875 gnd.n7107 gnd.n7106 585
R1876 gnd.n7108 gnd.n7107 585
R1877 gnd.n492 gnd.n491 585
R1878 gnd.n491 gnd.n490 585
R1879 gnd.n7102 gnd.n7101 585
R1880 gnd.n7101 gnd.n7100 585
R1881 gnd.n495 gnd.n494 585
R1882 gnd.n7099 gnd.n495 585
R1883 gnd.n7097 gnd.n7096 585
R1884 gnd.n7098 gnd.n7097 585
R1885 gnd.n498 gnd.n497 585
R1886 gnd.n497 gnd.n496 585
R1887 gnd.n7092 gnd.n7091 585
R1888 gnd.n7091 gnd.n7090 585
R1889 gnd.n501 gnd.n500 585
R1890 gnd.n7089 gnd.n501 585
R1891 gnd.n7087 gnd.n7086 585
R1892 gnd.n7088 gnd.n7087 585
R1893 gnd.n504 gnd.n503 585
R1894 gnd.n503 gnd.n502 585
R1895 gnd.n7082 gnd.n7081 585
R1896 gnd.n7081 gnd.n7080 585
R1897 gnd.n507 gnd.n506 585
R1898 gnd.n7079 gnd.n507 585
R1899 gnd.n7077 gnd.n7076 585
R1900 gnd.n7078 gnd.n7077 585
R1901 gnd.n510 gnd.n509 585
R1902 gnd.n509 gnd.n508 585
R1903 gnd.n7072 gnd.n7071 585
R1904 gnd.n7071 gnd.n7070 585
R1905 gnd.n513 gnd.n512 585
R1906 gnd.n7069 gnd.n513 585
R1907 gnd.n7067 gnd.n7066 585
R1908 gnd.n7068 gnd.n7067 585
R1909 gnd.n516 gnd.n515 585
R1910 gnd.n515 gnd.n514 585
R1911 gnd.n6400 gnd.n6399 585
R1912 gnd.n6399 gnd.n6398 585
R1913 gnd.n6401 gnd.n1060 585
R1914 gnd.n4694 gnd.n1060 585
R1915 gnd.n6403 gnd.n6402 585
R1916 gnd.n6404 gnd.n6403 585
R1917 gnd.n1045 gnd.n1044 585
R1918 gnd.n4687 gnd.n1045 585
R1919 gnd.n6412 gnd.n6411 585
R1920 gnd.n6411 gnd.n6410 585
R1921 gnd.n6413 gnd.n1040 585
R1922 gnd.n4678 gnd.n1040 585
R1923 gnd.n6415 gnd.n6414 585
R1924 gnd.n6416 gnd.n6415 585
R1925 gnd.n1025 gnd.n1024 585
R1926 gnd.n4672 gnd.n1025 585
R1927 gnd.n6424 gnd.n6423 585
R1928 gnd.n6423 gnd.n6422 585
R1929 gnd.n6425 gnd.n1020 585
R1930 gnd.n4607 gnd.n1020 585
R1931 gnd.n6427 gnd.n6426 585
R1932 gnd.n6428 gnd.n6427 585
R1933 gnd.n1005 gnd.n1004 585
R1934 gnd.n4601 gnd.n1005 585
R1935 gnd.n6436 gnd.n6435 585
R1936 gnd.n6435 gnd.n6434 585
R1937 gnd.n6437 gnd.n1000 585
R1938 gnd.n4595 gnd.n1000 585
R1939 gnd.n6439 gnd.n6438 585
R1940 gnd.n6440 gnd.n6439 585
R1941 gnd.n985 gnd.n984 585
R1942 gnd.n4624 gnd.n985 585
R1943 gnd.n6448 gnd.n6447 585
R1944 gnd.n6447 gnd.n6446 585
R1945 gnd.n6449 gnd.n980 585
R1946 gnd.n4588 gnd.n980 585
R1947 gnd.n6451 gnd.n6450 585
R1948 gnd.n6452 gnd.n6451 585
R1949 gnd.n966 gnd.n965 585
R1950 gnd.n4580 gnd.n966 585
R1951 gnd.n6460 gnd.n6459 585
R1952 gnd.n6459 gnd.n6458 585
R1953 gnd.n6461 gnd.n960 585
R1954 gnd.n4573 gnd.n960 585
R1955 gnd.n6463 gnd.n6462 585
R1956 gnd.n6464 gnd.n6463 585
R1957 gnd.n961 gnd.n959 585
R1958 gnd.n4565 gnd.n959 585
R1959 gnd.n4525 gnd.n2434 585
R1960 gnd.n4535 gnd.n2434 585
R1961 gnd.n4526 gnd.n2441 585
R1962 gnd.n2441 gnd.n2432 585
R1963 gnd.n4528 gnd.n4527 585
R1964 gnd.n4529 gnd.n4528 585
R1965 gnd.n2442 gnd.n2440 585
R1966 gnd.n4516 gnd.n2440 585
R1967 gnd.n4491 gnd.n941 585
R1968 gnd.n6471 gnd.n941 585
R1969 gnd.n4493 gnd.n4492 585
R1970 gnd.n4492 gnd.n938 585
R1971 gnd.n4494 gnd.n2453 585
R1972 gnd.n4501 gnd.n2453 585
R1973 gnd.n4496 gnd.n4495 585
R1974 gnd.n4497 gnd.n4496 585
R1975 gnd.n2459 gnd.n2458 585
R1976 gnd.n2458 gnd.n2456 585
R1977 gnd.n4468 gnd.n2466 585
R1978 gnd.n4481 gnd.n2466 585
R1979 gnd.n4469 gnd.n2476 585
R1980 gnd.n2476 gnd.n2474 585
R1981 gnd.n4471 gnd.n4470 585
R1982 gnd.n4472 gnd.n4471 585
R1983 gnd.n2477 gnd.n2475 585
R1984 gnd.n4461 gnd.n2475 585
R1985 gnd.n4426 gnd.n4425 585
R1986 gnd.n4425 gnd.n2482 585
R1987 gnd.n4427 gnd.n2489 585
R1988 gnd.n4441 gnd.n2489 585
R1989 gnd.n4428 gnd.n2501 585
R1990 gnd.n2501 gnd.n2499 585
R1991 gnd.n4430 gnd.n4429 585
R1992 gnd.n4431 gnd.n4430 585
R1993 gnd.n2502 gnd.n2500 585
R1994 gnd.n2500 gnd.n2496 585
R1995 gnd.n4403 gnd.n2510 585
R1996 gnd.n4415 gnd.n2510 585
R1997 gnd.n4404 gnd.n2520 585
R1998 gnd.n2520 gnd.n2508 585
R1999 gnd.n4406 gnd.n4405 585
R2000 gnd.n4407 gnd.n4406 585
R2001 gnd.n2521 gnd.n2519 585
R2002 gnd.n2519 gnd.n2516 585
R2003 gnd.n4383 gnd.n2527 585
R2004 gnd.n4395 gnd.n2527 585
R2005 gnd.n4384 gnd.n2538 585
R2006 gnd.n2538 gnd.n2536 585
R2007 gnd.n4386 gnd.n4385 585
R2008 gnd.n4387 gnd.n4386 585
R2009 gnd.n2539 gnd.n2537 585
R2010 gnd.n2537 gnd.n2533 585
R2011 gnd.n2560 gnd.n2546 585
R2012 gnd.n4375 gnd.n2546 585
R2013 gnd.n2558 gnd.n2556 585
R2014 gnd.n2556 gnd.n2544 585
R2015 gnd.n4366 gnd.n4365 585
R2016 gnd.n4367 gnd.n4366 585
R2017 gnd.n2557 gnd.n2555 585
R2018 gnd.n2555 gnd.n2552 585
R2019 gnd.n4237 gnd.n4236 585
R2020 gnd.n4235 gnd.n4234 585
R2021 gnd.n4233 gnd.n4232 585
R2022 gnd.n4231 gnd.n4230 585
R2023 gnd.n4229 gnd.n4228 585
R2024 gnd.n4227 gnd.n4226 585
R2025 gnd.n4225 gnd.n4224 585
R2026 gnd.n4223 gnd.n4222 585
R2027 gnd.n4221 gnd.n4220 585
R2028 gnd.n4219 gnd.n4218 585
R2029 gnd.n4217 gnd.n4216 585
R2030 gnd.n4215 gnd.n4214 585
R2031 gnd.n4213 gnd.n4212 585
R2032 gnd.n4211 gnd.n4210 585
R2033 gnd.n4209 gnd.n4208 585
R2034 gnd.n4207 gnd.n4206 585
R2035 gnd.n4205 gnd.n4204 585
R2036 gnd.n4164 gnd.n4161 585
R2037 gnd.n4200 gnd.n4080 585
R2038 gnd.n4357 gnd.n4080 585
R2039 gnd.n4711 gnd.n4710 585
R2040 gnd.n4712 gnd.n2379 585
R2041 gnd.n4713 gnd.n2375 585
R2042 gnd.n2373 gnd.n2364 585
R2043 gnd.n4720 gnd.n2363 585
R2044 gnd.n4721 gnd.n2361 585
R2045 gnd.n2360 gnd.n2353 585
R2046 gnd.n4728 gnd.n2352 585
R2047 gnd.n4729 gnd.n2351 585
R2048 gnd.n2349 gnd.n2341 585
R2049 gnd.n4736 gnd.n2340 585
R2050 gnd.n4737 gnd.n2338 585
R2051 gnd.n2337 gnd.n2330 585
R2052 gnd.n4744 gnd.n2329 585
R2053 gnd.n4745 gnd.n2328 585
R2054 gnd.n2326 gnd.n2318 585
R2055 gnd.n4752 gnd.n2317 585
R2056 gnd.n4753 gnd.n2315 585
R2057 gnd.n2314 gnd.n1064 585
R2058 gnd.n1073 gnd.n1064 585
R2059 gnd.n4697 gnd.n1067 585
R2060 gnd.n6398 gnd.n1067 585
R2061 gnd.n4696 gnd.n4695 585
R2062 gnd.n4695 gnd.n4694 585
R2063 gnd.n2382 gnd.n1059 585
R2064 gnd.n6404 gnd.n1059 585
R2065 gnd.n4686 gnd.n4685 585
R2066 gnd.n4687 gnd.n4686 585
R2067 gnd.n2386 gnd.n1048 585
R2068 gnd.n6410 gnd.n1048 585
R2069 gnd.n4680 gnd.n4679 585
R2070 gnd.n4679 gnd.n4678 585
R2071 gnd.n2388 gnd.n1038 585
R2072 gnd.n6416 gnd.n1038 585
R2073 gnd.n4610 gnd.n2391 585
R2074 gnd.n4672 gnd.n2391 585
R2075 gnd.n4611 gnd.n1028 585
R2076 gnd.n6422 gnd.n1028 585
R2077 gnd.n4612 gnd.n4608 585
R2078 gnd.n4608 gnd.n4607 585
R2079 gnd.n2410 gnd.n1018 585
R2080 gnd.n6428 gnd.n1018 585
R2081 gnd.n4616 gnd.n2409 585
R2082 gnd.n4601 gnd.n2409 585
R2083 gnd.n4617 gnd.n1008 585
R2084 gnd.n6434 gnd.n1008 585
R2085 gnd.n4618 gnd.n2408 585
R2086 gnd.n4595 gnd.n2408 585
R2087 gnd.n2405 gnd.n998 585
R2088 gnd.n6440 gnd.n998 585
R2089 gnd.n4623 gnd.n4622 585
R2090 gnd.n4624 gnd.n4623 585
R2091 gnd.n2404 gnd.n988 585
R2092 gnd.n6446 gnd.n988 585
R2093 gnd.n4587 gnd.n4586 585
R2094 gnd.n4588 gnd.n4587 585
R2095 gnd.n2413 gnd.n978 585
R2096 gnd.n6452 gnd.n978 585
R2097 gnd.n4582 gnd.n4581 585
R2098 gnd.n4581 gnd.n4580 585
R2099 gnd.n2415 gnd.n969 585
R2100 gnd.n6458 gnd.n969 585
R2101 gnd.n4572 gnd.n4571 585
R2102 gnd.n4573 gnd.n4572 585
R2103 gnd.n2418 gnd.n957 585
R2104 gnd.n6464 gnd.n957 585
R2105 gnd.n4567 gnd.n4566 585
R2106 gnd.n4566 gnd.n4565 585
R2107 gnd.n2421 gnd.n2420 585
R2108 gnd.n4535 gnd.n2421 585
R2109 gnd.n4509 gnd.n4508 585
R2110 gnd.n4508 gnd.n2432 585
R2111 gnd.n4513 gnd.n2438 585
R2112 gnd.n4529 gnd.n2438 585
R2113 gnd.n4515 gnd.n4514 585
R2114 gnd.n4516 gnd.n4515 585
R2115 gnd.n2448 gnd.n940 585
R2116 gnd.n6471 gnd.n940 585
R2117 gnd.n4504 gnd.n4503 585
R2118 gnd.n4503 gnd.n938 585
R2119 gnd.n4502 gnd.n2450 585
R2120 gnd.n4502 gnd.n4501 585
R2121 gnd.n4452 gnd.n2451 585
R2122 gnd.n4497 gnd.n2451 585
R2123 gnd.n4454 gnd.n4453 585
R2124 gnd.n4453 gnd.n2456 585
R2125 gnd.n4455 gnd.n2465 585
R2126 gnd.n4481 gnd.n2465 585
R2127 gnd.n4457 gnd.n4456 585
R2128 gnd.n4456 gnd.n2474 585
R2129 gnd.n4458 gnd.n2473 585
R2130 gnd.n4472 gnd.n2473 585
R2131 gnd.n4460 gnd.n4459 585
R2132 gnd.n4461 gnd.n4460 585
R2133 gnd.n2484 gnd.n2483 585
R2134 gnd.n2483 gnd.n2482 585
R2135 gnd.n4443 gnd.n4442 585
R2136 gnd.n4442 gnd.n4441 585
R2137 gnd.n2487 gnd.n2486 585
R2138 gnd.n2499 gnd.n2487 585
R2139 gnd.n4178 gnd.n2498 585
R2140 gnd.n4431 gnd.n2498 585
R2141 gnd.n4180 gnd.n4179 585
R2142 gnd.n4179 gnd.n2496 585
R2143 gnd.n4181 gnd.n2509 585
R2144 gnd.n4415 gnd.n2509 585
R2145 gnd.n4183 gnd.n4182 585
R2146 gnd.n4182 gnd.n2508 585
R2147 gnd.n4184 gnd.n2518 585
R2148 gnd.n4407 gnd.n2518 585
R2149 gnd.n4186 gnd.n4185 585
R2150 gnd.n4185 gnd.n2516 585
R2151 gnd.n4187 gnd.n2526 585
R2152 gnd.n4395 gnd.n2526 585
R2153 gnd.n4189 gnd.n4188 585
R2154 gnd.n4188 gnd.n2536 585
R2155 gnd.n4190 gnd.n2535 585
R2156 gnd.n4387 gnd.n2535 585
R2157 gnd.n4192 gnd.n4191 585
R2158 gnd.n4191 gnd.n2533 585
R2159 gnd.n4193 gnd.n2545 585
R2160 gnd.n4375 gnd.n2545 585
R2161 gnd.n4195 gnd.n4194 585
R2162 gnd.n4194 gnd.n2544 585
R2163 gnd.n4196 gnd.n2554 585
R2164 gnd.n4367 gnd.n2554 585
R2165 gnd.n4198 gnd.n4197 585
R2166 gnd.n4197 gnd.n2552 585
R2167 gnd.n3951 gnd.n3950 585
R2168 gnd.n3952 gnd.n3951 585
R2169 gnd.n2641 gnd.n2640 585
R2170 gnd.n2647 gnd.n2640 585
R2171 gnd.n3926 gnd.n2659 585
R2172 gnd.n2659 gnd.n2646 585
R2173 gnd.n3928 gnd.n3927 585
R2174 gnd.n3929 gnd.n3928 585
R2175 gnd.n2660 gnd.n2658 585
R2176 gnd.n2658 gnd.n2654 585
R2177 gnd.n3660 gnd.n3659 585
R2178 gnd.n3659 gnd.n3658 585
R2179 gnd.n2665 gnd.n2664 585
R2180 gnd.n3628 gnd.n2665 585
R2181 gnd.n3648 gnd.n3647 585
R2182 gnd.n3647 gnd.n3646 585
R2183 gnd.n2672 gnd.n2671 585
R2184 gnd.n3634 gnd.n2672 585
R2185 gnd.n3604 gnd.n2692 585
R2186 gnd.n2692 gnd.n2691 585
R2187 gnd.n3606 gnd.n3605 585
R2188 gnd.n3607 gnd.n3606 585
R2189 gnd.n2693 gnd.n2690 585
R2190 gnd.n2701 gnd.n2690 585
R2191 gnd.n3582 gnd.n2713 585
R2192 gnd.n2713 gnd.n2700 585
R2193 gnd.n3584 gnd.n3583 585
R2194 gnd.n3585 gnd.n3584 585
R2195 gnd.n2714 gnd.n2712 585
R2196 gnd.n2712 gnd.n2708 585
R2197 gnd.n3570 gnd.n3569 585
R2198 gnd.n3569 gnd.n3568 585
R2199 gnd.n2719 gnd.n2718 585
R2200 gnd.n2729 gnd.n2719 585
R2201 gnd.n3559 gnd.n3558 585
R2202 gnd.n3558 gnd.n3557 585
R2203 gnd.n2726 gnd.n2725 585
R2204 gnd.n3545 gnd.n2726 585
R2205 gnd.n3519 gnd.n2747 585
R2206 gnd.n2747 gnd.n2736 585
R2207 gnd.n3521 gnd.n3520 585
R2208 gnd.n3522 gnd.n3521 585
R2209 gnd.n2748 gnd.n2746 585
R2210 gnd.n2756 gnd.n2746 585
R2211 gnd.n3497 gnd.n2768 585
R2212 gnd.n2768 gnd.n2755 585
R2213 gnd.n3499 gnd.n3498 585
R2214 gnd.n3500 gnd.n3499 585
R2215 gnd.n2769 gnd.n2767 585
R2216 gnd.n2767 gnd.n2763 585
R2217 gnd.n3485 gnd.n3484 585
R2218 gnd.n3484 gnd.n3483 585
R2219 gnd.n2774 gnd.n2773 585
R2220 gnd.n2783 gnd.n2774 585
R2221 gnd.n3474 gnd.n3473 585
R2222 gnd.n3473 gnd.n3472 585
R2223 gnd.n2781 gnd.n2780 585
R2224 gnd.n3460 gnd.n2781 585
R2225 gnd.n2898 gnd.n2897 585
R2226 gnd.n2898 gnd.n2790 585
R2227 gnd.n3417 gnd.n3416 585
R2228 gnd.n3416 gnd.n3415 585
R2229 gnd.n3418 gnd.n2892 585
R2230 gnd.n2903 gnd.n2892 585
R2231 gnd.n3420 gnd.n3419 585
R2232 gnd.n3421 gnd.n3420 585
R2233 gnd.n2893 gnd.n2891 585
R2234 gnd.n2916 gnd.n2891 585
R2235 gnd.n2876 gnd.n2875 585
R2236 gnd.n2879 gnd.n2876 585
R2237 gnd.n3431 gnd.n3430 585
R2238 gnd.n3430 gnd.n3429 585
R2239 gnd.n3432 gnd.n2870 585
R2240 gnd.n3391 gnd.n2870 585
R2241 gnd.n3434 gnd.n3433 585
R2242 gnd.n3435 gnd.n3434 585
R2243 gnd.n2871 gnd.n2869 585
R2244 gnd.n2930 gnd.n2869 585
R2245 gnd.n3383 gnd.n3382 585
R2246 gnd.n3382 gnd.n3381 585
R2247 gnd.n2927 gnd.n2926 585
R2248 gnd.n3365 gnd.n2927 585
R2249 gnd.n3352 gnd.n2946 585
R2250 gnd.n2946 gnd.n2945 585
R2251 gnd.n3354 gnd.n3353 585
R2252 gnd.n3355 gnd.n3354 585
R2253 gnd.n2947 gnd.n2944 585
R2254 gnd.n2953 gnd.n2944 585
R2255 gnd.n3333 gnd.n3332 585
R2256 gnd.n3334 gnd.n3333 585
R2257 gnd.n2964 gnd.n2963 585
R2258 gnd.n2963 gnd.n2959 585
R2259 gnd.n3323 gnd.n3322 585
R2260 gnd.n3324 gnd.n3323 585
R2261 gnd.n2974 gnd.n2973 585
R2262 gnd.n2979 gnd.n2973 585
R2263 gnd.n3301 gnd.n2992 585
R2264 gnd.n2992 gnd.n2978 585
R2265 gnd.n3303 gnd.n3302 585
R2266 gnd.n3304 gnd.n3303 585
R2267 gnd.n2993 gnd.n2991 585
R2268 gnd.n2991 gnd.n2987 585
R2269 gnd.n3292 gnd.n3291 585
R2270 gnd.n3293 gnd.n3292 585
R2271 gnd.n3000 gnd.n2999 585
R2272 gnd.n3004 gnd.n2999 585
R2273 gnd.n3269 gnd.n3021 585
R2274 gnd.n3021 gnd.n3003 585
R2275 gnd.n3271 gnd.n3270 585
R2276 gnd.n3272 gnd.n3271 585
R2277 gnd.n3022 gnd.n3020 585
R2278 gnd.n3020 gnd.n3011 585
R2279 gnd.n3264 gnd.n3263 585
R2280 gnd.n3263 gnd.n3262 585
R2281 gnd.n3069 gnd.n3068 585
R2282 gnd.n3070 gnd.n3069 585
R2283 gnd.n3223 gnd.n3222 585
R2284 gnd.n3224 gnd.n3223 585
R2285 gnd.n3079 gnd.n3078 585
R2286 gnd.n3078 gnd.n3077 585
R2287 gnd.n3218 gnd.n3217 585
R2288 gnd.n3217 gnd.n3216 585
R2289 gnd.n3082 gnd.n3081 585
R2290 gnd.n3083 gnd.n3082 585
R2291 gnd.n3207 gnd.n3206 585
R2292 gnd.n3208 gnd.n3207 585
R2293 gnd.n3090 gnd.n3089 585
R2294 gnd.n3199 gnd.n3089 585
R2295 gnd.n3202 gnd.n3201 585
R2296 gnd.n3201 gnd.n3200 585
R2297 gnd.n3093 gnd.n3092 585
R2298 gnd.n3094 gnd.n3093 585
R2299 gnd.n3188 gnd.n3187 585
R2300 gnd.n3186 gnd.n3112 585
R2301 gnd.n3185 gnd.n3111 585
R2302 gnd.n3190 gnd.n3111 585
R2303 gnd.n3184 gnd.n3183 585
R2304 gnd.n3182 gnd.n3181 585
R2305 gnd.n3180 gnd.n3179 585
R2306 gnd.n3178 gnd.n3177 585
R2307 gnd.n3176 gnd.n3175 585
R2308 gnd.n3174 gnd.n3173 585
R2309 gnd.n3172 gnd.n3171 585
R2310 gnd.n3170 gnd.n3169 585
R2311 gnd.n3168 gnd.n3167 585
R2312 gnd.n3166 gnd.n3165 585
R2313 gnd.n3164 gnd.n3163 585
R2314 gnd.n3162 gnd.n3161 585
R2315 gnd.n3160 gnd.n3159 585
R2316 gnd.n3158 gnd.n3157 585
R2317 gnd.n3156 gnd.n3155 585
R2318 gnd.n3154 gnd.n3153 585
R2319 gnd.n3152 gnd.n3151 585
R2320 gnd.n3150 gnd.n3149 585
R2321 gnd.n3148 gnd.n3147 585
R2322 gnd.n3146 gnd.n3145 585
R2323 gnd.n3144 gnd.n3143 585
R2324 gnd.n3142 gnd.n3141 585
R2325 gnd.n3099 gnd.n3098 585
R2326 gnd.n3193 gnd.n3192 585
R2327 gnd.n3955 gnd.n3954 585
R2328 gnd.n3957 gnd.n3956 585
R2329 gnd.n3959 gnd.n3958 585
R2330 gnd.n3961 gnd.n3960 585
R2331 gnd.n3963 gnd.n3962 585
R2332 gnd.n3965 gnd.n3964 585
R2333 gnd.n3967 gnd.n3966 585
R2334 gnd.n3969 gnd.n3968 585
R2335 gnd.n3971 gnd.n3970 585
R2336 gnd.n3973 gnd.n3972 585
R2337 gnd.n3975 gnd.n3974 585
R2338 gnd.n3977 gnd.n3976 585
R2339 gnd.n3979 gnd.n3978 585
R2340 gnd.n3981 gnd.n3980 585
R2341 gnd.n3983 gnd.n3982 585
R2342 gnd.n3985 gnd.n3984 585
R2343 gnd.n3987 gnd.n3986 585
R2344 gnd.n3989 gnd.n3988 585
R2345 gnd.n3991 gnd.n3990 585
R2346 gnd.n3993 gnd.n3992 585
R2347 gnd.n3995 gnd.n3994 585
R2348 gnd.n3997 gnd.n3996 585
R2349 gnd.n3999 gnd.n3998 585
R2350 gnd.n4001 gnd.n4000 585
R2351 gnd.n4003 gnd.n4002 585
R2352 gnd.n4004 gnd.n2608 585
R2353 gnd.n4005 gnd.n2566 585
R2354 gnd.n4043 gnd.n2566 585
R2355 gnd.n3953 gnd.n2638 585
R2356 gnd.n3953 gnd.n3952 585
R2357 gnd.n3621 gnd.n2637 585
R2358 gnd.n2647 gnd.n2637 585
R2359 gnd.n3623 gnd.n3622 585
R2360 gnd.n3622 gnd.n2646 585
R2361 gnd.n3624 gnd.n2656 585
R2362 gnd.n3929 gnd.n2656 585
R2363 gnd.n3626 gnd.n3625 585
R2364 gnd.n3625 gnd.n2654 585
R2365 gnd.n3627 gnd.n2667 585
R2366 gnd.n3658 gnd.n2667 585
R2367 gnd.n3630 gnd.n3629 585
R2368 gnd.n3629 gnd.n3628 585
R2369 gnd.n3631 gnd.n2674 585
R2370 gnd.n3646 gnd.n2674 585
R2371 gnd.n3633 gnd.n3632 585
R2372 gnd.n3634 gnd.n3633 585
R2373 gnd.n2684 gnd.n2683 585
R2374 gnd.n2691 gnd.n2683 585
R2375 gnd.n3609 gnd.n3608 585
R2376 gnd.n3608 gnd.n3607 585
R2377 gnd.n2687 gnd.n2686 585
R2378 gnd.n2701 gnd.n2687 585
R2379 gnd.n3535 gnd.n3534 585
R2380 gnd.n3534 gnd.n2700 585
R2381 gnd.n3536 gnd.n2710 585
R2382 gnd.n3585 gnd.n2710 585
R2383 gnd.n3538 gnd.n3537 585
R2384 gnd.n3537 gnd.n2708 585
R2385 gnd.n3539 gnd.n2721 585
R2386 gnd.n3568 gnd.n2721 585
R2387 gnd.n3541 gnd.n3540 585
R2388 gnd.n3540 gnd.n2729 585
R2389 gnd.n3542 gnd.n2728 585
R2390 gnd.n3557 gnd.n2728 585
R2391 gnd.n3544 gnd.n3543 585
R2392 gnd.n3545 gnd.n3544 585
R2393 gnd.n2740 gnd.n2739 585
R2394 gnd.n2739 gnd.n2736 585
R2395 gnd.n3524 gnd.n3523 585
R2396 gnd.n3523 gnd.n3522 585
R2397 gnd.n2743 gnd.n2742 585
R2398 gnd.n2756 gnd.n2743 585
R2399 gnd.n3448 gnd.n3447 585
R2400 gnd.n3447 gnd.n2755 585
R2401 gnd.n3449 gnd.n2765 585
R2402 gnd.n3500 gnd.n2765 585
R2403 gnd.n3451 gnd.n3450 585
R2404 gnd.n3450 gnd.n2763 585
R2405 gnd.n3452 gnd.n2776 585
R2406 gnd.n3483 gnd.n2776 585
R2407 gnd.n3454 gnd.n3453 585
R2408 gnd.n3453 gnd.n2783 585
R2409 gnd.n3455 gnd.n2782 585
R2410 gnd.n3472 gnd.n2782 585
R2411 gnd.n3457 gnd.n3456 585
R2412 gnd.n3460 gnd.n3457 585
R2413 gnd.n2793 gnd.n2792 585
R2414 gnd.n2792 gnd.n2790 585
R2415 gnd.n2900 gnd.n2899 585
R2416 gnd.n3415 gnd.n2899 585
R2417 gnd.n2902 gnd.n2901 585
R2418 gnd.n2903 gnd.n2902 585
R2419 gnd.n2913 gnd.n2889 585
R2420 gnd.n3421 gnd.n2889 585
R2421 gnd.n2915 gnd.n2914 585
R2422 gnd.n2916 gnd.n2915 585
R2423 gnd.n2912 gnd.n2911 585
R2424 gnd.n2912 gnd.n2879 585
R2425 gnd.n2910 gnd.n2877 585
R2426 gnd.n3429 gnd.n2877 585
R2427 gnd.n2866 gnd.n2864 585
R2428 gnd.n3391 gnd.n2866 585
R2429 gnd.n3437 gnd.n3436 585
R2430 gnd.n3436 gnd.n3435 585
R2431 gnd.n2865 gnd.n2863 585
R2432 gnd.n2930 gnd.n2865 585
R2433 gnd.n3362 gnd.n2929 585
R2434 gnd.n3381 gnd.n2929 585
R2435 gnd.n3364 gnd.n3363 585
R2436 gnd.n3365 gnd.n3364 585
R2437 gnd.n2939 gnd.n2938 585
R2438 gnd.n2945 gnd.n2938 585
R2439 gnd.n3357 gnd.n3356 585
R2440 gnd.n3356 gnd.n3355 585
R2441 gnd.n2942 gnd.n2941 585
R2442 gnd.n2953 gnd.n2942 585
R2443 gnd.n3242 gnd.n2961 585
R2444 gnd.n3334 gnd.n2961 585
R2445 gnd.n3244 gnd.n3243 585
R2446 gnd.n3243 gnd.n2959 585
R2447 gnd.n3245 gnd.n2972 585
R2448 gnd.n3324 gnd.n2972 585
R2449 gnd.n3247 gnd.n3246 585
R2450 gnd.n3247 gnd.n2979 585
R2451 gnd.n3249 gnd.n3248 585
R2452 gnd.n3248 gnd.n2978 585
R2453 gnd.n3250 gnd.n2989 585
R2454 gnd.n3304 gnd.n2989 585
R2455 gnd.n3252 gnd.n3251 585
R2456 gnd.n3251 gnd.n2987 585
R2457 gnd.n3253 gnd.n2998 585
R2458 gnd.n3293 gnd.n2998 585
R2459 gnd.n3255 gnd.n3254 585
R2460 gnd.n3255 gnd.n3004 585
R2461 gnd.n3257 gnd.n3256 585
R2462 gnd.n3256 gnd.n3003 585
R2463 gnd.n3258 gnd.n3019 585
R2464 gnd.n3272 gnd.n3019 585
R2465 gnd.n3259 gnd.n3072 585
R2466 gnd.n3072 gnd.n3011 585
R2467 gnd.n3261 gnd.n3260 585
R2468 gnd.n3262 gnd.n3261 585
R2469 gnd.n3073 gnd.n3071 585
R2470 gnd.n3071 gnd.n3070 585
R2471 gnd.n3226 gnd.n3225 585
R2472 gnd.n3225 gnd.n3224 585
R2473 gnd.n3076 gnd.n3075 585
R2474 gnd.n3077 gnd.n3076 585
R2475 gnd.n3215 gnd.n3214 585
R2476 gnd.n3216 gnd.n3215 585
R2477 gnd.n3085 gnd.n3084 585
R2478 gnd.n3084 gnd.n3083 585
R2479 gnd.n3210 gnd.n3209 585
R2480 gnd.n3209 gnd.n3208 585
R2481 gnd.n3088 gnd.n3087 585
R2482 gnd.n3199 gnd.n3088 585
R2483 gnd.n3198 gnd.n3197 585
R2484 gnd.n3200 gnd.n3198 585
R2485 gnd.n3096 gnd.n3095 585
R2486 gnd.n3095 gnd.n3094 585
R2487 gnd.n7539 gnd.n7538 585
R2488 gnd.n7538 gnd.n7537 585
R2489 gnd.n7540 gnd.n204 585
R2490 gnd.n209 gnd.n204 585
R2491 gnd.n7542 gnd.n7541 585
R2492 gnd.n7543 gnd.n7542 585
R2493 gnd.n190 gnd.n189 585
R2494 gnd.n194 gnd.n190 585
R2495 gnd.n7551 gnd.n7550 585
R2496 gnd.n7550 gnd.n7549 585
R2497 gnd.n7552 gnd.n185 585
R2498 gnd.n191 gnd.n185 585
R2499 gnd.n7554 gnd.n7553 585
R2500 gnd.n7555 gnd.n7554 585
R2501 gnd.n170 gnd.n169 585
R2502 gnd.n174 gnd.n170 585
R2503 gnd.n7563 gnd.n7562 585
R2504 gnd.n7562 gnd.n7561 585
R2505 gnd.n7564 gnd.n165 585
R2506 gnd.n171 gnd.n165 585
R2507 gnd.n7566 gnd.n7565 585
R2508 gnd.n7567 gnd.n7566 585
R2509 gnd.n152 gnd.n151 585
R2510 gnd.n162 gnd.n152 585
R2511 gnd.n7575 gnd.n7574 585
R2512 gnd.n7574 gnd.n7573 585
R2513 gnd.n7576 gnd.n147 585
R2514 gnd.n147 gnd.n146 585
R2515 gnd.n7578 gnd.n7577 585
R2516 gnd.n7579 gnd.n7578 585
R2517 gnd.n132 gnd.n131 585
R2518 gnd.n136 gnd.n132 585
R2519 gnd.n7587 gnd.n7586 585
R2520 gnd.n7586 gnd.n7585 585
R2521 gnd.n7588 gnd.n127 585
R2522 gnd.n133 gnd.n127 585
R2523 gnd.n7590 gnd.n7589 585
R2524 gnd.n7591 gnd.n7590 585
R2525 gnd.n115 gnd.n114 585
R2526 gnd.n124 gnd.n115 585
R2527 gnd.n7599 gnd.n7598 585
R2528 gnd.n7598 gnd.n7597 585
R2529 gnd.n7600 gnd.n109 585
R2530 gnd.n109 gnd.n107 585
R2531 gnd.n7602 gnd.n7601 585
R2532 gnd.n7603 gnd.n7602 585
R2533 gnd.n110 gnd.n108 585
R2534 gnd.n7345 gnd.n108 585
R2535 gnd.n7301 gnd.n7300 585
R2536 gnd.n7300 gnd.n368 585
R2537 gnd.n7299 gnd.n91 585
R2538 gnd.n7611 gnd.n91 585
R2539 gnd.n7298 gnd.n7297 585
R2540 gnd.n7297 gnd.n7296 585
R2541 gnd.n374 gnd.n372 585
R2542 gnd.n7283 gnd.n374 585
R2543 gnd.n7289 gnd.n7288 585
R2544 gnd.n7288 gnd.n7287 585
R2545 gnd.n380 gnd.n379 585
R2546 gnd.n1597 gnd.n380 585
R2547 gnd.n1589 gnd.n1588 585
R2548 gnd.n5888 gnd.n1589 585
R2549 gnd.n5894 gnd.n5893 585
R2550 gnd.n5893 gnd.n5892 585
R2551 gnd.n5895 gnd.n1584 585
R2552 gnd.n5859 gnd.n1584 585
R2553 gnd.n5897 gnd.n5896 585
R2554 gnd.n5898 gnd.n5897 585
R2555 gnd.n1569 gnd.n1568 585
R2556 gnd.n5875 gnd.n1569 585
R2557 gnd.n5906 gnd.n5905 585
R2558 gnd.n5905 gnd.n5904 585
R2559 gnd.n5907 gnd.n1564 585
R2560 gnd.n5845 gnd.n1564 585
R2561 gnd.n5909 gnd.n5908 585
R2562 gnd.n5910 gnd.n5909 585
R2563 gnd.n1549 gnd.n1548 585
R2564 gnd.n5837 gnd.n1549 585
R2565 gnd.n5918 gnd.n5917 585
R2566 gnd.n5917 gnd.n5916 585
R2567 gnd.n5919 gnd.n1544 585
R2568 gnd.n5830 gnd.n1544 585
R2569 gnd.n5921 gnd.n5920 585
R2570 gnd.n5922 gnd.n5921 585
R2571 gnd.n1529 gnd.n1528 585
R2572 gnd.n5822 gnd.n1529 585
R2573 gnd.n5930 gnd.n5929 585
R2574 gnd.n5929 gnd.n5928 585
R2575 gnd.n5931 gnd.n1524 585
R2576 gnd.n5759 gnd.n1524 585
R2577 gnd.n5933 gnd.n5932 585
R2578 gnd.n5934 gnd.n5933 585
R2579 gnd.n1509 gnd.n1508 585
R2580 gnd.n5750 gnd.n1509 585
R2581 gnd.n5942 gnd.n5941 585
R2582 gnd.n5941 gnd.n5940 585
R2583 gnd.n5943 gnd.n1502 585
R2584 gnd.n5744 gnd.n1502 585
R2585 gnd.n5945 gnd.n5944 585
R2586 gnd.n5946 gnd.n5945 585
R2587 gnd.n1503 gnd.n1501 585
R2588 gnd.n5737 gnd.n1501 585
R2589 gnd.n1485 gnd.n1479 585
R2590 gnd.n5952 gnd.n1485 585
R2591 gnd.n5957 gnd.n1477 585
R2592 gnd.n5776 gnd.n1477 585
R2593 gnd.n5959 gnd.n5958 585
R2594 gnd.n5960 gnd.n5959 585
R2595 gnd.n1476 gnd.n1316 585
R2596 gnd.n6127 gnd.n1317 585
R2597 gnd.n6126 gnd.n1318 585
R2598 gnd.n1393 gnd.n1319 585
R2599 gnd.n6119 gnd.n1325 585
R2600 gnd.n6118 gnd.n1326 585
R2601 gnd.n1396 gnd.n1327 585
R2602 gnd.n6111 gnd.n1333 585
R2603 gnd.n6110 gnd.n1334 585
R2604 gnd.n1398 gnd.n1335 585
R2605 gnd.n6103 gnd.n1341 585
R2606 gnd.n6102 gnd.n1342 585
R2607 gnd.n1401 gnd.n1343 585
R2608 gnd.n6095 gnd.n1349 585
R2609 gnd.n6094 gnd.n1350 585
R2610 gnd.n1403 gnd.n1351 585
R2611 gnd.n6087 gnd.n1359 585
R2612 gnd.n6086 gnd.n6083 585
R2613 gnd.n1362 gnd.n1360 585
R2614 gnd.n6081 gnd.n1362 585
R2615 gnd.n349 gnd.n348 585
R2616 gnd.n7393 gnd.n344 585
R2617 gnd.n7395 gnd.n7394 585
R2618 gnd.n7397 gnd.n342 585
R2619 gnd.n7399 gnd.n7398 585
R2620 gnd.n7400 gnd.n337 585
R2621 gnd.n7402 gnd.n7401 585
R2622 gnd.n7404 gnd.n335 585
R2623 gnd.n7406 gnd.n7405 585
R2624 gnd.n7407 gnd.n330 585
R2625 gnd.n7409 gnd.n7408 585
R2626 gnd.n7411 gnd.n328 585
R2627 gnd.n7413 gnd.n7412 585
R2628 gnd.n7414 gnd.n323 585
R2629 gnd.n7416 gnd.n7415 585
R2630 gnd.n7418 gnd.n321 585
R2631 gnd.n7420 gnd.n7419 585
R2632 gnd.n7421 gnd.n319 585
R2633 gnd.n7422 gnd.n208 585
R2634 gnd.n212 gnd.n208 585
R2635 gnd.n7389 gnd.n211 585
R2636 gnd.n7537 gnd.n211 585
R2637 gnd.n7388 gnd.n7387 585
R2638 gnd.n7387 gnd.n209 585
R2639 gnd.n7386 gnd.n203 585
R2640 gnd.n7543 gnd.n203 585
R2641 gnd.n354 gnd.n353 585
R2642 gnd.n353 gnd.n194 585
R2643 gnd.n7382 gnd.n193 585
R2644 gnd.n7549 gnd.n193 585
R2645 gnd.n7381 gnd.n7380 585
R2646 gnd.n7380 gnd.n191 585
R2647 gnd.n7379 gnd.n183 585
R2648 gnd.n7555 gnd.n183 585
R2649 gnd.n357 gnd.n356 585
R2650 gnd.n356 gnd.n174 585
R2651 gnd.n7375 gnd.n173 585
R2652 gnd.n7561 gnd.n173 585
R2653 gnd.n7374 gnd.n7373 585
R2654 gnd.n7373 gnd.n171 585
R2655 gnd.n7372 gnd.n164 585
R2656 gnd.n7567 gnd.n164 585
R2657 gnd.n360 gnd.n359 585
R2658 gnd.n359 gnd.n162 585
R2659 gnd.n7368 gnd.n154 585
R2660 gnd.n7573 gnd.n154 585
R2661 gnd.n7367 gnd.n7366 585
R2662 gnd.n7366 gnd.n146 585
R2663 gnd.n7365 gnd.n145 585
R2664 gnd.n7579 gnd.n145 585
R2665 gnd.n363 gnd.n362 585
R2666 gnd.n362 gnd.n136 585
R2667 gnd.n7361 gnd.n135 585
R2668 gnd.n7585 gnd.n135 585
R2669 gnd.n7360 gnd.n7359 585
R2670 gnd.n7359 gnd.n133 585
R2671 gnd.n7358 gnd.n126 585
R2672 gnd.n7591 gnd.n126 585
R2673 gnd.n366 gnd.n365 585
R2674 gnd.n365 gnd.n124 585
R2675 gnd.n7354 gnd.n117 585
R2676 gnd.n7597 gnd.n117 585
R2677 gnd.n7353 gnd.n7352 585
R2678 gnd.n7352 gnd.n107 585
R2679 gnd.n7351 gnd.n106 585
R2680 gnd.n7603 gnd.n106 585
R2681 gnd.n7347 gnd.n7346 585
R2682 gnd.n7346 gnd.n7345 585
R2683 gnd.n88 gnd.n87 585
R2684 gnd.n368 gnd.n88 585
R2685 gnd.n7613 gnd.n7612 585
R2686 gnd.n7612 gnd.n7611 585
R2687 gnd.n7614 gnd.n86 585
R2688 gnd.n7296 gnd.n86 585
R2689 gnd.n7282 gnd.n85 585
R2690 gnd.n7283 gnd.n7282 585
R2691 gnd.n5863 gnd.n383 585
R2692 gnd.n7287 gnd.n383 585
R2693 gnd.n5862 gnd.n5861 585
R2694 gnd.n5861 gnd.n1597 585
R2695 gnd.n5867 gnd.n1596 585
R2696 gnd.n5888 gnd.n1596 585
R2697 gnd.n5868 gnd.n1592 585
R2698 gnd.n5892 gnd.n1592 585
R2699 gnd.n5869 gnd.n5860 585
R2700 gnd.n5860 gnd.n5859 585
R2701 gnd.n1606 gnd.n1582 585
R2702 gnd.n5898 gnd.n1582 585
R2703 gnd.n5874 gnd.n5873 585
R2704 gnd.n5875 gnd.n5874 585
R2705 gnd.n1605 gnd.n1572 585
R2706 gnd.n5904 gnd.n1572 585
R2707 gnd.n5844 gnd.n5843 585
R2708 gnd.n5845 gnd.n5844 585
R2709 gnd.n1610 gnd.n1562 585
R2710 gnd.n5910 gnd.n1562 585
R2711 gnd.n5839 gnd.n5838 585
R2712 gnd.n5838 gnd.n5837 585
R2713 gnd.n1612 gnd.n1552 585
R2714 gnd.n5916 gnd.n1552 585
R2715 gnd.n5829 gnd.n5828 585
R2716 gnd.n5830 gnd.n5829 585
R2717 gnd.n1615 gnd.n1542 585
R2718 gnd.n5922 gnd.n1542 585
R2719 gnd.n5824 gnd.n5823 585
R2720 gnd.n5823 gnd.n5822 585
R2721 gnd.n1617 gnd.n1532 585
R2722 gnd.n5928 gnd.n1532 585
R2723 gnd.n5762 gnd.n5760 585
R2724 gnd.n5760 gnd.n5759 585
R2725 gnd.n5763 gnd.n1522 585
R2726 gnd.n5934 gnd.n1522 585
R2727 gnd.n5764 gnd.n5742 585
R2728 gnd.n5750 gnd.n5742 585
R2729 gnd.n5740 gnd.n1512 585
R2730 gnd.n5940 gnd.n1512 585
R2731 gnd.n5768 gnd.n5739 585
R2732 gnd.n5744 gnd.n5739 585
R2733 gnd.n5769 gnd.n1499 585
R2734 gnd.n5946 gnd.n1499 585
R2735 gnd.n5770 gnd.n5738 585
R2736 gnd.n5738 gnd.n5737 585
R2737 gnd.n1634 gnd.n1483 585
R2738 gnd.n5952 gnd.n1483 585
R2739 gnd.n5775 gnd.n5774 585
R2740 gnd.n5776 gnd.n5775 585
R2741 gnd.n1633 gnd.n1474 585
R2742 gnd.n5960 gnd.n1474 585
R2743 gnd.n3938 gnd.n2588 585
R2744 gnd.n2588 gnd.n2565 585
R2745 gnd.n3939 gnd.n2649 585
R2746 gnd.n2649 gnd.n2639 585
R2747 gnd.n3941 gnd.n3940 585
R2748 gnd.n3942 gnd.n3941 585
R2749 gnd.n2650 gnd.n2648 585
R2750 gnd.n2657 gnd.n2648 585
R2751 gnd.n3932 gnd.n3931 585
R2752 gnd.n3931 gnd.n3930 585
R2753 gnd.n2653 gnd.n2652 585
R2754 gnd.n3657 gnd.n2653 585
R2755 gnd.n3642 gnd.n2676 585
R2756 gnd.n2676 gnd.n2666 585
R2757 gnd.n3644 gnd.n3643 585
R2758 gnd.n3645 gnd.n3644 585
R2759 gnd.n2677 gnd.n2675 585
R2760 gnd.n2675 gnd.n2673 585
R2761 gnd.n3637 gnd.n3636 585
R2762 gnd.n3636 gnd.n3635 585
R2763 gnd.n2680 gnd.n2679 585
R2764 gnd.n2689 gnd.n2680 585
R2765 gnd.n3593 gnd.n2703 585
R2766 gnd.n2703 gnd.n2688 585
R2767 gnd.n3595 gnd.n3594 585
R2768 gnd.n3596 gnd.n3595 585
R2769 gnd.n2704 gnd.n2702 585
R2770 gnd.n2711 gnd.n2702 585
R2771 gnd.n3588 gnd.n3587 585
R2772 gnd.n3587 gnd.n3586 585
R2773 gnd.n2707 gnd.n2706 585
R2774 gnd.n3567 gnd.n2707 585
R2775 gnd.n3553 gnd.n2731 585
R2776 gnd.n2731 gnd.n2720 585
R2777 gnd.n3555 gnd.n3554 585
R2778 gnd.n3556 gnd.n3555 585
R2779 gnd.n2732 gnd.n2730 585
R2780 gnd.n2730 gnd.n2727 585
R2781 gnd.n3548 gnd.n3547 585
R2782 gnd.n3547 gnd.n3546 585
R2783 gnd.n2735 gnd.n2734 585
R2784 gnd.n2745 gnd.n2735 585
R2785 gnd.n3508 gnd.n2758 585
R2786 gnd.n2758 gnd.n2744 585
R2787 gnd.n3510 gnd.n3509 585
R2788 gnd.n3511 gnd.n3510 585
R2789 gnd.n2759 gnd.n2757 585
R2790 gnd.n2766 gnd.n2757 585
R2791 gnd.n3503 gnd.n3502 585
R2792 gnd.n3502 gnd.n3501 585
R2793 gnd.n2762 gnd.n2761 585
R2794 gnd.n3482 gnd.n2762 585
R2795 gnd.n3468 gnd.n2785 585
R2796 gnd.n2785 gnd.n2775 585
R2797 gnd.n3470 gnd.n3469 585
R2798 gnd.n3471 gnd.n3470 585
R2799 gnd.n2786 gnd.n2784 585
R2800 gnd.n3459 gnd.n2784 585
R2801 gnd.n3463 gnd.n3462 585
R2802 gnd.n3462 gnd.n3461 585
R2803 gnd.n2789 gnd.n2788 585
R2804 gnd.n3414 gnd.n2789 585
R2805 gnd.n2907 gnd.n2906 585
R2806 gnd.n2908 gnd.n2907 585
R2807 gnd.n2887 gnd.n2886 585
R2808 gnd.n2890 gnd.n2887 585
R2809 gnd.n3424 gnd.n3423 585
R2810 gnd.n3423 gnd.n3422 585
R2811 gnd.n3425 gnd.n2881 585
R2812 gnd.n2917 gnd.n2881 585
R2813 gnd.n3427 gnd.n3426 585
R2814 gnd.n3428 gnd.n3427 585
R2815 gnd.n2882 gnd.n2880 585
R2816 gnd.n3392 gnd.n2880 585
R2817 gnd.n3376 gnd.n3375 585
R2818 gnd.n3375 gnd.n2868 585
R2819 gnd.n3377 gnd.n2932 585
R2820 gnd.n2932 gnd.n2867 585
R2821 gnd.n3379 gnd.n3378 585
R2822 gnd.n3380 gnd.n3379 585
R2823 gnd.n2933 gnd.n2931 585
R2824 gnd.n2931 gnd.n2928 585
R2825 gnd.n3368 gnd.n3367 585
R2826 gnd.n3367 gnd.n3366 585
R2827 gnd.n2936 gnd.n2935 585
R2828 gnd.n2943 gnd.n2936 585
R2829 gnd.n3342 gnd.n3341 585
R2830 gnd.n3343 gnd.n3342 585
R2831 gnd.n2955 gnd.n2954 585
R2832 gnd.n2962 gnd.n2954 585
R2833 gnd.n3337 gnd.n3336 585
R2834 gnd.n3336 gnd.n3335 585
R2835 gnd.n2958 gnd.n2957 585
R2836 gnd.n3325 gnd.n2958 585
R2837 gnd.n3312 gnd.n2982 585
R2838 gnd.n2982 gnd.n2981 585
R2839 gnd.n3314 gnd.n3313 585
R2840 gnd.n3315 gnd.n3314 585
R2841 gnd.n2983 gnd.n2980 585
R2842 gnd.n2990 gnd.n2980 585
R2843 gnd.n3307 gnd.n3306 585
R2844 gnd.n3306 gnd.n3305 585
R2845 gnd.n2986 gnd.n2985 585
R2846 gnd.n3294 gnd.n2986 585
R2847 gnd.n3281 gnd.n3007 585
R2848 gnd.n3007 gnd.n3006 585
R2849 gnd.n3283 gnd.n3282 585
R2850 gnd.n3284 gnd.n3283 585
R2851 gnd.n3277 gnd.n3005 585
R2852 gnd.n3276 gnd.n3275 585
R2853 gnd.n3010 gnd.n3009 585
R2854 gnd.n3273 gnd.n3010 585
R2855 gnd.n3032 gnd.n3031 585
R2856 gnd.n3035 gnd.n3034 585
R2857 gnd.n3033 gnd.n3028 585
R2858 gnd.n3040 gnd.n3039 585
R2859 gnd.n3042 gnd.n3041 585
R2860 gnd.n3045 gnd.n3044 585
R2861 gnd.n3043 gnd.n3026 585
R2862 gnd.n3050 gnd.n3049 585
R2863 gnd.n3052 gnd.n3051 585
R2864 gnd.n3055 gnd.n3054 585
R2865 gnd.n3053 gnd.n3024 585
R2866 gnd.n3060 gnd.n3059 585
R2867 gnd.n3064 gnd.n3061 585
R2868 gnd.n3065 gnd.n3002 585
R2869 gnd.n3944 gnd.n2603 585
R2870 gnd.n4011 gnd.n4010 585
R2871 gnd.n4013 gnd.n4012 585
R2872 gnd.n4015 gnd.n4014 585
R2873 gnd.n4017 gnd.n4016 585
R2874 gnd.n4019 gnd.n4018 585
R2875 gnd.n4021 gnd.n4020 585
R2876 gnd.n4023 gnd.n4022 585
R2877 gnd.n4025 gnd.n4024 585
R2878 gnd.n4027 gnd.n4026 585
R2879 gnd.n4029 gnd.n4028 585
R2880 gnd.n4031 gnd.n4030 585
R2881 gnd.n4033 gnd.n4032 585
R2882 gnd.n4036 gnd.n4035 585
R2883 gnd.n4034 gnd.n2591 585
R2884 gnd.n4040 gnd.n2589 585
R2885 gnd.n4042 gnd.n4041 585
R2886 gnd.n4043 gnd.n4042 585
R2887 gnd.n3945 gnd.n2644 585
R2888 gnd.n3945 gnd.n2565 585
R2889 gnd.n3947 gnd.n3946 585
R2890 gnd.n3946 gnd.n2639 585
R2891 gnd.n3943 gnd.n2643 585
R2892 gnd.n3943 gnd.n3942 585
R2893 gnd.n3922 gnd.n2645 585
R2894 gnd.n2657 gnd.n2645 585
R2895 gnd.n3921 gnd.n2655 585
R2896 gnd.n3930 gnd.n2655 585
R2897 gnd.n3655 gnd.n2662 585
R2898 gnd.n3657 gnd.n3655 585
R2899 gnd.n3654 gnd.n3653 585
R2900 gnd.n3654 gnd.n2666 585
R2901 gnd.n3652 gnd.n2668 585
R2902 gnd.n3645 gnd.n2668 585
R2903 gnd.n2681 gnd.n2669 585
R2904 gnd.n2681 gnd.n2673 585
R2905 gnd.n3601 gnd.n2682 585
R2906 gnd.n3635 gnd.n2682 585
R2907 gnd.n3600 gnd.n3599 585
R2908 gnd.n3599 gnd.n2689 585
R2909 gnd.n3598 gnd.n2697 585
R2910 gnd.n3598 gnd.n2688 585
R2911 gnd.n3597 gnd.n2699 585
R2912 gnd.n3597 gnd.n3596 585
R2913 gnd.n3576 gnd.n2698 585
R2914 gnd.n2711 gnd.n2698 585
R2915 gnd.n3575 gnd.n2709 585
R2916 gnd.n3586 gnd.n2709 585
R2917 gnd.n3566 gnd.n2716 585
R2918 gnd.n3567 gnd.n3566 585
R2919 gnd.n3565 gnd.n3564 585
R2920 gnd.n3565 gnd.n2720 585
R2921 gnd.n3563 gnd.n2722 585
R2922 gnd.n3556 gnd.n2722 585
R2923 gnd.n2737 gnd.n2723 585
R2924 gnd.n2737 gnd.n2727 585
R2925 gnd.n3516 gnd.n2738 585
R2926 gnd.n3546 gnd.n2738 585
R2927 gnd.n3515 gnd.n3514 585
R2928 gnd.n3514 gnd.n2745 585
R2929 gnd.n3513 gnd.n2752 585
R2930 gnd.n3513 gnd.n2744 585
R2931 gnd.n3512 gnd.n2754 585
R2932 gnd.n3512 gnd.n3511 585
R2933 gnd.n3491 gnd.n2753 585
R2934 gnd.n2766 gnd.n2753 585
R2935 gnd.n3490 gnd.n2764 585
R2936 gnd.n3501 gnd.n2764 585
R2937 gnd.n3481 gnd.n2771 585
R2938 gnd.n3482 gnd.n3481 585
R2939 gnd.n3480 gnd.n3479 585
R2940 gnd.n3480 gnd.n2775 585
R2941 gnd.n3478 gnd.n2777 585
R2942 gnd.n3471 gnd.n2777 585
R2943 gnd.n3458 gnd.n2778 585
R2944 gnd.n3459 gnd.n3458 585
R2945 gnd.n3411 gnd.n2791 585
R2946 gnd.n3461 gnd.n2791 585
R2947 gnd.n3413 gnd.n3412 585
R2948 gnd.n3414 gnd.n3413 585
R2949 gnd.n3406 gnd.n2909 585
R2950 gnd.n2909 gnd.n2908 585
R2951 gnd.n3404 gnd.n3403 585
R2952 gnd.n3403 gnd.n2890 585
R2953 gnd.n3401 gnd.n2888 585
R2954 gnd.n3422 gnd.n2888 585
R2955 gnd.n2919 gnd.n2918 585
R2956 gnd.n2918 gnd.n2917 585
R2957 gnd.n3395 gnd.n2878 585
R2958 gnd.n3428 gnd.n2878 585
R2959 gnd.n3394 gnd.n3393 585
R2960 gnd.n3393 gnd.n3392 585
R2961 gnd.n3390 gnd.n2921 585
R2962 gnd.n3390 gnd.n2868 585
R2963 gnd.n3389 gnd.n3388 585
R2964 gnd.n3389 gnd.n2867 585
R2965 gnd.n2924 gnd.n2923 585
R2966 gnd.n3380 gnd.n2923 585
R2967 gnd.n3348 gnd.n3347 585
R2968 gnd.n3347 gnd.n2928 585
R2969 gnd.n3349 gnd.n2937 585
R2970 gnd.n3366 gnd.n2937 585
R2971 gnd.n3346 gnd.n3345 585
R2972 gnd.n3345 gnd.n2943 585
R2973 gnd.n3344 gnd.n2951 585
R2974 gnd.n3344 gnd.n3343 585
R2975 gnd.n3329 gnd.n2952 585
R2976 gnd.n2962 gnd.n2952 585
R2977 gnd.n3328 gnd.n2960 585
R2978 gnd.n3335 gnd.n2960 585
R2979 gnd.n3327 gnd.n3326 585
R2980 gnd.n3326 gnd.n3325 585
R2981 gnd.n2971 gnd.n2968 585
R2982 gnd.n2981 gnd.n2971 585
R2983 gnd.n3317 gnd.n3316 585
R2984 gnd.n3316 gnd.n3315 585
R2985 gnd.n2977 gnd.n2976 585
R2986 gnd.n2990 gnd.n2977 585
R2987 gnd.n3297 gnd.n2988 585
R2988 gnd.n3305 gnd.n2988 585
R2989 gnd.n3296 gnd.n3295 585
R2990 gnd.n3295 gnd.n3294 585
R2991 gnd.n2997 gnd.n2995 585
R2992 gnd.n3006 gnd.n2997 585
R2993 gnd.n3286 gnd.n3285 585
R2994 gnd.n3285 gnd.n3284 585
R2995 gnd.n5544 gnd.n1772 585
R2996 gnd.n1772 gnd.n1728 585
R2997 gnd.n5546 gnd.n5545 585
R2998 gnd.n5547 gnd.n5546 585
R2999 gnd.n5455 gnd.n1771 585
R3000 gnd.n1776 gnd.n1771 585
R3001 gnd.n5454 gnd.n5453 585
R3002 gnd.n5453 gnd.n5452 585
R3003 gnd.n1774 gnd.n1773 585
R3004 gnd.n5428 gnd.n1774 585
R3005 gnd.n5440 gnd.n5439 585
R3006 gnd.n5441 gnd.n5440 585
R3007 gnd.n5438 gnd.n1787 585
R3008 gnd.n1787 gnd.n1784 585
R3009 gnd.n5437 gnd.n5436 585
R3010 gnd.n5436 gnd.n5435 585
R3011 gnd.n1789 gnd.n1788 585
R3012 gnd.n1802 gnd.n1789 585
R3013 gnd.n5394 gnd.n5393 585
R3014 gnd.n5393 gnd.n1801 585
R3015 gnd.n5395 gnd.n1814 585
R3016 gnd.n5382 gnd.n1814 585
R3017 gnd.n5397 gnd.n5396 585
R3018 gnd.n5398 gnd.n5397 585
R3019 gnd.n5392 gnd.n1813 585
R3020 gnd.n1813 gnd.n1808 585
R3021 gnd.n5391 gnd.n5390 585
R3022 gnd.n5390 gnd.n5389 585
R3023 gnd.n1816 gnd.n1815 585
R3024 gnd.n1822 gnd.n1816 585
R3025 gnd.n5375 gnd.n5374 585
R3026 gnd.n5376 gnd.n5375 585
R3027 gnd.n5373 gnd.n1824 585
R3028 gnd.n1830 gnd.n1824 585
R3029 gnd.n5372 gnd.n5371 585
R3030 gnd.n5371 gnd.n5370 585
R3031 gnd.n1826 gnd.n1825 585
R3032 gnd.n1841 gnd.n1826 585
R3033 gnd.n5358 gnd.n5357 585
R3034 gnd.t23 gnd.n5358 585
R3035 gnd.n5356 gnd.n1842 585
R3036 gnd.n1842 gnd.n1838 585
R3037 gnd.n5355 gnd.n5354 585
R3038 gnd.n5354 gnd.n5353 585
R3039 gnd.n1844 gnd.n1843 585
R3040 gnd.n1845 gnd.n1844 585
R3041 gnd.n5311 gnd.n1867 585
R3042 gnd.n5311 gnd.n5310 585
R3043 gnd.n5313 gnd.n5312 585
R3044 gnd.n5312 gnd.n1853 585
R3045 gnd.n5314 gnd.n1865 585
R3046 gnd.n5294 gnd.n1865 585
R3047 gnd.n5316 gnd.n5315 585
R3048 gnd.n5317 gnd.n5316 585
R3049 gnd.n1866 gnd.n1864 585
R3050 gnd.n1864 gnd.n1860 585
R3051 gnd.n1895 gnd.n1873 585
R3052 gnd.n5289 gnd.n1873 585
R3053 gnd.n1897 gnd.n1896 585
R3054 gnd.n1897 gnd.n1872 585
R3055 gnd.n5261 gnd.n1894 585
R3056 gnd.n5261 gnd.n5260 585
R3057 gnd.n5263 gnd.n5262 585
R3058 gnd.n5262 gnd.n1880 585
R3059 gnd.n5264 gnd.n1892 585
R3060 gnd.n5252 gnd.n1892 585
R3061 gnd.n5266 gnd.n5265 585
R3062 gnd.n5267 gnd.n5266 585
R3063 gnd.n1893 gnd.n1891 585
R3064 gnd.n1891 gnd.n1887 585
R3065 gnd.n5246 gnd.n5245 585
R3066 gnd.n5247 gnd.n5246 585
R3067 gnd.n5244 gnd.n1902 585
R3068 gnd.n1907 gnd.n1902 585
R3069 gnd.n5243 gnd.n5242 585
R3070 gnd.n5242 gnd.n5241 585
R3071 gnd.n1904 gnd.n1903 585
R3072 gnd.n5217 gnd.n1904 585
R3073 gnd.n5229 gnd.n5228 585
R3074 gnd.n5230 gnd.n5229 585
R3075 gnd.n5227 gnd.n1917 585
R3076 gnd.n1917 gnd.n1913 585
R3077 gnd.n5226 gnd.n5225 585
R3078 gnd.n5225 gnd.n5224 585
R3079 gnd.n1919 gnd.n1918 585
R3080 gnd.n1925 gnd.n1919 585
R3081 gnd.n5210 gnd.n5209 585
R3082 gnd.n5211 gnd.n5210 585
R3083 gnd.n5208 gnd.n1927 585
R3084 gnd.n1934 gnd.n1927 585
R3085 gnd.n5207 gnd.n5206 585
R3086 gnd.n5206 gnd.n5205 585
R3087 gnd.n1929 gnd.n1928 585
R3088 gnd.n1943 gnd.n1929 585
R3089 gnd.n5192 gnd.n5191 585
R3090 gnd.n5193 gnd.n5192 585
R3091 gnd.n5190 gnd.n1944 585
R3092 gnd.n5185 gnd.n1944 585
R3093 gnd.n5189 gnd.n5188 585
R3094 gnd.n5188 gnd.n5187 585
R3095 gnd.n1946 gnd.n1945 585
R3096 gnd.n1947 gnd.n1946 585
R3097 gnd.n5173 gnd.n5172 585
R3098 gnd.n5174 gnd.n5173 585
R3099 gnd.n5171 gnd.n1952 585
R3100 gnd.n1957 gnd.n1952 585
R3101 gnd.n5170 gnd.n5169 585
R3102 gnd.n5169 gnd.n5168 585
R3103 gnd.n1954 gnd.n1953 585
R3104 gnd.n1955 gnd.n1954 585
R3105 gnd.n5125 gnd.n5124 585
R3106 gnd.n5126 gnd.n5125 585
R3107 gnd.n5123 gnd.n1975 585
R3108 gnd.n5119 gnd.n1975 585
R3109 gnd.n5122 gnd.n5121 585
R3110 gnd.n5121 gnd.n5120 585
R3111 gnd.n1977 gnd.n1976 585
R3112 gnd.n5108 gnd.n1977 585
R3113 gnd.n5088 gnd.n5087 585
R3114 gnd.n5087 gnd.n1983 585
R3115 gnd.n5089 gnd.n1995 585
R3116 gnd.n5076 gnd.n1995 585
R3117 gnd.n5091 gnd.n5090 585
R3118 gnd.n5092 gnd.n5091 585
R3119 gnd.n5086 gnd.n1994 585
R3120 gnd.n1994 gnd.t58 585
R3121 gnd.n5085 gnd.n5084 585
R3122 gnd.n5084 gnd.n5083 585
R3123 gnd.n1997 gnd.n1996 585
R3124 gnd.n2004 gnd.n1997 585
R3125 gnd.n5071 gnd.n5070 585
R3126 gnd.n5072 gnd.n5071 585
R3127 gnd.n5069 gnd.n2006 585
R3128 gnd.n2012 gnd.n2006 585
R3129 gnd.n5068 gnd.n5067 585
R3130 gnd.n5067 gnd.n5066 585
R3131 gnd.n2008 gnd.n2007 585
R3132 gnd.n2021 gnd.n2008 585
R3133 gnd.n5052 gnd.n5051 585
R3134 gnd.n5053 gnd.n5052 585
R3135 gnd.n5050 gnd.n2022 585
R3136 gnd.n5045 gnd.n2022 585
R3137 gnd.n5049 gnd.n5048 585
R3138 gnd.n5048 gnd.n5047 585
R3139 gnd.n2024 gnd.n2023 585
R3140 gnd.n5035 gnd.n2024 585
R3141 gnd.n4978 gnd.n4977 585
R3142 gnd.n4978 gnd.n2029 585
R3143 gnd.n4980 gnd.n4979 585
R3144 gnd.n4979 gnd.n2031 585
R3145 gnd.n4981 gnd.n4974 585
R3146 gnd.n4974 gnd.n4973 585
R3147 gnd.n4983 gnd.n4982 585
R3148 gnd.n4984 gnd.n4983 585
R3149 gnd.n4976 gnd.n4972 585
R3150 gnd.n4972 gnd.n4971 585
R3151 gnd.n4975 gnd.n4893 585
R3152 gnd.n4990 gnd.n4893 585
R3153 gnd.n1182 gnd.n1181 585
R3154 gnd.n4892 gnd.n1182 585
R3155 gnd.n6275 gnd.n6274 585
R3156 gnd.n6274 gnd.n6273 585
R3157 gnd.n6276 gnd.n1160 585
R3158 gnd.n4961 gnd.n1160 585
R3159 gnd.n6341 gnd.n6340 585
R3160 gnd.n6339 gnd.n1159 585
R3161 gnd.n6338 gnd.n1158 585
R3162 gnd.n6343 gnd.n1158 585
R3163 gnd.n6337 gnd.n6336 585
R3164 gnd.n6335 gnd.n6334 585
R3165 gnd.n6333 gnd.n6332 585
R3166 gnd.n6331 gnd.n6330 585
R3167 gnd.n6329 gnd.n6328 585
R3168 gnd.n6327 gnd.n6326 585
R3169 gnd.n6325 gnd.n6324 585
R3170 gnd.n6323 gnd.n6322 585
R3171 gnd.n6321 gnd.n6320 585
R3172 gnd.n6319 gnd.n6318 585
R3173 gnd.n6317 gnd.n6316 585
R3174 gnd.n6315 gnd.n6314 585
R3175 gnd.n6313 gnd.n6312 585
R3176 gnd.n6311 gnd.n6310 585
R3177 gnd.n6309 gnd.n6308 585
R3178 gnd.n6307 gnd.n6306 585
R3179 gnd.n6305 gnd.n6304 585
R3180 gnd.n6303 gnd.n6302 585
R3181 gnd.n6301 gnd.n6300 585
R3182 gnd.n6299 gnd.n6298 585
R3183 gnd.n6297 gnd.n6296 585
R3184 gnd.n6295 gnd.n6294 585
R3185 gnd.n6293 gnd.n6292 585
R3186 gnd.n6291 gnd.n6290 585
R3187 gnd.n6289 gnd.n6288 585
R3188 gnd.n6287 gnd.n6286 585
R3189 gnd.n6285 gnd.n6284 585
R3190 gnd.n6283 gnd.n6282 585
R3191 gnd.n6281 gnd.n1122 585
R3192 gnd.n6346 gnd.n6345 585
R3193 gnd.n1124 gnd.n1121 585
R3194 gnd.n4899 gnd.n4898 585
R3195 gnd.n4901 gnd.n4900 585
R3196 gnd.n4904 gnd.n4903 585
R3197 gnd.n4906 gnd.n4905 585
R3198 gnd.n4908 gnd.n4907 585
R3199 gnd.n4910 gnd.n4909 585
R3200 gnd.n4912 gnd.n4911 585
R3201 gnd.n4914 gnd.n4913 585
R3202 gnd.n4916 gnd.n4915 585
R3203 gnd.n4918 gnd.n4917 585
R3204 gnd.n4920 gnd.n4919 585
R3205 gnd.n4922 gnd.n4921 585
R3206 gnd.n4924 gnd.n4923 585
R3207 gnd.n4926 gnd.n4925 585
R3208 gnd.n4928 gnd.n4927 585
R3209 gnd.n4930 gnd.n4929 585
R3210 gnd.n4932 gnd.n4931 585
R3211 gnd.n4934 gnd.n4933 585
R3212 gnd.n4936 gnd.n4935 585
R3213 gnd.n4938 gnd.n4937 585
R3214 gnd.n4940 gnd.n4939 585
R3215 gnd.n4942 gnd.n4941 585
R3216 gnd.n4944 gnd.n4943 585
R3217 gnd.n4946 gnd.n4945 585
R3218 gnd.n4948 gnd.n4947 585
R3219 gnd.n4950 gnd.n4949 585
R3220 gnd.n4952 gnd.n4951 585
R3221 gnd.n4954 gnd.n4953 585
R3222 gnd.n4956 gnd.n4955 585
R3223 gnd.n4958 gnd.n4957 585
R3224 gnd.n4960 gnd.n4959 585
R3225 gnd.n5551 gnd.n5550 585
R3226 gnd.n5553 gnd.n5552 585
R3227 gnd.n5555 gnd.n5554 585
R3228 gnd.n5557 gnd.n5556 585
R3229 gnd.n5559 gnd.n5558 585
R3230 gnd.n5561 gnd.n5560 585
R3231 gnd.n5563 gnd.n5562 585
R3232 gnd.n5565 gnd.n5564 585
R3233 gnd.n5567 gnd.n5566 585
R3234 gnd.n5569 gnd.n5568 585
R3235 gnd.n5571 gnd.n5570 585
R3236 gnd.n5573 gnd.n5572 585
R3237 gnd.n5575 gnd.n5574 585
R3238 gnd.n5577 gnd.n5576 585
R3239 gnd.n5579 gnd.n5578 585
R3240 gnd.n5581 gnd.n5580 585
R3241 gnd.n5583 gnd.n5582 585
R3242 gnd.n5585 gnd.n5584 585
R3243 gnd.n5587 gnd.n5586 585
R3244 gnd.n5589 gnd.n5588 585
R3245 gnd.n5591 gnd.n5590 585
R3246 gnd.n5593 gnd.n5592 585
R3247 gnd.n5595 gnd.n5594 585
R3248 gnd.n5597 gnd.n5596 585
R3249 gnd.n5599 gnd.n5598 585
R3250 gnd.n5601 gnd.n5600 585
R3251 gnd.n5603 gnd.n5602 585
R3252 gnd.n5605 gnd.n5604 585
R3253 gnd.n5607 gnd.n5606 585
R3254 gnd.n5610 gnd.n5609 585
R3255 gnd.n5612 gnd.n5611 585
R3256 gnd.n5614 gnd.n5613 585
R3257 gnd.n5616 gnd.n5615 585
R3258 gnd.n5477 gnd.n1437 585
R3259 gnd.n5479 gnd.n5478 585
R3260 gnd.n5481 gnd.n5480 585
R3261 gnd.n5483 gnd.n5482 585
R3262 gnd.n5486 gnd.n5485 585
R3263 gnd.n5488 gnd.n5487 585
R3264 gnd.n5490 gnd.n5489 585
R3265 gnd.n5492 gnd.n5491 585
R3266 gnd.n5494 gnd.n5493 585
R3267 gnd.n5496 gnd.n5495 585
R3268 gnd.n5498 gnd.n5497 585
R3269 gnd.n5500 gnd.n5499 585
R3270 gnd.n5502 gnd.n5501 585
R3271 gnd.n5504 gnd.n5503 585
R3272 gnd.n5506 gnd.n5505 585
R3273 gnd.n5508 gnd.n5507 585
R3274 gnd.n5510 gnd.n5509 585
R3275 gnd.n5512 gnd.n5511 585
R3276 gnd.n5514 gnd.n5513 585
R3277 gnd.n5516 gnd.n5515 585
R3278 gnd.n5518 gnd.n5517 585
R3279 gnd.n5520 gnd.n5519 585
R3280 gnd.n5522 gnd.n5521 585
R3281 gnd.n5524 gnd.n5523 585
R3282 gnd.n5526 gnd.n5525 585
R3283 gnd.n5528 gnd.n5527 585
R3284 gnd.n5530 gnd.n5529 585
R3285 gnd.n5532 gnd.n5531 585
R3286 gnd.n5534 gnd.n5533 585
R3287 gnd.n5536 gnd.n5535 585
R3288 gnd.n5538 gnd.n5537 585
R3289 gnd.n5540 gnd.n5539 585
R3290 gnd.n5542 gnd.n5541 585
R3291 gnd.n5549 gnd.n1767 585
R3292 gnd.n5549 gnd.n1728 585
R3293 gnd.n5548 gnd.n1769 585
R3294 gnd.n5548 gnd.n5547 585
R3295 gnd.n1794 gnd.n1768 585
R3296 gnd.n1776 gnd.n1768 585
R3297 gnd.n1795 gnd.n1777 585
R3298 gnd.n5452 gnd.n1777 585
R3299 gnd.n5430 gnd.n5429 585
R3300 gnd.n5429 gnd.n5428 585
R3301 gnd.n5431 gnd.n1786 585
R3302 gnd.n5441 gnd.n1786 585
R3303 gnd.n5432 gnd.n1792 585
R3304 gnd.n1792 gnd.n1784 585
R3305 gnd.n5434 gnd.n5433 585
R3306 gnd.n5435 gnd.n5434 585
R3307 gnd.n1793 gnd.n1791 585
R3308 gnd.n1802 gnd.n1791 585
R3309 gnd.n5381 gnd.n5380 585
R3310 gnd.n5381 gnd.n1801 585
R3311 gnd.n5384 gnd.n5383 585
R3312 gnd.n5383 gnd.n5382 585
R3313 gnd.n5385 gnd.n1810 585
R3314 gnd.n5398 gnd.n1810 585
R3315 gnd.n5386 gnd.n1819 585
R3316 gnd.n1819 gnd.n1808 585
R3317 gnd.n5388 gnd.n5387 585
R3318 gnd.n5389 gnd.n5388 585
R3319 gnd.n5379 gnd.n1818 585
R3320 gnd.n1822 gnd.n1818 585
R3321 gnd.n5378 gnd.n5377 585
R3322 gnd.n5377 gnd.n5376 585
R3323 gnd.n1821 gnd.n1820 585
R3324 gnd.n1830 gnd.n1821 585
R3325 gnd.n5298 gnd.n1828 585
R3326 gnd.n5370 gnd.n1828 585
R3327 gnd.n5300 gnd.n5299 585
R3328 gnd.n5299 gnd.n1841 585
R3329 gnd.n5301 gnd.n1840 585
R3330 gnd.t23 gnd.n1840 585
R3331 gnd.n5303 gnd.n5302 585
R3332 gnd.n5302 gnd.n1838 585
R3333 gnd.n5304 gnd.n1846 585
R3334 gnd.n5353 gnd.n1846 585
R3335 gnd.n5305 gnd.n1869 585
R3336 gnd.n1869 gnd.n1845 585
R3337 gnd.n5307 gnd.n5306 585
R3338 gnd.n5310 gnd.n5307 585
R3339 gnd.n5297 gnd.n1868 585
R3340 gnd.n1868 gnd.n1853 585
R3341 gnd.n5296 gnd.n5295 585
R3342 gnd.n5295 gnd.n5294 585
R3343 gnd.n5293 gnd.n1862 585
R3344 gnd.n5317 gnd.n1862 585
R3345 gnd.n5292 gnd.n5291 585
R3346 gnd.n5291 gnd.n1860 585
R3347 gnd.n5290 gnd.n1870 585
R3348 gnd.n5290 gnd.n5289 585
R3349 gnd.n5256 gnd.n1871 585
R3350 gnd.n1872 gnd.n1871 585
R3351 gnd.n5258 gnd.n5257 585
R3352 gnd.n5260 gnd.n5258 585
R3353 gnd.n5255 gnd.n1898 585
R3354 gnd.n1898 gnd.n1880 585
R3355 gnd.n5254 gnd.n5253 585
R3356 gnd.n5253 gnd.n5252 585
R3357 gnd.n5251 gnd.n1889 585
R3358 gnd.n5267 gnd.n1889 585
R3359 gnd.n5250 gnd.n5249 585
R3360 gnd.n5249 gnd.n1887 585
R3361 gnd.n5248 gnd.n1899 585
R3362 gnd.n5248 gnd.n5247 585
R3363 gnd.n5215 gnd.n1900 585
R3364 gnd.n1907 gnd.n1900 585
R3365 gnd.n5216 gnd.n1905 585
R3366 gnd.n5241 gnd.n1905 585
R3367 gnd.n5219 gnd.n5218 585
R3368 gnd.n5218 gnd.n5217 585
R3369 gnd.n5220 gnd.n1915 585
R3370 gnd.n5230 gnd.n1915 585
R3371 gnd.n5221 gnd.n1922 585
R3372 gnd.n1922 gnd.n1913 585
R3373 gnd.n5223 gnd.n5222 585
R3374 gnd.n5224 gnd.n5223 585
R3375 gnd.n5214 gnd.n1921 585
R3376 gnd.n1925 gnd.n1921 585
R3377 gnd.n5213 gnd.n5212 585
R3378 gnd.n5212 gnd.n5211 585
R3379 gnd.n1924 gnd.n1923 585
R3380 gnd.n1934 gnd.n1924 585
R3381 gnd.n5179 gnd.n1932 585
R3382 gnd.n5205 gnd.n1932 585
R3383 gnd.n5181 gnd.n5180 585
R3384 gnd.n5180 gnd.n1943 585
R3385 gnd.n5182 gnd.n1942 585
R3386 gnd.n5193 gnd.n1942 585
R3387 gnd.n5184 gnd.n5183 585
R3388 gnd.n5185 gnd.n5184 585
R3389 gnd.n5178 gnd.n1948 585
R3390 gnd.n5187 gnd.n1948 585
R3391 gnd.n5177 gnd.n5176 585
R3392 gnd.n5176 gnd.n1947 585
R3393 gnd.n5175 gnd.n1950 585
R3394 gnd.n5175 gnd.n5174 585
R3395 gnd.n5112 gnd.n1951 585
R3396 gnd.n1957 gnd.n1951 585
R3397 gnd.n5113 gnd.n1958 585
R3398 gnd.n5168 gnd.n1958 585
R3399 gnd.n5115 gnd.n5114 585
R3400 gnd.n5114 gnd.n1955 585
R3401 gnd.n5116 gnd.n1974 585
R3402 gnd.n5126 gnd.n1974 585
R3403 gnd.n5118 gnd.n5117 585
R3404 gnd.n5119 gnd.n5118 585
R3405 gnd.n5111 gnd.n1980 585
R3406 gnd.n5120 gnd.n1980 585
R3407 gnd.n5110 gnd.n5109 585
R3408 gnd.n5109 gnd.n5108 585
R3409 gnd.n1982 gnd.n1981 585
R3410 gnd.n1983 gnd.n1982 585
R3411 gnd.n5078 gnd.n5077 585
R3412 gnd.n5077 gnd.n5076 585
R3413 gnd.n5079 gnd.n1992 585
R3414 gnd.n5092 gnd.n1992 585
R3415 gnd.n5080 gnd.n2001 585
R3416 gnd.n2001 gnd.t58 585
R3417 gnd.n5082 gnd.n5081 585
R3418 gnd.n5083 gnd.n5082 585
R3419 gnd.n5075 gnd.n2000 585
R3420 gnd.n2004 gnd.n2000 585
R3421 gnd.n5074 gnd.n5073 585
R3422 gnd.n5073 gnd.n5072 585
R3423 gnd.n2003 gnd.n2002 585
R3424 gnd.n2012 gnd.n2003 585
R3425 gnd.n5039 gnd.n2010 585
R3426 gnd.n5066 gnd.n2010 585
R3427 gnd.n5041 gnd.n5040 585
R3428 gnd.n5040 gnd.n2021 585
R3429 gnd.n5042 gnd.n2020 585
R3430 gnd.n5053 gnd.n2020 585
R3431 gnd.n5044 gnd.n5043 585
R3432 gnd.n5045 gnd.n5044 585
R3433 gnd.n5038 gnd.n2025 585
R3434 gnd.n5047 gnd.n2025 585
R3435 gnd.n5037 gnd.n5036 585
R3436 gnd.n5036 gnd.n5035 585
R3437 gnd.n2028 gnd.n2027 585
R3438 gnd.n2029 gnd.n2028 585
R3439 gnd.n4968 gnd.n4967 585
R3440 gnd.n4968 gnd.n2031 585
R3441 gnd.n4969 gnd.n4966 585
R3442 gnd.n4973 gnd.n4969 585
R3443 gnd.n4986 gnd.n4985 585
R3444 gnd.n4985 gnd.n4984 585
R3445 gnd.n4987 gnd.n4895 585
R3446 gnd.n4971 gnd.n4895 585
R3447 gnd.n4989 gnd.n4988 585
R3448 gnd.n4990 gnd.n4989 585
R3449 gnd.n4965 gnd.n4894 585
R3450 gnd.n4894 gnd.n4892 585
R3451 gnd.n4964 gnd.n1184 585
R3452 gnd.n6273 gnd.n1184 585
R3453 gnd.n4963 gnd.n4962 585
R3454 gnd.n4962 gnd.n4961 585
R3455 gnd.n6397 gnd.n6396 585
R3456 gnd.n6398 gnd.n6397 585
R3457 gnd.n1056 gnd.n1055 585
R3458 gnd.n4694 gnd.n1056 585
R3459 gnd.n6406 gnd.n6405 585
R3460 gnd.n6405 gnd.n6404 585
R3461 gnd.n6407 gnd.n1050 585
R3462 gnd.n4687 gnd.n1050 585
R3463 gnd.n6409 gnd.n6408 585
R3464 gnd.n6410 gnd.n6409 585
R3465 gnd.n1036 gnd.n1035 585
R3466 gnd.n4678 gnd.n1036 585
R3467 gnd.n6418 gnd.n6417 585
R3468 gnd.n6417 gnd.n6416 585
R3469 gnd.n6419 gnd.n1030 585
R3470 gnd.n4672 gnd.n1030 585
R3471 gnd.n6421 gnd.n6420 585
R3472 gnd.n6422 gnd.n6421 585
R3473 gnd.n1015 gnd.n1014 585
R3474 gnd.n4607 gnd.n1015 585
R3475 gnd.n6430 gnd.n6429 585
R3476 gnd.n6429 gnd.n6428 585
R3477 gnd.n6431 gnd.n1009 585
R3478 gnd.n4601 gnd.n1009 585
R3479 gnd.n6433 gnd.n6432 585
R3480 gnd.n6434 gnd.n6433 585
R3481 gnd.n996 gnd.n995 585
R3482 gnd.n4595 gnd.n996 585
R3483 gnd.n6442 gnd.n6441 585
R3484 gnd.n6441 gnd.n6440 585
R3485 gnd.n6443 gnd.n990 585
R3486 gnd.n4624 gnd.n990 585
R3487 gnd.n6445 gnd.n6444 585
R3488 gnd.n6446 gnd.n6445 585
R3489 gnd.n975 gnd.n974 585
R3490 gnd.n4588 gnd.n975 585
R3491 gnd.n6454 gnd.n6453 585
R3492 gnd.n6453 gnd.n6452 585
R3493 gnd.n6455 gnd.n970 585
R3494 gnd.n4580 gnd.n970 585
R3495 gnd.n6457 gnd.n6456 585
R3496 gnd.n6458 gnd.n6457 585
R3497 gnd.n955 gnd.n953 585
R3498 gnd.n4573 gnd.n955 585
R3499 gnd.n6466 gnd.n6465 585
R3500 gnd.n6465 gnd.n6464 585
R3501 gnd.n954 gnd.n952 585
R3502 gnd.n4565 gnd.n954 585
R3503 gnd.n4534 gnd.n4533 585
R3504 gnd.n4535 gnd.n4534 585
R3505 gnd.n4532 gnd.n4531 585
R3506 gnd.n4531 gnd.n2432 585
R3507 gnd.n4530 gnd.n2435 585
R3508 gnd.n4530 gnd.n4529 585
R3509 gnd.n945 gnd.n943 585
R3510 gnd.n4516 gnd.n943 585
R3511 gnd.n6470 gnd.n6469 585
R3512 gnd.n6471 gnd.n6470 585
R3513 gnd.n944 gnd.n942 585
R3514 gnd.n942 gnd.n938 585
R3515 gnd.n4500 gnd.n4499 585
R3516 gnd.n4501 gnd.n4500 585
R3517 gnd.n4498 gnd.n2455 585
R3518 gnd.n4498 gnd.n4497 585
R3519 gnd.n4478 gnd.n2454 585
R3520 gnd.n2456 gnd.n2454 585
R3521 gnd.n4480 gnd.n4479 585
R3522 gnd.n4481 gnd.n4480 585
R3523 gnd.n2468 gnd.n2467 585
R3524 gnd.n2474 gnd.n2467 585
R3525 gnd.n4474 gnd.n4473 585
R3526 gnd.n4473 gnd.n4472 585
R3527 gnd.n2471 gnd.n2470 585
R3528 gnd.n4461 gnd.n2471 585
R3529 gnd.n4438 gnd.n2491 585
R3530 gnd.n2491 gnd.n2482 585
R3531 gnd.n4440 gnd.n4439 585
R3532 gnd.n4441 gnd.n4440 585
R3533 gnd.n2492 gnd.n2490 585
R3534 gnd.n2499 gnd.n2490 585
R3535 gnd.n4433 gnd.n4432 585
R3536 gnd.n4432 gnd.n4431 585
R3537 gnd.n2495 gnd.n2494 585
R3538 gnd.n2496 gnd.n2495 585
R3539 gnd.n4414 gnd.n4413 585
R3540 gnd.n4415 gnd.n4414 585
R3541 gnd.n2512 gnd.n2511 585
R3542 gnd.n2511 gnd.n2508 585
R3543 gnd.n4409 gnd.n4408 585
R3544 gnd.n4408 gnd.n4407 585
R3545 gnd.n2515 gnd.n2514 585
R3546 gnd.n2516 gnd.n2515 585
R3547 gnd.n4394 gnd.n4393 585
R3548 gnd.n4395 gnd.n4394 585
R3549 gnd.n2529 gnd.n2528 585
R3550 gnd.n2536 gnd.n2528 585
R3551 gnd.n4389 gnd.n4388 585
R3552 gnd.n4388 gnd.n4387 585
R3553 gnd.n2532 gnd.n2531 585
R3554 gnd.n2533 gnd.n2532 585
R3555 gnd.n4374 gnd.n4373 585
R3556 gnd.n4375 gnd.n4374 585
R3557 gnd.n2548 gnd.n2547 585
R3558 gnd.n2547 gnd.n2544 585
R3559 gnd.n4369 gnd.n4368 585
R3560 gnd.n4368 gnd.n4367 585
R3561 gnd.n2551 gnd.n2550 585
R3562 gnd.n2552 gnd.n2551 585
R3563 gnd.n4355 gnd.n4354 585
R3564 gnd.n4353 gnd.n4082 585
R3565 gnd.n4352 gnd.n4081 585
R3566 gnd.n4357 gnd.n4081 585
R3567 gnd.n4351 gnd.n4350 585
R3568 gnd.n4349 gnd.n4348 585
R3569 gnd.n4347 gnd.n4346 585
R3570 gnd.n4345 gnd.n4344 585
R3571 gnd.n4343 gnd.n4342 585
R3572 gnd.n4341 gnd.n4340 585
R3573 gnd.n4339 gnd.n4338 585
R3574 gnd.n4337 gnd.n4336 585
R3575 gnd.n4335 gnd.n4334 585
R3576 gnd.n4333 gnd.n4332 585
R3577 gnd.n4331 gnd.n4330 585
R3578 gnd.n4329 gnd.n4328 585
R3579 gnd.n4327 gnd.n4326 585
R3580 gnd.n4325 gnd.n4324 585
R3581 gnd.n4323 gnd.n4322 585
R3582 gnd.n4320 gnd.n4319 585
R3583 gnd.n4318 gnd.n4317 585
R3584 gnd.n4316 gnd.n4315 585
R3585 gnd.n4314 gnd.n4313 585
R3586 gnd.n4312 gnd.n4311 585
R3587 gnd.n4310 gnd.n4309 585
R3588 gnd.n4308 gnd.n4307 585
R3589 gnd.n4306 gnd.n4305 585
R3590 gnd.n4304 gnd.n4303 585
R3591 gnd.n4302 gnd.n4301 585
R3592 gnd.n4300 gnd.n4299 585
R3593 gnd.n4298 gnd.n4297 585
R3594 gnd.n4296 gnd.n4295 585
R3595 gnd.n4294 gnd.n4293 585
R3596 gnd.n4292 gnd.n4291 585
R3597 gnd.n4290 gnd.n4289 585
R3598 gnd.n4288 gnd.n4287 585
R3599 gnd.n4286 gnd.n4285 585
R3600 gnd.n4284 gnd.n4283 585
R3601 gnd.n4282 gnd.n4281 585
R3602 gnd.n4280 gnd.n4279 585
R3603 gnd.n4278 gnd.n4277 585
R3604 gnd.n4276 gnd.n4275 585
R3605 gnd.n4274 gnd.n4273 585
R3606 gnd.n4272 gnd.n4271 585
R3607 gnd.n4270 gnd.n4269 585
R3608 gnd.n4268 gnd.n4267 585
R3609 gnd.n4266 gnd.n4265 585
R3610 gnd.n4264 gnd.n4263 585
R3611 gnd.n4262 gnd.n4261 585
R3612 gnd.n4260 gnd.n4259 585
R3613 gnd.n4258 gnd.n4257 585
R3614 gnd.n4256 gnd.n4255 585
R3615 gnd.n4254 gnd.n4253 585
R3616 gnd.n4252 gnd.n4251 585
R3617 gnd.n4250 gnd.n4249 585
R3618 gnd.n4248 gnd.n4247 585
R3619 gnd.n4246 gnd.n4245 585
R3620 gnd.n4244 gnd.n4243 585
R3621 gnd.n4242 gnd.n2564 585
R3622 gnd.n4359 gnd.n2563 585
R3623 gnd.n2303 gnd.n2302 585
R3624 gnd.n2300 gnd.n2196 585
R3625 gnd.n2299 gnd.n2298 585
R3626 gnd.n2292 gnd.n2198 585
R3627 gnd.n2294 gnd.n2293 585
R3628 gnd.n2290 gnd.n2200 585
R3629 gnd.n2289 gnd.n2288 585
R3630 gnd.n2282 gnd.n2202 585
R3631 gnd.n2284 gnd.n2283 585
R3632 gnd.n2280 gnd.n2204 585
R3633 gnd.n2279 gnd.n2278 585
R3634 gnd.n2272 gnd.n2206 585
R3635 gnd.n2274 gnd.n2273 585
R3636 gnd.n2270 gnd.n2208 585
R3637 gnd.n2269 gnd.n2268 585
R3638 gnd.n2262 gnd.n2210 585
R3639 gnd.n2264 gnd.n2263 585
R3640 gnd.n2260 gnd.n2212 585
R3641 gnd.n2259 gnd.n2258 585
R3642 gnd.n2252 gnd.n2214 585
R3643 gnd.n2254 gnd.n2253 585
R3644 gnd.n2250 gnd.n2218 585
R3645 gnd.n2249 gnd.n2248 585
R3646 gnd.n2242 gnd.n2220 585
R3647 gnd.n2244 gnd.n2243 585
R3648 gnd.n2240 gnd.n2222 585
R3649 gnd.n2239 gnd.n2238 585
R3650 gnd.n2232 gnd.n2224 585
R3651 gnd.n2234 gnd.n2233 585
R3652 gnd.n2230 gnd.n2227 585
R3653 gnd.n2229 gnd.n1117 585
R3654 gnd.n6348 gnd.n1113 585
R3655 gnd.n6350 gnd.n6349 585
R3656 gnd.n6352 gnd.n1111 585
R3657 gnd.n6354 gnd.n6353 585
R3658 gnd.n6355 gnd.n1106 585
R3659 gnd.n6357 gnd.n6356 585
R3660 gnd.n6359 gnd.n1104 585
R3661 gnd.n6361 gnd.n6360 585
R3662 gnd.n6363 gnd.n1097 585
R3663 gnd.n6365 gnd.n6364 585
R3664 gnd.n6367 gnd.n1095 585
R3665 gnd.n6369 gnd.n6368 585
R3666 gnd.n6370 gnd.n1090 585
R3667 gnd.n6372 gnd.n6371 585
R3668 gnd.n6374 gnd.n1088 585
R3669 gnd.n6376 gnd.n6375 585
R3670 gnd.n6377 gnd.n1083 585
R3671 gnd.n6379 gnd.n6378 585
R3672 gnd.n6381 gnd.n1081 585
R3673 gnd.n6383 gnd.n6382 585
R3674 gnd.n6384 gnd.n1075 585
R3675 gnd.n6386 gnd.n6385 585
R3676 gnd.n6388 gnd.n1074 585
R3677 gnd.n6389 gnd.n1072 585
R3678 gnd.n6392 gnd.n6391 585
R3679 gnd.n6393 gnd.n1069 585
R3680 gnd.n1073 gnd.n1069 585
R3681 gnd.n4691 gnd.n1066 585
R3682 gnd.n6398 gnd.n1066 585
R3683 gnd.n4693 gnd.n4692 585
R3684 gnd.n4694 gnd.n4693 585
R3685 gnd.n4690 gnd.n1058 585
R3686 gnd.n6404 gnd.n1058 585
R3687 gnd.n4689 gnd.n4688 585
R3688 gnd.n4688 gnd.n4687 585
R3689 gnd.n2384 gnd.n1047 585
R3690 gnd.n6410 gnd.n1047 585
R3691 gnd.n4677 gnd.n4676 585
R3692 gnd.n4678 gnd.n4677 585
R3693 gnd.n4675 gnd.n1037 585
R3694 gnd.n6416 gnd.n1037 585
R3695 gnd.n4674 gnd.n4673 585
R3696 gnd.n4673 gnd.n4672 585
R3697 gnd.n2389 gnd.n1027 585
R3698 gnd.n6422 gnd.n1027 585
R3699 gnd.n4606 gnd.n4605 585
R3700 gnd.n4607 gnd.n4606 585
R3701 gnd.n4604 gnd.n1017 585
R3702 gnd.n6428 gnd.n1017 585
R3703 gnd.n4603 gnd.n4602 585
R3704 gnd.n4602 gnd.n4601 585
R3705 gnd.n4598 gnd.n1007 585
R3706 gnd.n6434 gnd.n1007 585
R3707 gnd.n4597 gnd.n4596 585
R3708 gnd.n4596 gnd.n4595 585
R3709 gnd.n4594 gnd.n997 585
R3710 gnd.n6440 gnd.n997 585
R3711 gnd.n4593 gnd.n2403 585
R3712 gnd.n4624 gnd.n2403 585
R3713 gnd.n4591 gnd.n987 585
R3714 gnd.n6446 gnd.n987 585
R3715 gnd.n4590 gnd.n4589 585
R3716 gnd.n4589 gnd.n4588 585
R3717 gnd.n2412 gnd.n977 585
R3718 gnd.n6452 gnd.n977 585
R3719 gnd.n4579 gnd.n4578 585
R3720 gnd.n4580 gnd.n4579 585
R3721 gnd.n4576 gnd.n968 585
R3722 gnd.n6458 gnd.n968 585
R3723 gnd.n4575 gnd.n4574 585
R3724 gnd.n4574 gnd.n4573 585
R3725 gnd.n2417 gnd.n956 585
R3726 gnd.n6464 gnd.n956 585
R3727 gnd.n4522 gnd.n2423 585
R3728 gnd.n4565 gnd.n2423 585
R3729 gnd.n4523 gnd.n2433 585
R3730 gnd.n4535 gnd.n2433 585
R3731 gnd.n4521 gnd.n4520 585
R3732 gnd.n4520 gnd.n2432 585
R3733 gnd.n4519 gnd.n2437 585
R3734 gnd.n4529 gnd.n2437 585
R3735 gnd.n4518 gnd.n4517 585
R3736 gnd.n4517 gnd.n4516 585
R3737 gnd.n2446 gnd.n939 585
R3738 gnd.n6471 gnd.n939 585
R3739 gnd.n4488 gnd.n4487 585
R3740 gnd.n4487 gnd.n938 585
R3741 gnd.n4486 gnd.n2452 585
R3742 gnd.n4501 gnd.n2452 585
R3743 gnd.n4485 gnd.n2457 585
R3744 gnd.n4497 gnd.n2457 585
R3745 gnd.n4484 gnd.n4483 585
R3746 gnd.n4483 gnd.n2456 585
R3747 gnd.n4482 gnd.n2462 585
R3748 gnd.n4482 gnd.n4481 585
R3749 gnd.n4465 gnd.n2464 585
R3750 gnd.n2474 gnd.n2464 585
R3751 gnd.n4464 gnd.n2472 585
R3752 gnd.n4472 gnd.n2472 585
R3753 gnd.n4463 gnd.n4462 585
R3754 gnd.n4462 gnd.n4461 585
R3755 gnd.n2481 gnd.n2479 585
R3756 gnd.n2482 gnd.n2481 585
R3757 gnd.n4422 gnd.n2488 585
R3758 gnd.n4441 gnd.n2488 585
R3759 gnd.n4421 gnd.n4420 585
R3760 gnd.n4420 gnd.n2499 585
R3761 gnd.n4419 gnd.n2497 585
R3762 gnd.n4431 gnd.n2497 585
R3763 gnd.n4418 gnd.n4417 585
R3764 gnd.n4417 gnd.n2496 585
R3765 gnd.n4416 gnd.n2505 585
R3766 gnd.n4416 gnd.n4415 585
R3767 gnd.n4400 gnd.n2507 585
R3768 gnd.n2508 gnd.n2507 585
R3769 gnd.n4399 gnd.n2517 585
R3770 gnd.n4407 gnd.n2517 585
R3771 gnd.n4398 gnd.n4397 585
R3772 gnd.n4397 gnd.n2516 585
R3773 gnd.n4396 gnd.n2523 585
R3774 gnd.n4396 gnd.n4395 585
R3775 gnd.n4380 gnd.n2525 585
R3776 gnd.n2536 gnd.n2525 585
R3777 gnd.n4379 gnd.n2534 585
R3778 gnd.n4387 gnd.n2534 585
R3779 gnd.n4378 gnd.n4377 585
R3780 gnd.n4377 gnd.n2533 585
R3781 gnd.n4376 gnd.n2541 585
R3782 gnd.n4376 gnd.n4375 585
R3783 gnd.n4362 gnd.n2543 585
R3784 gnd.n2544 gnd.n2543 585
R3785 gnd.n4363 gnd.n2553 585
R3786 gnd.n4367 gnd.n2553 585
R3787 gnd.n4361 gnd.n4360 585
R3788 gnd.n4360 gnd.n2552 585
R3789 gnd.n7536 gnd.n7535 585
R3790 gnd.n7537 gnd.n7536 585
R3791 gnd.n201 gnd.n200 585
R3792 gnd.n209 gnd.n201 585
R3793 gnd.n7545 gnd.n7544 585
R3794 gnd.n7544 gnd.n7543 585
R3795 gnd.n7546 gnd.n195 585
R3796 gnd.n195 gnd.n194 585
R3797 gnd.n7548 gnd.n7547 585
R3798 gnd.n7549 gnd.n7548 585
R3799 gnd.n181 gnd.n180 585
R3800 gnd.n191 gnd.n181 585
R3801 gnd.n7557 gnd.n7556 585
R3802 gnd.n7556 gnd.n7555 585
R3803 gnd.n7558 gnd.n175 585
R3804 gnd.n175 gnd.n174 585
R3805 gnd.n7560 gnd.n7559 585
R3806 gnd.n7561 gnd.n7560 585
R3807 gnd.n161 gnd.n160 585
R3808 gnd.n171 gnd.n161 585
R3809 gnd.n7569 gnd.n7568 585
R3810 gnd.n7568 gnd.n7567 585
R3811 gnd.n7570 gnd.n155 585
R3812 gnd.n162 gnd.n155 585
R3813 gnd.n7572 gnd.n7571 585
R3814 gnd.n7573 gnd.n7572 585
R3815 gnd.n143 gnd.n142 585
R3816 gnd.n146 gnd.n143 585
R3817 gnd.n7581 gnd.n7580 585
R3818 gnd.n7580 gnd.n7579 585
R3819 gnd.n7582 gnd.n137 585
R3820 gnd.n137 gnd.n136 585
R3821 gnd.n7584 gnd.n7583 585
R3822 gnd.n7585 gnd.n7584 585
R3823 gnd.n123 gnd.n122 585
R3824 gnd.n133 gnd.n123 585
R3825 gnd.n7593 gnd.n7592 585
R3826 gnd.n7592 gnd.n7591 585
R3827 gnd.n7594 gnd.n118 585
R3828 gnd.n124 gnd.n118 585
R3829 gnd.n7596 gnd.n7595 585
R3830 gnd.n7597 gnd.n7596 585
R3831 gnd.n104 gnd.n102 585
R3832 gnd.n107 gnd.n104 585
R3833 gnd.n7605 gnd.n7604 585
R3834 gnd.n7604 gnd.n7603 585
R3835 gnd.n103 gnd.n95 585
R3836 gnd.n7345 gnd.n103 585
R3837 gnd.n7608 gnd.n93 585
R3838 gnd.n368 gnd.n93 585
R3839 gnd.n7610 gnd.n7609 585
R3840 gnd.n7611 gnd.n7610 585
R3841 gnd.n385 gnd.n92 585
R3842 gnd.n7296 gnd.n92 585
R3843 gnd.n7284 gnd.n386 585
R3844 gnd.n7284 gnd.n7283 585
R3845 gnd.n7286 gnd.n7285 585
R3846 gnd.n7287 gnd.n7286 585
R3847 gnd.n384 gnd.n100 585
R3848 gnd.n1597 gnd.n384 585
R3849 gnd.n5889 gnd.n1593 585
R3850 gnd.n5889 gnd.n5888 585
R3851 gnd.n5891 gnd.n5890 585
R3852 gnd.n5892 gnd.n5891 585
R3853 gnd.n1580 gnd.n1579 585
R3854 gnd.n5859 gnd.n1580 585
R3855 gnd.n5900 gnd.n5899 585
R3856 gnd.n5899 gnd.n5898 585
R3857 gnd.n5901 gnd.n1574 585
R3858 gnd.n5875 gnd.n1574 585
R3859 gnd.n5903 gnd.n5902 585
R3860 gnd.n5904 gnd.n5903 585
R3861 gnd.n1559 gnd.n1558 585
R3862 gnd.n5845 gnd.n1559 585
R3863 gnd.n5912 gnd.n5911 585
R3864 gnd.n5911 gnd.n5910 585
R3865 gnd.n5913 gnd.n1553 585
R3866 gnd.n5837 gnd.n1553 585
R3867 gnd.n5915 gnd.n5914 585
R3868 gnd.n5916 gnd.n5915 585
R3869 gnd.n1540 gnd.n1539 585
R3870 gnd.n5830 gnd.n1540 585
R3871 gnd.n5924 gnd.n5923 585
R3872 gnd.n5923 gnd.n5922 585
R3873 gnd.n5925 gnd.n1534 585
R3874 gnd.n5822 gnd.n1534 585
R3875 gnd.n5927 gnd.n5926 585
R3876 gnd.n5928 gnd.n5927 585
R3877 gnd.n1519 gnd.n1518 585
R3878 gnd.n5759 gnd.n1519 585
R3879 gnd.n5936 gnd.n5935 585
R3880 gnd.n5935 gnd.n5934 585
R3881 gnd.n5937 gnd.n1513 585
R3882 gnd.n5750 gnd.n1513 585
R3883 gnd.n5939 gnd.n5938 585
R3884 gnd.n5940 gnd.n5939 585
R3885 gnd.n1496 gnd.n1495 585
R3886 gnd.n5744 gnd.n1496 585
R3887 gnd.n5948 gnd.n5947 585
R3888 gnd.n5947 gnd.n5946 585
R3889 gnd.n5949 gnd.n1487 585
R3890 gnd.n5737 gnd.n1487 585
R3891 gnd.n5951 gnd.n5950 585
R3892 gnd.n5952 gnd.n5951 585
R3893 gnd.n1488 gnd.n1486 585
R3894 gnd.n5776 gnd.n1486 585
R3895 gnd.n1489 gnd.n1408 585
R3896 gnd.n5960 gnd.n1408 585
R3897 gnd.n6079 gnd.n6078 585
R3898 gnd.n6077 gnd.n1407 585
R3899 gnd.n6076 gnd.n1406 585
R3900 gnd.n6081 gnd.n1406 585
R3901 gnd.n6075 gnd.n6074 585
R3902 gnd.n6073 gnd.n6072 585
R3903 gnd.n6071 gnd.n6070 585
R3904 gnd.n6069 gnd.n6068 585
R3905 gnd.n6067 gnd.n6066 585
R3906 gnd.n6065 gnd.n6064 585
R3907 gnd.n6063 gnd.n6062 585
R3908 gnd.n6061 gnd.n6060 585
R3909 gnd.n6059 gnd.n6058 585
R3910 gnd.n6057 gnd.n6056 585
R3911 gnd.n6055 gnd.n6054 585
R3912 gnd.n6053 gnd.n6052 585
R3913 gnd.n6051 gnd.n6050 585
R3914 gnd.n6049 gnd.n6048 585
R3915 gnd.n6047 gnd.n6046 585
R3916 gnd.n6044 gnd.n6043 585
R3917 gnd.n6042 gnd.n6041 585
R3918 gnd.n6040 gnd.n6039 585
R3919 gnd.n6038 gnd.n6037 585
R3920 gnd.n6036 gnd.n6035 585
R3921 gnd.n6034 gnd.n6033 585
R3922 gnd.n6032 gnd.n6031 585
R3923 gnd.n6030 gnd.n6029 585
R3924 gnd.n6027 gnd.n6026 585
R3925 gnd.n6025 gnd.n6024 585
R3926 gnd.n6023 gnd.n6022 585
R3927 gnd.n6021 gnd.n6020 585
R3928 gnd.n6019 gnd.n6018 585
R3929 gnd.n6017 gnd.n6016 585
R3930 gnd.n6015 gnd.n6014 585
R3931 gnd.n6013 gnd.n6012 585
R3932 gnd.n6011 gnd.n6010 585
R3933 gnd.n6009 gnd.n6008 585
R3934 gnd.n6007 gnd.n6006 585
R3935 gnd.n6005 gnd.n6004 585
R3936 gnd.n6003 gnd.n6002 585
R3937 gnd.n6001 gnd.n6000 585
R3938 gnd.n5999 gnd.n5998 585
R3939 gnd.n5997 gnd.n5996 585
R3940 gnd.n5995 gnd.n5994 585
R3941 gnd.n5993 gnd.n5992 585
R3942 gnd.n5991 gnd.n5990 585
R3943 gnd.n5989 gnd.n5988 585
R3944 gnd.n5987 gnd.n5986 585
R3945 gnd.n5985 gnd.n5984 585
R3946 gnd.n5983 gnd.n5982 585
R3947 gnd.n5981 gnd.n5980 585
R3948 gnd.n5979 gnd.n5978 585
R3949 gnd.n5977 gnd.n5976 585
R3950 gnd.n5975 gnd.n5974 585
R3951 gnd.n5973 gnd.n5972 585
R3952 gnd.n5971 gnd.n5970 585
R3953 gnd.n5969 gnd.n5968 585
R3954 gnd.n5963 gnd.n5962 585
R3955 gnd.n7427 gnd.n7426 585
R3956 gnd.n7429 gnd.n315 585
R3957 gnd.n7431 gnd.n7430 585
R3958 gnd.n7432 gnd.n308 585
R3959 gnd.n7434 gnd.n7433 585
R3960 gnd.n7436 gnd.n306 585
R3961 gnd.n7438 gnd.n7437 585
R3962 gnd.n7439 gnd.n301 585
R3963 gnd.n7441 gnd.n7440 585
R3964 gnd.n7443 gnd.n299 585
R3965 gnd.n7445 gnd.n7444 585
R3966 gnd.n7446 gnd.n294 585
R3967 gnd.n7448 gnd.n7447 585
R3968 gnd.n7450 gnd.n292 585
R3969 gnd.n7452 gnd.n7451 585
R3970 gnd.n7453 gnd.n287 585
R3971 gnd.n7455 gnd.n7454 585
R3972 gnd.n7457 gnd.n286 585
R3973 gnd.n7458 gnd.n283 585
R3974 gnd.n7461 gnd.n7460 585
R3975 gnd.n285 gnd.n279 585
R3976 gnd.n7465 gnd.n276 585
R3977 gnd.n7467 gnd.n7466 585
R3978 gnd.n7469 gnd.n274 585
R3979 gnd.n7471 gnd.n7470 585
R3980 gnd.n7472 gnd.n269 585
R3981 gnd.n7474 gnd.n7473 585
R3982 gnd.n7476 gnd.n267 585
R3983 gnd.n7478 gnd.n7477 585
R3984 gnd.n7479 gnd.n262 585
R3985 gnd.n7481 gnd.n7480 585
R3986 gnd.n7483 gnd.n260 585
R3987 gnd.n7485 gnd.n7484 585
R3988 gnd.n7486 gnd.n255 585
R3989 gnd.n7488 gnd.n7487 585
R3990 gnd.n7490 gnd.n253 585
R3991 gnd.n7492 gnd.n7491 585
R3992 gnd.n7493 gnd.n248 585
R3993 gnd.n7495 gnd.n7494 585
R3994 gnd.n7497 gnd.n246 585
R3995 gnd.n7499 gnd.n7498 585
R3996 gnd.n7503 gnd.n241 585
R3997 gnd.n7505 gnd.n7504 585
R3998 gnd.n7507 gnd.n239 585
R3999 gnd.n7509 gnd.n7508 585
R4000 gnd.n7510 gnd.n234 585
R4001 gnd.n7512 gnd.n7511 585
R4002 gnd.n7514 gnd.n232 585
R4003 gnd.n7516 gnd.n7515 585
R4004 gnd.n7517 gnd.n227 585
R4005 gnd.n7519 gnd.n7518 585
R4006 gnd.n7521 gnd.n225 585
R4007 gnd.n7523 gnd.n7522 585
R4008 gnd.n7524 gnd.n220 585
R4009 gnd.n7526 gnd.n7525 585
R4010 gnd.n7528 gnd.n218 585
R4011 gnd.n7530 gnd.n7529 585
R4012 gnd.n7531 gnd.n216 585
R4013 gnd.n7532 gnd.n213 585
R4014 gnd.n213 gnd.n212 585
R4015 gnd.n7309 gnd.n210 585
R4016 gnd.n7537 gnd.n210 585
R4017 gnd.n7311 gnd.n7310 585
R4018 gnd.n7310 gnd.n209 585
R4019 gnd.n7312 gnd.n202 585
R4020 gnd.n7543 gnd.n202 585
R4021 gnd.n7314 gnd.n7313 585
R4022 gnd.n7313 gnd.n194 585
R4023 gnd.n7315 gnd.n192 585
R4024 gnd.n7549 gnd.n192 585
R4025 gnd.n7317 gnd.n7316 585
R4026 gnd.n7316 gnd.n191 585
R4027 gnd.n7318 gnd.n182 585
R4028 gnd.n7555 gnd.n182 585
R4029 gnd.n7320 gnd.n7319 585
R4030 gnd.n7319 gnd.n174 585
R4031 gnd.n7321 gnd.n172 585
R4032 gnd.n7561 gnd.n172 585
R4033 gnd.n7323 gnd.n7322 585
R4034 gnd.n7322 gnd.n171 585
R4035 gnd.n7324 gnd.n163 585
R4036 gnd.n7567 gnd.n163 585
R4037 gnd.n7326 gnd.n7325 585
R4038 gnd.n7325 gnd.n162 585
R4039 gnd.n7327 gnd.n153 585
R4040 gnd.n7573 gnd.n153 585
R4041 gnd.n7329 gnd.n7328 585
R4042 gnd.n7328 gnd.n146 585
R4043 gnd.n7330 gnd.n144 585
R4044 gnd.n7579 gnd.n144 585
R4045 gnd.n7332 gnd.n7331 585
R4046 gnd.n7331 gnd.n136 585
R4047 gnd.n7333 gnd.n134 585
R4048 gnd.n7585 gnd.n134 585
R4049 gnd.n7335 gnd.n7334 585
R4050 gnd.n7334 gnd.n133 585
R4051 gnd.n7336 gnd.n125 585
R4052 gnd.n7591 gnd.n125 585
R4053 gnd.n7338 gnd.n7337 585
R4054 gnd.n7337 gnd.n124 585
R4055 gnd.n7339 gnd.n116 585
R4056 gnd.n7597 gnd.n116 585
R4057 gnd.n7341 gnd.n7340 585
R4058 gnd.n7340 gnd.n107 585
R4059 gnd.n7342 gnd.n105 585
R4060 gnd.n7603 gnd.n105 585
R4061 gnd.n7344 gnd.n7343 585
R4062 gnd.n7345 gnd.n7344 585
R4063 gnd.n370 gnd.n369 585
R4064 gnd.n369 gnd.n368 585
R4065 gnd.n7293 gnd.n89 585
R4066 gnd.n7611 gnd.n89 585
R4067 gnd.n7295 gnd.n7294 585
R4068 gnd.n7296 gnd.n7295 585
R4069 gnd.n7292 gnd.n376 585
R4070 gnd.n7283 gnd.n376 585
R4071 gnd.n382 gnd.n377 585
R4072 gnd.n7287 gnd.n382 585
R4073 gnd.n5854 gnd.n5853 585
R4074 gnd.n5853 gnd.n1597 585
R4075 gnd.n5855 gnd.n1595 585
R4076 gnd.n5888 gnd.n1595 585
R4077 gnd.n5856 gnd.n1591 585
R4078 gnd.n5892 gnd.n1591 585
R4079 gnd.n5858 gnd.n5857 585
R4080 gnd.n5859 gnd.n5858 585
R4081 gnd.n5851 gnd.n1581 585
R4082 gnd.n5898 gnd.n1581 585
R4083 gnd.n5850 gnd.n1604 585
R4084 gnd.n5875 gnd.n1604 585
R4085 gnd.n5848 gnd.n1571 585
R4086 gnd.n5904 gnd.n1571 585
R4087 gnd.n5847 gnd.n5846 585
R4088 gnd.n5846 gnd.n5845 585
R4089 gnd.n1609 gnd.n1561 585
R4090 gnd.n5910 gnd.n1561 585
R4091 gnd.n5836 gnd.n5835 585
R4092 gnd.n5837 gnd.n5836 585
R4093 gnd.n5833 gnd.n1551 585
R4094 gnd.n5916 gnd.n1551 585
R4095 gnd.n5832 gnd.n5831 585
R4096 gnd.n5831 gnd.n5830 585
R4097 gnd.n1614 gnd.n1541 585
R4098 gnd.n5922 gnd.n1541 585
R4099 gnd.n5755 gnd.n1618 585
R4100 gnd.n5822 gnd.n1618 585
R4101 gnd.n5756 gnd.n1531 585
R4102 gnd.n5928 gnd.n1531 585
R4103 gnd.n5758 gnd.n5757 585
R4104 gnd.n5759 gnd.n5758 585
R4105 gnd.n5753 gnd.n1521 585
R4106 gnd.n5934 gnd.n1521 585
R4107 gnd.n5752 gnd.n5751 585
R4108 gnd.n5751 gnd.n5750 585
R4109 gnd.n5747 gnd.n1511 585
R4110 gnd.n5940 gnd.n1511 585
R4111 gnd.n5746 gnd.n5745 585
R4112 gnd.n5745 gnd.n5744 585
R4113 gnd.n5743 gnd.n1498 585
R4114 gnd.n5946 gnd.n1498 585
R4115 gnd.n1482 gnd.n1481 585
R4116 gnd.n5737 gnd.n1482 585
R4117 gnd.n5954 gnd.n5953 585
R4118 gnd.n5953 gnd.n5952 585
R4119 gnd.n5955 gnd.n1471 585
R4120 gnd.n5776 gnd.n1471 585
R4121 gnd.n5961 gnd.n1472 585
R4122 gnd.n5961 gnd.n5960 585
R4123 gnd.n6474 gnd.n6473 585
R4124 gnd.n6473 gnd.n6472 585
R4125 gnd.n7275 gnd.n7274 585
R4126 gnd.n7274 gnd.n90 585
R4127 gnd.n7278 gnd.n388 585
R4128 gnd.n388 gnd.n375 585
R4129 gnd.n7280 gnd.n7279 585
R4130 gnd.n7281 gnd.n7280 585
R4131 gnd.n389 gnd.n387 585
R4132 gnd.n387 gnd.n381 585
R4133 gnd.n5886 gnd.n5885 585
R4134 gnd.n5887 gnd.n5886 585
R4135 gnd.n1599 gnd.n1598 585
R4136 gnd.n1598 gnd.n1594 585
R4137 gnd.n5880 gnd.n5879 585
R4138 gnd.n5879 gnd.n1590 585
R4139 gnd.n5878 gnd.n1601 585
R4140 gnd.n5878 gnd.n1583 585
R4141 gnd.n5877 gnd.n1603 585
R4142 gnd.n5877 gnd.n5876 585
R4143 gnd.n5809 gnd.n1602 585
R4144 gnd.n1602 gnd.n1573 585
R4145 gnd.n5811 gnd.n5810 585
R4146 gnd.n5810 gnd.n1570 585
R4147 gnd.n5812 gnd.n5802 585
R4148 gnd.n5802 gnd.n1563 585
R4149 gnd.n5814 gnd.n5813 585
R4150 gnd.n5814 gnd.n1560 585
R4151 gnd.n5815 gnd.n5801 585
R4152 gnd.n5815 gnd.n1613 585
R4153 gnd.n5817 gnd.n5816 585
R4154 gnd.n5816 gnd.n1550 585
R4155 gnd.n5818 gnd.n1620 585
R4156 gnd.n1620 gnd.n1543 585
R4157 gnd.n5820 gnd.n5819 585
R4158 gnd.n5821 gnd.n5820 585
R4159 gnd.n1621 gnd.n1619 585
R4160 gnd.n1619 gnd.n1533 585
R4161 gnd.n5795 gnd.n5794 585
R4162 gnd.n5794 gnd.n1530 585
R4163 gnd.n5793 gnd.n1623 585
R4164 gnd.n5793 gnd.n1523 585
R4165 gnd.n5792 gnd.n5791 585
R4166 gnd.n5792 gnd.n1520 585
R4167 gnd.n1625 gnd.n1624 585
R4168 gnd.n5749 gnd.n1624 585
R4169 gnd.n5787 gnd.n5786 585
R4170 gnd.n5786 gnd.n1510 585
R4171 gnd.n5785 gnd.n1627 585
R4172 gnd.n5785 gnd.n1500 585
R4173 gnd.n5784 gnd.n5783 585
R4174 gnd.n5784 gnd.n1497 585
R4175 gnd.n1629 gnd.n1628 585
R4176 gnd.n1628 gnd.n1484 585
R4177 gnd.n5779 gnd.n5778 585
R4178 gnd.n5778 gnd.n5777 585
R4179 gnd.n1632 gnd.n1631 585
R4180 gnd.n1632 gnd.n1475 585
R4181 gnd.n5720 gnd.n5719 585
R4182 gnd.n5720 gnd.n1473 585
R4183 gnd.n5721 gnd.n5716 585
R4184 gnd.n5721 gnd.n1405 585
R4185 gnd.n5723 gnd.n5722 585
R4186 gnd.n5722 gnd.n1363 585
R4187 gnd.n5724 gnd.n1664 585
R4188 gnd.n1664 gnd.n1662 585
R4189 gnd.n5726 gnd.n5725 585
R4190 gnd.n5727 gnd.n5726 585
R4191 gnd.n1665 gnd.n1663 585
R4192 gnd.n1663 gnd.n1296 585
R4193 gnd.n5710 gnd.n1295 585
R4194 gnd.n6149 gnd.n1295 585
R4195 gnd.n5709 gnd.n5708 585
R4196 gnd.n5708 gnd.n1294 585
R4197 gnd.n5707 gnd.n1667 585
R4198 gnd.n5707 gnd.n5706 585
R4199 gnd.n5694 gnd.n1668 585
R4200 gnd.n1669 gnd.n1668 585
R4201 gnd.n5696 gnd.n5695 585
R4202 gnd.n5697 gnd.n5696 585
R4203 gnd.n1677 gnd.n1676 585
R4204 gnd.n1676 gnd.n1675 585
R4205 gnd.n5688 gnd.n5687 585
R4206 gnd.n5687 gnd.n5686 585
R4207 gnd.n1680 gnd.n1679 585
R4208 gnd.n1687 gnd.n1680 585
R4209 gnd.n5676 gnd.n5675 585
R4210 gnd.n5677 gnd.n5676 585
R4211 gnd.n1689 gnd.n1688 585
R4212 gnd.n1688 gnd.n1686 585
R4213 gnd.n5671 gnd.n5670 585
R4214 gnd.n5670 gnd.n5669 585
R4215 gnd.n1692 gnd.n1691 585
R4216 gnd.n1693 gnd.n1692 585
R4217 gnd.n5659 gnd.n5658 585
R4218 gnd.n5660 gnd.n5659 585
R4219 gnd.n1701 gnd.n1700 585
R4220 gnd.n1700 gnd.n1699 585
R4221 gnd.n5654 gnd.n5653 585
R4222 gnd.n5653 gnd.n5652 585
R4223 gnd.n1704 gnd.n1703 585
R4224 gnd.n1705 gnd.n1704 585
R4225 gnd.n5642 gnd.n5641 585
R4226 gnd.n5643 gnd.n5642 585
R4227 gnd.n1713 gnd.n1712 585
R4228 gnd.n1712 gnd.n1711 585
R4229 gnd.n5637 gnd.n5636 585
R4230 gnd.n5636 gnd.n5635 585
R4231 gnd.n1716 gnd.n1715 585
R4232 gnd.n1717 gnd.n1716 585
R4233 gnd.n5625 gnd.n5624 585
R4234 gnd.n5626 gnd.n5625 585
R4235 gnd.n1724 gnd.n1723 585
R4236 gnd.n1747 gnd.n1723 585
R4237 gnd.n5620 gnd.n5619 585
R4238 gnd.n5619 gnd.n5618 585
R4239 gnd.n1727 gnd.n1726 585
R4240 gnd.n5415 gnd.n1727 585
R4241 gnd.n5449 gnd.n1779 585
R4242 gnd.n1779 gnd.n1770 585
R4243 gnd.n5451 gnd.n5450 585
R4244 gnd.n5452 gnd.n5451 585
R4245 gnd.n1780 gnd.n1778 585
R4246 gnd.n5427 gnd.n1778 585
R4247 gnd.n5444 gnd.n5443 585
R4248 gnd.n5443 gnd.n5442 585
R4249 gnd.n1783 gnd.n1782 585
R4250 gnd.n1790 gnd.n1783 585
R4251 gnd.n5406 gnd.n5405 585
R4252 gnd.n5407 gnd.n5406 585
R4253 gnd.n1804 gnd.n1803 585
R4254 gnd.n1812 gnd.n1803 585
R4255 gnd.n5401 gnd.n5400 585
R4256 gnd.n5400 gnd.n5399 585
R4257 gnd.n1807 gnd.n1806 585
R4258 gnd.n1817 gnd.n1807 585
R4259 gnd.n5366 gnd.n1833 585
R4260 gnd.n1833 gnd.n1823 585
R4261 gnd.n5368 gnd.n5367 585
R4262 gnd.n5369 gnd.n5368 585
R4263 gnd.n1834 gnd.n1832 585
R4264 gnd.n1832 gnd.n1827 585
R4265 gnd.n5361 gnd.n5360 585
R4266 gnd.n5360 gnd.n5359 585
R4267 gnd.n1837 gnd.n1836 585
R4268 gnd.n5352 gnd.n1837 585
R4269 gnd.n5325 gnd.n1855 585
R4270 gnd.n5309 gnd.n1855 585
R4271 gnd.n5327 gnd.n5326 585
R4272 gnd.n5328 gnd.n5327 585
R4273 gnd.n1856 gnd.n1854 585
R4274 gnd.n1863 gnd.n1854 585
R4275 gnd.n5320 gnd.n5319 585
R4276 gnd.n5319 gnd.n5318 585
R4277 gnd.n1859 gnd.n1858 585
R4278 gnd.n5289 gnd.n1859 585
R4279 gnd.n5276 gnd.n1882 585
R4280 gnd.n5259 gnd.n1882 585
R4281 gnd.n5278 gnd.n5277 585
R4282 gnd.n5279 gnd.n5278 585
R4283 gnd.n1883 gnd.n1881 585
R4284 gnd.n1890 gnd.n1881 585
R4285 gnd.n5271 gnd.n5270 585
R4286 gnd.n5270 gnd.n5269 585
R4287 gnd.n1886 gnd.n1885 585
R4288 gnd.n1901 gnd.n1886 585
R4289 gnd.n5239 gnd.n5238 585
R4290 gnd.n5240 gnd.n5239 585
R4291 gnd.n1909 gnd.n1908 585
R4292 gnd.n1916 gnd.n1908 585
R4293 gnd.n5234 gnd.n5233 585
R4294 gnd.n5233 gnd.n5232 585
R4295 gnd.n1912 gnd.n1911 585
R4296 gnd.n1920 gnd.n1912 585
R4297 gnd.n5201 gnd.n1936 585
R4298 gnd.n1936 gnd.n1926 585
R4299 gnd.n5203 gnd.n5202 585
R4300 gnd.n5204 gnd.n5203 585
R4301 gnd.n1937 gnd.n1935 585
R4302 gnd.n1935 gnd.n1931 585
R4303 gnd.n5196 gnd.n5195 585
R4304 gnd.n5195 gnd.n5194 585
R4305 gnd.n1940 gnd.n1939 585
R4306 gnd.n5186 gnd.n1940 585
R4307 gnd.n5164 gnd.n5163 585
R4308 gnd.n5163 gnd.n5162 585
R4309 gnd.n5165 gnd.n1960 585
R4310 gnd.n1966 gnd.n1960 585
R4311 gnd.n5167 gnd.n5166 585
R4312 gnd.n5168 gnd.n5167 585
R4313 gnd.n1961 gnd.n1959 585
R4314 gnd.n5127 gnd.n1959 585
R4315 gnd.n5103 gnd.n5102 585
R4316 gnd.n5102 gnd.n1973 585
R4317 gnd.n5104 gnd.n1986 585
R4318 gnd.n1986 gnd.n1979 585
R4319 gnd.n5106 gnd.n5105 585
R4320 gnd.n5107 gnd.n5106 585
R4321 gnd.n1987 gnd.n1985 585
R4322 gnd.n1993 gnd.n1985 585
R4323 gnd.n5095 gnd.n5094 585
R4324 gnd.n5094 gnd.n5093 585
R4325 gnd.n1990 gnd.n1989 585
R4326 gnd.n1999 gnd.n1990 585
R4327 gnd.n5062 gnd.n2014 585
R4328 gnd.n2014 gnd.n2005 585
R4329 gnd.n5064 gnd.n5063 585
R4330 gnd.n5065 gnd.n5064 585
R4331 gnd.n2015 gnd.n2013 585
R4332 gnd.n2013 gnd.n2009 585
R4333 gnd.n5057 gnd.n5056 585
R4334 gnd.n5056 gnd.n5055 585
R4335 gnd.n2018 gnd.n2017 585
R4336 gnd.n5046 gnd.n2018 585
R4337 gnd.n5033 gnd.n5032 585
R4338 gnd.n5034 gnd.n5033 585
R4339 gnd.n5028 gnd.n5027 585
R4340 gnd.n5027 gnd.n5026 585
R4341 gnd.n1194 gnd.n1193 585
R4342 gnd.n4970 gnd.n1194 585
R4343 gnd.n6268 gnd.n6267 585
R4344 gnd.n6267 gnd.n6266 585
R4345 gnd.n6269 gnd.n1188 585
R4346 gnd.n4990 gnd.n1188 585
R4347 gnd.n6271 gnd.n6270 585
R4348 gnd.n6272 gnd.n6271 585
R4349 gnd.n1189 gnd.n1187 585
R4350 gnd.n1187 gnd.n1183 585
R4351 gnd.n4878 gnd.n4877 585
R4352 gnd.n4877 gnd.n1157 585
R4353 gnd.n4879 gnd.n2044 585
R4354 gnd.n2044 gnd.n1125 585
R4355 gnd.n4881 gnd.n4880 585
R4356 gnd.n4882 gnd.n4881 585
R4357 gnd.n2045 gnd.n2043 585
R4358 gnd.n2043 gnd.n2041 585
R4359 gnd.n4870 gnd.n4869 585
R4360 gnd.n4869 gnd.n4868 585
R4361 gnd.n2048 gnd.n2047 585
R4362 gnd.n2049 gnd.n2048 585
R4363 gnd.n4845 gnd.n4844 585
R4364 gnd.n4846 gnd.n4845 585
R4365 gnd.n2060 gnd.n2059 585
R4366 gnd.n2066 gnd.n2059 585
R4367 gnd.n4840 gnd.n4839 585
R4368 gnd.n4839 gnd.n4838 585
R4369 gnd.n2063 gnd.n2062 585
R4370 gnd.n2064 gnd.n2063 585
R4371 gnd.n4829 gnd.n4828 585
R4372 gnd.n4830 gnd.n4829 585
R4373 gnd.n2074 gnd.n2073 585
R4374 gnd.n2080 gnd.n2073 585
R4375 gnd.n4824 gnd.n4823 585
R4376 gnd.n4823 gnd.n4822 585
R4377 gnd.n2077 gnd.n2076 585
R4378 gnd.n2078 gnd.n2077 585
R4379 gnd.n4813 gnd.n4812 585
R4380 gnd.n4814 gnd.n4813 585
R4381 gnd.n2089 gnd.n2088 585
R4382 gnd.n2088 gnd.n2086 585
R4383 gnd.n4808 gnd.n4807 585
R4384 gnd.n4807 gnd.n4806 585
R4385 gnd.n2092 gnd.n2091 585
R4386 gnd.n2093 gnd.n2092 585
R4387 gnd.n4797 gnd.n4796 585
R4388 gnd.n4798 gnd.n4797 585
R4389 gnd.n2103 gnd.n2102 585
R4390 gnd.n2102 gnd.n2100 585
R4391 gnd.n4792 gnd.n4791 585
R4392 gnd.n4791 gnd.n4790 585
R4393 gnd.n2106 gnd.n2105 585
R4394 gnd.n2114 gnd.n2106 585
R4395 gnd.n4781 gnd.n4780 585
R4396 gnd.n4782 gnd.n4781 585
R4397 gnd.n2116 gnd.n2115 585
R4398 gnd.n2115 gnd.n2112 585
R4399 gnd.n4776 gnd.n4775 585
R4400 gnd.n4775 gnd.n4774 585
R4401 gnd.n2119 gnd.n2118 585
R4402 gnd.n2120 gnd.n2119 585
R4403 gnd.n4655 gnd.n4651 585
R4404 gnd.n4651 gnd.n4650 585
R4405 gnd.n4658 gnd.n4656 585
R4406 gnd.n4658 gnd.n4657 585
R4407 gnd.n4659 gnd.n4649 585
R4408 gnd.n4659 gnd.n1068 585
R4409 gnd.n4661 gnd.n4660 585
R4410 gnd.n4660 gnd.n1065 585
R4411 gnd.n4662 gnd.n4644 585
R4412 gnd.n4644 gnd.n2383 585
R4413 gnd.n4664 gnd.n4663 585
R4414 gnd.n4664 gnd.n1057 585
R4415 gnd.n4665 gnd.n4643 585
R4416 gnd.n4665 gnd.n1049 585
R4417 gnd.n4667 gnd.n4666 585
R4418 gnd.n4666 gnd.n1046 585
R4419 gnd.n4668 gnd.n2393 585
R4420 gnd.n2393 gnd.n1039 585
R4421 gnd.n4670 gnd.n4669 585
R4422 gnd.n4671 gnd.n4670 585
R4423 gnd.n2394 gnd.n2392 585
R4424 gnd.n2392 gnd.n1029 585
R4425 gnd.n4637 gnd.n4636 585
R4426 gnd.n4636 gnd.n1026 585
R4427 gnd.n4635 gnd.n2396 585
R4428 gnd.n4635 gnd.n1019 585
R4429 gnd.n4634 gnd.n4633 585
R4430 gnd.n4634 gnd.n1016 585
R4431 gnd.n2398 gnd.n2397 585
R4432 gnd.n4600 gnd.n2397 585
R4433 gnd.n4629 gnd.n4628 585
R4434 gnd.n4628 gnd.n1006 585
R4435 gnd.n4627 gnd.n2400 585
R4436 gnd.n4627 gnd.n999 585
R4437 gnd.n4626 gnd.n2402 585
R4438 gnd.n4626 gnd.n4625 585
R4439 gnd.n4552 gnd.n2401 585
R4440 gnd.n2401 gnd.n989 585
R4441 gnd.n4554 gnd.n4553 585
R4442 gnd.n4553 gnd.n986 585
R4443 gnd.n4555 gnd.n4545 585
R4444 gnd.n4545 gnd.n979 585
R4445 gnd.n4557 gnd.n4556 585
R4446 gnd.n4557 gnd.n976 585
R4447 gnd.n4558 gnd.n4544 585
R4448 gnd.n4558 gnd.n2416 585
R4449 gnd.n4560 gnd.n4559 585
R4450 gnd.n4559 gnd.n967 585
R4451 gnd.n4561 gnd.n2425 585
R4452 gnd.n2425 gnd.n958 585
R4453 gnd.n4563 gnd.n4562 585
R4454 gnd.n4564 gnd.n4563 585
R4455 gnd.n2426 gnd.n2424 585
R4456 gnd.n2424 gnd.n2422 585
R4457 gnd.n4538 gnd.n4537 585
R4458 gnd.n4537 gnd.n4536 585
R4459 gnd.n2431 gnd.n2430 585
R4460 gnd.n2439 gnd.n2431 585
R4461 gnd.n2427 gnd.n937 585
R4462 gnd.n2436 gnd.n937 585
R4463 gnd.n6148 gnd.n6147 585
R4464 gnd.n6149 gnd.n6148 585
R4465 gnd.n1299 gnd.n1297 585
R4466 gnd.n1297 gnd.n1294 585
R4467 gnd.n5704 gnd.n5703 585
R4468 gnd.n5706 gnd.n5704 585
R4469 gnd.n1671 gnd.n1670 585
R4470 gnd.n1670 gnd.n1669 585
R4471 gnd.n5699 gnd.n5698 585
R4472 gnd.n5698 gnd.n5697 585
R4473 gnd.n1674 gnd.n1673 585
R4474 gnd.n1675 gnd.n1674 585
R4475 gnd.n5684 gnd.n5683 585
R4476 gnd.n5686 gnd.n5684 585
R4477 gnd.n1682 gnd.n1681 585
R4478 gnd.n1687 gnd.n1681 585
R4479 gnd.n5679 gnd.n5678 585
R4480 gnd.n5678 gnd.n5677 585
R4481 gnd.n1685 gnd.n1684 585
R4482 gnd.n1686 gnd.n1685 585
R4483 gnd.n5667 gnd.n5666 585
R4484 gnd.n5669 gnd.n5667 585
R4485 gnd.n1695 gnd.n1694 585
R4486 gnd.n1694 gnd.n1693 585
R4487 gnd.n5662 gnd.n5661 585
R4488 gnd.n5661 gnd.n5660 585
R4489 gnd.n1698 gnd.n1697 585
R4490 gnd.n1699 gnd.n1698 585
R4491 gnd.n5650 gnd.n5649 585
R4492 gnd.n5652 gnd.n5650 585
R4493 gnd.n1707 gnd.n1706 585
R4494 gnd.n1706 gnd.n1705 585
R4495 gnd.n5645 gnd.n5644 585
R4496 gnd.n5644 gnd.n5643 585
R4497 gnd.n1710 gnd.n1709 585
R4498 gnd.n1711 gnd.n1710 585
R4499 gnd.n5633 gnd.n5632 585
R4500 gnd.n5635 gnd.n5633 585
R4501 gnd.n1719 gnd.n1718 585
R4502 gnd.n1718 gnd.n1717 585
R4503 gnd.n5628 gnd.n5627 585
R4504 gnd.n5627 gnd.n5626 585
R4505 gnd.n1722 gnd.n1721 585
R4506 gnd.n1747 gnd.n1722 585
R4507 gnd.n5418 gnd.n1729 585
R4508 gnd.n5618 gnd.n1729 585
R4509 gnd.n5419 gnd.n5416 585
R4510 gnd.n5416 gnd.n5415 585
R4511 gnd.n5420 gnd.n5414 585
R4512 gnd.n5414 gnd.n1770 585
R4513 gnd.n1797 gnd.n1775 585
R4514 gnd.n5452 gnd.n1775 585
R4515 gnd.n5425 gnd.n5424 585
R4516 gnd.n5427 gnd.n5425 585
R4517 gnd.n1796 gnd.n1785 585
R4518 gnd.n5442 gnd.n1785 585
R4519 gnd.n5410 gnd.n5409 585
R4520 gnd.n5409 gnd.n1790 585
R4521 gnd.n5408 gnd.n1799 585
R4522 gnd.n5408 gnd.n5407 585
R4523 gnd.n5339 gnd.n1800 585
R4524 gnd.n1812 gnd.n1800 585
R4525 gnd.n5340 gnd.n1809 585
R4526 gnd.n5399 gnd.n1809 585
R4527 gnd.n5337 gnd.n5336 585
R4528 gnd.n5336 gnd.n1817 585
R4529 gnd.n5344 gnd.n5335 585
R4530 gnd.n5335 gnd.n1823 585
R4531 gnd.n5345 gnd.n1829 585
R4532 gnd.n5369 gnd.n1829 585
R4533 gnd.n5346 gnd.n5334 585
R4534 gnd.n5334 gnd.n1827 585
R4535 gnd.n1849 gnd.n1839 585
R4536 gnd.n5359 gnd.n1839 585
R4537 gnd.n5351 gnd.n5350 585
R4538 gnd.n5352 gnd.n5351 585
R4539 gnd.n1848 gnd.n1847 585
R4540 gnd.n5309 gnd.n1847 585
R4541 gnd.n5330 gnd.n5329 585
R4542 gnd.n5329 gnd.n5328 585
R4543 gnd.n1852 gnd.n1851 585
R4544 gnd.n1863 gnd.n1852 585
R4545 gnd.n1876 gnd.n1861 585
R4546 gnd.n5318 gnd.n1861 585
R4547 gnd.n5287 gnd.n5286 585
R4548 gnd.n5289 gnd.n5287 585
R4549 gnd.n1875 gnd.n1874 585
R4550 gnd.n5259 gnd.n1874 585
R4551 gnd.n5281 gnd.n5280 585
R4552 gnd.n5280 gnd.n5279 585
R4553 gnd.n1879 gnd.n1878 585
R4554 gnd.n1890 gnd.n1879 585
R4555 gnd.n5143 gnd.n1888 585
R4556 gnd.n5269 gnd.n1888 585
R4557 gnd.n5144 gnd.n5142 585
R4558 gnd.n5142 gnd.n1901 585
R4559 gnd.n5140 gnd.n1906 585
R4560 gnd.n5240 gnd.n1906 585
R4561 gnd.n5148 gnd.n5139 585
R4562 gnd.n5139 gnd.n1916 585
R4563 gnd.n5149 gnd.n1914 585
R4564 gnd.n5232 gnd.n1914 585
R4565 gnd.n5150 gnd.n5138 585
R4566 gnd.n5138 gnd.n1920 585
R4567 gnd.n5137 gnd.n5135 585
R4568 gnd.n5137 gnd.n1926 585
R4569 gnd.n5154 gnd.n1933 585
R4570 gnd.n5204 gnd.n1933 585
R4571 gnd.n5155 gnd.n5134 585
R4572 gnd.n5134 gnd.n1931 585
R4573 gnd.n5156 gnd.n1941 585
R4574 gnd.n5194 gnd.n1941 585
R4575 gnd.n1969 gnd.n1949 585
R4576 gnd.n5186 gnd.n1949 585
R4577 gnd.n5161 gnd.n5160 585
R4578 gnd.n5162 gnd.n5161 585
R4579 gnd.n1968 gnd.n1967 585
R4580 gnd.n1967 gnd.n1966 585
R4581 gnd.n5130 gnd.n1956 585
R4582 gnd.n5168 gnd.n1956 585
R4583 gnd.n5129 gnd.n5128 585
R4584 gnd.n5128 gnd.n5127 585
R4585 gnd.n1972 gnd.n1971 585
R4586 gnd.n1973 gnd.n1972 585
R4587 gnd.n5007 gnd.n5006 585
R4588 gnd.n5006 gnd.n1979 585
R4589 gnd.n5008 gnd.n1984 585
R4590 gnd.n5107 gnd.n1984 585
R4591 gnd.n5003 gnd.n5002 585
R4592 gnd.n5002 gnd.n1993 585
R4593 gnd.n5012 gnd.n1991 585
R4594 gnd.n5093 gnd.n1991 585
R4595 gnd.n5013 gnd.n5001 585
R4596 gnd.n5001 gnd.n1999 585
R4597 gnd.n5014 gnd.n5000 585
R4598 gnd.n5000 gnd.n2005 585
R4599 gnd.n4998 gnd.n2011 585
R4600 gnd.n5065 gnd.n2011 585
R4601 gnd.n5018 gnd.n4997 585
R4602 gnd.n4997 gnd.n2009 585
R4603 gnd.n5019 gnd.n2019 585
R4604 gnd.n5055 gnd.n2019 585
R4605 gnd.n5020 gnd.n2026 585
R4606 gnd.n5046 gnd.n2026 585
R4607 gnd.n2034 gnd.n2030 585
R4608 gnd.n5034 gnd.n2030 585
R4609 gnd.n5025 gnd.n5024 585
R4610 gnd.n5026 gnd.n5025 585
R4611 gnd.n2033 gnd.n2032 585
R4612 gnd.n4970 gnd.n2032 585
R4613 gnd.n4993 gnd.n1195 585
R4614 gnd.n6266 gnd.n1195 585
R4615 gnd.n4992 gnd.n4991 585
R4616 gnd.n4991 gnd.n4990 585
R4617 gnd.n4891 gnd.n1185 585
R4618 gnd.n6272 gnd.n1185 585
R4619 gnd.n4885 gnd.n2036 585
R4620 gnd.n4885 gnd.n1183 585
R4621 gnd.n4887 gnd.n4886 585
R4622 gnd.n4886 gnd.n1157 585
R4623 gnd.n4884 gnd.n2038 585
R4624 gnd.n4884 gnd.n1125 585
R4625 gnd.n4883 gnd.n2040 585
R4626 gnd.n4883 gnd.n4882 585
R4627 gnd.n2154 gnd.n2039 585
R4628 gnd.n2041 gnd.n2039 585
R4629 gnd.n2158 gnd.n2050 585
R4630 gnd.n4868 gnd.n2050 585
R4631 gnd.n2159 gnd.n2153 585
R4632 gnd.n2153 gnd.n2049 585
R4633 gnd.n2160 gnd.n2058 585
R4634 gnd.n4846 gnd.n2058 585
R4635 gnd.n2151 gnd.n2150 585
R4636 gnd.n2150 gnd.n2066 585
R4637 gnd.n2164 gnd.n2065 585
R4638 gnd.n4838 gnd.n2065 585
R4639 gnd.n2165 gnd.n2149 585
R4640 gnd.n2149 gnd.n2064 585
R4641 gnd.n2166 gnd.n2072 585
R4642 gnd.n4830 gnd.n2072 585
R4643 gnd.n2147 gnd.n2146 585
R4644 gnd.n2146 gnd.n2080 585
R4645 gnd.n2170 gnd.n2079 585
R4646 gnd.n4822 gnd.n2079 585
R4647 gnd.n2171 gnd.n2145 585
R4648 gnd.n2145 gnd.n2078 585
R4649 gnd.n2172 gnd.n2087 585
R4650 gnd.n4814 gnd.n2087 585
R4651 gnd.n2143 gnd.n2142 585
R4652 gnd.n2142 gnd.n2086 585
R4653 gnd.n2176 gnd.n2094 585
R4654 gnd.n4806 gnd.n2094 585
R4655 gnd.n2177 gnd.n2141 585
R4656 gnd.n2141 gnd.n2093 585
R4657 gnd.n2178 gnd.n2101 585
R4658 gnd.n4798 gnd.n2101 585
R4659 gnd.n2139 gnd.n2138 585
R4660 gnd.n2138 gnd.n2100 585
R4661 gnd.n2182 gnd.n2107 585
R4662 gnd.n4790 gnd.n2107 585
R4663 gnd.n2183 gnd.n2137 585
R4664 gnd.n2137 gnd.n2114 585
R4665 gnd.n2184 gnd.n2113 585
R4666 gnd.n4782 gnd.n2113 585
R4667 gnd.n4771 gnd.n4770 585
R4668 gnd.n4769 gnd.n2135 585
R4669 gnd.n2187 gnd.n2134 585
R4670 gnd.n4773 gnd.n2134 585
R4671 gnd.n4765 gnd.n2189 585
R4672 gnd.n4764 gnd.n2190 585
R4673 gnd.n4763 gnd.n2191 585
R4674 gnd.n2307 gnd.n2192 585
R4675 gnd.n4758 gnd.n2308 585
R4676 gnd.n4757 gnd.n2309 585
R4677 gnd.n4756 gnd.n2310 585
R4678 gnd.n2320 gnd.n2311 585
R4679 gnd.n4749 gnd.n2321 585
R4680 gnd.n4748 gnd.n2322 585
R4681 gnd.n2324 gnd.n2323 585
R4682 gnd.n4741 gnd.n2332 585
R4683 gnd.n4740 gnd.n2333 585
R4684 gnd.n2343 gnd.n2334 585
R4685 gnd.n4733 gnd.n2344 585
R4686 gnd.n4732 gnd.n2345 585
R4687 gnd.n2347 gnd.n2346 585
R4688 gnd.n4725 gnd.n2355 585
R4689 gnd.n4724 gnd.n2356 585
R4690 gnd.n2366 gnd.n2357 585
R4691 gnd.n4717 gnd.n2367 585
R4692 gnd.n4716 gnd.n2368 585
R4693 gnd.n4701 gnd.n4700 585
R4694 gnd.n4703 gnd.n4702 585
R4695 gnd.n4706 gnd.n4704 585
R4696 gnd.n4705 gnd.n2111 585
R4697 gnd.n6151 gnd.n6150 585
R4698 gnd.n6150 gnd.n6149 585
R4699 gnd.n6152 gnd.n1292 585
R4700 gnd.n1294 gnd.n1292 585
R4701 gnd.n5705 gnd.n1290 585
R4702 gnd.n5706 gnd.n5705 585
R4703 gnd.n6156 gnd.n1289 585
R4704 gnd.n1669 gnd.n1289 585
R4705 gnd.n6157 gnd.n1288 585
R4706 gnd.n5697 gnd.n1288 585
R4707 gnd.n6158 gnd.n1287 585
R4708 gnd.n1675 gnd.n1287 585
R4709 gnd.n5685 gnd.n1285 585
R4710 gnd.n5686 gnd.n5685 585
R4711 gnd.n6162 gnd.n1284 585
R4712 gnd.n1687 gnd.n1284 585
R4713 gnd.n6163 gnd.n1283 585
R4714 gnd.n5677 gnd.n1283 585
R4715 gnd.n6164 gnd.n1282 585
R4716 gnd.n1686 gnd.n1282 585
R4717 gnd.n5668 gnd.n1280 585
R4718 gnd.n5669 gnd.n5668 585
R4719 gnd.n6168 gnd.n1279 585
R4720 gnd.n1693 gnd.n1279 585
R4721 gnd.n6169 gnd.n1278 585
R4722 gnd.n5660 gnd.n1278 585
R4723 gnd.n6170 gnd.n1277 585
R4724 gnd.n1699 gnd.n1277 585
R4725 gnd.n5651 gnd.n1275 585
R4726 gnd.n5652 gnd.n5651 585
R4727 gnd.n6174 gnd.n1274 585
R4728 gnd.n1705 gnd.n1274 585
R4729 gnd.n6175 gnd.n1273 585
R4730 gnd.n5643 gnd.n1273 585
R4731 gnd.n6176 gnd.n1272 585
R4732 gnd.n1711 gnd.n1272 585
R4733 gnd.n5634 gnd.n1270 585
R4734 gnd.n5635 gnd.n5634 585
R4735 gnd.n6180 gnd.n1269 585
R4736 gnd.n1717 gnd.n1269 585
R4737 gnd.n6181 gnd.n1268 585
R4738 gnd.n5626 gnd.n1268 585
R4739 gnd.n6182 gnd.n1267 585
R4740 gnd.n1747 gnd.n1267 585
R4741 gnd.n5617 gnd.n1265 585
R4742 gnd.n5618 gnd.n5617 585
R4743 gnd.n6186 gnd.n1264 585
R4744 gnd.n5415 gnd.n1264 585
R4745 gnd.n6187 gnd.n1263 585
R4746 gnd.n1770 gnd.n1263 585
R4747 gnd.n6188 gnd.n1262 585
R4748 gnd.n5452 gnd.n1262 585
R4749 gnd.n5426 gnd.n1260 585
R4750 gnd.n5427 gnd.n5426 585
R4751 gnd.n6192 gnd.n1259 585
R4752 gnd.n5442 gnd.n1259 585
R4753 gnd.n6193 gnd.n1258 585
R4754 gnd.n1790 gnd.n1258 585
R4755 gnd.n6194 gnd.n1257 585
R4756 gnd.n5407 gnd.n1257 585
R4757 gnd.n1811 gnd.n1255 585
R4758 gnd.n1812 gnd.n1811 585
R4759 gnd.n6198 gnd.n1254 585
R4760 gnd.n5399 gnd.n1254 585
R4761 gnd.n6199 gnd.n1253 585
R4762 gnd.n1817 gnd.n1253 585
R4763 gnd.n6200 gnd.n1252 585
R4764 gnd.n1823 gnd.n1252 585
R4765 gnd.n1831 gnd.n1250 585
R4766 gnd.n5369 gnd.n1831 585
R4767 gnd.n6204 gnd.n1249 585
R4768 gnd.n1827 gnd.n1249 585
R4769 gnd.n6205 gnd.n1248 585
R4770 gnd.n5359 gnd.n1248 585
R4771 gnd.n6206 gnd.n1247 585
R4772 gnd.n5352 gnd.n1247 585
R4773 gnd.n5308 gnd.n1245 585
R4774 gnd.n5309 gnd.n5308 585
R4775 gnd.n6210 gnd.n1244 585
R4776 gnd.n5328 gnd.n1244 585
R4777 gnd.n6211 gnd.n1243 585
R4778 gnd.n1863 gnd.n1243 585
R4779 gnd.n6212 gnd.n1242 585
R4780 gnd.n5318 gnd.n1242 585
R4781 gnd.n5288 gnd.n1240 585
R4782 gnd.n5289 gnd.n5288 585
R4783 gnd.n6216 gnd.n1239 585
R4784 gnd.n5259 gnd.n1239 585
R4785 gnd.n6217 gnd.n1238 585
R4786 gnd.n5279 gnd.n1238 585
R4787 gnd.n6218 gnd.n1237 585
R4788 gnd.n1890 gnd.n1237 585
R4789 gnd.n5268 gnd.n1235 585
R4790 gnd.n5269 gnd.n5268 585
R4791 gnd.n6222 gnd.n1234 585
R4792 gnd.n1901 gnd.n1234 585
R4793 gnd.n6223 gnd.n1233 585
R4794 gnd.n5240 gnd.n1233 585
R4795 gnd.n6224 gnd.n1232 585
R4796 gnd.n1916 gnd.n1232 585
R4797 gnd.n5231 gnd.n1230 585
R4798 gnd.n5232 gnd.n5231 585
R4799 gnd.n6228 gnd.n1229 585
R4800 gnd.n1920 gnd.n1229 585
R4801 gnd.n6229 gnd.n1228 585
R4802 gnd.n1926 gnd.n1228 585
R4803 gnd.n6230 gnd.n1227 585
R4804 gnd.n5204 gnd.n1227 585
R4805 gnd.n1930 gnd.n1225 585
R4806 gnd.n1931 gnd.n1930 585
R4807 gnd.n6234 gnd.n1224 585
R4808 gnd.n5194 gnd.n1224 585
R4809 gnd.n6235 gnd.n1223 585
R4810 gnd.n5186 gnd.n1223 585
R4811 gnd.n6236 gnd.n1222 585
R4812 gnd.n5162 gnd.n1222 585
R4813 gnd.n1965 gnd.n1220 585
R4814 gnd.n1966 gnd.n1965 585
R4815 gnd.n6240 gnd.n1219 585
R4816 gnd.n5168 gnd.n1219 585
R4817 gnd.n6241 gnd.n1218 585
R4818 gnd.n5127 gnd.n1218 585
R4819 gnd.n6242 gnd.n1217 585
R4820 gnd.n1973 gnd.n1217 585
R4821 gnd.n1978 gnd.n1215 585
R4822 gnd.n1979 gnd.n1978 585
R4823 gnd.n6246 gnd.n1214 585
R4824 gnd.n5107 gnd.n1214 585
R4825 gnd.n6247 gnd.n1213 585
R4826 gnd.n1993 gnd.n1213 585
R4827 gnd.n6248 gnd.n1212 585
R4828 gnd.n5093 gnd.n1212 585
R4829 gnd.n1998 gnd.n1210 585
R4830 gnd.n1999 gnd.n1998 585
R4831 gnd.n6252 gnd.n1209 585
R4832 gnd.n2005 gnd.n1209 585
R4833 gnd.n6253 gnd.n1208 585
R4834 gnd.n5065 gnd.n1208 585
R4835 gnd.n6254 gnd.n1207 585
R4836 gnd.n2009 gnd.n1207 585
R4837 gnd.n5054 gnd.n1205 585
R4838 gnd.n5055 gnd.n5054 585
R4839 gnd.n6258 gnd.n1204 585
R4840 gnd.n5046 gnd.n1204 585
R4841 gnd.n6259 gnd.n1203 585
R4842 gnd.n5034 gnd.n1203 585
R4843 gnd.n6260 gnd.n1202 585
R4844 gnd.n5026 gnd.n1202 585
R4845 gnd.n1199 gnd.n1197 585
R4846 gnd.n4970 gnd.n1197 585
R4847 gnd.n6265 gnd.n6264 585
R4848 gnd.n6266 gnd.n6265 585
R4849 gnd.n1198 gnd.n1196 585
R4850 gnd.n4990 gnd.n1196 585
R4851 gnd.n4856 gnd.n1186 585
R4852 gnd.n6272 gnd.n1186 585
R4853 gnd.n4855 gnd.n4854 585
R4854 gnd.n4854 gnd.n1183 585
R4855 gnd.n4860 gnd.n4853 585
R4856 gnd.n4853 gnd.n1157 585
R4857 gnd.n4861 gnd.n4852 585
R4858 gnd.n4852 gnd.n1125 585
R4859 gnd.n4862 gnd.n2042 585
R4860 gnd.n4882 gnd.n2042 585
R4861 gnd.n2054 gnd.n2052 585
R4862 gnd.n2052 gnd.n2041 585
R4863 gnd.n4867 gnd.n4866 585
R4864 gnd.n4868 gnd.n4867 585
R4865 gnd.n2053 gnd.n2051 585
R4866 gnd.n2051 gnd.n2049 585
R4867 gnd.n4848 gnd.n4847 585
R4868 gnd.n4847 gnd.n4846 585
R4869 gnd.n2057 gnd.n2056 585
R4870 gnd.n2066 gnd.n2057 585
R4871 gnd.n4837 gnd.n4836 585
R4872 gnd.n4838 gnd.n4837 585
R4873 gnd.n2068 gnd.n2067 585
R4874 gnd.n2067 gnd.n2064 585
R4875 gnd.n4832 gnd.n4831 585
R4876 gnd.n4831 gnd.n4830 585
R4877 gnd.n2071 gnd.n2070 585
R4878 gnd.n2080 gnd.n2071 585
R4879 gnd.n4821 gnd.n4820 585
R4880 gnd.n4822 gnd.n4821 585
R4881 gnd.n2082 gnd.n2081 585
R4882 gnd.n2081 gnd.n2078 585
R4883 gnd.n4816 gnd.n4815 585
R4884 gnd.n4815 gnd.n4814 585
R4885 gnd.n2085 gnd.n2084 585
R4886 gnd.n2086 gnd.n2085 585
R4887 gnd.n4805 gnd.n4804 585
R4888 gnd.n4806 gnd.n4805 585
R4889 gnd.n2096 gnd.n2095 585
R4890 gnd.n2095 gnd.n2093 585
R4891 gnd.n4800 gnd.n4799 585
R4892 gnd.n4799 gnd.n4798 585
R4893 gnd.n2099 gnd.n2098 585
R4894 gnd.n2100 gnd.n2099 585
R4895 gnd.n4789 gnd.n4788 585
R4896 gnd.n4790 gnd.n4789 585
R4897 gnd.n2109 gnd.n2108 585
R4898 gnd.n2114 gnd.n2108 585
R4899 gnd.n4784 gnd.n4783 585
R4900 gnd.n4783 gnd.n4782 585
R4901 gnd.n6090 gnd.n1354 585
R4902 gnd.n5728 gnd.n1354 585
R4903 gnd.n6091 gnd.n1353 585
R4904 gnd.n1657 gnd.n1347 585
R4905 gnd.n6098 gnd.n1346 585
R4906 gnd.n6099 gnd.n1345 585
R4907 gnd.n1654 gnd.n1339 585
R4908 gnd.n6106 gnd.n1338 585
R4909 gnd.n6107 gnd.n1337 585
R4910 gnd.n1652 gnd.n1331 585
R4911 gnd.n6114 gnd.n1330 585
R4912 gnd.n6115 gnd.n1329 585
R4913 gnd.n1649 gnd.n1323 585
R4914 gnd.n6122 gnd.n1322 585
R4915 gnd.n6123 gnd.n1321 585
R4916 gnd.n1647 gnd.n1314 585
R4917 gnd.n6130 gnd.n1313 585
R4918 gnd.n6131 gnd.n1312 585
R4919 gnd.n1644 gnd.n1309 585
R4920 gnd.n6136 gnd.n1308 585
R4921 gnd.n6137 gnd.n1307 585
R4922 gnd.n6138 gnd.n1306 585
R4923 gnd.n1641 gnd.n1304 585
R4924 gnd.n6142 gnd.n1303 585
R4925 gnd.n6143 gnd.n1302 585
R4926 gnd.n6144 gnd.n1298 585
R4927 gnd.n5731 gnd.n1293 585
R4928 gnd.n5732 gnd.n5730 585
R4929 gnd.n1639 gnd.n1638 585
R4930 gnd.n1660 gnd.n1659 585
R4931 gnd.n5541 gnd.n1772 511.721
R4932 gnd.n5550 gnd.n5549 511.721
R4933 gnd.n4962 gnd.n4960 511.721
R4934 gnd.n6341 gnd.n1160 511.721
R4935 gnd.n6640 gnd.n766 466.675
R4936 gnd.n4896 gnd.t151 389.64
R4937 gnd.n1765 gnd.t101 389.64
R4938 gnd.n6278 gnd.t72 389.64
R4939 gnd.n5475 gnd.t157 389.64
R4940 gnd.n2369 gnd.t116 371.625
R4941 gnd.n6084 gnd.t76 371.625
R4942 gnd.n2376 gnd.t112 371.625
R4943 gnd.n1427 gnd.t173 371.625
R4944 gnd.n1450 gnd.t176 371.625
R4945 gnd.n5964 gnd.t126 371.625
R4946 gnd.n313 gnd.t154 371.625
R4947 gnd.n280 gnd.t105 371.625
R4948 gnd.n7500 gnd.t148 371.625
R4949 gnd.n350 gnd.t94 371.625
R4950 gnd.n4101 gnd.t129 371.625
R4951 gnd.n4123 gnd.t132 371.625
R4952 gnd.n4144 gnd.t80 371.625
R4953 gnd.n4162 gnd.t163 371.625
R4954 gnd.n1101 gnd.t141 371.625
R4955 gnd.n2194 gnd.t166 371.625
R4956 gnd.n2216 gnd.t186 371.625
R4957 gnd.n1355 gnd.t90 371.625
R4958 gnd.n3062 gnd.t108 323.425
R4959 gnd.n2604 gnd.t144 323.425
R4960 gnd.n3911 gnd.n3885 289.615
R4961 gnd.n3879 gnd.n3853 289.615
R4962 gnd.n3847 gnd.n3821 289.615
R4963 gnd.n3816 gnd.n3790 289.615
R4964 gnd.n3784 gnd.n3758 289.615
R4965 gnd.n3752 gnd.n3726 289.615
R4966 gnd.n3720 gnd.n3694 289.615
R4967 gnd.n3689 gnd.n3663 289.615
R4968 gnd.n3136 gnd.t182 279.217
R4969 gnd.n2630 gnd.t169 279.217
R4970 gnd.n1167 gnd.t89 260.649
R4971 gnd.n5467 gnd.t122 260.649
R4972 gnd.n6343 gnd.n6342 256.663
R4973 gnd.n6343 gnd.n1126 256.663
R4974 gnd.n6343 gnd.n1127 256.663
R4975 gnd.n6343 gnd.n1128 256.663
R4976 gnd.n6343 gnd.n1129 256.663
R4977 gnd.n6343 gnd.n1130 256.663
R4978 gnd.n6343 gnd.n1131 256.663
R4979 gnd.n6343 gnd.n1132 256.663
R4980 gnd.n6343 gnd.n1133 256.663
R4981 gnd.n6343 gnd.n1134 256.663
R4982 gnd.n6343 gnd.n1135 256.663
R4983 gnd.n6343 gnd.n1136 256.663
R4984 gnd.n6343 gnd.n1137 256.663
R4985 gnd.n6343 gnd.n1138 256.663
R4986 gnd.n6343 gnd.n1139 256.663
R4987 gnd.n6343 gnd.n1140 256.663
R4988 gnd.n6346 gnd.n1123 256.663
R4989 gnd.n6344 gnd.n6343 256.663
R4990 gnd.n6343 gnd.n1141 256.663
R4991 gnd.n6343 gnd.n1142 256.663
R4992 gnd.n6343 gnd.n1143 256.663
R4993 gnd.n6343 gnd.n1144 256.663
R4994 gnd.n6343 gnd.n1145 256.663
R4995 gnd.n6343 gnd.n1146 256.663
R4996 gnd.n6343 gnd.n1147 256.663
R4997 gnd.n6343 gnd.n1148 256.663
R4998 gnd.n6343 gnd.n1149 256.663
R4999 gnd.n6343 gnd.n1150 256.663
R5000 gnd.n6343 gnd.n1151 256.663
R5001 gnd.n6343 gnd.n1152 256.663
R5002 gnd.n6343 gnd.n1153 256.663
R5003 gnd.n6343 gnd.n1154 256.663
R5004 gnd.n6343 gnd.n1155 256.663
R5005 gnd.n6343 gnd.n1156 256.663
R5006 gnd.n5616 gnd.n1748 256.663
R5007 gnd.n5616 gnd.n1749 256.663
R5008 gnd.n5616 gnd.n1750 256.663
R5009 gnd.n5616 gnd.n1751 256.663
R5010 gnd.n5616 gnd.n1752 256.663
R5011 gnd.n5616 gnd.n1753 256.663
R5012 gnd.n5616 gnd.n1754 256.663
R5013 gnd.n5616 gnd.n1755 256.663
R5014 gnd.n5616 gnd.n1756 256.663
R5015 gnd.n5616 gnd.n1757 256.663
R5016 gnd.n5616 gnd.n1758 256.663
R5017 gnd.n5616 gnd.n1759 256.663
R5018 gnd.n5616 gnd.n1760 256.663
R5019 gnd.n5616 gnd.n1761 256.663
R5020 gnd.n5616 gnd.n1762 256.663
R5021 gnd.n5616 gnd.n1763 256.663
R5022 gnd.n1764 gnd.n1437 256.663
R5023 gnd.n5616 gnd.n1746 256.663
R5024 gnd.n5616 gnd.n1745 256.663
R5025 gnd.n5616 gnd.n1744 256.663
R5026 gnd.n5616 gnd.n1743 256.663
R5027 gnd.n5616 gnd.n1742 256.663
R5028 gnd.n5616 gnd.n1741 256.663
R5029 gnd.n5616 gnd.n1740 256.663
R5030 gnd.n5616 gnd.n1739 256.663
R5031 gnd.n5616 gnd.n1738 256.663
R5032 gnd.n5616 gnd.n1737 256.663
R5033 gnd.n5616 gnd.n1736 256.663
R5034 gnd.n5616 gnd.n1735 256.663
R5035 gnd.n5616 gnd.n1734 256.663
R5036 gnd.n5616 gnd.n1733 256.663
R5037 gnd.n5616 gnd.n1732 256.663
R5038 gnd.n5616 gnd.n1731 256.663
R5039 gnd.n5616 gnd.n1730 256.663
R5040 gnd.n4357 gnd.n4071 242.672
R5041 gnd.n4357 gnd.n4072 242.672
R5042 gnd.n4357 gnd.n4073 242.672
R5043 gnd.n4357 gnd.n4074 242.672
R5044 gnd.n4357 gnd.n4075 242.672
R5045 gnd.n4357 gnd.n4076 242.672
R5046 gnd.n4357 gnd.n4077 242.672
R5047 gnd.n4357 gnd.n4078 242.672
R5048 gnd.n4357 gnd.n4079 242.672
R5049 gnd.n4709 gnd.n1073 242.672
R5050 gnd.n2374 gnd.n1073 242.672
R5051 gnd.n2362 gnd.n1073 242.672
R5052 gnd.n2359 gnd.n1073 242.672
R5053 gnd.n2350 gnd.n1073 242.672
R5054 gnd.n2339 gnd.n1073 242.672
R5055 gnd.n2336 gnd.n1073 242.672
R5056 gnd.n2327 gnd.n1073 242.672
R5057 gnd.n2316 gnd.n1073 242.672
R5058 gnd.n3190 gnd.n3189 242.672
R5059 gnd.n3190 gnd.n3100 242.672
R5060 gnd.n3190 gnd.n3101 242.672
R5061 gnd.n3190 gnd.n3102 242.672
R5062 gnd.n3190 gnd.n3103 242.672
R5063 gnd.n3190 gnd.n3104 242.672
R5064 gnd.n3190 gnd.n3105 242.672
R5065 gnd.n3190 gnd.n3106 242.672
R5066 gnd.n3190 gnd.n3107 242.672
R5067 gnd.n3190 gnd.n3108 242.672
R5068 gnd.n3190 gnd.n3109 242.672
R5069 gnd.n3190 gnd.n3110 242.672
R5070 gnd.n3191 gnd.n3190 242.672
R5071 gnd.n4043 gnd.n2579 242.672
R5072 gnd.n4043 gnd.n2578 242.672
R5073 gnd.n4043 gnd.n2577 242.672
R5074 gnd.n4043 gnd.n2576 242.672
R5075 gnd.n4043 gnd.n2575 242.672
R5076 gnd.n4043 gnd.n2574 242.672
R5077 gnd.n4043 gnd.n2573 242.672
R5078 gnd.n4043 gnd.n2572 242.672
R5079 gnd.n4043 gnd.n2571 242.672
R5080 gnd.n4043 gnd.n2570 242.672
R5081 gnd.n4043 gnd.n2569 242.672
R5082 gnd.n4043 gnd.n2568 242.672
R5083 gnd.n4043 gnd.n2567 242.672
R5084 gnd.n6081 gnd.n1392 242.672
R5085 gnd.n6081 gnd.n1394 242.672
R5086 gnd.n6081 gnd.n1395 242.672
R5087 gnd.n6081 gnd.n1397 242.672
R5088 gnd.n6081 gnd.n1399 242.672
R5089 gnd.n6081 gnd.n1400 242.672
R5090 gnd.n6081 gnd.n1402 242.672
R5091 gnd.n6081 gnd.n1404 242.672
R5092 gnd.n6082 gnd.n6081 242.672
R5093 gnd.n347 gnd.n212 242.672
R5094 gnd.n7396 gnd.n212 242.672
R5095 gnd.n343 gnd.n212 242.672
R5096 gnd.n7403 gnd.n212 242.672
R5097 gnd.n336 gnd.n212 242.672
R5098 gnd.n7410 gnd.n212 242.672
R5099 gnd.n329 gnd.n212 242.672
R5100 gnd.n7417 gnd.n212 242.672
R5101 gnd.n322 gnd.n212 242.672
R5102 gnd.n3274 gnd.n3273 242.672
R5103 gnd.n3273 gnd.n3012 242.672
R5104 gnd.n3273 gnd.n3013 242.672
R5105 gnd.n3273 gnd.n3014 242.672
R5106 gnd.n3273 gnd.n3015 242.672
R5107 gnd.n3273 gnd.n3016 242.672
R5108 gnd.n3273 gnd.n3017 242.672
R5109 gnd.n3273 gnd.n3018 242.672
R5110 gnd.n4043 gnd.n2580 242.672
R5111 gnd.n4043 gnd.n2581 242.672
R5112 gnd.n4043 gnd.n2582 242.672
R5113 gnd.n4043 gnd.n2583 242.672
R5114 gnd.n4043 gnd.n2584 242.672
R5115 gnd.n4043 gnd.n2585 242.672
R5116 gnd.n4043 gnd.n2586 242.672
R5117 gnd.n4043 gnd.n2587 242.672
R5118 gnd.n4357 gnd.n4356 242.672
R5119 gnd.n4357 gnd.n4044 242.672
R5120 gnd.n4357 gnd.n4045 242.672
R5121 gnd.n4357 gnd.n4046 242.672
R5122 gnd.n4357 gnd.n4047 242.672
R5123 gnd.n4357 gnd.n4048 242.672
R5124 gnd.n4357 gnd.n4049 242.672
R5125 gnd.n4357 gnd.n4050 242.672
R5126 gnd.n4357 gnd.n4051 242.672
R5127 gnd.n4357 gnd.n4052 242.672
R5128 gnd.n4357 gnd.n4053 242.672
R5129 gnd.n4357 gnd.n4054 242.672
R5130 gnd.n4357 gnd.n4055 242.672
R5131 gnd.n4357 gnd.n4056 242.672
R5132 gnd.n4357 gnd.n4057 242.672
R5133 gnd.n4357 gnd.n4058 242.672
R5134 gnd.n4357 gnd.n4059 242.672
R5135 gnd.n4357 gnd.n4060 242.672
R5136 gnd.n4357 gnd.n4061 242.672
R5137 gnd.n4357 gnd.n4062 242.672
R5138 gnd.n4357 gnd.n4063 242.672
R5139 gnd.n4357 gnd.n4064 242.672
R5140 gnd.n4357 gnd.n4065 242.672
R5141 gnd.n4357 gnd.n4066 242.672
R5142 gnd.n4357 gnd.n4067 242.672
R5143 gnd.n4357 gnd.n4068 242.672
R5144 gnd.n4357 gnd.n4069 242.672
R5145 gnd.n4357 gnd.n4070 242.672
R5146 gnd.n4358 gnd.n4357 242.672
R5147 gnd.n2301 gnd.n1073 242.672
R5148 gnd.n2197 gnd.n1073 242.672
R5149 gnd.n2291 gnd.n1073 242.672
R5150 gnd.n2201 gnd.n1073 242.672
R5151 gnd.n2281 gnd.n1073 242.672
R5152 gnd.n2205 gnd.n1073 242.672
R5153 gnd.n2271 gnd.n1073 242.672
R5154 gnd.n2209 gnd.n1073 242.672
R5155 gnd.n2261 gnd.n1073 242.672
R5156 gnd.n2213 gnd.n1073 242.672
R5157 gnd.n2251 gnd.n1073 242.672
R5158 gnd.n2219 gnd.n1073 242.672
R5159 gnd.n2241 gnd.n1073 242.672
R5160 gnd.n2223 gnd.n1073 242.672
R5161 gnd.n2231 gnd.n1073 242.672
R5162 gnd.n2228 gnd.n1073 242.672
R5163 gnd.n6347 gnd.n1119 242.672
R5164 gnd.n1118 gnd.n1073 242.672
R5165 gnd.n6351 gnd.n1073 242.672
R5166 gnd.n1112 gnd.n1073 242.672
R5167 gnd.n6358 gnd.n1073 242.672
R5168 gnd.n1105 gnd.n1073 242.672
R5169 gnd.n6366 gnd.n1073 242.672
R5170 gnd.n1096 gnd.n1073 242.672
R5171 gnd.n6373 gnd.n1073 242.672
R5172 gnd.n1089 gnd.n1073 242.672
R5173 gnd.n6380 gnd.n1073 242.672
R5174 gnd.n1082 gnd.n1073 242.672
R5175 gnd.n6387 gnd.n1073 242.672
R5176 gnd.n6390 gnd.n1073 242.672
R5177 gnd.n6081 gnd.n6080 242.672
R5178 gnd.n6081 gnd.n1364 242.672
R5179 gnd.n6081 gnd.n1365 242.672
R5180 gnd.n6081 gnd.n1366 242.672
R5181 gnd.n6081 gnd.n1367 242.672
R5182 gnd.n6081 gnd.n1368 242.672
R5183 gnd.n6081 gnd.n1369 242.672
R5184 gnd.n6081 gnd.n1370 242.672
R5185 gnd.n6081 gnd.n1371 242.672
R5186 gnd.n6081 gnd.n1372 242.672
R5187 gnd.n6081 gnd.n1373 242.672
R5188 gnd.n6081 gnd.n1374 242.672
R5189 gnd.n6081 gnd.n1375 242.672
R5190 gnd.n6028 gnd.n1438 242.672
R5191 gnd.n6081 gnd.n1376 242.672
R5192 gnd.n6081 gnd.n1377 242.672
R5193 gnd.n6081 gnd.n1378 242.672
R5194 gnd.n6081 gnd.n1379 242.672
R5195 gnd.n6081 gnd.n1380 242.672
R5196 gnd.n6081 gnd.n1381 242.672
R5197 gnd.n6081 gnd.n1382 242.672
R5198 gnd.n6081 gnd.n1383 242.672
R5199 gnd.n6081 gnd.n1384 242.672
R5200 gnd.n6081 gnd.n1385 242.672
R5201 gnd.n6081 gnd.n1386 242.672
R5202 gnd.n6081 gnd.n1387 242.672
R5203 gnd.n6081 gnd.n1388 242.672
R5204 gnd.n6081 gnd.n1389 242.672
R5205 gnd.n6081 gnd.n1390 242.672
R5206 gnd.n6081 gnd.n1391 242.672
R5207 gnd.n7428 gnd.n212 242.672
R5208 gnd.n316 gnd.n212 242.672
R5209 gnd.n7435 gnd.n212 242.672
R5210 gnd.n307 gnd.n212 242.672
R5211 gnd.n7442 gnd.n212 242.672
R5212 gnd.n300 gnd.n212 242.672
R5213 gnd.n7449 gnd.n212 242.672
R5214 gnd.n293 gnd.n212 242.672
R5215 gnd.n7456 gnd.n212 242.672
R5216 gnd.n7459 gnd.n212 242.672
R5217 gnd.n284 gnd.n212 242.672
R5218 gnd.n7468 gnd.n212 242.672
R5219 gnd.n275 gnd.n212 242.672
R5220 gnd.n7475 gnd.n212 242.672
R5221 gnd.n268 gnd.n212 242.672
R5222 gnd.n7482 gnd.n212 242.672
R5223 gnd.n261 gnd.n212 242.672
R5224 gnd.n7489 gnd.n212 242.672
R5225 gnd.n254 gnd.n212 242.672
R5226 gnd.n7496 gnd.n212 242.672
R5227 gnd.n247 gnd.n212 242.672
R5228 gnd.n7506 gnd.n212 242.672
R5229 gnd.n240 gnd.n212 242.672
R5230 gnd.n7513 gnd.n212 242.672
R5231 gnd.n233 gnd.n212 242.672
R5232 gnd.n7520 gnd.n212 242.672
R5233 gnd.n226 gnd.n212 242.672
R5234 gnd.n7527 gnd.n212 242.672
R5235 gnd.n219 gnd.n212 242.672
R5236 gnd.n4773 gnd.n4772 242.672
R5237 gnd.n4773 gnd.n2121 242.672
R5238 gnd.n4773 gnd.n2122 242.672
R5239 gnd.n4773 gnd.n2123 242.672
R5240 gnd.n4773 gnd.n2124 242.672
R5241 gnd.n4773 gnd.n2125 242.672
R5242 gnd.n4773 gnd.n2126 242.672
R5243 gnd.n4773 gnd.n2127 242.672
R5244 gnd.n4773 gnd.n2128 242.672
R5245 gnd.n4773 gnd.n2129 242.672
R5246 gnd.n4773 gnd.n2130 242.672
R5247 gnd.n4773 gnd.n2131 242.672
R5248 gnd.n4773 gnd.n2132 242.672
R5249 gnd.n4773 gnd.n2133 242.672
R5250 gnd.n5728 gnd.n1658 242.672
R5251 gnd.n5728 gnd.n1656 242.672
R5252 gnd.n5728 gnd.n1655 242.672
R5253 gnd.n5728 gnd.n1653 242.672
R5254 gnd.n5728 gnd.n1651 242.672
R5255 gnd.n5728 gnd.n1650 242.672
R5256 gnd.n5728 gnd.n1648 242.672
R5257 gnd.n5728 gnd.n1646 242.672
R5258 gnd.n5728 gnd.n1645 242.672
R5259 gnd.n5728 gnd.n1643 242.672
R5260 gnd.n5728 gnd.n1642 242.672
R5261 gnd.n5728 gnd.n1640 242.672
R5262 gnd.n5729 gnd.n5728 242.672
R5263 gnd.n5728 gnd.n1661 242.672
R5264 gnd.n216 gnd.n213 240.244
R5265 gnd.n7529 gnd.n7528 240.244
R5266 gnd.n7526 gnd.n220 240.244
R5267 gnd.n7522 gnd.n7521 240.244
R5268 gnd.n7519 gnd.n227 240.244
R5269 gnd.n7515 gnd.n7514 240.244
R5270 gnd.n7512 gnd.n234 240.244
R5271 gnd.n7508 gnd.n7507 240.244
R5272 gnd.n7505 gnd.n241 240.244
R5273 gnd.n7498 gnd.n7497 240.244
R5274 gnd.n7495 gnd.n248 240.244
R5275 gnd.n7491 gnd.n7490 240.244
R5276 gnd.n7488 gnd.n255 240.244
R5277 gnd.n7484 gnd.n7483 240.244
R5278 gnd.n7481 gnd.n262 240.244
R5279 gnd.n7477 gnd.n7476 240.244
R5280 gnd.n7474 gnd.n269 240.244
R5281 gnd.n7470 gnd.n7469 240.244
R5282 gnd.n7467 gnd.n276 240.244
R5283 gnd.n7460 gnd.n285 240.244
R5284 gnd.n7458 gnd.n7457 240.244
R5285 gnd.n7455 gnd.n287 240.244
R5286 gnd.n7451 gnd.n7450 240.244
R5287 gnd.n7448 gnd.n294 240.244
R5288 gnd.n7444 gnd.n7443 240.244
R5289 gnd.n7441 gnd.n301 240.244
R5290 gnd.n7437 gnd.n7436 240.244
R5291 gnd.n7434 gnd.n308 240.244
R5292 gnd.n7430 gnd.n7429 240.244
R5293 gnd.n5961 gnd.n1471 240.244
R5294 gnd.n5953 gnd.n1471 240.244
R5295 gnd.n5953 gnd.n1482 240.244
R5296 gnd.n1498 gnd.n1482 240.244
R5297 gnd.n5745 gnd.n1498 240.244
R5298 gnd.n5745 gnd.n1511 240.244
R5299 gnd.n5751 gnd.n1511 240.244
R5300 gnd.n5751 gnd.n1521 240.244
R5301 gnd.n5758 gnd.n1521 240.244
R5302 gnd.n5758 gnd.n1531 240.244
R5303 gnd.n1618 gnd.n1531 240.244
R5304 gnd.n1618 gnd.n1541 240.244
R5305 gnd.n5831 gnd.n1541 240.244
R5306 gnd.n5831 gnd.n1551 240.244
R5307 gnd.n5836 gnd.n1551 240.244
R5308 gnd.n5836 gnd.n1561 240.244
R5309 gnd.n5846 gnd.n1561 240.244
R5310 gnd.n5846 gnd.n1571 240.244
R5311 gnd.n1604 gnd.n1571 240.244
R5312 gnd.n1604 gnd.n1581 240.244
R5313 gnd.n5858 gnd.n1581 240.244
R5314 gnd.n5858 gnd.n1591 240.244
R5315 gnd.n1595 gnd.n1591 240.244
R5316 gnd.n5853 gnd.n1595 240.244
R5317 gnd.n5853 gnd.n382 240.244
R5318 gnd.n382 gnd.n376 240.244
R5319 gnd.n7295 gnd.n376 240.244
R5320 gnd.n7295 gnd.n89 240.244
R5321 gnd.n369 gnd.n89 240.244
R5322 gnd.n7344 gnd.n369 240.244
R5323 gnd.n7344 gnd.n105 240.244
R5324 gnd.n7340 gnd.n105 240.244
R5325 gnd.n7340 gnd.n116 240.244
R5326 gnd.n7337 gnd.n116 240.244
R5327 gnd.n7337 gnd.n125 240.244
R5328 gnd.n7334 gnd.n125 240.244
R5329 gnd.n7334 gnd.n134 240.244
R5330 gnd.n7331 gnd.n134 240.244
R5331 gnd.n7331 gnd.n144 240.244
R5332 gnd.n7328 gnd.n144 240.244
R5333 gnd.n7328 gnd.n153 240.244
R5334 gnd.n7325 gnd.n153 240.244
R5335 gnd.n7325 gnd.n163 240.244
R5336 gnd.n7322 gnd.n163 240.244
R5337 gnd.n7322 gnd.n172 240.244
R5338 gnd.n7319 gnd.n172 240.244
R5339 gnd.n7319 gnd.n182 240.244
R5340 gnd.n7316 gnd.n182 240.244
R5341 gnd.n7316 gnd.n192 240.244
R5342 gnd.n7313 gnd.n192 240.244
R5343 gnd.n7313 gnd.n202 240.244
R5344 gnd.n7310 gnd.n202 240.244
R5345 gnd.n7310 gnd.n210 240.244
R5346 gnd.n1407 gnd.n1406 240.244
R5347 gnd.n6074 gnd.n1406 240.244
R5348 gnd.n6072 gnd.n6071 240.244
R5349 gnd.n6068 gnd.n6067 240.244
R5350 gnd.n6064 gnd.n6063 240.244
R5351 gnd.n6060 gnd.n6059 240.244
R5352 gnd.n6056 gnd.n6055 240.244
R5353 gnd.n6052 gnd.n6051 240.244
R5354 gnd.n6048 gnd.n6047 240.244
R5355 gnd.n6043 gnd.n6042 240.244
R5356 gnd.n6039 gnd.n6038 240.244
R5357 gnd.n6035 gnd.n6034 240.244
R5358 gnd.n6031 gnd.n6030 240.244
R5359 gnd.n6026 gnd.n6025 240.244
R5360 gnd.n6022 gnd.n6021 240.244
R5361 gnd.n6018 gnd.n6017 240.244
R5362 gnd.n6014 gnd.n6013 240.244
R5363 gnd.n6010 gnd.n6009 240.244
R5364 gnd.n6006 gnd.n6005 240.244
R5365 gnd.n6002 gnd.n6001 240.244
R5366 gnd.n5998 gnd.n5997 240.244
R5367 gnd.n5994 gnd.n5993 240.244
R5368 gnd.n5990 gnd.n5989 240.244
R5369 gnd.n5986 gnd.n5985 240.244
R5370 gnd.n5982 gnd.n5981 240.244
R5371 gnd.n5978 gnd.n5977 240.244
R5372 gnd.n5974 gnd.n5973 240.244
R5373 gnd.n5970 gnd.n5969 240.244
R5374 gnd.n1486 gnd.n1408 240.244
R5375 gnd.n5951 gnd.n1486 240.244
R5376 gnd.n5951 gnd.n1487 240.244
R5377 gnd.n5947 gnd.n1487 240.244
R5378 gnd.n5947 gnd.n1496 240.244
R5379 gnd.n5939 gnd.n1496 240.244
R5380 gnd.n5939 gnd.n1513 240.244
R5381 gnd.n5935 gnd.n1513 240.244
R5382 gnd.n5935 gnd.n1519 240.244
R5383 gnd.n5927 gnd.n1519 240.244
R5384 gnd.n5927 gnd.n1534 240.244
R5385 gnd.n5923 gnd.n1534 240.244
R5386 gnd.n5923 gnd.n1540 240.244
R5387 gnd.n5915 gnd.n1540 240.244
R5388 gnd.n5915 gnd.n1553 240.244
R5389 gnd.n5911 gnd.n1553 240.244
R5390 gnd.n5911 gnd.n1559 240.244
R5391 gnd.n5903 gnd.n1559 240.244
R5392 gnd.n5903 gnd.n1574 240.244
R5393 gnd.n5899 gnd.n1574 240.244
R5394 gnd.n5899 gnd.n1580 240.244
R5395 gnd.n5891 gnd.n1580 240.244
R5396 gnd.n5891 gnd.n5889 240.244
R5397 gnd.n5889 gnd.n384 240.244
R5398 gnd.n7286 gnd.n384 240.244
R5399 gnd.n7286 gnd.n7284 240.244
R5400 gnd.n7284 gnd.n92 240.244
R5401 gnd.n7610 gnd.n92 240.244
R5402 gnd.n7610 gnd.n93 240.244
R5403 gnd.n103 gnd.n93 240.244
R5404 gnd.n7604 gnd.n103 240.244
R5405 gnd.n7604 gnd.n104 240.244
R5406 gnd.n7596 gnd.n104 240.244
R5407 gnd.n7596 gnd.n118 240.244
R5408 gnd.n7592 gnd.n118 240.244
R5409 gnd.n7592 gnd.n123 240.244
R5410 gnd.n7584 gnd.n123 240.244
R5411 gnd.n7584 gnd.n137 240.244
R5412 gnd.n7580 gnd.n137 240.244
R5413 gnd.n7580 gnd.n143 240.244
R5414 gnd.n7572 gnd.n143 240.244
R5415 gnd.n7572 gnd.n155 240.244
R5416 gnd.n7568 gnd.n155 240.244
R5417 gnd.n7568 gnd.n161 240.244
R5418 gnd.n7560 gnd.n161 240.244
R5419 gnd.n7560 gnd.n175 240.244
R5420 gnd.n7556 gnd.n175 240.244
R5421 gnd.n7556 gnd.n181 240.244
R5422 gnd.n7548 gnd.n181 240.244
R5423 gnd.n7548 gnd.n195 240.244
R5424 gnd.n7544 gnd.n195 240.244
R5425 gnd.n7544 gnd.n201 240.244
R5426 gnd.n7536 gnd.n201 240.244
R5427 gnd.n6391 gnd.n1069 240.244
R5428 gnd.n6389 gnd.n6388 240.244
R5429 gnd.n6386 gnd.n1075 240.244
R5430 gnd.n6382 gnd.n6381 240.244
R5431 gnd.n6379 gnd.n1083 240.244
R5432 gnd.n6375 gnd.n6374 240.244
R5433 gnd.n6372 gnd.n1090 240.244
R5434 gnd.n6368 gnd.n6367 240.244
R5435 gnd.n6365 gnd.n1097 240.244
R5436 gnd.n6360 gnd.n6359 240.244
R5437 gnd.n6357 gnd.n1106 240.244
R5438 gnd.n6353 gnd.n6352 240.244
R5439 gnd.n6350 gnd.n1113 240.244
R5440 gnd.n2230 gnd.n2229 240.244
R5441 gnd.n2233 gnd.n2232 240.244
R5442 gnd.n2240 gnd.n2239 240.244
R5443 gnd.n2243 gnd.n2242 240.244
R5444 gnd.n2250 gnd.n2249 240.244
R5445 gnd.n2253 gnd.n2252 240.244
R5446 gnd.n2260 gnd.n2259 240.244
R5447 gnd.n2263 gnd.n2262 240.244
R5448 gnd.n2270 gnd.n2269 240.244
R5449 gnd.n2273 gnd.n2272 240.244
R5450 gnd.n2280 gnd.n2279 240.244
R5451 gnd.n2283 gnd.n2282 240.244
R5452 gnd.n2290 gnd.n2289 240.244
R5453 gnd.n2293 gnd.n2292 240.244
R5454 gnd.n2300 gnd.n2299 240.244
R5455 gnd.n4360 gnd.n2553 240.244
R5456 gnd.n2553 gnd.n2543 240.244
R5457 gnd.n4376 gnd.n2543 240.244
R5458 gnd.n4377 gnd.n4376 240.244
R5459 gnd.n4377 gnd.n2534 240.244
R5460 gnd.n2534 gnd.n2525 240.244
R5461 gnd.n4396 gnd.n2525 240.244
R5462 gnd.n4397 gnd.n4396 240.244
R5463 gnd.n4397 gnd.n2517 240.244
R5464 gnd.n2517 gnd.n2507 240.244
R5465 gnd.n4416 gnd.n2507 240.244
R5466 gnd.n4417 gnd.n4416 240.244
R5467 gnd.n4417 gnd.n2497 240.244
R5468 gnd.n4420 gnd.n2497 240.244
R5469 gnd.n4420 gnd.n2488 240.244
R5470 gnd.n2488 gnd.n2481 240.244
R5471 gnd.n4462 gnd.n2481 240.244
R5472 gnd.n4462 gnd.n2472 240.244
R5473 gnd.n2472 gnd.n2464 240.244
R5474 gnd.n4482 gnd.n2464 240.244
R5475 gnd.n4483 gnd.n4482 240.244
R5476 gnd.n4483 gnd.n2457 240.244
R5477 gnd.n2457 gnd.n2452 240.244
R5478 gnd.n4487 gnd.n2452 240.244
R5479 gnd.n4487 gnd.n939 240.244
R5480 gnd.n4517 gnd.n939 240.244
R5481 gnd.n4517 gnd.n2437 240.244
R5482 gnd.n4520 gnd.n2437 240.244
R5483 gnd.n4520 gnd.n2433 240.244
R5484 gnd.n2433 gnd.n2423 240.244
R5485 gnd.n2423 gnd.n956 240.244
R5486 gnd.n4574 gnd.n956 240.244
R5487 gnd.n4574 gnd.n968 240.244
R5488 gnd.n4579 gnd.n968 240.244
R5489 gnd.n4579 gnd.n977 240.244
R5490 gnd.n4589 gnd.n977 240.244
R5491 gnd.n4589 gnd.n987 240.244
R5492 gnd.n2403 gnd.n987 240.244
R5493 gnd.n2403 gnd.n997 240.244
R5494 gnd.n4596 gnd.n997 240.244
R5495 gnd.n4596 gnd.n1007 240.244
R5496 gnd.n4602 gnd.n1007 240.244
R5497 gnd.n4602 gnd.n1017 240.244
R5498 gnd.n4606 gnd.n1017 240.244
R5499 gnd.n4606 gnd.n1027 240.244
R5500 gnd.n4673 gnd.n1027 240.244
R5501 gnd.n4673 gnd.n1037 240.244
R5502 gnd.n4677 gnd.n1037 240.244
R5503 gnd.n4677 gnd.n1047 240.244
R5504 gnd.n4688 gnd.n1047 240.244
R5505 gnd.n4688 gnd.n1058 240.244
R5506 gnd.n4693 gnd.n1058 240.244
R5507 gnd.n4693 gnd.n1066 240.244
R5508 gnd.n4082 gnd.n4081 240.244
R5509 gnd.n4350 gnd.n4081 240.244
R5510 gnd.n4348 gnd.n4347 240.244
R5511 gnd.n4344 gnd.n4343 240.244
R5512 gnd.n4340 gnd.n4339 240.244
R5513 gnd.n4336 gnd.n4335 240.244
R5514 gnd.n4332 gnd.n4331 240.244
R5515 gnd.n4328 gnd.n4327 240.244
R5516 gnd.n4324 gnd.n4323 240.244
R5517 gnd.n4319 gnd.n4318 240.244
R5518 gnd.n4315 gnd.n4314 240.244
R5519 gnd.n4311 gnd.n4310 240.244
R5520 gnd.n4307 gnd.n4306 240.244
R5521 gnd.n4303 gnd.n4302 240.244
R5522 gnd.n4299 gnd.n4298 240.244
R5523 gnd.n4295 gnd.n4294 240.244
R5524 gnd.n4291 gnd.n4290 240.244
R5525 gnd.n4287 gnd.n4286 240.244
R5526 gnd.n4283 gnd.n4282 240.244
R5527 gnd.n4279 gnd.n4278 240.244
R5528 gnd.n4275 gnd.n4274 240.244
R5529 gnd.n4271 gnd.n4270 240.244
R5530 gnd.n4267 gnd.n4266 240.244
R5531 gnd.n4263 gnd.n4262 240.244
R5532 gnd.n4259 gnd.n4258 240.244
R5533 gnd.n4255 gnd.n4254 240.244
R5534 gnd.n4251 gnd.n4250 240.244
R5535 gnd.n4247 gnd.n4246 240.244
R5536 gnd.n4243 gnd.n2564 240.244
R5537 gnd.n4368 gnd.n2551 240.244
R5538 gnd.n4368 gnd.n2547 240.244
R5539 gnd.n4374 gnd.n2547 240.244
R5540 gnd.n4374 gnd.n2532 240.244
R5541 gnd.n4388 gnd.n2532 240.244
R5542 gnd.n4388 gnd.n2528 240.244
R5543 gnd.n4394 gnd.n2528 240.244
R5544 gnd.n4394 gnd.n2515 240.244
R5545 gnd.n4408 gnd.n2515 240.244
R5546 gnd.n4408 gnd.n2511 240.244
R5547 gnd.n4414 gnd.n2511 240.244
R5548 gnd.n4414 gnd.n2495 240.244
R5549 gnd.n4432 gnd.n2495 240.244
R5550 gnd.n4432 gnd.n2490 240.244
R5551 gnd.n4440 gnd.n2490 240.244
R5552 gnd.n4440 gnd.n2491 240.244
R5553 gnd.n2491 gnd.n2471 240.244
R5554 gnd.n4473 gnd.n2471 240.244
R5555 gnd.n4473 gnd.n2467 240.244
R5556 gnd.n4480 gnd.n2467 240.244
R5557 gnd.n4480 gnd.n2454 240.244
R5558 gnd.n4498 gnd.n2454 240.244
R5559 gnd.n4500 gnd.n4498 240.244
R5560 gnd.n4500 gnd.n942 240.244
R5561 gnd.n6470 gnd.n942 240.244
R5562 gnd.n6470 gnd.n943 240.244
R5563 gnd.n4530 gnd.n943 240.244
R5564 gnd.n4531 gnd.n4530 240.244
R5565 gnd.n4534 gnd.n4531 240.244
R5566 gnd.n4534 gnd.n954 240.244
R5567 gnd.n6465 gnd.n954 240.244
R5568 gnd.n6465 gnd.n955 240.244
R5569 gnd.n6457 gnd.n955 240.244
R5570 gnd.n6457 gnd.n970 240.244
R5571 gnd.n6453 gnd.n970 240.244
R5572 gnd.n6453 gnd.n975 240.244
R5573 gnd.n6445 gnd.n975 240.244
R5574 gnd.n6445 gnd.n990 240.244
R5575 gnd.n6441 gnd.n990 240.244
R5576 gnd.n6441 gnd.n996 240.244
R5577 gnd.n6433 gnd.n996 240.244
R5578 gnd.n6433 gnd.n1009 240.244
R5579 gnd.n6429 gnd.n1009 240.244
R5580 gnd.n6429 gnd.n1015 240.244
R5581 gnd.n6421 gnd.n1015 240.244
R5582 gnd.n6421 gnd.n1030 240.244
R5583 gnd.n6417 gnd.n1030 240.244
R5584 gnd.n6417 gnd.n1036 240.244
R5585 gnd.n6409 gnd.n1036 240.244
R5586 gnd.n6409 gnd.n1050 240.244
R5587 gnd.n6405 gnd.n1050 240.244
R5588 gnd.n6405 gnd.n1056 240.244
R5589 gnd.n6397 gnd.n1056 240.244
R5590 gnd.n4042 gnd.n2589 240.244
R5591 gnd.n4035 gnd.n4034 240.244
R5592 gnd.n4032 gnd.n4031 240.244
R5593 gnd.n4028 gnd.n4027 240.244
R5594 gnd.n4024 gnd.n4023 240.244
R5595 gnd.n4020 gnd.n4019 240.244
R5596 gnd.n4016 gnd.n4015 240.244
R5597 gnd.n4012 gnd.n4011 240.244
R5598 gnd.n3285 gnd.n2997 240.244
R5599 gnd.n3295 gnd.n2997 240.244
R5600 gnd.n3295 gnd.n2988 240.244
R5601 gnd.n2988 gnd.n2977 240.244
R5602 gnd.n3316 gnd.n2977 240.244
R5603 gnd.n3316 gnd.n2971 240.244
R5604 gnd.n3326 gnd.n2971 240.244
R5605 gnd.n3326 gnd.n2960 240.244
R5606 gnd.n2960 gnd.n2952 240.244
R5607 gnd.n3344 gnd.n2952 240.244
R5608 gnd.n3345 gnd.n3344 240.244
R5609 gnd.n3345 gnd.n2937 240.244
R5610 gnd.n3347 gnd.n2937 240.244
R5611 gnd.n3347 gnd.n2923 240.244
R5612 gnd.n3389 gnd.n2923 240.244
R5613 gnd.n3390 gnd.n3389 240.244
R5614 gnd.n3393 gnd.n3390 240.244
R5615 gnd.n3393 gnd.n2878 240.244
R5616 gnd.n2918 gnd.n2878 240.244
R5617 gnd.n2918 gnd.n2888 240.244
R5618 gnd.n3403 gnd.n2888 240.244
R5619 gnd.n3403 gnd.n2909 240.244
R5620 gnd.n3413 gnd.n2909 240.244
R5621 gnd.n3413 gnd.n2791 240.244
R5622 gnd.n3458 gnd.n2791 240.244
R5623 gnd.n3458 gnd.n2777 240.244
R5624 gnd.n3480 gnd.n2777 240.244
R5625 gnd.n3481 gnd.n3480 240.244
R5626 gnd.n3481 gnd.n2764 240.244
R5627 gnd.n2764 gnd.n2753 240.244
R5628 gnd.n3512 gnd.n2753 240.244
R5629 gnd.n3513 gnd.n3512 240.244
R5630 gnd.n3514 gnd.n3513 240.244
R5631 gnd.n3514 gnd.n2738 240.244
R5632 gnd.n2738 gnd.n2737 240.244
R5633 gnd.n2737 gnd.n2722 240.244
R5634 gnd.n3565 gnd.n2722 240.244
R5635 gnd.n3566 gnd.n3565 240.244
R5636 gnd.n3566 gnd.n2709 240.244
R5637 gnd.n2709 gnd.n2698 240.244
R5638 gnd.n3597 gnd.n2698 240.244
R5639 gnd.n3598 gnd.n3597 240.244
R5640 gnd.n3599 gnd.n3598 240.244
R5641 gnd.n3599 gnd.n2682 240.244
R5642 gnd.n2682 gnd.n2681 240.244
R5643 gnd.n2681 gnd.n2668 240.244
R5644 gnd.n3654 gnd.n2668 240.244
R5645 gnd.n3655 gnd.n3654 240.244
R5646 gnd.n3655 gnd.n2655 240.244
R5647 gnd.n2655 gnd.n2645 240.244
R5648 gnd.n3943 gnd.n2645 240.244
R5649 gnd.n3946 gnd.n3943 240.244
R5650 gnd.n3946 gnd.n3945 240.244
R5651 gnd.n3275 gnd.n3010 240.244
R5652 gnd.n3031 gnd.n3010 240.244
R5653 gnd.n3034 gnd.n3033 240.244
R5654 gnd.n3041 gnd.n3040 240.244
R5655 gnd.n3044 gnd.n3043 240.244
R5656 gnd.n3051 gnd.n3050 240.244
R5657 gnd.n3054 gnd.n3053 240.244
R5658 gnd.n3061 gnd.n3060 240.244
R5659 gnd.n3283 gnd.n3007 240.244
R5660 gnd.n3007 gnd.n2986 240.244
R5661 gnd.n3306 gnd.n2986 240.244
R5662 gnd.n3306 gnd.n2980 240.244
R5663 gnd.n3314 gnd.n2980 240.244
R5664 gnd.n3314 gnd.n2982 240.244
R5665 gnd.n2982 gnd.n2958 240.244
R5666 gnd.n3336 gnd.n2958 240.244
R5667 gnd.n3336 gnd.n2954 240.244
R5668 gnd.n3342 gnd.n2954 240.244
R5669 gnd.n3342 gnd.n2936 240.244
R5670 gnd.n3367 gnd.n2936 240.244
R5671 gnd.n3367 gnd.n2931 240.244
R5672 gnd.n3379 gnd.n2931 240.244
R5673 gnd.n3379 gnd.n2932 240.244
R5674 gnd.n3375 gnd.n2932 240.244
R5675 gnd.n3375 gnd.n2880 240.244
R5676 gnd.n3427 gnd.n2880 240.244
R5677 gnd.n3427 gnd.n2881 240.244
R5678 gnd.n3423 gnd.n2881 240.244
R5679 gnd.n3423 gnd.n2887 240.244
R5680 gnd.n2907 gnd.n2887 240.244
R5681 gnd.n2907 gnd.n2789 240.244
R5682 gnd.n3462 gnd.n2789 240.244
R5683 gnd.n3462 gnd.n2784 240.244
R5684 gnd.n3470 gnd.n2784 240.244
R5685 gnd.n3470 gnd.n2785 240.244
R5686 gnd.n2785 gnd.n2762 240.244
R5687 gnd.n3502 gnd.n2762 240.244
R5688 gnd.n3502 gnd.n2757 240.244
R5689 gnd.n3510 gnd.n2757 240.244
R5690 gnd.n3510 gnd.n2758 240.244
R5691 gnd.n2758 gnd.n2735 240.244
R5692 gnd.n3547 gnd.n2735 240.244
R5693 gnd.n3547 gnd.n2730 240.244
R5694 gnd.n3555 gnd.n2730 240.244
R5695 gnd.n3555 gnd.n2731 240.244
R5696 gnd.n2731 gnd.n2707 240.244
R5697 gnd.n3587 gnd.n2707 240.244
R5698 gnd.n3587 gnd.n2702 240.244
R5699 gnd.n3595 gnd.n2702 240.244
R5700 gnd.n3595 gnd.n2703 240.244
R5701 gnd.n2703 gnd.n2680 240.244
R5702 gnd.n3636 gnd.n2680 240.244
R5703 gnd.n3636 gnd.n2675 240.244
R5704 gnd.n3644 gnd.n2675 240.244
R5705 gnd.n3644 gnd.n2676 240.244
R5706 gnd.n2676 gnd.n2653 240.244
R5707 gnd.n3931 gnd.n2653 240.244
R5708 gnd.n3931 gnd.n2648 240.244
R5709 gnd.n3941 gnd.n2648 240.244
R5710 gnd.n3941 gnd.n2649 240.244
R5711 gnd.n2649 gnd.n2588 240.244
R5712 gnd.n319 gnd.n208 240.244
R5713 gnd.n7419 gnd.n7418 240.244
R5714 gnd.n7416 gnd.n323 240.244
R5715 gnd.n7412 gnd.n7411 240.244
R5716 gnd.n7409 gnd.n330 240.244
R5717 gnd.n7405 gnd.n7404 240.244
R5718 gnd.n7402 gnd.n337 240.244
R5719 gnd.n7398 gnd.n7397 240.244
R5720 gnd.n7395 gnd.n344 240.244
R5721 gnd.n5775 gnd.n1474 240.244
R5722 gnd.n5775 gnd.n1483 240.244
R5723 gnd.n5738 gnd.n1483 240.244
R5724 gnd.n5738 gnd.n1499 240.244
R5725 gnd.n5739 gnd.n1499 240.244
R5726 gnd.n5739 gnd.n1512 240.244
R5727 gnd.n5742 gnd.n1512 240.244
R5728 gnd.n5742 gnd.n1522 240.244
R5729 gnd.n5760 gnd.n1522 240.244
R5730 gnd.n5760 gnd.n1532 240.244
R5731 gnd.n5823 gnd.n1532 240.244
R5732 gnd.n5823 gnd.n1542 240.244
R5733 gnd.n5829 gnd.n1542 240.244
R5734 gnd.n5829 gnd.n1552 240.244
R5735 gnd.n5838 gnd.n1552 240.244
R5736 gnd.n5838 gnd.n1562 240.244
R5737 gnd.n5844 gnd.n1562 240.244
R5738 gnd.n5844 gnd.n1572 240.244
R5739 gnd.n5874 gnd.n1572 240.244
R5740 gnd.n5874 gnd.n1582 240.244
R5741 gnd.n5860 gnd.n1582 240.244
R5742 gnd.n5860 gnd.n1592 240.244
R5743 gnd.n1596 gnd.n1592 240.244
R5744 gnd.n5861 gnd.n1596 240.244
R5745 gnd.n5861 gnd.n383 240.244
R5746 gnd.n7282 gnd.n383 240.244
R5747 gnd.n7282 gnd.n86 240.244
R5748 gnd.n7612 gnd.n86 240.244
R5749 gnd.n7612 gnd.n88 240.244
R5750 gnd.n7346 gnd.n88 240.244
R5751 gnd.n7346 gnd.n106 240.244
R5752 gnd.n7352 gnd.n106 240.244
R5753 gnd.n7352 gnd.n117 240.244
R5754 gnd.n365 gnd.n117 240.244
R5755 gnd.n365 gnd.n126 240.244
R5756 gnd.n7359 gnd.n126 240.244
R5757 gnd.n7359 gnd.n135 240.244
R5758 gnd.n362 gnd.n135 240.244
R5759 gnd.n362 gnd.n145 240.244
R5760 gnd.n7366 gnd.n145 240.244
R5761 gnd.n7366 gnd.n154 240.244
R5762 gnd.n359 gnd.n154 240.244
R5763 gnd.n359 gnd.n164 240.244
R5764 gnd.n7373 gnd.n164 240.244
R5765 gnd.n7373 gnd.n173 240.244
R5766 gnd.n356 gnd.n173 240.244
R5767 gnd.n356 gnd.n183 240.244
R5768 gnd.n7380 gnd.n183 240.244
R5769 gnd.n7380 gnd.n193 240.244
R5770 gnd.n353 gnd.n193 240.244
R5771 gnd.n353 gnd.n203 240.244
R5772 gnd.n7387 gnd.n203 240.244
R5773 gnd.n7387 gnd.n211 240.244
R5774 gnd.n1318 gnd.n1317 240.244
R5775 gnd.n1393 gnd.n1325 240.244
R5776 gnd.n1396 gnd.n1326 240.244
R5777 gnd.n1334 gnd.n1333 240.244
R5778 gnd.n1398 gnd.n1341 240.244
R5779 gnd.n1401 gnd.n1342 240.244
R5780 gnd.n1350 gnd.n1349 240.244
R5781 gnd.n1403 gnd.n1359 240.244
R5782 gnd.n6083 gnd.n1362 240.244
R5783 gnd.n5959 gnd.n1477 240.244
R5784 gnd.n1485 gnd.n1477 240.244
R5785 gnd.n1501 gnd.n1485 240.244
R5786 gnd.n5945 gnd.n1501 240.244
R5787 gnd.n5945 gnd.n1502 240.244
R5788 gnd.n5941 gnd.n1502 240.244
R5789 gnd.n5941 gnd.n1509 240.244
R5790 gnd.n5933 gnd.n1509 240.244
R5791 gnd.n5933 gnd.n1524 240.244
R5792 gnd.n5929 gnd.n1524 240.244
R5793 gnd.n5929 gnd.n1529 240.244
R5794 gnd.n5921 gnd.n1529 240.244
R5795 gnd.n5921 gnd.n1544 240.244
R5796 gnd.n5917 gnd.n1544 240.244
R5797 gnd.n5917 gnd.n1549 240.244
R5798 gnd.n5909 gnd.n1549 240.244
R5799 gnd.n5909 gnd.n1564 240.244
R5800 gnd.n5905 gnd.n1564 240.244
R5801 gnd.n5905 gnd.n1569 240.244
R5802 gnd.n5897 gnd.n1569 240.244
R5803 gnd.n5897 gnd.n1584 240.244
R5804 gnd.n5893 gnd.n1584 240.244
R5805 gnd.n5893 gnd.n1589 240.244
R5806 gnd.n1589 gnd.n380 240.244
R5807 gnd.n7288 gnd.n380 240.244
R5808 gnd.n7288 gnd.n374 240.244
R5809 gnd.n7297 gnd.n374 240.244
R5810 gnd.n7297 gnd.n91 240.244
R5811 gnd.n7300 gnd.n91 240.244
R5812 gnd.n7300 gnd.n108 240.244
R5813 gnd.n7602 gnd.n108 240.244
R5814 gnd.n7602 gnd.n109 240.244
R5815 gnd.n7598 gnd.n109 240.244
R5816 gnd.n7598 gnd.n115 240.244
R5817 gnd.n7590 gnd.n115 240.244
R5818 gnd.n7590 gnd.n127 240.244
R5819 gnd.n7586 gnd.n127 240.244
R5820 gnd.n7586 gnd.n132 240.244
R5821 gnd.n7578 gnd.n132 240.244
R5822 gnd.n7578 gnd.n147 240.244
R5823 gnd.n7574 gnd.n147 240.244
R5824 gnd.n7574 gnd.n152 240.244
R5825 gnd.n7566 gnd.n152 240.244
R5826 gnd.n7566 gnd.n165 240.244
R5827 gnd.n7562 gnd.n165 240.244
R5828 gnd.n7562 gnd.n170 240.244
R5829 gnd.n7554 gnd.n170 240.244
R5830 gnd.n7554 gnd.n185 240.244
R5831 gnd.n7550 gnd.n185 240.244
R5832 gnd.n7550 gnd.n190 240.244
R5833 gnd.n7542 gnd.n190 240.244
R5834 gnd.n7542 gnd.n204 240.244
R5835 gnd.n7538 gnd.n204 240.244
R5836 gnd.n2608 gnd.n2566 240.244
R5837 gnd.n4002 gnd.n4001 240.244
R5838 gnd.n3998 gnd.n3997 240.244
R5839 gnd.n3994 gnd.n3993 240.244
R5840 gnd.n3990 gnd.n3989 240.244
R5841 gnd.n3986 gnd.n3985 240.244
R5842 gnd.n3982 gnd.n3981 240.244
R5843 gnd.n3978 gnd.n3977 240.244
R5844 gnd.n3974 gnd.n3973 240.244
R5845 gnd.n3970 gnd.n3969 240.244
R5846 gnd.n3966 gnd.n3965 240.244
R5847 gnd.n3962 gnd.n3961 240.244
R5848 gnd.n3958 gnd.n3957 240.244
R5849 gnd.n3198 gnd.n3095 240.244
R5850 gnd.n3198 gnd.n3088 240.244
R5851 gnd.n3209 gnd.n3088 240.244
R5852 gnd.n3209 gnd.n3084 240.244
R5853 gnd.n3215 gnd.n3084 240.244
R5854 gnd.n3215 gnd.n3076 240.244
R5855 gnd.n3225 gnd.n3076 240.244
R5856 gnd.n3225 gnd.n3071 240.244
R5857 gnd.n3261 gnd.n3071 240.244
R5858 gnd.n3261 gnd.n3072 240.244
R5859 gnd.n3072 gnd.n3019 240.244
R5860 gnd.n3256 gnd.n3019 240.244
R5861 gnd.n3256 gnd.n3255 240.244
R5862 gnd.n3255 gnd.n2998 240.244
R5863 gnd.n3251 gnd.n2998 240.244
R5864 gnd.n3251 gnd.n2989 240.244
R5865 gnd.n3248 gnd.n2989 240.244
R5866 gnd.n3248 gnd.n3247 240.244
R5867 gnd.n3247 gnd.n2972 240.244
R5868 gnd.n3243 gnd.n2972 240.244
R5869 gnd.n3243 gnd.n2961 240.244
R5870 gnd.n2961 gnd.n2942 240.244
R5871 gnd.n3356 gnd.n2942 240.244
R5872 gnd.n3356 gnd.n2938 240.244
R5873 gnd.n3364 gnd.n2938 240.244
R5874 gnd.n3364 gnd.n2929 240.244
R5875 gnd.n2929 gnd.n2865 240.244
R5876 gnd.n3436 gnd.n2865 240.244
R5877 gnd.n3436 gnd.n2866 240.244
R5878 gnd.n2877 gnd.n2866 240.244
R5879 gnd.n2912 gnd.n2877 240.244
R5880 gnd.n2915 gnd.n2912 240.244
R5881 gnd.n2915 gnd.n2889 240.244
R5882 gnd.n2902 gnd.n2889 240.244
R5883 gnd.n2902 gnd.n2899 240.244
R5884 gnd.n2899 gnd.n2792 240.244
R5885 gnd.n3457 gnd.n2792 240.244
R5886 gnd.n3457 gnd.n2782 240.244
R5887 gnd.n3453 gnd.n2782 240.244
R5888 gnd.n3453 gnd.n2776 240.244
R5889 gnd.n3450 gnd.n2776 240.244
R5890 gnd.n3450 gnd.n2765 240.244
R5891 gnd.n3447 gnd.n2765 240.244
R5892 gnd.n3447 gnd.n2743 240.244
R5893 gnd.n3523 gnd.n2743 240.244
R5894 gnd.n3523 gnd.n2739 240.244
R5895 gnd.n3544 gnd.n2739 240.244
R5896 gnd.n3544 gnd.n2728 240.244
R5897 gnd.n3540 gnd.n2728 240.244
R5898 gnd.n3540 gnd.n2721 240.244
R5899 gnd.n3537 gnd.n2721 240.244
R5900 gnd.n3537 gnd.n2710 240.244
R5901 gnd.n3534 gnd.n2710 240.244
R5902 gnd.n3534 gnd.n2687 240.244
R5903 gnd.n3608 gnd.n2687 240.244
R5904 gnd.n3608 gnd.n2683 240.244
R5905 gnd.n3633 gnd.n2683 240.244
R5906 gnd.n3633 gnd.n2674 240.244
R5907 gnd.n3629 gnd.n2674 240.244
R5908 gnd.n3629 gnd.n2667 240.244
R5909 gnd.n3625 gnd.n2667 240.244
R5910 gnd.n3625 gnd.n2656 240.244
R5911 gnd.n3622 gnd.n2656 240.244
R5912 gnd.n3622 gnd.n2637 240.244
R5913 gnd.n3953 gnd.n2637 240.244
R5914 gnd.n3112 gnd.n3111 240.244
R5915 gnd.n3183 gnd.n3111 240.244
R5916 gnd.n3181 gnd.n3180 240.244
R5917 gnd.n3177 gnd.n3176 240.244
R5918 gnd.n3173 gnd.n3172 240.244
R5919 gnd.n3169 gnd.n3168 240.244
R5920 gnd.n3165 gnd.n3164 240.244
R5921 gnd.n3161 gnd.n3160 240.244
R5922 gnd.n3157 gnd.n3156 240.244
R5923 gnd.n3153 gnd.n3152 240.244
R5924 gnd.n3149 gnd.n3148 240.244
R5925 gnd.n3145 gnd.n3144 240.244
R5926 gnd.n3141 gnd.n3099 240.244
R5927 gnd.n3201 gnd.n3093 240.244
R5928 gnd.n3201 gnd.n3089 240.244
R5929 gnd.n3207 gnd.n3089 240.244
R5930 gnd.n3207 gnd.n3082 240.244
R5931 gnd.n3217 gnd.n3082 240.244
R5932 gnd.n3217 gnd.n3078 240.244
R5933 gnd.n3223 gnd.n3078 240.244
R5934 gnd.n3223 gnd.n3069 240.244
R5935 gnd.n3263 gnd.n3069 240.244
R5936 gnd.n3263 gnd.n3020 240.244
R5937 gnd.n3271 gnd.n3020 240.244
R5938 gnd.n3271 gnd.n3021 240.244
R5939 gnd.n3021 gnd.n2999 240.244
R5940 gnd.n3292 gnd.n2999 240.244
R5941 gnd.n3292 gnd.n2991 240.244
R5942 gnd.n3303 gnd.n2991 240.244
R5943 gnd.n3303 gnd.n2992 240.244
R5944 gnd.n2992 gnd.n2973 240.244
R5945 gnd.n3323 gnd.n2973 240.244
R5946 gnd.n3323 gnd.n2963 240.244
R5947 gnd.n3333 gnd.n2963 240.244
R5948 gnd.n3333 gnd.n2944 240.244
R5949 gnd.n3354 gnd.n2944 240.244
R5950 gnd.n3354 gnd.n2946 240.244
R5951 gnd.n2946 gnd.n2927 240.244
R5952 gnd.n3382 gnd.n2927 240.244
R5953 gnd.n3382 gnd.n2869 240.244
R5954 gnd.n3434 gnd.n2869 240.244
R5955 gnd.n3434 gnd.n2870 240.244
R5956 gnd.n3430 gnd.n2870 240.244
R5957 gnd.n3430 gnd.n2876 240.244
R5958 gnd.n2891 gnd.n2876 240.244
R5959 gnd.n3420 gnd.n2891 240.244
R5960 gnd.n3420 gnd.n2892 240.244
R5961 gnd.n3416 gnd.n2892 240.244
R5962 gnd.n3416 gnd.n2898 240.244
R5963 gnd.n2898 gnd.n2781 240.244
R5964 gnd.n3473 gnd.n2781 240.244
R5965 gnd.n3473 gnd.n2774 240.244
R5966 gnd.n3484 gnd.n2774 240.244
R5967 gnd.n3484 gnd.n2767 240.244
R5968 gnd.n3499 gnd.n2767 240.244
R5969 gnd.n3499 gnd.n2768 240.244
R5970 gnd.n2768 gnd.n2746 240.244
R5971 gnd.n3521 gnd.n2746 240.244
R5972 gnd.n3521 gnd.n2747 240.244
R5973 gnd.n2747 gnd.n2726 240.244
R5974 gnd.n3558 gnd.n2726 240.244
R5975 gnd.n3558 gnd.n2719 240.244
R5976 gnd.n3569 gnd.n2719 240.244
R5977 gnd.n3569 gnd.n2712 240.244
R5978 gnd.n3584 gnd.n2712 240.244
R5979 gnd.n3584 gnd.n2713 240.244
R5980 gnd.n2713 gnd.n2690 240.244
R5981 gnd.n3606 gnd.n2690 240.244
R5982 gnd.n3606 gnd.n2692 240.244
R5983 gnd.n2692 gnd.n2672 240.244
R5984 gnd.n3647 gnd.n2672 240.244
R5985 gnd.n3647 gnd.n2665 240.244
R5986 gnd.n3659 gnd.n2665 240.244
R5987 gnd.n3659 gnd.n2658 240.244
R5988 gnd.n3928 gnd.n2658 240.244
R5989 gnd.n3928 gnd.n2659 240.244
R5990 gnd.n2659 gnd.n2640 240.244
R5991 gnd.n3951 gnd.n2640 240.244
R5992 gnd.n2315 gnd.n1064 240.244
R5993 gnd.n2326 gnd.n2317 240.244
R5994 gnd.n2329 gnd.n2328 240.244
R5995 gnd.n2338 gnd.n2337 240.244
R5996 gnd.n2349 gnd.n2340 240.244
R5997 gnd.n2352 gnd.n2351 240.244
R5998 gnd.n2361 gnd.n2360 240.244
R5999 gnd.n2373 gnd.n2363 240.244
R6000 gnd.n2379 gnd.n2375 240.244
R6001 gnd.n4197 gnd.n2554 240.244
R6002 gnd.n4194 gnd.n2554 240.244
R6003 gnd.n4194 gnd.n2545 240.244
R6004 gnd.n4191 gnd.n2545 240.244
R6005 gnd.n4191 gnd.n2535 240.244
R6006 gnd.n4188 gnd.n2535 240.244
R6007 gnd.n4188 gnd.n2526 240.244
R6008 gnd.n4185 gnd.n2526 240.244
R6009 gnd.n4185 gnd.n2518 240.244
R6010 gnd.n4182 gnd.n2518 240.244
R6011 gnd.n4182 gnd.n2509 240.244
R6012 gnd.n4179 gnd.n2509 240.244
R6013 gnd.n4179 gnd.n2498 240.244
R6014 gnd.n2498 gnd.n2487 240.244
R6015 gnd.n4442 gnd.n2487 240.244
R6016 gnd.n4442 gnd.n2483 240.244
R6017 gnd.n4460 gnd.n2483 240.244
R6018 gnd.n4460 gnd.n2473 240.244
R6019 gnd.n4456 gnd.n2473 240.244
R6020 gnd.n4456 gnd.n2465 240.244
R6021 gnd.n4453 gnd.n2465 240.244
R6022 gnd.n4453 gnd.n2451 240.244
R6023 gnd.n4502 gnd.n2451 240.244
R6024 gnd.n4503 gnd.n4502 240.244
R6025 gnd.n4503 gnd.n940 240.244
R6026 gnd.n4515 gnd.n940 240.244
R6027 gnd.n4515 gnd.n2438 240.244
R6028 gnd.n4508 gnd.n2438 240.244
R6029 gnd.n4508 gnd.n2421 240.244
R6030 gnd.n4566 gnd.n2421 240.244
R6031 gnd.n4566 gnd.n957 240.244
R6032 gnd.n4572 gnd.n957 240.244
R6033 gnd.n4572 gnd.n969 240.244
R6034 gnd.n4581 gnd.n969 240.244
R6035 gnd.n4581 gnd.n978 240.244
R6036 gnd.n4587 gnd.n978 240.244
R6037 gnd.n4587 gnd.n988 240.244
R6038 gnd.n4623 gnd.n988 240.244
R6039 gnd.n4623 gnd.n998 240.244
R6040 gnd.n2408 gnd.n998 240.244
R6041 gnd.n2408 gnd.n1008 240.244
R6042 gnd.n2409 gnd.n1008 240.244
R6043 gnd.n2409 gnd.n1018 240.244
R6044 gnd.n4608 gnd.n1018 240.244
R6045 gnd.n4608 gnd.n1028 240.244
R6046 gnd.n2391 gnd.n1028 240.244
R6047 gnd.n2391 gnd.n1038 240.244
R6048 gnd.n4679 gnd.n1038 240.244
R6049 gnd.n4679 gnd.n1048 240.244
R6050 gnd.n4686 gnd.n1048 240.244
R6051 gnd.n4686 gnd.n1059 240.244
R6052 gnd.n4695 gnd.n1059 240.244
R6053 gnd.n4695 gnd.n1067 240.244
R6054 gnd.n4234 gnd.n4233 240.244
R6055 gnd.n4230 gnd.n4229 240.244
R6056 gnd.n4226 gnd.n4225 240.244
R6057 gnd.n4222 gnd.n4221 240.244
R6058 gnd.n4218 gnd.n4217 240.244
R6059 gnd.n4214 gnd.n4213 240.244
R6060 gnd.n4210 gnd.n4209 240.244
R6061 gnd.n4206 gnd.n4205 240.244
R6062 gnd.n4161 gnd.n4080 240.244
R6063 gnd.n4366 gnd.n2555 240.244
R6064 gnd.n4366 gnd.n2556 240.244
R6065 gnd.n2556 gnd.n2546 240.244
R6066 gnd.n2546 gnd.n2537 240.244
R6067 gnd.n4386 gnd.n2537 240.244
R6068 gnd.n4386 gnd.n2538 240.244
R6069 gnd.n2538 gnd.n2527 240.244
R6070 gnd.n2527 gnd.n2519 240.244
R6071 gnd.n4406 gnd.n2519 240.244
R6072 gnd.n4406 gnd.n2520 240.244
R6073 gnd.n2520 gnd.n2510 240.244
R6074 gnd.n2510 gnd.n2500 240.244
R6075 gnd.n4430 gnd.n2500 240.244
R6076 gnd.n4430 gnd.n2501 240.244
R6077 gnd.n2501 gnd.n2489 240.244
R6078 gnd.n4425 gnd.n2489 240.244
R6079 gnd.n4425 gnd.n2475 240.244
R6080 gnd.n4471 gnd.n2475 240.244
R6081 gnd.n4471 gnd.n2476 240.244
R6082 gnd.n2476 gnd.n2466 240.244
R6083 gnd.n2466 gnd.n2458 240.244
R6084 gnd.n4496 gnd.n2458 240.244
R6085 gnd.n4496 gnd.n2453 240.244
R6086 gnd.n4492 gnd.n2453 240.244
R6087 gnd.n4492 gnd.n941 240.244
R6088 gnd.n2440 gnd.n941 240.244
R6089 gnd.n4528 gnd.n2440 240.244
R6090 gnd.n4528 gnd.n2441 240.244
R6091 gnd.n2441 gnd.n2434 240.244
R6092 gnd.n2434 gnd.n959 240.244
R6093 gnd.n6463 gnd.n959 240.244
R6094 gnd.n6463 gnd.n960 240.244
R6095 gnd.n6459 gnd.n960 240.244
R6096 gnd.n6459 gnd.n966 240.244
R6097 gnd.n6451 gnd.n966 240.244
R6098 gnd.n6451 gnd.n980 240.244
R6099 gnd.n6447 gnd.n980 240.244
R6100 gnd.n6447 gnd.n985 240.244
R6101 gnd.n6439 gnd.n985 240.244
R6102 gnd.n6439 gnd.n1000 240.244
R6103 gnd.n6435 gnd.n1000 240.244
R6104 gnd.n6435 gnd.n1005 240.244
R6105 gnd.n6427 gnd.n1005 240.244
R6106 gnd.n6427 gnd.n1020 240.244
R6107 gnd.n6423 gnd.n1020 240.244
R6108 gnd.n6423 gnd.n1025 240.244
R6109 gnd.n6415 gnd.n1025 240.244
R6110 gnd.n6415 gnd.n1040 240.244
R6111 gnd.n6411 gnd.n1040 240.244
R6112 gnd.n6411 gnd.n1045 240.244
R6113 gnd.n6403 gnd.n1045 240.244
R6114 gnd.n6403 gnd.n1060 240.244
R6115 gnd.n6399 gnd.n1060 240.244
R6116 gnd.n6647 gnd.n767 240.244
R6117 gnd.n6647 gnd.n765 240.244
R6118 gnd.n6651 gnd.n765 240.244
R6119 gnd.n6651 gnd.n761 240.244
R6120 gnd.n6657 gnd.n761 240.244
R6121 gnd.n6657 gnd.n759 240.244
R6122 gnd.n6661 gnd.n759 240.244
R6123 gnd.n6661 gnd.n755 240.244
R6124 gnd.n6667 gnd.n755 240.244
R6125 gnd.n6667 gnd.n753 240.244
R6126 gnd.n6671 gnd.n753 240.244
R6127 gnd.n6671 gnd.n749 240.244
R6128 gnd.n6677 gnd.n749 240.244
R6129 gnd.n6677 gnd.n747 240.244
R6130 gnd.n6681 gnd.n747 240.244
R6131 gnd.n6681 gnd.n743 240.244
R6132 gnd.n6687 gnd.n743 240.244
R6133 gnd.n6687 gnd.n741 240.244
R6134 gnd.n6691 gnd.n741 240.244
R6135 gnd.n6691 gnd.n737 240.244
R6136 gnd.n6697 gnd.n737 240.244
R6137 gnd.n6697 gnd.n735 240.244
R6138 gnd.n6701 gnd.n735 240.244
R6139 gnd.n6701 gnd.n731 240.244
R6140 gnd.n6707 gnd.n731 240.244
R6141 gnd.n6707 gnd.n729 240.244
R6142 gnd.n6711 gnd.n729 240.244
R6143 gnd.n6711 gnd.n725 240.244
R6144 gnd.n6717 gnd.n725 240.244
R6145 gnd.n6717 gnd.n723 240.244
R6146 gnd.n6721 gnd.n723 240.244
R6147 gnd.n6721 gnd.n719 240.244
R6148 gnd.n6727 gnd.n719 240.244
R6149 gnd.n6727 gnd.n717 240.244
R6150 gnd.n6731 gnd.n717 240.244
R6151 gnd.n6731 gnd.n713 240.244
R6152 gnd.n6737 gnd.n713 240.244
R6153 gnd.n6737 gnd.n711 240.244
R6154 gnd.n6741 gnd.n711 240.244
R6155 gnd.n6741 gnd.n707 240.244
R6156 gnd.n6747 gnd.n707 240.244
R6157 gnd.n6747 gnd.n705 240.244
R6158 gnd.n6751 gnd.n705 240.244
R6159 gnd.n6751 gnd.n701 240.244
R6160 gnd.n6757 gnd.n701 240.244
R6161 gnd.n6757 gnd.n699 240.244
R6162 gnd.n6761 gnd.n699 240.244
R6163 gnd.n6761 gnd.n695 240.244
R6164 gnd.n6767 gnd.n695 240.244
R6165 gnd.n6767 gnd.n693 240.244
R6166 gnd.n6771 gnd.n693 240.244
R6167 gnd.n6771 gnd.n689 240.244
R6168 gnd.n6777 gnd.n689 240.244
R6169 gnd.n6777 gnd.n687 240.244
R6170 gnd.n6781 gnd.n687 240.244
R6171 gnd.n6781 gnd.n683 240.244
R6172 gnd.n6787 gnd.n683 240.244
R6173 gnd.n6787 gnd.n681 240.244
R6174 gnd.n6791 gnd.n681 240.244
R6175 gnd.n6791 gnd.n677 240.244
R6176 gnd.n6797 gnd.n677 240.244
R6177 gnd.n6797 gnd.n675 240.244
R6178 gnd.n6801 gnd.n675 240.244
R6179 gnd.n6801 gnd.n671 240.244
R6180 gnd.n6807 gnd.n671 240.244
R6181 gnd.n6807 gnd.n669 240.244
R6182 gnd.n6811 gnd.n669 240.244
R6183 gnd.n6811 gnd.n665 240.244
R6184 gnd.n6817 gnd.n665 240.244
R6185 gnd.n6817 gnd.n663 240.244
R6186 gnd.n6821 gnd.n663 240.244
R6187 gnd.n6821 gnd.n659 240.244
R6188 gnd.n6827 gnd.n659 240.244
R6189 gnd.n6827 gnd.n657 240.244
R6190 gnd.n6831 gnd.n657 240.244
R6191 gnd.n6831 gnd.n653 240.244
R6192 gnd.n6837 gnd.n653 240.244
R6193 gnd.n6837 gnd.n651 240.244
R6194 gnd.n6841 gnd.n651 240.244
R6195 gnd.n6841 gnd.n647 240.244
R6196 gnd.n6847 gnd.n647 240.244
R6197 gnd.n6847 gnd.n645 240.244
R6198 gnd.n6851 gnd.n645 240.244
R6199 gnd.n6851 gnd.n641 240.244
R6200 gnd.n6857 gnd.n641 240.244
R6201 gnd.n6857 gnd.n639 240.244
R6202 gnd.n6861 gnd.n639 240.244
R6203 gnd.n6861 gnd.n635 240.244
R6204 gnd.n6867 gnd.n635 240.244
R6205 gnd.n6867 gnd.n633 240.244
R6206 gnd.n6871 gnd.n633 240.244
R6207 gnd.n6871 gnd.n629 240.244
R6208 gnd.n6877 gnd.n629 240.244
R6209 gnd.n6877 gnd.n627 240.244
R6210 gnd.n6881 gnd.n627 240.244
R6211 gnd.n6881 gnd.n623 240.244
R6212 gnd.n6887 gnd.n623 240.244
R6213 gnd.n6887 gnd.n621 240.244
R6214 gnd.n6891 gnd.n621 240.244
R6215 gnd.n6891 gnd.n617 240.244
R6216 gnd.n6897 gnd.n617 240.244
R6217 gnd.n6897 gnd.n615 240.244
R6218 gnd.n6901 gnd.n615 240.244
R6219 gnd.n6901 gnd.n611 240.244
R6220 gnd.n6907 gnd.n611 240.244
R6221 gnd.n6907 gnd.n609 240.244
R6222 gnd.n6911 gnd.n609 240.244
R6223 gnd.n6911 gnd.n605 240.244
R6224 gnd.n6917 gnd.n605 240.244
R6225 gnd.n6917 gnd.n603 240.244
R6226 gnd.n6921 gnd.n603 240.244
R6227 gnd.n6921 gnd.n599 240.244
R6228 gnd.n6927 gnd.n599 240.244
R6229 gnd.n6927 gnd.n597 240.244
R6230 gnd.n6931 gnd.n597 240.244
R6231 gnd.n6931 gnd.n593 240.244
R6232 gnd.n6937 gnd.n593 240.244
R6233 gnd.n6937 gnd.n591 240.244
R6234 gnd.n6941 gnd.n591 240.244
R6235 gnd.n6941 gnd.n587 240.244
R6236 gnd.n6947 gnd.n587 240.244
R6237 gnd.n6947 gnd.n585 240.244
R6238 gnd.n6951 gnd.n585 240.244
R6239 gnd.n6951 gnd.n581 240.244
R6240 gnd.n6957 gnd.n581 240.244
R6241 gnd.n6957 gnd.n579 240.244
R6242 gnd.n6961 gnd.n579 240.244
R6243 gnd.n6961 gnd.n575 240.244
R6244 gnd.n6967 gnd.n575 240.244
R6245 gnd.n6967 gnd.n573 240.244
R6246 gnd.n6971 gnd.n573 240.244
R6247 gnd.n6971 gnd.n569 240.244
R6248 gnd.n6977 gnd.n569 240.244
R6249 gnd.n6977 gnd.n567 240.244
R6250 gnd.n6981 gnd.n567 240.244
R6251 gnd.n6981 gnd.n563 240.244
R6252 gnd.n6987 gnd.n563 240.244
R6253 gnd.n6987 gnd.n561 240.244
R6254 gnd.n6991 gnd.n561 240.244
R6255 gnd.n6991 gnd.n557 240.244
R6256 gnd.n6997 gnd.n557 240.244
R6257 gnd.n6997 gnd.n555 240.244
R6258 gnd.n7001 gnd.n555 240.244
R6259 gnd.n7001 gnd.n551 240.244
R6260 gnd.n7007 gnd.n551 240.244
R6261 gnd.n7007 gnd.n549 240.244
R6262 gnd.n7011 gnd.n549 240.244
R6263 gnd.n7011 gnd.n545 240.244
R6264 gnd.n7017 gnd.n545 240.244
R6265 gnd.n7017 gnd.n543 240.244
R6266 gnd.n7021 gnd.n543 240.244
R6267 gnd.n7021 gnd.n539 240.244
R6268 gnd.n7027 gnd.n539 240.244
R6269 gnd.n7027 gnd.n537 240.244
R6270 gnd.n7031 gnd.n537 240.244
R6271 gnd.n7031 gnd.n533 240.244
R6272 gnd.n7037 gnd.n533 240.244
R6273 gnd.n7037 gnd.n531 240.244
R6274 gnd.n7041 gnd.n531 240.244
R6275 gnd.n7041 gnd.n527 240.244
R6276 gnd.n7047 gnd.n527 240.244
R6277 gnd.n7047 gnd.n525 240.244
R6278 gnd.n7051 gnd.n525 240.244
R6279 gnd.n7051 gnd.n521 240.244
R6280 gnd.n7057 gnd.n521 240.244
R6281 gnd.n7057 gnd.n519 240.244
R6282 gnd.n7061 gnd.n519 240.244
R6283 gnd.n7067 gnd.n515 240.244
R6284 gnd.n7067 gnd.n513 240.244
R6285 gnd.n7071 gnd.n513 240.244
R6286 gnd.n7071 gnd.n509 240.244
R6287 gnd.n7077 gnd.n509 240.244
R6288 gnd.n7077 gnd.n507 240.244
R6289 gnd.n7081 gnd.n507 240.244
R6290 gnd.n7081 gnd.n503 240.244
R6291 gnd.n7087 gnd.n503 240.244
R6292 gnd.n7087 gnd.n501 240.244
R6293 gnd.n7091 gnd.n501 240.244
R6294 gnd.n7091 gnd.n497 240.244
R6295 gnd.n7097 gnd.n497 240.244
R6296 gnd.n7097 gnd.n495 240.244
R6297 gnd.n7101 gnd.n495 240.244
R6298 gnd.n7101 gnd.n491 240.244
R6299 gnd.n7107 gnd.n491 240.244
R6300 gnd.n7107 gnd.n489 240.244
R6301 gnd.n7111 gnd.n489 240.244
R6302 gnd.n7111 gnd.n485 240.244
R6303 gnd.n7117 gnd.n485 240.244
R6304 gnd.n7117 gnd.n483 240.244
R6305 gnd.n7121 gnd.n483 240.244
R6306 gnd.n7121 gnd.n479 240.244
R6307 gnd.n7127 gnd.n479 240.244
R6308 gnd.n7127 gnd.n477 240.244
R6309 gnd.n7131 gnd.n477 240.244
R6310 gnd.n7131 gnd.n473 240.244
R6311 gnd.n7137 gnd.n473 240.244
R6312 gnd.n7137 gnd.n471 240.244
R6313 gnd.n7141 gnd.n471 240.244
R6314 gnd.n7141 gnd.n467 240.244
R6315 gnd.n7147 gnd.n467 240.244
R6316 gnd.n7147 gnd.n465 240.244
R6317 gnd.n7151 gnd.n465 240.244
R6318 gnd.n7151 gnd.n461 240.244
R6319 gnd.n7157 gnd.n461 240.244
R6320 gnd.n7157 gnd.n459 240.244
R6321 gnd.n7161 gnd.n459 240.244
R6322 gnd.n7161 gnd.n455 240.244
R6323 gnd.n7167 gnd.n455 240.244
R6324 gnd.n7167 gnd.n453 240.244
R6325 gnd.n7171 gnd.n453 240.244
R6326 gnd.n7171 gnd.n449 240.244
R6327 gnd.n7177 gnd.n449 240.244
R6328 gnd.n7177 gnd.n447 240.244
R6329 gnd.n7181 gnd.n447 240.244
R6330 gnd.n7181 gnd.n443 240.244
R6331 gnd.n7187 gnd.n443 240.244
R6332 gnd.n7187 gnd.n441 240.244
R6333 gnd.n7191 gnd.n441 240.244
R6334 gnd.n7191 gnd.n437 240.244
R6335 gnd.n7197 gnd.n437 240.244
R6336 gnd.n7197 gnd.n435 240.244
R6337 gnd.n7201 gnd.n435 240.244
R6338 gnd.n7201 gnd.n431 240.244
R6339 gnd.n7207 gnd.n431 240.244
R6340 gnd.n7207 gnd.n429 240.244
R6341 gnd.n7211 gnd.n429 240.244
R6342 gnd.n7211 gnd.n425 240.244
R6343 gnd.n7217 gnd.n425 240.244
R6344 gnd.n7217 gnd.n423 240.244
R6345 gnd.n7221 gnd.n423 240.244
R6346 gnd.n7221 gnd.n419 240.244
R6347 gnd.n7227 gnd.n419 240.244
R6348 gnd.n7227 gnd.n417 240.244
R6349 gnd.n7231 gnd.n417 240.244
R6350 gnd.n7231 gnd.n413 240.244
R6351 gnd.n7237 gnd.n413 240.244
R6352 gnd.n7237 gnd.n411 240.244
R6353 gnd.n7241 gnd.n411 240.244
R6354 gnd.n7241 gnd.n407 240.244
R6355 gnd.n7247 gnd.n407 240.244
R6356 gnd.n7247 gnd.n405 240.244
R6357 gnd.n7251 gnd.n405 240.244
R6358 gnd.n7251 gnd.n401 240.244
R6359 gnd.n7257 gnd.n401 240.244
R6360 gnd.n7257 gnd.n399 240.244
R6361 gnd.n7261 gnd.n399 240.244
R6362 gnd.n7261 gnd.n395 240.244
R6363 gnd.n7269 gnd.n395 240.244
R6364 gnd.n7269 gnd.n393 240.244
R6365 gnd.n7273 gnd.n393 240.244
R6366 gnd.n7274 gnd.n7273 240.244
R6367 gnd.n2431 gnd.n937 240.244
R6368 gnd.n4537 gnd.n2431 240.244
R6369 gnd.n4537 gnd.n2424 240.244
R6370 gnd.n4563 gnd.n2424 240.244
R6371 gnd.n4563 gnd.n2425 240.244
R6372 gnd.n4559 gnd.n2425 240.244
R6373 gnd.n4559 gnd.n4558 240.244
R6374 gnd.n4558 gnd.n4557 240.244
R6375 gnd.n4557 gnd.n4545 240.244
R6376 gnd.n4553 gnd.n4545 240.244
R6377 gnd.n4553 gnd.n2401 240.244
R6378 gnd.n4626 gnd.n2401 240.244
R6379 gnd.n4627 gnd.n4626 240.244
R6380 gnd.n4628 gnd.n4627 240.244
R6381 gnd.n4628 gnd.n2397 240.244
R6382 gnd.n4634 gnd.n2397 240.244
R6383 gnd.n4635 gnd.n4634 240.244
R6384 gnd.n4636 gnd.n4635 240.244
R6385 gnd.n4636 gnd.n2392 240.244
R6386 gnd.n4670 gnd.n2392 240.244
R6387 gnd.n4670 gnd.n2393 240.244
R6388 gnd.n4666 gnd.n2393 240.244
R6389 gnd.n4666 gnd.n4665 240.244
R6390 gnd.n4665 gnd.n4664 240.244
R6391 gnd.n4664 gnd.n4644 240.244
R6392 gnd.n4660 gnd.n4644 240.244
R6393 gnd.n4660 gnd.n4659 240.244
R6394 gnd.n4659 gnd.n4658 240.244
R6395 gnd.n4658 gnd.n4651 240.244
R6396 gnd.n4651 gnd.n2119 240.244
R6397 gnd.n4775 gnd.n2119 240.244
R6398 gnd.n4775 gnd.n2115 240.244
R6399 gnd.n4781 gnd.n2115 240.244
R6400 gnd.n4781 gnd.n2106 240.244
R6401 gnd.n4791 gnd.n2106 240.244
R6402 gnd.n4791 gnd.n2102 240.244
R6403 gnd.n4797 gnd.n2102 240.244
R6404 gnd.n4797 gnd.n2092 240.244
R6405 gnd.n4807 gnd.n2092 240.244
R6406 gnd.n4807 gnd.n2088 240.244
R6407 gnd.n4813 gnd.n2088 240.244
R6408 gnd.n4813 gnd.n2077 240.244
R6409 gnd.n4823 gnd.n2077 240.244
R6410 gnd.n4823 gnd.n2073 240.244
R6411 gnd.n4829 gnd.n2073 240.244
R6412 gnd.n4829 gnd.n2063 240.244
R6413 gnd.n4839 gnd.n2063 240.244
R6414 gnd.n4839 gnd.n2059 240.244
R6415 gnd.n4845 gnd.n2059 240.244
R6416 gnd.n4845 gnd.n2048 240.244
R6417 gnd.n4869 gnd.n2048 240.244
R6418 gnd.n4869 gnd.n2043 240.244
R6419 gnd.n4881 gnd.n2043 240.244
R6420 gnd.n4881 gnd.n2044 240.244
R6421 gnd.n4877 gnd.n2044 240.244
R6422 gnd.n4877 gnd.n1187 240.244
R6423 gnd.n6271 gnd.n1187 240.244
R6424 gnd.n6271 gnd.n1188 240.244
R6425 gnd.n6267 gnd.n1188 240.244
R6426 gnd.n6267 gnd.n1194 240.244
R6427 gnd.n5027 gnd.n1194 240.244
R6428 gnd.n5033 gnd.n5027 240.244
R6429 gnd.n5033 gnd.n2018 240.244
R6430 gnd.n5056 gnd.n2018 240.244
R6431 gnd.n5056 gnd.n2013 240.244
R6432 gnd.n5064 gnd.n2013 240.244
R6433 gnd.n5064 gnd.n2014 240.244
R6434 gnd.n2014 gnd.n1990 240.244
R6435 gnd.n5094 gnd.n1990 240.244
R6436 gnd.n5094 gnd.n1985 240.244
R6437 gnd.n5106 gnd.n1985 240.244
R6438 gnd.n5106 gnd.n1986 240.244
R6439 gnd.n5102 gnd.n1986 240.244
R6440 gnd.n5102 gnd.n1959 240.244
R6441 gnd.n5167 gnd.n1959 240.244
R6442 gnd.n5167 gnd.n1960 240.244
R6443 gnd.n5163 gnd.n1960 240.244
R6444 gnd.n5163 gnd.n1940 240.244
R6445 gnd.n5195 gnd.n1940 240.244
R6446 gnd.n5195 gnd.n1935 240.244
R6447 gnd.n5203 gnd.n1935 240.244
R6448 gnd.n5203 gnd.n1936 240.244
R6449 gnd.n1936 gnd.n1912 240.244
R6450 gnd.n5233 gnd.n1912 240.244
R6451 gnd.n5233 gnd.n1908 240.244
R6452 gnd.n5239 gnd.n1908 240.244
R6453 gnd.n5239 gnd.n1886 240.244
R6454 gnd.n5270 gnd.n1886 240.244
R6455 gnd.n5270 gnd.n1881 240.244
R6456 gnd.n5278 gnd.n1881 240.244
R6457 gnd.n5278 gnd.n1882 240.244
R6458 gnd.n1882 gnd.n1859 240.244
R6459 gnd.n5319 gnd.n1859 240.244
R6460 gnd.n5319 gnd.n1854 240.244
R6461 gnd.n5327 gnd.n1854 240.244
R6462 gnd.n5327 gnd.n1855 240.244
R6463 gnd.n1855 gnd.n1837 240.244
R6464 gnd.n5360 gnd.n1837 240.244
R6465 gnd.n5360 gnd.n1832 240.244
R6466 gnd.n5368 gnd.n1832 240.244
R6467 gnd.n5368 gnd.n1833 240.244
R6468 gnd.n1833 gnd.n1807 240.244
R6469 gnd.n5400 gnd.n1807 240.244
R6470 gnd.n5400 gnd.n1803 240.244
R6471 gnd.n5406 gnd.n1803 240.244
R6472 gnd.n5406 gnd.n1783 240.244
R6473 gnd.n5443 gnd.n1783 240.244
R6474 gnd.n5443 gnd.n1778 240.244
R6475 gnd.n5451 gnd.n1778 240.244
R6476 gnd.n5451 gnd.n1779 240.244
R6477 gnd.n1779 gnd.n1727 240.244
R6478 gnd.n5619 gnd.n1727 240.244
R6479 gnd.n5619 gnd.n1723 240.244
R6480 gnd.n5625 gnd.n1723 240.244
R6481 gnd.n5625 gnd.n1716 240.244
R6482 gnd.n5636 gnd.n1716 240.244
R6483 gnd.n5636 gnd.n1712 240.244
R6484 gnd.n5642 gnd.n1712 240.244
R6485 gnd.n5642 gnd.n1704 240.244
R6486 gnd.n5653 gnd.n1704 240.244
R6487 gnd.n5653 gnd.n1700 240.244
R6488 gnd.n5659 gnd.n1700 240.244
R6489 gnd.n5659 gnd.n1692 240.244
R6490 gnd.n5670 gnd.n1692 240.244
R6491 gnd.n5670 gnd.n1688 240.244
R6492 gnd.n5676 gnd.n1688 240.244
R6493 gnd.n5676 gnd.n1680 240.244
R6494 gnd.n5687 gnd.n1680 240.244
R6495 gnd.n5687 gnd.n1676 240.244
R6496 gnd.n5696 gnd.n1676 240.244
R6497 gnd.n5696 gnd.n1668 240.244
R6498 gnd.n5707 gnd.n1668 240.244
R6499 gnd.n5708 gnd.n5707 240.244
R6500 gnd.n5708 gnd.n1295 240.244
R6501 gnd.n1663 gnd.n1295 240.244
R6502 gnd.n5726 gnd.n1663 240.244
R6503 gnd.n5726 gnd.n1664 240.244
R6504 gnd.n5722 gnd.n1664 240.244
R6505 gnd.n5722 gnd.n5721 240.244
R6506 gnd.n5721 gnd.n5720 240.244
R6507 gnd.n5720 gnd.n1632 240.244
R6508 gnd.n5778 gnd.n1632 240.244
R6509 gnd.n5778 gnd.n1628 240.244
R6510 gnd.n5784 gnd.n1628 240.244
R6511 gnd.n5785 gnd.n5784 240.244
R6512 gnd.n5786 gnd.n5785 240.244
R6513 gnd.n5786 gnd.n1624 240.244
R6514 gnd.n5792 gnd.n1624 240.244
R6515 gnd.n5793 gnd.n5792 240.244
R6516 gnd.n5794 gnd.n5793 240.244
R6517 gnd.n5794 gnd.n1619 240.244
R6518 gnd.n5820 gnd.n1619 240.244
R6519 gnd.n5820 gnd.n1620 240.244
R6520 gnd.n5816 gnd.n1620 240.244
R6521 gnd.n5816 gnd.n5815 240.244
R6522 gnd.n5815 gnd.n5814 240.244
R6523 gnd.n5814 gnd.n5802 240.244
R6524 gnd.n5810 gnd.n5802 240.244
R6525 gnd.n5810 gnd.n1602 240.244
R6526 gnd.n5877 gnd.n1602 240.244
R6527 gnd.n5878 gnd.n5877 240.244
R6528 gnd.n5879 gnd.n5878 240.244
R6529 gnd.n5879 gnd.n1598 240.244
R6530 gnd.n5886 gnd.n1598 240.244
R6531 gnd.n5886 gnd.n387 240.244
R6532 gnd.n7280 gnd.n387 240.244
R6533 gnd.n7280 gnd.n388 240.244
R6534 gnd.n6641 gnd.n771 240.244
R6535 gnd.n6637 gnd.n771 240.244
R6536 gnd.n6637 gnd.n773 240.244
R6537 gnd.n6633 gnd.n773 240.244
R6538 gnd.n6633 gnd.n778 240.244
R6539 gnd.n6629 gnd.n778 240.244
R6540 gnd.n6629 gnd.n780 240.244
R6541 gnd.n6625 gnd.n780 240.244
R6542 gnd.n6625 gnd.n786 240.244
R6543 gnd.n6621 gnd.n786 240.244
R6544 gnd.n6621 gnd.n788 240.244
R6545 gnd.n6617 gnd.n788 240.244
R6546 gnd.n6617 gnd.n794 240.244
R6547 gnd.n6613 gnd.n794 240.244
R6548 gnd.n6613 gnd.n796 240.244
R6549 gnd.n6609 gnd.n796 240.244
R6550 gnd.n6609 gnd.n802 240.244
R6551 gnd.n6605 gnd.n802 240.244
R6552 gnd.n6605 gnd.n804 240.244
R6553 gnd.n6601 gnd.n804 240.244
R6554 gnd.n6601 gnd.n810 240.244
R6555 gnd.n6597 gnd.n810 240.244
R6556 gnd.n6597 gnd.n812 240.244
R6557 gnd.n6593 gnd.n812 240.244
R6558 gnd.n6593 gnd.n818 240.244
R6559 gnd.n6589 gnd.n818 240.244
R6560 gnd.n6589 gnd.n820 240.244
R6561 gnd.n6585 gnd.n820 240.244
R6562 gnd.n6585 gnd.n826 240.244
R6563 gnd.n6581 gnd.n826 240.244
R6564 gnd.n6581 gnd.n828 240.244
R6565 gnd.n6577 gnd.n828 240.244
R6566 gnd.n6577 gnd.n834 240.244
R6567 gnd.n6573 gnd.n834 240.244
R6568 gnd.n6573 gnd.n836 240.244
R6569 gnd.n6569 gnd.n836 240.244
R6570 gnd.n6569 gnd.n842 240.244
R6571 gnd.n6565 gnd.n842 240.244
R6572 gnd.n6565 gnd.n844 240.244
R6573 gnd.n6561 gnd.n844 240.244
R6574 gnd.n6561 gnd.n850 240.244
R6575 gnd.n6557 gnd.n850 240.244
R6576 gnd.n6557 gnd.n852 240.244
R6577 gnd.n6553 gnd.n852 240.244
R6578 gnd.n6553 gnd.n858 240.244
R6579 gnd.n6549 gnd.n858 240.244
R6580 gnd.n6549 gnd.n860 240.244
R6581 gnd.n6545 gnd.n860 240.244
R6582 gnd.n6545 gnd.n866 240.244
R6583 gnd.n6541 gnd.n866 240.244
R6584 gnd.n6541 gnd.n868 240.244
R6585 gnd.n6537 gnd.n868 240.244
R6586 gnd.n6537 gnd.n874 240.244
R6587 gnd.n6533 gnd.n874 240.244
R6588 gnd.n6533 gnd.n876 240.244
R6589 gnd.n6529 gnd.n876 240.244
R6590 gnd.n6529 gnd.n882 240.244
R6591 gnd.n6525 gnd.n882 240.244
R6592 gnd.n6525 gnd.n884 240.244
R6593 gnd.n6521 gnd.n884 240.244
R6594 gnd.n6521 gnd.n890 240.244
R6595 gnd.n6517 gnd.n890 240.244
R6596 gnd.n6517 gnd.n892 240.244
R6597 gnd.n6513 gnd.n892 240.244
R6598 gnd.n6513 gnd.n898 240.244
R6599 gnd.n6509 gnd.n898 240.244
R6600 gnd.n6509 gnd.n900 240.244
R6601 gnd.n6505 gnd.n900 240.244
R6602 gnd.n6505 gnd.n906 240.244
R6603 gnd.n6501 gnd.n906 240.244
R6604 gnd.n6501 gnd.n908 240.244
R6605 gnd.n6497 gnd.n908 240.244
R6606 gnd.n6497 gnd.n914 240.244
R6607 gnd.n6493 gnd.n914 240.244
R6608 gnd.n6493 gnd.n916 240.244
R6609 gnd.n6489 gnd.n916 240.244
R6610 gnd.n6489 gnd.n922 240.244
R6611 gnd.n6485 gnd.n922 240.244
R6612 gnd.n6485 gnd.n924 240.244
R6613 gnd.n6481 gnd.n924 240.244
R6614 gnd.n6481 gnd.n930 240.244
R6615 gnd.n6477 gnd.n930 240.244
R6616 gnd.n6477 gnd.n932 240.244
R6617 gnd.n6473 gnd.n932 240.244
R6618 gnd.n2137 gnd.n2113 240.244
R6619 gnd.n2137 gnd.n2107 240.244
R6620 gnd.n2138 gnd.n2107 240.244
R6621 gnd.n2138 gnd.n2101 240.244
R6622 gnd.n2141 gnd.n2101 240.244
R6623 gnd.n2141 gnd.n2094 240.244
R6624 gnd.n2142 gnd.n2094 240.244
R6625 gnd.n2142 gnd.n2087 240.244
R6626 gnd.n2145 gnd.n2087 240.244
R6627 gnd.n2145 gnd.n2079 240.244
R6628 gnd.n2146 gnd.n2079 240.244
R6629 gnd.n2146 gnd.n2072 240.244
R6630 gnd.n2149 gnd.n2072 240.244
R6631 gnd.n2149 gnd.n2065 240.244
R6632 gnd.n2150 gnd.n2065 240.244
R6633 gnd.n2150 gnd.n2058 240.244
R6634 gnd.n2153 gnd.n2058 240.244
R6635 gnd.n2153 gnd.n2050 240.244
R6636 gnd.n2050 gnd.n2039 240.244
R6637 gnd.n4883 gnd.n2039 240.244
R6638 gnd.n4884 gnd.n4883 240.244
R6639 gnd.n4886 gnd.n4884 240.244
R6640 gnd.n4886 gnd.n4885 240.244
R6641 gnd.n4885 gnd.n1185 240.244
R6642 gnd.n4991 gnd.n1185 240.244
R6643 gnd.n4991 gnd.n1195 240.244
R6644 gnd.n2032 gnd.n1195 240.244
R6645 gnd.n5025 gnd.n2032 240.244
R6646 gnd.n5025 gnd.n2030 240.244
R6647 gnd.n2030 gnd.n2026 240.244
R6648 gnd.n2026 gnd.n2019 240.244
R6649 gnd.n4997 gnd.n2019 240.244
R6650 gnd.n4997 gnd.n2011 240.244
R6651 gnd.n5000 gnd.n2011 240.244
R6652 gnd.n5001 gnd.n5000 240.244
R6653 gnd.n5001 gnd.n1991 240.244
R6654 gnd.n5002 gnd.n1991 240.244
R6655 gnd.n5002 gnd.n1984 240.244
R6656 gnd.n5006 gnd.n1984 240.244
R6657 gnd.n5006 gnd.n1972 240.244
R6658 gnd.n5128 gnd.n1972 240.244
R6659 gnd.n5128 gnd.n1956 240.244
R6660 gnd.n1967 gnd.n1956 240.244
R6661 gnd.n5161 gnd.n1967 240.244
R6662 gnd.n5161 gnd.n1949 240.244
R6663 gnd.n1949 gnd.n1941 240.244
R6664 gnd.n5134 gnd.n1941 240.244
R6665 gnd.n5134 gnd.n1933 240.244
R6666 gnd.n5137 gnd.n1933 240.244
R6667 gnd.n5138 gnd.n5137 240.244
R6668 gnd.n5138 gnd.n1914 240.244
R6669 gnd.n5139 gnd.n1914 240.244
R6670 gnd.n5139 gnd.n1906 240.244
R6671 gnd.n5142 gnd.n1906 240.244
R6672 gnd.n5142 gnd.n1888 240.244
R6673 gnd.n1888 gnd.n1879 240.244
R6674 gnd.n5280 gnd.n1879 240.244
R6675 gnd.n5280 gnd.n1874 240.244
R6676 gnd.n5287 gnd.n1874 240.244
R6677 gnd.n5287 gnd.n1861 240.244
R6678 gnd.n1861 gnd.n1852 240.244
R6679 gnd.n5329 gnd.n1852 240.244
R6680 gnd.n5329 gnd.n1847 240.244
R6681 gnd.n5351 gnd.n1847 240.244
R6682 gnd.n5351 gnd.n1839 240.244
R6683 gnd.n5334 gnd.n1839 240.244
R6684 gnd.n5334 gnd.n1829 240.244
R6685 gnd.n5335 gnd.n1829 240.244
R6686 gnd.n5336 gnd.n5335 240.244
R6687 gnd.n5336 gnd.n1809 240.244
R6688 gnd.n1809 gnd.n1800 240.244
R6689 gnd.n5408 gnd.n1800 240.244
R6690 gnd.n5409 gnd.n5408 240.244
R6691 gnd.n5409 gnd.n1785 240.244
R6692 gnd.n5425 gnd.n1785 240.244
R6693 gnd.n5425 gnd.n1775 240.244
R6694 gnd.n5414 gnd.n1775 240.244
R6695 gnd.n5416 gnd.n5414 240.244
R6696 gnd.n5416 gnd.n1729 240.244
R6697 gnd.n1729 gnd.n1722 240.244
R6698 gnd.n5627 gnd.n1722 240.244
R6699 gnd.n5627 gnd.n1718 240.244
R6700 gnd.n5633 gnd.n1718 240.244
R6701 gnd.n5633 gnd.n1710 240.244
R6702 gnd.n5644 gnd.n1710 240.244
R6703 gnd.n5644 gnd.n1706 240.244
R6704 gnd.n5650 gnd.n1706 240.244
R6705 gnd.n5650 gnd.n1698 240.244
R6706 gnd.n5661 gnd.n1698 240.244
R6707 gnd.n5661 gnd.n1694 240.244
R6708 gnd.n5667 gnd.n1694 240.244
R6709 gnd.n5667 gnd.n1685 240.244
R6710 gnd.n5678 gnd.n1685 240.244
R6711 gnd.n5678 gnd.n1681 240.244
R6712 gnd.n5684 gnd.n1681 240.244
R6713 gnd.n5684 gnd.n1674 240.244
R6714 gnd.n5698 gnd.n1674 240.244
R6715 gnd.n5698 gnd.n1670 240.244
R6716 gnd.n5704 gnd.n1670 240.244
R6717 gnd.n5704 gnd.n1297 240.244
R6718 gnd.n6148 gnd.n1297 240.244
R6719 gnd.n2135 gnd.n2134 240.244
R6720 gnd.n2189 gnd.n2134 240.244
R6721 gnd.n2191 gnd.n2190 240.244
R6722 gnd.n2308 gnd.n2307 240.244
R6723 gnd.n2310 gnd.n2309 240.244
R6724 gnd.n2321 gnd.n2320 240.244
R6725 gnd.n2323 gnd.n2322 240.244
R6726 gnd.n2333 gnd.n2332 240.244
R6727 gnd.n2344 gnd.n2343 240.244
R6728 gnd.n2346 gnd.n2345 240.244
R6729 gnd.n2356 gnd.n2355 240.244
R6730 gnd.n2367 gnd.n2366 240.244
R6731 gnd.n4700 gnd.n2368 240.244
R6732 gnd.n4704 gnd.n4703 240.244
R6733 gnd.n4783 gnd.n2108 240.244
R6734 gnd.n4789 gnd.n2108 240.244
R6735 gnd.n4789 gnd.n2099 240.244
R6736 gnd.n4799 gnd.n2099 240.244
R6737 gnd.n4799 gnd.n2095 240.244
R6738 gnd.n4805 gnd.n2095 240.244
R6739 gnd.n4805 gnd.n2085 240.244
R6740 gnd.n4815 gnd.n2085 240.244
R6741 gnd.n4815 gnd.n2081 240.244
R6742 gnd.n4821 gnd.n2081 240.244
R6743 gnd.n4821 gnd.n2071 240.244
R6744 gnd.n4831 gnd.n2071 240.244
R6745 gnd.n4831 gnd.n2067 240.244
R6746 gnd.n4837 gnd.n2067 240.244
R6747 gnd.n4837 gnd.n2057 240.244
R6748 gnd.n4847 gnd.n2057 240.244
R6749 gnd.n4847 gnd.n2051 240.244
R6750 gnd.n4867 gnd.n2051 240.244
R6751 gnd.n4867 gnd.n2052 240.244
R6752 gnd.n2052 gnd.n2042 240.244
R6753 gnd.n4852 gnd.n2042 240.244
R6754 gnd.n4853 gnd.n4852 240.244
R6755 gnd.n4854 gnd.n4853 240.244
R6756 gnd.n4854 gnd.n1186 240.244
R6757 gnd.n1196 gnd.n1186 240.244
R6758 gnd.n6265 gnd.n1196 240.244
R6759 gnd.n6265 gnd.n1197 240.244
R6760 gnd.n1202 gnd.n1197 240.244
R6761 gnd.n1203 gnd.n1202 240.244
R6762 gnd.n1204 gnd.n1203 240.244
R6763 gnd.n5054 gnd.n1204 240.244
R6764 gnd.n5054 gnd.n1207 240.244
R6765 gnd.n1208 gnd.n1207 240.244
R6766 gnd.n1209 gnd.n1208 240.244
R6767 gnd.n1998 gnd.n1209 240.244
R6768 gnd.n1998 gnd.n1212 240.244
R6769 gnd.n1213 gnd.n1212 240.244
R6770 gnd.n1214 gnd.n1213 240.244
R6771 gnd.n1978 gnd.n1214 240.244
R6772 gnd.n1978 gnd.n1217 240.244
R6773 gnd.n1218 gnd.n1217 240.244
R6774 gnd.n1219 gnd.n1218 240.244
R6775 gnd.n1965 gnd.n1219 240.244
R6776 gnd.n1965 gnd.n1222 240.244
R6777 gnd.n1223 gnd.n1222 240.244
R6778 gnd.n1224 gnd.n1223 240.244
R6779 gnd.n1930 gnd.n1224 240.244
R6780 gnd.n1930 gnd.n1227 240.244
R6781 gnd.n1228 gnd.n1227 240.244
R6782 gnd.n1229 gnd.n1228 240.244
R6783 gnd.n5231 gnd.n1229 240.244
R6784 gnd.n5231 gnd.n1232 240.244
R6785 gnd.n1233 gnd.n1232 240.244
R6786 gnd.n1234 gnd.n1233 240.244
R6787 gnd.n5268 gnd.n1234 240.244
R6788 gnd.n5268 gnd.n1237 240.244
R6789 gnd.n1238 gnd.n1237 240.244
R6790 gnd.n1239 gnd.n1238 240.244
R6791 gnd.n5288 gnd.n1239 240.244
R6792 gnd.n5288 gnd.n1242 240.244
R6793 gnd.n1243 gnd.n1242 240.244
R6794 gnd.n1244 gnd.n1243 240.244
R6795 gnd.n5308 gnd.n1244 240.244
R6796 gnd.n5308 gnd.n1247 240.244
R6797 gnd.n1248 gnd.n1247 240.244
R6798 gnd.n1249 gnd.n1248 240.244
R6799 gnd.n1831 gnd.n1249 240.244
R6800 gnd.n1831 gnd.n1252 240.244
R6801 gnd.n1253 gnd.n1252 240.244
R6802 gnd.n1254 gnd.n1253 240.244
R6803 gnd.n1811 gnd.n1254 240.244
R6804 gnd.n1811 gnd.n1257 240.244
R6805 gnd.n1258 gnd.n1257 240.244
R6806 gnd.n1259 gnd.n1258 240.244
R6807 gnd.n5426 gnd.n1259 240.244
R6808 gnd.n5426 gnd.n1262 240.244
R6809 gnd.n1263 gnd.n1262 240.244
R6810 gnd.n1264 gnd.n1263 240.244
R6811 gnd.n5617 gnd.n1264 240.244
R6812 gnd.n5617 gnd.n1267 240.244
R6813 gnd.n1268 gnd.n1267 240.244
R6814 gnd.n1269 gnd.n1268 240.244
R6815 gnd.n5634 gnd.n1269 240.244
R6816 gnd.n5634 gnd.n1272 240.244
R6817 gnd.n1273 gnd.n1272 240.244
R6818 gnd.n1274 gnd.n1273 240.244
R6819 gnd.n5651 gnd.n1274 240.244
R6820 gnd.n5651 gnd.n1277 240.244
R6821 gnd.n1278 gnd.n1277 240.244
R6822 gnd.n1279 gnd.n1278 240.244
R6823 gnd.n5668 gnd.n1279 240.244
R6824 gnd.n5668 gnd.n1282 240.244
R6825 gnd.n1283 gnd.n1282 240.244
R6826 gnd.n1284 gnd.n1283 240.244
R6827 gnd.n5685 gnd.n1284 240.244
R6828 gnd.n5685 gnd.n1287 240.244
R6829 gnd.n1288 gnd.n1287 240.244
R6830 gnd.n1289 gnd.n1288 240.244
R6831 gnd.n5705 gnd.n1289 240.244
R6832 gnd.n5705 gnd.n1292 240.244
R6833 gnd.n6150 gnd.n1292 240.244
R6834 gnd.n1303 gnd.n1302 240.244
R6835 gnd.n1641 gnd.n1306 240.244
R6836 gnd.n1308 gnd.n1307 240.244
R6837 gnd.n1644 gnd.n1312 240.244
R6838 gnd.n1647 gnd.n1313 240.244
R6839 gnd.n1322 gnd.n1321 240.244
R6840 gnd.n1649 gnd.n1329 240.244
R6841 gnd.n1652 gnd.n1330 240.244
R6842 gnd.n1338 gnd.n1337 240.244
R6843 gnd.n1654 gnd.n1345 240.244
R6844 gnd.n1657 gnd.n1346 240.244
R6845 gnd.n1354 gnd.n1353 240.244
R6846 gnd.n1660 gnd.n1354 240.244
R6847 gnd.n5730 gnd.n1639 240.244
R6848 gnd.n1167 gnd.n1166 240.132
R6849 gnd.n5467 gnd.n5466 240.132
R6850 gnd.n6648 gnd.n766 225.874
R6851 gnd.n6649 gnd.n6648 225.874
R6852 gnd.n6650 gnd.n6649 225.874
R6853 gnd.n6650 gnd.n760 225.874
R6854 gnd.n6658 gnd.n760 225.874
R6855 gnd.n6659 gnd.n6658 225.874
R6856 gnd.n6660 gnd.n6659 225.874
R6857 gnd.n6660 gnd.n754 225.874
R6858 gnd.n6668 gnd.n754 225.874
R6859 gnd.n6669 gnd.n6668 225.874
R6860 gnd.n6670 gnd.n6669 225.874
R6861 gnd.n6670 gnd.n748 225.874
R6862 gnd.n6678 gnd.n748 225.874
R6863 gnd.n6679 gnd.n6678 225.874
R6864 gnd.n6680 gnd.n6679 225.874
R6865 gnd.n6680 gnd.n742 225.874
R6866 gnd.n6688 gnd.n742 225.874
R6867 gnd.n6689 gnd.n6688 225.874
R6868 gnd.n6690 gnd.n6689 225.874
R6869 gnd.n6690 gnd.n736 225.874
R6870 gnd.n6698 gnd.n736 225.874
R6871 gnd.n6699 gnd.n6698 225.874
R6872 gnd.n6700 gnd.n6699 225.874
R6873 gnd.n6700 gnd.n730 225.874
R6874 gnd.n6708 gnd.n730 225.874
R6875 gnd.n6709 gnd.n6708 225.874
R6876 gnd.n6710 gnd.n6709 225.874
R6877 gnd.n6710 gnd.n724 225.874
R6878 gnd.n6718 gnd.n724 225.874
R6879 gnd.n6719 gnd.n6718 225.874
R6880 gnd.n6720 gnd.n6719 225.874
R6881 gnd.n6720 gnd.n718 225.874
R6882 gnd.n6728 gnd.n718 225.874
R6883 gnd.n6729 gnd.n6728 225.874
R6884 gnd.n6730 gnd.n6729 225.874
R6885 gnd.n6730 gnd.n712 225.874
R6886 gnd.n6738 gnd.n712 225.874
R6887 gnd.n6739 gnd.n6738 225.874
R6888 gnd.n6740 gnd.n6739 225.874
R6889 gnd.n6740 gnd.n706 225.874
R6890 gnd.n6748 gnd.n706 225.874
R6891 gnd.n6749 gnd.n6748 225.874
R6892 gnd.n6750 gnd.n6749 225.874
R6893 gnd.n6750 gnd.n700 225.874
R6894 gnd.n6758 gnd.n700 225.874
R6895 gnd.n6759 gnd.n6758 225.874
R6896 gnd.n6760 gnd.n6759 225.874
R6897 gnd.n6760 gnd.n694 225.874
R6898 gnd.n6768 gnd.n694 225.874
R6899 gnd.n6769 gnd.n6768 225.874
R6900 gnd.n6770 gnd.n6769 225.874
R6901 gnd.n6770 gnd.n688 225.874
R6902 gnd.n6778 gnd.n688 225.874
R6903 gnd.n6779 gnd.n6778 225.874
R6904 gnd.n6780 gnd.n6779 225.874
R6905 gnd.n6780 gnd.n682 225.874
R6906 gnd.n6788 gnd.n682 225.874
R6907 gnd.n6789 gnd.n6788 225.874
R6908 gnd.n6790 gnd.n6789 225.874
R6909 gnd.n6790 gnd.n676 225.874
R6910 gnd.n6798 gnd.n676 225.874
R6911 gnd.n6799 gnd.n6798 225.874
R6912 gnd.n6800 gnd.n6799 225.874
R6913 gnd.n6800 gnd.n670 225.874
R6914 gnd.n6808 gnd.n670 225.874
R6915 gnd.n6809 gnd.n6808 225.874
R6916 gnd.n6810 gnd.n6809 225.874
R6917 gnd.n6810 gnd.n664 225.874
R6918 gnd.n6818 gnd.n664 225.874
R6919 gnd.n6819 gnd.n6818 225.874
R6920 gnd.n6820 gnd.n6819 225.874
R6921 gnd.n6820 gnd.n658 225.874
R6922 gnd.n6828 gnd.n658 225.874
R6923 gnd.n6829 gnd.n6828 225.874
R6924 gnd.n6830 gnd.n6829 225.874
R6925 gnd.n6830 gnd.n652 225.874
R6926 gnd.n6838 gnd.n652 225.874
R6927 gnd.n6839 gnd.n6838 225.874
R6928 gnd.n6840 gnd.n6839 225.874
R6929 gnd.n6840 gnd.n646 225.874
R6930 gnd.n6848 gnd.n646 225.874
R6931 gnd.n6849 gnd.n6848 225.874
R6932 gnd.n6850 gnd.n6849 225.874
R6933 gnd.n6850 gnd.n640 225.874
R6934 gnd.n6858 gnd.n640 225.874
R6935 gnd.n6859 gnd.n6858 225.874
R6936 gnd.n6860 gnd.n6859 225.874
R6937 gnd.n6860 gnd.n634 225.874
R6938 gnd.n6868 gnd.n634 225.874
R6939 gnd.n6869 gnd.n6868 225.874
R6940 gnd.n6870 gnd.n6869 225.874
R6941 gnd.n6870 gnd.n628 225.874
R6942 gnd.n6878 gnd.n628 225.874
R6943 gnd.n6879 gnd.n6878 225.874
R6944 gnd.n6880 gnd.n6879 225.874
R6945 gnd.n6880 gnd.n622 225.874
R6946 gnd.n6888 gnd.n622 225.874
R6947 gnd.n6889 gnd.n6888 225.874
R6948 gnd.n6890 gnd.n6889 225.874
R6949 gnd.n6890 gnd.n616 225.874
R6950 gnd.n6898 gnd.n616 225.874
R6951 gnd.n6899 gnd.n6898 225.874
R6952 gnd.n6900 gnd.n6899 225.874
R6953 gnd.n6900 gnd.n610 225.874
R6954 gnd.n6908 gnd.n610 225.874
R6955 gnd.n6909 gnd.n6908 225.874
R6956 gnd.n6910 gnd.n6909 225.874
R6957 gnd.n6910 gnd.n604 225.874
R6958 gnd.n6918 gnd.n604 225.874
R6959 gnd.n6919 gnd.n6918 225.874
R6960 gnd.n6920 gnd.n6919 225.874
R6961 gnd.n6920 gnd.n598 225.874
R6962 gnd.n6928 gnd.n598 225.874
R6963 gnd.n6929 gnd.n6928 225.874
R6964 gnd.n6930 gnd.n6929 225.874
R6965 gnd.n6930 gnd.n592 225.874
R6966 gnd.n6938 gnd.n592 225.874
R6967 gnd.n6939 gnd.n6938 225.874
R6968 gnd.n6940 gnd.n6939 225.874
R6969 gnd.n6940 gnd.n586 225.874
R6970 gnd.n6948 gnd.n586 225.874
R6971 gnd.n6949 gnd.n6948 225.874
R6972 gnd.n6950 gnd.n6949 225.874
R6973 gnd.n6950 gnd.n580 225.874
R6974 gnd.n6958 gnd.n580 225.874
R6975 gnd.n6959 gnd.n6958 225.874
R6976 gnd.n6960 gnd.n6959 225.874
R6977 gnd.n6960 gnd.n574 225.874
R6978 gnd.n6968 gnd.n574 225.874
R6979 gnd.n6969 gnd.n6968 225.874
R6980 gnd.n6970 gnd.n6969 225.874
R6981 gnd.n6970 gnd.n568 225.874
R6982 gnd.n6978 gnd.n568 225.874
R6983 gnd.n6979 gnd.n6978 225.874
R6984 gnd.n6980 gnd.n6979 225.874
R6985 gnd.n6980 gnd.n562 225.874
R6986 gnd.n6988 gnd.n562 225.874
R6987 gnd.n6989 gnd.n6988 225.874
R6988 gnd.n6990 gnd.n6989 225.874
R6989 gnd.n6990 gnd.n556 225.874
R6990 gnd.n6998 gnd.n556 225.874
R6991 gnd.n6999 gnd.n6998 225.874
R6992 gnd.n7000 gnd.n6999 225.874
R6993 gnd.n7000 gnd.n550 225.874
R6994 gnd.n7008 gnd.n550 225.874
R6995 gnd.n7009 gnd.n7008 225.874
R6996 gnd.n7010 gnd.n7009 225.874
R6997 gnd.n7010 gnd.n544 225.874
R6998 gnd.n7018 gnd.n544 225.874
R6999 gnd.n7019 gnd.n7018 225.874
R7000 gnd.n7020 gnd.n7019 225.874
R7001 gnd.n7020 gnd.n538 225.874
R7002 gnd.n7028 gnd.n538 225.874
R7003 gnd.n7029 gnd.n7028 225.874
R7004 gnd.n7030 gnd.n7029 225.874
R7005 gnd.n7030 gnd.n532 225.874
R7006 gnd.n7038 gnd.n532 225.874
R7007 gnd.n7039 gnd.n7038 225.874
R7008 gnd.n7040 gnd.n7039 225.874
R7009 gnd.n7040 gnd.n526 225.874
R7010 gnd.n7048 gnd.n526 225.874
R7011 gnd.n7049 gnd.n7048 225.874
R7012 gnd.n7050 gnd.n7049 225.874
R7013 gnd.n7050 gnd.n520 225.874
R7014 gnd.n7058 gnd.n520 225.874
R7015 gnd.n7059 gnd.n7058 225.874
R7016 gnd.n7060 gnd.n7059 225.874
R7017 gnd.n3136 gnd.t185 224.174
R7018 gnd.n2630 gnd.t171 224.174
R7019 gnd.n1438 gnd.n1375 199.319
R7020 gnd.n1438 gnd.n1376 199.319
R7021 gnd.n1119 gnd.n1118 199.319
R7022 gnd.n2228 gnd.n1119 199.319
R7023 gnd.n1168 gnd.n1165 186.49
R7024 gnd.n5468 gnd.n5465 186.49
R7025 gnd.n3912 gnd.n3911 185
R7026 gnd.n3910 gnd.n3909 185
R7027 gnd.n3889 gnd.n3888 185
R7028 gnd.n3904 gnd.n3903 185
R7029 gnd.n3902 gnd.n3901 185
R7030 gnd.n3893 gnd.n3892 185
R7031 gnd.n3896 gnd.n3895 185
R7032 gnd.n3880 gnd.n3879 185
R7033 gnd.n3878 gnd.n3877 185
R7034 gnd.n3857 gnd.n3856 185
R7035 gnd.n3872 gnd.n3871 185
R7036 gnd.n3870 gnd.n3869 185
R7037 gnd.n3861 gnd.n3860 185
R7038 gnd.n3864 gnd.n3863 185
R7039 gnd.n3848 gnd.n3847 185
R7040 gnd.n3846 gnd.n3845 185
R7041 gnd.n3825 gnd.n3824 185
R7042 gnd.n3840 gnd.n3839 185
R7043 gnd.n3838 gnd.n3837 185
R7044 gnd.n3829 gnd.n3828 185
R7045 gnd.n3832 gnd.n3831 185
R7046 gnd.n3817 gnd.n3816 185
R7047 gnd.n3815 gnd.n3814 185
R7048 gnd.n3794 gnd.n3793 185
R7049 gnd.n3809 gnd.n3808 185
R7050 gnd.n3807 gnd.n3806 185
R7051 gnd.n3798 gnd.n3797 185
R7052 gnd.n3801 gnd.n3800 185
R7053 gnd.n3785 gnd.n3784 185
R7054 gnd.n3783 gnd.n3782 185
R7055 gnd.n3762 gnd.n3761 185
R7056 gnd.n3777 gnd.n3776 185
R7057 gnd.n3775 gnd.n3774 185
R7058 gnd.n3766 gnd.n3765 185
R7059 gnd.n3769 gnd.n3768 185
R7060 gnd.n3753 gnd.n3752 185
R7061 gnd.n3751 gnd.n3750 185
R7062 gnd.n3730 gnd.n3729 185
R7063 gnd.n3745 gnd.n3744 185
R7064 gnd.n3743 gnd.n3742 185
R7065 gnd.n3734 gnd.n3733 185
R7066 gnd.n3737 gnd.n3736 185
R7067 gnd.n3721 gnd.n3720 185
R7068 gnd.n3719 gnd.n3718 185
R7069 gnd.n3698 gnd.n3697 185
R7070 gnd.n3713 gnd.n3712 185
R7071 gnd.n3711 gnd.n3710 185
R7072 gnd.n3702 gnd.n3701 185
R7073 gnd.n3705 gnd.n3704 185
R7074 gnd.n3690 gnd.n3689 185
R7075 gnd.n3688 gnd.n3687 185
R7076 gnd.n3667 gnd.n3666 185
R7077 gnd.n3682 gnd.n3681 185
R7078 gnd.n3680 gnd.n3679 185
R7079 gnd.n3671 gnd.n3670 185
R7080 gnd.n3674 gnd.n3673 185
R7081 gnd.n3137 gnd.t184 178.987
R7082 gnd.n2631 gnd.t172 178.987
R7083 gnd.n1 gnd.t7 170.774
R7084 gnd.n9 gnd.t50 170.103
R7085 gnd.n8 gnd.t20 170.103
R7086 gnd.n7 gnd.t57 170.103
R7087 gnd.n6 gnd.t355 170.103
R7088 gnd.n5 gnd.t363 170.103
R7089 gnd.n4 gnd.t12 170.103
R7090 gnd.n3 gnd.t18 170.103
R7091 gnd.n2 gnd.t65 170.103
R7092 gnd.n1 gnd.t53 170.103
R7093 gnd.n6028 gnd.n1437 167.873
R7094 gnd.n6347 gnd.n6346 167.873
R7095 gnd.n5539 gnd.n5538 163.367
R7096 gnd.n5535 gnd.n5534 163.367
R7097 gnd.n5531 gnd.n5530 163.367
R7098 gnd.n5527 gnd.n5526 163.367
R7099 gnd.n5523 gnd.n5522 163.367
R7100 gnd.n5519 gnd.n5518 163.367
R7101 gnd.n5515 gnd.n5514 163.367
R7102 gnd.n5511 gnd.n5510 163.367
R7103 gnd.n5507 gnd.n5506 163.367
R7104 gnd.n5503 gnd.n5502 163.367
R7105 gnd.n5499 gnd.n5498 163.367
R7106 gnd.n5495 gnd.n5494 163.367
R7107 gnd.n5491 gnd.n5490 163.367
R7108 gnd.n5487 gnd.n5486 163.367
R7109 gnd.n5482 gnd.n5481 163.367
R7110 gnd.n5478 gnd.n5477 163.367
R7111 gnd.n5615 gnd.n5614 163.367
R7112 gnd.n5611 gnd.n5610 163.367
R7113 gnd.n5606 gnd.n5605 163.367
R7114 gnd.n5602 gnd.n5601 163.367
R7115 gnd.n5598 gnd.n5597 163.367
R7116 gnd.n5594 gnd.n5593 163.367
R7117 gnd.n5590 gnd.n5589 163.367
R7118 gnd.n5586 gnd.n5585 163.367
R7119 gnd.n5582 gnd.n5581 163.367
R7120 gnd.n5578 gnd.n5577 163.367
R7121 gnd.n5574 gnd.n5573 163.367
R7122 gnd.n5570 gnd.n5569 163.367
R7123 gnd.n5566 gnd.n5565 163.367
R7124 gnd.n5562 gnd.n5561 163.367
R7125 gnd.n5558 gnd.n5557 163.367
R7126 gnd.n5554 gnd.n5553 163.367
R7127 gnd.n4962 gnd.n1184 163.367
R7128 gnd.n4894 gnd.n1184 163.367
R7129 gnd.n4989 gnd.n4894 163.367
R7130 gnd.n4989 gnd.n4895 163.367
R7131 gnd.n4985 gnd.n4895 163.367
R7132 gnd.n4985 gnd.n4969 163.367
R7133 gnd.n4969 gnd.n4968 163.367
R7134 gnd.n4968 gnd.n2028 163.367
R7135 gnd.n5036 gnd.n2028 163.367
R7136 gnd.n5036 gnd.n2025 163.367
R7137 gnd.n5044 gnd.n2025 163.367
R7138 gnd.n5044 gnd.n2020 163.367
R7139 gnd.n5040 gnd.n2020 163.367
R7140 gnd.n5040 gnd.n2010 163.367
R7141 gnd.n2010 gnd.n2003 163.367
R7142 gnd.n5073 gnd.n2003 163.367
R7143 gnd.n5073 gnd.n2000 163.367
R7144 gnd.n5082 gnd.n2000 163.367
R7145 gnd.n5082 gnd.n2001 163.367
R7146 gnd.n2001 gnd.n1992 163.367
R7147 gnd.n5077 gnd.n1992 163.367
R7148 gnd.n5077 gnd.n1982 163.367
R7149 gnd.n5109 gnd.n1982 163.367
R7150 gnd.n5109 gnd.n1980 163.367
R7151 gnd.n5118 gnd.n1980 163.367
R7152 gnd.n5118 gnd.n1974 163.367
R7153 gnd.n5114 gnd.n1974 163.367
R7154 gnd.n5114 gnd.n1958 163.367
R7155 gnd.n1958 gnd.n1951 163.367
R7156 gnd.n5175 gnd.n1951 163.367
R7157 gnd.n5176 gnd.n5175 163.367
R7158 gnd.n5176 gnd.n1948 163.367
R7159 gnd.n5184 gnd.n1948 163.367
R7160 gnd.n5184 gnd.n1942 163.367
R7161 gnd.n5180 gnd.n1942 163.367
R7162 gnd.n5180 gnd.n1932 163.367
R7163 gnd.n1932 gnd.n1924 163.367
R7164 gnd.n5212 gnd.n1924 163.367
R7165 gnd.n5212 gnd.n1921 163.367
R7166 gnd.n5223 gnd.n1921 163.367
R7167 gnd.n5223 gnd.n1922 163.367
R7168 gnd.n1922 gnd.n1915 163.367
R7169 gnd.n5218 gnd.n1915 163.367
R7170 gnd.n5218 gnd.n1905 163.367
R7171 gnd.n1905 gnd.n1900 163.367
R7172 gnd.n5248 gnd.n1900 163.367
R7173 gnd.n5249 gnd.n5248 163.367
R7174 gnd.n5249 gnd.n1889 163.367
R7175 gnd.n5253 gnd.n1889 163.367
R7176 gnd.n5253 gnd.n1898 163.367
R7177 gnd.n5258 gnd.n1898 163.367
R7178 gnd.n5258 gnd.n1871 163.367
R7179 gnd.n5290 gnd.n1871 163.367
R7180 gnd.n5291 gnd.n5290 163.367
R7181 gnd.n5291 gnd.n1862 163.367
R7182 gnd.n5295 gnd.n1862 163.367
R7183 gnd.n5295 gnd.n1868 163.367
R7184 gnd.n5307 gnd.n1868 163.367
R7185 gnd.n5307 gnd.n1869 163.367
R7186 gnd.n1869 gnd.n1846 163.367
R7187 gnd.n5302 gnd.n1846 163.367
R7188 gnd.n5302 gnd.n1840 163.367
R7189 gnd.n5299 gnd.n1840 163.367
R7190 gnd.n5299 gnd.n1828 163.367
R7191 gnd.n1828 gnd.n1821 163.367
R7192 gnd.n5377 gnd.n1821 163.367
R7193 gnd.n5377 gnd.n1818 163.367
R7194 gnd.n5388 gnd.n1818 163.367
R7195 gnd.n5388 gnd.n1819 163.367
R7196 gnd.n1819 gnd.n1810 163.367
R7197 gnd.n5383 gnd.n1810 163.367
R7198 gnd.n5383 gnd.n5381 163.367
R7199 gnd.n5381 gnd.n1791 163.367
R7200 gnd.n5434 gnd.n1791 163.367
R7201 gnd.n5434 gnd.n1792 163.367
R7202 gnd.n1792 gnd.n1786 163.367
R7203 gnd.n5429 gnd.n1786 163.367
R7204 gnd.n5429 gnd.n1777 163.367
R7205 gnd.n1777 gnd.n1768 163.367
R7206 gnd.n5548 gnd.n1768 163.367
R7207 gnd.n5549 gnd.n5548 163.367
R7208 gnd.n1159 gnd.n1158 163.367
R7209 gnd.n6336 gnd.n1158 163.367
R7210 gnd.n6334 gnd.n6333 163.367
R7211 gnd.n6330 gnd.n6329 163.367
R7212 gnd.n6326 gnd.n6325 163.367
R7213 gnd.n6322 gnd.n6321 163.367
R7214 gnd.n6318 gnd.n6317 163.367
R7215 gnd.n6314 gnd.n6313 163.367
R7216 gnd.n6310 gnd.n6309 163.367
R7217 gnd.n6306 gnd.n6305 163.367
R7218 gnd.n6302 gnd.n6301 163.367
R7219 gnd.n6298 gnd.n6297 163.367
R7220 gnd.n6294 gnd.n6293 163.367
R7221 gnd.n6290 gnd.n6289 163.367
R7222 gnd.n6286 gnd.n6285 163.367
R7223 gnd.n6282 gnd.n6281 163.367
R7224 gnd.n6345 gnd.n1124 163.367
R7225 gnd.n4900 gnd.n4899 163.367
R7226 gnd.n4905 gnd.n4904 163.367
R7227 gnd.n4909 gnd.n4908 163.367
R7228 gnd.n4913 gnd.n4912 163.367
R7229 gnd.n4917 gnd.n4916 163.367
R7230 gnd.n4921 gnd.n4920 163.367
R7231 gnd.n4925 gnd.n4924 163.367
R7232 gnd.n4929 gnd.n4928 163.367
R7233 gnd.n4933 gnd.n4932 163.367
R7234 gnd.n4937 gnd.n4936 163.367
R7235 gnd.n4941 gnd.n4940 163.367
R7236 gnd.n4945 gnd.n4944 163.367
R7237 gnd.n4949 gnd.n4948 163.367
R7238 gnd.n4953 gnd.n4952 163.367
R7239 gnd.n4957 gnd.n4956 163.367
R7240 gnd.n6274 gnd.n1160 163.367
R7241 gnd.n6274 gnd.n1182 163.367
R7242 gnd.n4893 gnd.n1182 163.367
R7243 gnd.n4972 gnd.n4893 163.367
R7244 gnd.n4983 gnd.n4972 163.367
R7245 gnd.n4983 gnd.n4974 163.367
R7246 gnd.n4979 gnd.n4974 163.367
R7247 gnd.n4979 gnd.n4978 163.367
R7248 gnd.n4978 gnd.n2024 163.367
R7249 gnd.n5048 gnd.n2024 163.367
R7250 gnd.n5048 gnd.n2022 163.367
R7251 gnd.n5052 gnd.n2022 163.367
R7252 gnd.n5052 gnd.n2008 163.367
R7253 gnd.n5067 gnd.n2008 163.367
R7254 gnd.n5067 gnd.n2006 163.367
R7255 gnd.n5071 gnd.n2006 163.367
R7256 gnd.n5071 gnd.n1997 163.367
R7257 gnd.n5084 gnd.n1997 163.367
R7258 gnd.n5084 gnd.n1994 163.367
R7259 gnd.n5091 gnd.n1994 163.367
R7260 gnd.n5091 gnd.n1995 163.367
R7261 gnd.n5087 gnd.n1995 163.367
R7262 gnd.n5087 gnd.n1977 163.367
R7263 gnd.n5121 gnd.n1977 163.367
R7264 gnd.n5121 gnd.n1975 163.367
R7265 gnd.n5125 gnd.n1975 163.367
R7266 gnd.n5125 gnd.n1954 163.367
R7267 gnd.n5169 gnd.n1954 163.367
R7268 gnd.n5169 gnd.n1952 163.367
R7269 gnd.n5173 gnd.n1952 163.367
R7270 gnd.n5173 gnd.n1946 163.367
R7271 gnd.n5188 gnd.n1946 163.367
R7272 gnd.n5188 gnd.n1944 163.367
R7273 gnd.n5192 gnd.n1944 163.367
R7274 gnd.n5192 gnd.n1929 163.367
R7275 gnd.n5206 gnd.n1929 163.367
R7276 gnd.n5206 gnd.n1927 163.367
R7277 gnd.n5210 gnd.n1927 163.367
R7278 gnd.n5210 gnd.n1919 163.367
R7279 gnd.n5225 gnd.n1919 163.367
R7280 gnd.n5225 gnd.n1917 163.367
R7281 gnd.n5229 gnd.n1917 163.367
R7282 gnd.n5229 gnd.n1904 163.367
R7283 gnd.n5242 gnd.n1904 163.367
R7284 gnd.n5242 gnd.n1902 163.367
R7285 gnd.n5246 gnd.n1902 163.367
R7286 gnd.n5246 gnd.n1891 163.367
R7287 gnd.n5266 gnd.n1891 163.367
R7288 gnd.n5266 gnd.n1892 163.367
R7289 gnd.n5262 gnd.n1892 163.367
R7290 gnd.n5262 gnd.n5261 163.367
R7291 gnd.n5261 gnd.n1897 163.367
R7292 gnd.n1897 gnd.n1873 163.367
R7293 gnd.n1873 gnd.n1864 163.367
R7294 gnd.n5316 gnd.n1864 163.367
R7295 gnd.n5316 gnd.n1865 163.367
R7296 gnd.n5312 gnd.n1865 163.367
R7297 gnd.n5312 gnd.n5311 163.367
R7298 gnd.n5311 gnd.n1844 163.367
R7299 gnd.n5354 gnd.n1844 163.367
R7300 gnd.n5354 gnd.n1842 163.367
R7301 gnd.n5358 gnd.n1842 163.367
R7302 gnd.n5358 gnd.n1826 163.367
R7303 gnd.n5371 gnd.n1826 163.367
R7304 gnd.n5371 gnd.n1824 163.367
R7305 gnd.n5375 gnd.n1824 163.367
R7306 gnd.n5375 gnd.n1816 163.367
R7307 gnd.n5390 gnd.n1816 163.367
R7308 gnd.n5390 gnd.n1813 163.367
R7309 gnd.n5397 gnd.n1813 163.367
R7310 gnd.n5397 gnd.n1814 163.367
R7311 gnd.n5393 gnd.n1814 163.367
R7312 gnd.n5393 gnd.n1789 163.367
R7313 gnd.n5436 gnd.n1789 163.367
R7314 gnd.n5436 gnd.n1787 163.367
R7315 gnd.n5440 gnd.n1787 163.367
R7316 gnd.n5440 gnd.n1774 163.367
R7317 gnd.n5453 gnd.n1774 163.367
R7318 gnd.n5453 gnd.n1771 163.367
R7319 gnd.n5546 gnd.n1771 163.367
R7320 gnd.n5546 gnd.n1772 163.367
R7321 gnd.n5474 gnd.n5473 156.462
R7322 gnd.n3852 gnd.n3820 153.042
R7323 gnd.n3916 gnd.n3915 152.079
R7324 gnd.n3884 gnd.n3883 152.079
R7325 gnd.n3852 gnd.n3851 152.079
R7326 gnd.n1173 gnd.n1172 152
R7327 gnd.n1174 gnd.n1163 152
R7328 gnd.n1176 gnd.n1175 152
R7329 gnd.n1178 gnd.n1161 152
R7330 gnd.n1180 gnd.n1179 152
R7331 gnd.n5472 gnd.n5456 152
R7332 gnd.n5464 gnd.n5457 152
R7333 gnd.n5463 gnd.n5462 152
R7334 gnd.n5461 gnd.n5458 152
R7335 gnd.n5459 gnd.t120 150.546
R7336 gnd.t63 gnd.n3894 147.661
R7337 gnd.t357 gnd.n3862 147.661
R7338 gnd.t38 gnd.n3830 147.661
R7339 gnd.t46 gnd.n3799 147.661
R7340 gnd.t55 gnd.n3767 147.661
R7341 gnd.t26 gnd.n3735 147.661
R7342 gnd.t41 gnd.n3703 147.661
R7343 gnd.t359 gnd.n3672 147.661
R7344 gnd.n1764 gnd.n1746 143.351
R7345 gnd.n1140 gnd.n1123 143.351
R7346 gnd.n6344 gnd.n1123 143.351
R7347 gnd.n1170 gnd.t179 130.484
R7348 gnd.n1179 gnd.t87 126.766
R7349 gnd.n1177 gnd.t138 126.766
R7350 gnd.n1163 gnd.t98 126.766
R7351 gnd.n1171 gnd.t123 126.766
R7352 gnd.n5460 gnd.t189 126.766
R7353 gnd.n5462 gnd.t135 126.766
R7354 gnd.n5471 gnd.t84 126.766
R7355 gnd.n5473 gnd.t160 126.766
R7356 gnd.n7068 gnd.n514 106.77
R7357 gnd.n7069 gnd.n7068 106.77
R7358 gnd.n7070 gnd.n7069 106.77
R7359 gnd.n7070 gnd.n508 106.77
R7360 gnd.n7078 gnd.n508 106.77
R7361 gnd.n7079 gnd.n7078 106.77
R7362 gnd.n7080 gnd.n7079 106.77
R7363 gnd.n7080 gnd.n502 106.77
R7364 gnd.n7088 gnd.n502 106.77
R7365 gnd.n7089 gnd.n7088 106.77
R7366 gnd.n7090 gnd.n7089 106.77
R7367 gnd.n7090 gnd.n496 106.77
R7368 gnd.n7098 gnd.n496 106.77
R7369 gnd.n7099 gnd.n7098 106.77
R7370 gnd.n7100 gnd.n7099 106.77
R7371 gnd.n7100 gnd.n490 106.77
R7372 gnd.n7108 gnd.n490 106.77
R7373 gnd.n7109 gnd.n7108 106.77
R7374 gnd.n7110 gnd.n7109 106.77
R7375 gnd.n7110 gnd.n484 106.77
R7376 gnd.n7118 gnd.n484 106.77
R7377 gnd.n7119 gnd.n7118 106.77
R7378 gnd.n7120 gnd.n7119 106.77
R7379 gnd.n7120 gnd.n478 106.77
R7380 gnd.n7128 gnd.n478 106.77
R7381 gnd.n7129 gnd.n7128 106.77
R7382 gnd.n7130 gnd.n7129 106.77
R7383 gnd.n7130 gnd.n472 106.77
R7384 gnd.n7138 gnd.n472 106.77
R7385 gnd.n7139 gnd.n7138 106.77
R7386 gnd.n7140 gnd.n7139 106.77
R7387 gnd.n7140 gnd.n466 106.77
R7388 gnd.n7148 gnd.n466 106.77
R7389 gnd.n7149 gnd.n7148 106.77
R7390 gnd.n7150 gnd.n7149 106.77
R7391 gnd.n7150 gnd.n460 106.77
R7392 gnd.n7158 gnd.n460 106.77
R7393 gnd.n7159 gnd.n7158 106.77
R7394 gnd.n7160 gnd.n7159 106.77
R7395 gnd.n7160 gnd.n454 106.77
R7396 gnd.n7168 gnd.n454 106.77
R7397 gnd.n7169 gnd.n7168 106.77
R7398 gnd.n7170 gnd.n7169 106.77
R7399 gnd.n7170 gnd.n448 106.77
R7400 gnd.n7178 gnd.n448 106.77
R7401 gnd.n7179 gnd.n7178 106.77
R7402 gnd.n7180 gnd.n7179 106.77
R7403 gnd.n7180 gnd.n442 106.77
R7404 gnd.n7188 gnd.n442 106.77
R7405 gnd.n7189 gnd.n7188 106.77
R7406 gnd.n7190 gnd.n7189 106.77
R7407 gnd.n7190 gnd.n436 106.77
R7408 gnd.n7198 gnd.n436 106.77
R7409 gnd.n7199 gnd.n7198 106.77
R7410 gnd.n7200 gnd.n7199 106.77
R7411 gnd.n7200 gnd.n430 106.77
R7412 gnd.n7208 gnd.n430 106.77
R7413 gnd.n7209 gnd.n7208 106.77
R7414 gnd.n7210 gnd.n7209 106.77
R7415 gnd.n7210 gnd.n424 106.77
R7416 gnd.n7218 gnd.n424 106.77
R7417 gnd.n7219 gnd.n7218 106.77
R7418 gnd.n7220 gnd.n7219 106.77
R7419 gnd.n7220 gnd.n418 106.77
R7420 gnd.n7228 gnd.n418 106.77
R7421 gnd.n7229 gnd.n7228 106.77
R7422 gnd.n7230 gnd.n7229 106.77
R7423 gnd.n7230 gnd.n412 106.77
R7424 gnd.n7238 gnd.n412 106.77
R7425 gnd.n7239 gnd.n7238 106.77
R7426 gnd.n7240 gnd.n7239 106.77
R7427 gnd.n7240 gnd.n406 106.77
R7428 gnd.n7248 gnd.n406 106.77
R7429 gnd.n7249 gnd.n7248 106.77
R7430 gnd.n7250 gnd.n7249 106.77
R7431 gnd.n7250 gnd.n400 106.77
R7432 gnd.n7258 gnd.n400 106.77
R7433 gnd.n7259 gnd.n7258 106.77
R7434 gnd.n7260 gnd.n7259 106.77
R7435 gnd.n7260 gnd.n394 106.77
R7436 gnd.n7270 gnd.n394 106.77
R7437 gnd.n7271 gnd.n7270 106.77
R7438 gnd.n7272 gnd.n7271 106.77
R7439 gnd.n3911 gnd.n3910 104.615
R7440 gnd.n3910 gnd.n3888 104.615
R7441 gnd.n3903 gnd.n3888 104.615
R7442 gnd.n3903 gnd.n3902 104.615
R7443 gnd.n3902 gnd.n3892 104.615
R7444 gnd.n3895 gnd.n3892 104.615
R7445 gnd.n3879 gnd.n3878 104.615
R7446 gnd.n3878 gnd.n3856 104.615
R7447 gnd.n3871 gnd.n3856 104.615
R7448 gnd.n3871 gnd.n3870 104.615
R7449 gnd.n3870 gnd.n3860 104.615
R7450 gnd.n3863 gnd.n3860 104.615
R7451 gnd.n3847 gnd.n3846 104.615
R7452 gnd.n3846 gnd.n3824 104.615
R7453 gnd.n3839 gnd.n3824 104.615
R7454 gnd.n3839 gnd.n3838 104.615
R7455 gnd.n3838 gnd.n3828 104.615
R7456 gnd.n3831 gnd.n3828 104.615
R7457 gnd.n3816 gnd.n3815 104.615
R7458 gnd.n3815 gnd.n3793 104.615
R7459 gnd.n3808 gnd.n3793 104.615
R7460 gnd.n3808 gnd.n3807 104.615
R7461 gnd.n3807 gnd.n3797 104.615
R7462 gnd.n3800 gnd.n3797 104.615
R7463 gnd.n3784 gnd.n3783 104.615
R7464 gnd.n3783 gnd.n3761 104.615
R7465 gnd.n3776 gnd.n3761 104.615
R7466 gnd.n3776 gnd.n3775 104.615
R7467 gnd.n3775 gnd.n3765 104.615
R7468 gnd.n3768 gnd.n3765 104.615
R7469 gnd.n3752 gnd.n3751 104.615
R7470 gnd.n3751 gnd.n3729 104.615
R7471 gnd.n3744 gnd.n3729 104.615
R7472 gnd.n3744 gnd.n3743 104.615
R7473 gnd.n3743 gnd.n3733 104.615
R7474 gnd.n3736 gnd.n3733 104.615
R7475 gnd.n3720 gnd.n3719 104.615
R7476 gnd.n3719 gnd.n3697 104.615
R7477 gnd.n3712 gnd.n3697 104.615
R7478 gnd.n3712 gnd.n3711 104.615
R7479 gnd.n3711 gnd.n3701 104.615
R7480 gnd.n3704 gnd.n3701 104.615
R7481 gnd.n3689 gnd.n3688 104.615
R7482 gnd.n3688 gnd.n3666 104.615
R7483 gnd.n3681 gnd.n3666 104.615
R7484 gnd.n3681 gnd.n3680 104.615
R7485 gnd.n3680 gnd.n3670 104.615
R7486 gnd.n3673 gnd.n3670 104.615
R7487 gnd.n3062 gnd.t111 100.632
R7488 gnd.n2604 gnd.t146 100.632
R7489 gnd.n7529 gnd.n219 99.6594
R7490 gnd.n7527 gnd.n7526 99.6594
R7491 gnd.n7522 gnd.n226 99.6594
R7492 gnd.n7520 gnd.n7519 99.6594
R7493 gnd.n7515 gnd.n233 99.6594
R7494 gnd.n7513 gnd.n7512 99.6594
R7495 gnd.n7508 gnd.n240 99.6594
R7496 gnd.n7506 gnd.n7505 99.6594
R7497 gnd.n7498 gnd.n247 99.6594
R7498 gnd.n7496 gnd.n7495 99.6594
R7499 gnd.n7491 gnd.n254 99.6594
R7500 gnd.n7489 gnd.n7488 99.6594
R7501 gnd.n7484 gnd.n261 99.6594
R7502 gnd.n7482 gnd.n7481 99.6594
R7503 gnd.n7477 gnd.n268 99.6594
R7504 gnd.n7475 gnd.n7474 99.6594
R7505 gnd.n7470 gnd.n275 99.6594
R7506 gnd.n7468 gnd.n7467 99.6594
R7507 gnd.n285 gnd.n284 99.6594
R7508 gnd.n7459 gnd.n7458 99.6594
R7509 gnd.n7456 gnd.n7455 99.6594
R7510 gnd.n7451 gnd.n293 99.6594
R7511 gnd.n7449 gnd.n7448 99.6594
R7512 gnd.n7444 gnd.n300 99.6594
R7513 gnd.n7442 gnd.n7441 99.6594
R7514 gnd.n7437 gnd.n307 99.6594
R7515 gnd.n7435 gnd.n7434 99.6594
R7516 gnd.n7430 gnd.n316 99.6594
R7517 gnd.n7428 gnd.n7427 99.6594
R7518 gnd.n6080 gnd.n6079 99.6594
R7519 gnd.n6074 gnd.n1364 99.6594
R7520 gnd.n6071 gnd.n1365 99.6594
R7521 gnd.n6067 gnd.n1366 99.6594
R7522 gnd.n6063 gnd.n1367 99.6594
R7523 gnd.n6059 gnd.n1368 99.6594
R7524 gnd.n6055 gnd.n1369 99.6594
R7525 gnd.n6051 gnd.n1370 99.6594
R7526 gnd.n6047 gnd.n1371 99.6594
R7527 gnd.n6042 gnd.n1372 99.6594
R7528 gnd.n6038 gnd.n1373 99.6594
R7529 gnd.n6034 gnd.n1374 99.6594
R7530 gnd.n6030 gnd.n1375 99.6594
R7531 gnd.n6025 gnd.n1377 99.6594
R7532 gnd.n6021 gnd.n1378 99.6594
R7533 gnd.n6017 gnd.n1379 99.6594
R7534 gnd.n6013 gnd.n1380 99.6594
R7535 gnd.n6009 gnd.n1381 99.6594
R7536 gnd.n6005 gnd.n1382 99.6594
R7537 gnd.n6001 gnd.n1383 99.6594
R7538 gnd.n5997 gnd.n1384 99.6594
R7539 gnd.n5993 gnd.n1385 99.6594
R7540 gnd.n5989 gnd.n1386 99.6594
R7541 gnd.n5985 gnd.n1387 99.6594
R7542 gnd.n5981 gnd.n1388 99.6594
R7543 gnd.n5977 gnd.n1389 99.6594
R7544 gnd.n5973 gnd.n1390 99.6594
R7545 gnd.n5969 gnd.n1391 99.6594
R7546 gnd.n6390 gnd.n6389 99.6594
R7547 gnd.n6387 gnd.n6386 99.6594
R7548 gnd.n6382 gnd.n1082 99.6594
R7549 gnd.n6380 gnd.n6379 99.6594
R7550 gnd.n6375 gnd.n1089 99.6594
R7551 gnd.n6373 gnd.n6372 99.6594
R7552 gnd.n6368 gnd.n1096 99.6594
R7553 gnd.n6366 gnd.n6365 99.6594
R7554 gnd.n6360 gnd.n1105 99.6594
R7555 gnd.n6358 gnd.n6357 99.6594
R7556 gnd.n6353 gnd.n1112 99.6594
R7557 gnd.n6351 gnd.n6350 99.6594
R7558 gnd.n2229 gnd.n2228 99.6594
R7559 gnd.n2233 gnd.n2231 99.6594
R7560 gnd.n2239 gnd.n2223 99.6594
R7561 gnd.n2243 gnd.n2241 99.6594
R7562 gnd.n2249 gnd.n2219 99.6594
R7563 gnd.n2253 gnd.n2251 99.6594
R7564 gnd.n2259 gnd.n2213 99.6594
R7565 gnd.n2263 gnd.n2261 99.6594
R7566 gnd.n2269 gnd.n2209 99.6594
R7567 gnd.n2273 gnd.n2271 99.6594
R7568 gnd.n2279 gnd.n2205 99.6594
R7569 gnd.n2283 gnd.n2281 99.6594
R7570 gnd.n2289 gnd.n2201 99.6594
R7571 gnd.n2293 gnd.n2291 99.6594
R7572 gnd.n2299 gnd.n2197 99.6594
R7573 gnd.n2302 gnd.n2301 99.6594
R7574 gnd.n4356 gnd.n4355 99.6594
R7575 gnd.n4350 gnd.n4044 99.6594
R7576 gnd.n4347 gnd.n4045 99.6594
R7577 gnd.n4343 gnd.n4046 99.6594
R7578 gnd.n4339 gnd.n4047 99.6594
R7579 gnd.n4335 gnd.n4048 99.6594
R7580 gnd.n4331 gnd.n4049 99.6594
R7581 gnd.n4327 gnd.n4050 99.6594
R7582 gnd.n4323 gnd.n4051 99.6594
R7583 gnd.n4318 gnd.n4052 99.6594
R7584 gnd.n4314 gnd.n4053 99.6594
R7585 gnd.n4310 gnd.n4054 99.6594
R7586 gnd.n4306 gnd.n4055 99.6594
R7587 gnd.n4302 gnd.n4056 99.6594
R7588 gnd.n4298 gnd.n4057 99.6594
R7589 gnd.n4294 gnd.n4058 99.6594
R7590 gnd.n4290 gnd.n4059 99.6594
R7591 gnd.n4286 gnd.n4060 99.6594
R7592 gnd.n4282 gnd.n4061 99.6594
R7593 gnd.n4278 gnd.n4062 99.6594
R7594 gnd.n4274 gnd.n4063 99.6594
R7595 gnd.n4270 gnd.n4064 99.6594
R7596 gnd.n4266 gnd.n4065 99.6594
R7597 gnd.n4262 gnd.n4066 99.6594
R7598 gnd.n4258 gnd.n4067 99.6594
R7599 gnd.n4254 gnd.n4068 99.6594
R7600 gnd.n4250 gnd.n4069 99.6594
R7601 gnd.n4246 gnd.n4070 99.6594
R7602 gnd.n4358 gnd.n2564 99.6594
R7603 gnd.n4034 gnd.n2587 99.6594
R7604 gnd.n4032 gnd.n2586 99.6594
R7605 gnd.n4028 gnd.n2585 99.6594
R7606 gnd.n4024 gnd.n2584 99.6594
R7607 gnd.n4020 gnd.n2583 99.6594
R7608 gnd.n4016 gnd.n2582 99.6594
R7609 gnd.n4012 gnd.n2581 99.6594
R7610 gnd.n3944 gnd.n2580 99.6594
R7611 gnd.n3274 gnd.n3005 99.6594
R7612 gnd.n3031 gnd.n3012 99.6594
R7613 gnd.n3033 gnd.n3013 99.6594
R7614 gnd.n3041 gnd.n3014 99.6594
R7615 gnd.n3043 gnd.n3015 99.6594
R7616 gnd.n3051 gnd.n3016 99.6594
R7617 gnd.n3053 gnd.n3017 99.6594
R7618 gnd.n3061 gnd.n3018 99.6594
R7619 gnd.n7419 gnd.n322 99.6594
R7620 gnd.n7417 gnd.n7416 99.6594
R7621 gnd.n7412 gnd.n329 99.6594
R7622 gnd.n7410 gnd.n7409 99.6594
R7623 gnd.n7405 gnd.n336 99.6594
R7624 gnd.n7403 gnd.n7402 99.6594
R7625 gnd.n7398 gnd.n343 99.6594
R7626 gnd.n7396 gnd.n7395 99.6594
R7627 gnd.n348 gnd.n347 99.6594
R7628 gnd.n1476 gnd.n1392 99.6594
R7629 gnd.n1394 gnd.n1318 99.6594
R7630 gnd.n1395 gnd.n1325 99.6594
R7631 gnd.n1397 gnd.n1396 99.6594
R7632 gnd.n1399 gnd.n1334 99.6594
R7633 gnd.n1400 gnd.n1341 99.6594
R7634 gnd.n1402 gnd.n1401 99.6594
R7635 gnd.n1404 gnd.n1350 99.6594
R7636 gnd.n6082 gnd.n1359 99.6594
R7637 gnd.n4002 gnd.n2567 99.6594
R7638 gnd.n3998 gnd.n2568 99.6594
R7639 gnd.n3994 gnd.n2569 99.6594
R7640 gnd.n3990 gnd.n2570 99.6594
R7641 gnd.n3986 gnd.n2571 99.6594
R7642 gnd.n3982 gnd.n2572 99.6594
R7643 gnd.n3978 gnd.n2573 99.6594
R7644 gnd.n3974 gnd.n2574 99.6594
R7645 gnd.n3970 gnd.n2575 99.6594
R7646 gnd.n3966 gnd.n2576 99.6594
R7647 gnd.n3962 gnd.n2577 99.6594
R7648 gnd.n3958 gnd.n2578 99.6594
R7649 gnd.n3954 gnd.n2579 99.6594
R7650 gnd.n3189 gnd.n3188 99.6594
R7651 gnd.n3183 gnd.n3100 99.6594
R7652 gnd.n3180 gnd.n3101 99.6594
R7653 gnd.n3176 gnd.n3102 99.6594
R7654 gnd.n3172 gnd.n3103 99.6594
R7655 gnd.n3168 gnd.n3104 99.6594
R7656 gnd.n3164 gnd.n3105 99.6594
R7657 gnd.n3160 gnd.n3106 99.6594
R7658 gnd.n3156 gnd.n3107 99.6594
R7659 gnd.n3152 gnd.n3108 99.6594
R7660 gnd.n3148 gnd.n3109 99.6594
R7661 gnd.n3144 gnd.n3110 99.6594
R7662 gnd.n3191 gnd.n3099 99.6594
R7663 gnd.n2317 gnd.n2316 99.6594
R7664 gnd.n2328 gnd.n2327 99.6594
R7665 gnd.n2337 gnd.n2336 99.6594
R7666 gnd.n2340 gnd.n2339 99.6594
R7667 gnd.n2351 gnd.n2350 99.6594
R7668 gnd.n2360 gnd.n2359 99.6594
R7669 gnd.n2363 gnd.n2362 99.6594
R7670 gnd.n2375 gnd.n2374 99.6594
R7671 gnd.n4710 gnd.n4709 99.6594
R7672 gnd.n4236 gnd.n4071 99.6594
R7673 gnd.n4233 gnd.n4072 99.6594
R7674 gnd.n4229 gnd.n4073 99.6594
R7675 gnd.n4225 gnd.n4074 99.6594
R7676 gnd.n4221 gnd.n4075 99.6594
R7677 gnd.n4217 gnd.n4076 99.6594
R7678 gnd.n4213 gnd.n4077 99.6594
R7679 gnd.n4209 gnd.n4078 99.6594
R7680 gnd.n4205 gnd.n4079 99.6594
R7681 gnd.n4234 gnd.n4071 99.6594
R7682 gnd.n4230 gnd.n4072 99.6594
R7683 gnd.n4226 gnd.n4073 99.6594
R7684 gnd.n4222 gnd.n4074 99.6594
R7685 gnd.n4218 gnd.n4075 99.6594
R7686 gnd.n4214 gnd.n4076 99.6594
R7687 gnd.n4210 gnd.n4077 99.6594
R7688 gnd.n4206 gnd.n4078 99.6594
R7689 gnd.n4161 gnd.n4079 99.6594
R7690 gnd.n4709 gnd.n2379 99.6594
R7691 gnd.n2374 gnd.n2373 99.6594
R7692 gnd.n2362 gnd.n2361 99.6594
R7693 gnd.n2359 gnd.n2352 99.6594
R7694 gnd.n2350 gnd.n2349 99.6594
R7695 gnd.n2339 gnd.n2338 99.6594
R7696 gnd.n2336 gnd.n2329 99.6594
R7697 gnd.n2327 gnd.n2326 99.6594
R7698 gnd.n2316 gnd.n2315 99.6594
R7699 gnd.n3189 gnd.n3112 99.6594
R7700 gnd.n3181 gnd.n3100 99.6594
R7701 gnd.n3177 gnd.n3101 99.6594
R7702 gnd.n3173 gnd.n3102 99.6594
R7703 gnd.n3169 gnd.n3103 99.6594
R7704 gnd.n3165 gnd.n3104 99.6594
R7705 gnd.n3161 gnd.n3105 99.6594
R7706 gnd.n3157 gnd.n3106 99.6594
R7707 gnd.n3153 gnd.n3107 99.6594
R7708 gnd.n3149 gnd.n3108 99.6594
R7709 gnd.n3145 gnd.n3109 99.6594
R7710 gnd.n3141 gnd.n3110 99.6594
R7711 gnd.n3192 gnd.n3191 99.6594
R7712 gnd.n3957 gnd.n2579 99.6594
R7713 gnd.n3961 gnd.n2578 99.6594
R7714 gnd.n3965 gnd.n2577 99.6594
R7715 gnd.n3969 gnd.n2576 99.6594
R7716 gnd.n3973 gnd.n2575 99.6594
R7717 gnd.n3977 gnd.n2574 99.6594
R7718 gnd.n3981 gnd.n2573 99.6594
R7719 gnd.n3985 gnd.n2572 99.6594
R7720 gnd.n3989 gnd.n2571 99.6594
R7721 gnd.n3993 gnd.n2570 99.6594
R7722 gnd.n3997 gnd.n2569 99.6594
R7723 gnd.n4001 gnd.n2568 99.6594
R7724 gnd.n2608 gnd.n2567 99.6594
R7725 gnd.n1392 gnd.n1317 99.6594
R7726 gnd.n1394 gnd.n1393 99.6594
R7727 gnd.n1395 gnd.n1326 99.6594
R7728 gnd.n1397 gnd.n1333 99.6594
R7729 gnd.n1399 gnd.n1398 99.6594
R7730 gnd.n1400 gnd.n1342 99.6594
R7731 gnd.n1402 gnd.n1349 99.6594
R7732 gnd.n1404 gnd.n1403 99.6594
R7733 gnd.n6083 gnd.n6082 99.6594
R7734 gnd.n347 gnd.n344 99.6594
R7735 gnd.n7397 gnd.n7396 99.6594
R7736 gnd.n343 gnd.n337 99.6594
R7737 gnd.n7404 gnd.n7403 99.6594
R7738 gnd.n336 gnd.n330 99.6594
R7739 gnd.n7411 gnd.n7410 99.6594
R7740 gnd.n329 gnd.n323 99.6594
R7741 gnd.n7418 gnd.n7417 99.6594
R7742 gnd.n322 gnd.n319 99.6594
R7743 gnd.n3275 gnd.n3274 99.6594
R7744 gnd.n3034 gnd.n3012 99.6594
R7745 gnd.n3040 gnd.n3013 99.6594
R7746 gnd.n3044 gnd.n3014 99.6594
R7747 gnd.n3050 gnd.n3015 99.6594
R7748 gnd.n3054 gnd.n3016 99.6594
R7749 gnd.n3060 gnd.n3017 99.6594
R7750 gnd.n3018 gnd.n3002 99.6594
R7751 gnd.n4011 gnd.n2580 99.6594
R7752 gnd.n4015 gnd.n2581 99.6594
R7753 gnd.n4019 gnd.n2582 99.6594
R7754 gnd.n4023 gnd.n2583 99.6594
R7755 gnd.n4027 gnd.n2584 99.6594
R7756 gnd.n4031 gnd.n2585 99.6594
R7757 gnd.n4035 gnd.n2586 99.6594
R7758 gnd.n2589 gnd.n2587 99.6594
R7759 gnd.n4356 gnd.n4082 99.6594
R7760 gnd.n4348 gnd.n4044 99.6594
R7761 gnd.n4344 gnd.n4045 99.6594
R7762 gnd.n4340 gnd.n4046 99.6594
R7763 gnd.n4336 gnd.n4047 99.6594
R7764 gnd.n4332 gnd.n4048 99.6594
R7765 gnd.n4328 gnd.n4049 99.6594
R7766 gnd.n4324 gnd.n4050 99.6594
R7767 gnd.n4319 gnd.n4051 99.6594
R7768 gnd.n4315 gnd.n4052 99.6594
R7769 gnd.n4311 gnd.n4053 99.6594
R7770 gnd.n4307 gnd.n4054 99.6594
R7771 gnd.n4303 gnd.n4055 99.6594
R7772 gnd.n4299 gnd.n4056 99.6594
R7773 gnd.n4295 gnd.n4057 99.6594
R7774 gnd.n4291 gnd.n4058 99.6594
R7775 gnd.n4287 gnd.n4059 99.6594
R7776 gnd.n4283 gnd.n4060 99.6594
R7777 gnd.n4279 gnd.n4061 99.6594
R7778 gnd.n4275 gnd.n4062 99.6594
R7779 gnd.n4271 gnd.n4063 99.6594
R7780 gnd.n4267 gnd.n4064 99.6594
R7781 gnd.n4263 gnd.n4065 99.6594
R7782 gnd.n4259 gnd.n4066 99.6594
R7783 gnd.n4255 gnd.n4067 99.6594
R7784 gnd.n4251 gnd.n4068 99.6594
R7785 gnd.n4247 gnd.n4069 99.6594
R7786 gnd.n4243 gnd.n4070 99.6594
R7787 gnd.n4359 gnd.n4358 99.6594
R7788 gnd.n2301 gnd.n2300 99.6594
R7789 gnd.n2292 gnd.n2197 99.6594
R7790 gnd.n2291 gnd.n2290 99.6594
R7791 gnd.n2282 gnd.n2201 99.6594
R7792 gnd.n2281 gnd.n2280 99.6594
R7793 gnd.n2272 gnd.n2205 99.6594
R7794 gnd.n2271 gnd.n2270 99.6594
R7795 gnd.n2262 gnd.n2209 99.6594
R7796 gnd.n2261 gnd.n2260 99.6594
R7797 gnd.n2252 gnd.n2213 99.6594
R7798 gnd.n2251 gnd.n2250 99.6594
R7799 gnd.n2242 gnd.n2219 99.6594
R7800 gnd.n2241 gnd.n2240 99.6594
R7801 gnd.n2232 gnd.n2223 99.6594
R7802 gnd.n2231 gnd.n2230 99.6594
R7803 gnd.n1118 gnd.n1113 99.6594
R7804 gnd.n6352 gnd.n6351 99.6594
R7805 gnd.n1112 gnd.n1106 99.6594
R7806 gnd.n6359 gnd.n6358 99.6594
R7807 gnd.n1105 gnd.n1097 99.6594
R7808 gnd.n6367 gnd.n6366 99.6594
R7809 gnd.n1096 gnd.n1090 99.6594
R7810 gnd.n6374 gnd.n6373 99.6594
R7811 gnd.n1089 gnd.n1083 99.6594
R7812 gnd.n6381 gnd.n6380 99.6594
R7813 gnd.n1082 gnd.n1075 99.6594
R7814 gnd.n6388 gnd.n6387 99.6594
R7815 gnd.n6391 gnd.n6390 99.6594
R7816 gnd.n6080 gnd.n1407 99.6594
R7817 gnd.n6072 gnd.n1364 99.6594
R7818 gnd.n6068 gnd.n1365 99.6594
R7819 gnd.n6064 gnd.n1366 99.6594
R7820 gnd.n6060 gnd.n1367 99.6594
R7821 gnd.n6056 gnd.n1368 99.6594
R7822 gnd.n6052 gnd.n1369 99.6594
R7823 gnd.n6048 gnd.n1370 99.6594
R7824 gnd.n6043 gnd.n1371 99.6594
R7825 gnd.n6039 gnd.n1372 99.6594
R7826 gnd.n6035 gnd.n1373 99.6594
R7827 gnd.n6031 gnd.n1374 99.6594
R7828 gnd.n6026 gnd.n1376 99.6594
R7829 gnd.n6022 gnd.n1377 99.6594
R7830 gnd.n6018 gnd.n1378 99.6594
R7831 gnd.n6014 gnd.n1379 99.6594
R7832 gnd.n6010 gnd.n1380 99.6594
R7833 gnd.n6006 gnd.n1381 99.6594
R7834 gnd.n6002 gnd.n1382 99.6594
R7835 gnd.n5998 gnd.n1383 99.6594
R7836 gnd.n5994 gnd.n1384 99.6594
R7837 gnd.n5990 gnd.n1385 99.6594
R7838 gnd.n5986 gnd.n1386 99.6594
R7839 gnd.n5982 gnd.n1387 99.6594
R7840 gnd.n5978 gnd.n1388 99.6594
R7841 gnd.n5974 gnd.n1389 99.6594
R7842 gnd.n5970 gnd.n1390 99.6594
R7843 gnd.n5962 gnd.n1391 99.6594
R7844 gnd.n7429 gnd.n7428 99.6594
R7845 gnd.n316 gnd.n308 99.6594
R7846 gnd.n7436 gnd.n7435 99.6594
R7847 gnd.n307 gnd.n301 99.6594
R7848 gnd.n7443 gnd.n7442 99.6594
R7849 gnd.n300 gnd.n294 99.6594
R7850 gnd.n7450 gnd.n7449 99.6594
R7851 gnd.n293 gnd.n287 99.6594
R7852 gnd.n7457 gnd.n7456 99.6594
R7853 gnd.n7460 gnd.n7459 99.6594
R7854 gnd.n284 gnd.n276 99.6594
R7855 gnd.n7469 gnd.n7468 99.6594
R7856 gnd.n275 gnd.n269 99.6594
R7857 gnd.n7476 gnd.n7475 99.6594
R7858 gnd.n268 gnd.n262 99.6594
R7859 gnd.n7483 gnd.n7482 99.6594
R7860 gnd.n261 gnd.n255 99.6594
R7861 gnd.n7490 gnd.n7489 99.6594
R7862 gnd.n254 gnd.n248 99.6594
R7863 gnd.n7497 gnd.n7496 99.6594
R7864 gnd.n247 gnd.n241 99.6594
R7865 gnd.n7507 gnd.n7506 99.6594
R7866 gnd.n240 gnd.n234 99.6594
R7867 gnd.n7514 gnd.n7513 99.6594
R7868 gnd.n233 gnd.n227 99.6594
R7869 gnd.n7521 gnd.n7520 99.6594
R7870 gnd.n226 gnd.n220 99.6594
R7871 gnd.n7528 gnd.n7527 99.6594
R7872 gnd.n219 gnd.n216 99.6594
R7873 gnd.n4772 gnd.n4771 99.6594
R7874 gnd.n2189 gnd.n2121 99.6594
R7875 gnd.n2191 gnd.n2122 99.6594
R7876 gnd.n2308 gnd.n2123 99.6594
R7877 gnd.n2310 gnd.n2124 99.6594
R7878 gnd.n2321 gnd.n2125 99.6594
R7879 gnd.n2323 gnd.n2126 99.6594
R7880 gnd.n2333 gnd.n2127 99.6594
R7881 gnd.n2344 gnd.n2128 99.6594
R7882 gnd.n2346 gnd.n2129 99.6594
R7883 gnd.n2356 gnd.n2130 99.6594
R7884 gnd.n2367 gnd.n2131 99.6594
R7885 gnd.n4700 gnd.n2132 99.6594
R7886 gnd.n4704 gnd.n2133 99.6594
R7887 gnd.n4772 gnd.n2135 99.6594
R7888 gnd.n2190 gnd.n2121 99.6594
R7889 gnd.n2307 gnd.n2122 99.6594
R7890 gnd.n2309 gnd.n2123 99.6594
R7891 gnd.n2320 gnd.n2124 99.6594
R7892 gnd.n2322 gnd.n2125 99.6594
R7893 gnd.n2332 gnd.n2126 99.6594
R7894 gnd.n2343 gnd.n2127 99.6594
R7895 gnd.n2345 gnd.n2128 99.6594
R7896 gnd.n2355 gnd.n2129 99.6594
R7897 gnd.n2366 gnd.n2130 99.6594
R7898 gnd.n2368 gnd.n2131 99.6594
R7899 gnd.n4703 gnd.n2132 99.6594
R7900 gnd.n2133 gnd.n2111 99.6594
R7901 gnd.n1640 gnd.n1302 99.6594
R7902 gnd.n1642 gnd.n1641 99.6594
R7903 gnd.n1643 gnd.n1307 99.6594
R7904 gnd.n1645 gnd.n1644 99.6594
R7905 gnd.n1646 gnd.n1313 99.6594
R7906 gnd.n1648 gnd.n1321 99.6594
R7907 gnd.n1650 gnd.n1649 99.6594
R7908 gnd.n1651 gnd.n1330 99.6594
R7909 gnd.n1653 gnd.n1337 99.6594
R7910 gnd.n1655 gnd.n1654 99.6594
R7911 gnd.n1656 gnd.n1346 99.6594
R7912 gnd.n1658 gnd.n1353 99.6594
R7913 gnd.n1661 gnd.n1660 99.6594
R7914 gnd.n5730 gnd.n5729 99.6594
R7915 gnd.n1658 gnd.n1657 99.6594
R7916 gnd.n1656 gnd.n1345 99.6594
R7917 gnd.n1655 gnd.n1338 99.6594
R7918 gnd.n1653 gnd.n1652 99.6594
R7919 gnd.n1651 gnd.n1329 99.6594
R7920 gnd.n1650 gnd.n1322 99.6594
R7921 gnd.n1648 gnd.n1647 99.6594
R7922 gnd.n1646 gnd.n1312 99.6594
R7923 gnd.n1645 gnd.n1308 99.6594
R7924 gnd.n1643 gnd.n1306 99.6594
R7925 gnd.n1642 gnd.n1303 99.6594
R7926 gnd.n1640 gnd.n1298 99.6594
R7927 gnd.n5729 gnd.n1293 99.6594
R7928 gnd.n1661 gnd.n1639 99.6594
R7929 gnd.n2369 gnd.t119 98.63
R7930 gnd.n6084 gnd.t79 98.63
R7931 gnd.n2376 gnd.t114 98.63
R7932 gnd.n1427 gnd.t175 98.63
R7933 gnd.n1450 gnd.t178 98.63
R7934 gnd.n5964 gnd.t128 98.63
R7935 gnd.n313 gnd.t155 98.63
R7936 gnd.n280 gnd.t106 98.63
R7937 gnd.n7500 gnd.t149 98.63
R7938 gnd.n350 gnd.t96 98.63
R7939 gnd.n4101 gnd.t131 98.63
R7940 gnd.n4123 gnd.t134 98.63
R7941 gnd.n4144 gnd.t83 98.63
R7942 gnd.n4162 gnd.t165 98.63
R7943 gnd.n1101 gnd.t142 98.63
R7944 gnd.n2194 gnd.t167 98.63
R7945 gnd.n2216 gnd.t187 98.63
R7946 gnd.n1355 gnd.t92 98.63
R7947 gnd.n4896 gnd.t153 96.6984
R7948 gnd.n1765 gnd.t103 96.6984
R7949 gnd.n6278 gnd.t75 96.6906
R7950 gnd.n5475 gnd.t158 96.6906
R7951 gnd.n1170 gnd.n1169 81.8399
R7952 gnd.n3063 gnd.t110 74.8376
R7953 gnd.n2605 gnd.t147 74.8376
R7954 gnd.n4897 gnd.t152 72.8438
R7955 gnd.n1766 gnd.t104 72.8438
R7956 gnd.n1171 gnd.n1164 72.8411
R7957 gnd.n1177 gnd.n1162 72.8411
R7958 gnd.n5471 gnd.n5470 72.8411
R7959 gnd.n2370 gnd.t118 72.836
R7960 gnd.n6279 gnd.t74 72.836
R7961 gnd.n5476 gnd.t159 72.836
R7962 gnd.n6085 gnd.t78 72.836
R7963 gnd.n2377 gnd.t115 72.836
R7964 gnd.n1428 gnd.t174 72.836
R7965 gnd.n1451 gnd.t177 72.836
R7966 gnd.n5965 gnd.t127 72.836
R7967 gnd.n314 gnd.t156 72.836
R7968 gnd.n281 gnd.t107 72.836
R7969 gnd.n7501 gnd.t150 72.836
R7970 gnd.n351 gnd.t97 72.836
R7971 gnd.n4102 gnd.t130 72.836
R7972 gnd.n4124 gnd.t133 72.836
R7973 gnd.n4145 gnd.t82 72.836
R7974 gnd.n4163 gnd.t164 72.836
R7975 gnd.n1102 gnd.t143 72.836
R7976 gnd.n2195 gnd.t168 72.836
R7977 gnd.n2217 gnd.t188 72.836
R7978 gnd.n1356 gnd.t93 72.836
R7979 gnd.n5539 gnd.n1730 71.676
R7980 gnd.n5535 gnd.n1731 71.676
R7981 gnd.n5531 gnd.n1732 71.676
R7982 gnd.n5527 gnd.n1733 71.676
R7983 gnd.n5523 gnd.n1734 71.676
R7984 gnd.n5519 gnd.n1735 71.676
R7985 gnd.n5515 gnd.n1736 71.676
R7986 gnd.n5511 gnd.n1737 71.676
R7987 gnd.n5507 gnd.n1738 71.676
R7988 gnd.n5503 gnd.n1739 71.676
R7989 gnd.n5499 gnd.n1740 71.676
R7990 gnd.n5495 gnd.n1741 71.676
R7991 gnd.n5491 gnd.n1742 71.676
R7992 gnd.n5487 gnd.n1743 71.676
R7993 gnd.n5482 gnd.n1744 71.676
R7994 gnd.n5478 gnd.n1745 71.676
R7995 gnd.n5615 gnd.n1764 71.676
R7996 gnd.n5611 gnd.n1763 71.676
R7997 gnd.n5606 gnd.n1762 71.676
R7998 gnd.n5602 gnd.n1761 71.676
R7999 gnd.n5598 gnd.n1760 71.676
R8000 gnd.n5594 gnd.n1759 71.676
R8001 gnd.n5590 gnd.n1758 71.676
R8002 gnd.n5586 gnd.n1757 71.676
R8003 gnd.n5582 gnd.n1756 71.676
R8004 gnd.n5578 gnd.n1755 71.676
R8005 gnd.n5574 gnd.n1754 71.676
R8006 gnd.n5570 gnd.n1753 71.676
R8007 gnd.n5566 gnd.n1752 71.676
R8008 gnd.n5562 gnd.n1751 71.676
R8009 gnd.n5558 gnd.n1750 71.676
R8010 gnd.n5554 gnd.n1749 71.676
R8011 gnd.n5550 gnd.n1748 71.676
R8012 gnd.n6342 gnd.n6341 71.676
R8013 gnd.n6336 gnd.n1126 71.676
R8014 gnd.n6333 gnd.n1127 71.676
R8015 gnd.n6329 gnd.n1128 71.676
R8016 gnd.n6325 gnd.n1129 71.676
R8017 gnd.n6321 gnd.n1130 71.676
R8018 gnd.n6317 gnd.n1131 71.676
R8019 gnd.n6313 gnd.n1132 71.676
R8020 gnd.n6309 gnd.n1133 71.676
R8021 gnd.n6305 gnd.n1134 71.676
R8022 gnd.n6301 gnd.n1135 71.676
R8023 gnd.n6297 gnd.n1136 71.676
R8024 gnd.n6293 gnd.n1137 71.676
R8025 gnd.n6289 gnd.n1138 71.676
R8026 gnd.n6285 gnd.n1139 71.676
R8027 gnd.n6281 gnd.n1140 71.676
R8028 gnd.n1141 gnd.n1124 71.676
R8029 gnd.n4900 gnd.n1142 71.676
R8030 gnd.n4905 gnd.n1143 71.676
R8031 gnd.n4909 gnd.n1144 71.676
R8032 gnd.n4913 gnd.n1145 71.676
R8033 gnd.n4917 gnd.n1146 71.676
R8034 gnd.n4921 gnd.n1147 71.676
R8035 gnd.n4925 gnd.n1148 71.676
R8036 gnd.n4929 gnd.n1149 71.676
R8037 gnd.n4933 gnd.n1150 71.676
R8038 gnd.n4937 gnd.n1151 71.676
R8039 gnd.n4941 gnd.n1152 71.676
R8040 gnd.n4945 gnd.n1153 71.676
R8041 gnd.n4949 gnd.n1154 71.676
R8042 gnd.n4953 gnd.n1155 71.676
R8043 gnd.n4957 gnd.n1156 71.676
R8044 gnd.n6342 gnd.n1159 71.676
R8045 gnd.n6334 gnd.n1126 71.676
R8046 gnd.n6330 gnd.n1127 71.676
R8047 gnd.n6326 gnd.n1128 71.676
R8048 gnd.n6322 gnd.n1129 71.676
R8049 gnd.n6318 gnd.n1130 71.676
R8050 gnd.n6314 gnd.n1131 71.676
R8051 gnd.n6310 gnd.n1132 71.676
R8052 gnd.n6306 gnd.n1133 71.676
R8053 gnd.n6302 gnd.n1134 71.676
R8054 gnd.n6298 gnd.n1135 71.676
R8055 gnd.n6294 gnd.n1136 71.676
R8056 gnd.n6290 gnd.n1137 71.676
R8057 gnd.n6286 gnd.n1138 71.676
R8058 gnd.n6282 gnd.n1139 71.676
R8059 gnd.n6345 gnd.n6344 71.676
R8060 gnd.n4899 gnd.n1141 71.676
R8061 gnd.n4904 gnd.n1142 71.676
R8062 gnd.n4908 gnd.n1143 71.676
R8063 gnd.n4912 gnd.n1144 71.676
R8064 gnd.n4916 gnd.n1145 71.676
R8065 gnd.n4920 gnd.n1146 71.676
R8066 gnd.n4924 gnd.n1147 71.676
R8067 gnd.n4928 gnd.n1148 71.676
R8068 gnd.n4932 gnd.n1149 71.676
R8069 gnd.n4936 gnd.n1150 71.676
R8070 gnd.n4940 gnd.n1151 71.676
R8071 gnd.n4944 gnd.n1152 71.676
R8072 gnd.n4948 gnd.n1153 71.676
R8073 gnd.n4952 gnd.n1154 71.676
R8074 gnd.n4956 gnd.n1155 71.676
R8075 gnd.n4960 gnd.n1156 71.676
R8076 gnd.n5553 gnd.n1748 71.676
R8077 gnd.n5557 gnd.n1749 71.676
R8078 gnd.n5561 gnd.n1750 71.676
R8079 gnd.n5565 gnd.n1751 71.676
R8080 gnd.n5569 gnd.n1752 71.676
R8081 gnd.n5573 gnd.n1753 71.676
R8082 gnd.n5577 gnd.n1754 71.676
R8083 gnd.n5581 gnd.n1755 71.676
R8084 gnd.n5585 gnd.n1756 71.676
R8085 gnd.n5589 gnd.n1757 71.676
R8086 gnd.n5593 gnd.n1758 71.676
R8087 gnd.n5597 gnd.n1759 71.676
R8088 gnd.n5601 gnd.n1760 71.676
R8089 gnd.n5605 gnd.n1761 71.676
R8090 gnd.n5610 gnd.n1762 71.676
R8091 gnd.n5614 gnd.n1763 71.676
R8092 gnd.n5477 gnd.n1746 71.676
R8093 gnd.n5481 gnd.n1745 71.676
R8094 gnd.n5486 gnd.n1744 71.676
R8095 gnd.n5490 gnd.n1743 71.676
R8096 gnd.n5494 gnd.n1742 71.676
R8097 gnd.n5498 gnd.n1741 71.676
R8098 gnd.n5502 gnd.n1740 71.676
R8099 gnd.n5506 gnd.n1739 71.676
R8100 gnd.n5510 gnd.n1738 71.676
R8101 gnd.n5514 gnd.n1737 71.676
R8102 gnd.n5518 gnd.n1736 71.676
R8103 gnd.n5522 gnd.n1735 71.676
R8104 gnd.n5526 gnd.n1734 71.676
R8105 gnd.n5530 gnd.n1733 71.676
R8106 gnd.n5534 gnd.n1732 71.676
R8107 gnd.n5538 gnd.n1731 71.676
R8108 gnd.n5541 gnd.n1730 71.676
R8109 gnd.n10 gnd.t361 69.1507
R8110 gnd.n18 gnd.t353 68.4792
R8111 gnd.n17 gnd.t44 68.4792
R8112 gnd.n16 gnd.t28 68.4792
R8113 gnd.n15 gnd.t367 68.4792
R8114 gnd.n14 gnd.t48 68.4792
R8115 gnd.n13 gnd.t365 68.4792
R8116 gnd.n12 gnd.t68 68.4792
R8117 gnd.n11 gnd.t60 68.4792
R8118 gnd.n10 gnd.t70 68.4792
R8119 gnd.n3190 gnd.n3094 64.369
R8120 gnd.n7272 gnd.n184 64.0626
R8121 gnd.n4902 gnd.n4897 59.5399
R8122 gnd.n5608 gnd.n1766 59.5399
R8123 gnd.n6280 gnd.n6279 59.5399
R8124 gnd.n5484 gnd.n5476 59.5399
R8125 gnd.n6277 gnd.n1180 59.1804
R8126 gnd.n4043 gnd.n2565 57.3586
R8127 gnd.n4357 gnd.n2552 57.3586
R8128 gnd.n7537 gnd.n212 57.3586
R8129 gnd.n2845 gnd.t317 56.407
R8130 gnd.n2798 gnd.t335 56.407
R8131 gnd.n2813 gnd.t298 56.407
R8132 gnd.n2829 gnd.t207 56.407
R8133 gnd.n68 gnd.t291 56.407
R8134 gnd.n21 gnd.t218 56.407
R8135 gnd.n36 gnd.t278 56.407
R8136 gnd.n52 gnd.t328 56.407
R8137 gnd.n2858 gnd.t270 55.8337
R8138 gnd.n2811 gnd.t226 55.8337
R8139 gnd.n2826 gnd.t247 55.8337
R8140 gnd.n2842 gnd.t306 55.8337
R8141 gnd.n81 gnd.t331 55.8337
R8142 gnd.n34 gnd.t241 55.8337
R8143 gnd.n49 gnd.t350 55.8337
R8144 gnd.n65 gnd.t245 55.8337
R8145 gnd.n1168 gnd.n1167 54.358
R8146 gnd.n5468 gnd.n5467 54.358
R8147 gnd.n2845 gnd.n2844 53.0052
R8148 gnd.n2847 gnd.n2846 53.0052
R8149 gnd.n2849 gnd.n2848 53.0052
R8150 gnd.n2851 gnd.n2850 53.0052
R8151 gnd.n2853 gnd.n2852 53.0052
R8152 gnd.n2855 gnd.n2854 53.0052
R8153 gnd.n2857 gnd.n2856 53.0052
R8154 gnd.n2798 gnd.n2797 53.0052
R8155 gnd.n2800 gnd.n2799 53.0052
R8156 gnd.n2802 gnd.n2801 53.0052
R8157 gnd.n2804 gnd.n2803 53.0052
R8158 gnd.n2806 gnd.n2805 53.0052
R8159 gnd.n2808 gnd.n2807 53.0052
R8160 gnd.n2810 gnd.n2809 53.0052
R8161 gnd.n2813 gnd.n2812 53.0052
R8162 gnd.n2815 gnd.n2814 53.0052
R8163 gnd.n2817 gnd.n2816 53.0052
R8164 gnd.n2819 gnd.n2818 53.0052
R8165 gnd.n2821 gnd.n2820 53.0052
R8166 gnd.n2823 gnd.n2822 53.0052
R8167 gnd.n2825 gnd.n2824 53.0052
R8168 gnd.n2829 gnd.n2828 53.0052
R8169 gnd.n2831 gnd.n2830 53.0052
R8170 gnd.n2833 gnd.n2832 53.0052
R8171 gnd.n2835 gnd.n2834 53.0052
R8172 gnd.n2837 gnd.n2836 53.0052
R8173 gnd.n2839 gnd.n2838 53.0052
R8174 gnd.n2841 gnd.n2840 53.0052
R8175 gnd.n80 gnd.n79 53.0052
R8176 gnd.n78 gnd.n77 53.0052
R8177 gnd.n76 gnd.n75 53.0052
R8178 gnd.n74 gnd.n73 53.0052
R8179 gnd.n72 gnd.n71 53.0052
R8180 gnd.n70 gnd.n69 53.0052
R8181 gnd.n68 gnd.n67 53.0052
R8182 gnd.n33 gnd.n32 53.0052
R8183 gnd.n31 gnd.n30 53.0052
R8184 gnd.n29 gnd.n28 53.0052
R8185 gnd.n27 gnd.n26 53.0052
R8186 gnd.n25 gnd.n24 53.0052
R8187 gnd.n23 gnd.n22 53.0052
R8188 gnd.n21 gnd.n20 53.0052
R8189 gnd.n48 gnd.n47 53.0052
R8190 gnd.n46 gnd.n45 53.0052
R8191 gnd.n44 gnd.n43 53.0052
R8192 gnd.n42 gnd.n41 53.0052
R8193 gnd.n40 gnd.n39 53.0052
R8194 gnd.n38 gnd.n37 53.0052
R8195 gnd.n36 gnd.n35 53.0052
R8196 gnd.n64 gnd.n63 53.0052
R8197 gnd.n62 gnd.n61 53.0052
R8198 gnd.n60 gnd.n59 53.0052
R8199 gnd.n58 gnd.n57 53.0052
R8200 gnd.n56 gnd.n55 53.0052
R8201 gnd.n54 gnd.n53 53.0052
R8202 gnd.n52 gnd.n51 53.0052
R8203 gnd.n5459 gnd.n5458 52.4801
R8204 gnd.n3895 gnd.t63 52.3082
R8205 gnd.n3863 gnd.t357 52.3082
R8206 gnd.n3831 gnd.t38 52.3082
R8207 gnd.n3800 gnd.t46 52.3082
R8208 gnd.n3768 gnd.t55 52.3082
R8209 gnd.n3736 gnd.t26 52.3082
R8210 gnd.n3704 gnd.t41 52.3082
R8211 gnd.n3673 gnd.t359 52.3082
R8212 gnd.n3725 gnd.n3693 51.4173
R8213 gnd.n3789 gnd.n3788 50.455
R8214 gnd.n3757 gnd.n3756 50.455
R8215 gnd.n3725 gnd.n3724 50.455
R8216 gnd.n3137 gnd.n3136 45.1884
R8217 gnd.n2631 gnd.n2630 45.1884
R8218 gnd.n5543 gnd.n5474 44.3322
R8219 gnd.n1171 gnd.n1170 44.3189
R8220 gnd.n2371 gnd.n2370 42.4732
R8221 gnd.n1357 gnd.n1356 42.4732
R8222 gnd.n6086 gnd.n6085 42.2793
R8223 gnd.n3138 gnd.n3137 42.2793
R8224 gnd.n2632 gnd.n2631 42.2793
R8225 gnd.n3064 gnd.n3063 42.2793
R8226 gnd.n4010 gnd.n2605 42.2793
R8227 gnd.n4712 gnd.n2377 42.2793
R8228 gnd.n6045 gnd.n1428 42.2793
R8229 gnd.n6008 gnd.n1451 42.2793
R8230 gnd.n5968 gnd.n5965 42.2793
R8231 gnd.n315 gnd.n314 42.2793
R8232 gnd.n7465 gnd.n281 42.2793
R8233 gnd.n7502 gnd.n7501 42.2793
R8234 gnd.n7393 gnd.n351 42.2793
R8235 gnd.n4321 gnd.n4102 42.2793
R8236 gnd.n4281 gnd.n4124 42.2793
R8237 gnd.n4242 gnd.n4145 42.2793
R8238 gnd.n4164 gnd.n4163 42.2793
R8239 gnd.n6362 gnd.n1102 42.2793
R8240 gnd.n2196 gnd.n2195 42.2793
R8241 gnd.n2218 gnd.n2217 42.2793
R8242 gnd.n1169 gnd.n1168 41.6274
R8243 gnd.n5469 gnd.n5468 41.6274
R8244 gnd.n1178 gnd.n1177 40.8975
R8245 gnd.n5472 gnd.n5471 40.8975
R8246 gnd.n1177 gnd.n1176 35.055
R8247 gnd.n1172 gnd.n1171 35.055
R8248 gnd.n5461 gnd.n5460 35.055
R8249 gnd.n5471 gnd.n5457 35.055
R8250 gnd.n6640 gnd.n6639 34.6789
R8251 gnd.n6639 gnd.n6638 34.6789
R8252 gnd.n6638 gnd.n772 34.6789
R8253 gnd.n6632 gnd.n772 34.6789
R8254 gnd.n6632 gnd.n6631 34.6789
R8255 gnd.n6631 gnd.n6630 34.6789
R8256 gnd.n6630 gnd.n779 34.6789
R8257 gnd.n6624 gnd.n779 34.6789
R8258 gnd.n6624 gnd.n6623 34.6789
R8259 gnd.n6623 gnd.n6622 34.6789
R8260 gnd.n6622 gnd.n787 34.6789
R8261 gnd.n6616 gnd.n787 34.6789
R8262 gnd.n6616 gnd.n6615 34.6789
R8263 gnd.n6615 gnd.n6614 34.6789
R8264 gnd.n6614 gnd.n795 34.6789
R8265 gnd.n6608 gnd.n795 34.6789
R8266 gnd.n6608 gnd.n6607 34.6789
R8267 gnd.n6607 gnd.n6606 34.6789
R8268 gnd.n6606 gnd.n803 34.6789
R8269 gnd.n6600 gnd.n803 34.6789
R8270 gnd.n6600 gnd.n6599 34.6789
R8271 gnd.n6599 gnd.n6598 34.6789
R8272 gnd.n6598 gnd.n811 34.6789
R8273 gnd.n6592 gnd.n811 34.6789
R8274 gnd.n6592 gnd.n6591 34.6789
R8275 gnd.n6591 gnd.n6590 34.6789
R8276 gnd.n6590 gnd.n819 34.6789
R8277 gnd.n6584 gnd.n819 34.6789
R8278 gnd.n6584 gnd.n6583 34.6789
R8279 gnd.n6583 gnd.n6582 34.6789
R8280 gnd.n6582 gnd.n827 34.6789
R8281 gnd.n6576 gnd.n827 34.6789
R8282 gnd.n6576 gnd.n6575 34.6789
R8283 gnd.n6575 gnd.n6574 34.6789
R8284 gnd.n6574 gnd.n835 34.6789
R8285 gnd.n6568 gnd.n835 34.6789
R8286 gnd.n6568 gnd.n6567 34.6789
R8287 gnd.n6567 gnd.n6566 34.6789
R8288 gnd.n6566 gnd.n843 34.6789
R8289 gnd.n6560 gnd.n843 34.6789
R8290 gnd.n6560 gnd.n6559 34.6789
R8291 gnd.n6559 gnd.n6558 34.6789
R8292 gnd.n6558 gnd.n851 34.6789
R8293 gnd.n6552 gnd.n851 34.6789
R8294 gnd.n6552 gnd.n6551 34.6789
R8295 gnd.n6551 gnd.n6550 34.6789
R8296 gnd.n6550 gnd.n859 34.6789
R8297 gnd.n6544 gnd.n859 34.6789
R8298 gnd.n6544 gnd.n6543 34.6789
R8299 gnd.n6543 gnd.n6542 34.6789
R8300 gnd.n6542 gnd.n867 34.6789
R8301 gnd.n6536 gnd.n867 34.6789
R8302 gnd.n6536 gnd.n6535 34.6789
R8303 gnd.n6535 gnd.n6534 34.6789
R8304 gnd.n6534 gnd.n875 34.6789
R8305 gnd.n6528 gnd.n875 34.6789
R8306 gnd.n6528 gnd.n6527 34.6789
R8307 gnd.n6527 gnd.n6526 34.6789
R8308 gnd.n6526 gnd.n883 34.6789
R8309 gnd.n6520 gnd.n883 34.6789
R8310 gnd.n6520 gnd.n6519 34.6789
R8311 gnd.n6519 gnd.n6518 34.6789
R8312 gnd.n6518 gnd.n891 34.6789
R8313 gnd.n6512 gnd.n891 34.6789
R8314 gnd.n6512 gnd.n6511 34.6789
R8315 gnd.n6511 gnd.n6510 34.6789
R8316 gnd.n6510 gnd.n899 34.6789
R8317 gnd.n6504 gnd.n899 34.6789
R8318 gnd.n6504 gnd.n6503 34.6789
R8319 gnd.n6503 gnd.n6502 34.6789
R8320 gnd.n6502 gnd.n907 34.6789
R8321 gnd.n6496 gnd.n907 34.6789
R8322 gnd.n6496 gnd.n6495 34.6789
R8323 gnd.n6495 gnd.n6494 34.6789
R8324 gnd.n6494 gnd.n915 34.6789
R8325 gnd.n6488 gnd.n915 34.6789
R8326 gnd.n6488 gnd.n6487 34.6789
R8327 gnd.n6487 gnd.n6486 34.6789
R8328 gnd.n6486 gnd.n923 34.6789
R8329 gnd.n6480 gnd.n923 34.6789
R8330 gnd.n6480 gnd.n6479 34.6789
R8331 gnd.n6479 gnd.n6478 34.6789
R8332 gnd.n6478 gnd.n931 34.6789
R8333 gnd.n5551 gnd.n1767 33.2493
R8334 gnd.n4963 gnd.n4959 33.2493
R8335 gnd.n3200 gnd.n3094 31.8661
R8336 gnd.n3200 gnd.n3199 31.8661
R8337 gnd.n3208 gnd.n3083 31.8661
R8338 gnd.n3216 gnd.n3083 31.8661
R8339 gnd.n3216 gnd.n3077 31.8661
R8340 gnd.n3224 gnd.n3077 31.8661
R8341 gnd.n3224 gnd.n3070 31.8661
R8342 gnd.n3262 gnd.n3070 31.8661
R8343 gnd.n3272 gnd.n3003 31.8661
R8344 gnd.n4367 gnd.n2552 31.8661
R8345 gnd.n4375 gnd.n2544 31.8661
R8346 gnd.n4375 gnd.n2533 31.8661
R8347 gnd.n4387 gnd.n2533 31.8661
R8348 gnd.n4387 gnd.n2536 31.8661
R8349 gnd.n4395 gnd.n2516 31.8661
R8350 gnd.n4407 gnd.n2516 31.8661
R8351 gnd.n4415 gnd.n2508 31.8661
R8352 gnd.n4431 gnd.n2496 31.8661
R8353 gnd.n4431 gnd.n2499 31.8661
R8354 gnd.n4441 gnd.n2482 31.8661
R8355 gnd.n4461 gnd.n2482 31.8661
R8356 gnd.n4472 gnd.n2474 31.8661
R8357 gnd.n4481 gnd.n2456 31.8661
R8358 gnd.n4497 gnd.n2456 31.8661
R8359 gnd.n4501 gnd.n938 31.8661
R8360 gnd.n4657 gnd.n1068 31.8661
R8361 gnd.n4650 gnd.n2120 31.8661
R8362 gnd.n4774 gnd.n2120 31.8661
R8363 gnd.n4782 gnd.n2112 31.8661
R8364 gnd.n4782 gnd.n2114 31.8661
R8365 gnd.n4790 gnd.n2100 31.8661
R8366 gnd.n4798 gnd.n2100 31.8661
R8367 gnd.n4798 gnd.n2093 31.8661
R8368 gnd.n4806 gnd.n2093 31.8661
R8369 gnd.n4814 gnd.n2086 31.8661
R8370 gnd.n4814 gnd.n2078 31.8661
R8371 gnd.n4822 gnd.n2078 31.8661
R8372 gnd.n4822 gnd.n2080 31.8661
R8373 gnd.n4830 gnd.n2064 31.8661
R8374 gnd.n4838 gnd.n2064 31.8661
R8375 gnd.n4838 gnd.n2066 31.8661
R8376 gnd.n4846 gnd.n2049 31.8661
R8377 gnd.n4868 gnd.n2049 31.8661
R8378 gnd.n4868 gnd.n2041 31.8661
R8379 gnd.n4882 gnd.n2041 31.8661
R8380 gnd.n5626 gnd.n1717 31.8661
R8381 gnd.n5635 gnd.n1717 31.8661
R8382 gnd.n5635 gnd.n1711 31.8661
R8383 gnd.n5643 gnd.n1711 31.8661
R8384 gnd.n5652 gnd.n1705 31.8661
R8385 gnd.n5652 gnd.n1699 31.8661
R8386 gnd.n5660 gnd.n1699 31.8661
R8387 gnd.n5669 gnd.n1693 31.8661
R8388 gnd.n5669 gnd.n1686 31.8661
R8389 gnd.n5677 gnd.n1686 31.8661
R8390 gnd.n5677 gnd.n1687 31.8661
R8391 gnd.n5686 gnd.n1675 31.8661
R8392 gnd.n5697 gnd.n1675 31.8661
R8393 gnd.n5697 gnd.n1669 31.8661
R8394 gnd.n5706 gnd.n1669 31.8661
R8395 gnd.n6149 gnd.n1294 31.8661
R8396 gnd.n6149 gnd.n1296 31.8661
R8397 gnd.n5727 gnd.n1662 31.8661
R8398 gnd.n1662 gnd.n1363 31.8661
R8399 gnd.n1473 gnd.n1405 31.8661
R8400 gnd.n7345 gnd.n368 31.8661
R8401 gnd.n7603 gnd.n107 31.8661
R8402 gnd.n7597 gnd.n107 31.8661
R8403 gnd.n7591 gnd.n124 31.8661
R8404 gnd.n7585 gnd.n133 31.8661
R8405 gnd.n7585 gnd.n136 31.8661
R8406 gnd.n7579 gnd.n146 31.8661
R8407 gnd.n7573 gnd.n146 31.8661
R8408 gnd.n7567 gnd.n162 31.8661
R8409 gnd.n7561 gnd.n171 31.8661
R8410 gnd.n7561 gnd.n174 31.8661
R8411 gnd.n7549 gnd.n191 31.8661
R8412 gnd.n7549 gnd.n194 31.8661
R8413 gnd.n7543 gnd.n194 31.8661
R8414 gnd.n7537 gnd.n209 31.8661
R8415 gnd.n5618 gnd.n1728 30.5915
R8416 gnd.n4415 gnd.t200 27.7236
R8417 gnd.n162 gnd.t276 27.7236
R8418 gnd.n2474 gnd.t198 27.0862
R8419 gnd.n2066 gnd.t52 27.0862
R8420 gnd.t43 gnd.n1705 27.0862
R8421 gnd.n124 gnd.t223 27.0862
R8422 gnd.n4516 gnd.t273 26.4489
R8423 gnd.n7296 gnd.t204 26.4489
R8424 gnd.n4472 gnd.t234 25.8116
R8425 gnd.n7591 gnd.t194 25.8116
R8426 gnd.n2370 gnd.n2369 25.7944
R8427 gnd.n6085 gnd.n6084 25.7944
R8428 gnd.n3063 gnd.n3062 25.7944
R8429 gnd.n2605 gnd.n2604 25.7944
R8430 gnd.n2377 gnd.n2376 25.7944
R8431 gnd.n1428 gnd.n1427 25.7944
R8432 gnd.n1451 gnd.n1450 25.7944
R8433 gnd.n5965 gnd.n5964 25.7944
R8434 gnd.n314 gnd.n313 25.7944
R8435 gnd.n281 gnd.n280 25.7944
R8436 gnd.n7501 gnd.n7500 25.7944
R8437 gnd.n351 gnd.n350 25.7944
R8438 gnd.n4102 gnd.n4101 25.7944
R8439 gnd.n4124 gnd.n4123 25.7944
R8440 gnd.n4145 gnd.n4144 25.7944
R8441 gnd.n4163 gnd.n4162 25.7944
R8442 gnd.n1102 gnd.n1101 25.7944
R8443 gnd.n2195 gnd.n2194 25.7944
R8444 gnd.n2217 gnd.n2216 25.7944
R8445 gnd.n1356 gnd.n1355 25.7944
R8446 gnd.t228 gnd.n2508 25.1743
R8447 gnd.n7567 gnd.t212 25.1743
R8448 gnd.n3284 gnd.n3004 24.8557
R8449 gnd.n3294 gnd.n2987 24.8557
R8450 gnd.n2990 gnd.n2978 24.8557
R8451 gnd.n3315 gnd.n2979 24.8557
R8452 gnd.n3325 gnd.n2959 24.8557
R8453 gnd.n3335 gnd.n3334 24.8557
R8454 gnd.n2945 gnd.n2943 24.8557
R8455 gnd.n3366 gnd.n3365 24.8557
R8456 gnd.n3381 gnd.n2928 24.8557
R8457 gnd.n3435 gnd.n2867 24.8557
R8458 gnd.n3391 gnd.n2868 24.8557
R8459 gnd.n3428 gnd.n2879 24.8557
R8460 gnd.n2917 gnd.n2916 24.8557
R8461 gnd.n3422 gnd.n3421 24.8557
R8462 gnd.n2903 gnd.n2890 24.8557
R8463 gnd.n3461 gnd.n3460 24.8557
R8464 gnd.n3471 gnd.n2783 24.8557
R8465 gnd.n3483 gnd.n2775 24.8557
R8466 gnd.n3482 gnd.n2763 24.8557
R8467 gnd.n3501 gnd.n3500 24.8557
R8468 gnd.n3511 gnd.n2756 24.8557
R8469 gnd.n3522 gnd.n2744 24.8557
R8470 gnd.n3546 gnd.n3545 24.8557
R8471 gnd.n3557 gnd.n2727 24.8557
R8472 gnd.n3556 gnd.n2729 24.8557
R8473 gnd.n3568 gnd.n2720 24.8557
R8474 gnd.n3586 gnd.n3585 24.8557
R8475 gnd.n2711 gnd.n2700 24.8557
R8476 gnd.n3607 gnd.n2688 24.8557
R8477 gnd.n3635 gnd.n3634 24.8557
R8478 gnd.n3646 gnd.n2673 24.8557
R8479 gnd.n3658 gnd.n2666 24.8557
R8480 gnd.n3930 gnd.n3929 24.8557
R8481 gnd.n3952 gnd.n2639 24.8557
R8482 gnd.n2114 gnd.t117 24.537
R8483 gnd.n4830 gnd.t360 24.537
R8484 gnd.n5660 gnd.t49 24.537
R8485 gnd.t91 gnd.n1294 24.537
R8486 gnd.n4773 gnd.n2112 23.8997
R8487 gnd.n5728 gnd.n1296 23.8997
R8488 gnd.n4897 gnd.n4896 23.855
R8489 gnd.n1766 gnd.n1765 23.855
R8490 gnd.n6279 gnd.n6278 23.855
R8491 gnd.n5476 gnd.n5475 23.855
R8492 gnd.n3305 gnd.t358 23.2624
R8493 gnd.n7555 gnd.n184 23.2624
R8494 gnd.n3006 gnd.t109 22.6251
R8495 gnd.n4367 gnd.t81 22.6251
R8496 gnd.n209 gnd.t95 22.6251
R8497 gnd.n4990 gnd.n4892 21.6691
R8498 gnd.n5053 gnd.n2021 21.6691
R8499 gnd.n5083 gnd.t58 21.6691
R8500 gnd.n5076 gnd.n1983 21.6691
R8501 gnd.n5120 gnd.n5119 21.6691
R8502 gnd.n5168 gnd.n1955 21.6691
R8503 gnd.n5168 gnd.n1957 21.6691
R8504 gnd.n5187 gnd.n1947 21.6691
R8505 gnd.n5193 gnd.n1943 21.6691
R8506 gnd.n5224 gnd.n1913 21.6691
R8507 gnd.n5247 gnd.n1887 21.6691
R8508 gnd.n5252 gnd.n1880 21.6691
R8509 gnd.n5289 gnd.n1872 21.6691
R8510 gnd.n5289 gnd.n1860 21.6691
R8511 gnd.n5294 gnd.n1853 21.6691
R8512 gnd.n5353 gnd.n1845 21.6691
R8513 gnd.t23 gnd.n1841 21.6691
R8514 gnd.n5389 gnd.n1808 21.6691
R8515 gnd.n5435 gnd.n1784 21.6691
R8516 gnd.t45 gnd.n3011 21.3504
R8517 gnd.n6277 gnd.n6276 21.0737
R8518 gnd.n5544 gnd.n5543 21.0737
R8519 gnd.n3656 gnd.n931 20.8076
R8520 gnd.t33 gnd.n2701 20.7131
R8521 gnd.n6273 gnd.n1183 20.3945
R8522 gnd.n4984 gnd.n4970 20.3945
R8523 gnd.n5126 gnd.n1973 20.3945
R8524 gnd.n5317 gnd.n1863 20.3945
R8525 gnd.t31 gnd.n2736 20.0758
R8526 gnd.t56 gnd.n1801 20.0758
R8527 gnd.n1166 gnd.t140 19.8005
R8528 gnd.n1166 gnd.t100 19.8005
R8529 gnd.n1165 gnd.t125 19.8005
R8530 gnd.n1165 gnd.t181 19.8005
R8531 gnd.n5466 gnd.t191 19.8005
R8532 gnd.n5466 gnd.t137 19.8005
R8533 gnd.n5465 gnd.t86 19.8005
R8534 gnd.n5465 gnd.t162 19.8005
R8535 gnd.n4650 gnd.n1073 19.7572
R8536 gnd.n6081 gnd.n1363 19.7572
R8537 gnd.n1162 gnd.n1161 19.5087
R8538 gnd.n1175 gnd.n1162 19.5087
R8539 gnd.n1173 gnd.n1164 19.5087
R8540 gnd.n5470 gnd.n5464 19.5087
R8541 gnd.n3472 gnd.t24 19.4385
R8542 gnd.n4806 gnd.t6 19.4385
R8543 gnd.n6343 gnd.n1125 19.4385
R8544 gnd.n5211 gnd.t364 19.4385
R8545 gnd.n5217 gnd.t362 19.4385
R8546 gnd.n5686 gnd.t352 19.4385
R8547 gnd.n4784 gnd.n2109 19.3944
R8548 gnd.n4788 gnd.n2109 19.3944
R8549 gnd.n4788 gnd.n2098 19.3944
R8550 gnd.n4800 gnd.n2098 19.3944
R8551 gnd.n4800 gnd.n2096 19.3944
R8552 gnd.n4804 gnd.n2096 19.3944
R8553 gnd.n4804 gnd.n2084 19.3944
R8554 gnd.n4816 gnd.n2084 19.3944
R8555 gnd.n4816 gnd.n2082 19.3944
R8556 gnd.n4820 gnd.n2082 19.3944
R8557 gnd.n4820 gnd.n2070 19.3944
R8558 gnd.n4832 gnd.n2070 19.3944
R8559 gnd.n4832 gnd.n2068 19.3944
R8560 gnd.n4836 gnd.n2068 19.3944
R8561 gnd.n4836 gnd.n2056 19.3944
R8562 gnd.n4848 gnd.n2056 19.3944
R8563 gnd.n4848 gnd.n2053 19.3944
R8564 gnd.n4866 gnd.n2053 19.3944
R8565 gnd.n4866 gnd.n2054 19.3944
R8566 gnd.n4862 gnd.n2054 19.3944
R8567 gnd.n4862 gnd.n4861 19.3944
R8568 gnd.n4861 gnd.n4860 19.3944
R8569 gnd.n4860 gnd.n4855 19.3944
R8570 gnd.n4856 gnd.n4855 19.3944
R8571 gnd.n4856 gnd.n1198 19.3944
R8572 gnd.n6264 gnd.n1198 19.3944
R8573 gnd.n6264 gnd.n1199 19.3944
R8574 gnd.n6260 gnd.n1199 19.3944
R8575 gnd.n6260 gnd.n6259 19.3944
R8576 gnd.n6259 gnd.n6258 19.3944
R8577 gnd.n6258 gnd.n1205 19.3944
R8578 gnd.n6254 gnd.n1205 19.3944
R8579 gnd.n6254 gnd.n6253 19.3944
R8580 gnd.n6253 gnd.n6252 19.3944
R8581 gnd.n6252 gnd.n1210 19.3944
R8582 gnd.n6248 gnd.n1210 19.3944
R8583 gnd.n6248 gnd.n6247 19.3944
R8584 gnd.n6247 gnd.n6246 19.3944
R8585 gnd.n6246 gnd.n1215 19.3944
R8586 gnd.n6242 gnd.n1215 19.3944
R8587 gnd.n6242 gnd.n6241 19.3944
R8588 gnd.n6241 gnd.n6240 19.3944
R8589 gnd.n6240 gnd.n1220 19.3944
R8590 gnd.n6236 gnd.n1220 19.3944
R8591 gnd.n6236 gnd.n6235 19.3944
R8592 gnd.n6235 gnd.n6234 19.3944
R8593 gnd.n6234 gnd.n1225 19.3944
R8594 gnd.n6230 gnd.n1225 19.3944
R8595 gnd.n6230 gnd.n6229 19.3944
R8596 gnd.n6229 gnd.n6228 19.3944
R8597 gnd.n6228 gnd.n1230 19.3944
R8598 gnd.n6224 gnd.n1230 19.3944
R8599 gnd.n6224 gnd.n6223 19.3944
R8600 gnd.n6223 gnd.n6222 19.3944
R8601 gnd.n6222 gnd.n1235 19.3944
R8602 gnd.n6218 gnd.n1235 19.3944
R8603 gnd.n6218 gnd.n6217 19.3944
R8604 gnd.n6217 gnd.n6216 19.3944
R8605 gnd.n6216 gnd.n1240 19.3944
R8606 gnd.n6212 gnd.n1240 19.3944
R8607 gnd.n6212 gnd.n6211 19.3944
R8608 gnd.n6211 gnd.n6210 19.3944
R8609 gnd.n6210 gnd.n1245 19.3944
R8610 gnd.n6206 gnd.n1245 19.3944
R8611 gnd.n6206 gnd.n6205 19.3944
R8612 gnd.n6205 gnd.n6204 19.3944
R8613 gnd.n6204 gnd.n1250 19.3944
R8614 gnd.n6200 gnd.n1250 19.3944
R8615 gnd.n6200 gnd.n6199 19.3944
R8616 gnd.n6199 gnd.n6198 19.3944
R8617 gnd.n6198 gnd.n1255 19.3944
R8618 gnd.n6194 gnd.n1255 19.3944
R8619 gnd.n6194 gnd.n6193 19.3944
R8620 gnd.n6193 gnd.n6192 19.3944
R8621 gnd.n6192 gnd.n1260 19.3944
R8622 gnd.n6188 gnd.n1260 19.3944
R8623 gnd.n6188 gnd.n6187 19.3944
R8624 gnd.n6187 gnd.n6186 19.3944
R8625 gnd.n6186 gnd.n1265 19.3944
R8626 gnd.n6182 gnd.n1265 19.3944
R8627 gnd.n6182 gnd.n6181 19.3944
R8628 gnd.n6181 gnd.n6180 19.3944
R8629 gnd.n6180 gnd.n1270 19.3944
R8630 gnd.n6176 gnd.n1270 19.3944
R8631 gnd.n6176 gnd.n6175 19.3944
R8632 gnd.n6175 gnd.n6174 19.3944
R8633 gnd.n6174 gnd.n1275 19.3944
R8634 gnd.n6170 gnd.n1275 19.3944
R8635 gnd.n6170 gnd.n6169 19.3944
R8636 gnd.n6169 gnd.n6168 19.3944
R8637 gnd.n6168 gnd.n1280 19.3944
R8638 gnd.n6164 gnd.n1280 19.3944
R8639 gnd.n6164 gnd.n6163 19.3944
R8640 gnd.n6163 gnd.n6162 19.3944
R8641 gnd.n6162 gnd.n1285 19.3944
R8642 gnd.n6158 gnd.n1285 19.3944
R8643 gnd.n6158 gnd.n6157 19.3944
R8644 gnd.n6157 gnd.n6156 19.3944
R8645 gnd.n6156 gnd.n1290 19.3944
R8646 gnd.n6152 gnd.n1290 19.3944
R8647 gnd.n6152 gnd.n6151 19.3944
R8648 gnd.n4702 gnd.n4701 19.3944
R8649 gnd.n4706 gnd.n4702 19.3944
R8650 gnd.n4706 gnd.n4705 19.3944
R8651 gnd.n4770 gnd.n4769 19.3944
R8652 gnd.n4769 gnd.n2187 19.3944
R8653 gnd.n4765 gnd.n2187 19.3944
R8654 gnd.n4765 gnd.n4764 19.3944
R8655 gnd.n4764 gnd.n4763 19.3944
R8656 gnd.n4763 gnd.n2192 19.3944
R8657 gnd.n4758 gnd.n2192 19.3944
R8658 gnd.n4758 gnd.n4757 19.3944
R8659 gnd.n4757 gnd.n4756 19.3944
R8660 gnd.n4756 gnd.n2311 19.3944
R8661 gnd.n4749 gnd.n2311 19.3944
R8662 gnd.n4749 gnd.n4748 19.3944
R8663 gnd.n4748 gnd.n2324 19.3944
R8664 gnd.n4741 gnd.n2324 19.3944
R8665 gnd.n4741 gnd.n4740 19.3944
R8666 gnd.n4740 gnd.n2334 19.3944
R8667 gnd.n4733 gnd.n2334 19.3944
R8668 gnd.n4733 gnd.n4732 19.3944
R8669 gnd.n4732 gnd.n2347 19.3944
R8670 gnd.n4725 gnd.n2347 19.3944
R8671 gnd.n4725 gnd.n4724 19.3944
R8672 gnd.n4724 gnd.n2357 19.3944
R8673 gnd.n4717 gnd.n2357 19.3944
R8674 gnd.n4717 gnd.n4716 19.3944
R8675 gnd.n6127 gnd.n1316 19.3944
R8676 gnd.n6127 gnd.n6126 19.3944
R8677 gnd.n6126 gnd.n1319 19.3944
R8678 gnd.n6119 gnd.n1319 19.3944
R8679 gnd.n6119 gnd.n6118 19.3944
R8680 gnd.n6118 gnd.n1327 19.3944
R8681 gnd.n6111 gnd.n1327 19.3944
R8682 gnd.n6111 gnd.n6110 19.3944
R8683 gnd.n6110 gnd.n1335 19.3944
R8684 gnd.n6103 gnd.n1335 19.3944
R8685 gnd.n6103 gnd.n6102 19.3944
R8686 gnd.n6102 gnd.n1343 19.3944
R8687 gnd.n6095 gnd.n1343 19.3944
R8688 gnd.n6095 gnd.n6094 19.3944
R8689 gnd.n6094 gnd.n1351 19.3944
R8690 gnd.n6087 gnd.n1351 19.3944
R8691 gnd.n3187 gnd.n3186 19.3944
R8692 gnd.n3186 gnd.n3185 19.3944
R8693 gnd.n3185 gnd.n3184 19.3944
R8694 gnd.n3184 gnd.n3182 19.3944
R8695 gnd.n3182 gnd.n3179 19.3944
R8696 gnd.n3179 gnd.n3178 19.3944
R8697 gnd.n3178 gnd.n3175 19.3944
R8698 gnd.n3175 gnd.n3174 19.3944
R8699 gnd.n3174 gnd.n3171 19.3944
R8700 gnd.n3171 gnd.n3170 19.3944
R8701 gnd.n3170 gnd.n3167 19.3944
R8702 gnd.n3167 gnd.n3166 19.3944
R8703 gnd.n3166 gnd.n3163 19.3944
R8704 gnd.n3163 gnd.n3162 19.3944
R8705 gnd.n3162 gnd.n3159 19.3944
R8706 gnd.n3159 gnd.n3158 19.3944
R8707 gnd.n3158 gnd.n3155 19.3944
R8708 gnd.n3155 gnd.n3154 19.3944
R8709 gnd.n3154 gnd.n3151 19.3944
R8710 gnd.n3151 gnd.n3150 19.3944
R8711 gnd.n3150 gnd.n3147 19.3944
R8712 gnd.n3147 gnd.n3146 19.3944
R8713 gnd.n3143 gnd.n3142 19.3944
R8714 gnd.n3142 gnd.n3098 19.3944
R8715 gnd.n3193 gnd.n3098 19.3944
R8716 gnd.n3960 gnd.n3959 19.3944
R8717 gnd.n3959 gnd.n3956 19.3944
R8718 gnd.n3956 gnd.n3955 19.3944
R8719 gnd.n4005 gnd.n4004 19.3944
R8720 gnd.n4004 gnd.n4003 19.3944
R8721 gnd.n4003 gnd.n4000 19.3944
R8722 gnd.n4000 gnd.n3999 19.3944
R8723 gnd.n3999 gnd.n3996 19.3944
R8724 gnd.n3996 gnd.n3995 19.3944
R8725 gnd.n3995 gnd.n3992 19.3944
R8726 gnd.n3992 gnd.n3991 19.3944
R8727 gnd.n3991 gnd.n3988 19.3944
R8728 gnd.n3988 gnd.n3987 19.3944
R8729 gnd.n3987 gnd.n3984 19.3944
R8730 gnd.n3984 gnd.n3983 19.3944
R8731 gnd.n3983 gnd.n3980 19.3944
R8732 gnd.n3980 gnd.n3979 19.3944
R8733 gnd.n3979 gnd.n3976 19.3944
R8734 gnd.n3976 gnd.n3975 19.3944
R8735 gnd.n3975 gnd.n3972 19.3944
R8736 gnd.n3972 gnd.n3971 19.3944
R8737 gnd.n3971 gnd.n3968 19.3944
R8738 gnd.n3968 gnd.n3967 19.3944
R8739 gnd.n3967 gnd.n3964 19.3944
R8740 gnd.n3964 gnd.n3963 19.3944
R8741 gnd.n3286 gnd.n2995 19.3944
R8742 gnd.n3296 gnd.n2995 19.3944
R8743 gnd.n3297 gnd.n3296 19.3944
R8744 gnd.n3297 gnd.n2976 19.3944
R8745 gnd.n3317 gnd.n2976 19.3944
R8746 gnd.n3317 gnd.n2968 19.3944
R8747 gnd.n3327 gnd.n2968 19.3944
R8748 gnd.n3328 gnd.n3327 19.3944
R8749 gnd.n3329 gnd.n3328 19.3944
R8750 gnd.n3329 gnd.n2951 19.3944
R8751 gnd.n3346 gnd.n2951 19.3944
R8752 gnd.n3349 gnd.n3346 19.3944
R8753 gnd.n3349 gnd.n3348 19.3944
R8754 gnd.n3348 gnd.n2924 19.3944
R8755 gnd.n3388 gnd.n2924 19.3944
R8756 gnd.n3388 gnd.n2921 19.3944
R8757 gnd.n3394 gnd.n2921 19.3944
R8758 gnd.n3395 gnd.n3394 19.3944
R8759 gnd.n3395 gnd.n2919 19.3944
R8760 gnd.n3401 gnd.n2919 19.3944
R8761 gnd.n3404 gnd.n3401 19.3944
R8762 gnd.n3406 gnd.n3404 19.3944
R8763 gnd.n3412 gnd.n3406 19.3944
R8764 gnd.n3412 gnd.n3411 19.3944
R8765 gnd.n3411 gnd.n2778 19.3944
R8766 gnd.n3478 gnd.n2778 19.3944
R8767 gnd.n3479 gnd.n3478 19.3944
R8768 gnd.n3479 gnd.n2771 19.3944
R8769 gnd.n3490 gnd.n2771 19.3944
R8770 gnd.n3491 gnd.n3490 19.3944
R8771 gnd.n3491 gnd.n2754 19.3944
R8772 gnd.n2754 gnd.n2752 19.3944
R8773 gnd.n3515 gnd.n2752 19.3944
R8774 gnd.n3516 gnd.n3515 19.3944
R8775 gnd.n3516 gnd.n2723 19.3944
R8776 gnd.n3563 gnd.n2723 19.3944
R8777 gnd.n3564 gnd.n3563 19.3944
R8778 gnd.n3564 gnd.n2716 19.3944
R8779 gnd.n3575 gnd.n2716 19.3944
R8780 gnd.n3576 gnd.n3575 19.3944
R8781 gnd.n3576 gnd.n2699 19.3944
R8782 gnd.n2699 gnd.n2697 19.3944
R8783 gnd.n3600 gnd.n2697 19.3944
R8784 gnd.n3601 gnd.n3600 19.3944
R8785 gnd.n3601 gnd.n2669 19.3944
R8786 gnd.n3652 gnd.n2669 19.3944
R8787 gnd.n3653 gnd.n3652 19.3944
R8788 gnd.n3653 gnd.n2662 19.3944
R8789 gnd.n3921 gnd.n2662 19.3944
R8790 gnd.n3922 gnd.n3921 19.3944
R8791 gnd.n3922 gnd.n2643 19.3944
R8792 gnd.n3947 gnd.n2643 19.3944
R8793 gnd.n3947 gnd.n2644 19.3944
R8794 gnd.n3277 gnd.n3276 19.3944
R8795 gnd.n3276 gnd.n3009 19.3944
R8796 gnd.n3032 gnd.n3009 19.3944
R8797 gnd.n3035 gnd.n3032 19.3944
R8798 gnd.n3035 gnd.n3028 19.3944
R8799 gnd.n3039 gnd.n3028 19.3944
R8800 gnd.n3042 gnd.n3039 19.3944
R8801 gnd.n3045 gnd.n3042 19.3944
R8802 gnd.n3045 gnd.n3026 19.3944
R8803 gnd.n3049 gnd.n3026 19.3944
R8804 gnd.n3052 gnd.n3049 19.3944
R8805 gnd.n3055 gnd.n3052 19.3944
R8806 gnd.n3055 gnd.n3024 19.3944
R8807 gnd.n3059 gnd.n3024 19.3944
R8808 gnd.n3282 gnd.n3281 19.3944
R8809 gnd.n3281 gnd.n2985 19.3944
R8810 gnd.n3307 gnd.n2985 19.3944
R8811 gnd.n3307 gnd.n2983 19.3944
R8812 gnd.n3313 gnd.n2983 19.3944
R8813 gnd.n3313 gnd.n3312 19.3944
R8814 gnd.n3312 gnd.n2957 19.3944
R8815 gnd.n3337 gnd.n2957 19.3944
R8816 gnd.n3337 gnd.n2955 19.3944
R8817 gnd.n3341 gnd.n2955 19.3944
R8818 gnd.n3341 gnd.n2935 19.3944
R8819 gnd.n3368 gnd.n2935 19.3944
R8820 gnd.n3368 gnd.n2933 19.3944
R8821 gnd.n3378 gnd.n2933 19.3944
R8822 gnd.n3378 gnd.n3377 19.3944
R8823 gnd.n3377 gnd.n3376 19.3944
R8824 gnd.n3376 gnd.n2882 19.3944
R8825 gnd.n3426 gnd.n2882 19.3944
R8826 gnd.n3426 gnd.n3425 19.3944
R8827 gnd.n3425 gnd.n3424 19.3944
R8828 gnd.n3424 gnd.n2886 19.3944
R8829 gnd.n2906 gnd.n2886 19.3944
R8830 gnd.n2906 gnd.n2788 19.3944
R8831 gnd.n3463 gnd.n2788 19.3944
R8832 gnd.n3463 gnd.n2786 19.3944
R8833 gnd.n3469 gnd.n2786 19.3944
R8834 gnd.n3469 gnd.n3468 19.3944
R8835 gnd.n3468 gnd.n2761 19.3944
R8836 gnd.n3503 gnd.n2761 19.3944
R8837 gnd.n3503 gnd.n2759 19.3944
R8838 gnd.n3509 gnd.n2759 19.3944
R8839 gnd.n3509 gnd.n3508 19.3944
R8840 gnd.n3508 gnd.n2734 19.3944
R8841 gnd.n3548 gnd.n2734 19.3944
R8842 gnd.n3548 gnd.n2732 19.3944
R8843 gnd.n3554 gnd.n2732 19.3944
R8844 gnd.n3554 gnd.n3553 19.3944
R8845 gnd.n3553 gnd.n2706 19.3944
R8846 gnd.n3588 gnd.n2706 19.3944
R8847 gnd.n3588 gnd.n2704 19.3944
R8848 gnd.n3594 gnd.n2704 19.3944
R8849 gnd.n3594 gnd.n3593 19.3944
R8850 gnd.n3593 gnd.n2679 19.3944
R8851 gnd.n3637 gnd.n2679 19.3944
R8852 gnd.n3637 gnd.n2677 19.3944
R8853 gnd.n3643 gnd.n2677 19.3944
R8854 gnd.n3643 gnd.n3642 19.3944
R8855 gnd.n3642 gnd.n2652 19.3944
R8856 gnd.n3932 gnd.n2652 19.3944
R8857 gnd.n3932 gnd.n2650 19.3944
R8858 gnd.n3940 gnd.n2650 19.3944
R8859 gnd.n3940 gnd.n3939 19.3944
R8860 gnd.n3939 gnd.n3938 19.3944
R8861 gnd.n4041 gnd.n4040 19.3944
R8862 gnd.n4040 gnd.n2591 19.3944
R8863 gnd.n4036 gnd.n2591 19.3944
R8864 gnd.n4036 gnd.n4033 19.3944
R8865 gnd.n4033 gnd.n4030 19.3944
R8866 gnd.n4030 gnd.n4029 19.3944
R8867 gnd.n4029 gnd.n4026 19.3944
R8868 gnd.n4026 gnd.n4025 19.3944
R8869 gnd.n4025 gnd.n4022 19.3944
R8870 gnd.n4022 gnd.n4021 19.3944
R8871 gnd.n4021 gnd.n4018 19.3944
R8872 gnd.n4018 gnd.n4017 19.3944
R8873 gnd.n4017 gnd.n4014 19.3944
R8874 gnd.n4014 gnd.n4013 19.3944
R8875 gnd.n3197 gnd.n3096 19.3944
R8876 gnd.n3197 gnd.n3087 19.3944
R8877 gnd.n3210 gnd.n3087 19.3944
R8878 gnd.n3210 gnd.n3085 19.3944
R8879 gnd.n3214 gnd.n3085 19.3944
R8880 gnd.n3214 gnd.n3075 19.3944
R8881 gnd.n3226 gnd.n3075 19.3944
R8882 gnd.n3226 gnd.n3073 19.3944
R8883 gnd.n3260 gnd.n3073 19.3944
R8884 gnd.n3260 gnd.n3259 19.3944
R8885 gnd.n3259 gnd.n3258 19.3944
R8886 gnd.n3258 gnd.n3257 19.3944
R8887 gnd.n3257 gnd.n3254 19.3944
R8888 gnd.n3254 gnd.n3253 19.3944
R8889 gnd.n3253 gnd.n3252 19.3944
R8890 gnd.n3252 gnd.n3250 19.3944
R8891 gnd.n3250 gnd.n3249 19.3944
R8892 gnd.n3249 gnd.n3246 19.3944
R8893 gnd.n3246 gnd.n3245 19.3944
R8894 gnd.n3245 gnd.n3244 19.3944
R8895 gnd.n3244 gnd.n3242 19.3944
R8896 gnd.n3242 gnd.n2941 19.3944
R8897 gnd.n3357 gnd.n2941 19.3944
R8898 gnd.n3357 gnd.n2939 19.3944
R8899 gnd.n3363 gnd.n2939 19.3944
R8900 gnd.n3363 gnd.n3362 19.3944
R8901 gnd.n3362 gnd.n2863 19.3944
R8902 gnd.n3437 gnd.n2863 19.3944
R8903 gnd.n3437 gnd.n2864 19.3944
R8904 gnd.n2911 gnd.n2910 19.3944
R8905 gnd.n2914 gnd.n2913 19.3944
R8906 gnd.n2901 gnd.n2900 19.3944
R8907 gnd.n3456 gnd.n2793 19.3944
R8908 gnd.n3456 gnd.n3455 19.3944
R8909 gnd.n3455 gnd.n3454 19.3944
R8910 gnd.n3454 gnd.n3452 19.3944
R8911 gnd.n3452 gnd.n3451 19.3944
R8912 gnd.n3451 gnd.n3449 19.3944
R8913 gnd.n3449 gnd.n3448 19.3944
R8914 gnd.n3448 gnd.n2742 19.3944
R8915 gnd.n3524 gnd.n2742 19.3944
R8916 gnd.n3524 gnd.n2740 19.3944
R8917 gnd.n3543 gnd.n2740 19.3944
R8918 gnd.n3543 gnd.n3542 19.3944
R8919 gnd.n3542 gnd.n3541 19.3944
R8920 gnd.n3541 gnd.n3539 19.3944
R8921 gnd.n3539 gnd.n3538 19.3944
R8922 gnd.n3538 gnd.n3536 19.3944
R8923 gnd.n3536 gnd.n3535 19.3944
R8924 gnd.n3535 gnd.n2686 19.3944
R8925 gnd.n3609 gnd.n2686 19.3944
R8926 gnd.n3609 gnd.n2684 19.3944
R8927 gnd.n3632 gnd.n2684 19.3944
R8928 gnd.n3632 gnd.n3631 19.3944
R8929 gnd.n3631 gnd.n3630 19.3944
R8930 gnd.n3630 gnd.n3627 19.3944
R8931 gnd.n3627 gnd.n3626 19.3944
R8932 gnd.n3626 gnd.n3624 19.3944
R8933 gnd.n3624 gnd.n3623 19.3944
R8934 gnd.n3623 gnd.n3621 19.3944
R8935 gnd.n3621 gnd.n2638 19.3944
R8936 gnd.n3202 gnd.n3092 19.3944
R8937 gnd.n3202 gnd.n3090 19.3944
R8938 gnd.n3206 gnd.n3090 19.3944
R8939 gnd.n3206 gnd.n3081 19.3944
R8940 gnd.n3218 gnd.n3081 19.3944
R8941 gnd.n3218 gnd.n3079 19.3944
R8942 gnd.n3222 gnd.n3079 19.3944
R8943 gnd.n3222 gnd.n3068 19.3944
R8944 gnd.n3264 gnd.n3068 19.3944
R8945 gnd.n3264 gnd.n3022 19.3944
R8946 gnd.n3270 gnd.n3022 19.3944
R8947 gnd.n3270 gnd.n3269 19.3944
R8948 gnd.n3269 gnd.n3000 19.3944
R8949 gnd.n3291 gnd.n3000 19.3944
R8950 gnd.n3291 gnd.n2993 19.3944
R8951 gnd.n3302 gnd.n2993 19.3944
R8952 gnd.n3302 gnd.n3301 19.3944
R8953 gnd.n3301 gnd.n2974 19.3944
R8954 gnd.n3322 gnd.n2974 19.3944
R8955 gnd.n3322 gnd.n2964 19.3944
R8956 gnd.n3332 gnd.n2964 19.3944
R8957 gnd.n3332 gnd.n2947 19.3944
R8958 gnd.n3353 gnd.n2947 19.3944
R8959 gnd.n3353 gnd.n3352 19.3944
R8960 gnd.n3352 gnd.n2926 19.3944
R8961 gnd.n3383 gnd.n2926 19.3944
R8962 gnd.n3383 gnd.n2871 19.3944
R8963 gnd.n3433 gnd.n2871 19.3944
R8964 gnd.n3433 gnd.n3432 19.3944
R8965 gnd.n3432 gnd.n3431 19.3944
R8966 gnd.n3431 gnd.n2875 19.3944
R8967 gnd.n2893 gnd.n2875 19.3944
R8968 gnd.n3419 gnd.n2893 19.3944
R8969 gnd.n3419 gnd.n3418 19.3944
R8970 gnd.n3418 gnd.n3417 19.3944
R8971 gnd.n3417 gnd.n2897 19.3944
R8972 gnd.n2897 gnd.n2780 19.3944
R8973 gnd.n3474 gnd.n2780 19.3944
R8974 gnd.n3474 gnd.n2773 19.3944
R8975 gnd.n3485 gnd.n2773 19.3944
R8976 gnd.n3485 gnd.n2769 19.3944
R8977 gnd.n3498 gnd.n2769 19.3944
R8978 gnd.n3498 gnd.n3497 19.3944
R8979 gnd.n3497 gnd.n2748 19.3944
R8980 gnd.n3520 gnd.n2748 19.3944
R8981 gnd.n3520 gnd.n3519 19.3944
R8982 gnd.n3519 gnd.n2725 19.3944
R8983 gnd.n3559 gnd.n2725 19.3944
R8984 gnd.n3559 gnd.n2718 19.3944
R8985 gnd.n3570 gnd.n2718 19.3944
R8986 gnd.n3570 gnd.n2714 19.3944
R8987 gnd.n3583 gnd.n2714 19.3944
R8988 gnd.n3583 gnd.n3582 19.3944
R8989 gnd.n3582 gnd.n2693 19.3944
R8990 gnd.n3605 gnd.n2693 19.3944
R8991 gnd.n3605 gnd.n3604 19.3944
R8992 gnd.n3604 gnd.n2671 19.3944
R8993 gnd.n3648 gnd.n2671 19.3944
R8994 gnd.n3648 gnd.n2664 19.3944
R8995 gnd.n3660 gnd.n2664 19.3944
R8996 gnd.n3660 gnd.n2660 19.3944
R8997 gnd.n3927 gnd.n2660 19.3944
R8998 gnd.n3927 gnd.n3926 19.3944
R8999 gnd.n3926 gnd.n2641 19.3944
R9000 gnd.n3950 gnd.n2641 19.3944
R9001 gnd.n4753 gnd.n2314 19.3944
R9002 gnd.n4753 gnd.n4752 19.3944
R9003 gnd.n4752 gnd.n2318 19.3944
R9004 gnd.n4745 gnd.n2318 19.3944
R9005 gnd.n4745 gnd.n4744 19.3944
R9006 gnd.n4744 gnd.n2330 19.3944
R9007 gnd.n4737 gnd.n2330 19.3944
R9008 gnd.n4737 gnd.n4736 19.3944
R9009 gnd.n4736 gnd.n2341 19.3944
R9010 gnd.n4729 gnd.n2341 19.3944
R9011 gnd.n4729 gnd.n4728 19.3944
R9012 gnd.n4728 gnd.n2353 19.3944
R9013 gnd.n4721 gnd.n2353 19.3944
R9014 gnd.n4721 gnd.n4720 19.3944
R9015 gnd.n4720 gnd.n2364 19.3944
R9016 gnd.n4713 gnd.n2364 19.3944
R9017 gnd.n2430 gnd.n2427 19.3944
R9018 gnd.n4538 gnd.n2430 19.3944
R9019 gnd.n4538 gnd.n2426 19.3944
R9020 gnd.n4562 gnd.n2426 19.3944
R9021 gnd.n4562 gnd.n4561 19.3944
R9022 gnd.n4561 gnd.n4560 19.3944
R9023 gnd.n4560 gnd.n4544 19.3944
R9024 gnd.n4556 gnd.n4544 19.3944
R9025 gnd.n4556 gnd.n4555 19.3944
R9026 gnd.n4555 gnd.n4554 19.3944
R9027 gnd.n4554 gnd.n4552 19.3944
R9028 gnd.n4552 gnd.n2402 19.3944
R9029 gnd.n2402 gnd.n2400 19.3944
R9030 gnd.n4629 gnd.n2400 19.3944
R9031 gnd.n4629 gnd.n2398 19.3944
R9032 gnd.n4633 gnd.n2398 19.3944
R9033 gnd.n4633 gnd.n2396 19.3944
R9034 gnd.n4637 gnd.n2396 19.3944
R9035 gnd.n4637 gnd.n2394 19.3944
R9036 gnd.n4669 gnd.n2394 19.3944
R9037 gnd.n4669 gnd.n4668 19.3944
R9038 gnd.n4668 gnd.n4667 19.3944
R9039 gnd.n4667 gnd.n4643 19.3944
R9040 gnd.n4663 gnd.n4643 19.3944
R9041 gnd.n4663 gnd.n4662 19.3944
R9042 gnd.n4662 gnd.n4661 19.3944
R9043 gnd.n4661 gnd.n4649 19.3944
R9044 gnd.n4656 gnd.n4649 19.3944
R9045 gnd.n4656 gnd.n4655 19.3944
R9046 gnd.n4655 gnd.n2118 19.3944
R9047 gnd.n4776 gnd.n2118 19.3944
R9048 gnd.n4776 gnd.n2116 19.3944
R9049 gnd.n4780 gnd.n2116 19.3944
R9050 gnd.n4780 gnd.n2105 19.3944
R9051 gnd.n4792 gnd.n2105 19.3944
R9052 gnd.n4792 gnd.n2103 19.3944
R9053 gnd.n4796 gnd.n2103 19.3944
R9054 gnd.n4796 gnd.n2091 19.3944
R9055 gnd.n4808 gnd.n2091 19.3944
R9056 gnd.n4808 gnd.n2089 19.3944
R9057 gnd.n4812 gnd.n2089 19.3944
R9058 gnd.n4812 gnd.n2076 19.3944
R9059 gnd.n4824 gnd.n2076 19.3944
R9060 gnd.n4824 gnd.n2074 19.3944
R9061 gnd.n4828 gnd.n2074 19.3944
R9062 gnd.n4828 gnd.n2062 19.3944
R9063 gnd.n4840 gnd.n2062 19.3944
R9064 gnd.n4840 gnd.n2060 19.3944
R9065 gnd.n4844 gnd.n2060 19.3944
R9066 gnd.n4844 gnd.n2047 19.3944
R9067 gnd.n4870 gnd.n2047 19.3944
R9068 gnd.n4870 gnd.n2045 19.3944
R9069 gnd.n4880 gnd.n2045 19.3944
R9070 gnd.n4880 gnd.n4879 19.3944
R9071 gnd.n4879 gnd.n4878 19.3944
R9072 gnd.n4878 gnd.n1189 19.3944
R9073 gnd.n6270 gnd.n1189 19.3944
R9074 gnd.n6270 gnd.n6269 19.3944
R9075 gnd.n6269 gnd.n6268 19.3944
R9076 gnd.n6268 gnd.n1193 19.3944
R9077 gnd.n5028 gnd.n1193 19.3944
R9078 gnd.n5032 gnd.n5028 19.3944
R9079 gnd.n5032 gnd.n2017 19.3944
R9080 gnd.n5057 gnd.n2017 19.3944
R9081 gnd.n5057 gnd.n2015 19.3944
R9082 gnd.n5063 gnd.n2015 19.3944
R9083 gnd.n5063 gnd.n5062 19.3944
R9084 gnd.n5062 gnd.n1989 19.3944
R9085 gnd.n5095 gnd.n1989 19.3944
R9086 gnd.n5095 gnd.n1987 19.3944
R9087 gnd.n5105 gnd.n1987 19.3944
R9088 gnd.n5105 gnd.n5104 19.3944
R9089 gnd.n5104 gnd.n5103 19.3944
R9090 gnd.n5103 gnd.n1961 19.3944
R9091 gnd.n5166 gnd.n1961 19.3944
R9092 gnd.n5166 gnd.n5165 19.3944
R9093 gnd.n5165 gnd.n5164 19.3944
R9094 gnd.n5164 gnd.n1939 19.3944
R9095 gnd.n5196 gnd.n1939 19.3944
R9096 gnd.n5196 gnd.n1937 19.3944
R9097 gnd.n5202 gnd.n1937 19.3944
R9098 gnd.n5202 gnd.n5201 19.3944
R9099 gnd.n5201 gnd.n1911 19.3944
R9100 gnd.n5234 gnd.n1911 19.3944
R9101 gnd.n5234 gnd.n1909 19.3944
R9102 gnd.n5238 gnd.n1909 19.3944
R9103 gnd.n5238 gnd.n1885 19.3944
R9104 gnd.n5271 gnd.n1885 19.3944
R9105 gnd.n5271 gnd.n1883 19.3944
R9106 gnd.n5277 gnd.n1883 19.3944
R9107 gnd.n5277 gnd.n5276 19.3944
R9108 gnd.n5276 gnd.n1858 19.3944
R9109 gnd.n5320 gnd.n1858 19.3944
R9110 gnd.n5320 gnd.n1856 19.3944
R9111 gnd.n5326 gnd.n1856 19.3944
R9112 gnd.n5326 gnd.n5325 19.3944
R9113 gnd.n5325 gnd.n1836 19.3944
R9114 gnd.n5361 gnd.n1836 19.3944
R9115 gnd.n5361 gnd.n1834 19.3944
R9116 gnd.n5367 gnd.n1834 19.3944
R9117 gnd.n5367 gnd.n5366 19.3944
R9118 gnd.n5366 gnd.n1806 19.3944
R9119 gnd.n5401 gnd.n1806 19.3944
R9120 gnd.n5401 gnd.n1804 19.3944
R9121 gnd.n5405 gnd.n1804 19.3944
R9122 gnd.n5405 gnd.n1782 19.3944
R9123 gnd.n5444 gnd.n1782 19.3944
R9124 gnd.n5444 gnd.n1780 19.3944
R9125 gnd.n5450 gnd.n1780 19.3944
R9126 gnd.n5450 gnd.n5449 19.3944
R9127 gnd.n5449 gnd.n1726 19.3944
R9128 gnd.n5620 gnd.n1726 19.3944
R9129 gnd.n5620 gnd.n1724 19.3944
R9130 gnd.n5624 gnd.n1724 19.3944
R9131 gnd.n5624 gnd.n1715 19.3944
R9132 gnd.n5637 gnd.n1715 19.3944
R9133 gnd.n5637 gnd.n1713 19.3944
R9134 gnd.n5641 gnd.n1713 19.3944
R9135 gnd.n5641 gnd.n1703 19.3944
R9136 gnd.n5654 gnd.n1703 19.3944
R9137 gnd.n5654 gnd.n1701 19.3944
R9138 gnd.n5658 gnd.n1701 19.3944
R9139 gnd.n5658 gnd.n1691 19.3944
R9140 gnd.n5671 gnd.n1691 19.3944
R9141 gnd.n5671 gnd.n1689 19.3944
R9142 gnd.n5675 gnd.n1689 19.3944
R9143 gnd.n5675 gnd.n1679 19.3944
R9144 gnd.n5688 gnd.n1679 19.3944
R9145 gnd.n5688 gnd.n1677 19.3944
R9146 gnd.n5695 gnd.n1677 19.3944
R9147 gnd.n5695 gnd.n5694 19.3944
R9148 gnd.n5694 gnd.n1667 19.3944
R9149 gnd.n5709 gnd.n1667 19.3944
R9150 gnd.n5710 gnd.n5709 19.3944
R9151 gnd.n5710 gnd.n1665 19.3944
R9152 gnd.n5725 gnd.n1665 19.3944
R9153 gnd.n5725 gnd.n5724 19.3944
R9154 gnd.n5724 gnd.n5723 19.3944
R9155 gnd.n5723 gnd.n5716 19.3944
R9156 gnd.n5719 gnd.n5716 19.3944
R9157 gnd.n5719 gnd.n1631 19.3944
R9158 gnd.n5779 gnd.n1631 19.3944
R9159 gnd.n5779 gnd.n1629 19.3944
R9160 gnd.n5783 gnd.n1629 19.3944
R9161 gnd.n5783 gnd.n1627 19.3944
R9162 gnd.n5787 gnd.n1627 19.3944
R9163 gnd.n5787 gnd.n1625 19.3944
R9164 gnd.n5791 gnd.n1625 19.3944
R9165 gnd.n5791 gnd.n1623 19.3944
R9166 gnd.n5795 gnd.n1623 19.3944
R9167 gnd.n5795 gnd.n1621 19.3944
R9168 gnd.n5819 gnd.n1621 19.3944
R9169 gnd.n5819 gnd.n5818 19.3944
R9170 gnd.n5818 gnd.n5817 19.3944
R9171 gnd.n5817 gnd.n5801 19.3944
R9172 gnd.n5813 gnd.n5801 19.3944
R9173 gnd.n5813 gnd.n5812 19.3944
R9174 gnd.n5812 gnd.n5811 19.3944
R9175 gnd.n5811 gnd.n5809 19.3944
R9176 gnd.n5809 gnd.n1603 19.3944
R9177 gnd.n1603 gnd.n1601 19.3944
R9178 gnd.n5880 gnd.n1601 19.3944
R9179 gnd.n5880 gnd.n1599 19.3944
R9180 gnd.n5885 gnd.n1599 19.3944
R9181 gnd.n5885 gnd.n389 19.3944
R9182 gnd.n7279 gnd.n389 19.3944
R9183 gnd.n7279 gnd.n7278 19.3944
R9184 gnd.n7066 gnd.n516 19.3944
R9185 gnd.n7066 gnd.n512 19.3944
R9186 gnd.n7072 gnd.n512 19.3944
R9187 gnd.n7072 gnd.n510 19.3944
R9188 gnd.n7076 gnd.n510 19.3944
R9189 gnd.n7076 gnd.n506 19.3944
R9190 gnd.n7082 gnd.n506 19.3944
R9191 gnd.n7082 gnd.n504 19.3944
R9192 gnd.n7086 gnd.n504 19.3944
R9193 gnd.n7086 gnd.n500 19.3944
R9194 gnd.n7092 gnd.n500 19.3944
R9195 gnd.n7092 gnd.n498 19.3944
R9196 gnd.n7096 gnd.n498 19.3944
R9197 gnd.n7096 gnd.n494 19.3944
R9198 gnd.n7102 gnd.n494 19.3944
R9199 gnd.n7102 gnd.n492 19.3944
R9200 gnd.n7106 gnd.n492 19.3944
R9201 gnd.n7106 gnd.n488 19.3944
R9202 gnd.n7112 gnd.n488 19.3944
R9203 gnd.n7112 gnd.n486 19.3944
R9204 gnd.n7116 gnd.n486 19.3944
R9205 gnd.n7116 gnd.n482 19.3944
R9206 gnd.n7122 gnd.n482 19.3944
R9207 gnd.n7122 gnd.n480 19.3944
R9208 gnd.n7126 gnd.n480 19.3944
R9209 gnd.n7126 gnd.n476 19.3944
R9210 gnd.n7132 gnd.n476 19.3944
R9211 gnd.n7132 gnd.n474 19.3944
R9212 gnd.n7136 gnd.n474 19.3944
R9213 gnd.n7136 gnd.n470 19.3944
R9214 gnd.n7142 gnd.n470 19.3944
R9215 gnd.n7142 gnd.n468 19.3944
R9216 gnd.n7146 gnd.n468 19.3944
R9217 gnd.n7146 gnd.n464 19.3944
R9218 gnd.n7152 gnd.n464 19.3944
R9219 gnd.n7152 gnd.n462 19.3944
R9220 gnd.n7156 gnd.n462 19.3944
R9221 gnd.n7156 gnd.n458 19.3944
R9222 gnd.n7162 gnd.n458 19.3944
R9223 gnd.n7162 gnd.n456 19.3944
R9224 gnd.n7166 gnd.n456 19.3944
R9225 gnd.n7166 gnd.n452 19.3944
R9226 gnd.n7172 gnd.n452 19.3944
R9227 gnd.n7172 gnd.n450 19.3944
R9228 gnd.n7176 gnd.n450 19.3944
R9229 gnd.n7176 gnd.n446 19.3944
R9230 gnd.n7182 gnd.n446 19.3944
R9231 gnd.n7182 gnd.n444 19.3944
R9232 gnd.n7186 gnd.n444 19.3944
R9233 gnd.n7186 gnd.n440 19.3944
R9234 gnd.n7192 gnd.n440 19.3944
R9235 gnd.n7192 gnd.n438 19.3944
R9236 gnd.n7196 gnd.n438 19.3944
R9237 gnd.n7196 gnd.n434 19.3944
R9238 gnd.n7202 gnd.n434 19.3944
R9239 gnd.n7202 gnd.n432 19.3944
R9240 gnd.n7206 gnd.n432 19.3944
R9241 gnd.n7206 gnd.n428 19.3944
R9242 gnd.n7212 gnd.n428 19.3944
R9243 gnd.n7212 gnd.n426 19.3944
R9244 gnd.n7216 gnd.n426 19.3944
R9245 gnd.n7216 gnd.n422 19.3944
R9246 gnd.n7222 gnd.n422 19.3944
R9247 gnd.n7222 gnd.n420 19.3944
R9248 gnd.n7226 gnd.n420 19.3944
R9249 gnd.n7226 gnd.n416 19.3944
R9250 gnd.n7232 gnd.n416 19.3944
R9251 gnd.n7232 gnd.n414 19.3944
R9252 gnd.n7236 gnd.n414 19.3944
R9253 gnd.n7236 gnd.n410 19.3944
R9254 gnd.n7242 gnd.n410 19.3944
R9255 gnd.n7242 gnd.n408 19.3944
R9256 gnd.n7246 gnd.n408 19.3944
R9257 gnd.n7246 gnd.n404 19.3944
R9258 gnd.n7252 gnd.n404 19.3944
R9259 gnd.n7252 gnd.n402 19.3944
R9260 gnd.n7256 gnd.n402 19.3944
R9261 gnd.n7256 gnd.n398 19.3944
R9262 gnd.n7262 gnd.n398 19.3944
R9263 gnd.n7262 gnd.n396 19.3944
R9264 gnd.n7268 gnd.n396 19.3944
R9265 gnd.n7268 gnd.n7267 19.3944
R9266 gnd.n7267 gnd.n392 19.3944
R9267 gnd.n7275 gnd.n392 19.3944
R9268 gnd.n6646 gnd.n768 19.3944
R9269 gnd.n6646 gnd.n764 19.3944
R9270 gnd.n6652 gnd.n764 19.3944
R9271 gnd.n6652 gnd.n762 19.3944
R9272 gnd.n6656 gnd.n762 19.3944
R9273 gnd.n6656 gnd.n758 19.3944
R9274 gnd.n6662 gnd.n758 19.3944
R9275 gnd.n6662 gnd.n756 19.3944
R9276 gnd.n6666 gnd.n756 19.3944
R9277 gnd.n6666 gnd.n752 19.3944
R9278 gnd.n6672 gnd.n752 19.3944
R9279 gnd.n6672 gnd.n750 19.3944
R9280 gnd.n6676 gnd.n750 19.3944
R9281 gnd.n6676 gnd.n746 19.3944
R9282 gnd.n6682 gnd.n746 19.3944
R9283 gnd.n6682 gnd.n744 19.3944
R9284 gnd.n6686 gnd.n744 19.3944
R9285 gnd.n6686 gnd.n740 19.3944
R9286 gnd.n6692 gnd.n740 19.3944
R9287 gnd.n6692 gnd.n738 19.3944
R9288 gnd.n6696 gnd.n738 19.3944
R9289 gnd.n6696 gnd.n734 19.3944
R9290 gnd.n6702 gnd.n734 19.3944
R9291 gnd.n6702 gnd.n732 19.3944
R9292 gnd.n6706 gnd.n732 19.3944
R9293 gnd.n6706 gnd.n728 19.3944
R9294 gnd.n6712 gnd.n728 19.3944
R9295 gnd.n6712 gnd.n726 19.3944
R9296 gnd.n6716 gnd.n726 19.3944
R9297 gnd.n6716 gnd.n722 19.3944
R9298 gnd.n6722 gnd.n722 19.3944
R9299 gnd.n6722 gnd.n720 19.3944
R9300 gnd.n6726 gnd.n720 19.3944
R9301 gnd.n6726 gnd.n716 19.3944
R9302 gnd.n6732 gnd.n716 19.3944
R9303 gnd.n6732 gnd.n714 19.3944
R9304 gnd.n6736 gnd.n714 19.3944
R9305 gnd.n6736 gnd.n710 19.3944
R9306 gnd.n6742 gnd.n710 19.3944
R9307 gnd.n6742 gnd.n708 19.3944
R9308 gnd.n6746 gnd.n708 19.3944
R9309 gnd.n6746 gnd.n704 19.3944
R9310 gnd.n6752 gnd.n704 19.3944
R9311 gnd.n6752 gnd.n702 19.3944
R9312 gnd.n6756 gnd.n702 19.3944
R9313 gnd.n6756 gnd.n698 19.3944
R9314 gnd.n6762 gnd.n698 19.3944
R9315 gnd.n6762 gnd.n696 19.3944
R9316 gnd.n6766 gnd.n696 19.3944
R9317 gnd.n6766 gnd.n692 19.3944
R9318 gnd.n6772 gnd.n692 19.3944
R9319 gnd.n6772 gnd.n690 19.3944
R9320 gnd.n6776 gnd.n690 19.3944
R9321 gnd.n6776 gnd.n686 19.3944
R9322 gnd.n6782 gnd.n686 19.3944
R9323 gnd.n6782 gnd.n684 19.3944
R9324 gnd.n6786 gnd.n684 19.3944
R9325 gnd.n6786 gnd.n680 19.3944
R9326 gnd.n6792 gnd.n680 19.3944
R9327 gnd.n6792 gnd.n678 19.3944
R9328 gnd.n6796 gnd.n678 19.3944
R9329 gnd.n6796 gnd.n674 19.3944
R9330 gnd.n6802 gnd.n674 19.3944
R9331 gnd.n6802 gnd.n672 19.3944
R9332 gnd.n6806 gnd.n672 19.3944
R9333 gnd.n6806 gnd.n668 19.3944
R9334 gnd.n6812 gnd.n668 19.3944
R9335 gnd.n6812 gnd.n666 19.3944
R9336 gnd.n6816 gnd.n666 19.3944
R9337 gnd.n6816 gnd.n662 19.3944
R9338 gnd.n6822 gnd.n662 19.3944
R9339 gnd.n6822 gnd.n660 19.3944
R9340 gnd.n6826 gnd.n660 19.3944
R9341 gnd.n6826 gnd.n656 19.3944
R9342 gnd.n6832 gnd.n656 19.3944
R9343 gnd.n6832 gnd.n654 19.3944
R9344 gnd.n6836 gnd.n654 19.3944
R9345 gnd.n6836 gnd.n650 19.3944
R9346 gnd.n6842 gnd.n650 19.3944
R9347 gnd.n6842 gnd.n648 19.3944
R9348 gnd.n6846 gnd.n648 19.3944
R9349 gnd.n6846 gnd.n644 19.3944
R9350 gnd.n6852 gnd.n644 19.3944
R9351 gnd.n6852 gnd.n642 19.3944
R9352 gnd.n6856 gnd.n642 19.3944
R9353 gnd.n6856 gnd.n638 19.3944
R9354 gnd.n6862 gnd.n638 19.3944
R9355 gnd.n6862 gnd.n636 19.3944
R9356 gnd.n6866 gnd.n636 19.3944
R9357 gnd.n6866 gnd.n632 19.3944
R9358 gnd.n6872 gnd.n632 19.3944
R9359 gnd.n6872 gnd.n630 19.3944
R9360 gnd.n6876 gnd.n630 19.3944
R9361 gnd.n6876 gnd.n626 19.3944
R9362 gnd.n6882 gnd.n626 19.3944
R9363 gnd.n6882 gnd.n624 19.3944
R9364 gnd.n6886 gnd.n624 19.3944
R9365 gnd.n6886 gnd.n620 19.3944
R9366 gnd.n6892 gnd.n620 19.3944
R9367 gnd.n6892 gnd.n618 19.3944
R9368 gnd.n6896 gnd.n618 19.3944
R9369 gnd.n6896 gnd.n614 19.3944
R9370 gnd.n6902 gnd.n614 19.3944
R9371 gnd.n6902 gnd.n612 19.3944
R9372 gnd.n6906 gnd.n612 19.3944
R9373 gnd.n6906 gnd.n608 19.3944
R9374 gnd.n6912 gnd.n608 19.3944
R9375 gnd.n6912 gnd.n606 19.3944
R9376 gnd.n6916 gnd.n606 19.3944
R9377 gnd.n6916 gnd.n602 19.3944
R9378 gnd.n6922 gnd.n602 19.3944
R9379 gnd.n6922 gnd.n600 19.3944
R9380 gnd.n6926 gnd.n600 19.3944
R9381 gnd.n6926 gnd.n596 19.3944
R9382 gnd.n6932 gnd.n596 19.3944
R9383 gnd.n6932 gnd.n594 19.3944
R9384 gnd.n6936 gnd.n594 19.3944
R9385 gnd.n6936 gnd.n590 19.3944
R9386 gnd.n6942 gnd.n590 19.3944
R9387 gnd.n6942 gnd.n588 19.3944
R9388 gnd.n6946 gnd.n588 19.3944
R9389 gnd.n6946 gnd.n584 19.3944
R9390 gnd.n6952 gnd.n584 19.3944
R9391 gnd.n6952 gnd.n582 19.3944
R9392 gnd.n6956 gnd.n582 19.3944
R9393 gnd.n6956 gnd.n578 19.3944
R9394 gnd.n6962 gnd.n578 19.3944
R9395 gnd.n6962 gnd.n576 19.3944
R9396 gnd.n6966 gnd.n576 19.3944
R9397 gnd.n6966 gnd.n572 19.3944
R9398 gnd.n6972 gnd.n572 19.3944
R9399 gnd.n6972 gnd.n570 19.3944
R9400 gnd.n6976 gnd.n570 19.3944
R9401 gnd.n6976 gnd.n566 19.3944
R9402 gnd.n6982 gnd.n566 19.3944
R9403 gnd.n6982 gnd.n564 19.3944
R9404 gnd.n6986 gnd.n564 19.3944
R9405 gnd.n6986 gnd.n560 19.3944
R9406 gnd.n6992 gnd.n560 19.3944
R9407 gnd.n6992 gnd.n558 19.3944
R9408 gnd.n6996 gnd.n558 19.3944
R9409 gnd.n6996 gnd.n554 19.3944
R9410 gnd.n7002 gnd.n554 19.3944
R9411 gnd.n7002 gnd.n552 19.3944
R9412 gnd.n7006 gnd.n552 19.3944
R9413 gnd.n7006 gnd.n548 19.3944
R9414 gnd.n7012 gnd.n548 19.3944
R9415 gnd.n7012 gnd.n546 19.3944
R9416 gnd.n7016 gnd.n546 19.3944
R9417 gnd.n7016 gnd.n542 19.3944
R9418 gnd.n7022 gnd.n542 19.3944
R9419 gnd.n7022 gnd.n540 19.3944
R9420 gnd.n7026 gnd.n540 19.3944
R9421 gnd.n7026 gnd.n536 19.3944
R9422 gnd.n7032 gnd.n536 19.3944
R9423 gnd.n7032 gnd.n534 19.3944
R9424 gnd.n7036 gnd.n534 19.3944
R9425 gnd.n7036 gnd.n530 19.3944
R9426 gnd.n7042 gnd.n530 19.3944
R9427 gnd.n7042 gnd.n528 19.3944
R9428 gnd.n7046 gnd.n528 19.3944
R9429 gnd.n7046 gnd.n524 19.3944
R9430 gnd.n7052 gnd.n524 19.3944
R9431 gnd.n7052 gnd.n522 19.3944
R9432 gnd.n7056 gnd.n522 19.3944
R9433 gnd.n7056 gnd.n518 19.3944
R9434 gnd.n7062 gnd.n518 19.3944
R9435 gnd.n6078 gnd.n6077 19.3944
R9436 gnd.n6077 gnd.n6076 19.3944
R9437 gnd.n6076 gnd.n6075 19.3944
R9438 gnd.n6075 gnd.n6073 19.3944
R9439 gnd.n6073 gnd.n6070 19.3944
R9440 gnd.n6070 gnd.n6069 19.3944
R9441 gnd.n6069 gnd.n6066 19.3944
R9442 gnd.n6066 gnd.n6065 19.3944
R9443 gnd.n6065 gnd.n6062 19.3944
R9444 gnd.n6062 gnd.n6061 19.3944
R9445 gnd.n6061 gnd.n6058 19.3944
R9446 gnd.n6058 gnd.n6057 19.3944
R9447 gnd.n6057 gnd.n6054 19.3944
R9448 gnd.n6054 gnd.n6053 19.3944
R9449 gnd.n6053 gnd.n6050 19.3944
R9450 gnd.n6050 gnd.n6049 19.3944
R9451 gnd.n6049 gnd.n6046 19.3944
R9452 gnd.n6044 gnd.n6041 19.3944
R9453 gnd.n6041 gnd.n6040 19.3944
R9454 gnd.n6040 gnd.n6037 19.3944
R9455 gnd.n6037 gnd.n6036 19.3944
R9456 gnd.n6036 gnd.n6033 19.3944
R9457 gnd.n6033 gnd.n6032 19.3944
R9458 gnd.n6032 gnd.n6029 19.3944
R9459 gnd.n6027 gnd.n6024 19.3944
R9460 gnd.n6024 gnd.n6023 19.3944
R9461 gnd.n6023 gnd.n6020 19.3944
R9462 gnd.n6020 gnd.n6019 19.3944
R9463 gnd.n6019 gnd.n6016 19.3944
R9464 gnd.n6016 gnd.n6015 19.3944
R9465 gnd.n6015 gnd.n6012 19.3944
R9466 gnd.n6012 gnd.n6011 19.3944
R9467 gnd.n6007 gnd.n6004 19.3944
R9468 gnd.n6004 gnd.n6003 19.3944
R9469 gnd.n6003 gnd.n6000 19.3944
R9470 gnd.n6000 gnd.n5999 19.3944
R9471 gnd.n5999 gnd.n5996 19.3944
R9472 gnd.n5996 gnd.n5995 19.3944
R9473 gnd.n5995 gnd.n5992 19.3944
R9474 gnd.n5992 gnd.n5991 19.3944
R9475 gnd.n5991 gnd.n5988 19.3944
R9476 gnd.n5988 gnd.n5987 19.3944
R9477 gnd.n5987 gnd.n5984 19.3944
R9478 gnd.n5984 gnd.n5983 19.3944
R9479 gnd.n5983 gnd.n5980 19.3944
R9480 gnd.n5980 gnd.n5979 19.3944
R9481 gnd.n5979 gnd.n5976 19.3944
R9482 gnd.n5976 gnd.n5975 19.3944
R9483 gnd.n5975 gnd.n5972 19.3944
R9484 gnd.n5972 gnd.n5971 19.3944
R9485 gnd.n5955 gnd.n1472 19.3944
R9486 gnd.n5955 gnd.n5954 19.3944
R9487 gnd.n5954 gnd.n1481 19.3944
R9488 gnd.n5743 gnd.n1481 19.3944
R9489 gnd.n5746 gnd.n5743 19.3944
R9490 gnd.n5747 gnd.n5746 19.3944
R9491 gnd.n5752 gnd.n5747 19.3944
R9492 gnd.n5753 gnd.n5752 19.3944
R9493 gnd.n5757 gnd.n5753 19.3944
R9494 gnd.n5757 gnd.n5756 19.3944
R9495 gnd.n5756 gnd.n5755 19.3944
R9496 gnd.n5755 gnd.n1614 19.3944
R9497 gnd.n5832 gnd.n1614 19.3944
R9498 gnd.n5833 gnd.n5832 19.3944
R9499 gnd.n5835 gnd.n5833 19.3944
R9500 gnd.n5835 gnd.n1609 19.3944
R9501 gnd.n5847 gnd.n1609 19.3944
R9502 gnd.n5848 gnd.n5847 19.3944
R9503 gnd.n5850 gnd.n5848 19.3944
R9504 gnd.n5851 gnd.n5850 19.3944
R9505 gnd.n5857 gnd.n5851 19.3944
R9506 gnd.n5857 gnd.n5856 19.3944
R9507 gnd.n5856 gnd.n5855 19.3944
R9508 gnd.n5855 gnd.n5854 19.3944
R9509 gnd.n5854 gnd.n377 19.3944
R9510 gnd.n7292 gnd.n377 19.3944
R9511 gnd.n7294 gnd.n7292 19.3944
R9512 gnd.n7294 gnd.n7293 19.3944
R9513 gnd.n7293 gnd.n370 19.3944
R9514 gnd.n7343 gnd.n370 19.3944
R9515 gnd.n7343 gnd.n7342 19.3944
R9516 gnd.n7342 gnd.n7341 19.3944
R9517 gnd.n7341 gnd.n7339 19.3944
R9518 gnd.n7339 gnd.n7338 19.3944
R9519 gnd.n7338 gnd.n7336 19.3944
R9520 gnd.n7336 gnd.n7335 19.3944
R9521 gnd.n7335 gnd.n7333 19.3944
R9522 gnd.n7333 gnd.n7332 19.3944
R9523 gnd.n7332 gnd.n7330 19.3944
R9524 gnd.n7330 gnd.n7329 19.3944
R9525 gnd.n7329 gnd.n7327 19.3944
R9526 gnd.n7327 gnd.n7326 19.3944
R9527 gnd.n7326 gnd.n7324 19.3944
R9528 gnd.n7324 gnd.n7323 19.3944
R9529 gnd.n7323 gnd.n7321 19.3944
R9530 gnd.n7321 gnd.n7320 19.3944
R9531 gnd.n7320 gnd.n7318 19.3944
R9532 gnd.n7318 gnd.n7317 19.3944
R9533 gnd.n7317 gnd.n7315 19.3944
R9534 gnd.n7315 gnd.n7314 19.3944
R9535 gnd.n7314 gnd.n7312 19.3944
R9536 gnd.n7312 gnd.n7311 19.3944
R9537 gnd.n7311 gnd.n7309 19.3944
R9538 gnd.n5958 gnd.n5957 19.3944
R9539 gnd.n5957 gnd.n1479 19.3944
R9540 gnd.n1503 gnd.n1479 19.3944
R9541 gnd.n5944 gnd.n1503 19.3944
R9542 gnd.n5944 gnd.n5943 19.3944
R9543 gnd.n5943 gnd.n5942 19.3944
R9544 gnd.n5942 gnd.n1508 19.3944
R9545 gnd.n5932 gnd.n1508 19.3944
R9546 gnd.n5932 gnd.n5931 19.3944
R9547 gnd.n5931 gnd.n5930 19.3944
R9548 gnd.n5930 gnd.n1528 19.3944
R9549 gnd.n5920 gnd.n1528 19.3944
R9550 gnd.n5920 gnd.n5919 19.3944
R9551 gnd.n5919 gnd.n5918 19.3944
R9552 gnd.n5918 gnd.n1548 19.3944
R9553 gnd.n5908 gnd.n1548 19.3944
R9554 gnd.n5908 gnd.n5907 19.3944
R9555 gnd.n5907 gnd.n5906 19.3944
R9556 gnd.n5906 gnd.n1568 19.3944
R9557 gnd.n5896 gnd.n1568 19.3944
R9558 gnd.n5896 gnd.n5895 19.3944
R9559 gnd.n5895 gnd.n5894 19.3944
R9560 gnd.n5894 gnd.n1588 19.3944
R9561 gnd.n1588 gnd.n379 19.3944
R9562 gnd.n7289 gnd.n379 19.3944
R9563 gnd.n7289 gnd.n372 19.3944
R9564 gnd.n7298 gnd.n372 19.3944
R9565 gnd.n7299 gnd.n7298 19.3944
R9566 gnd.n7301 gnd.n7299 19.3944
R9567 gnd.n7301 gnd.n110 19.3944
R9568 gnd.n7601 gnd.n110 19.3944
R9569 gnd.n7601 gnd.n7600 19.3944
R9570 gnd.n7600 gnd.n7599 19.3944
R9571 gnd.n7599 gnd.n114 19.3944
R9572 gnd.n7589 gnd.n114 19.3944
R9573 gnd.n7589 gnd.n7588 19.3944
R9574 gnd.n7588 gnd.n7587 19.3944
R9575 gnd.n7587 gnd.n131 19.3944
R9576 gnd.n7577 gnd.n131 19.3944
R9577 gnd.n7577 gnd.n7576 19.3944
R9578 gnd.n7576 gnd.n7575 19.3944
R9579 gnd.n7575 gnd.n151 19.3944
R9580 gnd.n7565 gnd.n151 19.3944
R9581 gnd.n7565 gnd.n7564 19.3944
R9582 gnd.n7564 gnd.n7563 19.3944
R9583 gnd.n7563 gnd.n169 19.3944
R9584 gnd.n7553 gnd.n169 19.3944
R9585 gnd.n7553 gnd.n7552 19.3944
R9586 gnd.n7552 gnd.n7551 19.3944
R9587 gnd.n7551 gnd.n189 19.3944
R9588 gnd.n7541 gnd.n189 19.3944
R9589 gnd.n7541 gnd.n7540 19.3944
R9590 gnd.n7540 gnd.n7539 19.3944
R9591 gnd.n7461 gnd.n279 19.3944
R9592 gnd.n7461 gnd.n283 19.3944
R9593 gnd.n286 gnd.n283 19.3944
R9594 gnd.n7454 gnd.n286 19.3944
R9595 gnd.n7454 gnd.n7453 19.3944
R9596 gnd.n7453 gnd.n7452 19.3944
R9597 gnd.n7452 gnd.n292 19.3944
R9598 gnd.n7447 gnd.n292 19.3944
R9599 gnd.n7447 gnd.n7446 19.3944
R9600 gnd.n7446 gnd.n7445 19.3944
R9601 gnd.n7445 gnd.n299 19.3944
R9602 gnd.n7440 gnd.n299 19.3944
R9603 gnd.n7440 gnd.n7439 19.3944
R9604 gnd.n7439 gnd.n7438 19.3944
R9605 gnd.n7438 gnd.n306 19.3944
R9606 gnd.n7433 gnd.n306 19.3944
R9607 gnd.n7433 gnd.n7432 19.3944
R9608 gnd.n7432 gnd.n7431 19.3944
R9609 gnd.n7499 gnd.n246 19.3944
R9610 gnd.n7494 gnd.n246 19.3944
R9611 gnd.n7494 gnd.n7493 19.3944
R9612 gnd.n7493 gnd.n7492 19.3944
R9613 gnd.n7492 gnd.n253 19.3944
R9614 gnd.n7487 gnd.n253 19.3944
R9615 gnd.n7487 gnd.n7486 19.3944
R9616 gnd.n7486 gnd.n7485 19.3944
R9617 gnd.n7485 gnd.n260 19.3944
R9618 gnd.n7480 gnd.n260 19.3944
R9619 gnd.n7480 gnd.n7479 19.3944
R9620 gnd.n7479 gnd.n7478 19.3944
R9621 gnd.n7478 gnd.n267 19.3944
R9622 gnd.n7473 gnd.n267 19.3944
R9623 gnd.n7473 gnd.n7472 19.3944
R9624 gnd.n7472 gnd.n7471 19.3944
R9625 gnd.n7471 gnd.n274 19.3944
R9626 gnd.n7466 gnd.n274 19.3944
R9627 gnd.n7532 gnd.n7531 19.3944
R9628 gnd.n7531 gnd.n7530 19.3944
R9629 gnd.n7530 gnd.n218 19.3944
R9630 gnd.n7525 gnd.n218 19.3944
R9631 gnd.n7525 gnd.n7524 19.3944
R9632 gnd.n7524 gnd.n7523 19.3944
R9633 gnd.n7523 gnd.n225 19.3944
R9634 gnd.n7518 gnd.n225 19.3944
R9635 gnd.n7518 gnd.n7517 19.3944
R9636 gnd.n7517 gnd.n7516 19.3944
R9637 gnd.n7516 gnd.n232 19.3944
R9638 gnd.n7511 gnd.n232 19.3944
R9639 gnd.n7511 gnd.n7510 19.3944
R9640 gnd.n7510 gnd.n7509 19.3944
R9641 gnd.n7509 gnd.n239 19.3944
R9642 gnd.n7504 gnd.n239 19.3944
R9643 gnd.n7504 gnd.n7503 19.3944
R9644 gnd.n7422 gnd.n7421 19.3944
R9645 gnd.n7421 gnd.n7420 19.3944
R9646 gnd.n7420 gnd.n321 19.3944
R9647 gnd.n7415 gnd.n321 19.3944
R9648 gnd.n7415 gnd.n7414 19.3944
R9649 gnd.n7414 gnd.n7413 19.3944
R9650 gnd.n7413 gnd.n328 19.3944
R9651 gnd.n7408 gnd.n328 19.3944
R9652 gnd.n7408 gnd.n7407 19.3944
R9653 gnd.n7407 gnd.n7406 19.3944
R9654 gnd.n7406 gnd.n335 19.3944
R9655 gnd.n7401 gnd.n335 19.3944
R9656 gnd.n7401 gnd.n7400 19.3944
R9657 gnd.n7400 gnd.n7399 19.3944
R9658 gnd.n7399 gnd.n342 19.3944
R9659 gnd.n7394 gnd.n342 19.3944
R9660 gnd.n5774 gnd.n1633 19.3944
R9661 gnd.n5774 gnd.n1634 19.3944
R9662 gnd.n5770 gnd.n1634 19.3944
R9663 gnd.n5770 gnd.n5769 19.3944
R9664 gnd.n5769 gnd.n5768 19.3944
R9665 gnd.n5768 gnd.n5740 19.3944
R9666 gnd.n5764 gnd.n5740 19.3944
R9667 gnd.n5764 gnd.n5763 19.3944
R9668 gnd.n5763 gnd.n5762 19.3944
R9669 gnd.n5762 gnd.n1617 19.3944
R9670 gnd.n5824 gnd.n1617 19.3944
R9671 gnd.n5824 gnd.n1615 19.3944
R9672 gnd.n5828 gnd.n1615 19.3944
R9673 gnd.n5828 gnd.n1612 19.3944
R9674 gnd.n5839 gnd.n1612 19.3944
R9675 gnd.n5839 gnd.n1610 19.3944
R9676 gnd.n5843 gnd.n1610 19.3944
R9677 gnd.n5843 gnd.n1605 19.3944
R9678 gnd.n5873 gnd.n1605 19.3944
R9679 gnd.n5873 gnd.n1606 19.3944
R9680 gnd.n5869 gnd.n1606 19.3944
R9681 gnd.n5869 gnd.n5868 19.3944
R9682 gnd.n5868 gnd.n5867 19.3944
R9683 gnd.n5867 gnd.n5862 19.3944
R9684 gnd.n5863 gnd.n5862 19.3944
R9685 gnd.n5863 gnd.n85 19.3944
R9686 gnd.n7614 gnd.n85 19.3944
R9687 gnd.n7614 gnd.n7613 19.3944
R9688 gnd.n7613 gnd.n87 19.3944
R9689 gnd.n7347 gnd.n87 19.3944
R9690 gnd.n7351 gnd.n7347 19.3944
R9691 gnd.n7353 gnd.n7351 19.3944
R9692 gnd.n7354 gnd.n7353 19.3944
R9693 gnd.n7354 gnd.n366 19.3944
R9694 gnd.n7358 gnd.n366 19.3944
R9695 gnd.n7360 gnd.n7358 19.3944
R9696 gnd.n7361 gnd.n7360 19.3944
R9697 gnd.n7361 gnd.n363 19.3944
R9698 gnd.n7365 gnd.n363 19.3944
R9699 gnd.n7367 gnd.n7365 19.3944
R9700 gnd.n7368 gnd.n7367 19.3944
R9701 gnd.n7368 gnd.n360 19.3944
R9702 gnd.n7372 gnd.n360 19.3944
R9703 gnd.n7374 gnd.n7372 19.3944
R9704 gnd.n7375 gnd.n7374 19.3944
R9705 gnd.n7375 gnd.n357 19.3944
R9706 gnd.n7379 gnd.n357 19.3944
R9707 gnd.n7381 gnd.n7379 19.3944
R9708 gnd.n7382 gnd.n7381 19.3944
R9709 gnd.n7382 gnd.n354 19.3944
R9710 gnd.n7386 gnd.n354 19.3944
R9711 gnd.n7388 gnd.n7386 19.3944
R9712 gnd.n7389 gnd.n7388 19.3944
R9713 gnd.n1489 gnd.n1488 19.3944
R9714 gnd.n5950 gnd.n1488 19.3944
R9715 gnd.n5950 gnd.n5949 19.3944
R9716 gnd.n5949 gnd.n5948 19.3944
R9717 gnd.n5948 gnd.n1495 19.3944
R9718 gnd.n5938 gnd.n1495 19.3944
R9719 gnd.n5938 gnd.n5937 19.3944
R9720 gnd.n5937 gnd.n5936 19.3944
R9721 gnd.n5936 gnd.n1518 19.3944
R9722 gnd.n5926 gnd.n1518 19.3944
R9723 gnd.n5926 gnd.n5925 19.3944
R9724 gnd.n5925 gnd.n5924 19.3944
R9725 gnd.n5924 gnd.n1539 19.3944
R9726 gnd.n5914 gnd.n1539 19.3944
R9727 gnd.n5914 gnd.n5913 19.3944
R9728 gnd.n5913 gnd.n5912 19.3944
R9729 gnd.n5912 gnd.n1558 19.3944
R9730 gnd.n5902 gnd.n1558 19.3944
R9731 gnd.n5902 gnd.n5901 19.3944
R9732 gnd.n5901 gnd.n5900 19.3944
R9733 gnd.n5900 gnd.n1579 19.3944
R9734 gnd.n5890 gnd.n1579 19.3944
R9735 gnd.n1593 gnd.n100 19.3944
R9736 gnd.n7285 gnd.n100 19.3944
R9737 gnd.n386 gnd.n385 19.3944
R9738 gnd.n7609 gnd.n7608 19.3944
R9739 gnd.n7605 gnd.n95 19.3944
R9740 gnd.n7605 gnd.n102 19.3944
R9741 gnd.n7595 gnd.n102 19.3944
R9742 gnd.n7595 gnd.n7594 19.3944
R9743 gnd.n7594 gnd.n7593 19.3944
R9744 gnd.n7593 gnd.n122 19.3944
R9745 gnd.n7583 gnd.n122 19.3944
R9746 gnd.n7583 gnd.n7582 19.3944
R9747 gnd.n7582 gnd.n7581 19.3944
R9748 gnd.n7581 gnd.n142 19.3944
R9749 gnd.n7571 gnd.n142 19.3944
R9750 gnd.n7571 gnd.n7570 19.3944
R9751 gnd.n7570 gnd.n7569 19.3944
R9752 gnd.n7569 gnd.n160 19.3944
R9753 gnd.n7559 gnd.n160 19.3944
R9754 gnd.n7559 gnd.n7558 19.3944
R9755 gnd.n7558 gnd.n7557 19.3944
R9756 gnd.n7557 gnd.n180 19.3944
R9757 gnd.n7547 gnd.n180 19.3944
R9758 gnd.n7547 gnd.n7546 19.3944
R9759 gnd.n7546 gnd.n7545 19.3944
R9760 gnd.n7545 gnd.n200 19.3944
R9761 gnd.n7535 gnd.n200 19.3944
R9762 gnd.n4354 gnd.n4353 19.3944
R9763 gnd.n4353 gnd.n4352 19.3944
R9764 gnd.n4352 gnd.n4351 19.3944
R9765 gnd.n4351 gnd.n4349 19.3944
R9766 gnd.n4349 gnd.n4346 19.3944
R9767 gnd.n4346 gnd.n4345 19.3944
R9768 gnd.n4345 gnd.n4342 19.3944
R9769 gnd.n4342 gnd.n4341 19.3944
R9770 gnd.n4341 gnd.n4338 19.3944
R9771 gnd.n4338 gnd.n4337 19.3944
R9772 gnd.n4337 gnd.n4334 19.3944
R9773 gnd.n4334 gnd.n4333 19.3944
R9774 gnd.n4333 gnd.n4330 19.3944
R9775 gnd.n4330 gnd.n4329 19.3944
R9776 gnd.n4329 gnd.n4326 19.3944
R9777 gnd.n4326 gnd.n4325 19.3944
R9778 gnd.n4325 gnd.n4322 19.3944
R9779 gnd.n4320 gnd.n4317 19.3944
R9780 gnd.n4317 gnd.n4316 19.3944
R9781 gnd.n4316 gnd.n4313 19.3944
R9782 gnd.n4313 gnd.n4312 19.3944
R9783 gnd.n4312 gnd.n4309 19.3944
R9784 gnd.n4309 gnd.n4308 19.3944
R9785 gnd.n4308 gnd.n4305 19.3944
R9786 gnd.n4305 gnd.n4304 19.3944
R9787 gnd.n4304 gnd.n4301 19.3944
R9788 gnd.n4301 gnd.n4300 19.3944
R9789 gnd.n4300 gnd.n4297 19.3944
R9790 gnd.n4297 gnd.n4296 19.3944
R9791 gnd.n4296 gnd.n4293 19.3944
R9792 gnd.n4293 gnd.n4292 19.3944
R9793 gnd.n4292 gnd.n4289 19.3944
R9794 gnd.n4289 gnd.n4288 19.3944
R9795 gnd.n4288 gnd.n4285 19.3944
R9796 gnd.n4285 gnd.n4284 19.3944
R9797 gnd.n4280 gnd.n4277 19.3944
R9798 gnd.n4277 gnd.n4276 19.3944
R9799 gnd.n4276 gnd.n4273 19.3944
R9800 gnd.n4273 gnd.n4272 19.3944
R9801 gnd.n4272 gnd.n4269 19.3944
R9802 gnd.n4269 gnd.n4268 19.3944
R9803 gnd.n4268 gnd.n4265 19.3944
R9804 gnd.n4265 gnd.n4264 19.3944
R9805 gnd.n4264 gnd.n4261 19.3944
R9806 gnd.n4261 gnd.n4260 19.3944
R9807 gnd.n4260 gnd.n4257 19.3944
R9808 gnd.n4257 gnd.n4256 19.3944
R9809 gnd.n4256 gnd.n4253 19.3944
R9810 gnd.n4253 gnd.n4252 19.3944
R9811 gnd.n4252 gnd.n4249 19.3944
R9812 gnd.n4249 gnd.n4248 19.3944
R9813 gnd.n4248 gnd.n4245 19.3944
R9814 gnd.n4245 gnd.n4244 19.3944
R9815 gnd.n4237 gnd.n4235 19.3944
R9816 gnd.n4235 gnd.n4232 19.3944
R9817 gnd.n4232 gnd.n4231 19.3944
R9818 gnd.n4231 gnd.n4228 19.3944
R9819 gnd.n4228 gnd.n4227 19.3944
R9820 gnd.n4227 gnd.n4224 19.3944
R9821 gnd.n4224 gnd.n4223 19.3944
R9822 gnd.n4223 gnd.n4220 19.3944
R9823 gnd.n4220 gnd.n4219 19.3944
R9824 gnd.n4219 gnd.n4216 19.3944
R9825 gnd.n4216 gnd.n4215 19.3944
R9826 gnd.n4215 gnd.n4212 19.3944
R9827 gnd.n4212 gnd.n4211 19.3944
R9828 gnd.n4211 gnd.n4208 19.3944
R9829 gnd.n4208 gnd.n4207 19.3944
R9830 gnd.n4207 gnd.n4204 19.3944
R9831 gnd.n4198 gnd.n4196 19.3944
R9832 gnd.n4196 gnd.n4195 19.3944
R9833 gnd.n4195 gnd.n4193 19.3944
R9834 gnd.n4193 gnd.n4192 19.3944
R9835 gnd.n4192 gnd.n4190 19.3944
R9836 gnd.n4190 gnd.n4189 19.3944
R9837 gnd.n4189 gnd.n4187 19.3944
R9838 gnd.n4187 gnd.n4186 19.3944
R9839 gnd.n4186 gnd.n4184 19.3944
R9840 gnd.n4184 gnd.n4183 19.3944
R9841 gnd.n4183 gnd.n4181 19.3944
R9842 gnd.n4181 gnd.n4180 19.3944
R9843 gnd.n4180 gnd.n4178 19.3944
R9844 gnd.n4178 gnd.n2486 19.3944
R9845 gnd.n4443 gnd.n2486 19.3944
R9846 gnd.n4443 gnd.n2484 19.3944
R9847 gnd.n4459 gnd.n2484 19.3944
R9848 gnd.n4459 gnd.n4458 19.3944
R9849 gnd.n4458 gnd.n4457 19.3944
R9850 gnd.n4457 gnd.n4455 19.3944
R9851 gnd.n4455 gnd.n4454 19.3944
R9852 gnd.n4454 gnd.n4452 19.3944
R9853 gnd.n4452 gnd.n2450 19.3944
R9854 gnd.n4504 gnd.n2450 19.3944
R9855 gnd.n4504 gnd.n2448 19.3944
R9856 gnd.n4514 gnd.n2448 19.3944
R9857 gnd.n4514 gnd.n4513 19.3944
R9858 gnd.n4513 gnd.n4509 19.3944
R9859 gnd.n4509 gnd.n2420 19.3944
R9860 gnd.n4567 gnd.n2420 19.3944
R9861 gnd.n4567 gnd.n2418 19.3944
R9862 gnd.n4571 gnd.n2418 19.3944
R9863 gnd.n4571 gnd.n2415 19.3944
R9864 gnd.n4582 gnd.n2415 19.3944
R9865 gnd.n4582 gnd.n2413 19.3944
R9866 gnd.n4586 gnd.n2413 19.3944
R9867 gnd.n4586 gnd.n2404 19.3944
R9868 gnd.n4622 gnd.n2404 19.3944
R9869 gnd.n4622 gnd.n2405 19.3944
R9870 gnd.n4618 gnd.n2405 19.3944
R9871 gnd.n4618 gnd.n4617 19.3944
R9872 gnd.n4617 gnd.n4616 19.3944
R9873 gnd.n4616 gnd.n2410 19.3944
R9874 gnd.n4612 gnd.n2410 19.3944
R9875 gnd.n4612 gnd.n4611 19.3944
R9876 gnd.n4611 gnd.n4610 19.3944
R9877 gnd.n4610 gnd.n2388 19.3944
R9878 gnd.n4680 gnd.n2388 19.3944
R9879 gnd.n4680 gnd.n2386 19.3944
R9880 gnd.n4685 gnd.n2386 19.3944
R9881 gnd.n4685 gnd.n2382 19.3944
R9882 gnd.n4696 gnd.n2382 19.3944
R9883 gnd.n4697 gnd.n4696 19.3944
R9884 gnd.n4363 gnd.n4361 19.3944
R9885 gnd.n4363 gnd.n4362 19.3944
R9886 gnd.n4362 gnd.n2541 19.3944
R9887 gnd.n4378 gnd.n2541 19.3944
R9888 gnd.n4379 gnd.n4378 19.3944
R9889 gnd.n4380 gnd.n4379 19.3944
R9890 gnd.n4380 gnd.n2523 19.3944
R9891 gnd.n4398 gnd.n2523 19.3944
R9892 gnd.n4399 gnd.n4398 19.3944
R9893 gnd.n4400 gnd.n4399 19.3944
R9894 gnd.n4400 gnd.n2505 19.3944
R9895 gnd.n4418 gnd.n2505 19.3944
R9896 gnd.n4419 gnd.n4418 19.3944
R9897 gnd.n4421 gnd.n4419 19.3944
R9898 gnd.n4422 gnd.n4421 19.3944
R9899 gnd.n4422 gnd.n2479 19.3944
R9900 gnd.n4463 gnd.n2479 19.3944
R9901 gnd.n4464 gnd.n4463 19.3944
R9902 gnd.n4465 gnd.n4464 19.3944
R9903 gnd.n4465 gnd.n2462 19.3944
R9904 gnd.n4484 gnd.n2462 19.3944
R9905 gnd.n4485 gnd.n4484 19.3944
R9906 gnd.n4486 gnd.n4485 19.3944
R9907 gnd.n4488 gnd.n4486 19.3944
R9908 gnd.n4488 gnd.n2446 19.3944
R9909 gnd.n4518 gnd.n2446 19.3944
R9910 gnd.n4519 gnd.n4518 19.3944
R9911 gnd.n4521 gnd.n4519 19.3944
R9912 gnd.n4523 gnd.n4521 19.3944
R9913 gnd.n4523 gnd.n4522 19.3944
R9914 gnd.n4522 gnd.n2417 19.3944
R9915 gnd.n4575 gnd.n2417 19.3944
R9916 gnd.n4576 gnd.n4575 19.3944
R9917 gnd.n4578 gnd.n4576 19.3944
R9918 gnd.n4578 gnd.n2412 19.3944
R9919 gnd.n4590 gnd.n2412 19.3944
R9920 gnd.n4591 gnd.n4590 19.3944
R9921 gnd.n4593 gnd.n4591 19.3944
R9922 gnd.n4594 gnd.n4593 19.3944
R9923 gnd.n4597 gnd.n4594 19.3944
R9924 gnd.n4598 gnd.n4597 19.3944
R9925 gnd.n4603 gnd.n4598 19.3944
R9926 gnd.n4604 gnd.n4603 19.3944
R9927 gnd.n4605 gnd.n4604 19.3944
R9928 gnd.n4605 gnd.n2389 19.3944
R9929 gnd.n4674 gnd.n2389 19.3944
R9930 gnd.n4675 gnd.n4674 19.3944
R9931 gnd.n4676 gnd.n4675 19.3944
R9932 gnd.n4676 gnd.n2384 19.3944
R9933 gnd.n4689 gnd.n2384 19.3944
R9934 gnd.n4690 gnd.n4689 19.3944
R9935 gnd.n4692 gnd.n4690 19.3944
R9936 gnd.n4692 gnd.n4691 19.3944
R9937 gnd.n4365 gnd.n2557 19.3944
R9938 gnd.n4365 gnd.n2558 19.3944
R9939 gnd.n2560 gnd.n2558 19.3944
R9940 gnd.n2560 gnd.n2539 19.3944
R9941 gnd.n4385 gnd.n2539 19.3944
R9942 gnd.n4385 gnd.n4384 19.3944
R9943 gnd.n4384 gnd.n4383 19.3944
R9944 gnd.n4383 gnd.n2521 19.3944
R9945 gnd.n4405 gnd.n2521 19.3944
R9946 gnd.n4405 gnd.n4404 19.3944
R9947 gnd.n4404 gnd.n4403 19.3944
R9948 gnd.n4403 gnd.n2502 19.3944
R9949 gnd.n4429 gnd.n2502 19.3944
R9950 gnd.n4429 gnd.n4428 19.3944
R9951 gnd.n4428 gnd.n4427 19.3944
R9952 gnd.n4427 gnd.n4426 19.3944
R9953 gnd.n4426 gnd.n2477 19.3944
R9954 gnd.n4470 gnd.n2477 19.3944
R9955 gnd.n4470 gnd.n4469 19.3944
R9956 gnd.n4469 gnd.n4468 19.3944
R9957 gnd.n4468 gnd.n2459 19.3944
R9958 gnd.n4495 gnd.n2459 19.3944
R9959 gnd.n4495 gnd.n4494 19.3944
R9960 gnd.n4494 gnd.n4493 19.3944
R9961 gnd.n4493 gnd.n4491 19.3944
R9962 gnd.n4491 gnd.n2442 19.3944
R9963 gnd.n4527 gnd.n2442 19.3944
R9964 gnd.n4527 gnd.n4526 19.3944
R9965 gnd.n4526 gnd.n4525 19.3944
R9966 gnd.n4525 gnd.n961 19.3944
R9967 gnd.n6462 gnd.n961 19.3944
R9968 gnd.n6462 gnd.n6461 19.3944
R9969 gnd.n6461 gnd.n6460 19.3944
R9970 gnd.n6460 gnd.n965 19.3944
R9971 gnd.n6450 gnd.n965 19.3944
R9972 gnd.n6450 gnd.n6449 19.3944
R9973 gnd.n6449 gnd.n6448 19.3944
R9974 gnd.n6448 gnd.n984 19.3944
R9975 gnd.n6438 gnd.n984 19.3944
R9976 gnd.n6438 gnd.n6437 19.3944
R9977 gnd.n6437 gnd.n6436 19.3944
R9978 gnd.n6436 gnd.n1004 19.3944
R9979 gnd.n6426 gnd.n1004 19.3944
R9980 gnd.n6426 gnd.n6425 19.3944
R9981 gnd.n6425 gnd.n6424 19.3944
R9982 gnd.n6424 gnd.n1024 19.3944
R9983 gnd.n6414 gnd.n1024 19.3944
R9984 gnd.n6414 gnd.n6413 19.3944
R9985 gnd.n6413 gnd.n6412 19.3944
R9986 gnd.n6412 gnd.n1044 19.3944
R9987 gnd.n6402 gnd.n1044 19.3944
R9988 gnd.n6402 gnd.n6401 19.3944
R9989 gnd.n6401 gnd.n6400 19.3944
R9990 gnd.n6393 gnd.n6392 19.3944
R9991 gnd.n6392 gnd.n1072 19.3944
R9992 gnd.n1074 gnd.n1072 19.3944
R9993 gnd.n6385 gnd.n1074 19.3944
R9994 gnd.n6385 gnd.n6384 19.3944
R9995 gnd.n6384 gnd.n6383 19.3944
R9996 gnd.n6383 gnd.n1081 19.3944
R9997 gnd.n6378 gnd.n1081 19.3944
R9998 gnd.n6378 gnd.n6377 19.3944
R9999 gnd.n6377 gnd.n6376 19.3944
R10000 gnd.n6376 gnd.n1088 19.3944
R10001 gnd.n6371 gnd.n1088 19.3944
R10002 gnd.n6371 gnd.n6370 19.3944
R10003 gnd.n6370 gnd.n6369 19.3944
R10004 gnd.n6369 gnd.n1095 19.3944
R10005 gnd.n6364 gnd.n1095 19.3944
R10006 gnd.n6364 gnd.n6363 19.3944
R10007 gnd.n2254 gnd.n2214 19.3944
R10008 gnd.n2258 gnd.n2214 19.3944
R10009 gnd.n2258 gnd.n2212 19.3944
R10010 gnd.n2264 gnd.n2212 19.3944
R10011 gnd.n2264 gnd.n2210 19.3944
R10012 gnd.n2268 gnd.n2210 19.3944
R10013 gnd.n2268 gnd.n2208 19.3944
R10014 gnd.n2274 gnd.n2208 19.3944
R10015 gnd.n2274 gnd.n2206 19.3944
R10016 gnd.n2278 gnd.n2206 19.3944
R10017 gnd.n2278 gnd.n2204 19.3944
R10018 gnd.n2284 gnd.n2204 19.3944
R10019 gnd.n2284 gnd.n2202 19.3944
R10020 gnd.n2288 gnd.n2202 19.3944
R10021 gnd.n2288 gnd.n2200 19.3944
R10022 gnd.n2294 gnd.n2200 19.3944
R10023 gnd.n2294 gnd.n2198 19.3944
R10024 gnd.n2298 gnd.n2198 19.3944
R10025 gnd.n2227 gnd.n1117 19.3944
R10026 gnd.n2234 gnd.n2227 19.3944
R10027 gnd.n2234 gnd.n2224 19.3944
R10028 gnd.n2238 gnd.n2224 19.3944
R10029 gnd.n2238 gnd.n2222 19.3944
R10030 gnd.n2244 gnd.n2222 19.3944
R10031 gnd.n2244 gnd.n2220 19.3944
R10032 gnd.n2248 gnd.n2220 19.3944
R10033 gnd.n6361 gnd.n1104 19.3944
R10034 gnd.n6356 gnd.n1104 19.3944
R10035 gnd.n6356 gnd.n6355 19.3944
R10036 gnd.n6355 gnd.n6354 19.3944
R10037 gnd.n6354 gnd.n1111 19.3944
R10038 gnd.n6349 gnd.n1111 19.3944
R10039 gnd.n6349 gnd.n6348 19.3944
R10040 gnd.n4369 gnd.n2550 19.3944
R10041 gnd.n4369 gnd.n2548 19.3944
R10042 gnd.n4373 gnd.n2548 19.3944
R10043 gnd.n4373 gnd.n2531 19.3944
R10044 gnd.n4389 gnd.n2531 19.3944
R10045 gnd.n4389 gnd.n2529 19.3944
R10046 gnd.n4393 gnd.n2529 19.3944
R10047 gnd.n4393 gnd.n2514 19.3944
R10048 gnd.n4409 gnd.n2514 19.3944
R10049 gnd.n4409 gnd.n2512 19.3944
R10050 gnd.n4413 gnd.n2512 19.3944
R10051 gnd.n4413 gnd.n2494 19.3944
R10052 gnd.n4433 gnd.n2494 19.3944
R10053 gnd.n4433 gnd.n2492 19.3944
R10054 gnd.n4439 gnd.n2492 19.3944
R10055 gnd.n4439 gnd.n4438 19.3944
R10056 gnd.n4438 gnd.n2470 19.3944
R10057 gnd.n4474 gnd.n2470 19.3944
R10058 gnd.n4474 gnd.n2468 19.3944
R10059 gnd.n4479 gnd.n2468 19.3944
R10060 gnd.n4479 gnd.n4478 19.3944
R10061 gnd.n4478 gnd.n2455 19.3944
R10062 gnd.n4499 gnd.n944 19.3944
R10063 gnd.n6469 gnd.n944 19.3944
R10064 gnd.n2435 gnd.n945 19.3944
R10065 gnd.n4533 gnd.n4532 19.3944
R10066 gnd.n6466 gnd.n952 19.3944
R10067 gnd.n6466 gnd.n953 19.3944
R10068 gnd.n6456 gnd.n953 19.3944
R10069 gnd.n6456 gnd.n6455 19.3944
R10070 gnd.n6455 gnd.n6454 19.3944
R10071 gnd.n6454 gnd.n974 19.3944
R10072 gnd.n6444 gnd.n974 19.3944
R10073 gnd.n6444 gnd.n6443 19.3944
R10074 gnd.n6443 gnd.n6442 19.3944
R10075 gnd.n6442 gnd.n995 19.3944
R10076 gnd.n6432 gnd.n995 19.3944
R10077 gnd.n6432 gnd.n6431 19.3944
R10078 gnd.n6431 gnd.n6430 19.3944
R10079 gnd.n6430 gnd.n1014 19.3944
R10080 gnd.n6420 gnd.n1014 19.3944
R10081 gnd.n6420 gnd.n6419 19.3944
R10082 gnd.n6419 gnd.n6418 19.3944
R10083 gnd.n6418 gnd.n1035 19.3944
R10084 gnd.n6408 gnd.n1035 19.3944
R10085 gnd.n6408 gnd.n6407 19.3944
R10086 gnd.n6407 gnd.n6406 19.3944
R10087 gnd.n6406 gnd.n1055 19.3944
R10088 gnd.n6396 gnd.n1055 19.3944
R10089 gnd.n6642 gnd.n770 19.3944
R10090 gnd.n6636 gnd.n770 19.3944
R10091 gnd.n6636 gnd.n6635 19.3944
R10092 gnd.n6635 gnd.n6634 19.3944
R10093 gnd.n6634 gnd.n777 19.3944
R10094 gnd.n6628 gnd.n777 19.3944
R10095 gnd.n6628 gnd.n6627 19.3944
R10096 gnd.n6627 gnd.n6626 19.3944
R10097 gnd.n6626 gnd.n785 19.3944
R10098 gnd.n6620 gnd.n785 19.3944
R10099 gnd.n6620 gnd.n6619 19.3944
R10100 gnd.n6619 gnd.n6618 19.3944
R10101 gnd.n6618 gnd.n793 19.3944
R10102 gnd.n6612 gnd.n793 19.3944
R10103 gnd.n6612 gnd.n6611 19.3944
R10104 gnd.n6611 gnd.n6610 19.3944
R10105 gnd.n6610 gnd.n801 19.3944
R10106 gnd.n6604 gnd.n801 19.3944
R10107 gnd.n6604 gnd.n6603 19.3944
R10108 gnd.n6603 gnd.n6602 19.3944
R10109 gnd.n6602 gnd.n809 19.3944
R10110 gnd.n6596 gnd.n809 19.3944
R10111 gnd.n6596 gnd.n6595 19.3944
R10112 gnd.n6595 gnd.n6594 19.3944
R10113 gnd.n6594 gnd.n817 19.3944
R10114 gnd.n6588 gnd.n817 19.3944
R10115 gnd.n6588 gnd.n6587 19.3944
R10116 gnd.n6587 gnd.n6586 19.3944
R10117 gnd.n6586 gnd.n825 19.3944
R10118 gnd.n6580 gnd.n825 19.3944
R10119 gnd.n6580 gnd.n6579 19.3944
R10120 gnd.n6579 gnd.n6578 19.3944
R10121 gnd.n6578 gnd.n833 19.3944
R10122 gnd.n6572 gnd.n833 19.3944
R10123 gnd.n6572 gnd.n6571 19.3944
R10124 gnd.n6571 gnd.n6570 19.3944
R10125 gnd.n6570 gnd.n841 19.3944
R10126 gnd.n6564 gnd.n841 19.3944
R10127 gnd.n6564 gnd.n6563 19.3944
R10128 gnd.n6563 gnd.n6562 19.3944
R10129 gnd.n6562 gnd.n849 19.3944
R10130 gnd.n6556 gnd.n849 19.3944
R10131 gnd.n6556 gnd.n6555 19.3944
R10132 gnd.n6555 gnd.n6554 19.3944
R10133 gnd.n6554 gnd.n857 19.3944
R10134 gnd.n6548 gnd.n857 19.3944
R10135 gnd.n6548 gnd.n6547 19.3944
R10136 gnd.n6547 gnd.n6546 19.3944
R10137 gnd.n6546 gnd.n865 19.3944
R10138 gnd.n6540 gnd.n865 19.3944
R10139 gnd.n6540 gnd.n6539 19.3944
R10140 gnd.n6539 gnd.n6538 19.3944
R10141 gnd.n6538 gnd.n873 19.3944
R10142 gnd.n6532 gnd.n873 19.3944
R10143 gnd.n6532 gnd.n6531 19.3944
R10144 gnd.n6531 gnd.n6530 19.3944
R10145 gnd.n6530 gnd.n881 19.3944
R10146 gnd.n6524 gnd.n881 19.3944
R10147 gnd.n6524 gnd.n6523 19.3944
R10148 gnd.n6523 gnd.n6522 19.3944
R10149 gnd.n6522 gnd.n889 19.3944
R10150 gnd.n6516 gnd.n889 19.3944
R10151 gnd.n6516 gnd.n6515 19.3944
R10152 gnd.n6515 gnd.n6514 19.3944
R10153 gnd.n6514 gnd.n897 19.3944
R10154 gnd.n6508 gnd.n897 19.3944
R10155 gnd.n6508 gnd.n6507 19.3944
R10156 gnd.n6507 gnd.n6506 19.3944
R10157 gnd.n6506 gnd.n905 19.3944
R10158 gnd.n6500 gnd.n905 19.3944
R10159 gnd.n6500 gnd.n6499 19.3944
R10160 gnd.n6499 gnd.n6498 19.3944
R10161 gnd.n6498 gnd.n913 19.3944
R10162 gnd.n6492 gnd.n913 19.3944
R10163 gnd.n6492 gnd.n6491 19.3944
R10164 gnd.n6491 gnd.n6490 19.3944
R10165 gnd.n6490 gnd.n921 19.3944
R10166 gnd.n6484 gnd.n921 19.3944
R10167 gnd.n6484 gnd.n6483 19.3944
R10168 gnd.n6483 gnd.n6482 19.3944
R10169 gnd.n6482 gnd.n929 19.3944
R10170 gnd.n6476 gnd.n929 19.3944
R10171 gnd.n6476 gnd.n6475 19.3944
R10172 gnd.n6475 gnd.n6474 19.3944
R10173 gnd.n2184 gnd.n2183 19.3944
R10174 gnd.n2183 gnd.n2182 19.3944
R10175 gnd.n2182 gnd.n2139 19.3944
R10176 gnd.n2178 gnd.n2139 19.3944
R10177 gnd.n2178 gnd.n2177 19.3944
R10178 gnd.n2177 gnd.n2176 19.3944
R10179 gnd.n2176 gnd.n2143 19.3944
R10180 gnd.n2172 gnd.n2143 19.3944
R10181 gnd.n2172 gnd.n2171 19.3944
R10182 gnd.n2171 gnd.n2170 19.3944
R10183 gnd.n2170 gnd.n2147 19.3944
R10184 gnd.n2166 gnd.n2147 19.3944
R10185 gnd.n2166 gnd.n2165 19.3944
R10186 gnd.n2165 gnd.n2164 19.3944
R10187 gnd.n2164 gnd.n2151 19.3944
R10188 gnd.n2160 gnd.n2151 19.3944
R10189 gnd.n2160 gnd.n2159 19.3944
R10190 gnd.n2159 gnd.n2158 19.3944
R10191 gnd.n2158 gnd.n2154 19.3944
R10192 gnd.n2154 gnd.n2040 19.3944
R10193 gnd.n2040 gnd.n2038 19.3944
R10194 gnd.n4887 gnd.n2038 19.3944
R10195 gnd.n4887 gnd.n2036 19.3944
R10196 gnd.n4891 gnd.n2036 19.3944
R10197 gnd.n4992 gnd.n4891 19.3944
R10198 gnd.n4993 gnd.n4992 19.3944
R10199 gnd.n4993 gnd.n2033 19.3944
R10200 gnd.n5024 gnd.n2033 19.3944
R10201 gnd.n5024 gnd.n2034 19.3944
R10202 gnd.n5020 gnd.n2034 19.3944
R10203 gnd.n5020 gnd.n5019 19.3944
R10204 gnd.n5019 gnd.n5018 19.3944
R10205 gnd.n5018 gnd.n4998 19.3944
R10206 gnd.n5014 gnd.n4998 19.3944
R10207 gnd.n5014 gnd.n5013 19.3944
R10208 gnd.n5013 gnd.n5012 19.3944
R10209 gnd.n5012 gnd.n5003 19.3944
R10210 gnd.n5008 gnd.n5003 19.3944
R10211 gnd.n5008 gnd.n5007 19.3944
R10212 gnd.n5007 gnd.n1971 19.3944
R10213 gnd.n5129 gnd.n1971 19.3944
R10214 gnd.n5130 gnd.n5129 19.3944
R10215 gnd.n5130 gnd.n1968 19.3944
R10216 gnd.n5160 gnd.n1968 19.3944
R10217 gnd.n5160 gnd.n1969 19.3944
R10218 gnd.n5156 gnd.n1969 19.3944
R10219 gnd.n5156 gnd.n5155 19.3944
R10220 gnd.n5155 gnd.n5154 19.3944
R10221 gnd.n5154 gnd.n5135 19.3944
R10222 gnd.n5150 gnd.n5135 19.3944
R10223 gnd.n5150 gnd.n5149 19.3944
R10224 gnd.n5149 gnd.n5148 19.3944
R10225 gnd.n5148 gnd.n5140 19.3944
R10226 gnd.n5144 gnd.n5140 19.3944
R10227 gnd.n5144 gnd.n5143 19.3944
R10228 gnd.n5143 gnd.n1878 19.3944
R10229 gnd.n5281 gnd.n1878 19.3944
R10230 gnd.n5281 gnd.n1875 19.3944
R10231 gnd.n5286 gnd.n1875 19.3944
R10232 gnd.n5286 gnd.n1876 19.3944
R10233 gnd.n1876 gnd.n1851 19.3944
R10234 gnd.n5330 gnd.n1851 19.3944
R10235 gnd.n5330 gnd.n1848 19.3944
R10236 gnd.n5350 gnd.n1848 19.3944
R10237 gnd.n5350 gnd.n1849 19.3944
R10238 gnd.n5346 gnd.n1849 19.3944
R10239 gnd.n5346 gnd.n5345 19.3944
R10240 gnd.n5345 gnd.n5344 19.3944
R10241 gnd.n5344 gnd.n5337 19.3944
R10242 gnd.n5340 gnd.n5337 19.3944
R10243 gnd.n5340 gnd.n5339 19.3944
R10244 gnd.n5339 gnd.n1799 19.3944
R10245 gnd.n5410 gnd.n1799 19.3944
R10246 gnd.n5410 gnd.n1796 19.3944
R10247 gnd.n5424 gnd.n1796 19.3944
R10248 gnd.n5424 gnd.n1797 19.3944
R10249 gnd.n5420 gnd.n1797 19.3944
R10250 gnd.n5420 gnd.n5419 19.3944
R10251 gnd.n5419 gnd.n5418 19.3944
R10252 gnd.n5418 gnd.n1721 19.3944
R10253 gnd.n5628 gnd.n1721 19.3944
R10254 gnd.n5628 gnd.n1719 19.3944
R10255 gnd.n5632 gnd.n1719 19.3944
R10256 gnd.n5632 gnd.n1709 19.3944
R10257 gnd.n5645 gnd.n1709 19.3944
R10258 gnd.n5645 gnd.n1707 19.3944
R10259 gnd.n5649 gnd.n1707 19.3944
R10260 gnd.n5649 gnd.n1697 19.3944
R10261 gnd.n5662 gnd.n1697 19.3944
R10262 gnd.n5662 gnd.n1695 19.3944
R10263 gnd.n5666 gnd.n1695 19.3944
R10264 gnd.n5666 gnd.n1684 19.3944
R10265 gnd.n5679 gnd.n1684 19.3944
R10266 gnd.n5679 gnd.n1682 19.3944
R10267 gnd.n5683 gnd.n1682 19.3944
R10268 gnd.n5683 gnd.n1673 19.3944
R10269 gnd.n5699 gnd.n1673 19.3944
R10270 gnd.n5699 gnd.n1671 19.3944
R10271 gnd.n5703 gnd.n1671 19.3944
R10272 gnd.n5703 gnd.n1299 19.3944
R10273 gnd.n6147 gnd.n1299 19.3944
R10274 gnd.n6144 gnd.n6143 19.3944
R10275 gnd.n6143 gnd.n6142 19.3944
R10276 gnd.n6142 gnd.n1304 19.3944
R10277 gnd.n6138 gnd.n1304 19.3944
R10278 gnd.n6138 gnd.n6137 19.3944
R10279 gnd.n6137 gnd.n6136 19.3944
R10280 gnd.n6136 gnd.n1309 19.3944
R10281 gnd.n6131 gnd.n1309 19.3944
R10282 gnd.n6131 gnd.n6130 19.3944
R10283 gnd.n6130 gnd.n1314 19.3944
R10284 gnd.n6123 gnd.n1314 19.3944
R10285 gnd.n6123 gnd.n6122 19.3944
R10286 gnd.n6122 gnd.n1323 19.3944
R10287 gnd.n6115 gnd.n1323 19.3944
R10288 gnd.n6115 gnd.n6114 19.3944
R10289 gnd.n6114 gnd.n1331 19.3944
R10290 gnd.n6107 gnd.n1331 19.3944
R10291 gnd.n6107 gnd.n6106 19.3944
R10292 gnd.n6106 gnd.n1339 19.3944
R10293 gnd.n6099 gnd.n1339 19.3944
R10294 gnd.n6099 gnd.n6098 19.3944
R10295 gnd.n6098 gnd.n1347 19.3944
R10296 gnd.n6091 gnd.n1347 19.3944
R10297 gnd.n6091 gnd.n6090 19.3944
R10298 gnd.n1659 gnd.n1638 19.3944
R10299 gnd.n5732 gnd.n1638 19.3944
R10300 gnd.n5732 gnd.n5731 19.3944
R10301 gnd.t88 gnd.n1157 19.1199
R10302 gnd.n5034 gnd.n2029 19.1199
R10303 gnd.n5407 gnd.n1802 19.1199
R10304 gnd.n3429 gnd.t29 18.8012
R10305 gnd.n3414 gnd.t356 18.8012
R10306 gnd.n4971 gnd.t64 18.8012
R10307 gnd.n5428 gnd.t27 18.8012
R10308 gnd.n3273 gnd.n3272 18.4825
R10309 gnd.n4529 gnd.n2436 18.4825
R10310 gnd.n4536 gnd.n4535 18.4825
R10311 gnd.n4565 gnd.n2422 18.4825
R10312 gnd.n4573 gnd.n958 18.4825
R10313 gnd.n6458 gnd.n967 18.4825
R10314 gnd.n4580 gnd.n2416 18.4825
R10315 gnd.n6452 gnd.n976 18.4825
R10316 gnd.n6446 gnd.n986 18.4825
R10317 gnd.n4624 gnd.n989 18.4825
R10318 gnd.n4595 gnd.n999 18.4825
R10319 gnd.n6434 gnd.n1006 18.4825
R10320 gnd.n4601 gnd.n4600 18.4825
R10321 gnd.n6428 gnd.n1016 18.4825
R10322 gnd.n6422 gnd.n1026 18.4825
R10323 gnd.n4672 gnd.n1029 18.4825
R10324 gnd.n4678 gnd.n1039 18.4825
R10325 gnd.n6410 gnd.n1046 18.4825
R10326 gnd.n4687 gnd.n1049 18.4825
R10327 gnd.n6404 gnd.n1057 18.4825
R10328 gnd.n4694 gnd.n2383 18.4825
R10329 gnd.n6398 gnd.n1065 18.4825
R10330 gnd.n5960 gnd.n1475 18.4825
R10331 gnd.n5777 gnd.n5776 18.4825
R10332 gnd.n5952 gnd.n1484 18.4825
R10333 gnd.n5737 gnd.n1497 18.4825
R10334 gnd.n5946 gnd.n1500 18.4825
R10335 gnd.n5744 gnd.n1510 18.4825
R10336 gnd.n5750 gnd.n1520 18.4825
R10337 gnd.n5934 gnd.n1523 18.4825
R10338 gnd.n5928 gnd.n1533 18.4825
R10339 gnd.n5822 gnd.n5821 18.4825
R10340 gnd.n5922 gnd.n1543 18.4825
R10341 gnd.n5830 gnd.n1550 18.4825
R10342 gnd.n5837 gnd.n1560 18.4825
R10343 gnd.n5910 gnd.n1563 18.4825
R10344 gnd.n5904 gnd.n1573 18.4825
R10345 gnd.n5876 gnd.n5875 18.4825
R10346 gnd.n5898 gnd.n1583 18.4825
R10347 gnd.n5859 gnd.n1590 18.4825
R10348 gnd.n5888 gnd.n5887 18.4825
R10349 gnd.n1597 gnd.n381 18.4825
R10350 gnd.n7283 gnd.n375 18.4825
R10351 gnd.n6029 gnd.n6028 18.4247
R10352 gnd.n6348 gnd.n6347 18.4247
R10353 gnd.n6087 gnd.n6086 18.2308
R10354 gnd.n4713 gnd.n4712 18.2308
R10355 gnd.n7394 gnd.n7393 18.2308
R10356 gnd.n4204 gnd.n4164 18.2308
R10357 gnd.t36 gnd.n2953 18.1639
R10358 gnd.n5093 gnd.n5092 17.8452
R10359 gnd.n5205 gnd.n5204 17.8452
R10360 gnd.n5240 gnd.n1907 17.8452
R10361 gnd.n5359 gnd.n1838 17.8452
R10362 gnd.n5442 gnd.t190 17.8452
R10363 gnd.n2981 gnd.t34 17.5266
R10364 gnd.n2536 gnd.t225 17.5266
R10365 gnd.n6416 gnd.t206 17.5266
R10366 gnd.n5940 gnd.t217 17.5266
R10367 gnd.n7555 gnd.t240 17.5266
R10368 gnd.n4973 gnd.t124 17.2079
R10369 gnd.n3380 gnd.t2 16.8893
R10370 gnd.n3657 gnd.n3656 16.8893
R10371 gnd.n2499 gnd.t238 16.8893
R10372 gnd.n6472 gnd.n6471 16.8893
R10373 gnd.n6440 gnd.t257 16.8893
R10374 gnd.t69 gnd.n1125 16.8893
R10375 gnd.n1747 gnd.t19 16.8893
R10376 gnd.n5916 gnd.t196 16.8893
R10377 gnd.n7611 gnd.n90 16.8893
R10378 gnd.n7579 gnd.t208 16.8893
R10379 gnd.n6011 gnd.n6008 16.6793
R10380 gnd.n7466 gnd.n7465 16.6793
R10381 gnd.n4284 gnd.n4281 16.6793
R10382 gnd.n2248 gnd.n2218 16.6793
R10383 gnd.n5045 gnd.t39 16.5706
R10384 gnd.n5066 gnd.n5065 16.5706
R10385 gnd.n1925 gnd.n1920 16.5706
R10386 gnd.n5232 gnd.n5230 16.5706
R10387 gnd.n1823 gnd.n1822 16.5706
R10388 gnd.t16 gnd.n5398 16.5706
R10389 gnd.n5547 gnd.t85 16.5706
R10390 gnd.n3208 gnd.t183 16.2519
R10391 gnd.n2908 gnd.t9 16.2519
R10392 gnd.n4497 gnd.t249 16.2519
R10393 gnd.n6464 gnd.t202 16.2519
R10394 gnd.n5892 gnd.t253 16.2519
R10395 gnd.n7603 gnd.t215 16.2519
R10396 gnd.n3896 gnd.n3894 15.6674
R10397 gnd.n3864 gnd.n3862 15.6674
R10398 gnd.n3832 gnd.n3830 15.6674
R10399 gnd.n3801 gnd.n3799 15.6674
R10400 gnd.n3769 gnd.n3767 15.6674
R10401 gnd.n3737 gnd.n3735 15.6674
R10402 gnd.n3705 gnd.n3703 15.6674
R10403 gnd.n3674 gnd.n3672 15.6674
R10404 gnd.n3199 gnd.t183 15.6146
R10405 gnd.t170 gnd.n2646 15.6146
R10406 gnd.t145 gnd.n2647 15.6146
R10407 gnd.n4501 gnd.t249 15.6146
R10408 gnd.n7345 gnd.t215 15.6146
R10409 gnd.n5968 gnd.n5963 15.3217
R10410 gnd.n7426 gnd.n315 15.3217
R10411 gnd.n4242 gnd.n2563 15.3217
R10412 gnd.n2303 gnd.n2196 15.3217
R10413 gnd.n5066 gnd.n2009 15.296
R10414 gnd.n2004 gnd.n1999 15.296
R10415 gnd.n1926 gnd.n1925 15.296
R10416 gnd.n5230 gnd.n1916 15.296
R10417 gnd.n5370 gnd.n1827 15.296
R10418 gnd.n1822 gnd.n1817 15.296
R10419 gnd.n5460 gnd.n5459 15.0827
R10420 gnd.n1169 gnd.n1164 15.0481
R10421 gnd.n5470 gnd.n5469 15.0481
R10422 gnd.n3567 gnd.t1 14.9773
R10423 gnd.n4441 gnd.t238 14.9773
R10424 gnd.n6472 gnd.n938 14.9773
R10425 gnd.n4882 gnd.t69 14.9773
R10426 gnd.t180 gnd.t59 14.9773
R10427 gnd.n5626 gnd.t19 14.9773
R10428 gnd.n368 gnd.n90 14.9773
R10429 gnd.t208 gnd.n136 14.9773
R10430 gnd.t136 gnd.n1776 14.6587
R10431 gnd.t161 gnd.n1747 14.6587
R10432 gnd.t54 gnd.n2689 14.34
R10433 gnd.n3645 gnd.t35 14.34
R10434 gnd.n4395 gnd.t225 14.34
R10435 gnd.t240 gnd.n174 14.34
R10436 gnd.n5046 gnd.n5045 14.0214
R10437 gnd.n5092 gnd.n1993 14.0214
R10438 gnd.n5205 gnd.n1931 14.0214
R10439 gnd.n1907 gnd.n1901 14.0214
R10440 gnd.n5352 gnd.n1838 14.0214
R10441 gnd.n5398 gnd.n1812 14.0214
R10442 gnd.n3355 gnd.t37 13.7027
R10443 gnd.n5162 gnd.t11 13.7027
R10444 gnd.n5279 gnd.t47 13.7027
R10445 gnd.n3065 gnd.n3064 13.5763
R10446 gnd.n4010 gnd.n2603 13.5763
R10447 gnd.n3273 gnd.n3011 13.384
R10448 gnd.n4516 gnd.n2436 13.384
R10449 gnd.n4529 gnd.n2439 13.384
R10450 gnd.n4536 gnd.n2432 13.384
R10451 gnd.n4535 gnd.n2422 13.384
R10452 gnd.n4565 gnd.n4564 13.384
R10453 gnd.n6464 gnd.n958 13.384
R10454 gnd.n4573 gnd.n967 13.384
R10455 gnd.n4580 gnd.n976 13.384
R10456 gnd.n6452 gnd.n979 13.384
R10457 gnd.n4588 gnd.n986 13.384
R10458 gnd.n6446 gnd.n989 13.384
R10459 gnd.n4625 gnd.n4624 13.384
R10460 gnd.n6440 gnd.n999 13.384
R10461 gnd.n4595 gnd.n1006 13.384
R10462 gnd.n4601 gnd.n1016 13.384
R10463 gnd.n6428 gnd.n1019 13.384
R10464 gnd.n4607 gnd.n1026 13.384
R10465 gnd.n6422 gnd.n1029 13.384
R10466 gnd.n4672 gnd.n4671 13.384
R10467 gnd.n6416 gnd.n1039 13.384
R10468 gnd.n4678 gnd.n1046 13.384
R10469 gnd.n6410 gnd.n1049 13.384
R10470 gnd.n4687 gnd.n1057 13.384
R10471 gnd.n4694 gnd.n1065 13.384
R10472 gnd.n6398 gnd.n1068 13.384
R10473 gnd.n5072 gnd.t8 13.384
R10474 gnd.n1830 gnd.t13 13.384
R10475 gnd.n5960 gnd.n1473 13.384
R10476 gnd.n5776 gnd.n1475 13.384
R10477 gnd.n5737 gnd.n1484 13.384
R10478 gnd.n5946 gnd.n1497 13.384
R10479 gnd.n5744 gnd.n1500 13.384
R10480 gnd.n5940 gnd.n1510 13.384
R10481 gnd.n5750 gnd.n5749 13.384
R10482 gnd.n5934 gnd.n1520 13.384
R10483 gnd.n5759 gnd.n1523 13.384
R10484 gnd.n5928 gnd.n1530 13.384
R10485 gnd.n5822 gnd.n1533 13.384
R10486 gnd.n5830 gnd.n1543 13.384
R10487 gnd.n5916 gnd.n1550 13.384
R10488 gnd.n5837 gnd.n1613 13.384
R10489 gnd.n5910 gnd.n1560 13.384
R10490 gnd.n5845 gnd.n1563 13.384
R10491 gnd.n5904 gnd.n1570 13.384
R10492 gnd.n5875 gnd.n1573 13.384
R10493 gnd.n5859 gnd.n1583 13.384
R10494 gnd.n5892 gnd.n1590 13.384
R10495 gnd.n5888 gnd.n1594 13.384
R10496 gnd.n5887 gnd.n1597 13.384
R10497 gnd.n7287 gnd.n381 13.384
R10498 gnd.n7283 gnd.n7281 13.384
R10499 gnd.n7296 gnd.n375 13.384
R10500 gnd.n1180 gnd.n1161 13.1884
R10501 gnd.n1175 gnd.n1174 13.1884
R10502 gnd.n1174 gnd.n1173 13.1884
R10503 gnd.n5463 gnd.n5458 13.1884
R10504 gnd.n5464 gnd.n5463 13.1884
R10505 gnd.n1176 gnd.n1163 13.146
R10506 gnd.n1172 gnd.n1163 13.146
R10507 gnd.n5462 gnd.n5461 13.146
R10508 gnd.n5462 gnd.n5457 13.146
R10509 gnd.n2439 gnd.t221 13.0654
R10510 gnd.n7281 gnd.t230 13.0654
R10511 gnd.n3897 gnd.n3893 12.8005
R10512 gnd.n3865 gnd.n3861 12.8005
R10513 gnd.n3833 gnd.n3829 12.8005
R10514 gnd.n3802 gnd.n3798 12.8005
R10515 gnd.n3770 gnd.n3766 12.8005
R10516 gnd.n3738 gnd.n3734 12.8005
R10517 gnd.n3706 gnd.n3702 12.8005
R10518 gnd.n3675 gnd.n3671 12.8005
R10519 gnd.n5026 gnd.n2029 12.7467
R10520 gnd.n5186 gnd.n5185 12.7467
R10521 gnd.n5267 gnd.n1890 12.7467
R10522 gnd.t255 gnd.n979 12.4281
R10523 gnd.t6 gnd.n2086 12.4281
R10524 gnd.n6343 gnd.n1157 12.4281
R10525 gnd.n5618 gnd.n5616 12.4281
R10526 gnd.n1687 gnd.t352 12.4281
R10527 gnd.t192 gnd.n1570 12.4281
R10528 gnd.n3064 gnd.n3059 12.4126
R10529 gnd.n4013 gnd.n4010 12.4126
R10530 gnd.n6340 gnd.n6277 12.1761
R10531 gnd.n5543 gnd.n5542 12.1761
R10532 gnd.n4657 gnd.n1073 12.1094
R10533 gnd.n6081 gnd.n1405 12.1094
R10534 gnd.n3901 gnd.n3900 12.0247
R10535 gnd.n3869 gnd.n3868 12.0247
R10536 gnd.n3837 gnd.n3836 12.0247
R10537 gnd.n3806 gnd.n3805 12.0247
R10538 gnd.n3774 gnd.n3773 12.0247
R10539 gnd.n3742 gnd.n3741 12.0247
R10540 gnd.n3710 gnd.n3709 12.0247
R10541 gnd.n3679 gnd.n3678 12.0247
R10542 gnd.t271 gnd.n1019 11.7908
R10543 gnd.t219 gnd.n1530 11.7908
R10544 gnd.n4961 gnd.t88 11.4721
R10545 gnd.n6273 gnd.n6272 11.4721
R10546 gnd.n5547 gnd.n1770 11.4721
R10547 gnd.n3904 gnd.n3891 11.249
R10548 gnd.n3872 gnd.n3859 11.249
R10549 gnd.n3840 gnd.n3827 11.249
R10550 gnd.n3809 gnd.n3796 11.249
R10551 gnd.n3777 gnd.n3764 11.249
R10552 gnd.n3745 gnd.n3732 11.249
R10553 gnd.n3713 gnd.n3700 11.249
R10554 gnd.n3682 gnd.n3669 11.249
R10555 gnd.n3343 gnd.t37 11.1535
R10556 gnd.n5108 gnd.t67 11.1535
R10557 gnd.n5310 gnd.t354 11.1535
R10558 gnd.t15 gnd.n5107 10.8348
R10559 gnd.t42 gnd.n5309 10.8348
R10560 gnd.n5971 gnd.n5968 10.6672
R10561 gnd.n7431 gnd.n315 10.6672
R10562 gnd.n4244 gnd.n4242 10.6672
R10563 gnd.n2298 gnd.n2196 10.6672
R10564 gnd.n5613 gnd.n5612 10.6151
R10565 gnd.n5612 gnd.n5609 10.6151
R10566 gnd.n5607 gnd.n5604 10.6151
R10567 gnd.n5604 gnd.n5603 10.6151
R10568 gnd.n5603 gnd.n5600 10.6151
R10569 gnd.n5600 gnd.n5599 10.6151
R10570 gnd.n5599 gnd.n5596 10.6151
R10571 gnd.n5596 gnd.n5595 10.6151
R10572 gnd.n5595 gnd.n5592 10.6151
R10573 gnd.n5592 gnd.n5591 10.6151
R10574 gnd.n5591 gnd.n5588 10.6151
R10575 gnd.n5588 gnd.n5587 10.6151
R10576 gnd.n5587 gnd.n5584 10.6151
R10577 gnd.n5584 gnd.n5583 10.6151
R10578 gnd.n5583 gnd.n5580 10.6151
R10579 gnd.n5580 gnd.n5579 10.6151
R10580 gnd.n5579 gnd.n5576 10.6151
R10581 gnd.n5576 gnd.n5575 10.6151
R10582 gnd.n5575 gnd.n5572 10.6151
R10583 gnd.n5572 gnd.n5571 10.6151
R10584 gnd.n5571 gnd.n5568 10.6151
R10585 gnd.n5568 gnd.n5567 10.6151
R10586 gnd.n5567 gnd.n5564 10.6151
R10587 gnd.n5564 gnd.n5563 10.6151
R10588 gnd.n5563 gnd.n5560 10.6151
R10589 gnd.n5560 gnd.n5559 10.6151
R10590 gnd.n5559 gnd.n5556 10.6151
R10591 gnd.n5556 gnd.n5555 10.6151
R10592 gnd.n5555 gnd.n5552 10.6151
R10593 gnd.n5552 gnd.n5551 10.6151
R10594 gnd.n4964 gnd.n4963 10.6151
R10595 gnd.n4965 gnd.n4964 10.6151
R10596 gnd.n4988 gnd.n4965 10.6151
R10597 gnd.n4988 gnd.n4987 10.6151
R10598 gnd.n4987 gnd.n4986 10.6151
R10599 gnd.n4986 gnd.n4966 10.6151
R10600 gnd.n4967 gnd.n4966 10.6151
R10601 gnd.n4967 gnd.n2027 10.6151
R10602 gnd.n5037 gnd.n2027 10.6151
R10603 gnd.n5038 gnd.n5037 10.6151
R10604 gnd.n5043 gnd.n5038 10.6151
R10605 gnd.n5043 gnd.n5042 10.6151
R10606 gnd.n5042 gnd.n5041 10.6151
R10607 gnd.n5041 gnd.n5039 10.6151
R10608 gnd.n5039 gnd.n2002 10.6151
R10609 gnd.n5074 gnd.n2002 10.6151
R10610 gnd.n5075 gnd.n5074 10.6151
R10611 gnd.n5081 gnd.n5075 10.6151
R10612 gnd.n5081 gnd.n5080 10.6151
R10613 gnd.n5080 gnd.n5079 10.6151
R10614 gnd.n5079 gnd.n5078 10.6151
R10615 gnd.n5078 gnd.n1981 10.6151
R10616 gnd.n5110 gnd.n1981 10.6151
R10617 gnd.n5111 gnd.n5110 10.6151
R10618 gnd.n5117 gnd.n5111 10.6151
R10619 gnd.n5117 gnd.n5116 10.6151
R10620 gnd.n5116 gnd.n5115 10.6151
R10621 gnd.n5115 gnd.n5113 10.6151
R10622 gnd.n5113 gnd.n5112 10.6151
R10623 gnd.n5112 gnd.n1950 10.6151
R10624 gnd.n5177 gnd.n1950 10.6151
R10625 gnd.n5178 gnd.n5177 10.6151
R10626 gnd.n5183 gnd.n5178 10.6151
R10627 gnd.n5183 gnd.n5182 10.6151
R10628 gnd.n5182 gnd.n5181 10.6151
R10629 gnd.n5181 gnd.n5179 10.6151
R10630 gnd.n5179 gnd.n1923 10.6151
R10631 gnd.n5213 gnd.n1923 10.6151
R10632 gnd.n5214 gnd.n5213 10.6151
R10633 gnd.n5222 gnd.n5214 10.6151
R10634 gnd.n5222 gnd.n5221 10.6151
R10635 gnd.n5221 gnd.n5220 10.6151
R10636 gnd.n5220 gnd.n5219 10.6151
R10637 gnd.n5219 gnd.n5216 10.6151
R10638 gnd.n5216 gnd.n5215 10.6151
R10639 gnd.n5215 gnd.n1899 10.6151
R10640 gnd.n5250 gnd.n1899 10.6151
R10641 gnd.n5251 gnd.n5250 10.6151
R10642 gnd.n5254 gnd.n5251 10.6151
R10643 gnd.n5255 gnd.n5254 10.6151
R10644 gnd.n5257 gnd.n5255 10.6151
R10645 gnd.n5257 gnd.n5256 10.6151
R10646 gnd.n5256 gnd.n1870 10.6151
R10647 gnd.n5292 gnd.n1870 10.6151
R10648 gnd.n5293 gnd.n5292 10.6151
R10649 gnd.n5296 gnd.n5293 10.6151
R10650 gnd.n5297 gnd.n5296 10.6151
R10651 gnd.n5306 gnd.n5297 10.6151
R10652 gnd.n5306 gnd.n5305 10.6151
R10653 gnd.n5305 gnd.n5304 10.6151
R10654 gnd.n5304 gnd.n5303 10.6151
R10655 gnd.n5303 gnd.n5301 10.6151
R10656 gnd.n5301 gnd.n5300 10.6151
R10657 gnd.n5300 gnd.n5298 10.6151
R10658 gnd.n5298 gnd.n1820 10.6151
R10659 gnd.n5378 gnd.n1820 10.6151
R10660 gnd.n5379 gnd.n5378 10.6151
R10661 gnd.n5387 gnd.n5379 10.6151
R10662 gnd.n5387 gnd.n5386 10.6151
R10663 gnd.n5386 gnd.n5385 10.6151
R10664 gnd.n5385 gnd.n5384 10.6151
R10665 gnd.n5384 gnd.n5380 10.6151
R10666 gnd.n5380 gnd.n1793 10.6151
R10667 gnd.n5433 gnd.n1793 10.6151
R10668 gnd.n5433 gnd.n5432 10.6151
R10669 gnd.n5432 gnd.n5431 10.6151
R10670 gnd.n5431 gnd.n5430 10.6151
R10671 gnd.n5430 gnd.n1795 10.6151
R10672 gnd.n1795 gnd.n1794 10.6151
R10673 gnd.n1794 gnd.n1769 10.6151
R10674 gnd.n1769 gnd.n1767 10.6151
R10675 gnd.n4898 gnd.n1121 10.6151
R10676 gnd.n4901 gnd.n4898 10.6151
R10677 gnd.n4906 gnd.n4903 10.6151
R10678 gnd.n4907 gnd.n4906 10.6151
R10679 gnd.n4910 gnd.n4907 10.6151
R10680 gnd.n4911 gnd.n4910 10.6151
R10681 gnd.n4914 gnd.n4911 10.6151
R10682 gnd.n4915 gnd.n4914 10.6151
R10683 gnd.n4918 gnd.n4915 10.6151
R10684 gnd.n4919 gnd.n4918 10.6151
R10685 gnd.n4922 gnd.n4919 10.6151
R10686 gnd.n4923 gnd.n4922 10.6151
R10687 gnd.n4926 gnd.n4923 10.6151
R10688 gnd.n4927 gnd.n4926 10.6151
R10689 gnd.n4930 gnd.n4927 10.6151
R10690 gnd.n4931 gnd.n4930 10.6151
R10691 gnd.n4934 gnd.n4931 10.6151
R10692 gnd.n4935 gnd.n4934 10.6151
R10693 gnd.n4938 gnd.n4935 10.6151
R10694 gnd.n4939 gnd.n4938 10.6151
R10695 gnd.n4942 gnd.n4939 10.6151
R10696 gnd.n4943 gnd.n4942 10.6151
R10697 gnd.n4946 gnd.n4943 10.6151
R10698 gnd.n4947 gnd.n4946 10.6151
R10699 gnd.n4950 gnd.n4947 10.6151
R10700 gnd.n4951 gnd.n4950 10.6151
R10701 gnd.n4954 gnd.n4951 10.6151
R10702 gnd.n4955 gnd.n4954 10.6151
R10703 gnd.n4958 gnd.n4955 10.6151
R10704 gnd.n4959 gnd.n4958 10.6151
R10705 gnd.n6340 gnd.n6339 10.6151
R10706 gnd.n6339 gnd.n6338 10.6151
R10707 gnd.n6338 gnd.n6337 10.6151
R10708 gnd.n6337 gnd.n6335 10.6151
R10709 gnd.n6335 gnd.n6332 10.6151
R10710 gnd.n6332 gnd.n6331 10.6151
R10711 gnd.n6331 gnd.n6328 10.6151
R10712 gnd.n6328 gnd.n6327 10.6151
R10713 gnd.n6327 gnd.n6324 10.6151
R10714 gnd.n6324 gnd.n6323 10.6151
R10715 gnd.n6323 gnd.n6320 10.6151
R10716 gnd.n6320 gnd.n6319 10.6151
R10717 gnd.n6319 gnd.n6316 10.6151
R10718 gnd.n6316 gnd.n6315 10.6151
R10719 gnd.n6315 gnd.n6312 10.6151
R10720 gnd.n6312 gnd.n6311 10.6151
R10721 gnd.n6311 gnd.n6308 10.6151
R10722 gnd.n6308 gnd.n6307 10.6151
R10723 gnd.n6307 gnd.n6304 10.6151
R10724 gnd.n6304 gnd.n6303 10.6151
R10725 gnd.n6303 gnd.n6300 10.6151
R10726 gnd.n6300 gnd.n6299 10.6151
R10727 gnd.n6299 gnd.n6296 10.6151
R10728 gnd.n6296 gnd.n6295 10.6151
R10729 gnd.n6295 gnd.n6292 10.6151
R10730 gnd.n6292 gnd.n6291 10.6151
R10731 gnd.n6291 gnd.n6288 10.6151
R10732 gnd.n6288 gnd.n6287 10.6151
R10733 gnd.n6284 gnd.n6283 10.6151
R10734 gnd.n6283 gnd.n1122 10.6151
R10735 gnd.n5542 gnd.n5540 10.6151
R10736 gnd.n5540 gnd.n5537 10.6151
R10737 gnd.n5537 gnd.n5536 10.6151
R10738 gnd.n5536 gnd.n5533 10.6151
R10739 gnd.n5533 gnd.n5532 10.6151
R10740 gnd.n5532 gnd.n5529 10.6151
R10741 gnd.n5529 gnd.n5528 10.6151
R10742 gnd.n5528 gnd.n5525 10.6151
R10743 gnd.n5525 gnd.n5524 10.6151
R10744 gnd.n5524 gnd.n5521 10.6151
R10745 gnd.n5521 gnd.n5520 10.6151
R10746 gnd.n5520 gnd.n5517 10.6151
R10747 gnd.n5517 gnd.n5516 10.6151
R10748 gnd.n5516 gnd.n5513 10.6151
R10749 gnd.n5513 gnd.n5512 10.6151
R10750 gnd.n5512 gnd.n5509 10.6151
R10751 gnd.n5509 gnd.n5508 10.6151
R10752 gnd.n5508 gnd.n5505 10.6151
R10753 gnd.n5505 gnd.n5504 10.6151
R10754 gnd.n5504 gnd.n5501 10.6151
R10755 gnd.n5501 gnd.n5500 10.6151
R10756 gnd.n5500 gnd.n5497 10.6151
R10757 gnd.n5497 gnd.n5496 10.6151
R10758 gnd.n5496 gnd.n5493 10.6151
R10759 gnd.n5493 gnd.n5492 10.6151
R10760 gnd.n5492 gnd.n5489 10.6151
R10761 gnd.n5489 gnd.n5488 10.6151
R10762 gnd.n5488 gnd.n5485 10.6151
R10763 gnd.n5483 gnd.n5480 10.6151
R10764 gnd.n5480 gnd.n5479 10.6151
R10765 gnd.n6276 gnd.n6275 10.6151
R10766 gnd.n6275 gnd.n1181 10.6151
R10767 gnd.n4975 gnd.n1181 10.6151
R10768 gnd.n4976 gnd.n4975 10.6151
R10769 gnd.n4982 gnd.n4976 10.6151
R10770 gnd.n4982 gnd.n4981 10.6151
R10771 gnd.n4981 gnd.n4980 10.6151
R10772 gnd.n4980 gnd.n4977 10.6151
R10773 gnd.n4977 gnd.n2023 10.6151
R10774 gnd.n5049 gnd.n2023 10.6151
R10775 gnd.n5050 gnd.n5049 10.6151
R10776 gnd.n5051 gnd.n5050 10.6151
R10777 gnd.n5051 gnd.n2007 10.6151
R10778 gnd.n5068 gnd.n2007 10.6151
R10779 gnd.n5069 gnd.n5068 10.6151
R10780 gnd.n5070 gnd.n5069 10.6151
R10781 gnd.n5070 gnd.n1996 10.6151
R10782 gnd.n5085 gnd.n1996 10.6151
R10783 gnd.n5086 gnd.n5085 10.6151
R10784 gnd.n5090 gnd.n5086 10.6151
R10785 gnd.n5090 gnd.n5089 10.6151
R10786 gnd.n5089 gnd.n5088 10.6151
R10787 gnd.n5088 gnd.n1976 10.6151
R10788 gnd.n5122 gnd.n1976 10.6151
R10789 gnd.n5123 gnd.n5122 10.6151
R10790 gnd.n5124 gnd.n5123 10.6151
R10791 gnd.n5124 gnd.n1953 10.6151
R10792 gnd.n5170 gnd.n1953 10.6151
R10793 gnd.n5171 gnd.n5170 10.6151
R10794 gnd.n5172 gnd.n5171 10.6151
R10795 gnd.n5172 gnd.n1945 10.6151
R10796 gnd.n5189 gnd.n1945 10.6151
R10797 gnd.n5190 gnd.n5189 10.6151
R10798 gnd.n5191 gnd.n5190 10.6151
R10799 gnd.n5191 gnd.n1928 10.6151
R10800 gnd.n5207 gnd.n1928 10.6151
R10801 gnd.n5208 gnd.n5207 10.6151
R10802 gnd.n5209 gnd.n5208 10.6151
R10803 gnd.n5209 gnd.n1918 10.6151
R10804 gnd.n5226 gnd.n1918 10.6151
R10805 gnd.n5227 gnd.n5226 10.6151
R10806 gnd.n5228 gnd.n5227 10.6151
R10807 gnd.n5228 gnd.n1903 10.6151
R10808 gnd.n5243 gnd.n1903 10.6151
R10809 gnd.n5244 gnd.n5243 10.6151
R10810 gnd.n5245 gnd.n5244 10.6151
R10811 gnd.n5245 gnd.n1893 10.6151
R10812 gnd.n5265 gnd.n1893 10.6151
R10813 gnd.n5265 gnd.n5264 10.6151
R10814 gnd.n5264 gnd.n5263 10.6151
R10815 gnd.n5263 gnd.n1894 10.6151
R10816 gnd.n1896 gnd.n1894 10.6151
R10817 gnd.n1896 gnd.n1895 10.6151
R10818 gnd.n1895 gnd.n1866 10.6151
R10819 gnd.n5315 gnd.n1866 10.6151
R10820 gnd.n5315 gnd.n5314 10.6151
R10821 gnd.n5314 gnd.n5313 10.6151
R10822 gnd.n5313 gnd.n1867 10.6151
R10823 gnd.n1867 gnd.n1843 10.6151
R10824 gnd.n5355 gnd.n1843 10.6151
R10825 gnd.n5356 gnd.n5355 10.6151
R10826 gnd.n5357 gnd.n5356 10.6151
R10827 gnd.n5357 gnd.n1825 10.6151
R10828 gnd.n5372 gnd.n1825 10.6151
R10829 gnd.n5373 gnd.n5372 10.6151
R10830 gnd.n5374 gnd.n5373 10.6151
R10831 gnd.n5374 gnd.n1815 10.6151
R10832 gnd.n5391 gnd.n1815 10.6151
R10833 gnd.n5392 gnd.n5391 10.6151
R10834 gnd.n5396 gnd.n5392 10.6151
R10835 gnd.n5396 gnd.n5395 10.6151
R10836 gnd.n5395 gnd.n5394 10.6151
R10837 gnd.n5394 gnd.n1788 10.6151
R10838 gnd.n5437 gnd.n1788 10.6151
R10839 gnd.n5438 gnd.n5437 10.6151
R10840 gnd.n5439 gnd.n5438 10.6151
R10841 gnd.n5439 gnd.n1773 10.6151
R10842 gnd.n5454 gnd.n1773 10.6151
R10843 gnd.n5455 gnd.n5454 10.6151
R10844 gnd.n5545 gnd.n5455 10.6151
R10845 gnd.n5545 gnd.n5544 10.6151
R10846 gnd.n3262 gnd.t45 10.5161
R10847 gnd.n2691 gnd.t54 10.5161
R10848 gnd.n3628 gnd.t35 10.5161
R10849 gnd.n2005 gnd.t17 10.5161
R10850 gnd.t366 gnd.n5369 10.5161
R10851 gnd.n3905 gnd.n3889 10.4732
R10852 gnd.n3873 gnd.n3857 10.4732
R10853 gnd.n3841 gnd.n3825 10.4732
R10854 gnd.n3810 gnd.n3794 10.4732
R10855 gnd.n3778 gnd.n3762 10.4732
R10856 gnd.n3746 gnd.n3730 10.4732
R10857 gnd.n3714 gnd.n3698 10.4732
R10858 gnd.n3683 gnd.n3667 10.4732
R10859 gnd.n6266 gnd.t73 10.1975
R10860 gnd.n5127 gnd.n1955 10.1975
R10861 gnd.n1966 gnd.n1957 10.1975
R10862 gnd.n5185 gnd.t21 10.1975
R10863 gnd.t22 gnd.n5267 10.1975
R10864 gnd.n5259 gnd.n1872 10.1975
R10865 gnd.n5318 gnd.n1860 10.1975
R10866 gnd.n5427 gnd.t102 10.1975
R10867 gnd.n5428 gnd.n5427 10.1975
R10868 gnd.n1776 gnd.n1770 10.1975
R10869 gnd.t1 gnd.n2708 9.87883
R10870 gnd.n3909 gnd.n3908 9.69747
R10871 gnd.n3877 gnd.n3876 9.69747
R10872 gnd.n3845 gnd.n3844 9.69747
R10873 gnd.n3814 gnd.n3813 9.69747
R10874 gnd.n3782 gnd.n3781 9.69747
R10875 gnd.n3750 gnd.n3749 9.69747
R10876 gnd.n3718 gnd.n3717 9.69747
R10877 gnd.n3687 gnd.n3686 9.69747
R10878 gnd.n1802 gnd.t121 9.56018
R10879 gnd.n3915 gnd.n3914 9.45567
R10880 gnd.n3883 gnd.n3882 9.45567
R10881 gnd.n3851 gnd.n3850 9.45567
R10882 gnd.n3820 gnd.n3819 9.45567
R10883 gnd.n3788 gnd.n3787 9.45567
R10884 gnd.n3756 gnd.n3755 9.45567
R10885 gnd.n3724 gnd.n3723 9.45567
R10886 gnd.n3693 gnd.n3692 9.45567
R10887 gnd.n6008 gnd.n6007 9.30959
R10888 gnd.n7465 gnd.n279 9.30959
R10889 gnd.n4281 gnd.n4280 9.30959
R10890 gnd.n2254 gnd.n2218 9.30959
R10891 gnd.n3914 gnd.n3913 9.3005
R10892 gnd.n3887 gnd.n3886 9.3005
R10893 gnd.n3908 gnd.n3907 9.3005
R10894 gnd.n3906 gnd.n3905 9.3005
R10895 gnd.n3891 gnd.n3890 9.3005
R10896 gnd.n3900 gnd.n3899 9.3005
R10897 gnd.n3898 gnd.n3897 9.3005
R10898 gnd.n3882 gnd.n3881 9.3005
R10899 gnd.n3855 gnd.n3854 9.3005
R10900 gnd.n3876 gnd.n3875 9.3005
R10901 gnd.n3874 gnd.n3873 9.3005
R10902 gnd.n3859 gnd.n3858 9.3005
R10903 gnd.n3868 gnd.n3867 9.3005
R10904 gnd.n3866 gnd.n3865 9.3005
R10905 gnd.n3850 gnd.n3849 9.3005
R10906 gnd.n3823 gnd.n3822 9.3005
R10907 gnd.n3844 gnd.n3843 9.3005
R10908 gnd.n3842 gnd.n3841 9.3005
R10909 gnd.n3827 gnd.n3826 9.3005
R10910 gnd.n3836 gnd.n3835 9.3005
R10911 gnd.n3834 gnd.n3833 9.3005
R10912 gnd.n3819 gnd.n3818 9.3005
R10913 gnd.n3792 gnd.n3791 9.3005
R10914 gnd.n3813 gnd.n3812 9.3005
R10915 gnd.n3811 gnd.n3810 9.3005
R10916 gnd.n3796 gnd.n3795 9.3005
R10917 gnd.n3805 gnd.n3804 9.3005
R10918 gnd.n3803 gnd.n3802 9.3005
R10919 gnd.n3787 gnd.n3786 9.3005
R10920 gnd.n3760 gnd.n3759 9.3005
R10921 gnd.n3781 gnd.n3780 9.3005
R10922 gnd.n3779 gnd.n3778 9.3005
R10923 gnd.n3764 gnd.n3763 9.3005
R10924 gnd.n3773 gnd.n3772 9.3005
R10925 gnd.n3771 gnd.n3770 9.3005
R10926 gnd.n3755 gnd.n3754 9.3005
R10927 gnd.n3728 gnd.n3727 9.3005
R10928 gnd.n3749 gnd.n3748 9.3005
R10929 gnd.n3747 gnd.n3746 9.3005
R10930 gnd.n3732 gnd.n3731 9.3005
R10931 gnd.n3741 gnd.n3740 9.3005
R10932 gnd.n3739 gnd.n3738 9.3005
R10933 gnd.n3723 gnd.n3722 9.3005
R10934 gnd.n3696 gnd.n3695 9.3005
R10935 gnd.n3717 gnd.n3716 9.3005
R10936 gnd.n3715 gnd.n3714 9.3005
R10937 gnd.n3700 gnd.n3699 9.3005
R10938 gnd.n3709 gnd.n3708 9.3005
R10939 gnd.n3707 gnd.n3706 9.3005
R10940 gnd.n3692 gnd.n3691 9.3005
R10941 gnd.n3665 gnd.n3664 9.3005
R10942 gnd.n3686 gnd.n3685 9.3005
R10943 gnd.n3684 gnd.n3683 9.3005
R10944 gnd.n3669 gnd.n3668 9.3005
R10945 gnd.n3678 gnd.n3677 9.3005
R10946 gnd.n3676 gnd.n3675 9.3005
R10947 gnd.n4040 gnd.n4039 9.3005
R10948 gnd.n4038 gnd.n2591 9.3005
R10949 gnd.n4037 gnd.n4036 9.3005
R10950 gnd.n4033 gnd.n2592 9.3005
R10951 gnd.n4030 gnd.n2593 9.3005
R10952 gnd.n4029 gnd.n2594 9.3005
R10953 gnd.n4026 gnd.n2595 9.3005
R10954 gnd.n4025 gnd.n2596 9.3005
R10955 gnd.n4022 gnd.n2597 9.3005
R10956 gnd.n4021 gnd.n2598 9.3005
R10957 gnd.n4018 gnd.n2599 9.3005
R10958 gnd.n4017 gnd.n2600 9.3005
R10959 gnd.n4014 gnd.n2601 9.3005
R10960 gnd.n4013 gnd.n2602 9.3005
R10961 gnd.n4010 gnd.n4009 9.3005
R10962 gnd.n4008 gnd.n2603 9.3005
R10963 gnd.n4041 gnd.n2590 9.3005
R10964 gnd.n3281 gnd.n3280 9.3005
R10965 gnd.n2985 gnd.n2984 9.3005
R10966 gnd.n3308 gnd.n3307 9.3005
R10967 gnd.n3309 gnd.n2983 9.3005
R10968 gnd.n3313 gnd.n3310 9.3005
R10969 gnd.n3312 gnd.n3311 9.3005
R10970 gnd.n2957 gnd.n2956 9.3005
R10971 gnd.n3338 gnd.n3337 9.3005
R10972 gnd.n3339 gnd.n2955 9.3005
R10973 gnd.n3341 gnd.n3340 9.3005
R10974 gnd.n2935 gnd.n2934 9.3005
R10975 gnd.n3369 gnd.n3368 9.3005
R10976 gnd.n3370 gnd.n2933 9.3005
R10977 gnd.n3378 gnd.n3371 9.3005
R10978 gnd.n3377 gnd.n3372 9.3005
R10979 gnd.n3376 gnd.n3374 9.3005
R10980 gnd.n3373 gnd.n2882 9.3005
R10981 gnd.n3426 gnd.n2883 9.3005
R10982 gnd.n3425 gnd.n2884 9.3005
R10983 gnd.n3424 gnd.n2885 9.3005
R10984 gnd.n2904 gnd.n2886 9.3005
R10985 gnd.n2906 gnd.n2905 9.3005
R10986 gnd.n2788 gnd.n2787 9.3005
R10987 gnd.n3464 gnd.n3463 9.3005
R10988 gnd.n3465 gnd.n2786 9.3005
R10989 gnd.n3469 gnd.n3466 9.3005
R10990 gnd.n3468 gnd.n3467 9.3005
R10991 gnd.n2761 gnd.n2760 9.3005
R10992 gnd.n3504 gnd.n3503 9.3005
R10993 gnd.n3505 gnd.n2759 9.3005
R10994 gnd.n3509 gnd.n3506 9.3005
R10995 gnd.n3508 gnd.n3507 9.3005
R10996 gnd.n2734 gnd.n2733 9.3005
R10997 gnd.n3549 gnd.n3548 9.3005
R10998 gnd.n3550 gnd.n2732 9.3005
R10999 gnd.n3554 gnd.n3551 9.3005
R11000 gnd.n3553 gnd.n3552 9.3005
R11001 gnd.n2706 gnd.n2705 9.3005
R11002 gnd.n3589 gnd.n3588 9.3005
R11003 gnd.n3590 gnd.n2704 9.3005
R11004 gnd.n3594 gnd.n3591 9.3005
R11005 gnd.n3593 gnd.n3592 9.3005
R11006 gnd.n2679 gnd.n2678 9.3005
R11007 gnd.n3638 gnd.n3637 9.3005
R11008 gnd.n3639 gnd.n2677 9.3005
R11009 gnd.n3643 gnd.n3640 9.3005
R11010 gnd.n3642 gnd.n3641 9.3005
R11011 gnd.n2652 gnd.n2651 9.3005
R11012 gnd.n3933 gnd.n3932 9.3005
R11013 gnd.n3934 gnd.n2650 9.3005
R11014 gnd.n3940 gnd.n3935 9.3005
R11015 gnd.n3939 gnd.n3936 9.3005
R11016 gnd.n3938 gnd.n3937 9.3005
R11017 gnd.n3282 gnd.n3279 9.3005
R11018 gnd.n3064 gnd.n3023 9.3005
R11019 gnd.n3059 gnd.n3058 9.3005
R11020 gnd.n3057 gnd.n3024 9.3005
R11021 gnd.n3056 gnd.n3055 9.3005
R11022 gnd.n3052 gnd.n3025 9.3005
R11023 gnd.n3049 gnd.n3048 9.3005
R11024 gnd.n3047 gnd.n3026 9.3005
R11025 gnd.n3046 gnd.n3045 9.3005
R11026 gnd.n3042 gnd.n3027 9.3005
R11027 gnd.n3039 gnd.n3038 9.3005
R11028 gnd.n3037 gnd.n3028 9.3005
R11029 gnd.n3036 gnd.n3035 9.3005
R11030 gnd.n3032 gnd.n3030 9.3005
R11031 gnd.n3029 gnd.n3009 9.3005
R11032 gnd.n3276 gnd.n3008 9.3005
R11033 gnd.n3278 gnd.n3277 9.3005
R11034 gnd.n3066 gnd.n3065 9.3005
R11035 gnd.n3289 gnd.n2995 9.3005
R11036 gnd.n3296 gnd.n2996 9.3005
R11037 gnd.n3298 gnd.n3297 9.3005
R11038 gnd.n3299 gnd.n2976 9.3005
R11039 gnd.n3318 gnd.n3317 9.3005
R11040 gnd.n3320 gnd.n2968 9.3005
R11041 gnd.n3327 gnd.n2970 9.3005
R11042 gnd.n3328 gnd.n2965 9.3005
R11043 gnd.n3330 gnd.n3329 9.3005
R11044 gnd.n2966 gnd.n2951 9.3005
R11045 gnd.n3346 gnd.n2949 9.3005
R11046 gnd.n3350 gnd.n3349 9.3005
R11047 gnd.n3348 gnd.n2925 9.3005
R11048 gnd.n3385 gnd.n2924 9.3005
R11049 gnd.n3388 gnd.n3387 9.3005
R11050 gnd.n2921 gnd.n2920 9.3005
R11051 gnd.n3394 gnd.n2922 9.3005
R11052 gnd.n3396 gnd.n3395 9.3005
R11053 gnd.n3398 gnd.n2919 9.3005
R11054 gnd.n3401 gnd.n3400 9.3005
R11055 gnd.n3404 gnd.n3402 9.3005
R11056 gnd.n3406 gnd.n3405 9.3005
R11057 gnd.n3412 gnd.n3407 9.3005
R11058 gnd.n3411 gnd.n3410 9.3005
R11059 gnd.n2779 gnd.n2778 9.3005
R11060 gnd.n3478 gnd.n3477 9.3005
R11061 gnd.n3479 gnd.n2772 9.3005
R11062 gnd.n3487 gnd.n2771 9.3005
R11063 gnd.n3490 gnd.n3489 9.3005
R11064 gnd.n3492 gnd.n3491 9.3005
R11065 gnd.n3495 gnd.n2754 9.3005
R11066 gnd.n3493 gnd.n2752 9.3005
R11067 gnd.n3515 gnd.n2750 9.3005
R11068 gnd.n3517 gnd.n3516 9.3005
R11069 gnd.n2724 gnd.n2723 9.3005
R11070 gnd.n3563 gnd.n3562 9.3005
R11071 gnd.n3564 gnd.n2717 9.3005
R11072 gnd.n3572 gnd.n2716 9.3005
R11073 gnd.n3575 gnd.n3574 9.3005
R11074 gnd.n3577 gnd.n3576 9.3005
R11075 gnd.n3580 gnd.n2699 9.3005
R11076 gnd.n3578 gnd.n2697 9.3005
R11077 gnd.n3600 gnd.n2695 9.3005
R11078 gnd.n3602 gnd.n3601 9.3005
R11079 gnd.n2670 gnd.n2669 9.3005
R11080 gnd.n3652 gnd.n3651 9.3005
R11081 gnd.n3653 gnd.n2663 9.3005
R11082 gnd.n3662 gnd.n2662 9.3005
R11083 gnd.n3921 gnd.n3920 9.3005
R11084 gnd.n3923 gnd.n3922 9.3005
R11085 gnd.n3924 gnd.n2643 9.3005
R11086 gnd.n3948 gnd.n3947 9.3005
R11087 gnd.n2644 gnd.n2606 9.3005
R11088 gnd.n3287 gnd.n3286 9.3005
R11089 gnd.n4004 gnd.n2607 9.3005
R11090 gnd.n4003 gnd.n2609 9.3005
R11091 gnd.n4000 gnd.n2610 9.3005
R11092 gnd.n3999 gnd.n2611 9.3005
R11093 gnd.n3996 gnd.n2612 9.3005
R11094 gnd.n3995 gnd.n2613 9.3005
R11095 gnd.n3992 gnd.n2614 9.3005
R11096 gnd.n3991 gnd.n2615 9.3005
R11097 gnd.n3988 gnd.n2616 9.3005
R11098 gnd.n3987 gnd.n2617 9.3005
R11099 gnd.n3984 gnd.n2618 9.3005
R11100 gnd.n3983 gnd.n2619 9.3005
R11101 gnd.n3980 gnd.n2620 9.3005
R11102 gnd.n3979 gnd.n2621 9.3005
R11103 gnd.n3976 gnd.n2622 9.3005
R11104 gnd.n3975 gnd.n2623 9.3005
R11105 gnd.n3972 gnd.n2624 9.3005
R11106 gnd.n3971 gnd.n2625 9.3005
R11107 gnd.n3968 gnd.n2626 9.3005
R11108 gnd.n3967 gnd.n2627 9.3005
R11109 gnd.n3964 gnd.n2628 9.3005
R11110 gnd.n3963 gnd.n2629 9.3005
R11111 gnd.n3960 gnd.n2633 9.3005
R11112 gnd.n3959 gnd.n2634 9.3005
R11113 gnd.n3956 gnd.n2635 9.3005
R11114 gnd.n3955 gnd.n2636 9.3005
R11115 gnd.n4006 gnd.n4005 9.3005
R11116 gnd.n3456 gnd.n3440 9.3005
R11117 gnd.n3455 gnd.n3441 9.3005
R11118 gnd.n3454 gnd.n3442 9.3005
R11119 gnd.n3452 gnd.n3443 9.3005
R11120 gnd.n3451 gnd.n3444 9.3005
R11121 gnd.n3449 gnd.n3445 9.3005
R11122 gnd.n3448 gnd.n3446 9.3005
R11123 gnd.n2742 gnd.n2741 9.3005
R11124 gnd.n3525 gnd.n3524 9.3005
R11125 gnd.n3526 gnd.n2740 9.3005
R11126 gnd.n3543 gnd.n3527 9.3005
R11127 gnd.n3542 gnd.n3528 9.3005
R11128 gnd.n3541 gnd.n3529 9.3005
R11129 gnd.n3539 gnd.n3530 9.3005
R11130 gnd.n3538 gnd.n3531 9.3005
R11131 gnd.n3536 gnd.n3532 9.3005
R11132 gnd.n3535 gnd.n3533 9.3005
R11133 gnd.n2686 gnd.n2685 9.3005
R11134 gnd.n3610 gnd.n3609 9.3005
R11135 gnd.n3611 gnd.n2684 9.3005
R11136 gnd.n3632 gnd.n3612 9.3005
R11137 gnd.n3631 gnd.n3613 9.3005
R11138 gnd.n3630 gnd.n3614 9.3005
R11139 gnd.n3627 gnd.n3615 9.3005
R11140 gnd.n3626 gnd.n3616 9.3005
R11141 gnd.n3624 gnd.n3617 9.3005
R11142 gnd.n3623 gnd.n3618 9.3005
R11143 gnd.n3621 gnd.n3620 9.3005
R11144 gnd.n3619 gnd.n2638 9.3005
R11145 gnd.n3197 gnd.n3196 9.3005
R11146 gnd.n3087 gnd.n3086 9.3005
R11147 gnd.n3211 gnd.n3210 9.3005
R11148 gnd.n3212 gnd.n3085 9.3005
R11149 gnd.n3214 gnd.n3213 9.3005
R11150 gnd.n3075 gnd.n3074 9.3005
R11151 gnd.n3227 gnd.n3226 9.3005
R11152 gnd.n3228 gnd.n3073 9.3005
R11153 gnd.n3260 gnd.n3229 9.3005
R11154 gnd.n3259 gnd.n3230 9.3005
R11155 gnd.n3258 gnd.n3231 9.3005
R11156 gnd.n3257 gnd.n3232 9.3005
R11157 gnd.n3254 gnd.n3233 9.3005
R11158 gnd.n3253 gnd.n3234 9.3005
R11159 gnd.n3252 gnd.n3235 9.3005
R11160 gnd.n3250 gnd.n3236 9.3005
R11161 gnd.n3249 gnd.n3237 9.3005
R11162 gnd.n3246 gnd.n3238 9.3005
R11163 gnd.n3245 gnd.n3239 9.3005
R11164 gnd.n3244 gnd.n3240 9.3005
R11165 gnd.n3242 gnd.n3241 9.3005
R11166 gnd.n2941 gnd.n2940 9.3005
R11167 gnd.n3358 gnd.n3357 9.3005
R11168 gnd.n3359 gnd.n2939 9.3005
R11169 gnd.n3363 gnd.n3360 9.3005
R11170 gnd.n3362 gnd.n3361 9.3005
R11171 gnd.n2863 gnd.n2862 9.3005
R11172 gnd.n3438 gnd.n3437 9.3005
R11173 gnd.n3195 gnd.n3096 9.3005
R11174 gnd.n3098 gnd.n3097 9.3005
R11175 gnd.n3142 gnd.n3140 9.3005
R11176 gnd.n3143 gnd.n3139 9.3005
R11177 gnd.n3146 gnd.n3135 9.3005
R11178 gnd.n3147 gnd.n3134 9.3005
R11179 gnd.n3150 gnd.n3133 9.3005
R11180 gnd.n3151 gnd.n3132 9.3005
R11181 gnd.n3154 gnd.n3131 9.3005
R11182 gnd.n3155 gnd.n3130 9.3005
R11183 gnd.n3158 gnd.n3129 9.3005
R11184 gnd.n3159 gnd.n3128 9.3005
R11185 gnd.n3162 gnd.n3127 9.3005
R11186 gnd.n3163 gnd.n3126 9.3005
R11187 gnd.n3166 gnd.n3125 9.3005
R11188 gnd.n3167 gnd.n3124 9.3005
R11189 gnd.n3170 gnd.n3123 9.3005
R11190 gnd.n3171 gnd.n3122 9.3005
R11191 gnd.n3174 gnd.n3121 9.3005
R11192 gnd.n3175 gnd.n3120 9.3005
R11193 gnd.n3178 gnd.n3119 9.3005
R11194 gnd.n3179 gnd.n3118 9.3005
R11195 gnd.n3182 gnd.n3117 9.3005
R11196 gnd.n3184 gnd.n3116 9.3005
R11197 gnd.n3185 gnd.n3115 9.3005
R11198 gnd.n3186 gnd.n3114 9.3005
R11199 gnd.n3187 gnd.n3113 9.3005
R11200 gnd.n3194 gnd.n3193 9.3005
R11201 gnd.n3203 gnd.n3202 9.3005
R11202 gnd.n3204 gnd.n3090 9.3005
R11203 gnd.n3206 gnd.n3205 9.3005
R11204 gnd.n3081 gnd.n3080 9.3005
R11205 gnd.n3219 gnd.n3218 9.3005
R11206 gnd.n3220 gnd.n3079 9.3005
R11207 gnd.n3222 gnd.n3221 9.3005
R11208 gnd.n3068 gnd.n3067 9.3005
R11209 gnd.n3265 gnd.n3264 9.3005
R11210 gnd.n3266 gnd.n3022 9.3005
R11211 gnd.n3270 gnd.n3268 9.3005
R11212 gnd.n3269 gnd.n3001 9.3005
R11213 gnd.n3288 gnd.n3000 9.3005
R11214 gnd.n3291 gnd.n3290 9.3005
R11215 gnd.n2994 gnd.n2993 9.3005
R11216 gnd.n3302 gnd.n3300 9.3005
R11217 gnd.n3301 gnd.n2975 9.3005
R11218 gnd.n3319 gnd.n2974 9.3005
R11219 gnd.n3322 gnd.n3321 9.3005
R11220 gnd.n2969 gnd.n2964 9.3005
R11221 gnd.n3332 gnd.n3331 9.3005
R11222 gnd.n2967 gnd.n2947 9.3005
R11223 gnd.n3353 gnd.n2948 9.3005
R11224 gnd.n3352 gnd.n3351 9.3005
R11225 gnd.n2950 gnd.n2926 9.3005
R11226 gnd.n3384 gnd.n3383 9.3005
R11227 gnd.n3386 gnd.n2871 9.3005
R11228 gnd.n3433 gnd.n2872 9.3005
R11229 gnd.n3432 gnd.n2873 9.3005
R11230 gnd.n3431 gnd.n2874 9.3005
R11231 gnd.n3397 gnd.n2875 9.3005
R11232 gnd.n3399 gnd.n2893 9.3005
R11233 gnd.n3419 gnd.n2894 9.3005
R11234 gnd.n3418 gnd.n2895 9.3005
R11235 gnd.n3417 gnd.n2896 9.3005
R11236 gnd.n3408 gnd.n2897 9.3005
R11237 gnd.n3409 gnd.n2780 9.3005
R11238 gnd.n3475 gnd.n3474 9.3005
R11239 gnd.n3476 gnd.n2773 9.3005
R11240 gnd.n3486 gnd.n3485 9.3005
R11241 gnd.n3488 gnd.n2769 9.3005
R11242 gnd.n3498 gnd.n2770 9.3005
R11243 gnd.n3497 gnd.n3496 9.3005
R11244 gnd.n3494 gnd.n2748 9.3005
R11245 gnd.n3520 gnd.n2749 9.3005
R11246 gnd.n3519 gnd.n3518 9.3005
R11247 gnd.n2751 gnd.n2725 9.3005
R11248 gnd.n3560 gnd.n3559 9.3005
R11249 gnd.n3561 gnd.n2718 9.3005
R11250 gnd.n3571 gnd.n3570 9.3005
R11251 gnd.n3573 gnd.n2714 9.3005
R11252 gnd.n3583 gnd.n2715 9.3005
R11253 gnd.n3582 gnd.n3581 9.3005
R11254 gnd.n3579 gnd.n2693 9.3005
R11255 gnd.n3605 gnd.n2694 9.3005
R11256 gnd.n3604 gnd.n3603 9.3005
R11257 gnd.n2696 gnd.n2671 9.3005
R11258 gnd.n3649 gnd.n3648 9.3005
R11259 gnd.n3650 gnd.n2664 9.3005
R11260 gnd.n3661 gnd.n3660 9.3005
R11261 gnd.n3919 gnd.n2660 9.3005
R11262 gnd.n3927 gnd.n2661 9.3005
R11263 gnd.n3926 gnd.n3925 9.3005
R11264 gnd.n2642 gnd.n2641 9.3005
R11265 gnd.n3950 gnd.n3949 9.3005
R11266 gnd.n3092 gnd.n3091 9.3005
R11267 gnd.n6644 gnd.n768 9.3005
R11268 gnd.n6646 gnd.n6645 9.3005
R11269 gnd.n764 gnd.n763 9.3005
R11270 gnd.n6653 gnd.n6652 9.3005
R11271 gnd.n6654 gnd.n762 9.3005
R11272 gnd.n6656 gnd.n6655 9.3005
R11273 gnd.n758 gnd.n757 9.3005
R11274 gnd.n6663 gnd.n6662 9.3005
R11275 gnd.n6664 gnd.n756 9.3005
R11276 gnd.n6666 gnd.n6665 9.3005
R11277 gnd.n752 gnd.n751 9.3005
R11278 gnd.n6673 gnd.n6672 9.3005
R11279 gnd.n6674 gnd.n750 9.3005
R11280 gnd.n6676 gnd.n6675 9.3005
R11281 gnd.n746 gnd.n745 9.3005
R11282 gnd.n6683 gnd.n6682 9.3005
R11283 gnd.n6684 gnd.n744 9.3005
R11284 gnd.n6686 gnd.n6685 9.3005
R11285 gnd.n740 gnd.n739 9.3005
R11286 gnd.n6693 gnd.n6692 9.3005
R11287 gnd.n6694 gnd.n738 9.3005
R11288 gnd.n6696 gnd.n6695 9.3005
R11289 gnd.n734 gnd.n733 9.3005
R11290 gnd.n6703 gnd.n6702 9.3005
R11291 gnd.n6704 gnd.n732 9.3005
R11292 gnd.n6706 gnd.n6705 9.3005
R11293 gnd.n728 gnd.n727 9.3005
R11294 gnd.n6713 gnd.n6712 9.3005
R11295 gnd.n6714 gnd.n726 9.3005
R11296 gnd.n6716 gnd.n6715 9.3005
R11297 gnd.n722 gnd.n721 9.3005
R11298 gnd.n6723 gnd.n6722 9.3005
R11299 gnd.n6724 gnd.n720 9.3005
R11300 gnd.n6726 gnd.n6725 9.3005
R11301 gnd.n716 gnd.n715 9.3005
R11302 gnd.n6733 gnd.n6732 9.3005
R11303 gnd.n6734 gnd.n714 9.3005
R11304 gnd.n6736 gnd.n6735 9.3005
R11305 gnd.n710 gnd.n709 9.3005
R11306 gnd.n6743 gnd.n6742 9.3005
R11307 gnd.n6744 gnd.n708 9.3005
R11308 gnd.n6746 gnd.n6745 9.3005
R11309 gnd.n704 gnd.n703 9.3005
R11310 gnd.n6753 gnd.n6752 9.3005
R11311 gnd.n6754 gnd.n702 9.3005
R11312 gnd.n6756 gnd.n6755 9.3005
R11313 gnd.n698 gnd.n697 9.3005
R11314 gnd.n6763 gnd.n6762 9.3005
R11315 gnd.n6764 gnd.n696 9.3005
R11316 gnd.n6766 gnd.n6765 9.3005
R11317 gnd.n692 gnd.n691 9.3005
R11318 gnd.n6773 gnd.n6772 9.3005
R11319 gnd.n6774 gnd.n690 9.3005
R11320 gnd.n6776 gnd.n6775 9.3005
R11321 gnd.n686 gnd.n685 9.3005
R11322 gnd.n6783 gnd.n6782 9.3005
R11323 gnd.n6784 gnd.n684 9.3005
R11324 gnd.n6786 gnd.n6785 9.3005
R11325 gnd.n680 gnd.n679 9.3005
R11326 gnd.n6793 gnd.n6792 9.3005
R11327 gnd.n6794 gnd.n678 9.3005
R11328 gnd.n6796 gnd.n6795 9.3005
R11329 gnd.n674 gnd.n673 9.3005
R11330 gnd.n6803 gnd.n6802 9.3005
R11331 gnd.n6804 gnd.n672 9.3005
R11332 gnd.n6806 gnd.n6805 9.3005
R11333 gnd.n668 gnd.n667 9.3005
R11334 gnd.n6813 gnd.n6812 9.3005
R11335 gnd.n6814 gnd.n666 9.3005
R11336 gnd.n6816 gnd.n6815 9.3005
R11337 gnd.n662 gnd.n661 9.3005
R11338 gnd.n6823 gnd.n6822 9.3005
R11339 gnd.n6824 gnd.n660 9.3005
R11340 gnd.n6826 gnd.n6825 9.3005
R11341 gnd.n656 gnd.n655 9.3005
R11342 gnd.n6833 gnd.n6832 9.3005
R11343 gnd.n6834 gnd.n654 9.3005
R11344 gnd.n6836 gnd.n6835 9.3005
R11345 gnd.n650 gnd.n649 9.3005
R11346 gnd.n6843 gnd.n6842 9.3005
R11347 gnd.n6844 gnd.n648 9.3005
R11348 gnd.n6846 gnd.n6845 9.3005
R11349 gnd.n644 gnd.n643 9.3005
R11350 gnd.n6853 gnd.n6852 9.3005
R11351 gnd.n6854 gnd.n642 9.3005
R11352 gnd.n6856 gnd.n6855 9.3005
R11353 gnd.n638 gnd.n637 9.3005
R11354 gnd.n6863 gnd.n6862 9.3005
R11355 gnd.n6864 gnd.n636 9.3005
R11356 gnd.n6866 gnd.n6865 9.3005
R11357 gnd.n632 gnd.n631 9.3005
R11358 gnd.n6873 gnd.n6872 9.3005
R11359 gnd.n6874 gnd.n630 9.3005
R11360 gnd.n6876 gnd.n6875 9.3005
R11361 gnd.n626 gnd.n625 9.3005
R11362 gnd.n6883 gnd.n6882 9.3005
R11363 gnd.n6884 gnd.n624 9.3005
R11364 gnd.n6886 gnd.n6885 9.3005
R11365 gnd.n620 gnd.n619 9.3005
R11366 gnd.n6893 gnd.n6892 9.3005
R11367 gnd.n6894 gnd.n618 9.3005
R11368 gnd.n6896 gnd.n6895 9.3005
R11369 gnd.n614 gnd.n613 9.3005
R11370 gnd.n6903 gnd.n6902 9.3005
R11371 gnd.n6904 gnd.n612 9.3005
R11372 gnd.n6906 gnd.n6905 9.3005
R11373 gnd.n608 gnd.n607 9.3005
R11374 gnd.n6913 gnd.n6912 9.3005
R11375 gnd.n6914 gnd.n606 9.3005
R11376 gnd.n6916 gnd.n6915 9.3005
R11377 gnd.n602 gnd.n601 9.3005
R11378 gnd.n6923 gnd.n6922 9.3005
R11379 gnd.n6924 gnd.n600 9.3005
R11380 gnd.n6926 gnd.n6925 9.3005
R11381 gnd.n596 gnd.n595 9.3005
R11382 gnd.n6933 gnd.n6932 9.3005
R11383 gnd.n6934 gnd.n594 9.3005
R11384 gnd.n6936 gnd.n6935 9.3005
R11385 gnd.n590 gnd.n589 9.3005
R11386 gnd.n6943 gnd.n6942 9.3005
R11387 gnd.n6944 gnd.n588 9.3005
R11388 gnd.n6946 gnd.n6945 9.3005
R11389 gnd.n584 gnd.n583 9.3005
R11390 gnd.n6953 gnd.n6952 9.3005
R11391 gnd.n6954 gnd.n582 9.3005
R11392 gnd.n6956 gnd.n6955 9.3005
R11393 gnd.n578 gnd.n577 9.3005
R11394 gnd.n6963 gnd.n6962 9.3005
R11395 gnd.n6964 gnd.n576 9.3005
R11396 gnd.n6966 gnd.n6965 9.3005
R11397 gnd.n572 gnd.n571 9.3005
R11398 gnd.n6973 gnd.n6972 9.3005
R11399 gnd.n6974 gnd.n570 9.3005
R11400 gnd.n6976 gnd.n6975 9.3005
R11401 gnd.n566 gnd.n565 9.3005
R11402 gnd.n6983 gnd.n6982 9.3005
R11403 gnd.n6984 gnd.n564 9.3005
R11404 gnd.n6986 gnd.n6985 9.3005
R11405 gnd.n560 gnd.n559 9.3005
R11406 gnd.n6993 gnd.n6992 9.3005
R11407 gnd.n6994 gnd.n558 9.3005
R11408 gnd.n6996 gnd.n6995 9.3005
R11409 gnd.n554 gnd.n553 9.3005
R11410 gnd.n7003 gnd.n7002 9.3005
R11411 gnd.n7004 gnd.n552 9.3005
R11412 gnd.n7006 gnd.n7005 9.3005
R11413 gnd.n548 gnd.n547 9.3005
R11414 gnd.n7013 gnd.n7012 9.3005
R11415 gnd.n7014 gnd.n546 9.3005
R11416 gnd.n7016 gnd.n7015 9.3005
R11417 gnd.n542 gnd.n541 9.3005
R11418 gnd.n7023 gnd.n7022 9.3005
R11419 gnd.n7024 gnd.n540 9.3005
R11420 gnd.n7026 gnd.n7025 9.3005
R11421 gnd.n536 gnd.n535 9.3005
R11422 gnd.n7033 gnd.n7032 9.3005
R11423 gnd.n7034 gnd.n534 9.3005
R11424 gnd.n7036 gnd.n7035 9.3005
R11425 gnd.n530 gnd.n529 9.3005
R11426 gnd.n7043 gnd.n7042 9.3005
R11427 gnd.n7044 gnd.n528 9.3005
R11428 gnd.n7046 gnd.n7045 9.3005
R11429 gnd.n524 gnd.n523 9.3005
R11430 gnd.n7053 gnd.n7052 9.3005
R11431 gnd.n7054 gnd.n522 9.3005
R11432 gnd.n7056 gnd.n7055 9.3005
R11433 gnd.n518 gnd.n517 9.3005
R11434 gnd.n7063 gnd.n7062 9.3005
R11435 gnd.n7066 gnd.n7065 9.3005
R11436 gnd.n512 gnd.n511 9.3005
R11437 gnd.n7073 gnd.n7072 9.3005
R11438 gnd.n7074 gnd.n510 9.3005
R11439 gnd.n7076 gnd.n7075 9.3005
R11440 gnd.n506 gnd.n505 9.3005
R11441 gnd.n7083 gnd.n7082 9.3005
R11442 gnd.n7084 gnd.n504 9.3005
R11443 gnd.n7086 gnd.n7085 9.3005
R11444 gnd.n500 gnd.n499 9.3005
R11445 gnd.n7093 gnd.n7092 9.3005
R11446 gnd.n7094 gnd.n498 9.3005
R11447 gnd.n7096 gnd.n7095 9.3005
R11448 gnd.n494 gnd.n493 9.3005
R11449 gnd.n7103 gnd.n7102 9.3005
R11450 gnd.n7104 gnd.n492 9.3005
R11451 gnd.n7106 gnd.n7105 9.3005
R11452 gnd.n488 gnd.n487 9.3005
R11453 gnd.n7113 gnd.n7112 9.3005
R11454 gnd.n7114 gnd.n486 9.3005
R11455 gnd.n7116 gnd.n7115 9.3005
R11456 gnd.n482 gnd.n481 9.3005
R11457 gnd.n7123 gnd.n7122 9.3005
R11458 gnd.n7124 gnd.n480 9.3005
R11459 gnd.n7126 gnd.n7125 9.3005
R11460 gnd.n476 gnd.n475 9.3005
R11461 gnd.n7133 gnd.n7132 9.3005
R11462 gnd.n7134 gnd.n474 9.3005
R11463 gnd.n7136 gnd.n7135 9.3005
R11464 gnd.n470 gnd.n469 9.3005
R11465 gnd.n7143 gnd.n7142 9.3005
R11466 gnd.n7144 gnd.n468 9.3005
R11467 gnd.n7146 gnd.n7145 9.3005
R11468 gnd.n464 gnd.n463 9.3005
R11469 gnd.n7153 gnd.n7152 9.3005
R11470 gnd.n7154 gnd.n462 9.3005
R11471 gnd.n7156 gnd.n7155 9.3005
R11472 gnd.n458 gnd.n457 9.3005
R11473 gnd.n7163 gnd.n7162 9.3005
R11474 gnd.n7164 gnd.n456 9.3005
R11475 gnd.n7166 gnd.n7165 9.3005
R11476 gnd.n452 gnd.n451 9.3005
R11477 gnd.n7173 gnd.n7172 9.3005
R11478 gnd.n7174 gnd.n450 9.3005
R11479 gnd.n7176 gnd.n7175 9.3005
R11480 gnd.n446 gnd.n445 9.3005
R11481 gnd.n7183 gnd.n7182 9.3005
R11482 gnd.n7184 gnd.n444 9.3005
R11483 gnd.n7186 gnd.n7185 9.3005
R11484 gnd.n440 gnd.n439 9.3005
R11485 gnd.n7193 gnd.n7192 9.3005
R11486 gnd.n7194 gnd.n438 9.3005
R11487 gnd.n7196 gnd.n7195 9.3005
R11488 gnd.n434 gnd.n433 9.3005
R11489 gnd.n7203 gnd.n7202 9.3005
R11490 gnd.n7204 gnd.n432 9.3005
R11491 gnd.n7206 gnd.n7205 9.3005
R11492 gnd.n428 gnd.n427 9.3005
R11493 gnd.n7213 gnd.n7212 9.3005
R11494 gnd.n7214 gnd.n426 9.3005
R11495 gnd.n7216 gnd.n7215 9.3005
R11496 gnd.n422 gnd.n421 9.3005
R11497 gnd.n7223 gnd.n7222 9.3005
R11498 gnd.n7224 gnd.n420 9.3005
R11499 gnd.n7226 gnd.n7225 9.3005
R11500 gnd.n416 gnd.n415 9.3005
R11501 gnd.n7233 gnd.n7232 9.3005
R11502 gnd.n7234 gnd.n414 9.3005
R11503 gnd.n7236 gnd.n7235 9.3005
R11504 gnd.n410 gnd.n409 9.3005
R11505 gnd.n7243 gnd.n7242 9.3005
R11506 gnd.n7244 gnd.n408 9.3005
R11507 gnd.n7246 gnd.n7245 9.3005
R11508 gnd.n404 gnd.n403 9.3005
R11509 gnd.n7253 gnd.n7252 9.3005
R11510 gnd.n7254 gnd.n402 9.3005
R11511 gnd.n7256 gnd.n7255 9.3005
R11512 gnd.n398 gnd.n397 9.3005
R11513 gnd.n7263 gnd.n7262 9.3005
R11514 gnd.n7264 gnd.n396 9.3005
R11515 gnd.n7268 gnd.n7265 9.3005
R11516 gnd.n7267 gnd.n7266 9.3005
R11517 gnd.n392 gnd.n391 9.3005
R11518 gnd.n7276 gnd.n7275 9.3005
R11519 gnd.n7064 gnd.n516 9.3005
R11520 gnd.n7615 gnd.n7614 9.3005
R11521 gnd.n7613 gnd.n84 9.3005
R11522 gnd.n7348 gnd.n87 9.3005
R11523 gnd.n7349 gnd.n7347 9.3005
R11524 gnd.n7351 gnd.n7350 9.3005
R11525 gnd.n7353 gnd.n367 9.3005
R11526 gnd.n7355 gnd.n7354 9.3005
R11527 gnd.n7356 gnd.n366 9.3005
R11528 gnd.n7358 gnd.n7357 9.3005
R11529 gnd.n7360 gnd.n364 9.3005
R11530 gnd.n7362 gnd.n7361 9.3005
R11531 gnd.n7363 gnd.n363 9.3005
R11532 gnd.n7365 gnd.n7364 9.3005
R11533 gnd.n7367 gnd.n361 9.3005
R11534 gnd.n7369 gnd.n7368 9.3005
R11535 gnd.n7370 gnd.n360 9.3005
R11536 gnd.n7372 gnd.n7371 9.3005
R11537 gnd.n7374 gnd.n358 9.3005
R11538 gnd.n7376 gnd.n7375 9.3005
R11539 gnd.n7377 gnd.n357 9.3005
R11540 gnd.n7379 gnd.n7378 9.3005
R11541 gnd.n7381 gnd.n355 9.3005
R11542 gnd.n7383 gnd.n7382 9.3005
R11543 gnd.n7384 gnd.n354 9.3005
R11544 gnd.n7386 gnd.n7385 9.3005
R11545 gnd.n7388 gnd.n352 9.3005
R11546 gnd.n7390 gnd.n7389 9.3005
R11547 gnd.n7421 gnd.n318 9.3005
R11548 gnd.n7420 gnd.n320 9.3005
R11549 gnd.n324 gnd.n321 9.3005
R11550 gnd.n7415 gnd.n325 9.3005
R11551 gnd.n7414 gnd.n326 9.3005
R11552 gnd.n7413 gnd.n327 9.3005
R11553 gnd.n331 gnd.n328 9.3005
R11554 gnd.n7408 gnd.n332 9.3005
R11555 gnd.n7407 gnd.n333 9.3005
R11556 gnd.n7406 gnd.n334 9.3005
R11557 gnd.n338 gnd.n335 9.3005
R11558 gnd.n7401 gnd.n339 9.3005
R11559 gnd.n7400 gnd.n340 9.3005
R11560 gnd.n7399 gnd.n341 9.3005
R11561 gnd.n345 gnd.n342 9.3005
R11562 gnd.n7394 gnd.n346 9.3005
R11563 gnd.n7393 gnd.n7392 9.3005
R11564 gnd.n7391 gnd.n349 9.3005
R11565 gnd.n7423 gnd.n7422 9.3005
R11566 gnd.n7531 gnd.n215 9.3005
R11567 gnd.n7530 gnd.n217 9.3005
R11568 gnd.n221 gnd.n218 9.3005
R11569 gnd.n7525 gnd.n222 9.3005
R11570 gnd.n7524 gnd.n223 9.3005
R11571 gnd.n7523 gnd.n224 9.3005
R11572 gnd.n228 gnd.n225 9.3005
R11573 gnd.n7518 gnd.n229 9.3005
R11574 gnd.n7517 gnd.n230 9.3005
R11575 gnd.n7516 gnd.n231 9.3005
R11576 gnd.n235 gnd.n232 9.3005
R11577 gnd.n7511 gnd.n236 9.3005
R11578 gnd.n7510 gnd.n237 9.3005
R11579 gnd.n7509 gnd.n238 9.3005
R11580 gnd.n242 gnd.n239 9.3005
R11581 gnd.n7504 gnd.n243 9.3005
R11582 gnd.n7503 gnd.n244 9.3005
R11583 gnd.n7499 gnd.n245 9.3005
R11584 gnd.n249 gnd.n246 9.3005
R11585 gnd.n7494 gnd.n250 9.3005
R11586 gnd.n7493 gnd.n251 9.3005
R11587 gnd.n7492 gnd.n252 9.3005
R11588 gnd.n256 gnd.n253 9.3005
R11589 gnd.n7487 gnd.n257 9.3005
R11590 gnd.n7486 gnd.n258 9.3005
R11591 gnd.n7485 gnd.n259 9.3005
R11592 gnd.n263 gnd.n260 9.3005
R11593 gnd.n7480 gnd.n264 9.3005
R11594 gnd.n7479 gnd.n265 9.3005
R11595 gnd.n7478 gnd.n266 9.3005
R11596 gnd.n270 gnd.n267 9.3005
R11597 gnd.n7473 gnd.n271 9.3005
R11598 gnd.n7472 gnd.n272 9.3005
R11599 gnd.n7471 gnd.n273 9.3005
R11600 gnd.n277 gnd.n274 9.3005
R11601 gnd.n7466 gnd.n278 9.3005
R11602 gnd.n7465 gnd.n7464 9.3005
R11603 gnd.n7463 gnd.n279 9.3005
R11604 gnd.n7462 gnd.n7461 9.3005
R11605 gnd.n283 gnd.n282 9.3005
R11606 gnd.n288 gnd.n286 9.3005
R11607 gnd.n7454 gnd.n289 9.3005
R11608 gnd.n7453 gnd.n290 9.3005
R11609 gnd.n7452 gnd.n291 9.3005
R11610 gnd.n295 gnd.n292 9.3005
R11611 gnd.n7447 gnd.n296 9.3005
R11612 gnd.n7446 gnd.n297 9.3005
R11613 gnd.n7445 gnd.n298 9.3005
R11614 gnd.n302 gnd.n299 9.3005
R11615 gnd.n7440 gnd.n303 9.3005
R11616 gnd.n7439 gnd.n304 9.3005
R11617 gnd.n7438 gnd.n305 9.3005
R11618 gnd.n309 gnd.n306 9.3005
R11619 gnd.n7433 gnd.n310 9.3005
R11620 gnd.n7432 gnd.n311 9.3005
R11621 gnd.n7431 gnd.n312 9.3005
R11622 gnd.n317 gnd.n315 9.3005
R11623 gnd.n7426 gnd.n7425 9.3005
R11624 gnd.n7533 gnd.n7532 9.3005
R11625 gnd.n5957 gnd.n5956 9.3005
R11626 gnd.n1480 gnd.n1479 9.3005
R11627 gnd.n1504 gnd.n1503 9.3005
R11628 gnd.n5944 gnd.n1505 9.3005
R11629 gnd.n5943 gnd.n1506 9.3005
R11630 gnd.n5942 gnd.n1507 9.3005
R11631 gnd.n5748 gnd.n1508 9.3005
R11632 gnd.n5932 gnd.n1525 9.3005
R11633 gnd.n5931 gnd.n1526 9.3005
R11634 gnd.n5930 gnd.n1527 9.3005
R11635 gnd.n5754 gnd.n1528 9.3005
R11636 gnd.n5920 gnd.n1545 9.3005
R11637 gnd.n5919 gnd.n1546 9.3005
R11638 gnd.n5918 gnd.n1547 9.3005
R11639 gnd.n5834 gnd.n1548 9.3005
R11640 gnd.n5908 gnd.n1565 9.3005
R11641 gnd.n5907 gnd.n1566 9.3005
R11642 gnd.n5906 gnd.n1567 9.3005
R11643 gnd.n5849 gnd.n1568 9.3005
R11644 gnd.n5896 gnd.n1585 9.3005
R11645 gnd.n5895 gnd.n1586 9.3005
R11646 gnd.n5894 gnd.n1587 9.3005
R11647 gnd.n5852 gnd.n1588 9.3005
R11648 gnd.n379 gnd.n378 9.3005
R11649 gnd.n7290 gnd.n7289 9.3005
R11650 gnd.n7291 gnd.n372 9.3005
R11651 gnd.n7298 gnd.n373 9.3005
R11652 gnd.n7299 gnd.n371 9.3005
R11653 gnd.n7302 gnd.n7301 9.3005
R11654 gnd.n7303 gnd.n110 9.3005
R11655 gnd.n7601 gnd.n111 9.3005
R11656 gnd.n7600 gnd.n112 9.3005
R11657 gnd.n7599 gnd.n113 9.3005
R11658 gnd.n7304 gnd.n114 9.3005
R11659 gnd.n7589 gnd.n128 9.3005
R11660 gnd.n7588 gnd.n129 9.3005
R11661 gnd.n7587 gnd.n130 9.3005
R11662 gnd.n7305 gnd.n131 9.3005
R11663 gnd.n7577 gnd.n148 9.3005
R11664 gnd.n7576 gnd.n149 9.3005
R11665 gnd.n7575 gnd.n150 9.3005
R11666 gnd.n7306 gnd.n151 9.3005
R11667 gnd.n7565 gnd.n166 9.3005
R11668 gnd.n7564 gnd.n167 9.3005
R11669 gnd.n7563 gnd.n168 9.3005
R11670 gnd.n7307 gnd.n169 9.3005
R11671 gnd.n7553 gnd.n186 9.3005
R11672 gnd.n7552 gnd.n187 9.3005
R11673 gnd.n7551 gnd.n188 9.3005
R11674 gnd.n7308 gnd.n189 9.3005
R11675 gnd.n7541 gnd.n205 9.3005
R11676 gnd.n7540 gnd.n206 9.3005
R11677 gnd.n7539 gnd.n207 9.3005
R11678 gnd.n5958 gnd.n1478 9.3005
R11679 gnd.n5956 gnd.n5955 9.3005
R11680 gnd.n5954 gnd.n1480 9.3005
R11681 gnd.n1504 gnd.n1481 9.3005
R11682 gnd.n5743 gnd.n1505 9.3005
R11683 gnd.n5746 gnd.n1506 9.3005
R11684 gnd.n5747 gnd.n1507 9.3005
R11685 gnd.n5752 gnd.n5748 9.3005
R11686 gnd.n5753 gnd.n1525 9.3005
R11687 gnd.n5757 gnd.n1526 9.3005
R11688 gnd.n5756 gnd.n1527 9.3005
R11689 gnd.n5755 gnd.n5754 9.3005
R11690 gnd.n1614 gnd.n1545 9.3005
R11691 gnd.n5832 gnd.n1546 9.3005
R11692 gnd.n5833 gnd.n1547 9.3005
R11693 gnd.n5835 gnd.n5834 9.3005
R11694 gnd.n1609 gnd.n1565 9.3005
R11695 gnd.n5847 gnd.n1566 9.3005
R11696 gnd.n5848 gnd.n1567 9.3005
R11697 gnd.n5850 gnd.n5849 9.3005
R11698 gnd.n5851 gnd.n1585 9.3005
R11699 gnd.n5857 gnd.n1586 9.3005
R11700 gnd.n5856 gnd.n1587 9.3005
R11701 gnd.n5855 gnd.n5852 9.3005
R11702 gnd.n5854 gnd.n378 9.3005
R11703 gnd.n7290 gnd.n377 9.3005
R11704 gnd.n7292 gnd.n7291 9.3005
R11705 gnd.n7294 gnd.n373 9.3005
R11706 gnd.n7293 gnd.n371 9.3005
R11707 gnd.n7302 gnd.n370 9.3005
R11708 gnd.n7343 gnd.n7303 9.3005
R11709 gnd.n7342 gnd.n111 9.3005
R11710 gnd.n7341 gnd.n112 9.3005
R11711 gnd.n7339 gnd.n113 9.3005
R11712 gnd.n7338 gnd.n7304 9.3005
R11713 gnd.n7336 gnd.n128 9.3005
R11714 gnd.n7335 gnd.n129 9.3005
R11715 gnd.n7333 gnd.n130 9.3005
R11716 gnd.n7332 gnd.n7305 9.3005
R11717 gnd.n7330 gnd.n148 9.3005
R11718 gnd.n7329 gnd.n149 9.3005
R11719 gnd.n7327 gnd.n150 9.3005
R11720 gnd.n7326 gnd.n7306 9.3005
R11721 gnd.n7324 gnd.n166 9.3005
R11722 gnd.n7323 gnd.n167 9.3005
R11723 gnd.n7321 gnd.n168 9.3005
R11724 gnd.n7320 gnd.n7307 9.3005
R11725 gnd.n7318 gnd.n186 9.3005
R11726 gnd.n7317 gnd.n187 9.3005
R11727 gnd.n7315 gnd.n188 9.3005
R11728 gnd.n7314 gnd.n7308 9.3005
R11729 gnd.n7312 gnd.n205 9.3005
R11730 gnd.n7311 gnd.n206 9.3005
R11731 gnd.n7309 gnd.n207 9.3005
R11732 gnd.n1478 gnd.n1472 9.3005
R11733 gnd.n5968 gnd.n5967 9.3005
R11734 gnd.n5971 gnd.n1470 9.3005
R11735 gnd.n5972 gnd.n1469 9.3005
R11736 gnd.n5975 gnd.n1468 9.3005
R11737 gnd.n5976 gnd.n1467 9.3005
R11738 gnd.n5979 gnd.n1466 9.3005
R11739 gnd.n5980 gnd.n1465 9.3005
R11740 gnd.n5983 gnd.n1464 9.3005
R11741 gnd.n5984 gnd.n1463 9.3005
R11742 gnd.n5987 gnd.n1462 9.3005
R11743 gnd.n5988 gnd.n1461 9.3005
R11744 gnd.n5991 gnd.n1460 9.3005
R11745 gnd.n5992 gnd.n1459 9.3005
R11746 gnd.n5995 gnd.n1458 9.3005
R11747 gnd.n5996 gnd.n1457 9.3005
R11748 gnd.n5999 gnd.n1456 9.3005
R11749 gnd.n6000 gnd.n1455 9.3005
R11750 gnd.n6003 gnd.n1454 9.3005
R11751 gnd.n6004 gnd.n1453 9.3005
R11752 gnd.n6007 gnd.n1452 9.3005
R11753 gnd.n6011 gnd.n1448 9.3005
R11754 gnd.n6012 gnd.n1447 9.3005
R11755 gnd.n6015 gnd.n1446 9.3005
R11756 gnd.n6016 gnd.n1445 9.3005
R11757 gnd.n6019 gnd.n1444 9.3005
R11758 gnd.n6020 gnd.n1443 9.3005
R11759 gnd.n6023 gnd.n1442 9.3005
R11760 gnd.n6024 gnd.n1441 9.3005
R11761 gnd.n6027 gnd.n1440 9.3005
R11762 gnd.n6029 gnd.n1436 9.3005
R11763 gnd.n6032 gnd.n1435 9.3005
R11764 gnd.n6033 gnd.n1434 9.3005
R11765 gnd.n6036 gnd.n1433 9.3005
R11766 gnd.n6037 gnd.n1432 9.3005
R11767 gnd.n6040 gnd.n1431 9.3005
R11768 gnd.n6041 gnd.n1430 9.3005
R11769 gnd.n6044 gnd.n1429 9.3005
R11770 gnd.n6046 gnd.n1426 9.3005
R11771 gnd.n6049 gnd.n1425 9.3005
R11772 gnd.n6050 gnd.n1424 9.3005
R11773 gnd.n6053 gnd.n1423 9.3005
R11774 gnd.n6054 gnd.n1422 9.3005
R11775 gnd.n6057 gnd.n1421 9.3005
R11776 gnd.n6058 gnd.n1420 9.3005
R11777 gnd.n6061 gnd.n1419 9.3005
R11778 gnd.n6062 gnd.n1418 9.3005
R11779 gnd.n6065 gnd.n1417 9.3005
R11780 gnd.n6066 gnd.n1416 9.3005
R11781 gnd.n6069 gnd.n1415 9.3005
R11782 gnd.n6070 gnd.n1414 9.3005
R11783 gnd.n6073 gnd.n1413 9.3005
R11784 gnd.n6075 gnd.n1412 9.3005
R11785 gnd.n6076 gnd.n1411 9.3005
R11786 gnd.n6077 gnd.n1410 9.3005
R11787 gnd.n6078 gnd.n1409 9.3005
R11788 gnd.n6008 gnd.n1449 9.3005
R11789 gnd.n5966 gnd.n5963 9.3005
R11790 gnd.n1491 gnd.n1488 9.3005
R11791 gnd.n5950 gnd.n1492 9.3005
R11792 gnd.n5949 gnd.n1493 9.3005
R11793 gnd.n5948 gnd.n1494 9.3005
R11794 gnd.n1514 gnd.n1495 9.3005
R11795 gnd.n5938 gnd.n1515 9.3005
R11796 gnd.n5937 gnd.n1516 9.3005
R11797 gnd.n5936 gnd.n1517 9.3005
R11798 gnd.n1535 gnd.n1518 9.3005
R11799 gnd.n5926 gnd.n1536 9.3005
R11800 gnd.n5925 gnd.n1537 9.3005
R11801 gnd.n5924 gnd.n1538 9.3005
R11802 gnd.n1554 gnd.n1539 9.3005
R11803 gnd.n5914 gnd.n1555 9.3005
R11804 gnd.n5913 gnd.n1556 9.3005
R11805 gnd.n5912 gnd.n1557 9.3005
R11806 gnd.n1575 gnd.n1558 9.3005
R11807 gnd.n5902 gnd.n1576 9.3005
R11808 gnd.n5901 gnd.n1577 9.3005
R11809 gnd.n5900 gnd.n1578 9.3005
R11810 gnd.n1579 gnd.n97 9.3005
R11811 gnd.n102 gnd.n96 9.3005
R11812 gnd.n7595 gnd.n119 9.3005
R11813 gnd.n7594 gnd.n120 9.3005
R11814 gnd.n7593 gnd.n121 9.3005
R11815 gnd.n138 gnd.n122 9.3005
R11816 gnd.n7583 gnd.n139 9.3005
R11817 gnd.n7582 gnd.n140 9.3005
R11818 gnd.n7581 gnd.n141 9.3005
R11819 gnd.n156 gnd.n142 9.3005
R11820 gnd.n7571 gnd.n157 9.3005
R11821 gnd.n7570 gnd.n158 9.3005
R11822 gnd.n7569 gnd.n159 9.3005
R11823 gnd.n176 gnd.n160 9.3005
R11824 gnd.n7559 gnd.n177 9.3005
R11825 gnd.n7558 gnd.n178 9.3005
R11826 gnd.n7557 gnd.n179 9.3005
R11827 gnd.n196 gnd.n180 9.3005
R11828 gnd.n7547 gnd.n197 9.3005
R11829 gnd.n7546 gnd.n198 9.3005
R11830 gnd.n7545 gnd.n199 9.3005
R11831 gnd.n214 gnd.n200 9.3005
R11832 gnd.n7535 gnd.n7534 9.3005
R11833 gnd.n1490 gnd.n1489 9.3005
R11834 gnd.n7606 gnd.n100 9.3005
R11835 gnd.n7606 gnd.n7605 9.3005
R11836 gnd.n5881 gnd.n5880 9.3005
R11837 gnd.n5882 gnd.n1599 9.3005
R11838 gnd.n5885 gnd.n5884 9.3005
R11839 gnd.n5883 gnd.n389 9.3005
R11840 gnd.n7279 gnd.n390 9.3005
R11841 gnd.n7278 gnd.n7277 9.3005
R11842 gnd.n4560 gnd.n4543 9.3005
R11843 gnd.n4546 gnd.n4544 9.3005
R11844 gnd.n4556 gnd.n4547 9.3005
R11845 gnd.n4555 gnd.n4548 9.3005
R11846 gnd.n4554 gnd.n4549 9.3005
R11847 gnd.n4552 gnd.n4551 9.3005
R11848 gnd.n4550 gnd.n2402 9.3005
R11849 gnd.n2400 gnd.n2399 9.3005
R11850 gnd.n4630 gnd.n4629 9.3005
R11851 gnd.n4631 gnd.n2398 9.3005
R11852 gnd.n4633 gnd.n4632 9.3005
R11853 gnd.n2396 gnd.n2395 9.3005
R11854 gnd.n4638 gnd.n4637 9.3005
R11855 gnd.n4639 gnd.n2394 9.3005
R11856 gnd.n4669 gnd.n4640 9.3005
R11857 gnd.n4668 gnd.n4641 9.3005
R11858 gnd.n4667 gnd.n4642 9.3005
R11859 gnd.n4645 gnd.n4643 9.3005
R11860 gnd.n4663 gnd.n4646 9.3005
R11861 gnd.n4662 gnd.n4647 9.3005
R11862 gnd.n4661 gnd.n4648 9.3005
R11863 gnd.n4652 gnd.n4649 9.3005
R11864 gnd.n4656 gnd.n4653 9.3005
R11865 gnd.n4655 gnd.n4654 9.3005
R11866 gnd.n2118 gnd.n2117 9.3005
R11867 gnd.n4777 gnd.n4776 9.3005
R11868 gnd.n4778 gnd.n2116 9.3005
R11869 gnd.n4780 gnd.n4779 9.3005
R11870 gnd.n2105 gnd.n2104 9.3005
R11871 gnd.n4793 gnd.n4792 9.3005
R11872 gnd.n4794 gnd.n2103 9.3005
R11873 gnd.n4796 gnd.n4795 9.3005
R11874 gnd.n2091 gnd.n2090 9.3005
R11875 gnd.n4809 gnd.n4808 9.3005
R11876 gnd.n4810 gnd.n2089 9.3005
R11877 gnd.n4812 gnd.n4811 9.3005
R11878 gnd.n2076 gnd.n2075 9.3005
R11879 gnd.n4825 gnd.n4824 9.3005
R11880 gnd.n4826 gnd.n2074 9.3005
R11881 gnd.n4828 gnd.n4827 9.3005
R11882 gnd.n2062 gnd.n2061 9.3005
R11883 gnd.n4841 gnd.n4840 9.3005
R11884 gnd.n4842 gnd.n2060 9.3005
R11885 gnd.n4844 gnd.n4843 9.3005
R11886 gnd.n2047 gnd.n2046 9.3005
R11887 gnd.n4871 gnd.n4870 9.3005
R11888 gnd.n4872 gnd.n2045 9.3005
R11889 gnd.n4880 gnd.n4873 9.3005
R11890 gnd.n4879 gnd.n4874 9.3005
R11891 gnd.n4878 gnd.n4876 9.3005
R11892 gnd.n4875 gnd.n1189 9.3005
R11893 gnd.n6270 gnd.n1190 9.3005
R11894 gnd.n6269 gnd.n1191 9.3005
R11895 gnd.n6268 gnd.n1192 9.3005
R11896 gnd.n5029 gnd.n1193 9.3005
R11897 gnd.n5030 gnd.n5028 9.3005
R11898 gnd.n5032 gnd.n5031 9.3005
R11899 gnd.n2017 gnd.n2016 9.3005
R11900 gnd.n5058 gnd.n5057 9.3005
R11901 gnd.n5059 gnd.n2015 9.3005
R11902 gnd.n5063 gnd.n5060 9.3005
R11903 gnd.n5062 gnd.n5061 9.3005
R11904 gnd.n1989 gnd.n1988 9.3005
R11905 gnd.n5096 gnd.n5095 9.3005
R11906 gnd.n5097 gnd.n1987 9.3005
R11907 gnd.n5105 gnd.n5098 9.3005
R11908 gnd.n5104 gnd.n5099 9.3005
R11909 gnd.n5103 gnd.n5101 9.3005
R11910 gnd.n5100 gnd.n1961 9.3005
R11911 gnd.n5166 gnd.n1962 9.3005
R11912 gnd.n5165 gnd.n1963 9.3005
R11913 gnd.n5164 gnd.n1964 9.3005
R11914 gnd.n1939 gnd.n1938 9.3005
R11915 gnd.n5197 gnd.n5196 9.3005
R11916 gnd.n5198 gnd.n1937 9.3005
R11917 gnd.n5202 gnd.n5199 9.3005
R11918 gnd.n5201 gnd.n5200 9.3005
R11919 gnd.n1911 gnd.n1910 9.3005
R11920 gnd.n5235 gnd.n5234 9.3005
R11921 gnd.n5236 gnd.n1909 9.3005
R11922 gnd.n5238 gnd.n5237 9.3005
R11923 gnd.n1885 gnd.n1884 9.3005
R11924 gnd.n5272 gnd.n5271 9.3005
R11925 gnd.n5273 gnd.n1883 9.3005
R11926 gnd.n5277 gnd.n5274 9.3005
R11927 gnd.n5276 gnd.n5275 9.3005
R11928 gnd.n1858 gnd.n1857 9.3005
R11929 gnd.n5321 gnd.n5320 9.3005
R11930 gnd.n5322 gnd.n1856 9.3005
R11931 gnd.n5326 gnd.n5323 9.3005
R11932 gnd.n5325 gnd.n5324 9.3005
R11933 gnd.n1836 gnd.n1835 9.3005
R11934 gnd.n5362 gnd.n5361 9.3005
R11935 gnd.n5363 gnd.n1834 9.3005
R11936 gnd.n5367 gnd.n5364 9.3005
R11937 gnd.n5366 gnd.n5365 9.3005
R11938 gnd.n1806 gnd.n1805 9.3005
R11939 gnd.n5402 gnd.n5401 9.3005
R11940 gnd.n5403 gnd.n1804 9.3005
R11941 gnd.n5405 gnd.n5404 9.3005
R11942 gnd.n1782 gnd.n1781 9.3005
R11943 gnd.n5445 gnd.n5444 9.3005
R11944 gnd.n5446 gnd.n1780 9.3005
R11945 gnd.n5450 gnd.n5447 9.3005
R11946 gnd.n5449 gnd.n5448 9.3005
R11947 gnd.n1726 gnd.n1725 9.3005
R11948 gnd.n5621 gnd.n5620 9.3005
R11949 gnd.n5622 gnd.n1724 9.3005
R11950 gnd.n5624 gnd.n5623 9.3005
R11951 gnd.n1715 gnd.n1714 9.3005
R11952 gnd.n5638 gnd.n5637 9.3005
R11953 gnd.n5639 gnd.n1713 9.3005
R11954 gnd.n5641 gnd.n5640 9.3005
R11955 gnd.n1703 gnd.n1702 9.3005
R11956 gnd.n5655 gnd.n5654 9.3005
R11957 gnd.n5656 gnd.n1701 9.3005
R11958 gnd.n5658 gnd.n5657 9.3005
R11959 gnd.n1691 gnd.n1690 9.3005
R11960 gnd.n5672 gnd.n5671 9.3005
R11961 gnd.n5673 gnd.n1689 9.3005
R11962 gnd.n5675 gnd.n5674 9.3005
R11963 gnd.n1679 gnd.n1678 9.3005
R11964 gnd.n5689 gnd.n5688 9.3005
R11965 gnd.n5690 gnd.n1677 9.3005
R11966 gnd.n5695 gnd.n5691 9.3005
R11967 gnd.n5694 gnd.n5693 9.3005
R11968 gnd.n5692 gnd.n1667 9.3005
R11969 gnd.n5709 gnd.n1666 9.3005
R11970 gnd.n5711 gnd.n5710 9.3005
R11971 gnd.n5712 gnd.n1665 9.3005
R11972 gnd.n5725 gnd.n5713 9.3005
R11973 gnd.n5724 gnd.n5714 9.3005
R11974 gnd.n5723 gnd.n5715 9.3005
R11975 gnd.n5717 gnd.n5716 9.3005
R11976 gnd.n5719 gnd.n5718 9.3005
R11977 gnd.n1631 gnd.n1630 9.3005
R11978 gnd.n5780 gnd.n5779 9.3005
R11979 gnd.n5781 gnd.n1629 9.3005
R11980 gnd.n5783 gnd.n5782 9.3005
R11981 gnd.n1627 gnd.n1626 9.3005
R11982 gnd.n5788 gnd.n5787 9.3005
R11983 gnd.n5789 gnd.n1625 9.3005
R11984 gnd.n5791 gnd.n5790 9.3005
R11985 gnd.n1623 gnd.n1622 9.3005
R11986 gnd.n5796 gnd.n5795 9.3005
R11987 gnd.n5797 gnd.n1621 9.3005
R11988 gnd.n5819 gnd.n5798 9.3005
R11989 gnd.n5818 gnd.n5799 9.3005
R11990 gnd.n5817 gnd.n5800 9.3005
R11991 gnd.n5803 gnd.n5801 9.3005
R11992 gnd.n5813 gnd.n5804 9.3005
R11993 gnd.n5812 gnd.n5805 9.3005
R11994 gnd.n5811 gnd.n5806 9.3005
R11995 gnd.n5809 gnd.n5808 9.3005
R11996 gnd.n5807 gnd.n1603 9.3005
R11997 gnd.n1601 gnd.n1600 9.3005
R11998 gnd.n4196 gnd.n4165 9.3005
R11999 gnd.n4195 gnd.n4166 9.3005
R12000 gnd.n4193 gnd.n4167 9.3005
R12001 gnd.n4192 gnd.n4168 9.3005
R12002 gnd.n4190 gnd.n4169 9.3005
R12003 gnd.n4189 gnd.n4170 9.3005
R12004 gnd.n4187 gnd.n4171 9.3005
R12005 gnd.n4186 gnd.n4172 9.3005
R12006 gnd.n4184 gnd.n4173 9.3005
R12007 gnd.n4183 gnd.n4174 9.3005
R12008 gnd.n4181 gnd.n4175 9.3005
R12009 gnd.n4180 gnd.n4176 9.3005
R12010 gnd.n4178 gnd.n4177 9.3005
R12011 gnd.n2486 gnd.n2485 9.3005
R12012 gnd.n4444 gnd.n4443 9.3005
R12013 gnd.n4445 gnd.n2484 9.3005
R12014 gnd.n4459 gnd.n4446 9.3005
R12015 gnd.n4458 gnd.n4447 9.3005
R12016 gnd.n4457 gnd.n4448 9.3005
R12017 gnd.n4455 gnd.n4449 9.3005
R12018 gnd.n4454 gnd.n4450 9.3005
R12019 gnd.n4452 gnd.n4451 9.3005
R12020 gnd.n2450 gnd.n2449 9.3005
R12021 gnd.n4505 gnd.n4504 9.3005
R12022 gnd.n4506 gnd.n2448 9.3005
R12023 gnd.n4514 gnd.n4507 9.3005
R12024 gnd.n4199 gnd.n4198 9.3005
R12025 gnd.n4204 gnd.n4203 9.3005
R12026 gnd.n4207 gnd.n4160 9.3005
R12027 gnd.n4208 gnd.n4159 9.3005
R12028 gnd.n4211 gnd.n4158 9.3005
R12029 gnd.n4212 gnd.n4157 9.3005
R12030 gnd.n4215 gnd.n4156 9.3005
R12031 gnd.n4216 gnd.n4155 9.3005
R12032 gnd.n4219 gnd.n4154 9.3005
R12033 gnd.n4220 gnd.n4153 9.3005
R12034 gnd.n4223 gnd.n4152 9.3005
R12035 gnd.n4224 gnd.n4151 9.3005
R12036 gnd.n4227 gnd.n4150 9.3005
R12037 gnd.n4228 gnd.n4149 9.3005
R12038 gnd.n4231 gnd.n4148 9.3005
R12039 gnd.n4232 gnd.n4147 9.3005
R12040 gnd.n4235 gnd.n4146 9.3005
R12041 gnd.n4238 gnd.n4237 9.3005
R12042 gnd.n4202 gnd.n4164 9.3005
R12043 gnd.n4201 gnd.n4200 9.3005
R12044 gnd.n6348 gnd.n1116 9.3005
R12045 gnd.n6349 gnd.n1115 9.3005
R12046 gnd.n1114 gnd.n1111 9.3005
R12047 gnd.n6354 gnd.n1110 9.3005
R12048 gnd.n6355 gnd.n1109 9.3005
R12049 gnd.n6356 gnd.n1108 9.3005
R12050 gnd.n1107 gnd.n1104 9.3005
R12051 gnd.n6361 gnd.n1103 9.3005
R12052 gnd.n6363 gnd.n1100 9.3005
R12053 gnd.n6364 gnd.n1099 9.3005
R12054 gnd.n1098 gnd.n1095 9.3005
R12055 gnd.n6369 gnd.n1094 9.3005
R12056 gnd.n6370 gnd.n1093 9.3005
R12057 gnd.n6371 gnd.n1092 9.3005
R12058 gnd.n1091 gnd.n1088 9.3005
R12059 gnd.n6376 gnd.n1087 9.3005
R12060 gnd.n6377 gnd.n1086 9.3005
R12061 gnd.n6378 gnd.n1085 9.3005
R12062 gnd.n1084 gnd.n1081 9.3005
R12063 gnd.n6383 gnd.n1080 9.3005
R12064 gnd.n6384 gnd.n1079 9.3005
R12065 gnd.n6385 gnd.n1078 9.3005
R12066 gnd.n1077 gnd.n1074 9.3005
R12067 gnd.n1076 gnd.n1072 9.3005
R12068 gnd.n6392 gnd.n1071 9.3005
R12069 gnd.n6394 gnd.n6393 9.3005
R12070 gnd.n2227 gnd.n2226 9.3005
R12071 gnd.n2235 gnd.n2234 9.3005
R12072 gnd.n2236 gnd.n2224 9.3005
R12073 gnd.n2238 gnd.n2237 9.3005
R12074 gnd.n2222 gnd.n2221 9.3005
R12075 gnd.n2245 gnd.n2244 9.3005
R12076 gnd.n2246 gnd.n2220 9.3005
R12077 gnd.n2248 gnd.n2247 9.3005
R12078 gnd.n2218 gnd.n2215 9.3005
R12079 gnd.n2255 gnd.n2254 9.3005
R12080 gnd.n2256 gnd.n2214 9.3005
R12081 gnd.n2258 gnd.n2257 9.3005
R12082 gnd.n2212 gnd.n2211 9.3005
R12083 gnd.n2265 gnd.n2264 9.3005
R12084 gnd.n2266 gnd.n2210 9.3005
R12085 gnd.n2268 gnd.n2267 9.3005
R12086 gnd.n2208 gnd.n2207 9.3005
R12087 gnd.n2275 gnd.n2274 9.3005
R12088 gnd.n2276 gnd.n2206 9.3005
R12089 gnd.n2278 gnd.n2277 9.3005
R12090 gnd.n2204 gnd.n2203 9.3005
R12091 gnd.n2285 gnd.n2284 9.3005
R12092 gnd.n2286 gnd.n2202 9.3005
R12093 gnd.n2288 gnd.n2287 9.3005
R12094 gnd.n2200 gnd.n2199 9.3005
R12095 gnd.n2295 gnd.n2294 9.3005
R12096 gnd.n2296 gnd.n2198 9.3005
R12097 gnd.n2298 gnd.n2297 9.3005
R12098 gnd.n2196 gnd.n2193 9.3005
R12099 gnd.n2304 gnd.n2303 9.3005
R12100 gnd.n2225 gnd.n1117 9.3005
R12101 gnd.n4365 gnd.n4364 9.3005
R12102 gnd.n2562 gnd.n2558 9.3005
R12103 gnd.n2561 gnd.n2560 9.3005
R12104 gnd.n2542 gnd.n2539 9.3005
R12105 gnd.n4385 gnd.n2540 9.3005
R12106 gnd.n4384 gnd.n4381 9.3005
R12107 gnd.n4383 gnd.n4382 9.3005
R12108 gnd.n2524 gnd.n2521 9.3005
R12109 gnd.n4405 gnd.n2522 9.3005
R12110 gnd.n4404 gnd.n4401 9.3005
R12111 gnd.n4403 gnd.n4402 9.3005
R12112 gnd.n2506 gnd.n2502 9.3005
R12113 gnd.n4429 gnd.n2503 9.3005
R12114 gnd.n4428 gnd.n2504 9.3005
R12115 gnd.n4427 gnd.n4423 9.3005
R12116 gnd.n4426 gnd.n4424 9.3005
R12117 gnd.n2480 gnd.n2477 9.3005
R12118 gnd.n4470 gnd.n2478 9.3005
R12119 gnd.n4469 gnd.n4466 9.3005
R12120 gnd.n4468 gnd.n4467 9.3005
R12121 gnd.n2463 gnd.n2459 9.3005
R12122 gnd.n4495 gnd.n2460 9.3005
R12123 gnd.n4494 gnd.n2461 9.3005
R12124 gnd.n4493 gnd.n4489 9.3005
R12125 gnd.n4491 gnd.n4490 9.3005
R12126 gnd.n2447 gnd.n2442 9.3005
R12127 gnd.n4527 gnd.n2443 9.3005
R12128 gnd.n4526 gnd.n2444 9.3005
R12129 gnd.n4525 gnd.n4524 9.3005
R12130 gnd.n2445 gnd.n961 9.3005
R12131 gnd.n6462 gnd.n962 9.3005
R12132 gnd.n6461 gnd.n963 9.3005
R12133 gnd.n6460 gnd.n964 9.3005
R12134 gnd.n4577 gnd.n965 9.3005
R12135 gnd.n6450 gnd.n981 9.3005
R12136 gnd.n6449 gnd.n982 9.3005
R12137 gnd.n6448 gnd.n983 9.3005
R12138 gnd.n4592 gnd.n984 9.3005
R12139 gnd.n6438 gnd.n1001 9.3005
R12140 gnd.n6437 gnd.n1002 9.3005
R12141 gnd.n6436 gnd.n1003 9.3005
R12142 gnd.n4599 gnd.n1004 9.3005
R12143 gnd.n6426 gnd.n1021 9.3005
R12144 gnd.n6425 gnd.n1022 9.3005
R12145 gnd.n6424 gnd.n1023 9.3005
R12146 gnd.n2390 gnd.n1024 9.3005
R12147 gnd.n6414 gnd.n1041 9.3005
R12148 gnd.n6413 gnd.n1042 9.3005
R12149 gnd.n6412 gnd.n1043 9.3005
R12150 gnd.n2385 gnd.n1044 9.3005
R12151 gnd.n6402 gnd.n1061 9.3005
R12152 gnd.n6401 gnd.n1062 9.3005
R12153 gnd.n6400 gnd.n1063 9.3005
R12154 gnd.n2559 gnd.n2557 9.3005
R12155 gnd.n4364 gnd.n4363 9.3005
R12156 gnd.n4362 gnd.n2562 9.3005
R12157 gnd.n2561 gnd.n2541 9.3005
R12158 gnd.n4378 gnd.n2542 9.3005
R12159 gnd.n4379 gnd.n2540 9.3005
R12160 gnd.n4381 gnd.n4380 9.3005
R12161 gnd.n4382 gnd.n2523 9.3005
R12162 gnd.n4398 gnd.n2524 9.3005
R12163 gnd.n4399 gnd.n2522 9.3005
R12164 gnd.n4401 gnd.n4400 9.3005
R12165 gnd.n4402 gnd.n2505 9.3005
R12166 gnd.n4418 gnd.n2506 9.3005
R12167 gnd.n4419 gnd.n2503 9.3005
R12168 gnd.n4421 gnd.n2504 9.3005
R12169 gnd.n4423 gnd.n4422 9.3005
R12170 gnd.n4424 gnd.n2479 9.3005
R12171 gnd.n4463 gnd.n2480 9.3005
R12172 gnd.n4464 gnd.n2478 9.3005
R12173 gnd.n4466 gnd.n4465 9.3005
R12174 gnd.n4467 gnd.n2462 9.3005
R12175 gnd.n4484 gnd.n2463 9.3005
R12176 gnd.n4485 gnd.n2460 9.3005
R12177 gnd.n4486 gnd.n2461 9.3005
R12178 gnd.n4489 gnd.n4488 9.3005
R12179 gnd.n4490 gnd.n2446 9.3005
R12180 gnd.n4518 gnd.n2447 9.3005
R12181 gnd.n4519 gnd.n2443 9.3005
R12182 gnd.n4521 gnd.n2444 9.3005
R12183 gnd.n4524 gnd.n4523 9.3005
R12184 gnd.n4522 gnd.n2445 9.3005
R12185 gnd.n2417 gnd.n962 9.3005
R12186 gnd.n4575 gnd.n963 9.3005
R12187 gnd.n4576 gnd.n964 9.3005
R12188 gnd.n4578 gnd.n4577 9.3005
R12189 gnd.n2412 gnd.n981 9.3005
R12190 gnd.n4590 gnd.n982 9.3005
R12191 gnd.n4591 gnd.n983 9.3005
R12192 gnd.n4593 gnd.n4592 9.3005
R12193 gnd.n4594 gnd.n1001 9.3005
R12194 gnd.n4597 gnd.n1002 9.3005
R12195 gnd.n4598 gnd.n1003 9.3005
R12196 gnd.n4603 gnd.n4599 9.3005
R12197 gnd.n4604 gnd.n1021 9.3005
R12198 gnd.n4605 gnd.n1022 9.3005
R12199 gnd.n2389 gnd.n1023 9.3005
R12200 gnd.n4674 gnd.n2390 9.3005
R12201 gnd.n4675 gnd.n1041 9.3005
R12202 gnd.n4676 gnd.n1042 9.3005
R12203 gnd.n2384 gnd.n1043 9.3005
R12204 gnd.n4689 gnd.n2385 9.3005
R12205 gnd.n4690 gnd.n1061 9.3005
R12206 gnd.n4692 gnd.n1062 9.3005
R12207 gnd.n4691 gnd.n1063 9.3005
R12208 gnd.n4361 gnd.n2559 9.3005
R12209 gnd.n4242 gnd.n4241 9.3005
R12210 gnd.n4244 gnd.n4143 9.3005
R12211 gnd.n4245 gnd.n4142 9.3005
R12212 gnd.n4248 gnd.n4141 9.3005
R12213 gnd.n4249 gnd.n4140 9.3005
R12214 gnd.n4252 gnd.n4139 9.3005
R12215 gnd.n4253 gnd.n4138 9.3005
R12216 gnd.n4256 gnd.n4137 9.3005
R12217 gnd.n4257 gnd.n4136 9.3005
R12218 gnd.n4260 gnd.n4135 9.3005
R12219 gnd.n4261 gnd.n4134 9.3005
R12220 gnd.n4264 gnd.n4133 9.3005
R12221 gnd.n4265 gnd.n4132 9.3005
R12222 gnd.n4268 gnd.n4131 9.3005
R12223 gnd.n4269 gnd.n4130 9.3005
R12224 gnd.n4272 gnd.n4129 9.3005
R12225 gnd.n4273 gnd.n4128 9.3005
R12226 gnd.n4276 gnd.n4127 9.3005
R12227 gnd.n4277 gnd.n4126 9.3005
R12228 gnd.n4280 gnd.n4125 9.3005
R12229 gnd.n4284 gnd.n4121 9.3005
R12230 gnd.n4285 gnd.n4120 9.3005
R12231 gnd.n4288 gnd.n4119 9.3005
R12232 gnd.n4289 gnd.n4118 9.3005
R12233 gnd.n4292 gnd.n4117 9.3005
R12234 gnd.n4293 gnd.n4116 9.3005
R12235 gnd.n4296 gnd.n4115 9.3005
R12236 gnd.n4297 gnd.n4114 9.3005
R12237 gnd.n4300 gnd.n4113 9.3005
R12238 gnd.n4301 gnd.n4112 9.3005
R12239 gnd.n4304 gnd.n4111 9.3005
R12240 gnd.n4305 gnd.n4110 9.3005
R12241 gnd.n4308 gnd.n4109 9.3005
R12242 gnd.n4309 gnd.n4108 9.3005
R12243 gnd.n4312 gnd.n4107 9.3005
R12244 gnd.n4313 gnd.n4106 9.3005
R12245 gnd.n4316 gnd.n4105 9.3005
R12246 gnd.n4317 gnd.n4104 9.3005
R12247 gnd.n4320 gnd.n4103 9.3005
R12248 gnd.n4322 gnd.n4100 9.3005
R12249 gnd.n4325 gnd.n4099 9.3005
R12250 gnd.n4326 gnd.n4098 9.3005
R12251 gnd.n4329 gnd.n4097 9.3005
R12252 gnd.n4330 gnd.n4096 9.3005
R12253 gnd.n4333 gnd.n4095 9.3005
R12254 gnd.n4334 gnd.n4094 9.3005
R12255 gnd.n4337 gnd.n4093 9.3005
R12256 gnd.n4338 gnd.n4092 9.3005
R12257 gnd.n4341 gnd.n4091 9.3005
R12258 gnd.n4342 gnd.n4090 9.3005
R12259 gnd.n4345 gnd.n4089 9.3005
R12260 gnd.n4346 gnd.n4088 9.3005
R12261 gnd.n4349 gnd.n4087 9.3005
R12262 gnd.n4351 gnd.n4086 9.3005
R12263 gnd.n4352 gnd.n4085 9.3005
R12264 gnd.n4353 gnd.n4084 9.3005
R12265 gnd.n4354 gnd.n4083 9.3005
R12266 gnd.n4281 gnd.n4122 9.3005
R12267 gnd.n4240 gnd.n2563 9.3005
R12268 gnd.n4370 gnd.n4369 9.3005
R12269 gnd.n4371 gnd.n2548 9.3005
R12270 gnd.n4373 gnd.n4372 9.3005
R12271 gnd.n2531 gnd.n2530 9.3005
R12272 gnd.n4390 gnd.n4389 9.3005
R12273 gnd.n4391 gnd.n2529 9.3005
R12274 gnd.n4393 gnd.n4392 9.3005
R12275 gnd.n2514 gnd.n2513 9.3005
R12276 gnd.n4410 gnd.n4409 9.3005
R12277 gnd.n4411 gnd.n2512 9.3005
R12278 gnd.n4413 gnd.n4412 9.3005
R12279 gnd.n2494 gnd.n2493 9.3005
R12280 gnd.n4434 gnd.n4433 9.3005
R12281 gnd.n4435 gnd.n2492 9.3005
R12282 gnd.n4439 gnd.n4436 9.3005
R12283 gnd.n4438 gnd.n4437 9.3005
R12284 gnd.n2470 gnd.n2469 9.3005
R12285 gnd.n4475 gnd.n4474 9.3005
R12286 gnd.n4476 gnd.n2468 9.3005
R12287 gnd.n4479 gnd.n4477 9.3005
R12288 gnd.n4478 gnd.n947 9.3005
R12289 gnd.n953 gnd.n946 9.3005
R12290 gnd.n6456 gnd.n971 9.3005
R12291 gnd.n6455 gnd.n972 9.3005
R12292 gnd.n6454 gnd.n973 9.3005
R12293 gnd.n991 gnd.n974 9.3005
R12294 gnd.n6444 gnd.n992 9.3005
R12295 gnd.n6443 gnd.n993 9.3005
R12296 gnd.n6442 gnd.n994 9.3005
R12297 gnd.n1010 gnd.n995 9.3005
R12298 gnd.n6432 gnd.n1011 9.3005
R12299 gnd.n6431 gnd.n1012 9.3005
R12300 gnd.n6430 gnd.n1013 9.3005
R12301 gnd.n1031 gnd.n1014 9.3005
R12302 gnd.n6420 gnd.n1032 9.3005
R12303 gnd.n6419 gnd.n1033 9.3005
R12304 gnd.n6418 gnd.n1034 9.3005
R12305 gnd.n1051 gnd.n1035 9.3005
R12306 gnd.n6408 gnd.n1052 9.3005
R12307 gnd.n6407 gnd.n1053 9.3005
R12308 gnd.n6406 gnd.n1054 9.3005
R12309 gnd.n1070 gnd.n1055 9.3005
R12310 gnd.n6396 gnd.n6395 9.3005
R12311 gnd.n2550 gnd.n2549 9.3005
R12312 gnd.n6467 gnd.n944 9.3005
R12313 gnd.n6467 gnd.n6466 9.3005
R12314 gnd.n2430 gnd.n2429 9.3005
R12315 gnd.n4539 gnd.n4538 9.3005
R12316 gnd.n4540 gnd.n2426 9.3005
R12317 gnd.n4562 gnd.n4541 9.3005
R12318 gnd.n4561 gnd.n4542 9.3005
R12319 gnd.n2428 gnd.n2427 9.3005
R12320 gnd.n6475 gnd.n935 9.3005
R12321 gnd.n6476 gnd.n934 9.3005
R12322 gnd.n933 gnd.n929 9.3005
R12323 gnd.n6482 gnd.n928 9.3005
R12324 gnd.n6483 gnd.n927 9.3005
R12325 gnd.n6484 gnd.n926 9.3005
R12326 gnd.n925 gnd.n921 9.3005
R12327 gnd.n6490 gnd.n920 9.3005
R12328 gnd.n6491 gnd.n919 9.3005
R12329 gnd.n6492 gnd.n918 9.3005
R12330 gnd.n917 gnd.n913 9.3005
R12331 gnd.n6498 gnd.n912 9.3005
R12332 gnd.n6499 gnd.n911 9.3005
R12333 gnd.n6500 gnd.n910 9.3005
R12334 gnd.n909 gnd.n905 9.3005
R12335 gnd.n6506 gnd.n904 9.3005
R12336 gnd.n6507 gnd.n903 9.3005
R12337 gnd.n6508 gnd.n902 9.3005
R12338 gnd.n901 gnd.n897 9.3005
R12339 gnd.n6514 gnd.n896 9.3005
R12340 gnd.n6515 gnd.n895 9.3005
R12341 gnd.n6516 gnd.n894 9.3005
R12342 gnd.n893 gnd.n889 9.3005
R12343 gnd.n6522 gnd.n888 9.3005
R12344 gnd.n6523 gnd.n887 9.3005
R12345 gnd.n6524 gnd.n886 9.3005
R12346 gnd.n885 gnd.n881 9.3005
R12347 gnd.n6530 gnd.n880 9.3005
R12348 gnd.n6531 gnd.n879 9.3005
R12349 gnd.n6532 gnd.n878 9.3005
R12350 gnd.n877 gnd.n873 9.3005
R12351 gnd.n6538 gnd.n872 9.3005
R12352 gnd.n6539 gnd.n871 9.3005
R12353 gnd.n6540 gnd.n870 9.3005
R12354 gnd.n869 gnd.n865 9.3005
R12355 gnd.n6546 gnd.n864 9.3005
R12356 gnd.n6547 gnd.n863 9.3005
R12357 gnd.n6548 gnd.n862 9.3005
R12358 gnd.n861 gnd.n857 9.3005
R12359 gnd.n6554 gnd.n856 9.3005
R12360 gnd.n6555 gnd.n855 9.3005
R12361 gnd.n6556 gnd.n854 9.3005
R12362 gnd.n853 gnd.n849 9.3005
R12363 gnd.n6562 gnd.n848 9.3005
R12364 gnd.n6563 gnd.n847 9.3005
R12365 gnd.n6564 gnd.n846 9.3005
R12366 gnd.n845 gnd.n841 9.3005
R12367 gnd.n6570 gnd.n840 9.3005
R12368 gnd.n6571 gnd.n839 9.3005
R12369 gnd.n6572 gnd.n838 9.3005
R12370 gnd.n837 gnd.n833 9.3005
R12371 gnd.n6578 gnd.n832 9.3005
R12372 gnd.n6579 gnd.n831 9.3005
R12373 gnd.n6580 gnd.n830 9.3005
R12374 gnd.n829 gnd.n825 9.3005
R12375 gnd.n6586 gnd.n824 9.3005
R12376 gnd.n6587 gnd.n823 9.3005
R12377 gnd.n6588 gnd.n822 9.3005
R12378 gnd.n821 gnd.n817 9.3005
R12379 gnd.n6594 gnd.n816 9.3005
R12380 gnd.n6595 gnd.n815 9.3005
R12381 gnd.n6596 gnd.n814 9.3005
R12382 gnd.n813 gnd.n809 9.3005
R12383 gnd.n6602 gnd.n808 9.3005
R12384 gnd.n6603 gnd.n807 9.3005
R12385 gnd.n6604 gnd.n806 9.3005
R12386 gnd.n805 gnd.n801 9.3005
R12387 gnd.n6610 gnd.n800 9.3005
R12388 gnd.n6611 gnd.n799 9.3005
R12389 gnd.n6612 gnd.n798 9.3005
R12390 gnd.n797 gnd.n793 9.3005
R12391 gnd.n6618 gnd.n792 9.3005
R12392 gnd.n6619 gnd.n791 9.3005
R12393 gnd.n6620 gnd.n790 9.3005
R12394 gnd.n789 gnd.n785 9.3005
R12395 gnd.n6626 gnd.n784 9.3005
R12396 gnd.n6627 gnd.n783 9.3005
R12397 gnd.n6628 gnd.n782 9.3005
R12398 gnd.n781 gnd.n777 9.3005
R12399 gnd.n6634 gnd.n776 9.3005
R12400 gnd.n6635 gnd.n775 9.3005
R12401 gnd.n6636 gnd.n774 9.3005
R12402 gnd.n770 gnd.n769 9.3005
R12403 gnd.n6643 gnd.n6642 9.3005
R12404 gnd.n6474 gnd.n936 9.3005
R12405 gnd.n5731 gnd.n1635 9.3005
R12406 gnd.n4786 gnd.n2109 9.3005
R12407 gnd.n4788 gnd.n4787 9.3005
R12408 gnd.n2098 gnd.n2097 9.3005
R12409 gnd.n4801 gnd.n4800 9.3005
R12410 gnd.n4802 gnd.n2096 9.3005
R12411 gnd.n4804 gnd.n4803 9.3005
R12412 gnd.n2084 gnd.n2083 9.3005
R12413 gnd.n4817 gnd.n4816 9.3005
R12414 gnd.n4818 gnd.n2082 9.3005
R12415 gnd.n4820 gnd.n4819 9.3005
R12416 gnd.n2070 gnd.n2069 9.3005
R12417 gnd.n4833 gnd.n4832 9.3005
R12418 gnd.n4834 gnd.n2068 9.3005
R12419 gnd.n4836 gnd.n4835 9.3005
R12420 gnd.n2056 gnd.n2055 9.3005
R12421 gnd.n4849 gnd.n4848 9.3005
R12422 gnd.n4850 gnd.n2053 9.3005
R12423 gnd.n4866 gnd.n4865 9.3005
R12424 gnd.n4864 gnd.n2054 9.3005
R12425 gnd.n4863 gnd.n4862 9.3005
R12426 gnd.n4861 gnd.n4851 9.3005
R12427 gnd.n4860 gnd.n4859 9.3005
R12428 gnd.n4858 gnd.n4855 9.3005
R12429 gnd.n4857 gnd.n4856 9.3005
R12430 gnd.n1200 gnd.n1198 9.3005
R12431 gnd.n6264 gnd.n6263 9.3005
R12432 gnd.n6262 gnd.n1199 9.3005
R12433 gnd.n6261 gnd.n6260 9.3005
R12434 gnd.n6259 gnd.n1201 9.3005
R12435 gnd.n6258 gnd.n6257 9.3005
R12436 gnd.n6256 gnd.n1205 9.3005
R12437 gnd.n6255 gnd.n6254 9.3005
R12438 gnd.n6253 gnd.n1206 9.3005
R12439 gnd.n6252 gnd.n6251 9.3005
R12440 gnd.n6250 gnd.n1210 9.3005
R12441 gnd.n6249 gnd.n6248 9.3005
R12442 gnd.n6247 gnd.n1211 9.3005
R12443 gnd.n6246 gnd.n6245 9.3005
R12444 gnd.n6244 gnd.n1215 9.3005
R12445 gnd.n6243 gnd.n6242 9.3005
R12446 gnd.n6241 gnd.n1216 9.3005
R12447 gnd.n6240 gnd.n6239 9.3005
R12448 gnd.n6238 gnd.n1220 9.3005
R12449 gnd.n6237 gnd.n6236 9.3005
R12450 gnd.n6235 gnd.n1221 9.3005
R12451 gnd.n6234 gnd.n6233 9.3005
R12452 gnd.n6232 gnd.n1225 9.3005
R12453 gnd.n6231 gnd.n6230 9.3005
R12454 gnd.n6229 gnd.n1226 9.3005
R12455 gnd.n6228 gnd.n6227 9.3005
R12456 gnd.n6226 gnd.n1230 9.3005
R12457 gnd.n6225 gnd.n6224 9.3005
R12458 gnd.n6223 gnd.n1231 9.3005
R12459 gnd.n6222 gnd.n6221 9.3005
R12460 gnd.n6220 gnd.n1235 9.3005
R12461 gnd.n6219 gnd.n6218 9.3005
R12462 gnd.n6217 gnd.n1236 9.3005
R12463 gnd.n6216 gnd.n6215 9.3005
R12464 gnd.n6214 gnd.n1240 9.3005
R12465 gnd.n6213 gnd.n6212 9.3005
R12466 gnd.n6211 gnd.n1241 9.3005
R12467 gnd.n6210 gnd.n6209 9.3005
R12468 gnd.n6208 gnd.n1245 9.3005
R12469 gnd.n6207 gnd.n6206 9.3005
R12470 gnd.n6205 gnd.n1246 9.3005
R12471 gnd.n6204 gnd.n6203 9.3005
R12472 gnd.n6202 gnd.n1250 9.3005
R12473 gnd.n6201 gnd.n6200 9.3005
R12474 gnd.n6199 gnd.n1251 9.3005
R12475 gnd.n6198 gnd.n6197 9.3005
R12476 gnd.n6196 gnd.n1255 9.3005
R12477 gnd.n6195 gnd.n6194 9.3005
R12478 gnd.n6193 gnd.n1256 9.3005
R12479 gnd.n6192 gnd.n6191 9.3005
R12480 gnd.n6190 gnd.n1260 9.3005
R12481 gnd.n6189 gnd.n6188 9.3005
R12482 gnd.n6187 gnd.n1261 9.3005
R12483 gnd.n6186 gnd.n6185 9.3005
R12484 gnd.n6184 gnd.n1265 9.3005
R12485 gnd.n6183 gnd.n6182 9.3005
R12486 gnd.n6181 gnd.n1266 9.3005
R12487 gnd.n6180 gnd.n6179 9.3005
R12488 gnd.n6178 gnd.n1270 9.3005
R12489 gnd.n6177 gnd.n6176 9.3005
R12490 gnd.n6175 gnd.n1271 9.3005
R12491 gnd.n6174 gnd.n6173 9.3005
R12492 gnd.n6172 gnd.n1275 9.3005
R12493 gnd.n6171 gnd.n6170 9.3005
R12494 gnd.n6169 gnd.n1276 9.3005
R12495 gnd.n6168 gnd.n6167 9.3005
R12496 gnd.n6166 gnd.n1280 9.3005
R12497 gnd.n6165 gnd.n6164 9.3005
R12498 gnd.n6163 gnd.n1281 9.3005
R12499 gnd.n6162 gnd.n6161 9.3005
R12500 gnd.n6160 gnd.n1285 9.3005
R12501 gnd.n6159 gnd.n6158 9.3005
R12502 gnd.n6157 gnd.n1286 9.3005
R12503 gnd.n6156 gnd.n6155 9.3005
R12504 gnd.n6154 gnd.n1290 9.3005
R12505 gnd.n6153 gnd.n6152 9.3005
R12506 gnd.n6151 gnd.n1291 9.3005
R12507 gnd.n4785 gnd.n4784 9.3005
R12508 gnd.n4705 gnd.n2110 9.3005
R12509 gnd.n4513 gnd.n4512 9.3005
R12510 gnd.n4511 gnd.n4509 9.3005
R12511 gnd.n2420 gnd.n2419 9.3005
R12512 gnd.n4568 gnd.n4567 9.3005
R12513 gnd.n4569 gnd.n2418 9.3005
R12514 gnd.n4571 gnd.n4570 9.3005
R12515 gnd.n2415 gnd.n2414 9.3005
R12516 gnd.n4583 gnd.n4582 9.3005
R12517 gnd.n4584 gnd.n2413 9.3005
R12518 gnd.n4586 gnd.n4585 9.3005
R12519 gnd.n2406 gnd.n2404 9.3005
R12520 gnd.n4622 gnd.n4621 9.3005
R12521 gnd.n4620 gnd.n2405 9.3005
R12522 gnd.n4619 gnd.n4618 9.3005
R12523 gnd.n4617 gnd.n2407 9.3005
R12524 gnd.n4616 gnd.n4615 9.3005
R12525 gnd.n4614 gnd.n2410 9.3005
R12526 gnd.n4613 gnd.n4612 9.3005
R12527 gnd.n4611 gnd.n2411 9.3005
R12528 gnd.n4610 gnd.n4609 9.3005
R12529 gnd.n2388 gnd.n2387 9.3005
R12530 gnd.n4681 gnd.n4680 9.3005
R12531 gnd.n4682 gnd.n2386 9.3005
R12532 gnd.n4685 gnd.n4684 9.3005
R12533 gnd.n4683 gnd.n2382 9.3005
R12534 gnd.n4696 gnd.n2381 9.3005
R12535 gnd.n4698 gnd.n4697 9.3005
R12536 gnd.n4754 gnd.n4753 9.3005
R12537 gnd.n4752 gnd.n4751 9.3005
R12538 gnd.n2319 gnd.n2318 9.3005
R12539 gnd.n4746 gnd.n4745 9.3005
R12540 gnd.n4744 gnd.n4743 9.3005
R12541 gnd.n2331 gnd.n2330 9.3005
R12542 gnd.n4738 gnd.n4737 9.3005
R12543 gnd.n4736 gnd.n4735 9.3005
R12544 gnd.n2342 gnd.n2341 9.3005
R12545 gnd.n4730 gnd.n4729 9.3005
R12546 gnd.n4728 gnd.n4727 9.3005
R12547 gnd.n2354 gnd.n2353 9.3005
R12548 gnd.n4722 gnd.n4721 9.3005
R12549 gnd.n4720 gnd.n4719 9.3005
R12550 gnd.n2365 gnd.n2364 9.3005
R12551 gnd.n4714 gnd.n4713 9.3005
R12552 gnd.n4712 gnd.n2378 9.3005
R12553 gnd.n4711 gnd.n4708 9.3005
R12554 gnd.n2314 gnd.n2312 9.3005
R12555 gnd.n4707 gnd.n4706 9.3005
R12556 gnd.n4702 gnd.n2380 9.3005
R12557 gnd.n4701 gnd.n2372 9.3005
R12558 gnd.n4716 gnd.n4715 9.3005
R12559 gnd.n4718 gnd.n4717 9.3005
R12560 gnd.n2358 gnd.n2357 9.3005
R12561 gnd.n4724 gnd.n4723 9.3005
R12562 gnd.n4726 gnd.n4725 9.3005
R12563 gnd.n2348 gnd.n2347 9.3005
R12564 gnd.n4732 gnd.n4731 9.3005
R12565 gnd.n4734 gnd.n4733 9.3005
R12566 gnd.n2335 gnd.n2334 9.3005
R12567 gnd.n4740 gnd.n4739 9.3005
R12568 gnd.n4742 gnd.n4741 9.3005
R12569 gnd.n2325 gnd.n2324 9.3005
R12570 gnd.n4748 gnd.n4747 9.3005
R12571 gnd.n4750 gnd.n4749 9.3005
R12572 gnd.n2313 gnd.n2311 9.3005
R12573 gnd.n4756 gnd.n4755 9.3005
R12574 gnd.n4757 gnd.n2306 9.3005
R12575 gnd.n4759 gnd.n4758 9.3005
R12576 gnd.n4761 gnd.n2192 9.3005
R12577 gnd.n4763 gnd.n4762 9.3005
R12578 gnd.n4764 gnd.n2188 9.3005
R12579 gnd.n4766 gnd.n4765 9.3005
R12580 gnd.n4767 gnd.n2187 9.3005
R12581 gnd.n4769 gnd.n4768 9.3005
R12582 gnd.n4770 gnd.n2186 9.3005
R12583 gnd.n2183 gnd.n2136 9.3005
R12584 gnd.n2182 gnd.n2181 9.3005
R12585 gnd.n2180 gnd.n2139 9.3005
R12586 gnd.n2179 gnd.n2178 9.3005
R12587 gnd.n2177 gnd.n2140 9.3005
R12588 gnd.n2176 gnd.n2175 9.3005
R12589 gnd.n2174 gnd.n2143 9.3005
R12590 gnd.n2173 gnd.n2172 9.3005
R12591 gnd.n2171 gnd.n2144 9.3005
R12592 gnd.n2170 gnd.n2169 9.3005
R12593 gnd.n2168 gnd.n2147 9.3005
R12594 gnd.n2167 gnd.n2166 9.3005
R12595 gnd.n2165 gnd.n2148 9.3005
R12596 gnd.n2164 gnd.n2163 9.3005
R12597 gnd.n2162 gnd.n2151 9.3005
R12598 gnd.n2161 gnd.n2160 9.3005
R12599 gnd.n2159 gnd.n2152 9.3005
R12600 gnd.n2158 gnd.n2157 9.3005
R12601 gnd.n2156 gnd.n2154 9.3005
R12602 gnd.n2155 gnd.n2040 9.3005
R12603 gnd.n2038 gnd.n2037 9.3005
R12604 gnd.n4888 gnd.n4887 9.3005
R12605 gnd.n4889 gnd.n2036 9.3005
R12606 gnd.n4891 gnd.n4890 9.3005
R12607 gnd.n4992 gnd.n2035 9.3005
R12608 gnd.n4994 gnd.n4993 9.3005
R12609 gnd.n4995 gnd.n2033 9.3005
R12610 gnd.n5024 gnd.n5023 9.3005
R12611 gnd.n5022 gnd.n2034 9.3005
R12612 gnd.n5021 gnd.n5020 9.3005
R12613 gnd.n5019 gnd.n4996 9.3005
R12614 gnd.n5018 gnd.n5017 9.3005
R12615 gnd.n5016 gnd.n4998 9.3005
R12616 gnd.n5015 gnd.n5014 9.3005
R12617 gnd.n5013 gnd.n4999 9.3005
R12618 gnd.n5012 gnd.n5011 9.3005
R12619 gnd.n5010 gnd.n5003 9.3005
R12620 gnd.n5009 gnd.n5008 9.3005
R12621 gnd.n5007 gnd.n5005 9.3005
R12622 gnd.n5004 gnd.n1971 9.3005
R12623 gnd.n5129 gnd.n1970 9.3005
R12624 gnd.n5131 gnd.n5130 9.3005
R12625 gnd.n5132 gnd.n1968 9.3005
R12626 gnd.n5160 gnd.n5159 9.3005
R12627 gnd.n5158 gnd.n1969 9.3005
R12628 gnd.n5157 gnd.n5156 9.3005
R12629 gnd.n5155 gnd.n5133 9.3005
R12630 gnd.n5154 gnd.n5153 9.3005
R12631 gnd.n5152 gnd.n5135 9.3005
R12632 gnd.n5151 gnd.n5150 9.3005
R12633 gnd.n5149 gnd.n5136 9.3005
R12634 gnd.n5148 gnd.n5147 9.3005
R12635 gnd.n5146 gnd.n5140 9.3005
R12636 gnd.n5145 gnd.n5144 9.3005
R12637 gnd.n5143 gnd.n5141 9.3005
R12638 gnd.n1878 gnd.n1877 9.3005
R12639 gnd.n5282 gnd.n5281 9.3005
R12640 gnd.n5283 gnd.n1875 9.3005
R12641 gnd.n5286 gnd.n5285 9.3005
R12642 gnd.n5284 gnd.n1876 9.3005
R12643 gnd.n1851 gnd.n1850 9.3005
R12644 gnd.n5331 gnd.n5330 9.3005
R12645 gnd.n5332 gnd.n1848 9.3005
R12646 gnd.n5350 gnd.n5349 9.3005
R12647 gnd.n5348 gnd.n1849 9.3005
R12648 gnd.n5347 gnd.n5346 9.3005
R12649 gnd.n5345 gnd.n5333 9.3005
R12650 gnd.n5344 gnd.n5343 9.3005
R12651 gnd.n5342 gnd.n5337 9.3005
R12652 gnd.n5341 gnd.n5340 9.3005
R12653 gnd.n5339 gnd.n5338 9.3005
R12654 gnd.n1799 gnd.n1798 9.3005
R12655 gnd.n5411 gnd.n5410 9.3005
R12656 gnd.n5412 gnd.n1796 9.3005
R12657 gnd.n5424 gnd.n5423 9.3005
R12658 gnd.n5422 gnd.n1797 9.3005
R12659 gnd.n5421 gnd.n5420 9.3005
R12660 gnd.n5419 gnd.n5413 9.3005
R12661 gnd.n5418 gnd.n5417 9.3005
R12662 gnd.n1721 gnd.n1720 9.3005
R12663 gnd.n5629 gnd.n5628 9.3005
R12664 gnd.n5630 gnd.n1719 9.3005
R12665 gnd.n5632 gnd.n5631 9.3005
R12666 gnd.n1709 gnd.n1708 9.3005
R12667 gnd.n5646 gnd.n5645 9.3005
R12668 gnd.n5647 gnd.n1707 9.3005
R12669 gnd.n5649 gnd.n5648 9.3005
R12670 gnd.n1697 gnd.n1696 9.3005
R12671 gnd.n5663 gnd.n5662 9.3005
R12672 gnd.n5664 gnd.n1695 9.3005
R12673 gnd.n5666 gnd.n5665 9.3005
R12674 gnd.n1684 gnd.n1683 9.3005
R12675 gnd.n5680 gnd.n5679 9.3005
R12676 gnd.n5681 gnd.n1682 9.3005
R12677 gnd.n5683 gnd.n5682 9.3005
R12678 gnd.n1673 gnd.n1672 9.3005
R12679 gnd.n5700 gnd.n5699 9.3005
R12680 gnd.n5701 gnd.n1671 9.3005
R12681 gnd.n5703 gnd.n5702 9.3005
R12682 gnd.n1300 gnd.n1299 9.3005
R12683 gnd.n6147 gnd.n6146 9.3005
R12684 gnd.n2185 gnd.n2184 9.3005
R12685 gnd.n6143 gnd.n1301 9.3005
R12686 gnd.n6142 gnd.n6141 9.3005
R12687 gnd.n6140 gnd.n1304 9.3005
R12688 gnd.n6139 gnd.n6138 9.3005
R12689 gnd.n6137 gnd.n1305 9.3005
R12690 gnd.n6136 gnd.n6135 9.3005
R12691 gnd.n6145 gnd.n6144 9.3005
R12692 gnd.n6088 gnd.n6087 9.3005
R12693 gnd.n1352 gnd.n1351 9.3005
R12694 gnd.n6094 gnd.n6093 9.3005
R12695 gnd.n6096 gnd.n6095 9.3005
R12696 gnd.n1344 gnd.n1343 9.3005
R12697 gnd.n6102 gnd.n6101 9.3005
R12698 gnd.n6104 gnd.n6103 9.3005
R12699 gnd.n1336 gnd.n1335 9.3005
R12700 gnd.n6110 gnd.n6109 9.3005
R12701 gnd.n6112 gnd.n6111 9.3005
R12702 gnd.n1328 gnd.n1327 9.3005
R12703 gnd.n6118 gnd.n6117 9.3005
R12704 gnd.n6120 gnd.n6119 9.3005
R12705 gnd.n1320 gnd.n1319 9.3005
R12706 gnd.n6126 gnd.n6125 9.3005
R12707 gnd.n6128 gnd.n6127 9.3005
R12708 gnd.n1316 gnd.n1311 9.3005
R12709 gnd.n6086 gnd.n1361 9.3005
R12710 gnd.n1636 gnd.n1360 9.3005
R12711 gnd.n6133 gnd.n1309 9.3005
R12712 gnd.n6132 gnd.n6131 9.3005
R12713 gnd.n6130 gnd.n6129 9.3005
R12714 gnd.n1315 gnd.n1314 9.3005
R12715 gnd.n6124 gnd.n6123 9.3005
R12716 gnd.n6122 gnd.n6121 9.3005
R12717 gnd.n1324 gnd.n1323 9.3005
R12718 gnd.n6116 gnd.n6115 9.3005
R12719 gnd.n6114 gnd.n6113 9.3005
R12720 gnd.n1332 gnd.n1331 9.3005
R12721 gnd.n6108 gnd.n6107 9.3005
R12722 gnd.n6106 gnd.n6105 9.3005
R12723 gnd.n1340 gnd.n1339 9.3005
R12724 gnd.n6100 gnd.n6099 9.3005
R12725 gnd.n6098 gnd.n6097 9.3005
R12726 gnd.n1348 gnd.n1347 9.3005
R12727 gnd.n6092 gnd.n6091 9.3005
R12728 gnd.n6090 gnd.n6089 9.3005
R12729 gnd.n1659 gnd.n1358 9.3005
R12730 gnd.n1638 gnd.n1637 9.3005
R12731 gnd.n5733 gnd.n5732 9.3005
R12732 gnd.n5774 gnd.n5773 9.3005
R12733 gnd.n5772 gnd.n1634 9.3005
R12734 gnd.n5771 gnd.n5770 9.3005
R12735 gnd.n5769 gnd.n5736 9.3005
R12736 gnd.n5768 gnd.n5767 9.3005
R12737 gnd.n5766 gnd.n5740 9.3005
R12738 gnd.n5765 gnd.n5764 9.3005
R12739 gnd.n5763 gnd.n5741 9.3005
R12740 gnd.n5762 gnd.n5761 9.3005
R12741 gnd.n1617 gnd.n1616 9.3005
R12742 gnd.n5825 gnd.n5824 9.3005
R12743 gnd.n5826 gnd.n1615 9.3005
R12744 gnd.n5828 gnd.n5827 9.3005
R12745 gnd.n1612 gnd.n1611 9.3005
R12746 gnd.n5840 gnd.n5839 9.3005
R12747 gnd.n5841 gnd.n1610 9.3005
R12748 gnd.n5843 gnd.n5842 9.3005
R12749 gnd.n1607 gnd.n1605 9.3005
R12750 gnd.n5873 gnd.n5872 9.3005
R12751 gnd.n5871 gnd.n1606 9.3005
R12752 gnd.n5870 gnd.n5869 9.3005
R12753 gnd.n5868 gnd.n1608 9.3005
R12754 gnd.n5867 gnd.n5866 9.3005
R12755 gnd.n5865 gnd.n5862 9.3005
R12756 gnd.n5864 gnd.n5863 9.3005
R12757 gnd.n85 gnd.n83 9.3005
R12758 gnd.n5735 gnd.n1633 9.3005
R12759 gnd.t0 gnd.n2755 9.24152
R12760 gnd.n2657 gnd.t170 9.24152
R12761 gnd.n3942 gnd.t145 9.24152
R12762 gnd.t81 gnd.n2544 9.24152
R12763 gnd.n4600 gnd.t285 9.24152
R12764 gnd.n6404 gnd.t113 9.24152
R12765 gnd.n5952 gnd.t77 9.24152
R12766 gnd.n5821 gnd.t232 9.24152
R12767 gnd.n7543 gnd.t95 9.24152
R12768 gnd.t25 gnd.t0 8.92286
R12769 gnd.n5026 gnd.n2031 8.92286
R12770 gnd.n5120 gnd.n1979 8.92286
R12771 gnd.n5187 gnd.n5186 8.92286
R12772 gnd.n5194 gnd.t21 8.92286
R12773 gnd.n5269 gnd.t22 8.92286
R12774 gnd.n5252 gnd.n1890 8.92286
R12775 gnd.n5328 gnd.n1853 8.92286
R12776 gnd.n5435 gnd.n1790 8.92286
R12777 gnd.n3912 gnd.n3887 8.92171
R12778 gnd.n3880 gnd.n3855 8.92171
R12779 gnd.n3848 gnd.n3823 8.92171
R12780 gnd.n3817 gnd.n3792 8.92171
R12781 gnd.n3785 gnd.n3760 8.92171
R12782 gnd.n3753 gnd.n3728 8.92171
R12783 gnd.n3721 gnd.n3696 8.92171
R12784 gnd.n3690 gnd.n3665 8.92171
R12785 gnd.n5474 gnd.n5456 8.72777
R12786 gnd.n3415 gnd.t9 8.60421
R12787 gnd.n2416 gnd.t210 8.60421
R12788 gnd.n5876 gnd.t261 8.60421
R12789 gnd.n191 gnd.n184 8.60421
R12790 gnd.n2827 gnd.n2811 8.43656
R12791 gnd.n50 gnd.n34 8.43656
R12792 gnd.n6272 gnd.t139 8.28555
R12793 gnd.n2012 gnd.t8 8.28555
R12794 gnd.n5108 gnd.t15 8.28555
R12795 gnd.n1966 gnd.t66 8.28555
R12796 gnd.t5 gnd.n5259 8.28555
R12797 gnd.n5310 gnd.t42 8.28555
R12798 gnd.n5376 gnd.t13 8.28555
R12799 gnd.n3913 gnd.n3885 8.14595
R12800 gnd.n3881 gnd.n3853 8.14595
R12801 gnd.n3849 gnd.n3821 8.14595
R12802 gnd.n3818 gnd.n3790 8.14595
R12803 gnd.n3786 gnd.n3758 8.14595
R12804 gnd.n3754 gnd.n3726 8.14595
R12805 gnd.n3722 gnd.n3694 8.14595
R12806 gnd.n3691 gnd.n3663 8.14595
R12807 gnd.n4510 gnd.n0 8.10675
R12808 gnd.n7617 gnd.n7616 8.10675
R12809 gnd.n3918 gnd.n3917 7.97301
R12810 gnd.t2 gnd.n2930 7.9669
R12811 gnd.n3656 gnd.n2654 7.9669
R12812 gnd.n4774 gnd.n4773 7.9669
R12813 gnd.n5728 gnd.n5727 7.9669
R12814 gnd.n7617 gnd.n82 7.86902
R12815 gnd.n6086 gnd.n1360 7.75808
R12816 gnd.n4712 gnd.n4711 7.75808
R12817 gnd.n7393 gnd.n349 7.75808
R12818 gnd.n4200 gnd.n4164 7.75808
R12819 gnd.n4971 gnd.t99 7.64824
R12820 gnd.n5047 gnd.n5046 7.64824
R12821 gnd.n5076 gnd.n1993 7.64824
R12822 gnd.n1943 gnd.n1931 7.64824
R12823 gnd.n5247 gnd.n1901 7.64824
R12824 gnd.n5353 gnd.n5352 7.64824
R12825 gnd.n5382 gnd.n1812 7.64824
R12826 gnd.n2860 gnd.n2859 7.53171
R12827 gnd.n3324 gnd.t34 7.32958
R12828 gnd.n4790 gnd.t117 7.32958
R12829 gnd.n2080 gnd.t360 7.32958
R12830 gnd.t49 gnd.n1693 7.32958
R12831 gnd.n5706 gnd.t91 7.32958
R12832 gnd.n1179 gnd.n1178 7.30353
R12833 gnd.n5473 gnd.n5472 7.30353
R12834 gnd.n3284 gnd.n3003 7.01093
R12835 gnd.n3006 gnd.n3004 7.01093
R12836 gnd.n3294 gnd.n3293 7.01093
R12837 gnd.n3305 gnd.n2987 7.01093
R12838 gnd.n3304 gnd.n2990 7.01093
R12839 gnd.n3315 gnd.n2978 7.01093
R12840 gnd.n2981 gnd.n2979 7.01093
R12841 gnd.n3325 gnd.n3324 7.01093
R12842 gnd.n3335 gnd.n2959 7.01093
R12843 gnd.n3334 gnd.n2962 7.01093
R12844 gnd.n3343 gnd.n2953 7.01093
R12845 gnd.n3355 gnd.n2943 7.01093
R12846 gnd.n3365 gnd.n2928 7.01093
R12847 gnd.n3381 gnd.n3380 7.01093
R12848 gnd.n2930 gnd.n2867 7.01093
R12849 gnd.n3435 gnd.n2868 7.01093
R12850 gnd.n3429 gnd.n3428 7.01093
R12851 gnd.n2917 gnd.n2879 7.01093
R12852 gnd.n3421 gnd.n2890 7.01093
R12853 gnd.n2908 gnd.n2903 7.01093
R12854 gnd.n3415 gnd.n3414 7.01093
R12855 gnd.n3461 gnd.n2790 7.01093
R12856 gnd.n3460 gnd.n3459 7.01093
R12857 gnd.n3472 gnd.n3471 7.01093
R12858 gnd.n2783 gnd.n2775 7.01093
R12859 gnd.n3501 gnd.n2763 7.01093
R12860 gnd.n3500 gnd.n2766 7.01093
R12861 gnd.n3511 gnd.n2755 7.01093
R12862 gnd.n2756 gnd.n2744 7.01093
R12863 gnd.n3522 gnd.n2745 7.01093
R12864 gnd.n3546 gnd.n2736 7.01093
R12865 gnd.n3545 gnd.n2727 7.01093
R12866 gnd.n3568 gnd.n3567 7.01093
R12867 gnd.n3586 gnd.n2708 7.01093
R12868 gnd.n3585 gnd.n2711 7.01093
R12869 gnd.n3596 gnd.n2700 7.01093
R12870 gnd.n2701 gnd.n2688 7.01093
R12871 gnd.n3607 gnd.n2689 7.01093
R12872 gnd.n3634 gnd.n2673 7.01093
R12873 gnd.n3646 gnd.n3645 7.01093
R12874 gnd.n3628 gnd.n2666 7.01093
R12875 gnd.n3658 gnd.n3657 7.01093
R12876 gnd.n3930 gnd.n2654 7.01093
R12877 gnd.n3929 gnd.n2657 7.01093
R12878 gnd.n3942 gnd.n2646 7.01093
R12879 gnd.n2647 gnd.n2639 7.01093
R12880 gnd.n3952 gnd.n2565 7.01093
R12881 gnd.n5452 gnd.t136 7.01093
R12882 gnd.n2962 gnd.t36 6.69227
R12883 gnd.n2766 gnd.t25 6.69227
R12884 gnd.n3635 gnd.t3 6.69227
R12885 gnd.n4407 gnd.t228 6.69227
R12886 gnd.n4607 gnd.t271 6.69227
R12887 gnd.n5174 gnd.t11 6.69227
R12888 gnd.n5260 gnd.t47 6.69227
R12889 gnd.n5759 gnd.t219 6.69227
R12890 gnd.n171 gnd.t212 6.69227
R12891 gnd.n5609 gnd.n5608 6.5566
R12892 gnd.n4902 gnd.n4901 6.5566
R12893 gnd.n6284 gnd.n6280 6.5566
R12894 gnd.n5484 gnd.n5483 6.5566
R12895 gnd.n2021 gnd.n2009 6.37362
R12896 gnd.n5083 gnd.n1999 6.37362
R12897 gnd.n5127 gnd.t71 6.37362
R12898 gnd.n5211 gnd.n1926 6.37362
R12899 gnd.n5217 gnd.n1916 6.37362
R12900 gnd.n5318 gnd.t51 6.37362
R12901 gnd.n1841 gnd.n1827 6.37362
R12902 gnd.n5389 gnd.n1817 6.37362
R12903 gnd.n4701 gnd.n2371 6.20656
R12904 gnd.n1659 gnd.n1357 6.20656
R12905 gnd.t40 gnd.n3391 6.05496
R12906 gnd.n3392 gnd.t29 6.05496
R12907 gnd.t356 gnd.n2790 6.05496
R12908 gnd.t30 gnd.n3556 6.05496
R12909 gnd.n4461 gnd.t234 6.05496
R12910 gnd.n4588 gnd.t255 6.05496
R12911 gnd.t17 gnd.n2004 6.05496
R12912 gnd.n5370 gnd.t366 6.05496
R12913 gnd.n5845 gnd.t192 6.05496
R12914 gnd.n133 gnd.t194 6.05496
R12915 gnd.n3915 gnd.n3885 5.81868
R12916 gnd.n3883 gnd.n3853 5.81868
R12917 gnd.n3851 gnd.n3821 5.81868
R12918 gnd.n3820 gnd.n3790 5.81868
R12919 gnd.n3788 gnd.n3758 5.81868
R12920 gnd.n3756 gnd.n3726 5.81868
R12921 gnd.n3724 gnd.n3694 5.81868
R12922 gnd.n3693 gnd.n3663 5.81868
R12923 gnd.n5613 gnd.n1437 5.62001
R12924 gnd.n6346 gnd.n1121 5.62001
R12925 gnd.n6346 gnd.n1122 5.62001
R12926 gnd.n5479 gnd.n1437 5.62001
R12927 gnd.n3143 gnd.n3138 5.4308
R12928 gnd.n3960 gnd.n2632 5.4308
R12929 gnd.n3459 gnd.t24 5.41765
R12930 gnd.t10 gnd.n3482 5.41765
R12931 gnd.t62 gnd.n2720 5.41765
R12932 gnd.n6471 gnd.t273 5.41765
R12933 gnd.t221 gnd.n2432 5.41765
R12934 gnd.n7287 gnd.t230 5.41765
R12935 gnd.n7611 gnd.t204 5.41765
R12936 gnd.n5035 gnd.t180 5.09899
R12937 gnd.n5065 gnd.n2012 5.09899
R12938 gnd.n5072 gnd.n2005 5.09899
R12939 gnd.t71 gnd.n5126 5.09899
R12940 gnd.n5224 gnd.n1920 5.09899
R12941 gnd.n5232 gnd.n1913 5.09899
R12942 gnd.t51 gnd.n5317 5.09899
R12943 gnd.n5369 gnd.n1830 5.09899
R12944 gnd.n5376 gnd.n1823 5.09899
R12945 gnd.n3913 gnd.n3912 5.04292
R12946 gnd.n3881 gnd.n3880 5.04292
R12947 gnd.n3849 gnd.n3848 5.04292
R12948 gnd.n3818 gnd.n3817 5.04292
R12949 gnd.n3786 gnd.n3785 5.04292
R12950 gnd.n3754 gnd.n3753 5.04292
R12951 gnd.n3722 gnd.n3721 5.04292
R12952 gnd.n3691 gnd.n3690 5.04292
R12953 gnd.n3422 gnd.t32 4.78034
R12954 gnd.n2745 gnd.t31 4.78034
R12955 gnd.n4481 gnd.t198 4.78034
R12956 gnd.n6458 gnd.t210 4.78034
R12957 gnd.n4846 gnd.t52 4.78034
R12958 gnd.n5616 gnd.t161 4.78034
R12959 gnd.n5643 gnd.t43 4.78034
R12960 gnd.n5898 gnd.t261 4.78034
R12961 gnd.n7597 gnd.t223 4.78034
R12962 gnd.n2864 gnd.n2861 4.74817
R12963 gnd.n2914 gnd.n2796 4.74817
R12964 gnd.n2901 gnd.n2795 4.74817
R12965 gnd.n2794 gnd.n2793 4.74817
R12966 gnd.n2910 gnd.n2861 4.74817
R12967 gnd.n2911 gnd.n2796 4.74817
R12968 gnd.n2913 gnd.n2795 4.74817
R12969 gnd.n2900 gnd.n2794 4.74817
R12970 gnd.n5890 gnd.n101 4.74817
R12971 gnd.n386 gnd.n99 4.74817
R12972 gnd.n7609 gnd.n94 4.74817
R12973 gnd.n7607 gnd.n95 4.74817
R12974 gnd.n1593 gnd.n101 4.74817
R12975 gnd.n7285 gnd.n99 4.74817
R12976 gnd.n385 gnd.n94 4.74817
R12977 gnd.n7608 gnd.n7607 4.74817
R12978 gnd.n2455 gnd.n951 4.74817
R12979 gnd.n6468 gnd.n945 4.74817
R12980 gnd.n4532 gnd.n950 4.74817
R12981 gnd.n952 gnd.n949 4.74817
R12982 gnd.n4499 gnd.n951 4.74817
R12983 gnd.n6469 gnd.n6468 4.74817
R12984 gnd.n2435 gnd.n950 4.74817
R12985 gnd.n4533 gnd.n949 4.74817
R12986 gnd.n2859 gnd.n2858 4.74296
R12987 gnd.n82 gnd.n81 4.74296
R12988 gnd.n2827 gnd.n2826 4.7074
R12989 gnd.n2843 gnd.n2842 4.7074
R12990 gnd.n50 gnd.n49 4.7074
R12991 gnd.n66 gnd.n65 4.7074
R12992 gnd.n2859 gnd.n2843 4.65959
R12993 gnd.n82 gnd.n66 4.65959
R12994 gnd.n6028 gnd.n1439 4.6132
R12995 gnd.n6347 gnd.n1120 4.6132
R12996 gnd.t124 gnd.n2031 4.46168
R12997 gnd.n5469 gnd.n5456 4.46111
R12998 gnd.n3898 gnd.n3894 4.38594
R12999 gnd.n3866 gnd.n3862 4.38594
R13000 gnd.n3834 gnd.n3830 4.38594
R13001 gnd.n3803 gnd.n3799 4.38594
R13002 gnd.n3771 gnd.n3767 4.38594
R13003 gnd.n3739 gnd.n3735 4.38594
R13004 gnd.n3707 gnd.n3703 4.38594
R13005 gnd.n3676 gnd.n3672 4.38594
R13006 gnd.n3909 gnd.n3887 4.26717
R13007 gnd.n3877 gnd.n3855 4.26717
R13008 gnd.n3845 gnd.n3823 4.26717
R13009 gnd.n3814 gnd.n3792 4.26717
R13010 gnd.n3782 gnd.n3760 4.26717
R13011 gnd.n3750 gnd.n3728 4.26717
R13012 gnd.n3718 gnd.n3696 4.26717
R13013 gnd.n3687 gnd.n3665 4.26717
R13014 gnd.n3366 gnd.t4 4.14303
R13015 gnd.n3596 gnd.t33 4.14303
R13016 gnd.t200 gnd.n2496 4.14303
R13017 gnd.n6434 gnd.t285 4.14303
R13018 gnd.n2383 gnd.t113 4.14303
R13019 gnd.n5777 gnd.t77 4.14303
R13020 gnd.n5922 gnd.t232 4.14303
R13021 gnd.n7573 gnd.t276 4.14303
R13022 gnd.n3917 gnd.n3916 4.08274
R13023 gnd.n5608 gnd.n5607 4.05904
R13024 gnd.n4903 gnd.n4902 4.05904
R13025 gnd.n6287 gnd.n6280 4.05904
R13026 gnd.n5485 gnd.n5484 4.05904
R13027 gnd.n19 gnd.n9 3.99943
R13028 gnd.n5055 gnd.n5053 3.82437
R13029 gnd.n5093 gnd.t58 3.82437
R13030 gnd.n5204 gnd.n1934 3.82437
R13031 gnd.n5241 gnd.n5240 3.82437
R13032 gnd.n5359 gnd.t23 3.82437
R13033 gnd.n5399 gnd.n1808 3.82437
R13034 gnd.n5415 gnd.t85 3.82437
R13035 gnd.n3439 gnd.n2860 3.81325
R13036 gnd.n2843 gnd.n2827 3.72967
R13037 gnd.n66 gnd.n50 3.72967
R13038 gnd.n3917 gnd.n3789 3.70378
R13039 gnd.n19 gnd.n18 3.60163
R13040 gnd.n3908 gnd.n3889 3.49141
R13041 gnd.n3876 gnd.n3857 3.49141
R13042 gnd.n3844 gnd.n3825 3.49141
R13043 gnd.n3813 gnd.n3794 3.49141
R13044 gnd.n3781 gnd.n3762 3.49141
R13045 gnd.n3749 gnd.n3730 3.49141
R13046 gnd.n3717 gnd.n3698 3.49141
R13047 gnd.n3686 gnd.n3667 3.49141
R13048 gnd.n6046 gnd.n6045 3.29747
R13049 gnd.n6045 gnd.n6044 3.29747
R13050 gnd.n7502 gnd.n7499 3.29747
R13051 gnd.n7503 gnd.n7502 3.29747
R13052 gnd.n4322 gnd.n4321 3.29747
R13053 gnd.n4321 gnd.n4320 3.29747
R13054 gnd.n6363 gnd.n6362 3.29747
R13055 gnd.n6362 gnd.n6361 3.29747
R13056 gnd.n5174 gnd.t66 3.18706
R13057 gnd.n5260 gnd.t5 3.18706
R13058 gnd.t121 gnd.n1790 3.18706
R13059 gnd.n2945 gnd.t4 2.8684
R13060 gnd.n4990 gnd.t64 2.8684
R13061 gnd.n5452 gnd.t27 2.8684
R13062 gnd.n2844 gnd.t296 2.82907
R13063 gnd.n2844 gnd.t351 2.82907
R13064 gnd.n2846 gnd.t256 2.82907
R13065 gnd.n2846 gnd.t340 2.82907
R13066 gnd.n2848 gnd.t203 2.82907
R13067 gnd.n2848 gnd.t321 2.82907
R13068 gnd.n2850 gnd.t343 2.82907
R13069 gnd.n2850 gnd.t251 2.82907
R13070 gnd.n2852 gnd.t283 2.82907
R13071 gnd.n2852 gnd.t267 2.82907
R13072 gnd.n2854 gnd.t265 2.82907
R13073 gnd.n2854 gnd.t235 2.82907
R13074 gnd.n2856 gnd.t269 2.82907
R13075 gnd.n2856 gnd.t311 2.82907
R13076 gnd.n2797 gnd.t302 2.82907
R13077 gnd.n2797 gnd.t318 2.82907
R13078 gnd.n2799 gnd.t299 2.82907
R13079 gnd.n2799 gnd.t344 2.82907
R13080 gnd.n2801 gnd.t293 2.82907
R13081 gnd.n2801 gnd.t307 2.82907
R13082 gnd.n2803 gnd.t319 2.82907
R13083 gnd.n2803 gnd.t222 2.82907
R13084 gnd.n2805 gnd.t305 2.82907
R13085 gnd.n2805 gnd.t301 2.82907
R13086 gnd.n2807 gnd.t334 2.82907
R13087 gnd.n2807 gnd.t329 2.82907
R13088 gnd.n2809 gnd.t244 2.82907
R13089 gnd.n2809 gnd.t314 2.82907
R13090 gnd.n2812 gnd.t286 2.82907
R13091 gnd.n2812 gnd.t272 2.82907
R13092 gnd.n2814 gnd.t275 2.82907
R13093 gnd.n2814 gnd.t300 2.82907
R13094 gnd.n2816 gnd.t248 2.82907
R13095 gnd.n2816 gnd.t287 2.82907
R13096 gnd.n2818 gnd.t288 2.82907
R13097 gnd.n2818 gnd.t268 2.82907
R13098 gnd.n2820 gnd.t199 2.82907
R13099 gnd.n2820 gnd.t250 2.82907
R13100 gnd.n2822 gnd.t239 2.82907
R13101 gnd.n2822 gnd.t290 2.82907
R13102 gnd.n2824 gnd.t229 2.82907
R13103 gnd.n2824 gnd.t201 2.82907
R13104 gnd.n2828 gnd.t333 2.82907
R13105 gnd.n2828 gnd.t292 2.82907
R13106 gnd.n2830 gnd.t309 2.82907
R13107 gnd.n2830 gnd.t258 2.82907
R13108 gnd.n2832 gnd.t295 2.82907
R13109 gnd.n2832 gnd.t211 2.82907
R13110 gnd.n2834 gnd.t274 2.82907
R13111 gnd.n2834 gnd.t312 2.82907
R13112 gnd.n2836 gnd.t327 2.82907
R13113 gnd.n2836 gnd.t308 2.82907
R13114 gnd.n2838 gnd.t315 2.82907
R13115 gnd.n2838 gnd.t304 2.82907
R13116 gnd.n2840 gnd.t320 2.82907
R13117 gnd.n2840 gnd.t348 2.82907
R13118 gnd.n79 gnd.t277 2.82907
R13119 gnd.n79 gnd.t323 2.82907
R13120 gnd.n77 gnd.t338 2.82907
R13121 gnd.n77 gnd.t347 2.82907
R13122 gnd.n75 gnd.t349 2.82907
R13123 gnd.n75 gnd.t246 2.82907
R13124 gnd.n73 gnd.t345 2.82907
R13125 gnd.n73 gnd.t316 2.82907
R13126 gnd.n71 gnd.t294 2.82907
R13127 gnd.n71 gnd.t336 2.82907
R13128 gnd.n69 gnd.t313 2.82907
R13129 gnd.n69 gnd.t346 2.82907
R13130 gnd.n67 gnd.t326 2.82907
R13131 gnd.n67 gnd.t233 2.82907
R13132 gnd.n32 gnd.t337 2.82907
R13133 gnd.n32 gnd.t227 2.82907
R13134 gnd.n30 gnd.t195 2.82907
R13135 gnd.n30 gnd.t214 2.82907
R13136 gnd.n28 gnd.t324 2.82907
R13137 gnd.n28 gnd.t297 2.82907
R13138 gnd.n26 gnd.t282 2.82907
R13139 gnd.n26 gnd.t342 2.82907
R13140 gnd.n24 gnd.t332 2.82907
R13141 gnd.n24 gnd.t259 2.82907
R13142 gnd.n22 gnd.t243 2.82907
R13143 gnd.n22 gnd.t193 2.82907
R13144 gnd.n20 gnd.t341 2.82907
R13145 gnd.n20 gnd.t325 2.82907
R13146 gnd.n47 gnd.t339 2.82907
R13147 gnd.n47 gnd.t242 2.82907
R13148 gnd.n45 gnd.t264 2.82907
R13149 gnd.n45 gnd.t209 2.82907
R13150 gnd.n43 gnd.t216 2.82907
R13151 gnd.n43 gnd.t224 2.82907
R13152 gnd.n41 gnd.t231 2.82907
R13153 gnd.n41 gnd.t260 2.82907
R13154 gnd.n39 gnd.t262 2.82907
R13155 gnd.n39 gnd.t254 2.82907
R13156 gnd.n37 gnd.t279 2.82907
R13157 gnd.n37 gnd.t236 2.82907
R13158 gnd.n35 gnd.t237 2.82907
R13159 gnd.n35 gnd.t252 2.82907
R13160 gnd.n63 gnd.t322 2.82907
R13161 gnd.n63 gnd.t213 2.82907
R13162 gnd.n61 gnd.t266 2.82907
R13163 gnd.n61 gnd.t284 2.82907
R13164 gnd.n59 gnd.t289 2.82907
R13165 gnd.n59 gnd.t310 2.82907
R13166 gnd.n57 gnd.t280 2.82907
R13167 gnd.n57 gnd.t205 2.82907
R13168 gnd.n55 gnd.t330 2.82907
R13169 gnd.n55 gnd.t263 2.82907
R13170 gnd.n53 gnd.t197 2.82907
R13171 gnd.n53 gnd.t281 2.82907
R13172 gnd.n51 gnd.t220 2.82907
R13173 gnd.n51 gnd.t303 2.82907
R13174 gnd.n3905 gnd.n3904 2.71565
R13175 gnd.n3873 gnd.n3872 2.71565
R13176 gnd.n3841 gnd.n3840 2.71565
R13177 gnd.n3810 gnd.n3809 2.71565
R13178 gnd.n3778 gnd.n3777 2.71565
R13179 gnd.n3746 gnd.n3745 2.71565
R13180 gnd.n3714 gnd.n3713 2.71565
R13181 gnd.n3683 gnd.n3682 2.71565
R13182 gnd.n6266 gnd.t99 2.54975
R13183 gnd.n5035 gnd.n5034 2.54975
R13184 gnd.n5107 gnd.n1983 2.54975
R13185 gnd.n5194 gnd.n5193 2.54975
R13186 gnd.n5269 gnd.n1887 2.54975
R13187 gnd.n5309 gnd.n1845 2.54975
R13188 gnd.n5407 gnd.n1801 2.54975
R13189 gnd.t190 gnd.n5441 2.54975
R13190 gnd.n3439 gnd.n2861 2.27742
R13191 gnd.n3439 gnd.n2796 2.27742
R13192 gnd.n3439 gnd.n2795 2.27742
R13193 gnd.n3439 gnd.n2794 2.27742
R13194 gnd.n7606 gnd.n101 2.27742
R13195 gnd.n7606 gnd.n99 2.27742
R13196 gnd.n7606 gnd.n94 2.27742
R13197 gnd.n7607 gnd.n7606 2.27742
R13198 gnd.n6467 gnd.n951 2.27742
R13199 gnd.n6468 gnd.n6467 2.27742
R13200 gnd.n6467 gnd.n950 2.27742
R13201 gnd.n6467 gnd.n949 2.27742
R13202 gnd.n3293 gnd.t109 2.23109
R13203 gnd.n2916 gnd.t32 2.23109
R13204 gnd.n4564 gnd.t202 2.23109
R13205 gnd.n1594 gnd.t253 2.23109
R13206 gnd.n3901 gnd.n3891 1.93989
R13207 gnd.n3869 gnd.n3859 1.93989
R13208 gnd.n3837 gnd.n3827 1.93989
R13209 gnd.n3806 gnd.n3796 1.93989
R13210 gnd.n3774 gnd.n3764 1.93989
R13211 gnd.n3742 gnd.n3732 1.93989
R13212 gnd.n3710 gnd.n3700 1.93989
R13213 gnd.n3679 gnd.n3669 1.93989
R13214 gnd.n4892 gnd.t139 1.91244
R13215 gnd.n1934 gnd.t61 1.91244
R13216 gnd.n5241 gnd.t14 1.91244
R13217 gnd.t358 gnd.n3304 1.59378
R13218 gnd.n3483 gnd.t10 1.59378
R13219 gnd.n2729 gnd.t62 1.59378
R13220 gnd.n4625 gnd.t257 1.59378
R13221 gnd.n5047 gnd.t59 1.59378
R13222 gnd.t67 gnd.n1979 1.59378
R13223 gnd.n5328 gnd.t354 1.59378
R13224 gnd.n5382 gnd.t56 1.59378
R13225 gnd.n1613 gnd.t196 1.59378
R13226 gnd.n4961 gnd.n1183 1.27512
R13227 gnd.n4984 gnd.t73 1.27512
R13228 gnd.n4973 gnd.n4970 1.27512
R13229 gnd.n5055 gnd.t39 1.27512
R13230 gnd.n5119 gnd.n1973 1.27512
R13231 gnd.n5162 gnd.n1947 1.27512
R13232 gnd.n5279 gnd.n1880 1.27512
R13233 gnd.n5294 gnd.n1863 1.27512
R13234 gnd.n5399 gnd.t16 1.27512
R13235 gnd.n5442 gnd.n1784 1.27512
R13236 gnd.n5441 gnd.t102 1.27512
R13237 gnd.n5415 gnd.n1728 1.27512
R13238 gnd.n3146 gnd.n3138 1.16414
R13239 gnd.n3963 gnd.n2632 1.16414
R13240 gnd.n3900 gnd.n3893 1.16414
R13241 gnd.n3868 gnd.n3861 1.16414
R13242 gnd.n3836 gnd.n3829 1.16414
R13243 gnd.n3805 gnd.n3798 1.16414
R13244 gnd.n3773 gnd.n3766 1.16414
R13245 gnd.n3741 gnd.n3734 1.16414
R13246 gnd.n3709 gnd.n3702 1.16414
R13247 gnd.n3678 gnd.n3671 1.16414
R13248 gnd.n6028 gnd.n6027 0.970197
R13249 gnd.n6347 gnd.n1117 0.970197
R13250 gnd.n3884 gnd.n3852 0.962709
R13251 gnd.n3916 gnd.n3884 0.962709
R13252 gnd.n3757 gnd.n3725 0.962709
R13253 gnd.n3789 gnd.n3757 0.962709
R13254 gnd.n3392 gnd.t40 0.956468
R13255 gnd.n3557 gnd.t30 0.956468
R13256 gnd.n4671 gnd.t206 0.956468
R13257 gnd.n5749 gnd.t217 0.956468
R13258 gnd.n2 gnd.n1 0.672012
R13259 gnd.n3 gnd.n2 0.672012
R13260 gnd.n4 gnd.n3 0.672012
R13261 gnd.n5 gnd.n4 0.672012
R13262 gnd.n6 gnd.n5 0.672012
R13263 gnd.n7 gnd.n6 0.672012
R13264 gnd.n8 gnd.n7 0.672012
R13265 gnd.n9 gnd.n8 0.672012
R13266 gnd.n11 gnd.n10 0.672012
R13267 gnd.n12 gnd.n11 0.672012
R13268 gnd.n13 gnd.n12 0.672012
R13269 gnd.n14 gnd.n13 0.672012
R13270 gnd.n15 gnd.n14 0.672012
R13271 gnd.n16 gnd.n15 0.672012
R13272 gnd.n17 gnd.n16 0.672012
R13273 gnd.n18 gnd.n17 0.672012
R13274 gnd gnd.n0 0.665707
R13275 gnd.n2858 gnd.n2857 0.573776
R13276 gnd.n2857 gnd.n2855 0.573776
R13277 gnd.n2855 gnd.n2853 0.573776
R13278 gnd.n2853 gnd.n2851 0.573776
R13279 gnd.n2851 gnd.n2849 0.573776
R13280 gnd.n2849 gnd.n2847 0.573776
R13281 gnd.n2847 gnd.n2845 0.573776
R13282 gnd.n2811 gnd.n2810 0.573776
R13283 gnd.n2810 gnd.n2808 0.573776
R13284 gnd.n2808 gnd.n2806 0.573776
R13285 gnd.n2806 gnd.n2804 0.573776
R13286 gnd.n2804 gnd.n2802 0.573776
R13287 gnd.n2802 gnd.n2800 0.573776
R13288 gnd.n2800 gnd.n2798 0.573776
R13289 gnd.n2826 gnd.n2825 0.573776
R13290 gnd.n2825 gnd.n2823 0.573776
R13291 gnd.n2823 gnd.n2821 0.573776
R13292 gnd.n2821 gnd.n2819 0.573776
R13293 gnd.n2819 gnd.n2817 0.573776
R13294 gnd.n2817 gnd.n2815 0.573776
R13295 gnd.n2815 gnd.n2813 0.573776
R13296 gnd.n2842 gnd.n2841 0.573776
R13297 gnd.n2841 gnd.n2839 0.573776
R13298 gnd.n2839 gnd.n2837 0.573776
R13299 gnd.n2837 gnd.n2835 0.573776
R13300 gnd.n2835 gnd.n2833 0.573776
R13301 gnd.n2833 gnd.n2831 0.573776
R13302 gnd.n2831 gnd.n2829 0.573776
R13303 gnd.n70 gnd.n68 0.573776
R13304 gnd.n72 gnd.n70 0.573776
R13305 gnd.n74 gnd.n72 0.573776
R13306 gnd.n76 gnd.n74 0.573776
R13307 gnd.n78 gnd.n76 0.573776
R13308 gnd.n80 gnd.n78 0.573776
R13309 gnd.n81 gnd.n80 0.573776
R13310 gnd.n23 gnd.n21 0.573776
R13311 gnd.n25 gnd.n23 0.573776
R13312 gnd.n27 gnd.n25 0.573776
R13313 gnd.n29 gnd.n27 0.573776
R13314 gnd.n31 gnd.n29 0.573776
R13315 gnd.n33 gnd.n31 0.573776
R13316 gnd.n34 gnd.n33 0.573776
R13317 gnd.n38 gnd.n36 0.573776
R13318 gnd.n40 gnd.n38 0.573776
R13319 gnd.n42 gnd.n40 0.573776
R13320 gnd.n44 gnd.n42 0.573776
R13321 gnd.n46 gnd.n44 0.573776
R13322 gnd.n48 gnd.n46 0.573776
R13323 gnd.n49 gnd.n48 0.573776
R13324 gnd.n54 gnd.n52 0.573776
R13325 gnd.n56 gnd.n54 0.573776
R13326 gnd.n58 gnd.n56 0.573776
R13327 gnd.n60 gnd.n58 0.573776
R13328 gnd.n62 gnd.n60 0.573776
R13329 gnd.n64 gnd.n62 0.573776
R13330 gnd.n65 gnd.n64 0.573776
R13331 gnd.n7618 gnd.n7617 0.553847
R13332 gnd.n7391 gnd.n7390 0.505073
R13333 gnd.n4201 gnd.n4199 0.505073
R13334 gnd.n3619 gnd.n2636 0.486781
R13335 gnd.n3195 gnd.n3194 0.48678
R13336 gnd.n3937 gnd.n2590 0.480683
R13337 gnd.n3279 gnd.n3278 0.480683
R13338 gnd.n6644 gnd.n6643 0.480683
R13339 gnd.n7064 gnd.n7063 0.480683
R13340 gnd.n7277 gnd.n7276 0.480683
R13341 gnd.n2428 gnd.n936 0.480683
R13342 gnd.n7534 gnd.n7533 0.470012
R13343 gnd.n1490 gnd.n1409 0.470012
R13344 gnd.n6395 gnd.n6394 0.470012
R13345 gnd.n4083 gnd.n2549 0.470012
R13346 gnd.n1635 gnd.n1291 0.451719
R13347 gnd.n4785 gnd.n2110 0.451719
R13348 gnd.n2186 gnd.n2185 0.451719
R13349 gnd.n6146 gnd.n6145 0.451719
R13350 gnd.n7606 gnd.n98 0.420375
R13351 gnd.n6467 gnd.n948 0.420375
R13352 gnd.n4716 gnd.n2371 0.388379
R13353 gnd.n3897 gnd.n3896 0.388379
R13354 gnd.n3865 gnd.n3864 0.388379
R13355 gnd.n3833 gnd.n3832 0.388379
R13356 gnd.n3802 gnd.n3801 0.388379
R13357 gnd.n3770 gnd.n3769 0.388379
R13358 gnd.n3738 gnd.n3737 0.388379
R13359 gnd.n3706 gnd.n3705 0.388379
R13360 gnd.n3675 gnd.n3674 0.388379
R13361 gnd.n6090 gnd.n1357 0.388379
R13362 gnd.n7618 gnd.n19 0.374463
R13363 gnd gnd.n7618 0.367492
R13364 gnd.n2691 gnd.t3 0.319156
R13365 gnd.t61 gnd.t364 0.319156
R13366 gnd.t362 gnd.t14 0.319156
R13367 gnd.n3113 gnd.n3091 0.311721
R13368 gnd.n7424 gnd.n7423 0.293183
R13369 gnd.n4239 gnd.n4238 0.293183
R13370 gnd.n4699 gnd.n4698 0.27489
R13371 gnd.n5735 gnd.n5734 0.27489
R13372 gnd.n4008 gnd.n4007 0.268793
R13373 gnd.n7425 gnd.n7424 0.258122
R13374 gnd.n5966 gnd.n1310 0.258122
R13375 gnd.n2305 gnd.n2304 0.258122
R13376 gnd.n4240 gnd.n4239 0.258122
R13377 gnd.n4007 gnd.n4006 0.241354
R13378 gnd.n1439 gnd.n1436 0.229039
R13379 gnd.n1440 gnd.n1439 0.229039
R13380 gnd.n1120 gnd.n1116 0.229039
R13381 gnd.n2225 gnd.n1120 0.229039
R13382 gnd.n3267 gnd.n3066 0.206293
R13383 gnd.n2860 gnd.n0 0.169152
R13384 gnd.n3914 gnd.n3886 0.155672
R13385 gnd.n3907 gnd.n3886 0.155672
R13386 gnd.n3907 gnd.n3906 0.155672
R13387 gnd.n3906 gnd.n3890 0.155672
R13388 gnd.n3899 gnd.n3890 0.155672
R13389 gnd.n3899 gnd.n3898 0.155672
R13390 gnd.n3882 gnd.n3854 0.155672
R13391 gnd.n3875 gnd.n3854 0.155672
R13392 gnd.n3875 gnd.n3874 0.155672
R13393 gnd.n3874 gnd.n3858 0.155672
R13394 gnd.n3867 gnd.n3858 0.155672
R13395 gnd.n3867 gnd.n3866 0.155672
R13396 gnd.n3850 gnd.n3822 0.155672
R13397 gnd.n3843 gnd.n3822 0.155672
R13398 gnd.n3843 gnd.n3842 0.155672
R13399 gnd.n3842 gnd.n3826 0.155672
R13400 gnd.n3835 gnd.n3826 0.155672
R13401 gnd.n3835 gnd.n3834 0.155672
R13402 gnd.n3819 gnd.n3791 0.155672
R13403 gnd.n3812 gnd.n3791 0.155672
R13404 gnd.n3812 gnd.n3811 0.155672
R13405 gnd.n3811 gnd.n3795 0.155672
R13406 gnd.n3804 gnd.n3795 0.155672
R13407 gnd.n3804 gnd.n3803 0.155672
R13408 gnd.n3787 gnd.n3759 0.155672
R13409 gnd.n3780 gnd.n3759 0.155672
R13410 gnd.n3780 gnd.n3779 0.155672
R13411 gnd.n3779 gnd.n3763 0.155672
R13412 gnd.n3772 gnd.n3763 0.155672
R13413 gnd.n3772 gnd.n3771 0.155672
R13414 gnd.n3755 gnd.n3727 0.155672
R13415 gnd.n3748 gnd.n3727 0.155672
R13416 gnd.n3748 gnd.n3747 0.155672
R13417 gnd.n3747 gnd.n3731 0.155672
R13418 gnd.n3740 gnd.n3731 0.155672
R13419 gnd.n3740 gnd.n3739 0.155672
R13420 gnd.n3723 gnd.n3695 0.155672
R13421 gnd.n3716 gnd.n3695 0.155672
R13422 gnd.n3716 gnd.n3715 0.155672
R13423 gnd.n3715 gnd.n3699 0.155672
R13424 gnd.n3708 gnd.n3699 0.155672
R13425 gnd.n3708 gnd.n3707 0.155672
R13426 gnd.n3692 gnd.n3664 0.155672
R13427 gnd.n3685 gnd.n3664 0.155672
R13428 gnd.n3685 gnd.n3684 0.155672
R13429 gnd.n3684 gnd.n3668 0.155672
R13430 gnd.n3677 gnd.n3668 0.155672
R13431 gnd.n3677 gnd.n3676 0.155672
R13432 gnd.n4039 gnd.n2590 0.152939
R13433 gnd.n4039 gnd.n4038 0.152939
R13434 gnd.n4038 gnd.n4037 0.152939
R13435 gnd.n4037 gnd.n2592 0.152939
R13436 gnd.n2593 gnd.n2592 0.152939
R13437 gnd.n2594 gnd.n2593 0.152939
R13438 gnd.n2595 gnd.n2594 0.152939
R13439 gnd.n2596 gnd.n2595 0.152939
R13440 gnd.n2597 gnd.n2596 0.152939
R13441 gnd.n2598 gnd.n2597 0.152939
R13442 gnd.n2599 gnd.n2598 0.152939
R13443 gnd.n2600 gnd.n2599 0.152939
R13444 gnd.n2601 gnd.n2600 0.152939
R13445 gnd.n2602 gnd.n2601 0.152939
R13446 gnd.n4009 gnd.n2602 0.152939
R13447 gnd.n4009 gnd.n4008 0.152939
R13448 gnd.n3280 gnd.n3279 0.152939
R13449 gnd.n3280 gnd.n2984 0.152939
R13450 gnd.n3308 gnd.n2984 0.152939
R13451 gnd.n3309 gnd.n3308 0.152939
R13452 gnd.n3310 gnd.n3309 0.152939
R13453 gnd.n3311 gnd.n3310 0.152939
R13454 gnd.n3311 gnd.n2956 0.152939
R13455 gnd.n3338 gnd.n2956 0.152939
R13456 gnd.n3339 gnd.n3338 0.152939
R13457 gnd.n3340 gnd.n3339 0.152939
R13458 gnd.n3340 gnd.n2934 0.152939
R13459 gnd.n3369 gnd.n2934 0.152939
R13460 gnd.n3370 gnd.n3369 0.152939
R13461 gnd.n3371 gnd.n3370 0.152939
R13462 gnd.n3372 gnd.n3371 0.152939
R13463 gnd.n3374 gnd.n3372 0.152939
R13464 gnd.n3374 gnd.n3373 0.152939
R13465 gnd.n3373 gnd.n2883 0.152939
R13466 gnd.n2884 gnd.n2883 0.152939
R13467 gnd.n2885 gnd.n2884 0.152939
R13468 gnd.n2904 gnd.n2885 0.152939
R13469 gnd.n2905 gnd.n2904 0.152939
R13470 gnd.n2905 gnd.n2787 0.152939
R13471 gnd.n3464 gnd.n2787 0.152939
R13472 gnd.n3465 gnd.n3464 0.152939
R13473 gnd.n3466 gnd.n3465 0.152939
R13474 gnd.n3467 gnd.n3466 0.152939
R13475 gnd.n3467 gnd.n2760 0.152939
R13476 gnd.n3504 gnd.n2760 0.152939
R13477 gnd.n3505 gnd.n3504 0.152939
R13478 gnd.n3506 gnd.n3505 0.152939
R13479 gnd.n3507 gnd.n3506 0.152939
R13480 gnd.n3507 gnd.n2733 0.152939
R13481 gnd.n3549 gnd.n2733 0.152939
R13482 gnd.n3550 gnd.n3549 0.152939
R13483 gnd.n3551 gnd.n3550 0.152939
R13484 gnd.n3552 gnd.n3551 0.152939
R13485 gnd.n3552 gnd.n2705 0.152939
R13486 gnd.n3589 gnd.n2705 0.152939
R13487 gnd.n3590 gnd.n3589 0.152939
R13488 gnd.n3591 gnd.n3590 0.152939
R13489 gnd.n3592 gnd.n3591 0.152939
R13490 gnd.n3592 gnd.n2678 0.152939
R13491 gnd.n3638 gnd.n2678 0.152939
R13492 gnd.n3639 gnd.n3638 0.152939
R13493 gnd.n3640 gnd.n3639 0.152939
R13494 gnd.n3641 gnd.n3640 0.152939
R13495 gnd.n3641 gnd.n2651 0.152939
R13496 gnd.n3933 gnd.n2651 0.152939
R13497 gnd.n3934 gnd.n3933 0.152939
R13498 gnd.n3935 gnd.n3934 0.152939
R13499 gnd.n3936 gnd.n3935 0.152939
R13500 gnd.n3937 gnd.n3936 0.152939
R13501 gnd.n3278 gnd.n3008 0.152939
R13502 gnd.n3029 gnd.n3008 0.152939
R13503 gnd.n3030 gnd.n3029 0.152939
R13504 gnd.n3036 gnd.n3030 0.152939
R13505 gnd.n3037 gnd.n3036 0.152939
R13506 gnd.n3038 gnd.n3037 0.152939
R13507 gnd.n3038 gnd.n3027 0.152939
R13508 gnd.n3046 gnd.n3027 0.152939
R13509 gnd.n3047 gnd.n3046 0.152939
R13510 gnd.n3048 gnd.n3047 0.152939
R13511 gnd.n3048 gnd.n3025 0.152939
R13512 gnd.n3056 gnd.n3025 0.152939
R13513 gnd.n3057 gnd.n3056 0.152939
R13514 gnd.n3058 gnd.n3057 0.152939
R13515 gnd.n3058 gnd.n3023 0.152939
R13516 gnd.n3066 gnd.n3023 0.152939
R13517 gnd.n4006 gnd.n2607 0.152939
R13518 gnd.n2609 gnd.n2607 0.152939
R13519 gnd.n2610 gnd.n2609 0.152939
R13520 gnd.n2611 gnd.n2610 0.152939
R13521 gnd.n2612 gnd.n2611 0.152939
R13522 gnd.n2613 gnd.n2612 0.152939
R13523 gnd.n2614 gnd.n2613 0.152939
R13524 gnd.n2615 gnd.n2614 0.152939
R13525 gnd.n2616 gnd.n2615 0.152939
R13526 gnd.n2617 gnd.n2616 0.152939
R13527 gnd.n2618 gnd.n2617 0.152939
R13528 gnd.n2619 gnd.n2618 0.152939
R13529 gnd.n2620 gnd.n2619 0.152939
R13530 gnd.n2621 gnd.n2620 0.152939
R13531 gnd.n2622 gnd.n2621 0.152939
R13532 gnd.n2623 gnd.n2622 0.152939
R13533 gnd.n2624 gnd.n2623 0.152939
R13534 gnd.n2625 gnd.n2624 0.152939
R13535 gnd.n2626 gnd.n2625 0.152939
R13536 gnd.n2627 gnd.n2626 0.152939
R13537 gnd.n2628 gnd.n2627 0.152939
R13538 gnd.n2629 gnd.n2628 0.152939
R13539 gnd.n2633 gnd.n2629 0.152939
R13540 gnd.n2634 gnd.n2633 0.152939
R13541 gnd.n2635 gnd.n2634 0.152939
R13542 gnd.n2636 gnd.n2635 0.152939
R13543 gnd.n3441 gnd.n3440 0.152939
R13544 gnd.n3442 gnd.n3441 0.152939
R13545 gnd.n3443 gnd.n3442 0.152939
R13546 gnd.n3444 gnd.n3443 0.152939
R13547 gnd.n3445 gnd.n3444 0.152939
R13548 gnd.n3446 gnd.n3445 0.152939
R13549 gnd.n3446 gnd.n2741 0.152939
R13550 gnd.n3525 gnd.n2741 0.152939
R13551 gnd.n3526 gnd.n3525 0.152939
R13552 gnd.n3527 gnd.n3526 0.152939
R13553 gnd.n3528 gnd.n3527 0.152939
R13554 gnd.n3529 gnd.n3528 0.152939
R13555 gnd.n3530 gnd.n3529 0.152939
R13556 gnd.n3531 gnd.n3530 0.152939
R13557 gnd.n3532 gnd.n3531 0.152939
R13558 gnd.n3533 gnd.n3532 0.152939
R13559 gnd.n3533 gnd.n2685 0.152939
R13560 gnd.n3610 gnd.n2685 0.152939
R13561 gnd.n3611 gnd.n3610 0.152939
R13562 gnd.n3612 gnd.n3611 0.152939
R13563 gnd.n3613 gnd.n3612 0.152939
R13564 gnd.n3614 gnd.n3613 0.152939
R13565 gnd.n3615 gnd.n3614 0.152939
R13566 gnd.n3616 gnd.n3615 0.152939
R13567 gnd.n3617 gnd.n3616 0.152939
R13568 gnd.n3618 gnd.n3617 0.152939
R13569 gnd.n3620 gnd.n3618 0.152939
R13570 gnd.n3620 gnd.n3619 0.152939
R13571 gnd.n3196 gnd.n3195 0.152939
R13572 gnd.n3196 gnd.n3086 0.152939
R13573 gnd.n3211 gnd.n3086 0.152939
R13574 gnd.n3212 gnd.n3211 0.152939
R13575 gnd.n3213 gnd.n3212 0.152939
R13576 gnd.n3213 gnd.n3074 0.152939
R13577 gnd.n3227 gnd.n3074 0.152939
R13578 gnd.n3228 gnd.n3227 0.152939
R13579 gnd.n3229 gnd.n3228 0.152939
R13580 gnd.n3230 gnd.n3229 0.152939
R13581 gnd.n3231 gnd.n3230 0.152939
R13582 gnd.n3232 gnd.n3231 0.152939
R13583 gnd.n3233 gnd.n3232 0.152939
R13584 gnd.n3234 gnd.n3233 0.152939
R13585 gnd.n3235 gnd.n3234 0.152939
R13586 gnd.n3236 gnd.n3235 0.152939
R13587 gnd.n3237 gnd.n3236 0.152939
R13588 gnd.n3238 gnd.n3237 0.152939
R13589 gnd.n3239 gnd.n3238 0.152939
R13590 gnd.n3240 gnd.n3239 0.152939
R13591 gnd.n3241 gnd.n3240 0.152939
R13592 gnd.n3241 gnd.n2940 0.152939
R13593 gnd.n3358 gnd.n2940 0.152939
R13594 gnd.n3359 gnd.n3358 0.152939
R13595 gnd.n3360 gnd.n3359 0.152939
R13596 gnd.n3361 gnd.n3360 0.152939
R13597 gnd.n3361 gnd.n2862 0.152939
R13598 gnd.n3438 gnd.n2862 0.152939
R13599 gnd.n3114 gnd.n3113 0.152939
R13600 gnd.n3115 gnd.n3114 0.152939
R13601 gnd.n3116 gnd.n3115 0.152939
R13602 gnd.n3117 gnd.n3116 0.152939
R13603 gnd.n3118 gnd.n3117 0.152939
R13604 gnd.n3119 gnd.n3118 0.152939
R13605 gnd.n3120 gnd.n3119 0.152939
R13606 gnd.n3121 gnd.n3120 0.152939
R13607 gnd.n3122 gnd.n3121 0.152939
R13608 gnd.n3123 gnd.n3122 0.152939
R13609 gnd.n3124 gnd.n3123 0.152939
R13610 gnd.n3125 gnd.n3124 0.152939
R13611 gnd.n3126 gnd.n3125 0.152939
R13612 gnd.n3127 gnd.n3126 0.152939
R13613 gnd.n3128 gnd.n3127 0.152939
R13614 gnd.n3129 gnd.n3128 0.152939
R13615 gnd.n3130 gnd.n3129 0.152939
R13616 gnd.n3131 gnd.n3130 0.152939
R13617 gnd.n3132 gnd.n3131 0.152939
R13618 gnd.n3133 gnd.n3132 0.152939
R13619 gnd.n3134 gnd.n3133 0.152939
R13620 gnd.n3135 gnd.n3134 0.152939
R13621 gnd.n3139 gnd.n3135 0.152939
R13622 gnd.n3140 gnd.n3139 0.152939
R13623 gnd.n3140 gnd.n3097 0.152939
R13624 gnd.n3194 gnd.n3097 0.152939
R13625 gnd.n6645 gnd.n6644 0.152939
R13626 gnd.n6645 gnd.n763 0.152939
R13627 gnd.n6653 gnd.n763 0.152939
R13628 gnd.n6654 gnd.n6653 0.152939
R13629 gnd.n6655 gnd.n6654 0.152939
R13630 gnd.n6655 gnd.n757 0.152939
R13631 gnd.n6663 gnd.n757 0.152939
R13632 gnd.n6664 gnd.n6663 0.152939
R13633 gnd.n6665 gnd.n6664 0.152939
R13634 gnd.n6665 gnd.n751 0.152939
R13635 gnd.n6673 gnd.n751 0.152939
R13636 gnd.n6674 gnd.n6673 0.152939
R13637 gnd.n6675 gnd.n6674 0.152939
R13638 gnd.n6675 gnd.n745 0.152939
R13639 gnd.n6683 gnd.n745 0.152939
R13640 gnd.n6684 gnd.n6683 0.152939
R13641 gnd.n6685 gnd.n6684 0.152939
R13642 gnd.n6685 gnd.n739 0.152939
R13643 gnd.n6693 gnd.n739 0.152939
R13644 gnd.n6694 gnd.n6693 0.152939
R13645 gnd.n6695 gnd.n6694 0.152939
R13646 gnd.n6695 gnd.n733 0.152939
R13647 gnd.n6703 gnd.n733 0.152939
R13648 gnd.n6704 gnd.n6703 0.152939
R13649 gnd.n6705 gnd.n6704 0.152939
R13650 gnd.n6705 gnd.n727 0.152939
R13651 gnd.n6713 gnd.n727 0.152939
R13652 gnd.n6714 gnd.n6713 0.152939
R13653 gnd.n6715 gnd.n6714 0.152939
R13654 gnd.n6715 gnd.n721 0.152939
R13655 gnd.n6723 gnd.n721 0.152939
R13656 gnd.n6724 gnd.n6723 0.152939
R13657 gnd.n6725 gnd.n6724 0.152939
R13658 gnd.n6725 gnd.n715 0.152939
R13659 gnd.n6733 gnd.n715 0.152939
R13660 gnd.n6734 gnd.n6733 0.152939
R13661 gnd.n6735 gnd.n6734 0.152939
R13662 gnd.n6735 gnd.n709 0.152939
R13663 gnd.n6743 gnd.n709 0.152939
R13664 gnd.n6744 gnd.n6743 0.152939
R13665 gnd.n6745 gnd.n6744 0.152939
R13666 gnd.n6745 gnd.n703 0.152939
R13667 gnd.n6753 gnd.n703 0.152939
R13668 gnd.n6754 gnd.n6753 0.152939
R13669 gnd.n6755 gnd.n6754 0.152939
R13670 gnd.n6755 gnd.n697 0.152939
R13671 gnd.n6763 gnd.n697 0.152939
R13672 gnd.n6764 gnd.n6763 0.152939
R13673 gnd.n6765 gnd.n6764 0.152939
R13674 gnd.n6765 gnd.n691 0.152939
R13675 gnd.n6773 gnd.n691 0.152939
R13676 gnd.n6774 gnd.n6773 0.152939
R13677 gnd.n6775 gnd.n6774 0.152939
R13678 gnd.n6775 gnd.n685 0.152939
R13679 gnd.n6783 gnd.n685 0.152939
R13680 gnd.n6784 gnd.n6783 0.152939
R13681 gnd.n6785 gnd.n6784 0.152939
R13682 gnd.n6785 gnd.n679 0.152939
R13683 gnd.n6793 gnd.n679 0.152939
R13684 gnd.n6794 gnd.n6793 0.152939
R13685 gnd.n6795 gnd.n6794 0.152939
R13686 gnd.n6795 gnd.n673 0.152939
R13687 gnd.n6803 gnd.n673 0.152939
R13688 gnd.n6804 gnd.n6803 0.152939
R13689 gnd.n6805 gnd.n6804 0.152939
R13690 gnd.n6805 gnd.n667 0.152939
R13691 gnd.n6813 gnd.n667 0.152939
R13692 gnd.n6814 gnd.n6813 0.152939
R13693 gnd.n6815 gnd.n6814 0.152939
R13694 gnd.n6815 gnd.n661 0.152939
R13695 gnd.n6823 gnd.n661 0.152939
R13696 gnd.n6824 gnd.n6823 0.152939
R13697 gnd.n6825 gnd.n6824 0.152939
R13698 gnd.n6825 gnd.n655 0.152939
R13699 gnd.n6833 gnd.n655 0.152939
R13700 gnd.n6834 gnd.n6833 0.152939
R13701 gnd.n6835 gnd.n6834 0.152939
R13702 gnd.n6835 gnd.n649 0.152939
R13703 gnd.n6843 gnd.n649 0.152939
R13704 gnd.n6844 gnd.n6843 0.152939
R13705 gnd.n6845 gnd.n6844 0.152939
R13706 gnd.n6845 gnd.n643 0.152939
R13707 gnd.n6853 gnd.n643 0.152939
R13708 gnd.n6854 gnd.n6853 0.152939
R13709 gnd.n6855 gnd.n6854 0.152939
R13710 gnd.n6855 gnd.n637 0.152939
R13711 gnd.n6863 gnd.n637 0.152939
R13712 gnd.n6864 gnd.n6863 0.152939
R13713 gnd.n6865 gnd.n6864 0.152939
R13714 gnd.n6865 gnd.n631 0.152939
R13715 gnd.n6873 gnd.n631 0.152939
R13716 gnd.n6874 gnd.n6873 0.152939
R13717 gnd.n6875 gnd.n6874 0.152939
R13718 gnd.n6875 gnd.n625 0.152939
R13719 gnd.n6883 gnd.n625 0.152939
R13720 gnd.n6884 gnd.n6883 0.152939
R13721 gnd.n6885 gnd.n6884 0.152939
R13722 gnd.n6885 gnd.n619 0.152939
R13723 gnd.n6893 gnd.n619 0.152939
R13724 gnd.n6894 gnd.n6893 0.152939
R13725 gnd.n6895 gnd.n6894 0.152939
R13726 gnd.n6895 gnd.n613 0.152939
R13727 gnd.n6903 gnd.n613 0.152939
R13728 gnd.n6904 gnd.n6903 0.152939
R13729 gnd.n6905 gnd.n6904 0.152939
R13730 gnd.n6905 gnd.n607 0.152939
R13731 gnd.n6913 gnd.n607 0.152939
R13732 gnd.n6914 gnd.n6913 0.152939
R13733 gnd.n6915 gnd.n6914 0.152939
R13734 gnd.n6915 gnd.n601 0.152939
R13735 gnd.n6923 gnd.n601 0.152939
R13736 gnd.n6924 gnd.n6923 0.152939
R13737 gnd.n6925 gnd.n6924 0.152939
R13738 gnd.n6925 gnd.n595 0.152939
R13739 gnd.n6933 gnd.n595 0.152939
R13740 gnd.n6934 gnd.n6933 0.152939
R13741 gnd.n6935 gnd.n6934 0.152939
R13742 gnd.n6935 gnd.n589 0.152939
R13743 gnd.n6943 gnd.n589 0.152939
R13744 gnd.n6944 gnd.n6943 0.152939
R13745 gnd.n6945 gnd.n6944 0.152939
R13746 gnd.n6945 gnd.n583 0.152939
R13747 gnd.n6953 gnd.n583 0.152939
R13748 gnd.n6954 gnd.n6953 0.152939
R13749 gnd.n6955 gnd.n6954 0.152939
R13750 gnd.n6955 gnd.n577 0.152939
R13751 gnd.n6963 gnd.n577 0.152939
R13752 gnd.n6964 gnd.n6963 0.152939
R13753 gnd.n6965 gnd.n6964 0.152939
R13754 gnd.n6965 gnd.n571 0.152939
R13755 gnd.n6973 gnd.n571 0.152939
R13756 gnd.n6974 gnd.n6973 0.152939
R13757 gnd.n6975 gnd.n6974 0.152939
R13758 gnd.n6975 gnd.n565 0.152939
R13759 gnd.n6983 gnd.n565 0.152939
R13760 gnd.n6984 gnd.n6983 0.152939
R13761 gnd.n6985 gnd.n6984 0.152939
R13762 gnd.n6985 gnd.n559 0.152939
R13763 gnd.n6993 gnd.n559 0.152939
R13764 gnd.n6994 gnd.n6993 0.152939
R13765 gnd.n6995 gnd.n6994 0.152939
R13766 gnd.n6995 gnd.n553 0.152939
R13767 gnd.n7003 gnd.n553 0.152939
R13768 gnd.n7004 gnd.n7003 0.152939
R13769 gnd.n7005 gnd.n7004 0.152939
R13770 gnd.n7005 gnd.n547 0.152939
R13771 gnd.n7013 gnd.n547 0.152939
R13772 gnd.n7014 gnd.n7013 0.152939
R13773 gnd.n7015 gnd.n7014 0.152939
R13774 gnd.n7015 gnd.n541 0.152939
R13775 gnd.n7023 gnd.n541 0.152939
R13776 gnd.n7024 gnd.n7023 0.152939
R13777 gnd.n7025 gnd.n7024 0.152939
R13778 gnd.n7025 gnd.n535 0.152939
R13779 gnd.n7033 gnd.n535 0.152939
R13780 gnd.n7034 gnd.n7033 0.152939
R13781 gnd.n7035 gnd.n7034 0.152939
R13782 gnd.n7035 gnd.n529 0.152939
R13783 gnd.n7043 gnd.n529 0.152939
R13784 gnd.n7044 gnd.n7043 0.152939
R13785 gnd.n7045 gnd.n7044 0.152939
R13786 gnd.n7045 gnd.n523 0.152939
R13787 gnd.n7053 gnd.n523 0.152939
R13788 gnd.n7054 gnd.n7053 0.152939
R13789 gnd.n7055 gnd.n7054 0.152939
R13790 gnd.n7055 gnd.n517 0.152939
R13791 gnd.n7063 gnd.n517 0.152939
R13792 gnd.n7065 gnd.n7064 0.152939
R13793 gnd.n7065 gnd.n511 0.152939
R13794 gnd.n7073 gnd.n511 0.152939
R13795 gnd.n7074 gnd.n7073 0.152939
R13796 gnd.n7075 gnd.n7074 0.152939
R13797 gnd.n7075 gnd.n505 0.152939
R13798 gnd.n7083 gnd.n505 0.152939
R13799 gnd.n7084 gnd.n7083 0.152939
R13800 gnd.n7085 gnd.n7084 0.152939
R13801 gnd.n7085 gnd.n499 0.152939
R13802 gnd.n7093 gnd.n499 0.152939
R13803 gnd.n7094 gnd.n7093 0.152939
R13804 gnd.n7095 gnd.n7094 0.152939
R13805 gnd.n7095 gnd.n493 0.152939
R13806 gnd.n7103 gnd.n493 0.152939
R13807 gnd.n7104 gnd.n7103 0.152939
R13808 gnd.n7105 gnd.n7104 0.152939
R13809 gnd.n7105 gnd.n487 0.152939
R13810 gnd.n7113 gnd.n487 0.152939
R13811 gnd.n7114 gnd.n7113 0.152939
R13812 gnd.n7115 gnd.n7114 0.152939
R13813 gnd.n7115 gnd.n481 0.152939
R13814 gnd.n7123 gnd.n481 0.152939
R13815 gnd.n7124 gnd.n7123 0.152939
R13816 gnd.n7125 gnd.n7124 0.152939
R13817 gnd.n7125 gnd.n475 0.152939
R13818 gnd.n7133 gnd.n475 0.152939
R13819 gnd.n7134 gnd.n7133 0.152939
R13820 gnd.n7135 gnd.n7134 0.152939
R13821 gnd.n7135 gnd.n469 0.152939
R13822 gnd.n7143 gnd.n469 0.152939
R13823 gnd.n7144 gnd.n7143 0.152939
R13824 gnd.n7145 gnd.n7144 0.152939
R13825 gnd.n7145 gnd.n463 0.152939
R13826 gnd.n7153 gnd.n463 0.152939
R13827 gnd.n7154 gnd.n7153 0.152939
R13828 gnd.n7155 gnd.n7154 0.152939
R13829 gnd.n7155 gnd.n457 0.152939
R13830 gnd.n7163 gnd.n457 0.152939
R13831 gnd.n7164 gnd.n7163 0.152939
R13832 gnd.n7165 gnd.n7164 0.152939
R13833 gnd.n7165 gnd.n451 0.152939
R13834 gnd.n7173 gnd.n451 0.152939
R13835 gnd.n7174 gnd.n7173 0.152939
R13836 gnd.n7175 gnd.n7174 0.152939
R13837 gnd.n7175 gnd.n445 0.152939
R13838 gnd.n7183 gnd.n445 0.152939
R13839 gnd.n7184 gnd.n7183 0.152939
R13840 gnd.n7185 gnd.n7184 0.152939
R13841 gnd.n7185 gnd.n439 0.152939
R13842 gnd.n7193 gnd.n439 0.152939
R13843 gnd.n7194 gnd.n7193 0.152939
R13844 gnd.n7195 gnd.n7194 0.152939
R13845 gnd.n7195 gnd.n433 0.152939
R13846 gnd.n7203 gnd.n433 0.152939
R13847 gnd.n7204 gnd.n7203 0.152939
R13848 gnd.n7205 gnd.n7204 0.152939
R13849 gnd.n7205 gnd.n427 0.152939
R13850 gnd.n7213 gnd.n427 0.152939
R13851 gnd.n7214 gnd.n7213 0.152939
R13852 gnd.n7215 gnd.n7214 0.152939
R13853 gnd.n7215 gnd.n421 0.152939
R13854 gnd.n7223 gnd.n421 0.152939
R13855 gnd.n7224 gnd.n7223 0.152939
R13856 gnd.n7225 gnd.n7224 0.152939
R13857 gnd.n7225 gnd.n415 0.152939
R13858 gnd.n7233 gnd.n415 0.152939
R13859 gnd.n7234 gnd.n7233 0.152939
R13860 gnd.n7235 gnd.n7234 0.152939
R13861 gnd.n7235 gnd.n409 0.152939
R13862 gnd.n7243 gnd.n409 0.152939
R13863 gnd.n7244 gnd.n7243 0.152939
R13864 gnd.n7245 gnd.n7244 0.152939
R13865 gnd.n7245 gnd.n403 0.152939
R13866 gnd.n7253 gnd.n403 0.152939
R13867 gnd.n7254 gnd.n7253 0.152939
R13868 gnd.n7255 gnd.n7254 0.152939
R13869 gnd.n7255 gnd.n397 0.152939
R13870 gnd.n7263 gnd.n397 0.152939
R13871 gnd.n7264 gnd.n7263 0.152939
R13872 gnd.n7265 gnd.n7264 0.152939
R13873 gnd.n7266 gnd.n7265 0.152939
R13874 gnd.n7266 gnd.n391 0.152939
R13875 gnd.n7276 gnd.n391 0.152939
R13876 gnd.n119 gnd.n96 0.152939
R13877 gnd.n120 gnd.n119 0.152939
R13878 gnd.n121 gnd.n120 0.152939
R13879 gnd.n138 gnd.n121 0.152939
R13880 gnd.n139 gnd.n138 0.152939
R13881 gnd.n140 gnd.n139 0.152939
R13882 gnd.n141 gnd.n140 0.152939
R13883 gnd.n156 gnd.n141 0.152939
R13884 gnd.n157 gnd.n156 0.152939
R13885 gnd.n158 gnd.n157 0.152939
R13886 gnd.n159 gnd.n158 0.152939
R13887 gnd.n176 gnd.n159 0.152939
R13888 gnd.n177 gnd.n176 0.152939
R13889 gnd.n178 gnd.n177 0.152939
R13890 gnd.n179 gnd.n178 0.152939
R13891 gnd.n196 gnd.n179 0.152939
R13892 gnd.n197 gnd.n196 0.152939
R13893 gnd.n198 gnd.n197 0.152939
R13894 gnd.n199 gnd.n198 0.152939
R13895 gnd.n214 gnd.n199 0.152939
R13896 gnd.n7534 gnd.n214 0.152939
R13897 gnd.n7615 gnd.n84 0.152939
R13898 gnd.n7348 gnd.n84 0.152939
R13899 gnd.n7349 gnd.n7348 0.152939
R13900 gnd.n7350 gnd.n7349 0.152939
R13901 gnd.n7350 gnd.n367 0.152939
R13902 gnd.n7355 gnd.n367 0.152939
R13903 gnd.n7356 gnd.n7355 0.152939
R13904 gnd.n7357 gnd.n7356 0.152939
R13905 gnd.n7357 gnd.n364 0.152939
R13906 gnd.n7362 gnd.n364 0.152939
R13907 gnd.n7363 gnd.n7362 0.152939
R13908 gnd.n7364 gnd.n7363 0.152939
R13909 gnd.n7364 gnd.n361 0.152939
R13910 gnd.n7369 gnd.n361 0.152939
R13911 gnd.n7370 gnd.n7369 0.152939
R13912 gnd.n7371 gnd.n7370 0.152939
R13913 gnd.n7371 gnd.n358 0.152939
R13914 gnd.n7376 gnd.n358 0.152939
R13915 gnd.n7377 gnd.n7376 0.152939
R13916 gnd.n7378 gnd.n7377 0.152939
R13917 gnd.n7378 gnd.n355 0.152939
R13918 gnd.n7383 gnd.n355 0.152939
R13919 gnd.n7384 gnd.n7383 0.152939
R13920 gnd.n7385 gnd.n7384 0.152939
R13921 gnd.n7385 gnd.n352 0.152939
R13922 gnd.n7390 gnd.n352 0.152939
R13923 gnd.n7423 gnd.n318 0.152939
R13924 gnd.n320 gnd.n318 0.152939
R13925 gnd.n324 gnd.n320 0.152939
R13926 gnd.n325 gnd.n324 0.152939
R13927 gnd.n326 gnd.n325 0.152939
R13928 gnd.n327 gnd.n326 0.152939
R13929 gnd.n331 gnd.n327 0.152939
R13930 gnd.n332 gnd.n331 0.152939
R13931 gnd.n333 gnd.n332 0.152939
R13932 gnd.n334 gnd.n333 0.152939
R13933 gnd.n338 gnd.n334 0.152939
R13934 gnd.n339 gnd.n338 0.152939
R13935 gnd.n340 gnd.n339 0.152939
R13936 gnd.n341 gnd.n340 0.152939
R13937 gnd.n345 gnd.n341 0.152939
R13938 gnd.n346 gnd.n345 0.152939
R13939 gnd.n7392 gnd.n346 0.152939
R13940 gnd.n7392 gnd.n7391 0.152939
R13941 gnd.n7533 gnd.n215 0.152939
R13942 gnd.n217 gnd.n215 0.152939
R13943 gnd.n221 gnd.n217 0.152939
R13944 gnd.n222 gnd.n221 0.152939
R13945 gnd.n223 gnd.n222 0.152939
R13946 gnd.n224 gnd.n223 0.152939
R13947 gnd.n228 gnd.n224 0.152939
R13948 gnd.n229 gnd.n228 0.152939
R13949 gnd.n230 gnd.n229 0.152939
R13950 gnd.n231 gnd.n230 0.152939
R13951 gnd.n235 gnd.n231 0.152939
R13952 gnd.n236 gnd.n235 0.152939
R13953 gnd.n237 gnd.n236 0.152939
R13954 gnd.n238 gnd.n237 0.152939
R13955 gnd.n242 gnd.n238 0.152939
R13956 gnd.n243 gnd.n242 0.152939
R13957 gnd.n244 gnd.n243 0.152939
R13958 gnd.n245 gnd.n244 0.152939
R13959 gnd.n249 gnd.n245 0.152939
R13960 gnd.n250 gnd.n249 0.152939
R13961 gnd.n251 gnd.n250 0.152939
R13962 gnd.n252 gnd.n251 0.152939
R13963 gnd.n256 gnd.n252 0.152939
R13964 gnd.n257 gnd.n256 0.152939
R13965 gnd.n258 gnd.n257 0.152939
R13966 gnd.n259 gnd.n258 0.152939
R13967 gnd.n263 gnd.n259 0.152939
R13968 gnd.n264 gnd.n263 0.152939
R13969 gnd.n265 gnd.n264 0.152939
R13970 gnd.n266 gnd.n265 0.152939
R13971 gnd.n270 gnd.n266 0.152939
R13972 gnd.n271 gnd.n270 0.152939
R13973 gnd.n272 gnd.n271 0.152939
R13974 gnd.n273 gnd.n272 0.152939
R13975 gnd.n277 gnd.n273 0.152939
R13976 gnd.n278 gnd.n277 0.152939
R13977 gnd.n7464 gnd.n278 0.152939
R13978 gnd.n7464 gnd.n7463 0.152939
R13979 gnd.n7463 gnd.n7462 0.152939
R13980 gnd.n7462 gnd.n282 0.152939
R13981 gnd.n288 gnd.n282 0.152939
R13982 gnd.n289 gnd.n288 0.152939
R13983 gnd.n290 gnd.n289 0.152939
R13984 gnd.n291 gnd.n290 0.152939
R13985 gnd.n295 gnd.n291 0.152939
R13986 gnd.n296 gnd.n295 0.152939
R13987 gnd.n297 gnd.n296 0.152939
R13988 gnd.n298 gnd.n297 0.152939
R13989 gnd.n302 gnd.n298 0.152939
R13990 gnd.n303 gnd.n302 0.152939
R13991 gnd.n304 gnd.n303 0.152939
R13992 gnd.n305 gnd.n304 0.152939
R13993 gnd.n309 gnd.n305 0.152939
R13994 gnd.n310 gnd.n309 0.152939
R13995 gnd.n311 gnd.n310 0.152939
R13996 gnd.n312 gnd.n311 0.152939
R13997 gnd.n317 gnd.n312 0.152939
R13998 gnd.n7425 gnd.n317 0.152939
R13999 gnd.n1410 gnd.n1409 0.152939
R14000 gnd.n1411 gnd.n1410 0.152939
R14001 gnd.n1412 gnd.n1411 0.152939
R14002 gnd.n1413 gnd.n1412 0.152939
R14003 gnd.n1414 gnd.n1413 0.152939
R14004 gnd.n1415 gnd.n1414 0.152939
R14005 gnd.n1416 gnd.n1415 0.152939
R14006 gnd.n1417 gnd.n1416 0.152939
R14007 gnd.n1418 gnd.n1417 0.152939
R14008 gnd.n1419 gnd.n1418 0.152939
R14009 gnd.n1420 gnd.n1419 0.152939
R14010 gnd.n1421 gnd.n1420 0.152939
R14011 gnd.n1422 gnd.n1421 0.152939
R14012 gnd.n1423 gnd.n1422 0.152939
R14013 gnd.n1424 gnd.n1423 0.152939
R14014 gnd.n1425 gnd.n1424 0.152939
R14015 gnd.n1426 gnd.n1425 0.152939
R14016 gnd.n1429 gnd.n1426 0.152939
R14017 gnd.n1430 gnd.n1429 0.152939
R14018 gnd.n1431 gnd.n1430 0.152939
R14019 gnd.n1432 gnd.n1431 0.152939
R14020 gnd.n1433 gnd.n1432 0.152939
R14021 gnd.n1434 gnd.n1433 0.152939
R14022 gnd.n1435 gnd.n1434 0.152939
R14023 gnd.n1436 gnd.n1435 0.152939
R14024 gnd.n1441 gnd.n1440 0.152939
R14025 gnd.n1442 gnd.n1441 0.152939
R14026 gnd.n1443 gnd.n1442 0.152939
R14027 gnd.n1444 gnd.n1443 0.152939
R14028 gnd.n1445 gnd.n1444 0.152939
R14029 gnd.n1446 gnd.n1445 0.152939
R14030 gnd.n1447 gnd.n1446 0.152939
R14031 gnd.n1448 gnd.n1447 0.152939
R14032 gnd.n1449 gnd.n1448 0.152939
R14033 gnd.n1452 gnd.n1449 0.152939
R14034 gnd.n1453 gnd.n1452 0.152939
R14035 gnd.n1454 gnd.n1453 0.152939
R14036 gnd.n1455 gnd.n1454 0.152939
R14037 gnd.n1456 gnd.n1455 0.152939
R14038 gnd.n1457 gnd.n1456 0.152939
R14039 gnd.n1458 gnd.n1457 0.152939
R14040 gnd.n1459 gnd.n1458 0.152939
R14041 gnd.n1460 gnd.n1459 0.152939
R14042 gnd.n1461 gnd.n1460 0.152939
R14043 gnd.n1462 gnd.n1461 0.152939
R14044 gnd.n1463 gnd.n1462 0.152939
R14045 gnd.n1464 gnd.n1463 0.152939
R14046 gnd.n1465 gnd.n1464 0.152939
R14047 gnd.n1466 gnd.n1465 0.152939
R14048 gnd.n1467 gnd.n1466 0.152939
R14049 gnd.n1468 gnd.n1467 0.152939
R14050 gnd.n1469 gnd.n1468 0.152939
R14051 gnd.n1470 gnd.n1469 0.152939
R14052 gnd.n5967 gnd.n1470 0.152939
R14053 gnd.n5967 gnd.n5966 0.152939
R14054 gnd.n1491 gnd.n1490 0.152939
R14055 gnd.n1492 gnd.n1491 0.152939
R14056 gnd.n1493 gnd.n1492 0.152939
R14057 gnd.n1494 gnd.n1493 0.152939
R14058 gnd.n1514 gnd.n1494 0.152939
R14059 gnd.n1515 gnd.n1514 0.152939
R14060 gnd.n1516 gnd.n1515 0.152939
R14061 gnd.n1517 gnd.n1516 0.152939
R14062 gnd.n1535 gnd.n1517 0.152939
R14063 gnd.n1536 gnd.n1535 0.152939
R14064 gnd.n1537 gnd.n1536 0.152939
R14065 gnd.n1538 gnd.n1537 0.152939
R14066 gnd.n1554 gnd.n1538 0.152939
R14067 gnd.n1555 gnd.n1554 0.152939
R14068 gnd.n1556 gnd.n1555 0.152939
R14069 gnd.n1557 gnd.n1556 0.152939
R14070 gnd.n1575 gnd.n1557 0.152939
R14071 gnd.n1576 gnd.n1575 0.152939
R14072 gnd.n1577 gnd.n1576 0.152939
R14073 gnd.n1578 gnd.n1577 0.152939
R14074 gnd.n1578 gnd.n97 0.152939
R14075 gnd.n5881 gnd.n1600 0.152939
R14076 gnd.n5882 gnd.n5881 0.152939
R14077 gnd.n5884 gnd.n5882 0.152939
R14078 gnd.n5884 gnd.n5883 0.152939
R14079 gnd.n7277 gnd.n390 0.152939
R14080 gnd.n4543 gnd.n4542 0.152939
R14081 gnd.n4546 gnd.n4543 0.152939
R14082 gnd.n4547 gnd.n4546 0.152939
R14083 gnd.n4548 gnd.n4547 0.152939
R14084 gnd.n4549 gnd.n4548 0.152939
R14085 gnd.n4551 gnd.n4549 0.152939
R14086 gnd.n4551 gnd.n4550 0.152939
R14087 gnd.n4550 gnd.n2399 0.152939
R14088 gnd.n4630 gnd.n2399 0.152939
R14089 gnd.n4631 gnd.n4630 0.152939
R14090 gnd.n4632 gnd.n4631 0.152939
R14091 gnd.n4632 gnd.n2395 0.152939
R14092 gnd.n4638 gnd.n2395 0.152939
R14093 gnd.n4639 gnd.n4638 0.152939
R14094 gnd.n4640 gnd.n4639 0.152939
R14095 gnd.n4641 gnd.n4640 0.152939
R14096 gnd.n4642 gnd.n4641 0.152939
R14097 gnd.n4645 gnd.n4642 0.152939
R14098 gnd.n4646 gnd.n4645 0.152939
R14099 gnd.n4647 gnd.n4646 0.152939
R14100 gnd.n4648 gnd.n4647 0.152939
R14101 gnd.n4652 gnd.n4648 0.152939
R14102 gnd.n4653 gnd.n4652 0.152939
R14103 gnd.n4654 gnd.n4653 0.152939
R14104 gnd.n4654 gnd.n2117 0.152939
R14105 gnd.n4777 gnd.n2117 0.152939
R14106 gnd.n4778 gnd.n4777 0.152939
R14107 gnd.n4779 gnd.n4778 0.152939
R14108 gnd.n4779 gnd.n2104 0.152939
R14109 gnd.n4793 gnd.n2104 0.152939
R14110 gnd.n4794 gnd.n4793 0.152939
R14111 gnd.n4795 gnd.n4794 0.152939
R14112 gnd.n4795 gnd.n2090 0.152939
R14113 gnd.n4809 gnd.n2090 0.152939
R14114 gnd.n4810 gnd.n4809 0.152939
R14115 gnd.n4811 gnd.n4810 0.152939
R14116 gnd.n4811 gnd.n2075 0.152939
R14117 gnd.n4825 gnd.n2075 0.152939
R14118 gnd.n4826 gnd.n4825 0.152939
R14119 gnd.n4827 gnd.n4826 0.152939
R14120 gnd.n4827 gnd.n2061 0.152939
R14121 gnd.n4841 gnd.n2061 0.152939
R14122 gnd.n4842 gnd.n4841 0.152939
R14123 gnd.n4843 gnd.n4842 0.152939
R14124 gnd.n4843 gnd.n2046 0.152939
R14125 gnd.n4871 gnd.n2046 0.152939
R14126 gnd.n4872 gnd.n4871 0.152939
R14127 gnd.n4873 gnd.n4872 0.152939
R14128 gnd.n4874 gnd.n4873 0.152939
R14129 gnd.n4876 gnd.n4874 0.152939
R14130 gnd.n4876 gnd.n4875 0.152939
R14131 gnd.n4875 gnd.n1190 0.152939
R14132 gnd.n1191 gnd.n1190 0.152939
R14133 gnd.n1192 gnd.n1191 0.152939
R14134 gnd.n5029 gnd.n1192 0.152939
R14135 gnd.n5030 gnd.n5029 0.152939
R14136 gnd.n5031 gnd.n5030 0.152939
R14137 gnd.n5031 gnd.n2016 0.152939
R14138 gnd.n5058 gnd.n2016 0.152939
R14139 gnd.n5059 gnd.n5058 0.152939
R14140 gnd.n5060 gnd.n5059 0.152939
R14141 gnd.n5061 gnd.n5060 0.152939
R14142 gnd.n5061 gnd.n1988 0.152939
R14143 gnd.n5096 gnd.n1988 0.152939
R14144 gnd.n5097 gnd.n5096 0.152939
R14145 gnd.n5098 gnd.n5097 0.152939
R14146 gnd.n5099 gnd.n5098 0.152939
R14147 gnd.n5101 gnd.n5099 0.152939
R14148 gnd.n5101 gnd.n5100 0.152939
R14149 gnd.n5100 gnd.n1962 0.152939
R14150 gnd.n1963 gnd.n1962 0.152939
R14151 gnd.n1964 gnd.n1963 0.152939
R14152 gnd.n1964 gnd.n1938 0.152939
R14153 gnd.n5197 gnd.n1938 0.152939
R14154 gnd.n5198 gnd.n5197 0.152939
R14155 gnd.n5199 gnd.n5198 0.152939
R14156 gnd.n5200 gnd.n5199 0.152939
R14157 gnd.n5200 gnd.n1910 0.152939
R14158 gnd.n5235 gnd.n1910 0.152939
R14159 gnd.n5236 gnd.n5235 0.152939
R14160 gnd.n5237 gnd.n5236 0.152939
R14161 gnd.n5237 gnd.n1884 0.152939
R14162 gnd.n5272 gnd.n1884 0.152939
R14163 gnd.n5273 gnd.n5272 0.152939
R14164 gnd.n5274 gnd.n5273 0.152939
R14165 gnd.n5275 gnd.n5274 0.152939
R14166 gnd.n5275 gnd.n1857 0.152939
R14167 gnd.n5321 gnd.n1857 0.152939
R14168 gnd.n5322 gnd.n5321 0.152939
R14169 gnd.n5323 gnd.n5322 0.152939
R14170 gnd.n5324 gnd.n5323 0.152939
R14171 gnd.n5324 gnd.n1835 0.152939
R14172 gnd.n5362 gnd.n1835 0.152939
R14173 gnd.n5363 gnd.n5362 0.152939
R14174 gnd.n5364 gnd.n5363 0.152939
R14175 gnd.n5365 gnd.n5364 0.152939
R14176 gnd.n5365 gnd.n1805 0.152939
R14177 gnd.n5402 gnd.n1805 0.152939
R14178 gnd.n5403 gnd.n5402 0.152939
R14179 gnd.n5404 gnd.n5403 0.152939
R14180 gnd.n5404 gnd.n1781 0.152939
R14181 gnd.n5445 gnd.n1781 0.152939
R14182 gnd.n5446 gnd.n5445 0.152939
R14183 gnd.n5447 gnd.n5446 0.152939
R14184 gnd.n5448 gnd.n5447 0.152939
R14185 gnd.n5448 gnd.n1725 0.152939
R14186 gnd.n5621 gnd.n1725 0.152939
R14187 gnd.n5622 gnd.n5621 0.152939
R14188 gnd.n5623 gnd.n5622 0.152939
R14189 gnd.n5623 gnd.n1714 0.152939
R14190 gnd.n5638 gnd.n1714 0.152939
R14191 gnd.n5639 gnd.n5638 0.152939
R14192 gnd.n5640 gnd.n5639 0.152939
R14193 gnd.n5640 gnd.n1702 0.152939
R14194 gnd.n5655 gnd.n1702 0.152939
R14195 gnd.n5656 gnd.n5655 0.152939
R14196 gnd.n5657 gnd.n5656 0.152939
R14197 gnd.n5657 gnd.n1690 0.152939
R14198 gnd.n5672 gnd.n1690 0.152939
R14199 gnd.n5673 gnd.n5672 0.152939
R14200 gnd.n5674 gnd.n5673 0.152939
R14201 gnd.n5674 gnd.n1678 0.152939
R14202 gnd.n5689 gnd.n1678 0.152939
R14203 gnd.n5690 gnd.n5689 0.152939
R14204 gnd.n5691 gnd.n5690 0.152939
R14205 gnd.n5693 gnd.n5691 0.152939
R14206 gnd.n5693 gnd.n5692 0.152939
R14207 gnd.n5692 gnd.n1666 0.152939
R14208 gnd.n5711 gnd.n1666 0.152939
R14209 gnd.n5712 gnd.n5711 0.152939
R14210 gnd.n5713 gnd.n5712 0.152939
R14211 gnd.n5714 gnd.n5713 0.152939
R14212 gnd.n5715 gnd.n5714 0.152939
R14213 gnd.n5717 gnd.n5715 0.152939
R14214 gnd.n5718 gnd.n5717 0.152939
R14215 gnd.n5718 gnd.n1630 0.152939
R14216 gnd.n5780 gnd.n1630 0.152939
R14217 gnd.n5781 gnd.n5780 0.152939
R14218 gnd.n5782 gnd.n5781 0.152939
R14219 gnd.n5782 gnd.n1626 0.152939
R14220 gnd.n5788 gnd.n1626 0.152939
R14221 gnd.n5789 gnd.n5788 0.152939
R14222 gnd.n5790 gnd.n5789 0.152939
R14223 gnd.n5790 gnd.n1622 0.152939
R14224 gnd.n5796 gnd.n1622 0.152939
R14225 gnd.n5797 gnd.n5796 0.152939
R14226 gnd.n5798 gnd.n5797 0.152939
R14227 gnd.n5799 gnd.n5798 0.152939
R14228 gnd.n5800 gnd.n5799 0.152939
R14229 gnd.n5803 gnd.n5800 0.152939
R14230 gnd.n5804 gnd.n5803 0.152939
R14231 gnd.n5805 gnd.n5804 0.152939
R14232 gnd.n5806 gnd.n5805 0.152939
R14233 gnd.n5808 gnd.n5806 0.152939
R14234 gnd.n5808 gnd.n5807 0.152939
R14235 gnd.n5807 gnd.n1600 0.152939
R14236 gnd.n4199 gnd.n4165 0.152939
R14237 gnd.n4166 gnd.n4165 0.152939
R14238 gnd.n4167 gnd.n4166 0.152939
R14239 gnd.n4168 gnd.n4167 0.152939
R14240 gnd.n4169 gnd.n4168 0.152939
R14241 gnd.n4170 gnd.n4169 0.152939
R14242 gnd.n4171 gnd.n4170 0.152939
R14243 gnd.n4172 gnd.n4171 0.152939
R14244 gnd.n4173 gnd.n4172 0.152939
R14245 gnd.n4174 gnd.n4173 0.152939
R14246 gnd.n4175 gnd.n4174 0.152939
R14247 gnd.n4176 gnd.n4175 0.152939
R14248 gnd.n4177 gnd.n4176 0.152939
R14249 gnd.n4177 gnd.n2485 0.152939
R14250 gnd.n4444 gnd.n2485 0.152939
R14251 gnd.n4445 gnd.n4444 0.152939
R14252 gnd.n4446 gnd.n4445 0.152939
R14253 gnd.n4447 gnd.n4446 0.152939
R14254 gnd.n4448 gnd.n4447 0.152939
R14255 gnd.n4449 gnd.n4448 0.152939
R14256 gnd.n4450 gnd.n4449 0.152939
R14257 gnd.n4451 gnd.n4450 0.152939
R14258 gnd.n4451 gnd.n2449 0.152939
R14259 gnd.n4505 gnd.n2449 0.152939
R14260 gnd.n4506 gnd.n4505 0.152939
R14261 gnd.n4507 gnd.n4506 0.152939
R14262 gnd.n4238 gnd.n4146 0.152939
R14263 gnd.n4147 gnd.n4146 0.152939
R14264 gnd.n4148 gnd.n4147 0.152939
R14265 gnd.n4149 gnd.n4148 0.152939
R14266 gnd.n4150 gnd.n4149 0.152939
R14267 gnd.n4151 gnd.n4150 0.152939
R14268 gnd.n4152 gnd.n4151 0.152939
R14269 gnd.n4153 gnd.n4152 0.152939
R14270 gnd.n4154 gnd.n4153 0.152939
R14271 gnd.n4155 gnd.n4154 0.152939
R14272 gnd.n4156 gnd.n4155 0.152939
R14273 gnd.n4157 gnd.n4156 0.152939
R14274 gnd.n4158 gnd.n4157 0.152939
R14275 gnd.n4159 gnd.n4158 0.152939
R14276 gnd.n4160 gnd.n4159 0.152939
R14277 gnd.n4203 gnd.n4160 0.152939
R14278 gnd.n4203 gnd.n4202 0.152939
R14279 gnd.n4202 gnd.n4201 0.152939
R14280 gnd.n971 gnd.n946 0.152939
R14281 gnd.n972 gnd.n971 0.152939
R14282 gnd.n973 gnd.n972 0.152939
R14283 gnd.n991 gnd.n973 0.152939
R14284 gnd.n992 gnd.n991 0.152939
R14285 gnd.n993 gnd.n992 0.152939
R14286 gnd.n994 gnd.n993 0.152939
R14287 gnd.n1010 gnd.n994 0.152939
R14288 gnd.n1011 gnd.n1010 0.152939
R14289 gnd.n1012 gnd.n1011 0.152939
R14290 gnd.n1013 gnd.n1012 0.152939
R14291 gnd.n1031 gnd.n1013 0.152939
R14292 gnd.n1032 gnd.n1031 0.152939
R14293 gnd.n1033 gnd.n1032 0.152939
R14294 gnd.n1034 gnd.n1033 0.152939
R14295 gnd.n1051 gnd.n1034 0.152939
R14296 gnd.n1052 gnd.n1051 0.152939
R14297 gnd.n1053 gnd.n1052 0.152939
R14298 gnd.n1054 gnd.n1053 0.152939
R14299 gnd.n1070 gnd.n1054 0.152939
R14300 gnd.n6395 gnd.n1070 0.152939
R14301 gnd.n6394 gnd.n1071 0.152939
R14302 gnd.n1076 gnd.n1071 0.152939
R14303 gnd.n1077 gnd.n1076 0.152939
R14304 gnd.n1078 gnd.n1077 0.152939
R14305 gnd.n1079 gnd.n1078 0.152939
R14306 gnd.n1080 gnd.n1079 0.152939
R14307 gnd.n1084 gnd.n1080 0.152939
R14308 gnd.n1085 gnd.n1084 0.152939
R14309 gnd.n1086 gnd.n1085 0.152939
R14310 gnd.n1087 gnd.n1086 0.152939
R14311 gnd.n1091 gnd.n1087 0.152939
R14312 gnd.n1092 gnd.n1091 0.152939
R14313 gnd.n1093 gnd.n1092 0.152939
R14314 gnd.n1094 gnd.n1093 0.152939
R14315 gnd.n1098 gnd.n1094 0.152939
R14316 gnd.n1099 gnd.n1098 0.152939
R14317 gnd.n1100 gnd.n1099 0.152939
R14318 gnd.n1103 gnd.n1100 0.152939
R14319 gnd.n1107 gnd.n1103 0.152939
R14320 gnd.n1108 gnd.n1107 0.152939
R14321 gnd.n1109 gnd.n1108 0.152939
R14322 gnd.n1110 gnd.n1109 0.152939
R14323 gnd.n1114 gnd.n1110 0.152939
R14324 gnd.n1115 gnd.n1114 0.152939
R14325 gnd.n1116 gnd.n1115 0.152939
R14326 gnd.n2226 gnd.n2225 0.152939
R14327 gnd.n2235 gnd.n2226 0.152939
R14328 gnd.n2236 gnd.n2235 0.152939
R14329 gnd.n2237 gnd.n2236 0.152939
R14330 gnd.n2237 gnd.n2221 0.152939
R14331 gnd.n2245 gnd.n2221 0.152939
R14332 gnd.n2246 gnd.n2245 0.152939
R14333 gnd.n2247 gnd.n2246 0.152939
R14334 gnd.n2247 gnd.n2215 0.152939
R14335 gnd.n2255 gnd.n2215 0.152939
R14336 gnd.n2256 gnd.n2255 0.152939
R14337 gnd.n2257 gnd.n2256 0.152939
R14338 gnd.n2257 gnd.n2211 0.152939
R14339 gnd.n2265 gnd.n2211 0.152939
R14340 gnd.n2266 gnd.n2265 0.152939
R14341 gnd.n2267 gnd.n2266 0.152939
R14342 gnd.n2267 gnd.n2207 0.152939
R14343 gnd.n2275 gnd.n2207 0.152939
R14344 gnd.n2276 gnd.n2275 0.152939
R14345 gnd.n2277 gnd.n2276 0.152939
R14346 gnd.n2277 gnd.n2203 0.152939
R14347 gnd.n2285 gnd.n2203 0.152939
R14348 gnd.n2286 gnd.n2285 0.152939
R14349 gnd.n2287 gnd.n2286 0.152939
R14350 gnd.n2287 gnd.n2199 0.152939
R14351 gnd.n2295 gnd.n2199 0.152939
R14352 gnd.n2296 gnd.n2295 0.152939
R14353 gnd.n2297 gnd.n2296 0.152939
R14354 gnd.n2297 gnd.n2193 0.152939
R14355 gnd.n2304 gnd.n2193 0.152939
R14356 gnd.n4084 gnd.n4083 0.152939
R14357 gnd.n4085 gnd.n4084 0.152939
R14358 gnd.n4086 gnd.n4085 0.152939
R14359 gnd.n4087 gnd.n4086 0.152939
R14360 gnd.n4088 gnd.n4087 0.152939
R14361 gnd.n4089 gnd.n4088 0.152939
R14362 gnd.n4090 gnd.n4089 0.152939
R14363 gnd.n4091 gnd.n4090 0.152939
R14364 gnd.n4092 gnd.n4091 0.152939
R14365 gnd.n4093 gnd.n4092 0.152939
R14366 gnd.n4094 gnd.n4093 0.152939
R14367 gnd.n4095 gnd.n4094 0.152939
R14368 gnd.n4096 gnd.n4095 0.152939
R14369 gnd.n4097 gnd.n4096 0.152939
R14370 gnd.n4098 gnd.n4097 0.152939
R14371 gnd.n4099 gnd.n4098 0.152939
R14372 gnd.n4100 gnd.n4099 0.152939
R14373 gnd.n4103 gnd.n4100 0.152939
R14374 gnd.n4104 gnd.n4103 0.152939
R14375 gnd.n4105 gnd.n4104 0.152939
R14376 gnd.n4106 gnd.n4105 0.152939
R14377 gnd.n4107 gnd.n4106 0.152939
R14378 gnd.n4108 gnd.n4107 0.152939
R14379 gnd.n4109 gnd.n4108 0.152939
R14380 gnd.n4110 gnd.n4109 0.152939
R14381 gnd.n4111 gnd.n4110 0.152939
R14382 gnd.n4112 gnd.n4111 0.152939
R14383 gnd.n4113 gnd.n4112 0.152939
R14384 gnd.n4114 gnd.n4113 0.152939
R14385 gnd.n4115 gnd.n4114 0.152939
R14386 gnd.n4116 gnd.n4115 0.152939
R14387 gnd.n4117 gnd.n4116 0.152939
R14388 gnd.n4118 gnd.n4117 0.152939
R14389 gnd.n4119 gnd.n4118 0.152939
R14390 gnd.n4120 gnd.n4119 0.152939
R14391 gnd.n4121 gnd.n4120 0.152939
R14392 gnd.n4122 gnd.n4121 0.152939
R14393 gnd.n4125 gnd.n4122 0.152939
R14394 gnd.n4126 gnd.n4125 0.152939
R14395 gnd.n4127 gnd.n4126 0.152939
R14396 gnd.n4128 gnd.n4127 0.152939
R14397 gnd.n4129 gnd.n4128 0.152939
R14398 gnd.n4130 gnd.n4129 0.152939
R14399 gnd.n4131 gnd.n4130 0.152939
R14400 gnd.n4132 gnd.n4131 0.152939
R14401 gnd.n4133 gnd.n4132 0.152939
R14402 gnd.n4134 gnd.n4133 0.152939
R14403 gnd.n4135 gnd.n4134 0.152939
R14404 gnd.n4136 gnd.n4135 0.152939
R14405 gnd.n4137 gnd.n4136 0.152939
R14406 gnd.n4138 gnd.n4137 0.152939
R14407 gnd.n4139 gnd.n4138 0.152939
R14408 gnd.n4140 gnd.n4139 0.152939
R14409 gnd.n4141 gnd.n4140 0.152939
R14410 gnd.n4142 gnd.n4141 0.152939
R14411 gnd.n4143 gnd.n4142 0.152939
R14412 gnd.n4241 gnd.n4143 0.152939
R14413 gnd.n4241 gnd.n4240 0.152939
R14414 gnd.n4370 gnd.n2549 0.152939
R14415 gnd.n4371 gnd.n4370 0.152939
R14416 gnd.n4372 gnd.n4371 0.152939
R14417 gnd.n4372 gnd.n2530 0.152939
R14418 gnd.n4390 gnd.n2530 0.152939
R14419 gnd.n4391 gnd.n4390 0.152939
R14420 gnd.n4392 gnd.n4391 0.152939
R14421 gnd.n4392 gnd.n2513 0.152939
R14422 gnd.n4410 gnd.n2513 0.152939
R14423 gnd.n4411 gnd.n4410 0.152939
R14424 gnd.n4412 gnd.n4411 0.152939
R14425 gnd.n4412 gnd.n2493 0.152939
R14426 gnd.n4434 gnd.n2493 0.152939
R14427 gnd.n4435 gnd.n4434 0.152939
R14428 gnd.n4436 gnd.n4435 0.152939
R14429 gnd.n4437 gnd.n4436 0.152939
R14430 gnd.n4437 gnd.n2469 0.152939
R14431 gnd.n4475 gnd.n2469 0.152939
R14432 gnd.n4476 gnd.n4475 0.152939
R14433 gnd.n4477 gnd.n4476 0.152939
R14434 gnd.n4477 gnd.n947 0.152939
R14435 gnd.n2429 gnd.n2428 0.152939
R14436 gnd.n4540 gnd.n4539 0.152939
R14437 gnd.n4541 gnd.n4540 0.152939
R14438 gnd.n4542 gnd.n4541 0.152939
R14439 gnd.n6643 gnd.n769 0.152939
R14440 gnd.n774 gnd.n769 0.152939
R14441 gnd.n775 gnd.n774 0.152939
R14442 gnd.n776 gnd.n775 0.152939
R14443 gnd.n781 gnd.n776 0.152939
R14444 gnd.n782 gnd.n781 0.152939
R14445 gnd.n783 gnd.n782 0.152939
R14446 gnd.n784 gnd.n783 0.152939
R14447 gnd.n789 gnd.n784 0.152939
R14448 gnd.n790 gnd.n789 0.152939
R14449 gnd.n791 gnd.n790 0.152939
R14450 gnd.n792 gnd.n791 0.152939
R14451 gnd.n797 gnd.n792 0.152939
R14452 gnd.n798 gnd.n797 0.152939
R14453 gnd.n799 gnd.n798 0.152939
R14454 gnd.n800 gnd.n799 0.152939
R14455 gnd.n805 gnd.n800 0.152939
R14456 gnd.n806 gnd.n805 0.152939
R14457 gnd.n807 gnd.n806 0.152939
R14458 gnd.n808 gnd.n807 0.152939
R14459 gnd.n813 gnd.n808 0.152939
R14460 gnd.n814 gnd.n813 0.152939
R14461 gnd.n815 gnd.n814 0.152939
R14462 gnd.n816 gnd.n815 0.152939
R14463 gnd.n821 gnd.n816 0.152939
R14464 gnd.n822 gnd.n821 0.152939
R14465 gnd.n823 gnd.n822 0.152939
R14466 gnd.n824 gnd.n823 0.152939
R14467 gnd.n829 gnd.n824 0.152939
R14468 gnd.n830 gnd.n829 0.152939
R14469 gnd.n831 gnd.n830 0.152939
R14470 gnd.n832 gnd.n831 0.152939
R14471 gnd.n837 gnd.n832 0.152939
R14472 gnd.n838 gnd.n837 0.152939
R14473 gnd.n839 gnd.n838 0.152939
R14474 gnd.n840 gnd.n839 0.152939
R14475 gnd.n845 gnd.n840 0.152939
R14476 gnd.n846 gnd.n845 0.152939
R14477 gnd.n847 gnd.n846 0.152939
R14478 gnd.n848 gnd.n847 0.152939
R14479 gnd.n853 gnd.n848 0.152939
R14480 gnd.n854 gnd.n853 0.152939
R14481 gnd.n855 gnd.n854 0.152939
R14482 gnd.n856 gnd.n855 0.152939
R14483 gnd.n861 gnd.n856 0.152939
R14484 gnd.n862 gnd.n861 0.152939
R14485 gnd.n863 gnd.n862 0.152939
R14486 gnd.n864 gnd.n863 0.152939
R14487 gnd.n869 gnd.n864 0.152939
R14488 gnd.n870 gnd.n869 0.152939
R14489 gnd.n871 gnd.n870 0.152939
R14490 gnd.n872 gnd.n871 0.152939
R14491 gnd.n877 gnd.n872 0.152939
R14492 gnd.n878 gnd.n877 0.152939
R14493 gnd.n879 gnd.n878 0.152939
R14494 gnd.n880 gnd.n879 0.152939
R14495 gnd.n885 gnd.n880 0.152939
R14496 gnd.n886 gnd.n885 0.152939
R14497 gnd.n887 gnd.n886 0.152939
R14498 gnd.n888 gnd.n887 0.152939
R14499 gnd.n893 gnd.n888 0.152939
R14500 gnd.n894 gnd.n893 0.152939
R14501 gnd.n895 gnd.n894 0.152939
R14502 gnd.n896 gnd.n895 0.152939
R14503 gnd.n901 gnd.n896 0.152939
R14504 gnd.n902 gnd.n901 0.152939
R14505 gnd.n903 gnd.n902 0.152939
R14506 gnd.n904 gnd.n903 0.152939
R14507 gnd.n909 gnd.n904 0.152939
R14508 gnd.n910 gnd.n909 0.152939
R14509 gnd.n911 gnd.n910 0.152939
R14510 gnd.n912 gnd.n911 0.152939
R14511 gnd.n917 gnd.n912 0.152939
R14512 gnd.n918 gnd.n917 0.152939
R14513 gnd.n919 gnd.n918 0.152939
R14514 gnd.n920 gnd.n919 0.152939
R14515 gnd.n925 gnd.n920 0.152939
R14516 gnd.n926 gnd.n925 0.152939
R14517 gnd.n927 gnd.n926 0.152939
R14518 gnd.n928 gnd.n927 0.152939
R14519 gnd.n933 gnd.n928 0.152939
R14520 gnd.n934 gnd.n933 0.152939
R14521 gnd.n935 gnd.n934 0.152939
R14522 gnd.n936 gnd.n935 0.152939
R14523 gnd.n4786 gnd.n4785 0.152939
R14524 gnd.n4787 gnd.n4786 0.152939
R14525 gnd.n4787 gnd.n2097 0.152939
R14526 gnd.n4801 gnd.n2097 0.152939
R14527 gnd.n4802 gnd.n4801 0.152939
R14528 gnd.n4803 gnd.n4802 0.152939
R14529 gnd.n4803 gnd.n2083 0.152939
R14530 gnd.n4817 gnd.n2083 0.152939
R14531 gnd.n4818 gnd.n4817 0.152939
R14532 gnd.n4819 gnd.n4818 0.152939
R14533 gnd.n4819 gnd.n2069 0.152939
R14534 gnd.n4833 gnd.n2069 0.152939
R14535 gnd.n4834 gnd.n4833 0.152939
R14536 gnd.n4835 gnd.n4834 0.152939
R14537 gnd.n4835 gnd.n2055 0.152939
R14538 gnd.n4849 gnd.n2055 0.152939
R14539 gnd.n4850 gnd.n4849 0.152939
R14540 gnd.n4865 gnd.n4850 0.152939
R14541 gnd.n4865 gnd.n4864 0.152939
R14542 gnd.n4864 gnd.n4863 0.152939
R14543 gnd.n4863 gnd.n4851 0.152939
R14544 gnd.n4859 gnd.n4851 0.152939
R14545 gnd.n4859 gnd.n4858 0.152939
R14546 gnd.n4858 gnd.n4857 0.152939
R14547 gnd.n4857 gnd.n1200 0.152939
R14548 gnd.n6263 gnd.n1200 0.152939
R14549 gnd.n6263 gnd.n6262 0.152939
R14550 gnd.n6262 gnd.n6261 0.152939
R14551 gnd.n6261 gnd.n1201 0.152939
R14552 gnd.n6257 gnd.n1201 0.152939
R14553 gnd.n6257 gnd.n6256 0.152939
R14554 gnd.n6256 gnd.n6255 0.152939
R14555 gnd.n6255 gnd.n1206 0.152939
R14556 gnd.n6251 gnd.n1206 0.152939
R14557 gnd.n6251 gnd.n6250 0.152939
R14558 gnd.n6250 gnd.n6249 0.152939
R14559 gnd.n6249 gnd.n1211 0.152939
R14560 gnd.n6245 gnd.n1211 0.152939
R14561 gnd.n6245 gnd.n6244 0.152939
R14562 gnd.n6244 gnd.n6243 0.152939
R14563 gnd.n6243 gnd.n1216 0.152939
R14564 gnd.n6239 gnd.n1216 0.152939
R14565 gnd.n6239 gnd.n6238 0.152939
R14566 gnd.n6238 gnd.n6237 0.152939
R14567 gnd.n6237 gnd.n1221 0.152939
R14568 gnd.n6233 gnd.n1221 0.152939
R14569 gnd.n6233 gnd.n6232 0.152939
R14570 gnd.n6232 gnd.n6231 0.152939
R14571 gnd.n6231 gnd.n1226 0.152939
R14572 gnd.n6227 gnd.n1226 0.152939
R14573 gnd.n6227 gnd.n6226 0.152939
R14574 gnd.n6226 gnd.n6225 0.152939
R14575 gnd.n6225 gnd.n1231 0.152939
R14576 gnd.n6221 gnd.n1231 0.152939
R14577 gnd.n6221 gnd.n6220 0.152939
R14578 gnd.n6220 gnd.n6219 0.152939
R14579 gnd.n6219 gnd.n1236 0.152939
R14580 gnd.n6215 gnd.n1236 0.152939
R14581 gnd.n6215 gnd.n6214 0.152939
R14582 gnd.n6214 gnd.n6213 0.152939
R14583 gnd.n6213 gnd.n1241 0.152939
R14584 gnd.n6209 gnd.n1241 0.152939
R14585 gnd.n6209 gnd.n6208 0.152939
R14586 gnd.n6208 gnd.n6207 0.152939
R14587 gnd.n6207 gnd.n1246 0.152939
R14588 gnd.n6203 gnd.n1246 0.152939
R14589 gnd.n6203 gnd.n6202 0.152939
R14590 gnd.n6202 gnd.n6201 0.152939
R14591 gnd.n6201 gnd.n1251 0.152939
R14592 gnd.n6197 gnd.n1251 0.152939
R14593 gnd.n6197 gnd.n6196 0.152939
R14594 gnd.n6196 gnd.n6195 0.152939
R14595 gnd.n6195 gnd.n1256 0.152939
R14596 gnd.n6191 gnd.n1256 0.152939
R14597 gnd.n6191 gnd.n6190 0.152939
R14598 gnd.n6190 gnd.n6189 0.152939
R14599 gnd.n6189 gnd.n1261 0.152939
R14600 gnd.n6185 gnd.n1261 0.152939
R14601 gnd.n6185 gnd.n6184 0.152939
R14602 gnd.n6184 gnd.n6183 0.152939
R14603 gnd.n6183 gnd.n1266 0.152939
R14604 gnd.n6179 gnd.n1266 0.152939
R14605 gnd.n6179 gnd.n6178 0.152939
R14606 gnd.n6178 gnd.n6177 0.152939
R14607 gnd.n6177 gnd.n1271 0.152939
R14608 gnd.n6173 gnd.n1271 0.152939
R14609 gnd.n6173 gnd.n6172 0.152939
R14610 gnd.n6172 gnd.n6171 0.152939
R14611 gnd.n6171 gnd.n1276 0.152939
R14612 gnd.n6167 gnd.n1276 0.152939
R14613 gnd.n6167 gnd.n6166 0.152939
R14614 gnd.n6166 gnd.n6165 0.152939
R14615 gnd.n6165 gnd.n1281 0.152939
R14616 gnd.n6161 gnd.n1281 0.152939
R14617 gnd.n6161 gnd.n6160 0.152939
R14618 gnd.n6160 gnd.n6159 0.152939
R14619 gnd.n6159 gnd.n1286 0.152939
R14620 gnd.n6155 gnd.n1286 0.152939
R14621 gnd.n6155 gnd.n6154 0.152939
R14622 gnd.n6154 gnd.n6153 0.152939
R14623 gnd.n6153 gnd.n1291 0.152939
R14624 gnd.n4512 gnd.n4511 0.152939
R14625 gnd.n4511 gnd.n2419 0.152939
R14626 gnd.n4568 gnd.n2419 0.152939
R14627 gnd.n4569 gnd.n4568 0.152939
R14628 gnd.n4570 gnd.n4569 0.152939
R14629 gnd.n4570 gnd.n2414 0.152939
R14630 gnd.n4583 gnd.n2414 0.152939
R14631 gnd.n4584 gnd.n4583 0.152939
R14632 gnd.n4585 gnd.n4584 0.152939
R14633 gnd.n4585 gnd.n2406 0.152939
R14634 gnd.n4621 gnd.n2406 0.152939
R14635 gnd.n4621 gnd.n4620 0.152939
R14636 gnd.n4620 gnd.n4619 0.152939
R14637 gnd.n4619 gnd.n2407 0.152939
R14638 gnd.n4615 gnd.n2407 0.152939
R14639 gnd.n4615 gnd.n4614 0.152939
R14640 gnd.n4614 gnd.n4613 0.152939
R14641 gnd.n4613 gnd.n2411 0.152939
R14642 gnd.n4609 gnd.n2411 0.152939
R14643 gnd.n4609 gnd.n2387 0.152939
R14644 gnd.n4681 gnd.n2387 0.152939
R14645 gnd.n4682 gnd.n4681 0.152939
R14646 gnd.n4684 gnd.n4682 0.152939
R14647 gnd.n4684 gnd.n4683 0.152939
R14648 gnd.n4683 gnd.n2381 0.152939
R14649 gnd.n4698 gnd.n2381 0.152939
R14650 gnd.n4768 gnd.n2186 0.152939
R14651 gnd.n4768 gnd.n4767 0.152939
R14652 gnd.n4767 gnd.n4766 0.152939
R14653 gnd.n4766 gnd.n2188 0.152939
R14654 gnd.n4762 gnd.n2188 0.152939
R14655 gnd.n4762 gnd.n4761 0.152939
R14656 gnd.n2185 gnd.n2136 0.152939
R14657 gnd.n2181 gnd.n2136 0.152939
R14658 gnd.n2181 gnd.n2180 0.152939
R14659 gnd.n2180 gnd.n2179 0.152939
R14660 gnd.n2179 gnd.n2140 0.152939
R14661 gnd.n2175 gnd.n2140 0.152939
R14662 gnd.n2175 gnd.n2174 0.152939
R14663 gnd.n2174 gnd.n2173 0.152939
R14664 gnd.n2173 gnd.n2144 0.152939
R14665 gnd.n2169 gnd.n2144 0.152939
R14666 gnd.n2169 gnd.n2168 0.152939
R14667 gnd.n2168 gnd.n2167 0.152939
R14668 gnd.n2167 gnd.n2148 0.152939
R14669 gnd.n2163 gnd.n2148 0.152939
R14670 gnd.n2163 gnd.n2162 0.152939
R14671 gnd.n2162 gnd.n2161 0.152939
R14672 gnd.n2161 gnd.n2152 0.152939
R14673 gnd.n2157 gnd.n2152 0.152939
R14674 gnd.n2157 gnd.n2156 0.152939
R14675 gnd.n2156 gnd.n2155 0.152939
R14676 gnd.n2155 gnd.n2037 0.152939
R14677 gnd.n4888 gnd.n2037 0.152939
R14678 gnd.n4889 gnd.n4888 0.152939
R14679 gnd.n4890 gnd.n4889 0.152939
R14680 gnd.n4890 gnd.n2035 0.152939
R14681 gnd.n4994 gnd.n2035 0.152939
R14682 gnd.n4995 gnd.n4994 0.152939
R14683 gnd.n5023 gnd.n4995 0.152939
R14684 gnd.n5023 gnd.n5022 0.152939
R14685 gnd.n5022 gnd.n5021 0.152939
R14686 gnd.n5021 gnd.n4996 0.152939
R14687 gnd.n5017 gnd.n4996 0.152939
R14688 gnd.n5017 gnd.n5016 0.152939
R14689 gnd.n5016 gnd.n5015 0.152939
R14690 gnd.n5015 gnd.n4999 0.152939
R14691 gnd.n5011 gnd.n4999 0.152939
R14692 gnd.n5011 gnd.n5010 0.152939
R14693 gnd.n5010 gnd.n5009 0.152939
R14694 gnd.n5009 gnd.n5005 0.152939
R14695 gnd.n5005 gnd.n5004 0.152939
R14696 gnd.n5004 gnd.n1970 0.152939
R14697 gnd.n5131 gnd.n1970 0.152939
R14698 gnd.n5132 gnd.n5131 0.152939
R14699 gnd.n5159 gnd.n5132 0.152939
R14700 gnd.n5159 gnd.n5158 0.152939
R14701 gnd.n5158 gnd.n5157 0.152939
R14702 gnd.n5157 gnd.n5133 0.152939
R14703 gnd.n5153 gnd.n5133 0.152939
R14704 gnd.n5153 gnd.n5152 0.152939
R14705 gnd.n5152 gnd.n5151 0.152939
R14706 gnd.n5151 gnd.n5136 0.152939
R14707 gnd.n5147 gnd.n5136 0.152939
R14708 gnd.n5147 gnd.n5146 0.152939
R14709 gnd.n5146 gnd.n5145 0.152939
R14710 gnd.n5145 gnd.n5141 0.152939
R14711 gnd.n5141 gnd.n1877 0.152939
R14712 gnd.n5282 gnd.n1877 0.152939
R14713 gnd.n5283 gnd.n5282 0.152939
R14714 gnd.n5285 gnd.n5283 0.152939
R14715 gnd.n5285 gnd.n5284 0.152939
R14716 gnd.n5284 gnd.n1850 0.152939
R14717 gnd.n5331 gnd.n1850 0.152939
R14718 gnd.n5332 gnd.n5331 0.152939
R14719 gnd.n5349 gnd.n5332 0.152939
R14720 gnd.n5349 gnd.n5348 0.152939
R14721 gnd.n5348 gnd.n5347 0.152939
R14722 gnd.n5347 gnd.n5333 0.152939
R14723 gnd.n5343 gnd.n5333 0.152939
R14724 gnd.n5343 gnd.n5342 0.152939
R14725 gnd.n5342 gnd.n5341 0.152939
R14726 gnd.n5341 gnd.n5338 0.152939
R14727 gnd.n5338 gnd.n1798 0.152939
R14728 gnd.n5411 gnd.n1798 0.152939
R14729 gnd.n5412 gnd.n5411 0.152939
R14730 gnd.n5423 gnd.n5412 0.152939
R14731 gnd.n5423 gnd.n5422 0.152939
R14732 gnd.n5422 gnd.n5421 0.152939
R14733 gnd.n5421 gnd.n5413 0.152939
R14734 gnd.n5417 gnd.n5413 0.152939
R14735 gnd.n5417 gnd.n1720 0.152939
R14736 gnd.n5629 gnd.n1720 0.152939
R14737 gnd.n5630 gnd.n5629 0.152939
R14738 gnd.n5631 gnd.n5630 0.152939
R14739 gnd.n5631 gnd.n1708 0.152939
R14740 gnd.n5646 gnd.n1708 0.152939
R14741 gnd.n5647 gnd.n5646 0.152939
R14742 gnd.n5648 gnd.n5647 0.152939
R14743 gnd.n5648 gnd.n1696 0.152939
R14744 gnd.n5663 gnd.n1696 0.152939
R14745 gnd.n5664 gnd.n5663 0.152939
R14746 gnd.n5665 gnd.n5664 0.152939
R14747 gnd.n5665 gnd.n1683 0.152939
R14748 gnd.n5680 gnd.n1683 0.152939
R14749 gnd.n5681 gnd.n5680 0.152939
R14750 gnd.n5682 gnd.n5681 0.152939
R14751 gnd.n5682 gnd.n1672 0.152939
R14752 gnd.n5700 gnd.n1672 0.152939
R14753 gnd.n5701 gnd.n5700 0.152939
R14754 gnd.n5702 gnd.n5701 0.152939
R14755 gnd.n5702 gnd.n1300 0.152939
R14756 gnd.n6146 gnd.n1300 0.152939
R14757 gnd.n6145 gnd.n1301 0.152939
R14758 gnd.n6141 gnd.n1301 0.152939
R14759 gnd.n6141 gnd.n6140 0.152939
R14760 gnd.n6140 gnd.n6139 0.152939
R14761 gnd.n6139 gnd.n1305 0.152939
R14762 gnd.n6135 gnd.n1305 0.152939
R14763 gnd.n5773 gnd.n5735 0.152939
R14764 gnd.n5773 gnd.n5772 0.152939
R14765 gnd.n5772 gnd.n5771 0.152939
R14766 gnd.n5771 gnd.n5736 0.152939
R14767 gnd.n5767 gnd.n5736 0.152939
R14768 gnd.n5767 gnd.n5766 0.152939
R14769 gnd.n5766 gnd.n5765 0.152939
R14770 gnd.n5765 gnd.n5741 0.152939
R14771 gnd.n5761 gnd.n5741 0.152939
R14772 gnd.n5761 gnd.n1616 0.152939
R14773 gnd.n5825 gnd.n1616 0.152939
R14774 gnd.n5826 gnd.n5825 0.152939
R14775 gnd.n5827 gnd.n5826 0.152939
R14776 gnd.n5827 gnd.n1611 0.152939
R14777 gnd.n5840 gnd.n1611 0.152939
R14778 gnd.n5841 gnd.n5840 0.152939
R14779 gnd.n5842 gnd.n5841 0.152939
R14780 gnd.n5842 gnd.n1607 0.152939
R14781 gnd.n5872 gnd.n1607 0.152939
R14782 gnd.n5872 gnd.n5871 0.152939
R14783 gnd.n5871 gnd.n5870 0.152939
R14784 gnd.n5870 gnd.n1608 0.152939
R14785 gnd.n5866 gnd.n1608 0.152939
R14786 gnd.n5866 gnd.n5865 0.152939
R14787 gnd.n5865 gnd.n5864 0.152939
R14788 gnd.n5864 gnd.n83 0.152939
R14789 gnd.n4761 gnd.n4760 0.128549
R14790 gnd.n6135 gnd.n6134 0.128549
R14791 gnd.n5883 gnd.n98 0.098061
R14792 gnd.n4539 gnd.n948 0.098061
R14793 gnd.n3440 gnd.n3439 0.0767195
R14794 gnd.n3439 gnd.n3438 0.0767195
R14795 gnd.n7606 gnd.n96 0.0767195
R14796 gnd.n7606 gnd.n97 0.0767195
R14797 gnd.n6467 gnd.n946 0.0767195
R14798 gnd.n6467 gnd.n947 0.0767195
R14799 gnd.n7616 gnd.n7615 0.0695946
R14800 gnd.n4510 gnd.n4507 0.0695946
R14801 gnd.n4512 gnd.n4510 0.0695946
R14802 gnd.n7616 gnd.n83 0.0695946
R14803 gnd.n4760 gnd.n2305 0.063
R14804 gnd.n6134 gnd.n1310 0.063
R14805 gnd.n390 gnd.n98 0.055378
R14806 gnd.n2429 gnd.n948 0.055378
R14807 gnd.n4007 gnd.n2606 0.0477147
R14808 gnd.n1478 gnd.n1310 0.0477147
R14809 gnd.n7424 gnd.n207 0.0477147
R14810 gnd.n4239 gnd.n2559 0.0477147
R14811 gnd.n2305 gnd.n1063 0.0477147
R14812 gnd.n3203 gnd.n3091 0.0442063
R14813 gnd.n3204 gnd.n3203 0.0442063
R14814 gnd.n3205 gnd.n3204 0.0442063
R14815 gnd.n3205 gnd.n3080 0.0442063
R14816 gnd.n3219 gnd.n3080 0.0442063
R14817 gnd.n3220 gnd.n3219 0.0442063
R14818 gnd.n3221 gnd.n3220 0.0442063
R14819 gnd.n3221 gnd.n3067 0.0442063
R14820 gnd.n3265 gnd.n3067 0.0442063
R14821 gnd.n3266 gnd.n3265 0.0442063
R14822 gnd.n3268 gnd.n3001 0.0344674
R14823 gnd.n5956 gnd.n1478 0.0344674
R14824 gnd.n5956 gnd.n1480 0.0344674
R14825 gnd.n1504 gnd.n1480 0.0344674
R14826 gnd.n1505 gnd.n1504 0.0344674
R14827 gnd.n1506 gnd.n1505 0.0344674
R14828 gnd.n1507 gnd.n1506 0.0344674
R14829 gnd.n5748 gnd.n1507 0.0344674
R14830 gnd.n5748 gnd.n1525 0.0344674
R14831 gnd.n1526 gnd.n1525 0.0344674
R14832 gnd.n1527 gnd.n1526 0.0344674
R14833 gnd.n5754 gnd.n1527 0.0344674
R14834 gnd.n5754 gnd.n1545 0.0344674
R14835 gnd.n1546 gnd.n1545 0.0344674
R14836 gnd.n1547 gnd.n1546 0.0344674
R14837 gnd.n5834 gnd.n1547 0.0344674
R14838 gnd.n5834 gnd.n1565 0.0344674
R14839 gnd.n1566 gnd.n1565 0.0344674
R14840 gnd.n1567 gnd.n1566 0.0344674
R14841 gnd.n5849 gnd.n1567 0.0344674
R14842 gnd.n5849 gnd.n1585 0.0344674
R14843 gnd.n1586 gnd.n1585 0.0344674
R14844 gnd.n1587 gnd.n1586 0.0344674
R14845 gnd.n5852 gnd.n1587 0.0344674
R14846 gnd.n5852 gnd.n378 0.0344674
R14847 gnd.n7290 gnd.n378 0.0344674
R14848 gnd.n7291 gnd.n7290 0.0344674
R14849 gnd.n7291 gnd.n373 0.0344674
R14850 gnd.n373 gnd.n371 0.0344674
R14851 gnd.n7302 gnd.n371 0.0344674
R14852 gnd.n7303 gnd.n7302 0.0344674
R14853 gnd.n7303 gnd.n111 0.0344674
R14854 gnd.n112 gnd.n111 0.0344674
R14855 gnd.n113 gnd.n112 0.0344674
R14856 gnd.n7304 gnd.n113 0.0344674
R14857 gnd.n7304 gnd.n128 0.0344674
R14858 gnd.n129 gnd.n128 0.0344674
R14859 gnd.n130 gnd.n129 0.0344674
R14860 gnd.n7305 gnd.n130 0.0344674
R14861 gnd.n7305 gnd.n148 0.0344674
R14862 gnd.n149 gnd.n148 0.0344674
R14863 gnd.n150 gnd.n149 0.0344674
R14864 gnd.n7306 gnd.n150 0.0344674
R14865 gnd.n7306 gnd.n166 0.0344674
R14866 gnd.n167 gnd.n166 0.0344674
R14867 gnd.n168 gnd.n167 0.0344674
R14868 gnd.n7307 gnd.n168 0.0344674
R14869 gnd.n7307 gnd.n186 0.0344674
R14870 gnd.n187 gnd.n186 0.0344674
R14871 gnd.n188 gnd.n187 0.0344674
R14872 gnd.n7308 gnd.n188 0.0344674
R14873 gnd.n7308 gnd.n205 0.0344674
R14874 gnd.n206 gnd.n205 0.0344674
R14875 gnd.n207 gnd.n206 0.0344674
R14876 gnd.n4364 gnd.n2559 0.0344674
R14877 gnd.n4364 gnd.n2562 0.0344674
R14878 gnd.n2562 gnd.n2561 0.0344674
R14879 gnd.n2561 gnd.n2542 0.0344674
R14880 gnd.n2542 gnd.n2540 0.0344674
R14881 gnd.n4381 gnd.n2540 0.0344674
R14882 gnd.n4382 gnd.n4381 0.0344674
R14883 gnd.n4382 gnd.n2524 0.0344674
R14884 gnd.n2524 gnd.n2522 0.0344674
R14885 gnd.n4401 gnd.n2522 0.0344674
R14886 gnd.n4402 gnd.n4401 0.0344674
R14887 gnd.n4402 gnd.n2506 0.0344674
R14888 gnd.n2506 gnd.n2503 0.0344674
R14889 gnd.n2504 gnd.n2503 0.0344674
R14890 gnd.n4423 gnd.n2504 0.0344674
R14891 gnd.n4424 gnd.n4423 0.0344674
R14892 gnd.n4424 gnd.n2480 0.0344674
R14893 gnd.n2480 gnd.n2478 0.0344674
R14894 gnd.n4466 gnd.n2478 0.0344674
R14895 gnd.n4467 gnd.n4466 0.0344674
R14896 gnd.n4467 gnd.n2463 0.0344674
R14897 gnd.n2463 gnd.n2460 0.0344674
R14898 gnd.n2461 gnd.n2460 0.0344674
R14899 gnd.n4489 gnd.n2461 0.0344674
R14900 gnd.n4490 gnd.n4489 0.0344674
R14901 gnd.n4490 gnd.n2447 0.0344674
R14902 gnd.n2447 gnd.n2443 0.0344674
R14903 gnd.n2444 gnd.n2443 0.0344674
R14904 gnd.n4524 gnd.n2444 0.0344674
R14905 gnd.n4524 gnd.n2445 0.0344674
R14906 gnd.n2445 gnd.n962 0.0344674
R14907 gnd.n963 gnd.n962 0.0344674
R14908 gnd.n964 gnd.n963 0.0344674
R14909 gnd.n4577 gnd.n964 0.0344674
R14910 gnd.n4577 gnd.n981 0.0344674
R14911 gnd.n982 gnd.n981 0.0344674
R14912 gnd.n983 gnd.n982 0.0344674
R14913 gnd.n4592 gnd.n983 0.0344674
R14914 gnd.n4592 gnd.n1001 0.0344674
R14915 gnd.n1002 gnd.n1001 0.0344674
R14916 gnd.n1003 gnd.n1002 0.0344674
R14917 gnd.n4599 gnd.n1003 0.0344674
R14918 gnd.n4599 gnd.n1021 0.0344674
R14919 gnd.n1022 gnd.n1021 0.0344674
R14920 gnd.n1023 gnd.n1022 0.0344674
R14921 gnd.n2390 gnd.n1023 0.0344674
R14922 gnd.n2390 gnd.n1041 0.0344674
R14923 gnd.n1042 gnd.n1041 0.0344674
R14924 gnd.n1043 gnd.n1042 0.0344674
R14925 gnd.n2385 gnd.n1043 0.0344674
R14926 gnd.n2385 gnd.n1061 0.0344674
R14927 gnd.n1062 gnd.n1061 0.0344674
R14928 gnd.n1063 gnd.n1062 0.0344674
R14929 gnd.n4759 gnd.n2306 0.0343753
R14930 gnd.n6133 gnd.n6132 0.0343753
R14931 gnd.n4707 gnd.n4699 0.0296328
R14932 gnd.n5734 gnd.n5733 0.0296328
R14933 gnd.n3288 gnd.n3287 0.0269946
R14934 gnd.n3290 gnd.n3289 0.0269946
R14935 gnd.n2996 gnd.n2994 0.0269946
R14936 gnd.n3300 gnd.n3298 0.0269946
R14937 gnd.n3299 gnd.n2975 0.0269946
R14938 gnd.n3319 gnd.n3318 0.0269946
R14939 gnd.n3321 gnd.n3320 0.0269946
R14940 gnd.n2970 gnd.n2969 0.0269946
R14941 gnd.n3331 gnd.n2965 0.0269946
R14942 gnd.n3330 gnd.n2967 0.0269946
R14943 gnd.n2966 gnd.n2948 0.0269946
R14944 gnd.n3351 gnd.n2949 0.0269946
R14945 gnd.n3350 gnd.n2950 0.0269946
R14946 gnd.n3384 gnd.n2925 0.0269946
R14947 gnd.n3386 gnd.n3385 0.0269946
R14948 gnd.n3387 gnd.n2872 0.0269946
R14949 gnd.n2920 gnd.n2873 0.0269946
R14950 gnd.n2922 gnd.n2874 0.0269946
R14951 gnd.n3397 gnd.n3396 0.0269946
R14952 gnd.n3399 gnd.n3398 0.0269946
R14953 gnd.n3400 gnd.n2894 0.0269946
R14954 gnd.n3402 gnd.n2895 0.0269946
R14955 gnd.n3405 gnd.n2896 0.0269946
R14956 gnd.n3408 gnd.n3407 0.0269946
R14957 gnd.n3410 gnd.n3409 0.0269946
R14958 gnd.n3475 gnd.n2779 0.0269946
R14959 gnd.n3477 gnd.n3476 0.0269946
R14960 gnd.n3486 gnd.n2772 0.0269946
R14961 gnd.n3488 gnd.n3487 0.0269946
R14962 gnd.n3489 gnd.n2770 0.0269946
R14963 gnd.n3496 gnd.n3492 0.0269946
R14964 gnd.n3495 gnd.n3494 0.0269946
R14965 gnd.n3493 gnd.n2749 0.0269946
R14966 gnd.n3518 gnd.n2750 0.0269946
R14967 gnd.n3517 gnd.n2751 0.0269946
R14968 gnd.n3560 gnd.n2724 0.0269946
R14969 gnd.n3562 gnd.n3561 0.0269946
R14970 gnd.n3571 gnd.n2717 0.0269946
R14971 gnd.n3573 gnd.n3572 0.0269946
R14972 gnd.n3574 gnd.n2715 0.0269946
R14973 gnd.n3581 gnd.n3577 0.0269946
R14974 gnd.n3580 gnd.n3579 0.0269946
R14975 gnd.n3578 gnd.n2694 0.0269946
R14976 gnd.n3603 gnd.n2695 0.0269946
R14977 gnd.n3602 gnd.n2696 0.0269946
R14978 gnd.n3649 gnd.n2670 0.0269946
R14979 gnd.n3651 gnd.n3650 0.0269946
R14980 gnd.n3661 gnd.n2663 0.0269946
R14981 gnd.n3920 gnd.n2661 0.0269946
R14982 gnd.n3925 gnd.n3923 0.0269946
R14983 gnd.n3924 gnd.n2642 0.0269946
R14984 gnd.n3949 gnd.n3948 0.0269946
R14985 gnd.n4755 gnd.n2312 0.022519
R14986 gnd.n4754 gnd.n2313 0.022519
R14987 gnd.n4751 gnd.n4750 0.022519
R14988 gnd.n4747 gnd.n2319 0.022519
R14989 gnd.n4746 gnd.n2325 0.022519
R14990 gnd.n4743 gnd.n4742 0.022519
R14991 gnd.n4739 gnd.n2331 0.022519
R14992 gnd.n4738 gnd.n2335 0.022519
R14993 gnd.n4735 gnd.n4734 0.022519
R14994 gnd.n4731 gnd.n2342 0.022519
R14995 gnd.n4730 gnd.n2348 0.022519
R14996 gnd.n4727 gnd.n4726 0.022519
R14997 gnd.n4723 gnd.n2354 0.022519
R14998 gnd.n4722 gnd.n2358 0.022519
R14999 gnd.n4719 gnd.n4718 0.022519
R15000 gnd.n4715 gnd.n2365 0.022519
R15001 gnd.n4714 gnd.n2372 0.022519
R15002 gnd.n2380 gnd.n2378 0.022519
R15003 gnd.n4708 gnd.n4707 0.022519
R15004 gnd.n6129 gnd.n1311 0.022519
R15005 gnd.n6128 gnd.n1315 0.022519
R15006 gnd.n6125 gnd.n6124 0.022519
R15007 gnd.n6121 gnd.n1320 0.022519
R15008 gnd.n6120 gnd.n1324 0.022519
R15009 gnd.n6117 gnd.n6116 0.022519
R15010 gnd.n6113 gnd.n1328 0.022519
R15011 gnd.n6112 gnd.n1332 0.022519
R15012 gnd.n6109 gnd.n6108 0.022519
R15013 gnd.n6105 gnd.n1336 0.022519
R15014 gnd.n6104 gnd.n1340 0.022519
R15015 gnd.n6101 gnd.n6100 0.022519
R15016 gnd.n6097 gnd.n1344 0.022519
R15017 gnd.n6096 gnd.n1348 0.022519
R15018 gnd.n6093 gnd.n6092 0.022519
R15019 gnd.n6089 gnd.n1352 0.022519
R15020 gnd.n6088 gnd.n1358 0.022519
R15021 gnd.n1637 gnd.n1361 0.022519
R15022 gnd.n5733 gnd.n1636 0.022519
R15023 gnd.n5734 gnd.n1635 0.0218415
R15024 gnd.n4699 gnd.n2110 0.0218415
R15025 gnd.n3268 gnd.n3267 0.0202011
R15026 gnd.n3267 gnd.n3266 0.0148637
R15027 gnd.n3918 gnd.n3662 0.0144266
R15028 gnd.n3919 gnd.n3918 0.0130679
R15029 gnd.n2312 gnd.n2306 0.0123564
R15030 gnd.n4755 gnd.n4754 0.0123564
R15031 gnd.n4751 gnd.n2313 0.0123564
R15032 gnd.n4750 gnd.n2319 0.0123564
R15033 gnd.n4747 gnd.n4746 0.0123564
R15034 gnd.n4743 gnd.n2325 0.0123564
R15035 gnd.n4742 gnd.n2331 0.0123564
R15036 gnd.n4739 gnd.n4738 0.0123564
R15037 gnd.n4735 gnd.n2335 0.0123564
R15038 gnd.n4734 gnd.n2342 0.0123564
R15039 gnd.n4731 gnd.n4730 0.0123564
R15040 gnd.n4727 gnd.n2348 0.0123564
R15041 gnd.n4726 gnd.n2354 0.0123564
R15042 gnd.n4723 gnd.n4722 0.0123564
R15043 gnd.n4719 gnd.n2358 0.0123564
R15044 gnd.n4718 gnd.n2365 0.0123564
R15045 gnd.n4715 gnd.n4714 0.0123564
R15046 gnd.n2378 gnd.n2372 0.0123564
R15047 gnd.n4708 gnd.n2380 0.0123564
R15048 gnd.n6132 gnd.n1311 0.0123564
R15049 gnd.n6129 gnd.n6128 0.0123564
R15050 gnd.n6125 gnd.n1315 0.0123564
R15051 gnd.n6124 gnd.n1320 0.0123564
R15052 gnd.n6121 gnd.n6120 0.0123564
R15053 gnd.n6117 gnd.n1324 0.0123564
R15054 gnd.n6116 gnd.n1328 0.0123564
R15055 gnd.n6113 gnd.n6112 0.0123564
R15056 gnd.n6109 gnd.n1332 0.0123564
R15057 gnd.n6108 gnd.n1336 0.0123564
R15058 gnd.n6105 gnd.n6104 0.0123564
R15059 gnd.n6101 gnd.n1340 0.0123564
R15060 gnd.n6100 gnd.n1344 0.0123564
R15061 gnd.n6097 gnd.n6096 0.0123564
R15062 gnd.n6093 gnd.n1348 0.0123564
R15063 gnd.n6092 gnd.n1352 0.0123564
R15064 gnd.n6089 gnd.n6088 0.0123564
R15065 gnd.n1361 gnd.n1358 0.0123564
R15066 gnd.n1637 gnd.n1636 0.0123564
R15067 gnd.n3287 gnd.n3001 0.00797283
R15068 gnd.n3289 gnd.n3288 0.00797283
R15069 gnd.n3290 gnd.n2996 0.00797283
R15070 gnd.n3298 gnd.n2994 0.00797283
R15071 gnd.n3300 gnd.n3299 0.00797283
R15072 gnd.n3318 gnd.n2975 0.00797283
R15073 gnd.n3320 gnd.n3319 0.00797283
R15074 gnd.n3321 gnd.n2970 0.00797283
R15075 gnd.n2969 gnd.n2965 0.00797283
R15076 gnd.n3331 gnd.n3330 0.00797283
R15077 gnd.n2967 gnd.n2966 0.00797283
R15078 gnd.n2949 gnd.n2948 0.00797283
R15079 gnd.n3351 gnd.n3350 0.00797283
R15080 gnd.n2950 gnd.n2925 0.00797283
R15081 gnd.n3385 gnd.n3384 0.00797283
R15082 gnd.n3387 gnd.n3386 0.00797283
R15083 gnd.n2920 gnd.n2872 0.00797283
R15084 gnd.n2922 gnd.n2873 0.00797283
R15085 gnd.n3396 gnd.n2874 0.00797283
R15086 gnd.n3398 gnd.n3397 0.00797283
R15087 gnd.n3400 gnd.n3399 0.00797283
R15088 gnd.n3402 gnd.n2894 0.00797283
R15089 gnd.n3405 gnd.n2895 0.00797283
R15090 gnd.n3407 gnd.n2896 0.00797283
R15091 gnd.n3410 gnd.n3408 0.00797283
R15092 gnd.n3409 gnd.n2779 0.00797283
R15093 gnd.n3477 gnd.n3475 0.00797283
R15094 gnd.n3476 gnd.n2772 0.00797283
R15095 gnd.n3487 gnd.n3486 0.00797283
R15096 gnd.n3489 gnd.n3488 0.00797283
R15097 gnd.n3492 gnd.n2770 0.00797283
R15098 gnd.n3496 gnd.n3495 0.00797283
R15099 gnd.n3494 gnd.n3493 0.00797283
R15100 gnd.n2750 gnd.n2749 0.00797283
R15101 gnd.n3518 gnd.n3517 0.00797283
R15102 gnd.n2751 gnd.n2724 0.00797283
R15103 gnd.n3562 gnd.n3560 0.00797283
R15104 gnd.n3561 gnd.n2717 0.00797283
R15105 gnd.n3572 gnd.n3571 0.00797283
R15106 gnd.n3574 gnd.n3573 0.00797283
R15107 gnd.n3577 gnd.n2715 0.00797283
R15108 gnd.n3581 gnd.n3580 0.00797283
R15109 gnd.n3579 gnd.n3578 0.00797283
R15110 gnd.n2695 gnd.n2694 0.00797283
R15111 gnd.n3603 gnd.n3602 0.00797283
R15112 gnd.n2696 gnd.n2670 0.00797283
R15113 gnd.n3651 gnd.n3649 0.00797283
R15114 gnd.n3650 gnd.n2663 0.00797283
R15115 gnd.n3662 gnd.n3661 0.00797283
R15116 gnd.n3920 gnd.n3919 0.00797283
R15117 gnd.n3923 gnd.n2661 0.00797283
R15118 gnd.n3925 gnd.n3924 0.00797283
R15119 gnd.n3948 gnd.n2642 0.00797283
R15120 gnd.n3949 gnd.n2606 0.00797283
R15121 gnd.n4760 gnd.n4759 0.00592005
R15122 gnd.n6134 gnd.n6133 0.00592005
R15123 a_n7636_8799.n175 a_n7636_8799.t52 485.149
R15124 a_n7636_8799.n191 a_n7636_8799.t61 485.149
R15125 a_n7636_8799.n208 a_n7636_8799.t91 485.149
R15126 a_n7636_8799.n124 a_n7636_8799.t111 485.149
R15127 a_n7636_8799.n140 a_n7636_8799.t124 485.149
R15128 a_n7636_8799.n157 a_n7636_8799.t90 485.149
R15129 a_n7636_8799.n185 a_n7636_8799.t71 464.166
R15130 a_n7636_8799.n184 a_n7636_8799.t53 464.166
R15131 a_n7636_8799.n170 a_n7636_8799.t116 464.166
R15132 a_n7636_8799.n183 a_n7636_8799.t84 464.166
R15133 a_n7636_8799.n182 a_n7636_8799.t82 464.166
R15134 a_n7636_8799.n171 a_n7636_8799.t34 464.166
R15135 a_n7636_8799.n181 a_n7636_8799.t88 464.166
R15136 a_n7636_8799.n180 a_n7636_8799.t87 464.166
R15137 a_n7636_8799.n172 a_n7636_8799.t36 464.166
R15138 a_n7636_8799.n179 a_n7636_8799.t35 464.166
R15139 a_n7636_8799.n178 a_n7636_8799.t104 464.166
R15140 a_n7636_8799.n173 a_n7636_8799.t48 464.166
R15141 a_n7636_8799.n177 a_n7636_8799.t39 464.166
R15142 a_n7636_8799.n176 a_n7636_8799.t108 464.166
R15143 a_n7636_8799.n174 a_n7636_8799.t70 464.166
R15144 a_n7636_8799.n201 a_n7636_8799.t80 464.166
R15145 a_n7636_8799.n200 a_n7636_8799.t60 464.166
R15146 a_n7636_8799.n186 a_n7636_8799.t127 464.166
R15147 a_n7636_8799.n199 a_n7636_8799.t97 464.166
R15148 a_n7636_8799.n198 a_n7636_8799.t96 464.166
R15149 a_n7636_8799.n187 a_n7636_8799.t42 464.166
R15150 a_n7636_8799.n197 a_n7636_8799.t100 464.166
R15151 a_n7636_8799.n196 a_n7636_8799.t99 464.166
R15152 a_n7636_8799.n188 a_n7636_8799.t44 464.166
R15153 a_n7636_8799.n195 a_n7636_8799.t43 464.166
R15154 a_n7636_8799.n194 a_n7636_8799.t119 464.166
R15155 a_n7636_8799.n189 a_n7636_8799.t59 464.166
R15156 a_n7636_8799.n193 a_n7636_8799.t47 464.166
R15157 a_n7636_8799.n192 a_n7636_8799.t120 464.166
R15158 a_n7636_8799.n190 a_n7636_8799.t81 464.166
R15159 a_n7636_8799.n218 a_n7636_8799.t103 464.166
R15160 a_n7636_8799.n217 a_n7636_8799.t50 464.166
R15161 a_n7636_8799.n203 a_n7636_8799.t86 464.166
R15162 a_n7636_8799.n216 a_n7636_8799.t38 464.166
R15163 a_n7636_8799.n215 a_n7636_8799.t55 464.166
R15164 a_n7636_8799.n204 a_n7636_8799.t123 464.166
R15165 a_n7636_8799.n214 a_n7636_8799.t95 464.166
R15166 a_n7636_8799.n213 a_n7636_8799.t118 464.166
R15167 a_n7636_8799.n205 a_n7636_8799.t79 464.166
R15168 a_n7636_8799.n212 a_n7636_8799.t98 464.166
R15169 a_n7636_8799.n211 a_n7636_8799.t46 464.166
R15170 a_n7636_8799.n206 a_n7636_8799.t115 464.166
R15171 a_n7636_8799.n210 a_n7636_8799.t64 464.166
R15172 a_n7636_8799.n209 a_n7636_8799.t109 464.166
R15173 a_n7636_8799.n207 a_n7636_8799.t54 464.166
R15174 a_n7636_8799.n123 a_n7636_8799.t113 464.166
R15175 a_n7636_8799.n126 a_n7636_8799.t69 464.166
R15176 a_n7636_8799.n122 a_n7636_8799.t94 464.166
R15177 a_n7636_8799.n127 a_n7636_8799.t110 464.166
R15178 a_n7636_8799.n128 a_n7636_8799.t67 464.166
R15179 a_n7636_8799.n129 a_n7636_8799.t68 464.166
R15180 a_n7636_8799.n130 a_n7636_8799.t92 464.166
R15181 a_n7636_8799.n121 a_n7636_8799.t57 464.166
R15182 a_n7636_8799.n131 a_n7636_8799.t58 464.166
R15183 a_n7636_8799.n132 a_n7636_8799.t89 464.166
R15184 a_n7636_8799.n133 a_n7636_8799.t32 464.166
R15185 a_n7636_8799.n134 a_n7636_8799.t56 464.166
R15186 a_n7636_8799.n120 a_n7636_8799.t74 464.166
R15187 a_n7636_8799.n135 a_n7636_8799.t112 464.166
R15188 a_n7636_8799.n139 a_n7636_8799.t126 464.166
R15189 a_n7636_8799.n142 a_n7636_8799.t77 464.166
R15190 a_n7636_8799.n138 a_n7636_8799.t107 464.166
R15191 a_n7636_8799.n143 a_n7636_8799.t122 464.166
R15192 a_n7636_8799.n144 a_n7636_8799.t75 464.166
R15193 a_n7636_8799.n145 a_n7636_8799.t76 464.166
R15194 a_n7636_8799.n146 a_n7636_8799.t105 464.166
R15195 a_n7636_8799.n137 a_n7636_8799.t65 464.166
R15196 a_n7636_8799.n147 a_n7636_8799.t66 464.166
R15197 a_n7636_8799.n148 a_n7636_8799.t101 464.166
R15198 a_n7636_8799.n149 a_n7636_8799.t40 464.166
R15199 a_n7636_8799.n150 a_n7636_8799.t62 464.166
R15200 a_n7636_8799.n136 a_n7636_8799.t83 464.166
R15201 a_n7636_8799.n151 a_n7636_8799.t125 464.166
R15202 a_n7636_8799.n156 a_n7636_8799.t72 464.166
R15203 a_n7636_8799.n159 a_n7636_8799.t106 464.166
R15204 a_n7636_8799.n155 a_n7636_8799.t63 464.166
R15205 a_n7636_8799.n160 a_n7636_8799.t114 464.166
R15206 a_n7636_8799.n161 a_n7636_8799.t45 464.166
R15207 a_n7636_8799.n162 a_n7636_8799.t33 464.166
R15208 a_n7636_8799.n163 a_n7636_8799.t78 464.166
R15209 a_n7636_8799.n154 a_n7636_8799.t117 464.166
R15210 a_n7636_8799.n164 a_n7636_8799.t93 464.166
R15211 a_n7636_8799.n165 a_n7636_8799.t121 464.166
R15212 a_n7636_8799.n166 a_n7636_8799.t73 464.166
R15213 a_n7636_8799.n167 a_n7636_8799.t37 464.166
R15214 a_n7636_8799.n153 a_n7636_8799.t85 464.166
R15215 a_n7636_8799.n168 a_n7636_8799.t49 464.166
R15216 a_n7636_8799.n52 a_n7636_8799.n33 74.4178
R15217 a_n7636_8799.n176 a_n7636_8799.n52 12.4674
R15218 a_n7636_8799.n51 a_n7636_8799.n33 80.107
R15219 a_n7636_8799.n51 a_n7636_8799.n177 1.08907
R15220 a_n7636_8799.n34 a_n7636_8799.n50 75.3623
R15221 a_n7636_8799.n49 a_n7636_8799.n34 70.3058
R15222 a_n7636_8799.n36 a_n7636_8799.n48 70.1674
R15223 a_n7636_8799.n48 a_n7636_8799.n172 20.9683
R15224 a_n7636_8799.n47 a_n7636_8799.n36 75.0448
R15225 a_n7636_8799.n180 a_n7636_8799.n47 11.2134
R15226 a_n7636_8799.n46 a_n7636_8799.n35 80.4688
R15227 a_n7636_8799.n35 a_n7636_8799.n45 74.73
R15228 a_n7636_8799.n44 a_n7636_8799.n37 70.1674
R15229 a_n7636_8799.n183 a_n7636_8799.n44 20.9683
R15230 a_n7636_8799.n37 a_n7636_8799.n43 70.5844
R15231 a_n7636_8799.n43 a_n7636_8799.n170 20.1342
R15232 a_n7636_8799.n42 a_n7636_8799.n38 75.6825
R15233 a_n7636_8799.n184 a_n7636_8799.n42 9.93802
R15234 a_n7636_8799.n38 a_n7636_8799.n185 161.3
R15235 a_n7636_8799.n63 a_n7636_8799.n27 74.4178
R15236 a_n7636_8799.n192 a_n7636_8799.n63 12.4674
R15237 a_n7636_8799.n62 a_n7636_8799.n27 80.107
R15238 a_n7636_8799.n62 a_n7636_8799.n193 1.08907
R15239 a_n7636_8799.n28 a_n7636_8799.n61 75.3623
R15240 a_n7636_8799.n60 a_n7636_8799.n28 70.3058
R15241 a_n7636_8799.n30 a_n7636_8799.n59 70.1674
R15242 a_n7636_8799.n59 a_n7636_8799.n188 20.9683
R15243 a_n7636_8799.n58 a_n7636_8799.n30 75.0448
R15244 a_n7636_8799.n196 a_n7636_8799.n58 11.2134
R15245 a_n7636_8799.n57 a_n7636_8799.n29 80.4688
R15246 a_n7636_8799.n29 a_n7636_8799.n56 74.73
R15247 a_n7636_8799.n55 a_n7636_8799.n31 70.1674
R15248 a_n7636_8799.n199 a_n7636_8799.n55 20.9683
R15249 a_n7636_8799.n31 a_n7636_8799.n54 70.5844
R15250 a_n7636_8799.n54 a_n7636_8799.n186 20.1342
R15251 a_n7636_8799.n53 a_n7636_8799.n32 75.6825
R15252 a_n7636_8799.n200 a_n7636_8799.n53 9.93802
R15253 a_n7636_8799.n32 a_n7636_8799.n201 161.3
R15254 a_n7636_8799.n74 a_n7636_8799.n21 74.4178
R15255 a_n7636_8799.n209 a_n7636_8799.n74 12.4674
R15256 a_n7636_8799.n73 a_n7636_8799.n21 80.107
R15257 a_n7636_8799.n73 a_n7636_8799.n210 1.08907
R15258 a_n7636_8799.n22 a_n7636_8799.n72 75.3623
R15259 a_n7636_8799.n71 a_n7636_8799.n22 70.3058
R15260 a_n7636_8799.n24 a_n7636_8799.n70 70.1674
R15261 a_n7636_8799.n70 a_n7636_8799.n205 20.9683
R15262 a_n7636_8799.n69 a_n7636_8799.n24 75.0448
R15263 a_n7636_8799.n213 a_n7636_8799.n69 11.2134
R15264 a_n7636_8799.n68 a_n7636_8799.n23 80.4688
R15265 a_n7636_8799.n23 a_n7636_8799.n67 74.73
R15266 a_n7636_8799.n66 a_n7636_8799.n25 70.1674
R15267 a_n7636_8799.n216 a_n7636_8799.n66 20.9683
R15268 a_n7636_8799.n25 a_n7636_8799.n65 70.5844
R15269 a_n7636_8799.n65 a_n7636_8799.n203 20.1342
R15270 a_n7636_8799.n64 a_n7636_8799.n26 75.6825
R15271 a_n7636_8799.n217 a_n7636_8799.n64 9.93802
R15272 a_n7636_8799.n26 a_n7636_8799.n218 161.3
R15273 a_n7636_8799.n16 a_n7636_8799.n85 70.1674
R15274 a_n7636_8799.n135 a_n7636_8799.n85 20.9683
R15275 a_n7636_8799.n84 a_n7636_8799.n16 74.4178
R15276 a_n7636_8799.n84 a_n7636_8799.n120 12.4674
R15277 a_n7636_8799.n15 a_n7636_8799.n83 80.107
R15278 a_n7636_8799.n134 a_n7636_8799.n83 1.08907
R15279 a_n7636_8799.n82 a_n7636_8799.n15 75.3623
R15280 a_n7636_8799.n17 a_n7636_8799.n81 70.3058
R15281 a_n7636_8799.n80 a_n7636_8799.n17 70.1674
R15282 a_n7636_8799.n80 a_n7636_8799.n121 20.9683
R15283 a_n7636_8799.n18 a_n7636_8799.n79 75.0448
R15284 a_n7636_8799.n130 a_n7636_8799.n79 11.2134
R15285 a_n7636_8799.n78 a_n7636_8799.n18 80.4688
R15286 a_n7636_8799.n19 a_n7636_8799.n77 74.73
R15287 a_n7636_8799.n76 a_n7636_8799.n19 70.1674
R15288 a_n7636_8799.n76 a_n7636_8799.n122 20.9683
R15289 a_n7636_8799.n20 a_n7636_8799.n75 70.5844
R15290 a_n7636_8799.n126 a_n7636_8799.n75 20.1342
R15291 a_n7636_8799.n125 a_n7636_8799.n20 161.3
R15292 a_n7636_8799.n10 a_n7636_8799.n96 70.1674
R15293 a_n7636_8799.n151 a_n7636_8799.n96 20.9683
R15294 a_n7636_8799.n95 a_n7636_8799.n10 74.4178
R15295 a_n7636_8799.n95 a_n7636_8799.n136 12.4674
R15296 a_n7636_8799.n9 a_n7636_8799.n94 80.107
R15297 a_n7636_8799.n150 a_n7636_8799.n94 1.08907
R15298 a_n7636_8799.n93 a_n7636_8799.n9 75.3623
R15299 a_n7636_8799.n11 a_n7636_8799.n92 70.3058
R15300 a_n7636_8799.n91 a_n7636_8799.n11 70.1674
R15301 a_n7636_8799.n91 a_n7636_8799.n137 20.9683
R15302 a_n7636_8799.n12 a_n7636_8799.n90 75.0448
R15303 a_n7636_8799.n146 a_n7636_8799.n90 11.2134
R15304 a_n7636_8799.n89 a_n7636_8799.n12 80.4688
R15305 a_n7636_8799.n13 a_n7636_8799.n88 74.73
R15306 a_n7636_8799.n87 a_n7636_8799.n13 70.1674
R15307 a_n7636_8799.n87 a_n7636_8799.n138 20.9683
R15308 a_n7636_8799.n14 a_n7636_8799.n86 70.5844
R15309 a_n7636_8799.n142 a_n7636_8799.n86 20.1342
R15310 a_n7636_8799.n141 a_n7636_8799.n14 161.3
R15311 a_n7636_8799.n4 a_n7636_8799.n107 70.1674
R15312 a_n7636_8799.n168 a_n7636_8799.n107 20.9683
R15313 a_n7636_8799.n106 a_n7636_8799.n4 74.4178
R15314 a_n7636_8799.n106 a_n7636_8799.n153 12.4674
R15315 a_n7636_8799.n3 a_n7636_8799.n105 80.107
R15316 a_n7636_8799.n167 a_n7636_8799.n105 1.08907
R15317 a_n7636_8799.n104 a_n7636_8799.n3 75.3623
R15318 a_n7636_8799.n5 a_n7636_8799.n103 70.3058
R15319 a_n7636_8799.n102 a_n7636_8799.n5 70.1674
R15320 a_n7636_8799.n102 a_n7636_8799.n154 20.9683
R15321 a_n7636_8799.n6 a_n7636_8799.n101 75.0448
R15322 a_n7636_8799.n163 a_n7636_8799.n101 11.2134
R15323 a_n7636_8799.n100 a_n7636_8799.n6 80.4688
R15324 a_n7636_8799.n7 a_n7636_8799.n99 74.73
R15325 a_n7636_8799.n98 a_n7636_8799.n7 70.1674
R15326 a_n7636_8799.n98 a_n7636_8799.n155 20.9683
R15327 a_n7636_8799.n8 a_n7636_8799.n97 70.5844
R15328 a_n7636_8799.n159 a_n7636_8799.n97 20.1342
R15329 a_n7636_8799.n158 a_n7636_8799.n8 161.3
R15330 a_n7636_8799.n39 a_n7636_8799.n108 98.9633
R15331 a_n7636_8799.n41 a_n7636_8799.n223 98.9631
R15332 a_n7636_8799.n41 a_n7636_8799.n224 98.6055
R15333 a_n7636_8799.n41 a_n7636_8799.n225 98.6055
R15334 a_n7636_8799.n40 a_n7636_8799.n111 98.6055
R15335 a_n7636_8799.n40 a_n7636_8799.n110 98.6055
R15336 a_n7636_8799.n39 a_n7636_8799.n109 98.6055
R15337 a_n7636_8799.n227 a_n7636_8799.n226 98.6054
R15338 a_n7636_8799.n1 a_n7636_8799.n112 81.4626
R15339 a_n7636_8799.n2 a_n7636_8799.n116 81.4626
R15340 a_n7636_8799.n2 a_n7636_8799.n114 81.4626
R15341 a_n7636_8799.n0 a_n7636_8799.n118 80.9324
R15342 a_n7636_8799.n1 a_n7636_8799.n119 80.9324
R15343 a_n7636_8799.n1 a_n7636_8799.n113 80.9324
R15344 a_n7636_8799.n2 a_n7636_8799.n117 80.9324
R15345 a_n7636_8799.n2 a_n7636_8799.n115 80.9324
R15346 a_n7636_8799.n33 a_n7636_8799.n175 70.4033
R15347 a_n7636_8799.n27 a_n7636_8799.n191 70.4033
R15348 a_n7636_8799.n21 a_n7636_8799.n208 70.4033
R15349 a_n7636_8799.n20 a_n7636_8799.n124 70.4033
R15350 a_n7636_8799.n14 a_n7636_8799.n140 70.4033
R15351 a_n7636_8799.n8 a_n7636_8799.n157 70.4033
R15352 a_n7636_8799.n185 a_n7636_8799.n184 48.2005
R15353 a_n7636_8799.n44 a_n7636_8799.n182 20.9683
R15354 a_n7636_8799.n181 a_n7636_8799.n180 48.2005
R15355 a_n7636_8799.n179 a_n7636_8799.n48 20.9683
R15356 a_n7636_8799.n177 a_n7636_8799.n173 48.2005
R15357 a_n7636_8799.n201 a_n7636_8799.n200 48.2005
R15358 a_n7636_8799.n55 a_n7636_8799.n198 20.9683
R15359 a_n7636_8799.n197 a_n7636_8799.n196 48.2005
R15360 a_n7636_8799.n195 a_n7636_8799.n59 20.9683
R15361 a_n7636_8799.n193 a_n7636_8799.n189 48.2005
R15362 a_n7636_8799.n218 a_n7636_8799.n217 48.2005
R15363 a_n7636_8799.n66 a_n7636_8799.n215 20.9683
R15364 a_n7636_8799.n214 a_n7636_8799.n213 48.2005
R15365 a_n7636_8799.n212 a_n7636_8799.n70 20.9683
R15366 a_n7636_8799.n210 a_n7636_8799.n206 48.2005
R15367 a_n7636_8799.n127 a_n7636_8799.n76 20.9683
R15368 a_n7636_8799.n130 a_n7636_8799.n129 48.2005
R15369 a_n7636_8799.n131 a_n7636_8799.n80 20.9683
R15370 a_n7636_8799.n134 a_n7636_8799.n133 48.2005
R15371 a_n7636_8799.t41 a_n7636_8799.n85 485.135
R15372 a_n7636_8799.n143 a_n7636_8799.n87 20.9683
R15373 a_n7636_8799.n146 a_n7636_8799.n145 48.2005
R15374 a_n7636_8799.n147 a_n7636_8799.n91 20.9683
R15375 a_n7636_8799.n150 a_n7636_8799.n149 48.2005
R15376 a_n7636_8799.t51 a_n7636_8799.n96 485.135
R15377 a_n7636_8799.n160 a_n7636_8799.n98 20.9683
R15378 a_n7636_8799.n163 a_n7636_8799.n162 48.2005
R15379 a_n7636_8799.n164 a_n7636_8799.n102 20.9683
R15380 a_n7636_8799.n167 a_n7636_8799.n166 48.2005
R15381 a_n7636_8799.t102 a_n7636_8799.n107 485.135
R15382 a_n7636_8799.n46 a_n7636_8799.n171 47.835
R15383 a_n7636_8799.n49 a_n7636_8799.n178 20.6913
R15384 a_n7636_8799.n57 a_n7636_8799.n187 47.835
R15385 a_n7636_8799.n60 a_n7636_8799.n194 20.6913
R15386 a_n7636_8799.n68 a_n7636_8799.n204 47.835
R15387 a_n7636_8799.n71 a_n7636_8799.n211 20.6913
R15388 a_n7636_8799.n128 a_n7636_8799.n78 47.835
R15389 a_n7636_8799.n132 a_n7636_8799.n81 20.6913
R15390 a_n7636_8799.n144 a_n7636_8799.n89 47.835
R15391 a_n7636_8799.n148 a_n7636_8799.n92 20.6913
R15392 a_n7636_8799.n161 a_n7636_8799.n100 47.835
R15393 a_n7636_8799.n165 a_n7636_8799.n103 20.6913
R15394 a_n7636_8799.n183 a_n7636_8799.n43 22.3251
R15395 a_n7636_8799.n199 a_n7636_8799.n54 22.3251
R15396 a_n7636_8799.n216 a_n7636_8799.n65 22.3251
R15397 a_n7636_8799.n122 a_n7636_8799.n75 22.3251
R15398 a_n7636_8799.n138 a_n7636_8799.n86 22.3251
R15399 a_n7636_8799.n155 a_n7636_8799.n97 22.3251
R15400 a_n7636_8799.n226 a_n7636_8799.n222 31.7372
R15401 a_n7636_8799.n52 a_n7636_8799.n174 33.6462
R15402 a_n7636_8799.n63 a_n7636_8799.n190 33.6462
R15403 a_n7636_8799.n74 a_n7636_8799.n207 33.6462
R15404 a_n7636_8799.n126 a_n7636_8799.n125 27.0217
R15405 a_n7636_8799.n135 a_n7636_8799.n84 33.6462
R15406 a_n7636_8799.n142 a_n7636_8799.n141 27.0217
R15407 a_n7636_8799.n151 a_n7636_8799.n95 33.6462
R15408 a_n7636_8799.n159 a_n7636_8799.n158 27.0217
R15409 a_n7636_8799.n168 a_n7636_8799.n106 33.6462
R15410 a_n7636_8799.n45 a_n7636_8799.n171 11.843
R15411 a_n7636_8799.n178 a_n7636_8799.n50 36.139
R15412 a_n7636_8799.n56 a_n7636_8799.n187 11.843
R15413 a_n7636_8799.n194 a_n7636_8799.n61 36.139
R15414 a_n7636_8799.n67 a_n7636_8799.n204 11.843
R15415 a_n7636_8799.n211 a_n7636_8799.n72 36.139
R15416 a_n7636_8799.n128 a_n7636_8799.n77 11.843
R15417 a_n7636_8799.n132 a_n7636_8799.n82 36.139
R15418 a_n7636_8799.n144 a_n7636_8799.n88 11.843
R15419 a_n7636_8799.n148 a_n7636_8799.n93 36.139
R15420 a_n7636_8799.n161 a_n7636_8799.n99 11.843
R15421 a_n7636_8799.n165 a_n7636_8799.n104 36.139
R15422 a_n7636_8799.n47 a_n7636_8799.n172 35.3134
R15423 a_n7636_8799.n58 a_n7636_8799.n188 35.3134
R15424 a_n7636_8799.n69 a_n7636_8799.n205 35.3134
R15425 a_n7636_8799.n121 a_n7636_8799.n79 35.3134
R15426 a_n7636_8799.n137 a_n7636_8799.n90 35.3134
R15427 a_n7636_8799.n154 a_n7636_8799.n101 35.3134
R15428 a_n7636_8799.n182 a_n7636_8799.n45 34.4824
R15429 a_n7636_8799.n50 a_n7636_8799.n173 10.5784
R15430 a_n7636_8799.n198 a_n7636_8799.n56 34.4824
R15431 a_n7636_8799.n61 a_n7636_8799.n189 10.5784
R15432 a_n7636_8799.n215 a_n7636_8799.n67 34.4824
R15433 a_n7636_8799.n72 a_n7636_8799.n206 10.5784
R15434 a_n7636_8799.n77 a_n7636_8799.n127 34.4824
R15435 a_n7636_8799.n133 a_n7636_8799.n82 10.5784
R15436 a_n7636_8799.n88 a_n7636_8799.n143 34.4824
R15437 a_n7636_8799.n149 a_n7636_8799.n93 10.5784
R15438 a_n7636_8799.n99 a_n7636_8799.n160 34.4824
R15439 a_n7636_8799.n166 a_n7636_8799.n104 10.5784
R15440 a_n7636_8799.n42 a_n7636_8799.n170 36.9592
R15441 a_n7636_8799.n53 a_n7636_8799.n186 36.9592
R15442 a_n7636_8799.n64 a_n7636_8799.n203 36.9592
R15443 a_n7636_8799.n125 a_n7636_8799.n123 21.1793
R15444 a_n7636_8799.n141 a_n7636_8799.n139 21.1793
R15445 a_n7636_8799.n158 a_n7636_8799.n156 21.1793
R15446 a_n7636_8799.n175 a_n7636_8799.n174 20.9576
R15447 a_n7636_8799.n191 a_n7636_8799.n190 20.9576
R15448 a_n7636_8799.n208 a_n7636_8799.n207 20.9576
R15449 a_n7636_8799.n124 a_n7636_8799.n123 20.9576
R15450 a_n7636_8799.n140 a_n7636_8799.n139 20.9576
R15451 a_n7636_8799.n157 a_n7636_8799.n156 20.9576
R15452 a_n7636_8799.n222 a_n7636_8799.n40 18.8589
R15453 a_n7636_8799.n221 a_n7636_8799.n1 12.3339
R15454 a_n7636_8799.n222 a_n7636_8799.n221 11.4887
R15455 a_n7636_8799.n202 a_n7636_8799.n38 9.07815
R15456 a_n7636_8799.n152 a_n7636_8799.n16 9.07815
R15457 a_n7636_8799.n220 a_n7636_8799.n169 6.96667
R15458 a_n7636_8799.n220 a_n7636_8799.n219 6.62419
R15459 a_n7636_8799.n202 a_n7636_8799.n32 4.9702
R15460 a_n7636_8799.n219 a_n7636_8799.n26 4.9702
R15461 a_n7636_8799.n152 a_n7636_8799.n10 4.9702
R15462 a_n7636_8799.n169 a_n7636_8799.n4 4.9702
R15463 a_n7636_8799.n219 a_n7636_8799.n202 4.10845
R15464 a_n7636_8799.n169 a_n7636_8799.n152 4.10845
R15465 a_n7636_8799.n223 a_n7636_8799.t27 3.61217
R15466 a_n7636_8799.n223 a_n7636_8799.t10 3.61217
R15467 a_n7636_8799.n224 a_n7636_8799.t8 3.61217
R15468 a_n7636_8799.n224 a_n7636_8799.t18 3.61217
R15469 a_n7636_8799.n225 a_n7636_8799.t28 3.61217
R15470 a_n7636_8799.n225 a_n7636_8799.t31 3.61217
R15471 a_n7636_8799.n111 a_n7636_8799.t17 3.61217
R15472 a_n7636_8799.n111 a_n7636_8799.t9 3.61217
R15473 a_n7636_8799.n110 a_n7636_8799.t26 3.61217
R15474 a_n7636_8799.n110 a_n7636_8799.t22 3.61217
R15475 a_n7636_8799.n109 a_n7636_8799.t16 3.61217
R15476 a_n7636_8799.n109 a_n7636_8799.t7 3.61217
R15477 a_n7636_8799.n108 a_n7636_8799.t14 3.61217
R15478 a_n7636_8799.n108 a_n7636_8799.t19 3.61217
R15479 a_n7636_8799.n227 a_n7636_8799.t21 3.61217
R15480 a_n7636_8799.t6 a_n7636_8799.n227 3.61217
R15481 a_n7636_8799.n221 a_n7636_8799.n220 3.4105
R15482 a_n7636_8799.n118 a_n7636_8799.t25 2.82907
R15483 a_n7636_8799.n118 a_n7636_8799.t3 2.82907
R15484 a_n7636_8799.n119 a_n7636_8799.t13 2.82907
R15485 a_n7636_8799.n119 a_n7636_8799.t29 2.82907
R15486 a_n7636_8799.n113 a_n7636_8799.t0 2.82907
R15487 a_n7636_8799.n113 a_n7636_8799.t15 2.82907
R15488 a_n7636_8799.n112 a_n7636_8799.t11 2.82907
R15489 a_n7636_8799.n112 a_n7636_8799.t5 2.82907
R15490 a_n7636_8799.n116 a_n7636_8799.t4 2.82907
R15491 a_n7636_8799.n116 a_n7636_8799.t23 2.82907
R15492 a_n7636_8799.n117 a_n7636_8799.t30 2.82907
R15493 a_n7636_8799.n117 a_n7636_8799.t24 2.82907
R15494 a_n7636_8799.n115 a_n7636_8799.t20 2.82907
R15495 a_n7636_8799.n115 a_n7636_8799.t2 2.82907
R15496 a_n7636_8799.n114 a_n7636_8799.t12 2.82907
R15497 a_n7636_8799.n114 a_n7636_8799.t1 2.82907
R15498 a_n7636_8799.n51 a_n7636_8799.n176 47.0982
R15499 a_n7636_8799.n62 a_n7636_8799.n192 47.0982
R15500 a_n7636_8799.n73 a_n7636_8799.n209 47.0982
R15501 a_n7636_8799.n120 a_n7636_8799.n83 47.0982
R15502 a_n7636_8799.n136 a_n7636_8799.n94 47.0982
R15503 a_n7636_8799.n153 a_n7636_8799.n105 47.0982
R15504 a_n7636_8799.n0 a_n7636_8799.n2 33.2634
R15505 a_n7636_8799.n46 a_n7636_8799.n181 0.365327
R15506 a_n7636_8799.n179 a_n7636_8799.n49 21.4216
R15507 a_n7636_8799.n57 a_n7636_8799.n197 0.365327
R15508 a_n7636_8799.n195 a_n7636_8799.n60 21.4216
R15509 a_n7636_8799.n68 a_n7636_8799.n214 0.365327
R15510 a_n7636_8799.n212 a_n7636_8799.n71 21.4216
R15511 a_n7636_8799.n129 a_n7636_8799.n78 0.365327
R15512 a_n7636_8799.n81 a_n7636_8799.n131 21.4216
R15513 a_n7636_8799.n145 a_n7636_8799.n89 0.365327
R15514 a_n7636_8799.n92 a_n7636_8799.n147 21.4216
R15515 a_n7636_8799.n162 a_n7636_8799.n100 0.365327
R15516 a_n7636_8799.n103 a_n7636_8799.n164 21.4216
R15517 a_n7636_8799.n34 a_n7636_8799.n33 1.13686
R15518 a_n7636_8799.n28 a_n7636_8799.n27 1.13686
R15519 a_n7636_8799.n22 a_n7636_8799.n21 1.13686
R15520 a_n7636_8799.n16 a_n7636_8799.n15 1.13686
R15521 a_n7636_8799.n10 a_n7636_8799.n9 1.13686
R15522 a_n7636_8799.n4 a_n7636_8799.n3 1.13686
R15523 a_n7636_8799.n1 a_n7636_8799.n0 1.06084
R15524 a_n7636_8799.n38 a_n7636_8799.n37 0.758076
R15525 a_n7636_8799.n35 a_n7636_8799.n37 0.758076
R15526 a_n7636_8799.n36 a_n7636_8799.n35 0.758076
R15527 a_n7636_8799.n36 a_n7636_8799.n34 0.758076
R15528 a_n7636_8799.n32 a_n7636_8799.n31 0.758076
R15529 a_n7636_8799.n29 a_n7636_8799.n31 0.758076
R15530 a_n7636_8799.n30 a_n7636_8799.n29 0.758076
R15531 a_n7636_8799.n30 a_n7636_8799.n28 0.758076
R15532 a_n7636_8799.n26 a_n7636_8799.n25 0.758076
R15533 a_n7636_8799.n23 a_n7636_8799.n25 0.758076
R15534 a_n7636_8799.n24 a_n7636_8799.n23 0.758076
R15535 a_n7636_8799.n24 a_n7636_8799.n22 0.758076
R15536 a_n7636_8799.n19 a_n7636_8799.n20 0.758076
R15537 a_n7636_8799.n18 a_n7636_8799.n19 0.758076
R15538 a_n7636_8799.n17 a_n7636_8799.n18 0.758076
R15539 a_n7636_8799.n15 a_n7636_8799.n17 0.758076
R15540 a_n7636_8799.n13 a_n7636_8799.n14 0.758076
R15541 a_n7636_8799.n12 a_n7636_8799.n13 0.758076
R15542 a_n7636_8799.n11 a_n7636_8799.n12 0.758076
R15543 a_n7636_8799.n9 a_n7636_8799.n11 0.758076
R15544 a_n7636_8799.n7 a_n7636_8799.n8 0.758076
R15545 a_n7636_8799.n6 a_n7636_8799.n7 0.758076
R15546 a_n7636_8799.n5 a_n7636_8799.n6 0.758076
R15547 a_n7636_8799.n3 a_n7636_8799.n5 0.758076
R15548 a_n7636_8799.n226 a_n7636_8799.n41 0.716017
R15549 a_n7636_8799.n40 a_n7636_8799.n39 0.716017
R15550 vdd.n315 vdd.n279 756.745
R15551 vdd.n260 vdd.n224 756.745
R15552 vdd.n217 vdd.n181 756.745
R15553 vdd.n162 vdd.n126 756.745
R15554 vdd.n120 vdd.n84 756.745
R15555 vdd.n65 vdd.n29 756.745
R15556 vdd.n2046 vdd.n2010 756.745
R15557 vdd.n2101 vdd.n2065 756.745
R15558 vdd.n1948 vdd.n1912 756.745
R15559 vdd.n2003 vdd.n1967 756.745
R15560 vdd.n1851 vdd.n1815 756.745
R15561 vdd.n1906 vdd.n1870 756.745
R15562 vdd.n1224 vdd.t53 640.208
R15563 vdd.n952 vdd.t95 640.208
R15564 vdd.n1244 vdd.t68 640.208
R15565 vdd.n943 vdd.t113 640.208
R15566 vdd.n843 vdd.t71 640.208
R15567 vdd.n2621 vdd.t110 640.208
R15568 vdd.n804 vdd.t119 640.208
R15569 vdd.n2618 vdd.t99 640.208
R15570 vdd.n768 vdd.t49 640.208
R15571 vdd.n1014 vdd.t103 640.208
R15572 vdd.n1510 vdd.t86 592.009
R15573 vdd.n1666 vdd.t78 592.009
R15574 vdd.n1702 vdd.t89 592.009
R15575 vdd.n2186 vdd.t61 592.009
R15576 vdd.n1161 vdd.t92 592.009
R15577 vdd.n1121 vdd.t107 592.009
R15578 vdd.n405 vdd.t82 592.009
R15579 vdd.n419 vdd.t116 592.009
R15580 vdd.n431 vdd.t122 592.009
R15581 vdd.n723 vdd.t65 592.009
R15582 vdd.n686 vdd.t75 592.009
R15583 vdd.n3105 vdd.t57 592.009
R15584 vdd.n316 vdd.n315 585
R15585 vdd.n314 vdd.n281 585
R15586 vdd.n313 vdd.n312 585
R15587 vdd.n284 vdd.n282 585
R15588 vdd.n307 vdd.n306 585
R15589 vdd.n305 vdd.n304 585
R15590 vdd.n288 vdd.n287 585
R15591 vdd.n299 vdd.n298 585
R15592 vdd.n297 vdd.n296 585
R15593 vdd.n292 vdd.n291 585
R15594 vdd.n261 vdd.n260 585
R15595 vdd.n259 vdd.n226 585
R15596 vdd.n258 vdd.n257 585
R15597 vdd.n229 vdd.n227 585
R15598 vdd.n252 vdd.n251 585
R15599 vdd.n250 vdd.n249 585
R15600 vdd.n233 vdd.n232 585
R15601 vdd.n244 vdd.n243 585
R15602 vdd.n242 vdd.n241 585
R15603 vdd.n237 vdd.n236 585
R15604 vdd.n218 vdd.n217 585
R15605 vdd.n216 vdd.n183 585
R15606 vdd.n215 vdd.n214 585
R15607 vdd.n186 vdd.n184 585
R15608 vdd.n209 vdd.n208 585
R15609 vdd.n207 vdd.n206 585
R15610 vdd.n190 vdd.n189 585
R15611 vdd.n201 vdd.n200 585
R15612 vdd.n199 vdd.n198 585
R15613 vdd.n194 vdd.n193 585
R15614 vdd.n163 vdd.n162 585
R15615 vdd.n161 vdd.n128 585
R15616 vdd.n160 vdd.n159 585
R15617 vdd.n131 vdd.n129 585
R15618 vdd.n154 vdd.n153 585
R15619 vdd.n152 vdd.n151 585
R15620 vdd.n135 vdd.n134 585
R15621 vdd.n146 vdd.n145 585
R15622 vdd.n144 vdd.n143 585
R15623 vdd.n139 vdd.n138 585
R15624 vdd.n121 vdd.n120 585
R15625 vdd.n119 vdd.n86 585
R15626 vdd.n118 vdd.n117 585
R15627 vdd.n89 vdd.n87 585
R15628 vdd.n112 vdd.n111 585
R15629 vdd.n110 vdd.n109 585
R15630 vdd.n93 vdd.n92 585
R15631 vdd.n104 vdd.n103 585
R15632 vdd.n102 vdd.n101 585
R15633 vdd.n97 vdd.n96 585
R15634 vdd.n66 vdd.n65 585
R15635 vdd.n64 vdd.n31 585
R15636 vdd.n63 vdd.n62 585
R15637 vdd.n34 vdd.n32 585
R15638 vdd.n57 vdd.n56 585
R15639 vdd.n55 vdd.n54 585
R15640 vdd.n38 vdd.n37 585
R15641 vdd.n49 vdd.n48 585
R15642 vdd.n47 vdd.n46 585
R15643 vdd.n42 vdd.n41 585
R15644 vdd.n2047 vdd.n2046 585
R15645 vdd.n2045 vdd.n2012 585
R15646 vdd.n2044 vdd.n2043 585
R15647 vdd.n2015 vdd.n2013 585
R15648 vdd.n2038 vdd.n2037 585
R15649 vdd.n2036 vdd.n2035 585
R15650 vdd.n2019 vdd.n2018 585
R15651 vdd.n2030 vdd.n2029 585
R15652 vdd.n2028 vdd.n2027 585
R15653 vdd.n2023 vdd.n2022 585
R15654 vdd.n2102 vdd.n2101 585
R15655 vdd.n2100 vdd.n2067 585
R15656 vdd.n2099 vdd.n2098 585
R15657 vdd.n2070 vdd.n2068 585
R15658 vdd.n2093 vdd.n2092 585
R15659 vdd.n2091 vdd.n2090 585
R15660 vdd.n2074 vdd.n2073 585
R15661 vdd.n2085 vdd.n2084 585
R15662 vdd.n2083 vdd.n2082 585
R15663 vdd.n2078 vdd.n2077 585
R15664 vdd.n1949 vdd.n1948 585
R15665 vdd.n1947 vdd.n1914 585
R15666 vdd.n1946 vdd.n1945 585
R15667 vdd.n1917 vdd.n1915 585
R15668 vdd.n1940 vdd.n1939 585
R15669 vdd.n1938 vdd.n1937 585
R15670 vdd.n1921 vdd.n1920 585
R15671 vdd.n1932 vdd.n1931 585
R15672 vdd.n1930 vdd.n1929 585
R15673 vdd.n1925 vdd.n1924 585
R15674 vdd.n2004 vdd.n2003 585
R15675 vdd.n2002 vdd.n1969 585
R15676 vdd.n2001 vdd.n2000 585
R15677 vdd.n1972 vdd.n1970 585
R15678 vdd.n1995 vdd.n1994 585
R15679 vdd.n1993 vdd.n1992 585
R15680 vdd.n1976 vdd.n1975 585
R15681 vdd.n1987 vdd.n1986 585
R15682 vdd.n1985 vdd.n1984 585
R15683 vdd.n1980 vdd.n1979 585
R15684 vdd.n1852 vdd.n1851 585
R15685 vdd.n1850 vdd.n1817 585
R15686 vdd.n1849 vdd.n1848 585
R15687 vdd.n1820 vdd.n1818 585
R15688 vdd.n1843 vdd.n1842 585
R15689 vdd.n1841 vdd.n1840 585
R15690 vdd.n1824 vdd.n1823 585
R15691 vdd.n1835 vdd.n1834 585
R15692 vdd.n1833 vdd.n1832 585
R15693 vdd.n1828 vdd.n1827 585
R15694 vdd.n1907 vdd.n1906 585
R15695 vdd.n1905 vdd.n1872 585
R15696 vdd.n1904 vdd.n1903 585
R15697 vdd.n1875 vdd.n1873 585
R15698 vdd.n1898 vdd.n1897 585
R15699 vdd.n1896 vdd.n1895 585
R15700 vdd.n1879 vdd.n1878 585
R15701 vdd.n1890 vdd.n1889 585
R15702 vdd.n1888 vdd.n1887 585
R15703 vdd.n1883 vdd.n1882 585
R15704 vdd.n445 vdd.n370 462.44
R15705 vdd.n3343 vdd.n372 462.44
R15706 vdd.n3238 vdd.n657 462.44
R15707 vdd.n3236 vdd.n660 462.44
R15708 vdd.n2181 vdd.n1409 462.44
R15709 vdd.n2184 vdd.n2183 462.44
R15710 vdd.n1737 vdd.n1507 462.44
R15711 vdd.n1734 vdd.n1505 462.44
R15712 vdd.n293 vdd.t243 329.043
R15713 vdd.n238 vdd.t220 329.043
R15714 vdd.n195 vdd.t233 329.043
R15715 vdd.n140 vdd.t210 329.043
R15716 vdd.n98 vdd.t195 329.043
R15717 vdd.n43 vdd.t178 329.043
R15718 vdd.n2024 vdd.t254 329.043
R15719 vdd.n2079 vdd.t166 329.043
R15720 vdd.n1926 vdd.t246 329.043
R15721 vdd.n1981 vdd.t143 329.043
R15722 vdd.n1829 vdd.t173 329.043
R15723 vdd.n1884 vdd.t196 329.043
R15724 vdd.n1510 vdd.t88 319.788
R15725 vdd.n1666 vdd.t81 319.788
R15726 vdd.n1702 vdd.t91 319.788
R15727 vdd.n2186 vdd.t63 319.788
R15728 vdd.n1161 vdd.t93 319.788
R15729 vdd.n1121 vdd.t108 319.788
R15730 vdd.n405 vdd.t84 319.788
R15731 vdd.n419 vdd.t117 319.788
R15732 vdd.n431 vdd.t123 319.788
R15733 vdd.n723 vdd.t67 319.788
R15734 vdd.n686 vdd.t77 319.788
R15735 vdd.n3105 vdd.t60 319.788
R15736 vdd.n1511 vdd.t87 303.69
R15737 vdd.n1667 vdd.t80 303.69
R15738 vdd.n1703 vdd.t90 303.69
R15739 vdd.n2187 vdd.t64 303.69
R15740 vdd.n1162 vdd.t94 303.69
R15741 vdd.n1122 vdd.t109 303.69
R15742 vdd.n406 vdd.t85 303.69
R15743 vdd.n420 vdd.t118 303.69
R15744 vdd.n432 vdd.t124 303.69
R15745 vdd.n724 vdd.t66 303.69
R15746 vdd.n687 vdd.t76 303.69
R15747 vdd.n3106 vdd.t59 303.69
R15748 vdd.n2853 vdd.n898 291.221
R15749 vdd.n3067 vdd.n778 291.221
R15750 vdd.n3004 vdd.n775 291.221
R15751 vdd.n2785 vdd.n2784 291.221
R15752 vdd.n2581 vdd.n940 291.221
R15753 vdd.n2512 vdd.n2511 291.221
R15754 vdd.n1280 vdd.n1279 291.221
R15755 vdd.n2332 vdd.n1046 291.221
R15756 vdd.n2983 vdd.n776 291.221
R15757 vdd.n3070 vdd.n3069 291.221
R15758 vdd.n2689 vdd.n2615 291.221
R15759 vdd.n2857 vdd.n902 291.221
R15760 vdd.n2509 vdd.n950 291.221
R15761 vdd.n948 vdd.n922 291.221
R15762 vdd.n1358 vdd.n1087 291.221
R15763 vdd.n2336 vdd.n1051 291.221
R15764 vdd.n2985 vdd.n776 185
R15765 vdd.n3068 vdd.n776 185
R15766 vdd.n2987 vdd.n2986 185
R15767 vdd.n2986 vdd.n774 185
R15768 vdd.n2988 vdd.n810 185
R15769 vdd.n2998 vdd.n810 185
R15770 vdd.n2989 vdd.n819 185
R15771 vdd.n819 vdd.n817 185
R15772 vdd.n2991 vdd.n2990 185
R15773 vdd.n2992 vdd.n2991 185
R15774 vdd.n2944 vdd.n818 185
R15775 vdd.n818 vdd.n814 185
R15776 vdd.n2943 vdd.n2942 185
R15777 vdd.n2942 vdd.n2941 185
R15778 vdd.n821 vdd.n820 185
R15779 vdd.n822 vdd.n821 185
R15780 vdd.n2934 vdd.n2933 185
R15781 vdd.n2935 vdd.n2934 185
R15782 vdd.n2932 vdd.n831 185
R15783 vdd.n831 vdd.n828 185
R15784 vdd.n2931 vdd.n2930 185
R15785 vdd.n2930 vdd.n2929 185
R15786 vdd.n833 vdd.n832 185
R15787 vdd.n841 vdd.n833 185
R15788 vdd.n2922 vdd.n2921 185
R15789 vdd.n2923 vdd.n2922 185
R15790 vdd.n2919 vdd.n842 185
R15791 vdd.n849 vdd.n842 185
R15792 vdd.n2918 vdd.n2917 185
R15793 vdd.n2917 vdd.n2916 185
R15794 vdd.n845 vdd.n844 185
R15795 vdd.n846 vdd.n845 185
R15796 vdd.n2909 vdd.n2908 185
R15797 vdd.n2910 vdd.n2909 185
R15798 vdd.n2907 vdd.n856 185
R15799 vdd.n856 vdd.n853 185
R15800 vdd.n2906 vdd.n2905 185
R15801 vdd.n2905 vdd.n2904 185
R15802 vdd.n858 vdd.n857 185
R15803 vdd.n866 vdd.n858 185
R15804 vdd.n2897 vdd.n2896 185
R15805 vdd.n2898 vdd.n2897 185
R15806 vdd.n2895 vdd.n867 185
R15807 vdd.n872 vdd.n867 185
R15808 vdd.n2894 vdd.n2893 185
R15809 vdd.n2893 vdd.n2892 185
R15810 vdd.n869 vdd.n868 185
R15811 vdd.n2764 vdd.n869 185
R15812 vdd.n2885 vdd.n2884 185
R15813 vdd.n2886 vdd.n2885 185
R15814 vdd.n2883 vdd.n879 185
R15815 vdd.n879 vdd.n876 185
R15816 vdd.n2882 vdd.n2881 185
R15817 vdd.n2881 vdd.n2880 185
R15818 vdd.n881 vdd.n880 185
R15819 vdd.n882 vdd.n881 185
R15820 vdd.n2873 vdd.n2872 185
R15821 vdd.n2874 vdd.n2873 185
R15822 vdd.n2871 vdd.n891 185
R15823 vdd.n891 vdd.n888 185
R15824 vdd.n2870 vdd.n2869 185
R15825 vdd.n2869 vdd.n2868 185
R15826 vdd.n893 vdd.n892 185
R15827 vdd.n2779 vdd.n893 185
R15828 vdd.n2861 vdd.n2860 185
R15829 vdd.n2862 vdd.n2861 185
R15830 vdd.n2859 vdd.n902 185
R15831 vdd.n902 vdd.n899 185
R15832 vdd.n2858 vdd.n2857 185
R15833 vdd.n904 vdd.n903 185
R15834 vdd.n2625 vdd.n2624 185
R15835 vdd.n2627 vdd.n2626 185
R15836 vdd.n2629 vdd.n2628 185
R15837 vdd.n2631 vdd.n2630 185
R15838 vdd.n2633 vdd.n2632 185
R15839 vdd.n2635 vdd.n2634 185
R15840 vdd.n2637 vdd.n2636 185
R15841 vdd.n2639 vdd.n2638 185
R15842 vdd.n2641 vdd.n2640 185
R15843 vdd.n2643 vdd.n2642 185
R15844 vdd.n2645 vdd.n2644 185
R15845 vdd.n2647 vdd.n2646 185
R15846 vdd.n2649 vdd.n2648 185
R15847 vdd.n2651 vdd.n2650 185
R15848 vdd.n2653 vdd.n2652 185
R15849 vdd.n2655 vdd.n2654 185
R15850 vdd.n2657 vdd.n2656 185
R15851 vdd.n2659 vdd.n2658 185
R15852 vdd.n2661 vdd.n2660 185
R15853 vdd.n2663 vdd.n2662 185
R15854 vdd.n2665 vdd.n2664 185
R15855 vdd.n2667 vdd.n2666 185
R15856 vdd.n2669 vdd.n2668 185
R15857 vdd.n2671 vdd.n2670 185
R15858 vdd.n2673 vdd.n2672 185
R15859 vdd.n2675 vdd.n2674 185
R15860 vdd.n2677 vdd.n2676 185
R15861 vdd.n2679 vdd.n2678 185
R15862 vdd.n2681 vdd.n2680 185
R15863 vdd.n2683 vdd.n2682 185
R15864 vdd.n2685 vdd.n2684 185
R15865 vdd.n2687 vdd.n2686 185
R15866 vdd.n2688 vdd.n2615 185
R15867 vdd.n2855 vdd.n2615 185
R15868 vdd.n3071 vdd.n3070 185
R15869 vdd.n3072 vdd.n767 185
R15870 vdd.n3074 vdd.n3073 185
R15871 vdd.n3076 vdd.n765 185
R15872 vdd.n3078 vdd.n3077 185
R15873 vdd.n3079 vdd.n764 185
R15874 vdd.n3081 vdd.n3080 185
R15875 vdd.n3083 vdd.n762 185
R15876 vdd.n3085 vdd.n3084 185
R15877 vdd.n3086 vdd.n761 185
R15878 vdd.n3088 vdd.n3087 185
R15879 vdd.n3090 vdd.n759 185
R15880 vdd.n3092 vdd.n3091 185
R15881 vdd.n3093 vdd.n758 185
R15882 vdd.n3095 vdd.n3094 185
R15883 vdd.n3097 vdd.n757 185
R15884 vdd.n3098 vdd.n754 185
R15885 vdd.n3101 vdd.n3100 185
R15886 vdd.n755 vdd.n753 185
R15887 vdd.n2957 vdd.n2956 185
R15888 vdd.n2959 vdd.n2958 185
R15889 vdd.n2961 vdd.n2953 185
R15890 vdd.n2963 vdd.n2962 185
R15891 vdd.n2964 vdd.n2952 185
R15892 vdd.n2966 vdd.n2965 185
R15893 vdd.n2968 vdd.n2950 185
R15894 vdd.n2970 vdd.n2969 185
R15895 vdd.n2971 vdd.n2949 185
R15896 vdd.n2973 vdd.n2972 185
R15897 vdd.n2975 vdd.n2947 185
R15898 vdd.n2977 vdd.n2976 185
R15899 vdd.n2978 vdd.n2946 185
R15900 vdd.n2980 vdd.n2979 185
R15901 vdd.n2982 vdd.n2945 185
R15902 vdd.n2984 vdd.n2983 185
R15903 vdd.n2983 vdd.n756 185
R15904 vdd.n3069 vdd.n771 185
R15905 vdd.n3069 vdd.n3068 185
R15906 vdd.n2692 vdd.n773 185
R15907 vdd.n774 vdd.n773 185
R15908 vdd.n2693 vdd.n809 185
R15909 vdd.n2998 vdd.n809 185
R15910 vdd.n2695 vdd.n2694 185
R15911 vdd.n2694 vdd.n817 185
R15912 vdd.n2696 vdd.n816 185
R15913 vdd.n2992 vdd.n816 185
R15914 vdd.n2698 vdd.n2697 185
R15915 vdd.n2697 vdd.n814 185
R15916 vdd.n2699 vdd.n824 185
R15917 vdd.n2941 vdd.n824 185
R15918 vdd.n2701 vdd.n2700 185
R15919 vdd.n2700 vdd.n822 185
R15920 vdd.n2702 vdd.n830 185
R15921 vdd.n2935 vdd.n830 185
R15922 vdd.n2704 vdd.n2703 185
R15923 vdd.n2703 vdd.n828 185
R15924 vdd.n2705 vdd.n835 185
R15925 vdd.n2929 vdd.n835 185
R15926 vdd.n2707 vdd.n2706 185
R15927 vdd.n2706 vdd.n841 185
R15928 vdd.n2708 vdd.n840 185
R15929 vdd.n2923 vdd.n840 185
R15930 vdd.n2710 vdd.n2709 185
R15931 vdd.n2709 vdd.n849 185
R15932 vdd.n2711 vdd.n848 185
R15933 vdd.n2916 vdd.n848 185
R15934 vdd.n2713 vdd.n2712 185
R15935 vdd.n2712 vdd.n846 185
R15936 vdd.n2714 vdd.n855 185
R15937 vdd.n2910 vdd.n855 185
R15938 vdd.n2716 vdd.n2715 185
R15939 vdd.n2715 vdd.n853 185
R15940 vdd.n2717 vdd.n860 185
R15941 vdd.n2904 vdd.n860 185
R15942 vdd.n2719 vdd.n2718 185
R15943 vdd.n2718 vdd.n866 185
R15944 vdd.n2720 vdd.n865 185
R15945 vdd.n2898 vdd.n865 185
R15946 vdd.n2722 vdd.n2721 185
R15947 vdd.n2721 vdd.n872 185
R15948 vdd.n2723 vdd.n871 185
R15949 vdd.n2892 vdd.n871 185
R15950 vdd.n2766 vdd.n2765 185
R15951 vdd.n2765 vdd.n2764 185
R15952 vdd.n2767 vdd.n878 185
R15953 vdd.n2886 vdd.n878 185
R15954 vdd.n2769 vdd.n2768 185
R15955 vdd.n2768 vdd.n876 185
R15956 vdd.n2770 vdd.n884 185
R15957 vdd.n2880 vdd.n884 185
R15958 vdd.n2772 vdd.n2771 185
R15959 vdd.n2771 vdd.n882 185
R15960 vdd.n2773 vdd.n890 185
R15961 vdd.n2874 vdd.n890 185
R15962 vdd.n2775 vdd.n2774 185
R15963 vdd.n2774 vdd.n888 185
R15964 vdd.n2776 vdd.n895 185
R15965 vdd.n2868 vdd.n895 185
R15966 vdd.n2778 vdd.n2777 185
R15967 vdd.n2779 vdd.n2778 185
R15968 vdd.n2691 vdd.n901 185
R15969 vdd.n2862 vdd.n901 185
R15970 vdd.n2690 vdd.n2689 185
R15971 vdd.n2689 vdd.n899 185
R15972 vdd.n2181 vdd.n2180 185
R15973 vdd.n2182 vdd.n2181 185
R15974 vdd.n1410 vdd.n1408 185
R15975 vdd.n1408 vdd.n1407 185
R15976 vdd.n2176 vdd.n2175 185
R15977 vdd.n2175 vdd.n2174 185
R15978 vdd.n1413 vdd.n1412 185
R15979 vdd.n1414 vdd.n1413 185
R15980 vdd.n2163 vdd.n2162 185
R15981 vdd.n2164 vdd.n2163 185
R15982 vdd.n1422 vdd.n1421 185
R15983 vdd.n2155 vdd.n1421 185
R15984 vdd.n2158 vdd.n2157 185
R15985 vdd.n2157 vdd.n2156 185
R15986 vdd.n1425 vdd.n1424 185
R15987 vdd.n1431 vdd.n1425 185
R15988 vdd.n2146 vdd.n2145 185
R15989 vdd.n2147 vdd.n2146 185
R15990 vdd.n1433 vdd.n1432 185
R15991 vdd.n2138 vdd.n1432 185
R15992 vdd.n2141 vdd.n2140 185
R15993 vdd.n2140 vdd.n2139 185
R15994 vdd.n1436 vdd.n1435 185
R15995 vdd.n1437 vdd.n1436 185
R15996 vdd.n2129 vdd.n2128 185
R15997 vdd.n2130 vdd.n2129 185
R15998 vdd.n1445 vdd.n1444 185
R15999 vdd.n1444 vdd.n1443 185
R16000 vdd.n2124 vdd.n2123 185
R16001 vdd.n2123 vdd.n2122 185
R16002 vdd.n1448 vdd.n1447 185
R16003 vdd.n1454 vdd.n1448 185
R16004 vdd.n2113 vdd.n2112 185
R16005 vdd.n2114 vdd.n2113 185
R16006 vdd.n1456 vdd.n1455 185
R16007 vdd.n1810 vdd.n1455 185
R16008 vdd.n1813 vdd.n1812 185
R16009 vdd.n1812 vdd.n1811 185
R16010 vdd.n1459 vdd.n1458 185
R16011 vdd.n1466 vdd.n1459 185
R16012 vdd.n1801 vdd.n1800 185
R16013 vdd.n1802 vdd.n1801 185
R16014 vdd.n1468 vdd.n1467 185
R16015 vdd.n1467 vdd.n1465 185
R16016 vdd.n1796 vdd.n1795 185
R16017 vdd.n1795 vdd.n1794 185
R16018 vdd.n1471 vdd.n1470 185
R16019 vdd.n1472 vdd.n1471 185
R16020 vdd.n1785 vdd.n1784 185
R16021 vdd.n1786 vdd.n1785 185
R16022 vdd.n1479 vdd.n1478 185
R16023 vdd.n1777 vdd.n1478 185
R16024 vdd.n1780 vdd.n1779 185
R16025 vdd.n1779 vdd.n1778 185
R16026 vdd.n1482 vdd.n1481 185
R16027 vdd.n1488 vdd.n1482 185
R16028 vdd.n1768 vdd.n1767 185
R16029 vdd.n1769 vdd.n1768 185
R16030 vdd.n1490 vdd.n1489 185
R16031 vdd.n1760 vdd.n1489 185
R16032 vdd.n1763 vdd.n1762 185
R16033 vdd.n1762 vdd.n1761 185
R16034 vdd.n1493 vdd.n1492 185
R16035 vdd.n1494 vdd.n1493 185
R16036 vdd.n1751 vdd.n1750 185
R16037 vdd.n1752 vdd.n1751 185
R16038 vdd.n1502 vdd.n1501 185
R16039 vdd.n1501 vdd.n1500 185
R16040 vdd.n1746 vdd.n1745 185
R16041 vdd.n1745 vdd.n1744 185
R16042 vdd.n1505 vdd.n1504 185
R16043 vdd.n1506 vdd.n1505 185
R16044 vdd.n1734 vdd.n1733 185
R16045 vdd.n1732 vdd.n1545 185
R16046 vdd.n1547 vdd.n1544 185
R16047 vdd.n1736 vdd.n1544 185
R16048 vdd.n1728 vdd.n1549 185
R16049 vdd.n1727 vdd.n1550 185
R16050 vdd.n1726 vdd.n1551 185
R16051 vdd.n1554 vdd.n1552 185
R16052 vdd.n1722 vdd.n1555 185
R16053 vdd.n1721 vdd.n1556 185
R16054 vdd.n1720 vdd.n1557 185
R16055 vdd.n1560 vdd.n1558 185
R16056 vdd.n1716 vdd.n1561 185
R16057 vdd.n1715 vdd.n1562 185
R16058 vdd.n1714 vdd.n1563 185
R16059 vdd.n1566 vdd.n1564 185
R16060 vdd.n1710 vdd.n1567 185
R16061 vdd.n1709 vdd.n1568 185
R16062 vdd.n1708 vdd.n1569 185
R16063 vdd.n1700 vdd.n1570 185
R16064 vdd.n1704 vdd.n1701 185
R16065 vdd.n1699 vdd.n1572 185
R16066 vdd.n1698 vdd.n1573 185
R16067 vdd.n1576 vdd.n1574 185
R16068 vdd.n1694 vdd.n1577 185
R16069 vdd.n1693 vdd.n1578 185
R16070 vdd.n1692 vdd.n1579 185
R16071 vdd.n1582 vdd.n1580 185
R16072 vdd.n1688 vdd.n1583 185
R16073 vdd.n1687 vdd.n1584 185
R16074 vdd.n1686 vdd.n1585 185
R16075 vdd.n1588 vdd.n1586 185
R16076 vdd.n1682 vdd.n1589 185
R16077 vdd.n1681 vdd.n1590 185
R16078 vdd.n1680 vdd.n1591 185
R16079 vdd.n1594 vdd.n1592 185
R16080 vdd.n1676 vdd.n1595 185
R16081 vdd.n1675 vdd.n1596 185
R16082 vdd.n1674 vdd.n1597 185
R16083 vdd.n1600 vdd.n1598 185
R16084 vdd.n1670 vdd.n1601 185
R16085 vdd.n1669 vdd.n1602 185
R16086 vdd.n1668 vdd.n1665 185
R16087 vdd.n1605 vdd.n1603 185
R16088 vdd.n1661 vdd.n1606 185
R16089 vdd.n1660 vdd.n1607 185
R16090 vdd.n1659 vdd.n1608 185
R16091 vdd.n1611 vdd.n1609 185
R16092 vdd.n1655 vdd.n1612 185
R16093 vdd.n1654 vdd.n1613 185
R16094 vdd.n1653 vdd.n1614 185
R16095 vdd.n1617 vdd.n1615 185
R16096 vdd.n1649 vdd.n1618 185
R16097 vdd.n1648 vdd.n1619 185
R16098 vdd.n1647 vdd.n1620 185
R16099 vdd.n1623 vdd.n1621 185
R16100 vdd.n1643 vdd.n1624 185
R16101 vdd.n1642 vdd.n1625 185
R16102 vdd.n1641 vdd.n1626 185
R16103 vdd.n1629 vdd.n1627 185
R16104 vdd.n1637 vdd.n1630 185
R16105 vdd.n1636 vdd.n1631 185
R16106 vdd.n1635 vdd.n1632 185
R16107 vdd.n1633 vdd.n1513 185
R16108 vdd.n1738 vdd.n1737 185
R16109 vdd.n1737 vdd.n1736 185
R16110 vdd.n2185 vdd.n2184 185
R16111 vdd.n2189 vdd.n1403 185
R16112 vdd.n1402 vdd.n1396 185
R16113 vdd.n1400 vdd.n1399 185
R16114 vdd.n1398 vdd.n1192 185
R16115 vdd.n2193 vdd.n1189 185
R16116 vdd.n2195 vdd.n2194 185
R16117 vdd.n2197 vdd.n1187 185
R16118 vdd.n2199 vdd.n2198 185
R16119 vdd.n2200 vdd.n1182 185
R16120 vdd.n2202 vdd.n2201 185
R16121 vdd.n2204 vdd.n1180 185
R16122 vdd.n2206 vdd.n2205 185
R16123 vdd.n2207 vdd.n1175 185
R16124 vdd.n2209 vdd.n2208 185
R16125 vdd.n2211 vdd.n1173 185
R16126 vdd.n2213 vdd.n2212 185
R16127 vdd.n2214 vdd.n1169 185
R16128 vdd.n2216 vdd.n2215 185
R16129 vdd.n2218 vdd.n1166 185
R16130 vdd.n2220 vdd.n2219 185
R16131 vdd.n1167 vdd.n1160 185
R16132 vdd.n2224 vdd.n1164 185
R16133 vdd.n2225 vdd.n1156 185
R16134 vdd.n2227 vdd.n2226 185
R16135 vdd.n2229 vdd.n1154 185
R16136 vdd.n2231 vdd.n2230 185
R16137 vdd.n2232 vdd.n1149 185
R16138 vdd.n2234 vdd.n2233 185
R16139 vdd.n2236 vdd.n1147 185
R16140 vdd.n2238 vdd.n2237 185
R16141 vdd.n2239 vdd.n1142 185
R16142 vdd.n2241 vdd.n2240 185
R16143 vdd.n2243 vdd.n1140 185
R16144 vdd.n2245 vdd.n2244 185
R16145 vdd.n2246 vdd.n1135 185
R16146 vdd.n2248 vdd.n2247 185
R16147 vdd.n2250 vdd.n1133 185
R16148 vdd.n2252 vdd.n2251 185
R16149 vdd.n2253 vdd.n1129 185
R16150 vdd.n2255 vdd.n2254 185
R16151 vdd.n2257 vdd.n1126 185
R16152 vdd.n2259 vdd.n2258 185
R16153 vdd.n1127 vdd.n1120 185
R16154 vdd.n2263 vdd.n1124 185
R16155 vdd.n2264 vdd.n1116 185
R16156 vdd.n2266 vdd.n2265 185
R16157 vdd.n2268 vdd.n1114 185
R16158 vdd.n2270 vdd.n2269 185
R16159 vdd.n2271 vdd.n1109 185
R16160 vdd.n2273 vdd.n2272 185
R16161 vdd.n2275 vdd.n1107 185
R16162 vdd.n2277 vdd.n2276 185
R16163 vdd.n2278 vdd.n1102 185
R16164 vdd.n2280 vdd.n2279 185
R16165 vdd.n2282 vdd.n1100 185
R16166 vdd.n2284 vdd.n2283 185
R16167 vdd.n2285 vdd.n1098 185
R16168 vdd.n2287 vdd.n2286 185
R16169 vdd.n2290 vdd.n2289 185
R16170 vdd.n2292 vdd.n2291 185
R16171 vdd.n2294 vdd.n1096 185
R16172 vdd.n2296 vdd.n2295 185
R16173 vdd.n1409 vdd.n1095 185
R16174 vdd.n2183 vdd.n1406 185
R16175 vdd.n2183 vdd.n2182 185
R16176 vdd.n1417 vdd.n1405 185
R16177 vdd.n1407 vdd.n1405 185
R16178 vdd.n2173 vdd.n2172 185
R16179 vdd.n2174 vdd.n2173 185
R16180 vdd.n1416 vdd.n1415 185
R16181 vdd.n1415 vdd.n1414 185
R16182 vdd.n2166 vdd.n2165 185
R16183 vdd.n2165 vdd.n2164 185
R16184 vdd.n1420 vdd.n1419 185
R16185 vdd.n2155 vdd.n1420 185
R16186 vdd.n2154 vdd.n2153 185
R16187 vdd.n2156 vdd.n2154 185
R16188 vdd.n1427 vdd.n1426 185
R16189 vdd.n1431 vdd.n1426 185
R16190 vdd.n2149 vdd.n2148 185
R16191 vdd.n2148 vdd.n2147 185
R16192 vdd.n1430 vdd.n1429 185
R16193 vdd.n2138 vdd.n1430 185
R16194 vdd.n2137 vdd.n2136 185
R16195 vdd.n2139 vdd.n2137 185
R16196 vdd.n1439 vdd.n1438 185
R16197 vdd.n1438 vdd.n1437 185
R16198 vdd.n2132 vdd.n2131 185
R16199 vdd.n2131 vdd.n2130 185
R16200 vdd.n1442 vdd.n1441 185
R16201 vdd.n1443 vdd.n1442 185
R16202 vdd.n2121 vdd.n2120 185
R16203 vdd.n2122 vdd.n2121 185
R16204 vdd.n1450 vdd.n1449 185
R16205 vdd.n1454 vdd.n1449 185
R16206 vdd.n2116 vdd.n2115 185
R16207 vdd.n2115 vdd.n2114 185
R16208 vdd.n1453 vdd.n1452 185
R16209 vdd.n1810 vdd.n1453 185
R16210 vdd.n1809 vdd.n1808 185
R16211 vdd.n1811 vdd.n1809 185
R16212 vdd.n1461 vdd.n1460 185
R16213 vdd.n1466 vdd.n1460 185
R16214 vdd.n1804 vdd.n1803 185
R16215 vdd.n1803 vdd.n1802 185
R16216 vdd.n1464 vdd.n1463 185
R16217 vdd.n1465 vdd.n1464 185
R16218 vdd.n1793 vdd.n1792 185
R16219 vdd.n1794 vdd.n1793 185
R16220 vdd.n1474 vdd.n1473 185
R16221 vdd.n1473 vdd.n1472 185
R16222 vdd.n1788 vdd.n1787 185
R16223 vdd.n1787 vdd.n1786 185
R16224 vdd.n1477 vdd.n1476 185
R16225 vdd.n1777 vdd.n1477 185
R16226 vdd.n1776 vdd.n1775 185
R16227 vdd.n1778 vdd.n1776 185
R16228 vdd.n1484 vdd.n1483 185
R16229 vdd.n1488 vdd.n1483 185
R16230 vdd.n1771 vdd.n1770 185
R16231 vdd.n1770 vdd.n1769 185
R16232 vdd.n1487 vdd.n1486 185
R16233 vdd.n1760 vdd.n1487 185
R16234 vdd.n1759 vdd.n1758 185
R16235 vdd.n1761 vdd.n1759 185
R16236 vdd.n1496 vdd.n1495 185
R16237 vdd.n1495 vdd.n1494 185
R16238 vdd.n1754 vdd.n1753 185
R16239 vdd.n1753 vdd.n1752 185
R16240 vdd.n1499 vdd.n1498 185
R16241 vdd.n1500 vdd.n1499 185
R16242 vdd.n1743 vdd.n1742 185
R16243 vdd.n1744 vdd.n1743 185
R16244 vdd.n1508 vdd.n1507 185
R16245 vdd.n1507 vdd.n1506 185
R16246 vdd.n942 vdd.n940 185
R16247 vdd.n2510 vdd.n940 185
R16248 vdd.n2432 vdd.n960 185
R16249 vdd.n960 vdd.n947 185
R16250 vdd.n2434 vdd.n2433 185
R16251 vdd.n2435 vdd.n2434 185
R16252 vdd.n2431 vdd.n959 185
R16253 vdd.n1309 vdd.n959 185
R16254 vdd.n2430 vdd.n2429 185
R16255 vdd.n2429 vdd.n2428 185
R16256 vdd.n962 vdd.n961 185
R16257 vdd.n963 vdd.n962 185
R16258 vdd.n2419 vdd.n2418 185
R16259 vdd.n2420 vdd.n2419 185
R16260 vdd.n2417 vdd.n973 185
R16261 vdd.n973 vdd.n970 185
R16262 vdd.n2416 vdd.n2415 185
R16263 vdd.n2415 vdd.n2414 185
R16264 vdd.n975 vdd.n974 185
R16265 vdd.n976 vdd.n975 185
R16266 vdd.n2407 vdd.n2406 185
R16267 vdd.n2408 vdd.n2407 185
R16268 vdd.n2405 vdd.n984 185
R16269 vdd.n989 vdd.n984 185
R16270 vdd.n2404 vdd.n2403 185
R16271 vdd.n2403 vdd.n2402 185
R16272 vdd.n986 vdd.n985 185
R16273 vdd.n995 vdd.n986 185
R16274 vdd.n2395 vdd.n2394 185
R16275 vdd.n2396 vdd.n2395 185
R16276 vdd.n2393 vdd.n996 185
R16277 vdd.n1330 vdd.n996 185
R16278 vdd.n2392 vdd.n2391 185
R16279 vdd.n2391 vdd.n2390 185
R16280 vdd.n998 vdd.n997 185
R16281 vdd.n999 vdd.n998 185
R16282 vdd.n2383 vdd.n2382 185
R16283 vdd.n2384 vdd.n2383 185
R16284 vdd.n2381 vdd.n1008 185
R16285 vdd.n1008 vdd.n1005 185
R16286 vdd.n2380 vdd.n2379 185
R16287 vdd.n2379 vdd.n2378 185
R16288 vdd.n1010 vdd.n1009 185
R16289 vdd.n1019 vdd.n1010 185
R16290 vdd.n2370 vdd.n2369 185
R16291 vdd.n2371 vdd.n2370 185
R16292 vdd.n2368 vdd.n1020 185
R16293 vdd.n1026 vdd.n1020 185
R16294 vdd.n2367 vdd.n2366 185
R16295 vdd.n2366 vdd.n2365 185
R16296 vdd.n1022 vdd.n1021 185
R16297 vdd.n1023 vdd.n1022 185
R16298 vdd.n2358 vdd.n2357 185
R16299 vdd.n2359 vdd.n2358 185
R16300 vdd.n2356 vdd.n1033 185
R16301 vdd.n1033 vdd.n1030 185
R16302 vdd.n2355 vdd.n2354 185
R16303 vdd.n2354 vdd.n2353 185
R16304 vdd.n1035 vdd.n1034 185
R16305 vdd.n1036 vdd.n1035 185
R16306 vdd.n2346 vdd.n2345 185
R16307 vdd.n2347 vdd.n2346 185
R16308 vdd.n2344 vdd.n1044 185
R16309 vdd.n1050 vdd.n1044 185
R16310 vdd.n2343 vdd.n2342 185
R16311 vdd.n2342 vdd.n2341 185
R16312 vdd.n1046 vdd.n1045 185
R16313 vdd.n1047 vdd.n1046 185
R16314 vdd.n2332 vdd.n2331 185
R16315 vdd.n2330 vdd.n1089 185
R16316 vdd.n2329 vdd.n1088 185
R16317 vdd.n2334 vdd.n1088 185
R16318 vdd.n2328 vdd.n2327 185
R16319 vdd.n2326 vdd.n2325 185
R16320 vdd.n2324 vdd.n2323 185
R16321 vdd.n2322 vdd.n2321 185
R16322 vdd.n2320 vdd.n2319 185
R16323 vdd.n2318 vdd.n2317 185
R16324 vdd.n2316 vdd.n2315 185
R16325 vdd.n2314 vdd.n2313 185
R16326 vdd.n2312 vdd.n2311 185
R16327 vdd.n2310 vdd.n2309 185
R16328 vdd.n2308 vdd.n2307 185
R16329 vdd.n2306 vdd.n2305 185
R16330 vdd.n2304 vdd.n2303 185
R16331 vdd.n2302 vdd.n2301 185
R16332 vdd.n2300 vdd.n2299 185
R16333 vdd.n1246 vdd.n1090 185
R16334 vdd.n1248 vdd.n1247 185
R16335 vdd.n1250 vdd.n1249 185
R16336 vdd.n1252 vdd.n1251 185
R16337 vdd.n1254 vdd.n1253 185
R16338 vdd.n1256 vdd.n1255 185
R16339 vdd.n1258 vdd.n1257 185
R16340 vdd.n1260 vdd.n1259 185
R16341 vdd.n1262 vdd.n1261 185
R16342 vdd.n1264 vdd.n1263 185
R16343 vdd.n1266 vdd.n1265 185
R16344 vdd.n1268 vdd.n1267 185
R16345 vdd.n1270 vdd.n1269 185
R16346 vdd.n1272 vdd.n1271 185
R16347 vdd.n1275 vdd.n1274 185
R16348 vdd.n1277 vdd.n1276 185
R16349 vdd.n1279 vdd.n1278 185
R16350 vdd.n2513 vdd.n2512 185
R16351 vdd.n2515 vdd.n2514 185
R16352 vdd.n2517 vdd.n2516 185
R16353 vdd.n2520 vdd.n2519 185
R16354 vdd.n2522 vdd.n2521 185
R16355 vdd.n2524 vdd.n2523 185
R16356 vdd.n2526 vdd.n2525 185
R16357 vdd.n2528 vdd.n2527 185
R16358 vdd.n2530 vdd.n2529 185
R16359 vdd.n2532 vdd.n2531 185
R16360 vdd.n2534 vdd.n2533 185
R16361 vdd.n2536 vdd.n2535 185
R16362 vdd.n2538 vdd.n2537 185
R16363 vdd.n2540 vdd.n2539 185
R16364 vdd.n2542 vdd.n2541 185
R16365 vdd.n2544 vdd.n2543 185
R16366 vdd.n2546 vdd.n2545 185
R16367 vdd.n2548 vdd.n2547 185
R16368 vdd.n2550 vdd.n2549 185
R16369 vdd.n2552 vdd.n2551 185
R16370 vdd.n2554 vdd.n2553 185
R16371 vdd.n2556 vdd.n2555 185
R16372 vdd.n2558 vdd.n2557 185
R16373 vdd.n2560 vdd.n2559 185
R16374 vdd.n2562 vdd.n2561 185
R16375 vdd.n2564 vdd.n2563 185
R16376 vdd.n2566 vdd.n2565 185
R16377 vdd.n2568 vdd.n2567 185
R16378 vdd.n2570 vdd.n2569 185
R16379 vdd.n2572 vdd.n2571 185
R16380 vdd.n2574 vdd.n2573 185
R16381 vdd.n2576 vdd.n2575 185
R16382 vdd.n2578 vdd.n2577 185
R16383 vdd.n2579 vdd.n941 185
R16384 vdd.n2581 vdd.n2580 185
R16385 vdd.n2582 vdd.n2581 185
R16386 vdd.n2511 vdd.n945 185
R16387 vdd.n2511 vdd.n2510 185
R16388 vdd.n1307 vdd.n946 185
R16389 vdd.n947 vdd.n946 185
R16390 vdd.n1308 vdd.n957 185
R16391 vdd.n2435 vdd.n957 185
R16392 vdd.n1311 vdd.n1310 185
R16393 vdd.n1310 vdd.n1309 185
R16394 vdd.n1312 vdd.n964 185
R16395 vdd.n2428 vdd.n964 185
R16396 vdd.n1314 vdd.n1313 185
R16397 vdd.n1313 vdd.n963 185
R16398 vdd.n1315 vdd.n971 185
R16399 vdd.n2420 vdd.n971 185
R16400 vdd.n1317 vdd.n1316 185
R16401 vdd.n1316 vdd.n970 185
R16402 vdd.n1318 vdd.n977 185
R16403 vdd.n2414 vdd.n977 185
R16404 vdd.n1320 vdd.n1319 185
R16405 vdd.n1319 vdd.n976 185
R16406 vdd.n1321 vdd.n982 185
R16407 vdd.n2408 vdd.n982 185
R16408 vdd.n1323 vdd.n1322 185
R16409 vdd.n1322 vdd.n989 185
R16410 vdd.n1324 vdd.n987 185
R16411 vdd.n2402 vdd.n987 185
R16412 vdd.n1326 vdd.n1325 185
R16413 vdd.n1325 vdd.n995 185
R16414 vdd.n1327 vdd.n993 185
R16415 vdd.n2396 vdd.n993 185
R16416 vdd.n1329 vdd.n1328 185
R16417 vdd.n1330 vdd.n1329 185
R16418 vdd.n1306 vdd.n1000 185
R16419 vdd.n2390 vdd.n1000 185
R16420 vdd.n1305 vdd.n1304 185
R16421 vdd.n1304 vdd.n999 185
R16422 vdd.n1303 vdd.n1006 185
R16423 vdd.n2384 vdd.n1006 185
R16424 vdd.n1302 vdd.n1301 185
R16425 vdd.n1301 vdd.n1005 185
R16426 vdd.n1300 vdd.n1011 185
R16427 vdd.n2378 vdd.n1011 185
R16428 vdd.n1299 vdd.n1298 185
R16429 vdd.n1298 vdd.n1019 185
R16430 vdd.n1297 vdd.n1017 185
R16431 vdd.n2371 vdd.n1017 185
R16432 vdd.n1296 vdd.n1295 185
R16433 vdd.n1295 vdd.n1026 185
R16434 vdd.n1294 vdd.n1024 185
R16435 vdd.n2365 vdd.n1024 185
R16436 vdd.n1293 vdd.n1292 185
R16437 vdd.n1292 vdd.n1023 185
R16438 vdd.n1291 vdd.n1031 185
R16439 vdd.n2359 vdd.n1031 185
R16440 vdd.n1290 vdd.n1289 185
R16441 vdd.n1289 vdd.n1030 185
R16442 vdd.n1288 vdd.n1037 185
R16443 vdd.n2353 vdd.n1037 185
R16444 vdd.n1287 vdd.n1286 185
R16445 vdd.n1286 vdd.n1036 185
R16446 vdd.n1285 vdd.n1042 185
R16447 vdd.n2347 vdd.n1042 185
R16448 vdd.n1284 vdd.n1283 185
R16449 vdd.n1283 vdd.n1050 185
R16450 vdd.n1282 vdd.n1048 185
R16451 vdd.n2341 vdd.n1048 185
R16452 vdd.n1281 vdd.n1280 185
R16453 vdd.n1280 vdd.n1047 185
R16454 vdd.n370 vdd.n369 185
R16455 vdd.n3346 vdd.n370 185
R16456 vdd.n3349 vdd.n3348 185
R16457 vdd.n3348 vdd.n3347 185
R16458 vdd.n3350 vdd.n364 185
R16459 vdd.n364 vdd.n363 185
R16460 vdd.n3352 vdd.n3351 185
R16461 vdd.n3353 vdd.n3352 185
R16462 vdd.n359 vdd.n358 185
R16463 vdd.n3354 vdd.n359 185
R16464 vdd.n3357 vdd.n3356 185
R16465 vdd.n3356 vdd.n3355 185
R16466 vdd.n3358 vdd.n353 185
R16467 vdd.n3328 vdd.n353 185
R16468 vdd.n3360 vdd.n3359 185
R16469 vdd.n3361 vdd.n3360 185
R16470 vdd.n348 vdd.n347 185
R16471 vdd.n3362 vdd.n348 185
R16472 vdd.n3365 vdd.n3364 185
R16473 vdd.n3364 vdd.n3363 185
R16474 vdd.n3366 vdd.n342 185
R16475 vdd.n349 vdd.n342 185
R16476 vdd.n3368 vdd.n3367 185
R16477 vdd.n3369 vdd.n3368 185
R16478 vdd.n338 vdd.n337 185
R16479 vdd.n3370 vdd.n338 185
R16480 vdd.n3373 vdd.n3372 185
R16481 vdd.n3372 vdd.n3371 185
R16482 vdd.n3374 vdd.n333 185
R16483 vdd.n333 vdd.n332 185
R16484 vdd.n3376 vdd.n3375 185
R16485 vdd.n3377 vdd.n3376 185
R16486 vdd.n327 vdd.n325 185
R16487 vdd.n3378 vdd.n327 185
R16488 vdd.n3381 vdd.n3380 185
R16489 vdd.n3380 vdd.n3379 185
R16490 vdd.n326 vdd.n324 185
R16491 vdd.n328 vdd.n326 185
R16492 vdd.n3304 vdd.n3303 185
R16493 vdd.n3305 vdd.n3304 185
R16494 vdd.n615 vdd.n614 185
R16495 vdd.n614 vdd.n613 185
R16496 vdd.n3299 vdd.n3298 185
R16497 vdd.n3298 vdd.n3297 185
R16498 vdd.n618 vdd.n617 185
R16499 vdd.n624 vdd.n618 185
R16500 vdd.n3285 vdd.n3284 185
R16501 vdd.n3286 vdd.n3285 185
R16502 vdd.n626 vdd.n625 185
R16503 vdd.n3277 vdd.n625 185
R16504 vdd.n3280 vdd.n3279 185
R16505 vdd.n3279 vdd.n3278 185
R16506 vdd.n629 vdd.n628 185
R16507 vdd.n636 vdd.n629 185
R16508 vdd.n3268 vdd.n3267 185
R16509 vdd.n3269 vdd.n3268 185
R16510 vdd.n638 vdd.n637 185
R16511 vdd.n637 vdd.n635 185
R16512 vdd.n3263 vdd.n3262 185
R16513 vdd.n3262 vdd.n3261 185
R16514 vdd.n641 vdd.n640 185
R16515 vdd.n642 vdd.n641 185
R16516 vdd.n3252 vdd.n3251 185
R16517 vdd.n3253 vdd.n3252 185
R16518 vdd.n650 vdd.n649 185
R16519 vdd.n649 vdd.n648 185
R16520 vdd.n3247 vdd.n3246 185
R16521 vdd.n3246 vdd.n3245 185
R16522 vdd.n653 vdd.n652 185
R16523 vdd.n659 vdd.n653 185
R16524 vdd.n3236 vdd.n3235 185
R16525 vdd.n3237 vdd.n3236 185
R16526 vdd.n3232 vdd.n660 185
R16527 vdd.n3231 vdd.n3230 185
R16528 vdd.n3228 vdd.n662 185
R16529 vdd.n3228 vdd.n658 185
R16530 vdd.n3227 vdd.n3226 185
R16531 vdd.n3225 vdd.n3224 185
R16532 vdd.n3223 vdd.n3222 185
R16533 vdd.n3221 vdd.n3220 185
R16534 vdd.n3219 vdd.n668 185
R16535 vdd.n3217 vdd.n3216 185
R16536 vdd.n3215 vdd.n669 185
R16537 vdd.n3214 vdd.n3213 185
R16538 vdd.n3211 vdd.n674 185
R16539 vdd.n3209 vdd.n3208 185
R16540 vdd.n3207 vdd.n675 185
R16541 vdd.n3206 vdd.n3205 185
R16542 vdd.n3203 vdd.n680 185
R16543 vdd.n3201 vdd.n3200 185
R16544 vdd.n3199 vdd.n681 185
R16545 vdd.n3198 vdd.n3197 185
R16546 vdd.n3195 vdd.n688 185
R16547 vdd.n3193 vdd.n3192 185
R16548 vdd.n3191 vdd.n689 185
R16549 vdd.n3190 vdd.n3189 185
R16550 vdd.n3187 vdd.n694 185
R16551 vdd.n3185 vdd.n3184 185
R16552 vdd.n3183 vdd.n695 185
R16553 vdd.n3182 vdd.n3181 185
R16554 vdd.n3179 vdd.n700 185
R16555 vdd.n3177 vdd.n3176 185
R16556 vdd.n3175 vdd.n701 185
R16557 vdd.n3174 vdd.n3173 185
R16558 vdd.n3171 vdd.n706 185
R16559 vdd.n3169 vdd.n3168 185
R16560 vdd.n3167 vdd.n707 185
R16561 vdd.n3166 vdd.n3165 185
R16562 vdd.n3163 vdd.n712 185
R16563 vdd.n3161 vdd.n3160 185
R16564 vdd.n3159 vdd.n713 185
R16565 vdd.n3158 vdd.n3157 185
R16566 vdd.n3155 vdd.n718 185
R16567 vdd.n3153 vdd.n3152 185
R16568 vdd.n3151 vdd.n719 185
R16569 vdd.n728 vdd.n722 185
R16570 vdd.n3147 vdd.n3146 185
R16571 vdd.n3144 vdd.n726 185
R16572 vdd.n3143 vdd.n3142 185
R16573 vdd.n3141 vdd.n3140 185
R16574 vdd.n3139 vdd.n732 185
R16575 vdd.n3137 vdd.n3136 185
R16576 vdd.n3135 vdd.n733 185
R16577 vdd.n3134 vdd.n3133 185
R16578 vdd.n3131 vdd.n738 185
R16579 vdd.n3129 vdd.n3128 185
R16580 vdd.n3127 vdd.n739 185
R16581 vdd.n3126 vdd.n3125 185
R16582 vdd.n3123 vdd.n744 185
R16583 vdd.n3121 vdd.n3120 185
R16584 vdd.n3119 vdd.n745 185
R16585 vdd.n3118 vdd.n3117 185
R16586 vdd.n3115 vdd.n3114 185
R16587 vdd.n3113 vdd.n3112 185
R16588 vdd.n3111 vdd.n3110 185
R16589 vdd.n3109 vdd.n3108 185
R16590 vdd.n3104 vdd.n657 185
R16591 vdd.n658 vdd.n657 185
R16592 vdd.n3343 vdd.n3342 185
R16593 vdd.n599 vdd.n404 185
R16594 vdd.n598 vdd.n597 185
R16595 vdd.n596 vdd.n595 185
R16596 vdd.n594 vdd.n409 185
R16597 vdd.n590 vdd.n589 185
R16598 vdd.n588 vdd.n587 185
R16599 vdd.n586 vdd.n585 185
R16600 vdd.n584 vdd.n411 185
R16601 vdd.n580 vdd.n579 185
R16602 vdd.n578 vdd.n577 185
R16603 vdd.n576 vdd.n575 185
R16604 vdd.n574 vdd.n413 185
R16605 vdd.n570 vdd.n569 185
R16606 vdd.n568 vdd.n567 185
R16607 vdd.n566 vdd.n565 185
R16608 vdd.n564 vdd.n415 185
R16609 vdd.n560 vdd.n559 185
R16610 vdd.n558 vdd.n557 185
R16611 vdd.n556 vdd.n555 185
R16612 vdd.n554 vdd.n417 185
R16613 vdd.n550 vdd.n549 185
R16614 vdd.n548 vdd.n547 185
R16615 vdd.n546 vdd.n545 185
R16616 vdd.n544 vdd.n421 185
R16617 vdd.n540 vdd.n539 185
R16618 vdd.n538 vdd.n537 185
R16619 vdd.n536 vdd.n535 185
R16620 vdd.n534 vdd.n423 185
R16621 vdd.n530 vdd.n529 185
R16622 vdd.n528 vdd.n527 185
R16623 vdd.n526 vdd.n525 185
R16624 vdd.n524 vdd.n425 185
R16625 vdd.n520 vdd.n519 185
R16626 vdd.n518 vdd.n517 185
R16627 vdd.n516 vdd.n515 185
R16628 vdd.n514 vdd.n427 185
R16629 vdd.n510 vdd.n509 185
R16630 vdd.n508 vdd.n507 185
R16631 vdd.n506 vdd.n505 185
R16632 vdd.n504 vdd.n429 185
R16633 vdd.n500 vdd.n499 185
R16634 vdd.n498 vdd.n497 185
R16635 vdd.n496 vdd.n495 185
R16636 vdd.n494 vdd.n433 185
R16637 vdd.n490 vdd.n489 185
R16638 vdd.n488 vdd.n487 185
R16639 vdd.n486 vdd.n485 185
R16640 vdd.n484 vdd.n435 185
R16641 vdd.n480 vdd.n479 185
R16642 vdd.n478 vdd.n477 185
R16643 vdd.n476 vdd.n475 185
R16644 vdd.n474 vdd.n437 185
R16645 vdd.n470 vdd.n469 185
R16646 vdd.n468 vdd.n467 185
R16647 vdd.n466 vdd.n465 185
R16648 vdd.n464 vdd.n439 185
R16649 vdd.n460 vdd.n459 185
R16650 vdd.n458 vdd.n457 185
R16651 vdd.n456 vdd.n455 185
R16652 vdd.n454 vdd.n441 185
R16653 vdd.n450 vdd.n449 185
R16654 vdd.n448 vdd.n447 185
R16655 vdd.n446 vdd.n445 185
R16656 vdd.n3339 vdd.n372 185
R16657 vdd.n3346 vdd.n372 185
R16658 vdd.n3338 vdd.n371 185
R16659 vdd.n3347 vdd.n371 185
R16660 vdd.n3337 vdd.n3336 185
R16661 vdd.n3336 vdd.n363 185
R16662 vdd.n602 vdd.n362 185
R16663 vdd.n3353 vdd.n362 185
R16664 vdd.n3332 vdd.n361 185
R16665 vdd.n3354 vdd.n361 185
R16666 vdd.n3331 vdd.n360 185
R16667 vdd.n3355 vdd.n360 185
R16668 vdd.n3330 vdd.n3329 185
R16669 vdd.n3329 vdd.n3328 185
R16670 vdd.n604 vdd.n352 185
R16671 vdd.n3361 vdd.n352 185
R16672 vdd.n3324 vdd.n351 185
R16673 vdd.n3362 vdd.n351 185
R16674 vdd.n3323 vdd.n350 185
R16675 vdd.n3363 vdd.n350 185
R16676 vdd.n3322 vdd.n3321 185
R16677 vdd.n3321 vdd.n349 185
R16678 vdd.n606 vdd.n341 185
R16679 vdd.n3369 vdd.n341 185
R16680 vdd.n3317 vdd.n340 185
R16681 vdd.n3370 vdd.n340 185
R16682 vdd.n3316 vdd.n339 185
R16683 vdd.n3371 vdd.n339 185
R16684 vdd.n3315 vdd.n3314 185
R16685 vdd.n3314 vdd.n332 185
R16686 vdd.n608 vdd.n331 185
R16687 vdd.n3377 vdd.n331 185
R16688 vdd.n3310 vdd.n330 185
R16689 vdd.n3378 vdd.n330 185
R16690 vdd.n3309 vdd.n329 185
R16691 vdd.n3379 vdd.n329 185
R16692 vdd.n3308 vdd.n3307 185
R16693 vdd.n3307 vdd.n328 185
R16694 vdd.n3306 vdd.n610 185
R16695 vdd.n3306 vdd.n3305 185
R16696 vdd.n3294 vdd.n612 185
R16697 vdd.n613 vdd.n612 185
R16698 vdd.n3296 vdd.n3295 185
R16699 vdd.n3297 vdd.n3296 185
R16700 vdd.n620 vdd.n619 185
R16701 vdd.n624 vdd.n619 185
R16702 vdd.n3288 vdd.n3287 185
R16703 vdd.n3287 vdd.n3286 185
R16704 vdd.n623 vdd.n622 185
R16705 vdd.n3277 vdd.n623 185
R16706 vdd.n3276 vdd.n3275 185
R16707 vdd.n3278 vdd.n3276 185
R16708 vdd.n631 vdd.n630 185
R16709 vdd.n636 vdd.n630 185
R16710 vdd.n3271 vdd.n3270 185
R16711 vdd.n3270 vdd.n3269 185
R16712 vdd.n634 vdd.n633 185
R16713 vdd.n635 vdd.n634 185
R16714 vdd.n3260 vdd.n3259 185
R16715 vdd.n3261 vdd.n3260 185
R16716 vdd.n644 vdd.n643 185
R16717 vdd.n643 vdd.n642 185
R16718 vdd.n3255 vdd.n3254 185
R16719 vdd.n3254 vdd.n3253 185
R16720 vdd.n647 vdd.n646 185
R16721 vdd.n648 vdd.n647 185
R16722 vdd.n3244 vdd.n3243 185
R16723 vdd.n3245 vdd.n3244 185
R16724 vdd.n655 vdd.n654 185
R16725 vdd.n659 vdd.n654 185
R16726 vdd.n3239 vdd.n3238 185
R16727 vdd.n3238 vdd.n3237 185
R16728 vdd.n2853 vdd.n2852 185
R16729 vdd.n2851 vdd.n2617 185
R16730 vdd.n2850 vdd.n2616 185
R16731 vdd.n2855 vdd.n2616 185
R16732 vdd.n2849 vdd.n2848 185
R16733 vdd.n2847 vdd.n2846 185
R16734 vdd.n2845 vdd.n2844 185
R16735 vdd.n2843 vdd.n2842 185
R16736 vdd.n2841 vdd.n2840 185
R16737 vdd.n2839 vdd.n2838 185
R16738 vdd.n2837 vdd.n2836 185
R16739 vdd.n2835 vdd.n2834 185
R16740 vdd.n2833 vdd.n2832 185
R16741 vdd.n2831 vdd.n2830 185
R16742 vdd.n2829 vdd.n2828 185
R16743 vdd.n2827 vdd.n2826 185
R16744 vdd.n2825 vdd.n2824 185
R16745 vdd.n2823 vdd.n2822 185
R16746 vdd.n2821 vdd.n2820 185
R16747 vdd.n2819 vdd.n2818 185
R16748 vdd.n2817 vdd.n2816 185
R16749 vdd.n2815 vdd.n2814 185
R16750 vdd.n2813 vdd.n2812 185
R16751 vdd.n2811 vdd.n2810 185
R16752 vdd.n2809 vdd.n2808 185
R16753 vdd.n2807 vdd.n2806 185
R16754 vdd.n2805 vdd.n2804 185
R16755 vdd.n2803 vdd.n2802 185
R16756 vdd.n2801 vdd.n2800 185
R16757 vdd.n2799 vdd.n2798 185
R16758 vdd.n2797 vdd.n2796 185
R16759 vdd.n2795 vdd.n2794 185
R16760 vdd.n2793 vdd.n2792 185
R16761 vdd.n2790 vdd.n2789 185
R16762 vdd.n2788 vdd.n2787 185
R16763 vdd.n2786 vdd.n2785 185
R16764 vdd.n3005 vdd.n3004 185
R16765 vdd.n3006 vdd.n803 185
R16766 vdd.n3008 vdd.n3007 185
R16767 vdd.n3010 vdd.n801 185
R16768 vdd.n3012 vdd.n3011 185
R16769 vdd.n3013 vdd.n800 185
R16770 vdd.n3015 vdd.n3014 185
R16771 vdd.n3017 vdd.n798 185
R16772 vdd.n3019 vdd.n3018 185
R16773 vdd.n3020 vdd.n797 185
R16774 vdd.n3022 vdd.n3021 185
R16775 vdd.n3024 vdd.n795 185
R16776 vdd.n3026 vdd.n3025 185
R16777 vdd.n3027 vdd.n794 185
R16778 vdd.n3029 vdd.n3028 185
R16779 vdd.n3031 vdd.n792 185
R16780 vdd.n3033 vdd.n3032 185
R16781 vdd.n3035 vdd.n791 185
R16782 vdd.n3037 vdd.n3036 185
R16783 vdd.n3039 vdd.n789 185
R16784 vdd.n3041 vdd.n3040 185
R16785 vdd.n3042 vdd.n788 185
R16786 vdd.n3044 vdd.n3043 185
R16787 vdd.n3046 vdd.n786 185
R16788 vdd.n3048 vdd.n3047 185
R16789 vdd.n3049 vdd.n785 185
R16790 vdd.n3051 vdd.n3050 185
R16791 vdd.n3053 vdd.n783 185
R16792 vdd.n3055 vdd.n3054 185
R16793 vdd.n3056 vdd.n782 185
R16794 vdd.n3058 vdd.n3057 185
R16795 vdd.n3060 vdd.n781 185
R16796 vdd.n3061 vdd.n780 185
R16797 vdd.n3064 vdd.n3063 185
R16798 vdd.n3065 vdd.n778 185
R16799 vdd.n778 vdd.n756 185
R16800 vdd.n3002 vdd.n775 185
R16801 vdd.n3068 vdd.n775 185
R16802 vdd.n3001 vdd.n3000 185
R16803 vdd.n3000 vdd.n774 185
R16804 vdd.n2999 vdd.n807 185
R16805 vdd.n2999 vdd.n2998 185
R16806 vdd.n2733 vdd.n808 185
R16807 vdd.n817 vdd.n808 185
R16808 vdd.n2734 vdd.n815 185
R16809 vdd.n2992 vdd.n815 185
R16810 vdd.n2736 vdd.n2735 185
R16811 vdd.n2735 vdd.n814 185
R16812 vdd.n2737 vdd.n823 185
R16813 vdd.n2941 vdd.n823 185
R16814 vdd.n2739 vdd.n2738 185
R16815 vdd.n2738 vdd.n822 185
R16816 vdd.n2740 vdd.n829 185
R16817 vdd.n2935 vdd.n829 185
R16818 vdd.n2742 vdd.n2741 185
R16819 vdd.n2741 vdd.n828 185
R16820 vdd.n2743 vdd.n834 185
R16821 vdd.n2929 vdd.n834 185
R16822 vdd.n2745 vdd.n2744 185
R16823 vdd.n2744 vdd.n841 185
R16824 vdd.n2746 vdd.n839 185
R16825 vdd.n2923 vdd.n839 185
R16826 vdd.n2748 vdd.n2747 185
R16827 vdd.n2747 vdd.n849 185
R16828 vdd.n2749 vdd.n847 185
R16829 vdd.n2916 vdd.n847 185
R16830 vdd.n2751 vdd.n2750 185
R16831 vdd.n2750 vdd.n846 185
R16832 vdd.n2752 vdd.n854 185
R16833 vdd.n2910 vdd.n854 185
R16834 vdd.n2754 vdd.n2753 185
R16835 vdd.n2753 vdd.n853 185
R16836 vdd.n2755 vdd.n859 185
R16837 vdd.n2904 vdd.n859 185
R16838 vdd.n2757 vdd.n2756 185
R16839 vdd.n2756 vdd.n866 185
R16840 vdd.n2758 vdd.n864 185
R16841 vdd.n2898 vdd.n864 185
R16842 vdd.n2760 vdd.n2759 185
R16843 vdd.n2759 vdd.n872 185
R16844 vdd.n2761 vdd.n870 185
R16845 vdd.n2892 vdd.n870 185
R16846 vdd.n2763 vdd.n2762 185
R16847 vdd.n2764 vdd.n2763 185
R16848 vdd.n2732 vdd.n877 185
R16849 vdd.n2886 vdd.n877 185
R16850 vdd.n2731 vdd.n2730 185
R16851 vdd.n2730 vdd.n876 185
R16852 vdd.n2729 vdd.n883 185
R16853 vdd.n2880 vdd.n883 185
R16854 vdd.n2728 vdd.n2727 185
R16855 vdd.n2727 vdd.n882 185
R16856 vdd.n2726 vdd.n889 185
R16857 vdd.n2874 vdd.n889 185
R16858 vdd.n2725 vdd.n2724 185
R16859 vdd.n2724 vdd.n888 185
R16860 vdd.n2620 vdd.n894 185
R16861 vdd.n2868 vdd.n894 185
R16862 vdd.n2781 vdd.n2780 185
R16863 vdd.n2780 vdd.n2779 185
R16864 vdd.n2782 vdd.n900 185
R16865 vdd.n2862 vdd.n900 185
R16866 vdd.n2784 vdd.n2783 185
R16867 vdd.n2784 vdd.n899 185
R16868 vdd.n898 vdd.n897 185
R16869 vdd.n899 vdd.n898 185
R16870 vdd.n2864 vdd.n2863 185
R16871 vdd.n2863 vdd.n2862 185
R16872 vdd.n2865 vdd.n896 185
R16873 vdd.n2779 vdd.n896 185
R16874 vdd.n2867 vdd.n2866 185
R16875 vdd.n2868 vdd.n2867 185
R16876 vdd.n887 vdd.n886 185
R16877 vdd.n888 vdd.n887 185
R16878 vdd.n2876 vdd.n2875 185
R16879 vdd.n2875 vdd.n2874 185
R16880 vdd.n2877 vdd.n885 185
R16881 vdd.n885 vdd.n882 185
R16882 vdd.n2879 vdd.n2878 185
R16883 vdd.n2880 vdd.n2879 185
R16884 vdd.n875 vdd.n874 185
R16885 vdd.n876 vdd.n875 185
R16886 vdd.n2888 vdd.n2887 185
R16887 vdd.n2887 vdd.n2886 185
R16888 vdd.n2889 vdd.n873 185
R16889 vdd.n2764 vdd.n873 185
R16890 vdd.n2891 vdd.n2890 185
R16891 vdd.n2892 vdd.n2891 185
R16892 vdd.n863 vdd.n862 185
R16893 vdd.n872 vdd.n863 185
R16894 vdd.n2900 vdd.n2899 185
R16895 vdd.n2899 vdd.n2898 185
R16896 vdd.n2901 vdd.n861 185
R16897 vdd.n866 vdd.n861 185
R16898 vdd.n2903 vdd.n2902 185
R16899 vdd.n2904 vdd.n2903 185
R16900 vdd.n852 vdd.n851 185
R16901 vdd.n853 vdd.n852 185
R16902 vdd.n2912 vdd.n2911 185
R16903 vdd.n2911 vdd.n2910 185
R16904 vdd.n2913 vdd.n850 185
R16905 vdd.n850 vdd.n846 185
R16906 vdd.n2915 vdd.n2914 185
R16907 vdd.n2916 vdd.n2915 185
R16908 vdd.n838 vdd.n837 185
R16909 vdd.n849 vdd.n838 185
R16910 vdd.n2925 vdd.n2924 185
R16911 vdd.n2924 vdd.n2923 185
R16912 vdd.n2926 vdd.n836 185
R16913 vdd.n841 vdd.n836 185
R16914 vdd.n2928 vdd.n2927 185
R16915 vdd.n2929 vdd.n2928 185
R16916 vdd.n827 vdd.n826 185
R16917 vdd.n828 vdd.n827 185
R16918 vdd.n2937 vdd.n2936 185
R16919 vdd.n2936 vdd.n2935 185
R16920 vdd.n2938 vdd.n825 185
R16921 vdd.n825 vdd.n822 185
R16922 vdd.n2940 vdd.n2939 185
R16923 vdd.n2941 vdd.n2940 185
R16924 vdd.n813 vdd.n812 185
R16925 vdd.n814 vdd.n813 185
R16926 vdd.n2994 vdd.n2993 185
R16927 vdd.n2993 vdd.n2992 185
R16928 vdd.n2995 vdd.n811 185
R16929 vdd.n817 vdd.n811 185
R16930 vdd.n2997 vdd.n2996 185
R16931 vdd.n2998 vdd.n2997 185
R16932 vdd.n779 vdd.n777 185
R16933 vdd.n777 vdd.n774 185
R16934 vdd.n3067 vdd.n3066 185
R16935 vdd.n3068 vdd.n3067 185
R16936 vdd.n2509 vdd.n2508 185
R16937 vdd.n2510 vdd.n2509 185
R16938 vdd.n951 vdd.n949 185
R16939 vdd.n949 vdd.n947 185
R16940 vdd.n2424 vdd.n958 185
R16941 vdd.n2435 vdd.n958 185
R16942 vdd.n2425 vdd.n967 185
R16943 vdd.n1309 vdd.n967 185
R16944 vdd.n2427 vdd.n2426 185
R16945 vdd.n2428 vdd.n2427 185
R16946 vdd.n2423 vdd.n966 185
R16947 vdd.n966 vdd.n963 185
R16948 vdd.n2422 vdd.n2421 185
R16949 vdd.n2421 vdd.n2420 185
R16950 vdd.n969 vdd.n968 185
R16951 vdd.n970 vdd.n969 185
R16952 vdd.n2413 vdd.n2412 185
R16953 vdd.n2414 vdd.n2413 185
R16954 vdd.n2411 vdd.n979 185
R16955 vdd.n979 vdd.n976 185
R16956 vdd.n2410 vdd.n2409 185
R16957 vdd.n2409 vdd.n2408 185
R16958 vdd.n981 vdd.n980 185
R16959 vdd.n989 vdd.n981 185
R16960 vdd.n2401 vdd.n2400 185
R16961 vdd.n2402 vdd.n2401 185
R16962 vdd.n2399 vdd.n990 185
R16963 vdd.n995 vdd.n990 185
R16964 vdd.n2398 vdd.n2397 185
R16965 vdd.n2397 vdd.n2396 185
R16966 vdd.n992 vdd.n991 185
R16967 vdd.n1330 vdd.n992 185
R16968 vdd.n2389 vdd.n2388 185
R16969 vdd.n2390 vdd.n2389 185
R16970 vdd.n2387 vdd.n1002 185
R16971 vdd.n1002 vdd.n999 185
R16972 vdd.n2386 vdd.n2385 185
R16973 vdd.n2385 vdd.n2384 185
R16974 vdd.n1004 vdd.n1003 185
R16975 vdd.n1005 vdd.n1004 185
R16976 vdd.n2377 vdd.n2376 185
R16977 vdd.n2378 vdd.n2377 185
R16978 vdd.n2374 vdd.n1013 185
R16979 vdd.n1019 vdd.n1013 185
R16980 vdd.n2373 vdd.n2372 185
R16981 vdd.n2372 vdd.n2371 185
R16982 vdd.n1016 vdd.n1015 185
R16983 vdd.n1026 vdd.n1016 185
R16984 vdd.n2364 vdd.n2363 185
R16985 vdd.n2365 vdd.n2364 185
R16986 vdd.n2362 vdd.n1027 185
R16987 vdd.n1027 vdd.n1023 185
R16988 vdd.n2361 vdd.n2360 185
R16989 vdd.n2360 vdd.n2359 185
R16990 vdd.n1029 vdd.n1028 185
R16991 vdd.n1030 vdd.n1029 185
R16992 vdd.n2352 vdd.n2351 185
R16993 vdd.n2353 vdd.n2352 185
R16994 vdd.n2350 vdd.n1039 185
R16995 vdd.n1039 vdd.n1036 185
R16996 vdd.n2349 vdd.n2348 185
R16997 vdd.n2348 vdd.n2347 185
R16998 vdd.n1041 vdd.n1040 185
R16999 vdd.n1050 vdd.n1041 185
R17000 vdd.n2340 vdd.n2339 185
R17001 vdd.n2341 vdd.n2340 185
R17002 vdd.n2338 vdd.n1051 185
R17003 vdd.n1051 vdd.n1047 185
R17004 vdd.n2440 vdd.n922 185
R17005 vdd.n2582 vdd.n922 185
R17006 vdd.n2442 vdd.n2441 185
R17007 vdd.n2444 vdd.n2443 185
R17008 vdd.n2446 vdd.n2445 185
R17009 vdd.n2448 vdd.n2447 185
R17010 vdd.n2450 vdd.n2449 185
R17011 vdd.n2452 vdd.n2451 185
R17012 vdd.n2454 vdd.n2453 185
R17013 vdd.n2456 vdd.n2455 185
R17014 vdd.n2458 vdd.n2457 185
R17015 vdd.n2460 vdd.n2459 185
R17016 vdd.n2462 vdd.n2461 185
R17017 vdd.n2464 vdd.n2463 185
R17018 vdd.n2466 vdd.n2465 185
R17019 vdd.n2468 vdd.n2467 185
R17020 vdd.n2470 vdd.n2469 185
R17021 vdd.n2472 vdd.n2471 185
R17022 vdd.n2474 vdd.n2473 185
R17023 vdd.n2476 vdd.n2475 185
R17024 vdd.n2478 vdd.n2477 185
R17025 vdd.n2480 vdd.n2479 185
R17026 vdd.n2482 vdd.n2481 185
R17027 vdd.n2484 vdd.n2483 185
R17028 vdd.n2486 vdd.n2485 185
R17029 vdd.n2488 vdd.n2487 185
R17030 vdd.n2490 vdd.n2489 185
R17031 vdd.n2492 vdd.n2491 185
R17032 vdd.n2494 vdd.n2493 185
R17033 vdd.n2496 vdd.n2495 185
R17034 vdd.n2498 vdd.n2497 185
R17035 vdd.n2500 vdd.n2499 185
R17036 vdd.n2502 vdd.n2501 185
R17037 vdd.n2504 vdd.n2503 185
R17038 vdd.n2506 vdd.n2505 185
R17039 vdd.n2507 vdd.n950 185
R17040 vdd.n2439 vdd.n948 185
R17041 vdd.n2510 vdd.n948 185
R17042 vdd.n2438 vdd.n2437 185
R17043 vdd.n2437 vdd.n947 185
R17044 vdd.n2436 vdd.n955 185
R17045 vdd.n2436 vdd.n2435 185
R17046 vdd.n1227 vdd.n956 185
R17047 vdd.n1309 vdd.n956 185
R17048 vdd.n1228 vdd.n965 185
R17049 vdd.n2428 vdd.n965 185
R17050 vdd.n1230 vdd.n1229 185
R17051 vdd.n1229 vdd.n963 185
R17052 vdd.n1231 vdd.n972 185
R17053 vdd.n2420 vdd.n972 185
R17054 vdd.n1233 vdd.n1232 185
R17055 vdd.n1232 vdd.n970 185
R17056 vdd.n1234 vdd.n978 185
R17057 vdd.n2414 vdd.n978 185
R17058 vdd.n1236 vdd.n1235 185
R17059 vdd.n1235 vdd.n976 185
R17060 vdd.n1237 vdd.n983 185
R17061 vdd.n2408 vdd.n983 185
R17062 vdd.n1239 vdd.n1238 185
R17063 vdd.n1238 vdd.n989 185
R17064 vdd.n1240 vdd.n988 185
R17065 vdd.n2402 vdd.n988 185
R17066 vdd.n1242 vdd.n1241 185
R17067 vdd.n1241 vdd.n995 185
R17068 vdd.n1243 vdd.n994 185
R17069 vdd.n2396 vdd.n994 185
R17070 vdd.n1332 vdd.n1331 185
R17071 vdd.n1331 vdd.n1330 185
R17072 vdd.n1333 vdd.n1001 185
R17073 vdd.n2390 vdd.n1001 185
R17074 vdd.n1335 vdd.n1334 185
R17075 vdd.n1334 vdd.n999 185
R17076 vdd.n1336 vdd.n1007 185
R17077 vdd.n2384 vdd.n1007 185
R17078 vdd.n1338 vdd.n1337 185
R17079 vdd.n1337 vdd.n1005 185
R17080 vdd.n1339 vdd.n1012 185
R17081 vdd.n2378 vdd.n1012 185
R17082 vdd.n1341 vdd.n1340 185
R17083 vdd.n1340 vdd.n1019 185
R17084 vdd.n1342 vdd.n1018 185
R17085 vdd.n2371 vdd.n1018 185
R17086 vdd.n1344 vdd.n1343 185
R17087 vdd.n1343 vdd.n1026 185
R17088 vdd.n1345 vdd.n1025 185
R17089 vdd.n2365 vdd.n1025 185
R17090 vdd.n1347 vdd.n1346 185
R17091 vdd.n1346 vdd.n1023 185
R17092 vdd.n1348 vdd.n1032 185
R17093 vdd.n2359 vdd.n1032 185
R17094 vdd.n1350 vdd.n1349 185
R17095 vdd.n1349 vdd.n1030 185
R17096 vdd.n1351 vdd.n1038 185
R17097 vdd.n2353 vdd.n1038 185
R17098 vdd.n1353 vdd.n1352 185
R17099 vdd.n1352 vdd.n1036 185
R17100 vdd.n1354 vdd.n1043 185
R17101 vdd.n2347 vdd.n1043 185
R17102 vdd.n1356 vdd.n1355 185
R17103 vdd.n1355 vdd.n1050 185
R17104 vdd.n1357 vdd.n1049 185
R17105 vdd.n2341 vdd.n1049 185
R17106 vdd.n1359 vdd.n1358 185
R17107 vdd.n1358 vdd.n1047 185
R17108 vdd.n2337 vdd.n2336 185
R17109 vdd.n1053 vdd.n1052 185
R17110 vdd.n1194 vdd.n1193 185
R17111 vdd.n1196 vdd.n1195 185
R17112 vdd.n1198 vdd.n1197 185
R17113 vdd.n1200 vdd.n1199 185
R17114 vdd.n1202 vdd.n1201 185
R17115 vdd.n1204 vdd.n1203 185
R17116 vdd.n1206 vdd.n1205 185
R17117 vdd.n1208 vdd.n1207 185
R17118 vdd.n1210 vdd.n1209 185
R17119 vdd.n1212 vdd.n1211 185
R17120 vdd.n1214 vdd.n1213 185
R17121 vdd.n1216 vdd.n1215 185
R17122 vdd.n1218 vdd.n1217 185
R17123 vdd.n1220 vdd.n1219 185
R17124 vdd.n1222 vdd.n1221 185
R17125 vdd.n1393 vdd.n1223 185
R17126 vdd.n1392 vdd.n1391 185
R17127 vdd.n1390 vdd.n1389 185
R17128 vdd.n1388 vdd.n1387 185
R17129 vdd.n1386 vdd.n1385 185
R17130 vdd.n1384 vdd.n1383 185
R17131 vdd.n1382 vdd.n1381 185
R17132 vdd.n1380 vdd.n1379 185
R17133 vdd.n1378 vdd.n1377 185
R17134 vdd.n1376 vdd.n1375 185
R17135 vdd.n1374 vdd.n1373 185
R17136 vdd.n1372 vdd.n1371 185
R17137 vdd.n1370 vdd.n1369 185
R17138 vdd.n1368 vdd.n1367 185
R17139 vdd.n1366 vdd.n1365 185
R17140 vdd.n1364 vdd.n1363 185
R17141 vdd.n1362 vdd.n1361 185
R17142 vdd.n1360 vdd.n1087 185
R17143 vdd.n2334 vdd.n1087 185
R17144 vdd.n2334 vdd.n1054 179.345
R17145 vdd.n756 vdd.n658 179.345
R17146 vdd.n315 vdd.n314 171.744
R17147 vdd.n314 vdd.n313 171.744
R17148 vdd.n313 vdd.n282 171.744
R17149 vdd.n306 vdd.n282 171.744
R17150 vdd.n306 vdd.n305 171.744
R17151 vdd.n305 vdd.n287 171.744
R17152 vdd.n298 vdd.n287 171.744
R17153 vdd.n298 vdd.n297 171.744
R17154 vdd.n297 vdd.n291 171.744
R17155 vdd.n260 vdd.n259 171.744
R17156 vdd.n259 vdd.n258 171.744
R17157 vdd.n258 vdd.n227 171.744
R17158 vdd.n251 vdd.n227 171.744
R17159 vdd.n251 vdd.n250 171.744
R17160 vdd.n250 vdd.n232 171.744
R17161 vdd.n243 vdd.n232 171.744
R17162 vdd.n243 vdd.n242 171.744
R17163 vdd.n242 vdd.n236 171.744
R17164 vdd.n217 vdd.n216 171.744
R17165 vdd.n216 vdd.n215 171.744
R17166 vdd.n215 vdd.n184 171.744
R17167 vdd.n208 vdd.n184 171.744
R17168 vdd.n208 vdd.n207 171.744
R17169 vdd.n207 vdd.n189 171.744
R17170 vdd.n200 vdd.n189 171.744
R17171 vdd.n200 vdd.n199 171.744
R17172 vdd.n199 vdd.n193 171.744
R17173 vdd.n162 vdd.n161 171.744
R17174 vdd.n161 vdd.n160 171.744
R17175 vdd.n160 vdd.n129 171.744
R17176 vdd.n153 vdd.n129 171.744
R17177 vdd.n153 vdd.n152 171.744
R17178 vdd.n152 vdd.n134 171.744
R17179 vdd.n145 vdd.n134 171.744
R17180 vdd.n145 vdd.n144 171.744
R17181 vdd.n144 vdd.n138 171.744
R17182 vdd.n120 vdd.n119 171.744
R17183 vdd.n119 vdd.n118 171.744
R17184 vdd.n118 vdd.n87 171.744
R17185 vdd.n111 vdd.n87 171.744
R17186 vdd.n111 vdd.n110 171.744
R17187 vdd.n110 vdd.n92 171.744
R17188 vdd.n103 vdd.n92 171.744
R17189 vdd.n103 vdd.n102 171.744
R17190 vdd.n102 vdd.n96 171.744
R17191 vdd.n65 vdd.n64 171.744
R17192 vdd.n64 vdd.n63 171.744
R17193 vdd.n63 vdd.n32 171.744
R17194 vdd.n56 vdd.n32 171.744
R17195 vdd.n56 vdd.n55 171.744
R17196 vdd.n55 vdd.n37 171.744
R17197 vdd.n48 vdd.n37 171.744
R17198 vdd.n48 vdd.n47 171.744
R17199 vdd.n47 vdd.n41 171.744
R17200 vdd.n2046 vdd.n2045 171.744
R17201 vdd.n2045 vdd.n2044 171.744
R17202 vdd.n2044 vdd.n2013 171.744
R17203 vdd.n2037 vdd.n2013 171.744
R17204 vdd.n2037 vdd.n2036 171.744
R17205 vdd.n2036 vdd.n2018 171.744
R17206 vdd.n2029 vdd.n2018 171.744
R17207 vdd.n2029 vdd.n2028 171.744
R17208 vdd.n2028 vdd.n2022 171.744
R17209 vdd.n2101 vdd.n2100 171.744
R17210 vdd.n2100 vdd.n2099 171.744
R17211 vdd.n2099 vdd.n2068 171.744
R17212 vdd.n2092 vdd.n2068 171.744
R17213 vdd.n2092 vdd.n2091 171.744
R17214 vdd.n2091 vdd.n2073 171.744
R17215 vdd.n2084 vdd.n2073 171.744
R17216 vdd.n2084 vdd.n2083 171.744
R17217 vdd.n2083 vdd.n2077 171.744
R17218 vdd.n1948 vdd.n1947 171.744
R17219 vdd.n1947 vdd.n1946 171.744
R17220 vdd.n1946 vdd.n1915 171.744
R17221 vdd.n1939 vdd.n1915 171.744
R17222 vdd.n1939 vdd.n1938 171.744
R17223 vdd.n1938 vdd.n1920 171.744
R17224 vdd.n1931 vdd.n1920 171.744
R17225 vdd.n1931 vdd.n1930 171.744
R17226 vdd.n1930 vdd.n1924 171.744
R17227 vdd.n2003 vdd.n2002 171.744
R17228 vdd.n2002 vdd.n2001 171.744
R17229 vdd.n2001 vdd.n1970 171.744
R17230 vdd.n1994 vdd.n1970 171.744
R17231 vdd.n1994 vdd.n1993 171.744
R17232 vdd.n1993 vdd.n1975 171.744
R17233 vdd.n1986 vdd.n1975 171.744
R17234 vdd.n1986 vdd.n1985 171.744
R17235 vdd.n1985 vdd.n1979 171.744
R17236 vdd.n1851 vdd.n1850 171.744
R17237 vdd.n1850 vdd.n1849 171.744
R17238 vdd.n1849 vdd.n1818 171.744
R17239 vdd.n1842 vdd.n1818 171.744
R17240 vdd.n1842 vdd.n1841 171.744
R17241 vdd.n1841 vdd.n1823 171.744
R17242 vdd.n1834 vdd.n1823 171.744
R17243 vdd.n1834 vdd.n1833 171.744
R17244 vdd.n1833 vdd.n1827 171.744
R17245 vdd.n1906 vdd.n1905 171.744
R17246 vdd.n1905 vdd.n1904 171.744
R17247 vdd.n1904 vdd.n1873 171.744
R17248 vdd.n1897 vdd.n1873 171.744
R17249 vdd.n1897 vdd.n1896 171.744
R17250 vdd.n1896 vdd.n1878 171.744
R17251 vdd.n1889 vdd.n1878 171.744
R17252 vdd.n1889 vdd.n1888 171.744
R17253 vdd.n1888 vdd.n1882 171.744
R17254 vdd.n449 vdd.n448 146.341
R17255 vdd.n455 vdd.n454 146.341
R17256 vdd.n459 vdd.n458 146.341
R17257 vdd.n465 vdd.n464 146.341
R17258 vdd.n469 vdd.n468 146.341
R17259 vdd.n475 vdd.n474 146.341
R17260 vdd.n479 vdd.n478 146.341
R17261 vdd.n485 vdd.n484 146.341
R17262 vdd.n489 vdd.n488 146.341
R17263 vdd.n495 vdd.n494 146.341
R17264 vdd.n499 vdd.n498 146.341
R17265 vdd.n505 vdd.n504 146.341
R17266 vdd.n509 vdd.n508 146.341
R17267 vdd.n515 vdd.n514 146.341
R17268 vdd.n519 vdd.n518 146.341
R17269 vdd.n525 vdd.n524 146.341
R17270 vdd.n529 vdd.n528 146.341
R17271 vdd.n535 vdd.n534 146.341
R17272 vdd.n539 vdd.n538 146.341
R17273 vdd.n545 vdd.n544 146.341
R17274 vdd.n549 vdd.n548 146.341
R17275 vdd.n555 vdd.n554 146.341
R17276 vdd.n559 vdd.n558 146.341
R17277 vdd.n565 vdd.n564 146.341
R17278 vdd.n569 vdd.n568 146.341
R17279 vdd.n575 vdd.n574 146.341
R17280 vdd.n579 vdd.n578 146.341
R17281 vdd.n585 vdd.n584 146.341
R17282 vdd.n589 vdd.n588 146.341
R17283 vdd.n595 vdd.n594 146.341
R17284 vdd.n597 vdd.n404 146.341
R17285 vdd.n3238 vdd.n654 146.341
R17286 vdd.n3244 vdd.n654 146.341
R17287 vdd.n3244 vdd.n647 146.341
R17288 vdd.n3254 vdd.n647 146.341
R17289 vdd.n3254 vdd.n643 146.341
R17290 vdd.n3260 vdd.n643 146.341
R17291 vdd.n3260 vdd.n634 146.341
R17292 vdd.n3270 vdd.n634 146.341
R17293 vdd.n3270 vdd.n630 146.341
R17294 vdd.n3276 vdd.n630 146.341
R17295 vdd.n3276 vdd.n623 146.341
R17296 vdd.n3287 vdd.n623 146.341
R17297 vdd.n3287 vdd.n619 146.341
R17298 vdd.n3296 vdd.n619 146.341
R17299 vdd.n3296 vdd.n612 146.341
R17300 vdd.n3306 vdd.n612 146.341
R17301 vdd.n3307 vdd.n3306 146.341
R17302 vdd.n3307 vdd.n329 146.341
R17303 vdd.n330 vdd.n329 146.341
R17304 vdd.n331 vdd.n330 146.341
R17305 vdd.n3314 vdd.n331 146.341
R17306 vdd.n3314 vdd.n339 146.341
R17307 vdd.n340 vdd.n339 146.341
R17308 vdd.n341 vdd.n340 146.341
R17309 vdd.n3321 vdd.n341 146.341
R17310 vdd.n3321 vdd.n350 146.341
R17311 vdd.n351 vdd.n350 146.341
R17312 vdd.n352 vdd.n351 146.341
R17313 vdd.n3329 vdd.n352 146.341
R17314 vdd.n3329 vdd.n360 146.341
R17315 vdd.n361 vdd.n360 146.341
R17316 vdd.n362 vdd.n361 146.341
R17317 vdd.n3336 vdd.n362 146.341
R17318 vdd.n3336 vdd.n371 146.341
R17319 vdd.n372 vdd.n371 146.341
R17320 vdd.n3230 vdd.n3228 146.341
R17321 vdd.n3228 vdd.n3227 146.341
R17322 vdd.n3224 vdd.n3223 146.341
R17323 vdd.n3220 vdd.n3219 146.341
R17324 vdd.n3217 vdd.n669 146.341
R17325 vdd.n3213 vdd.n3211 146.341
R17326 vdd.n3209 vdd.n675 146.341
R17327 vdd.n3205 vdd.n3203 146.341
R17328 vdd.n3201 vdd.n681 146.341
R17329 vdd.n3197 vdd.n3195 146.341
R17330 vdd.n3193 vdd.n689 146.341
R17331 vdd.n3189 vdd.n3187 146.341
R17332 vdd.n3185 vdd.n695 146.341
R17333 vdd.n3181 vdd.n3179 146.341
R17334 vdd.n3177 vdd.n701 146.341
R17335 vdd.n3173 vdd.n3171 146.341
R17336 vdd.n3169 vdd.n707 146.341
R17337 vdd.n3165 vdd.n3163 146.341
R17338 vdd.n3161 vdd.n713 146.341
R17339 vdd.n3157 vdd.n3155 146.341
R17340 vdd.n3153 vdd.n719 146.341
R17341 vdd.n3146 vdd.n728 146.341
R17342 vdd.n3144 vdd.n3143 146.341
R17343 vdd.n3140 vdd.n3139 146.341
R17344 vdd.n3137 vdd.n733 146.341
R17345 vdd.n3133 vdd.n3131 146.341
R17346 vdd.n3129 vdd.n739 146.341
R17347 vdd.n3125 vdd.n3123 146.341
R17348 vdd.n3121 vdd.n745 146.341
R17349 vdd.n3117 vdd.n3115 146.341
R17350 vdd.n3112 vdd.n3111 146.341
R17351 vdd.n3108 vdd.n657 146.341
R17352 vdd.n3236 vdd.n653 146.341
R17353 vdd.n3246 vdd.n653 146.341
R17354 vdd.n3246 vdd.n649 146.341
R17355 vdd.n3252 vdd.n649 146.341
R17356 vdd.n3252 vdd.n641 146.341
R17357 vdd.n3262 vdd.n641 146.341
R17358 vdd.n3262 vdd.n637 146.341
R17359 vdd.n3268 vdd.n637 146.341
R17360 vdd.n3268 vdd.n629 146.341
R17361 vdd.n3279 vdd.n629 146.341
R17362 vdd.n3279 vdd.n625 146.341
R17363 vdd.n3285 vdd.n625 146.341
R17364 vdd.n3285 vdd.n618 146.341
R17365 vdd.n3298 vdd.n618 146.341
R17366 vdd.n3298 vdd.n614 146.341
R17367 vdd.n3304 vdd.n614 146.341
R17368 vdd.n3304 vdd.n326 146.341
R17369 vdd.n3380 vdd.n326 146.341
R17370 vdd.n3380 vdd.n327 146.341
R17371 vdd.n3376 vdd.n327 146.341
R17372 vdd.n3376 vdd.n333 146.341
R17373 vdd.n3372 vdd.n333 146.341
R17374 vdd.n3372 vdd.n338 146.341
R17375 vdd.n3368 vdd.n338 146.341
R17376 vdd.n3368 vdd.n342 146.341
R17377 vdd.n3364 vdd.n342 146.341
R17378 vdd.n3364 vdd.n348 146.341
R17379 vdd.n3360 vdd.n348 146.341
R17380 vdd.n3360 vdd.n353 146.341
R17381 vdd.n3356 vdd.n353 146.341
R17382 vdd.n3356 vdd.n359 146.341
R17383 vdd.n3352 vdd.n359 146.341
R17384 vdd.n3352 vdd.n364 146.341
R17385 vdd.n3348 vdd.n364 146.341
R17386 vdd.n3348 vdd.n370 146.341
R17387 vdd.n2295 vdd.n2294 146.341
R17388 vdd.n2292 vdd.n2289 146.341
R17389 vdd.n2287 vdd.n1098 146.341
R17390 vdd.n2283 vdd.n2282 146.341
R17391 vdd.n2280 vdd.n1102 146.341
R17392 vdd.n2276 vdd.n2275 146.341
R17393 vdd.n2273 vdd.n1109 146.341
R17394 vdd.n2269 vdd.n2268 146.341
R17395 vdd.n2266 vdd.n1116 146.341
R17396 vdd.n1127 vdd.n1124 146.341
R17397 vdd.n2258 vdd.n2257 146.341
R17398 vdd.n2255 vdd.n1129 146.341
R17399 vdd.n2251 vdd.n2250 146.341
R17400 vdd.n2248 vdd.n1135 146.341
R17401 vdd.n2244 vdd.n2243 146.341
R17402 vdd.n2241 vdd.n1142 146.341
R17403 vdd.n2237 vdd.n2236 146.341
R17404 vdd.n2234 vdd.n1149 146.341
R17405 vdd.n2230 vdd.n2229 146.341
R17406 vdd.n2227 vdd.n1156 146.341
R17407 vdd.n1167 vdd.n1164 146.341
R17408 vdd.n2219 vdd.n2218 146.341
R17409 vdd.n2216 vdd.n1169 146.341
R17410 vdd.n2212 vdd.n2211 146.341
R17411 vdd.n2209 vdd.n1175 146.341
R17412 vdd.n2205 vdd.n2204 146.341
R17413 vdd.n2202 vdd.n1182 146.341
R17414 vdd.n2198 vdd.n2197 146.341
R17415 vdd.n2195 vdd.n1189 146.341
R17416 vdd.n1400 vdd.n1398 146.341
R17417 vdd.n1403 vdd.n1402 146.341
R17418 vdd.n1743 vdd.n1507 146.341
R17419 vdd.n1743 vdd.n1499 146.341
R17420 vdd.n1753 vdd.n1499 146.341
R17421 vdd.n1753 vdd.n1495 146.341
R17422 vdd.n1759 vdd.n1495 146.341
R17423 vdd.n1759 vdd.n1487 146.341
R17424 vdd.n1770 vdd.n1487 146.341
R17425 vdd.n1770 vdd.n1483 146.341
R17426 vdd.n1776 vdd.n1483 146.341
R17427 vdd.n1776 vdd.n1477 146.341
R17428 vdd.n1787 vdd.n1477 146.341
R17429 vdd.n1787 vdd.n1473 146.341
R17430 vdd.n1793 vdd.n1473 146.341
R17431 vdd.n1793 vdd.n1464 146.341
R17432 vdd.n1803 vdd.n1464 146.341
R17433 vdd.n1803 vdd.n1460 146.341
R17434 vdd.n1809 vdd.n1460 146.341
R17435 vdd.n1809 vdd.n1453 146.341
R17436 vdd.n2115 vdd.n1453 146.341
R17437 vdd.n2115 vdd.n1449 146.341
R17438 vdd.n2121 vdd.n1449 146.341
R17439 vdd.n2121 vdd.n1442 146.341
R17440 vdd.n2131 vdd.n1442 146.341
R17441 vdd.n2131 vdd.n1438 146.341
R17442 vdd.n2137 vdd.n1438 146.341
R17443 vdd.n2137 vdd.n1430 146.341
R17444 vdd.n2148 vdd.n1430 146.341
R17445 vdd.n2148 vdd.n1426 146.341
R17446 vdd.n2154 vdd.n1426 146.341
R17447 vdd.n2154 vdd.n1420 146.341
R17448 vdd.n2165 vdd.n1420 146.341
R17449 vdd.n2165 vdd.n1415 146.341
R17450 vdd.n2173 vdd.n1415 146.341
R17451 vdd.n2173 vdd.n1405 146.341
R17452 vdd.n2183 vdd.n1405 146.341
R17453 vdd.n1545 vdd.n1544 146.341
R17454 vdd.n1549 vdd.n1544 146.341
R17455 vdd.n1551 vdd.n1550 146.341
R17456 vdd.n1555 vdd.n1554 146.341
R17457 vdd.n1557 vdd.n1556 146.341
R17458 vdd.n1561 vdd.n1560 146.341
R17459 vdd.n1563 vdd.n1562 146.341
R17460 vdd.n1567 vdd.n1566 146.341
R17461 vdd.n1569 vdd.n1568 146.341
R17462 vdd.n1701 vdd.n1700 146.341
R17463 vdd.n1573 vdd.n1572 146.341
R17464 vdd.n1577 vdd.n1576 146.341
R17465 vdd.n1579 vdd.n1578 146.341
R17466 vdd.n1583 vdd.n1582 146.341
R17467 vdd.n1585 vdd.n1584 146.341
R17468 vdd.n1589 vdd.n1588 146.341
R17469 vdd.n1591 vdd.n1590 146.341
R17470 vdd.n1595 vdd.n1594 146.341
R17471 vdd.n1597 vdd.n1596 146.341
R17472 vdd.n1601 vdd.n1600 146.341
R17473 vdd.n1665 vdd.n1602 146.341
R17474 vdd.n1606 vdd.n1605 146.341
R17475 vdd.n1608 vdd.n1607 146.341
R17476 vdd.n1612 vdd.n1611 146.341
R17477 vdd.n1614 vdd.n1613 146.341
R17478 vdd.n1618 vdd.n1617 146.341
R17479 vdd.n1620 vdd.n1619 146.341
R17480 vdd.n1624 vdd.n1623 146.341
R17481 vdd.n1626 vdd.n1625 146.341
R17482 vdd.n1630 vdd.n1629 146.341
R17483 vdd.n1632 vdd.n1631 146.341
R17484 vdd.n1737 vdd.n1513 146.341
R17485 vdd.n1745 vdd.n1505 146.341
R17486 vdd.n1745 vdd.n1501 146.341
R17487 vdd.n1751 vdd.n1501 146.341
R17488 vdd.n1751 vdd.n1493 146.341
R17489 vdd.n1762 vdd.n1493 146.341
R17490 vdd.n1762 vdd.n1489 146.341
R17491 vdd.n1768 vdd.n1489 146.341
R17492 vdd.n1768 vdd.n1482 146.341
R17493 vdd.n1779 vdd.n1482 146.341
R17494 vdd.n1779 vdd.n1478 146.341
R17495 vdd.n1785 vdd.n1478 146.341
R17496 vdd.n1785 vdd.n1471 146.341
R17497 vdd.n1795 vdd.n1471 146.341
R17498 vdd.n1795 vdd.n1467 146.341
R17499 vdd.n1801 vdd.n1467 146.341
R17500 vdd.n1801 vdd.n1459 146.341
R17501 vdd.n1812 vdd.n1459 146.341
R17502 vdd.n1812 vdd.n1455 146.341
R17503 vdd.n2113 vdd.n1455 146.341
R17504 vdd.n2113 vdd.n1448 146.341
R17505 vdd.n2123 vdd.n1448 146.341
R17506 vdd.n2123 vdd.n1444 146.341
R17507 vdd.n2129 vdd.n1444 146.341
R17508 vdd.n2129 vdd.n1436 146.341
R17509 vdd.n2140 vdd.n1436 146.341
R17510 vdd.n2140 vdd.n1432 146.341
R17511 vdd.n2146 vdd.n1432 146.341
R17512 vdd.n2146 vdd.n1425 146.341
R17513 vdd.n2157 vdd.n1425 146.341
R17514 vdd.n2157 vdd.n1421 146.341
R17515 vdd.n2163 vdd.n1421 146.341
R17516 vdd.n2163 vdd.n1413 146.341
R17517 vdd.n2175 vdd.n1413 146.341
R17518 vdd.n2175 vdd.n1408 146.341
R17519 vdd.n2181 vdd.n1408 146.341
R17520 vdd.n1224 vdd.t56 127.284
R17521 vdd.n952 vdd.t97 127.284
R17522 vdd.n1244 vdd.t70 127.284
R17523 vdd.n943 vdd.t114 127.284
R17524 vdd.n843 vdd.t73 127.284
R17525 vdd.n843 vdd.t74 127.284
R17526 vdd.n2621 vdd.t112 127.284
R17527 vdd.n804 vdd.t120 127.284
R17528 vdd.n2618 vdd.t102 127.284
R17529 vdd.n768 vdd.t51 127.284
R17530 vdd.n1014 vdd.t105 127.284
R17531 vdd.n1014 vdd.t106 127.284
R17532 vdd.n22 vdd.n20 117.314
R17533 vdd.n17 vdd.n15 117.314
R17534 vdd.n27 vdd.n26 116.927
R17535 vdd.n24 vdd.n23 116.927
R17536 vdd.n22 vdd.n21 116.927
R17537 vdd.n17 vdd.n16 116.927
R17538 vdd.n19 vdd.n18 116.927
R17539 vdd.n27 vdd.n25 116.927
R17540 vdd.n1225 vdd.t55 111.188
R17541 vdd.n953 vdd.t98 111.188
R17542 vdd.n1245 vdd.t69 111.188
R17543 vdd.n944 vdd.t115 111.188
R17544 vdd.n2622 vdd.t111 111.188
R17545 vdd.n805 vdd.t121 111.188
R17546 vdd.n2619 vdd.t101 111.188
R17547 vdd.n769 vdd.t52 111.188
R17548 vdd.n2863 vdd.n898 99.5127
R17549 vdd.n2863 vdd.n896 99.5127
R17550 vdd.n2867 vdd.n896 99.5127
R17551 vdd.n2867 vdd.n887 99.5127
R17552 vdd.n2875 vdd.n887 99.5127
R17553 vdd.n2875 vdd.n885 99.5127
R17554 vdd.n2879 vdd.n885 99.5127
R17555 vdd.n2879 vdd.n875 99.5127
R17556 vdd.n2887 vdd.n875 99.5127
R17557 vdd.n2887 vdd.n873 99.5127
R17558 vdd.n2891 vdd.n873 99.5127
R17559 vdd.n2891 vdd.n863 99.5127
R17560 vdd.n2899 vdd.n863 99.5127
R17561 vdd.n2899 vdd.n861 99.5127
R17562 vdd.n2903 vdd.n861 99.5127
R17563 vdd.n2903 vdd.n852 99.5127
R17564 vdd.n2911 vdd.n852 99.5127
R17565 vdd.n2911 vdd.n850 99.5127
R17566 vdd.n2915 vdd.n850 99.5127
R17567 vdd.n2915 vdd.n838 99.5127
R17568 vdd.n2924 vdd.n838 99.5127
R17569 vdd.n2924 vdd.n836 99.5127
R17570 vdd.n2928 vdd.n836 99.5127
R17571 vdd.n2928 vdd.n827 99.5127
R17572 vdd.n2936 vdd.n827 99.5127
R17573 vdd.n2936 vdd.n825 99.5127
R17574 vdd.n2940 vdd.n825 99.5127
R17575 vdd.n2940 vdd.n813 99.5127
R17576 vdd.n2993 vdd.n813 99.5127
R17577 vdd.n2993 vdd.n811 99.5127
R17578 vdd.n2997 vdd.n811 99.5127
R17579 vdd.n2997 vdd.n777 99.5127
R17580 vdd.n3067 vdd.n777 99.5127
R17581 vdd.n3063 vdd.n778 99.5127
R17582 vdd.n3061 vdd.n3060 99.5127
R17583 vdd.n3058 vdd.n782 99.5127
R17584 vdd.n3054 vdd.n3053 99.5127
R17585 vdd.n3051 vdd.n785 99.5127
R17586 vdd.n3047 vdd.n3046 99.5127
R17587 vdd.n3044 vdd.n788 99.5127
R17588 vdd.n3040 vdd.n3039 99.5127
R17589 vdd.n3037 vdd.n791 99.5127
R17590 vdd.n3032 vdd.n3031 99.5127
R17591 vdd.n3029 vdd.n794 99.5127
R17592 vdd.n3025 vdd.n3024 99.5127
R17593 vdd.n3022 vdd.n797 99.5127
R17594 vdd.n3018 vdd.n3017 99.5127
R17595 vdd.n3015 vdd.n800 99.5127
R17596 vdd.n3011 vdd.n3010 99.5127
R17597 vdd.n3008 vdd.n803 99.5127
R17598 vdd.n2784 vdd.n900 99.5127
R17599 vdd.n2780 vdd.n900 99.5127
R17600 vdd.n2780 vdd.n894 99.5127
R17601 vdd.n2724 vdd.n894 99.5127
R17602 vdd.n2724 vdd.n889 99.5127
R17603 vdd.n2727 vdd.n889 99.5127
R17604 vdd.n2727 vdd.n883 99.5127
R17605 vdd.n2730 vdd.n883 99.5127
R17606 vdd.n2730 vdd.n877 99.5127
R17607 vdd.n2763 vdd.n877 99.5127
R17608 vdd.n2763 vdd.n870 99.5127
R17609 vdd.n2759 vdd.n870 99.5127
R17610 vdd.n2759 vdd.n864 99.5127
R17611 vdd.n2756 vdd.n864 99.5127
R17612 vdd.n2756 vdd.n859 99.5127
R17613 vdd.n2753 vdd.n859 99.5127
R17614 vdd.n2753 vdd.n854 99.5127
R17615 vdd.n2750 vdd.n854 99.5127
R17616 vdd.n2750 vdd.n847 99.5127
R17617 vdd.n2747 vdd.n847 99.5127
R17618 vdd.n2747 vdd.n839 99.5127
R17619 vdd.n2744 vdd.n839 99.5127
R17620 vdd.n2744 vdd.n834 99.5127
R17621 vdd.n2741 vdd.n834 99.5127
R17622 vdd.n2741 vdd.n829 99.5127
R17623 vdd.n2738 vdd.n829 99.5127
R17624 vdd.n2738 vdd.n823 99.5127
R17625 vdd.n2735 vdd.n823 99.5127
R17626 vdd.n2735 vdd.n815 99.5127
R17627 vdd.n815 vdd.n808 99.5127
R17628 vdd.n2999 vdd.n808 99.5127
R17629 vdd.n3000 vdd.n2999 99.5127
R17630 vdd.n3000 vdd.n775 99.5127
R17631 vdd.n2617 vdd.n2616 99.5127
R17632 vdd.n2848 vdd.n2616 99.5127
R17633 vdd.n2846 vdd.n2845 99.5127
R17634 vdd.n2842 vdd.n2841 99.5127
R17635 vdd.n2838 vdd.n2837 99.5127
R17636 vdd.n2834 vdd.n2833 99.5127
R17637 vdd.n2830 vdd.n2829 99.5127
R17638 vdd.n2826 vdd.n2825 99.5127
R17639 vdd.n2822 vdd.n2821 99.5127
R17640 vdd.n2818 vdd.n2817 99.5127
R17641 vdd.n2814 vdd.n2813 99.5127
R17642 vdd.n2810 vdd.n2809 99.5127
R17643 vdd.n2806 vdd.n2805 99.5127
R17644 vdd.n2802 vdd.n2801 99.5127
R17645 vdd.n2798 vdd.n2797 99.5127
R17646 vdd.n2794 vdd.n2793 99.5127
R17647 vdd.n2789 vdd.n2788 99.5127
R17648 vdd.n2581 vdd.n941 99.5127
R17649 vdd.n2577 vdd.n2576 99.5127
R17650 vdd.n2573 vdd.n2572 99.5127
R17651 vdd.n2569 vdd.n2568 99.5127
R17652 vdd.n2565 vdd.n2564 99.5127
R17653 vdd.n2561 vdd.n2560 99.5127
R17654 vdd.n2557 vdd.n2556 99.5127
R17655 vdd.n2553 vdd.n2552 99.5127
R17656 vdd.n2549 vdd.n2548 99.5127
R17657 vdd.n2545 vdd.n2544 99.5127
R17658 vdd.n2541 vdd.n2540 99.5127
R17659 vdd.n2537 vdd.n2536 99.5127
R17660 vdd.n2533 vdd.n2532 99.5127
R17661 vdd.n2529 vdd.n2528 99.5127
R17662 vdd.n2525 vdd.n2524 99.5127
R17663 vdd.n2521 vdd.n2520 99.5127
R17664 vdd.n2516 vdd.n2515 99.5127
R17665 vdd.n1280 vdd.n1048 99.5127
R17666 vdd.n1283 vdd.n1048 99.5127
R17667 vdd.n1283 vdd.n1042 99.5127
R17668 vdd.n1286 vdd.n1042 99.5127
R17669 vdd.n1286 vdd.n1037 99.5127
R17670 vdd.n1289 vdd.n1037 99.5127
R17671 vdd.n1289 vdd.n1031 99.5127
R17672 vdd.n1292 vdd.n1031 99.5127
R17673 vdd.n1292 vdd.n1024 99.5127
R17674 vdd.n1295 vdd.n1024 99.5127
R17675 vdd.n1295 vdd.n1017 99.5127
R17676 vdd.n1298 vdd.n1017 99.5127
R17677 vdd.n1298 vdd.n1011 99.5127
R17678 vdd.n1301 vdd.n1011 99.5127
R17679 vdd.n1301 vdd.n1006 99.5127
R17680 vdd.n1304 vdd.n1006 99.5127
R17681 vdd.n1304 vdd.n1000 99.5127
R17682 vdd.n1329 vdd.n1000 99.5127
R17683 vdd.n1329 vdd.n993 99.5127
R17684 vdd.n1325 vdd.n993 99.5127
R17685 vdd.n1325 vdd.n987 99.5127
R17686 vdd.n1322 vdd.n987 99.5127
R17687 vdd.n1322 vdd.n982 99.5127
R17688 vdd.n1319 vdd.n982 99.5127
R17689 vdd.n1319 vdd.n977 99.5127
R17690 vdd.n1316 vdd.n977 99.5127
R17691 vdd.n1316 vdd.n971 99.5127
R17692 vdd.n1313 vdd.n971 99.5127
R17693 vdd.n1313 vdd.n964 99.5127
R17694 vdd.n1310 vdd.n964 99.5127
R17695 vdd.n1310 vdd.n957 99.5127
R17696 vdd.n957 vdd.n946 99.5127
R17697 vdd.n2511 vdd.n946 99.5127
R17698 vdd.n1089 vdd.n1088 99.5127
R17699 vdd.n2327 vdd.n1088 99.5127
R17700 vdd.n2325 vdd.n2324 99.5127
R17701 vdd.n2321 vdd.n2320 99.5127
R17702 vdd.n2317 vdd.n2316 99.5127
R17703 vdd.n2313 vdd.n2312 99.5127
R17704 vdd.n2309 vdd.n2308 99.5127
R17705 vdd.n2305 vdd.n2304 99.5127
R17706 vdd.n2301 vdd.n2300 99.5127
R17707 vdd.n1247 vdd.n1246 99.5127
R17708 vdd.n1251 vdd.n1250 99.5127
R17709 vdd.n1255 vdd.n1254 99.5127
R17710 vdd.n1259 vdd.n1258 99.5127
R17711 vdd.n1263 vdd.n1262 99.5127
R17712 vdd.n1267 vdd.n1266 99.5127
R17713 vdd.n1271 vdd.n1270 99.5127
R17714 vdd.n1276 vdd.n1275 99.5127
R17715 vdd.n2342 vdd.n1046 99.5127
R17716 vdd.n2342 vdd.n1044 99.5127
R17717 vdd.n2346 vdd.n1044 99.5127
R17718 vdd.n2346 vdd.n1035 99.5127
R17719 vdd.n2354 vdd.n1035 99.5127
R17720 vdd.n2354 vdd.n1033 99.5127
R17721 vdd.n2358 vdd.n1033 99.5127
R17722 vdd.n2358 vdd.n1022 99.5127
R17723 vdd.n2366 vdd.n1022 99.5127
R17724 vdd.n2366 vdd.n1020 99.5127
R17725 vdd.n2370 vdd.n1020 99.5127
R17726 vdd.n2370 vdd.n1010 99.5127
R17727 vdd.n2379 vdd.n1010 99.5127
R17728 vdd.n2379 vdd.n1008 99.5127
R17729 vdd.n2383 vdd.n1008 99.5127
R17730 vdd.n2383 vdd.n998 99.5127
R17731 vdd.n2391 vdd.n998 99.5127
R17732 vdd.n2391 vdd.n996 99.5127
R17733 vdd.n2395 vdd.n996 99.5127
R17734 vdd.n2395 vdd.n986 99.5127
R17735 vdd.n2403 vdd.n986 99.5127
R17736 vdd.n2403 vdd.n984 99.5127
R17737 vdd.n2407 vdd.n984 99.5127
R17738 vdd.n2407 vdd.n975 99.5127
R17739 vdd.n2415 vdd.n975 99.5127
R17740 vdd.n2415 vdd.n973 99.5127
R17741 vdd.n2419 vdd.n973 99.5127
R17742 vdd.n2419 vdd.n962 99.5127
R17743 vdd.n2429 vdd.n962 99.5127
R17744 vdd.n2429 vdd.n959 99.5127
R17745 vdd.n2434 vdd.n959 99.5127
R17746 vdd.n2434 vdd.n960 99.5127
R17747 vdd.n960 vdd.n940 99.5127
R17748 vdd.n2983 vdd.n2982 99.5127
R17749 vdd.n2980 vdd.n2946 99.5127
R17750 vdd.n2976 vdd.n2975 99.5127
R17751 vdd.n2973 vdd.n2949 99.5127
R17752 vdd.n2969 vdd.n2968 99.5127
R17753 vdd.n2966 vdd.n2952 99.5127
R17754 vdd.n2962 vdd.n2961 99.5127
R17755 vdd.n2959 vdd.n2956 99.5127
R17756 vdd.n3100 vdd.n755 99.5127
R17757 vdd.n3098 vdd.n3097 99.5127
R17758 vdd.n3095 vdd.n758 99.5127
R17759 vdd.n3091 vdd.n3090 99.5127
R17760 vdd.n3088 vdd.n761 99.5127
R17761 vdd.n3084 vdd.n3083 99.5127
R17762 vdd.n3081 vdd.n764 99.5127
R17763 vdd.n3077 vdd.n3076 99.5127
R17764 vdd.n3074 vdd.n767 99.5127
R17765 vdd.n2689 vdd.n901 99.5127
R17766 vdd.n2778 vdd.n901 99.5127
R17767 vdd.n2778 vdd.n895 99.5127
R17768 vdd.n2774 vdd.n895 99.5127
R17769 vdd.n2774 vdd.n890 99.5127
R17770 vdd.n2771 vdd.n890 99.5127
R17771 vdd.n2771 vdd.n884 99.5127
R17772 vdd.n2768 vdd.n884 99.5127
R17773 vdd.n2768 vdd.n878 99.5127
R17774 vdd.n2765 vdd.n878 99.5127
R17775 vdd.n2765 vdd.n871 99.5127
R17776 vdd.n2721 vdd.n871 99.5127
R17777 vdd.n2721 vdd.n865 99.5127
R17778 vdd.n2718 vdd.n865 99.5127
R17779 vdd.n2718 vdd.n860 99.5127
R17780 vdd.n2715 vdd.n860 99.5127
R17781 vdd.n2715 vdd.n855 99.5127
R17782 vdd.n2712 vdd.n855 99.5127
R17783 vdd.n2712 vdd.n848 99.5127
R17784 vdd.n2709 vdd.n848 99.5127
R17785 vdd.n2709 vdd.n840 99.5127
R17786 vdd.n2706 vdd.n840 99.5127
R17787 vdd.n2706 vdd.n835 99.5127
R17788 vdd.n2703 vdd.n835 99.5127
R17789 vdd.n2703 vdd.n830 99.5127
R17790 vdd.n2700 vdd.n830 99.5127
R17791 vdd.n2700 vdd.n824 99.5127
R17792 vdd.n2697 vdd.n824 99.5127
R17793 vdd.n2697 vdd.n816 99.5127
R17794 vdd.n2694 vdd.n816 99.5127
R17795 vdd.n2694 vdd.n809 99.5127
R17796 vdd.n809 vdd.n773 99.5127
R17797 vdd.n3069 vdd.n773 99.5127
R17798 vdd.n2624 vdd.n904 99.5127
R17799 vdd.n2628 vdd.n2627 99.5127
R17800 vdd.n2632 vdd.n2631 99.5127
R17801 vdd.n2636 vdd.n2635 99.5127
R17802 vdd.n2640 vdd.n2639 99.5127
R17803 vdd.n2644 vdd.n2643 99.5127
R17804 vdd.n2648 vdd.n2647 99.5127
R17805 vdd.n2652 vdd.n2651 99.5127
R17806 vdd.n2656 vdd.n2655 99.5127
R17807 vdd.n2660 vdd.n2659 99.5127
R17808 vdd.n2664 vdd.n2663 99.5127
R17809 vdd.n2668 vdd.n2667 99.5127
R17810 vdd.n2672 vdd.n2671 99.5127
R17811 vdd.n2676 vdd.n2675 99.5127
R17812 vdd.n2680 vdd.n2679 99.5127
R17813 vdd.n2684 vdd.n2683 99.5127
R17814 vdd.n2686 vdd.n2615 99.5127
R17815 vdd.n2861 vdd.n902 99.5127
R17816 vdd.n2861 vdd.n893 99.5127
R17817 vdd.n2869 vdd.n893 99.5127
R17818 vdd.n2869 vdd.n891 99.5127
R17819 vdd.n2873 vdd.n891 99.5127
R17820 vdd.n2873 vdd.n881 99.5127
R17821 vdd.n2881 vdd.n881 99.5127
R17822 vdd.n2881 vdd.n879 99.5127
R17823 vdd.n2885 vdd.n879 99.5127
R17824 vdd.n2885 vdd.n869 99.5127
R17825 vdd.n2893 vdd.n869 99.5127
R17826 vdd.n2893 vdd.n867 99.5127
R17827 vdd.n2897 vdd.n867 99.5127
R17828 vdd.n2897 vdd.n858 99.5127
R17829 vdd.n2905 vdd.n858 99.5127
R17830 vdd.n2905 vdd.n856 99.5127
R17831 vdd.n2909 vdd.n856 99.5127
R17832 vdd.n2909 vdd.n845 99.5127
R17833 vdd.n2917 vdd.n845 99.5127
R17834 vdd.n2917 vdd.n842 99.5127
R17835 vdd.n2922 vdd.n842 99.5127
R17836 vdd.n2922 vdd.n833 99.5127
R17837 vdd.n2930 vdd.n833 99.5127
R17838 vdd.n2930 vdd.n831 99.5127
R17839 vdd.n2934 vdd.n831 99.5127
R17840 vdd.n2934 vdd.n821 99.5127
R17841 vdd.n2942 vdd.n821 99.5127
R17842 vdd.n2942 vdd.n818 99.5127
R17843 vdd.n2991 vdd.n818 99.5127
R17844 vdd.n2991 vdd.n819 99.5127
R17845 vdd.n819 vdd.n810 99.5127
R17846 vdd.n2986 vdd.n810 99.5127
R17847 vdd.n2986 vdd.n776 99.5127
R17848 vdd.n2505 vdd.n2504 99.5127
R17849 vdd.n2501 vdd.n2500 99.5127
R17850 vdd.n2497 vdd.n2496 99.5127
R17851 vdd.n2493 vdd.n2492 99.5127
R17852 vdd.n2489 vdd.n2488 99.5127
R17853 vdd.n2485 vdd.n2484 99.5127
R17854 vdd.n2481 vdd.n2480 99.5127
R17855 vdd.n2477 vdd.n2476 99.5127
R17856 vdd.n2473 vdd.n2472 99.5127
R17857 vdd.n2469 vdd.n2468 99.5127
R17858 vdd.n2465 vdd.n2464 99.5127
R17859 vdd.n2461 vdd.n2460 99.5127
R17860 vdd.n2457 vdd.n2456 99.5127
R17861 vdd.n2453 vdd.n2452 99.5127
R17862 vdd.n2449 vdd.n2448 99.5127
R17863 vdd.n2445 vdd.n2444 99.5127
R17864 vdd.n2441 vdd.n922 99.5127
R17865 vdd.n1358 vdd.n1049 99.5127
R17866 vdd.n1355 vdd.n1049 99.5127
R17867 vdd.n1355 vdd.n1043 99.5127
R17868 vdd.n1352 vdd.n1043 99.5127
R17869 vdd.n1352 vdd.n1038 99.5127
R17870 vdd.n1349 vdd.n1038 99.5127
R17871 vdd.n1349 vdd.n1032 99.5127
R17872 vdd.n1346 vdd.n1032 99.5127
R17873 vdd.n1346 vdd.n1025 99.5127
R17874 vdd.n1343 vdd.n1025 99.5127
R17875 vdd.n1343 vdd.n1018 99.5127
R17876 vdd.n1340 vdd.n1018 99.5127
R17877 vdd.n1340 vdd.n1012 99.5127
R17878 vdd.n1337 vdd.n1012 99.5127
R17879 vdd.n1337 vdd.n1007 99.5127
R17880 vdd.n1334 vdd.n1007 99.5127
R17881 vdd.n1334 vdd.n1001 99.5127
R17882 vdd.n1331 vdd.n1001 99.5127
R17883 vdd.n1331 vdd.n994 99.5127
R17884 vdd.n1241 vdd.n994 99.5127
R17885 vdd.n1241 vdd.n988 99.5127
R17886 vdd.n1238 vdd.n988 99.5127
R17887 vdd.n1238 vdd.n983 99.5127
R17888 vdd.n1235 vdd.n983 99.5127
R17889 vdd.n1235 vdd.n978 99.5127
R17890 vdd.n1232 vdd.n978 99.5127
R17891 vdd.n1232 vdd.n972 99.5127
R17892 vdd.n1229 vdd.n972 99.5127
R17893 vdd.n1229 vdd.n965 99.5127
R17894 vdd.n965 vdd.n956 99.5127
R17895 vdd.n2436 vdd.n956 99.5127
R17896 vdd.n2437 vdd.n2436 99.5127
R17897 vdd.n2437 vdd.n948 99.5127
R17898 vdd.n1193 vdd.n1053 99.5127
R17899 vdd.n1197 vdd.n1196 99.5127
R17900 vdd.n1201 vdd.n1200 99.5127
R17901 vdd.n1205 vdd.n1204 99.5127
R17902 vdd.n1209 vdd.n1208 99.5127
R17903 vdd.n1213 vdd.n1212 99.5127
R17904 vdd.n1217 vdd.n1216 99.5127
R17905 vdd.n1221 vdd.n1220 99.5127
R17906 vdd.n1391 vdd.n1223 99.5127
R17907 vdd.n1389 vdd.n1388 99.5127
R17908 vdd.n1385 vdd.n1384 99.5127
R17909 vdd.n1381 vdd.n1380 99.5127
R17910 vdd.n1377 vdd.n1376 99.5127
R17911 vdd.n1373 vdd.n1372 99.5127
R17912 vdd.n1369 vdd.n1368 99.5127
R17913 vdd.n1365 vdd.n1364 99.5127
R17914 vdd.n1361 vdd.n1087 99.5127
R17915 vdd.n2340 vdd.n1051 99.5127
R17916 vdd.n2340 vdd.n1041 99.5127
R17917 vdd.n2348 vdd.n1041 99.5127
R17918 vdd.n2348 vdd.n1039 99.5127
R17919 vdd.n2352 vdd.n1039 99.5127
R17920 vdd.n2352 vdd.n1029 99.5127
R17921 vdd.n2360 vdd.n1029 99.5127
R17922 vdd.n2360 vdd.n1027 99.5127
R17923 vdd.n2364 vdd.n1027 99.5127
R17924 vdd.n2364 vdd.n1016 99.5127
R17925 vdd.n2372 vdd.n1016 99.5127
R17926 vdd.n2372 vdd.n1013 99.5127
R17927 vdd.n2377 vdd.n1013 99.5127
R17928 vdd.n2377 vdd.n1004 99.5127
R17929 vdd.n2385 vdd.n1004 99.5127
R17930 vdd.n2385 vdd.n1002 99.5127
R17931 vdd.n2389 vdd.n1002 99.5127
R17932 vdd.n2389 vdd.n992 99.5127
R17933 vdd.n2397 vdd.n992 99.5127
R17934 vdd.n2397 vdd.n990 99.5127
R17935 vdd.n2401 vdd.n990 99.5127
R17936 vdd.n2401 vdd.n981 99.5127
R17937 vdd.n2409 vdd.n981 99.5127
R17938 vdd.n2409 vdd.n979 99.5127
R17939 vdd.n2413 vdd.n979 99.5127
R17940 vdd.n2413 vdd.n969 99.5127
R17941 vdd.n2421 vdd.n969 99.5127
R17942 vdd.n2421 vdd.n966 99.5127
R17943 vdd.n2427 vdd.n966 99.5127
R17944 vdd.n2427 vdd.n967 99.5127
R17945 vdd.n967 vdd.n958 99.5127
R17946 vdd.n958 vdd.n949 99.5127
R17947 vdd.n2509 vdd.n949 99.5127
R17948 vdd.n9 vdd.n7 98.9633
R17949 vdd.n2 vdd.n0 98.9633
R17950 vdd.n9 vdd.n8 98.6055
R17951 vdd.n11 vdd.n10 98.6055
R17952 vdd.n13 vdd.n12 98.6055
R17953 vdd.n6 vdd.n5 98.6055
R17954 vdd.n4 vdd.n3 98.6055
R17955 vdd.n2 vdd.n1 98.6055
R17956 vdd.t243 vdd.n291 85.8723
R17957 vdd.t220 vdd.n236 85.8723
R17958 vdd.t233 vdd.n193 85.8723
R17959 vdd.t210 vdd.n138 85.8723
R17960 vdd.t195 vdd.n96 85.8723
R17961 vdd.t178 vdd.n41 85.8723
R17962 vdd.t254 vdd.n2022 85.8723
R17963 vdd.t166 vdd.n2077 85.8723
R17964 vdd.t246 vdd.n1924 85.8723
R17965 vdd.t143 vdd.n1979 85.8723
R17966 vdd.t173 vdd.n1827 85.8723
R17967 vdd.t196 vdd.n1882 85.8723
R17968 vdd.n2920 vdd.n843 78.546
R17969 vdd.n2375 vdd.n1014 78.546
R17970 vdd.n278 vdd.n277 75.1835
R17971 vdd.n276 vdd.n275 75.1835
R17972 vdd.n274 vdd.n273 75.1835
R17973 vdd.n272 vdd.n271 75.1835
R17974 vdd.n270 vdd.n269 75.1835
R17975 vdd.n268 vdd.n267 75.1835
R17976 vdd.n266 vdd.n265 75.1835
R17977 vdd.n180 vdd.n179 75.1835
R17978 vdd.n178 vdd.n177 75.1835
R17979 vdd.n176 vdd.n175 75.1835
R17980 vdd.n174 vdd.n173 75.1835
R17981 vdd.n172 vdd.n171 75.1835
R17982 vdd.n170 vdd.n169 75.1835
R17983 vdd.n168 vdd.n167 75.1835
R17984 vdd.n83 vdd.n82 75.1835
R17985 vdd.n81 vdd.n80 75.1835
R17986 vdd.n79 vdd.n78 75.1835
R17987 vdd.n77 vdd.n76 75.1835
R17988 vdd.n75 vdd.n74 75.1835
R17989 vdd.n73 vdd.n72 75.1835
R17990 vdd.n71 vdd.n70 75.1835
R17991 vdd.n2052 vdd.n2051 75.1835
R17992 vdd.n2054 vdd.n2053 75.1835
R17993 vdd.n2056 vdd.n2055 75.1835
R17994 vdd.n2058 vdd.n2057 75.1835
R17995 vdd.n2060 vdd.n2059 75.1835
R17996 vdd.n2062 vdd.n2061 75.1835
R17997 vdd.n2064 vdd.n2063 75.1835
R17998 vdd.n1954 vdd.n1953 75.1835
R17999 vdd.n1956 vdd.n1955 75.1835
R18000 vdd.n1958 vdd.n1957 75.1835
R18001 vdd.n1960 vdd.n1959 75.1835
R18002 vdd.n1962 vdd.n1961 75.1835
R18003 vdd.n1964 vdd.n1963 75.1835
R18004 vdd.n1966 vdd.n1965 75.1835
R18005 vdd.n1857 vdd.n1856 75.1835
R18006 vdd.n1859 vdd.n1858 75.1835
R18007 vdd.n1861 vdd.n1860 75.1835
R18008 vdd.n1863 vdd.n1862 75.1835
R18009 vdd.n1865 vdd.n1864 75.1835
R18010 vdd.n1867 vdd.n1866 75.1835
R18011 vdd.n1869 vdd.n1868 75.1835
R18012 vdd.n2856 vdd.n2855 72.8958
R18013 vdd.n2855 vdd.n2599 72.8958
R18014 vdd.n2855 vdd.n2600 72.8958
R18015 vdd.n2855 vdd.n2601 72.8958
R18016 vdd.n2855 vdd.n2602 72.8958
R18017 vdd.n2855 vdd.n2603 72.8958
R18018 vdd.n2855 vdd.n2604 72.8958
R18019 vdd.n2855 vdd.n2605 72.8958
R18020 vdd.n2855 vdd.n2606 72.8958
R18021 vdd.n2855 vdd.n2607 72.8958
R18022 vdd.n2855 vdd.n2608 72.8958
R18023 vdd.n2855 vdd.n2609 72.8958
R18024 vdd.n2855 vdd.n2610 72.8958
R18025 vdd.n2855 vdd.n2611 72.8958
R18026 vdd.n2855 vdd.n2612 72.8958
R18027 vdd.n2855 vdd.n2613 72.8958
R18028 vdd.n2855 vdd.n2614 72.8958
R18029 vdd.n772 vdd.n756 72.8958
R18030 vdd.n3075 vdd.n756 72.8958
R18031 vdd.n766 vdd.n756 72.8958
R18032 vdd.n3082 vdd.n756 72.8958
R18033 vdd.n763 vdd.n756 72.8958
R18034 vdd.n3089 vdd.n756 72.8958
R18035 vdd.n760 vdd.n756 72.8958
R18036 vdd.n3096 vdd.n756 72.8958
R18037 vdd.n3099 vdd.n756 72.8958
R18038 vdd.n2955 vdd.n756 72.8958
R18039 vdd.n2960 vdd.n756 72.8958
R18040 vdd.n2954 vdd.n756 72.8958
R18041 vdd.n2967 vdd.n756 72.8958
R18042 vdd.n2951 vdd.n756 72.8958
R18043 vdd.n2974 vdd.n756 72.8958
R18044 vdd.n2948 vdd.n756 72.8958
R18045 vdd.n2981 vdd.n756 72.8958
R18046 vdd.n2334 vdd.n2333 72.8958
R18047 vdd.n2334 vdd.n1055 72.8958
R18048 vdd.n2334 vdd.n1056 72.8958
R18049 vdd.n2334 vdd.n1057 72.8958
R18050 vdd.n2334 vdd.n1058 72.8958
R18051 vdd.n2334 vdd.n1059 72.8958
R18052 vdd.n2334 vdd.n1060 72.8958
R18053 vdd.n2334 vdd.n1061 72.8958
R18054 vdd.n2334 vdd.n1062 72.8958
R18055 vdd.n2334 vdd.n1063 72.8958
R18056 vdd.n2334 vdd.n1064 72.8958
R18057 vdd.n2334 vdd.n1065 72.8958
R18058 vdd.n2334 vdd.n1066 72.8958
R18059 vdd.n2334 vdd.n1067 72.8958
R18060 vdd.n2334 vdd.n1068 72.8958
R18061 vdd.n2334 vdd.n1069 72.8958
R18062 vdd.n2334 vdd.n1070 72.8958
R18063 vdd.n2582 vdd.n923 72.8958
R18064 vdd.n2582 vdd.n924 72.8958
R18065 vdd.n2582 vdd.n925 72.8958
R18066 vdd.n2582 vdd.n926 72.8958
R18067 vdd.n2582 vdd.n927 72.8958
R18068 vdd.n2582 vdd.n928 72.8958
R18069 vdd.n2582 vdd.n929 72.8958
R18070 vdd.n2582 vdd.n930 72.8958
R18071 vdd.n2582 vdd.n931 72.8958
R18072 vdd.n2582 vdd.n932 72.8958
R18073 vdd.n2582 vdd.n933 72.8958
R18074 vdd.n2582 vdd.n934 72.8958
R18075 vdd.n2582 vdd.n935 72.8958
R18076 vdd.n2582 vdd.n936 72.8958
R18077 vdd.n2582 vdd.n937 72.8958
R18078 vdd.n2582 vdd.n938 72.8958
R18079 vdd.n2582 vdd.n939 72.8958
R18080 vdd.n2855 vdd.n2854 72.8958
R18081 vdd.n2855 vdd.n2583 72.8958
R18082 vdd.n2855 vdd.n2584 72.8958
R18083 vdd.n2855 vdd.n2585 72.8958
R18084 vdd.n2855 vdd.n2586 72.8958
R18085 vdd.n2855 vdd.n2587 72.8958
R18086 vdd.n2855 vdd.n2588 72.8958
R18087 vdd.n2855 vdd.n2589 72.8958
R18088 vdd.n2855 vdd.n2590 72.8958
R18089 vdd.n2855 vdd.n2591 72.8958
R18090 vdd.n2855 vdd.n2592 72.8958
R18091 vdd.n2855 vdd.n2593 72.8958
R18092 vdd.n2855 vdd.n2594 72.8958
R18093 vdd.n2855 vdd.n2595 72.8958
R18094 vdd.n2855 vdd.n2596 72.8958
R18095 vdd.n2855 vdd.n2597 72.8958
R18096 vdd.n2855 vdd.n2598 72.8958
R18097 vdd.n3003 vdd.n756 72.8958
R18098 vdd.n3009 vdd.n756 72.8958
R18099 vdd.n802 vdd.n756 72.8958
R18100 vdd.n3016 vdd.n756 72.8958
R18101 vdd.n799 vdd.n756 72.8958
R18102 vdd.n3023 vdd.n756 72.8958
R18103 vdd.n796 vdd.n756 72.8958
R18104 vdd.n3030 vdd.n756 72.8958
R18105 vdd.n793 vdd.n756 72.8958
R18106 vdd.n3038 vdd.n756 72.8958
R18107 vdd.n790 vdd.n756 72.8958
R18108 vdd.n3045 vdd.n756 72.8958
R18109 vdd.n787 vdd.n756 72.8958
R18110 vdd.n3052 vdd.n756 72.8958
R18111 vdd.n784 vdd.n756 72.8958
R18112 vdd.n3059 vdd.n756 72.8958
R18113 vdd.n3062 vdd.n756 72.8958
R18114 vdd.n2582 vdd.n921 72.8958
R18115 vdd.n2582 vdd.n920 72.8958
R18116 vdd.n2582 vdd.n919 72.8958
R18117 vdd.n2582 vdd.n918 72.8958
R18118 vdd.n2582 vdd.n917 72.8958
R18119 vdd.n2582 vdd.n916 72.8958
R18120 vdd.n2582 vdd.n915 72.8958
R18121 vdd.n2582 vdd.n914 72.8958
R18122 vdd.n2582 vdd.n913 72.8958
R18123 vdd.n2582 vdd.n912 72.8958
R18124 vdd.n2582 vdd.n911 72.8958
R18125 vdd.n2582 vdd.n910 72.8958
R18126 vdd.n2582 vdd.n909 72.8958
R18127 vdd.n2582 vdd.n908 72.8958
R18128 vdd.n2582 vdd.n907 72.8958
R18129 vdd.n2582 vdd.n906 72.8958
R18130 vdd.n2582 vdd.n905 72.8958
R18131 vdd.n2335 vdd.n2334 72.8958
R18132 vdd.n2334 vdd.n1071 72.8958
R18133 vdd.n2334 vdd.n1072 72.8958
R18134 vdd.n2334 vdd.n1073 72.8958
R18135 vdd.n2334 vdd.n1074 72.8958
R18136 vdd.n2334 vdd.n1075 72.8958
R18137 vdd.n2334 vdd.n1076 72.8958
R18138 vdd.n2334 vdd.n1077 72.8958
R18139 vdd.n2334 vdd.n1078 72.8958
R18140 vdd.n2334 vdd.n1079 72.8958
R18141 vdd.n2334 vdd.n1080 72.8958
R18142 vdd.n2334 vdd.n1081 72.8958
R18143 vdd.n2334 vdd.n1082 72.8958
R18144 vdd.n2334 vdd.n1083 72.8958
R18145 vdd.n2334 vdd.n1084 72.8958
R18146 vdd.n2334 vdd.n1085 72.8958
R18147 vdd.n2334 vdd.n1086 72.8958
R18148 vdd.n1736 vdd.n1735 66.2847
R18149 vdd.n1736 vdd.n1514 66.2847
R18150 vdd.n1736 vdd.n1515 66.2847
R18151 vdd.n1736 vdd.n1516 66.2847
R18152 vdd.n1736 vdd.n1517 66.2847
R18153 vdd.n1736 vdd.n1518 66.2847
R18154 vdd.n1736 vdd.n1519 66.2847
R18155 vdd.n1736 vdd.n1520 66.2847
R18156 vdd.n1736 vdd.n1521 66.2847
R18157 vdd.n1736 vdd.n1522 66.2847
R18158 vdd.n1736 vdd.n1523 66.2847
R18159 vdd.n1736 vdd.n1524 66.2847
R18160 vdd.n1736 vdd.n1525 66.2847
R18161 vdd.n1736 vdd.n1526 66.2847
R18162 vdd.n1736 vdd.n1527 66.2847
R18163 vdd.n1736 vdd.n1528 66.2847
R18164 vdd.n1736 vdd.n1529 66.2847
R18165 vdd.n1736 vdd.n1530 66.2847
R18166 vdd.n1736 vdd.n1531 66.2847
R18167 vdd.n1736 vdd.n1532 66.2847
R18168 vdd.n1736 vdd.n1533 66.2847
R18169 vdd.n1736 vdd.n1534 66.2847
R18170 vdd.n1736 vdd.n1535 66.2847
R18171 vdd.n1736 vdd.n1536 66.2847
R18172 vdd.n1736 vdd.n1537 66.2847
R18173 vdd.n1736 vdd.n1538 66.2847
R18174 vdd.n1736 vdd.n1539 66.2847
R18175 vdd.n1736 vdd.n1540 66.2847
R18176 vdd.n1736 vdd.n1541 66.2847
R18177 vdd.n1736 vdd.n1542 66.2847
R18178 vdd.n1736 vdd.n1543 66.2847
R18179 vdd.n1404 vdd.n1054 66.2847
R18180 vdd.n1401 vdd.n1054 66.2847
R18181 vdd.n1397 vdd.n1054 66.2847
R18182 vdd.n2196 vdd.n1054 66.2847
R18183 vdd.n1188 vdd.n1054 66.2847
R18184 vdd.n2203 vdd.n1054 66.2847
R18185 vdd.n1181 vdd.n1054 66.2847
R18186 vdd.n2210 vdd.n1054 66.2847
R18187 vdd.n1174 vdd.n1054 66.2847
R18188 vdd.n2217 vdd.n1054 66.2847
R18189 vdd.n1168 vdd.n1054 66.2847
R18190 vdd.n1163 vdd.n1054 66.2847
R18191 vdd.n2228 vdd.n1054 66.2847
R18192 vdd.n1155 vdd.n1054 66.2847
R18193 vdd.n2235 vdd.n1054 66.2847
R18194 vdd.n1148 vdd.n1054 66.2847
R18195 vdd.n2242 vdd.n1054 66.2847
R18196 vdd.n1141 vdd.n1054 66.2847
R18197 vdd.n2249 vdd.n1054 66.2847
R18198 vdd.n1134 vdd.n1054 66.2847
R18199 vdd.n2256 vdd.n1054 66.2847
R18200 vdd.n1128 vdd.n1054 66.2847
R18201 vdd.n1123 vdd.n1054 66.2847
R18202 vdd.n2267 vdd.n1054 66.2847
R18203 vdd.n1115 vdd.n1054 66.2847
R18204 vdd.n2274 vdd.n1054 66.2847
R18205 vdd.n1108 vdd.n1054 66.2847
R18206 vdd.n2281 vdd.n1054 66.2847
R18207 vdd.n1101 vdd.n1054 66.2847
R18208 vdd.n2288 vdd.n1054 66.2847
R18209 vdd.n2293 vdd.n1054 66.2847
R18210 vdd.n1097 vdd.n1054 66.2847
R18211 vdd.n3229 vdd.n658 66.2847
R18212 vdd.n663 vdd.n658 66.2847
R18213 vdd.n666 vdd.n658 66.2847
R18214 vdd.n3218 vdd.n658 66.2847
R18215 vdd.n3212 vdd.n658 66.2847
R18216 vdd.n3210 vdd.n658 66.2847
R18217 vdd.n3204 vdd.n658 66.2847
R18218 vdd.n3202 vdd.n658 66.2847
R18219 vdd.n3196 vdd.n658 66.2847
R18220 vdd.n3194 vdd.n658 66.2847
R18221 vdd.n3188 vdd.n658 66.2847
R18222 vdd.n3186 vdd.n658 66.2847
R18223 vdd.n3180 vdd.n658 66.2847
R18224 vdd.n3178 vdd.n658 66.2847
R18225 vdd.n3172 vdd.n658 66.2847
R18226 vdd.n3170 vdd.n658 66.2847
R18227 vdd.n3164 vdd.n658 66.2847
R18228 vdd.n3162 vdd.n658 66.2847
R18229 vdd.n3156 vdd.n658 66.2847
R18230 vdd.n3154 vdd.n658 66.2847
R18231 vdd.n727 vdd.n658 66.2847
R18232 vdd.n3145 vdd.n658 66.2847
R18233 vdd.n729 vdd.n658 66.2847
R18234 vdd.n3138 vdd.n658 66.2847
R18235 vdd.n3132 vdd.n658 66.2847
R18236 vdd.n3130 vdd.n658 66.2847
R18237 vdd.n3124 vdd.n658 66.2847
R18238 vdd.n3122 vdd.n658 66.2847
R18239 vdd.n3116 vdd.n658 66.2847
R18240 vdd.n750 vdd.n658 66.2847
R18241 vdd.n752 vdd.n658 66.2847
R18242 vdd.n3345 vdd.n3344 66.2847
R18243 vdd.n3345 vdd.n403 66.2847
R18244 vdd.n3345 vdd.n402 66.2847
R18245 vdd.n3345 vdd.n401 66.2847
R18246 vdd.n3345 vdd.n400 66.2847
R18247 vdd.n3345 vdd.n399 66.2847
R18248 vdd.n3345 vdd.n398 66.2847
R18249 vdd.n3345 vdd.n397 66.2847
R18250 vdd.n3345 vdd.n396 66.2847
R18251 vdd.n3345 vdd.n395 66.2847
R18252 vdd.n3345 vdd.n394 66.2847
R18253 vdd.n3345 vdd.n393 66.2847
R18254 vdd.n3345 vdd.n392 66.2847
R18255 vdd.n3345 vdd.n391 66.2847
R18256 vdd.n3345 vdd.n390 66.2847
R18257 vdd.n3345 vdd.n389 66.2847
R18258 vdd.n3345 vdd.n388 66.2847
R18259 vdd.n3345 vdd.n387 66.2847
R18260 vdd.n3345 vdd.n386 66.2847
R18261 vdd.n3345 vdd.n385 66.2847
R18262 vdd.n3345 vdd.n384 66.2847
R18263 vdd.n3345 vdd.n383 66.2847
R18264 vdd.n3345 vdd.n382 66.2847
R18265 vdd.n3345 vdd.n381 66.2847
R18266 vdd.n3345 vdd.n380 66.2847
R18267 vdd.n3345 vdd.n379 66.2847
R18268 vdd.n3345 vdd.n378 66.2847
R18269 vdd.n3345 vdd.n377 66.2847
R18270 vdd.n3345 vdd.n376 66.2847
R18271 vdd.n3345 vdd.n375 66.2847
R18272 vdd.n3345 vdd.n374 66.2847
R18273 vdd.n3345 vdd.n373 66.2847
R18274 vdd.n448 vdd.n373 52.4337
R18275 vdd.n454 vdd.n374 52.4337
R18276 vdd.n458 vdd.n375 52.4337
R18277 vdd.n464 vdd.n376 52.4337
R18278 vdd.n468 vdd.n377 52.4337
R18279 vdd.n474 vdd.n378 52.4337
R18280 vdd.n478 vdd.n379 52.4337
R18281 vdd.n484 vdd.n380 52.4337
R18282 vdd.n488 vdd.n381 52.4337
R18283 vdd.n494 vdd.n382 52.4337
R18284 vdd.n498 vdd.n383 52.4337
R18285 vdd.n504 vdd.n384 52.4337
R18286 vdd.n508 vdd.n385 52.4337
R18287 vdd.n514 vdd.n386 52.4337
R18288 vdd.n518 vdd.n387 52.4337
R18289 vdd.n524 vdd.n388 52.4337
R18290 vdd.n528 vdd.n389 52.4337
R18291 vdd.n534 vdd.n390 52.4337
R18292 vdd.n538 vdd.n391 52.4337
R18293 vdd.n544 vdd.n392 52.4337
R18294 vdd.n548 vdd.n393 52.4337
R18295 vdd.n554 vdd.n394 52.4337
R18296 vdd.n558 vdd.n395 52.4337
R18297 vdd.n564 vdd.n396 52.4337
R18298 vdd.n568 vdd.n397 52.4337
R18299 vdd.n574 vdd.n398 52.4337
R18300 vdd.n578 vdd.n399 52.4337
R18301 vdd.n584 vdd.n400 52.4337
R18302 vdd.n588 vdd.n401 52.4337
R18303 vdd.n594 vdd.n402 52.4337
R18304 vdd.n597 vdd.n403 52.4337
R18305 vdd.n3344 vdd.n3343 52.4337
R18306 vdd.n3229 vdd.n660 52.4337
R18307 vdd.n3227 vdd.n663 52.4337
R18308 vdd.n3223 vdd.n666 52.4337
R18309 vdd.n3219 vdd.n3218 52.4337
R18310 vdd.n3212 vdd.n669 52.4337
R18311 vdd.n3211 vdd.n3210 52.4337
R18312 vdd.n3204 vdd.n675 52.4337
R18313 vdd.n3203 vdd.n3202 52.4337
R18314 vdd.n3196 vdd.n681 52.4337
R18315 vdd.n3195 vdd.n3194 52.4337
R18316 vdd.n3188 vdd.n689 52.4337
R18317 vdd.n3187 vdd.n3186 52.4337
R18318 vdd.n3180 vdd.n695 52.4337
R18319 vdd.n3179 vdd.n3178 52.4337
R18320 vdd.n3172 vdd.n701 52.4337
R18321 vdd.n3171 vdd.n3170 52.4337
R18322 vdd.n3164 vdd.n707 52.4337
R18323 vdd.n3163 vdd.n3162 52.4337
R18324 vdd.n3156 vdd.n713 52.4337
R18325 vdd.n3155 vdd.n3154 52.4337
R18326 vdd.n727 vdd.n719 52.4337
R18327 vdd.n3146 vdd.n3145 52.4337
R18328 vdd.n3143 vdd.n729 52.4337
R18329 vdd.n3139 vdd.n3138 52.4337
R18330 vdd.n3132 vdd.n733 52.4337
R18331 vdd.n3131 vdd.n3130 52.4337
R18332 vdd.n3124 vdd.n739 52.4337
R18333 vdd.n3123 vdd.n3122 52.4337
R18334 vdd.n3116 vdd.n745 52.4337
R18335 vdd.n3115 vdd.n750 52.4337
R18336 vdd.n3111 vdd.n752 52.4337
R18337 vdd.n2295 vdd.n1097 52.4337
R18338 vdd.n2293 vdd.n2292 52.4337
R18339 vdd.n2288 vdd.n2287 52.4337
R18340 vdd.n2283 vdd.n1101 52.4337
R18341 vdd.n2281 vdd.n2280 52.4337
R18342 vdd.n2276 vdd.n1108 52.4337
R18343 vdd.n2274 vdd.n2273 52.4337
R18344 vdd.n2269 vdd.n1115 52.4337
R18345 vdd.n2267 vdd.n2266 52.4337
R18346 vdd.n1124 vdd.n1123 52.4337
R18347 vdd.n2258 vdd.n1128 52.4337
R18348 vdd.n2256 vdd.n2255 52.4337
R18349 vdd.n2251 vdd.n1134 52.4337
R18350 vdd.n2249 vdd.n2248 52.4337
R18351 vdd.n2244 vdd.n1141 52.4337
R18352 vdd.n2242 vdd.n2241 52.4337
R18353 vdd.n2237 vdd.n1148 52.4337
R18354 vdd.n2235 vdd.n2234 52.4337
R18355 vdd.n2230 vdd.n1155 52.4337
R18356 vdd.n2228 vdd.n2227 52.4337
R18357 vdd.n1164 vdd.n1163 52.4337
R18358 vdd.n2219 vdd.n1168 52.4337
R18359 vdd.n2217 vdd.n2216 52.4337
R18360 vdd.n2212 vdd.n1174 52.4337
R18361 vdd.n2210 vdd.n2209 52.4337
R18362 vdd.n2205 vdd.n1181 52.4337
R18363 vdd.n2203 vdd.n2202 52.4337
R18364 vdd.n2198 vdd.n1188 52.4337
R18365 vdd.n2196 vdd.n2195 52.4337
R18366 vdd.n1398 vdd.n1397 52.4337
R18367 vdd.n1402 vdd.n1401 52.4337
R18368 vdd.n2184 vdd.n1404 52.4337
R18369 vdd.n1735 vdd.n1734 52.4337
R18370 vdd.n1549 vdd.n1514 52.4337
R18371 vdd.n1551 vdd.n1515 52.4337
R18372 vdd.n1555 vdd.n1516 52.4337
R18373 vdd.n1557 vdd.n1517 52.4337
R18374 vdd.n1561 vdd.n1518 52.4337
R18375 vdd.n1563 vdd.n1519 52.4337
R18376 vdd.n1567 vdd.n1520 52.4337
R18377 vdd.n1569 vdd.n1521 52.4337
R18378 vdd.n1701 vdd.n1522 52.4337
R18379 vdd.n1573 vdd.n1523 52.4337
R18380 vdd.n1577 vdd.n1524 52.4337
R18381 vdd.n1579 vdd.n1525 52.4337
R18382 vdd.n1583 vdd.n1526 52.4337
R18383 vdd.n1585 vdd.n1527 52.4337
R18384 vdd.n1589 vdd.n1528 52.4337
R18385 vdd.n1591 vdd.n1529 52.4337
R18386 vdd.n1595 vdd.n1530 52.4337
R18387 vdd.n1597 vdd.n1531 52.4337
R18388 vdd.n1601 vdd.n1532 52.4337
R18389 vdd.n1665 vdd.n1533 52.4337
R18390 vdd.n1606 vdd.n1534 52.4337
R18391 vdd.n1608 vdd.n1535 52.4337
R18392 vdd.n1612 vdd.n1536 52.4337
R18393 vdd.n1614 vdd.n1537 52.4337
R18394 vdd.n1618 vdd.n1538 52.4337
R18395 vdd.n1620 vdd.n1539 52.4337
R18396 vdd.n1624 vdd.n1540 52.4337
R18397 vdd.n1626 vdd.n1541 52.4337
R18398 vdd.n1630 vdd.n1542 52.4337
R18399 vdd.n1632 vdd.n1543 52.4337
R18400 vdd.n1735 vdd.n1545 52.4337
R18401 vdd.n1550 vdd.n1514 52.4337
R18402 vdd.n1554 vdd.n1515 52.4337
R18403 vdd.n1556 vdd.n1516 52.4337
R18404 vdd.n1560 vdd.n1517 52.4337
R18405 vdd.n1562 vdd.n1518 52.4337
R18406 vdd.n1566 vdd.n1519 52.4337
R18407 vdd.n1568 vdd.n1520 52.4337
R18408 vdd.n1700 vdd.n1521 52.4337
R18409 vdd.n1572 vdd.n1522 52.4337
R18410 vdd.n1576 vdd.n1523 52.4337
R18411 vdd.n1578 vdd.n1524 52.4337
R18412 vdd.n1582 vdd.n1525 52.4337
R18413 vdd.n1584 vdd.n1526 52.4337
R18414 vdd.n1588 vdd.n1527 52.4337
R18415 vdd.n1590 vdd.n1528 52.4337
R18416 vdd.n1594 vdd.n1529 52.4337
R18417 vdd.n1596 vdd.n1530 52.4337
R18418 vdd.n1600 vdd.n1531 52.4337
R18419 vdd.n1602 vdd.n1532 52.4337
R18420 vdd.n1605 vdd.n1533 52.4337
R18421 vdd.n1607 vdd.n1534 52.4337
R18422 vdd.n1611 vdd.n1535 52.4337
R18423 vdd.n1613 vdd.n1536 52.4337
R18424 vdd.n1617 vdd.n1537 52.4337
R18425 vdd.n1619 vdd.n1538 52.4337
R18426 vdd.n1623 vdd.n1539 52.4337
R18427 vdd.n1625 vdd.n1540 52.4337
R18428 vdd.n1629 vdd.n1541 52.4337
R18429 vdd.n1631 vdd.n1542 52.4337
R18430 vdd.n1543 vdd.n1513 52.4337
R18431 vdd.n1404 vdd.n1403 52.4337
R18432 vdd.n1401 vdd.n1400 52.4337
R18433 vdd.n1397 vdd.n1189 52.4337
R18434 vdd.n2197 vdd.n2196 52.4337
R18435 vdd.n1188 vdd.n1182 52.4337
R18436 vdd.n2204 vdd.n2203 52.4337
R18437 vdd.n1181 vdd.n1175 52.4337
R18438 vdd.n2211 vdd.n2210 52.4337
R18439 vdd.n1174 vdd.n1169 52.4337
R18440 vdd.n2218 vdd.n2217 52.4337
R18441 vdd.n1168 vdd.n1167 52.4337
R18442 vdd.n1163 vdd.n1156 52.4337
R18443 vdd.n2229 vdd.n2228 52.4337
R18444 vdd.n1155 vdd.n1149 52.4337
R18445 vdd.n2236 vdd.n2235 52.4337
R18446 vdd.n1148 vdd.n1142 52.4337
R18447 vdd.n2243 vdd.n2242 52.4337
R18448 vdd.n1141 vdd.n1135 52.4337
R18449 vdd.n2250 vdd.n2249 52.4337
R18450 vdd.n1134 vdd.n1129 52.4337
R18451 vdd.n2257 vdd.n2256 52.4337
R18452 vdd.n1128 vdd.n1127 52.4337
R18453 vdd.n1123 vdd.n1116 52.4337
R18454 vdd.n2268 vdd.n2267 52.4337
R18455 vdd.n1115 vdd.n1109 52.4337
R18456 vdd.n2275 vdd.n2274 52.4337
R18457 vdd.n1108 vdd.n1102 52.4337
R18458 vdd.n2282 vdd.n2281 52.4337
R18459 vdd.n1101 vdd.n1098 52.4337
R18460 vdd.n2289 vdd.n2288 52.4337
R18461 vdd.n2294 vdd.n2293 52.4337
R18462 vdd.n1409 vdd.n1097 52.4337
R18463 vdd.n3230 vdd.n3229 52.4337
R18464 vdd.n3224 vdd.n663 52.4337
R18465 vdd.n3220 vdd.n666 52.4337
R18466 vdd.n3218 vdd.n3217 52.4337
R18467 vdd.n3213 vdd.n3212 52.4337
R18468 vdd.n3210 vdd.n3209 52.4337
R18469 vdd.n3205 vdd.n3204 52.4337
R18470 vdd.n3202 vdd.n3201 52.4337
R18471 vdd.n3197 vdd.n3196 52.4337
R18472 vdd.n3194 vdd.n3193 52.4337
R18473 vdd.n3189 vdd.n3188 52.4337
R18474 vdd.n3186 vdd.n3185 52.4337
R18475 vdd.n3181 vdd.n3180 52.4337
R18476 vdd.n3178 vdd.n3177 52.4337
R18477 vdd.n3173 vdd.n3172 52.4337
R18478 vdd.n3170 vdd.n3169 52.4337
R18479 vdd.n3165 vdd.n3164 52.4337
R18480 vdd.n3162 vdd.n3161 52.4337
R18481 vdd.n3157 vdd.n3156 52.4337
R18482 vdd.n3154 vdd.n3153 52.4337
R18483 vdd.n728 vdd.n727 52.4337
R18484 vdd.n3145 vdd.n3144 52.4337
R18485 vdd.n3140 vdd.n729 52.4337
R18486 vdd.n3138 vdd.n3137 52.4337
R18487 vdd.n3133 vdd.n3132 52.4337
R18488 vdd.n3130 vdd.n3129 52.4337
R18489 vdd.n3125 vdd.n3124 52.4337
R18490 vdd.n3122 vdd.n3121 52.4337
R18491 vdd.n3117 vdd.n3116 52.4337
R18492 vdd.n3112 vdd.n750 52.4337
R18493 vdd.n3108 vdd.n752 52.4337
R18494 vdd.n3344 vdd.n404 52.4337
R18495 vdd.n595 vdd.n403 52.4337
R18496 vdd.n589 vdd.n402 52.4337
R18497 vdd.n585 vdd.n401 52.4337
R18498 vdd.n579 vdd.n400 52.4337
R18499 vdd.n575 vdd.n399 52.4337
R18500 vdd.n569 vdd.n398 52.4337
R18501 vdd.n565 vdd.n397 52.4337
R18502 vdd.n559 vdd.n396 52.4337
R18503 vdd.n555 vdd.n395 52.4337
R18504 vdd.n549 vdd.n394 52.4337
R18505 vdd.n545 vdd.n393 52.4337
R18506 vdd.n539 vdd.n392 52.4337
R18507 vdd.n535 vdd.n391 52.4337
R18508 vdd.n529 vdd.n390 52.4337
R18509 vdd.n525 vdd.n389 52.4337
R18510 vdd.n519 vdd.n388 52.4337
R18511 vdd.n515 vdd.n387 52.4337
R18512 vdd.n509 vdd.n386 52.4337
R18513 vdd.n505 vdd.n385 52.4337
R18514 vdd.n499 vdd.n384 52.4337
R18515 vdd.n495 vdd.n383 52.4337
R18516 vdd.n489 vdd.n382 52.4337
R18517 vdd.n485 vdd.n381 52.4337
R18518 vdd.n479 vdd.n380 52.4337
R18519 vdd.n475 vdd.n379 52.4337
R18520 vdd.n469 vdd.n378 52.4337
R18521 vdd.n465 vdd.n377 52.4337
R18522 vdd.n459 vdd.n376 52.4337
R18523 vdd.n455 vdd.n375 52.4337
R18524 vdd.n449 vdd.n374 52.4337
R18525 vdd.n445 vdd.n373 52.4337
R18526 vdd.t266 vdd.t132 51.4683
R18527 vdd.n266 vdd.n264 42.0461
R18528 vdd.n168 vdd.n166 42.0461
R18529 vdd.n71 vdd.n69 42.0461
R18530 vdd.n2052 vdd.n2050 42.0461
R18531 vdd.n1954 vdd.n1952 42.0461
R18532 vdd.n1857 vdd.n1855 42.0461
R18533 vdd.n320 vdd.n319 41.6884
R18534 vdd.n222 vdd.n221 41.6884
R18535 vdd.n125 vdd.n124 41.6884
R18536 vdd.n2106 vdd.n2105 41.6884
R18537 vdd.n2008 vdd.n2007 41.6884
R18538 vdd.n1911 vdd.n1910 41.6884
R18539 vdd.n1512 vdd.n1511 41.1157
R18540 vdd.n1668 vdd.n1667 41.1157
R18541 vdd.n1704 vdd.n1703 41.1157
R18542 vdd.n407 vdd.n406 41.1157
R18543 vdd.n547 vdd.n420 41.1157
R18544 vdd.n433 vdd.n432 41.1157
R18545 vdd.n3062 vdd.n3061 39.2114
R18546 vdd.n3059 vdd.n3058 39.2114
R18547 vdd.n3054 vdd.n784 39.2114
R18548 vdd.n3052 vdd.n3051 39.2114
R18549 vdd.n3047 vdd.n787 39.2114
R18550 vdd.n3045 vdd.n3044 39.2114
R18551 vdd.n3040 vdd.n790 39.2114
R18552 vdd.n3038 vdd.n3037 39.2114
R18553 vdd.n3032 vdd.n793 39.2114
R18554 vdd.n3030 vdd.n3029 39.2114
R18555 vdd.n3025 vdd.n796 39.2114
R18556 vdd.n3023 vdd.n3022 39.2114
R18557 vdd.n3018 vdd.n799 39.2114
R18558 vdd.n3016 vdd.n3015 39.2114
R18559 vdd.n3011 vdd.n802 39.2114
R18560 vdd.n3009 vdd.n3008 39.2114
R18561 vdd.n3004 vdd.n3003 39.2114
R18562 vdd.n2854 vdd.n2853 39.2114
R18563 vdd.n2848 vdd.n2583 39.2114
R18564 vdd.n2845 vdd.n2584 39.2114
R18565 vdd.n2841 vdd.n2585 39.2114
R18566 vdd.n2837 vdd.n2586 39.2114
R18567 vdd.n2833 vdd.n2587 39.2114
R18568 vdd.n2829 vdd.n2588 39.2114
R18569 vdd.n2825 vdd.n2589 39.2114
R18570 vdd.n2821 vdd.n2590 39.2114
R18571 vdd.n2817 vdd.n2591 39.2114
R18572 vdd.n2813 vdd.n2592 39.2114
R18573 vdd.n2809 vdd.n2593 39.2114
R18574 vdd.n2805 vdd.n2594 39.2114
R18575 vdd.n2801 vdd.n2595 39.2114
R18576 vdd.n2797 vdd.n2596 39.2114
R18577 vdd.n2793 vdd.n2597 39.2114
R18578 vdd.n2788 vdd.n2598 39.2114
R18579 vdd.n2577 vdd.n939 39.2114
R18580 vdd.n2573 vdd.n938 39.2114
R18581 vdd.n2569 vdd.n937 39.2114
R18582 vdd.n2565 vdd.n936 39.2114
R18583 vdd.n2561 vdd.n935 39.2114
R18584 vdd.n2557 vdd.n934 39.2114
R18585 vdd.n2553 vdd.n933 39.2114
R18586 vdd.n2549 vdd.n932 39.2114
R18587 vdd.n2545 vdd.n931 39.2114
R18588 vdd.n2541 vdd.n930 39.2114
R18589 vdd.n2537 vdd.n929 39.2114
R18590 vdd.n2533 vdd.n928 39.2114
R18591 vdd.n2529 vdd.n927 39.2114
R18592 vdd.n2525 vdd.n926 39.2114
R18593 vdd.n2521 vdd.n925 39.2114
R18594 vdd.n2516 vdd.n924 39.2114
R18595 vdd.n2512 vdd.n923 39.2114
R18596 vdd.n2333 vdd.n2332 39.2114
R18597 vdd.n2327 vdd.n1055 39.2114
R18598 vdd.n2324 vdd.n1056 39.2114
R18599 vdd.n2320 vdd.n1057 39.2114
R18600 vdd.n2316 vdd.n1058 39.2114
R18601 vdd.n2312 vdd.n1059 39.2114
R18602 vdd.n2308 vdd.n1060 39.2114
R18603 vdd.n2304 vdd.n1061 39.2114
R18604 vdd.n2300 vdd.n1062 39.2114
R18605 vdd.n1247 vdd.n1063 39.2114
R18606 vdd.n1251 vdd.n1064 39.2114
R18607 vdd.n1255 vdd.n1065 39.2114
R18608 vdd.n1259 vdd.n1066 39.2114
R18609 vdd.n1263 vdd.n1067 39.2114
R18610 vdd.n1267 vdd.n1068 39.2114
R18611 vdd.n1271 vdd.n1069 39.2114
R18612 vdd.n1276 vdd.n1070 39.2114
R18613 vdd.n2981 vdd.n2980 39.2114
R18614 vdd.n2976 vdd.n2948 39.2114
R18615 vdd.n2974 vdd.n2973 39.2114
R18616 vdd.n2969 vdd.n2951 39.2114
R18617 vdd.n2967 vdd.n2966 39.2114
R18618 vdd.n2962 vdd.n2954 39.2114
R18619 vdd.n2960 vdd.n2959 39.2114
R18620 vdd.n2955 vdd.n755 39.2114
R18621 vdd.n3099 vdd.n3098 39.2114
R18622 vdd.n3096 vdd.n3095 39.2114
R18623 vdd.n3091 vdd.n760 39.2114
R18624 vdd.n3089 vdd.n3088 39.2114
R18625 vdd.n3084 vdd.n763 39.2114
R18626 vdd.n3082 vdd.n3081 39.2114
R18627 vdd.n3077 vdd.n766 39.2114
R18628 vdd.n3075 vdd.n3074 39.2114
R18629 vdd.n3070 vdd.n772 39.2114
R18630 vdd.n2857 vdd.n2856 39.2114
R18631 vdd.n2624 vdd.n2599 39.2114
R18632 vdd.n2628 vdd.n2600 39.2114
R18633 vdd.n2632 vdd.n2601 39.2114
R18634 vdd.n2636 vdd.n2602 39.2114
R18635 vdd.n2640 vdd.n2603 39.2114
R18636 vdd.n2644 vdd.n2604 39.2114
R18637 vdd.n2648 vdd.n2605 39.2114
R18638 vdd.n2652 vdd.n2606 39.2114
R18639 vdd.n2656 vdd.n2607 39.2114
R18640 vdd.n2660 vdd.n2608 39.2114
R18641 vdd.n2664 vdd.n2609 39.2114
R18642 vdd.n2668 vdd.n2610 39.2114
R18643 vdd.n2672 vdd.n2611 39.2114
R18644 vdd.n2676 vdd.n2612 39.2114
R18645 vdd.n2680 vdd.n2613 39.2114
R18646 vdd.n2684 vdd.n2614 39.2114
R18647 vdd.n2856 vdd.n904 39.2114
R18648 vdd.n2627 vdd.n2599 39.2114
R18649 vdd.n2631 vdd.n2600 39.2114
R18650 vdd.n2635 vdd.n2601 39.2114
R18651 vdd.n2639 vdd.n2602 39.2114
R18652 vdd.n2643 vdd.n2603 39.2114
R18653 vdd.n2647 vdd.n2604 39.2114
R18654 vdd.n2651 vdd.n2605 39.2114
R18655 vdd.n2655 vdd.n2606 39.2114
R18656 vdd.n2659 vdd.n2607 39.2114
R18657 vdd.n2663 vdd.n2608 39.2114
R18658 vdd.n2667 vdd.n2609 39.2114
R18659 vdd.n2671 vdd.n2610 39.2114
R18660 vdd.n2675 vdd.n2611 39.2114
R18661 vdd.n2679 vdd.n2612 39.2114
R18662 vdd.n2683 vdd.n2613 39.2114
R18663 vdd.n2686 vdd.n2614 39.2114
R18664 vdd.n772 vdd.n767 39.2114
R18665 vdd.n3076 vdd.n3075 39.2114
R18666 vdd.n766 vdd.n764 39.2114
R18667 vdd.n3083 vdd.n3082 39.2114
R18668 vdd.n763 vdd.n761 39.2114
R18669 vdd.n3090 vdd.n3089 39.2114
R18670 vdd.n760 vdd.n758 39.2114
R18671 vdd.n3097 vdd.n3096 39.2114
R18672 vdd.n3100 vdd.n3099 39.2114
R18673 vdd.n2956 vdd.n2955 39.2114
R18674 vdd.n2961 vdd.n2960 39.2114
R18675 vdd.n2954 vdd.n2952 39.2114
R18676 vdd.n2968 vdd.n2967 39.2114
R18677 vdd.n2951 vdd.n2949 39.2114
R18678 vdd.n2975 vdd.n2974 39.2114
R18679 vdd.n2948 vdd.n2946 39.2114
R18680 vdd.n2982 vdd.n2981 39.2114
R18681 vdd.n2333 vdd.n1089 39.2114
R18682 vdd.n2325 vdd.n1055 39.2114
R18683 vdd.n2321 vdd.n1056 39.2114
R18684 vdd.n2317 vdd.n1057 39.2114
R18685 vdd.n2313 vdd.n1058 39.2114
R18686 vdd.n2309 vdd.n1059 39.2114
R18687 vdd.n2305 vdd.n1060 39.2114
R18688 vdd.n2301 vdd.n1061 39.2114
R18689 vdd.n1246 vdd.n1062 39.2114
R18690 vdd.n1250 vdd.n1063 39.2114
R18691 vdd.n1254 vdd.n1064 39.2114
R18692 vdd.n1258 vdd.n1065 39.2114
R18693 vdd.n1262 vdd.n1066 39.2114
R18694 vdd.n1266 vdd.n1067 39.2114
R18695 vdd.n1270 vdd.n1068 39.2114
R18696 vdd.n1275 vdd.n1069 39.2114
R18697 vdd.n1279 vdd.n1070 39.2114
R18698 vdd.n2515 vdd.n923 39.2114
R18699 vdd.n2520 vdd.n924 39.2114
R18700 vdd.n2524 vdd.n925 39.2114
R18701 vdd.n2528 vdd.n926 39.2114
R18702 vdd.n2532 vdd.n927 39.2114
R18703 vdd.n2536 vdd.n928 39.2114
R18704 vdd.n2540 vdd.n929 39.2114
R18705 vdd.n2544 vdd.n930 39.2114
R18706 vdd.n2548 vdd.n931 39.2114
R18707 vdd.n2552 vdd.n932 39.2114
R18708 vdd.n2556 vdd.n933 39.2114
R18709 vdd.n2560 vdd.n934 39.2114
R18710 vdd.n2564 vdd.n935 39.2114
R18711 vdd.n2568 vdd.n936 39.2114
R18712 vdd.n2572 vdd.n937 39.2114
R18713 vdd.n2576 vdd.n938 39.2114
R18714 vdd.n941 vdd.n939 39.2114
R18715 vdd.n2854 vdd.n2617 39.2114
R18716 vdd.n2846 vdd.n2583 39.2114
R18717 vdd.n2842 vdd.n2584 39.2114
R18718 vdd.n2838 vdd.n2585 39.2114
R18719 vdd.n2834 vdd.n2586 39.2114
R18720 vdd.n2830 vdd.n2587 39.2114
R18721 vdd.n2826 vdd.n2588 39.2114
R18722 vdd.n2822 vdd.n2589 39.2114
R18723 vdd.n2818 vdd.n2590 39.2114
R18724 vdd.n2814 vdd.n2591 39.2114
R18725 vdd.n2810 vdd.n2592 39.2114
R18726 vdd.n2806 vdd.n2593 39.2114
R18727 vdd.n2802 vdd.n2594 39.2114
R18728 vdd.n2798 vdd.n2595 39.2114
R18729 vdd.n2794 vdd.n2596 39.2114
R18730 vdd.n2789 vdd.n2597 39.2114
R18731 vdd.n2785 vdd.n2598 39.2114
R18732 vdd.n3003 vdd.n803 39.2114
R18733 vdd.n3010 vdd.n3009 39.2114
R18734 vdd.n802 vdd.n800 39.2114
R18735 vdd.n3017 vdd.n3016 39.2114
R18736 vdd.n799 vdd.n797 39.2114
R18737 vdd.n3024 vdd.n3023 39.2114
R18738 vdd.n796 vdd.n794 39.2114
R18739 vdd.n3031 vdd.n3030 39.2114
R18740 vdd.n793 vdd.n791 39.2114
R18741 vdd.n3039 vdd.n3038 39.2114
R18742 vdd.n790 vdd.n788 39.2114
R18743 vdd.n3046 vdd.n3045 39.2114
R18744 vdd.n787 vdd.n785 39.2114
R18745 vdd.n3053 vdd.n3052 39.2114
R18746 vdd.n784 vdd.n782 39.2114
R18747 vdd.n3060 vdd.n3059 39.2114
R18748 vdd.n3063 vdd.n3062 39.2114
R18749 vdd.n950 vdd.n905 39.2114
R18750 vdd.n2504 vdd.n906 39.2114
R18751 vdd.n2500 vdd.n907 39.2114
R18752 vdd.n2496 vdd.n908 39.2114
R18753 vdd.n2492 vdd.n909 39.2114
R18754 vdd.n2488 vdd.n910 39.2114
R18755 vdd.n2484 vdd.n911 39.2114
R18756 vdd.n2480 vdd.n912 39.2114
R18757 vdd.n2476 vdd.n913 39.2114
R18758 vdd.n2472 vdd.n914 39.2114
R18759 vdd.n2468 vdd.n915 39.2114
R18760 vdd.n2464 vdd.n916 39.2114
R18761 vdd.n2460 vdd.n917 39.2114
R18762 vdd.n2456 vdd.n918 39.2114
R18763 vdd.n2452 vdd.n919 39.2114
R18764 vdd.n2448 vdd.n920 39.2114
R18765 vdd.n2444 vdd.n921 39.2114
R18766 vdd.n2336 vdd.n2335 39.2114
R18767 vdd.n1193 vdd.n1071 39.2114
R18768 vdd.n1197 vdd.n1072 39.2114
R18769 vdd.n1201 vdd.n1073 39.2114
R18770 vdd.n1205 vdd.n1074 39.2114
R18771 vdd.n1209 vdd.n1075 39.2114
R18772 vdd.n1213 vdd.n1076 39.2114
R18773 vdd.n1217 vdd.n1077 39.2114
R18774 vdd.n1221 vdd.n1078 39.2114
R18775 vdd.n1391 vdd.n1079 39.2114
R18776 vdd.n1388 vdd.n1080 39.2114
R18777 vdd.n1384 vdd.n1081 39.2114
R18778 vdd.n1380 vdd.n1082 39.2114
R18779 vdd.n1376 vdd.n1083 39.2114
R18780 vdd.n1372 vdd.n1084 39.2114
R18781 vdd.n1368 vdd.n1085 39.2114
R18782 vdd.n1364 vdd.n1086 39.2114
R18783 vdd.n2441 vdd.n921 39.2114
R18784 vdd.n2445 vdd.n920 39.2114
R18785 vdd.n2449 vdd.n919 39.2114
R18786 vdd.n2453 vdd.n918 39.2114
R18787 vdd.n2457 vdd.n917 39.2114
R18788 vdd.n2461 vdd.n916 39.2114
R18789 vdd.n2465 vdd.n915 39.2114
R18790 vdd.n2469 vdd.n914 39.2114
R18791 vdd.n2473 vdd.n913 39.2114
R18792 vdd.n2477 vdd.n912 39.2114
R18793 vdd.n2481 vdd.n911 39.2114
R18794 vdd.n2485 vdd.n910 39.2114
R18795 vdd.n2489 vdd.n909 39.2114
R18796 vdd.n2493 vdd.n908 39.2114
R18797 vdd.n2497 vdd.n907 39.2114
R18798 vdd.n2501 vdd.n906 39.2114
R18799 vdd.n2505 vdd.n905 39.2114
R18800 vdd.n2335 vdd.n1053 39.2114
R18801 vdd.n1196 vdd.n1071 39.2114
R18802 vdd.n1200 vdd.n1072 39.2114
R18803 vdd.n1204 vdd.n1073 39.2114
R18804 vdd.n1208 vdd.n1074 39.2114
R18805 vdd.n1212 vdd.n1075 39.2114
R18806 vdd.n1216 vdd.n1076 39.2114
R18807 vdd.n1220 vdd.n1077 39.2114
R18808 vdd.n1223 vdd.n1078 39.2114
R18809 vdd.n1389 vdd.n1079 39.2114
R18810 vdd.n1385 vdd.n1080 39.2114
R18811 vdd.n1381 vdd.n1081 39.2114
R18812 vdd.n1377 vdd.n1082 39.2114
R18813 vdd.n1373 vdd.n1083 39.2114
R18814 vdd.n1369 vdd.n1084 39.2114
R18815 vdd.n1365 vdd.n1085 39.2114
R18816 vdd.n1361 vdd.n1086 39.2114
R18817 vdd.n2188 vdd.n2187 37.2369
R18818 vdd.n2224 vdd.n1162 37.2369
R18819 vdd.n2263 vdd.n1122 37.2369
R18820 vdd.n3151 vdd.n724 37.2369
R18821 vdd.n688 vdd.n687 37.2369
R18822 vdd.n3107 vdd.n3106 37.2369
R18823 vdd.n2331 vdd.n1045 31.0639
R18824 vdd.n2580 vdd.n942 31.0639
R18825 vdd.n2513 vdd.n945 31.0639
R18826 vdd.n1281 vdd.n1278 31.0639
R18827 vdd.n2786 vdd.n2783 31.0639
R18828 vdd.n3005 vdd.n3002 31.0639
R18829 vdd.n2852 vdd.n897 31.0639
R18830 vdd.n3066 vdd.n3065 31.0639
R18831 vdd.n2985 vdd.n2984 31.0639
R18832 vdd.n3071 vdd.n771 31.0639
R18833 vdd.n2690 vdd.n2688 31.0639
R18834 vdd.n2859 vdd.n2858 31.0639
R18835 vdd.n2338 vdd.n2337 31.0639
R18836 vdd.n2508 vdd.n2507 31.0639
R18837 vdd.n2440 vdd.n2439 31.0639
R18838 vdd.n1360 vdd.n1359 31.0639
R18839 vdd.n1226 vdd.n1225 30.449
R18840 vdd.n954 vdd.n953 30.449
R18841 vdd.n1273 vdd.n1245 30.449
R18842 vdd.n2518 vdd.n944 30.449
R18843 vdd.n2623 vdd.n2622 30.449
R18844 vdd.n806 vdd.n805 30.449
R18845 vdd.n2791 vdd.n2619 30.449
R18846 vdd.n770 vdd.n769 30.449
R18847 vdd.n1742 vdd.n1508 19.3944
R18848 vdd.n1742 vdd.n1498 19.3944
R18849 vdd.n1754 vdd.n1498 19.3944
R18850 vdd.n1754 vdd.n1496 19.3944
R18851 vdd.n1758 vdd.n1496 19.3944
R18852 vdd.n1758 vdd.n1486 19.3944
R18853 vdd.n1771 vdd.n1486 19.3944
R18854 vdd.n1771 vdd.n1484 19.3944
R18855 vdd.n1775 vdd.n1484 19.3944
R18856 vdd.n1775 vdd.n1476 19.3944
R18857 vdd.n1788 vdd.n1476 19.3944
R18858 vdd.n1788 vdd.n1474 19.3944
R18859 vdd.n1792 vdd.n1474 19.3944
R18860 vdd.n1792 vdd.n1463 19.3944
R18861 vdd.n1804 vdd.n1463 19.3944
R18862 vdd.n1804 vdd.n1461 19.3944
R18863 vdd.n1808 vdd.n1461 19.3944
R18864 vdd.n1808 vdd.n1452 19.3944
R18865 vdd.n2116 vdd.n1452 19.3944
R18866 vdd.n2116 vdd.n1450 19.3944
R18867 vdd.n2120 vdd.n1450 19.3944
R18868 vdd.n2120 vdd.n1441 19.3944
R18869 vdd.n2132 vdd.n1441 19.3944
R18870 vdd.n2132 vdd.n1439 19.3944
R18871 vdd.n2136 vdd.n1439 19.3944
R18872 vdd.n2136 vdd.n1429 19.3944
R18873 vdd.n2149 vdd.n1429 19.3944
R18874 vdd.n2149 vdd.n1427 19.3944
R18875 vdd.n2153 vdd.n1427 19.3944
R18876 vdd.n2153 vdd.n1419 19.3944
R18877 vdd.n2166 vdd.n1419 19.3944
R18878 vdd.n2166 vdd.n1416 19.3944
R18879 vdd.n2172 vdd.n1416 19.3944
R18880 vdd.n2172 vdd.n1417 19.3944
R18881 vdd.n1417 vdd.n1406 19.3944
R18882 vdd.n1661 vdd.n1603 19.3944
R18883 vdd.n1661 vdd.n1660 19.3944
R18884 vdd.n1660 vdd.n1659 19.3944
R18885 vdd.n1659 vdd.n1609 19.3944
R18886 vdd.n1655 vdd.n1609 19.3944
R18887 vdd.n1655 vdd.n1654 19.3944
R18888 vdd.n1654 vdd.n1653 19.3944
R18889 vdd.n1653 vdd.n1615 19.3944
R18890 vdd.n1649 vdd.n1615 19.3944
R18891 vdd.n1649 vdd.n1648 19.3944
R18892 vdd.n1648 vdd.n1647 19.3944
R18893 vdd.n1647 vdd.n1621 19.3944
R18894 vdd.n1643 vdd.n1621 19.3944
R18895 vdd.n1643 vdd.n1642 19.3944
R18896 vdd.n1642 vdd.n1641 19.3944
R18897 vdd.n1641 vdd.n1627 19.3944
R18898 vdd.n1637 vdd.n1627 19.3944
R18899 vdd.n1637 vdd.n1636 19.3944
R18900 vdd.n1636 vdd.n1635 19.3944
R18901 vdd.n1635 vdd.n1633 19.3944
R18902 vdd.n1699 vdd.n1698 19.3944
R18903 vdd.n1698 vdd.n1574 19.3944
R18904 vdd.n1694 vdd.n1574 19.3944
R18905 vdd.n1694 vdd.n1693 19.3944
R18906 vdd.n1693 vdd.n1692 19.3944
R18907 vdd.n1692 vdd.n1580 19.3944
R18908 vdd.n1688 vdd.n1580 19.3944
R18909 vdd.n1688 vdd.n1687 19.3944
R18910 vdd.n1687 vdd.n1686 19.3944
R18911 vdd.n1686 vdd.n1586 19.3944
R18912 vdd.n1682 vdd.n1586 19.3944
R18913 vdd.n1682 vdd.n1681 19.3944
R18914 vdd.n1681 vdd.n1680 19.3944
R18915 vdd.n1680 vdd.n1592 19.3944
R18916 vdd.n1676 vdd.n1592 19.3944
R18917 vdd.n1676 vdd.n1675 19.3944
R18918 vdd.n1675 vdd.n1674 19.3944
R18919 vdd.n1674 vdd.n1598 19.3944
R18920 vdd.n1670 vdd.n1598 19.3944
R18921 vdd.n1670 vdd.n1669 19.3944
R18922 vdd.n1733 vdd.n1732 19.3944
R18923 vdd.n1732 vdd.n1547 19.3944
R18924 vdd.n1728 vdd.n1547 19.3944
R18925 vdd.n1728 vdd.n1727 19.3944
R18926 vdd.n1727 vdd.n1726 19.3944
R18927 vdd.n1726 vdd.n1552 19.3944
R18928 vdd.n1722 vdd.n1552 19.3944
R18929 vdd.n1722 vdd.n1721 19.3944
R18930 vdd.n1721 vdd.n1720 19.3944
R18931 vdd.n1720 vdd.n1558 19.3944
R18932 vdd.n1716 vdd.n1558 19.3944
R18933 vdd.n1716 vdd.n1715 19.3944
R18934 vdd.n1715 vdd.n1714 19.3944
R18935 vdd.n1714 vdd.n1564 19.3944
R18936 vdd.n1710 vdd.n1564 19.3944
R18937 vdd.n1710 vdd.n1709 19.3944
R18938 vdd.n1709 vdd.n1708 19.3944
R18939 vdd.n1708 vdd.n1570 19.3944
R18940 vdd.n2220 vdd.n1160 19.3944
R18941 vdd.n2220 vdd.n1166 19.3944
R18942 vdd.n2215 vdd.n1166 19.3944
R18943 vdd.n2215 vdd.n2214 19.3944
R18944 vdd.n2214 vdd.n2213 19.3944
R18945 vdd.n2213 vdd.n1173 19.3944
R18946 vdd.n2208 vdd.n1173 19.3944
R18947 vdd.n2208 vdd.n2207 19.3944
R18948 vdd.n2207 vdd.n2206 19.3944
R18949 vdd.n2206 vdd.n1180 19.3944
R18950 vdd.n2201 vdd.n1180 19.3944
R18951 vdd.n2201 vdd.n2200 19.3944
R18952 vdd.n2200 vdd.n2199 19.3944
R18953 vdd.n2199 vdd.n1187 19.3944
R18954 vdd.n2194 vdd.n1187 19.3944
R18955 vdd.n2194 vdd.n2193 19.3944
R18956 vdd.n1399 vdd.n1192 19.3944
R18957 vdd.n2189 vdd.n1396 19.3944
R18958 vdd.n2259 vdd.n1120 19.3944
R18959 vdd.n2259 vdd.n1126 19.3944
R18960 vdd.n2254 vdd.n1126 19.3944
R18961 vdd.n2254 vdd.n2253 19.3944
R18962 vdd.n2253 vdd.n2252 19.3944
R18963 vdd.n2252 vdd.n1133 19.3944
R18964 vdd.n2247 vdd.n1133 19.3944
R18965 vdd.n2247 vdd.n2246 19.3944
R18966 vdd.n2246 vdd.n2245 19.3944
R18967 vdd.n2245 vdd.n1140 19.3944
R18968 vdd.n2240 vdd.n1140 19.3944
R18969 vdd.n2240 vdd.n2239 19.3944
R18970 vdd.n2239 vdd.n2238 19.3944
R18971 vdd.n2238 vdd.n1147 19.3944
R18972 vdd.n2233 vdd.n1147 19.3944
R18973 vdd.n2233 vdd.n2232 19.3944
R18974 vdd.n2232 vdd.n2231 19.3944
R18975 vdd.n2231 vdd.n1154 19.3944
R18976 vdd.n2226 vdd.n1154 19.3944
R18977 vdd.n2226 vdd.n2225 19.3944
R18978 vdd.n2296 vdd.n1095 19.3944
R18979 vdd.n2296 vdd.n1096 19.3944
R18980 vdd.n2291 vdd.n2290 19.3944
R18981 vdd.n2286 vdd.n2285 19.3944
R18982 vdd.n2285 vdd.n2284 19.3944
R18983 vdd.n2284 vdd.n1100 19.3944
R18984 vdd.n2279 vdd.n1100 19.3944
R18985 vdd.n2279 vdd.n2278 19.3944
R18986 vdd.n2278 vdd.n2277 19.3944
R18987 vdd.n2277 vdd.n1107 19.3944
R18988 vdd.n2272 vdd.n1107 19.3944
R18989 vdd.n2272 vdd.n2271 19.3944
R18990 vdd.n2271 vdd.n2270 19.3944
R18991 vdd.n2270 vdd.n1114 19.3944
R18992 vdd.n2265 vdd.n1114 19.3944
R18993 vdd.n2265 vdd.n2264 19.3944
R18994 vdd.n1746 vdd.n1504 19.3944
R18995 vdd.n1746 vdd.n1502 19.3944
R18996 vdd.n1750 vdd.n1502 19.3944
R18997 vdd.n1750 vdd.n1492 19.3944
R18998 vdd.n1763 vdd.n1492 19.3944
R18999 vdd.n1763 vdd.n1490 19.3944
R19000 vdd.n1767 vdd.n1490 19.3944
R19001 vdd.n1767 vdd.n1481 19.3944
R19002 vdd.n1780 vdd.n1481 19.3944
R19003 vdd.n1780 vdd.n1479 19.3944
R19004 vdd.n1784 vdd.n1479 19.3944
R19005 vdd.n1784 vdd.n1470 19.3944
R19006 vdd.n1796 vdd.n1470 19.3944
R19007 vdd.n1796 vdd.n1468 19.3944
R19008 vdd.n1800 vdd.n1468 19.3944
R19009 vdd.n1800 vdd.n1458 19.3944
R19010 vdd.n1813 vdd.n1458 19.3944
R19011 vdd.n1813 vdd.n1456 19.3944
R19012 vdd.n2112 vdd.n1456 19.3944
R19013 vdd.n2112 vdd.n1447 19.3944
R19014 vdd.n2124 vdd.n1447 19.3944
R19015 vdd.n2124 vdd.n1445 19.3944
R19016 vdd.n2128 vdd.n1445 19.3944
R19017 vdd.n2128 vdd.n1435 19.3944
R19018 vdd.n2141 vdd.n1435 19.3944
R19019 vdd.n2141 vdd.n1433 19.3944
R19020 vdd.n2145 vdd.n1433 19.3944
R19021 vdd.n2145 vdd.n1424 19.3944
R19022 vdd.n2158 vdd.n1424 19.3944
R19023 vdd.n2158 vdd.n1422 19.3944
R19024 vdd.n2162 vdd.n1422 19.3944
R19025 vdd.n2162 vdd.n1412 19.3944
R19026 vdd.n2176 vdd.n1412 19.3944
R19027 vdd.n2176 vdd.n1410 19.3944
R19028 vdd.n2180 vdd.n1410 19.3944
R19029 vdd.n3239 vdd.n655 19.3944
R19030 vdd.n3243 vdd.n655 19.3944
R19031 vdd.n3243 vdd.n646 19.3944
R19032 vdd.n3255 vdd.n646 19.3944
R19033 vdd.n3255 vdd.n644 19.3944
R19034 vdd.n3259 vdd.n644 19.3944
R19035 vdd.n3259 vdd.n633 19.3944
R19036 vdd.n3271 vdd.n633 19.3944
R19037 vdd.n3271 vdd.n631 19.3944
R19038 vdd.n3275 vdd.n631 19.3944
R19039 vdd.n3275 vdd.n622 19.3944
R19040 vdd.n3288 vdd.n622 19.3944
R19041 vdd.n3288 vdd.n620 19.3944
R19042 vdd.n3295 vdd.n620 19.3944
R19043 vdd.n3295 vdd.n3294 19.3944
R19044 vdd.n3294 vdd.n610 19.3944
R19045 vdd.n3308 vdd.n610 19.3944
R19046 vdd.n3309 vdd.n3308 19.3944
R19047 vdd.n3310 vdd.n3309 19.3944
R19048 vdd.n3310 vdd.n608 19.3944
R19049 vdd.n3315 vdd.n608 19.3944
R19050 vdd.n3316 vdd.n3315 19.3944
R19051 vdd.n3317 vdd.n3316 19.3944
R19052 vdd.n3317 vdd.n606 19.3944
R19053 vdd.n3322 vdd.n606 19.3944
R19054 vdd.n3323 vdd.n3322 19.3944
R19055 vdd.n3324 vdd.n3323 19.3944
R19056 vdd.n3324 vdd.n604 19.3944
R19057 vdd.n3330 vdd.n604 19.3944
R19058 vdd.n3331 vdd.n3330 19.3944
R19059 vdd.n3332 vdd.n3331 19.3944
R19060 vdd.n3332 vdd.n602 19.3944
R19061 vdd.n3337 vdd.n602 19.3944
R19062 vdd.n3338 vdd.n3337 19.3944
R19063 vdd.n3339 vdd.n3338 19.3944
R19064 vdd.n550 vdd.n417 19.3944
R19065 vdd.n556 vdd.n417 19.3944
R19066 vdd.n557 vdd.n556 19.3944
R19067 vdd.n560 vdd.n557 19.3944
R19068 vdd.n560 vdd.n415 19.3944
R19069 vdd.n566 vdd.n415 19.3944
R19070 vdd.n567 vdd.n566 19.3944
R19071 vdd.n570 vdd.n567 19.3944
R19072 vdd.n570 vdd.n413 19.3944
R19073 vdd.n576 vdd.n413 19.3944
R19074 vdd.n577 vdd.n576 19.3944
R19075 vdd.n580 vdd.n577 19.3944
R19076 vdd.n580 vdd.n411 19.3944
R19077 vdd.n586 vdd.n411 19.3944
R19078 vdd.n587 vdd.n586 19.3944
R19079 vdd.n590 vdd.n587 19.3944
R19080 vdd.n590 vdd.n409 19.3944
R19081 vdd.n596 vdd.n409 19.3944
R19082 vdd.n598 vdd.n596 19.3944
R19083 vdd.n599 vdd.n598 19.3944
R19084 vdd.n497 vdd.n496 19.3944
R19085 vdd.n500 vdd.n497 19.3944
R19086 vdd.n500 vdd.n429 19.3944
R19087 vdd.n506 vdd.n429 19.3944
R19088 vdd.n507 vdd.n506 19.3944
R19089 vdd.n510 vdd.n507 19.3944
R19090 vdd.n510 vdd.n427 19.3944
R19091 vdd.n516 vdd.n427 19.3944
R19092 vdd.n517 vdd.n516 19.3944
R19093 vdd.n520 vdd.n517 19.3944
R19094 vdd.n520 vdd.n425 19.3944
R19095 vdd.n526 vdd.n425 19.3944
R19096 vdd.n527 vdd.n526 19.3944
R19097 vdd.n530 vdd.n527 19.3944
R19098 vdd.n530 vdd.n423 19.3944
R19099 vdd.n536 vdd.n423 19.3944
R19100 vdd.n537 vdd.n536 19.3944
R19101 vdd.n540 vdd.n537 19.3944
R19102 vdd.n540 vdd.n421 19.3944
R19103 vdd.n546 vdd.n421 19.3944
R19104 vdd.n447 vdd.n446 19.3944
R19105 vdd.n450 vdd.n447 19.3944
R19106 vdd.n450 vdd.n441 19.3944
R19107 vdd.n456 vdd.n441 19.3944
R19108 vdd.n457 vdd.n456 19.3944
R19109 vdd.n460 vdd.n457 19.3944
R19110 vdd.n460 vdd.n439 19.3944
R19111 vdd.n466 vdd.n439 19.3944
R19112 vdd.n467 vdd.n466 19.3944
R19113 vdd.n470 vdd.n467 19.3944
R19114 vdd.n470 vdd.n437 19.3944
R19115 vdd.n476 vdd.n437 19.3944
R19116 vdd.n477 vdd.n476 19.3944
R19117 vdd.n480 vdd.n477 19.3944
R19118 vdd.n480 vdd.n435 19.3944
R19119 vdd.n486 vdd.n435 19.3944
R19120 vdd.n487 vdd.n486 19.3944
R19121 vdd.n490 vdd.n487 19.3944
R19122 vdd.n3235 vdd.n652 19.3944
R19123 vdd.n3247 vdd.n652 19.3944
R19124 vdd.n3247 vdd.n650 19.3944
R19125 vdd.n3251 vdd.n650 19.3944
R19126 vdd.n3251 vdd.n640 19.3944
R19127 vdd.n3263 vdd.n640 19.3944
R19128 vdd.n3263 vdd.n638 19.3944
R19129 vdd.n3267 vdd.n638 19.3944
R19130 vdd.n3267 vdd.n628 19.3944
R19131 vdd.n3280 vdd.n628 19.3944
R19132 vdd.n3280 vdd.n626 19.3944
R19133 vdd.n3284 vdd.n626 19.3944
R19134 vdd.n3284 vdd.n617 19.3944
R19135 vdd.n3299 vdd.n617 19.3944
R19136 vdd.n3299 vdd.n615 19.3944
R19137 vdd.n3303 vdd.n615 19.3944
R19138 vdd.n3303 vdd.n324 19.3944
R19139 vdd.n3381 vdd.n324 19.3944
R19140 vdd.n3381 vdd.n325 19.3944
R19141 vdd.n3375 vdd.n325 19.3944
R19142 vdd.n3375 vdd.n3374 19.3944
R19143 vdd.n3374 vdd.n3373 19.3944
R19144 vdd.n3373 vdd.n337 19.3944
R19145 vdd.n3367 vdd.n337 19.3944
R19146 vdd.n3367 vdd.n3366 19.3944
R19147 vdd.n3366 vdd.n3365 19.3944
R19148 vdd.n3365 vdd.n347 19.3944
R19149 vdd.n3359 vdd.n347 19.3944
R19150 vdd.n3359 vdd.n3358 19.3944
R19151 vdd.n3358 vdd.n3357 19.3944
R19152 vdd.n3357 vdd.n358 19.3944
R19153 vdd.n3351 vdd.n358 19.3944
R19154 vdd.n3351 vdd.n3350 19.3944
R19155 vdd.n3350 vdd.n3349 19.3944
R19156 vdd.n3349 vdd.n369 19.3944
R19157 vdd.n3192 vdd.n3191 19.3944
R19158 vdd.n3191 vdd.n3190 19.3944
R19159 vdd.n3190 vdd.n694 19.3944
R19160 vdd.n3184 vdd.n694 19.3944
R19161 vdd.n3184 vdd.n3183 19.3944
R19162 vdd.n3183 vdd.n3182 19.3944
R19163 vdd.n3182 vdd.n700 19.3944
R19164 vdd.n3176 vdd.n700 19.3944
R19165 vdd.n3176 vdd.n3175 19.3944
R19166 vdd.n3175 vdd.n3174 19.3944
R19167 vdd.n3174 vdd.n706 19.3944
R19168 vdd.n3168 vdd.n706 19.3944
R19169 vdd.n3168 vdd.n3167 19.3944
R19170 vdd.n3167 vdd.n3166 19.3944
R19171 vdd.n3166 vdd.n712 19.3944
R19172 vdd.n3160 vdd.n712 19.3944
R19173 vdd.n3160 vdd.n3159 19.3944
R19174 vdd.n3159 vdd.n3158 19.3944
R19175 vdd.n3158 vdd.n718 19.3944
R19176 vdd.n3152 vdd.n718 19.3944
R19177 vdd.n3232 vdd.n3231 19.3944
R19178 vdd.n3231 vdd.n662 19.3944
R19179 vdd.n3226 vdd.n3225 19.3944
R19180 vdd.n3222 vdd.n3221 19.3944
R19181 vdd.n3221 vdd.n668 19.3944
R19182 vdd.n3216 vdd.n668 19.3944
R19183 vdd.n3216 vdd.n3215 19.3944
R19184 vdd.n3215 vdd.n3214 19.3944
R19185 vdd.n3214 vdd.n674 19.3944
R19186 vdd.n3208 vdd.n674 19.3944
R19187 vdd.n3208 vdd.n3207 19.3944
R19188 vdd.n3207 vdd.n3206 19.3944
R19189 vdd.n3206 vdd.n680 19.3944
R19190 vdd.n3200 vdd.n680 19.3944
R19191 vdd.n3200 vdd.n3199 19.3944
R19192 vdd.n3199 vdd.n3198 19.3944
R19193 vdd.n3147 vdd.n722 19.3944
R19194 vdd.n3147 vdd.n726 19.3944
R19195 vdd.n3142 vdd.n726 19.3944
R19196 vdd.n3142 vdd.n3141 19.3944
R19197 vdd.n3141 vdd.n732 19.3944
R19198 vdd.n3136 vdd.n732 19.3944
R19199 vdd.n3136 vdd.n3135 19.3944
R19200 vdd.n3135 vdd.n3134 19.3944
R19201 vdd.n3134 vdd.n738 19.3944
R19202 vdd.n3128 vdd.n738 19.3944
R19203 vdd.n3128 vdd.n3127 19.3944
R19204 vdd.n3127 vdd.n3126 19.3944
R19205 vdd.n3126 vdd.n744 19.3944
R19206 vdd.n3120 vdd.n744 19.3944
R19207 vdd.n3120 vdd.n3119 19.3944
R19208 vdd.n3119 vdd.n3118 19.3944
R19209 vdd.n3114 vdd.n3113 19.3944
R19210 vdd.n3110 vdd.n3109 19.3944
R19211 vdd.n1668 vdd.n1603 19.0066
R19212 vdd.n2224 vdd.n1160 19.0066
R19213 vdd.n550 vdd.n547 19.0066
R19214 vdd.n3151 vdd.n722 19.0066
R19215 vdd.n1736 vdd.n1506 18.5924
R19216 vdd.n2182 vdd.n1054 18.5924
R19217 vdd.n3237 vdd.n658 18.5924
R19218 vdd.n3346 vdd.n3345 18.5924
R19219 vdd.n1225 vdd.n1224 16.0975
R19220 vdd.n953 vdd.n952 16.0975
R19221 vdd.n1511 vdd.n1510 16.0975
R19222 vdd.n1667 vdd.n1666 16.0975
R19223 vdd.n1703 vdd.n1702 16.0975
R19224 vdd.n2187 vdd.n2186 16.0975
R19225 vdd.n1162 vdd.n1161 16.0975
R19226 vdd.n1122 vdd.n1121 16.0975
R19227 vdd.n1245 vdd.n1244 16.0975
R19228 vdd.n944 vdd.n943 16.0975
R19229 vdd.n2622 vdd.n2621 16.0975
R19230 vdd.n406 vdd.n405 16.0975
R19231 vdd.n420 vdd.n419 16.0975
R19232 vdd.n432 vdd.n431 16.0975
R19233 vdd.n724 vdd.n723 16.0975
R19234 vdd.n687 vdd.n686 16.0975
R19235 vdd.n805 vdd.n804 16.0975
R19236 vdd.n2619 vdd.n2618 16.0975
R19237 vdd.n3106 vdd.n3105 16.0975
R19238 vdd.n769 vdd.n768 16.0975
R19239 vdd.t132 vdd.n2582 15.4182
R19240 vdd.n2855 vdd.t266 15.4182
R19241 vdd.n28 vdd.n27 14.7125
R19242 vdd.n2334 vdd.n1047 14.0578
R19243 vdd.n3068 vdd.n756 14.0578
R19244 vdd.n316 vdd.n281 13.1884
R19245 vdd.n261 vdd.n226 13.1884
R19246 vdd.n218 vdd.n183 13.1884
R19247 vdd.n163 vdd.n128 13.1884
R19248 vdd.n121 vdd.n86 13.1884
R19249 vdd.n66 vdd.n31 13.1884
R19250 vdd.n2047 vdd.n2012 13.1884
R19251 vdd.n2102 vdd.n2067 13.1884
R19252 vdd.n1949 vdd.n1914 13.1884
R19253 vdd.n2004 vdd.n1969 13.1884
R19254 vdd.n1852 vdd.n1817 13.1884
R19255 vdd.n1907 vdd.n1872 13.1884
R19256 vdd.n1704 vdd.n1699 12.9944
R19257 vdd.n1704 vdd.n1570 12.9944
R19258 vdd.n2263 vdd.n1120 12.9944
R19259 vdd.n2264 vdd.n2263 12.9944
R19260 vdd.n496 vdd.n433 12.9944
R19261 vdd.n490 vdd.n433 12.9944
R19262 vdd.n3192 vdd.n688 12.9944
R19263 vdd.n3198 vdd.n688 12.9944
R19264 vdd.n317 vdd.n279 12.8005
R19265 vdd.n312 vdd.n283 12.8005
R19266 vdd.n262 vdd.n224 12.8005
R19267 vdd.n257 vdd.n228 12.8005
R19268 vdd.n219 vdd.n181 12.8005
R19269 vdd.n214 vdd.n185 12.8005
R19270 vdd.n164 vdd.n126 12.8005
R19271 vdd.n159 vdd.n130 12.8005
R19272 vdd.n122 vdd.n84 12.8005
R19273 vdd.n117 vdd.n88 12.8005
R19274 vdd.n67 vdd.n29 12.8005
R19275 vdd.n62 vdd.n33 12.8005
R19276 vdd.n2048 vdd.n2010 12.8005
R19277 vdd.n2043 vdd.n2014 12.8005
R19278 vdd.n2103 vdd.n2065 12.8005
R19279 vdd.n2098 vdd.n2069 12.8005
R19280 vdd.n1950 vdd.n1912 12.8005
R19281 vdd.n1945 vdd.n1916 12.8005
R19282 vdd.n2005 vdd.n1967 12.8005
R19283 vdd.n2000 vdd.n1971 12.8005
R19284 vdd.n1853 vdd.n1815 12.8005
R19285 vdd.n1848 vdd.n1819 12.8005
R19286 vdd.n1908 vdd.n1870 12.8005
R19287 vdd.n1903 vdd.n1874 12.8005
R19288 vdd.n311 vdd.n284 12.0247
R19289 vdd.n256 vdd.n229 12.0247
R19290 vdd.n213 vdd.n186 12.0247
R19291 vdd.n158 vdd.n131 12.0247
R19292 vdd.n116 vdd.n89 12.0247
R19293 vdd.n61 vdd.n34 12.0247
R19294 vdd.n2042 vdd.n2015 12.0247
R19295 vdd.n2097 vdd.n2070 12.0247
R19296 vdd.n1944 vdd.n1917 12.0247
R19297 vdd.n1999 vdd.n1972 12.0247
R19298 vdd.n1847 vdd.n1820 12.0247
R19299 vdd.n1902 vdd.n1875 12.0247
R19300 vdd.n1744 vdd.n1506 11.337
R19301 vdd.n1752 vdd.n1500 11.337
R19302 vdd.n1752 vdd.n1494 11.337
R19303 vdd.n1761 vdd.n1494 11.337
R19304 vdd.n1769 vdd.n1488 11.337
R19305 vdd.n1778 vdd.n1777 11.337
R19306 vdd.n1794 vdd.n1472 11.337
R19307 vdd.n1802 vdd.n1465 11.337
R19308 vdd.n1811 vdd.n1810 11.337
R19309 vdd.n2114 vdd.n1454 11.337
R19310 vdd.n2130 vdd.n1443 11.337
R19311 vdd.n2139 vdd.n1437 11.337
R19312 vdd.n2147 vdd.n1431 11.337
R19313 vdd.n2156 vdd.n2155 11.337
R19314 vdd.n2164 vdd.n1414 11.337
R19315 vdd.n2174 vdd.n1414 11.337
R19316 vdd.n2182 vdd.n1407 11.337
R19317 vdd.n3237 vdd.n659 11.337
R19318 vdd.n3245 vdd.n648 11.337
R19319 vdd.n3253 vdd.n648 11.337
R19320 vdd.n3261 vdd.n642 11.337
R19321 vdd.n3269 vdd.n635 11.337
R19322 vdd.n3278 vdd.n3277 11.337
R19323 vdd.n3286 vdd.n624 11.337
R19324 vdd.n3305 vdd.n613 11.337
R19325 vdd.n3379 vdd.n328 11.337
R19326 vdd.n3377 vdd.n332 11.337
R19327 vdd.n3371 vdd.n3370 11.337
R19328 vdd.n3363 vdd.n349 11.337
R19329 vdd.n3362 vdd.n3361 11.337
R19330 vdd.n3355 vdd.n3354 11.337
R19331 vdd.n3354 vdd.n3353 11.337
R19332 vdd.n3353 vdd.n363 11.337
R19333 vdd.n3347 vdd.n3346 11.337
R19334 vdd.n308 vdd.n307 11.249
R19335 vdd.n253 vdd.n252 11.249
R19336 vdd.n210 vdd.n209 11.249
R19337 vdd.n155 vdd.n154 11.249
R19338 vdd.n113 vdd.n112 11.249
R19339 vdd.n58 vdd.n57 11.249
R19340 vdd.n2039 vdd.n2038 11.249
R19341 vdd.n2094 vdd.n2093 11.249
R19342 vdd.n1941 vdd.n1940 11.249
R19343 vdd.n1996 vdd.n1995 11.249
R19344 vdd.n1844 vdd.n1843 11.249
R19345 vdd.n1899 vdd.n1898 11.249
R19346 vdd.n2164 vdd.t172 10.7702
R19347 vdd.n3253 vdd.t177 10.7702
R19348 vdd.n293 vdd.n292 10.7238
R19349 vdd.n238 vdd.n237 10.7238
R19350 vdd.n195 vdd.n194 10.7238
R19351 vdd.n140 vdd.n139 10.7238
R19352 vdd.n98 vdd.n97 10.7238
R19353 vdd.n43 vdd.n42 10.7238
R19354 vdd.n2024 vdd.n2023 10.7238
R19355 vdd.n2079 vdd.n2078 10.7238
R19356 vdd.n1926 vdd.n1925 10.7238
R19357 vdd.n1981 vdd.n1980 10.7238
R19358 vdd.n1829 vdd.n1828 10.7238
R19359 vdd.n1884 vdd.n1883 10.7238
R19360 vdd.n2510 vdd.t19 10.6568
R19361 vdd.t38 vdd.n899 10.6568
R19362 vdd.n2343 vdd.n1045 10.6151
R19363 vdd.n2344 vdd.n2343 10.6151
R19364 vdd.n2345 vdd.n2344 10.6151
R19365 vdd.n2345 vdd.n1034 10.6151
R19366 vdd.n2355 vdd.n1034 10.6151
R19367 vdd.n2356 vdd.n2355 10.6151
R19368 vdd.n2357 vdd.n2356 10.6151
R19369 vdd.n2357 vdd.n1021 10.6151
R19370 vdd.n2367 vdd.n1021 10.6151
R19371 vdd.n2368 vdd.n2367 10.6151
R19372 vdd.n2369 vdd.n2368 10.6151
R19373 vdd.n2369 vdd.n1009 10.6151
R19374 vdd.n2380 vdd.n1009 10.6151
R19375 vdd.n2381 vdd.n2380 10.6151
R19376 vdd.n2382 vdd.n2381 10.6151
R19377 vdd.n2382 vdd.n997 10.6151
R19378 vdd.n2392 vdd.n997 10.6151
R19379 vdd.n2393 vdd.n2392 10.6151
R19380 vdd.n2394 vdd.n2393 10.6151
R19381 vdd.n2394 vdd.n985 10.6151
R19382 vdd.n2404 vdd.n985 10.6151
R19383 vdd.n2405 vdd.n2404 10.6151
R19384 vdd.n2406 vdd.n2405 10.6151
R19385 vdd.n2406 vdd.n974 10.6151
R19386 vdd.n2416 vdd.n974 10.6151
R19387 vdd.n2417 vdd.n2416 10.6151
R19388 vdd.n2418 vdd.n2417 10.6151
R19389 vdd.n2418 vdd.n961 10.6151
R19390 vdd.n2430 vdd.n961 10.6151
R19391 vdd.n2431 vdd.n2430 10.6151
R19392 vdd.n2433 vdd.n2431 10.6151
R19393 vdd.n2433 vdd.n2432 10.6151
R19394 vdd.n2432 vdd.n942 10.6151
R19395 vdd.n2580 vdd.n2579 10.6151
R19396 vdd.n2579 vdd.n2578 10.6151
R19397 vdd.n2578 vdd.n2575 10.6151
R19398 vdd.n2575 vdd.n2574 10.6151
R19399 vdd.n2574 vdd.n2571 10.6151
R19400 vdd.n2571 vdd.n2570 10.6151
R19401 vdd.n2570 vdd.n2567 10.6151
R19402 vdd.n2567 vdd.n2566 10.6151
R19403 vdd.n2566 vdd.n2563 10.6151
R19404 vdd.n2563 vdd.n2562 10.6151
R19405 vdd.n2562 vdd.n2559 10.6151
R19406 vdd.n2559 vdd.n2558 10.6151
R19407 vdd.n2558 vdd.n2555 10.6151
R19408 vdd.n2555 vdd.n2554 10.6151
R19409 vdd.n2554 vdd.n2551 10.6151
R19410 vdd.n2551 vdd.n2550 10.6151
R19411 vdd.n2550 vdd.n2547 10.6151
R19412 vdd.n2547 vdd.n2546 10.6151
R19413 vdd.n2546 vdd.n2543 10.6151
R19414 vdd.n2543 vdd.n2542 10.6151
R19415 vdd.n2542 vdd.n2539 10.6151
R19416 vdd.n2539 vdd.n2538 10.6151
R19417 vdd.n2538 vdd.n2535 10.6151
R19418 vdd.n2535 vdd.n2534 10.6151
R19419 vdd.n2534 vdd.n2531 10.6151
R19420 vdd.n2531 vdd.n2530 10.6151
R19421 vdd.n2530 vdd.n2527 10.6151
R19422 vdd.n2527 vdd.n2526 10.6151
R19423 vdd.n2526 vdd.n2523 10.6151
R19424 vdd.n2523 vdd.n2522 10.6151
R19425 vdd.n2522 vdd.n2519 10.6151
R19426 vdd.n2517 vdd.n2514 10.6151
R19427 vdd.n2514 vdd.n2513 10.6151
R19428 vdd.n1282 vdd.n1281 10.6151
R19429 vdd.n1284 vdd.n1282 10.6151
R19430 vdd.n1285 vdd.n1284 10.6151
R19431 vdd.n1287 vdd.n1285 10.6151
R19432 vdd.n1288 vdd.n1287 10.6151
R19433 vdd.n1290 vdd.n1288 10.6151
R19434 vdd.n1291 vdd.n1290 10.6151
R19435 vdd.n1293 vdd.n1291 10.6151
R19436 vdd.n1294 vdd.n1293 10.6151
R19437 vdd.n1296 vdd.n1294 10.6151
R19438 vdd.n1297 vdd.n1296 10.6151
R19439 vdd.n1299 vdd.n1297 10.6151
R19440 vdd.n1300 vdd.n1299 10.6151
R19441 vdd.n1302 vdd.n1300 10.6151
R19442 vdd.n1303 vdd.n1302 10.6151
R19443 vdd.n1305 vdd.n1303 10.6151
R19444 vdd.n1306 vdd.n1305 10.6151
R19445 vdd.n1328 vdd.n1306 10.6151
R19446 vdd.n1328 vdd.n1327 10.6151
R19447 vdd.n1327 vdd.n1326 10.6151
R19448 vdd.n1326 vdd.n1324 10.6151
R19449 vdd.n1324 vdd.n1323 10.6151
R19450 vdd.n1323 vdd.n1321 10.6151
R19451 vdd.n1321 vdd.n1320 10.6151
R19452 vdd.n1320 vdd.n1318 10.6151
R19453 vdd.n1318 vdd.n1317 10.6151
R19454 vdd.n1317 vdd.n1315 10.6151
R19455 vdd.n1315 vdd.n1314 10.6151
R19456 vdd.n1314 vdd.n1312 10.6151
R19457 vdd.n1312 vdd.n1311 10.6151
R19458 vdd.n1311 vdd.n1308 10.6151
R19459 vdd.n1308 vdd.n1307 10.6151
R19460 vdd.n1307 vdd.n945 10.6151
R19461 vdd.n2331 vdd.n2330 10.6151
R19462 vdd.n2330 vdd.n2329 10.6151
R19463 vdd.n2329 vdd.n2328 10.6151
R19464 vdd.n2328 vdd.n2326 10.6151
R19465 vdd.n2326 vdd.n2323 10.6151
R19466 vdd.n2323 vdd.n2322 10.6151
R19467 vdd.n2322 vdd.n2319 10.6151
R19468 vdd.n2319 vdd.n2318 10.6151
R19469 vdd.n2318 vdd.n2315 10.6151
R19470 vdd.n2315 vdd.n2314 10.6151
R19471 vdd.n2314 vdd.n2311 10.6151
R19472 vdd.n2311 vdd.n2310 10.6151
R19473 vdd.n2310 vdd.n2307 10.6151
R19474 vdd.n2307 vdd.n2306 10.6151
R19475 vdd.n2306 vdd.n2303 10.6151
R19476 vdd.n2303 vdd.n2302 10.6151
R19477 vdd.n2302 vdd.n2299 10.6151
R19478 vdd.n2299 vdd.n1090 10.6151
R19479 vdd.n1248 vdd.n1090 10.6151
R19480 vdd.n1249 vdd.n1248 10.6151
R19481 vdd.n1252 vdd.n1249 10.6151
R19482 vdd.n1253 vdd.n1252 10.6151
R19483 vdd.n1256 vdd.n1253 10.6151
R19484 vdd.n1257 vdd.n1256 10.6151
R19485 vdd.n1260 vdd.n1257 10.6151
R19486 vdd.n1261 vdd.n1260 10.6151
R19487 vdd.n1264 vdd.n1261 10.6151
R19488 vdd.n1265 vdd.n1264 10.6151
R19489 vdd.n1268 vdd.n1265 10.6151
R19490 vdd.n1269 vdd.n1268 10.6151
R19491 vdd.n1272 vdd.n1269 10.6151
R19492 vdd.n1277 vdd.n1274 10.6151
R19493 vdd.n1278 vdd.n1277 10.6151
R19494 vdd.n2783 vdd.n2782 10.6151
R19495 vdd.n2782 vdd.n2781 10.6151
R19496 vdd.n2781 vdd.n2620 10.6151
R19497 vdd.n2725 vdd.n2620 10.6151
R19498 vdd.n2726 vdd.n2725 10.6151
R19499 vdd.n2728 vdd.n2726 10.6151
R19500 vdd.n2729 vdd.n2728 10.6151
R19501 vdd.n2731 vdd.n2729 10.6151
R19502 vdd.n2732 vdd.n2731 10.6151
R19503 vdd.n2762 vdd.n2732 10.6151
R19504 vdd.n2762 vdd.n2761 10.6151
R19505 vdd.n2761 vdd.n2760 10.6151
R19506 vdd.n2760 vdd.n2758 10.6151
R19507 vdd.n2758 vdd.n2757 10.6151
R19508 vdd.n2757 vdd.n2755 10.6151
R19509 vdd.n2755 vdd.n2754 10.6151
R19510 vdd.n2754 vdd.n2752 10.6151
R19511 vdd.n2752 vdd.n2751 10.6151
R19512 vdd.n2751 vdd.n2749 10.6151
R19513 vdd.n2749 vdd.n2748 10.6151
R19514 vdd.n2748 vdd.n2746 10.6151
R19515 vdd.n2746 vdd.n2745 10.6151
R19516 vdd.n2745 vdd.n2743 10.6151
R19517 vdd.n2743 vdd.n2742 10.6151
R19518 vdd.n2742 vdd.n2740 10.6151
R19519 vdd.n2740 vdd.n2739 10.6151
R19520 vdd.n2739 vdd.n2737 10.6151
R19521 vdd.n2737 vdd.n2736 10.6151
R19522 vdd.n2736 vdd.n2734 10.6151
R19523 vdd.n2734 vdd.n2733 10.6151
R19524 vdd.n2733 vdd.n807 10.6151
R19525 vdd.n3001 vdd.n807 10.6151
R19526 vdd.n3002 vdd.n3001 10.6151
R19527 vdd.n2852 vdd.n2851 10.6151
R19528 vdd.n2851 vdd.n2850 10.6151
R19529 vdd.n2850 vdd.n2849 10.6151
R19530 vdd.n2849 vdd.n2847 10.6151
R19531 vdd.n2847 vdd.n2844 10.6151
R19532 vdd.n2844 vdd.n2843 10.6151
R19533 vdd.n2843 vdd.n2840 10.6151
R19534 vdd.n2840 vdd.n2839 10.6151
R19535 vdd.n2839 vdd.n2836 10.6151
R19536 vdd.n2836 vdd.n2835 10.6151
R19537 vdd.n2835 vdd.n2832 10.6151
R19538 vdd.n2832 vdd.n2831 10.6151
R19539 vdd.n2831 vdd.n2828 10.6151
R19540 vdd.n2828 vdd.n2827 10.6151
R19541 vdd.n2827 vdd.n2824 10.6151
R19542 vdd.n2824 vdd.n2823 10.6151
R19543 vdd.n2823 vdd.n2820 10.6151
R19544 vdd.n2820 vdd.n2819 10.6151
R19545 vdd.n2819 vdd.n2816 10.6151
R19546 vdd.n2816 vdd.n2815 10.6151
R19547 vdd.n2815 vdd.n2812 10.6151
R19548 vdd.n2812 vdd.n2811 10.6151
R19549 vdd.n2811 vdd.n2808 10.6151
R19550 vdd.n2808 vdd.n2807 10.6151
R19551 vdd.n2807 vdd.n2804 10.6151
R19552 vdd.n2804 vdd.n2803 10.6151
R19553 vdd.n2803 vdd.n2800 10.6151
R19554 vdd.n2800 vdd.n2799 10.6151
R19555 vdd.n2799 vdd.n2796 10.6151
R19556 vdd.n2796 vdd.n2795 10.6151
R19557 vdd.n2795 vdd.n2792 10.6151
R19558 vdd.n2790 vdd.n2787 10.6151
R19559 vdd.n2787 vdd.n2786 10.6151
R19560 vdd.n2864 vdd.n897 10.6151
R19561 vdd.n2865 vdd.n2864 10.6151
R19562 vdd.n2866 vdd.n2865 10.6151
R19563 vdd.n2866 vdd.n886 10.6151
R19564 vdd.n2876 vdd.n886 10.6151
R19565 vdd.n2877 vdd.n2876 10.6151
R19566 vdd.n2878 vdd.n2877 10.6151
R19567 vdd.n2878 vdd.n874 10.6151
R19568 vdd.n2888 vdd.n874 10.6151
R19569 vdd.n2889 vdd.n2888 10.6151
R19570 vdd.n2890 vdd.n2889 10.6151
R19571 vdd.n2890 vdd.n862 10.6151
R19572 vdd.n2900 vdd.n862 10.6151
R19573 vdd.n2901 vdd.n2900 10.6151
R19574 vdd.n2902 vdd.n2901 10.6151
R19575 vdd.n2902 vdd.n851 10.6151
R19576 vdd.n2912 vdd.n851 10.6151
R19577 vdd.n2913 vdd.n2912 10.6151
R19578 vdd.n2914 vdd.n2913 10.6151
R19579 vdd.n2914 vdd.n837 10.6151
R19580 vdd.n2925 vdd.n837 10.6151
R19581 vdd.n2926 vdd.n2925 10.6151
R19582 vdd.n2927 vdd.n2926 10.6151
R19583 vdd.n2927 vdd.n826 10.6151
R19584 vdd.n2937 vdd.n826 10.6151
R19585 vdd.n2938 vdd.n2937 10.6151
R19586 vdd.n2939 vdd.n2938 10.6151
R19587 vdd.n2939 vdd.n812 10.6151
R19588 vdd.n2994 vdd.n812 10.6151
R19589 vdd.n2995 vdd.n2994 10.6151
R19590 vdd.n2996 vdd.n2995 10.6151
R19591 vdd.n2996 vdd.n779 10.6151
R19592 vdd.n3066 vdd.n779 10.6151
R19593 vdd.n3065 vdd.n3064 10.6151
R19594 vdd.n3064 vdd.n780 10.6151
R19595 vdd.n781 vdd.n780 10.6151
R19596 vdd.n3057 vdd.n781 10.6151
R19597 vdd.n3057 vdd.n3056 10.6151
R19598 vdd.n3056 vdd.n3055 10.6151
R19599 vdd.n3055 vdd.n783 10.6151
R19600 vdd.n3050 vdd.n783 10.6151
R19601 vdd.n3050 vdd.n3049 10.6151
R19602 vdd.n3049 vdd.n3048 10.6151
R19603 vdd.n3048 vdd.n786 10.6151
R19604 vdd.n3043 vdd.n786 10.6151
R19605 vdd.n3043 vdd.n3042 10.6151
R19606 vdd.n3042 vdd.n3041 10.6151
R19607 vdd.n3041 vdd.n789 10.6151
R19608 vdd.n3036 vdd.n789 10.6151
R19609 vdd.n3036 vdd.n3035 10.6151
R19610 vdd.n3035 vdd.n3033 10.6151
R19611 vdd.n3033 vdd.n792 10.6151
R19612 vdd.n3028 vdd.n792 10.6151
R19613 vdd.n3028 vdd.n3027 10.6151
R19614 vdd.n3027 vdd.n3026 10.6151
R19615 vdd.n3026 vdd.n795 10.6151
R19616 vdd.n3021 vdd.n795 10.6151
R19617 vdd.n3021 vdd.n3020 10.6151
R19618 vdd.n3020 vdd.n3019 10.6151
R19619 vdd.n3019 vdd.n798 10.6151
R19620 vdd.n3014 vdd.n798 10.6151
R19621 vdd.n3014 vdd.n3013 10.6151
R19622 vdd.n3013 vdd.n3012 10.6151
R19623 vdd.n3012 vdd.n801 10.6151
R19624 vdd.n3007 vdd.n3006 10.6151
R19625 vdd.n3006 vdd.n3005 10.6151
R19626 vdd.n2984 vdd.n2945 10.6151
R19627 vdd.n2979 vdd.n2945 10.6151
R19628 vdd.n2979 vdd.n2978 10.6151
R19629 vdd.n2978 vdd.n2977 10.6151
R19630 vdd.n2977 vdd.n2947 10.6151
R19631 vdd.n2972 vdd.n2947 10.6151
R19632 vdd.n2972 vdd.n2971 10.6151
R19633 vdd.n2971 vdd.n2970 10.6151
R19634 vdd.n2970 vdd.n2950 10.6151
R19635 vdd.n2965 vdd.n2950 10.6151
R19636 vdd.n2965 vdd.n2964 10.6151
R19637 vdd.n2964 vdd.n2963 10.6151
R19638 vdd.n2963 vdd.n2953 10.6151
R19639 vdd.n2958 vdd.n2953 10.6151
R19640 vdd.n2958 vdd.n2957 10.6151
R19641 vdd.n2957 vdd.n753 10.6151
R19642 vdd.n3101 vdd.n753 10.6151
R19643 vdd.n3101 vdd.n754 10.6151
R19644 vdd.n757 vdd.n754 10.6151
R19645 vdd.n3094 vdd.n757 10.6151
R19646 vdd.n3094 vdd.n3093 10.6151
R19647 vdd.n3093 vdd.n3092 10.6151
R19648 vdd.n3092 vdd.n759 10.6151
R19649 vdd.n3087 vdd.n759 10.6151
R19650 vdd.n3087 vdd.n3086 10.6151
R19651 vdd.n3086 vdd.n3085 10.6151
R19652 vdd.n3085 vdd.n762 10.6151
R19653 vdd.n3080 vdd.n762 10.6151
R19654 vdd.n3080 vdd.n3079 10.6151
R19655 vdd.n3079 vdd.n3078 10.6151
R19656 vdd.n3078 vdd.n765 10.6151
R19657 vdd.n3073 vdd.n3072 10.6151
R19658 vdd.n3072 vdd.n3071 10.6151
R19659 vdd.n2691 vdd.n2690 10.6151
R19660 vdd.n2777 vdd.n2691 10.6151
R19661 vdd.n2777 vdd.n2776 10.6151
R19662 vdd.n2776 vdd.n2775 10.6151
R19663 vdd.n2775 vdd.n2773 10.6151
R19664 vdd.n2773 vdd.n2772 10.6151
R19665 vdd.n2772 vdd.n2770 10.6151
R19666 vdd.n2770 vdd.n2769 10.6151
R19667 vdd.n2769 vdd.n2767 10.6151
R19668 vdd.n2767 vdd.n2766 10.6151
R19669 vdd.n2766 vdd.n2723 10.6151
R19670 vdd.n2723 vdd.n2722 10.6151
R19671 vdd.n2722 vdd.n2720 10.6151
R19672 vdd.n2720 vdd.n2719 10.6151
R19673 vdd.n2719 vdd.n2717 10.6151
R19674 vdd.n2717 vdd.n2716 10.6151
R19675 vdd.n2716 vdd.n2714 10.6151
R19676 vdd.n2714 vdd.n2713 10.6151
R19677 vdd.n2713 vdd.n2711 10.6151
R19678 vdd.n2711 vdd.n2710 10.6151
R19679 vdd.n2710 vdd.n2708 10.6151
R19680 vdd.n2708 vdd.n2707 10.6151
R19681 vdd.n2707 vdd.n2705 10.6151
R19682 vdd.n2705 vdd.n2704 10.6151
R19683 vdd.n2704 vdd.n2702 10.6151
R19684 vdd.n2702 vdd.n2701 10.6151
R19685 vdd.n2701 vdd.n2699 10.6151
R19686 vdd.n2699 vdd.n2698 10.6151
R19687 vdd.n2698 vdd.n2696 10.6151
R19688 vdd.n2696 vdd.n2695 10.6151
R19689 vdd.n2695 vdd.n2693 10.6151
R19690 vdd.n2693 vdd.n2692 10.6151
R19691 vdd.n2692 vdd.n771 10.6151
R19692 vdd.n2858 vdd.n903 10.6151
R19693 vdd.n2625 vdd.n903 10.6151
R19694 vdd.n2626 vdd.n2625 10.6151
R19695 vdd.n2629 vdd.n2626 10.6151
R19696 vdd.n2630 vdd.n2629 10.6151
R19697 vdd.n2633 vdd.n2630 10.6151
R19698 vdd.n2634 vdd.n2633 10.6151
R19699 vdd.n2637 vdd.n2634 10.6151
R19700 vdd.n2638 vdd.n2637 10.6151
R19701 vdd.n2641 vdd.n2638 10.6151
R19702 vdd.n2642 vdd.n2641 10.6151
R19703 vdd.n2645 vdd.n2642 10.6151
R19704 vdd.n2646 vdd.n2645 10.6151
R19705 vdd.n2649 vdd.n2646 10.6151
R19706 vdd.n2650 vdd.n2649 10.6151
R19707 vdd.n2653 vdd.n2650 10.6151
R19708 vdd.n2654 vdd.n2653 10.6151
R19709 vdd.n2657 vdd.n2654 10.6151
R19710 vdd.n2658 vdd.n2657 10.6151
R19711 vdd.n2661 vdd.n2658 10.6151
R19712 vdd.n2662 vdd.n2661 10.6151
R19713 vdd.n2665 vdd.n2662 10.6151
R19714 vdd.n2666 vdd.n2665 10.6151
R19715 vdd.n2669 vdd.n2666 10.6151
R19716 vdd.n2670 vdd.n2669 10.6151
R19717 vdd.n2673 vdd.n2670 10.6151
R19718 vdd.n2674 vdd.n2673 10.6151
R19719 vdd.n2677 vdd.n2674 10.6151
R19720 vdd.n2678 vdd.n2677 10.6151
R19721 vdd.n2681 vdd.n2678 10.6151
R19722 vdd.n2682 vdd.n2681 10.6151
R19723 vdd.n2687 vdd.n2685 10.6151
R19724 vdd.n2688 vdd.n2687 10.6151
R19725 vdd.n2860 vdd.n2859 10.6151
R19726 vdd.n2860 vdd.n892 10.6151
R19727 vdd.n2870 vdd.n892 10.6151
R19728 vdd.n2871 vdd.n2870 10.6151
R19729 vdd.n2872 vdd.n2871 10.6151
R19730 vdd.n2872 vdd.n880 10.6151
R19731 vdd.n2882 vdd.n880 10.6151
R19732 vdd.n2883 vdd.n2882 10.6151
R19733 vdd.n2884 vdd.n2883 10.6151
R19734 vdd.n2884 vdd.n868 10.6151
R19735 vdd.n2894 vdd.n868 10.6151
R19736 vdd.n2895 vdd.n2894 10.6151
R19737 vdd.n2896 vdd.n2895 10.6151
R19738 vdd.n2896 vdd.n857 10.6151
R19739 vdd.n2906 vdd.n857 10.6151
R19740 vdd.n2907 vdd.n2906 10.6151
R19741 vdd.n2908 vdd.n2907 10.6151
R19742 vdd.n2908 vdd.n844 10.6151
R19743 vdd.n2918 vdd.n844 10.6151
R19744 vdd.n2919 vdd.n2918 10.6151
R19745 vdd.n2921 vdd.n832 10.6151
R19746 vdd.n2931 vdd.n832 10.6151
R19747 vdd.n2932 vdd.n2931 10.6151
R19748 vdd.n2933 vdd.n2932 10.6151
R19749 vdd.n2933 vdd.n820 10.6151
R19750 vdd.n2943 vdd.n820 10.6151
R19751 vdd.n2944 vdd.n2943 10.6151
R19752 vdd.n2990 vdd.n2944 10.6151
R19753 vdd.n2990 vdd.n2989 10.6151
R19754 vdd.n2989 vdd.n2988 10.6151
R19755 vdd.n2988 vdd.n2987 10.6151
R19756 vdd.n2987 vdd.n2985 10.6151
R19757 vdd.n2339 vdd.n2338 10.6151
R19758 vdd.n2339 vdd.n1040 10.6151
R19759 vdd.n2349 vdd.n1040 10.6151
R19760 vdd.n2350 vdd.n2349 10.6151
R19761 vdd.n2351 vdd.n2350 10.6151
R19762 vdd.n2351 vdd.n1028 10.6151
R19763 vdd.n2361 vdd.n1028 10.6151
R19764 vdd.n2362 vdd.n2361 10.6151
R19765 vdd.n2363 vdd.n2362 10.6151
R19766 vdd.n2363 vdd.n1015 10.6151
R19767 vdd.n2373 vdd.n1015 10.6151
R19768 vdd.n2374 vdd.n2373 10.6151
R19769 vdd.n2376 vdd.n1003 10.6151
R19770 vdd.n2386 vdd.n1003 10.6151
R19771 vdd.n2387 vdd.n2386 10.6151
R19772 vdd.n2388 vdd.n2387 10.6151
R19773 vdd.n2388 vdd.n991 10.6151
R19774 vdd.n2398 vdd.n991 10.6151
R19775 vdd.n2399 vdd.n2398 10.6151
R19776 vdd.n2400 vdd.n2399 10.6151
R19777 vdd.n2400 vdd.n980 10.6151
R19778 vdd.n2410 vdd.n980 10.6151
R19779 vdd.n2411 vdd.n2410 10.6151
R19780 vdd.n2412 vdd.n2411 10.6151
R19781 vdd.n2412 vdd.n968 10.6151
R19782 vdd.n2422 vdd.n968 10.6151
R19783 vdd.n2423 vdd.n2422 10.6151
R19784 vdd.n2426 vdd.n2423 10.6151
R19785 vdd.n2426 vdd.n2425 10.6151
R19786 vdd.n2425 vdd.n2424 10.6151
R19787 vdd.n2424 vdd.n951 10.6151
R19788 vdd.n2508 vdd.n951 10.6151
R19789 vdd.n2507 vdd.n2506 10.6151
R19790 vdd.n2506 vdd.n2503 10.6151
R19791 vdd.n2503 vdd.n2502 10.6151
R19792 vdd.n2502 vdd.n2499 10.6151
R19793 vdd.n2499 vdd.n2498 10.6151
R19794 vdd.n2498 vdd.n2495 10.6151
R19795 vdd.n2495 vdd.n2494 10.6151
R19796 vdd.n2494 vdd.n2491 10.6151
R19797 vdd.n2491 vdd.n2490 10.6151
R19798 vdd.n2490 vdd.n2487 10.6151
R19799 vdd.n2487 vdd.n2486 10.6151
R19800 vdd.n2486 vdd.n2483 10.6151
R19801 vdd.n2483 vdd.n2482 10.6151
R19802 vdd.n2482 vdd.n2479 10.6151
R19803 vdd.n2479 vdd.n2478 10.6151
R19804 vdd.n2478 vdd.n2475 10.6151
R19805 vdd.n2475 vdd.n2474 10.6151
R19806 vdd.n2474 vdd.n2471 10.6151
R19807 vdd.n2471 vdd.n2470 10.6151
R19808 vdd.n2470 vdd.n2467 10.6151
R19809 vdd.n2467 vdd.n2466 10.6151
R19810 vdd.n2466 vdd.n2463 10.6151
R19811 vdd.n2463 vdd.n2462 10.6151
R19812 vdd.n2462 vdd.n2459 10.6151
R19813 vdd.n2459 vdd.n2458 10.6151
R19814 vdd.n2458 vdd.n2455 10.6151
R19815 vdd.n2455 vdd.n2454 10.6151
R19816 vdd.n2454 vdd.n2451 10.6151
R19817 vdd.n2451 vdd.n2450 10.6151
R19818 vdd.n2450 vdd.n2447 10.6151
R19819 vdd.n2447 vdd.n2446 10.6151
R19820 vdd.n2443 vdd.n2442 10.6151
R19821 vdd.n2442 vdd.n2440 10.6151
R19822 vdd.n1359 vdd.n1357 10.6151
R19823 vdd.n1357 vdd.n1356 10.6151
R19824 vdd.n1356 vdd.n1354 10.6151
R19825 vdd.n1354 vdd.n1353 10.6151
R19826 vdd.n1353 vdd.n1351 10.6151
R19827 vdd.n1351 vdd.n1350 10.6151
R19828 vdd.n1350 vdd.n1348 10.6151
R19829 vdd.n1348 vdd.n1347 10.6151
R19830 vdd.n1347 vdd.n1345 10.6151
R19831 vdd.n1345 vdd.n1344 10.6151
R19832 vdd.n1344 vdd.n1342 10.6151
R19833 vdd.n1342 vdd.n1341 10.6151
R19834 vdd.n1341 vdd.n1339 10.6151
R19835 vdd.n1339 vdd.n1338 10.6151
R19836 vdd.n1338 vdd.n1336 10.6151
R19837 vdd.n1336 vdd.n1335 10.6151
R19838 vdd.n1335 vdd.n1333 10.6151
R19839 vdd.n1333 vdd.n1332 10.6151
R19840 vdd.n1332 vdd.n1243 10.6151
R19841 vdd.n1243 vdd.n1242 10.6151
R19842 vdd.n1242 vdd.n1240 10.6151
R19843 vdd.n1240 vdd.n1239 10.6151
R19844 vdd.n1239 vdd.n1237 10.6151
R19845 vdd.n1237 vdd.n1236 10.6151
R19846 vdd.n1236 vdd.n1234 10.6151
R19847 vdd.n1234 vdd.n1233 10.6151
R19848 vdd.n1233 vdd.n1231 10.6151
R19849 vdd.n1231 vdd.n1230 10.6151
R19850 vdd.n1230 vdd.n1228 10.6151
R19851 vdd.n1228 vdd.n1227 10.6151
R19852 vdd.n1227 vdd.n955 10.6151
R19853 vdd.n2438 vdd.n955 10.6151
R19854 vdd.n2439 vdd.n2438 10.6151
R19855 vdd.n2337 vdd.n1052 10.6151
R19856 vdd.n1194 vdd.n1052 10.6151
R19857 vdd.n1195 vdd.n1194 10.6151
R19858 vdd.n1198 vdd.n1195 10.6151
R19859 vdd.n1199 vdd.n1198 10.6151
R19860 vdd.n1202 vdd.n1199 10.6151
R19861 vdd.n1203 vdd.n1202 10.6151
R19862 vdd.n1206 vdd.n1203 10.6151
R19863 vdd.n1207 vdd.n1206 10.6151
R19864 vdd.n1210 vdd.n1207 10.6151
R19865 vdd.n1211 vdd.n1210 10.6151
R19866 vdd.n1214 vdd.n1211 10.6151
R19867 vdd.n1215 vdd.n1214 10.6151
R19868 vdd.n1218 vdd.n1215 10.6151
R19869 vdd.n1219 vdd.n1218 10.6151
R19870 vdd.n1222 vdd.n1219 10.6151
R19871 vdd.n1393 vdd.n1222 10.6151
R19872 vdd.n1393 vdd.n1392 10.6151
R19873 vdd.n1392 vdd.n1390 10.6151
R19874 vdd.n1390 vdd.n1387 10.6151
R19875 vdd.n1387 vdd.n1386 10.6151
R19876 vdd.n1386 vdd.n1383 10.6151
R19877 vdd.n1383 vdd.n1382 10.6151
R19878 vdd.n1382 vdd.n1379 10.6151
R19879 vdd.n1379 vdd.n1378 10.6151
R19880 vdd.n1378 vdd.n1375 10.6151
R19881 vdd.n1375 vdd.n1374 10.6151
R19882 vdd.n1374 vdd.n1371 10.6151
R19883 vdd.n1371 vdd.n1370 10.6151
R19884 vdd.n1370 vdd.n1367 10.6151
R19885 vdd.n1367 vdd.n1366 10.6151
R19886 vdd.n1363 vdd.n1362 10.6151
R19887 vdd.n1362 vdd.n1360 10.6151
R19888 vdd.t231 vdd.n2138 10.5435
R19889 vdd.n636 vdd.t185 10.5435
R19890 vdd.n304 vdd.n286 10.4732
R19891 vdd.n249 vdd.n231 10.4732
R19892 vdd.n206 vdd.n188 10.4732
R19893 vdd.n151 vdd.n133 10.4732
R19894 vdd.n109 vdd.n91 10.4732
R19895 vdd.n54 vdd.n36 10.4732
R19896 vdd.n2035 vdd.n2017 10.4732
R19897 vdd.n2090 vdd.n2072 10.4732
R19898 vdd.n1937 vdd.n1919 10.4732
R19899 vdd.n1992 vdd.n1974 10.4732
R19900 vdd.n1840 vdd.n1822 10.4732
R19901 vdd.n1895 vdd.n1877 10.4732
R19902 vdd.n2122 vdd.t191 10.3167
R19903 vdd.n3297 vdd.t180 10.3167
R19904 vdd.t213 vdd.n1466 10.09
R19905 vdd.n2174 vdd.t62 10.09
R19906 vdd.n3245 vdd.t58 10.09
R19907 vdd.n3378 vdd.t183 10.09
R19908 vdd.n1786 vdd.t168 9.86327
R19909 vdd.n3369 vdd.t228 9.86327
R19910 vdd.n2299 vdd.n2298 9.78206
R19911 vdd.n3035 vdd.n3034 9.78206
R19912 vdd.n3102 vdd.n3101 9.78206
R19913 vdd.n2191 vdd.n1393 9.78206
R19914 vdd.n303 vdd.n288 9.69747
R19915 vdd.n248 vdd.n233 9.69747
R19916 vdd.n205 vdd.n190 9.69747
R19917 vdd.n150 vdd.n135 9.69747
R19918 vdd.n108 vdd.n93 9.69747
R19919 vdd.n53 vdd.n38 9.69747
R19920 vdd.n2034 vdd.n2019 9.69747
R19921 vdd.n2089 vdd.n2074 9.69747
R19922 vdd.n1936 vdd.n1921 9.69747
R19923 vdd.n1991 vdd.n1976 9.69747
R19924 vdd.n1839 vdd.n1824 9.69747
R19925 vdd.n1894 vdd.n1879 9.69747
R19926 vdd.t142 vdd.n1760 9.63654
R19927 vdd.n3328 vdd.t194 9.63654
R19928 vdd.n319 vdd.n318 9.45567
R19929 vdd.n264 vdd.n263 9.45567
R19930 vdd.n221 vdd.n220 9.45567
R19931 vdd.n166 vdd.n165 9.45567
R19932 vdd.n124 vdd.n123 9.45567
R19933 vdd.n69 vdd.n68 9.45567
R19934 vdd.n2050 vdd.n2049 9.45567
R19935 vdd.n2105 vdd.n2104 9.45567
R19936 vdd.n1952 vdd.n1951 9.45567
R19937 vdd.n2007 vdd.n2006 9.45567
R19938 vdd.n1855 vdd.n1854 9.45567
R19939 vdd.n1910 vdd.n1909 9.45567
R19940 vdd.n2261 vdd.n1120 9.3005
R19941 vdd.n2260 vdd.n2259 9.3005
R19942 vdd.n1126 vdd.n1125 9.3005
R19943 vdd.n2254 vdd.n1130 9.3005
R19944 vdd.n2253 vdd.n1131 9.3005
R19945 vdd.n2252 vdd.n1132 9.3005
R19946 vdd.n1136 vdd.n1133 9.3005
R19947 vdd.n2247 vdd.n1137 9.3005
R19948 vdd.n2246 vdd.n1138 9.3005
R19949 vdd.n2245 vdd.n1139 9.3005
R19950 vdd.n1143 vdd.n1140 9.3005
R19951 vdd.n2240 vdd.n1144 9.3005
R19952 vdd.n2239 vdd.n1145 9.3005
R19953 vdd.n2238 vdd.n1146 9.3005
R19954 vdd.n1150 vdd.n1147 9.3005
R19955 vdd.n2233 vdd.n1151 9.3005
R19956 vdd.n2232 vdd.n1152 9.3005
R19957 vdd.n2231 vdd.n1153 9.3005
R19958 vdd.n1157 vdd.n1154 9.3005
R19959 vdd.n2226 vdd.n1158 9.3005
R19960 vdd.n2225 vdd.n1159 9.3005
R19961 vdd.n2224 vdd.n2223 9.3005
R19962 vdd.n2222 vdd.n1160 9.3005
R19963 vdd.n2221 vdd.n2220 9.3005
R19964 vdd.n1166 vdd.n1165 9.3005
R19965 vdd.n2215 vdd.n1170 9.3005
R19966 vdd.n2214 vdd.n1171 9.3005
R19967 vdd.n2213 vdd.n1172 9.3005
R19968 vdd.n1176 vdd.n1173 9.3005
R19969 vdd.n2208 vdd.n1177 9.3005
R19970 vdd.n2207 vdd.n1178 9.3005
R19971 vdd.n2206 vdd.n1179 9.3005
R19972 vdd.n1183 vdd.n1180 9.3005
R19973 vdd.n2201 vdd.n1184 9.3005
R19974 vdd.n2200 vdd.n1185 9.3005
R19975 vdd.n2199 vdd.n1186 9.3005
R19976 vdd.n1190 vdd.n1187 9.3005
R19977 vdd.n2194 vdd.n1191 9.3005
R19978 vdd.n2263 vdd.n2262 9.3005
R19979 vdd.n2285 vdd.n1091 9.3005
R19980 vdd.n2284 vdd.n1099 9.3005
R19981 vdd.n1103 vdd.n1100 9.3005
R19982 vdd.n2279 vdd.n1104 9.3005
R19983 vdd.n2278 vdd.n1105 9.3005
R19984 vdd.n2277 vdd.n1106 9.3005
R19985 vdd.n1110 vdd.n1107 9.3005
R19986 vdd.n2272 vdd.n1111 9.3005
R19987 vdd.n2271 vdd.n1112 9.3005
R19988 vdd.n2270 vdd.n1113 9.3005
R19989 vdd.n1117 vdd.n1114 9.3005
R19990 vdd.n2265 vdd.n1118 9.3005
R19991 vdd.n2264 vdd.n1119 9.3005
R19992 vdd.n2297 vdd.n2296 9.3005
R19993 vdd.n1095 vdd.n1094 9.3005
R19994 vdd.n2110 vdd.n1456 9.3005
R19995 vdd.n2112 vdd.n2111 9.3005
R19996 vdd.n1447 vdd.n1446 9.3005
R19997 vdd.n2125 vdd.n2124 9.3005
R19998 vdd.n2126 vdd.n1445 9.3005
R19999 vdd.n2128 vdd.n2127 9.3005
R20000 vdd.n1435 vdd.n1434 9.3005
R20001 vdd.n2142 vdd.n2141 9.3005
R20002 vdd.n2143 vdd.n1433 9.3005
R20003 vdd.n2145 vdd.n2144 9.3005
R20004 vdd.n1424 vdd.n1423 9.3005
R20005 vdd.n2159 vdd.n2158 9.3005
R20006 vdd.n2160 vdd.n1422 9.3005
R20007 vdd.n2162 vdd.n2161 9.3005
R20008 vdd.n1412 vdd.n1411 9.3005
R20009 vdd.n2177 vdd.n2176 9.3005
R20010 vdd.n2178 vdd.n1410 9.3005
R20011 vdd.n2180 vdd.n2179 9.3005
R20012 vdd.n295 vdd.n294 9.3005
R20013 vdd.n290 vdd.n289 9.3005
R20014 vdd.n301 vdd.n300 9.3005
R20015 vdd.n303 vdd.n302 9.3005
R20016 vdd.n286 vdd.n285 9.3005
R20017 vdd.n309 vdd.n308 9.3005
R20018 vdd.n311 vdd.n310 9.3005
R20019 vdd.n283 vdd.n280 9.3005
R20020 vdd.n318 vdd.n317 9.3005
R20021 vdd.n240 vdd.n239 9.3005
R20022 vdd.n235 vdd.n234 9.3005
R20023 vdd.n246 vdd.n245 9.3005
R20024 vdd.n248 vdd.n247 9.3005
R20025 vdd.n231 vdd.n230 9.3005
R20026 vdd.n254 vdd.n253 9.3005
R20027 vdd.n256 vdd.n255 9.3005
R20028 vdd.n228 vdd.n225 9.3005
R20029 vdd.n263 vdd.n262 9.3005
R20030 vdd.n197 vdd.n196 9.3005
R20031 vdd.n192 vdd.n191 9.3005
R20032 vdd.n203 vdd.n202 9.3005
R20033 vdd.n205 vdd.n204 9.3005
R20034 vdd.n188 vdd.n187 9.3005
R20035 vdd.n211 vdd.n210 9.3005
R20036 vdd.n213 vdd.n212 9.3005
R20037 vdd.n185 vdd.n182 9.3005
R20038 vdd.n220 vdd.n219 9.3005
R20039 vdd.n142 vdd.n141 9.3005
R20040 vdd.n137 vdd.n136 9.3005
R20041 vdd.n148 vdd.n147 9.3005
R20042 vdd.n150 vdd.n149 9.3005
R20043 vdd.n133 vdd.n132 9.3005
R20044 vdd.n156 vdd.n155 9.3005
R20045 vdd.n158 vdd.n157 9.3005
R20046 vdd.n130 vdd.n127 9.3005
R20047 vdd.n165 vdd.n164 9.3005
R20048 vdd.n100 vdd.n99 9.3005
R20049 vdd.n95 vdd.n94 9.3005
R20050 vdd.n106 vdd.n105 9.3005
R20051 vdd.n108 vdd.n107 9.3005
R20052 vdd.n91 vdd.n90 9.3005
R20053 vdd.n114 vdd.n113 9.3005
R20054 vdd.n116 vdd.n115 9.3005
R20055 vdd.n88 vdd.n85 9.3005
R20056 vdd.n123 vdd.n122 9.3005
R20057 vdd.n45 vdd.n44 9.3005
R20058 vdd.n40 vdd.n39 9.3005
R20059 vdd.n51 vdd.n50 9.3005
R20060 vdd.n53 vdd.n52 9.3005
R20061 vdd.n36 vdd.n35 9.3005
R20062 vdd.n59 vdd.n58 9.3005
R20063 vdd.n61 vdd.n60 9.3005
R20064 vdd.n33 vdd.n30 9.3005
R20065 vdd.n68 vdd.n67 9.3005
R20066 vdd.n3151 vdd.n3150 9.3005
R20067 vdd.n3152 vdd.n721 9.3005
R20068 vdd.n720 vdd.n718 9.3005
R20069 vdd.n3158 vdd.n717 9.3005
R20070 vdd.n3159 vdd.n716 9.3005
R20071 vdd.n3160 vdd.n715 9.3005
R20072 vdd.n714 vdd.n712 9.3005
R20073 vdd.n3166 vdd.n711 9.3005
R20074 vdd.n3167 vdd.n710 9.3005
R20075 vdd.n3168 vdd.n709 9.3005
R20076 vdd.n708 vdd.n706 9.3005
R20077 vdd.n3174 vdd.n705 9.3005
R20078 vdd.n3175 vdd.n704 9.3005
R20079 vdd.n3176 vdd.n703 9.3005
R20080 vdd.n702 vdd.n700 9.3005
R20081 vdd.n3182 vdd.n699 9.3005
R20082 vdd.n3183 vdd.n698 9.3005
R20083 vdd.n3184 vdd.n697 9.3005
R20084 vdd.n696 vdd.n694 9.3005
R20085 vdd.n3190 vdd.n693 9.3005
R20086 vdd.n3191 vdd.n692 9.3005
R20087 vdd.n3192 vdd.n691 9.3005
R20088 vdd.n690 vdd.n688 9.3005
R20089 vdd.n3198 vdd.n685 9.3005
R20090 vdd.n3199 vdd.n684 9.3005
R20091 vdd.n3200 vdd.n683 9.3005
R20092 vdd.n682 vdd.n680 9.3005
R20093 vdd.n3206 vdd.n679 9.3005
R20094 vdd.n3207 vdd.n678 9.3005
R20095 vdd.n3208 vdd.n677 9.3005
R20096 vdd.n676 vdd.n674 9.3005
R20097 vdd.n3214 vdd.n673 9.3005
R20098 vdd.n3215 vdd.n672 9.3005
R20099 vdd.n3216 vdd.n671 9.3005
R20100 vdd.n670 vdd.n668 9.3005
R20101 vdd.n3221 vdd.n667 9.3005
R20102 vdd.n3231 vdd.n661 9.3005
R20103 vdd.n3233 vdd.n3232 9.3005
R20104 vdd.n652 vdd.n651 9.3005
R20105 vdd.n3248 vdd.n3247 9.3005
R20106 vdd.n3249 vdd.n650 9.3005
R20107 vdd.n3251 vdd.n3250 9.3005
R20108 vdd.n640 vdd.n639 9.3005
R20109 vdd.n3264 vdd.n3263 9.3005
R20110 vdd.n3265 vdd.n638 9.3005
R20111 vdd.n3267 vdd.n3266 9.3005
R20112 vdd.n628 vdd.n627 9.3005
R20113 vdd.n3281 vdd.n3280 9.3005
R20114 vdd.n3282 vdd.n626 9.3005
R20115 vdd.n3284 vdd.n3283 9.3005
R20116 vdd.n617 vdd.n616 9.3005
R20117 vdd.n3300 vdd.n3299 9.3005
R20118 vdd.n3301 vdd.n615 9.3005
R20119 vdd.n3303 vdd.n3302 9.3005
R20120 vdd.n324 vdd.n322 9.3005
R20121 vdd.n3235 vdd.n3234 9.3005
R20122 vdd.n3382 vdd.n3381 9.3005
R20123 vdd.n325 vdd.n323 9.3005
R20124 vdd.n3375 vdd.n334 9.3005
R20125 vdd.n3374 vdd.n335 9.3005
R20126 vdd.n3373 vdd.n336 9.3005
R20127 vdd.n343 vdd.n337 9.3005
R20128 vdd.n3367 vdd.n344 9.3005
R20129 vdd.n3366 vdd.n345 9.3005
R20130 vdd.n3365 vdd.n346 9.3005
R20131 vdd.n354 vdd.n347 9.3005
R20132 vdd.n3359 vdd.n355 9.3005
R20133 vdd.n3358 vdd.n356 9.3005
R20134 vdd.n3357 vdd.n357 9.3005
R20135 vdd.n365 vdd.n358 9.3005
R20136 vdd.n3351 vdd.n366 9.3005
R20137 vdd.n3350 vdd.n367 9.3005
R20138 vdd.n3349 vdd.n368 9.3005
R20139 vdd.n443 vdd.n369 9.3005
R20140 vdd.n447 vdd.n442 9.3005
R20141 vdd.n451 vdd.n450 9.3005
R20142 vdd.n452 vdd.n441 9.3005
R20143 vdd.n456 vdd.n453 9.3005
R20144 vdd.n457 vdd.n440 9.3005
R20145 vdd.n461 vdd.n460 9.3005
R20146 vdd.n462 vdd.n439 9.3005
R20147 vdd.n466 vdd.n463 9.3005
R20148 vdd.n467 vdd.n438 9.3005
R20149 vdd.n471 vdd.n470 9.3005
R20150 vdd.n472 vdd.n437 9.3005
R20151 vdd.n476 vdd.n473 9.3005
R20152 vdd.n477 vdd.n436 9.3005
R20153 vdd.n481 vdd.n480 9.3005
R20154 vdd.n482 vdd.n435 9.3005
R20155 vdd.n486 vdd.n483 9.3005
R20156 vdd.n487 vdd.n434 9.3005
R20157 vdd.n491 vdd.n490 9.3005
R20158 vdd.n492 vdd.n433 9.3005
R20159 vdd.n496 vdd.n493 9.3005
R20160 vdd.n497 vdd.n430 9.3005
R20161 vdd.n501 vdd.n500 9.3005
R20162 vdd.n502 vdd.n429 9.3005
R20163 vdd.n506 vdd.n503 9.3005
R20164 vdd.n507 vdd.n428 9.3005
R20165 vdd.n511 vdd.n510 9.3005
R20166 vdd.n512 vdd.n427 9.3005
R20167 vdd.n516 vdd.n513 9.3005
R20168 vdd.n517 vdd.n426 9.3005
R20169 vdd.n521 vdd.n520 9.3005
R20170 vdd.n522 vdd.n425 9.3005
R20171 vdd.n526 vdd.n523 9.3005
R20172 vdd.n527 vdd.n424 9.3005
R20173 vdd.n531 vdd.n530 9.3005
R20174 vdd.n532 vdd.n423 9.3005
R20175 vdd.n536 vdd.n533 9.3005
R20176 vdd.n537 vdd.n422 9.3005
R20177 vdd.n541 vdd.n540 9.3005
R20178 vdd.n542 vdd.n421 9.3005
R20179 vdd.n546 vdd.n543 9.3005
R20180 vdd.n547 vdd.n418 9.3005
R20181 vdd.n551 vdd.n550 9.3005
R20182 vdd.n552 vdd.n417 9.3005
R20183 vdd.n556 vdd.n553 9.3005
R20184 vdd.n557 vdd.n416 9.3005
R20185 vdd.n561 vdd.n560 9.3005
R20186 vdd.n562 vdd.n415 9.3005
R20187 vdd.n566 vdd.n563 9.3005
R20188 vdd.n567 vdd.n414 9.3005
R20189 vdd.n571 vdd.n570 9.3005
R20190 vdd.n572 vdd.n413 9.3005
R20191 vdd.n576 vdd.n573 9.3005
R20192 vdd.n577 vdd.n412 9.3005
R20193 vdd.n581 vdd.n580 9.3005
R20194 vdd.n582 vdd.n411 9.3005
R20195 vdd.n586 vdd.n583 9.3005
R20196 vdd.n587 vdd.n410 9.3005
R20197 vdd.n591 vdd.n590 9.3005
R20198 vdd.n592 vdd.n409 9.3005
R20199 vdd.n596 vdd.n593 9.3005
R20200 vdd.n598 vdd.n408 9.3005
R20201 vdd.n600 vdd.n599 9.3005
R20202 vdd.n3342 vdd.n3341 9.3005
R20203 vdd.n446 vdd.n444 9.3005
R20204 vdd.n3241 vdd.n655 9.3005
R20205 vdd.n3243 vdd.n3242 9.3005
R20206 vdd.n646 vdd.n645 9.3005
R20207 vdd.n3256 vdd.n3255 9.3005
R20208 vdd.n3257 vdd.n644 9.3005
R20209 vdd.n3259 vdd.n3258 9.3005
R20210 vdd.n633 vdd.n632 9.3005
R20211 vdd.n3272 vdd.n3271 9.3005
R20212 vdd.n3273 vdd.n631 9.3005
R20213 vdd.n3275 vdd.n3274 9.3005
R20214 vdd.n622 vdd.n621 9.3005
R20215 vdd.n3289 vdd.n3288 9.3005
R20216 vdd.n3290 vdd.n620 9.3005
R20217 vdd.n3295 vdd.n3291 9.3005
R20218 vdd.n3294 vdd.n3293 9.3005
R20219 vdd.n3292 vdd.n610 9.3005
R20220 vdd.n3308 vdd.n611 9.3005
R20221 vdd.n3309 vdd.n609 9.3005
R20222 vdd.n3311 vdd.n3310 9.3005
R20223 vdd.n3312 vdd.n608 9.3005
R20224 vdd.n3315 vdd.n3313 9.3005
R20225 vdd.n3316 vdd.n607 9.3005
R20226 vdd.n3318 vdd.n3317 9.3005
R20227 vdd.n3319 vdd.n606 9.3005
R20228 vdd.n3322 vdd.n3320 9.3005
R20229 vdd.n3323 vdd.n605 9.3005
R20230 vdd.n3325 vdd.n3324 9.3005
R20231 vdd.n3326 vdd.n604 9.3005
R20232 vdd.n3330 vdd.n3327 9.3005
R20233 vdd.n3331 vdd.n603 9.3005
R20234 vdd.n3333 vdd.n3332 9.3005
R20235 vdd.n3334 vdd.n602 9.3005
R20236 vdd.n3337 vdd.n3335 9.3005
R20237 vdd.n3338 vdd.n601 9.3005
R20238 vdd.n3340 vdd.n3339 9.3005
R20239 vdd.n3240 vdd.n3239 9.3005
R20240 vdd.n3104 vdd.n656 9.3005
R20241 vdd.n3109 vdd.n3103 9.3005
R20242 vdd.n3119 vdd.n748 9.3005
R20243 vdd.n3120 vdd.n747 9.3005
R20244 vdd.n746 vdd.n744 9.3005
R20245 vdd.n3126 vdd.n743 9.3005
R20246 vdd.n3127 vdd.n742 9.3005
R20247 vdd.n3128 vdd.n741 9.3005
R20248 vdd.n740 vdd.n738 9.3005
R20249 vdd.n3134 vdd.n737 9.3005
R20250 vdd.n3135 vdd.n736 9.3005
R20251 vdd.n3136 vdd.n735 9.3005
R20252 vdd.n734 vdd.n732 9.3005
R20253 vdd.n3141 vdd.n731 9.3005
R20254 vdd.n3142 vdd.n730 9.3005
R20255 vdd.n726 vdd.n725 9.3005
R20256 vdd.n3148 vdd.n3147 9.3005
R20257 vdd.n3149 vdd.n722 9.3005
R20258 vdd.n2190 vdd.n2189 9.3005
R20259 vdd.n2185 vdd.n1395 9.3005
R20260 vdd.n1742 vdd.n1741 9.3005
R20261 vdd.n1498 vdd.n1497 9.3005
R20262 vdd.n1755 vdd.n1754 9.3005
R20263 vdd.n1756 vdd.n1496 9.3005
R20264 vdd.n1758 vdd.n1757 9.3005
R20265 vdd.n1486 vdd.n1485 9.3005
R20266 vdd.n1772 vdd.n1771 9.3005
R20267 vdd.n1773 vdd.n1484 9.3005
R20268 vdd.n1775 vdd.n1774 9.3005
R20269 vdd.n1476 vdd.n1475 9.3005
R20270 vdd.n1789 vdd.n1788 9.3005
R20271 vdd.n1790 vdd.n1474 9.3005
R20272 vdd.n1792 vdd.n1791 9.3005
R20273 vdd.n1463 vdd.n1462 9.3005
R20274 vdd.n1805 vdd.n1804 9.3005
R20275 vdd.n1806 vdd.n1461 9.3005
R20276 vdd.n1808 vdd.n1807 9.3005
R20277 vdd.n1452 vdd.n1451 9.3005
R20278 vdd.n2117 vdd.n2116 9.3005
R20279 vdd.n2118 vdd.n1450 9.3005
R20280 vdd.n2120 vdd.n2119 9.3005
R20281 vdd.n1441 vdd.n1440 9.3005
R20282 vdd.n2133 vdd.n2132 9.3005
R20283 vdd.n2134 vdd.n1439 9.3005
R20284 vdd.n2136 vdd.n2135 9.3005
R20285 vdd.n1429 vdd.n1428 9.3005
R20286 vdd.n2150 vdd.n2149 9.3005
R20287 vdd.n2151 vdd.n1427 9.3005
R20288 vdd.n2153 vdd.n2152 9.3005
R20289 vdd.n1419 vdd.n1418 9.3005
R20290 vdd.n2167 vdd.n2166 9.3005
R20291 vdd.n2168 vdd.n1416 9.3005
R20292 vdd.n2172 vdd.n2171 9.3005
R20293 vdd.n2170 vdd.n1417 9.3005
R20294 vdd.n2169 vdd.n1406 9.3005
R20295 vdd.n1740 vdd.n1508 9.3005
R20296 vdd.n1633 vdd.n1509 9.3005
R20297 vdd.n1635 vdd.n1634 9.3005
R20298 vdd.n1636 vdd.n1628 9.3005
R20299 vdd.n1638 vdd.n1637 9.3005
R20300 vdd.n1639 vdd.n1627 9.3005
R20301 vdd.n1641 vdd.n1640 9.3005
R20302 vdd.n1642 vdd.n1622 9.3005
R20303 vdd.n1644 vdd.n1643 9.3005
R20304 vdd.n1645 vdd.n1621 9.3005
R20305 vdd.n1647 vdd.n1646 9.3005
R20306 vdd.n1648 vdd.n1616 9.3005
R20307 vdd.n1650 vdd.n1649 9.3005
R20308 vdd.n1651 vdd.n1615 9.3005
R20309 vdd.n1653 vdd.n1652 9.3005
R20310 vdd.n1654 vdd.n1610 9.3005
R20311 vdd.n1656 vdd.n1655 9.3005
R20312 vdd.n1657 vdd.n1609 9.3005
R20313 vdd.n1659 vdd.n1658 9.3005
R20314 vdd.n1660 vdd.n1604 9.3005
R20315 vdd.n1662 vdd.n1661 9.3005
R20316 vdd.n1663 vdd.n1603 9.3005
R20317 vdd.n1668 vdd.n1664 9.3005
R20318 vdd.n1669 vdd.n1599 9.3005
R20319 vdd.n1671 vdd.n1670 9.3005
R20320 vdd.n1672 vdd.n1598 9.3005
R20321 vdd.n1674 vdd.n1673 9.3005
R20322 vdd.n1675 vdd.n1593 9.3005
R20323 vdd.n1677 vdd.n1676 9.3005
R20324 vdd.n1678 vdd.n1592 9.3005
R20325 vdd.n1680 vdd.n1679 9.3005
R20326 vdd.n1681 vdd.n1587 9.3005
R20327 vdd.n1683 vdd.n1682 9.3005
R20328 vdd.n1684 vdd.n1586 9.3005
R20329 vdd.n1686 vdd.n1685 9.3005
R20330 vdd.n1687 vdd.n1581 9.3005
R20331 vdd.n1689 vdd.n1688 9.3005
R20332 vdd.n1690 vdd.n1580 9.3005
R20333 vdd.n1692 vdd.n1691 9.3005
R20334 vdd.n1693 vdd.n1575 9.3005
R20335 vdd.n1695 vdd.n1694 9.3005
R20336 vdd.n1696 vdd.n1574 9.3005
R20337 vdd.n1698 vdd.n1697 9.3005
R20338 vdd.n1699 vdd.n1571 9.3005
R20339 vdd.n1705 vdd.n1704 9.3005
R20340 vdd.n1706 vdd.n1570 9.3005
R20341 vdd.n1708 vdd.n1707 9.3005
R20342 vdd.n1709 vdd.n1565 9.3005
R20343 vdd.n1711 vdd.n1710 9.3005
R20344 vdd.n1712 vdd.n1564 9.3005
R20345 vdd.n1714 vdd.n1713 9.3005
R20346 vdd.n1715 vdd.n1559 9.3005
R20347 vdd.n1717 vdd.n1716 9.3005
R20348 vdd.n1718 vdd.n1558 9.3005
R20349 vdd.n1720 vdd.n1719 9.3005
R20350 vdd.n1721 vdd.n1553 9.3005
R20351 vdd.n1723 vdd.n1722 9.3005
R20352 vdd.n1724 vdd.n1552 9.3005
R20353 vdd.n1726 vdd.n1725 9.3005
R20354 vdd.n1727 vdd.n1548 9.3005
R20355 vdd.n1729 vdd.n1728 9.3005
R20356 vdd.n1730 vdd.n1547 9.3005
R20357 vdd.n1732 vdd.n1731 9.3005
R20358 vdd.n1733 vdd.n1546 9.3005
R20359 vdd.n1739 vdd.n1738 9.3005
R20360 vdd.n1747 vdd.n1746 9.3005
R20361 vdd.n1748 vdd.n1502 9.3005
R20362 vdd.n1750 vdd.n1749 9.3005
R20363 vdd.n1492 vdd.n1491 9.3005
R20364 vdd.n1764 vdd.n1763 9.3005
R20365 vdd.n1765 vdd.n1490 9.3005
R20366 vdd.n1767 vdd.n1766 9.3005
R20367 vdd.n1481 vdd.n1480 9.3005
R20368 vdd.n1781 vdd.n1780 9.3005
R20369 vdd.n1782 vdd.n1479 9.3005
R20370 vdd.n1784 vdd.n1783 9.3005
R20371 vdd.n1470 vdd.n1469 9.3005
R20372 vdd.n1797 vdd.n1796 9.3005
R20373 vdd.n1798 vdd.n1468 9.3005
R20374 vdd.n1800 vdd.n1799 9.3005
R20375 vdd.n1458 vdd.n1457 9.3005
R20376 vdd.n1814 vdd.n1813 9.3005
R20377 vdd.n1504 vdd.n1503 9.3005
R20378 vdd.n2026 vdd.n2025 9.3005
R20379 vdd.n2021 vdd.n2020 9.3005
R20380 vdd.n2032 vdd.n2031 9.3005
R20381 vdd.n2034 vdd.n2033 9.3005
R20382 vdd.n2017 vdd.n2016 9.3005
R20383 vdd.n2040 vdd.n2039 9.3005
R20384 vdd.n2042 vdd.n2041 9.3005
R20385 vdd.n2014 vdd.n2011 9.3005
R20386 vdd.n2049 vdd.n2048 9.3005
R20387 vdd.n2081 vdd.n2080 9.3005
R20388 vdd.n2076 vdd.n2075 9.3005
R20389 vdd.n2087 vdd.n2086 9.3005
R20390 vdd.n2089 vdd.n2088 9.3005
R20391 vdd.n2072 vdd.n2071 9.3005
R20392 vdd.n2095 vdd.n2094 9.3005
R20393 vdd.n2097 vdd.n2096 9.3005
R20394 vdd.n2069 vdd.n2066 9.3005
R20395 vdd.n2104 vdd.n2103 9.3005
R20396 vdd.n1928 vdd.n1927 9.3005
R20397 vdd.n1923 vdd.n1922 9.3005
R20398 vdd.n1934 vdd.n1933 9.3005
R20399 vdd.n1936 vdd.n1935 9.3005
R20400 vdd.n1919 vdd.n1918 9.3005
R20401 vdd.n1942 vdd.n1941 9.3005
R20402 vdd.n1944 vdd.n1943 9.3005
R20403 vdd.n1916 vdd.n1913 9.3005
R20404 vdd.n1951 vdd.n1950 9.3005
R20405 vdd.n1983 vdd.n1982 9.3005
R20406 vdd.n1978 vdd.n1977 9.3005
R20407 vdd.n1989 vdd.n1988 9.3005
R20408 vdd.n1991 vdd.n1990 9.3005
R20409 vdd.n1974 vdd.n1973 9.3005
R20410 vdd.n1997 vdd.n1996 9.3005
R20411 vdd.n1999 vdd.n1998 9.3005
R20412 vdd.n1971 vdd.n1968 9.3005
R20413 vdd.n2006 vdd.n2005 9.3005
R20414 vdd.n1831 vdd.n1830 9.3005
R20415 vdd.n1826 vdd.n1825 9.3005
R20416 vdd.n1837 vdd.n1836 9.3005
R20417 vdd.n1839 vdd.n1838 9.3005
R20418 vdd.n1822 vdd.n1821 9.3005
R20419 vdd.n1845 vdd.n1844 9.3005
R20420 vdd.n1847 vdd.n1846 9.3005
R20421 vdd.n1819 vdd.n1816 9.3005
R20422 vdd.n1854 vdd.n1853 9.3005
R20423 vdd.n1886 vdd.n1885 9.3005
R20424 vdd.n1881 vdd.n1880 9.3005
R20425 vdd.n1892 vdd.n1891 9.3005
R20426 vdd.n1894 vdd.n1893 9.3005
R20427 vdd.n1877 vdd.n1876 9.3005
R20428 vdd.n1900 vdd.n1899 9.3005
R20429 vdd.n1902 vdd.n1901 9.3005
R20430 vdd.n1874 vdd.n1871 9.3005
R20431 vdd.n1909 vdd.n1908 9.3005
R20432 vdd.n1760 vdd.t138 9.18308
R20433 vdd.n3328 vdd.t206 9.18308
R20434 vdd.n1786 vdd.t146 8.95635
R20435 vdd.t159 vdd.n3369 8.95635
R20436 vdd.n300 vdd.n299 8.92171
R20437 vdd.n245 vdd.n244 8.92171
R20438 vdd.n202 vdd.n201 8.92171
R20439 vdd.n147 vdd.n146 8.92171
R20440 vdd.n105 vdd.n104 8.92171
R20441 vdd.n50 vdd.n49 8.92171
R20442 vdd.n2031 vdd.n2030 8.92171
R20443 vdd.n2086 vdd.n2085 8.92171
R20444 vdd.n1933 vdd.n1932 8.92171
R20445 vdd.n1988 vdd.n1987 8.92171
R20446 vdd.n1836 vdd.n1835 8.92171
R20447 vdd.n1891 vdd.n1890 8.92171
R20448 vdd.n223 vdd.n125 8.81535
R20449 vdd.n2009 vdd.n1911 8.81535
R20450 vdd.n1466 vdd.t174 8.72962
R20451 vdd.t204 vdd.n3378 8.72962
R20452 vdd.n2122 vdd.t148 8.50289
R20453 vdd.n3297 vdd.t144 8.50289
R20454 vdd.n28 vdd.n14 8.42249
R20455 vdd.n2138 vdd.t199 8.27616
R20456 vdd.t136 vdd.n636 8.27616
R20457 vdd.n3384 vdd.n3383 8.16225
R20458 vdd.n2109 vdd.n2108 8.16225
R20459 vdd.n296 vdd.n290 8.14595
R20460 vdd.n241 vdd.n235 8.14595
R20461 vdd.n198 vdd.n192 8.14595
R20462 vdd.n143 vdd.n137 8.14595
R20463 vdd.n101 vdd.n95 8.14595
R20464 vdd.n46 vdd.n40 8.14595
R20465 vdd.n2027 vdd.n2021 8.14595
R20466 vdd.n2082 vdd.n2076 8.14595
R20467 vdd.n1929 vdd.n1923 8.14595
R20468 vdd.n1984 vdd.n1978 8.14595
R20469 vdd.n1832 vdd.n1826 8.14595
R20470 vdd.n1887 vdd.n1881 8.14595
R20471 vdd.t79 vdd.n1500 7.8227
R20472 vdd.t83 vdd.n363 7.8227
R20473 vdd.n2341 vdd.n1047 7.70933
R20474 vdd.n2341 vdd.n1050 7.70933
R20475 vdd.n2347 vdd.n1036 7.70933
R20476 vdd.n2353 vdd.n1036 7.70933
R20477 vdd.n2353 vdd.n1030 7.70933
R20478 vdd.n2359 vdd.n1030 7.70933
R20479 vdd.n2365 vdd.n1023 7.70933
R20480 vdd.n2365 vdd.n1026 7.70933
R20481 vdd.n2371 vdd.n1019 7.70933
R20482 vdd.n2378 vdd.n1005 7.70933
R20483 vdd.n2384 vdd.n1005 7.70933
R20484 vdd.n2390 vdd.n999 7.70933
R20485 vdd.n2396 vdd.n995 7.70933
R20486 vdd.n2402 vdd.n989 7.70933
R20487 vdd.n2414 vdd.n976 7.70933
R20488 vdd.n2420 vdd.n970 7.70933
R20489 vdd.n2420 vdd.n963 7.70933
R20490 vdd.n2428 vdd.n963 7.70933
R20491 vdd.n2510 vdd.n947 7.70933
R20492 vdd.n2862 vdd.n899 7.70933
R20493 vdd.n2874 vdd.n888 7.70933
R20494 vdd.n2874 vdd.n882 7.70933
R20495 vdd.n2880 vdd.n882 7.70933
R20496 vdd.n2886 vdd.n876 7.70933
R20497 vdd.n2892 vdd.n872 7.70933
R20498 vdd.n2898 vdd.n866 7.70933
R20499 vdd.n2910 vdd.n853 7.70933
R20500 vdd.n2916 vdd.n846 7.70933
R20501 vdd.n2916 vdd.n849 7.70933
R20502 vdd.n2923 vdd.n841 7.70933
R20503 vdd.n2929 vdd.n828 7.70933
R20504 vdd.n2935 vdd.n828 7.70933
R20505 vdd.n2941 vdd.n822 7.70933
R20506 vdd.n2941 vdd.n814 7.70933
R20507 vdd.n2992 vdd.n814 7.70933
R20508 vdd.n2992 vdd.n817 7.70933
R20509 vdd.n2998 vdd.n774 7.70933
R20510 vdd.n3068 vdd.n774 7.70933
R20511 vdd.n2921 vdd.n2920 7.49318
R20512 vdd.n2375 vdd.n2374 7.49318
R20513 vdd.n295 vdd.n292 7.3702
R20514 vdd.n240 vdd.n237 7.3702
R20515 vdd.n197 vdd.n194 7.3702
R20516 vdd.n142 vdd.n139 7.3702
R20517 vdd.n100 vdd.n97 7.3702
R20518 vdd.n45 vdd.n42 7.3702
R20519 vdd.n2026 vdd.n2023 7.3702
R20520 vdd.n2081 vdd.n2078 7.3702
R20521 vdd.n1928 vdd.n1925 7.3702
R20522 vdd.n1983 vdd.n1980 7.3702
R20523 vdd.n1831 vdd.n1828 7.3702
R20524 vdd.n1886 vdd.n1883 7.3702
R20525 vdd.n2359 vdd.t125 7.36923
R20526 vdd.t21 vdd.n822 7.36923
R20527 vdd.n2435 vdd.t17 7.25587
R20528 vdd.n2779 vdd.t47 7.25587
R20529 vdd.n1669 vdd.n1668 6.98232
R20530 vdd.n2225 vdd.n2224 6.98232
R20531 vdd.n547 vdd.n546 6.98232
R20532 vdd.n3152 vdd.n3151 6.98232
R20533 vdd.n2156 vdd.t140 6.91577
R20534 vdd.n3261 vdd.t234 6.91577
R20535 vdd.t218 vdd.n1437 6.68904
R20536 vdd.n3277 vdd.t187 6.68904
R20537 vdd.n2114 vdd.t156 6.46231
R20538 vdd.n3305 vdd.t154 6.46231
R20539 vdd.n3384 vdd.n321 6.32949
R20540 vdd.n2108 vdd.n2107 6.32949
R20541 vdd.t215 vdd.n1465 6.23558
R20542 vdd.t152 vdd.n332 6.23558
R20543 vdd.n1778 vdd.t170 6.00885
R20544 vdd.n3363 vdd.t150 6.00885
R20545 vdd.t32 vdd.n976 5.89549
R20546 vdd.n2886 vdd.t9 5.89549
R20547 vdd.n296 vdd.n295 5.81868
R20548 vdd.n241 vdd.n240 5.81868
R20549 vdd.n198 vdd.n197 5.81868
R20550 vdd.n143 vdd.n142 5.81868
R20551 vdd.n101 vdd.n100 5.81868
R20552 vdd.n46 vdd.n45 5.81868
R20553 vdd.n2027 vdd.n2026 5.81868
R20554 vdd.n2082 vdd.n2081 5.81868
R20555 vdd.n1929 vdd.n1928 5.81868
R20556 vdd.n1984 vdd.n1983 5.81868
R20557 vdd.n1832 vdd.n1831 5.81868
R20558 vdd.n1887 vdd.n1886 5.81868
R20559 vdd.n2518 vdd.n2517 5.77611
R20560 vdd.n1274 vdd.n1273 5.77611
R20561 vdd.n2791 vdd.n2790 5.77611
R20562 vdd.n3007 vdd.n806 5.77611
R20563 vdd.n3073 vdd.n770 5.77611
R20564 vdd.n2685 vdd.n2623 5.77611
R20565 vdd.n2443 vdd.n954 5.77611
R20566 vdd.n1363 vdd.n1226 5.77611
R20567 vdd.n1738 vdd.n1512 5.62474
R20568 vdd.n2188 vdd.n2185 5.62474
R20569 vdd.n3342 vdd.n407 5.62474
R20570 vdd.n3107 vdd.n3104 5.62474
R20571 vdd.t35 vdd.n999 5.55539
R20572 vdd.n2390 vdd.t5 5.55539
R20573 vdd.t14 vdd.n853 5.55539
R20574 vdd.n2910 vdd.t126 5.55539
R20575 vdd.n1019 vdd.t104 5.44203
R20576 vdd.n2923 vdd.t72 5.44203
R20577 vdd.n1488 vdd.t170 5.32866
R20578 vdd.n2347 vdd.t54 5.32866
R20579 vdd.n1309 vdd.t96 5.32866
R20580 vdd.n2868 vdd.t100 5.32866
R20581 vdd.n817 vdd.t50 5.32866
R20582 vdd.t150 vdd.n3362 5.32866
R20583 vdd.n1794 vdd.t215 5.10193
R20584 vdd.n3371 vdd.t152 5.10193
R20585 vdd.n299 vdd.n290 5.04292
R20586 vdd.n244 vdd.n235 5.04292
R20587 vdd.n201 vdd.n192 5.04292
R20588 vdd.n146 vdd.n137 5.04292
R20589 vdd.n104 vdd.n95 5.04292
R20590 vdd.n49 vdd.n40 5.04292
R20591 vdd.n2030 vdd.n2021 5.04292
R20592 vdd.n2085 vdd.n2076 5.04292
R20593 vdd.n1932 vdd.n1923 5.04292
R20594 vdd.n1987 vdd.n1978 5.04292
R20595 vdd.n1835 vdd.n1826 5.04292
R20596 vdd.n1890 vdd.n1881 5.04292
R20597 vdd.n2396 vdd.t11 4.98857
R20598 vdd.n866 vdd.t264 4.98857
R20599 vdd.n1810 vdd.t156 4.8752
R20600 vdd.t44 vdd.t129 4.8752
R20601 vdd.t22 vdd.t45 4.8752
R20602 vdd.t134 vdd.t8 4.8752
R20603 vdd.t15 vdd.t40 4.8752
R20604 vdd.t154 vdd.n328 4.8752
R20605 vdd.n2519 vdd.n2518 4.83952
R20606 vdd.n1273 vdd.n1272 4.83952
R20607 vdd.n2792 vdd.n2791 4.83952
R20608 vdd.n806 vdd.n801 4.83952
R20609 vdd.n770 vdd.n765 4.83952
R20610 vdd.n2682 vdd.n2623 4.83952
R20611 vdd.n2446 vdd.n954 4.83952
R20612 vdd.n1366 vdd.n1226 4.83952
R20613 vdd.n2193 vdd.n2192 4.74817
R20614 vdd.n1399 vdd.n1394 4.74817
R20615 vdd.n1096 vdd.n1093 4.74817
R20616 vdd.n2286 vdd.n1092 4.74817
R20617 vdd.n2291 vdd.n1093 4.74817
R20618 vdd.n2290 vdd.n1092 4.74817
R20619 vdd.n664 vdd.n662 4.74817
R20620 vdd.n3222 vdd.n665 4.74817
R20621 vdd.n3225 vdd.n665 4.74817
R20622 vdd.n3226 vdd.n664 4.74817
R20623 vdd.n3114 vdd.n749 4.74817
R20624 vdd.n3110 vdd.n751 4.74817
R20625 vdd.n3113 vdd.n751 4.74817
R20626 vdd.n3118 vdd.n749 4.74817
R20627 vdd.n2192 vdd.n1192 4.74817
R20628 vdd.n1396 vdd.n1394 4.74817
R20629 vdd.n321 vdd.n320 4.7074
R20630 vdd.n223 vdd.n222 4.7074
R20631 vdd.n2107 vdd.n2106 4.7074
R20632 vdd.n2009 vdd.n2008 4.7074
R20633 vdd.n2130 vdd.t218 4.64847
R20634 vdd.n2371 vdd.t13 4.64847
R20635 vdd.n989 vdd.t131 4.64847
R20636 vdd.n2892 vdd.t37 4.64847
R20637 vdd.n841 vdd.t41 4.64847
R20638 vdd.n3286 vdd.t187 4.64847
R20639 vdd.n1431 vdd.t140 4.42174
R20640 vdd.t234 vdd.n635 4.42174
R20641 vdd.n300 vdd.n288 4.26717
R20642 vdd.n245 vdd.n233 4.26717
R20643 vdd.n202 vdd.n190 4.26717
R20644 vdd.n147 vdd.n135 4.26717
R20645 vdd.n105 vdd.n93 4.26717
R20646 vdd.n50 vdd.n38 4.26717
R20647 vdd.n2031 vdd.n2019 4.26717
R20648 vdd.n2086 vdd.n2074 4.26717
R20649 vdd.n1933 vdd.n1921 4.26717
R20650 vdd.n1988 vdd.n1976 4.26717
R20651 vdd.n1836 vdd.n1824 4.26717
R20652 vdd.n1891 vdd.n1879 4.26717
R20653 vdd.n321 vdd.n223 4.10845
R20654 vdd.n2107 vdd.n2009 4.10845
R20655 vdd.n277 vdd.t162 4.06363
R20656 vdd.n277 vdd.t222 4.06363
R20657 vdd.n275 vdd.t248 4.06363
R20658 vdd.n275 vdd.t256 4.06363
R20659 vdd.n273 vdd.t260 4.06363
R20660 vdd.n273 vdd.t176 4.06363
R20661 vdd.n271 vdd.t201 4.06363
R20662 vdd.n271 vdd.t259 4.06363
R20663 vdd.n269 vdd.t261 4.06363
R20664 vdd.n269 vdd.t198 4.06363
R20665 vdd.n267 vdd.t203 4.06363
R20666 vdd.n267 vdd.t209 4.06363
R20667 vdd.n265 vdd.t242 4.06363
R20668 vdd.n265 vdd.t158 4.06363
R20669 vdd.n179 vdd.t151 4.06363
R20670 vdd.n179 vdd.t207 4.06363
R20671 vdd.n177 vdd.t236 4.06363
R20672 vdd.n177 vdd.t244 4.06363
R20673 vdd.n175 vdd.t252 4.06363
R20674 vdd.n175 vdd.t153 4.06363
R20675 vdd.n173 vdd.t182 4.06363
R20676 vdd.n173 vdd.t251 4.06363
R20677 vdd.n171 vdd.t253 4.06363
R20678 vdd.n171 vdd.t181 4.06363
R20679 vdd.n169 vdd.t186 4.06363
R20680 vdd.n169 vdd.t188 4.06363
R20681 vdd.n167 vdd.t235 4.06363
R20682 vdd.n167 vdd.t137 4.06363
R20683 vdd.n82 vdd.t164 4.06363
R20684 vdd.n82 vdd.t241 4.06363
R20685 vdd.n80 vdd.t160 4.06363
R20686 vdd.n80 vdd.t229 4.06363
R20687 vdd.n78 vdd.t184 4.06363
R20688 vdd.n78 vdd.t249 4.06363
R20689 vdd.n76 vdd.t155 4.06363
R20690 vdd.n76 vdd.t205 4.06363
R20691 vdd.n74 vdd.t145 4.06363
R20692 vdd.n74 vdd.t189 4.06363
R20693 vdd.n72 vdd.t257 4.06363
R20694 vdd.n72 vdd.t240 4.06363
R20695 vdd.n70 vdd.t245 4.06363
R20696 vdd.n70 vdd.t202 4.06363
R20697 vdd.n2051 vdd.t217 4.06363
R20698 vdd.n2051 vdd.t165 4.06363
R20699 vdd.n2053 vdd.t263 4.06363
R20700 vdd.n2053 vdd.t239 4.06363
R20701 vdd.n2055 vdd.t237 4.06363
R20702 vdd.n2055 vdd.t197 4.06363
R20703 vdd.n2057 vdd.t193 4.06363
R20704 vdd.n2057 vdd.t238 4.06363
R20705 vdd.n2059 vdd.t225 4.06363
R20706 vdd.n2059 vdd.t224 4.06363
R20707 vdd.n2061 vdd.t190 4.06363
R20708 vdd.n2061 vdd.t167 4.06363
R20709 vdd.n2063 vdd.t163 4.06363
R20710 vdd.n2063 vdd.t223 4.06363
R20711 vdd.n1953 vdd.t208 4.06363
R20712 vdd.n1953 vdd.t141 4.06363
R20713 vdd.n1955 vdd.t255 4.06363
R20714 vdd.n1955 vdd.t232 4.06363
R20715 vdd.n1957 vdd.t226 4.06363
R20716 vdd.n1957 vdd.t179 4.06363
R20717 vdd.n1959 vdd.t175 4.06363
R20718 vdd.n1959 vdd.t227 4.06363
R20719 vdd.n1961 vdd.t216 4.06363
R20720 vdd.n1961 vdd.t214 4.06363
R20721 vdd.n1963 vdd.t169 4.06363
R20722 vdd.n1963 vdd.t147 4.06363
R20723 vdd.n1965 vdd.t139 4.06363
R20724 vdd.n1965 vdd.t212 4.06363
R20725 vdd.n1856 vdd.t200 4.06363
R20726 vdd.n1856 vdd.t247 4.06363
R20727 vdd.n1858 vdd.t219 4.06363
R20728 vdd.n1858 vdd.t258 4.06363
R20729 vdd.n1860 vdd.t192 4.06363
R20730 vdd.n1860 vdd.t149 4.06363
R20731 vdd.n1862 vdd.t211 4.06363
R20732 vdd.n1862 vdd.t157 4.06363
R20733 vdd.n1864 vdd.t250 4.06363
R20734 vdd.n1864 vdd.t262 4.06363
R20735 vdd.n1866 vdd.t230 4.06363
R20736 vdd.n1866 vdd.t161 4.06363
R20737 vdd.n1868 vdd.t221 4.06363
R20738 vdd.n1868 vdd.t171 4.06363
R20739 vdd.n26 vdd.t7 3.9605
R20740 vdd.n26 vdd.t0 3.9605
R20741 vdd.n23 vdd.t24 3.9605
R20742 vdd.n23 vdd.t27 3.9605
R20743 vdd.n21 vdd.t4 3.9605
R20744 vdd.n21 vdd.t2 3.9605
R20745 vdd.n20 vdd.t29 3.9605
R20746 vdd.n20 vdd.t31 3.9605
R20747 vdd.n15 vdd.t3 3.9605
R20748 vdd.n15 vdd.t30 3.9605
R20749 vdd.n16 vdd.t1 3.9605
R20750 vdd.n16 vdd.t28 3.9605
R20751 vdd.n18 vdd.t26 3.9605
R20752 vdd.n18 vdd.t25 3.9605
R20753 vdd.n25 vdd.t6 3.9605
R20754 vdd.n25 vdd.t23 3.9605
R20755 vdd.n2428 vdd.t127 3.85492
R20756 vdd.n1309 vdd.t127 3.85492
R20757 vdd.n2868 vdd.t42 3.85492
R20758 vdd.t42 vdd.n888 3.85492
R20759 vdd.n7 vdd.t16 3.61217
R20760 vdd.n7 vdd.t265 3.61217
R20761 vdd.n8 vdd.t135 3.61217
R20762 vdd.n8 vdd.t10 3.61217
R20763 vdd.n10 vdd.t48 3.61217
R20764 vdd.n10 vdd.t43 3.61217
R20765 vdd.n12 vdd.t267 3.61217
R20766 vdd.n12 vdd.t39 3.61217
R20767 vdd.n5 vdd.t20 3.61217
R20768 vdd.n5 vdd.t133 3.61217
R20769 vdd.n3 vdd.t128 3.61217
R20770 vdd.n3 vdd.t18 3.61217
R20771 vdd.n1 vdd.t33 3.61217
R20772 vdd.n1 vdd.t46 3.61217
R20773 vdd.n0 vdd.t12 3.61217
R20774 vdd.n0 vdd.t130 3.61217
R20775 vdd.n1744 vdd.t79 3.51482
R20776 vdd.n3347 vdd.t83 3.51482
R20777 vdd.n304 vdd.n303 3.49141
R20778 vdd.n249 vdd.n248 3.49141
R20779 vdd.n206 vdd.n205 3.49141
R20780 vdd.n151 vdd.n150 3.49141
R20781 vdd.n109 vdd.n108 3.49141
R20782 vdd.n54 vdd.n53 3.49141
R20783 vdd.n2035 vdd.n2034 3.49141
R20784 vdd.n2090 vdd.n2089 3.49141
R20785 vdd.n1937 vdd.n1936 3.49141
R20786 vdd.n1992 vdd.n1991 3.49141
R20787 vdd.n1840 vdd.n1839 3.49141
R20788 vdd.n1895 vdd.n1894 3.49141
R20789 vdd.n2582 vdd.t19 3.40145
R20790 vdd.n2855 vdd.t38 3.40145
R20791 vdd.n2920 vdd.n2919 3.12245
R20792 vdd.n2376 vdd.n2375 3.12245
R20793 vdd.n2147 vdd.t199 3.06136
R20794 vdd.n1026 vdd.t13 3.06136
R20795 vdd.n2408 vdd.t131 3.06136
R20796 vdd.n2764 vdd.t37 3.06136
R20797 vdd.n2929 vdd.t41 3.06136
R20798 vdd.n3269 vdd.t136 3.06136
R20799 vdd.t148 vdd.n1443 2.83463
R20800 vdd.n624 vdd.t144 2.83463
R20801 vdd.n1330 vdd.t11 2.72126
R20802 vdd.n2904 vdd.t264 2.72126
R20803 vdd.n307 vdd.n286 2.71565
R20804 vdd.n252 vdd.n231 2.71565
R20805 vdd.n209 vdd.n188 2.71565
R20806 vdd.n154 vdd.n133 2.71565
R20807 vdd.n112 vdd.n91 2.71565
R20808 vdd.n57 vdd.n36 2.71565
R20809 vdd.n2038 vdd.n2017 2.71565
R20810 vdd.n2093 vdd.n2072 2.71565
R20811 vdd.n1940 vdd.n1919 2.71565
R20812 vdd.n1995 vdd.n1974 2.71565
R20813 vdd.n1843 vdd.n1822 2.71565
R20814 vdd.n1898 vdd.n1877 2.71565
R20815 vdd.n1811 vdd.t174 2.6079
R20816 vdd.n3379 vdd.t204 2.6079
R20817 vdd.t45 vdd.n970 2.49453
R20818 vdd.n2880 vdd.t134 2.49453
R20819 vdd.n294 vdd.n293 2.4129
R20820 vdd.n239 vdd.n238 2.4129
R20821 vdd.n196 vdd.n195 2.4129
R20822 vdd.n141 vdd.n140 2.4129
R20823 vdd.n99 vdd.n98 2.4129
R20824 vdd.n44 vdd.n43 2.4129
R20825 vdd.n2025 vdd.n2024 2.4129
R20826 vdd.n2080 vdd.n2079 2.4129
R20827 vdd.n1927 vdd.n1926 2.4129
R20828 vdd.n1982 vdd.n1981 2.4129
R20829 vdd.n1830 vdd.n1829 2.4129
R20830 vdd.n1885 vdd.n1884 2.4129
R20831 vdd.t146 vdd.n1472 2.38117
R20832 vdd.n1050 vdd.t54 2.38117
R20833 vdd.n2435 vdd.t96 2.38117
R20834 vdd.n2779 vdd.t100 2.38117
R20835 vdd.n2998 vdd.t50 2.38117
R20836 vdd.n3370 vdd.t159 2.38117
R20837 vdd.n2298 vdd.n1093 2.27742
R20838 vdd.n2298 vdd.n1092 2.27742
R20839 vdd.n3034 vdd.n665 2.27742
R20840 vdd.n3034 vdd.n664 2.27742
R20841 vdd.n3102 vdd.n751 2.27742
R20842 vdd.n3102 vdd.n749 2.27742
R20843 vdd.n2192 vdd.n2191 2.27742
R20844 vdd.n2191 vdd.n1394 2.27742
R20845 vdd.n1769 vdd.t138 2.15444
R20846 vdd.n2384 vdd.t35 2.15444
R20847 vdd.n1330 vdd.t5 2.15444
R20848 vdd.n2904 vdd.t14 2.15444
R20849 vdd.t126 vdd.n846 2.15444
R20850 vdd.n3361 vdd.t206 2.15444
R20851 vdd.n308 vdd.n284 1.93989
R20852 vdd.n253 vdd.n229 1.93989
R20853 vdd.n210 vdd.n186 1.93989
R20854 vdd.n155 vdd.n131 1.93989
R20855 vdd.n113 vdd.n89 1.93989
R20856 vdd.n58 vdd.n34 1.93989
R20857 vdd.n2039 vdd.n2015 1.93989
R20858 vdd.n2094 vdd.n2070 1.93989
R20859 vdd.n1941 vdd.n1917 1.93989
R20860 vdd.n1996 vdd.n1972 1.93989
R20861 vdd.n1844 vdd.n1820 1.93989
R20862 vdd.n1899 vdd.n1875 1.93989
R20863 vdd.n2408 vdd.t32 1.81434
R20864 vdd.n2764 vdd.t9 1.81434
R20865 vdd.n1761 vdd.t142 1.70098
R20866 vdd.n3355 vdd.t194 1.70098
R20867 vdd.n2402 vdd.t129 1.58761
R20868 vdd.n872 vdd.t15 1.58761
R20869 vdd.n1777 vdd.t168 1.47425
R20870 vdd.n349 vdd.t228 1.47425
R20871 vdd.n1802 vdd.t213 1.24752
R20872 vdd.t62 vdd.n1407 1.24752
R20873 vdd.n2378 vdd.t36 1.24752
R20874 vdd.n995 vdd.t44 1.24752
R20875 vdd.n2898 vdd.t40 1.24752
R20876 vdd.n849 vdd.t34 1.24752
R20877 vdd.n659 vdd.t58 1.24752
R20878 vdd.t183 vdd.n3377 1.24752
R20879 vdd.n319 vdd.n279 1.16414
R20880 vdd.n312 vdd.n311 1.16414
R20881 vdd.n264 vdd.n224 1.16414
R20882 vdd.n257 vdd.n256 1.16414
R20883 vdd.n221 vdd.n181 1.16414
R20884 vdd.n214 vdd.n213 1.16414
R20885 vdd.n166 vdd.n126 1.16414
R20886 vdd.n159 vdd.n158 1.16414
R20887 vdd.n124 vdd.n84 1.16414
R20888 vdd.n117 vdd.n116 1.16414
R20889 vdd.n69 vdd.n29 1.16414
R20890 vdd.n62 vdd.n61 1.16414
R20891 vdd.n2050 vdd.n2010 1.16414
R20892 vdd.n2043 vdd.n2042 1.16414
R20893 vdd.n2105 vdd.n2065 1.16414
R20894 vdd.n2098 vdd.n2097 1.16414
R20895 vdd.n1952 vdd.n1912 1.16414
R20896 vdd.n1945 vdd.n1944 1.16414
R20897 vdd.n2007 vdd.n1967 1.16414
R20898 vdd.n2000 vdd.n1999 1.16414
R20899 vdd.n1855 vdd.n1815 1.16414
R20900 vdd.n1848 vdd.n1847 1.16414
R20901 vdd.n1910 vdd.n1870 1.16414
R20902 vdd.n1903 vdd.n1902 1.16414
R20903 vdd.n1454 vdd.t191 1.02079
R20904 vdd.t104 vdd.t36 1.02079
R20905 vdd.t34 vdd.t72 1.02079
R20906 vdd.t180 vdd.n613 1.02079
R20907 vdd.n1633 vdd.n1512 0.970197
R20908 vdd.n2189 vdd.n2188 0.970197
R20909 vdd.n599 vdd.n407 0.970197
R20910 vdd.n3109 vdd.n3107 0.970197
R20911 vdd.n2108 vdd.n28 0.956323
R20912 vdd vdd.n3384 0.94849
R20913 vdd.n2139 vdd.t231 0.794056
R20914 vdd.n3278 vdd.t185 0.794056
R20915 vdd.n2155 vdd.t172 0.567326
R20916 vdd.t177 vdd.n642 0.567326
R20917 vdd.n2179 vdd.n1094 0.482207
R20918 vdd.n3234 vdd.n3233 0.482207
R20919 vdd.n444 vdd.n443 0.482207
R20920 vdd.n3341 vdd.n3340 0.482207
R20921 vdd.n3240 vdd.n656 0.482207
R20922 vdd.n2169 vdd.n1395 0.482207
R20923 vdd.n1740 vdd.n1739 0.482207
R20924 vdd.n1546 vdd.n1503 0.482207
R20925 vdd.n4 vdd.n2 0.459552
R20926 vdd.n11 vdd.n9 0.459552
R20927 vdd.t17 vdd.n947 0.453961
R20928 vdd.n2862 vdd.t47 0.453961
R20929 vdd.n317 vdd.n316 0.388379
R20930 vdd.n283 vdd.n281 0.388379
R20931 vdd.n262 vdd.n261 0.388379
R20932 vdd.n228 vdd.n226 0.388379
R20933 vdd.n219 vdd.n218 0.388379
R20934 vdd.n185 vdd.n183 0.388379
R20935 vdd.n164 vdd.n163 0.388379
R20936 vdd.n130 vdd.n128 0.388379
R20937 vdd.n122 vdd.n121 0.388379
R20938 vdd.n88 vdd.n86 0.388379
R20939 vdd.n67 vdd.n66 0.388379
R20940 vdd.n33 vdd.n31 0.388379
R20941 vdd.n2048 vdd.n2047 0.388379
R20942 vdd.n2014 vdd.n2012 0.388379
R20943 vdd.n2103 vdd.n2102 0.388379
R20944 vdd.n2069 vdd.n2067 0.388379
R20945 vdd.n1950 vdd.n1949 0.388379
R20946 vdd.n1916 vdd.n1914 0.388379
R20947 vdd.n2005 vdd.n2004 0.388379
R20948 vdd.n1971 vdd.n1969 0.388379
R20949 vdd.n1853 vdd.n1852 0.388379
R20950 vdd.n1819 vdd.n1817 0.388379
R20951 vdd.n1908 vdd.n1907 0.388379
R20952 vdd.n1874 vdd.n1872 0.388379
R20953 vdd.n19 vdd.n17 0.387128
R20954 vdd.n24 vdd.n22 0.387128
R20955 vdd.n6 vdd.n4 0.358259
R20956 vdd.n13 vdd.n11 0.358259
R20957 vdd.n268 vdd.n266 0.358259
R20958 vdd.n270 vdd.n268 0.358259
R20959 vdd.n272 vdd.n270 0.358259
R20960 vdd.n274 vdd.n272 0.358259
R20961 vdd.n276 vdd.n274 0.358259
R20962 vdd.n278 vdd.n276 0.358259
R20963 vdd.n320 vdd.n278 0.358259
R20964 vdd.n170 vdd.n168 0.358259
R20965 vdd.n172 vdd.n170 0.358259
R20966 vdd.n174 vdd.n172 0.358259
R20967 vdd.n176 vdd.n174 0.358259
R20968 vdd.n178 vdd.n176 0.358259
R20969 vdd.n180 vdd.n178 0.358259
R20970 vdd.n222 vdd.n180 0.358259
R20971 vdd.n73 vdd.n71 0.358259
R20972 vdd.n75 vdd.n73 0.358259
R20973 vdd.n77 vdd.n75 0.358259
R20974 vdd.n79 vdd.n77 0.358259
R20975 vdd.n81 vdd.n79 0.358259
R20976 vdd.n83 vdd.n81 0.358259
R20977 vdd.n125 vdd.n83 0.358259
R20978 vdd.n2106 vdd.n2064 0.358259
R20979 vdd.n2064 vdd.n2062 0.358259
R20980 vdd.n2062 vdd.n2060 0.358259
R20981 vdd.n2060 vdd.n2058 0.358259
R20982 vdd.n2058 vdd.n2056 0.358259
R20983 vdd.n2056 vdd.n2054 0.358259
R20984 vdd.n2054 vdd.n2052 0.358259
R20985 vdd.n2008 vdd.n1966 0.358259
R20986 vdd.n1966 vdd.n1964 0.358259
R20987 vdd.n1964 vdd.n1962 0.358259
R20988 vdd.n1962 vdd.n1960 0.358259
R20989 vdd.n1960 vdd.n1958 0.358259
R20990 vdd.n1958 vdd.n1956 0.358259
R20991 vdd.n1956 vdd.n1954 0.358259
R20992 vdd.n1911 vdd.n1869 0.358259
R20993 vdd.n1869 vdd.n1867 0.358259
R20994 vdd.n1867 vdd.n1865 0.358259
R20995 vdd.n1865 vdd.n1863 0.358259
R20996 vdd.n1863 vdd.n1861 0.358259
R20997 vdd.n1861 vdd.n1859 0.358259
R20998 vdd.n1859 vdd.n1857 0.358259
R20999 vdd.t125 vdd.n1023 0.340595
R21000 vdd.n2414 vdd.t22 0.340595
R21001 vdd.t8 vdd.n876 0.340595
R21002 vdd.n2935 vdd.t21 0.340595
R21003 vdd.n14 vdd.n6 0.334552
R21004 vdd.n14 vdd.n13 0.334552
R21005 vdd.n27 vdd.n19 0.21707
R21006 vdd.n27 vdd.n24 0.21707
R21007 vdd.n318 vdd.n280 0.155672
R21008 vdd.n310 vdd.n280 0.155672
R21009 vdd.n310 vdd.n309 0.155672
R21010 vdd.n309 vdd.n285 0.155672
R21011 vdd.n302 vdd.n285 0.155672
R21012 vdd.n302 vdd.n301 0.155672
R21013 vdd.n301 vdd.n289 0.155672
R21014 vdd.n294 vdd.n289 0.155672
R21015 vdd.n263 vdd.n225 0.155672
R21016 vdd.n255 vdd.n225 0.155672
R21017 vdd.n255 vdd.n254 0.155672
R21018 vdd.n254 vdd.n230 0.155672
R21019 vdd.n247 vdd.n230 0.155672
R21020 vdd.n247 vdd.n246 0.155672
R21021 vdd.n246 vdd.n234 0.155672
R21022 vdd.n239 vdd.n234 0.155672
R21023 vdd.n220 vdd.n182 0.155672
R21024 vdd.n212 vdd.n182 0.155672
R21025 vdd.n212 vdd.n211 0.155672
R21026 vdd.n211 vdd.n187 0.155672
R21027 vdd.n204 vdd.n187 0.155672
R21028 vdd.n204 vdd.n203 0.155672
R21029 vdd.n203 vdd.n191 0.155672
R21030 vdd.n196 vdd.n191 0.155672
R21031 vdd.n165 vdd.n127 0.155672
R21032 vdd.n157 vdd.n127 0.155672
R21033 vdd.n157 vdd.n156 0.155672
R21034 vdd.n156 vdd.n132 0.155672
R21035 vdd.n149 vdd.n132 0.155672
R21036 vdd.n149 vdd.n148 0.155672
R21037 vdd.n148 vdd.n136 0.155672
R21038 vdd.n141 vdd.n136 0.155672
R21039 vdd.n123 vdd.n85 0.155672
R21040 vdd.n115 vdd.n85 0.155672
R21041 vdd.n115 vdd.n114 0.155672
R21042 vdd.n114 vdd.n90 0.155672
R21043 vdd.n107 vdd.n90 0.155672
R21044 vdd.n107 vdd.n106 0.155672
R21045 vdd.n106 vdd.n94 0.155672
R21046 vdd.n99 vdd.n94 0.155672
R21047 vdd.n68 vdd.n30 0.155672
R21048 vdd.n60 vdd.n30 0.155672
R21049 vdd.n60 vdd.n59 0.155672
R21050 vdd.n59 vdd.n35 0.155672
R21051 vdd.n52 vdd.n35 0.155672
R21052 vdd.n52 vdd.n51 0.155672
R21053 vdd.n51 vdd.n39 0.155672
R21054 vdd.n44 vdd.n39 0.155672
R21055 vdd.n2049 vdd.n2011 0.155672
R21056 vdd.n2041 vdd.n2011 0.155672
R21057 vdd.n2041 vdd.n2040 0.155672
R21058 vdd.n2040 vdd.n2016 0.155672
R21059 vdd.n2033 vdd.n2016 0.155672
R21060 vdd.n2033 vdd.n2032 0.155672
R21061 vdd.n2032 vdd.n2020 0.155672
R21062 vdd.n2025 vdd.n2020 0.155672
R21063 vdd.n2104 vdd.n2066 0.155672
R21064 vdd.n2096 vdd.n2066 0.155672
R21065 vdd.n2096 vdd.n2095 0.155672
R21066 vdd.n2095 vdd.n2071 0.155672
R21067 vdd.n2088 vdd.n2071 0.155672
R21068 vdd.n2088 vdd.n2087 0.155672
R21069 vdd.n2087 vdd.n2075 0.155672
R21070 vdd.n2080 vdd.n2075 0.155672
R21071 vdd.n1951 vdd.n1913 0.155672
R21072 vdd.n1943 vdd.n1913 0.155672
R21073 vdd.n1943 vdd.n1942 0.155672
R21074 vdd.n1942 vdd.n1918 0.155672
R21075 vdd.n1935 vdd.n1918 0.155672
R21076 vdd.n1935 vdd.n1934 0.155672
R21077 vdd.n1934 vdd.n1922 0.155672
R21078 vdd.n1927 vdd.n1922 0.155672
R21079 vdd.n2006 vdd.n1968 0.155672
R21080 vdd.n1998 vdd.n1968 0.155672
R21081 vdd.n1998 vdd.n1997 0.155672
R21082 vdd.n1997 vdd.n1973 0.155672
R21083 vdd.n1990 vdd.n1973 0.155672
R21084 vdd.n1990 vdd.n1989 0.155672
R21085 vdd.n1989 vdd.n1977 0.155672
R21086 vdd.n1982 vdd.n1977 0.155672
R21087 vdd.n1854 vdd.n1816 0.155672
R21088 vdd.n1846 vdd.n1816 0.155672
R21089 vdd.n1846 vdd.n1845 0.155672
R21090 vdd.n1845 vdd.n1821 0.155672
R21091 vdd.n1838 vdd.n1821 0.155672
R21092 vdd.n1838 vdd.n1837 0.155672
R21093 vdd.n1837 vdd.n1825 0.155672
R21094 vdd.n1830 vdd.n1825 0.155672
R21095 vdd.n1909 vdd.n1871 0.155672
R21096 vdd.n1901 vdd.n1871 0.155672
R21097 vdd.n1901 vdd.n1900 0.155672
R21098 vdd.n1900 vdd.n1876 0.155672
R21099 vdd.n1893 vdd.n1876 0.155672
R21100 vdd.n1893 vdd.n1892 0.155672
R21101 vdd.n1892 vdd.n1880 0.155672
R21102 vdd.n1885 vdd.n1880 0.155672
R21103 vdd.n1099 vdd.n1091 0.152939
R21104 vdd.n1103 vdd.n1099 0.152939
R21105 vdd.n1104 vdd.n1103 0.152939
R21106 vdd.n1105 vdd.n1104 0.152939
R21107 vdd.n1106 vdd.n1105 0.152939
R21108 vdd.n1110 vdd.n1106 0.152939
R21109 vdd.n1111 vdd.n1110 0.152939
R21110 vdd.n1112 vdd.n1111 0.152939
R21111 vdd.n1113 vdd.n1112 0.152939
R21112 vdd.n1117 vdd.n1113 0.152939
R21113 vdd.n1118 vdd.n1117 0.152939
R21114 vdd.n1119 vdd.n1118 0.152939
R21115 vdd.n2262 vdd.n1119 0.152939
R21116 vdd.n2262 vdd.n2261 0.152939
R21117 vdd.n2261 vdd.n2260 0.152939
R21118 vdd.n2260 vdd.n1125 0.152939
R21119 vdd.n1130 vdd.n1125 0.152939
R21120 vdd.n1131 vdd.n1130 0.152939
R21121 vdd.n1132 vdd.n1131 0.152939
R21122 vdd.n1136 vdd.n1132 0.152939
R21123 vdd.n1137 vdd.n1136 0.152939
R21124 vdd.n1138 vdd.n1137 0.152939
R21125 vdd.n1139 vdd.n1138 0.152939
R21126 vdd.n1143 vdd.n1139 0.152939
R21127 vdd.n1144 vdd.n1143 0.152939
R21128 vdd.n1145 vdd.n1144 0.152939
R21129 vdd.n1146 vdd.n1145 0.152939
R21130 vdd.n1150 vdd.n1146 0.152939
R21131 vdd.n1151 vdd.n1150 0.152939
R21132 vdd.n1152 vdd.n1151 0.152939
R21133 vdd.n1153 vdd.n1152 0.152939
R21134 vdd.n1157 vdd.n1153 0.152939
R21135 vdd.n1158 vdd.n1157 0.152939
R21136 vdd.n1159 vdd.n1158 0.152939
R21137 vdd.n2223 vdd.n1159 0.152939
R21138 vdd.n2223 vdd.n2222 0.152939
R21139 vdd.n2222 vdd.n2221 0.152939
R21140 vdd.n2221 vdd.n1165 0.152939
R21141 vdd.n1170 vdd.n1165 0.152939
R21142 vdd.n1171 vdd.n1170 0.152939
R21143 vdd.n1172 vdd.n1171 0.152939
R21144 vdd.n1176 vdd.n1172 0.152939
R21145 vdd.n1177 vdd.n1176 0.152939
R21146 vdd.n1178 vdd.n1177 0.152939
R21147 vdd.n1179 vdd.n1178 0.152939
R21148 vdd.n1183 vdd.n1179 0.152939
R21149 vdd.n1184 vdd.n1183 0.152939
R21150 vdd.n1185 vdd.n1184 0.152939
R21151 vdd.n1186 vdd.n1185 0.152939
R21152 vdd.n1190 vdd.n1186 0.152939
R21153 vdd.n1191 vdd.n1190 0.152939
R21154 vdd.n2297 vdd.n1094 0.152939
R21155 vdd.n2111 vdd.n2110 0.152939
R21156 vdd.n2111 vdd.n1446 0.152939
R21157 vdd.n2125 vdd.n1446 0.152939
R21158 vdd.n2126 vdd.n2125 0.152939
R21159 vdd.n2127 vdd.n2126 0.152939
R21160 vdd.n2127 vdd.n1434 0.152939
R21161 vdd.n2142 vdd.n1434 0.152939
R21162 vdd.n2143 vdd.n2142 0.152939
R21163 vdd.n2144 vdd.n2143 0.152939
R21164 vdd.n2144 vdd.n1423 0.152939
R21165 vdd.n2159 vdd.n1423 0.152939
R21166 vdd.n2160 vdd.n2159 0.152939
R21167 vdd.n2161 vdd.n2160 0.152939
R21168 vdd.n2161 vdd.n1411 0.152939
R21169 vdd.n2177 vdd.n1411 0.152939
R21170 vdd.n2178 vdd.n2177 0.152939
R21171 vdd.n2179 vdd.n2178 0.152939
R21172 vdd.n670 vdd.n667 0.152939
R21173 vdd.n671 vdd.n670 0.152939
R21174 vdd.n672 vdd.n671 0.152939
R21175 vdd.n673 vdd.n672 0.152939
R21176 vdd.n676 vdd.n673 0.152939
R21177 vdd.n677 vdd.n676 0.152939
R21178 vdd.n678 vdd.n677 0.152939
R21179 vdd.n679 vdd.n678 0.152939
R21180 vdd.n682 vdd.n679 0.152939
R21181 vdd.n683 vdd.n682 0.152939
R21182 vdd.n684 vdd.n683 0.152939
R21183 vdd.n685 vdd.n684 0.152939
R21184 vdd.n690 vdd.n685 0.152939
R21185 vdd.n691 vdd.n690 0.152939
R21186 vdd.n692 vdd.n691 0.152939
R21187 vdd.n693 vdd.n692 0.152939
R21188 vdd.n696 vdd.n693 0.152939
R21189 vdd.n697 vdd.n696 0.152939
R21190 vdd.n698 vdd.n697 0.152939
R21191 vdd.n699 vdd.n698 0.152939
R21192 vdd.n702 vdd.n699 0.152939
R21193 vdd.n703 vdd.n702 0.152939
R21194 vdd.n704 vdd.n703 0.152939
R21195 vdd.n705 vdd.n704 0.152939
R21196 vdd.n708 vdd.n705 0.152939
R21197 vdd.n709 vdd.n708 0.152939
R21198 vdd.n710 vdd.n709 0.152939
R21199 vdd.n711 vdd.n710 0.152939
R21200 vdd.n714 vdd.n711 0.152939
R21201 vdd.n715 vdd.n714 0.152939
R21202 vdd.n716 vdd.n715 0.152939
R21203 vdd.n717 vdd.n716 0.152939
R21204 vdd.n720 vdd.n717 0.152939
R21205 vdd.n721 vdd.n720 0.152939
R21206 vdd.n3150 vdd.n721 0.152939
R21207 vdd.n3150 vdd.n3149 0.152939
R21208 vdd.n3149 vdd.n3148 0.152939
R21209 vdd.n3148 vdd.n725 0.152939
R21210 vdd.n730 vdd.n725 0.152939
R21211 vdd.n731 vdd.n730 0.152939
R21212 vdd.n734 vdd.n731 0.152939
R21213 vdd.n735 vdd.n734 0.152939
R21214 vdd.n736 vdd.n735 0.152939
R21215 vdd.n737 vdd.n736 0.152939
R21216 vdd.n740 vdd.n737 0.152939
R21217 vdd.n741 vdd.n740 0.152939
R21218 vdd.n742 vdd.n741 0.152939
R21219 vdd.n743 vdd.n742 0.152939
R21220 vdd.n746 vdd.n743 0.152939
R21221 vdd.n747 vdd.n746 0.152939
R21222 vdd.n748 vdd.n747 0.152939
R21223 vdd.n3233 vdd.n661 0.152939
R21224 vdd.n3234 vdd.n651 0.152939
R21225 vdd.n3248 vdd.n651 0.152939
R21226 vdd.n3249 vdd.n3248 0.152939
R21227 vdd.n3250 vdd.n3249 0.152939
R21228 vdd.n3250 vdd.n639 0.152939
R21229 vdd.n3264 vdd.n639 0.152939
R21230 vdd.n3265 vdd.n3264 0.152939
R21231 vdd.n3266 vdd.n3265 0.152939
R21232 vdd.n3266 vdd.n627 0.152939
R21233 vdd.n3281 vdd.n627 0.152939
R21234 vdd.n3282 vdd.n3281 0.152939
R21235 vdd.n3283 vdd.n3282 0.152939
R21236 vdd.n3283 vdd.n616 0.152939
R21237 vdd.n3300 vdd.n616 0.152939
R21238 vdd.n3301 vdd.n3300 0.152939
R21239 vdd.n3302 vdd.n3301 0.152939
R21240 vdd.n3302 vdd.n322 0.152939
R21241 vdd.n3382 vdd.n323 0.152939
R21242 vdd.n334 vdd.n323 0.152939
R21243 vdd.n335 vdd.n334 0.152939
R21244 vdd.n336 vdd.n335 0.152939
R21245 vdd.n343 vdd.n336 0.152939
R21246 vdd.n344 vdd.n343 0.152939
R21247 vdd.n345 vdd.n344 0.152939
R21248 vdd.n346 vdd.n345 0.152939
R21249 vdd.n354 vdd.n346 0.152939
R21250 vdd.n355 vdd.n354 0.152939
R21251 vdd.n356 vdd.n355 0.152939
R21252 vdd.n357 vdd.n356 0.152939
R21253 vdd.n365 vdd.n357 0.152939
R21254 vdd.n366 vdd.n365 0.152939
R21255 vdd.n367 vdd.n366 0.152939
R21256 vdd.n368 vdd.n367 0.152939
R21257 vdd.n443 vdd.n368 0.152939
R21258 vdd.n444 vdd.n442 0.152939
R21259 vdd.n451 vdd.n442 0.152939
R21260 vdd.n452 vdd.n451 0.152939
R21261 vdd.n453 vdd.n452 0.152939
R21262 vdd.n453 vdd.n440 0.152939
R21263 vdd.n461 vdd.n440 0.152939
R21264 vdd.n462 vdd.n461 0.152939
R21265 vdd.n463 vdd.n462 0.152939
R21266 vdd.n463 vdd.n438 0.152939
R21267 vdd.n471 vdd.n438 0.152939
R21268 vdd.n472 vdd.n471 0.152939
R21269 vdd.n473 vdd.n472 0.152939
R21270 vdd.n473 vdd.n436 0.152939
R21271 vdd.n481 vdd.n436 0.152939
R21272 vdd.n482 vdd.n481 0.152939
R21273 vdd.n483 vdd.n482 0.152939
R21274 vdd.n483 vdd.n434 0.152939
R21275 vdd.n491 vdd.n434 0.152939
R21276 vdd.n492 vdd.n491 0.152939
R21277 vdd.n493 vdd.n492 0.152939
R21278 vdd.n493 vdd.n430 0.152939
R21279 vdd.n501 vdd.n430 0.152939
R21280 vdd.n502 vdd.n501 0.152939
R21281 vdd.n503 vdd.n502 0.152939
R21282 vdd.n503 vdd.n428 0.152939
R21283 vdd.n511 vdd.n428 0.152939
R21284 vdd.n512 vdd.n511 0.152939
R21285 vdd.n513 vdd.n512 0.152939
R21286 vdd.n513 vdd.n426 0.152939
R21287 vdd.n521 vdd.n426 0.152939
R21288 vdd.n522 vdd.n521 0.152939
R21289 vdd.n523 vdd.n522 0.152939
R21290 vdd.n523 vdd.n424 0.152939
R21291 vdd.n531 vdd.n424 0.152939
R21292 vdd.n532 vdd.n531 0.152939
R21293 vdd.n533 vdd.n532 0.152939
R21294 vdd.n533 vdd.n422 0.152939
R21295 vdd.n541 vdd.n422 0.152939
R21296 vdd.n542 vdd.n541 0.152939
R21297 vdd.n543 vdd.n542 0.152939
R21298 vdd.n543 vdd.n418 0.152939
R21299 vdd.n551 vdd.n418 0.152939
R21300 vdd.n552 vdd.n551 0.152939
R21301 vdd.n553 vdd.n552 0.152939
R21302 vdd.n553 vdd.n416 0.152939
R21303 vdd.n561 vdd.n416 0.152939
R21304 vdd.n562 vdd.n561 0.152939
R21305 vdd.n563 vdd.n562 0.152939
R21306 vdd.n563 vdd.n414 0.152939
R21307 vdd.n571 vdd.n414 0.152939
R21308 vdd.n572 vdd.n571 0.152939
R21309 vdd.n573 vdd.n572 0.152939
R21310 vdd.n573 vdd.n412 0.152939
R21311 vdd.n581 vdd.n412 0.152939
R21312 vdd.n582 vdd.n581 0.152939
R21313 vdd.n583 vdd.n582 0.152939
R21314 vdd.n583 vdd.n410 0.152939
R21315 vdd.n591 vdd.n410 0.152939
R21316 vdd.n592 vdd.n591 0.152939
R21317 vdd.n593 vdd.n592 0.152939
R21318 vdd.n593 vdd.n408 0.152939
R21319 vdd.n600 vdd.n408 0.152939
R21320 vdd.n3341 vdd.n600 0.152939
R21321 vdd.n3241 vdd.n3240 0.152939
R21322 vdd.n3242 vdd.n3241 0.152939
R21323 vdd.n3242 vdd.n645 0.152939
R21324 vdd.n3256 vdd.n645 0.152939
R21325 vdd.n3257 vdd.n3256 0.152939
R21326 vdd.n3258 vdd.n3257 0.152939
R21327 vdd.n3258 vdd.n632 0.152939
R21328 vdd.n3272 vdd.n632 0.152939
R21329 vdd.n3273 vdd.n3272 0.152939
R21330 vdd.n3274 vdd.n3273 0.152939
R21331 vdd.n3274 vdd.n621 0.152939
R21332 vdd.n3289 vdd.n621 0.152939
R21333 vdd.n3290 vdd.n3289 0.152939
R21334 vdd.n3291 vdd.n3290 0.152939
R21335 vdd.n3293 vdd.n3291 0.152939
R21336 vdd.n3293 vdd.n3292 0.152939
R21337 vdd.n3292 vdd.n611 0.152939
R21338 vdd.n611 vdd.n609 0.152939
R21339 vdd.n3311 vdd.n609 0.152939
R21340 vdd.n3312 vdd.n3311 0.152939
R21341 vdd.n3313 vdd.n3312 0.152939
R21342 vdd.n3313 vdd.n607 0.152939
R21343 vdd.n3318 vdd.n607 0.152939
R21344 vdd.n3319 vdd.n3318 0.152939
R21345 vdd.n3320 vdd.n3319 0.152939
R21346 vdd.n3320 vdd.n605 0.152939
R21347 vdd.n3325 vdd.n605 0.152939
R21348 vdd.n3326 vdd.n3325 0.152939
R21349 vdd.n3327 vdd.n3326 0.152939
R21350 vdd.n3327 vdd.n603 0.152939
R21351 vdd.n3333 vdd.n603 0.152939
R21352 vdd.n3334 vdd.n3333 0.152939
R21353 vdd.n3335 vdd.n3334 0.152939
R21354 vdd.n3335 vdd.n601 0.152939
R21355 vdd.n3340 vdd.n601 0.152939
R21356 vdd.n3103 vdd.n656 0.152939
R21357 vdd.n2190 vdd.n1395 0.152939
R21358 vdd.n1741 vdd.n1740 0.152939
R21359 vdd.n1741 vdd.n1497 0.152939
R21360 vdd.n1755 vdd.n1497 0.152939
R21361 vdd.n1756 vdd.n1755 0.152939
R21362 vdd.n1757 vdd.n1756 0.152939
R21363 vdd.n1757 vdd.n1485 0.152939
R21364 vdd.n1772 vdd.n1485 0.152939
R21365 vdd.n1773 vdd.n1772 0.152939
R21366 vdd.n1774 vdd.n1773 0.152939
R21367 vdd.n1774 vdd.n1475 0.152939
R21368 vdd.n1789 vdd.n1475 0.152939
R21369 vdd.n1790 vdd.n1789 0.152939
R21370 vdd.n1791 vdd.n1790 0.152939
R21371 vdd.n1791 vdd.n1462 0.152939
R21372 vdd.n1805 vdd.n1462 0.152939
R21373 vdd.n1806 vdd.n1805 0.152939
R21374 vdd.n1807 vdd.n1806 0.152939
R21375 vdd.n1807 vdd.n1451 0.152939
R21376 vdd.n2117 vdd.n1451 0.152939
R21377 vdd.n2118 vdd.n2117 0.152939
R21378 vdd.n2119 vdd.n2118 0.152939
R21379 vdd.n2119 vdd.n1440 0.152939
R21380 vdd.n2133 vdd.n1440 0.152939
R21381 vdd.n2134 vdd.n2133 0.152939
R21382 vdd.n2135 vdd.n2134 0.152939
R21383 vdd.n2135 vdd.n1428 0.152939
R21384 vdd.n2150 vdd.n1428 0.152939
R21385 vdd.n2151 vdd.n2150 0.152939
R21386 vdd.n2152 vdd.n2151 0.152939
R21387 vdd.n2152 vdd.n1418 0.152939
R21388 vdd.n2167 vdd.n1418 0.152939
R21389 vdd.n2168 vdd.n2167 0.152939
R21390 vdd.n2171 vdd.n2168 0.152939
R21391 vdd.n2171 vdd.n2170 0.152939
R21392 vdd.n2170 vdd.n2169 0.152939
R21393 vdd.n1731 vdd.n1546 0.152939
R21394 vdd.n1731 vdd.n1730 0.152939
R21395 vdd.n1730 vdd.n1729 0.152939
R21396 vdd.n1729 vdd.n1548 0.152939
R21397 vdd.n1725 vdd.n1548 0.152939
R21398 vdd.n1725 vdd.n1724 0.152939
R21399 vdd.n1724 vdd.n1723 0.152939
R21400 vdd.n1723 vdd.n1553 0.152939
R21401 vdd.n1719 vdd.n1553 0.152939
R21402 vdd.n1719 vdd.n1718 0.152939
R21403 vdd.n1718 vdd.n1717 0.152939
R21404 vdd.n1717 vdd.n1559 0.152939
R21405 vdd.n1713 vdd.n1559 0.152939
R21406 vdd.n1713 vdd.n1712 0.152939
R21407 vdd.n1712 vdd.n1711 0.152939
R21408 vdd.n1711 vdd.n1565 0.152939
R21409 vdd.n1707 vdd.n1565 0.152939
R21410 vdd.n1707 vdd.n1706 0.152939
R21411 vdd.n1706 vdd.n1705 0.152939
R21412 vdd.n1705 vdd.n1571 0.152939
R21413 vdd.n1697 vdd.n1571 0.152939
R21414 vdd.n1697 vdd.n1696 0.152939
R21415 vdd.n1696 vdd.n1695 0.152939
R21416 vdd.n1695 vdd.n1575 0.152939
R21417 vdd.n1691 vdd.n1575 0.152939
R21418 vdd.n1691 vdd.n1690 0.152939
R21419 vdd.n1690 vdd.n1689 0.152939
R21420 vdd.n1689 vdd.n1581 0.152939
R21421 vdd.n1685 vdd.n1581 0.152939
R21422 vdd.n1685 vdd.n1684 0.152939
R21423 vdd.n1684 vdd.n1683 0.152939
R21424 vdd.n1683 vdd.n1587 0.152939
R21425 vdd.n1679 vdd.n1587 0.152939
R21426 vdd.n1679 vdd.n1678 0.152939
R21427 vdd.n1678 vdd.n1677 0.152939
R21428 vdd.n1677 vdd.n1593 0.152939
R21429 vdd.n1673 vdd.n1593 0.152939
R21430 vdd.n1673 vdd.n1672 0.152939
R21431 vdd.n1672 vdd.n1671 0.152939
R21432 vdd.n1671 vdd.n1599 0.152939
R21433 vdd.n1664 vdd.n1599 0.152939
R21434 vdd.n1664 vdd.n1663 0.152939
R21435 vdd.n1663 vdd.n1662 0.152939
R21436 vdd.n1662 vdd.n1604 0.152939
R21437 vdd.n1658 vdd.n1604 0.152939
R21438 vdd.n1658 vdd.n1657 0.152939
R21439 vdd.n1657 vdd.n1656 0.152939
R21440 vdd.n1656 vdd.n1610 0.152939
R21441 vdd.n1652 vdd.n1610 0.152939
R21442 vdd.n1652 vdd.n1651 0.152939
R21443 vdd.n1651 vdd.n1650 0.152939
R21444 vdd.n1650 vdd.n1616 0.152939
R21445 vdd.n1646 vdd.n1616 0.152939
R21446 vdd.n1646 vdd.n1645 0.152939
R21447 vdd.n1645 vdd.n1644 0.152939
R21448 vdd.n1644 vdd.n1622 0.152939
R21449 vdd.n1640 vdd.n1622 0.152939
R21450 vdd.n1640 vdd.n1639 0.152939
R21451 vdd.n1639 vdd.n1638 0.152939
R21452 vdd.n1638 vdd.n1628 0.152939
R21453 vdd.n1634 vdd.n1628 0.152939
R21454 vdd.n1634 vdd.n1509 0.152939
R21455 vdd.n1739 vdd.n1509 0.152939
R21456 vdd.n1747 vdd.n1503 0.152939
R21457 vdd.n1748 vdd.n1747 0.152939
R21458 vdd.n1749 vdd.n1748 0.152939
R21459 vdd.n1749 vdd.n1491 0.152939
R21460 vdd.n1764 vdd.n1491 0.152939
R21461 vdd.n1765 vdd.n1764 0.152939
R21462 vdd.n1766 vdd.n1765 0.152939
R21463 vdd.n1766 vdd.n1480 0.152939
R21464 vdd.n1781 vdd.n1480 0.152939
R21465 vdd.n1782 vdd.n1781 0.152939
R21466 vdd.n1783 vdd.n1782 0.152939
R21467 vdd.n1783 vdd.n1469 0.152939
R21468 vdd.n1797 vdd.n1469 0.152939
R21469 vdd.n1798 vdd.n1797 0.152939
R21470 vdd.n1799 vdd.n1798 0.152939
R21471 vdd.n1799 vdd.n1457 0.152939
R21472 vdd.n1814 vdd.n1457 0.152939
R21473 vdd.n2298 vdd.n2297 0.110256
R21474 vdd.n3034 vdd.n661 0.110256
R21475 vdd.n3103 vdd.n3102 0.110256
R21476 vdd.n2191 vdd.n2190 0.110256
R21477 vdd.n2110 vdd.n2109 0.0695946
R21478 vdd.n3383 vdd.n322 0.0695946
R21479 vdd.n3383 vdd.n3382 0.0695946
R21480 vdd.n2109 vdd.n1814 0.0695946
R21481 vdd.n2298 vdd.n1091 0.0431829
R21482 vdd.n2191 vdd.n1191 0.0431829
R21483 vdd.n3034 vdd.n667 0.0431829
R21484 vdd.n3102 vdd.n748 0.0431829
R21485 vdd vdd.n28 0.00833333
R21486 CSoutput.n19 CSoutput.t206 184.661
R21487 CSoutput.n78 CSoutput.n77 165.8
R21488 CSoutput.n76 CSoutput.n0 165.8
R21489 CSoutput.n75 CSoutput.n74 165.8
R21490 CSoutput.n73 CSoutput.n72 165.8
R21491 CSoutput.n71 CSoutput.n2 165.8
R21492 CSoutput.n69 CSoutput.n68 165.8
R21493 CSoutput.n67 CSoutput.n3 165.8
R21494 CSoutput.n66 CSoutput.n65 165.8
R21495 CSoutput.n63 CSoutput.n4 165.8
R21496 CSoutput.n61 CSoutput.n60 165.8
R21497 CSoutput.n59 CSoutput.n5 165.8
R21498 CSoutput.n58 CSoutput.n57 165.8
R21499 CSoutput.n55 CSoutput.n6 165.8
R21500 CSoutput.n54 CSoutput.n53 165.8
R21501 CSoutput.n52 CSoutput.n51 165.8
R21502 CSoutput.n50 CSoutput.n8 165.8
R21503 CSoutput.n48 CSoutput.n47 165.8
R21504 CSoutput.n46 CSoutput.n9 165.8
R21505 CSoutput.n45 CSoutput.n44 165.8
R21506 CSoutput.n42 CSoutput.n10 165.8
R21507 CSoutput.n41 CSoutput.n40 165.8
R21508 CSoutput.n39 CSoutput.n38 165.8
R21509 CSoutput.n37 CSoutput.n12 165.8
R21510 CSoutput.n35 CSoutput.n34 165.8
R21511 CSoutput.n33 CSoutput.n13 165.8
R21512 CSoutput.n32 CSoutput.n31 165.8
R21513 CSoutput.n29 CSoutput.n14 165.8
R21514 CSoutput.n28 CSoutput.n27 165.8
R21515 CSoutput.n26 CSoutput.n25 165.8
R21516 CSoutput.n24 CSoutput.n16 165.8
R21517 CSoutput.n22 CSoutput.n21 165.8
R21518 CSoutput.n20 CSoutput.n17 165.8
R21519 CSoutput.n77 CSoutput.t207 162.194
R21520 CSoutput.n18 CSoutput.t208 120.501
R21521 CSoutput.n23 CSoutput.t196 120.501
R21522 CSoutput.n15 CSoutput.t194 120.501
R21523 CSoutput.n30 CSoutput.t210 120.501
R21524 CSoutput.n36 CSoutput.t198 120.501
R21525 CSoutput.n11 CSoutput.t200 120.501
R21526 CSoutput.n43 CSoutput.t213 120.501
R21527 CSoutput.n49 CSoutput.t201 120.501
R21528 CSoutput.n7 CSoutput.t203 120.501
R21529 CSoutput.n56 CSoutput.t197 120.501
R21530 CSoutput.n62 CSoutput.t211 120.501
R21531 CSoutput.n64 CSoutput.t205 120.501
R21532 CSoutput.n70 CSoutput.t199 120.501
R21533 CSoutput.n1 CSoutput.t195 120.501
R21534 CSoutput.n310 CSoutput.n308 103.469
R21535 CSoutput.n294 CSoutput.n292 103.469
R21536 CSoutput.n279 CSoutput.n277 103.469
R21537 CSoutput.n112 CSoutput.n110 103.469
R21538 CSoutput.n96 CSoutput.n94 103.469
R21539 CSoutput.n81 CSoutput.n79 103.469
R21540 CSoutput.n320 CSoutput.n319 103.111
R21541 CSoutput.n318 CSoutput.n317 103.111
R21542 CSoutput.n316 CSoutput.n315 103.111
R21543 CSoutput.n314 CSoutput.n313 103.111
R21544 CSoutput.n312 CSoutput.n311 103.111
R21545 CSoutput.n310 CSoutput.n309 103.111
R21546 CSoutput.n306 CSoutput.n305 103.111
R21547 CSoutput.n304 CSoutput.n303 103.111
R21548 CSoutput.n302 CSoutput.n301 103.111
R21549 CSoutput.n300 CSoutput.n299 103.111
R21550 CSoutput.n298 CSoutput.n297 103.111
R21551 CSoutput.n296 CSoutput.n295 103.111
R21552 CSoutput.n294 CSoutput.n293 103.111
R21553 CSoutput.n291 CSoutput.n290 103.111
R21554 CSoutput.n289 CSoutput.n288 103.111
R21555 CSoutput.n287 CSoutput.n286 103.111
R21556 CSoutput.n285 CSoutput.n284 103.111
R21557 CSoutput.n283 CSoutput.n282 103.111
R21558 CSoutput.n281 CSoutput.n280 103.111
R21559 CSoutput.n279 CSoutput.n278 103.111
R21560 CSoutput.n112 CSoutput.n111 103.111
R21561 CSoutput.n114 CSoutput.n113 103.111
R21562 CSoutput.n116 CSoutput.n115 103.111
R21563 CSoutput.n118 CSoutput.n117 103.111
R21564 CSoutput.n120 CSoutput.n119 103.111
R21565 CSoutput.n122 CSoutput.n121 103.111
R21566 CSoutput.n124 CSoutput.n123 103.111
R21567 CSoutput.n96 CSoutput.n95 103.111
R21568 CSoutput.n98 CSoutput.n97 103.111
R21569 CSoutput.n100 CSoutput.n99 103.111
R21570 CSoutput.n102 CSoutput.n101 103.111
R21571 CSoutput.n104 CSoutput.n103 103.111
R21572 CSoutput.n106 CSoutput.n105 103.111
R21573 CSoutput.n108 CSoutput.n107 103.111
R21574 CSoutput.n81 CSoutput.n80 103.111
R21575 CSoutput.n83 CSoutput.n82 103.111
R21576 CSoutput.n85 CSoutput.n84 103.111
R21577 CSoutput.n87 CSoutput.n86 103.111
R21578 CSoutput.n89 CSoutput.n88 103.111
R21579 CSoutput.n91 CSoutput.n90 103.111
R21580 CSoutput.n93 CSoutput.n92 103.111
R21581 CSoutput.n322 CSoutput.n321 103.111
R21582 CSoutput.n358 CSoutput.n356 81.5057
R21583 CSoutput.n342 CSoutput.n340 81.5057
R21584 CSoutput.n327 CSoutput.n325 81.5057
R21585 CSoutput.n406 CSoutput.n404 81.5057
R21586 CSoutput.n390 CSoutput.n388 81.5057
R21587 CSoutput.n375 CSoutput.n373 81.5057
R21588 CSoutput.n370 CSoutput.n369 80.9324
R21589 CSoutput.n368 CSoutput.n367 80.9324
R21590 CSoutput.n366 CSoutput.n365 80.9324
R21591 CSoutput.n364 CSoutput.n363 80.9324
R21592 CSoutput.n362 CSoutput.n361 80.9324
R21593 CSoutput.n360 CSoutput.n359 80.9324
R21594 CSoutput.n358 CSoutput.n357 80.9324
R21595 CSoutput.n354 CSoutput.n353 80.9324
R21596 CSoutput.n352 CSoutput.n351 80.9324
R21597 CSoutput.n350 CSoutput.n349 80.9324
R21598 CSoutput.n348 CSoutput.n347 80.9324
R21599 CSoutput.n346 CSoutput.n345 80.9324
R21600 CSoutput.n344 CSoutput.n343 80.9324
R21601 CSoutput.n342 CSoutput.n341 80.9324
R21602 CSoutput.n339 CSoutput.n338 80.9324
R21603 CSoutput.n337 CSoutput.n336 80.9324
R21604 CSoutput.n335 CSoutput.n334 80.9324
R21605 CSoutput.n333 CSoutput.n332 80.9324
R21606 CSoutput.n331 CSoutput.n330 80.9324
R21607 CSoutput.n329 CSoutput.n328 80.9324
R21608 CSoutput.n327 CSoutput.n326 80.9324
R21609 CSoutput.n406 CSoutput.n405 80.9324
R21610 CSoutput.n408 CSoutput.n407 80.9324
R21611 CSoutput.n410 CSoutput.n409 80.9324
R21612 CSoutput.n412 CSoutput.n411 80.9324
R21613 CSoutput.n414 CSoutput.n413 80.9324
R21614 CSoutput.n416 CSoutput.n415 80.9324
R21615 CSoutput.n418 CSoutput.n417 80.9324
R21616 CSoutput.n390 CSoutput.n389 80.9324
R21617 CSoutput.n392 CSoutput.n391 80.9324
R21618 CSoutput.n394 CSoutput.n393 80.9324
R21619 CSoutput.n396 CSoutput.n395 80.9324
R21620 CSoutput.n398 CSoutput.n397 80.9324
R21621 CSoutput.n400 CSoutput.n399 80.9324
R21622 CSoutput.n402 CSoutput.n401 80.9324
R21623 CSoutput.n375 CSoutput.n374 80.9324
R21624 CSoutput.n377 CSoutput.n376 80.9324
R21625 CSoutput.n379 CSoutput.n378 80.9324
R21626 CSoutput.n381 CSoutput.n380 80.9324
R21627 CSoutput.n383 CSoutput.n382 80.9324
R21628 CSoutput.n385 CSoutput.n384 80.9324
R21629 CSoutput.n387 CSoutput.n386 80.9324
R21630 CSoutput.n25 CSoutput.n24 48.1486
R21631 CSoutput.n69 CSoutput.n3 48.1486
R21632 CSoutput.n38 CSoutput.n37 48.1486
R21633 CSoutput.n42 CSoutput.n41 48.1486
R21634 CSoutput.n51 CSoutput.n50 48.1486
R21635 CSoutput.n55 CSoutput.n54 48.1486
R21636 CSoutput.n22 CSoutput.n17 46.462
R21637 CSoutput.n72 CSoutput.n71 46.462
R21638 CSoutput.n20 CSoutput.n19 44.9055
R21639 CSoutput.n29 CSoutput.n28 43.7635
R21640 CSoutput.n65 CSoutput.n63 43.7635
R21641 CSoutput.n35 CSoutput.n13 41.7396
R21642 CSoutput.n57 CSoutput.n5 41.7396
R21643 CSoutput.n44 CSoutput.n9 37.0171
R21644 CSoutput.n48 CSoutput.n9 37.0171
R21645 CSoutput.n76 CSoutput.n75 34.9932
R21646 CSoutput.n31 CSoutput.n13 32.2947
R21647 CSoutput.n61 CSoutput.n5 32.2947
R21648 CSoutput.n30 CSoutput.n29 29.6014
R21649 CSoutput.n63 CSoutput.n62 29.6014
R21650 CSoutput.n19 CSoutput.n18 28.4085
R21651 CSoutput.n18 CSoutput.n17 25.1176
R21652 CSoutput.n72 CSoutput.n1 25.1176
R21653 CSoutput.n43 CSoutput.n42 22.0922
R21654 CSoutput.n50 CSoutput.n49 22.0922
R21655 CSoutput.n77 CSoutput.n76 21.8586
R21656 CSoutput.n37 CSoutput.n36 18.9681
R21657 CSoutput.n56 CSoutput.n55 18.9681
R21658 CSoutput.n25 CSoutput.n15 17.6292
R21659 CSoutput.n64 CSoutput.n3 17.6292
R21660 CSoutput.n24 CSoutput.n23 15.844
R21661 CSoutput.n70 CSoutput.n69 15.844
R21662 CSoutput.n38 CSoutput.n11 14.5051
R21663 CSoutput.n54 CSoutput.n7 14.5051
R21664 CSoutput.n421 CSoutput.n78 11.4982
R21665 CSoutput.n41 CSoutput.n11 11.3811
R21666 CSoutput.n51 CSoutput.n7 11.3811
R21667 CSoutput.n23 CSoutput.n22 10.0422
R21668 CSoutput.n71 CSoutput.n70 10.0422
R21669 CSoutput.n307 CSoutput.n291 9.25285
R21670 CSoutput.n109 CSoutput.n93 9.25285
R21671 CSoutput.n355 CSoutput.n339 8.98182
R21672 CSoutput.n403 CSoutput.n387 8.98182
R21673 CSoutput.n372 CSoutput.n324 8.92798
R21674 CSoutput.n28 CSoutput.n15 8.25698
R21675 CSoutput.n65 CSoutput.n64 8.25698
R21676 CSoutput.n324 CSoutput.n323 7.12641
R21677 CSoutput.n126 CSoutput.n125 7.12641
R21678 CSoutput.n36 CSoutput.n35 6.91809
R21679 CSoutput.n57 CSoutput.n56 6.91809
R21680 CSoutput.n372 CSoutput.n371 6.02792
R21681 CSoutput.n420 CSoutput.n419 6.02792
R21682 CSoutput.n421 CSoutput.n126 5.33554
R21683 CSoutput.n371 CSoutput.n370 5.25266
R21684 CSoutput.n355 CSoutput.n354 5.25266
R21685 CSoutput.n419 CSoutput.n418 5.25266
R21686 CSoutput.n403 CSoutput.n402 5.25266
R21687 CSoutput.n323 CSoutput.n322 5.1449
R21688 CSoutput.n307 CSoutput.n306 5.1449
R21689 CSoutput.n125 CSoutput.n124 5.1449
R21690 CSoutput.n109 CSoutput.n108 5.1449
R21691 CSoutput.n217 CSoutput.n170 4.5005
R21692 CSoutput.n186 CSoutput.n170 4.5005
R21693 CSoutput.n181 CSoutput.n165 4.5005
R21694 CSoutput.n181 CSoutput.n167 4.5005
R21695 CSoutput.n181 CSoutput.n164 4.5005
R21696 CSoutput.n181 CSoutput.n168 4.5005
R21697 CSoutput.n181 CSoutput.n163 4.5005
R21698 CSoutput.n181 CSoutput.t209 4.5005
R21699 CSoutput.n181 CSoutput.n162 4.5005
R21700 CSoutput.n181 CSoutput.n169 4.5005
R21701 CSoutput.n181 CSoutput.n170 4.5005
R21702 CSoutput.n179 CSoutput.n165 4.5005
R21703 CSoutput.n179 CSoutput.n167 4.5005
R21704 CSoutput.n179 CSoutput.n164 4.5005
R21705 CSoutput.n179 CSoutput.n168 4.5005
R21706 CSoutput.n179 CSoutput.n163 4.5005
R21707 CSoutput.n179 CSoutput.t209 4.5005
R21708 CSoutput.n179 CSoutput.n162 4.5005
R21709 CSoutput.n179 CSoutput.n169 4.5005
R21710 CSoutput.n179 CSoutput.n170 4.5005
R21711 CSoutput.n178 CSoutput.n165 4.5005
R21712 CSoutput.n178 CSoutput.n167 4.5005
R21713 CSoutput.n178 CSoutput.n164 4.5005
R21714 CSoutput.n178 CSoutput.n168 4.5005
R21715 CSoutput.n178 CSoutput.n163 4.5005
R21716 CSoutput.n178 CSoutput.t209 4.5005
R21717 CSoutput.n178 CSoutput.n162 4.5005
R21718 CSoutput.n178 CSoutput.n169 4.5005
R21719 CSoutput.n178 CSoutput.n170 4.5005
R21720 CSoutput.n263 CSoutput.n165 4.5005
R21721 CSoutput.n263 CSoutput.n167 4.5005
R21722 CSoutput.n263 CSoutput.n164 4.5005
R21723 CSoutput.n263 CSoutput.n168 4.5005
R21724 CSoutput.n263 CSoutput.n163 4.5005
R21725 CSoutput.n263 CSoutput.t209 4.5005
R21726 CSoutput.n263 CSoutput.n162 4.5005
R21727 CSoutput.n263 CSoutput.n169 4.5005
R21728 CSoutput.n263 CSoutput.n170 4.5005
R21729 CSoutput.n261 CSoutput.n165 4.5005
R21730 CSoutput.n261 CSoutput.n167 4.5005
R21731 CSoutput.n261 CSoutput.n164 4.5005
R21732 CSoutput.n261 CSoutput.n168 4.5005
R21733 CSoutput.n261 CSoutput.n163 4.5005
R21734 CSoutput.n261 CSoutput.t209 4.5005
R21735 CSoutput.n261 CSoutput.n162 4.5005
R21736 CSoutput.n261 CSoutput.n169 4.5005
R21737 CSoutput.n259 CSoutput.n165 4.5005
R21738 CSoutput.n259 CSoutput.n167 4.5005
R21739 CSoutput.n259 CSoutput.n164 4.5005
R21740 CSoutput.n259 CSoutput.n168 4.5005
R21741 CSoutput.n259 CSoutput.n163 4.5005
R21742 CSoutput.n259 CSoutput.t209 4.5005
R21743 CSoutput.n259 CSoutput.n162 4.5005
R21744 CSoutput.n259 CSoutput.n169 4.5005
R21745 CSoutput.n189 CSoutput.n165 4.5005
R21746 CSoutput.n189 CSoutput.n167 4.5005
R21747 CSoutput.n189 CSoutput.n164 4.5005
R21748 CSoutput.n189 CSoutput.n168 4.5005
R21749 CSoutput.n189 CSoutput.n163 4.5005
R21750 CSoutput.n189 CSoutput.t209 4.5005
R21751 CSoutput.n189 CSoutput.n162 4.5005
R21752 CSoutput.n189 CSoutput.n169 4.5005
R21753 CSoutput.n189 CSoutput.n170 4.5005
R21754 CSoutput.n188 CSoutput.n165 4.5005
R21755 CSoutput.n188 CSoutput.n167 4.5005
R21756 CSoutput.n188 CSoutput.n164 4.5005
R21757 CSoutput.n188 CSoutput.n168 4.5005
R21758 CSoutput.n188 CSoutput.n163 4.5005
R21759 CSoutput.n188 CSoutput.t209 4.5005
R21760 CSoutput.n188 CSoutput.n162 4.5005
R21761 CSoutput.n188 CSoutput.n169 4.5005
R21762 CSoutput.n188 CSoutput.n170 4.5005
R21763 CSoutput.n192 CSoutput.n165 4.5005
R21764 CSoutput.n192 CSoutput.n167 4.5005
R21765 CSoutput.n192 CSoutput.n164 4.5005
R21766 CSoutput.n192 CSoutput.n168 4.5005
R21767 CSoutput.n192 CSoutput.n163 4.5005
R21768 CSoutput.n192 CSoutput.t209 4.5005
R21769 CSoutput.n192 CSoutput.n162 4.5005
R21770 CSoutput.n192 CSoutput.n169 4.5005
R21771 CSoutput.n192 CSoutput.n170 4.5005
R21772 CSoutput.n191 CSoutput.n165 4.5005
R21773 CSoutput.n191 CSoutput.n167 4.5005
R21774 CSoutput.n191 CSoutput.n164 4.5005
R21775 CSoutput.n191 CSoutput.n168 4.5005
R21776 CSoutput.n191 CSoutput.n163 4.5005
R21777 CSoutput.n191 CSoutput.t209 4.5005
R21778 CSoutput.n191 CSoutput.n162 4.5005
R21779 CSoutput.n191 CSoutput.n169 4.5005
R21780 CSoutput.n191 CSoutput.n170 4.5005
R21781 CSoutput.n174 CSoutput.n165 4.5005
R21782 CSoutput.n174 CSoutput.n167 4.5005
R21783 CSoutput.n174 CSoutput.n164 4.5005
R21784 CSoutput.n174 CSoutput.n168 4.5005
R21785 CSoutput.n174 CSoutput.n163 4.5005
R21786 CSoutput.n174 CSoutput.t209 4.5005
R21787 CSoutput.n174 CSoutput.n162 4.5005
R21788 CSoutput.n174 CSoutput.n169 4.5005
R21789 CSoutput.n174 CSoutput.n170 4.5005
R21790 CSoutput.n266 CSoutput.n165 4.5005
R21791 CSoutput.n266 CSoutput.n167 4.5005
R21792 CSoutput.n266 CSoutput.n164 4.5005
R21793 CSoutput.n266 CSoutput.n168 4.5005
R21794 CSoutput.n266 CSoutput.n163 4.5005
R21795 CSoutput.n266 CSoutput.t209 4.5005
R21796 CSoutput.n266 CSoutput.n162 4.5005
R21797 CSoutput.n266 CSoutput.n169 4.5005
R21798 CSoutput.n266 CSoutput.n170 4.5005
R21799 CSoutput.n253 CSoutput.n224 4.5005
R21800 CSoutput.n253 CSoutput.n230 4.5005
R21801 CSoutput.n211 CSoutput.n200 4.5005
R21802 CSoutput.n211 CSoutput.n202 4.5005
R21803 CSoutput.n211 CSoutput.n199 4.5005
R21804 CSoutput.n211 CSoutput.n203 4.5005
R21805 CSoutput.n211 CSoutput.n198 4.5005
R21806 CSoutput.n211 CSoutput.t202 4.5005
R21807 CSoutput.n211 CSoutput.n197 4.5005
R21808 CSoutput.n211 CSoutput.n204 4.5005
R21809 CSoutput.n253 CSoutput.n211 4.5005
R21810 CSoutput.n232 CSoutput.n200 4.5005
R21811 CSoutput.n232 CSoutput.n202 4.5005
R21812 CSoutput.n232 CSoutput.n199 4.5005
R21813 CSoutput.n232 CSoutput.n203 4.5005
R21814 CSoutput.n232 CSoutput.n198 4.5005
R21815 CSoutput.n232 CSoutput.t202 4.5005
R21816 CSoutput.n232 CSoutput.n197 4.5005
R21817 CSoutput.n232 CSoutput.n204 4.5005
R21818 CSoutput.n253 CSoutput.n232 4.5005
R21819 CSoutput.n210 CSoutput.n200 4.5005
R21820 CSoutput.n210 CSoutput.n202 4.5005
R21821 CSoutput.n210 CSoutput.n199 4.5005
R21822 CSoutput.n210 CSoutput.n203 4.5005
R21823 CSoutput.n210 CSoutput.n198 4.5005
R21824 CSoutput.n210 CSoutput.t202 4.5005
R21825 CSoutput.n210 CSoutput.n197 4.5005
R21826 CSoutput.n210 CSoutput.n204 4.5005
R21827 CSoutput.n253 CSoutput.n210 4.5005
R21828 CSoutput.n234 CSoutput.n200 4.5005
R21829 CSoutput.n234 CSoutput.n202 4.5005
R21830 CSoutput.n234 CSoutput.n199 4.5005
R21831 CSoutput.n234 CSoutput.n203 4.5005
R21832 CSoutput.n234 CSoutput.n198 4.5005
R21833 CSoutput.n234 CSoutput.t202 4.5005
R21834 CSoutput.n234 CSoutput.n197 4.5005
R21835 CSoutput.n234 CSoutput.n204 4.5005
R21836 CSoutput.n253 CSoutput.n234 4.5005
R21837 CSoutput.n200 CSoutput.n195 4.5005
R21838 CSoutput.n202 CSoutput.n195 4.5005
R21839 CSoutput.n199 CSoutput.n195 4.5005
R21840 CSoutput.n203 CSoutput.n195 4.5005
R21841 CSoutput.n198 CSoutput.n195 4.5005
R21842 CSoutput.t202 CSoutput.n195 4.5005
R21843 CSoutput.n197 CSoutput.n195 4.5005
R21844 CSoutput.n204 CSoutput.n195 4.5005
R21845 CSoutput.n256 CSoutput.n200 4.5005
R21846 CSoutput.n256 CSoutput.n202 4.5005
R21847 CSoutput.n256 CSoutput.n199 4.5005
R21848 CSoutput.n256 CSoutput.n203 4.5005
R21849 CSoutput.n256 CSoutput.n198 4.5005
R21850 CSoutput.n256 CSoutput.t202 4.5005
R21851 CSoutput.n256 CSoutput.n197 4.5005
R21852 CSoutput.n256 CSoutput.n204 4.5005
R21853 CSoutput.n254 CSoutput.n200 4.5005
R21854 CSoutput.n254 CSoutput.n202 4.5005
R21855 CSoutput.n254 CSoutput.n199 4.5005
R21856 CSoutput.n254 CSoutput.n203 4.5005
R21857 CSoutput.n254 CSoutput.n198 4.5005
R21858 CSoutput.n254 CSoutput.t202 4.5005
R21859 CSoutput.n254 CSoutput.n197 4.5005
R21860 CSoutput.n254 CSoutput.n204 4.5005
R21861 CSoutput.n254 CSoutput.n253 4.5005
R21862 CSoutput.n236 CSoutput.n200 4.5005
R21863 CSoutput.n236 CSoutput.n202 4.5005
R21864 CSoutput.n236 CSoutput.n199 4.5005
R21865 CSoutput.n236 CSoutput.n203 4.5005
R21866 CSoutput.n236 CSoutput.n198 4.5005
R21867 CSoutput.n236 CSoutput.t202 4.5005
R21868 CSoutput.n236 CSoutput.n197 4.5005
R21869 CSoutput.n236 CSoutput.n204 4.5005
R21870 CSoutput.n253 CSoutput.n236 4.5005
R21871 CSoutput.n208 CSoutput.n200 4.5005
R21872 CSoutput.n208 CSoutput.n202 4.5005
R21873 CSoutput.n208 CSoutput.n199 4.5005
R21874 CSoutput.n208 CSoutput.n203 4.5005
R21875 CSoutput.n208 CSoutput.n198 4.5005
R21876 CSoutput.n208 CSoutput.t202 4.5005
R21877 CSoutput.n208 CSoutput.n197 4.5005
R21878 CSoutput.n208 CSoutput.n204 4.5005
R21879 CSoutput.n253 CSoutput.n208 4.5005
R21880 CSoutput.n238 CSoutput.n200 4.5005
R21881 CSoutput.n238 CSoutput.n202 4.5005
R21882 CSoutput.n238 CSoutput.n199 4.5005
R21883 CSoutput.n238 CSoutput.n203 4.5005
R21884 CSoutput.n238 CSoutput.n198 4.5005
R21885 CSoutput.n238 CSoutput.t202 4.5005
R21886 CSoutput.n238 CSoutput.n197 4.5005
R21887 CSoutput.n238 CSoutput.n204 4.5005
R21888 CSoutput.n253 CSoutput.n238 4.5005
R21889 CSoutput.n207 CSoutput.n200 4.5005
R21890 CSoutput.n207 CSoutput.n202 4.5005
R21891 CSoutput.n207 CSoutput.n199 4.5005
R21892 CSoutput.n207 CSoutput.n203 4.5005
R21893 CSoutput.n207 CSoutput.n198 4.5005
R21894 CSoutput.n207 CSoutput.t202 4.5005
R21895 CSoutput.n207 CSoutput.n197 4.5005
R21896 CSoutput.n207 CSoutput.n204 4.5005
R21897 CSoutput.n253 CSoutput.n207 4.5005
R21898 CSoutput.n252 CSoutput.n200 4.5005
R21899 CSoutput.n252 CSoutput.n202 4.5005
R21900 CSoutput.n252 CSoutput.n199 4.5005
R21901 CSoutput.n252 CSoutput.n203 4.5005
R21902 CSoutput.n252 CSoutput.n198 4.5005
R21903 CSoutput.n252 CSoutput.t202 4.5005
R21904 CSoutput.n252 CSoutput.n197 4.5005
R21905 CSoutput.n252 CSoutput.n204 4.5005
R21906 CSoutput.n253 CSoutput.n252 4.5005
R21907 CSoutput.n251 CSoutput.n136 4.5005
R21908 CSoutput.n152 CSoutput.n136 4.5005
R21909 CSoutput.n147 CSoutput.n131 4.5005
R21910 CSoutput.n147 CSoutput.n133 4.5005
R21911 CSoutput.n147 CSoutput.n130 4.5005
R21912 CSoutput.n147 CSoutput.n134 4.5005
R21913 CSoutput.n147 CSoutput.n129 4.5005
R21914 CSoutput.n147 CSoutput.t192 4.5005
R21915 CSoutput.n147 CSoutput.n128 4.5005
R21916 CSoutput.n147 CSoutput.n135 4.5005
R21917 CSoutput.n147 CSoutput.n136 4.5005
R21918 CSoutput.n145 CSoutput.n131 4.5005
R21919 CSoutput.n145 CSoutput.n133 4.5005
R21920 CSoutput.n145 CSoutput.n130 4.5005
R21921 CSoutput.n145 CSoutput.n134 4.5005
R21922 CSoutput.n145 CSoutput.n129 4.5005
R21923 CSoutput.n145 CSoutput.t192 4.5005
R21924 CSoutput.n145 CSoutput.n128 4.5005
R21925 CSoutput.n145 CSoutput.n135 4.5005
R21926 CSoutput.n145 CSoutput.n136 4.5005
R21927 CSoutput.n144 CSoutput.n131 4.5005
R21928 CSoutput.n144 CSoutput.n133 4.5005
R21929 CSoutput.n144 CSoutput.n130 4.5005
R21930 CSoutput.n144 CSoutput.n134 4.5005
R21931 CSoutput.n144 CSoutput.n129 4.5005
R21932 CSoutput.n144 CSoutput.t192 4.5005
R21933 CSoutput.n144 CSoutput.n128 4.5005
R21934 CSoutput.n144 CSoutput.n135 4.5005
R21935 CSoutput.n144 CSoutput.n136 4.5005
R21936 CSoutput.n273 CSoutput.n131 4.5005
R21937 CSoutput.n273 CSoutput.n133 4.5005
R21938 CSoutput.n273 CSoutput.n130 4.5005
R21939 CSoutput.n273 CSoutput.n134 4.5005
R21940 CSoutput.n273 CSoutput.n129 4.5005
R21941 CSoutput.n273 CSoutput.t192 4.5005
R21942 CSoutput.n273 CSoutput.n128 4.5005
R21943 CSoutput.n273 CSoutput.n135 4.5005
R21944 CSoutput.n273 CSoutput.n136 4.5005
R21945 CSoutput.n271 CSoutput.n131 4.5005
R21946 CSoutput.n271 CSoutput.n133 4.5005
R21947 CSoutput.n271 CSoutput.n130 4.5005
R21948 CSoutput.n271 CSoutput.n134 4.5005
R21949 CSoutput.n271 CSoutput.n129 4.5005
R21950 CSoutput.n271 CSoutput.t192 4.5005
R21951 CSoutput.n271 CSoutput.n128 4.5005
R21952 CSoutput.n271 CSoutput.n135 4.5005
R21953 CSoutput.n269 CSoutput.n131 4.5005
R21954 CSoutput.n269 CSoutput.n133 4.5005
R21955 CSoutput.n269 CSoutput.n130 4.5005
R21956 CSoutput.n269 CSoutput.n134 4.5005
R21957 CSoutput.n269 CSoutput.n129 4.5005
R21958 CSoutput.n269 CSoutput.t192 4.5005
R21959 CSoutput.n269 CSoutput.n128 4.5005
R21960 CSoutput.n269 CSoutput.n135 4.5005
R21961 CSoutput.n155 CSoutput.n131 4.5005
R21962 CSoutput.n155 CSoutput.n133 4.5005
R21963 CSoutput.n155 CSoutput.n130 4.5005
R21964 CSoutput.n155 CSoutput.n134 4.5005
R21965 CSoutput.n155 CSoutput.n129 4.5005
R21966 CSoutput.n155 CSoutput.t192 4.5005
R21967 CSoutput.n155 CSoutput.n128 4.5005
R21968 CSoutput.n155 CSoutput.n135 4.5005
R21969 CSoutput.n155 CSoutput.n136 4.5005
R21970 CSoutput.n154 CSoutput.n131 4.5005
R21971 CSoutput.n154 CSoutput.n133 4.5005
R21972 CSoutput.n154 CSoutput.n130 4.5005
R21973 CSoutput.n154 CSoutput.n134 4.5005
R21974 CSoutput.n154 CSoutput.n129 4.5005
R21975 CSoutput.n154 CSoutput.t192 4.5005
R21976 CSoutput.n154 CSoutput.n128 4.5005
R21977 CSoutput.n154 CSoutput.n135 4.5005
R21978 CSoutput.n154 CSoutput.n136 4.5005
R21979 CSoutput.n158 CSoutput.n131 4.5005
R21980 CSoutput.n158 CSoutput.n133 4.5005
R21981 CSoutput.n158 CSoutput.n130 4.5005
R21982 CSoutput.n158 CSoutput.n134 4.5005
R21983 CSoutput.n158 CSoutput.n129 4.5005
R21984 CSoutput.n158 CSoutput.t192 4.5005
R21985 CSoutput.n158 CSoutput.n128 4.5005
R21986 CSoutput.n158 CSoutput.n135 4.5005
R21987 CSoutput.n158 CSoutput.n136 4.5005
R21988 CSoutput.n157 CSoutput.n131 4.5005
R21989 CSoutput.n157 CSoutput.n133 4.5005
R21990 CSoutput.n157 CSoutput.n130 4.5005
R21991 CSoutput.n157 CSoutput.n134 4.5005
R21992 CSoutput.n157 CSoutput.n129 4.5005
R21993 CSoutput.n157 CSoutput.t192 4.5005
R21994 CSoutput.n157 CSoutput.n128 4.5005
R21995 CSoutput.n157 CSoutput.n135 4.5005
R21996 CSoutput.n157 CSoutput.n136 4.5005
R21997 CSoutput.n140 CSoutput.n131 4.5005
R21998 CSoutput.n140 CSoutput.n133 4.5005
R21999 CSoutput.n140 CSoutput.n130 4.5005
R22000 CSoutput.n140 CSoutput.n134 4.5005
R22001 CSoutput.n140 CSoutput.n129 4.5005
R22002 CSoutput.n140 CSoutput.t192 4.5005
R22003 CSoutput.n140 CSoutput.n128 4.5005
R22004 CSoutput.n140 CSoutput.n135 4.5005
R22005 CSoutput.n140 CSoutput.n136 4.5005
R22006 CSoutput.n276 CSoutput.n131 4.5005
R22007 CSoutput.n276 CSoutput.n133 4.5005
R22008 CSoutput.n276 CSoutput.n130 4.5005
R22009 CSoutput.n276 CSoutput.n134 4.5005
R22010 CSoutput.n276 CSoutput.n129 4.5005
R22011 CSoutput.n276 CSoutput.t192 4.5005
R22012 CSoutput.n276 CSoutput.n128 4.5005
R22013 CSoutput.n276 CSoutput.n135 4.5005
R22014 CSoutput.n276 CSoutput.n136 4.5005
R22015 CSoutput.n323 CSoutput.n307 4.10845
R22016 CSoutput.n125 CSoutput.n109 4.10845
R22017 CSoutput.n321 CSoutput.t57 4.06363
R22018 CSoutput.n321 CSoutput.t75 4.06363
R22019 CSoutput.n319 CSoutput.t88 4.06363
R22020 CSoutput.n319 CSoutput.t19 4.06363
R22021 CSoutput.n317 CSoutput.t23 4.06363
R22022 CSoutput.n317 CSoutput.t79 4.06363
R22023 CSoutput.n315 CSoutput.t91 4.06363
R22024 CSoutput.n315 CSoutput.t92 4.06363
R22025 CSoutput.n313 CSoutput.t39 4.06363
R22026 CSoutput.n313 CSoutput.t40 4.06363
R22027 CSoutput.n311 CSoutput.t45 4.06363
R22028 CSoutput.n311 CSoutput.t93 4.06363
R22029 CSoutput.n309 CSoutput.t11 4.06363
R22030 CSoutput.n309 CSoutput.t43 4.06363
R22031 CSoutput.n308 CSoutput.t56 4.06363
R22032 CSoutput.n308 CSoutput.t74 4.06363
R22033 CSoutput.n305 CSoutput.t46 4.06363
R22034 CSoutput.n305 CSoutput.t66 4.06363
R22035 CSoutput.n303 CSoutput.t80 4.06363
R22036 CSoutput.n303 CSoutput.t7 4.06363
R22037 CSoutput.n301 CSoutput.t8 4.06363
R22038 CSoutput.n301 CSoutput.t68 4.06363
R22039 CSoutput.n299 CSoutput.t83 4.06363
R22040 CSoutput.n299 CSoutput.t84 4.06363
R22041 CSoutput.n297 CSoutput.t27 4.06363
R22042 CSoutput.n297 CSoutput.t28 4.06363
R22043 CSoutput.n295 CSoutput.t31 4.06363
R22044 CSoutput.n295 CSoutput.t85 4.06363
R22045 CSoutput.n293 CSoutput.t0 4.06363
R22046 CSoutput.n293 CSoutput.t30 4.06363
R22047 CSoutput.n292 CSoutput.t47 4.06363
R22048 CSoutput.n292 CSoutput.t67 4.06363
R22049 CSoutput.n290 CSoutput.t73 4.06363
R22050 CSoutput.n290 CSoutput.t36 4.06363
R22051 CSoutput.n288 CSoutput.t63 4.06363
R22052 CSoutput.n288 CSoutput.t18 4.06363
R22053 CSoutput.n286 CSoutput.t81 4.06363
R22054 CSoutput.n286 CSoutput.t12 4.06363
R22055 CSoutput.n284 CSoutput.t48 4.06363
R22056 CSoutput.n284 CSoutput.t29 4.06363
R22057 CSoutput.n282 CSoutput.t32 4.06363
R22058 CSoutput.n282 CSoutput.t9 4.06363
R22059 CSoutput.n280 CSoutput.t72 4.06363
R22060 CSoutput.n280 CSoutput.t4 4.06363
R22061 CSoutput.n278 CSoutput.t41 4.06363
R22062 CSoutput.n278 CSoutput.t89 4.06363
R22063 CSoutput.n277 CSoutput.t24 4.06363
R22064 CSoutput.n277 CSoutput.t77 4.06363
R22065 CSoutput.n110 CSoutput.t15 4.06363
R22066 CSoutput.n110 CSoutput.t86 4.06363
R22067 CSoutput.n111 CSoutput.t71 4.06363
R22068 CSoutput.n111 CSoutput.t53 4.06363
R22069 CSoutput.n113 CSoutput.t38 4.06363
R22070 CSoutput.n113 CSoutput.t95 4.06363
R22071 CSoutput.n115 CSoutput.t70 4.06363
R22072 CSoutput.n115 CSoutput.t69 4.06363
R22073 CSoutput.n117 CSoutput.t59 4.06363
R22074 CSoutput.n117 CSoutput.t35 4.06363
R22075 CSoutput.n119 CSoutput.t17 4.06363
R22076 CSoutput.n119 CSoutput.t60 4.06363
R22077 CSoutput.n121 CSoutput.t58 4.06363
R22078 CSoutput.n121 CSoutput.t33 4.06363
R22079 CSoutput.n123 CSoutput.t16 4.06363
R22080 CSoutput.n123 CSoutput.t14 4.06363
R22081 CSoutput.n94 CSoutput.t2 4.06363
R22082 CSoutput.n94 CSoutput.t76 4.06363
R22083 CSoutput.n95 CSoutput.t65 4.06363
R22084 CSoutput.n95 CSoutput.t44 4.06363
R22085 CSoutput.n97 CSoutput.t26 4.06363
R22086 CSoutput.n97 CSoutput.t87 4.06363
R22087 CSoutput.n99 CSoutput.t62 4.06363
R22088 CSoutput.n99 CSoutput.t61 4.06363
R22089 CSoutput.n101 CSoutput.t51 4.06363
R22090 CSoutput.n101 CSoutput.t22 4.06363
R22091 CSoutput.n103 CSoutput.t5 4.06363
R22092 CSoutput.n103 CSoutput.t52 4.06363
R22093 CSoutput.n105 CSoutput.t50 4.06363
R22094 CSoutput.n105 CSoutput.t20 4.06363
R22095 CSoutput.n107 CSoutput.t3 4.06363
R22096 CSoutput.n107 CSoutput.t1 4.06363
R22097 CSoutput.n79 CSoutput.t78 4.06363
R22098 CSoutput.n79 CSoutput.t25 4.06363
R22099 CSoutput.n80 CSoutput.t90 4.06363
R22100 CSoutput.n80 CSoutput.t42 4.06363
R22101 CSoutput.n82 CSoutput.t6 4.06363
R22102 CSoutput.n82 CSoutput.t54 4.06363
R22103 CSoutput.n84 CSoutput.t10 4.06363
R22104 CSoutput.n84 CSoutput.t34 4.06363
R22105 CSoutput.n86 CSoutput.t94 4.06363
R22106 CSoutput.n86 CSoutput.t49 4.06363
R22107 CSoutput.n88 CSoutput.t13 4.06363
R22108 CSoutput.n88 CSoutput.t82 4.06363
R22109 CSoutput.n90 CSoutput.t21 4.06363
R22110 CSoutput.n90 CSoutput.t64 4.06363
R22111 CSoutput.n92 CSoutput.t37 4.06363
R22112 CSoutput.n92 CSoutput.t55 4.06363
R22113 CSoutput.n44 CSoutput.n43 3.79402
R22114 CSoutput.n49 CSoutput.n48 3.79402
R22115 CSoutput.n371 CSoutput.n355 3.72967
R22116 CSoutput.n419 CSoutput.n403 3.72967
R22117 CSoutput.n421 CSoutput.n420 3.57343
R22118 CSoutput.n420 CSoutput.n372 3.3798
R22119 CSoutput.n369 CSoutput.t112 2.82907
R22120 CSoutput.n369 CSoutput.t119 2.82907
R22121 CSoutput.n367 CSoutput.t105 2.82907
R22122 CSoutput.n367 CSoutput.t185 2.82907
R22123 CSoutput.n365 CSoutput.t154 2.82907
R22124 CSoutput.n365 CSoutput.t97 2.82907
R22125 CSoutput.n363 CSoutput.t188 2.82907
R22126 CSoutput.n363 CSoutput.t174 2.82907
R22127 CSoutput.n361 CSoutput.t135 2.82907
R22128 CSoutput.n361 CSoutput.t144 2.82907
R22129 CSoutput.n359 CSoutput.t96 2.82907
R22130 CSoutput.n359 CSoutput.t181 2.82907
R22131 CSoutput.n357 CSoutput.t175 2.82907
R22132 CSoutput.n357 CSoutput.t121 2.82907
R22133 CSoutput.n356 CSoutput.t107 2.82907
R22134 CSoutput.n356 CSoutput.t187 2.82907
R22135 CSoutput.n353 CSoutput.t120 2.82907
R22136 CSoutput.n353 CSoutput.t191 2.82907
R22137 CSoutput.n351 CSoutput.t103 2.82907
R22138 CSoutput.n351 CSoutput.t186 2.82907
R22139 CSoutput.n349 CSoutput.t114 2.82907
R22140 CSoutput.n349 CSoutput.t130 2.82907
R22141 CSoutput.n347 CSoutput.t128 2.82907
R22142 CSoutput.n347 CSoutput.t106 2.82907
R22143 CSoutput.n345 CSoutput.t141 2.82907
R22144 CSoutput.n345 CSoutput.t115 2.82907
R22145 CSoutput.n343 CSoutput.t116 2.82907
R22146 CSoutput.n343 CSoutput.t129 2.82907
R22147 CSoutput.n341 CSoutput.t127 2.82907
R22148 CSoutput.n341 CSoutput.t139 2.82907
R22149 CSoutput.n340 CSoutput.t140 2.82907
R22150 CSoutput.n340 CSoutput.t117 2.82907
R22151 CSoutput.n338 CSoutput.t108 2.82907
R22152 CSoutput.n338 CSoutput.t123 2.82907
R22153 CSoutput.n336 CSoutput.t145 2.82907
R22154 CSoutput.n336 CSoutput.t173 2.82907
R22155 CSoutput.n334 CSoutput.t163 2.82907
R22156 CSoutput.n334 CSoutput.t132 2.82907
R22157 CSoutput.n332 CSoutput.t101 2.82907
R22158 CSoutput.n332 CSoutput.t149 2.82907
R22159 CSoutput.n330 CSoutput.t131 2.82907
R22160 CSoutput.n330 CSoutput.t142 2.82907
R22161 CSoutput.n328 CSoutput.t143 2.82907
R22162 CSoutput.n328 CSoutput.t180 2.82907
R22163 CSoutput.n326 CSoutput.t159 2.82907
R22164 CSoutput.n326 CSoutput.t98 2.82907
R22165 CSoutput.n325 CSoutput.t177 2.82907
R22166 CSoutput.n325 CSoutput.t109 2.82907
R22167 CSoutput.n404 CSoutput.t169 2.82907
R22168 CSoutput.n404 CSoutput.t184 2.82907
R22169 CSoutput.n405 CSoutput.t189 2.82907
R22170 CSoutput.n405 CSoutput.t158 2.82907
R22171 CSoutput.n407 CSoutput.t162 2.82907
R22172 CSoutput.n407 CSoutput.t178 2.82907
R22173 CSoutput.n409 CSoutput.t110 2.82907
R22174 CSoutput.n409 CSoutput.t152 2.82907
R22175 CSoutput.n411 CSoutput.t157 2.82907
R22176 CSoutput.n411 CSoutput.t170 2.82907
R22177 CSoutput.n413 CSoutput.t179 2.82907
R22178 CSoutput.n413 CSoutput.t161 2.82907
R22179 CSoutput.n415 CSoutput.t166 2.82907
R22180 CSoutput.n415 CSoutput.t183 2.82907
R22181 CSoutput.n417 CSoutput.t111 2.82907
R22182 CSoutput.n417 CSoutput.t122 2.82907
R22183 CSoutput.n388 CSoutput.t137 2.82907
R22184 CSoutput.n388 CSoutput.t155 2.82907
R22185 CSoutput.n389 CSoutput.t156 2.82907
R22186 CSoutput.n389 CSoutput.t146 2.82907
R22187 CSoutput.n391 CSoutput.t147 2.82907
R22188 CSoutput.n391 CSoutput.t138 2.82907
R22189 CSoutput.n393 CSoutput.t133 2.82907
R22190 CSoutput.n393 CSoutput.t125 2.82907
R22191 CSoutput.n395 CSoutput.t126 2.82907
R22192 CSoutput.n395 CSoutput.t148 2.82907
R22193 CSoutput.n397 CSoutput.t150 2.82907
R22194 CSoutput.n397 CSoutput.t99 2.82907
R22195 CSoutput.n399 CSoutput.t100 2.82907
R22196 CSoutput.n399 CSoutput.t118 2.82907
R22197 CSoutput.n401 CSoutput.t124 2.82907
R22198 CSoutput.n401 CSoutput.t113 2.82907
R22199 CSoutput.n373 CSoutput.t151 2.82907
R22200 CSoutput.n373 CSoutput.t102 2.82907
R22201 CSoutput.n374 CSoutput.t134 2.82907
R22202 CSoutput.n374 CSoutput.t182 2.82907
R22203 CSoutput.n376 CSoutput.t104 2.82907
R22204 CSoutput.n376 CSoutput.t165 2.82907
R22205 CSoutput.n378 CSoutput.t164 2.82907
R22206 CSoutput.n378 CSoutput.t153 2.82907
R22207 CSoutput.n380 CSoutput.t168 2.82907
R22208 CSoutput.n380 CSoutput.t136 2.82907
R22209 CSoutput.n382 CSoutput.t160 2.82907
R22210 CSoutput.n382 CSoutput.t176 2.82907
R22211 CSoutput.n384 CSoutput.t190 2.82907
R22212 CSoutput.n384 CSoutput.t167 2.82907
R22213 CSoutput.n386 CSoutput.t172 2.82907
R22214 CSoutput.n386 CSoutput.t171 2.82907
R22215 CSoutput.n324 CSoutput.n126 2.57547
R22216 CSoutput.n75 CSoutput.n1 2.45513
R22217 CSoutput.n217 CSoutput.n215 2.251
R22218 CSoutput.n217 CSoutput.n214 2.251
R22219 CSoutput.n217 CSoutput.n213 2.251
R22220 CSoutput.n217 CSoutput.n212 2.251
R22221 CSoutput.n186 CSoutput.n185 2.251
R22222 CSoutput.n186 CSoutput.n184 2.251
R22223 CSoutput.n186 CSoutput.n183 2.251
R22224 CSoutput.n186 CSoutput.n182 2.251
R22225 CSoutput.n259 CSoutput.n258 2.251
R22226 CSoutput.n224 CSoutput.n222 2.251
R22227 CSoutput.n224 CSoutput.n221 2.251
R22228 CSoutput.n224 CSoutput.n220 2.251
R22229 CSoutput.n242 CSoutput.n224 2.251
R22230 CSoutput.n230 CSoutput.n229 2.251
R22231 CSoutput.n230 CSoutput.n228 2.251
R22232 CSoutput.n230 CSoutput.n227 2.251
R22233 CSoutput.n230 CSoutput.n226 2.251
R22234 CSoutput.n256 CSoutput.n196 2.251
R22235 CSoutput.n251 CSoutput.n249 2.251
R22236 CSoutput.n251 CSoutput.n248 2.251
R22237 CSoutput.n251 CSoutput.n247 2.251
R22238 CSoutput.n251 CSoutput.n246 2.251
R22239 CSoutput.n152 CSoutput.n151 2.251
R22240 CSoutput.n152 CSoutput.n150 2.251
R22241 CSoutput.n152 CSoutput.n149 2.251
R22242 CSoutput.n152 CSoutput.n148 2.251
R22243 CSoutput.n269 CSoutput.n268 2.251
R22244 CSoutput.n186 CSoutput.n166 2.2505
R22245 CSoutput.n181 CSoutput.n166 2.2505
R22246 CSoutput.n179 CSoutput.n166 2.2505
R22247 CSoutput.n178 CSoutput.n166 2.2505
R22248 CSoutput.n263 CSoutput.n166 2.2505
R22249 CSoutput.n261 CSoutput.n166 2.2505
R22250 CSoutput.n259 CSoutput.n166 2.2505
R22251 CSoutput.n189 CSoutput.n166 2.2505
R22252 CSoutput.n188 CSoutput.n166 2.2505
R22253 CSoutput.n192 CSoutput.n166 2.2505
R22254 CSoutput.n191 CSoutput.n166 2.2505
R22255 CSoutput.n174 CSoutput.n166 2.2505
R22256 CSoutput.n266 CSoutput.n166 2.2505
R22257 CSoutput.n266 CSoutput.n265 2.2505
R22258 CSoutput.n230 CSoutput.n201 2.2505
R22259 CSoutput.n211 CSoutput.n201 2.2505
R22260 CSoutput.n232 CSoutput.n201 2.2505
R22261 CSoutput.n210 CSoutput.n201 2.2505
R22262 CSoutput.n234 CSoutput.n201 2.2505
R22263 CSoutput.n201 CSoutput.n195 2.2505
R22264 CSoutput.n256 CSoutput.n201 2.2505
R22265 CSoutput.n254 CSoutput.n201 2.2505
R22266 CSoutput.n236 CSoutput.n201 2.2505
R22267 CSoutput.n208 CSoutput.n201 2.2505
R22268 CSoutput.n238 CSoutput.n201 2.2505
R22269 CSoutput.n207 CSoutput.n201 2.2505
R22270 CSoutput.n252 CSoutput.n201 2.2505
R22271 CSoutput.n252 CSoutput.n205 2.2505
R22272 CSoutput.n152 CSoutput.n132 2.2505
R22273 CSoutput.n147 CSoutput.n132 2.2505
R22274 CSoutput.n145 CSoutput.n132 2.2505
R22275 CSoutput.n144 CSoutput.n132 2.2505
R22276 CSoutput.n273 CSoutput.n132 2.2505
R22277 CSoutput.n271 CSoutput.n132 2.2505
R22278 CSoutput.n269 CSoutput.n132 2.2505
R22279 CSoutput.n155 CSoutput.n132 2.2505
R22280 CSoutput.n154 CSoutput.n132 2.2505
R22281 CSoutput.n158 CSoutput.n132 2.2505
R22282 CSoutput.n157 CSoutput.n132 2.2505
R22283 CSoutput.n140 CSoutput.n132 2.2505
R22284 CSoutput.n276 CSoutput.n132 2.2505
R22285 CSoutput.n276 CSoutput.n275 2.2505
R22286 CSoutput.n194 CSoutput.n187 2.25024
R22287 CSoutput.n194 CSoutput.n180 2.25024
R22288 CSoutput.n262 CSoutput.n194 2.25024
R22289 CSoutput.n194 CSoutput.n190 2.25024
R22290 CSoutput.n194 CSoutput.n193 2.25024
R22291 CSoutput.n194 CSoutput.n161 2.25024
R22292 CSoutput.n244 CSoutput.n241 2.25024
R22293 CSoutput.n244 CSoutput.n240 2.25024
R22294 CSoutput.n244 CSoutput.n239 2.25024
R22295 CSoutput.n244 CSoutput.n206 2.25024
R22296 CSoutput.n244 CSoutput.n243 2.25024
R22297 CSoutput.n245 CSoutput.n244 2.25024
R22298 CSoutput.n160 CSoutput.n153 2.25024
R22299 CSoutput.n160 CSoutput.n146 2.25024
R22300 CSoutput.n272 CSoutput.n160 2.25024
R22301 CSoutput.n160 CSoutput.n156 2.25024
R22302 CSoutput.n160 CSoutput.n159 2.25024
R22303 CSoutput.n160 CSoutput.n127 2.25024
R22304 CSoutput.n261 CSoutput.n171 1.50111
R22305 CSoutput.n209 CSoutput.n195 1.50111
R22306 CSoutput.n271 CSoutput.n137 1.50111
R22307 CSoutput.n217 CSoutput.n216 1.501
R22308 CSoutput.n224 CSoutput.n223 1.501
R22309 CSoutput.n251 CSoutput.n250 1.501
R22310 CSoutput.n265 CSoutput.n176 1.12536
R22311 CSoutput.n265 CSoutput.n177 1.12536
R22312 CSoutput.n265 CSoutput.n264 1.12536
R22313 CSoutput.n225 CSoutput.n205 1.12536
R22314 CSoutput.n231 CSoutput.n205 1.12536
R22315 CSoutput.n233 CSoutput.n205 1.12536
R22316 CSoutput.n275 CSoutput.n142 1.12536
R22317 CSoutput.n275 CSoutput.n143 1.12536
R22318 CSoutput.n275 CSoutput.n274 1.12536
R22319 CSoutput.n265 CSoutput.n172 1.12536
R22320 CSoutput.n265 CSoutput.n173 1.12536
R22321 CSoutput.n265 CSoutput.n175 1.12536
R22322 CSoutput.n255 CSoutput.n205 1.12536
R22323 CSoutput.n235 CSoutput.n205 1.12536
R22324 CSoutput.n237 CSoutput.n205 1.12536
R22325 CSoutput.n275 CSoutput.n138 1.12536
R22326 CSoutput.n275 CSoutput.n139 1.12536
R22327 CSoutput.n275 CSoutput.n141 1.12536
R22328 CSoutput.n31 CSoutput.n30 0.669944
R22329 CSoutput.n62 CSoutput.n61 0.669944
R22330 CSoutput.n360 CSoutput.n358 0.573776
R22331 CSoutput.n362 CSoutput.n360 0.573776
R22332 CSoutput.n364 CSoutput.n362 0.573776
R22333 CSoutput.n366 CSoutput.n364 0.573776
R22334 CSoutput.n368 CSoutput.n366 0.573776
R22335 CSoutput.n370 CSoutput.n368 0.573776
R22336 CSoutput.n344 CSoutput.n342 0.573776
R22337 CSoutput.n346 CSoutput.n344 0.573776
R22338 CSoutput.n348 CSoutput.n346 0.573776
R22339 CSoutput.n350 CSoutput.n348 0.573776
R22340 CSoutput.n352 CSoutput.n350 0.573776
R22341 CSoutput.n354 CSoutput.n352 0.573776
R22342 CSoutput.n329 CSoutput.n327 0.573776
R22343 CSoutput.n331 CSoutput.n329 0.573776
R22344 CSoutput.n333 CSoutput.n331 0.573776
R22345 CSoutput.n335 CSoutput.n333 0.573776
R22346 CSoutput.n337 CSoutput.n335 0.573776
R22347 CSoutput.n339 CSoutput.n337 0.573776
R22348 CSoutput.n418 CSoutput.n416 0.573776
R22349 CSoutput.n416 CSoutput.n414 0.573776
R22350 CSoutput.n414 CSoutput.n412 0.573776
R22351 CSoutput.n412 CSoutput.n410 0.573776
R22352 CSoutput.n410 CSoutput.n408 0.573776
R22353 CSoutput.n408 CSoutput.n406 0.573776
R22354 CSoutput.n402 CSoutput.n400 0.573776
R22355 CSoutput.n400 CSoutput.n398 0.573776
R22356 CSoutput.n398 CSoutput.n396 0.573776
R22357 CSoutput.n396 CSoutput.n394 0.573776
R22358 CSoutput.n394 CSoutput.n392 0.573776
R22359 CSoutput.n392 CSoutput.n390 0.573776
R22360 CSoutput.n387 CSoutput.n385 0.573776
R22361 CSoutput.n385 CSoutput.n383 0.573776
R22362 CSoutput.n383 CSoutput.n381 0.573776
R22363 CSoutput.n381 CSoutput.n379 0.573776
R22364 CSoutput.n379 CSoutput.n377 0.573776
R22365 CSoutput.n377 CSoutput.n375 0.573776
R22366 CSoutput.n421 CSoutput.n276 0.53442
R22367 CSoutput.n312 CSoutput.n310 0.358259
R22368 CSoutput.n314 CSoutput.n312 0.358259
R22369 CSoutput.n316 CSoutput.n314 0.358259
R22370 CSoutput.n318 CSoutput.n316 0.358259
R22371 CSoutput.n320 CSoutput.n318 0.358259
R22372 CSoutput.n322 CSoutput.n320 0.358259
R22373 CSoutput.n296 CSoutput.n294 0.358259
R22374 CSoutput.n298 CSoutput.n296 0.358259
R22375 CSoutput.n300 CSoutput.n298 0.358259
R22376 CSoutput.n302 CSoutput.n300 0.358259
R22377 CSoutput.n304 CSoutput.n302 0.358259
R22378 CSoutput.n306 CSoutput.n304 0.358259
R22379 CSoutput.n281 CSoutput.n279 0.358259
R22380 CSoutput.n283 CSoutput.n281 0.358259
R22381 CSoutput.n285 CSoutput.n283 0.358259
R22382 CSoutput.n287 CSoutput.n285 0.358259
R22383 CSoutput.n289 CSoutput.n287 0.358259
R22384 CSoutput.n291 CSoutput.n289 0.358259
R22385 CSoutput.n124 CSoutput.n122 0.358259
R22386 CSoutput.n122 CSoutput.n120 0.358259
R22387 CSoutput.n120 CSoutput.n118 0.358259
R22388 CSoutput.n118 CSoutput.n116 0.358259
R22389 CSoutput.n116 CSoutput.n114 0.358259
R22390 CSoutput.n114 CSoutput.n112 0.358259
R22391 CSoutput.n108 CSoutput.n106 0.358259
R22392 CSoutput.n106 CSoutput.n104 0.358259
R22393 CSoutput.n104 CSoutput.n102 0.358259
R22394 CSoutput.n102 CSoutput.n100 0.358259
R22395 CSoutput.n100 CSoutput.n98 0.358259
R22396 CSoutput.n98 CSoutput.n96 0.358259
R22397 CSoutput.n93 CSoutput.n91 0.358259
R22398 CSoutput.n91 CSoutput.n89 0.358259
R22399 CSoutput.n89 CSoutput.n87 0.358259
R22400 CSoutput.n87 CSoutput.n85 0.358259
R22401 CSoutput.n85 CSoutput.n83 0.358259
R22402 CSoutput.n83 CSoutput.n81 0.358259
R22403 CSoutput.n21 CSoutput.n20 0.169105
R22404 CSoutput.n21 CSoutput.n16 0.169105
R22405 CSoutput.n26 CSoutput.n16 0.169105
R22406 CSoutput.n27 CSoutput.n26 0.169105
R22407 CSoutput.n27 CSoutput.n14 0.169105
R22408 CSoutput.n32 CSoutput.n14 0.169105
R22409 CSoutput.n33 CSoutput.n32 0.169105
R22410 CSoutput.n34 CSoutput.n33 0.169105
R22411 CSoutput.n34 CSoutput.n12 0.169105
R22412 CSoutput.n39 CSoutput.n12 0.169105
R22413 CSoutput.n40 CSoutput.n39 0.169105
R22414 CSoutput.n40 CSoutput.n10 0.169105
R22415 CSoutput.n45 CSoutput.n10 0.169105
R22416 CSoutput.n46 CSoutput.n45 0.169105
R22417 CSoutput.n47 CSoutput.n46 0.169105
R22418 CSoutput.n47 CSoutput.n8 0.169105
R22419 CSoutput.n52 CSoutput.n8 0.169105
R22420 CSoutput.n53 CSoutput.n52 0.169105
R22421 CSoutput.n53 CSoutput.n6 0.169105
R22422 CSoutput.n58 CSoutput.n6 0.169105
R22423 CSoutput.n59 CSoutput.n58 0.169105
R22424 CSoutput.n60 CSoutput.n59 0.169105
R22425 CSoutput.n60 CSoutput.n4 0.169105
R22426 CSoutput.n66 CSoutput.n4 0.169105
R22427 CSoutput.n67 CSoutput.n66 0.169105
R22428 CSoutput.n68 CSoutput.n67 0.169105
R22429 CSoutput.n68 CSoutput.n2 0.169105
R22430 CSoutput.n73 CSoutput.n2 0.169105
R22431 CSoutput.n74 CSoutput.n73 0.169105
R22432 CSoutput.n74 CSoutput.n0 0.169105
R22433 CSoutput.n78 CSoutput.n0 0.169105
R22434 CSoutput.n219 CSoutput.n218 0.0910737
R22435 CSoutput.n270 CSoutput.n267 0.0723685
R22436 CSoutput.n224 CSoutput.n219 0.0522944
R22437 CSoutput.n267 CSoutput.n266 0.0499135
R22438 CSoutput.n218 CSoutput.n217 0.0499135
R22439 CSoutput.n252 CSoutput.n251 0.0464294
R22440 CSoutput.n260 CSoutput.n257 0.0391444
R22441 CSoutput.n219 CSoutput.t212 0.023435
R22442 CSoutput.n267 CSoutput.t204 0.02262
R22443 CSoutput.n218 CSoutput.t193 0.02262
R22444 CSoutput CSoutput.n421 0.0052
R22445 CSoutput.n189 CSoutput.n172 0.00365111
R22446 CSoutput.n192 CSoutput.n173 0.00365111
R22447 CSoutput.n175 CSoutput.n174 0.00365111
R22448 CSoutput.n217 CSoutput.n176 0.00365111
R22449 CSoutput.n181 CSoutput.n177 0.00365111
R22450 CSoutput.n264 CSoutput.n178 0.00365111
R22451 CSoutput.n255 CSoutput.n254 0.00365111
R22452 CSoutput.n235 CSoutput.n208 0.00365111
R22453 CSoutput.n237 CSoutput.n207 0.00365111
R22454 CSoutput.n225 CSoutput.n224 0.00365111
R22455 CSoutput.n231 CSoutput.n211 0.00365111
R22456 CSoutput.n233 CSoutput.n210 0.00365111
R22457 CSoutput.n155 CSoutput.n138 0.00365111
R22458 CSoutput.n158 CSoutput.n139 0.00365111
R22459 CSoutput.n141 CSoutput.n140 0.00365111
R22460 CSoutput.n251 CSoutput.n142 0.00365111
R22461 CSoutput.n147 CSoutput.n143 0.00365111
R22462 CSoutput.n274 CSoutput.n144 0.00365111
R22463 CSoutput.n186 CSoutput.n176 0.00340054
R22464 CSoutput.n179 CSoutput.n177 0.00340054
R22465 CSoutput.n264 CSoutput.n263 0.00340054
R22466 CSoutput.n259 CSoutput.n172 0.00340054
R22467 CSoutput.n188 CSoutput.n173 0.00340054
R22468 CSoutput.n191 CSoutput.n175 0.00340054
R22469 CSoutput.n230 CSoutput.n225 0.00340054
R22470 CSoutput.n232 CSoutput.n231 0.00340054
R22471 CSoutput.n234 CSoutput.n233 0.00340054
R22472 CSoutput.n256 CSoutput.n255 0.00340054
R22473 CSoutput.n236 CSoutput.n235 0.00340054
R22474 CSoutput.n238 CSoutput.n237 0.00340054
R22475 CSoutput.n152 CSoutput.n142 0.00340054
R22476 CSoutput.n145 CSoutput.n143 0.00340054
R22477 CSoutput.n274 CSoutput.n273 0.00340054
R22478 CSoutput.n269 CSoutput.n138 0.00340054
R22479 CSoutput.n154 CSoutput.n139 0.00340054
R22480 CSoutput.n157 CSoutput.n141 0.00340054
R22481 CSoutput.n187 CSoutput.n181 0.00252698
R22482 CSoutput.n180 CSoutput.n178 0.00252698
R22483 CSoutput.n262 CSoutput.n261 0.00252698
R22484 CSoutput.n190 CSoutput.n188 0.00252698
R22485 CSoutput.n193 CSoutput.n191 0.00252698
R22486 CSoutput.n266 CSoutput.n161 0.00252698
R22487 CSoutput.n187 CSoutput.n186 0.00252698
R22488 CSoutput.n180 CSoutput.n179 0.00252698
R22489 CSoutput.n263 CSoutput.n262 0.00252698
R22490 CSoutput.n190 CSoutput.n189 0.00252698
R22491 CSoutput.n193 CSoutput.n192 0.00252698
R22492 CSoutput.n174 CSoutput.n161 0.00252698
R22493 CSoutput.n241 CSoutput.n211 0.00252698
R22494 CSoutput.n240 CSoutput.n210 0.00252698
R22495 CSoutput.n239 CSoutput.n195 0.00252698
R22496 CSoutput.n236 CSoutput.n206 0.00252698
R22497 CSoutput.n243 CSoutput.n238 0.00252698
R22498 CSoutput.n252 CSoutput.n245 0.00252698
R22499 CSoutput.n241 CSoutput.n230 0.00252698
R22500 CSoutput.n240 CSoutput.n232 0.00252698
R22501 CSoutput.n239 CSoutput.n234 0.00252698
R22502 CSoutput.n254 CSoutput.n206 0.00252698
R22503 CSoutput.n243 CSoutput.n208 0.00252698
R22504 CSoutput.n245 CSoutput.n207 0.00252698
R22505 CSoutput.n153 CSoutput.n147 0.00252698
R22506 CSoutput.n146 CSoutput.n144 0.00252698
R22507 CSoutput.n272 CSoutput.n271 0.00252698
R22508 CSoutput.n156 CSoutput.n154 0.00252698
R22509 CSoutput.n159 CSoutput.n157 0.00252698
R22510 CSoutput.n276 CSoutput.n127 0.00252698
R22511 CSoutput.n153 CSoutput.n152 0.00252698
R22512 CSoutput.n146 CSoutput.n145 0.00252698
R22513 CSoutput.n273 CSoutput.n272 0.00252698
R22514 CSoutput.n156 CSoutput.n155 0.00252698
R22515 CSoutput.n159 CSoutput.n158 0.00252698
R22516 CSoutput.n140 CSoutput.n127 0.00252698
R22517 CSoutput.n261 CSoutput.n260 0.0020275
R22518 CSoutput.n260 CSoutput.n259 0.0020275
R22519 CSoutput.n257 CSoutput.n195 0.0020275
R22520 CSoutput.n257 CSoutput.n256 0.0020275
R22521 CSoutput.n271 CSoutput.n270 0.0020275
R22522 CSoutput.n270 CSoutput.n269 0.0020275
R22523 CSoutput.n171 CSoutput.n170 0.00166668
R22524 CSoutput.n253 CSoutput.n209 0.00166668
R22525 CSoutput.n137 CSoutput.n136 0.00166668
R22526 CSoutput.n275 CSoutput.n137 0.00133328
R22527 CSoutput.n209 CSoutput.n205 0.00133328
R22528 CSoutput.n265 CSoutput.n171 0.00133328
R22529 CSoutput.n268 CSoutput.n160 0.001
R22530 CSoutput.n246 CSoutput.n160 0.001
R22531 CSoutput.n148 CSoutput.n128 0.001
R22532 CSoutput.n247 CSoutput.n128 0.001
R22533 CSoutput.n149 CSoutput.n129 0.001
R22534 CSoutput.n248 CSoutput.n129 0.001
R22535 CSoutput.n150 CSoutput.n130 0.001
R22536 CSoutput.n249 CSoutput.n130 0.001
R22537 CSoutput.n151 CSoutput.n131 0.001
R22538 CSoutput.n250 CSoutput.n131 0.001
R22539 CSoutput.n244 CSoutput.n196 0.001
R22540 CSoutput.n244 CSoutput.n242 0.001
R22541 CSoutput.n226 CSoutput.n197 0.001
R22542 CSoutput.n220 CSoutput.n197 0.001
R22543 CSoutput.n227 CSoutput.n198 0.001
R22544 CSoutput.n221 CSoutput.n198 0.001
R22545 CSoutput.n228 CSoutput.n199 0.001
R22546 CSoutput.n222 CSoutput.n199 0.001
R22547 CSoutput.n229 CSoutput.n200 0.001
R22548 CSoutput.n223 CSoutput.n200 0.001
R22549 CSoutput.n258 CSoutput.n194 0.001
R22550 CSoutput.n212 CSoutput.n194 0.001
R22551 CSoutput.n182 CSoutput.n162 0.001
R22552 CSoutput.n213 CSoutput.n162 0.001
R22553 CSoutput.n183 CSoutput.n163 0.001
R22554 CSoutput.n214 CSoutput.n163 0.001
R22555 CSoutput.n184 CSoutput.n164 0.001
R22556 CSoutput.n215 CSoutput.n164 0.001
R22557 CSoutput.n185 CSoutput.n165 0.001
R22558 CSoutput.n216 CSoutput.n165 0.001
R22559 CSoutput.n216 CSoutput.n166 0.001
R22560 CSoutput.n215 CSoutput.n167 0.001
R22561 CSoutput.n214 CSoutput.n168 0.001
R22562 CSoutput.n213 CSoutput.t209 0.001
R22563 CSoutput.n212 CSoutput.n169 0.001
R22564 CSoutput.n185 CSoutput.n167 0.001
R22565 CSoutput.n184 CSoutput.n168 0.001
R22566 CSoutput.n183 CSoutput.t209 0.001
R22567 CSoutput.n182 CSoutput.n169 0.001
R22568 CSoutput.n258 CSoutput.n170 0.001
R22569 CSoutput.n223 CSoutput.n201 0.001
R22570 CSoutput.n222 CSoutput.n202 0.001
R22571 CSoutput.n221 CSoutput.n203 0.001
R22572 CSoutput.n220 CSoutput.t202 0.001
R22573 CSoutput.n242 CSoutput.n204 0.001
R22574 CSoutput.n229 CSoutput.n202 0.001
R22575 CSoutput.n228 CSoutput.n203 0.001
R22576 CSoutput.n227 CSoutput.t202 0.001
R22577 CSoutput.n226 CSoutput.n204 0.001
R22578 CSoutput.n253 CSoutput.n196 0.001
R22579 CSoutput.n250 CSoutput.n132 0.001
R22580 CSoutput.n249 CSoutput.n133 0.001
R22581 CSoutput.n248 CSoutput.n134 0.001
R22582 CSoutput.n247 CSoutput.t192 0.001
R22583 CSoutput.n246 CSoutput.n135 0.001
R22584 CSoutput.n151 CSoutput.n133 0.001
R22585 CSoutput.n150 CSoutput.n134 0.001
R22586 CSoutput.n149 CSoutput.t192 0.001
R22587 CSoutput.n148 CSoutput.n135 0.001
R22588 CSoutput.n268 CSoutput.n136 0.001
R22589 a_n2318_13878.n57 a_n2318_13878.t31 533.335
R22590 a_n2318_13878.n112 a_n2318_13878.t15 512.366
R22591 a_n2318_13878.n64 a_n2318_13878.t17 512.366
R22592 a_n2318_13878.n111 a_n2318_13878.t27 512.366
R22593 a_n2318_13878.n110 a_n2318_13878.t3 512.366
R22594 a_n2318_13878.n65 a_n2318_13878.t9 512.366
R22595 a_n2318_13878.n109 a_n2318_13878.t5 512.366
R22596 a_n2318_13878.n51 a_n2318_13878.t78 533.335
R22597 a_n2318_13878.n108 a_n2318_13878.t59 512.366
R22598 a_n2318_13878.n74 a_n2318_13878.t63 512.366
R22599 a_n2318_13878.n107 a_n2318_13878.t53 512.366
R22600 a_n2318_13878.n106 a_n2318_13878.t68 512.366
R22601 a_n2318_13878.n75 a_n2318_13878.t75 512.366
R22602 a_n2318_13878.n105 a_n2318_13878.t76 512.366
R22603 a_n2318_13878.n36 a_n2318_13878.t11 533.335
R22604 a_n2318_13878.n86 a_n2318_13878.t7 512.366
R22605 a_n2318_13878.n87 a_n2318_13878.t13 512.366
R22606 a_n2318_13878.n88 a_n2318_13878.t21 512.366
R22607 a_n2318_13878.n89 a_n2318_13878.t33 512.366
R22608 a_n2318_13878.n79 a_n2318_13878.t29 512.366
R22609 a_n2318_13878.n90 a_n2318_13878.t19 512.366
R22610 a_n2318_13878.n29 a_n2318_13878.t74 533.335
R22611 a_n2318_13878.n81 a_n2318_13878.t52 512.366
R22612 a_n2318_13878.n82 a_n2318_13878.t71 512.366
R22613 a_n2318_13878.n83 a_n2318_13878.t72 512.366
R22614 a_n2318_13878.n84 a_n2318_13878.t49 512.366
R22615 a_n2318_13878.n80 a_n2318_13878.t58 512.366
R22616 a_n2318_13878.n85 a_n2318_13878.t67 512.366
R22617 a_n2318_13878.n102 a_n2318_13878.t65 512.366
R22618 a_n2318_13878.n92 a_n2318_13878.t56 512.366
R22619 a_n2318_13878.n103 a_n2318_13878.t48 512.366
R22620 a_n2318_13878.n100 a_n2318_13878.t73 512.366
R22621 a_n2318_13878.n93 a_n2318_13878.t62 512.366
R22622 a_n2318_13878.n101 a_n2318_13878.t61 512.366
R22623 a_n2318_13878.n98 a_n2318_13878.t69 512.366
R22624 a_n2318_13878.n94 a_n2318_13878.t54 512.366
R22625 a_n2318_13878.n99 a_n2318_13878.t55 512.366
R22626 a_n2318_13878.n96 a_n2318_13878.t57 512.366
R22627 a_n2318_13878.n95 a_n2318_13878.t66 512.366
R22628 a_n2318_13878.n97 a_n2318_13878.t79 512.366
R22629 a_n2318_13878.n63 a_n2318_13878.n28 70.1674
R22630 a_n2318_13878.n56 a_n2318_13878.n6 70.1674
R22631 a_n2318_13878.n18 a_n2318_13878.n42 70.1674
R22632 a_n2318_13878.n21 a_n2318_13878.n35 70.1674
R22633 a_n2318_13878.n85 a_n2318_13878.n35 20.9683
R22634 a_n2318_13878.n34 a_n2318_13878.n22 72.3034
R22635 a_n2318_13878.n34 a_n2318_13878.n80 16.6962
R22636 a_n2318_13878.n22 a_n2318_13878.n33 77.6622
R22637 a_n2318_13878.n84 a_n2318_13878.n33 5.97853
R22638 a_n2318_13878.n32 a_n2318_13878.n23 77.6622
R22639 a_n2318_13878.n23 a_n2318_13878.n31 72.3034
R22640 a_n2318_13878.n81 a_n2318_13878.n29 20.9683
R22641 a_n2318_13878.n30 a_n2318_13878.n29 70.1674
R22642 a_n2318_13878.n90 a_n2318_13878.n42 20.9683
R22643 a_n2318_13878.n41 a_n2318_13878.n19 72.3034
R22644 a_n2318_13878.n41 a_n2318_13878.n79 16.6962
R22645 a_n2318_13878.n19 a_n2318_13878.n40 77.6622
R22646 a_n2318_13878.n89 a_n2318_13878.n40 5.97853
R22647 a_n2318_13878.n39 a_n2318_13878.n20 77.6622
R22648 a_n2318_13878.n20 a_n2318_13878.n38 72.3034
R22649 a_n2318_13878.n86 a_n2318_13878.n36 20.9683
R22650 a_n2318_13878.n37 a_n2318_13878.n36 70.1674
R22651 a_n2318_13878.n9 a_n2318_13878.n50 70.1674
R22652 a_n2318_13878.n11 a_n2318_13878.n48 70.1674
R22653 a_n2318_13878.n13 a_n2318_13878.n46 70.1674
R22654 a_n2318_13878.n16 a_n2318_13878.n44 70.1674
R22655 a_n2318_13878.n97 a_n2318_13878.n44 20.9683
R22656 a_n2318_13878.n43 a_n2318_13878.n17 75.0448
R22657 a_n2318_13878.n43 a_n2318_13878.n95 11.2134
R22658 a_n2318_13878.n17 a_n2318_13878.n96 161.3
R22659 a_n2318_13878.n99 a_n2318_13878.n46 20.9683
R22660 a_n2318_13878.n45 a_n2318_13878.n14 75.0448
R22661 a_n2318_13878.n45 a_n2318_13878.n94 11.2134
R22662 a_n2318_13878.n14 a_n2318_13878.n98 161.3
R22663 a_n2318_13878.n101 a_n2318_13878.n48 20.9683
R22664 a_n2318_13878.n47 a_n2318_13878.n12 75.0448
R22665 a_n2318_13878.n47 a_n2318_13878.n93 11.2134
R22666 a_n2318_13878.n12 a_n2318_13878.n100 161.3
R22667 a_n2318_13878.n103 a_n2318_13878.n50 20.9683
R22668 a_n2318_13878.n49 a_n2318_13878.n10 75.0448
R22669 a_n2318_13878.n49 a_n2318_13878.n92 11.2134
R22670 a_n2318_13878.n10 a_n2318_13878.n102 161.3
R22671 a_n2318_13878.n105 a_n2318_13878.n56 20.9683
R22672 a_n2318_13878.n7 a_n2318_13878.n55 72.3034
R22673 a_n2318_13878.n55 a_n2318_13878.n75 16.6962
R22674 a_n2318_13878.n54 a_n2318_13878.n7 77.6622
R22675 a_n2318_13878.n106 a_n2318_13878.n54 5.97853
R22676 a_n2318_13878.n53 a_n2318_13878.n5 77.6622
R22677 a_n2318_13878.n5 a_n2318_13878.n52 72.3034
R22678 a_n2318_13878.n108 a_n2318_13878.n51 20.9683
R22679 a_n2318_13878.n8 a_n2318_13878.n51 70.1674
R22680 a_n2318_13878.n109 a_n2318_13878.n63 20.9683
R22681 a_n2318_13878.n28 a_n2318_13878.n62 72.3034
R22682 a_n2318_13878.n62 a_n2318_13878.n65 16.6962
R22683 a_n2318_13878.n61 a_n2318_13878.n60 77.6622
R22684 a_n2318_13878.n110 a_n2318_13878.n61 5.97853
R22685 a_n2318_13878.n59 a_n2318_13878.n4 77.6622
R22686 a_n2318_13878.n4 a_n2318_13878.n58 72.3034
R22687 a_n2318_13878.n112 a_n2318_13878.n57 20.9683
R22688 a_n2318_13878.n3 a_n2318_13878.n57 70.1674
R22689 a_n2318_13878.n1 a_n2318_13878.n72 81.4626
R22690 a_n2318_13878.n2 a_n2318_13878.n68 81.4626
R22691 a_n2318_13878.n2 a_n2318_13878.n66 81.4626
R22692 a_n2318_13878.n1 a_n2318_13878.n73 80.9324
R22693 a_n2318_13878.n1 a_n2318_13878.n71 80.9324
R22694 a_n2318_13878.n0 a_n2318_13878.n70 80.9324
R22695 a_n2318_13878.n2 a_n2318_13878.n69 80.9324
R22696 a_n2318_13878.n2 a_n2318_13878.n67 80.9324
R22697 a_n2318_13878.n27 a_n2318_13878.t26 74.6477
R22698 a_n2318_13878.n24 a_n2318_13878.t12 74.6477
R22699 a_n2318_13878.n26 a_n2318_13878.t32 74.2899
R22700 a_n2318_13878.n25 a_n2318_13878.t24 74.2897
R22701 a_n2318_13878.n27 a_n2318_13878.n115 70.6783
R22702 a_n2318_13878.n26 a_n2318_13878.n114 70.6783
R22703 a_n2318_13878.n25 a_n2318_13878.n78 70.6783
R22704 a_n2318_13878.n24 a_n2318_13878.n77 70.6783
R22705 a_n2318_13878.n24 a_n2318_13878.n76 70.6783
R22706 a_n2318_13878.n116 a_n2318_13878.n27 70.6782
R22707 a_n2318_13878.n111 a_n2318_13878.n110 48.2005
R22708 a_n2318_13878.n63 a_n2318_13878.t25 533.335
R22709 a_n2318_13878.n107 a_n2318_13878.n106 48.2005
R22710 a_n2318_13878.n56 a_n2318_13878.t50 533.335
R22711 a_n2318_13878.n89 a_n2318_13878.n88 48.2005
R22712 a_n2318_13878.t23 a_n2318_13878.n42 533.335
R22713 a_n2318_13878.n84 a_n2318_13878.n83 48.2005
R22714 a_n2318_13878.t51 a_n2318_13878.n35 533.335
R22715 a_n2318_13878.n102 a_n2318_13878.n92 48.2005
R22716 a_n2318_13878.t70 a_n2318_13878.n50 533.335
R22717 a_n2318_13878.n100 a_n2318_13878.n93 48.2005
R22718 a_n2318_13878.t77 a_n2318_13878.n48 533.335
R22719 a_n2318_13878.n98 a_n2318_13878.n94 48.2005
R22720 a_n2318_13878.t64 a_n2318_13878.n46 533.335
R22721 a_n2318_13878.n96 a_n2318_13878.n95 48.2005
R22722 a_n2318_13878.t60 a_n2318_13878.n44 533.335
R22723 a_n2318_13878.n58 a_n2318_13878.n64 16.6962
R22724 a_n2318_13878.n109 a_n2318_13878.n62 27.6507
R22725 a_n2318_13878.n52 a_n2318_13878.n74 16.6962
R22726 a_n2318_13878.n105 a_n2318_13878.n55 27.6507
R22727 a_n2318_13878.n87 a_n2318_13878.n38 16.6962
R22728 a_n2318_13878.n90 a_n2318_13878.n41 27.6507
R22729 a_n2318_13878.n82 a_n2318_13878.n31 16.6962
R22730 a_n2318_13878.n85 a_n2318_13878.n34 27.6507
R22731 a_n2318_13878.n59 a_n2318_13878.n64 41.7634
R22732 a_n2318_13878.n53 a_n2318_13878.n74 41.7634
R22733 a_n2318_13878.n87 a_n2318_13878.n39 41.7634
R22734 a_n2318_13878.n82 a_n2318_13878.n32 41.7634
R22735 a_n2318_13878.n103 a_n2318_13878.n49 35.3134
R22736 a_n2318_13878.n101 a_n2318_13878.n47 35.3134
R22737 a_n2318_13878.n99 a_n2318_13878.n45 35.3134
R22738 a_n2318_13878.n97 a_n2318_13878.n43 35.3134
R22739 a_n2318_13878.n28 a_n2318_13878.n1 23.891
R22740 a_n2318_13878.n30 a_n2318_13878.n15 12.705
R22741 a_n2318_13878.n6 a_n2318_13878.n104 12.5005
R22742 a_n2318_13878.n59 a_n2318_13878.n111 5.97853
R22743 a_n2318_13878.n61 a_n2318_13878.n65 41.7634
R22744 a_n2318_13878.n53 a_n2318_13878.n107 5.97853
R22745 a_n2318_13878.n54 a_n2318_13878.n75 41.7634
R22746 a_n2318_13878.n88 a_n2318_13878.n39 5.97853
R22747 a_n2318_13878.n79 a_n2318_13878.n40 41.7634
R22748 a_n2318_13878.n83 a_n2318_13878.n32 5.97853
R22749 a_n2318_13878.n80 a_n2318_13878.n33 41.7634
R22750 a_n2318_13878.n0 a_n2318_13878.n2 32.5247
R22751 a_n2318_13878.n113 a_n2318_13878.n3 11.1956
R22752 a_n2318_13878.n112 a_n2318_13878.n58 27.6507
R22753 a_n2318_13878.n108 a_n2318_13878.n52 27.6507
R22754 a_n2318_13878.n38 a_n2318_13878.n86 27.6507
R22755 a_n2318_13878.n31 a_n2318_13878.n81 27.6507
R22756 a_n2318_13878.n91 a_n2318_13878.n25 9.85898
R22757 a_n2318_13878.n17 a_n2318_13878.n15 8.73345
R22758 a_n2318_13878.n104 a_n2318_13878.n9 8.73345
R22759 a_n2318_13878.n91 a_n2318_13878.n18 7.36035
R22760 a_n2318_13878.n26 a_n2318_13878.n113 6.01559
R22761 a_n2318_13878.n104 a_n2318_13878.n91 5.3452
R22762 a_n2318_13878.n37 a_n2318_13878.n21 4.01186
R22763 a_n2318_13878.n28 a_n2318_13878.n8 4.0079
R22764 a_n2318_13878.n115 a_n2318_13878.t10 3.61217
R22765 a_n2318_13878.n115 a_n2318_13878.t6 3.61217
R22766 a_n2318_13878.n114 a_n2318_13878.t16 3.61217
R22767 a_n2318_13878.n114 a_n2318_13878.t18 3.61217
R22768 a_n2318_13878.n78 a_n2318_13878.t30 3.61217
R22769 a_n2318_13878.n78 a_n2318_13878.t20 3.61217
R22770 a_n2318_13878.n77 a_n2318_13878.t22 3.61217
R22771 a_n2318_13878.n77 a_n2318_13878.t34 3.61217
R22772 a_n2318_13878.n76 a_n2318_13878.t8 3.61217
R22773 a_n2318_13878.n76 a_n2318_13878.t14 3.61217
R22774 a_n2318_13878.n116 a_n2318_13878.t28 3.61217
R22775 a_n2318_13878.t4 a_n2318_13878.n116 3.61217
R22776 a_n2318_13878.n72 a_n2318_13878.t41 2.82907
R22777 a_n2318_13878.n72 a_n2318_13878.t44 2.82907
R22778 a_n2318_13878.n73 a_n2318_13878.t43 2.82907
R22779 a_n2318_13878.n73 a_n2318_13878.t47 2.82907
R22780 a_n2318_13878.n71 a_n2318_13878.t38 2.82907
R22781 a_n2318_13878.n71 a_n2318_13878.t2 2.82907
R22782 a_n2318_13878.n70 a_n2318_13878.t36 2.82907
R22783 a_n2318_13878.n70 a_n2318_13878.t42 2.82907
R22784 a_n2318_13878.n68 a_n2318_13878.t0 2.82907
R22785 a_n2318_13878.n68 a_n2318_13878.t39 2.82907
R22786 a_n2318_13878.n69 a_n2318_13878.t40 2.82907
R22787 a_n2318_13878.n69 a_n2318_13878.t35 2.82907
R22788 a_n2318_13878.n67 a_n2318_13878.t46 2.82907
R22789 a_n2318_13878.n67 a_n2318_13878.t45 2.82907
R22790 a_n2318_13878.n66 a_n2318_13878.t1 2.82907
R22791 a_n2318_13878.n66 a_n2318_13878.t37 2.82907
R22792 a_n2318_13878.n113 a_n2318_13878.n15 1.30542
R22793 a_n2318_13878.n27 a_n2318_13878.n26 1.07378
R22794 a_n2318_13878.n25 a_n2318_13878.n24 1.07378
R22795 a_n2318_13878.n1 a_n2318_13878.n0 1.06084
R22796 a_n2318_13878.n12 a_n2318_13878.n13 1.04595
R22797 a_n2318_13878.n23 a_n2318_13878.n22 0.758076
R22798 a_n2318_13878.n22 a_n2318_13878.n21 0.758076
R22799 a_n2318_13878.n20 a_n2318_13878.n19 0.758076
R22800 a_n2318_13878.n19 a_n2318_13878.n18 0.758076
R22801 a_n2318_13878.n17 a_n2318_13878.n16 0.758076
R22802 a_n2318_13878.n14 a_n2318_13878.n13 0.758076
R22803 a_n2318_13878.n12 a_n2318_13878.n11 0.758076
R22804 a_n2318_13878.n10 a_n2318_13878.n9 0.758076
R22805 a_n2318_13878.n7 a_n2318_13878.n5 0.758076
R22806 a_n2318_13878.n7 a_n2318_13878.n6 0.758076
R22807 a_n2318_13878.n60 a_n2318_13878.n4 0.758076
R22808 a_n2318_13878.n60 a_n2318_13878.n28 0.724161
R22809 a_n2318_13878.n14 a_n2318_13878.n16 0.67853
R22810 a_n2318_13878.n10 a_n2318_13878.n11 0.67853
R22811 a_n2318_13878.n4 a_n2318_13878.n3 0.568682
R22812 a_n2318_13878.n5 a_n2318_13878.n8 0.568682
R22813 a_n2318_13878.n37 a_n2318_13878.n20 0.568682
R22814 a_n2318_13878.n30 a_n2318_13878.n23 0.568682
R22815 a_n2140_13878.n21 a_n2140_13878.n20 98.9632
R22816 a_n2140_13878.n2 a_n2140_13878.n0 98.7517
R22817 a_n2140_13878.n18 a_n2140_13878.n17 98.6055
R22818 a_n2140_13878.n20 a_n2140_13878.n19 98.6055
R22819 a_n2140_13878.n6 a_n2140_13878.n5 98.6055
R22820 a_n2140_13878.n4 a_n2140_13878.n3 98.6055
R22821 a_n2140_13878.n2 a_n2140_13878.n1 98.6055
R22822 a_n2140_13878.n16 a_n2140_13878.n15 98.6054
R22823 a_n2140_13878.n8 a_n2140_13878.t17 74.6477
R22824 a_n2140_13878.n13 a_n2140_13878.t18 74.2899
R22825 a_n2140_13878.n10 a_n2140_13878.t19 74.2899
R22826 a_n2140_13878.n9 a_n2140_13878.t16 74.2899
R22827 a_n2140_13878.n12 a_n2140_13878.n11 70.6783
R22828 a_n2140_13878.n8 a_n2140_13878.n7 70.6783
R22829 a_n2140_13878.n14 a_n2140_13878.n6 14.2849
R22830 a_n2140_13878.n16 a_n2140_13878.n14 11.9339
R22831 a_n2140_13878.n14 a_n2140_13878.n13 6.95632
R22832 a_n2140_13878.n15 a_n2140_13878.t6 3.61217
R22833 a_n2140_13878.n15 a_n2140_13878.t7 3.61217
R22834 a_n2140_13878.n17 a_n2140_13878.t13 3.61217
R22835 a_n2140_13878.n17 a_n2140_13878.t14 3.61217
R22836 a_n2140_13878.n19 a_n2140_13878.t0 3.61217
R22837 a_n2140_13878.n19 a_n2140_13878.t8 3.61217
R22838 a_n2140_13878.n11 a_n2140_13878.t22 3.61217
R22839 a_n2140_13878.n11 a_n2140_13878.t23 3.61217
R22840 a_n2140_13878.n7 a_n2140_13878.t20 3.61217
R22841 a_n2140_13878.n7 a_n2140_13878.t21 3.61217
R22842 a_n2140_13878.n5 a_n2140_13878.t9 3.61217
R22843 a_n2140_13878.n5 a_n2140_13878.t1 3.61217
R22844 a_n2140_13878.n3 a_n2140_13878.t12 3.61217
R22845 a_n2140_13878.n3 a_n2140_13878.t3 3.61217
R22846 a_n2140_13878.n1 a_n2140_13878.t2 3.61217
R22847 a_n2140_13878.n1 a_n2140_13878.t4 3.61217
R22848 a_n2140_13878.n0 a_n2140_13878.t10 3.61217
R22849 a_n2140_13878.n0 a_n2140_13878.t5 3.61217
R22850 a_n2140_13878.n21 a_n2140_13878.t11 3.61217
R22851 a_n2140_13878.t15 a_n2140_13878.n21 3.61217
R22852 a_n2140_13878.n9 a_n2140_13878.n8 0.358259
R22853 a_n2140_13878.n12 a_n2140_13878.n10 0.358259
R22854 a_n2140_13878.n13 a_n2140_13878.n12 0.358259
R22855 a_n2140_13878.n20 a_n2140_13878.n18 0.358259
R22856 a_n2140_13878.n18 a_n2140_13878.n16 0.358259
R22857 a_n2140_13878.n4 a_n2140_13878.n2 0.146627
R22858 a_n2140_13878.n6 a_n2140_13878.n4 0.146627
R22859 a_n2140_13878.n10 a_n2140_13878.n9 0.101793
R22860 plus.n46 plus.t9 252.611
R22861 plus.n9 plus.t11 252.611
R22862 plus.n76 plus.t4 243.97
R22863 plus.n72 plus.t12 231.093
R22864 plus.n35 plus.t7 231.093
R22865 plus.n76 plus.n75 223.454
R22866 plus.n78 plus.n77 223.454
R22867 plus.n47 plus.t5 187.445
R22868 plus.n44 plus.t18 187.445
R22869 plus.n42 plus.t17 187.445
R22870 plus.n59 plus.t13 187.445
R22871 plus.n65 plus.t14 187.445
R22872 plus.n38 plus.t10 187.445
R22873 plus.n1 plus.t6 187.445
R22874 plus.n28 plus.t16 187.445
R22875 plus.n22 plus.t15 187.445
R22876 plus.n5 plus.t20 187.445
R22877 plus.n7 plus.t19 187.445
R22878 plus.n10 plus.t8 187.445
R22879 plus.n73 plus.n72 161.3
R22880 plus.n71 plus.n37 161.3
R22881 plus.n70 plus.n69 161.3
R22882 plus.n68 plus.n67 161.3
R22883 plus.n66 plus.n39 161.3
R22884 plus.n64 plus.n63 161.3
R22885 plus.n62 plus.n40 161.3
R22886 plus.n61 plus.n60 161.3
R22887 plus.n58 plus.n41 161.3
R22888 plus.n57 plus.n56 161.3
R22889 plus.n55 plus.n54 161.3
R22890 plus.n53 plus.n43 161.3
R22891 plus.n52 plus.n51 161.3
R22892 plus.n50 plus.n49 161.3
R22893 plus.n48 plus.n45 161.3
R22894 plus.n11 plus.n8 161.3
R22895 plus.n13 plus.n12 161.3
R22896 plus.n15 plus.n14 161.3
R22897 plus.n16 plus.n6 161.3
R22898 plus.n18 plus.n17 161.3
R22899 plus.n20 plus.n19 161.3
R22900 plus.n21 plus.n4 161.3
R22901 plus.n24 plus.n23 161.3
R22902 plus.n25 plus.n3 161.3
R22903 plus.n27 plus.n26 161.3
R22904 plus.n29 plus.n2 161.3
R22905 plus.n31 plus.n30 161.3
R22906 plus.n33 plus.n32 161.3
R22907 plus.n34 plus.n0 161.3
R22908 plus.n36 plus.n35 161.3
R22909 plus.n49 plus.n48 56.5617
R22910 plus.n58 plus.n57 56.5617
R22911 plus.n67 plus.n66 56.5617
R22912 plus.n30 plus.n29 56.5617
R22913 plus.n21 plus.n20 56.5617
R22914 plus.n12 plus.n11 56.5617
R22915 plus.n71 plus.n70 46.3896
R22916 plus.n34 plus.n33 46.3896
R22917 plus.n46 plus.n45 42.8164
R22918 plus.n9 plus.n8 42.8164
R22919 plus.n54 plus.n53 42.5146
R22920 plus.n60 plus.n40 42.5146
R22921 plus.n23 plus.n3 42.5146
R22922 plus.n17 plus.n16 42.5146
R22923 plus.n53 plus.n52 38.6395
R22924 plus.n64 plus.n40 38.6395
R22925 plus.n27 plus.n3 38.6395
R22926 plus.n16 plus.n15 38.6395
R22927 plus.n47 plus.n46 38.2514
R22928 plus.n10 plus.n9 38.2514
R22929 plus.n74 plus.n73 31.491
R22930 plus.n49 plus.n44 19.9199
R22931 plus.n66 plus.n65 19.9199
R22932 plus.n29 plus.n28 19.9199
R22933 plus.n12 plus.n7 19.9199
R22934 plus.n75 plus.t1 19.8005
R22935 plus.n75 plus.t2 19.8005
R22936 plus.n77 plus.t0 19.8005
R22937 plus.n77 plus.t3 19.8005
R22938 plus.n57 plus.n42 17.9525
R22939 plus.n59 plus.n58 17.9525
R22940 plus.n22 plus.n21 17.9525
R22941 plus.n20 plus.n5 17.9525
R22942 plus.n48 plus.n47 15.9852
R22943 plus.n67 plus.n38 15.9852
R22944 plus.n30 plus.n1 15.9852
R22945 plus.n11 plus.n10 15.9852
R22946 plus.n72 plus.n71 15.3369
R22947 plus.n35 plus.n34 15.3369
R22948 plus plus.n79 14.7178
R22949 plus.n74 plus.n36 11.9494
R22950 plus.n70 plus.n38 8.60764
R22951 plus.n33 plus.n1 8.60764
R22952 plus.n54 plus.n42 6.6403
R22953 plus.n60 plus.n59 6.6403
R22954 plus.n23 plus.n22 6.6403
R22955 plus.n17 plus.n5 6.6403
R22956 plus.n79 plus.n78 5.40567
R22957 plus.n52 plus.n44 4.67295
R22958 plus.n65 plus.n64 4.67295
R22959 plus.n28 plus.n27 4.67295
R22960 plus.n15 plus.n7 4.67295
R22961 plus.n79 plus.n74 1.188
R22962 plus.n78 plus.n76 0.716017
R22963 plus.n50 plus.n45 0.189894
R22964 plus.n51 plus.n50 0.189894
R22965 plus.n51 plus.n43 0.189894
R22966 plus.n55 plus.n43 0.189894
R22967 plus.n56 plus.n55 0.189894
R22968 plus.n56 plus.n41 0.189894
R22969 plus.n61 plus.n41 0.189894
R22970 plus.n62 plus.n61 0.189894
R22971 plus.n63 plus.n62 0.189894
R22972 plus.n63 plus.n39 0.189894
R22973 plus.n68 plus.n39 0.189894
R22974 plus.n69 plus.n68 0.189894
R22975 plus.n69 plus.n37 0.189894
R22976 plus.n73 plus.n37 0.189894
R22977 plus.n36 plus.n0 0.189894
R22978 plus.n32 plus.n0 0.189894
R22979 plus.n32 plus.n31 0.189894
R22980 plus.n31 plus.n2 0.189894
R22981 plus.n26 plus.n2 0.189894
R22982 plus.n26 plus.n25 0.189894
R22983 plus.n25 plus.n24 0.189894
R22984 plus.n24 plus.n4 0.189894
R22985 plus.n19 plus.n4 0.189894
R22986 plus.n19 plus.n18 0.189894
R22987 plus.n18 plus.n6 0.189894
R22988 plus.n14 plus.n6 0.189894
R22989 plus.n14 plus.n13 0.189894
R22990 plus.n13 plus.n8 0.189894
R22991 a_n3827_n3924.n2 a_n3827_n3924.t10 214.994
R22992 a_n3827_n3924.n12 a_n3827_n3924.t0 214.994
R22993 a_n3827_n3924.n2 a_n3827_n3924.t6 214.321
R22994 a_n3827_n3924.n13 a_n3827_n3924.t12 214.321
R22995 a_n3827_n3924.n14 a_n3827_n3924.t37 214.321
R22996 a_n3827_n3924.n15 a_n3827_n3924.t38 214.321
R22997 a_n3827_n3924.n16 a_n3827_n3924.t1 214.321
R22998 a_n3827_n3924.n17 a_n3827_n3924.t5 214.321
R22999 a_n3827_n3924.n0 a_n3827_n3924.t30 214.321
R23000 a_n3827_n3924.n12 a_n3827_n3924.t11 214.321
R23001 a_n3827_n3924.n1 a_n3827_n3924.t25 55.8337
R23002 a_n3827_n3924.n4 a_n3827_n3924.t36 55.8337
R23003 a_n3827_n3924.n11 a_n3827_n3924.t8 55.8337
R23004 a_n3827_n3924.n36 a_n3827_n3924.t22 55.8335
R23005 a_n3827_n3924.n34 a_n3827_n3924.t31 55.8335
R23006 a_n3827_n3924.n27 a_n3827_n3924.t3 55.8335
R23007 a_n3827_n3924.n26 a_n3827_n3924.t23 55.8335
R23008 a_n3827_n3924.n19 a_n3827_n3924.t27 55.8335
R23009 a_n3827_n3924.n38 a_n3827_n3924.n37 53.0052
R23010 a_n3827_n3924.n40 a_n3827_n3924.n39 53.0052
R23011 a_n3827_n3924.n6 a_n3827_n3924.n5 53.0052
R23012 a_n3827_n3924.n8 a_n3827_n3924.n7 53.0052
R23013 a_n3827_n3924.n10 a_n3827_n3924.n9 53.0052
R23014 a_n3827_n3924.n33 a_n3827_n3924.n32 53.0051
R23015 a_n3827_n3924.n31 a_n3827_n3924.n30 53.0051
R23016 a_n3827_n3924.n29 a_n3827_n3924.n28 53.0051
R23017 a_n3827_n3924.n25 a_n3827_n3924.n24 53.0051
R23018 a_n3827_n3924.n23 a_n3827_n3924.n22 53.0051
R23019 a_n3827_n3924.n21 a_n3827_n3924.n20 53.0051
R23020 a_n3827_n3924.n42 a_n3827_n3924.n41 53.0051
R23021 a_n3827_n3924.n18 a_n3827_n3924.n11 12.2417
R23022 a_n3827_n3924.n36 a_n3827_n3924.n35 12.2417
R23023 a_n3827_n3924.n19 a_n3827_n3924.n18 5.16214
R23024 a_n3827_n3924.n35 a_n3827_n3924.n34 5.16214
R23025 a_n3827_n3924.n37 a_n3827_n3924.t20 2.82907
R23026 a_n3827_n3924.n37 a_n3827_n3924.t24 2.82907
R23027 a_n3827_n3924.n39 a_n3827_n3924.t17 2.82907
R23028 a_n3827_n3924.n39 a_n3827_n3924.t21 2.82907
R23029 a_n3827_n3924.n5 a_n3827_n3924.t41 2.82907
R23030 a_n3827_n3924.n5 a_n3827_n3924.t33 2.82907
R23031 a_n3827_n3924.n7 a_n3827_n3924.t4 2.82907
R23032 a_n3827_n3924.n7 a_n3827_n3924.t35 2.82907
R23033 a_n3827_n3924.n9 a_n3827_n3924.t34 2.82907
R23034 a_n3827_n3924.n9 a_n3827_n3924.t13 2.82907
R23035 a_n3827_n3924.n32 a_n3827_n3924.t7 2.82907
R23036 a_n3827_n3924.n32 a_n3827_n3924.t2 2.82907
R23037 a_n3827_n3924.n30 a_n3827_n3924.t39 2.82907
R23038 a_n3827_n3924.n30 a_n3827_n3924.t32 2.82907
R23039 a_n3827_n3924.n28 a_n3827_n3924.t9 2.82907
R23040 a_n3827_n3924.n28 a_n3827_n3924.t40 2.82907
R23041 a_n3827_n3924.n24 a_n3827_n3924.t15 2.82907
R23042 a_n3827_n3924.n24 a_n3827_n3924.t26 2.82907
R23043 a_n3827_n3924.n22 a_n3827_n3924.t19 2.82907
R23044 a_n3827_n3924.n22 a_n3827_n3924.t14 2.82907
R23045 a_n3827_n3924.n20 a_n3827_n3924.t28 2.82907
R23046 a_n3827_n3924.n20 a_n3827_n3924.t18 2.82907
R23047 a_n3827_n3924.t29 a_n3827_n3924.n42 2.82907
R23048 a_n3827_n3924.n42 a_n3827_n3924.t16 2.82907
R23049 a_n3827_n3924.n35 a_n3827_n3924.n3 1.95694
R23050 a_n3827_n3924.n18 a_n3827_n3924.n0 1.95694
R23051 a_n3827_n3924.n0 a_n3827_n3924.n17 0.672012
R23052 a_n3827_n3924.n17 a_n3827_n3924.n16 0.672012
R23053 a_n3827_n3924.n16 a_n3827_n3924.n15 0.672012
R23054 a_n3827_n3924.n15 a_n3827_n3924.n14 0.672012
R23055 a_n3827_n3924.n14 a_n3827_n3924.n13 0.672012
R23056 a_n3827_n3924.n0 a_n3827_n3924.n12 0.672012
R23057 a_n3827_n3924.n13 a_n3827_n3924.n3 0.541924
R23058 a_n3827_n3924.n21 a_n3827_n3924.n19 0.530672
R23059 a_n3827_n3924.n23 a_n3827_n3924.n21 0.530672
R23060 a_n3827_n3924.n25 a_n3827_n3924.n23 0.530672
R23061 a_n3827_n3924.n26 a_n3827_n3924.n25 0.530672
R23062 a_n3827_n3924.n29 a_n3827_n3924.n27 0.530672
R23063 a_n3827_n3924.n31 a_n3827_n3924.n29 0.530672
R23064 a_n3827_n3924.n33 a_n3827_n3924.n31 0.530672
R23065 a_n3827_n3924.n34 a_n3827_n3924.n33 0.530672
R23066 a_n3827_n3924.n11 a_n3827_n3924.n10 0.530672
R23067 a_n3827_n3924.n10 a_n3827_n3924.n8 0.530672
R23068 a_n3827_n3924.n8 a_n3827_n3924.n6 0.530672
R23069 a_n3827_n3924.n6 a_n3827_n3924.n4 0.530672
R23070 a_n3827_n3924.n41 a_n3827_n3924.n1 0.530672
R23071 a_n3827_n3924.n41 a_n3827_n3924.n40 0.530672
R23072 a_n3827_n3924.n40 a_n3827_n3924.n38 0.530672
R23073 a_n3827_n3924.n38 a_n3827_n3924.n36 0.530672
R23074 a_n3827_n3924.n27 a_n3827_n3924.n26 0.235414
R23075 a_n3827_n3924.n4 a_n3827_n3924.n1 0.235414
R23076 a_n3827_n3924.n3 a_n3827_n3924.n2 0.130587
R23077 diffpairibias.n0 diffpairibias.t27 436.822
R23078 diffpairibias.n27 diffpairibias.t24 435.479
R23079 diffpairibias.n26 diffpairibias.t21 435.479
R23080 diffpairibias.n25 diffpairibias.t22 435.479
R23081 diffpairibias.n24 diffpairibias.t26 435.479
R23082 diffpairibias.n23 diffpairibias.t20 435.479
R23083 diffpairibias.n0 diffpairibias.t23 435.479
R23084 diffpairibias.n1 diffpairibias.t28 435.479
R23085 diffpairibias.n2 diffpairibias.t25 435.479
R23086 diffpairibias.n3 diffpairibias.t29 435.479
R23087 diffpairibias.n13 diffpairibias.t14 377.536
R23088 diffpairibias.n13 diffpairibias.t0 376.193
R23089 diffpairibias.n14 diffpairibias.t10 376.193
R23090 diffpairibias.n15 diffpairibias.t12 376.193
R23091 diffpairibias.n16 diffpairibias.t6 376.193
R23092 diffpairibias.n17 diffpairibias.t2 376.193
R23093 diffpairibias.n18 diffpairibias.t16 376.193
R23094 diffpairibias.n19 diffpairibias.t4 376.193
R23095 diffpairibias.n20 diffpairibias.t18 376.193
R23096 diffpairibias.n21 diffpairibias.t8 376.193
R23097 diffpairibias.n4 diffpairibias.t15 113.368
R23098 diffpairibias.n4 diffpairibias.t1 112.698
R23099 diffpairibias.n5 diffpairibias.t11 112.698
R23100 diffpairibias.n6 diffpairibias.t13 112.698
R23101 diffpairibias.n7 diffpairibias.t7 112.698
R23102 diffpairibias.n8 diffpairibias.t3 112.698
R23103 diffpairibias.n9 diffpairibias.t17 112.698
R23104 diffpairibias.n10 diffpairibias.t5 112.698
R23105 diffpairibias.n11 diffpairibias.t19 112.698
R23106 diffpairibias.n12 diffpairibias.t9 112.698
R23107 diffpairibias.n22 diffpairibias.n21 4.77242
R23108 diffpairibias.n22 diffpairibias.n12 4.30807
R23109 diffpairibias.n23 diffpairibias.n22 4.13945
R23110 diffpairibias.n21 diffpairibias.n20 1.34352
R23111 diffpairibias.n20 diffpairibias.n19 1.34352
R23112 diffpairibias.n19 diffpairibias.n18 1.34352
R23113 diffpairibias.n18 diffpairibias.n17 1.34352
R23114 diffpairibias.n17 diffpairibias.n16 1.34352
R23115 diffpairibias.n16 diffpairibias.n15 1.34352
R23116 diffpairibias.n15 diffpairibias.n14 1.34352
R23117 diffpairibias.n14 diffpairibias.n13 1.34352
R23118 diffpairibias.n3 diffpairibias.n2 1.34352
R23119 diffpairibias.n2 diffpairibias.n1 1.34352
R23120 diffpairibias.n1 diffpairibias.n0 1.34352
R23121 diffpairibias.n24 diffpairibias.n23 1.34352
R23122 diffpairibias.n25 diffpairibias.n24 1.34352
R23123 diffpairibias.n26 diffpairibias.n25 1.34352
R23124 diffpairibias.n27 diffpairibias.n26 1.34352
R23125 diffpairibias.n28 diffpairibias.n27 0.862419
R23126 diffpairibias diffpairibias.n28 0.684875
R23127 diffpairibias.n12 diffpairibias.n11 0.672012
R23128 diffpairibias.n11 diffpairibias.n10 0.672012
R23129 diffpairibias.n10 diffpairibias.n9 0.672012
R23130 diffpairibias.n9 diffpairibias.n8 0.672012
R23131 diffpairibias.n8 diffpairibias.n7 0.672012
R23132 diffpairibias.n7 diffpairibias.n6 0.672012
R23133 diffpairibias.n6 diffpairibias.n5 0.672012
R23134 diffpairibias.n5 diffpairibias.n4 0.672012
R23135 diffpairibias.n28 diffpairibias.n3 0.190907
R23136 minus.n46 minus.t20 252.611
R23137 minus.n9 minus.t13 252.611
R23138 minus.n78 minus.t3 243.255
R23139 minus.n72 minus.t15 231.093
R23140 minus.n35 minus.t17 231.093
R23141 minus.n77 minus.n75 224.169
R23142 minus.n77 minus.n76 223.454
R23143 minus.n38 minus.t12 187.445
R23144 minus.n65 minus.t7 187.445
R23145 minus.n59 minus.t6 187.445
R23146 minus.n42 minus.t11 187.445
R23147 minus.n44 minus.t10 187.445
R23148 minus.n47 minus.t16 187.445
R23149 minus.n10 minus.t9 187.445
R23150 minus.n7 minus.t8 187.445
R23151 minus.n5 minus.t5 187.445
R23152 minus.n22 minus.t18 187.445
R23153 minus.n28 minus.t19 187.445
R23154 minus.n1 minus.t14 187.445
R23155 minus.n48 minus.n45 161.3
R23156 minus.n50 minus.n49 161.3
R23157 minus.n52 minus.n51 161.3
R23158 minus.n53 minus.n43 161.3
R23159 minus.n55 minus.n54 161.3
R23160 minus.n57 minus.n56 161.3
R23161 minus.n58 minus.n41 161.3
R23162 minus.n61 minus.n60 161.3
R23163 minus.n62 minus.n40 161.3
R23164 minus.n64 minus.n63 161.3
R23165 minus.n66 minus.n39 161.3
R23166 minus.n68 minus.n67 161.3
R23167 minus.n70 minus.n69 161.3
R23168 minus.n71 minus.n37 161.3
R23169 minus.n73 minus.n72 161.3
R23170 minus.n36 minus.n35 161.3
R23171 minus.n34 minus.n0 161.3
R23172 minus.n33 minus.n32 161.3
R23173 minus.n31 minus.n30 161.3
R23174 minus.n29 minus.n2 161.3
R23175 minus.n27 minus.n26 161.3
R23176 minus.n25 minus.n3 161.3
R23177 minus.n24 minus.n23 161.3
R23178 minus.n21 minus.n4 161.3
R23179 minus.n20 minus.n19 161.3
R23180 minus.n18 minus.n17 161.3
R23181 minus.n16 minus.n6 161.3
R23182 minus.n15 minus.n14 161.3
R23183 minus.n13 minus.n12 161.3
R23184 minus.n11 minus.n8 161.3
R23185 minus.n67 minus.n66 56.5617
R23186 minus.n58 minus.n57 56.5617
R23187 minus.n49 minus.n48 56.5617
R23188 minus.n12 minus.n11 56.5617
R23189 minus.n21 minus.n20 56.5617
R23190 minus.n30 minus.n29 56.5617
R23191 minus.n71 minus.n70 46.3896
R23192 minus.n34 minus.n33 46.3896
R23193 minus.n46 minus.n45 42.8164
R23194 minus.n9 minus.n8 42.8164
R23195 minus.n60 minus.n40 42.5146
R23196 minus.n54 minus.n53 42.5146
R23197 minus.n17 minus.n16 42.5146
R23198 minus.n23 minus.n3 42.5146
R23199 minus.n64 minus.n40 38.6395
R23200 minus.n53 minus.n52 38.6395
R23201 minus.n16 minus.n15 38.6395
R23202 minus.n27 minus.n3 38.6395
R23203 minus.n47 minus.n46 38.2514
R23204 minus.n10 minus.n9 38.2514
R23205 minus.n74 minus.n73 31.7069
R23206 minus.n66 minus.n65 19.9199
R23207 minus.n49 minus.n44 19.9199
R23208 minus.n12 minus.n7 19.9199
R23209 minus.n29 minus.n28 19.9199
R23210 minus.n76 minus.t2 19.8005
R23211 minus.n76 minus.t0 19.8005
R23212 minus.n75 minus.t1 19.8005
R23213 minus.n75 minus.t4 19.8005
R23214 minus.n59 minus.n58 17.9525
R23215 minus.n57 minus.n42 17.9525
R23216 minus.n20 minus.n5 17.9525
R23217 minus.n22 minus.n21 17.9525
R23218 minus.n67 minus.n38 15.9852
R23219 minus.n48 minus.n47 15.9852
R23220 minus.n11 minus.n10 15.9852
R23221 minus.n30 minus.n1 15.9852
R23222 minus.n72 minus.n71 15.3369
R23223 minus.n35 minus.n34 15.3369
R23224 minus.n74 minus.n36 12.1653
R23225 minus minus.n79 11.8456
R23226 minus.n70 minus.n38 8.60764
R23227 minus.n33 minus.n1 8.60764
R23228 minus.n60 minus.n59 6.6403
R23229 minus.n54 minus.n42 6.6403
R23230 minus.n17 minus.n5 6.6403
R23231 minus.n23 minus.n22 6.6403
R23232 minus.n79 minus.n78 4.80222
R23233 minus.n65 minus.n64 4.67295
R23234 minus.n52 minus.n44 4.67295
R23235 minus.n15 minus.n7 4.67295
R23236 minus.n28 minus.n27 4.67295
R23237 minus.n79 minus.n74 0.972091
R23238 minus.n78 minus.n77 0.716017
R23239 minus.n73 minus.n37 0.189894
R23240 minus.n69 minus.n37 0.189894
R23241 minus.n69 minus.n68 0.189894
R23242 minus.n68 minus.n39 0.189894
R23243 minus.n63 minus.n39 0.189894
R23244 minus.n63 minus.n62 0.189894
R23245 minus.n62 minus.n61 0.189894
R23246 minus.n61 minus.n41 0.189894
R23247 minus.n56 minus.n41 0.189894
R23248 minus.n56 minus.n55 0.189894
R23249 minus.n55 minus.n43 0.189894
R23250 minus.n51 minus.n43 0.189894
R23251 minus.n51 minus.n50 0.189894
R23252 minus.n50 minus.n45 0.189894
R23253 minus.n13 minus.n8 0.189894
R23254 minus.n14 minus.n13 0.189894
R23255 minus.n14 minus.n6 0.189894
R23256 minus.n18 minus.n6 0.189894
R23257 minus.n19 minus.n18 0.189894
R23258 minus.n19 minus.n4 0.189894
R23259 minus.n24 minus.n4 0.189894
R23260 minus.n25 minus.n24 0.189894
R23261 minus.n26 minus.n25 0.189894
R23262 minus.n26 minus.n2 0.189894
R23263 minus.n31 minus.n2 0.189894
R23264 minus.n32 minus.n31 0.189894
R23265 minus.n32 minus.n0 0.189894
R23266 minus.n36 minus.n0 0.189894
R23267 a_n2318_8322.n8 a_n2318_8322.t3 74.6477
R23268 a_n2318_8322.n1 a_n2318_8322.t22 74.6477
R23269 a_n2318_8322.n20 a_n2318_8322.t21 74.6474
R23270 a_n2318_8322.n16 a_n2318_8322.t11 74.2899
R23271 a_n2318_8322.n9 a_n2318_8322.t1 74.2899
R23272 a_n2318_8322.n10 a_n2318_8322.t4 74.2899
R23273 a_n2318_8322.n13 a_n2318_8322.t5 74.2899
R23274 a_n2318_8322.n6 a_n2318_8322.t8 74.2899
R23275 a_n2318_8322.n20 a_n2318_8322.n19 70.6783
R23276 a_n2318_8322.n18 a_n2318_8322.n17 70.6783
R23277 a_n2318_8322.n8 a_n2318_8322.n7 70.6783
R23278 a_n2318_8322.n12 a_n2318_8322.n11 70.6783
R23279 a_n2318_8322.n1 a_n2318_8322.n0 70.6783
R23280 a_n2318_8322.n3 a_n2318_8322.n2 70.6783
R23281 a_n2318_8322.n5 a_n2318_8322.n4 70.6783
R23282 a_n2318_8322.n22 a_n2318_8322.n21 70.6782
R23283 a_n2318_8322.n14 a_n2318_8322.n6 23.4712
R23284 a_n2318_8322.n15 a_n2318_8322.t24 10.0049
R23285 a_n2318_8322.n14 a_n2318_8322.n13 6.95632
R23286 a_n2318_8322.n16 a_n2318_8322.n15 6.19447
R23287 a_n2318_8322.n15 a_n2318_8322.n14 5.3452
R23288 a_n2318_8322.n19 a_n2318_8322.t18 3.61217
R23289 a_n2318_8322.n19 a_n2318_8322.t15 3.61217
R23290 a_n2318_8322.n17 a_n2318_8322.t20 3.61217
R23291 a_n2318_8322.n17 a_n2318_8322.t13 3.61217
R23292 a_n2318_8322.n7 a_n2318_8322.t7 3.61217
R23293 a_n2318_8322.n7 a_n2318_8322.t6 3.61217
R23294 a_n2318_8322.n11 a_n2318_8322.t2 3.61217
R23295 a_n2318_8322.n11 a_n2318_8322.t0 3.61217
R23296 a_n2318_8322.n0 a_n2318_8322.t10 3.61217
R23297 a_n2318_8322.n0 a_n2318_8322.t9 3.61217
R23298 a_n2318_8322.n2 a_n2318_8322.t19 3.61217
R23299 a_n2318_8322.n2 a_n2318_8322.t14 3.61217
R23300 a_n2318_8322.n4 a_n2318_8322.t17 3.61217
R23301 a_n2318_8322.n4 a_n2318_8322.t16 3.61217
R23302 a_n2318_8322.n22 a_n2318_8322.t12 3.61217
R23303 a_n2318_8322.t23 a_n2318_8322.n22 3.61217
R23304 a_n2318_8322.n13 a_n2318_8322.n12 0.358259
R23305 a_n2318_8322.n12 a_n2318_8322.n10 0.358259
R23306 a_n2318_8322.n9 a_n2318_8322.n8 0.358259
R23307 a_n2318_8322.n6 a_n2318_8322.n5 0.358259
R23308 a_n2318_8322.n5 a_n2318_8322.n3 0.358259
R23309 a_n2318_8322.n3 a_n2318_8322.n1 0.358259
R23310 a_n2318_8322.n18 a_n2318_8322.n16 0.358259
R23311 a_n2318_8322.n21 a_n2318_8322.n18 0.358259
R23312 a_n2318_8322.n21 a_n2318_8322.n20 0.358259
R23313 a_n2318_8322.n10 a_n2318_8322.n9 0.101793
R23314 a_n2318_8322.t26 a_n2318_8322.t27 0.0788333
R23315 a_n2318_8322.t25 a_n2318_8322.t26 0.0631667
R23316 a_n2318_8322.t24 a_n2318_8322.t25 0.0471944
R23317 a_n2318_8322.t24 a_n2318_8322.t27 0.0453889
R23318 outputibias.n27 outputibias.n1 289.615
R23319 outputibias.n58 outputibias.n32 289.615
R23320 outputibias.n90 outputibias.n64 289.615
R23321 outputibias.n122 outputibias.n96 289.615
R23322 outputibias.n28 outputibias.n27 185
R23323 outputibias.n26 outputibias.n25 185
R23324 outputibias.n5 outputibias.n4 185
R23325 outputibias.n20 outputibias.n19 185
R23326 outputibias.n18 outputibias.n17 185
R23327 outputibias.n9 outputibias.n8 185
R23328 outputibias.n12 outputibias.n11 185
R23329 outputibias.n59 outputibias.n58 185
R23330 outputibias.n57 outputibias.n56 185
R23331 outputibias.n36 outputibias.n35 185
R23332 outputibias.n51 outputibias.n50 185
R23333 outputibias.n49 outputibias.n48 185
R23334 outputibias.n40 outputibias.n39 185
R23335 outputibias.n43 outputibias.n42 185
R23336 outputibias.n91 outputibias.n90 185
R23337 outputibias.n89 outputibias.n88 185
R23338 outputibias.n68 outputibias.n67 185
R23339 outputibias.n83 outputibias.n82 185
R23340 outputibias.n81 outputibias.n80 185
R23341 outputibias.n72 outputibias.n71 185
R23342 outputibias.n75 outputibias.n74 185
R23343 outputibias.n123 outputibias.n122 185
R23344 outputibias.n121 outputibias.n120 185
R23345 outputibias.n100 outputibias.n99 185
R23346 outputibias.n115 outputibias.n114 185
R23347 outputibias.n113 outputibias.n112 185
R23348 outputibias.n104 outputibias.n103 185
R23349 outputibias.n107 outputibias.n106 185
R23350 outputibias.n0 outputibias.t9 178.945
R23351 outputibias.n133 outputibias.t8 177.018
R23352 outputibias.n132 outputibias.t11 177.018
R23353 outputibias.n0 outputibias.t10 177.018
R23354 outputibias.t5 outputibias.n10 147.661
R23355 outputibias.t7 outputibias.n41 147.661
R23356 outputibias.t1 outputibias.n73 147.661
R23357 outputibias.t3 outputibias.n105 147.661
R23358 outputibias.n128 outputibias.t4 132.363
R23359 outputibias.n128 outputibias.t6 130.436
R23360 outputibias.n129 outputibias.t0 130.436
R23361 outputibias.n130 outputibias.t2 130.436
R23362 outputibias.n27 outputibias.n26 104.615
R23363 outputibias.n26 outputibias.n4 104.615
R23364 outputibias.n19 outputibias.n4 104.615
R23365 outputibias.n19 outputibias.n18 104.615
R23366 outputibias.n18 outputibias.n8 104.615
R23367 outputibias.n11 outputibias.n8 104.615
R23368 outputibias.n58 outputibias.n57 104.615
R23369 outputibias.n57 outputibias.n35 104.615
R23370 outputibias.n50 outputibias.n35 104.615
R23371 outputibias.n50 outputibias.n49 104.615
R23372 outputibias.n49 outputibias.n39 104.615
R23373 outputibias.n42 outputibias.n39 104.615
R23374 outputibias.n90 outputibias.n89 104.615
R23375 outputibias.n89 outputibias.n67 104.615
R23376 outputibias.n82 outputibias.n67 104.615
R23377 outputibias.n82 outputibias.n81 104.615
R23378 outputibias.n81 outputibias.n71 104.615
R23379 outputibias.n74 outputibias.n71 104.615
R23380 outputibias.n122 outputibias.n121 104.615
R23381 outputibias.n121 outputibias.n99 104.615
R23382 outputibias.n114 outputibias.n99 104.615
R23383 outputibias.n114 outputibias.n113 104.615
R23384 outputibias.n113 outputibias.n103 104.615
R23385 outputibias.n106 outputibias.n103 104.615
R23386 outputibias.n63 outputibias.n31 95.6354
R23387 outputibias.n63 outputibias.n62 94.6732
R23388 outputibias.n95 outputibias.n94 94.6732
R23389 outputibias.n127 outputibias.n126 94.6732
R23390 outputibias.n11 outputibias.t5 52.3082
R23391 outputibias.n42 outputibias.t7 52.3082
R23392 outputibias.n74 outputibias.t1 52.3082
R23393 outputibias.n106 outputibias.t3 52.3082
R23394 outputibias.n12 outputibias.n10 15.6674
R23395 outputibias.n43 outputibias.n41 15.6674
R23396 outputibias.n75 outputibias.n73 15.6674
R23397 outputibias.n107 outputibias.n105 15.6674
R23398 outputibias.n13 outputibias.n9 12.8005
R23399 outputibias.n44 outputibias.n40 12.8005
R23400 outputibias.n76 outputibias.n72 12.8005
R23401 outputibias.n108 outputibias.n104 12.8005
R23402 outputibias.n17 outputibias.n16 12.0247
R23403 outputibias.n48 outputibias.n47 12.0247
R23404 outputibias.n80 outputibias.n79 12.0247
R23405 outputibias.n112 outputibias.n111 12.0247
R23406 outputibias.n20 outputibias.n7 11.249
R23407 outputibias.n51 outputibias.n38 11.249
R23408 outputibias.n83 outputibias.n70 11.249
R23409 outputibias.n115 outputibias.n102 11.249
R23410 outputibias.n21 outputibias.n5 10.4732
R23411 outputibias.n52 outputibias.n36 10.4732
R23412 outputibias.n84 outputibias.n68 10.4732
R23413 outputibias.n116 outputibias.n100 10.4732
R23414 outputibias.n25 outputibias.n24 9.69747
R23415 outputibias.n56 outputibias.n55 9.69747
R23416 outputibias.n88 outputibias.n87 9.69747
R23417 outputibias.n120 outputibias.n119 9.69747
R23418 outputibias.n31 outputibias.n30 9.45567
R23419 outputibias.n62 outputibias.n61 9.45567
R23420 outputibias.n94 outputibias.n93 9.45567
R23421 outputibias.n126 outputibias.n125 9.45567
R23422 outputibias.n30 outputibias.n29 9.3005
R23423 outputibias.n3 outputibias.n2 9.3005
R23424 outputibias.n24 outputibias.n23 9.3005
R23425 outputibias.n22 outputibias.n21 9.3005
R23426 outputibias.n7 outputibias.n6 9.3005
R23427 outputibias.n16 outputibias.n15 9.3005
R23428 outputibias.n14 outputibias.n13 9.3005
R23429 outputibias.n61 outputibias.n60 9.3005
R23430 outputibias.n34 outputibias.n33 9.3005
R23431 outputibias.n55 outputibias.n54 9.3005
R23432 outputibias.n53 outputibias.n52 9.3005
R23433 outputibias.n38 outputibias.n37 9.3005
R23434 outputibias.n47 outputibias.n46 9.3005
R23435 outputibias.n45 outputibias.n44 9.3005
R23436 outputibias.n93 outputibias.n92 9.3005
R23437 outputibias.n66 outputibias.n65 9.3005
R23438 outputibias.n87 outputibias.n86 9.3005
R23439 outputibias.n85 outputibias.n84 9.3005
R23440 outputibias.n70 outputibias.n69 9.3005
R23441 outputibias.n79 outputibias.n78 9.3005
R23442 outputibias.n77 outputibias.n76 9.3005
R23443 outputibias.n125 outputibias.n124 9.3005
R23444 outputibias.n98 outputibias.n97 9.3005
R23445 outputibias.n119 outputibias.n118 9.3005
R23446 outputibias.n117 outputibias.n116 9.3005
R23447 outputibias.n102 outputibias.n101 9.3005
R23448 outputibias.n111 outputibias.n110 9.3005
R23449 outputibias.n109 outputibias.n108 9.3005
R23450 outputibias.n28 outputibias.n3 8.92171
R23451 outputibias.n59 outputibias.n34 8.92171
R23452 outputibias.n91 outputibias.n66 8.92171
R23453 outputibias.n123 outputibias.n98 8.92171
R23454 outputibias.n29 outputibias.n1 8.14595
R23455 outputibias.n60 outputibias.n32 8.14595
R23456 outputibias.n92 outputibias.n64 8.14595
R23457 outputibias.n124 outputibias.n96 8.14595
R23458 outputibias.n31 outputibias.n1 5.81868
R23459 outputibias.n62 outputibias.n32 5.81868
R23460 outputibias.n94 outputibias.n64 5.81868
R23461 outputibias.n126 outputibias.n96 5.81868
R23462 outputibias.n131 outputibias.n130 5.20947
R23463 outputibias.n29 outputibias.n28 5.04292
R23464 outputibias.n60 outputibias.n59 5.04292
R23465 outputibias.n92 outputibias.n91 5.04292
R23466 outputibias.n124 outputibias.n123 5.04292
R23467 outputibias.n131 outputibias.n127 4.42209
R23468 outputibias.n14 outputibias.n10 4.38594
R23469 outputibias.n45 outputibias.n41 4.38594
R23470 outputibias.n77 outputibias.n73 4.38594
R23471 outputibias.n109 outputibias.n105 4.38594
R23472 outputibias.n132 outputibias.n131 4.28454
R23473 outputibias.n25 outputibias.n3 4.26717
R23474 outputibias.n56 outputibias.n34 4.26717
R23475 outputibias.n88 outputibias.n66 4.26717
R23476 outputibias.n120 outputibias.n98 4.26717
R23477 outputibias.n24 outputibias.n5 3.49141
R23478 outputibias.n55 outputibias.n36 3.49141
R23479 outputibias.n87 outputibias.n68 3.49141
R23480 outputibias.n119 outputibias.n100 3.49141
R23481 outputibias.n21 outputibias.n20 2.71565
R23482 outputibias.n52 outputibias.n51 2.71565
R23483 outputibias.n84 outputibias.n83 2.71565
R23484 outputibias.n116 outputibias.n115 2.71565
R23485 outputibias.n17 outputibias.n7 1.93989
R23486 outputibias.n48 outputibias.n38 1.93989
R23487 outputibias.n80 outputibias.n70 1.93989
R23488 outputibias.n112 outputibias.n102 1.93989
R23489 outputibias.n130 outputibias.n129 1.9266
R23490 outputibias.n129 outputibias.n128 1.9266
R23491 outputibias.n133 outputibias.n132 1.92658
R23492 outputibias.n134 outputibias.n133 1.29913
R23493 outputibias.n16 outputibias.n9 1.16414
R23494 outputibias.n47 outputibias.n40 1.16414
R23495 outputibias.n79 outputibias.n72 1.16414
R23496 outputibias.n111 outputibias.n104 1.16414
R23497 outputibias.n127 outputibias.n95 0.962709
R23498 outputibias.n95 outputibias.n63 0.962709
R23499 outputibias.n13 outputibias.n12 0.388379
R23500 outputibias.n44 outputibias.n43 0.388379
R23501 outputibias.n76 outputibias.n75 0.388379
R23502 outputibias.n108 outputibias.n107 0.388379
R23503 outputibias.n134 outputibias.n0 0.337251
R23504 outputibias outputibias.n134 0.302375
R23505 outputibias.n30 outputibias.n2 0.155672
R23506 outputibias.n23 outputibias.n2 0.155672
R23507 outputibias.n23 outputibias.n22 0.155672
R23508 outputibias.n22 outputibias.n6 0.155672
R23509 outputibias.n15 outputibias.n6 0.155672
R23510 outputibias.n15 outputibias.n14 0.155672
R23511 outputibias.n61 outputibias.n33 0.155672
R23512 outputibias.n54 outputibias.n33 0.155672
R23513 outputibias.n54 outputibias.n53 0.155672
R23514 outputibias.n53 outputibias.n37 0.155672
R23515 outputibias.n46 outputibias.n37 0.155672
R23516 outputibias.n46 outputibias.n45 0.155672
R23517 outputibias.n93 outputibias.n65 0.155672
R23518 outputibias.n86 outputibias.n65 0.155672
R23519 outputibias.n86 outputibias.n85 0.155672
R23520 outputibias.n85 outputibias.n69 0.155672
R23521 outputibias.n78 outputibias.n69 0.155672
R23522 outputibias.n78 outputibias.n77 0.155672
R23523 outputibias.n125 outputibias.n97 0.155672
R23524 outputibias.n118 outputibias.n97 0.155672
R23525 outputibias.n118 outputibias.n117 0.155672
R23526 outputibias.n117 outputibias.n101 0.155672
R23527 outputibias.n110 outputibias.n101 0.155672
R23528 outputibias.n110 outputibias.n109 0.155672
R23529 output.n41 output.n15 289.615
R23530 output.n72 output.n46 289.615
R23531 output.n104 output.n78 289.615
R23532 output.n136 output.n110 289.615
R23533 output.n77 output.n45 197.26
R23534 output.n77 output.n76 196.298
R23535 output.n109 output.n108 196.298
R23536 output.n141 output.n140 196.298
R23537 output.n42 output.n41 185
R23538 output.n40 output.n39 185
R23539 output.n19 output.n18 185
R23540 output.n34 output.n33 185
R23541 output.n32 output.n31 185
R23542 output.n23 output.n22 185
R23543 output.n26 output.n25 185
R23544 output.n73 output.n72 185
R23545 output.n71 output.n70 185
R23546 output.n50 output.n49 185
R23547 output.n65 output.n64 185
R23548 output.n63 output.n62 185
R23549 output.n54 output.n53 185
R23550 output.n57 output.n56 185
R23551 output.n105 output.n104 185
R23552 output.n103 output.n102 185
R23553 output.n82 output.n81 185
R23554 output.n97 output.n96 185
R23555 output.n95 output.n94 185
R23556 output.n86 output.n85 185
R23557 output.n89 output.n88 185
R23558 output.n137 output.n136 185
R23559 output.n135 output.n134 185
R23560 output.n114 output.n113 185
R23561 output.n129 output.n128 185
R23562 output.n127 output.n126 185
R23563 output.n118 output.n117 185
R23564 output.n121 output.n120 185
R23565 output.t2 output.n24 147.661
R23566 output.t1 output.n55 147.661
R23567 output.t3 output.n87 147.661
R23568 output.t0 output.n119 147.661
R23569 output.n41 output.n40 104.615
R23570 output.n40 output.n18 104.615
R23571 output.n33 output.n18 104.615
R23572 output.n33 output.n32 104.615
R23573 output.n32 output.n22 104.615
R23574 output.n25 output.n22 104.615
R23575 output.n72 output.n71 104.615
R23576 output.n71 output.n49 104.615
R23577 output.n64 output.n49 104.615
R23578 output.n64 output.n63 104.615
R23579 output.n63 output.n53 104.615
R23580 output.n56 output.n53 104.615
R23581 output.n104 output.n103 104.615
R23582 output.n103 output.n81 104.615
R23583 output.n96 output.n81 104.615
R23584 output.n96 output.n95 104.615
R23585 output.n95 output.n85 104.615
R23586 output.n88 output.n85 104.615
R23587 output.n136 output.n135 104.615
R23588 output.n135 output.n113 104.615
R23589 output.n128 output.n113 104.615
R23590 output.n128 output.n127 104.615
R23591 output.n127 output.n117 104.615
R23592 output.n120 output.n117 104.615
R23593 output.n1 output.t8 77.056
R23594 output.n14 output.t9 76.6694
R23595 output.n1 output.n0 72.7095
R23596 output.n3 output.n2 72.7095
R23597 output.n5 output.n4 72.7095
R23598 output.n7 output.n6 72.7095
R23599 output.n9 output.n8 72.7095
R23600 output.n11 output.n10 72.7095
R23601 output.n13 output.n12 72.7095
R23602 output.n25 output.t2 52.3082
R23603 output.n56 output.t1 52.3082
R23604 output.n88 output.t3 52.3082
R23605 output.n120 output.t0 52.3082
R23606 output.n26 output.n24 15.6674
R23607 output.n57 output.n55 15.6674
R23608 output.n89 output.n87 15.6674
R23609 output.n121 output.n119 15.6674
R23610 output.n27 output.n23 12.8005
R23611 output.n58 output.n54 12.8005
R23612 output.n90 output.n86 12.8005
R23613 output.n122 output.n118 12.8005
R23614 output.n31 output.n30 12.0247
R23615 output.n62 output.n61 12.0247
R23616 output.n94 output.n93 12.0247
R23617 output.n126 output.n125 12.0247
R23618 output.n34 output.n21 11.249
R23619 output.n65 output.n52 11.249
R23620 output.n97 output.n84 11.249
R23621 output.n129 output.n116 11.249
R23622 output.n35 output.n19 10.4732
R23623 output.n66 output.n50 10.4732
R23624 output.n98 output.n82 10.4732
R23625 output.n130 output.n114 10.4732
R23626 output.n39 output.n38 9.69747
R23627 output.n70 output.n69 9.69747
R23628 output.n102 output.n101 9.69747
R23629 output.n134 output.n133 9.69747
R23630 output.n45 output.n44 9.45567
R23631 output.n76 output.n75 9.45567
R23632 output.n108 output.n107 9.45567
R23633 output.n140 output.n139 9.45567
R23634 output.n44 output.n43 9.3005
R23635 output.n17 output.n16 9.3005
R23636 output.n38 output.n37 9.3005
R23637 output.n36 output.n35 9.3005
R23638 output.n21 output.n20 9.3005
R23639 output.n30 output.n29 9.3005
R23640 output.n28 output.n27 9.3005
R23641 output.n75 output.n74 9.3005
R23642 output.n48 output.n47 9.3005
R23643 output.n69 output.n68 9.3005
R23644 output.n67 output.n66 9.3005
R23645 output.n52 output.n51 9.3005
R23646 output.n61 output.n60 9.3005
R23647 output.n59 output.n58 9.3005
R23648 output.n107 output.n106 9.3005
R23649 output.n80 output.n79 9.3005
R23650 output.n101 output.n100 9.3005
R23651 output.n99 output.n98 9.3005
R23652 output.n84 output.n83 9.3005
R23653 output.n93 output.n92 9.3005
R23654 output.n91 output.n90 9.3005
R23655 output.n139 output.n138 9.3005
R23656 output.n112 output.n111 9.3005
R23657 output.n133 output.n132 9.3005
R23658 output.n131 output.n130 9.3005
R23659 output.n116 output.n115 9.3005
R23660 output.n125 output.n124 9.3005
R23661 output.n123 output.n122 9.3005
R23662 output.n42 output.n17 8.92171
R23663 output.n73 output.n48 8.92171
R23664 output.n105 output.n80 8.92171
R23665 output.n137 output.n112 8.92171
R23666 output output.n141 8.15037
R23667 output.n43 output.n15 8.14595
R23668 output.n74 output.n46 8.14595
R23669 output.n106 output.n78 8.14595
R23670 output.n138 output.n110 8.14595
R23671 output.n45 output.n15 5.81868
R23672 output.n76 output.n46 5.81868
R23673 output.n108 output.n78 5.81868
R23674 output.n140 output.n110 5.81868
R23675 output.n43 output.n42 5.04292
R23676 output.n74 output.n73 5.04292
R23677 output.n106 output.n105 5.04292
R23678 output.n138 output.n137 5.04292
R23679 output.n28 output.n24 4.38594
R23680 output.n59 output.n55 4.38594
R23681 output.n91 output.n87 4.38594
R23682 output.n123 output.n119 4.38594
R23683 output.n39 output.n17 4.26717
R23684 output.n70 output.n48 4.26717
R23685 output.n102 output.n80 4.26717
R23686 output.n134 output.n112 4.26717
R23687 output.n0 output.t14 3.9605
R23688 output.n0 output.t18 3.9605
R23689 output.n2 output.t5 3.9605
R23690 output.n2 output.t10 3.9605
R23691 output.n4 output.t11 3.9605
R23692 output.n4 output.t16 3.9605
R23693 output.n6 output.t4 3.9605
R23694 output.n6 output.t12 3.9605
R23695 output.n8 output.t15 3.9605
R23696 output.n8 output.t13 3.9605
R23697 output.n10 output.t19 3.9605
R23698 output.n10 output.t6 3.9605
R23699 output.n12 output.t7 3.9605
R23700 output.n12 output.t17 3.9605
R23701 output.n38 output.n19 3.49141
R23702 output.n69 output.n50 3.49141
R23703 output.n101 output.n82 3.49141
R23704 output.n133 output.n114 3.49141
R23705 output.n35 output.n34 2.71565
R23706 output.n66 output.n65 2.71565
R23707 output.n98 output.n97 2.71565
R23708 output.n130 output.n129 2.71565
R23709 output.n31 output.n21 1.93989
R23710 output.n62 output.n52 1.93989
R23711 output.n94 output.n84 1.93989
R23712 output.n126 output.n116 1.93989
R23713 output.n30 output.n23 1.16414
R23714 output.n61 output.n54 1.16414
R23715 output.n93 output.n86 1.16414
R23716 output.n125 output.n118 1.16414
R23717 output.n141 output.n109 0.962709
R23718 output.n109 output.n77 0.962709
R23719 output.n27 output.n26 0.388379
R23720 output.n58 output.n57 0.388379
R23721 output.n90 output.n89 0.388379
R23722 output.n122 output.n121 0.388379
R23723 output.n14 output.n13 0.387128
R23724 output.n13 output.n11 0.387128
R23725 output.n11 output.n9 0.387128
R23726 output.n9 output.n7 0.387128
R23727 output.n7 output.n5 0.387128
R23728 output.n5 output.n3 0.387128
R23729 output.n3 output.n1 0.387128
R23730 output.n44 output.n16 0.155672
R23731 output.n37 output.n16 0.155672
R23732 output.n37 output.n36 0.155672
R23733 output.n36 output.n20 0.155672
R23734 output.n29 output.n20 0.155672
R23735 output.n29 output.n28 0.155672
R23736 output.n75 output.n47 0.155672
R23737 output.n68 output.n47 0.155672
R23738 output.n68 output.n67 0.155672
R23739 output.n67 output.n51 0.155672
R23740 output.n60 output.n51 0.155672
R23741 output.n60 output.n59 0.155672
R23742 output.n107 output.n79 0.155672
R23743 output.n100 output.n79 0.155672
R23744 output.n100 output.n99 0.155672
R23745 output.n99 output.n83 0.155672
R23746 output.n92 output.n83 0.155672
R23747 output.n92 output.n91 0.155672
R23748 output.n139 output.n111 0.155672
R23749 output.n132 output.n111 0.155672
R23750 output.n132 output.n131 0.155672
R23751 output.n131 output.n115 0.155672
R23752 output.n124 output.n115 0.155672
R23753 output.n124 output.n123 0.155672
R23754 output output.n14 0.126227
C0 output outputibias 2.34152f
C1 vdd output 7.23429f
C2 CSoutput output 6.13881f
C3 CSoutput outputibias 0.032386f
C4 vdd CSoutput 0.116623p
C5 commonsourceibias output 0.006808f
C6 minus diffpairibias 3.46e-19
C7 CSoutput minus 3.01338f
C8 vdd plus 0.085153f
C9 plus diffpairibias 2.47e-19
C10 commonsourceibias outputibias 0.003832f
C11 vdd commonsourceibias 0.004218f
C12 CSoutput plus 0.874205f
C13 commonsourceibias diffpairibias 0.064336f
C14 CSoutput commonsourceibias 54.554f
C15 minus plus 9.502349f
C16 minus commonsourceibias 0.331977f
C17 plus commonsourceibias 0.277692f
C18 diffpairibias gnd 60.00283f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.184151p
C22 plus gnd 33.4439f
C23 minus gnd 28.02365f
C24 CSoutput gnd 0.126253p
C25 vdd gnd 0.442313p
C26 output.t8 gnd 0.464308f
C27 output.t14 gnd 0.044422f
C28 output.t18 gnd 0.044422f
C29 output.n0 gnd 0.364624f
C30 output.n1 gnd 0.614102f
C31 output.t5 gnd 0.044422f
C32 output.t10 gnd 0.044422f
C33 output.n2 gnd 0.364624f
C34 output.n3 gnd 0.350265f
C35 output.t11 gnd 0.044422f
C36 output.t16 gnd 0.044422f
C37 output.n4 gnd 0.364624f
C38 output.n5 gnd 0.350265f
C39 output.t4 gnd 0.044422f
C40 output.t12 gnd 0.044422f
C41 output.n6 gnd 0.364624f
C42 output.n7 gnd 0.350265f
C43 output.t15 gnd 0.044422f
C44 output.t13 gnd 0.044422f
C45 output.n8 gnd 0.364624f
C46 output.n9 gnd 0.350265f
C47 output.t19 gnd 0.044422f
C48 output.t6 gnd 0.044422f
C49 output.n10 gnd 0.364624f
C50 output.n11 gnd 0.350265f
C51 output.t7 gnd 0.044422f
C52 output.t17 gnd 0.044422f
C53 output.n12 gnd 0.364624f
C54 output.n13 gnd 0.350265f
C55 output.t9 gnd 0.462979f
C56 output.n14 gnd 0.28994f
C57 output.n15 gnd 0.015803f
C58 output.n16 gnd 0.011243f
C59 output.n17 gnd 0.006041f
C60 output.n18 gnd 0.01428f
C61 output.n19 gnd 0.006397f
C62 output.n20 gnd 0.011243f
C63 output.n21 gnd 0.006041f
C64 output.n22 gnd 0.01428f
C65 output.n23 gnd 0.006397f
C66 output.n24 gnd 0.048111f
C67 output.t2 gnd 0.023274f
C68 output.n25 gnd 0.01071f
C69 output.n26 gnd 0.008435f
C70 output.n27 gnd 0.006041f
C71 output.n28 gnd 0.267512f
C72 output.n29 gnd 0.011243f
C73 output.n30 gnd 0.006041f
C74 output.n31 gnd 0.006397f
C75 output.n32 gnd 0.01428f
C76 output.n33 gnd 0.01428f
C77 output.n34 gnd 0.006397f
C78 output.n35 gnd 0.006041f
C79 output.n36 gnd 0.011243f
C80 output.n37 gnd 0.011243f
C81 output.n38 gnd 0.006041f
C82 output.n39 gnd 0.006397f
C83 output.n40 gnd 0.01428f
C84 output.n41 gnd 0.030913f
C85 output.n42 gnd 0.006397f
C86 output.n43 gnd 0.006041f
C87 output.n44 gnd 0.025987f
C88 output.n45 gnd 0.097665f
C89 output.n46 gnd 0.015803f
C90 output.n47 gnd 0.011243f
C91 output.n48 gnd 0.006041f
C92 output.n49 gnd 0.01428f
C93 output.n50 gnd 0.006397f
C94 output.n51 gnd 0.011243f
C95 output.n52 gnd 0.006041f
C96 output.n53 gnd 0.01428f
C97 output.n54 gnd 0.006397f
C98 output.n55 gnd 0.048111f
C99 output.t1 gnd 0.023274f
C100 output.n56 gnd 0.01071f
C101 output.n57 gnd 0.008435f
C102 output.n58 gnd 0.006041f
C103 output.n59 gnd 0.267512f
C104 output.n60 gnd 0.011243f
C105 output.n61 gnd 0.006041f
C106 output.n62 gnd 0.006397f
C107 output.n63 gnd 0.01428f
C108 output.n64 gnd 0.01428f
C109 output.n65 gnd 0.006397f
C110 output.n66 gnd 0.006041f
C111 output.n67 gnd 0.011243f
C112 output.n68 gnd 0.011243f
C113 output.n69 gnd 0.006041f
C114 output.n70 gnd 0.006397f
C115 output.n71 gnd 0.01428f
C116 output.n72 gnd 0.030913f
C117 output.n73 gnd 0.006397f
C118 output.n74 gnd 0.006041f
C119 output.n75 gnd 0.025987f
C120 output.n76 gnd 0.09306f
C121 output.n77 gnd 1.65264f
C122 output.n78 gnd 0.015803f
C123 output.n79 gnd 0.011243f
C124 output.n80 gnd 0.006041f
C125 output.n81 gnd 0.01428f
C126 output.n82 gnd 0.006397f
C127 output.n83 gnd 0.011243f
C128 output.n84 gnd 0.006041f
C129 output.n85 gnd 0.01428f
C130 output.n86 gnd 0.006397f
C131 output.n87 gnd 0.048111f
C132 output.t3 gnd 0.023274f
C133 output.n88 gnd 0.01071f
C134 output.n89 gnd 0.008435f
C135 output.n90 gnd 0.006041f
C136 output.n91 gnd 0.267512f
C137 output.n92 gnd 0.011243f
C138 output.n93 gnd 0.006041f
C139 output.n94 gnd 0.006397f
C140 output.n95 gnd 0.01428f
C141 output.n96 gnd 0.01428f
C142 output.n97 gnd 0.006397f
C143 output.n98 gnd 0.006041f
C144 output.n99 gnd 0.011243f
C145 output.n100 gnd 0.011243f
C146 output.n101 gnd 0.006041f
C147 output.n102 gnd 0.006397f
C148 output.n103 gnd 0.01428f
C149 output.n104 gnd 0.030913f
C150 output.n105 gnd 0.006397f
C151 output.n106 gnd 0.006041f
C152 output.n107 gnd 0.025987f
C153 output.n108 gnd 0.09306f
C154 output.n109 gnd 0.713089f
C155 output.n110 gnd 0.015803f
C156 output.n111 gnd 0.011243f
C157 output.n112 gnd 0.006041f
C158 output.n113 gnd 0.01428f
C159 output.n114 gnd 0.006397f
C160 output.n115 gnd 0.011243f
C161 output.n116 gnd 0.006041f
C162 output.n117 gnd 0.01428f
C163 output.n118 gnd 0.006397f
C164 output.n119 gnd 0.048111f
C165 output.t0 gnd 0.023274f
C166 output.n120 gnd 0.01071f
C167 output.n121 gnd 0.008435f
C168 output.n122 gnd 0.006041f
C169 output.n123 gnd 0.267512f
C170 output.n124 gnd 0.011243f
C171 output.n125 gnd 0.006041f
C172 output.n126 gnd 0.006397f
C173 output.n127 gnd 0.01428f
C174 output.n128 gnd 0.01428f
C175 output.n129 gnd 0.006397f
C176 output.n130 gnd 0.006041f
C177 output.n131 gnd 0.011243f
C178 output.n132 gnd 0.011243f
C179 output.n133 gnd 0.006041f
C180 output.n134 gnd 0.006397f
C181 output.n135 gnd 0.01428f
C182 output.n136 gnd 0.030913f
C183 output.n137 gnd 0.006397f
C184 output.n138 gnd 0.006041f
C185 output.n139 gnd 0.025987f
C186 output.n140 gnd 0.09306f
C187 output.n141 gnd 1.67353f
C188 outputibias.t10 gnd 0.11477f
C189 outputibias.t9 gnd 0.115567f
C190 outputibias.n0 gnd 0.130108f
C191 outputibias.n1 gnd 0.001372f
C192 outputibias.n2 gnd 9.76e-19
C193 outputibias.n3 gnd 5.24e-19
C194 outputibias.n4 gnd 0.001239f
C195 outputibias.n5 gnd 5.55e-19
C196 outputibias.n6 gnd 9.76e-19
C197 outputibias.n7 gnd 5.24e-19
C198 outputibias.n8 gnd 0.001239f
C199 outputibias.n9 gnd 5.55e-19
C200 outputibias.n10 gnd 0.004176f
C201 outputibias.t5 gnd 0.00202f
C202 outputibias.n11 gnd 9.3e-19
C203 outputibias.n12 gnd 7.32e-19
C204 outputibias.n13 gnd 5.24e-19
C205 outputibias.n14 gnd 0.02322f
C206 outputibias.n15 gnd 9.76e-19
C207 outputibias.n16 gnd 5.24e-19
C208 outputibias.n17 gnd 5.55e-19
C209 outputibias.n18 gnd 0.001239f
C210 outputibias.n19 gnd 0.001239f
C211 outputibias.n20 gnd 5.55e-19
C212 outputibias.n21 gnd 5.24e-19
C213 outputibias.n22 gnd 9.76e-19
C214 outputibias.n23 gnd 9.76e-19
C215 outputibias.n24 gnd 5.24e-19
C216 outputibias.n25 gnd 5.55e-19
C217 outputibias.n26 gnd 0.001239f
C218 outputibias.n27 gnd 0.002683f
C219 outputibias.n28 gnd 5.55e-19
C220 outputibias.n29 gnd 5.24e-19
C221 outputibias.n30 gnd 0.002256f
C222 outputibias.n31 gnd 0.005781f
C223 outputibias.n32 gnd 0.001372f
C224 outputibias.n33 gnd 9.76e-19
C225 outputibias.n34 gnd 5.24e-19
C226 outputibias.n35 gnd 0.001239f
C227 outputibias.n36 gnd 5.55e-19
C228 outputibias.n37 gnd 9.76e-19
C229 outputibias.n38 gnd 5.24e-19
C230 outputibias.n39 gnd 0.001239f
C231 outputibias.n40 gnd 5.55e-19
C232 outputibias.n41 gnd 0.004176f
C233 outputibias.t7 gnd 0.00202f
C234 outputibias.n42 gnd 9.3e-19
C235 outputibias.n43 gnd 7.32e-19
C236 outputibias.n44 gnd 5.24e-19
C237 outputibias.n45 gnd 0.02322f
C238 outputibias.n46 gnd 9.76e-19
C239 outputibias.n47 gnd 5.24e-19
C240 outputibias.n48 gnd 5.55e-19
C241 outputibias.n49 gnd 0.001239f
C242 outputibias.n50 gnd 0.001239f
C243 outputibias.n51 gnd 5.55e-19
C244 outputibias.n52 gnd 5.24e-19
C245 outputibias.n53 gnd 9.76e-19
C246 outputibias.n54 gnd 9.76e-19
C247 outputibias.n55 gnd 5.24e-19
C248 outputibias.n56 gnd 5.55e-19
C249 outputibias.n57 gnd 0.001239f
C250 outputibias.n58 gnd 0.002683f
C251 outputibias.n59 gnd 5.55e-19
C252 outputibias.n60 gnd 5.24e-19
C253 outputibias.n61 gnd 0.002256f
C254 outputibias.n62 gnd 0.005197f
C255 outputibias.n63 gnd 0.121892f
C256 outputibias.n64 gnd 0.001372f
C257 outputibias.n65 gnd 9.76e-19
C258 outputibias.n66 gnd 5.24e-19
C259 outputibias.n67 gnd 0.001239f
C260 outputibias.n68 gnd 5.55e-19
C261 outputibias.n69 gnd 9.76e-19
C262 outputibias.n70 gnd 5.24e-19
C263 outputibias.n71 gnd 0.001239f
C264 outputibias.n72 gnd 5.55e-19
C265 outputibias.n73 gnd 0.004176f
C266 outputibias.t1 gnd 0.00202f
C267 outputibias.n74 gnd 9.3e-19
C268 outputibias.n75 gnd 7.32e-19
C269 outputibias.n76 gnd 5.24e-19
C270 outputibias.n77 gnd 0.02322f
C271 outputibias.n78 gnd 9.76e-19
C272 outputibias.n79 gnd 5.24e-19
C273 outputibias.n80 gnd 5.55e-19
C274 outputibias.n81 gnd 0.001239f
C275 outputibias.n82 gnd 0.001239f
C276 outputibias.n83 gnd 5.55e-19
C277 outputibias.n84 gnd 5.24e-19
C278 outputibias.n85 gnd 9.76e-19
C279 outputibias.n86 gnd 9.76e-19
C280 outputibias.n87 gnd 5.24e-19
C281 outputibias.n88 gnd 5.55e-19
C282 outputibias.n89 gnd 0.001239f
C283 outputibias.n90 gnd 0.002683f
C284 outputibias.n91 gnd 5.55e-19
C285 outputibias.n92 gnd 5.24e-19
C286 outputibias.n93 gnd 0.002256f
C287 outputibias.n94 gnd 0.005197f
C288 outputibias.n95 gnd 0.064513f
C289 outputibias.n96 gnd 0.001372f
C290 outputibias.n97 gnd 9.76e-19
C291 outputibias.n98 gnd 5.24e-19
C292 outputibias.n99 gnd 0.001239f
C293 outputibias.n100 gnd 5.55e-19
C294 outputibias.n101 gnd 9.76e-19
C295 outputibias.n102 gnd 5.24e-19
C296 outputibias.n103 gnd 0.001239f
C297 outputibias.n104 gnd 5.55e-19
C298 outputibias.n105 gnd 0.004176f
C299 outputibias.t3 gnd 0.00202f
C300 outputibias.n106 gnd 9.3e-19
C301 outputibias.n107 gnd 7.32e-19
C302 outputibias.n108 gnd 5.24e-19
C303 outputibias.n109 gnd 0.02322f
C304 outputibias.n110 gnd 9.76e-19
C305 outputibias.n111 gnd 5.24e-19
C306 outputibias.n112 gnd 5.55e-19
C307 outputibias.n113 gnd 0.001239f
C308 outputibias.n114 gnd 0.001239f
C309 outputibias.n115 gnd 5.55e-19
C310 outputibias.n116 gnd 5.24e-19
C311 outputibias.n117 gnd 9.76e-19
C312 outputibias.n118 gnd 9.76e-19
C313 outputibias.n119 gnd 5.24e-19
C314 outputibias.n120 gnd 5.55e-19
C315 outputibias.n121 gnd 0.001239f
C316 outputibias.n122 gnd 0.002683f
C317 outputibias.n123 gnd 5.55e-19
C318 outputibias.n124 gnd 5.24e-19
C319 outputibias.n125 gnd 0.002256f
C320 outputibias.n126 gnd 0.005197f
C321 outputibias.n127 gnd 0.084814f
C322 outputibias.t2 gnd 0.108319f
C323 outputibias.t0 gnd 0.108319f
C324 outputibias.t6 gnd 0.108319f
C325 outputibias.t4 gnd 0.109238f
C326 outputibias.n128 gnd 0.134674f
C327 outputibias.n129 gnd 0.07244f
C328 outputibias.n130 gnd 0.079818f
C329 outputibias.n131 gnd 0.164901f
C330 outputibias.t11 gnd 0.11477f
C331 outputibias.n132 gnd 0.067481f
C332 outputibias.t8 gnd 0.11477f
C333 outputibias.n133 gnd 0.065115f
C334 outputibias.n134 gnd 0.029159f
C335 a_n2318_8322.t27 gnd 39.5861f
C336 a_n2318_8322.t24 gnd 29.0796f
C337 a_n2318_8322.t26 gnd 19.7234f
C338 a_n2318_8322.t25 gnd 39.5861f
C339 a_n2318_8322.t12 gnd 0.095743f
C340 a_n2318_8322.t22 gnd 0.896485f
C341 a_n2318_8322.t10 gnd 0.095743f
C342 a_n2318_8322.t9 gnd 0.095743f
C343 a_n2318_8322.n0 gnd 0.674411f
C344 a_n2318_8322.n1 gnd 0.753555f
C345 a_n2318_8322.t19 gnd 0.095743f
C346 a_n2318_8322.t14 gnd 0.095743f
C347 a_n2318_8322.n2 gnd 0.674411f
C348 a_n2318_8322.n3 gnd 0.382872f
C349 a_n2318_8322.t17 gnd 0.095743f
C350 a_n2318_8322.t16 gnd 0.095743f
C351 a_n2318_8322.n4 gnd 0.674411f
C352 a_n2318_8322.n5 gnd 0.382872f
C353 a_n2318_8322.t8 gnd 0.8947f
C354 a_n2318_8322.n6 gnd 1.55065f
C355 a_n2318_8322.t3 gnd 0.896485f
C356 a_n2318_8322.t7 gnd 0.095743f
C357 a_n2318_8322.t6 gnd 0.095743f
C358 a_n2318_8322.n7 gnd 0.674411f
C359 a_n2318_8322.n8 gnd 0.753555f
C360 a_n2318_8322.t1 gnd 0.8947f
C361 a_n2318_8322.n9 gnd 0.379199f
C362 a_n2318_8322.t4 gnd 0.8947f
C363 a_n2318_8322.n10 gnd 0.379199f
C364 a_n2318_8322.t2 gnd 0.095743f
C365 a_n2318_8322.t0 gnd 0.095743f
C366 a_n2318_8322.n11 gnd 0.674411f
C367 a_n2318_8322.n12 gnd 0.382872f
C368 a_n2318_8322.t5 gnd 0.8947f
C369 a_n2318_8322.n13 gnd 1.0738f
C370 a_n2318_8322.n14 gnd 1.82539f
C371 a_n2318_8322.n15 gnd 3.67064f
C372 a_n2318_8322.t11 gnd 0.8947f
C373 a_n2318_8322.n16 gnd 0.880763f
C374 a_n2318_8322.t20 gnd 0.095743f
C375 a_n2318_8322.t13 gnd 0.095743f
C376 a_n2318_8322.n17 gnd 0.674411f
C377 a_n2318_8322.n18 gnd 0.382872f
C378 a_n2318_8322.t21 gnd 0.896483f
C379 a_n2318_8322.t18 gnd 0.095743f
C380 a_n2318_8322.t15 gnd 0.095743f
C381 a_n2318_8322.n19 gnd 0.674411f
C382 a_n2318_8322.n20 gnd 0.753557f
C383 a_n2318_8322.n21 gnd 0.38287f
C384 a_n2318_8322.n22 gnd 0.674413f
C385 a_n2318_8322.t23 gnd 0.095743f
C386 minus.n0 gnd 0.029476f
C387 minus.t14 gnd 0.495627f
C388 minus.n1 gnd 0.200454f
C389 minus.n2 gnd 0.029476f
C390 minus.t19 gnd 0.495627f
C391 minus.n3 gnd 0.023957f
C392 minus.n4 gnd 0.029476f
C393 minus.t18 gnd 0.495627f
C394 minus.t5 gnd 0.495627f
C395 minus.n5 gnd 0.200454f
C396 minus.n6 gnd 0.029476f
C397 minus.t8 gnd 0.495627f
C398 minus.n7 gnd 0.200454f
C399 minus.n8 gnd 0.126527f
C400 minus.t9 gnd 0.495627f
C401 minus.t13 gnd 0.556459f
C402 minus.n9 gnd 0.232581f
C403 minus.n10 gnd 0.231493f
C404 minus.n11 gnd 0.036665f
C405 minus.n12 gnd 0.034458f
C406 minus.n13 gnd 0.029476f
C407 minus.n14 gnd 0.029476f
C408 minus.n15 gnd 0.036923f
C409 minus.n16 gnd 0.023957f
C410 minus.n17 gnd 0.037919f
C411 minus.n18 gnd 0.029476f
C412 minus.n19 gnd 0.029476f
C413 minus.n20 gnd 0.035562f
C414 minus.n21 gnd 0.035562f
C415 minus.n22 gnd 0.200454f
C416 minus.n23 gnd 0.037919f
C417 minus.n24 gnd 0.029476f
C418 minus.n25 gnd 0.029476f
C419 minus.n26 gnd 0.029476f
C420 minus.n27 gnd 0.036923f
C421 minus.n28 gnd 0.200454f
C422 minus.n29 gnd 0.034458f
C423 minus.n30 gnd 0.036665f
C424 minus.n31 gnd 0.029476f
C425 minus.n32 gnd 0.029476f
C426 minus.n33 gnd 0.038388f
C427 minus.n34 gnd 0.012208f
C428 minus.t17 gnd 0.536021f
C429 minus.n35 gnd 0.232818f
C430 minus.n36 gnd 0.346343f
C431 minus.n37 gnd 0.029476f
C432 minus.t15 gnd 0.536021f
C433 minus.t12 gnd 0.495627f
C434 minus.n38 gnd 0.200454f
C435 minus.n39 gnd 0.029476f
C436 minus.t7 gnd 0.495627f
C437 minus.n40 gnd 0.023957f
C438 minus.n41 gnd 0.029476f
C439 minus.t6 gnd 0.495627f
C440 minus.t11 gnd 0.495627f
C441 minus.n42 gnd 0.200454f
C442 minus.n43 gnd 0.029476f
C443 minus.t10 gnd 0.495627f
C444 minus.n44 gnd 0.200454f
C445 minus.n45 gnd 0.126527f
C446 minus.t16 gnd 0.495627f
C447 minus.t20 gnd 0.556459f
C448 minus.n46 gnd 0.232581f
C449 minus.n47 gnd 0.231493f
C450 minus.n48 gnd 0.036665f
C451 minus.n49 gnd 0.034458f
C452 minus.n50 gnd 0.029476f
C453 minus.n51 gnd 0.029476f
C454 minus.n52 gnd 0.036923f
C455 minus.n53 gnd 0.023957f
C456 minus.n54 gnd 0.037919f
C457 minus.n55 gnd 0.029476f
C458 minus.n56 gnd 0.029476f
C459 minus.n57 gnd 0.035562f
C460 minus.n58 gnd 0.035562f
C461 minus.n59 gnd 0.200454f
C462 minus.n60 gnd 0.037919f
C463 minus.n61 gnd 0.029476f
C464 minus.n62 gnd 0.029476f
C465 minus.n63 gnd 0.029476f
C466 minus.n64 gnd 0.036923f
C467 minus.n65 gnd 0.200454f
C468 minus.n66 gnd 0.034458f
C469 minus.n67 gnd 0.036665f
C470 minus.n68 gnd 0.029476f
C471 minus.n69 gnd 0.029476f
C472 minus.n70 gnd 0.038388f
C473 minus.n71 gnd 0.012208f
C474 minus.n72 gnd 0.232818f
C475 minus.n73 gnd 0.918445f
C476 minus.n74 gnd 1.3805f
C477 minus.t1 gnd 0.009087f
C478 minus.t4 gnd 0.009087f
C479 minus.n75 gnd 0.029878f
C480 minus.t2 gnd 0.009087f
C481 minus.t0 gnd 0.009087f
C482 minus.n76 gnd 0.029469f
C483 minus.n77 gnd 0.251504f
C484 minus.t3 gnd 0.050574f
C485 minus.n78 gnd 0.137244f
C486 minus.n79 gnd 2.05319f
C487 diffpairibias.t27 gnd 0.090128f
C488 diffpairibias.t23 gnd 0.08996f
C489 diffpairibias.n0 gnd 0.105991f
C490 diffpairibias.t28 gnd 0.08996f
C491 diffpairibias.n1 gnd 0.051736f
C492 diffpairibias.t25 gnd 0.08996f
C493 diffpairibias.n2 gnd 0.051736f
C494 diffpairibias.t29 gnd 0.08996f
C495 diffpairibias.n3 gnd 0.041084f
C496 diffpairibias.t15 gnd 0.086371f
C497 diffpairibias.t1 gnd 0.085993f
C498 diffpairibias.n4 gnd 0.13579f
C499 diffpairibias.t11 gnd 0.085993f
C500 diffpairibias.n5 gnd 0.072463f
C501 diffpairibias.t13 gnd 0.085993f
C502 diffpairibias.n6 gnd 0.072463f
C503 diffpairibias.t7 gnd 0.085993f
C504 diffpairibias.n7 gnd 0.072463f
C505 diffpairibias.t3 gnd 0.085993f
C506 diffpairibias.n8 gnd 0.072463f
C507 diffpairibias.t17 gnd 0.085993f
C508 diffpairibias.n9 gnd 0.072463f
C509 diffpairibias.t5 gnd 0.085993f
C510 diffpairibias.n10 gnd 0.072463f
C511 diffpairibias.t19 gnd 0.085993f
C512 diffpairibias.n11 gnd 0.072463f
C513 diffpairibias.t9 gnd 0.085993f
C514 diffpairibias.n12 gnd 0.102883f
C515 diffpairibias.t14 gnd 0.086899f
C516 diffpairibias.t0 gnd 0.086748f
C517 diffpairibias.n13 gnd 0.094648f
C518 diffpairibias.t10 gnd 0.086748f
C519 diffpairibias.n14 gnd 0.052262f
C520 diffpairibias.t12 gnd 0.086748f
C521 diffpairibias.n15 gnd 0.052262f
C522 diffpairibias.t6 gnd 0.086748f
C523 diffpairibias.n16 gnd 0.052262f
C524 diffpairibias.t2 gnd 0.086748f
C525 diffpairibias.n17 gnd 0.052262f
C526 diffpairibias.t16 gnd 0.086748f
C527 diffpairibias.n18 gnd 0.052262f
C528 diffpairibias.t4 gnd 0.086748f
C529 diffpairibias.n19 gnd 0.052262f
C530 diffpairibias.t18 gnd 0.086748f
C531 diffpairibias.n20 gnd 0.052262f
C532 diffpairibias.t8 gnd 0.086748f
C533 diffpairibias.n21 gnd 0.061849f
C534 diffpairibias.n22 gnd 0.233513f
C535 diffpairibias.t20 gnd 0.08996f
C536 diffpairibias.n23 gnd 0.051747f
C537 diffpairibias.t26 gnd 0.08996f
C538 diffpairibias.n24 gnd 0.051736f
C539 diffpairibias.t22 gnd 0.08996f
C540 diffpairibias.n25 gnd 0.051736f
C541 diffpairibias.t21 gnd 0.08996f
C542 diffpairibias.n26 gnd 0.051736f
C543 diffpairibias.t24 gnd 0.08996f
C544 diffpairibias.n27 gnd 0.04729f
C545 diffpairibias.n28 gnd 0.047711f
C546 a_n3827_n3924.n0 gnd 0.8843f
C547 a_n3827_n3924.t16 gnd 0.083157f
C548 a_n3827_n3924.t25 gnd 0.864269f
C549 a_n3827_n3924.n1 gnd 0.326732f
C550 a_n3827_n3924.t10 gnd 1.07678f
C551 a_n3827_n3924.t6 gnd 1.07383f
C552 a_n3827_n3924.n2 gnd 1.46419f
C553 a_n3827_n3924.n3 gnd 0.408778f
C554 a_n3827_n3924.t36 gnd 0.864269f
C555 a_n3827_n3924.n4 gnd 0.326732f
C556 a_n3827_n3924.t41 gnd 0.083157f
C557 a_n3827_n3924.t33 gnd 0.083157f
C558 a_n3827_n3924.n5 gnd 0.67916f
C559 a_n3827_n3924.n6 gnd 0.342258f
C560 a_n3827_n3924.t4 gnd 0.083157f
C561 a_n3827_n3924.t35 gnd 0.083157f
C562 a_n3827_n3924.n7 gnd 0.67916f
C563 a_n3827_n3924.n8 gnd 0.342258f
C564 a_n3827_n3924.t34 gnd 0.083157f
C565 a_n3827_n3924.t13 gnd 0.083157f
C566 a_n3827_n3924.n9 gnd 0.67916f
C567 a_n3827_n3924.n10 gnd 0.342258f
C568 a_n3827_n3924.t8 gnd 0.864269f
C569 a_n3827_n3924.n11 gnd 0.809022f
C570 a_n3827_n3924.t0 gnd 1.07537f
C571 a_n3827_n3924.t11 gnd 1.07383f
C572 a_n3827_n3924.n12 gnd 1.24022f
C573 a_n3827_n3924.t12 gnd 1.07383f
C574 a_n3827_n3924.n13 gnd 0.700903f
C575 a_n3827_n3924.t37 gnd 1.07383f
C576 a_n3827_n3924.n14 gnd 0.75632f
C577 a_n3827_n3924.t38 gnd 1.07383f
C578 a_n3827_n3924.n15 gnd 0.75632f
C579 a_n3827_n3924.t1 gnd 1.07383f
C580 a_n3827_n3924.n16 gnd 0.75632f
C581 a_n3827_n3924.t5 gnd 1.07383f
C582 a_n3827_n3924.n17 gnd 0.75632f
C583 a_n3827_n3924.t30 gnd 1.07383f
C584 a_n3827_n3924.n18 gnd 0.783961f
C585 a_n3827_n3924.t27 gnd 0.864266f
C586 a_n3827_n3924.n19 gnd 0.536839f
C587 a_n3827_n3924.t28 gnd 0.083157f
C588 a_n3827_n3924.t18 gnd 0.083157f
C589 a_n3827_n3924.n20 gnd 0.679159f
C590 a_n3827_n3924.n21 gnd 0.342259f
C591 a_n3827_n3924.t19 gnd 0.083157f
C592 a_n3827_n3924.t14 gnd 0.083157f
C593 a_n3827_n3924.n22 gnd 0.679159f
C594 a_n3827_n3924.n23 gnd 0.342259f
C595 a_n3827_n3924.t15 gnd 0.083157f
C596 a_n3827_n3924.t26 gnd 0.083157f
C597 a_n3827_n3924.n24 gnd 0.679159f
C598 a_n3827_n3924.n25 gnd 0.342259f
C599 a_n3827_n3924.t23 gnd 0.864266f
C600 a_n3827_n3924.n26 gnd 0.326736f
C601 a_n3827_n3924.t3 gnd 0.864266f
C602 a_n3827_n3924.n27 gnd 0.326736f
C603 a_n3827_n3924.t9 gnd 0.083157f
C604 a_n3827_n3924.t40 gnd 0.083157f
C605 a_n3827_n3924.n28 gnd 0.679159f
C606 a_n3827_n3924.n29 gnd 0.342259f
C607 a_n3827_n3924.t39 gnd 0.083157f
C608 a_n3827_n3924.t32 gnd 0.083157f
C609 a_n3827_n3924.n30 gnd 0.679159f
C610 a_n3827_n3924.n31 gnd 0.342259f
C611 a_n3827_n3924.t7 gnd 0.083157f
C612 a_n3827_n3924.t2 gnd 0.083157f
C613 a_n3827_n3924.n32 gnd 0.679159f
C614 a_n3827_n3924.n33 gnd 0.342259f
C615 a_n3827_n3924.t31 gnd 0.864266f
C616 a_n3827_n3924.n34 gnd 0.536839f
C617 a_n3827_n3924.n35 gnd 0.783961f
C618 a_n3827_n3924.t22 gnd 0.864266f
C619 a_n3827_n3924.n36 gnd 0.809025f
C620 a_n3827_n3924.t20 gnd 0.083157f
C621 a_n3827_n3924.t24 gnd 0.083157f
C622 a_n3827_n3924.n37 gnd 0.67916f
C623 a_n3827_n3924.n38 gnd 0.342258f
C624 a_n3827_n3924.t17 gnd 0.083157f
C625 a_n3827_n3924.t21 gnd 0.083157f
C626 a_n3827_n3924.n39 gnd 0.67916f
C627 a_n3827_n3924.n40 gnd 0.342258f
C628 a_n3827_n3924.n41 gnd 0.342257f
C629 a_n3827_n3924.n42 gnd 0.679161f
C630 a_n3827_n3924.t29 gnd 0.083157f
C631 plus.n0 gnd 0.021653f
C632 plus.t7 gnd 0.393769f
C633 plus.t6 gnd 0.364095f
C634 plus.n1 gnd 0.147256f
C635 plus.n2 gnd 0.021653f
C636 plus.t16 gnd 0.364095f
C637 plus.n3 gnd 0.017599f
C638 plus.n4 gnd 0.021653f
C639 plus.t15 gnd 0.364095f
C640 plus.t20 gnd 0.364095f
C641 plus.n5 gnd 0.147256f
C642 plus.n6 gnd 0.021653f
C643 plus.t19 gnd 0.364095f
C644 plus.n7 gnd 0.147256f
C645 plus.n8 gnd 0.092948f
C646 plus.t8 gnd 0.364095f
C647 plus.t11 gnd 0.408783f
C648 plus.n9 gnd 0.170858f
C649 plus.n10 gnd 0.170058f
C650 plus.n11 gnd 0.026935f
C651 plus.n12 gnd 0.025314f
C652 plus.n13 gnd 0.021653f
C653 plus.n14 gnd 0.021653f
C654 plus.n15 gnd 0.027124f
C655 plus.n16 gnd 0.017599f
C656 plus.n17 gnd 0.027856f
C657 plus.n18 gnd 0.021653f
C658 plus.n19 gnd 0.021653f
C659 plus.n20 gnd 0.026124f
C660 plus.n21 gnd 0.026124f
C661 plus.n22 gnd 0.147256f
C662 plus.n23 gnd 0.027856f
C663 plus.n24 gnd 0.021653f
C664 plus.n25 gnd 0.021653f
C665 plus.n26 gnd 0.021653f
C666 plus.n27 gnd 0.027124f
C667 plus.n28 gnd 0.147256f
C668 plus.n29 gnd 0.025314f
C669 plus.n30 gnd 0.026935f
C670 plus.n31 gnd 0.021653f
C671 plus.n32 gnd 0.021653f
C672 plus.n33 gnd 0.0282f
C673 plus.n34 gnd 0.008968f
C674 plus.n35 gnd 0.171032f
C675 plus.n36 gnd 0.24886f
C676 plus.n37 gnd 0.021653f
C677 plus.t10 gnd 0.364095f
C678 plus.n38 gnd 0.147256f
C679 plus.n39 gnd 0.021653f
C680 plus.t14 gnd 0.364095f
C681 plus.n40 gnd 0.017599f
C682 plus.n41 gnd 0.021653f
C683 plus.t13 gnd 0.364095f
C684 plus.t17 gnd 0.364095f
C685 plus.n42 gnd 0.147256f
C686 plus.n43 gnd 0.021653f
C687 plus.t18 gnd 0.364095f
C688 plus.n44 gnd 0.147256f
C689 plus.n45 gnd 0.092948f
C690 plus.t5 gnd 0.364095f
C691 plus.t9 gnd 0.408783f
C692 plus.n46 gnd 0.170858f
C693 plus.n47 gnd 0.170058f
C694 plus.n48 gnd 0.026935f
C695 plus.n49 gnd 0.025314f
C696 plus.n50 gnd 0.021653f
C697 plus.n51 gnd 0.021653f
C698 plus.n52 gnd 0.027124f
C699 plus.n53 gnd 0.017599f
C700 plus.n54 gnd 0.027856f
C701 plus.n55 gnd 0.021653f
C702 plus.n56 gnd 0.021653f
C703 plus.n57 gnd 0.026124f
C704 plus.n58 gnd 0.026124f
C705 plus.n59 gnd 0.147256f
C706 plus.n60 gnd 0.027856f
C707 plus.n61 gnd 0.021653f
C708 plus.n62 gnd 0.021653f
C709 plus.n63 gnd 0.021653f
C710 plus.n64 gnd 0.027124f
C711 plus.n65 gnd 0.147256f
C712 plus.n66 gnd 0.025314f
C713 plus.n67 gnd 0.026935f
C714 plus.n68 gnd 0.021653f
C715 plus.n69 gnd 0.021653f
C716 plus.n70 gnd 0.0282f
C717 plus.n71 gnd 0.008968f
C718 plus.t12 gnd 0.393769f
C719 plus.n72 gnd 0.171032f
C720 plus.n73 gnd 0.666028f
C721 plus.n74 gnd 1.00555f
C722 plus.t4 gnd 0.03738f
C723 plus.t1 gnd 0.006675f
C724 plus.t2 gnd 0.006675f
C725 plus.n75 gnd 0.021648f
C726 plus.n76 gnd 0.168058f
C727 plus.t0 gnd 0.006675f
C728 plus.t3 gnd 0.006675f
C729 plus.n77 gnd 0.021648f
C730 plus.n78 gnd 0.126148f
C731 plus.n79 gnd 2.62972f
C732 a_n2140_13878.t11 gnd 0.186868f
C733 a_n2140_13878.t10 gnd 0.186868f
C734 a_n2140_13878.t5 gnd 0.186868f
C735 a_n2140_13878.n0 gnd 1.47299f
C736 a_n2140_13878.t2 gnd 0.186868f
C737 a_n2140_13878.t4 gnd 0.186868f
C738 a_n2140_13878.n1 gnd 1.47143f
C739 a_n2140_13878.n2 gnd 2.05603f
C740 a_n2140_13878.t12 gnd 0.186868f
C741 a_n2140_13878.t3 gnd 0.186868f
C742 a_n2140_13878.n3 gnd 1.47143f
C743 a_n2140_13878.n4 gnd 1.00289f
C744 a_n2140_13878.t9 gnd 0.186868f
C745 a_n2140_13878.t1 gnd 0.186868f
C746 a_n2140_13878.n5 gnd 1.47143f
C747 a_n2140_13878.n6 gnd 4.06212f
C748 a_n2140_13878.t17 gnd 1.74974f
C749 a_n2140_13878.t20 gnd 0.186868f
C750 a_n2140_13878.t21 gnd 0.186868f
C751 a_n2140_13878.n7 gnd 1.3163f
C752 a_n2140_13878.n8 gnd 1.47077f
C753 a_n2140_13878.t16 gnd 1.74626f
C754 a_n2140_13878.n9 gnd 0.740113f
C755 a_n2140_13878.t19 gnd 1.74626f
C756 a_n2140_13878.n10 gnd 0.740113f
C757 a_n2140_13878.t22 gnd 0.186868f
C758 a_n2140_13878.t23 gnd 0.186868f
C759 a_n2140_13878.n11 gnd 1.3163f
C760 a_n2140_13878.n12 gnd 0.74728f
C761 a_n2140_13878.t18 gnd 1.74626f
C762 a_n2140_13878.n13 gnd 2.09583f
C763 a_n2140_13878.n14 gnd 2.85974f
C764 a_n2140_13878.t6 gnd 0.186868f
C765 a_n2140_13878.t7 gnd 0.186868f
C766 a_n2140_13878.n15 gnd 1.47142f
C767 a_n2140_13878.n16 gnd 2.01665f
C768 a_n2140_13878.t13 gnd 0.186868f
C769 a_n2140_13878.t14 gnd 0.186868f
C770 a_n2140_13878.n17 gnd 1.47143f
C771 a_n2140_13878.n18 gnd 0.651951f
C772 a_n2140_13878.t0 gnd 0.186868f
C773 a_n2140_13878.t8 gnd 0.186868f
C774 a_n2140_13878.n19 gnd 1.47143f
C775 a_n2140_13878.n20 gnd 1.32263f
C776 a_n2140_13878.n21 gnd 1.47386f
C777 a_n2140_13878.t15 gnd 0.186868f
C778 a_n2318_13878.n0 gnd 2.73227f
C779 a_n2318_13878.n1 gnd 3.94723f
C780 a_n2318_13878.n2 gnd 3.81658f
C781 a_n2318_13878.n3 gnd 0.652811f
C782 a_n2318_13878.n4 gnd 0.210856f
C783 a_n2318_13878.n5 gnd 0.210856f
C784 a_n2318_13878.n6 gnd 0.729399f
C785 a_n2318_13878.n7 gnd 0.210856f
C786 a_n2318_13878.n8 gnd 0.433021f
C787 a_n2318_13878.n9 gnd 0.652788f
C788 a_n2318_13878.n10 gnd 0.200068f
C789 a_n2318_13878.n11 gnd 0.147354f
C790 a_n2318_13878.n12 gnd 0.231593f
C791 a_n2318_13878.n13 gnd 0.178879f
C792 a_n2318_13878.n14 gnd 0.200068f
C793 a_n2318_13878.n15 gnd 1.09189f
C794 a_n2318_13878.n16 gnd 0.147354f
C795 a_n2318_13878.n17 gnd 0.705502f
C796 a_n2318_13878.n18 gnd 0.50033f
C797 a_n2318_13878.n19 gnd 0.210856f
C798 a_n2318_13878.n20 gnd 0.210856f
C799 a_n2318_13878.n21 gnd 0.433358f
C800 a_n2318_13878.n22 gnd 0.210856f
C801 a_n2318_13878.n23 gnd 0.210856f
C802 a_n2318_13878.n24 gnd 1.73596f
C803 a_n2318_13878.n25 gnd 2.03016f
C804 a_n2318_13878.n26 gnd 1.85287f
C805 a_n2318_13878.n27 gnd 1.73595f
C806 a_n2318_13878.n28 gnd 3.14412f
C807 a_n2318_13878.n29 gnd 0.278541f
C808 a_n2318_13878.n30 gnd 0.742063f
C809 a_n2318_13878.n31 gnd 0.004739f
C810 a_n2318_13878.n32 gnd 0.01025f
C811 a_n2318_13878.n33 gnd 0.01025f
C812 a_n2318_13878.n34 gnd 0.004739f
C813 a_n2318_13878.n35 gnd 0.278541f
C814 a_n2318_13878.n36 gnd 0.278541f
C815 a_n2318_13878.n37 gnd 0.433358f
C816 a_n2318_13878.n38 gnd 0.004739f
C817 a_n2318_13878.n39 gnd 0.01025f
C818 a_n2318_13878.n40 gnd 0.01025f
C819 a_n2318_13878.n41 gnd 0.004739f
C820 a_n2318_13878.n42 gnd 0.278541f
C821 a_n2318_13878.n43 gnd 0.008164f
C822 a_n2318_13878.n44 gnd 0.278541f
C823 a_n2318_13878.n45 gnd 0.008164f
C824 a_n2318_13878.n46 gnd 0.278541f
C825 a_n2318_13878.n47 gnd 0.008164f
C826 a_n2318_13878.n48 gnd 0.278541f
C827 a_n2318_13878.n49 gnd 0.008164f
C828 a_n2318_13878.n50 gnd 0.278541f
C829 a_n2318_13878.n51 gnd 0.278541f
C830 a_n2318_13878.n52 gnd 0.004739f
C831 a_n2318_13878.n53 gnd 0.01025f
C832 a_n2318_13878.n54 gnd 0.01025f
C833 a_n2318_13878.n55 gnd 0.004739f
C834 a_n2318_13878.n56 gnd 0.278541f
C835 a_n2318_13878.n57 gnd 0.278541f
C836 a_n2318_13878.n58 gnd 0.004739f
C837 a_n2318_13878.n59 gnd 0.01025f
C838 a_n2318_13878.n60 gnd 0.105428f
C839 a_n2318_13878.n61 gnd 0.01025f
C840 a_n2318_13878.n62 gnd 0.004739f
C841 a_n2318_13878.n63 gnd 0.278541f
C842 a_n2318_13878.t28 gnd 0.146252f
C843 a_n2318_13878.t31 gnd 0.691694f
C844 a_n2318_13878.t15 gnd 0.680295f
C845 a_n2318_13878.t17 gnd 0.680295f
C846 a_n2318_13878.n64 gnd 0.297177f
C847 a_n2318_13878.t27 gnd 0.680295f
C848 a_n2318_13878.t3 gnd 0.680295f
C849 a_n2318_13878.t9 gnd 0.680295f
C850 a_n2318_13878.n65 gnd 0.297177f
C851 a_n2318_13878.t5 gnd 0.680295f
C852 a_n2318_13878.t25 gnd 0.691694f
C853 a_n2318_13878.t1 gnd 0.113752f
C854 a_n2318_13878.t37 gnd 0.113752f
C855 a_n2318_13878.n66 gnd 1.00811f
C856 a_n2318_13878.t46 gnd 0.113752f
C857 a_n2318_13878.t45 gnd 0.113752f
C858 a_n2318_13878.n67 gnd 1.00515f
C859 a_n2318_13878.t0 gnd 0.113752f
C860 a_n2318_13878.t39 gnd 0.113752f
C861 a_n2318_13878.n68 gnd 1.00811f
C862 a_n2318_13878.t40 gnd 0.113752f
C863 a_n2318_13878.t35 gnd 0.113752f
C864 a_n2318_13878.n69 gnd 1.00515f
C865 a_n2318_13878.t36 gnd 0.113752f
C866 a_n2318_13878.t42 gnd 0.113752f
C867 a_n2318_13878.n70 gnd 1.00515f
C868 a_n2318_13878.t38 gnd 0.113752f
C869 a_n2318_13878.t2 gnd 0.113752f
C870 a_n2318_13878.n71 gnd 1.00515f
C871 a_n2318_13878.t41 gnd 0.113752f
C872 a_n2318_13878.t44 gnd 0.113752f
C873 a_n2318_13878.n72 gnd 1.00811f
C874 a_n2318_13878.t43 gnd 0.113752f
C875 a_n2318_13878.t47 gnd 0.113752f
C876 a_n2318_13878.n73 gnd 1.00515f
C877 a_n2318_13878.t78 gnd 0.691694f
C878 a_n2318_13878.t59 gnd 0.680295f
C879 a_n2318_13878.t63 gnd 0.680295f
C880 a_n2318_13878.n74 gnd 0.297177f
C881 a_n2318_13878.t53 gnd 0.680295f
C882 a_n2318_13878.t68 gnd 0.680295f
C883 a_n2318_13878.t75 gnd 0.680295f
C884 a_n2318_13878.n75 gnd 0.297177f
C885 a_n2318_13878.t76 gnd 0.680295f
C886 a_n2318_13878.t50 gnd 0.691694f
C887 a_n2318_13878.t12 gnd 1.36943f
C888 a_n2318_13878.t8 gnd 0.146252f
C889 a_n2318_13878.t14 gnd 0.146252f
C890 a_n2318_13878.n76 gnd 1.0302f
C891 a_n2318_13878.t22 gnd 0.146252f
C892 a_n2318_13878.t34 gnd 0.146252f
C893 a_n2318_13878.n77 gnd 1.0302f
C894 a_n2318_13878.t30 gnd 0.146252f
C895 a_n2318_13878.t20 gnd 0.146252f
C896 a_n2318_13878.n78 gnd 1.0302f
C897 a_n2318_13878.t24 gnd 1.3667f
C898 a_n2318_13878.t29 gnd 0.680295f
C899 a_n2318_13878.n79 gnd 0.297177f
C900 a_n2318_13878.t21 gnd 0.680295f
C901 a_n2318_13878.t11 gnd 0.691694f
C902 a_n2318_13878.t7 gnd 0.680295f
C903 a_n2318_13878.t58 gnd 0.680295f
C904 a_n2318_13878.n80 gnd 0.297177f
C905 a_n2318_13878.t72 gnd 0.680295f
C906 a_n2318_13878.t74 gnd 0.691694f
C907 a_n2318_13878.t52 gnd 0.680295f
C908 a_n2318_13878.n81 gnd 0.2996f
C909 a_n2318_13878.t71 gnd 0.680295f
C910 a_n2318_13878.n82 gnd 0.297177f
C911 a_n2318_13878.n83 gnd 0.292702f
C912 a_n2318_13878.t49 gnd 0.680295f
C913 a_n2318_13878.n84 gnd 0.292702f
C914 a_n2318_13878.t67 gnd 0.680295f
C915 a_n2318_13878.n85 gnd 0.2996f
C916 a_n2318_13878.t51 gnd 0.691694f
C917 a_n2318_13878.n86 gnd 0.2996f
C918 a_n2318_13878.t13 gnd 0.680295f
C919 a_n2318_13878.n87 gnd 0.297177f
C920 a_n2318_13878.n88 gnd 0.292702f
C921 a_n2318_13878.t33 gnd 0.680295f
C922 a_n2318_13878.n89 gnd 0.292702f
C923 a_n2318_13878.t19 gnd 0.680295f
C924 a_n2318_13878.n90 gnd 0.2996f
C925 a_n2318_13878.t23 gnd 0.691694f
C926 a_n2318_13878.n91 gnd 1.17031f
C927 a_n2318_13878.t56 gnd 0.680295f
C928 a_n2318_13878.n92 gnd 0.295302f
C929 a_n2318_13878.t62 gnd 0.680295f
C930 a_n2318_13878.n93 gnd 0.295302f
C931 a_n2318_13878.t54 gnd 0.680295f
C932 a_n2318_13878.n94 gnd 0.295302f
C933 a_n2318_13878.t66 gnd 0.680295f
C934 a_n2318_13878.n95 gnd 0.295302f
C935 a_n2318_13878.t57 gnd 0.680295f
C936 a_n2318_13878.n96 gnd 0.28994f
C937 a_n2318_13878.t79 gnd 0.680295f
C938 a_n2318_13878.n97 gnd 0.299101f
C939 a_n2318_13878.t60 gnd 0.691694f
C940 a_n2318_13878.t69 gnd 0.680295f
C941 a_n2318_13878.n98 gnd 0.28994f
C942 a_n2318_13878.t55 gnd 0.680295f
C943 a_n2318_13878.n99 gnd 0.299101f
C944 a_n2318_13878.t64 gnd 0.691694f
C945 a_n2318_13878.t73 gnd 0.680295f
C946 a_n2318_13878.n100 gnd 0.28994f
C947 a_n2318_13878.t61 gnd 0.680295f
C948 a_n2318_13878.n101 gnd 0.299101f
C949 a_n2318_13878.t77 gnd 0.691694f
C950 a_n2318_13878.t65 gnd 0.680295f
C951 a_n2318_13878.n102 gnd 0.28994f
C952 a_n2318_13878.t48 gnd 0.680295f
C953 a_n2318_13878.n103 gnd 0.299101f
C954 a_n2318_13878.t70 gnd 0.691694f
C955 a_n2318_13878.n104 gnd 1.41607f
C956 a_n2318_13878.n105 gnd 0.2996f
C957 a_n2318_13878.n106 gnd 0.292702f
C958 a_n2318_13878.n107 gnd 0.292702f
C959 a_n2318_13878.n108 gnd 0.2996f
C960 a_n2318_13878.n109 gnd 0.2996f
C961 a_n2318_13878.n110 gnd 0.292702f
C962 a_n2318_13878.n111 gnd 0.292702f
C963 a_n2318_13878.n112 gnd 0.2996f
C964 a_n2318_13878.n113 gnd 0.839379f
C965 a_n2318_13878.t32 gnd 1.36671f
C966 a_n2318_13878.t16 gnd 0.146252f
C967 a_n2318_13878.t18 gnd 0.146252f
C968 a_n2318_13878.n114 gnd 1.0302f
C969 a_n2318_13878.t26 gnd 1.36943f
C970 a_n2318_13878.t10 gnd 0.146252f
C971 a_n2318_13878.t6 gnd 0.146252f
C972 a_n2318_13878.n115 gnd 1.0302f
C973 a_n2318_13878.n116 gnd 1.0302f
C974 a_n2318_13878.t4 gnd 0.146252f
C975 CSoutput.n0 gnd 0.045471f
C976 CSoutput.t195 gnd 0.300781f
C977 CSoutput.n1 gnd 0.135818f
C978 CSoutput.n2 gnd 0.045471f
C979 CSoutput.t199 gnd 0.300781f
C980 CSoutput.n3 gnd 0.03604f
C981 CSoutput.n4 gnd 0.045471f
C982 CSoutput.t211 gnd 0.300781f
C983 CSoutput.n5 gnd 0.031077f
C984 CSoutput.n6 gnd 0.045471f
C985 CSoutput.t197 gnd 0.300781f
C986 CSoutput.t203 gnd 0.300781f
C987 CSoutput.n7 gnd 0.134337f
C988 CSoutput.n8 gnd 0.045471f
C989 CSoutput.t201 gnd 0.300781f
C990 CSoutput.n9 gnd 0.02963f
C991 CSoutput.n10 gnd 0.045471f
C992 CSoutput.t213 gnd 0.300781f
C993 CSoutput.t200 gnd 0.300781f
C994 CSoutput.n11 gnd 0.134337f
C995 CSoutput.n12 gnd 0.045471f
C996 CSoutput.t198 gnd 0.300781f
C997 CSoutput.n13 gnd 0.031077f
C998 CSoutput.n14 gnd 0.045471f
C999 CSoutput.t210 gnd 0.300781f
C1000 CSoutput.t194 gnd 0.300781f
C1001 CSoutput.n15 gnd 0.134337f
C1002 CSoutput.n16 gnd 0.045471f
C1003 CSoutput.t196 gnd 0.300781f
C1004 CSoutput.n17 gnd 0.033192f
C1005 CSoutput.t206 gnd 0.359441f
C1006 CSoutput.t208 gnd 0.300781f
C1007 CSoutput.n18 gnd 0.171497f
C1008 CSoutput.n19 gnd 0.166411f
C1009 CSoutput.n20 gnd 0.193057f
C1010 CSoutput.n21 gnd 0.045471f
C1011 CSoutput.n22 gnd 0.037951f
C1012 CSoutput.n23 gnd 0.134337f
C1013 CSoutput.n24 gnd 0.036583f
C1014 CSoutput.n25 gnd 0.03604f
C1015 CSoutput.n26 gnd 0.045471f
C1016 CSoutput.n27 gnd 0.045471f
C1017 CSoutput.n28 gnd 0.037659f
C1018 CSoutput.n29 gnd 0.031973f
C1019 CSoutput.n30 gnd 0.137328f
C1020 CSoutput.n31 gnd 0.032414f
C1021 CSoutput.n32 gnd 0.045471f
C1022 CSoutput.n33 gnd 0.045471f
C1023 CSoutput.n34 gnd 0.045471f
C1024 CSoutput.n35 gnd 0.037258f
C1025 CSoutput.n36 gnd 0.134337f
C1026 CSoutput.n37 gnd 0.035632f
C1027 CSoutput.n38 gnd 0.036991f
C1028 CSoutput.n39 gnd 0.045471f
C1029 CSoutput.n40 gnd 0.045471f
C1030 CSoutput.n41 gnd 0.037943f
C1031 CSoutput.n42 gnd 0.03468f
C1032 CSoutput.n43 gnd 0.134337f
C1033 CSoutput.n44 gnd 0.035559f
C1034 CSoutput.n45 gnd 0.045471f
C1035 CSoutput.n46 gnd 0.045471f
C1036 CSoutput.n47 gnd 0.045471f
C1037 CSoutput.n48 gnd 0.035559f
C1038 CSoutput.n49 gnd 0.134337f
C1039 CSoutput.n50 gnd 0.03468f
C1040 CSoutput.n51 gnd 0.037943f
C1041 CSoutput.n52 gnd 0.045471f
C1042 CSoutput.n53 gnd 0.045471f
C1043 CSoutput.n54 gnd 0.036991f
C1044 CSoutput.n55 gnd 0.035632f
C1045 CSoutput.n56 gnd 0.134337f
C1046 CSoutput.n57 gnd 0.037258f
C1047 CSoutput.n58 gnd 0.045471f
C1048 CSoutput.n59 gnd 0.045471f
C1049 CSoutput.n60 gnd 0.045471f
C1050 CSoutput.n61 gnd 0.032414f
C1051 CSoutput.n62 gnd 0.137328f
C1052 CSoutput.n63 gnd 0.031973f
C1053 CSoutput.t205 gnd 0.300781f
C1054 CSoutput.n64 gnd 0.134337f
C1055 CSoutput.n65 gnd 0.037659f
C1056 CSoutput.n66 gnd 0.045471f
C1057 CSoutput.n67 gnd 0.045471f
C1058 CSoutput.n68 gnd 0.045471f
C1059 CSoutput.n69 gnd 0.036583f
C1060 CSoutput.n70 gnd 0.134337f
C1061 CSoutput.n71 gnd 0.037951f
C1062 CSoutput.n72 gnd 0.033192f
C1063 CSoutput.n73 gnd 0.045471f
C1064 CSoutput.n74 gnd 0.045471f
C1065 CSoutput.n75 gnd 0.034422f
C1066 CSoutput.n76 gnd 0.020444f
C1067 CSoutput.t207 gnd 0.337949f
C1068 CSoutput.n77 gnd 0.167879f
C1069 CSoutput.n78 gnd 0.686787f
C1070 CSoutput.t78 gnd 0.056719f
C1071 CSoutput.t25 gnd 0.056719f
C1072 CSoutput.n79 gnd 0.439135f
C1073 CSoutput.t90 gnd 0.056719f
C1074 CSoutput.t42 gnd 0.056719f
C1075 CSoutput.n80 gnd 0.438352f
C1076 CSoutput.n81 gnd 0.444927f
C1077 CSoutput.t6 gnd 0.056719f
C1078 CSoutput.t54 gnd 0.056719f
C1079 CSoutput.n82 gnd 0.438352f
C1080 CSoutput.n83 gnd 0.219241f
C1081 CSoutput.t10 gnd 0.056719f
C1082 CSoutput.t34 gnd 0.056719f
C1083 CSoutput.n84 gnd 0.438352f
C1084 CSoutput.n85 gnd 0.219241f
C1085 CSoutput.t94 gnd 0.056719f
C1086 CSoutput.t49 gnd 0.056719f
C1087 CSoutput.n86 gnd 0.438352f
C1088 CSoutput.n87 gnd 0.219241f
C1089 CSoutput.t13 gnd 0.056719f
C1090 CSoutput.t82 gnd 0.056719f
C1091 CSoutput.n88 gnd 0.438352f
C1092 CSoutput.n89 gnd 0.219241f
C1093 CSoutput.t21 gnd 0.056719f
C1094 CSoutput.t64 gnd 0.056719f
C1095 CSoutput.n90 gnd 0.438352f
C1096 CSoutput.n91 gnd 0.219241f
C1097 CSoutput.t37 gnd 0.056719f
C1098 CSoutput.t55 gnd 0.056719f
C1099 CSoutput.n92 gnd 0.438352f
C1100 CSoutput.n93 gnd 0.402038f
C1101 CSoutput.t2 gnd 0.056719f
C1102 CSoutput.t76 gnd 0.056719f
C1103 CSoutput.n94 gnd 0.439135f
C1104 CSoutput.t65 gnd 0.056719f
C1105 CSoutput.t44 gnd 0.056719f
C1106 CSoutput.n95 gnd 0.438352f
C1107 CSoutput.n96 gnd 0.444927f
C1108 CSoutput.t26 gnd 0.056719f
C1109 CSoutput.t87 gnd 0.056719f
C1110 CSoutput.n97 gnd 0.438352f
C1111 CSoutput.n98 gnd 0.219241f
C1112 CSoutput.t62 gnd 0.056719f
C1113 CSoutput.t61 gnd 0.056719f
C1114 CSoutput.n99 gnd 0.438352f
C1115 CSoutput.n100 gnd 0.219241f
C1116 CSoutput.t51 gnd 0.056719f
C1117 CSoutput.t22 gnd 0.056719f
C1118 CSoutput.n101 gnd 0.438352f
C1119 CSoutput.n102 gnd 0.219241f
C1120 CSoutput.t5 gnd 0.056719f
C1121 CSoutput.t52 gnd 0.056719f
C1122 CSoutput.n103 gnd 0.438352f
C1123 CSoutput.n104 gnd 0.219241f
C1124 CSoutput.t50 gnd 0.056719f
C1125 CSoutput.t20 gnd 0.056719f
C1126 CSoutput.n105 gnd 0.438352f
C1127 CSoutput.n106 gnd 0.219241f
C1128 CSoutput.t3 gnd 0.056719f
C1129 CSoutput.t1 gnd 0.056719f
C1130 CSoutput.n107 gnd 0.438352f
C1131 CSoutput.n108 gnd 0.326944f
C1132 CSoutput.n109 gnd 0.412274f
C1133 CSoutput.t15 gnd 0.056719f
C1134 CSoutput.t86 gnd 0.056719f
C1135 CSoutput.n110 gnd 0.439135f
C1136 CSoutput.t71 gnd 0.056719f
C1137 CSoutput.t53 gnd 0.056719f
C1138 CSoutput.n111 gnd 0.438352f
C1139 CSoutput.n112 gnd 0.444927f
C1140 CSoutput.t38 gnd 0.056719f
C1141 CSoutput.t95 gnd 0.056719f
C1142 CSoutput.n113 gnd 0.438352f
C1143 CSoutput.n114 gnd 0.219241f
C1144 CSoutput.t70 gnd 0.056719f
C1145 CSoutput.t69 gnd 0.056719f
C1146 CSoutput.n115 gnd 0.438352f
C1147 CSoutput.n116 gnd 0.219241f
C1148 CSoutput.t59 gnd 0.056719f
C1149 CSoutput.t35 gnd 0.056719f
C1150 CSoutput.n117 gnd 0.438352f
C1151 CSoutput.n118 gnd 0.219241f
C1152 CSoutput.t17 gnd 0.056719f
C1153 CSoutput.t60 gnd 0.056719f
C1154 CSoutput.n119 gnd 0.438352f
C1155 CSoutput.n120 gnd 0.219241f
C1156 CSoutput.t58 gnd 0.056719f
C1157 CSoutput.t33 gnd 0.056719f
C1158 CSoutput.n121 gnd 0.438352f
C1159 CSoutput.n122 gnd 0.219241f
C1160 CSoutput.t16 gnd 0.056719f
C1161 CSoutput.t14 gnd 0.056719f
C1162 CSoutput.n123 gnd 0.438352f
C1163 CSoutput.n124 gnd 0.326944f
C1164 CSoutput.n125 gnd 0.460817f
C1165 CSoutput.n126 gnd 9.030571f
C1166 CSoutput.n128 gnd 0.804375f
C1167 CSoutput.n129 gnd 0.603281f
C1168 CSoutput.n130 gnd 0.804375f
C1169 CSoutput.n131 gnd 0.804375f
C1170 CSoutput.n132 gnd 2.16562f
C1171 CSoutput.n133 gnd 0.804375f
C1172 CSoutput.n134 gnd 0.804375f
C1173 CSoutput.t192 gnd 1.00547f
C1174 CSoutput.n135 gnd 0.804375f
C1175 CSoutput.n136 gnd 0.804375f
C1176 CSoutput.n140 gnd 0.804375f
C1177 CSoutput.n144 gnd 0.804375f
C1178 CSoutput.n145 gnd 0.804375f
C1179 CSoutput.n147 gnd 0.804375f
C1180 CSoutput.n152 gnd 0.804375f
C1181 CSoutput.n154 gnd 0.804375f
C1182 CSoutput.n155 gnd 0.804375f
C1183 CSoutput.n157 gnd 0.804375f
C1184 CSoutput.n158 gnd 0.804375f
C1185 CSoutput.n160 gnd 0.804375f
C1186 CSoutput.t204 gnd 13.441f
C1187 CSoutput.n162 gnd 0.804375f
C1188 CSoutput.n163 gnd 0.603281f
C1189 CSoutput.n164 gnd 0.804375f
C1190 CSoutput.n165 gnd 0.804375f
C1191 CSoutput.n166 gnd 2.16562f
C1192 CSoutput.n167 gnd 0.804375f
C1193 CSoutput.n168 gnd 0.804375f
C1194 CSoutput.t209 gnd 1.00547f
C1195 CSoutput.n169 gnd 0.804375f
C1196 CSoutput.n170 gnd 0.804375f
C1197 CSoutput.n174 gnd 0.804375f
C1198 CSoutput.n178 gnd 0.804375f
C1199 CSoutput.n179 gnd 0.804375f
C1200 CSoutput.n181 gnd 0.804375f
C1201 CSoutput.n186 gnd 0.804375f
C1202 CSoutput.n188 gnd 0.804375f
C1203 CSoutput.n189 gnd 0.804375f
C1204 CSoutput.n191 gnd 0.804375f
C1205 CSoutput.n192 gnd 0.804375f
C1206 CSoutput.n194 gnd 0.804375f
C1207 CSoutput.n195 gnd 0.603281f
C1208 CSoutput.n197 gnd 0.804375f
C1209 CSoutput.n198 gnd 0.603281f
C1210 CSoutput.n199 gnd 0.804375f
C1211 CSoutput.n200 gnd 0.804375f
C1212 CSoutput.n201 gnd 2.16562f
C1213 CSoutput.n202 gnd 0.804375f
C1214 CSoutput.n203 gnd 0.804375f
C1215 CSoutput.t202 gnd 1.00547f
C1216 CSoutput.n204 gnd 0.804375f
C1217 CSoutput.n205 gnd 2.16562f
C1218 CSoutput.n207 gnd 0.804375f
C1219 CSoutput.n208 gnd 0.804375f
C1220 CSoutput.n210 gnd 0.804375f
C1221 CSoutput.n211 gnd 0.804375f
C1222 CSoutput.t212 gnd 13.222f
C1223 CSoutput.t193 gnd 13.441f
C1224 CSoutput.n217 gnd 2.52344f
C1225 CSoutput.n218 gnd 10.279599f
C1226 CSoutput.n219 gnd 10.7097f
C1227 CSoutput.n224 gnd 2.73357f
C1228 CSoutput.n230 gnd 0.804375f
C1229 CSoutput.n232 gnd 0.804375f
C1230 CSoutput.n234 gnd 0.804375f
C1231 CSoutput.n236 gnd 0.804375f
C1232 CSoutput.n238 gnd 0.804375f
C1233 CSoutput.n244 gnd 0.804375f
C1234 CSoutput.n251 gnd 1.47572f
C1235 CSoutput.n252 gnd 1.47572f
C1236 CSoutput.n253 gnd 0.804375f
C1237 CSoutput.n254 gnd 0.804375f
C1238 CSoutput.n256 gnd 0.603281f
C1239 CSoutput.n257 gnd 0.516656f
C1240 CSoutput.n259 gnd 0.603281f
C1241 CSoutput.n260 gnd 0.516656f
C1242 CSoutput.n261 gnd 0.603281f
C1243 CSoutput.n263 gnd 0.804375f
C1244 CSoutput.n265 gnd 2.16562f
C1245 CSoutput.n266 gnd 2.52344f
C1246 CSoutput.n267 gnd 9.45457f
C1247 CSoutput.n269 gnd 0.603281f
C1248 CSoutput.n270 gnd 1.55228f
C1249 CSoutput.n271 gnd 0.603281f
C1250 CSoutput.n273 gnd 0.804375f
C1251 CSoutput.n275 gnd 2.16562f
C1252 CSoutput.n276 gnd 4.71708f
C1253 CSoutput.t24 gnd 0.056719f
C1254 CSoutput.t77 gnd 0.056719f
C1255 CSoutput.n277 gnd 0.439135f
C1256 CSoutput.t41 gnd 0.056719f
C1257 CSoutput.t89 gnd 0.056719f
C1258 CSoutput.n278 gnd 0.438352f
C1259 CSoutput.n279 gnd 0.444927f
C1260 CSoutput.t72 gnd 0.056719f
C1261 CSoutput.t4 gnd 0.056719f
C1262 CSoutput.n280 gnd 0.438352f
C1263 CSoutput.n281 gnd 0.219241f
C1264 CSoutput.t32 gnd 0.056719f
C1265 CSoutput.t9 gnd 0.056719f
C1266 CSoutput.n282 gnd 0.438352f
C1267 CSoutput.n283 gnd 0.219241f
C1268 CSoutput.t48 gnd 0.056719f
C1269 CSoutput.t29 gnd 0.056719f
C1270 CSoutput.n284 gnd 0.438352f
C1271 CSoutput.n285 gnd 0.219241f
C1272 CSoutput.t81 gnd 0.056719f
C1273 CSoutput.t12 gnd 0.056719f
C1274 CSoutput.n286 gnd 0.438352f
C1275 CSoutput.n287 gnd 0.219241f
C1276 CSoutput.t63 gnd 0.056719f
C1277 CSoutput.t18 gnd 0.056719f
C1278 CSoutput.n288 gnd 0.438352f
C1279 CSoutput.n289 gnd 0.219241f
C1280 CSoutput.t73 gnd 0.056719f
C1281 CSoutput.t36 gnd 0.056719f
C1282 CSoutput.n290 gnd 0.438352f
C1283 CSoutput.n291 gnd 0.402038f
C1284 CSoutput.t47 gnd 0.056719f
C1285 CSoutput.t67 gnd 0.056719f
C1286 CSoutput.n292 gnd 0.439135f
C1287 CSoutput.t0 gnd 0.056719f
C1288 CSoutput.t30 gnd 0.056719f
C1289 CSoutput.n293 gnd 0.438352f
C1290 CSoutput.n294 gnd 0.444927f
C1291 CSoutput.t31 gnd 0.056719f
C1292 CSoutput.t85 gnd 0.056719f
C1293 CSoutput.n295 gnd 0.438352f
C1294 CSoutput.n296 gnd 0.219241f
C1295 CSoutput.t27 gnd 0.056719f
C1296 CSoutput.t28 gnd 0.056719f
C1297 CSoutput.n297 gnd 0.438352f
C1298 CSoutput.n298 gnd 0.219241f
C1299 CSoutput.t83 gnd 0.056719f
C1300 CSoutput.t84 gnd 0.056719f
C1301 CSoutput.n299 gnd 0.438352f
C1302 CSoutput.n300 gnd 0.219241f
C1303 CSoutput.t8 gnd 0.056719f
C1304 CSoutput.t68 gnd 0.056719f
C1305 CSoutput.n301 gnd 0.438352f
C1306 CSoutput.n302 gnd 0.219241f
C1307 CSoutput.t80 gnd 0.056719f
C1308 CSoutput.t7 gnd 0.056719f
C1309 CSoutput.n303 gnd 0.438352f
C1310 CSoutput.n304 gnd 0.219241f
C1311 CSoutput.t46 gnd 0.056719f
C1312 CSoutput.t66 gnd 0.056719f
C1313 CSoutput.n305 gnd 0.438352f
C1314 CSoutput.n306 gnd 0.326944f
C1315 CSoutput.n307 gnd 0.412274f
C1316 CSoutput.t56 gnd 0.056719f
C1317 CSoutput.t74 gnd 0.056719f
C1318 CSoutput.n308 gnd 0.439135f
C1319 CSoutput.t11 gnd 0.056719f
C1320 CSoutput.t43 gnd 0.056719f
C1321 CSoutput.n309 gnd 0.438352f
C1322 CSoutput.n310 gnd 0.444927f
C1323 CSoutput.t45 gnd 0.056719f
C1324 CSoutput.t93 gnd 0.056719f
C1325 CSoutput.n311 gnd 0.438352f
C1326 CSoutput.n312 gnd 0.219241f
C1327 CSoutput.t39 gnd 0.056719f
C1328 CSoutput.t40 gnd 0.056719f
C1329 CSoutput.n313 gnd 0.438352f
C1330 CSoutput.n314 gnd 0.219241f
C1331 CSoutput.t91 gnd 0.056719f
C1332 CSoutput.t92 gnd 0.056719f
C1333 CSoutput.n315 gnd 0.438352f
C1334 CSoutput.n316 gnd 0.219241f
C1335 CSoutput.t23 gnd 0.056719f
C1336 CSoutput.t79 gnd 0.056719f
C1337 CSoutput.n317 gnd 0.438352f
C1338 CSoutput.n318 gnd 0.219241f
C1339 CSoutput.t88 gnd 0.056719f
C1340 CSoutput.t19 gnd 0.056719f
C1341 CSoutput.n319 gnd 0.438352f
C1342 CSoutput.n320 gnd 0.219241f
C1343 CSoutput.t57 gnd 0.056719f
C1344 CSoutput.t75 gnd 0.056719f
C1345 CSoutput.n321 gnd 0.438351f
C1346 CSoutput.n322 gnd 0.326945f
C1347 CSoutput.n323 gnd 0.460817f
C1348 CSoutput.n324 gnd 12.6621f
C1349 CSoutput.t177 gnd 0.049629f
C1350 CSoutput.t109 gnd 0.049629f
C1351 CSoutput.n325 gnd 0.440006f
C1352 CSoutput.t159 gnd 0.049629f
C1353 CSoutput.t98 gnd 0.049629f
C1354 CSoutput.n326 gnd 0.438538f
C1355 CSoutput.n327 gnd 0.408636f
C1356 CSoutput.t143 gnd 0.049629f
C1357 CSoutput.t180 gnd 0.049629f
C1358 CSoutput.n328 gnd 0.438538f
C1359 CSoutput.n329 gnd 0.201438f
C1360 CSoutput.t131 gnd 0.049629f
C1361 CSoutput.t142 gnd 0.049629f
C1362 CSoutput.n330 gnd 0.438538f
C1363 CSoutput.n331 gnd 0.201438f
C1364 CSoutput.t101 gnd 0.049629f
C1365 CSoutput.t149 gnd 0.049629f
C1366 CSoutput.n332 gnd 0.438538f
C1367 CSoutput.n333 gnd 0.201438f
C1368 CSoutput.t163 gnd 0.049629f
C1369 CSoutput.t132 gnd 0.049629f
C1370 CSoutput.n334 gnd 0.438538f
C1371 CSoutput.n335 gnd 0.201438f
C1372 CSoutput.t145 gnd 0.049629f
C1373 CSoutput.t173 gnd 0.049629f
C1374 CSoutput.n336 gnd 0.438538f
C1375 CSoutput.n337 gnd 0.201438f
C1376 CSoutput.t108 gnd 0.049629f
C1377 CSoutput.t123 gnd 0.049629f
C1378 CSoutput.n338 gnd 0.438538f
C1379 CSoutput.n339 gnd 0.371542f
C1380 CSoutput.t140 gnd 0.049629f
C1381 CSoutput.t117 gnd 0.049629f
C1382 CSoutput.n340 gnd 0.440006f
C1383 CSoutput.t127 gnd 0.049629f
C1384 CSoutput.t139 gnd 0.049629f
C1385 CSoutput.n341 gnd 0.438538f
C1386 CSoutput.n342 gnd 0.408636f
C1387 CSoutput.t116 gnd 0.049629f
C1388 CSoutput.t129 gnd 0.049629f
C1389 CSoutput.n343 gnd 0.438538f
C1390 CSoutput.n344 gnd 0.201438f
C1391 CSoutput.t141 gnd 0.049629f
C1392 CSoutput.t115 gnd 0.049629f
C1393 CSoutput.n345 gnd 0.438538f
C1394 CSoutput.n346 gnd 0.201438f
C1395 CSoutput.t128 gnd 0.049629f
C1396 CSoutput.t106 gnd 0.049629f
C1397 CSoutput.n347 gnd 0.438538f
C1398 CSoutput.n348 gnd 0.201438f
C1399 CSoutput.t114 gnd 0.049629f
C1400 CSoutput.t130 gnd 0.049629f
C1401 CSoutput.n349 gnd 0.438538f
C1402 CSoutput.n350 gnd 0.201438f
C1403 CSoutput.t103 gnd 0.049629f
C1404 CSoutput.t186 gnd 0.049629f
C1405 CSoutput.n351 gnd 0.438538f
C1406 CSoutput.n352 gnd 0.201438f
C1407 CSoutput.t120 gnd 0.049629f
C1408 CSoutput.t191 gnd 0.049629f
C1409 CSoutput.n353 gnd 0.438538f
C1410 CSoutput.n354 gnd 0.305826f
C1411 CSoutput.n355 gnd 0.385742f
C1412 CSoutput.t107 gnd 0.049629f
C1413 CSoutput.t187 gnd 0.049629f
C1414 CSoutput.n356 gnd 0.440006f
C1415 CSoutput.t175 gnd 0.049629f
C1416 CSoutput.t121 gnd 0.049629f
C1417 CSoutput.n357 gnd 0.438538f
C1418 CSoutput.n358 gnd 0.408636f
C1419 CSoutput.t96 gnd 0.049629f
C1420 CSoutput.t181 gnd 0.049629f
C1421 CSoutput.n359 gnd 0.438538f
C1422 CSoutput.n360 gnd 0.201438f
C1423 CSoutput.t135 gnd 0.049629f
C1424 CSoutput.t144 gnd 0.049629f
C1425 CSoutput.n361 gnd 0.438538f
C1426 CSoutput.n362 gnd 0.201438f
C1427 CSoutput.t188 gnd 0.049629f
C1428 CSoutput.t174 gnd 0.049629f
C1429 CSoutput.n363 gnd 0.438538f
C1430 CSoutput.n364 gnd 0.201438f
C1431 CSoutput.t154 gnd 0.049629f
C1432 CSoutput.t97 gnd 0.049629f
C1433 CSoutput.n365 gnd 0.438538f
C1434 CSoutput.n366 gnd 0.201438f
C1435 CSoutput.t105 gnd 0.049629f
C1436 CSoutput.t185 gnd 0.049629f
C1437 CSoutput.n367 gnd 0.438538f
C1438 CSoutput.n368 gnd 0.201438f
C1439 CSoutput.t112 gnd 0.049629f
C1440 CSoutput.t119 gnd 0.049629f
C1441 CSoutput.n369 gnd 0.438538f
C1442 CSoutput.n370 gnd 0.305826f
C1443 CSoutput.n371 gnd 0.414226f
C1444 CSoutput.n372 gnd 13.216401f
C1445 CSoutput.t151 gnd 0.049629f
C1446 CSoutput.t102 gnd 0.049629f
C1447 CSoutput.n373 gnd 0.440006f
C1448 CSoutput.t134 gnd 0.049629f
C1449 CSoutput.t182 gnd 0.049629f
C1450 CSoutput.n374 gnd 0.438538f
C1451 CSoutput.n375 gnd 0.408636f
C1452 CSoutput.t104 gnd 0.049629f
C1453 CSoutput.t165 gnd 0.049629f
C1454 CSoutput.n376 gnd 0.438538f
C1455 CSoutput.n377 gnd 0.201438f
C1456 CSoutput.t164 gnd 0.049629f
C1457 CSoutput.t153 gnd 0.049629f
C1458 CSoutput.n378 gnd 0.438538f
C1459 CSoutput.n379 gnd 0.201438f
C1460 CSoutput.t168 gnd 0.049629f
C1461 CSoutput.t136 gnd 0.049629f
C1462 CSoutput.n380 gnd 0.438538f
C1463 CSoutput.n381 gnd 0.201438f
C1464 CSoutput.t160 gnd 0.049629f
C1465 CSoutput.t176 gnd 0.049629f
C1466 CSoutput.n382 gnd 0.438538f
C1467 CSoutput.n383 gnd 0.201438f
C1468 CSoutput.t190 gnd 0.049629f
C1469 CSoutput.t167 gnd 0.049629f
C1470 CSoutput.n384 gnd 0.438538f
C1471 CSoutput.n385 gnd 0.201438f
C1472 CSoutput.t172 gnd 0.049629f
C1473 CSoutput.t171 gnd 0.049629f
C1474 CSoutput.n386 gnd 0.438538f
C1475 CSoutput.n387 gnd 0.371542f
C1476 CSoutput.t137 gnd 0.049629f
C1477 CSoutput.t155 gnd 0.049629f
C1478 CSoutput.n388 gnd 0.440006f
C1479 CSoutput.t156 gnd 0.049629f
C1480 CSoutput.t146 gnd 0.049629f
C1481 CSoutput.n389 gnd 0.438538f
C1482 CSoutput.n390 gnd 0.408636f
C1483 CSoutput.t147 gnd 0.049629f
C1484 CSoutput.t138 gnd 0.049629f
C1485 CSoutput.n391 gnd 0.438538f
C1486 CSoutput.n392 gnd 0.201438f
C1487 CSoutput.t133 gnd 0.049629f
C1488 CSoutput.t125 gnd 0.049629f
C1489 CSoutput.n393 gnd 0.438538f
C1490 CSoutput.n394 gnd 0.201438f
C1491 CSoutput.t126 gnd 0.049629f
C1492 CSoutput.t148 gnd 0.049629f
C1493 CSoutput.n395 gnd 0.438538f
C1494 CSoutput.n396 gnd 0.201438f
C1495 CSoutput.t150 gnd 0.049629f
C1496 CSoutput.t99 gnd 0.049629f
C1497 CSoutput.n397 gnd 0.438538f
C1498 CSoutput.n398 gnd 0.201438f
C1499 CSoutput.t100 gnd 0.049629f
C1500 CSoutput.t118 gnd 0.049629f
C1501 CSoutput.n399 gnd 0.438538f
C1502 CSoutput.n400 gnd 0.201438f
C1503 CSoutput.t124 gnd 0.049629f
C1504 CSoutput.t113 gnd 0.049629f
C1505 CSoutput.n401 gnd 0.438538f
C1506 CSoutput.n402 gnd 0.305826f
C1507 CSoutput.n403 gnd 0.385742f
C1508 CSoutput.t169 gnd 0.049629f
C1509 CSoutput.t184 gnd 0.049629f
C1510 CSoutput.n404 gnd 0.440006f
C1511 CSoutput.t189 gnd 0.049629f
C1512 CSoutput.t158 gnd 0.049629f
C1513 CSoutput.n405 gnd 0.438538f
C1514 CSoutput.n406 gnd 0.408636f
C1515 CSoutput.t162 gnd 0.049629f
C1516 CSoutput.t178 gnd 0.049629f
C1517 CSoutput.n407 gnd 0.438538f
C1518 CSoutput.n408 gnd 0.201438f
C1519 CSoutput.t110 gnd 0.049629f
C1520 CSoutput.t152 gnd 0.049629f
C1521 CSoutput.n409 gnd 0.438538f
C1522 CSoutput.n410 gnd 0.201438f
C1523 CSoutput.t157 gnd 0.049629f
C1524 CSoutput.t170 gnd 0.049629f
C1525 CSoutput.n411 gnd 0.438538f
C1526 CSoutput.n412 gnd 0.201438f
C1527 CSoutput.t179 gnd 0.049629f
C1528 CSoutput.t161 gnd 0.049629f
C1529 CSoutput.n413 gnd 0.438538f
C1530 CSoutput.n414 gnd 0.201438f
C1531 CSoutput.t166 gnd 0.049629f
C1532 CSoutput.t183 gnd 0.049629f
C1533 CSoutput.n415 gnd 0.438538f
C1534 CSoutput.n416 gnd 0.201438f
C1535 CSoutput.t111 gnd 0.049629f
C1536 CSoutput.t122 gnd 0.049629f
C1537 CSoutput.n417 gnd 0.438538f
C1538 CSoutput.n418 gnd 0.305826f
C1539 CSoutput.n419 gnd 0.414226f
C1540 CSoutput.n420 gnd 7.822569f
C1541 CSoutput.n421 gnd 13.8894f
C1542 vdd.t12 gnd 0.037171f
C1543 vdd.t130 gnd 0.037171f
C1544 vdd.n0 gnd 0.293176f
C1545 vdd.t33 gnd 0.037171f
C1546 vdd.t46 gnd 0.037171f
C1547 vdd.n1 gnd 0.292692f
C1548 vdd.n2 gnd 0.269918f
C1549 vdd.t128 gnd 0.037171f
C1550 vdd.t18 gnd 0.037171f
C1551 vdd.n3 gnd 0.292692f
C1552 vdd.n4 gnd 0.136508f
C1553 vdd.t20 gnd 0.037171f
C1554 vdd.t133 gnd 0.037171f
C1555 vdd.n5 gnd 0.292692f
C1556 vdd.n6 gnd 0.128087f
C1557 vdd.t16 gnd 0.037171f
C1558 vdd.t265 gnd 0.037171f
C1559 vdd.n7 gnd 0.293176f
C1560 vdd.t135 gnd 0.037171f
C1561 vdd.t10 gnd 0.037171f
C1562 vdd.n8 gnd 0.292692f
C1563 vdd.n9 gnd 0.269918f
C1564 vdd.t48 gnd 0.037171f
C1565 vdd.t43 gnd 0.037171f
C1566 vdd.n10 gnd 0.292692f
C1567 vdd.n11 gnd 0.136508f
C1568 vdd.t267 gnd 0.037171f
C1569 vdd.t39 gnd 0.037171f
C1570 vdd.n12 gnd 0.292692f
C1571 vdd.n13 gnd 0.128087f
C1572 vdd.n14 gnd 0.090555f
C1573 vdd.t3 gnd 0.020651f
C1574 vdd.t30 gnd 0.020651f
C1575 vdd.n15 gnd 0.190081f
C1576 vdd.t1 gnd 0.020651f
C1577 vdd.t28 gnd 0.020651f
C1578 vdd.n16 gnd 0.189525f
C1579 vdd.n17 gnd 0.329833f
C1580 vdd.t26 gnd 0.020651f
C1581 vdd.t25 gnd 0.020651f
C1582 vdd.n18 gnd 0.189525f
C1583 vdd.n19 gnd 0.136456f
C1584 vdd.t29 gnd 0.020651f
C1585 vdd.t31 gnd 0.020651f
C1586 vdd.n20 gnd 0.190081f
C1587 vdd.t4 gnd 0.020651f
C1588 vdd.t2 gnd 0.020651f
C1589 vdd.n21 gnd 0.189525f
C1590 vdd.n22 gnd 0.329833f
C1591 vdd.t24 gnd 0.020651f
C1592 vdd.t27 gnd 0.020651f
C1593 vdd.n23 gnd 0.189525f
C1594 vdd.n24 gnd 0.136456f
C1595 vdd.t6 gnd 0.020651f
C1596 vdd.t23 gnd 0.020651f
C1597 vdd.n25 gnd 0.189525f
C1598 vdd.t7 gnd 0.020651f
C1599 vdd.t0 gnd 0.020651f
C1600 vdd.n26 gnd 0.189525f
C1601 vdd.n27 gnd 20.9766f
C1602 vdd.n28 gnd 8.16153f
C1603 vdd.n29 gnd 0.005632f
C1604 vdd.n30 gnd 0.005227f
C1605 vdd.n31 gnd 0.002891f
C1606 vdd.n32 gnd 0.006638f
C1607 vdd.n33 gnd 0.002809f
C1608 vdd.n34 gnd 0.002974f
C1609 vdd.n35 gnd 0.005227f
C1610 vdd.n36 gnd 0.002809f
C1611 vdd.n37 gnd 0.006638f
C1612 vdd.n38 gnd 0.002974f
C1613 vdd.n39 gnd 0.005227f
C1614 vdd.n40 gnd 0.002809f
C1615 vdd.n41 gnd 0.004979f
C1616 vdd.n42 gnd 0.004994f
C1617 vdd.t178 gnd 0.014262f
C1618 vdd.n43 gnd 0.031732f
C1619 vdd.n44 gnd 0.165142f
C1620 vdd.n45 gnd 0.002809f
C1621 vdd.n46 gnd 0.002974f
C1622 vdd.n47 gnd 0.006638f
C1623 vdd.n48 gnd 0.006638f
C1624 vdd.n49 gnd 0.002974f
C1625 vdd.n50 gnd 0.002809f
C1626 vdd.n51 gnd 0.005227f
C1627 vdd.n52 gnd 0.005227f
C1628 vdd.n53 gnd 0.002809f
C1629 vdd.n54 gnd 0.002974f
C1630 vdd.n55 gnd 0.006638f
C1631 vdd.n56 gnd 0.006638f
C1632 vdd.n57 gnd 0.002974f
C1633 vdd.n58 gnd 0.002809f
C1634 vdd.n59 gnd 0.005227f
C1635 vdd.n60 gnd 0.005227f
C1636 vdd.n61 gnd 0.002809f
C1637 vdd.n62 gnd 0.002974f
C1638 vdd.n63 gnd 0.006638f
C1639 vdd.n64 gnd 0.006638f
C1640 vdd.n65 gnd 0.015694f
C1641 vdd.n66 gnd 0.002891f
C1642 vdd.n67 gnd 0.002809f
C1643 vdd.n68 gnd 0.013509f
C1644 vdd.n69 gnd 0.009431f
C1645 vdd.t245 gnd 0.033041f
C1646 vdd.t202 gnd 0.033041f
C1647 vdd.n70 gnd 0.227082f
C1648 vdd.n71 gnd 0.178565f
C1649 vdd.t257 gnd 0.033041f
C1650 vdd.t240 gnd 0.033041f
C1651 vdd.n72 gnd 0.227082f
C1652 vdd.n73 gnd 0.144101f
C1653 vdd.t145 gnd 0.033041f
C1654 vdd.t189 gnd 0.033041f
C1655 vdd.n74 gnd 0.227082f
C1656 vdd.n75 gnd 0.144101f
C1657 vdd.t155 gnd 0.033041f
C1658 vdd.t205 gnd 0.033041f
C1659 vdd.n76 gnd 0.227082f
C1660 vdd.n77 gnd 0.144101f
C1661 vdd.t184 gnd 0.033041f
C1662 vdd.t249 gnd 0.033041f
C1663 vdd.n78 gnd 0.227082f
C1664 vdd.n79 gnd 0.144101f
C1665 vdd.t160 gnd 0.033041f
C1666 vdd.t229 gnd 0.033041f
C1667 vdd.n80 gnd 0.227082f
C1668 vdd.n81 gnd 0.144101f
C1669 vdd.t164 gnd 0.033041f
C1670 vdd.t241 gnd 0.033041f
C1671 vdd.n82 gnd 0.227082f
C1672 vdd.n83 gnd 0.144101f
C1673 vdd.n84 gnd 0.005632f
C1674 vdd.n85 gnd 0.005227f
C1675 vdd.n86 gnd 0.002891f
C1676 vdd.n87 gnd 0.006638f
C1677 vdd.n88 gnd 0.002809f
C1678 vdd.n89 gnd 0.002974f
C1679 vdd.n90 gnd 0.005227f
C1680 vdd.n91 gnd 0.002809f
C1681 vdd.n92 gnd 0.006638f
C1682 vdd.n93 gnd 0.002974f
C1683 vdd.n94 gnd 0.005227f
C1684 vdd.n95 gnd 0.002809f
C1685 vdd.n96 gnd 0.004979f
C1686 vdd.n97 gnd 0.004994f
C1687 vdd.t195 gnd 0.014262f
C1688 vdd.n98 gnd 0.031732f
C1689 vdd.n99 gnd 0.165142f
C1690 vdd.n100 gnd 0.002809f
C1691 vdd.n101 gnd 0.002974f
C1692 vdd.n102 gnd 0.006638f
C1693 vdd.n103 gnd 0.006638f
C1694 vdd.n104 gnd 0.002974f
C1695 vdd.n105 gnd 0.002809f
C1696 vdd.n106 gnd 0.005227f
C1697 vdd.n107 gnd 0.005227f
C1698 vdd.n108 gnd 0.002809f
C1699 vdd.n109 gnd 0.002974f
C1700 vdd.n110 gnd 0.006638f
C1701 vdd.n111 gnd 0.006638f
C1702 vdd.n112 gnd 0.002974f
C1703 vdd.n113 gnd 0.002809f
C1704 vdd.n114 gnd 0.005227f
C1705 vdd.n115 gnd 0.005227f
C1706 vdd.n116 gnd 0.002809f
C1707 vdd.n117 gnd 0.002974f
C1708 vdd.n118 gnd 0.006638f
C1709 vdd.n119 gnd 0.006638f
C1710 vdd.n120 gnd 0.015694f
C1711 vdd.n121 gnd 0.002891f
C1712 vdd.n122 gnd 0.002809f
C1713 vdd.n123 gnd 0.013509f
C1714 vdd.n124 gnd 0.009135f
C1715 vdd.n125 gnd 0.107212f
C1716 vdd.n126 gnd 0.005632f
C1717 vdd.n127 gnd 0.005227f
C1718 vdd.n128 gnd 0.002891f
C1719 vdd.n129 gnd 0.006638f
C1720 vdd.n130 gnd 0.002809f
C1721 vdd.n131 gnd 0.002974f
C1722 vdd.n132 gnd 0.005227f
C1723 vdd.n133 gnd 0.002809f
C1724 vdd.n134 gnd 0.006638f
C1725 vdd.n135 gnd 0.002974f
C1726 vdd.n136 gnd 0.005227f
C1727 vdd.n137 gnd 0.002809f
C1728 vdd.n138 gnd 0.004979f
C1729 vdd.n139 gnd 0.004994f
C1730 vdd.t210 gnd 0.014262f
C1731 vdd.n140 gnd 0.031732f
C1732 vdd.n141 gnd 0.165142f
C1733 vdd.n142 gnd 0.002809f
C1734 vdd.n143 gnd 0.002974f
C1735 vdd.n144 gnd 0.006638f
C1736 vdd.n145 gnd 0.006638f
C1737 vdd.n146 gnd 0.002974f
C1738 vdd.n147 gnd 0.002809f
C1739 vdd.n148 gnd 0.005227f
C1740 vdd.n149 gnd 0.005227f
C1741 vdd.n150 gnd 0.002809f
C1742 vdd.n151 gnd 0.002974f
C1743 vdd.n152 gnd 0.006638f
C1744 vdd.n153 gnd 0.006638f
C1745 vdd.n154 gnd 0.002974f
C1746 vdd.n155 gnd 0.002809f
C1747 vdd.n156 gnd 0.005227f
C1748 vdd.n157 gnd 0.005227f
C1749 vdd.n158 gnd 0.002809f
C1750 vdd.n159 gnd 0.002974f
C1751 vdd.n160 gnd 0.006638f
C1752 vdd.n161 gnd 0.006638f
C1753 vdd.n162 gnd 0.015694f
C1754 vdd.n163 gnd 0.002891f
C1755 vdd.n164 gnd 0.002809f
C1756 vdd.n165 gnd 0.013509f
C1757 vdd.n166 gnd 0.009431f
C1758 vdd.t235 gnd 0.033041f
C1759 vdd.t137 gnd 0.033041f
C1760 vdd.n167 gnd 0.227082f
C1761 vdd.n168 gnd 0.178565f
C1762 vdd.t186 gnd 0.033041f
C1763 vdd.t188 gnd 0.033041f
C1764 vdd.n169 gnd 0.227082f
C1765 vdd.n170 gnd 0.144101f
C1766 vdd.t253 gnd 0.033041f
C1767 vdd.t181 gnd 0.033041f
C1768 vdd.n171 gnd 0.227082f
C1769 vdd.n172 gnd 0.144101f
C1770 vdd.t182 gnd 0.033041f
C1771 vdd.t251 gnd 0.033041f
C1772 vdd.n173 gnd 0.227082f
C1773 vdd.n174 gnd 0.144101f
C1774 vdd.t252 gnd 0.033041f
C1775 vdd.t153 gnd 0.033041f
C1776 vdd.n175 gnd 0.227082f
C1777 vdd.n176 gnd 0.144101f
C1778 vdd.t236 gnd 0.033041f
C1779 vdd.t244 gnd 0.033041f
C1780 vdd.n177 gnd 0.227082f
C1781 vdd.n178 gnd 0.144101f
C1782 vdd.t151 gnd 0.033041f
C1783 vdd.t207 gnd 0.033041f
C1784 vdd.n179 gnd 0.227082f
C1785 vdd.n180 gnd 0.144101f
C1786 vdd.n181 gnd 0.005632f
C1787 vdd.n182 gnd 0.005227f
C1788 vdd.n183 gnd 0.002891f
C1789 vdd.n184 gnd 0.006638f
C1790 vdd.n185 gnd 0.002809f
C1791 vdd.n186 gnd 0.002974f
C1792 vdd.n187 gnd 0.005227f
C1793 vdd.n188 gnd 0.002809f
C1794 vdd.n189 gnd 0.006638f
C1795 vdd.n190 gnd 0.002974f
C1796 vdd.n191 gnd 0.005227f
C1797 vdd.n192 gnd 0.002809f
C1798 vdd.n193 gnd 0.004979f
C1799 vdd.n194 gnd 0.004994f
C1800 vdd.t233 gnd 0.014262f
C1801 vdd.n195 gnd 0.031732f
C1802 vdd.n196 gnd 0.165142f
C1803 vdd.n197 gnd 0.002809f
C1804 vdd.n198 gnd 0.002974f
C1805 vdd.n199 gnd 0.006638f
C1806 vdd.n200 gnd 0.006638f
C1807 vdd.n201 gnd 0.002974f
C1808 vdd.n202 gnd 0.002809f
C1809 vdd.n203 gnd 0.005227f
C1810 vdd.n204 gnd 0.005227f
C1811 vdd.n205 gnd 0.002809f
C1812 vdd.n206 gnd 0.002974f
C1813 vdd.n207 gnd 0.006638f
C1814 vdd.n208 gnd 0.006638f
C1815 vdd.n209 gnd 0.002974f
C1816 vdd.n210 gnd 0.002809f
C1817 vdd.n211 gnd 0.005227f
C1818 vdd.n212 gnd 0.005227f
C1819 vdd.n213 gnd 0.002809f
C1820 vdd.n214 gnd 0.002974f
C1821 vdd.n215 gnd 0.006638f
C1822 vdd.n216 gnd 0.006638f
C1823 vdd.n217 gnd 0.015694f
C1824 vdd.n218 gnd 0.002891f
C1825 vdd.n219 gnd 0.002809f
C1826 vdd.n220 gnd 0.013509f
C1827 vdd.n221 gnd 0.009135f
C1828 vdd.n222 gnd 0.06378f
C1829 vdd.n223 gnd 0.229817f
C1830 vdd.n224 gnd 0.005632f
C1831 vdd.n225 gnd 0.005227f
C1832 vdd.n226 gnd 0.002891f
C1833 vdd.n227 gnd 0.006638f
C1834 vdd.n228 gnd 0.002809f
C1835 vdd.n229 gnd 0.002974f
C1836 vdd.n230 gnd 0.005227f
C1837 vdd.n231 gnd 0.002809f
C1838 vdd.n232 gnd 0.006638f
C1839 vdd.n233 gnd 0.002974f
C1840 vdd.n234 gnd 0.005227f
C1841 vdd.n235 gnd 0.002809f
C1842 vdd.n236 gnd 0.004979f
C1843 vdd.n237 gnd 0.004994f
C1844 vdd.t220 gnd 0.014262f
C1845 vdd.n238 gnd 0.031732f
C1846 vdd.n239 gnd 0.165142f
C1847 vdd.n240 gnd 0.002809f
C1848 vdd.n241 gnd 0.002974f
C1849 vdd.n242 gnd 0.006638f
C1850 vdd.n243 gnd 0.006638f
C1851 vdd.n244 gnd 0.002974f
C1852 vdd.n245 gnd 0.002809f
C1853 vdd.n246 gnd 0.005227f
C1854 vdd.n247 gnd 0.005227f
C1855 vdd.n248 gnd 0.002809f
C1856 vdd.n249 gnd 0.002974f
C1857 vdd.n250 gnd 0.006638f
C1858 vdd.n251 gnd 0.006638f
C1859 vdd.n252 gnd 0.002974f
C1860 vdd.n253 gnd 0.002809f
C1861 vdd.n254 gnd 0.005227f
C1862 vdd.n255 gnd 0.005227f
C1863 vdd.n256 gnd 0.002809f
C1864 vdd.n257 gnd 0.002974f
C1865 vdd.n258 gnd 0.006638f
C1866 vdd.n259 gnd 0.006638f
C1867 vdd.n260 gnd 0.015694f
C1868 vdd.n261 gnd 0.002891f
C1869 vdd.n262 gnd 0.002809f
C1870 vdd.n263 gnd 0.013509f
C1871 vdd.n264 gnd 0.009431f
C1872 vdd.t242 gnd 0.033041f
C1873 vdd.t158 gnd 0.033041f
C1874 vdd.n265 gnd 0.227082f
C1875 vdd.n266 gnd 0.178565f
C1876 vdd.t203 gnd 0.033041f
C1877 vdd.t209 gnd 0.033041f
C1878 vdd.n267 gnd 0.227082f
C1879 vdd.n268 gnd 0.144101f
C1880 vdd.t261 gnd 0.033041f
C1881 vdd.t198 gnd 0.033041f
C1882 vdd.n269 gnd 0.227082f
C1883 vdd.n270 gnd 0.144101f
C1884 vdd.t201 gnd 0.033041f
C1885 vdd.t259 gnd 0.033041f
C1886 vdd.n271 gnd 0.227082f
C1887 vdd.n272 gnd 0.144101f
C1888 vdd.t260 gnd 0.033041f
C1889 vdd.t176 gnd 0.033041f
C1890 vdd.n273 gnd 0.227082f
C1891 vdd.n274 gnd 0.144101f
C1892 vdd.t248 gnd 0.033041f
C1893 vdd.t256 gnd 0.033041f
C1894 vdd.n275 gnd 0.227082f
C1895 vdd.n276 gnd 0.144101f
C1896 vdd.t162 gnd 0.033041f
C1897 vdd.t222 gnd 0.033041f
C1898 vdd.n277 gnd 0.227082f
C1899 vdd.n278 gnd 0.144101f
C1900 vdd.n279 gnd 0.005632f
C1901 vdd.n280 gnd 0.005227f
C1902 vdd.n281 gnd 0.002891f
C1903 vdd.n282 gnd 0.006638f
C1904 vdd.n283 gnd 0.002809f
C1905 vdd.n284 gnd 0.002974f
C1906 vdd.n285 gnd 0.005227f
C1907 vdd.n286 gnd 0.002809f
C1908 vdd.n287 gnd 0.006638f
C1909 vdd.n288 gnd 0.002974f
C1910 vdd.n289 gnd 0.005227f
C1911 vdd.n290 gnd 0.002809f
C1912 vdd.n291 gnd 0.004979f
C1913 vdd.n292 gnd 0.004994f
C1914 vdd.t243 gnd 0.014262f
C1915 vdd.n293 gnd 0.031732f
C1916 vdd.n294 gnd 0.165142f
C1917 vdd.n295 gnd 0.002809f
C1918 vdd.n296 gnd 0.002974f
C1919 vdd.n297 gnd 0.006638f
C1920 vdd.n298 gnd 0.006638f
C1921 vdd.n299 gnd 0.002974f
C1922 vdd.n300 gnd 0.002809f
C1923 vdd.n301 gnd 0.005227f
C1924 vdd.n302 gnd 0.005227f
C1925 vdd.n303 gnd 0.002809f
C1926 vdd.n304 gnd 0.002974f
C1927 vdd.n305 gnd 0.006638f
C1928 vdd.n306 gnd 0.006638f
C1929 vdd.n307 gnd 0.002974f
C1930 vdd.n308 gnd 0.002809f
C1931 vdd.n309 gnd 0.005227f
C1932 vdd.n310 gnd 0.005227f
C1933 vdd.n311 gnd 0.002809f
C1934 vdd.n312 gnd 0.002974f
C1935 vdd.n313 gnd 0.006638f
C1936 vdd.n314 gnd 0.006638f
C1937 vdd.n315 gnd 0.015694f
C1938 vdd.n316 gnd 0.002891f
C1939 vdd.n317 gnd 0.002809f
C1940 vdd.n318 gnd 0.013509f
C1941 vdd.n319 gnd 0.009135f
C1942 vdd.n320 gnd 0.06378f
C1943 vdd.n321 gnd 0.257364f
C1944 vdd.n322 gnd 0.007888f
C1945 vdd.n323 gnd 0.010263f
C1946 vdd.n324 gnd 0.00826f
C1947 vdd.n325 gnd 0.00826f
C1948 vdd.n326 gnd 0.010263f
C1949 vdd.n327 gnd 0.010263f
C1950 vdd.n328 gnd 0.749897f
C1951 vdd.n329 gnd 0.010263f
C1952 vdd.n330 gnd 0.010263f
C1953 vdd.n331 gnd 0.010263f
C1954 vdd.n332 gnd 0.812826f
C1955 vdd.n333 gnd 0.010263f
C1956 vdd.n334 gnd 0.010263f
C1957 vdd.n335 gnd 0.010263f
C1958 vdd.n336 gnd 0.010263f
C1959 vdd.n337 gnd 0.00826f
C1960 vdd.n338 gnd 0.010263f
C1961 vdd.t152 gnd 0.524404f
C1962 vdd.n339 gnd 0.010263f
C1963 vdd.n340 gnd 0.010263f
C1964 vdd.n341 gnd 0.010263f
C1965 vdd.t228 gnd 0.524404f
C1966 vdd.n342 gnd 0.010263f
C1967 vdd.n343 gnd 0.010263f
C1968 vdd.n344 gnd 0.010263f
C1969 vdd.n345 gnd 0.010263f
C1970 vdd.n346 gnd 0.010263f
C1971 vdd.n347 gnd 0.00826f
C1972 vdd.n348 gnd 0.010263f
C1973 vdd.n349 gnd 0.592576f
C1974 vdd.n350 gnd 0.010263f
C1975 vdd.n351 gnd 0.010263f
C1976 vdd.n352 gnd 0.010263f
C1977 vdd.t206 gnd 0.524404f
C1978 vdd.n353 gnd 0.010263f
C1979 vdd.n354 gnd 0.010263f
C1980 vdd.n355 gnd 0.010263f
C1981 vdd.n356 gnd 0.010263f
C1982 vdd.n357 gnd 0.010263f
C1983 vdd.n358 gnd 0.00826f
C1984 vdd.n359 gnd 0.010263f
C1985 vdd.t194 gnd 0.524404f
C1986 vdd.n360 gnd 0.010263f
C1987 vdd.n361 gnd 0.010263f
C1988 vdd.n362 gnd 0.010263f
C1989 vdd.n363 gnd 0.886242f
C1990 vdd.n364 gnd 0.010263f
C1991 vdd.n365 gnd 0.010263f
C1992 vdd.n366 gnd 0.010263f
C1993 vdd.n367 gnd 0.010263f
C1994 vdd.n368 gnd 0.010263f
C1995 vdd.n369 gnd 0.006856f
C1996 vdd.n370 gnd 0.023371f
C1997 vdd.t83 gnd 0.524404f
C1998 vdd.n371 gnd 0.010263f
C1999 vdd.n372 gnd 0.023371f
C2000 vdd.n404 gnd 0.010263f
C2001 vdd.t85 gnd 0.126259f
C2002 vdd.t84 gnd 0.134936f
C2003 vdd.t82 gnd 0.164893f
C2004 vdd.n405 gnd 0.211369f
C2005 vdd.n406 gnd 0.178414f
C2006 vdd.n407 gnd 0.013547f
C2007 vdd.n408 gnd 0.010263f
C2008 vdd.n409 gnd 0.00826f
C2009 vdd.n410 gnd 0.010263f
C2010 vdd.n411 gnd 0.00826f
C2011 vdd.n412 gnd 0.010263f
C2012 vdd.n413 gnd 0.00826f
C2013 vdd.n414 gnd 0.010263f
C2014 vdd.n415 gnd 0.00826f
C2015 vdd.n416 gnd 0.010263f
C2016 vdd.n417 gnd 0.00826f
C2017 vdd.n418 gnd 0.010263f
C2018 vdd.t118 gnd 0.126259f
C2019 vdd.t117 gnd 0.134936f
C2020 vdd.t116 gnd 0.164893f
C2021 vdd.n419 gnd 0.211369f
C2022 vdd.n420 gnd 0.178414f
C2023 vdd.n421 gnd 0.00826f
C2024 vdd.n422 gnd 0.010263f
C2025 vdd.n423 gnd 0.00826f
C2026 vdd.n424 gnd 0.010263f
C2027 vdd.n425 gnd 0.00826f
C2028 vdd.n426 gnd 0.010263f
C2029 vdd.n427 gnd 0.00826f
C2030 vdd.n428 gnd 0.010263f
C2031 vdd.n429 gnd 0.00826f
C2032 vdd.n430 gnd 0.010263f
C2033 vdd.t124 gnd 0.126259f
C2034 vdd.t123 gnd 0.134936f
C2035 vdd.t122 gnd 0.164893f
C2036 vdd.n431 gnd 0.211369f
C2037 vdd.n432 gnd 0.178414f
C2038 vdd.n433 gnd 0.017677f
C2039 vdd.n434 gnd 0.010263f
C2040 vdd.n435 gnd 0.00826f
C2041 vdd.n436 gnd 0.010263f
C2042 vdd.n437 gnd 0.00826f
C2043 vdd.n438 gnd 0.010263f
C2044 vdd.n439 gnd 0.00826f
C2045 vdd.n440 gnd 0.010263f
C2046 vdd.n441 gnd 0.00826f
C2047 vdd.n442 gnd 0.010263f
C2048 vdd.n443 gnd 0.023371f
C2049 vdd.n444 gnd 0.02353f
C2050 vdd.n445 gnd 0.02353f
C2051 vdd.n446 gnd 0.006856f
C2052 vdd.n447 gnd 0.00826f
C2053 vdd.n448 gnd 0.010263f
C2054 vdd.n449 gnd 0.010263f
C2055 vdd.n450 gnd 0.00826f
C2056 vdd.n451 gnd 0.010263f
C2057 vdd.n452 gnd 0.010263f
C2058 vdd.n453 gnd 0.010263f
C2059 vdd.n454 gnd 0.010263f
C2060 vdd.n455 gnd 0.010263f
C2061 vdd.n456 gnd 0.00826f
C2062 vdd.n457 gnd 0.00826f
C2063 vdd.n458 gnd 0.010263f
C2064 vdd.n459 gnd 0.010263f
C2065 vdd.n460 gnd 0.00826f
C2066 vdd.n461 gnd 0.010263f
C2067 vdd.n462 gnd 0.010263f
C2068 vdd.n463 gnd 0.010263f
C2069 vdd.n464 gnd 0.010263f
C2070 vdd.n465 gnd 0.010263f
C2071 vdd.n466 gnd 0.00826f
C2072 vdd.n467 gnd 0.00826f
C2073 vdd.n468 gnd 0.010263f
C2074 vdd.n469 gnd 0.010263f
C2075 vdd.n470 gnd 0.00826f
C2076 vdd.n471 gnd 0.010263f
C2077 vdd.n472 gnd 0.010263f
C2078 vdd.n473 gnd 0.010263f
C2079 vdd.n474 gnd 0.010263f
C2080 vdd.n475 gnd 0.010263f
C2081 vdd.n476 gnd 0.00826f
C2082 vdd.n477 gnd 0.00826f
C2083 vdd.n478 gnd 0.010263f
C2084 vdd.n479 gnd 0.010263f
C2085 vdd.n480 gnd 0.00826f
C2086 vdd.n481 gnd 0.010263f
C2087 vdd.n482 gnd 0.010263f
C2088 vdd.n483 gnd 0.010263f
C2089 vdd.n484 gnd 0.010263f
C2090 vdd.n485 gnd 0.010263f
C2091 vdd.n486 gnd 0.00826f
C2092 vdd.n487 gnd 0.00826f
C2093 vdd.n488 gnd 0.010263f
C2094 vdd.n489 gnd 0.010263f
C2095 vdd.n490 gnd 0.006897f
C2096 vdd.n491 gnd 0.010263f
C2097 vdd.n492 gnd 0.010263f
C2098 vdd.n493 gnd 0.010263f
C2099 vdd.n494 gnd 0.010263f
C2100 vdd.n495 gnd 0.010263f
C2101 vdd.n496 gnd 0.006897f
C2102 vdd.n497 gnd 0.00826f
C2103 vdd.n498 gnd 0.010263f
C2104 vdd.n499 gnd 0.010263f
C2105 vdd.n500 gnd 0.00826f
C2106 vdd.n501 gnd 0.010263f
C2107 vdd.n502 gnd 0.010263f
C2108 vdd.n503 gnd 0.010263f
C2109 vdd.n504 gnd 0.010263f
C2110 vdd.n505 gnd 0.010263f
C2111 vdd.n506 gnd 0.00826f
C2112 vdd.n507 gnd 0.00826f
C2113 vdd.n508 gnd 0.010263f
C2114 vdd.n509 gnd 0.010263f
C2115 vdd.n510 gnd 0.00826f
C2116 vdd.n511 gnd 0.010263f
C2117 vdd.n512 gnd 0.010263f
C2118 vdd.n513 gnd 0.010263f
C2119 vdd.n514 gnd 0.010263f
C2120 vdd.n515 gnd 0.010263f
C2121 vdd.n516 gnd 0.00826f
C2122 vdd.n517 gnd 0.00826f
C2123 vdd.n518 gnd 0.010263f
C2124 vdd.n519 gnd 0.010263f
C2125 vdd.n520 gnd 0.00826f
C2126 vdd.n521 gnd 0.010263f
C2127 vdd.n522 gnd 0.010263f
C2128 vdd.n523 gnd 0.010263f
C2129 vdd.n524 gnd 0.010263f
C2130 vdd.n525 gnd 0.010263f
C2131 vdd.n526 gnd 0.00826f
C2132 vdd.n527 gnd 0.00826f
C2133 vdd.n528 gnd 0.010263f
C2134 vdd.n529 gnd 0.010263f
C2135 vdd.n530 gnd 0.00826f
C2136 vdd.n531 gnd 0.010263f
C2137 vdd.n532 gnd 0.010263f
C2138 vdd.n533 gnd 0.010263f
C2139 vdd.n534 gnd 0.010263f
C2140 vdd.n535 gnd 0.010263f
C2141 vdd.n536 gnd 0.00826f
C2142 vdd.n537 gnd 0.00826f
C2143 vdd.n538 gnd 0.010263f
C2144 vdd.n539 gnd 0.010263f
C2145 vdd.n540 gnd 0.00826f
C2146 vdd.n541 gnd 0.010263f
C2147 vdd.n542 gnd 0.010263f
C2148 vdd.n543 gnd 0.010263f
C2149 vdd.n544 gnd 0.010263f
C2150 vdd.n545 gnd 0.010263f
C2151 vdd.n546 gnd 0.005617f
C2152 vdd.n547 gnd 0.017677f
C2153 vdd.n548 gnd 0.010263f
C2154 vdd.n549 gnd 0.010263f
C2155 vdd.n550 gnd 0.008178f
C2156 vdd.n551 gnd 0.010263f
C2157 vdd.n552 gnd 0.010263f
C2158 vdd.n553 gnd 0.010263f
C2159 vdd.n554 gnd 0.010263f
C2160 vdd.n555 gnd 0.010263f
C2161 vdd.n556 gnd 0.00826f
C2162 vdd.n557 gnd 0.00826f
C2163 vdd.n558 gnd 0.010263f
C2164 vdd.n559 gnd 0.010263f
C2165 vdd.n560 gnd 0.00826f
C2166 vdd.n561 gnd 0.010263f
C2167 vdd.n562 gnd 0.010263f
C2168 vdd.n563 gnd 0.010263f
C2169 vdd.n564 gnd 0.010263f
C2170 vdd.n565 gnd 0.010263f
C2171 vdd.n566 gnd 0.00826f
C2172 vdd.n567 gnd 0.00826f
C2173 vdd.n568 gnd 0.010263f
C2174 vdd.n569 gnd 0.010263f
C2175 vdd.n570 gnd 0.00826f
C2176 vdd.n571 gnd 0.010263f
C2177 vdd.n572 gnd 0.010263f
C2178 vdd.n573 gnd 0.010263f
C2179 vdd.n574 gnd 0.010263f
C2180 vdd.n575 gnd 0.010263f
C2181 vdd.n576 gnd 0.00826f
C2182 vdd.n577 gnd 0.00826f
C2183 vdd.n578 gnd 0.010263f
C2184 vdd.n579 gnd 0.010263f
C2185 vdd.n580 gnd 0.00826f
C2186 vdd.n581 gnd 0.010263f
C2187 vdd.n582 gnd 0.010263f
C2188 vdd.n583 gnd 0.010263f
C2189 vdd.n584 gnd 0.010263f
C2190 vdd.n585 gnd 0.010263f
C2191 vdd.n586 gnd 0.00826f
C2192 vdd.n587 gnd 0.00826f
C2193 vdd.n588 gnd 0.010263f
C2194 vdd.n589 gnd 0.010263f
C2195 vdd.n590 gnd 0.00826f
C2196 vdd.n591 gnd 0.010263f
C2197 vdd.n592 gnd 0.010263f
C2198 vdd.n593 gnd 0.010263f
C2199 vdd.n594 gnd 0.010263f
C2200 vdd.n595 gnd 0.010263f
C2201 vdd.n596 gnd 0.00826f
C2202 vdd.n597 gnd 0.010263f
C2203 vdd.n598 gnd 0.00826f
C2204 vdd.n599 gnd 0.004337f
C2205 vdd.n600 gnd 0.010263f
C2206 vdd.n601 gnd 0.010263f
C2207 vdd.n602 gnd 0.00826f
C2208 vdd.n603 gnd 0.010263f
C2209 vdd.n604 gnd 0.00826f
C2210 vdd.n605 gnd 0.010263f
C2211 vdd.n606 gnd 0.00826f
C2212 vdd.n607 gnd 0.010263f
C2213 vdd.n608 gnd 0.00826f
C2214 vdd.n609 gnd 0.010263f
C2215 vdd.n610 gnd 0.00826f
C2216 vdd.n611 gnd 0.010263f
C2217 vdd.n612 gnd 0.010263f
C2218 vdd.n613 gnd 0.5716f
C2219 vdd.t154 gnd 0.524404f
C2220 vdd.n614 gnd 0.010263f
C2221 vdd.n615 gnd 0.00826f
C2222 vdd.n616 gnd 0.010263f
C2223 vdd.n617 gnd 0.00826f
C2224 vdd.n618 gnd 0.010263f
C2225 vdd.t144 gnd 0.524404f
C2226 vdd.n619 gnd 0.010263f
C2227 vdd.n620 gnd 0.00826f
C2228 vdd.n621 gnd 0.010263f
C2229 vdd.n622 gnd 0.00826f
C2230 vdd.n623 gnd 0.010263f
C2231 vdd.t187 gnd 0.524404f
C2232 vdd.n624 gnd 0.655505f
C2233 vdd.n625 gnd 0.010263f
C2234 vdd.n626 gnd 0.00826f
C2235 vdd.n627 gnd 0.010263f
C2236 vdd.n628 gnd 0.00826f
C2237 vdd.n629 gnd 0.010263f
C2238 vdd.t185 gnd 0.524404f
C2239 vdd.n630 gnd 0.010263f
C2240 vdd.n631 gnd 0.00826f
C2241 vdd.n632 gnd 0.010263f
C2242 vdd.n633 gnd 0.00826f
C2243 vdd.n634 gnd 0.010263f
C2244 vdd.n635 gnd 0.728921f
C2245 vdd.n636 gnd 0.87051f
C2246 vdd.t136 gnd 0.524404f
C2247 vdd.n637 gnd 0.010263f
C2248 vdd.n638 gnd 0.00826f
C2249 vdd.n639 gnd 0.010263f
C2250 vdd.n640 gnd 0.00826f
C2251 vdd.n641 gnd 0.010263f
C2252 vdd.n642 gnd 0.550624f
C2253 vdd.n643 gnd 0.010263f
C2254 vdd.n644 gnd 0.00826f
C2255 vdd.n645 gnd 0.010263f
C2256 vdd.n646 gnd 0.00826f
C2257 vdd.n647 gnd 0.010263f
C2258 vdd.n648 gnd 1.04881f
C2259 vdd.t177 gnd 0.524404f
C2260 vdd.n649 gnd 0.010263f
C2261 vdd.n650 gnd 0.00826f
C2262 vdd.n651 gnd 0.010263f
C2263 vdd.n652 gnd 0.00826f
C2264 vdd.n653 gnd 0.010263f
C2265 vdd.t58 gnd 0.524404f
C2266 vdd.n654 gnd 0.010263f
C2267 vdd.n655 gnd 0.00826f
C2268 vdd.n656 gnd 0.02353f
C2269 vdd.n657 gnd 0.02353f
C2270 vdd.n658 gnd 9.15609f
C2271 vdd.n659 gnd 0.582088f
C2272 vdd.n660 gnd 0.02353f
C2273 vdd.n661 gnd 0.008826f
C2274 vdd.n662 gnd 0.00826f
C2275 vdd.n667 gnd 0.006568f
C2276 vdd.n668 gnd 0.00826f
C2277 vdd.n669 gnd 0.010263f
C2278 vdd.n670 gnd 0.010263f
C2279 vdd.n671 gnd 0.010263f
C2280 vdd.n672 gnd 0.010263f
C2281 vdd.n673 gnd 0.010263f
C2282 vdd.n674 gnd 0.00826f
C2283 vdd.n675 gnd 0.010263f
C2284 vdd.n676 gnd 0.010263f
C2285 vdd.n677 gnd 0.010263f
C2286 vdd.n678 gnd 0.010263f
C2287 vdd.n679 gnd 0.010263f
C2288 vdd.n680 gnd 0.00826f
C2289 vdd.n681 gnd 0.010263f
C2290 vdd.n682 gnd 0.010263f
C2291 vdd.n683 gnd 0.010263f
C2292 vdd.n684 gnd 0.010263f
C2293 vdd.n685 gnd 0.010263f
C2294 vdd.t76 gnd 0.126259f
C2295 vdd.t77 gnd 0.134936f
C2296 vdd.t75 gnd 0.164893f
C2297 vdd.n686 gnd 0.211369f
C2298 vdd.n687 gnd 0.177588f
C2299 vdd.n688 gnd 0.016851f
C2300 vdd.n689 gnd 0.010263f
C2301 vdd.n690 gnd 0.010263f
C2302 vdd.n691 gnd 0.010263f
C2303 vdd.n692 gnd 0.010263f
C2304 vdd.n693 gnd 0.010263f
C2305 vdd.n694 gnd 0.00826f
C2306 vdd.n695 gnd 0.010263f
C2307 vdd.n696 gnd 0.010263f
C2308 vdd.n697 gnd 0.010263f
C2309 vdd.n698 gnd 0.010263f
C2310 vdd.n699 gnd 0.010263f
C2311 vdd.n700 gnd 0.00826f
C2312 vdd.n701 gnd 0.010263f
C2313 vdd.n702 gnd 0.010263f
C2314 vdd.n703 gnd 0.010263f
C2315 vdd.n704 gnd 0.010263f
C2316 vdd.n705 gnd 0.010263f
C2317 vdd.n706 gnd 0.00826f
C2318 vdd.n707 gnd 0.010263f
C2319 vdd.n708 gnd 0.010263f
C2320 vdd.n709 gnd 0.010263f
C2321 vdd.n710 gnd 0.010263f
C2322 vdd.n711 gnd 0.010263f
C2323 vdd.n712 gnd 0.00826f
C2324 vdd.n713 gnd 0.010263f
C2325 vdd.n714 gnd 0.010263f
C2326 vdd.n715 gnd 0.010263f
C2327 vdd.n716 gnd 0.010263f
C2328 vdd.n717 gnd 0.010263f
C2329 vdd.n718 gnd 0.00826f
C2330 vdd.n719 gnd 0.010263f
C2331 vdd.n720 gnd 0.010263f
C2332 vdd.n721 gnd 0.010263f
C2333 vdd.n722 gnd 0.008178f
C2334 vdd.t66 gnd 0.126259f
C2335 vdd.t67 gnd 0.134936f
C2336 vdd.t65 gnd 0.164893f
C2337 vdd.n723 gnd 0.211369f
C2338 vdd.n724 gnd 0.177588f
C2339 vdd.n725 gnd 0.010263f
C2340 vdd.n726 gnd 0.00826f
C2341 vdd.n728 gnd 0.010263f
C2342 vdd.n730 gnd 0.010263f
C2343 vdd.n731 gnd 0.010263f
C2344 vdd.n732 gnd 0.00826f
C2345 vdd.n733 gnd 0.010263f
C2346 vdd.n734 gnd 0.010263f
C2347 vdd.n735 gnd 0.010263f
C2348 vdd.n736 gnd 0.010263f
C2349 vdd.n737 gnd 0.010263f
C2350 vdd.n738 gnd 0.00826f
C2351 vdd.n739 gnd 0.010263f
C2352 vdd.n740 gnd 0.010263f
C2353 vdd.n741 gnd 0.010263f
C2354 vdd.n742 gnd 0.010263f
C2355 vdd.n743 gnd 0.010263f
C2356 vdd.n744 gnd 0.00826f
C2357 vdd.n745 gnd 0.010263f
C2358 vdd.n746 gnd 0.010263f
C2359 vdd.n747 gnd 0.010263f
C2360 vdd.n748 gnd 0.006568f
C2361 vdd.n753 gnd 0.006979f
C2362 vdd.n754 gnd 0.006979f
C2363 vdd.n755 gnd 0.006979f
C2364 vdd.n756 gnd 8.94633f
C2365 vdd.n757 gnd 0.006979f
C2366 vdd.n758 gnd 0.006979f
C2367 vdd.n759 gnd 0.006979f
C2368 vdd.n761 gnd 0.006979f
C2369 vdd.n762 gnd 0.006979f
C2370 vdd.n764 gnd 0.006979f
C2371 vdd.n765 gnd 0.00508f
C2372 vdd.n767 gnd 0.006979f
C2373 vdd.t52 gnd 0.282008f
C2374 vdd.t51 gnd 0.28867f
C2375 vdd.t49 gnd 0.184106f
C2376 vdd.n768 gnd 0.099499f
C2377 vdd.n769 gnd 0.056439f
C2378 vdd.n770 gnd 0.009974f
C2379 vdd.n771 gnd 0.016154f
C2380 vdd.n773 gnd 0.006979f
C2381 vdd.n774 gnd 0.713189f
C2382 vdd.n775 gnd 0.015287f
C2383 vdd.n776 gnd 0.015287f
C2384 vdd.n777 gnd 0.006979f
C2385 vdd.n778 gnd 0.016323f
C2386 vdd.n779 gnd 0.006979f
C2387 vdd.n780 gnd 0.006979f
C2388 vdd.n781 gnd 0.006979f
C2389 vdd.n782 gnd 0.006979f
C2390 vdd.n783 gnd 0.006979f
C2391 vdd.n785 gnd 0.006979f
C2392 vdd.n786 gnd 0.006979f
C2393 vdd.n788 gnd 0.006979f
C2394 vdd.n789 gnd 0.006979f
C2395 vdd.n791 gnd 0.006979f
C2396 vdd.n792 gnd 0.006979f
C2397 vdd.n794 gnd 0.006979f
C2398 vdd.n795 gnd 0.006979f
C2399 vdd.n797 gnd 0.006979f
C2400 vdd.n798 gnd 0.006979f
C2401 vdd.n800 gnd 0.006979f
C2402 vdd.n801 gnd 0.00508f
C2403 vdd.n803 gnd 0.006979f
C2404 vdd.t121 gnd 0.282008f
C2405 vdd.t120 gnd 0.28867f
C2406 vdd.t119 gnd 0.184106f
C2407 vdd.n804 gnd 0.099499f
C2408 vdd.n805 gnd 0.056439f
C2409 vdd.n806 gnd 0.009974f
C2410 vdd.n807 gnd 0.006979f
C2411 vdd.n808 gnd 0.006979f
C2412 vdd.t50 gnd 0.356594f
C2413 vdd.n809 gnd 0.006979f
C2414 vdd.n810 gnd 0.006979f
C2415 vdd.n811 gnd 0.006979f
C2416 vdd.n812 gnd 0.006979f
C2417 vdd.n813 gnd 0.006979f
C2418 vdd.n814 gnd 0.713189f
C2419 vdd.n815 gnd 0.006979f
C2420 vdd.n816 gnd 0.006979f
C2421 vdd.n817 gnd 0.603064f
C2422 vdd.n818 gnd 0.006979f
C2423 vdd.n819 gnd 0.006979f
C2424 vdd.n820 gnd 0.006979f
C2425 vdd.n821 gnd 0.006979f
C2426 vdd.n822 gnd 0.697457f
C2427 vdd.n823 gnd 0.006979f
C2428 vdd.n824 gnd 0.006979f
C2429 vdd.n825 gnd 0.006979f
C2430 vdd.n826 gnd 0.006979f
C2431 vdd.n827 gnd 0.006979f
C2432 vdd.n828 gnd 0.713189f
C2433 vdd.n829 gnd 0.006979f
C2434 vdd.n830 gnd 0.006979f
C2435 vdd.t21 gnd 0.356594f
C2436 vdd.n831 gnd 0.006979f
C2437 vdd.n832 gnd 0.006979f
C2438 vdd.n833 gnd 0.006979f
C2439 vdd.t41 gnd 0.356594f
C2440 vdd.n834 gnd 0.006979f
C2441 vdd.n835 gnd 0.006979f
C2442 vdd.n836 gnd 0.006979f
C2443 vdd.n837 gnd 0.006979f
C2444 vdd.n838 gnd 0.006979f
C2445 vdd.t72 gnd 0.29891f
C2446 vdd.n839 gnd 0.006979f
C2447 vdd.n840 gnd 0.006979f
C2448 vdd.n841 gnd 0.5716f
C2449 vdd.n842 gnd 0.006979f
C2450 vdd.t73 gnd 0.28867f
C2451 vdd.t71 gnd 0.184106f
C2452 vdd.t74 gnd 0.28867f
C2453 vdd.n843 gnd 0.162244f
C2454 vdd.n844 gnd 0.006979f
C2455 vdd.n845 gnd 0.006979f
C2456 vdd.n846 gnd 0.456231f
C2457 vdd.n847 gnd 0.006979f
C2458 vdd.n848 gnd 0.006979f
C2459 vdd.t34 gnd 0.104881f
C2460 vdd.n849 gnd 0.414279f
C2461 vdd.n850 gnd 0.006979f
C2462 vdd.n851 gnd 0.006979f
C2463 vdd.n852 gnd 0.006979f
C2464 vdd.n853 gnd 0.613552f
C2465 vdd.n854 gnd 0.006979f
C2466 vdd.n855 gnd 0.006979f
C2467 vdd.t126 gnd 0.356594f
C2468 vdd.n856 gnd 0.006979f
C2469 vdd.n857 gnd 0.006979f
C2470 vdd.n858 gnd 0.006979f
C2471 vdd.t264 gnd 0.356594f
C2472 vdd.n859 gnd 0.006979f
C2473 vdd.n860 gnd 0.006979f
C2474 vdd.t14 gnd 0.356594f
C2475 vdd.n861 gnd 0.006979f
C2476 vdd.n862 gnd 0.006979f
C2477 vdd.n863 gnd 0.006979f
C2478 vdd.t40 gnd 0.283178f
C2479 vdd.n864 gnd 0.006979f
C2480 vdd.n865 gnd 0.006979f
C2481 vdd.n866 gnd 0.587332f
C2482 vdd.n867 gnd 0.006979f
C2483 vdd.n868 gnd 0.006979f
C2484 vdd.n869 gnd 0.006979f
C2485 vdd.t37 gnd 0.356594f
C2486 vdd.n870 gnd 0.006979f
C2487 vdd.n871 gnd 0.006979f
C2488 vdd.t15 gnd 0.29891f
C2489 vdd.n872 gnd 0.430011f
C2490 vdd.n873 gnd 0.006979f
C2491 vdd.n874 gnd 0.006979f
C2492 vdd.n875 gnd 0.006979f
C2493 vdd.n876 gnd 0.372327f
C2494 vdd.n877 gnd 0.006979f
C2495 vdd.n878 gnd 0.006979f
C2496 vdd.t9 gnd 0.356594f
C2497 vdd.n879 gnd 0.006979f
C2498 vdd.n880 gnd 0.006979f
C2499 vdd.n881 gnd 0.006979f
C2500 vdd.n882 gnd 0.713189f
C2501 vdd.n883 gnd 0.006979f
C2502 vdd.n884 gnd 0.006979f
C2503 vdd.t8 gnd 0.241226f
C2504 vdd.t134 gnd 0.340862f
C2505 vdd.n885 gnd 0.006979f
C2506 vdd.n886 gnd 0.006979f
C2507 vdd.n887 gnd 0.006979f
C2508 vdd.n888 gnd 0.534892f
C2509 vdd.n889 gnd 0.006979f
C2510 vdd.n890 gnd 0.006979f
C2511 vdd.n891 gnd 0.006979f
C2512 vdd.n892 gnd 0.006979f
C2513 vdd.n893 gnd 0.006979f
C2514 vdd.t100 gnd 0.356594f
C2515 vdd.n894 gnd 0.006979f
C2516 vdd.n895 gnd 0.006979f
C2517 vdd.t42 gnd 0.356594f
C2518 vdd.n896 gnd 0.006979f
C2519 vdd.n897 gnd 0.015287f
C2520 vdd.n898 gnd 0.015287f
C2521 vdd.n899 gnd 0.849534f
C2522 vdd.n900 gnd 0.006979f
C2523 vdd.n901 gnd 0.006979f
C2524 vdd.t47 gnd 0.356594f
C2525 vdd.n902 gnd 0.015287f
C2526 vdd.n903 gnd 0.006979f
C2527 vdd.n904 gnd 0.006979f
C2528 vdd.t19 gnd 0.650261f
C2529 vdd.n922 gnd 0.016323f
C2530 vdd.n940 gnd 0.015287f
C2531 vdd.n941 gnd 0.006979f
C2532 vdd.n942 gnd 0.015287f
C2533 vdd.t115 gnd 0.282008f
C2534 vdd.t114 gnd 0.28867f
C2535 vdd.t113 gnd 0.184106f
C2536 vdd.n943 gnd 0.099499f
C2537 vdd.n944 gnd 0.056439f
C2538 vdd.n945 gnd 0.016154f
C2539 vdd.n946 gnd 0.006979f
C2540 vdd.n947 gnd 0.377571f
C2541 vdd.n948 gnd 0.015287f
C2542 vdd.n949 gnd 0.006979f
C2543 vdd.n950 gnd 0.016323f
C2544 vdd.n951 gnd 0.006979f
C2545 vdd.t98 gnd 0.282008f
C2546 vdd.t97 gnd 0.28867f
C2547 vdd.t95 gnd 0.184106f
C2548 vdd.n952 gnd 0.099499f
C2549 vdd.n953 gnd 0.056439f
C2550 vdd.n954 gnd 0.009974f
C2551 vdd.n955 gnd 0.006979f
C2552 vdd.n956 gnd 0.006979f
C2553 vdd.t96 gnd 0.356594f
C2554 vdd.n957 gnd 0.006979f
C2555 vdd.t17 gnd 0.356594f
C2556 vdd.n958 gnd 0.006979f
C2557 vdd.n959 gnd 0.006979f
C2558 vdd.n960 gnd 0.006979f
C2559 vdd.n961 gnd 0.006979f
C2560 vdd.n962 gnd 0.006979f
C2561 vdd.n963 gnd 0.713189f
C2562 vdd.n964 gnd 0.006979f
C2563 vdd.n965 gnd 0.006979f
C2564 vdd.t127 gnd 0.356594f
C2565 vdd.n966 gnd 0.006979f
C2566 vdd.n967 gnd 0.006979f
C2567 vdd.n968 gnd 0.006979f
C2568 vdd.n969 gnd 0.006979f
C2569 vdd.n970 gnd 0.471963f
C2570 vdd.n971 gnd 0.006979f
C2571 vdd.n972 gnd 0.006979f
C2572 vdd.n973 gnd 0.006979f
C2573 vdd.n974 gnd 0.006979f
C2574 vdd.n975 gnd 0.006979f
C2575 vdd.n976 gnd 0.629284f
C2576 vdd.n977 gnd 0.006979f
C2577 vdd.n978 gnd 0.006979f
C2578 vdd.t45 gnd 0.340862f
C2579 vdd.t22 gnd 0.241226f
C2580 vdd.n979 gnd 0.006979f
C2581 vdd.n980 gnd 0.006979f
C2582 vdd.n981 gnd 0.006979f
C2583 vdd.t131 gnd 0.356594f
C2584 vdd.n982 gnd 0.006979f
C2585 vdd.n983 gnd 0.006979f
C2586 vdd.t32 gnd 0.356594f
C2587 vdd.n984 gnd 0.006979f
C2588 vdd.n985 gnd 0.006979f
C2589 vdd.n986 gnd 0.006979f
C2590 vdd.t129 gnd 0.29891f
C2591 vdd.n987 gnd 0.006979f
C2592 vdd.n988 gnd 0.006979f
C2593 vdd.n989 gnd 0.5716f
C2594 vdd.n990 gnd 0.006979f
C2595 vdd.n991 gnd 0.006979f
C2596 vdd.n992 gnd 0.006979f
C2597 vdd.t11 gnd 0.356594f
C2598 vdd.n993 gnd 0.006979f
C2599 vdd.n994 gnd 0.006979f
C2600 vdd.t44 gnd 0.283178f
C2601 vdd.n995 gnd 0.414279f
C2602 vdd.n996 gnd 0.006979f
C2603 vdd.n997 gnd 0.006979f
C2604 vdd.n998 gnd 0.006979f
C2605 vdd.n999 gnd 0.613552f
C2606 vdd.n1000 gnd 0.006979f
C2607 vdd.n1001 gnd 0.006979f
C2608 vdd.t5 gnd 0.356594f
C2609 vdd.n1002 gnd 0.006979f
C2610 vdd.n1003 gnd 0.006979f
C2611 vdd.n1004 gnd 0.006979f
C2612 vdd.n1005 gnd 0.713189f
C2613 vdd.n1006 gnd 0.006979f
C2614 vdd.n1007 gnd 0.006979f
C2615 vdd.t35 gnd 0.356594f
C2616 vdd.n1008 gnd 0.006979f
C2617 vdd.n1009 gnd 0.006979f
C2618 vdd.n1010 gnd 0.006979f
C2619 vdd.t36 gnd 0.104881f
C2620 vdd.n1011 gnd 0.006979f
C2621 vdd.n1012 gnd 0.006979f
C2622 vdd.n1013 gnd 0.006979f
C2623 vdd.t105 gnd 0.28867f
C2624 vdd.t103 gnd 0.184106f
C2625 vdd.t106 gnd 0.28867f
C2626 vdd.n1014 gnd 0.162244f
C2627 vdd.n1015 gnd 0.006979f
C2628 vdd.n1016 gnd 0.006979f
C2629 vdd.t13 gnd 0.356594f
C2630 vdd.n1017 gnd 0.006979f
C2631 vdd.n1018 gnd 0.006979f
C2632 vdd.t104 gnd 0.29891f
C2633 vdd.n1019 gnd 0.608308f
C2634 vdd.n1020 gnd 0.006979f
C2635 vdd.n1021 gnd 0.006979f
C2636 vdd.n1022 gnd 0.006979f
C2637 vdd.n1023 gnd 0.372327f
C2638 vdd.n1024 gnd 0.006979f
C2639 vdd.n1025 gnd 0.006979f
C2640 vdd.n1026 gnd 0.498183f
C2641 vdd.n1027 gnd 0.006979f
C2642 vdd.n1028 gnd 0.006979f
C2643 vdd.n1029 gnd 0.006979f
C2644 vdd.n1030 gnd 0.713189f
C2645 vdd.n1031 gnd 0.006979f
C2646 vdd.n1032 gnd 0.006979f
C2647 vdd.t125 gnd 0.356594f
C2648 vdd.n1033 gnd 0.006979f
C2649 vdd.n1034 gnd 0.006979f
C2650 vdd.n1035 gnd 0.006979f
C2651 vdd.n1036 gnd 0.713189f
C2652 vdd.n1037 gnd 0.006979f
C2653 vdd.n1038 gnd 0.006979f
C2654 vdd.n1039 gnd 0.006979f
C2655 vdd.n1040 gnd 0.006979f
C2656 vdd.n1041 gnd 0.006979f
C2657 vdd.t54 gnd 0.356594f
C2658 vdd.n1042 gnd 0.006979f
C2659 vdd.n1043 gnd 0.006979f
C2660 vdd.n1044 gnd 0.006979f
C2661 vdd.n1045 gnd 0.015287f
C2662 vdd.n1046 gnd 0.015287f
C2663 vdd.n1047 gnd 1.00686f
C2664 vdd.n1048 gnd 0.006979f
C2665 vdd.n1049 gnd 0.006979f
C2666 vdd.n1050 gnd 0.466719f
C2667 vdd.n1051 gnd 0.015287f
C2668 vdd.n1052 gnd 0.006979f
C2669 vdd.n1053 gnd 0.006979f
C2670 vdd.n1054 gnd 9.15609f
C2671 vdd.n1087 gnd 0.016323f
C2672 vdd.n1088 gnd 0.006979f
C2673 vdd.n1089 gnd 0.006979f
C2674 vdd.n1090 gnd 0.006979f
C2675 vdd.n1091 gnd 0.006568f
C2676 vdd.n1094 gnd 0.02353f
C2677 vdd.n1095 gnd 0.006856f
C2678 vdd.n1096 gnd 0.00826f
C2679 vdd.n1098 gnd 0.010263f
C2680 vdd.n1099 gnd 0.010263f
C2681 vdd.n1100 gnd 0.00826f
C2682 vdd.n1102 gnd 0.010263f
C2683 vdd.n1103 gnd 0.010263f
C2684 vdd.n1104 gnd 0.010263f
C2685 vdd.n1105 gnd 0.010263f
C2686 vdd.n1106 gnd 0.010263f
C2687 vdd.n1107 gnd 0.00826f
C2688 vdd.n1109 gnd 0.010263f
C2689 vdd.n1110 gnd 0.010263f
C2690 vdd.n1111 gnd 0.010263f
C2691 vdd.n1112 gnd 0.010263f
C2692 vdd.n1113 gnd 0.010263f
C2693 vdd.n1114 gnd 0.00826f
C2694 vdd.n1116 gnd 0.010263f
C2695 vdd.n1117 gnd 0.010263f
C2696 vdd.n1118 gnd 0.010263f
C2697 vdd.n1119 gnd 0.010263f
C2698 vdd.n1120 gnd 0.006897f
C2699 vdd.t109 gnd 0.126259f
C2700 vdd.t108 gnd 0.134936f
C2701 vdd.t107 gnd 0.164893f
C2702 vdd.n1121 gnd 0.211369f
C2703 vdd.n1122 gnd 0.177588f
C2704 vdd.n1124 gnd 0.010263f
C2705 vdd.n1125 gnd 0.010263f
C2706 vdd.n1126 gnd 0.00826f
C2707 vdd.n1127 gnd 0.010263f
C2708 vdd.n1129 gnd 0.010263f
C2709 vdd.n1130 gnd 0.010263f
C2710 vdd.n1131 gnd 0.010263f
C2711 vdd.n1132 gnd 0.010263f
C2712 vdd.n1133 gnd 0.00826f
C2713 vdd.n1135 gnd 0.010263f
C2714 vdd.n1136 gnd 0.010263f
C2715 vdd.n1137 gnd 0.010263f
C2716 vdd.n1138 gnd 0.010263f
C2717 vdd.n1139 gnd 0.010263f
C2718 vdd.n1140 gnd 0.00826f
C2719 vdd.n1142 gnd 0.010263f
C2720 vdd.n1143 gnd 0.010263f
C2721 vdd.n1144 gnd 0.010263f
C2722 vdd.n1145 gnd 0.010263f
C2723 vdd.n1146 gnd 0.010263f
C2724 vdd.n1147 gnd 0.00826f
C2725 vdd.n1149 gnd 0.010263f
C2726 vdd.n1150 gnd 0.010263f
C2727 vdd.n1151 gnd 0.010263f
C2728 vdd.n1152 gnd 0.010263f
C2729 vdd.n1153 gnd 0.010263f
C2730 vdd.n1154 gnd 0.00826f
C2731 vdd.n1156 gnd 0.010263f
C2732 vdd.n1157 gnd 0.010263f
C2733 vdd.n1158 gnd 0.010263f
C2734 vdd.n1159 gnd 0.010263f
C2735 vdd.n1160 gnd 0.008178f
C2736 vdd.t94 gnd 0.126259f
C2737 vdd.t93 gnd 0.134936f
C2738 vdd.t92 gnd 0.164893f
C2739 vdd.n1161 gnd 0.211369f
C2740 vdd.n1162 gnd 0.177588f
C2741 vdd.n1164 gnd 0.010263f
C2742 vdd.n1165 gnd 0.010263f
C2743 vdd.n1166 gnd 0.00826f
C2744 vdd.n1167 gnd 0.010263f
C2745 vdd.n1169 gnd 0.010263f
C2746 vdd.n1170 gnd 0.010263f
C2747 vdd.n1171 gnd 0.010263f
C2748 vdd.n1172 gnd 0.010263f
C2749 vdd.n1173 gnd 0.00826f
C2750 vdd.n1175 gnd 0.010263f
C2751 vdd.n1176 gnd 0.010263f
C2752 vdd.n1177 gnd 0.010263f
C2753 vdd.n1178 gnd 0.010263f
C2754 vdd.n1179 gnd 0.010263f
C2755 vdd.n1180 gnd 0.00826f
C2756 vdd.n1182 gnd 0.010263f
C2757 vdd.n1183 gnd 0.010263f
C2758 vdd.n1184 gnd 0.010263f
C2759 vdd.n1185 gnd 0.010263f
C2760 vdd.n1186 gnd 0.010263f
C2761 vdd.n1187 gnd 0.00826f
C2762 vdd.n1189 gnd 0.010263f
C2763 vdd.n1190 gnd 0.010263f
C2764 vdd.n1191 gnd 0.006568f
C2765 vdd.n1192 gnd 0.00826f
C2766 vdd.n1193 gnd 0.006979f
C2767 vdd.n1194 gnd 0.006979f
C2768 vdd.n1195 gnd 0.006979f
C2769 vdd.n1196 gnd 0.006979f
C2770 vdd.n1197 gnd 0.006979f
C2771 vdd.n1198 gnd 0.006979f
C2772 vdd.n1199 gnd 0.006979f
C2773 vdd.n1200 gnd 0.006979f
C2774 vdd.n1201 gnd 0.006979f
C2775 vdd.n1202 gnd 0.006979f
C2776 vdd.n1203 gnd 0.006979f
C2777 vdd.n1204 gnd 0.006979f
C2778 vdd.n1205 gnd 0.006979f
C2779 vdd.n1206 gnd 0.006979f
C2780 vdd.n1207 gnd 0.006979f
C2781 vdd.n1208 gnd 0.006979f
C2782 vdd.n1209 gnd 0.006979f
C2783 vdd.n1210 gnd 0.006979f
C2784 vdd.n1211 gnd 0.006979f
C2785 vdd.n1212 gnd 0.006979f
C2786 vdd.n1213 gnd 0.006979f
C2787 vdd.n1214 gnd 0.006979f
C2788 vdd.n1215 gnd 0.006979f
C2789 vdd.n1216 gnd 0.006979f
C2790 vdd.n1217 gnd 0.006979f
C2791 vdd.n1218 gnd 0.006979f
C2792 vdd.n1219 gnd 0.006979f
C2793 vdd.n1220 gnd 0.006979f
C2794 vdd.n1221 gnd 0.006979f
C2795 vdd.n1222 gnd 0.006979f
C2796 vdd.n1223 gnd 0.006979f
C2797 vdd.t55 gnd 0.282008f
C2798 vdd.t56 gnd 0.28867f
C2799 vdd.t53 gnd 0.184106f
C2800 vdd.n1224 gnd 0.099499f
C2801 vdd.n1225 gnd 0.056439f
C2802 vdd.n1226 gnd 0.009974f
C2803 vdd.n1227 gnd 0.006979f
C2804 vdd.n1228 gnd 0.006979f
C2805 vdd.n1229 gnd 0.006979f
C2806 vdd.n1230 gnd 0.006979f
C2807 vdd.n1231 gnd 0.006979f
C2808 vdd.n1232 gnd 0.006979f
C2809 vdd.n1233 gnd 0.006979f
C2810 vdd.n1234 gnd 0.006979f
C2811 vdd.n1235 gnd 0.006979f
C2812 vdd.n1236 gnd 0.006979f
C2813 vdd.n1237 gnd 0.006979f
C2814 vdd.n1238 gnd 0.006979f
C2815 vdd.n1239 gnd 0.006979f
C2816 vdd.n1240 gnd 0.006979f
C2817 vdd.n1241 gnd 0.006979f
C2818 vdd.n1242 gnd 0.006979f
C2819 vdd.n1243 gnd 0.006979f
C2820 vdd.t69 gnd 0.282008f
C2821 vdd.t70 gnd 0.28867f
C2822 vdd.t68 gnd 0.184106f
C2823 vdd.n1244 gnd 0.099499f
C2824 vdd.n1245 gnd 0.056439f
C2825 vdd.n1246 gnd 0.006979f
C2826 vdd.n1247 gnd 0.006979f
C2827 vdd.n1248 gnd 0.006979f
C2828 vdd.n1249 gnd 0.006979f
C2829 vdd.n1250 gnd 0.006979f
C2830 vdd.n1251 gnd 0.006979f
C2831 vdd.n1252 gnd 0.006979f
C2832 vdd.n1253 gnd 0.006979f
C2833 vdd.n1254 gnd 0.006979f
C2834 vdd.n1255 gnd 0.006979f
C2835 vdd.n1256 gnd 0.006979f
C2836 vdd.n1257 gnd 0.006979f
C2837 vdd.n1258 gnd 0.006979f
C2838 vdd.n1259 gnd 0.006979f
C2839 vdd.n1260 gnd 0.006979f
C2840 vdd.n1261 gnd 0.006979f
C2841 vdd.n1262 gnd 0.006979f
C2842 vdd.n1263 gnd 0.006979f
C2843 vdd.n1264 gnd 0.006979f
C2844 vdd.n1265 gnd 0.006979f
C2845 vdd.n1266 gnd 0.006979f
C2846 vdd.n1267 gnd 0.006979f
C2847 vdd.n1268 gnd 0.006979f
C2848 vdd.n1269 gnd 0.006979f
C2849 vdd.n1270 gnd 0.006979f
C2850 vdd.n1271 gnd 0.006979f
C2851 vdd.n1272 gnd 0.00508f
C2852 vdd.n1273 gnd 0.009974f
C2853 vdd.n1274 gnd 0.005388f
C2854 vdd.n1275 gnd 0.006979f
C2855 vdd.n1276 gnd 0.006979f
C2856 vdd.n1277 gnd 0.006979f
C2857 vdd.n1278 gnd 0.016323f
C2858 vdd.n1279 gnd 0.016323f
C2859 vdd.n1280 gnd 0.015287f
C2860 vdd.n1281 gnd 0.015287f
C2861 vdd.n1282 gnd 0.006979f
C2862 vdd.n1283 gnd 0.006979f
C2863 vdd.n1284 gnd 0.006979f
C2864 vdd.n1285 gnd 0.006979f
C2865 vdd.n1286 gnd 0.006979f
C2866 vdd.n1287 gnd 0.006979f
C2867 vdd.n1288 gnd 0.006979f
C2868 vdd.n1289 gnd 0.006979f
C2869 vdd.n1290 gnd 0.006979f
C2870 vdd.n1291 gnd 0.006979f
C2871 vdd.n1292 gnd 0.006979f
C2872 vdd.n1293 gnd 0.006979f
C2873 vdd.n1294 gnd 0.006979f
C2874 vdd.n1295 gnd 0.006979f
C2875 vdd.n1296 gnd 0.006979f
C2876 vdd.n1297 gnd 0.006979f
C2877 vdd.n1298 gnd 0.006979f
C2878 vdd.n1299 gnd 0.006979f
C2879 vdd.n1300 gnd 0.006979f
C2880 vdd.n1301 gnd 0.006979f
C2881 vdd.n1302 gnd 0.006979f
C2882 vdd.n1303 gnd 0.006979f
C2883 vdd.n1304 gnd 0.006979f
C2884 vdd.n1305 gnd 0.006979f
C2885 vdd.n1306 gnd 0.006979f
C2886 vdd.n1307 gnd 0.006979f
C2887 vdd.n1308 gnd 0.006979f
C2888 vdd.n1309 gnd 0.424767f
C2889 vdd.n1310 gnd 0.006979f
C2890 vdd.n1311 gnd 0.006979f
C2891 vdd.n1312 gnd 0.006979f
C2892 vdd.n1313 gnd 0.006979f
C2893 vdd.n1314 gnd 0.006979f
C2894 vdd.n1315 gnd 0.006979f
C2895 vdd.n1316 gnd 0.006979f
C2896 vdd.n1317 gnd 0.006979f
C2897 vdd.n1318 gnd 0.006979f
C2898 vdd.n1319 gnd 0.006979f
C2899 vdd.n1320 gnd 0.006979f
C2900 vdd.n1321 gnd 0.006979f
C2901 vdd.n1322 gnd 0.006979f
C2902 vdd.n1323 gnd 0.006979f
C2903 vdd.n1324 gnd 0.006979f
C2904 vdd.n1325 gnd 0.006979f
C2905 vdd.n1326 gnd 0.006979f
C2906 vdd.n1327 gnd 0.006979f
C2907 vdd.n1328 gnd 0.006979f
C2908 vdd.n1329 gnd 0.006979f
C2909 vdd.n1330 gnd 0.225494f
C2910 vdd.n1331 gnd 0.006979f
C2911 vdd.n1332 gnd 0.006979f
C2912 vdd.n1333 gnd 0.006979f
C2913 vdd.n1334 gnd 0.006979f
C2914 vdd.n1335 gnd 0.006979f
C2915 vdd.n1336 gnd 0.006979f
C2916 vdd.n1337 gnd 0.006979f
C2917 vdd.n1338 gnd 0.006979f
C2918 vdd.n1339 gnd 0.006979f
C2919 vdd.n1340 gnd 0.006979f
C2920 vdd.n1341 gnd 0.006979f
C2921 vdd.n1342 gnd 0.006979f
C2922 vdd.n1343 gnd 0.006979f
C2923 vdd.n1344 gnd 0.006979f
C2924 vdd.n1345 gnd 0.006979f
C2925 vdd.n1346 gnd 0.006979f
C2926 vdd.n1347 gnd 0.006979f
C2927 vdd.n1348 gnd 0.006979f
C2928 vdd.n1349 gnd 0.006979f
C2929 vdd.n1350 gnd 0.006979f
C2930 vdd.n1351 gnd 0.006979f
C2931 vdd.n1352 gnd 0.006979f
C2932 vdd.n1353 gnd 0.006979f
C2933 vdd.n1354 gnd 0.006979f
C2934 vdd.n1355 gnd 0.006979f
C2935 vdd.n1356 gnd 0.006979f
C2936 vdd.n1357 gnd 0.006979f
C2937 vdd.n1358 gnd 0.015287f
C2938 vdd.n1359 gnd 0.015287f
C2939 vdd.n1360 gnd 0.016323f
C2940 vdd.n1361 gnd 0.006979f
C2941 vdd.n1362 gnd 0.006979f
C2942 vdd.n1363 gnd 0.005388f
C2943 vdd.n1364 gnd 0.006979f
C2944 vdd.n1365 gnd 0.006979f
C2945 vdd.n1366 gnd 0.00508f
C2946 vdd.n1367 gnd 0.006979f
C2947 vdd.n1368 gnd 0.006979f
C2948 vdd.n1369 gnd 0.006979f
C2949 vdd.n1370 gnd 0.006979f
C2950 vdd.n1371 gnd 0.006979f
C2951 vdd.n1372 gnd 0.006979f
C2952 vdd.n1373 gnd 0.006979f
C2953 vdd.n1374 gnd 0.006979f
C2954 vdd.n1375 gnd 0.006979f
C2955 vdd.n1376 gnd 0.006979f
C2956 vdd.n1377 gnd 0.006979f
C2957 vdd.n1378 gnd 0.006979f
C2958 vdd.n1379 gnd 0.006979f
C2959 vdd.n1380 gnd 0.006979f
C2960 vdd.n1381 gnd 0.006979f
C2961 vdd.n1382 gnd 0.006979f
C2962 vdd.n1383 gnd 0.006979f
C2963 vdd.n1384 gnd 0.006979f
C2964 vdd.n1385 gnd 0.006979f
C2965 vdd.n1386 gnd 0.006979f
C2966 vdd.n1387 gnd 0.006979f
C2967 vdd.n1388 gnd 0.006979f
C2968 vdd.n1389 gnd 0.006979f
C2969 vdd.n1390 gnd 0.006979f
C2970 vdd.n1391 gnd 0.006979f
C2971 vdd.n1392 gnd 0.006979f
C2972 vdd.n1393 gnd 0.02797f
C2973 vdd.n1395 gnd 0.02353f
C2974 vdd.n1396 gnd 0.00826f
C2975 vdd.n1398 gnd 0.010263f
C2976 vdd.n1399 gnd 0.00826f
C2977 vdd.n1400 gnd 0.010263f
C2978 vdd.n1402 gnd 0.010263f
C2979 vdd.n1403 gnd 0.010263f
C2980 vdd.n1405 gnd 0.010263f
C2981 vdd.n1406 gnd 0.006856f
C2982 vdd.n1407 gnd 0.582088f
C2983 vdd.n1408 gnd 0.010263f
C2984 vdd.n1409 gnd 0.02353f
C2985 vdd.n1410 gnd 0.00826f
C2986 vdd.n1411 gnd 0.010263f
C2987 vdd.n1412 gnd 0.00826f
C2988 vdd.n1413 gnd 0.010263f
C2989 vdd.n1414 gnd 1.04881f
C2990 vdd.n1415 gnd 0.010263f
C2991 vdd.n1416 gnd 0.00826f
C2992 vdd.n1417 gnd 0.00826f
C2993 vdd.n1418 gnd 0.010263f
C2994 vdd.n1419 gnd 0.00826f
C2995 vdd.n1420 gnd 0.010263f
C2996 vdd.t172 gnd 0.524404f
C2997 vdd.n1421 gnd 0.010263f
C2998 vdd.n1422 gnd 0.00826f
C2999 vdd.n1423 gnd 0.010263f
C3000 vdd.n1424 gnd 0.00826f
C3001 vdd.n1425 gnd 0.010263f
C3002 vdd.t140 gnd 0.524404f
C3003 vdd.n1426 gnd 0.010263f
C3004 vdd.n1427 gnd 0.00826f
C3005 vdd.n1428 gnd 0.010263f
C3006 vdd.n1429 gnd 0.00826f
C3007 vdd.n1430 gnd 0.010263f
C3008 vdd.t199 gnd 0.524404f
C3009 vdd.n1431 gnd 0.728921f
C3010 vdd.n1432 gnd 0.010263f
C3011 vdd.n1433 gnd 0.00826f
C3012 vdd.n1434 gnd 0.010263f
C3013 vdd.n1435 gnd 0.00826f
C3014 vdd.n1436 gnd 0.010263f
C3015 vdd.n1437 gnd 0.833802f
C3016 vdd.n1438 gnd 0.010263f
C3017 vdd.n1439 gnd 0.00826f
C3018 vdd.n1440 gnd 0.010263f
C3019 vdd.n1441 gnd 0.00826f
C3020 vdd.n1442 gnd 0.010263f
C3021 vdd.n1443 gnd 0.655505f
C3022 vdd.t218 gnd 0.524404f
C3023 vdd.n1444 gnd 0.010263f
C3024 vdd.n1445 gnd 0.00826f
C3025 vdd.n1446 gnd 0.010263f
C3026 vdd.n1447 gnd 0.00826f
C3027 vdd.n1448 gnd 0.010263f
C3028 vdd.t191 gnd 0.524404f
C3029 vdd.n1449 gnd 0.010263f
C3030 vdd.n1450 gnd 0.00826f
C3031 vdd.n1451 gnd 0.010263f
C3032 vdd.n1452 gnd 0.00826f
C3033 vdd.n1453 gnd 0.010263f
C3034 vdd.t156 gnd 0.524404f
C3035 vdd.n1454 gnd 0.5716f
C3036 vdd.n1455 gnd 0.010263f
C3037 vdd.n1456 gnd 0.00826f
C3038 vdd.n1457 gnd 0.010263f
C3039 vdd.n1458 gnd 0.00826f
C3040 vdd.n1459 gnd 0.010263f
C3041 vdd.t174 gnd 0.524404f
C3042 vdd.n1460 gnd 0.010263f
C3043 vdd.n1461 gnd 0.00826f
C3044 vdd.n1462 gnd 0.010263f
C3045 vdd.n1463 gnd 0.00826f
C3046 vdd.n1464 gnd 0.010263f
C3047 vdd.n1465 gnd 0.812826f
C3048 vdd.n1466 gnd 0.87051f
C3049 vdd.t213 gnd 0.524404f
C3050 vdd.n1467 gnd 0.010263f
C3051 vdd.n1468 gnd 0.00826f
C3052 vdd.n1469 gnd 0.010263f
C3053 vdd.n1470 gnd 0.00826f
C3054 vdd.n1471 gnd 0.010263f
C3055 vdd.n1472 gnd 0.634528f
C3056 vdd.n1473 gnd 0.010263f
C3057 vdd.n1474 gnd 0.00826f
C3058 vdd.n1475 gnd 0.010263f
C3059 vdd.n1476 gnd 0.00826f
C3060 vdd.n1477 gnd 0.010263f
C3061 vdd.t168 gnd 0.524404f
C3062 vdd.t146 gnd 0.524404f
C3063 vdd.n1478 gnd 0.010263f
C3064 vdd.n1479 gnd 0.00826f
C3065 vdd.n1480 gnd 0.010263f
C3066 vdd.n1481 gnd 0.00826f
C3067 vdd.n1482 gnd 0.010263f
C3068 vdd.t170 gnd 0.524404f
C3069 vdd.n1483 gnd 0.010263f
C3070 vdd.n1484 gnd 0.00826f
C3071 vdd.n1485 gnd 0.010263f
C3072 vdd.n1486 gnd 0.00826f
C3073 vdd.n1487 gnd 0.010263f
C3074 vdd.t138 gnd 0.524404f
C3075 vdd.n1488 gnd 0.770873f
C3076 vdd.n1489 gnd 0.010263f
C3077 vdd.n1490 gnd 0.00826f
C3078 vdd.n1491 gnd 0.010263f
C3079 vdd.n1492 gnd 0.00826f
C3080 vdd.n1493 gnd 0.010263f
C3081 vdd.n1494 gnd 1.04881f
C3082 vdd.n1495 gnd 0.010263f
C3083 vdd.n1496 gnd 0.00826f
C3084 vdd.n1497 gnd 0.010263f
C3085 vdd.n1498 gnd 0.00826f
C3086 vdd.n1499 gnd 0.010263f
C3087 vdd.n1500 gnd 0.886242f
C3088 vdd.n1501 gnd 0.010263f
C3089 vdd.n1502 gnd 0.00826f
C3090 vdd.n1503 gnd 0.023371f
C3091 vdd.n1504 gnd 0.006856f
C3092 vdd.n1505 gnd 0.023371f
C3093 vdd.n1506 gnd 1.38443f
C3094 vdd.n1507 gnd 0.023371f
C3095 vdd.n1508 gnd 0.006856f
C3096 vdd.n1509 gnd 0.010263f
C3097 vdd.t87 gnd 0.126259f
C3098 vdd.t88 gnd 0.134936f
C3099 vdd.t86 gnd 0.164893f
C3100 vdd.n1510 gnd 0.211369f
C3101 vdd.n1511 gnd 0.178414f
C3102 vdd.n1512 gnd 0.013547f
C3103 vdd.n1513 gnd 0.010263f
C3104 vdd.n1544 gnd 0.010263f
C3105 vdd.n1545 gnd 0.010263f
C3106 vdd.n1546 gnd 0.02353f
C3107 vdd.n1547 gnd 0.00826f
C3108 vdd.n1548 gnd 0.010263f
C3109 vdd.n1549 gnd 0.010263f
C3110 vdd.n1550 gnd 0.010263f
C3111 vdd.n1551 gnd 0.010263f
C3112 vdd.n1552 gnd 0.00826f
C3113 vdd.n1553 gnd 0.010263f
C3114 vdd.n1554 gnd 0.010263f
C3115 vdd.n1555 gnd 0.010263f
C3116 vdd.n1556 gnd 0.010263f
C3117 vdd.n1557 gnd 0.010263f
C3118 vdd.n1558 gnd 0.00826f
C3119 vdd.n1559 gnd 0.010263f
C3120 vdd.n1560 gnd 0.010263f
C3121 vdd.n1561 gnd 0.010263f
C3122 vdd.n1562 gnd 0.010263f
C3123 vdd.n1563 gnd 0.010263f
C3124 vdd.n1564 gnd 0.00826f
C3125 vdd.n1565 gnd 0.010263f
C3126 vdd.n1566 gnd 0.010263f
C3127 vdd.n1567 gnd 0.010263f
C3128 vdd.n1568 gnd 0.010263f
C3129 vdd.n1569 gnd 0.010263f
C3130 vdd.n1570 gnd 0.006897f
C3131 vdd.n1571 gnd 0.010263f
C3132 vdd.n1572 gnd 0.010263f
C3133 vdd.n1573 gnd 0.010263f
C3134 vdd.n1574 gnd 0.00826f
C3135 vdd.n1575 gnd 0.010263f
C3136 vdd.n1576 gnd 0.010263f
C3137 vdd.n1577 gnd 0.010263f
C3138 vdd.n1578 gnd 0.010263f
C3139 vdd.n1579 gnd 0.010263f
C3140 vdd.n1580 gnd 0.00826f
C3141 vdd.n1581 gnd 0.010263f
C3142 vdd.n1582 gnd 0.010263f
C3143 vdd.n1583 gnd 0.010263f
C3144 vdd.n1584 gnd 0.010263f
C3145 vdd.n1585 gnd 0.010263f
C3146 vdd.n1586 gnd 0.00826f
C3147 vdd.n1587 gnd 0.010263f
C3148 vdd.n1588 gnd 0.010263f
C3149 vdd.n1589 gnd 0.010263f
C3150 vdd.n1590 gnd 0.010263f
C3151 vdd.n1591 gnd 0.010263f
C3152 vdd.n1592 gnd 0.00826f
C3153 vdd.n1593 gnd 0.010263f
C3154 vdd.n1594 gnd 0.010263f
C3155 vdd.n1595 gnd 0.010263f
C3156 vdd.n1596 gnd 0.010263f
C3157 vdd.n1597 gnd 0.010263f
C3158 vdd.n1598 gnd 0.00826f
C3159 vdd.n1599 gnd 0.010263f
C3160 vdd.n1600 gnd 0.010263f
C3161 vdd.n1601 gnd 0.010263f
C3162 vdd.n1602 gnd 0.010263f
C3163 vdd.n1603 gnd 0.008178f
C3164 vdd.n1604 gnd 0.010263f
C3165 vdd.n1605 gnd 0.010263f
C3166 vdd.n1606 gnd 0.010263f
C3167 vdd.n1607 gnd 0.010263f
C3168 vdd.n1608 gnd 0.010263f
C3169 vdd.n1609 gnd 0.00826f
C3170 vdd.n1610 gnd 0.010263f
C3171 vdd.n1611 gnd 0.010263f
C3172 vdd.n1612 gnd 0.010263f
C3173 vdd.n1613 gnd 0.010263f
C3174 vdd.n1614 gnd 0.010263f
C3175 vdd.n1615 gnd 0.00826f
C3176 vdd.n1616 gnd 0.010263f
C3177 vdd.n1617 gnd 0.010263f
C3178 vdd.n1618 gnd 0.010263f
C3179 vdd.n1619 gnd 0.010263f
C3180 vdd.n1620 gnd 0.010263f
C3181 vdd.n1621 gnd 0.00826f
C3182 vdd.n1622 gnd 0.010263f
C3183 vdd.n1623 gnd 0.010263f
C3184 vdd.n1624 gnd 0.010263f
C3185 vdd.n1625 gnd 0.010263f
C3186 vdd.n1626 gnd 0.010263f
C3187 vdd.n1627 gnd 0.00826f
C3188 vdd.n1628 gnd 0.010263f
C3189 vdd.n1629 gnd 0.010263f
C3190 vdd.n1630 gnd 0.010263f
C3191 vdd.n1631 gnd 0.010263f
C3192 vdd.n1632 gnd 0.010263f
C3193 vdd.n1633 gnd 0.004337f
C3194 vdd.n1634 gnd 0.010263f
C3195 vdd.n1635 gnd 0.00826f
C3196 vdd.n1636 gnd 0.00826f
C3197 vdd.n1637 gnd 0.00826f
C3198 vdd.n1638 gnd 0.010263f
C3199 vdd.n1639 gnd 0.010263f
C3200 vdd.n1640 gnd 0.010263f
C3201 vdd.n1641 gnd 0.00826f
C3202 vdd.n1642 gnd 0.00826f
C3203 vdd.n1643 gnd 0.00826f
C3204 vdd.n1644 gnd 0.010263f
C3205 vdd.n1645 gnd 0.010263f
C3206 vdd.n1646 gnd 0.010263f
C3207 vdd.n1647 gnd 0.00826f
C3208 vdd.n1648 gnd 0.00826f
C3209 vdd.n1649 gnd 0.00826f
C3210 vdd.n1650 gnd 0.010263f
C3211 vdd.n1651 gnd 0.010263f
C3212 vdd.n1652 gnd 0.010263f
C3213 vdd.n1653 gnd 0.00826f
C3214 vdd.n1654 gnd 0.00826f
C3215 vdd.n1655 gnd 0.00826f
C3216 vdd.n1656 gnd 0.010263f
C3217 vdd.n1657 gnd 0.010263f
C3218 vdd.n1658 gnd 0.010263f
C3219 vdd.n1659 gnd 0.00826f
C3220 vdd.n1660 gnd 0.00826f
C3221 vdd.n1661 gnd 0.00826f
C3222 vdd.n1662 gnd 0.010263f
C3223 vdd.n1663 gnd 0.010263f
C3224 vdd.n1664 gnd 0.010263f
C3225 vdd.n1665 gnd 0.010263f
C3226 vdd.t80 gnd 0.126259f
C3227 vdd.t81 gnd 0.134936f
C3228 vdd.t78 gnd 0.164893f
C3229 vdd.n1666 gnd 0.211369f
C3230 vdd.n1667 gnd 0.178414f
C3231 vdd.n1668 gnd 0.017677f
C3232 vdd.n1669 gnd 0.005617f
C3233 vdd.n1670 gnd 0.00826f
C3234 vdd.n1671 gnd 0.010263f
C3235 vdd.n1672 gnd 0.010263f
C3236 vdd.n1673 gnd 0.010263f
C3237 vdd.n1674 gnd 0.00826f
C3238 vdd.n1675 gnd 0.00826f
C3239 vdd.n1676 gnd 0.00826f
C3240 vdd.n1677 gnd 0.010263f
C3241 vdd.n1678 gnd 0.010263f
C3242 vdd.n1679 gnd 0.010263f
C3243 vdd.n1680 gnd 0.00826f
C3244 vdd.n1681 gnd 0.00826f
C3245 vdd.n1682 gnd 0.00826f
C3246 vdd.n1683 gnd 0.010263f
C3247 vdd.n1684 gnd 0.010263f
C3248 vdd.n1685 gnd 0.010263f
C3249 vdd.n1686 gnd 0.00826f
C3250 vdd.n1687 gnd 0.00826f
C3251 vdd.n1688 gnd 0.00826f
C3252 vdd.n1689 gnd 0.010263f
C3253 vdd.n1690 gnd 0.010263f
C3254 vdd.n1691 gnd 0.010263f
C3255 vdd.n1692 gnd 0.00826f
C3256 vdd.n1693 gnd 0.00826f
C3257 vdd.n1694 gnd 0.00826f
C3258 vdd.n1695 gnd 0.010263f
C3259 vdd.n1696 gnd 0.010263f
C3260 vdd.n1697 gnd 0.010263f
C3261 vdd.n1698 gnd 0.00826f
C3262 vdd.n1699 gnd 0.006897f
C3263 vdd.n1700 gnd 0.010263f
C3264 vdd.n1701 gnd 0.010263f
C3265 vdd.t90 gnd 0.126259f
C3266 vdd.t91 gnd 0.134936f
C3267 vdd.t89 gnd 0.164893f
C3268 vdd.n1702 gnd 0.211369f
C3269 vdd.n1703 gnd 0.178414f
C3270 vdd.n1704 gnd 0.017677f
C3271 vdd.n1705 gnd 0.010263f
C3272 vdd.n1706 gnd 0.010263f
C3273 vdd.n1707 gnd 0.010263f
C3274 vdd.n1708 gnd 0.00826f
C3275 vdd.n1709 gnd 0.00826f
C3276 vdd.n1710 gnd 0.00826f
C3277 vdd.n1711 gnd 0.010263f
C3278 vdd.n1712 gnd 0.010263f
C3279 vdd.n1713 gnd 0.010263f
C3280 vdd.n1714 gnd 0.00826f
C3281 vdd.n1715 gnd 0.00826f
C3282 vdd.n1716 gnd 0.00826f
C3283 vdd.n1717 gnd 0.010263f
C3284 vdd.n1718 gnd 0.010263f
C3285 vdd.n1719 gnd 0.010263f
C3286 vdd.n1720 gnd 0.00826f
C3287 vdd.n1721 gnd 0.00826f
C3288 vdd.n1722 gnd 0.00826f
C3289 vdd.n1723 gnd 0.010263f
C3290 vdd.n1724 gnd 0.010263f
C3291 vdd.n1725 gnd 0.010263f
C3292 vdd.n1726 gnd 0.00826f
C3293 vdd.n1727 gnd 0.00826f
C3294 vdd.n1728 gnd 0.00826f
C3295 vdd.n1729 gnd 0.010263f
C3296 vdd.n1730 gnd 0.010263f
C3297 vdd.n1731 gnd 0.010263f
C3298 vdd.n1732 gnd 0.00826f
C3299 vdd.n1733 gnd 0.006856f
C3300 vdd.n1734 gnd 0.02353f
C3301 vdd.n1736 gnd 2.31786f
C3302 vdd.n1737 gnd 0.02353f
C3303 vdd.n1738 gnd 0.003924f
C3304 vdd.n1739 gnd 0.02353f
C3305 vdd.n1740 gnd 0.023371f
C3306 vdd.n1741 gnd 0.010263f
C3307 vdd.n1742 gnd 0.00826f
C3308 vdd.n1743 gnd 0.010263f
C3309 vdd.t79 gnd 0.524404f
C3310 vdd.n1744 gnd 0.686969f
C3311 vdd.n1745 gnd 0.010263f
C3312 vdd.n1746 gnd 0.00826f
C3313 vdd.n1747 gnd 0.010263f
C3314 vdd.n1748 gnd 0.010263f
C3315 vdd.n1749 gnd 0.010263f
C3316 vdd.n1750 gnd 0.00826f
C3317 vdd.n1751 gnd 0.010263f
C3318 vdd.n1752 gnd 1.04881f
C3319 vdd.n1753 gnd 0.010263f
C3320 vdd.n1754 gnd 0.00826f
C3321 vdd.n1755 gnd 0.010263f
C3322 vdd.n1756 gnd 0.010263f
C3323 vdd.n1757 gnd 0.010263f
C3324 vdd.n1758 gnd 0.00826f
C3325 vdd.n1759 gnd 0.010263f
C3326 vdd.n1760 gnd 0.87051f
C3327 vdd.t142 gnd 0.524404f
C3328 vdd.n1761 gnd 0.603064f
C3329 vdd.n1762 gnd 0.010263f
C3330 vdd.n1763 gnd 0.00826f
C3331 vdd.n1764 gnd 0.010263f
C3332 vdd.n1765 gnd 0.010263f
C3333 vdd.n1766 gnd 0.010263f
C3334 vdd.n1767 gnd 0.00826f
C3335 vdd.n1768 gnd 0.010263f
C3336 vdd.n1769 gnd 0.62404f
C3337 vdd.n1770 gnd 0.010263f
C3338 vdd.n1771 gnd 0.00826f
C3339 vdd.n1772 gnd 0.010263f
C3340 vdd.n1773 gnd 0.010263f
C3341 vdd.n1774 gnd 0.010263f
C3342 vdd.n1775 gnd 0.00826f
C3343 vdd.n1776 gnd 0.010263f
C3344 vdd.n1777 gnd 0.592576f
C3345 vdd.n1778 gnd 0.802338f
C3346 vdd.n1779 gnd 0.010263f
C3347 vdd.n1780 gnd 0.00826f
C3348 vdd.n1781 gnd 0.010263f
C3349 vdd.n1782 gnd 0.010263f
C3350 vdd.n1783 gnd 0.010263f
C3351 vdd.n1784 gnd 0.00826f
C3352 vdd.n1785 gnd 0.010263f
C3353 vdd.n1786 gnd 0.87051f
C3354 vdd.n1787 gnd 0.010263f
C3355 vdd.n1788 gnd 0.00826f
C3356 vdd.n1789 gnd 0.010263f
C3357 vdd.n1790 gnd 0.010263f
C3358 vdd.n1791 gnd 0.010263f
C3359 vdd.n1792 gnd 0.00826f
C3360 vdd.n1793 gnd 0.010263f
C3361 vdd.t215 gnd 0.524404f
C3362 vdd.n1794 gnd 0.760385f
C3363 vdd.n1795 gnd 0.010263f
C3364 vdd.n1796 gnd 0.00826f
C3365 vdd.n1797 gnd 0.010263f
C3366 vdd.n1798 gnd 0.010263f
C3367 vdd.n1799 gnd 0.010263f
C3368 vdd.n1800 gnd 0.00826f
C3369 vdd.n1801 gnd 0.010263f
C3370 vdd.n1802 gnd 0.582088f
C3371 vdd.n1803 gnd 0.010263f
C3372 vdd.n1804 gnd 0.00826f
C3373 vdd.n1805 gnd 0.010263f
C3374 vdd.n1806 gnd 0.010263f
C3375 vdd.n1807 gnd 0.010263f
C3376 vdd.n1808 gnd 0.00826f
C3377 vdd.n1809 gnd 0.010263f
C3378 vdd.n1810 gnd 0.749897f
C3379 vdd.n1811 gnd 0.645016f
C3380 vdd.n1812 gnd 0.010263f
C3381 vdd.n1813 gnd 0.00826f
C3382 vdd.n1814 gnd 0.007888f
C3383 vdd.n1815 gnd 0.005632f
C3384 vdd.n1816 gnd 0.005227f
C3385 vdd.n1817 gnd 0.002891f
C3386 vdd.n1818 gnd 0.006638f
C3387 vdd.n1819 gnd 0.002809f
C3388 vdd.n1820 gnd 0.002974f
C3389 vdd.n1821 gnd 0.005227f
C3390 vdd.n1822 gnd 0.002809f
C3391 vdd.n1823 gnd 0.006638f
C3392 vdd.n1824 gnd 0.002974f
C3393 vdd.n1825 gnd 0.005227f
C3394 vdd.n1826 gnd 0.002809f
C3395 vdd.n1827 gnd 0.004979f
C3396 vdd.n1828 gnd 0.004994f
C3397 vdd.t173 gnd 0.014262f
C3398 vdd.n1829 gnd 0.031732f
C3399 vdd.n1830 gnd 0.165142f
C3400 vdd.n1831 gnd 0.002809f
C3401 vdd.n1832 gnd 0.002974f
C3402 vdd.n1833 gnd 0.006638f
C3403 vdd.n1834 gnd 0.006638f
C3404 vdd.n1835 gnd 0.002974f
C3405 vdd.n1836 gnd 0.002809f
C3406 vdd.n1837 gnd 0.005227f
C3407 vdd.n1838 gnd 0.005227f
C3408 vdd.n1839 gnd 0.002809f
C3409 vdd.n1840 gnd 0.002974f
C3410 vdd.n1841 gnd 0.006638f
C3411 vdd.n1842 gnd 0.006638f
C3412 vdd.n1843 gnd 0.002974f
C3413 vdd.n1844 gnd 0.002809f
C3414 vdd.n1845 gnd 0.005227f
C3415 vdd.n1846 gnd 0.005227f
C3416 vdd.n1847 gnd 0.002809f
C3417 vdd.n1848 gnd 0.002974f
C3418 vdd.n1849 gnd 0.006638f
C3419 vdd.n1850 gnd 0.006638f
C3420 vdd.n1851 gnd 0.015694f
C3421 vdd.n1852 gnd 0.002891f
C3422 vdd.n1853 gnd 0.002809f
C3423 vdd.n1854 gnd 0.013509f
C3424 vdd.n1855 gnd 0.009431f
C3425 vdd.t200 gnd 0.033041f
C3426 vdd.t247 gnd 0.033041f
C3427 vdd.n1856 gnd 0.227082f
C3428 vdd.n1857 gnd 0.178565f
C3429 vdd.t219 gnd 0.033041f
C3430 vdd.t258 gnd 0.033041f
C3431 vdd.n1858 gnd 0.227082f
C3432 vdd.n1859 gnd 0.144101f
C3433 vdd.t192 gnd 0.033041f
C3434 vdd.t149 gnd 0.033041f
C3435 vdd.n1860 gnd 0.227082f
C3436 vdd.n1861 gnd 0.144101f
C3437 vdd.t211 gnd 0.033041f
C3438 vdd.t157 gnd 0.033041f
C3439 vdd.n1862 gnd 0.227082f
C3440 vdd.n1863 gnd 0.144101f
C3441 vdd.t250 gnd 0.033041f
C3442 vdd.t262 gnd 0.033041f
C3443 vdd.n1864 gnd 0.227082f
C3444 vdd.n1865 gnd 0.144101f
C3445 vdd.t230 gnd 0.033041f
C3446 vdd.t161 gnd 0.033041f
C3447 vdd.n1866 gnd 0.227082f
C3448 vdd.n1867 gnd 0.144101f
C3449 vdd.t221 gnd 0.033041f
C3450 vdd.t171 gnd 0.033041f
C3451 vdd.n1868 gnd 0.227082f
C3452 vdd.n1869 gnd 0.144101f
C3453 vdd.n1870 gnd 0.005632f
C3454 vdd.n1871 gnd 0.005227f
C3455 vdd.n1872 gnd 0.002891f
C3456 vdd.n1873 gnd 0.006638f
C3457 vdd.n1874 gnd 0.002809f
C3458 vdd.n1875 gnd 0.002974f
C3459 vdd.n1876 gnd 0.005227f
C3460 vdd.n1877 gnd 0.002809f
C3461 vdd.n1878 gnd 0.006638f
C3462 vdd.n1879 gnd 0.002974f
C3463 vdd.n1880 gnd 0.005227f
C3464 vdd.n1881 gnd 0.002809f
C3465 vdd.n1882 gnd 0.004979f
C3466 vdd.n1883 gnd 0.004994f
C3467 vdd.t196 gnd 0.014262f
C3468 vdd.n1884 gnd 0.031732f
C3469 vdd.n1885 gnd 0.165142f
C3470 vdd.n1886 gnd 0.002809f
C3471 vdd.n1887 gnd 0.002974f
C3472 vdd.n1888 gnd 0.006638f
C3473 vdd.n1889 gnd 0.006638f
C3474 vdd.n1890 gnd 0.002974f
C3475 vdd.n1891 gnd 0.002809f
C3476 vdd.n1892 gnd 0.005227f
C3477 vdd.n1893 gnd 0.005227f
C3478 vdd.n1894 gnd 0.002809f
C3479 vdd.n1895 gnd 0.002974f
C3480 vdd.n1896 gnd 0.006638f
C3481 vdd.n1897 gnd 0.006638f
C3482 vdd.n1898 gnd 0.002974f
C3483 vdd.n1899 gnd 0.002809f
C3484 vdd.n1900 gnd 0.005227f
C3485 vdd.n1901 gnd 0.005227f
C3486 vdd.n1902 gnd 0.002809f
C3487 vdd.n1903 gnd 0.002974f
C3488 vdd.n1904 gnd 0.006638f
C3489 vdd.n1905 gnd 0.006638f
C3490 vdd.n1906 gnd 0.015694f
C3491 vdd.n1907 gnd 0.002891f
C3492 vdd.n1908 gnd 0.002809f
C3493 vdd.n1909 gnd 0.013509f
C3494 vdd.n1910 gnd 0.009135f
C3495 vdd.n1911 gnd 0.107212f
C3496 vdd.n1912 gnd 0.005632f
C3497 vdd.n1913 gnd 0.005227f
C3498 vdd.n1914 gnd 0.002891f
C3499 vdd.n1915 gnd 0.006638f
C3500 vdd.n1916 gnd 0.002809f
C3501 vdd.n1917 gnd 0.002974f
C3502 vdd.n1918 gnd 0.005227f
C3503 vdd.n1919 gnd 0.002809f
C3504 vdd.n1920 gnd 0.006638f
C3505 vdd.n1921 gnd 0.002974f
C3506 vdd.n1922 gnd 0.005227f
C3507 vdd.n1923 gnd 0.002809f
C3508 vdd.n1924 gnd 0.004979f
C3509 vdd.n1925 gnd 0.004994f
C3510 vdd.t246 gnd 0.014262f
C3511 vdd.n1926 gnd 0.031732f
C3512 vdd.n1927 gnd 0.165142f
C3513 vdd.n1928 gnd 0.002809f
C3514 vdd.n1929 gnd 0.002974f
C3515 vdd.n1930 gnd 0.006638f
C3516 vdd.n1931 gnd 0.006638f
C3517 vdd.n1932 gnd 0.002974f
C3518 vdd.n1933 gnd 0.002809f
C3519 vdd.n1934 gnd 0.005227f
C3520 vdd.n1935 gnd 0.005227f
C3521 vdd.n1936 gnd 0.002809f
C3522 vdd.n1937 gnd 0.002974f
C3523 vdd.n1938 gnd 0.006638f
C3524 vdd.n1939 gnd 0.006638f
C3525 vdd.n1940 gnd 0.002974f
C3526 vdd.n1941 gnd 0.002809f
C3527 vdd.n1942 gnd 0.005227f
C3528 vdd.n1943 gnd 0.005227f
C3529 vdd.n1944 gnd 0.002809f
C3530 vdd.n1945 gnd 0.002974f
C3531 vdd.n1946 gnd 0.006638f
C3532 vdd.n1947 gnd 0.006638f
C3533 vdd.n1948 gnd 0.015694f
C3534 vdd.n1949 gnd 0.002891f
C3535 vdd.n1950 gnd 0.002809f
C3536 vdd.n1951 gnd 0.013509f
C3537 vdd.n1952 gnd 0.009431f
C3538 vdd.t208 gnd 0.033041f
C3539 vdd.t141 gnd 0.033041f
C3540 vdd.n1953 gnd 0.227082f
C3541 vdd.n1954 gnd 0.178565f
C3542 vdd.t255 gnd 0.033041f
C3543 vdd.t232 gnd 0.033041f
C3544 vdd.n1955 gnd 0.227082f
C3545 vdd.n1956 gnd 0.144101f
C3546 vdd.t226 gnd 0.033041f
C3547 vdd.t179 gnd 0.033041f
C3548 vdd.n1957 gnd 0.227082f
C3549 vdd.n1958 gnd 0.144101f
C3550 vdd.t175 gnd 0.033041f
C3551 vdd.t227 gnd 0.033041f
C3552 vdd.n1959 gnd 0.227082f
C3553 vdd.n1960 gnd 0.144101f
C3554 vdd.t216 gnd 0.033041f
C3555 vdd.t214 gnd 0.033041f
C3556 vdd.n1961 gnd 0.227082f
C3557 vdd.n1962 gnd 0.144101f
C3558 vdd.t169 gnd 0.033041f
C3559 vdd.t147 gnd 0.033041f
C3560 vdd.n1963 gnd 0.227082f
C3561 vdd.n1964 gnd 0.144101f
C3562 vdd.t139 gnd 0.033041f
C3563 vdd.t212 gnd 0.033041f
C3564 vdd.n1965 gnd 0.227082f
C3565 vdd.n1966 gnd 0.144101f
C3566 vdd.n1967 gnd 0.005632f
C3567 vdd.n1968 gnd 0.005227f
C3568 vdd.n1969 gnd 0.002891f
C3569 vdd.n1970 gnd 0.006638f
C3570 vdd.n1971 gnd 0.002809f
C3571 vdd.n1972 gnd 0.002974f
C3572 vdd.n1973 gnd 0.005227f
C3573 vdd.n1974 gnd 0.002809f
C3574 vdd.n1975 gnd 0.006638f
C3575 vdd.n1976 gnd 0.002974f
C3576 vdd.n1977 gnd 0.005227f
C3577 vdd.n1978 gnd 0.002809f
C3578 vdd.n1979 gnd 0.004979f
C3579 vdd.n1980 gnd 0.004994f
C3580 vdd.t143 gnd 0.014262f
C3581 vdd.n1981 gnd 0.031732f
C3582 vdd.n1982 gnd 0.165142f
C3583 vdd.n1983 gnd 0.002809f
C3584 vdd.n1984 gnd 0.002974f
C3585 vdd.n1985 gnd 0.006638f
C3586 vdd.n1986 gnd 0.006638f
C3587 vdd.n1987 gnd 0.002974f
C3588 vdd.n1988 gnd 0.002809f
C3589 vdd.n1989 gnd 0.005227f
C3590 vdd.n1990 gnd 0.005227f
C3591 vdd.n1991 gnd 0.002809f
C3592 vdd.n1992 gnd 0.002974f
C3593 vdd.n1993 gnd 0.006638f
C3594 vdd.n1994 gnd 0.006638f
C3595 vdd.n1995 gnd 0.002974f
C3596 vdd.n1996 gnd 0.002809f
C3597 vdd.n1997 gnd 0.005227f
C3598 vdd.n1998 gnd 0.005227f
C3599 vdd.n1999 gnd 0.002809f
C3600 vdd.n2000 gnd 0.002974f
C3601 vdd.n2001 gnd 0.006638f
C3602 vdd.n2002 gnd 0.006638f
C3603 vdd.n2003 gnd 0.015694f
C3604 vdd.n2004 gnd 0.002891f
C3605 vdd.n2005 gnd 0.002809f
C3606 vdd.n2006 gnd 0.013509f
C3607 vdd.n2007 gnd 0.009135f
C3608 vdd.n2008 gnd 0.06378f
C3609 vdd.n2009 gnd 0.229817f
C3610 vdd.n2010 gnd 0.005632f
C3611 vdd.n2011 gnd 0.005227f
C3612 vdd.n2012 gnd 0.002891f
C3613 vdd.n2013 gnd 0.006638f
C3614 vdd.n2014 gnd 0.002809f
C3615 vdd.n2015 gnd 0.002974f
C3616 vdd.n2016 gnd 0.005227f
C3617 vdd.n2017 gnd 0.002809f
C3618 vdd.n2018 gnd 0.006638f
C3619 vdd.n2019 gnd 0.002974f
C3620 vdd.n2020 gnd 0.005227f
C3621 vdd.n2021 gnd 0.002809f
C3622 vdd.n2022 gnd 0.004979f
C3623 vdd.n2023 gnd 0.004994f
C3624 vdd.t254 gnd 0.014262f
C3625 vdd.n2024 gnd 0.031732f
C3626 vdd.n2025 gnd 0.165142f
C3627 vdd.n2026 gnd 0.002809f
C3628 vdd.n2027 gnd 0.002974f
C3629 vdd.n2028 gnd 0.006638f
C3630 vdd.n2029 gnd 0.006638f
C3631 vdd.n2030 gnd 0.002974f
C3632 vdd.n2031 gnd 0.002809f
C3633 vdd.n2032 gnd 0.005227f
C3634 vdd.n2033 gnd 0.005227f
C3635 vdd.n2034 gnd 0.002809f
C3636 vdd.n2035 gnd 0.002974f
C3637 vdd.n2036 gnd 0.006638f
C3638 vdd.n2037 gnd 0.006638f
C3639 vdd.n2038 gnd 0.002974f
C3640 vdd.n2039 gnd 0.002809f
C3641 vdd.n2040 gnd 0.005227f
C3642 vdd.n2041 gnd 0.005227f
C3643 vdd.n2042 gnd 0.002809f
C3644 vdd.n2043 gnd 0.002974f
C3645 vdd.n2044 gnd 0.006638f
C3646 vdd.n2045 gnd 0.006638f
C3647 vdd.n2046 gnd 0.015694f
C3648 vdd.n2047 gnd 0.002891f
C3649 vdd.n2048 gnd 0.002809f
C3650 vdd.n2049 gnd 0.013509f
C3651 vdd.n2050 gnd 0.009431f
C3652 vdd.t217 gnd 0.033041f
C3653 vdd.t165 gnd 0.033041f
C3654 vdd.n2051 gnd 0.227082f
C3655 vdd.n2052 gnd 0.178565f
C3656 vdd.t263 gnd 0.033041f
C3657 vdd.t239 gnd 0.033041f
C3658 vdd.n2053 gnd 0.227082f
C3659 vdd.n2054 gnd 0.144101f
C3660 vdd.t237 gnd 0.033041f
C3661 vdd.t197 gnd 0.033041f
C3662 vdd.n2055 gnd 0.227082f
C3663 vdd.n2056 gnd 0.144101f
C3664 vdd.t193 gnd 0.033041f
C3665 vdd.t238 gnd 0.033041f
C3666 vdd.n2057 gnd 0.227082f
C3667 vdd.n2058 gnd 0.144101f
C3668 vdd.t225 gnd 0.033041f
C3669 vdd.t224 gnd 0.033041f
C3670 vdd.n2059 gnd 0.227082f
C3671 vdd.n2060 gnd 0.144101f
C3672 vdd.t190 gnd 0.033041f
C3673 vdd.t167 gnd 0.033041f
C3674 vdd.n2061 gnd 0.227082f
C3675 vdd.n2062 gnd 0.144101f
C3676 vdd.t163 gnd 0.033041f
C3677 vdd.t223 gnd 0.033041f
C3678 vdd.n2063 gnd 0.227082f
C3679 vdd.n2064 gnd 0.144101f
C3680 vdd.n2065 gnd 0.005632f
C3681 vdd.n2066 gnd 0.005227f
C3682 vdd.n2067 gnd 0.002891f
C3683 vdd.n2068 gnd 0.006638f
C3684 vdd.n2069 gnd 0.002809f
C3685 vdd.n2070 gnd 0.002974f
C3686 vdd.n2071 gnd 0.005227f
C3687 vdd.n2072 gnd 0.002809f
C3688 vdd.n2073 gnd 0.006638f
C3689 vdd.n2074 gnd 0.002974f
C3690 vdd.n2075 gnd 0.005227f
C3691 vdd.n2076 gnd 0.002809f
C3692 vdd.n2077 gnd 0.004979f
C3693 vdd.n2078 gnd 0.004994f
C3694 vdd.t166 gnd 0.014262f
C3695 vdd.n2079 gnd 0.031732f
C3696 vdd.n2080 gnd 0.165142f
C3697 vdd.n2081 gnd 0.002809f
C3698 vdd.n2082 gnd 0.002974f
C3699 vdd.n2083 gnd 0.006638f
C3700 vdd.n2084 gnd 0.006638f
C3701 vdd.n2085 gnd 0.002974f
C3702 vdd.n2086 gnd 0.002809f
C3703 vdd.n2087 gnd 0.005227f
C3704 vdd.n2088 gnd 0.005227f
C3705 vdd.n2089 gnd 0.002809f
C3706 vdd.n2090 gnd 0.002974f
C3707 vdd.n2091 gnd 0.006638f
C3708 vdd.n2092 gnd 0.006638f
C3709 vdd.n2093 gnd 0.002974f
C3710 vdd.n2094 gnd 0.002809f
C3711 vdd.n2095 gnd 0.005227f
C3712 vdd.n2096 gnd 0.005227f
C3713 vdd.n2097 gnd 0.002809f
C3714 vdd.n2098 gnd 0.002974f
C3715 vdd.n2099 gnd 0.006638f
C3716 vdd.n2100 gnd 0.006638f
C3717 vdd.n2101 gnd 0.015694f
C3718 vdd.n2102 gnd 0.002891f
C3719 vdd.n2103 gnd 0.002809f
C3720 vdd.n2104 gnd 0.013509f
C3721 vdd.n2105 gnd 0.009135f
C3722 vdd.n2106 gnd 0.06378f
C3723 vdd.n2107 gnd 0.257364f
C3724 vdd.n2108 gnd 2.57896f
C3725 vdd.n2109 gnd 0.605338f
C3726 vdd.n2110 gnd 0.007888f
C3727 vdd.n2111 gnd 0.010263f
C3728 vdd.n2112 gnd 0.00826f
C3729 vdd.n2113 gnd 0.010263f
C3730 vdd.n2114 gnd 0.823314f
C3731 vdd.n2115 gnd 0.010263f
C3732 vdd.n2116 gnd 0.00826f
C3733 vdd.n2117 gnd 0.010263f
C3734 vdd.n2118 gnd 0.010263f
C3735 vdd.n2119 gnd 0.010263f
C3736 vdd.n2120 gnd 0.00826f
C3737 vdd.n2121 gnd 0.010263f
C3738 vdd.t148 gnd 0.524404f
C3739 vdd.n2122 gnd 0.87051f
C3740 vdd.n2123 gnd 0.010263f
C3741 vdd.n2124 gnd 0.00826f
C3742 vdd.n2125 gnd 0.010263f
C3743 vdd.n2126 gnd 0.010263f
C3744 vdd.n2127 gnd 0.010263f
C3745 vdd.n2128 gnd 0.00826f
C3746 vdd.n2129 gnd 0.010263f
C3747 vdd.n2130 gnd 0.739409f
C3748 vdd.n2131 gnd 0.010263f
C3749 vdd.n2132 gnd 0.00826f
C3750 vdd.n2133 gnd 0.010263f
C3751 vdd.n2134 gnd 0.010263f
C3752 vdd.n2135 gnd 0.010263f
C3753 vdd.n2136 gnd 0.00826f
C3754 vdd.n2137 gnd 0.010263f
C3755 vdd.n2138 gnd 0.87051f
C3756 vdd.t231 gnd 0.524404f
C3757 vdd.n2139 gnd 0.561112f
C3758 vdd.n2140 gnd 0.010263f
C3759 vdd.n2141 gnd 0.00826f
C3760 vdd.n2142 gnd 0.010263f
C3761 vdd.n2143 gnd 0.010263f
C3762 vdd.n2144 gnd 0.010263f
C3763 vdd.n2145 gnd 0.00826f
C3764 vdd.n2146 gnd 0.010263f
C3765 vdd.n2147 gnd 0.665993f
C3766 vdd.n2148 gnd 0.010263f
C3767 vdd.n2149 gnd 0.00826f
C3768 vdd.n2150 gnd 0.010263f
C3769 vdd.n2151 gnd 0.010263f
C3770 vdd.n2152 gnd 0.010263f
C3771 vdd.n2153 gnd 0.00826f
C3772 vdd.n2154 gnd 0.010263f
C3773 vdd.n2155 gnd 0.550624f
C3774 vdd.n2156 gnd 0.84429f
C3775 vdd.n2157 gnd 0.010263f
C3776 vdd.n2158 gnd 0.00826f
C3777 vdd.n2159 gnd 0.010263f
C3778 vdd.n2160 gnd 0.010263f
C3779 vdd.n2161 gnd 0.010263f
C3780 vdd.n2162 gnd 0.00826f
C3781 vdd.n2163 gnd 0.010263f
C3782 vdd.n2164 gnd 1.02259f
C3783 vdd.n2165 gnd 0.010263f
C3784 vdd.n2166 gnd 0.00826f
C3785 vdd.n2167 gnd 0.010263f
C3786 vdd.n2168 gnd 0.010263f
C3787 vdd.n2169 gnd 0.023371f
C3788 vdd.n2170 gnd 0.010263f
C3789 vdd.n2171 gnd 0.010263f
C3790 vdd.n2172 gnd 0.00826f
C3791 vdd.n2173 gnd 0.010263f
C3792 vdd.t62 gnd 0.524404f
C3793 vdd.n2174 gnd 0.991123f
C3794 vdd.n2175 gnd 0.010263f
C3795 vdd.n2176 gnd 0.00826f
C3796 vdd.n2177 gnd 0.010263f
C3797 vdd.n2178 gnd 0.010263f
C3798 vdd.n2179 gnd 0.023371f
C3799 vdd.n2180 gnd 0.006856f
C3800 vdd.n2181 gnd 0.023371f
C3801 vdd.n2182 gnd 1.38443f
C3802 vdd.n2183 gnd 0.023371f
C3803 vdd.n2184 gnd 0.02353f
C3804 vdd.n2185 gnd 0.003924f
C3805 vdd.t64 gnd 0.126259f
C3806 vdd.t63 gnd 0.134936f
C3807 vdd.t61 gnd 0.164893f
C3808 vdd.n2186 gnd 0.211369f
C3809 vdd.n2187 gnd 0.177588f
C3810 vdd.n2188 gnd 0.012721f
C3811 vdd.n2189 gnd 0.004337f
C3812 vdd.n2190 gnd 0.008826f
C3813 vdd.n2191 gnd 0.776127f
C3814 vdd.n2193 gnd 0.00826f
C3815 vdd.n2194 gnd 0.00826f
C3816 vdd.n2195 gnd 0.010263f
C3817 vdd.n2197 gnd 0.010263f
C3818 vdd.n2198 gnd 0.010263f
C3819 vdd.n2199 gnd 0.00826f
C3820 vdd.n2200 gnd 0.00826f
C3821 vdd.n2201 gnd 0.00826f
C3822 vdd.n2202 gnd 0.010263f
C3823 vdd.n2204 gnd 0.010263f
C3824 vdd.n2205 gnd 0.010263f
C3825 vdd.n2206 gnd 0.00826f
C3826 vdd.n2207 gnd 0.00826f
C3827 vdd.n2208 gnd 0.00826f
C3828 vdd.n2209 gnd 0.010263f
C3829 vdd.n2211 gnd 0.010263f
C3830 vdd.n2212 gnd 0.010263f
C3831 vdd.n2213 gnd 0.00826f
C3832 vdd.n2214 gnd 0.00826f
C3833 vdd.n2215 gnd 0.00826f
C3834 vdd.n2216 gnd 0.010263f
C3835 vdd.n2218 gnd 0.010263f
C3836 vdd.n2219 gnd 0.010263f
C3837 vdd.n2220 gnd 0.00826f
C3838 vdd.n2221 gnd 0.010263f
C3839 vdd.n2222 gnd 0.010263f
C3840 vdd.n2223 gnd 0.010263f
C3841 vdd.n2224 gnd 0.016851f
C3842 vdd.n2225 gnd 0.005617f
C3843 vdd.n2226 gnd 0.00826f
C3844 vdd.n2227 gnd 0.010263f
C3845 vdd.n2229 gnd 0.010263f
C3846 vdd.n2230 gnd 0.010263f
C3847 vdd.n2231 gnd 0.00826f
C3848 vdd.n2232 gnd 0.00826f
C3849 vdd.n2233 gnd 0.00826f
C3850 vdd.n2234 gnd 0.010263f
C3851 vdd.n2236 gnd 0.010263f
C3852 vdd.n2237 gnd 0.010263f
C3853 vdd.n2238 gnd 0.00826f
C3854 vdd.n2239 gnd 0.00826f
C3855 vdd.n2240 gnd 0.00826f
C3856 vdd.n2241 gnd 0.010263f
C3857 vdd.n2243 gnd 0.010263f
C3858 vdd.n2244 gnd 0.010263f
C3859 vdd.n2245 gnd 0.00826f
C3860 vdd.n2246 gnd 0.00826f
C3861 vdd.n2247 gnd 0.00826f
C3862 vdd.n2248 gnd 0.010263f
C3863 vdd.n2250 gnd 0.010263f
C3864 vdd.n2251 gnd 0.010263f
C3865 vdd.n2252 gnd 0.00826f
C3866 vdd.n2253 gnd 0.00826f
C3867 vdd.n2254 gnd 0.00826f
C3868 vdd.n2255 gnd 0.010263f
C3869 vdd.n2257 gnd 0.010263f
C3870 vdd.n2258 gnd 0.010263f
C3871 vdd.n2259 gnd 0.00826f
C3872 vdd.n2260 gnd 0.010263f
C3873 vdd.n2261 gnd 0.010263f
C3874 vdd.n2262 gnd 0.010263f
C3875 vdd.n2263 gnd 0.016851f
C3876 vdd.n2264 gnd 0.006897f
C3877 vdd.n2265 gnd 0.00826f
C3878 vdd.n2266 gnd 0.010263f
C3879 vdd.n2268 gnd 0.010263f
C3880 vdd.n2269 gnd 0.010263f
C3881 vdd.n2270 gnd 0.00826f
C3882 vdd.n2271 gnd 0.00826f
C3883 vdd.n2272 gnd 0.00826f
C3884 vdd.n2273 gnd 0.010263f
C3885 vdd.n2275 gnd 0.010263f
C3886 vdd.n2276 gnd 0.010263f
C3887 vdd.n2277 gnd 0.00826f
C3888 vdd.n2278 gnd 0.00826f
C3889 vdd.n2279 gnd 0.00826f
C3890 vdd.n2280 gnd 0.010263f
C3891 vdd.n2282 gnd 0.010263f
C3892 vdd.n2283 gnd 0.010263f
C3893 vdd.n2284 gnd 0.00826f
C3894 vdd.n2285 gnd 0.00826f
C3895 vdd.n2286 gnd 0.00826f
C3896 vdd.n2287 gnd 0.010263f
C3897 vdd.n2289 gnd 0.010263f
C3898 vdd.n2290 gnd 0.00826f
C3899 vdd.n2291 gnd 0.00826f
C3900 vdd.n2292 gnd 0.010263f
C3901 vdd.n2294 gnd 0.010263f
C3902 vdd.n2295 gnd 0.010263f
C3903 vdd.n2296 gnd 0.00826f
C3904 vdd.n2297 gnd 0.008826f
C3905 vdd.n2298 gnd 0.776127f
C3906 vdd.n2299 gnd 0.02797f
C3907 vdd.n2300 gnd 0.006979f
C3908 vdd.n2301 gnd 0.006979f
C3909 vdd.n2302 gnd 0.006979f
C3910 vdd.n2303 gnd 0.006979f
C3911 vdd.n2304 gnd 0.006979f
C3912 vdd.n2305 gnd 0.006979f
C3913 vdd.n2306 gnd 0.006979f
C3914 vdd.n2307 gnd 0.006979f
C3915 vdd.n2308 gnd 0.006979f
C3916 vdd.n2309 gnd 0.006979f
C3917 vdd.n2310 gnd 0.006979f
C3918 vdd.n2311 gnd 0.006979f
C3919 vdd.n2312 gnd 0.006979f
C3920 vdd.n2313 gnd 0.006979f
C3921 vdd.n2314 gnd 0.006979f
C3922 vdd.n2315 gnd 0.006979f
C3923 vdd.n2316 gnd 0.006979f
C3924 vdd.n2317 gnd 0.006979f
C3925 vdd.n2318 gnd 0.006979f
C3926 vdd.n2319 gnd 0.006979f
C3927 vdd.n2320 gnd 0.006979f
C3928 vdd.n2321 gnd 0.006979f
C3929 vdd.n2322 gnd 0.006979f
C3930 vdd.n2323 gnd 0.006979f
C3931 vdd.n2324 gnd 0.006979f
C3932 vdd.n2325 gnd 0.006979f
C3933 vdd.n2326 gnd 0.006979f
C3934 vdd.n2327 gnd 0.006979f
C3935 vdd.n2328 gnd 0.006979f
C3936 vdd.n2329 gnd 0.006979f
C3937 vdd.n2330 gnd 0.006979f
C3938 vdd.n2331 gnd 0.016323f
C3939 vdd.n2332 gnd 0.016323f
C3940 vdd.n2334 gnd 8.94633f
C3941 vdd.n2336 gnd 0.016323f
C3942 vdd.n2337 gnd 0.016323f
C3943 vdd.n2338 gnd 0.015287f
C3944 vdd.n2339 gnd 0.006979f
C3945 vdd.n2340 gnd 0.006979f
C3946 vdd.n2341 gnd 0.713189f
C3947 vdd.n2342 gnd 0.006979f
C3948 vdd.n2343 gnd 0.006979f
C3949 vdd.n2344 gnd 0.006979f
C3950 vdd.n2345 gnd 0.006979f
C3951 vdd.n2346 gnd 0.006979f
C3952 vdd.n2347 gnd 0.603064f
C3953 vdd.n2348 gnd 0.006979f
C3954 vdd.n2349 gnd 0.006979f
C3955 vdd.n2350 gnd 0.006979f
C3956 vdd.n2351 gnd 0.006979f
C3957 vdd.n2352 gnd 0.006979f
C3958 vdd.n2353 gnd 0.713189f
C3959 vdd.n2354 gnd 0.006979f
C3960 vdd.n2355 gnd 0.006979f
C3961 vdd.n2356 gnd 0.006979f
C3962 vdd.n2357 gnd 0.006979f
C3963 vdd.n2358 gnd 0.006979f
C3964 vdd.n2359 gnd 0.697457f
C3965 vdd.n2360 gnd 0.006979f
C3966 vdd.n2361 gnd 0.006979f
C3967 vdd.n2362 gnd 0.006979f
C3968 vdd.n2363 gnd 0.006979f
C3969 vdd.n2364 gnd 0.006979f
C3970 vdd.n2365 gnd 0.713189f
C3971 vdd.n2366 gnd 0.006979f
C3972 vdd.n2367 gnd 0.006979f
C3973 vdd.n2368 gnd 0.006979f
C3974 vdd.n2369 gnd 0.006979f
C3975 vdd.n2370 gnd 0.006979f
C3976 vdd.n2371 gnd 0.5716f
C3977 vdd.n2372 gnd 0.006979f
C3978 vdd.n2373 gnd 0.006979f
C3979 vdd.n2374 gnd 0.005952f
C3980 vdd.n2375 gnd 0.020216f
C3981 vdd.n2376 gnd 0.004516f
C3982 vdd.n2377 gnd 0.006979f
C3983 vdd.n2378 gnd 0.414279f
C3984 vdd.n2379 gnd 0.006979f
C3985 vdd.n2380 gnd 0.006979f
C3986 vdd.n2381 gnd 0.006979f
C3987 vdd.n2382 gnd 0.006979f
C3988 vdd.n2383 gnd 0.006979f
C3989 vdd.n2384 gnd 0.456231f
C3990 vdd.n2385 gnd 0.006979f
C3991 vdd.n2386 gnd 0.006979f
C3992 vdd.n2387 gnd 0.006979f
C3993 vdd.n2388 gnd 0.006979f
C3994 vdd.n2389 gnd 0.006979f
C3995 vdd.n2390 gnd 0.613552f
C3996 vdd.n2391 gnd 0.006979f
C3997 vdd.n2392 gnd 0.006979f
C3998 vdd.n2393 gnd 0.006979f
C3999 vdd.n2394 gnd 0.006979f
C4000 vdd.n2395 gnd 0.006979f
C4001 vdd.n2396 gnd 0.587332f
C4002 vdd.n2397 gnd 0.006979f
C4003 vdd.n2398 gnd 0.006979f
C4004 vdd.n2399 gnd 0.006979f
C4005 vdd.n2400 gnd 0.006979f
C4006 vdd.n2401 gnd 0.006979f
C4007 vdd.n2402 gnd 0.430011f
C4008 vdd.n2403 gnd 0.006979f
C4009 vdd.n2404 gnd 0.006979f
C4010 vdd.n2405 gnd 0.006979f
C4011 vdd.n2406 gnd 0.006979f
C4012 vdd.n2407 gnd 0.006979f
C4013 vdd.n2408 gnd 0.225494f
C4014 vdd.n2409 gnd 0.006979f
C4015 vdd.n2410 gnd 0.006979f
C4016 vdd.n2411 gnd 0.006979f
C4017 vdd.n2412 gnd 0.006979f
C4018 vdd.n2413 gnd 0.006979f
C4019 vdd.n2414 gnd 0.372327f
C4020 vdd.n2415 gnd 0.006979f
C4021 vdd.n2416 gnd 0.006979f
C4022 vdd.n2417 gnd 0.006979f
C4023 vdd.n2418 gnd 0.006979f
C4024 vdd.n2419 gnd 0.006979f
C4025 vdd.n2420 gnd 0.713189f
C4026 vdd.n2421 gnd 0.006979f
C4027 vdd.n2422 gnd 0.006979f
C4028 vdd.n2423 gnd 0.006979f
C4029 vdd.n2424 gnd 0.006979f
C4030 vdd.n2425 gnd 0.006979f
C4031 vdd.n2426 gnd 0.006979f
C4032 vdd.n2427 gnd 0.006979f
C4033 vdd.n2428 gnd 0.534892f
C4034 vdd.n2429 gnd 0.006979f
C4035 vdd.n2430 gnd 0.006979f
C4036 vdd.n2431 gnd 0.006979f
C4037 vdd.n2432 gnd 0.006979f
C4038 vdd.n2433 gnd 0.006979f
C4039 vdd.n2434 gnd 0.006979f
C4040 vdd.n2435 gnd 0.445743f
C4041 vdd.n2436 gnd 0.006979f
C4042 vdd.n2437 gnd 0.006979f
C4043 vdd.n2438 gnd 0.006979f
C4044 vdd.n2439 gnd 0.016154f
C4045 vdd.n2440 gnd 0.015456f
C4046 vdd.n2441 gnd 0.006979f
C4047 vdd.n2442 gnd 0.006979f
C4048 vdd.n2443 gnd 0.005388f
C4049 vdd.n2444 gnd 0.006979f
C4050 vdd.n2445 gnd 0.006979f
C4051 vdd.n2446 gnd 0.00508f
C4052 vdd.n2447 gnd 0.006979f
C4053 vdd.n2448 gnd 0.006979f
C4054 vdd.n2449 gnd 0.006979f
C4055 vdd.n2450 gnd 0.006979f
C4056 vdd.n2451 gnd 0.006979f
C4057 vdd.n2452 gnd 0.006979f
C4058 vdd.n2453 gnd 0.006979f
C4059 vdd.n2454 gnd 0.006979f
C4060 vdd.n2455 gnd 0.006979f
C4061 vdd.n2456 gnd 0.006979f
C4062 vdd.n2457 gnd 0.006979f
C4063 vdd.n2458 gnd 0.006979f
C4064 vdd.n2459 gnd 0.006979f
C4065 vdd.n2460 gnd 0.006979f
C4066 vdd.n2461 gnd 0.006979f
C4067 vdd.n2462 gnd 0.006979f
C4068 vdd.n2463 gnd 0.006979f
C4069 vdd.n2464 gnd 0.006979f
C4070 vdd.n2465 gnd 0.006979f
C4071 vdd.n2466 gnd 0.006979f
C4072 vdd.n2467 gnd 0.006979f
C4073 vdd.n2468 gnd 0.006979f
C4074 vdd.n2469 gnd 0.006979f
C4075 vdd.n2470 gnd 0.006979f
C4076 vdd.n2471 gnd 0.006979f
C4077 vdd.n2472 gnd 0.006979f
C4078 vdd.n2473 gnd 0.006979f
C4079 vdd.n2474 gnd 0.006979f
C4080 vdd.n2475 gnd 0.006979f
C4081 vdd.n2476 gnd 0.006979f
C4082 vdd.n2477 gnd 0.006979f
C4083 vdd.n2478 gnd 0.006979f
C4084 vdd.n2479 gnd 0.006979f
C4085 vdd.n2480 gnd 0.006979f
C4086 vdd.n2481 gnd 0.006979f
C4087 vdd.n2482 gnd 0.006979f
C4088 vdd.n2483 gnd 0.006979f
C4089 vdd.n2484 gnd 0.006979f
C4090 vdd.n2485 gnd 0.006979f
C4091 vdd.n2486 gnd 0.006979f
C4092 vdd.n2487 gnd 0.006979f
C4093 vdd.n2488 gnd 0.006979f
C4094 vdd.n2489 gnd 0.006979f
C4095 vdd.n2490 gnd 0.006979f
C4096 vdd.n2491 gnd 0.006979f
C4097 vdd.n2492 gnd 0.006979f
C4098 vdd.n2493 gnd 0.006979f
C4099 vdd.n2494 gnd 0.006979f
C4100 vdd.n2495 gnd 0.006979f
C4101 vdd.n2496 gnd 0.006979f
C4102 vdd.n2497 gnd 0.006979f
C4103 vdd.n2498 gnd 0.006979f
C4104 vdd.n2499 gnd 0.006979f
C4105 vdd.n2500 gnd 0.006979f
C4106 vdd.n2501 gnd 0.006979f
C4107 vdd.n2502 gnd 0.006979f
C4108 vdd.n2503 gnd 0.006979f
C4109 vdd.n2504 gnd 0.006979f
C4110 vdd.n2505 gnd 0.006979f
C4111 vdd.n2506 gnd 0.006979f
C4112 vdd.n2507 gnd 0.016323f
C4113 vdd.n2508 gnd 0.015287f
C4114 vdd.n2509 gnd 0.015287f
C4115 vdd.n2510 gnd 0.849534f
C4116 vdd.n2511 gnd 0.015287f
C4117 vdd.n2512 gnd 0.016323f
C4118 vdd.n2513 gnd 0.015456f
C4119 vdd.n2514 gnd 0.006979f
C4120 vdd.n2515 gnd 0.006979f
C4121 vdd.n2516 gnd 0.006979f
C4122 vdd.n2517 gnd 0.005388f
C4123 vdd.n2518 gnd 0.009974f
C4124 vdd.n2519 gnd 0.00508f
C4125 vdd.n2520 gnd 0.006979f
C4126 vdd.n2521 gnd 0.006979f
C4127 vdd.n2522 gnd 0.006979f
C4128 vdd.n2523 gnd 0.006979f
C4129 vdd.n2524 gnd 0.006979f
C4130 vdd.n2525 gnd 0.006979f
C4131 vdd.n2526 gnd 0.006979f
C4132 vdd.n2527 gnd 0.006979f
C4133 vdd.n2528 gnd 0.006979f
C4134 vdd.n2529 gnd 0.006979f
C4135 vdd.n2530 gnd 0.006979f
C4136 vdd.n2531 gnd 0.006979f
C4137 vdd.n2532 gnd 0.006979f
C4138 vdd.n2533 gnd 0.006979f
C4139 vdd.n2534 gnd 0.006979f
C4140 vdd.n2535 gnd 0.006979f
C4141 vdd.n2536 gnd 0.006979f
C4142 vdd.n2537 gnd 0.006979f
C4143 vdd.n2538 gnd 0.006979f
C4144 vdd.n2539 gnd 0.006979f
C4145 vdd.n2540 gnd 0.006979f
C4146 vdd.n2541 gnd 0.006979f
C4147 vdd.n2542 gnd 0.006979f
C4148 vdd.n2543 gnd 0.006979f
C4149 vdd.n2544 gnd 0.006979f
C4150 vdd.n2545 gnd 0.006979f
C4151 vdd.n2546 gnd 0.006979f
C4152 vdd.n2547 gnd 0.006979f
C4153 vdd.n2548 gnd 0.006979f
C4154 vdd.n2549 gnd 0.006979f
C4155 vdd.n2550 gnd 0.006979f
C4156 vdd.n2551 gnd 0.006979f
C4157 vdd.n2552 gnd 0.006979f
C4158 vdd.n2553 gnd 0.006979f
C4159 vdd.n2554 gnd 0.006979f
C4160 vdd.n2555 gnd 0.006979f
C4161 vdd.n2556 gnd 0.006979f
C4162 vdd.n2557 gnd 0.006979f
C4163 vdd.n2558 gnd 0.006979f
C4164 vdd.n2559 gnd 0.006979f
C4165 vdd.n2560 gnd 0.006979f
C4166 vdd.n2561 gnd 0.006979f
C4167 vdd.n2562 gnd 0.006979f
C4168 vdd.n2563 gnd 0.006979f
C4169 vdd.n2564 gnd 0.006979f
C4170 vdd.n2565 gnd 0.006979f
C4171 vdd.n2566 gnd 0.006979f
C4172 vdd.n2567 gnd 0.006979f
C4173 vdd.n2568 gnd 0.006979f
C4174 vdd.n2569 gnd 0.006979f
C4175 vdd.n2570 gnd 0.006979f
C4176 vdd.n2571 gnd 0.006979f
C4177 vdd.n2572 gnd 0.006979f
C4178 vdd.n2573 gnd 0.006979f
C4179 vdd.n2574 gnd 0.006979f
C4180 vdd.n2575 gnd 0.006979f
C4181 vdd.n2576 gnd 0.006979f
C4182 vdd.n2577 gnd 0.006979f
C4183 vdd.n2578 gnd 0.006979f
C4184 vdd.n2579 gnd 0.006979f
C4185 vdd.n2580 gnd 0.016323f
C4186 vdd.n2581 gnd 0.016323f
C4187 vdd.n2582 gnd 0.87051f
C4188 vdd.t132 gnd 3.09398f
C4189 vdd.t266 gnd 3.09398f
C4190 vdd.n2615 gnd 0.016323f
C4191 vdd.t38 gnd 0.650261f
C4192 vdd.n2616 gnd 0.006979f
C4193 vdd.n2617 gnd 0.006979f
C4194 vdd.t101 gnd 0.282008f
C4195 vdd.t102 gnd 0.28867f
C4196 vdd.t99 gnd 0.184106f
C4197 vdd.n2618 gnd 0.099499f
C4198 vdd.n2619 gnd 0.056439f
C4199 vdd.n2620 gnd 0.006979f
C4200 vdd.t111 gnd 0.282008f
C4201 vdd.t112 gnd 0.28867f
C4202 vdd.t110 gnd 0.184106f
C4203 vdd.n2621 gnd 0.099499f
C4204 vdd.n2622 gnd 0.056439f
C4205 vdd.n2623 gnd 0.009974f
C4206 vdd.n2624 gnd 0.006979f
C4207 vdd.n2625 gnd 0.006979f
C4208 vdd.n2626 gnd 0.006979f
C4209 vdd.n2627 gnd 0.006979f
C4210 vdd.n2628 gnd 0.006979f
C4211 vdd.n2629 gnd 0.006979f
C4212 vdd.n2630 gnd 0.006979f
C4213 vdd.n2631 gnd 0.006979f
C4214 vdd.n2632 gnd 0.006979f
C4215 vdd.n2633 gnd 0.006979f
C4216 vdd.n2634 gnd 0.006979f
C4217 vdd.n2635 gnd 0.006979f
C4218 vdd.n2636 gnd 0.006979f
C4219 vdd.n2637 gnd 0.006979f
C4220 vdd.n2638 gnd 0.006979f
C4221 vdd.n2639 gnd 0.006979f
C4222 vdd.n2640 gnd 0.006979f
C4223 vdd.n2641 gnd 0.006979f
C4224 vdd.n2642 gnd 0.006979f
C4225 vdd.n2643 gnd 0.006979f
C4226 vdd.n2644 gnd 0.006979f
C4227 vdd.n2645 gnd 0.006979f
C4228 vdd.n2646 gnd 0.006979f
C4229 vdd.n2647 gnd 0.006979f
C4230 vdd.n2648 gnd 0.006979f
C4231 vdd.n2649 gnd 0.006979f
C4232 vdd.n2650 gnd 0.006979f
C4233 vdd.n2651 gnd 0.006979f
C4234 vdd.n2652 gnd 0.006979f
C4235 vdd.n2653 gnd 0.006979f
C4236 vdd.n2654 gnd 0.006979f
C4237 vdd.n2655 gnd 0.006979f
C4238 vdd.n2656 gnd 0.006979f
C4239 vdd.n2657 gnd 0.006979f
C4240 vdd.n2658 gnd 0.006979f
C4241 vdd.n2659 gnd 0.006979f
C4242 vdd.n2660 gnd 0.006979f
C4243 vdd.n2661 gnd 0.006979f
C4244 vdd.n2662 gnd 0.006979f
C4245 vdd.n2663 gnd 0.006979f
C4246 vdd.n2664 gnd 0.006979f
C4247 vdd.n2665 gnd 0.006979f
C4248 vdd.n2666 gnd 0.006979f
C4249 vdd.n2667 gnd 0.006979f
C4250 vdd.n2668 gnd 0.006979f
C4251 vdd.n2669 gnd 0.006979f
C4252 vdd.n2670 gnd 0.006979f
C4253 vdd.n2671 gnd 0.006979f
C4254 vdd.n2672 gnd 0.006979f
C4255 vdd.n2673 gnd 0.006979f
C4256 vdd.n2674 gnd 0.006979f
C4257 vdd.n2675 gnd 0.006979f
C4258 vdd.n2676 gnd 0.006979f
C4259 vdd.n2677 gnd 0.006979f
C4260 vdd.n2678 gnd 0.006979f
C4261 vdd.n2679 gnd 0.006979f
C4262 vdd.n2680 gnd 0.006979f
C4263 vdd.n2681 gnd 0.006979f
C4264 vdd.n2682 gnd 0.00508f
C4265 vdd.n2683 gnd 0.006979f
C4266 vdd.n2684 gnd 0.006979f
C4267 vdd.n2685 gnd 0.005388f
C4268 vdd.n2686 gnd 0.006979f
C4269 vdd.n2687 gnd 0.006979f
C4270 vdd.n2688 gnd 0.016323f
C4271 vdd.n2689 gnd 0.015287f
C4272 vdd.n2690 gnd 0.015287f
C4273 vdd.n2691 gnd 0.006979f
C4274 vdd.n2692 gnd 0.006979f
C4275 vdd.n2693 gnd 0.006979f
C4276 vdd.n2694 gnd 0.006979f
C4277 vdd.n2695 gnd 0.006979f
C4278 vdd.n2696 gnd 0.006979f
C4279 vdd.n2697 gnd 0.006979f
C4280 vdd.n2698 gnd 0.006979f
C4281 vdd.n2699 gnd 0.006979f
C4282 vdd.n2700 gnd 0.006979f
C4283 vdd.n2701 gnd 0.006979f
C4284 vdd.n2702 gnd 0.006979f
C4285 vdd.n2703 gnd 0.006979f
C4286 vdd.n2704 gnd 0.006979f
C4287 vdd.n2705 gnd 0.006979f
C4288 vdd.n2706 gnd 0.006979f
C4289 vdd.n2707 gnd 0.006979f
C4290 vdd.n2708 gnd 0.006979f
C4291 vdd.n2709 gnd 0.006979f
C4292 vdd.n2710 gnd 0.006979f
C4293 vdd.n2711 gnd 0.006979f
C4294 vdd.n2712 gnd 0.006979f
C4295 vdd.n2713 gnd 0.006979f
C4296 vdd.n2714 gnd 0.006979f
C4297 vdd.n2715 gnd 0.006979f
C4298 vdd.n2716 gnd 0.006979f
C4299 vdd.n2717 gnd 0.006979f
C4300 vdd.n2718 gnd 0.006979f
C4301 vdd.n2719 gnd 0.006979f
C4302 vdd.n2720 gnd 0.006979f
C4303 vdd.n2721 gnd 0.006979f
C4304 vdd.n2722 gnd 0.006979f
C4305 vdd.n2723 gnd 0.006979f
C4306 vdd.n2724 gnd 0.006979f
C4307 vdd.n2725 gnd 0.006979f
C4308 vdd.n2726 gnd 0.006979f
C4309 vdd.n2727 gnd 0.006979f
C4310 vdd.n2728 gnd 0.006979f
C4311 vdd.n2729 gnd 0.006979f
C4312 vdd.n2730 gnd 0.006979f
C4313 vdd.n2731 gnd 0.006979f
C4314 vdd.n2732 gnd 0.006979f
C4315 vdd.n2733 gnd 0.006979f
C4316 vdd.n2734 gnd 0.006979f
C4317 vdd.n2735 gnd 0.006979f
C4318 vdd.n2736 gnd 0.006979f
C4319 vdd.n2737 gnd 0.006979f
C4320 vdd.n2738 gnd 0.006979f
C4321 vdd.n2739 gnd 0.006979f
C4322 vdd.n2740 gnd 0.006979f
C4323 vdd.n2741 gnd 0.006979f
C4324 vdd.n2742 gnd 0.006979f
C4325 vdd.n2743 gnd 0.006979f
C4326 vdd.n2744 gnd 0.006979f
C4327 vdd.n2745 gnd 0.006979f
C4328 vdd.n2746 gnd 0.006979f
C4329 vdd.n2747 gnd 0.006979f
C4330 vdd.n2748 gnd 0.006979f
C4331 vdd.n2749 gnd 0.006979f
C4332 vdd.n2750 gnd 0.006979f
C4333 vdd.n2751 gnd 0.006979f
C4334 vdd.n2752 gnd 0.006979f
C4335 vdd.n2753 gnd 0.006979f
C4336 vdd.n2754 gnd 0.006979f
C4337 vdd.n2755 gnd 0.006979f
C4338 vdd.n2756 gnd 0.006979f
C4339 vdd.n2757 gnd 0.006979f
C4340 vdd.n2758 gnd 0.006979f
C4341 vdd.n2759 gnd 0.006979f
C4342 vdd.n2760 gnd 0.006979f
C4343 vdd.n2761 gnd 0.006979f
C4344 vdd.n2762 gnd 0.006979f
C4345 vdd.n2763 gnd 0.006979f
C4346 vdd.n2764 gnd 0.225494f
C4347 vdd.n2765 gnd 0.006979f
C4348 vdd.n2766 gnd 0.006979f
C4349 vdd.n2767 gnd 0.006979f
C4350 vdd.n2768 gnd 0.006979f
C4351 vdd.n2769 gnd 0.006979f
C4352 vdd.n2770 gnd 0.006979f
C4353 vdd.n2771 gnd 0.006979f
C4354 vdd.n2772 gnd 0.006979f
C4355 vdd.n2773 gnd 0.006979f
C4356 vdd.n2774 gnd 0.006979f
C4357 vdd.n2775 gnd 0.006979f
C4358 vdd.n2776 gnd 0.006979f
C4359 vdd.n2777 gnd 0.006979f
C4360 vdd.n2778 gnd 0.006979f
C4361 vdd.n2779 gnd 0.445743f
C4362 vdd.n2780 gnd 0.006979f
C4363 vdd.n2781 gnd 0.006979f
C4364 vdd.n2782 gnd 0.006979f
C4365 vdd.n2783 gnd 0.015287f
C4366 vdd.n2784 gnd 0.015287f
C4367 vdd.n2785 gnd 0.016323f
C4368 vdd.n2786 gnd 0.016323f
C4369 vdd.n2787 gnd 0.006979f
C4370 vdd.n2788 gnd 0.006979f
C4371 vdd.n2789 gnd 0.006979f
C4372 vdd.n2790 gnd 0.005388f
C4373 vdd.n2791 gnd 0.009974f
C4374 vdd.n2792 gnd 0.00508f
C4375 vdd.n2793 gnd 0.006979f
C4376 vdd.n2794 gnd 0.006979f
C4377 vdd.n2795 gnd 0.006979f
C4378 vdd.n2796 gnd 0.006979f
C4379 vdd.n2797 gnd 0.006979f
C4380 vdd.n2798 gnd 0.006979f
C4381 vdd.n2799 gnd 0.006979f
C4382 vdd.n2800 gnd 0.006979f
C4383 vdd.n2801 gnd 0.006979f
C4384 vdd.n2802 gnd 0.006979f
C4385 vdd.n2803 gnd 0.006979f
C4386 vdd.n2804 gnd 0.006979f
C4387 vdd.n2805 gnd 0.006979f
C4388 vdd.n2806 gnd 0.006979f
C4389 vdd.n2807 gnd 0.006979f
C4390 vdd.n2808 gnd 0.006979f
C4391 vdd.n2809 gnd 0.006979f
C4392 vdd.n2810 gnd 0.006979f
C4393 vdd.n2811 gnd 0.006979f
C4394 vdd.n2812 gnd 0.006979f
C4395 vdd.n2813 gnd 0.006979f
C4396 vdd.n2814 gnd 0.006979f
C4397 vdd.n2815 gnd 0.006979f
C4398 vdd.n2816 gnd 0.006979f
C4399 vdd.n2817 gnd 0.006979f
C4400 vdd.n2818 gnd 0.006979f
C4401 vdd.n2819 gnd 0.006979f
C4402 vdd.n2820 gnd 0.006979f
C4403 vdd.n2821 gnd 0.006979f
C4404 vdd.n2822 gnd 0.006979f
C4405 vdd.n2823 gnd 0.006979f
C4406 vdd.n2824 gnd 0.006979f
C4407 vdd.n2825 gnd 0.006979f
C4408 vdd.n2826 gnd 0.006979f
C4409 vdd.n2827 gnd 0.006979f
C4410 vdd.n2828 gnd 0.006979f
C4411 vdd.n2829 gnd 0.006979f
C4412 vdd.n2830 gnd 0.006979f
C4413 vdd.n2831 gnd 0.006979f
C4414 vdd.n2832 gnd 0.006979f
C4415 vdd.n2833 gnd 0.006979f
C4416 vdd.n2834 gnd 0.006979f
C4417 vdd.n2835 gnd 0.006979f
C4418 vdd.n2836 gnd 0.006979f
C4419 vdd.n2837 gnd 0.006979f
C4420 vdd.n2838 gnd 0.006979f
C4421 vdd.n2839 gnd 0.006979f
C4422 vdd.n2840 gnd 0.006979f
C4423 vdd.n2841 gnd 0.006979f
C4424 vdd.n2842 gnd 0.006979f
C4425 vdd.n2843 gnd 0.006979f
C4426 vdd.n2844 gnd 0.006979f
C4427 vdd.n2845 gnd 0.006979f
C4428 vdd.n2846 gnd 0.006979f
C4429 vdd.n2847 gnd 0.006979f
C4430 vdd.n2848 gnd 0.006979f
C4431 vdd.n2849 gnd 0.006979f
C4432 vdd.n2850 gnd 0.006979f
C4433 vdd.n2851 gnd 0.006979f
C4434 vdd.n2852 gnd 0.016323f
C4435 vdd.n2853 gnd 0.016323f
C4436 vdd.n2855 gnd 0.87051f
C4437 vdd.n2857 gnd 0.016323f
C4438 vdd.n2858 gnd 0.016323f
C4439 vdd.n2859 gnd 0.015287f
C4440 vdd.n2860 gnd 0.006979f
C4441 vdd.n2861 gnd 0.006979f
C4442 vdd.n2862 gnd 0.377571f
C4443 vdd.n2863 gnd 0.006979f
C4444 vdd.n2864 gnd 0.006979f
C4445 vdd.n2865 gnd 0.006979f
C4446 vdd.n2866 gnd 0.006979f
C4447 vdd.n2867 gnd 0.006979f
C4448 vdd.n2868 gnd 0.424767f
C4449 vdd.n2869 gnd 0.006979f
C4450 vdd.n2870 gnd 0.006979f
C4451 vdd.n2871 gnd 0.006979f
C4452 vdd.n2872 gnd 0.006979f
C4453 vdd.n2873 gnd 0.006979f
C4454 vdd.n2874 gnd 0.713189f
C4455 vdd.n2875 gnd 0.006979f
C4456 vdd.n2876 gnd 0.006979f
C4457 vdd.n2877 gnd 0.006979f
C4458 vdd.n2878 gnd 0.006979f
C4459 vdd.n2879 gnd 0.006979f
C4460 vdd.n2880 gnd 0.471963f
C4461 vdd.n2881 gnd 0.006979f
C4462 vdd.n2882 gnd 0.006979f
C4463 vdd.n2883 gnd 0.006979f
C4464 vdd.n2884 gnd 0.006979f
C4465 vdd.n2885 gnd 0.006979f
C4466 vdd.n2886 gnd 0.629284f
C4467 vdd.n2887 gnd 0.006979f
C4468 vdd.n2888 gnd 0.006979f
C4469 vdd.n2889 gnd 0.006979f
C4470 vdd.n2890 gnd 0.006979f
C4471 vdd.n2891 gnd 0.006979f
C4472 vdd.n2892 gnd 0.5716f
C4473 vdd.n2893 gnd 0.006979f
C4474 vdd.n2894 gnd 0.006979f
C4475 vdd.n2895 gnd 0.006979f
C4476 vdd.n2896 gnd 0.006979f
C4477 vdd.n2897 gnd 0.006979f
C4478 vdd.n2898 gnd 0.414279f
C4479 vdd.n2899 gnd 0.006979f
C4480 vdd.n2900 gnd 0.006979f
C4481 vdd.n2901 gnd 0.006979f
C4482 vdd.n2902 gnd 0.006979f
C4483 vdd.n2903 gnd 0.006979f
C4484 vdd.n2904 gnd 0.225494f
C4485 vdd.n2905 gnd 0.006979f
C4486 vdd.n2906 gnd 0.006979f
C4487 vdd.n2907 gnd 0.006979f
C4488 vdd.n2908 gnd 0.006979f
C4489 vdd.n2909 gnd 0.006979f
C4490 vdd.n2910 gnd 0.613552f
C4491 vdd.n2911 gnd 0.006979f
C4492 vdd.n2912 gnd 0.006979f
C4493 vdd.n2913 gnd 0.006979f
C4494 vdd.n2914 gnd 0.006979f
C4495 vdd.n2915 gnd 0.006979f
C4496 vdd.n2916 gnd 0.713189f
C4497 vdd.n2917 gnd 0.006979f
C4498 vdd.n2918 gnd 0.006979f
C4499 vdd.n2919 gnd 0.004516f
C4500 vdd.n2920 gnd 0.020216f
C4501 vdd.n2921 gnd 0.005952f
C4502 vdd.n2922 gnd 0.006979f
C4503 vdd.n2923 gnd 0.608308f
C4504 vdd.n2924 gnd 0.006979f
C4505 vdd.n2925 gnd 0.006979f
C4506 vdd.n2926 gnd 0.006979f
C4507 vdd.n2927 gnd 0.006979f
C4508 vdd.n2928 gnd 0.006979f
C4509 vdd.n2929 gnd 0.498183f
C4510 vdd.n2930 gnd 0.006979f
C4511 vdd.n2931 gnd 0.006979f
C4512 vdd.n2932 gnd 0.006979f
C4513 vdd.n2933 gnd 0.006979f
C4514 vdd.n2934 gnd 0.006979f
C4515 vdd.n2935 gnd 0.372327f
C4516 vdd.n2936 gnd 0.006979f
C4517 vdd.n2937 gnd 0.006979f
C4518 vdd.n2938 gnd 0.006979f
C4519 vdd.n2939 gnd 0.006979f
C4520 vdd.n2940 gnd 0.006979f
C4521 vdd.n2941 gnd 0.713189f
C4522 vdd.n2942 gnd 0.006979f
C4523 vdd.n2943 gnd 0.006979f
C4524 vdd.n2944 gnd 0.006979f
C4525 vdd.n2945 gnd 0.006979f
C4526 vdd.n2946 gnd 0.006979f
C4527 vdd.n2947 gnd 0.006979f
C4528 vdd.n2949 gnd 0.006979f
C4529 vdd.n2950 gnd 0.006979f
C4530 vdd.n2952 gnd 0.006979f
C4531 vdd.n2953 gnd 0.006979f
C4532 vdd.n2956 gnd 0.006979f
C4533 vdd.n2957 gnd 0.006979f
C4534 vdd.n2958 gnd 0.006979f
C4535 vdd.n2959 gnd 0.006979f
C4536 vdd.n2961 gnd 0.006979f
C4537 vdd.n2962 gnd 0.006979f
C4538 vdd.n2963 gnd 0.006979f
C4539 vdd.n2964 gnd 0.006979f
C4540 vdd.n2965 gnd 0.006979f
C4541 vdd.n2966 gnd 0.006979f
C4542 vdd.n2968 gnd 0.006979f
C4543 vdd.n2969 gnd 0.006979f
C4544 vdd.n2970 gnd 0.006979f
C4545 vdd.n2971 gnd 0.006979f
C4546 vdd.n2972 gnd 0.006979f
C4547 vdd.n2973 gnd 0.006979f
C4548 vdd.n2975 gnd 0.006979f
C4549 vdd.n2976 gnd 0.006979f
C4550 vdd.n2977 gnd 0.006979f
C4551 vdd.n2978 gnd 0.006979f
C4552 vdd.n2979 gnd 0.006979f
C4553 vdd.n2980 gnd 0.006979f
C4554 vdd.n2982 gnd 0.006979f
C4555 vdd.n2983 gnd 0.016323f
C4556 vdd.n2984 gnd 0.016323f
C4557 vdd.n2985 gnd 0.015287f
C4558 vdd.n2986 gnd 0.006979f
C4559 vdd.n2987 gnd 0.006979f
C4560 vdd.n2988 gnd 0.006979f
C4561 vdd.n2989 gnd 0.006979f
C4562 vdd.n2990 gnd 0.006979f
C4563 vdd.n2991 gnd 0.006979f
C4564 vdd.n2992 gnd 0.713189f
C4565 vdd.n2993 gnd 0.006979f
C4566 vdd.n2994 gnd 0.006979f
C4567 vdd.n2995 gnd 0.006979f
C4568 vdd.n2996 gnd 0.006979f
C4569 vdd.n2997 gnd 0.006979f
C4570 vdd.n2998 gnd 0.466719f
C4571 vdd.n2999 gnd 0.006979f
C4572 vdd.n3000 gnd 0.006979f
C4573 vdd.n3001 gnd 0.006979f
C4574 vdd.n3002 gnd 0.016154f
C4575 vdd.n3004 gnd 0.016323f
C4576 vdd.n3005 gnd 0.015456f
C4577 vdd.n3006 gnd 0.006979f
C4578 vdd.n3007 gnd 0.005388f
C4579 vdd.n3008 gnd 0.006979f
C4580 vdd.n3010 gnd 0.006979f
C4581 vdd.n3011 gnd 0.006979f
C4582 vdd.n3012 gnd 0.006979f
C4583 vdd.n3013 gnd 0.006979f
C4584 vdd.n3014 gnd 0.006979f
C4585 vdd.n3015 gnd 0.006979f
C4586 vdd.n3017 gnd 0.006979f
C4587 vdd.n3018 gnd 0.006979f
C4588 vdd.n3019 gnd 0.006979f
C4589 vdd.n3020 gnd 0.006979f
C4590 vdd.n3021 gnd 0.006979f
C4591 vdd.n3022 gnd 0.006979f
C4592 vdd.n3024 gnd 0.006979f
C4593 vdd.n3025 gnd 0.006979f
C4594 vdd.n3026 gnd 0.006979f
C4595 vdd.n3027 gnd 0.006979f
C4596 vdd.n3028 gnd 0.006979f
C4597 vdd.n3029 gnd 0.006979f
C4598 vdd.n3031 gnd 0.006979f
C4599 vdd.n3032 gnd 0.006979f
C4600 vdd.n3033 gnd 0.006979f
C4601 vdd.n3034 gnd 0.78013f
C4602 vdd.n3035 gnd 0.023967f
C4603 vdd.n3036 gnd 0.006979f
C4604 vdd.n3037 gnd 0.006979f
C4605 vdd.n3039 gnd 0.006979f
C4606 vdd.n3040 gnd 0.006979f
C4607 vdd.n3041 gnd 0.006979f
C4608 vdd.n3042 gnd 0.006979f
C4609 vdd.n3043 gnd 0.006979f
C4610 vdd.n3044 gnd 0.006979f
C4611 vdd.n3046 gnd 0.006979f
C4612 vdd.n3047 gnd 0.006979f
C4613 vdd.n3048 gnd 0.006979f
C4614 vdd.n3049 gnd 0.006979f
C4615 vdd.n3050 gnd 0.006979f
C4616 vdd.n3051 gnd 0.006979f
C4617 vdd.n3053 gnd 0.006979f
C4618 vdd.n3054 gnd 0.006979f
C4619 vdd.n3055 gnd 0.006979f
C4620 vdd.n3056 gnd 0.006979f
C4621 vdd.n3057 gnd 0.006979f
C4622 vdd.n3058 gnd 0.006979f
C4623 vdd.n3060 gnd 0.006979f
C4624 vdd.n3061 gnd 0.006979f
C4625 vdd.n3063 gnd 0.006979f
C4626 vdd.n3064 gnd 0.006979f
C4627 vdd.n3065 gnd 0.016323f
C4628 vdd.n3066 gnd 0.015287f
C4629 vdd.n3067 gnd 0.015287f
C4630 vdd.n3068 gnd 1.00686f
C4631 vdd.n3069 gnd 0.015287f
C4632 vdd.n3070 gnd 0.016323f
C4633 vdd.n3071 gnd 0.015456f
C4634 vdd.n3072 gnd 0.006979f
C4635 vdd.n3073 gnd 0.005388f
C4636 vdd.n3074 gnd 0.006979f
C4637 vdd.n3076 gnd 0.006979f
C4638 vdd.n3077 gnd 0.006979f
C4639 vdd.n3078 gnd 0.006979f
C4640 vdd.n3079 gnd 0.006979f
C4641 vdd.n3080 gnd 0.006979f
C4642 vdd.n3081 gnd 0.006979f
C4643 vdd.n3083 gnd 0.006979f
C4644 vdd.n3084 gnd 0.006979f
C4645 vdd.n3085 gnd 0.006979f
C4646 vdd.n3086 gnd 0.006979f
C4647 vdd.n3087 gnd 0.006979f
C4648 vdd.n3088 gnd 0.006979f
C4649 vdd.n3090 gnd 0.006979f
C4650 vdd.n3091 gnd 0.006979f
C4651 vdd.n3092 gnd 0.006979f
C4652 vdd.n3093 gnd 0.006979f
C4653 vdd.n3094 gnd 0.006979f
C4654 vdd.n3095 gnd 0.006979f
C4655 vdd.n3097 gnd 0.006979f
C4656 vdd.n3098 gnd 0.006979f
C4657 vdd.n3100 gnd 0.006979f
C4658 vdd.n3101 gnd 0.023967f
C4659 vdd.n3102 gnd 0.78013f
C4660 vdd.n3103 gnd 0.008826f
C4661 vdd.n3104 gnd 0.003924f
C4662 vdd.t59 gnd 0.126259f
C4663 vdd.t60 gnd 0.134936f
C4664 vdd.t57 gnd 0.164893f
C4665 vdd.n3105 gnd 0.211369f
C4666 vdd.n3106 gnd 0.177588f
C4667 vdd.n3107 gnd 0.012721f
C4668 vdd.n3108 gnd 0.010263f
C4669 vdd.n3109 gnd 0.004337f
C4670 vdd.n3110 gnd 0.00826f
C4671 vdd.n3111 gnd 0.010263f
C4672 vdd.n3112 gnd 0.010263f
C4673 vdd.n3113 gnd 0.00826f
C4674 vdd.n3114 gnd 0.00826f
C4675 vdd.n3115 gnd 0.010263f
C4676 vdd.n3117 gnd 0.010263f
C4677 vdd.n3118 gnd 0.00826f
C4678 vdd.n3119 gnd 0.00826f
C4679 vdd.n3120 gnd 0.00826f
C4680 vdd.n3121 gnd 0.010263f
C4681 vdd.n3123 gnd 0.010263f
C4682 vdd.n3125 gnd 0.010263f
C4683 vdd.n3126 gnd 0.00826f
C4684 vdd.n3127 gnd 0.00826f
C4685 vdd.n3128 gnd 0.00826f
C4686 vdd.n3129 gnd 0.010263f
C4687 vdd.n3131 gnd 0.010263f
C4688 vdd.n3133 gnd 0.010263f
C4689 vdd.n3134 gnd 0.00826f
C4690 vdd.n3135 gnd 0.00826f
C4691 vdd.n3136 gnd 0.00826f
C4692 vdd.n3137 gnd 0.010263f
C4693 vdd.n3139 gnd 0.010263f
C4694 vdd.n3140 gnd 0.010263f
C4695 vdd.n3141 gnd 0.00826f
C4696 vdd.n3142 gnd 0.00826f
C4697 vdd.n3143 gnd 0.010263f
C4698 vdd.n3144 gnd 0.010263f
C4699 vdd.n3146 gnd 0.010263f
C4700 vdd.n3147 gnd 0.00826f
C4701 vdd.n3148 gnd 0.010263f
C4702 vdd.n3149 gnd 0.010263f
C4703 vdd.n3150 gnd 0.010263f
C4704 vdd.n3151 gnd 0.016851f
C4705 vdd.n3152 gnd 0.005617f
C4706 vdd.n3153 gnd 0.010263f
C4707 vdd.n3155 gnd 0.010263f
C4708 vdd.n3157 gnd 0.010263f
C4709 vdd.n3158 gnd 0.00826f
C4710 vdd.n3159 gnd 0.00826f
C4711 vdd.n3160 gnd 0.00826f
C4712 vdd.n3161 gnd 0.010263f
C4713 vdd.n3163 gnd 0.010263f
C4714 vdd.n3165 gnd 0.010263f
C4715 vdd.n3166 gnd 0.00826f
C4716 vdd.n3167 gnd 0.00826f
C4717 vdd.n3168 gnd 0.00826f
C4718 vdd.n3169 gnd 0.010263f
C4719 vdd.n3171 gnd 0.010263f
C4720 vdd.n3173 gnd 0.010263f
C4721 vdd.n3174 gnd 0.00826f
C4722 vdd.n3175 gnd 0.00826f
C4723 vdd.n3176 gnd 0.00826f
C4724 vdd.n3177 gnd 0.010263f
C4725 vdd.n3179 gnd 0.010263f
C4726 vdd.n3181 gnd 0.010263f
C4727 vdd.n3182 gnd 0.00826f
C4728 vdd.n3183 gnd 0.00826f
C4729 vdd.n3184 gnd 0.00826f
C4730 vdd.n3185 gnd 0.010263f
C4731 vdd.n3187 gnd 0.010263f
C4732 vdd.n3189 gnd 0.010263f
C4733 vdd.n3190 gnd 0.00826f
C4734 vdd.n3191 gnd 0.00826f
C4735 vdd.n3192 gnd 0.006897f
C4736 vdd.n3193 gnd 0.010263f
C4737 vdd.n3195 gnd 0.010263f
C4738 vdd.n3197 gnd 0.010263f
C4739 vdd.n3198 gnd 0.006897f
C4740 vdd.n3199 gnd 0.00826f
C4741 vdd.n3200 gnd 0.00826f
C4742 vdd.n3201 gnd 0.010263f
C4743 vdd.n3203 gnd 0.010263f
C4744 vdd.n3205 gnd 0.010263f
C4745 vdd.n3206 gnd 0.00826f
C4746 vdd.n3207 gnd 0.00826f
C4747 vdd.n3208 gnd 0.00826f
C4748 vdd.n3209 gnd 0.010263f
C4749 vdd.n3211 gnd 0.010263f
C4750 vdd.n3213 gnd 0.010263f
C4751 vdd.n3214 gnd 0.00826f
C4752 vdd.n3215 gnd 0.00826f
C4753 vdd.n3216 gnd 0.00826f
C4754 vdd.n3217 gnd 0.010263f
C4755 vdd.n3219 gnd 0.010263f
C4756 vdd.n3220 gnd 0.010263f
C4757 vdd.n3221 gnd 0.00826f
C4758 vdd.n3222 gnd 0.00826f
C4759 vdd.n3223 gnd 0.010263f
C4760 vdd.n3224 gnd 0.010263f
C4761 vdd.n3225 gnd 0.00826f
C4762 vdd.n3226 gnd 0.00826f
C4763 vdd.n3227 gnd 0.010263f
C4764 vdd.n3228 gnd 0.010263f
C4765 vdd.n3230 gnd 0.010263f
C4766 vdd.n3231 gnd 0.00826f
C4767 vdd.n3232 gnd 0.006856f
C4768 vdd.n3233 gnd 0.02353f
C4769 vdd.n3234 gnd 0.023371f
C4770 vdd.n3235 gnd 0.006856f
C4771 vdd.n3236 gnd 0.023371f
C4772 vdd.n3237 gnd 1.38443f
C4773 vdd.n3238 gnd 0.023371f
C4774 vdd.n3239 gnd 0.006856f
C4775 vdd.n3240 gnd 0.023371f
C4776 vdd.n3241 gnd 0.010263f
C4777 vdd.n3242 gnd 0.010263f
C4778 vdd.n3243 gnd 0.00826f
C4779 vdd.n3244 gnd 0.010263f
C4780 vdd.n3245 gnd 0.991123f
C4781 vdd.n3246 gnd 0.010263f
C4782 vdd.n3247 gnd 0.00826f
C4783 vdd.n3248 gnd 0.010263f
C4784 vdd.n3249 gnd 0.010263f
C4785 vdd.n3250 gnd 0.010263f
C4786 vdd.n3251 gnd 0.00826f
C4787 vdd.n3252 gnd 0.010263f
C4788 vdd.n3253 gnd 1.02259f
C4789 vdd.n3254 gnd 0.010263f
C4790 vdd.n3255 gnd 0.00826f
C4791 vdd.n3256 gnd 0.010263f
C4792 vdd.n3257 gnd 0.010263f
C4793 vdd.n3258 gnd 0.010263f
C4794 vdd.n3259 gnd 0.00826f
C4795 vdd.n3260 gnd 0.010263f
C4796 vdd.t234 gnd 0.524404f
C4797 vdd.n3261 gnd 0.84429f
C4798 vdd.n3262 gnd 0.010263f
C4799 vdd.n3263 gnd 0.00826f
C4800 vdd.n3264 gnd 0.010263f
C4801 vdd.n3265 gnd 0.010263f
C4802 vdd.n3266 gnd 0.010263f
C4803 vdd.n3267 gnd 0.00826f
C4804 vdd.n3268 gnd 0.010263f
C4805 vdd.n3269 gnd 0.665993f
C4806 vdd.n3270 gnd 0.010263f
C4807 vdd.n3271 gnd 0.00826f
C4808 vdd.n3272 gnd 0.010263f
C4809 vdd.n3273 gnd 0.010263f
C4810 vdd.n3274 gnd 0.010263f
C4811 vdd.n3275 gnd 0.00826f
C4812 vdd.n3276 gnd 0.010263f
C4813 vdd.n3277 gnd 0.833802f
C4814 vdd.n3278 gnd 0.561112f
C4815 vdd.n3279 gnd 0.010263f
C4816 vdd.n3280 gnd 0.00826f
C4817 vdd.n3281 gnd 0.010263f
C4818 vdd.n3282 gnd 0.010263f
C4819 vdd.n3283 gnd 0.010263f
C4820 vdd.n3284 gnd 0.00826f
C4821 vdd.n3285 gnd 0.010263f
C4822 vdd.n3286 gnd 0.739409f
C4823 vdd.n3287 gnd 0.010263f
C4824 vdd.n3288 gnd 0.00826f
C4825 vdd.n3289 gnd 0.010263f
C4826 vdd.n3290 gnd 0.010263f
C4827 vdd.n3291 gnd 0.010263f
C4828 vdd.n3292 gnd 0.010263f
C4829 vdd.n3293 gnd 0.010263f
C4830 vdd.n3294 gnd 0.00826f
C4831 vdd.n3295 gnd 0.00826f
C4832 vdd.n3296 gnd 0.010263f
C4833 vdd.t180 gnd 0.524404f
C4834 vdd.n3297 gnd 0.87051f
C4835 vdd.n3298 gnd 0.010263f
C4836 vdd.n3299 gnd 0.00826f
C4837 vdd.n3300 gnd 0.010263f
C4838 vdd.n3301 gnd 0.010263f
C4839 vdd.n3302 gnd 0.010263f
C4840 vdd.n3303 gnd 0.00826f
C4841 vdd.n3304 gnd 0.010263f
C4842 vdd.n3305 gnd 0.823314f
C4843 vdd.n3306 gnd 0.010263f
C4844 vdd.n3307 gnd 0.010263f
C4845 vdd.n3308 gnd 0.00826f
C4846 vdd.n3309 gnd 0.00826f
C4847 vdd.n3310 gnd 0.00826f
C4848 vdd.n3311 gnd 0.010263f
C4849 vdd.n3312 gnd 0.010263f
C4850 vdd.n3313 gnd 0.010263f
C4851 vdd.n3314 gnd 0.010263f
C4852 vdd.n3315 gnd 0.00826f
C4853 vdd.n3316 gnd 0.00826f
C4854 vdd.n3317 gnd 0.00826f
C4855 vdd.n3318 gnd 0.010263f
C4856 vdd.n3319 gnd 0.010263f
C4857 vdd.n3320 gnd 0.010263f
C4858 vdd.n3321 gnd 0.010263f
C4859 vdd.n3322 gnd 0.00826f
C4860 vdd.n3323 gnd 0.00826f
C4861 vdd.n3324 gnd 0.00826f
C4862 vdd.n3325 gnd 0.010263f
C4863 vdd.n3326 gnd 0.010263f
C4864 vdd.n3327 gnd 0.010263f
C4865 vdd.n3328 gnd 0.87051f
C4866 vdd.n3329 gnd 0.010263f
C4867 vdd.n3330 gnd 0.00826f
C4868 vdd.n3331 gnd 0.00826f
C4869 vdd.n3332 gnd 0.00826f
C4870 vdd.n3333 gnd 0.010263f
C4871 vdd.n3334 gnd 0.010263f
C4872 vdd.n3335 gnd 0.010263f
C4873 vdd.n3336 gnd 0.010263f
C4874 vdd.n3337 gnd 0.00826f
C4875 vdd.n3338 gnd 0.00826f
C4876 vdd.n3339 gnd 0.006856f
C4877 vdd.n3340 gnd 0.023371f
C4878 vdd.n3341 gnd 0.02353f
C4879 vdd.n3342 gnd 0.003924f
C4880 vdd.n3343 gnd 0.02353f
C4881 vdd.n3345 gnd 2.31786f
C4882 vdd.n3346 gnd 1.38443f
C4883 vdd.n3347 gnd 0.686969f
C4884 vdd.n3348 gnd 0.010263f
C4885 vdd.n3349 gnd 0.00826f
C4886 vdd.n3350 gnd 0.00826f
C4887 vdd.n3351 gnd 0.00826f
C4888 vdd.n3352 gnd 0.010263f
C4889 vdd.n3353 gnd 1.04881f
C4890 vdd.n3354 gnd 1.04881f
C4891 vdd.n3355 gnd 0.603064f
C4892 vdd.n3356 gnd 0.010263f
C4893 vdd.n3357 gnd 0.00826f
C4894 vdd.n3358 gnd 0.00826f
C4895 vdd.n3359 gnd 0.00826f
C4896 vdd.n3360 gnd 0.010263f
C4897 vdd.n3361 gnd 0.62404f
C4898 vdd.n3362 gnd 0.770873f
C4899 vdd.t150 gnd 0.524404f
C4900 vdd.n3363 gnd 0.802338f
C4901 vdd.n3364 gnd 0.010263f
C4902 vdd.n3365 gnd 0.00826f
C4903 vdd.n3366 gnd 0.00826f
C4904 vdd.n3367 gnd 0.00826f
C4905 vdd.n3368 gnd 0.010263f
C4906 vdd.n3369 gnd 0.87051f
C4907 vdd.t159 gnd 0.524404f
C4908 vdd.n3370 gnd 0.634528f
C4909 vdd.n3371 gnd 0.760385f
C4910 vdd.n3372 gnd 0.010263f
C4911 vdd.n3373 gnd 0.00826f
C4912 vdd.n3374 gnd 0.00826f
C4913 vdd.n3375 gnd 0.00826f
C4914 vdd.n3376 gnd 0.010263f
C4915 vdd.n3377 gnd 0.582088f
C4916 vdd.t183 gnd 0.524404f
C4917 vdd.n3378 gnd 0.87051f
C4918 vdd.t204 gnd 0.524404f
C4919 vdd.n3379 gnd 0.645016f
C4920 vdd.n3380 gnd 0.010263f
C4921 vdd.n3381 gnd 0.00826f
C4922 vdd.n3382 gnd 0.007888f
C4923 vdd.n3383 gnd 0.605337f
C4924 vdd.n3384 gnd 2.56752f
C4925 a_n7636_8799.n0 gnd 2.71862f
C4926 a_n7636_8799.n1 gnd 1.64714f
C4927 a_n7636_8799.n2 gnd 3.76848f
C4928 a_n7636_8799.n3 gnd 0.205533f
C4929 a_n7636_8799.n4 gnd 0.287271f
C4930 a_n7636_8799.n5 gnd 0.205533f
C4931 a_n7636_8799.n6 gnd 0.205533f
C4932 a_n7636_8799.n7 gnd 0.205533f
C4933 a_n7636_8799.n8 gnd 0.27078f
C4934 a_n7636_8799.n9 gnd 0.205533f
C4935 a_n7636_8799.n10 gnd 0.287271f
C4936 a_n7636_8799.n11 gnd 0.205533f
C4937 a_n7636_8799.n12 gnd 0.205533f
C4938 a_n7636_8799.n13 gnd 0.205533f
C4939 a_n7636_8799.n14 gnd 0.27078f
C4940 a_n7636_8799.n15 gnd 0.205533f
C4941 a_n7636_8799.n16 gnd 0.45021f
C4942 a_n7636_8799.n17 gnd 0.205533f
C4943 a_n7636_8799.n18 gnd 0.205533f
C4944 a_n7636_8799.n19 gnd 0.205533f
C4945 a_n7636_8799.n20 gnd 0.27078f
C4946 a_n7636_8799.n21 gnd 0.322163f
C4947 a_n7636_8799.n22 gnd 0.205533f
C4948 a_n7636_8799.n23 gnd 0.205533f
C4949 a_n7636_8799.n24 gnd 0.205533f
C4950 a_n7636_8799.n25 gnd 0.205533f
C4951 a_n7636_8799.n26 gnd 0.235888f
C4952 a_n7636_8799.n27 gnd 0.322163f
C4953 a_n7636_8799.n28 gnd 0.205533f
C4954 a_n7636_8799.n29 gnd 0.205533f
C4955 a_n7636_8799.n30 gnd 0.205533f
C4956 a_n7636_8799.n31 gnd 0.205533f
C4957 a_n7636_8799.n32 gnd 0.235888f
C4958 a_n7636_8799.n33 gnd 0.322163f
C4959 a_n7636_8799.n34 gnd 0.205533f
C4960 a_n7636_8799.n35 gnd 0.205533f
C4961 a_n7636_8799.n36 gnd 0.205533f
C4962 a_n7636_8799.n37 gnd 0.205533f
C4963 a_n7636_8799.n38 gnd 0.398827f
C4964 a_n7636_8799.n39 gnd 1.00902f
C4965 a_n7636_8799.n40 gnd 2.51925f
C4966 a_n7636_8799.n41 gnd 1.50639f
C4967 a_n7636_8799.n42 gnd 0.008525f
C4968 a_n7636_8799.n43 gnd 0.001144f
C4969 a_n7636_8799.n45 gnd 0.007655f
C4970 a_n7636_8799.n46 gnd 0.011571f
C4971 a_n7636_8799.n47 gnd 0.007958f
C4972 a_n7636_8799.n49 gnd 3.98e-19
C4973 a_n7636_8799.n50 gnd 0.008247f
C4974 a_n7636_8799.n51 gnd 0.01139f
C4975 a_n7636_8799.n52 gnd 0.007339f
C4976 a_n7636_8799.n53 gnd 0.008525f
C4977 a_n7636_8799.n54 gnd 0.001144f
C4978 a_n7636_8799.n56 gnd 0.007655f
C4979 a_n7636_8799.n57 gnd 0.011571f
C4980 a_n7636_8799.n58 gnd 0.007958f
C4981 a_n7636_8799.n60 gnd 3.98e-19
C4982 a_n7636_8799.n61 gnd 0.008247f
C4983 a_n7636_8799.n62 gnd 0.01139f
C4984 a_n7636_8799.n63 gnd 0.007339f
C4985 a_n7636_8799.n64 gnd 0.008525f
C4986 a_n7636_8799.n65 gnd 0.001144f
C4987 a_n7636_8799.n67 gnd 0.007655f
C4988 a_n7636_8799.n68 gnd 0.011571f
C4989 a_n7636_8799.n69 gnd 0.007958f
C4990 a_n7636_8799.n71 gnd 3.98e-19
C4991 a_n7636_8799.n72 gnd 0.008247f
C4992 a_n7636_8799.n73 gnd 0.01139f
C4993 a_n7636_8799.n74 gnd 0.007339f
C4994 a_n7636_8799.n75 gnd 0.001144f
C4995 a_n7636_8799.n77 gnd 0.007655f
C4996 a_n7636_8799.n78 gnd 0.011571f
C4997 a_n7636_8799.n79 gnd 0.007958f
C4998 a_n7636_8799.n81 gnd 3.98e-19
C4999 a_n7636_8799.n82 gnd 0.008247f
C5000 a_n7636_8799.n83 gnd 0.01139f
C5001 a_n7636_8799.n84 gnd 0.007339f
C5002 a_n7636_8799.n85 gnd 0.247442f
C5003 a_n7636_8799.n86 gnd 0.001144f
C5004 a_n7636_8799.n88 gnd 0.007655f
C5005 a_n7636_8799.n89 gnd 0.011571f
C5006 a_n7636_8799.n90 gnd 0.007958f
C5007 a_n7636_8799.n92 gnd 3.98e-19
C5008 a_n7636_8799.n93 gnd 0.008247f
C5009 a_n7636_8799.n94 gnd 0.01139f
C5010 a_n7636_8799.n95 gnd 0.007339f
C5011 a_n7636_8799.n96 gnd 0.247442f
C5012 a_n7636_8799.n97 gnd 0.001144f
C5013 a_n7636_8799.n99 gnd 0.007655f
C5014 a_n7636_8799.n100 gnd 0.011571f
C5015 a_n7636_8799.n101 gnd 0.007958f
C5016 a_n7636_8799.n103 gnd 3.98e-19
C5017 a_n7636_8799.n104 gnd 0.008247f
C5018 a_n7636_8799.n105 gnd 0.01139f
C5019 a_n7636_8799.n106 gnd 0.007339f
C5020 a_n7636_8799.n107 gnd 0.247442f
C5021 a_n7636_8799.t21 gnd 0.14256f
C5022 a_n7636_8799.t14 gnd 0.14256f
C5023 a_n7636_8799.t19 gnd 0.14256f
C5024 a_n7636_8799.n108 gnd 1.12439f
C5025 a_n7636_8799.t16 gnd 0.14256f
C5026 a_n7636_8799.t7 gnd 0.14256f
C5027 a_n7636_8799.n109 gnd 1.12254f
C5028 a_n7636_8799.t26 gnd 0.14256f
C5029 a_n7636_8799.t22 gnd 0.14256f
C5030 a_n7636_8799.n110 gnd 1.12254f
C5031 a_n7636_8799.t17 gnd 0.14256f
C5032 a_n7636_8799.t9 gnd 0.14256f
C5033 a_n7636_8799.n111 gnd 1.12254f
C5034 a_n7636_8799.t11 gnd 0.11088f
C5035 a_n7636_8799.t5 gnd 0.11088f
C5036 a_n7636_8799.n112 gnd 0.982662f
C5037 a_n7636_8799.t0 gnd 0.11088f
C5038 a_n7636_8799.t15 gnd 0.11088f
C5039 a_n7636_8799.n113 gnd 0.979773f
C5040 a_n7636_8799.t12 gnd 0.11088f
C5041 a_n7636_8799.t1 gnd 0.11088f
C5042 a_n7636_8799.n114 gnd 0.982661f
C5043 a_n7636_8799.t20 gnd 0.11088f
C5044 a_n7636_8799.t2 gnd 0.11088f
C5045 a_n7636_8799.n115 gnd 0.979772f
C5046 a_n7636_8799.t4 gnd 0.11088f
C5047 a_n7636_8799.t23 gnd 0.11088f
C5048 a_n7636_8799.n116 gnd 0.982661f
C5049 a_n7636_8799.t30 gnd 0.11088f
C5050 a_n7636_8799.t24 gnd 0.11088f
C5051 a_n7636_8799.n117 gnd 0.979772f
C5052 a_n7636_8799.t25 gnd 0.11088f
C5053 a_n7636_8799.t3 gnd 0.11088f
C5054 a_n7636_8799.n118 gnd 0.979773f
C5055 a_n7636_8799.t13 gnd 0.11088f
C5056 a_n7636_8799.t29 gnd 0.11088f
C5057 a_n7636_8799.n119 gnd 0.979773f
C5058 a_n7636_8799.t74 gnd 0.591119f
C5059 a_n7636_8799.n120 gnd 0.264275f
C5060 a_n7636_8799.t32 gnd 0.591119f
C5061 a_n7636_8799.t57 gnd 0.591119f
C5062 a_n7636_8799.n121 gnd 0.267549f
C5063 a_n7636_8799.t58 gnd 0.591119f
C5064 a_n7636_8799.t68 gnd 0.591119f
C5065 a_n7636_8799.t94 gnd 0.591119f
C5066 a_n7636_8799.n122 gnd 0.26961f
C5067 a_n7636_8799.t110 gnd 0.591119f
C5068 a_n7636_8799.t113 gnd 0.591119f
C5069 a_n7636_8799.n123 gnd 0.263213f
C5070 a_n7636_8799.t111 gnd 0.602307f
C5071 a_n7636_8799.n124 gnd 0.247823f
C5072 a_n7636_8799.n125 gnd 0.01166f
C5073 a_n7636_8799.t69 gnd 0.591119f
C5074 a_n7636_8799.n126 gnd 0.264005f
C5075 a_n7636_8799.n127 gnd 0.267534f
C5076 a_n7636_8799.t67 gnd 0.591119f
C5077 a_n7636_8799.n128 gnd 0.264094f
C5078 a_n7636_8799.n129 gnd 0.258778f
C5079 a_n7636_8799.t92 gnd 0.591119f
C5080 a_n7636_8799.n130 gnd 0.263847f
C5081 a_n7636_8799.n131 gnd 0.27004f
C5082 a_n7636_8799.t89 gnd 0.591119f
C5083 a_n7636_8799.n132 gnd 0.267418f
C5084 a_n7636_8799.n133 gnd 0.26353f
C5085 a_n7636_8799.t56 gnd 0.591119f
C5086 a_n7636_8799.n134 gnd 0.259095f
C5087 a_n7636_8799.t112 gnd 0.591119f
C5088 a_n7636_8799.n135 gnd 0.267533f
C5089 a_n7636_8799.t41 gnd 0.602297f
C5090 a_n7636_8799.t83 gnd 0.591119f
C5091 a_n7636_8799.n136 gnd 0.264275f
C5092 a_n7636_8799.t40 gnd 0.591119f
C5093 a_n7636_8799.t65 gnd 0.591119f
C5094 a_n7636_8799.n137 gnd 0.267549f
C5095 a_n7636_8799.t66 gnd 0.591119f
C5096 a_n7636_8799.t76 gnd 0.591119f
C5097 a_n7636_8799.t107 gnd 0.591119f
C5098 a_n7636_8799.n138 gnd 0.26961f
C5099 a_n7636_8799.t122 gnd 0.591119f
C5100 a_n7636_8799.t126 gnd 0.591119f
C5101 a_n7636_8799.n139 gnd 0.263213f
C5102 a_n7636_8799.t124 gnd 0.602307f
C5103 a_n7636_8799.n140 gnd 0.247823f
C5104 a_n7636_8799.n141 gnd 0.01166f
C5105 a_n7636_8799.t77 gnd 0.591119f
C5106 a_n7636_8799.n142 gnd 0.264005f
C5107 a_n7636_8799.n143 gnd 0.267534f
C5108 a_n7636_8799.t75 gnd 0.591119f
C5109 a_n7636_8799.n144 gnd 0.264094f
C5110 a_n7636_8799.n145 gnd 0.258778f
C5111 a_n7636_8799.t105 gnd 0.591119f
C5112 a_n7636_8799.n146 gnd 0.263847f
C5113 a_n7636_8799.n147 gnd 0.27004f
C5114 a_n7636_8799.t101 gnd 0.591119f
C5115 a_n7636_8799.n148 gnd 0.267418f
C5116 a_n7636_8799.n149 gnd 0.26353f
C5117 a_n7636_8799.t62 gnd 0.591119f
C5118 a_n7636_8799.n150 gnd 0.259095f
C5119 a_n7636_8799.t125 gnd 0.591119f
C5120 a_n7636_8799.n151 gnd 0.267533f
C5121 a_n7636_8799.t51 gnd 0.602297f
C5122 a_n7636_8799.n152 gnd 0.890291f
C5123 a_n7636_8799.t85 gnd 0.591119f
C5124 a_n7636_8799.n153 gnd 0.264275f
C5125 a_n7636_8799.t73 gnd 0.591119f
C5126 a_n7636_8799.t117 gnd 0.591119f
C5127 a_n7636_8799.n154 gnd 0.267549f
C5128 a_n7636_8799.t93 gnd 0.591119f
C5129 a_n7636_8799.t33 gnd 0.591119f
C5130 a_n7636_8799.t63 gnd 0.591119f
C5131 a_n7636_8799.n155 gnd 0.26961f
C5132 a_n7636_8799.t114 gnd 0.591119f
C5133 a_n7636_8799.t72 gnd 0.591119f
C5134 a_n7636_8799.n156 gnd 0.263213f
C5135 a_n7636_8799.t90 gnd 0.602307f
C5136 a_n7636_8799.n157 gnd 0.247823f
C5137 a_n7636_8799.n158 gnd 0.01166f
C5138 a_n7636_8799.t106 gnd 0.591119f
C5139 a_n7636_8799.n159 gnd 0.264005f
C5140 a_n7636_8799.n160 gnd 0.267534f
C5141 a_n7636_8799.t45 gnd 0.591119f
C5142 a_n7636_8799.n161 gnd 0.264094f
C5143 a_n7636_8799.n162 gnd 0.258778f
C5144 a_n7636_8799.t78 gnd 0.591119f
C5145 a_n7636_8799.n163 gnd 0.263847f
C5146 a_n7636_8799.n164 gnd 0.27004f
C5147 a_n7636_8799.t121 gnd 0.591119f
C5148 a_n7636_8799.n165 gnd 0.267418f
C5149 a_n7636_8799.n166 gnd 0.26353f
C5150 a_n7636_8799.t37 gnd 0.591119f
C5151 a_n7636_8799.n167 gnd 0.259095f
C5152 a_n7636_8799.t49 gnd 0.591119f
C5153 a_n7636_8799.n168 gnd 0.267533f
C5154 a_n7636_8799.t102 gnd 0.602297f
C5155 a_n7636_8799.n169 gnd 1.55447f
C5156 a_n7636_8799.t71 gnd 0.591119f
C5157 a_n7636_8799.t53 gnd 0.591119f
C5158 a_n7636_8799.t116 gnd 0.591119f
C5159 a_n7636_8799.n170 gnd 0.26714f
C5160 a_n7636_8799.t84 gnd 0.591119f
C5161 a_n7636_8799.t82 gnd 0.591119f
C5162 a_n7636_8799.t34 gnd 0.591119f
C5163 a_n7636_8799.n171 gnd 0.264094f
C5164 a_n7636_8799.t88 gnd 0.591119f
C5165 a_n7636_8799.t87 gnd 0.591119f
C5166 a_n7636_8799.t36 gnd 0.591119f
C5167 a_n7636_8799.n172 gnd 0.267549f
C5168 a_n7636_8799.t35 gnd 0.591119f
C5169 a_n7636_8799.t104 gnd 0.591119f
C5170 a_n7636_8799.t48 gnd 0.591119f
C5171 a_n7636_8799.n173 gnd 0.26353f
C5172 a_n7636_8799.t39 gnd 0.591119f
C5173 a_n7636_8799.t108 gnd 0.591119f
C5174 a_n7636_8799.t70 gnd 0.591119f
C5175 a_n7636_8799.n174 gnd 0.267533f
C5176 a_n7636_8799.t52 gnd 0.602307f
C5177 a_n7636_8799.n175 gnd 0.247823f
C5178 a_n7636_8799.n176 gnd 0.264275f
C5179 a_n7636_8799.n177 gnd 0.259095f
C5180 a_n7636_8799.n178 gnd 0.267418f
C5181 a_n7636_8799.n179 gnd 0.27004f
C5182 a_n7636_8799.n180 gnd 0.263847f
C5183 a_n7636_8799.n181 gnd 0.258778f
C5184 a_n7636_8799.n182 gnd 0.267534f
C5185 a_n7636_8799.n183 gnd 0.26961f
C5186 a_n7636_8799.n184 gnd 0.263213f
C5187 a_n7636_8799.n185 gnd 0.258619f
C5188 a_n7636_8799.t80 gnd 0.591119f
C5189 a_n7636_8799.t60 gnd 0.591119f
C5190 a_n7636_8799.t127 gnd 0.591119f
C5191 a_n7636_8799.n186 gnd 0.26714f
C5192 a_n7636_8799.t97 gnd 0.591119f
C5193 a_n7636_8799.t96 gnd 0.591119f
C5194 a_n7636_8799.t42 gnd 0.591119f
C5195 a_n7636_8799.n187 gnd 0.264094f
C5196 a_n7636_8799.t100 gnd 0.591119f
C5197 a_n7636_8799.t99 gnd 0.591119f
C5198 a_n7636_8799.t44 gnd 0.591119f
C5199 a_n7636_8799.n188 gnd 0.267549f
C5200 a_n7636_8799.t43 gnd 0.591119f
C5201 a_n7636_8799.t119 gnd 0.591119f
C5202 a_n7636_8799.t59 gnd 0.591119f
C5203 a_n7636_8799.n189 gnd 0.26353f
C5204 a_n7636_8799.t47 gnd 0.591119f
C5205 a_n7636_8799.t120 gnd 0.591119f
C5206 a_n7636_8799.t81 gnd 0.591119f
C5207 a_n7636_8799.n190 gnd 0.267533f
C5208 a_n7636_8799.t61 gnd 0.602307f
C5209 a_n7636_8799.n191 gnd 0.247823f
C5210 a_n7636_8799.n192 gnd 0.264275f
C5211 a_n7636_8799.n193 gnd 0.259095f
C5212 a_n7636_8799.n194 gnd 0.267418f
C5213 a_n7636_8799.n195 gnd 0.27004f
C5214 a_n7636_8799.n196 gnd 0.263847f
C5215 a_n7636_8799.n197 gnd 0.258778f
C5216 a_n7636_8799.n198 gnd 0.267534f
C5217 a_n7636_8799.n199 gnd 0.26961f
C5218 a_n7636_8799.n200 gnd 0.263213f
C5219 a_n7636_8799.n201 gnd 0.258619f
C5220 a_n7636_8799.n202 gnd 0.890291f
C5221 a_n7636_8799.t103 gnd 0.591119f
C5222 a_n7636_8799.t50 gnd 0.591119f
C5223 a_n7636_8799.t86 gnd 0.591119f
C5224 a_n7636_8799.n203 gnd 0.26714f
C5225 a_n7636_8799.t38 gnd 0.591119f
C5226 a_n7636_8799.t55 gnd 0.591119f
C5227 a_n7636_8799.t123 gnd 0.591119f
C5228 a_n7636_8799.n204 gnd 0.264094f
C5229 a_n7636_8799.t95 gnd 0.591119f
C5230 a_n7636_8799.t118 gnd 0.591119f
C5231 a_n7636_8799.t79 gnd 0.591119f
C5232 a_n7636_8799.n205 gnd 0.267549f
C5233 a_n7636_8799.t98 gnd 0.591119f
C5234 a_n7636_8799.t46 gnd 0.591119f
C5235 a_n7636_8799.t115 gnd 0.591119f
C5236 a_n7636_8799.n206 gnd 0.26353f
C5237 a_n7636_8799.t64 gnd 0.591119f
C5238 a_n7636_8799.t109 gnd 0.591119f
C5239 a_n7636_8799.t54 gnd 0.591119f
C5240 a_n7636_8799.n207 gnd 0.267533f
C5241 a_n7636_8799.t91 gnd 0.602307f
C5242 a_n7636_8799.n208 gnd 0.247823f
C5243 a_n7636_8799.n209 gnd 0.264275f
C5244 a_n7636_8799.n210 gnd 0.259095f
C5245 a_n7636_8799.n211 gnd 0.267418f
C5246 a_n7636_8799.n212 gnd 0.27004f
C5247 a_n7636_8799.n213 gnd 0.263847f
C5248 a_n7636_8799.n214 gnd 0.258778f
C5249 a_n7636_8799.n215 gnd 0.267534f
C5250 a_n7636_8799.n216 gnd 0.26961f
C5251 a_n7636_8799.n217 gnd 0.263213f
C5252 a_n7636_8799.n218 gnd 0.258619f
C5253 a_n7636_8799.n219 gnd 1.20614f
C5254 a_n7636_8799.n220 gnd 13.8223f
C5255 a_n7636_8799.n221 gnd 4.32613f
C5256 a_n7636_8799.n222 gnd 6.27519f
C5257 a_n7636_8799.t27 gnd 0.14256f
C5258 a_n7636_8799.t10 gnd 0.14256f
C5259 a_n7636_8799.n223 gnd 1.12439f
C5260 a_n7636_8799.t8 gnd 0.14256f
C5261 a_n7636_8799.t18 gnd 0.14256f
C5262 a_n7636_8799.n224 gnd 1.12254f
C5263 a_n7636_8799.t28 gnd 0.14256f
C5264 a_n7636_8799.t31 gnd 0.14256f
C5265 a_n7636_8799.n225 gnd 1.12254f
C5266 a_n7636_8799.n226 gnd 3.15296f
C5267 a_n7636_8799.n227 gnd 1.12254f
C5268 a_n7636_8799.t6 gnd 0.14256f
C5269 commonsourceibias.n0 gnd 0.012626f
C5270 commonsourceibias.t78 gnd 0.191194f
C5271 commonsourceibias.t146 gnd 0.176786f
C5272 commonsourceibias.n1 gnd 0.007691f
C5273 commonsourceibias.n2 gnd 0.009462f
C5274 commonsourceibias.t96 gnd 0.176786f
C5275 commonsourceibias.n3 gnd 0.009599f
C5276 commonsourceibias.n4 gnd 0.009462f
C5277 commonsourceibias.t157 gnd 0.176786f
C5278 commonsourceibias.n5 gnd 0.070538f
C5279 commonsourceibias.t112 gnd 0.176786f
C5280 commonsourceibias.n6 gnd 0.007654f
C5281 commonsourceibias.n7 gnd 0.009462f
C5282 commonsourceibias.t75 gnd 0.176786f
C5283 commonsourceibias.n8 gnd 0.009135f
C5284 commonsourceibias.n9 gnd 0.009462f
C5285 commonsourceibias.t124 gnd 0.176786f
C5286 commonsourceibias.n10 gnd 0.070538f
C5287 commonsourceibias.t113 gnd 0.176786f
C5288 commonsourceibias.n11 gnd 0.007642f
C5289 commonsourceibias.n12 gnd 0.012626f
C5290 commonsourceibias.t36 gnd 0.191194f
C5291 commonsourceibias.t32 gnd 0.176786f
C5292 commonsourceibias.n13 gnd 0.007691f
C5293 commonsourceibias.n14 gnd 0.009462f
C5294 commonsourceibias.t42 gnd 0.176786f
C5295 commonsourceibias.n15 gnd 0.009599f
C5296 commonsourceibias.n16 gnd 0.009462f
C5297 commonsourceibias.t20 gnd 0.176786f
C5298 commonsourceibias.n17 gnd 0.070538f
C5299 commonsourceibias.t0 gnd 0.176786f
C5300 commonsourceibias.n18 gnd 0.007654f
C5301 commonsourceibias.n19 gnd 0.009462f
C5302 commonsourceibias.t38 gnd 0.176786f
C5303 commonsourceibias.n20 gnd 0.009135f
C5304 commonsourceibias.n21 gnd 0.009462f
C5305 commonsourceibias.t50 gnd 0.176786f
C5306 commonsourceibias.n22 gnd 0.070538f
C5307 commonsourceibias.t58 gnd 0.176786f
C5308 commonsourceibias.n23 gnd 0.007642f
C5309 commonsourceibias.n24 gnd 0.009462f
C5310 commonsourceibias.t24 gnd 0.176786f
C5311 commonsourceibias.t4 gnd 0.176786f
C5312 commonsourceibias.n25 gnd 0.070538f
C5313 commonsourceibias.n26 gnd 0.009462f
C5314 commonsourceibias.t46 gnd 0.176786f
C5315 commonsourceibias.n27 gnd 0.070538f
C5316 commonsourceibias.n28 gnd 0.009462f
C5317 commonsourceibias.t52 gnd 0.176786f
C5318 commonsourceibias.n29 gnd 0.070538f
C5319 commonsourceibias.n30 gnd 0.009462f
C5320 commonsourceibias.t2 gnd 0.176786f
C5321 commonsourceibias.n31 gnd 0.010756f
C5322 commonsourceibias.n32 gnd 0.009462f
C5323 commonsourceibias.t16 gnd 0.176786f
C5324 commonsourceibias.n33 gnd 0.012719f
C5325 commonsourceibias.t48 gnd 0.196936f
C5326 commonsourceibias.t30 gnd 0.176786f
C5327 commonsourceibias.n34 gnd 0.078597f
C5328 commonsourceibias.n35 gnd 0.084205f
C5329 commonsourceibias.n36 gnd 0.040277f
C5330 commonsourceibias.n37 gnd 0.009462f
C5331 commonsourceibias.n38 gnd 0.007691f
C5332 commonsourceibias.n39 gnd 0.013039f
C5333 commonsourceibias.n40 gnd 0.070538f
C5334 commonsourceibias.n41 gnd 0.013095f
C5335 commonsourceibias.n42 gnd 0.009462f
C5336 commonsourceibias.n43 gnd 0.009462f
C5337 commonsourceibias.n44 gnd 0.009462f
C5338 commonsourceibias.n45 gnd 0.009599f
C5339 commonsourceibias.n46 gnd 0.070538f
C5340 commonsourceibias.n47 gnd 0.011663f
C5341 commonsourceibias.n48 gnd 0.012902f
C5342 commonsourceibias.n49 gnd 0.009462f
C5343 commonsourceibias.n50 gnd 0.009462f
C5344 commonsourceibias.n51 gnd 0.012818f
C5345 commonsourceibias.n52 gnd 0.007654f
C5346 commonsourceibias.n53 gnd 0.012977f
C5347 commonsourceibias.n54 gnd 0.009462f
C5348 commonsourceibias.n55 gnd 0.009462f
C5349 commonsourceibias.n56 gnd 0.013056f
C5350 commonsourceibias.n57 gnd 0.011258f
C5351 commonsourceibias.n58 gnd 0.009135f
C5352 commonsourceibias.n59 gnd 0.009462f
C5353 commonsourceibias.n60 gnd 0.009462f
C5354 commonsourceibias.n61 gnd 0.011574f
C5355 commonsourceibias.n62 gnd 0.012991f
C5356 commonsourceibias.n63 gnd 0.070538f
C5357 commonsourceibias.n64 gnd 0.012903f
C5358 commonsourceibias.n65 gnd 0.009462f
C5359 commonsourceibias.n66 gnd 0.009462f
C5360 commonsourceibias.n67 gnd 0.009462f
C5361 commonsourceibias.n68 gnd 0.012903f
C5362 commonsourceibias.n69 gnd 0.070538f
C5363 commonsourceibias.n70 gnd 0.012991f
C5364 commonsourceibias.n71 gnd 0.011574f
C5365 commonsourceibias.n72 gnd 0.009462f
C5366 commonsourceibias.n73 gnd 0.009462f
C5367 commonsourceibias.n74 gnd 0.009462f
C5368 commonsourceibias.n75 gnd 0.011258f
C5369 commonsourceibias.n76 gnd 0.013056f
C5370 commonsourceibias.n77 gnd 0.070538f
C5371 commonsourceibias.n78 gnd 0.012977f
C5372 commonsourceibias.n79 gnd 0.009462f
C5373 commonsourceibias.n80 gnd 0.009462f
C5374 commonsourceibias.n81 gnd 0.009462f
C5375 commonsourceibias.n82 gnd 0.012818f
C5376 commonsourceibias.n83 gnd 0.070538f
C5377 commonsourceibias.n84 gnd 0.012902f
C5378 commonsourceibias.n85 gnd 0.011663f
C5379 commonsourceibias.n86 gnd 0.009462f
C5380 commonsourceibias.n87 gnd 0.009462f
C5381 commonsourceibias.n88 gnd 0.009462f
C5382 commonsourceibias.n89 gnd 0.010756f
C5383 commonsourceibias.n90 gnd 0.013095f
C5384 commonsourceibias.n91 gnd 0.070538f
C5385 commonsourceibias.n92 gnd 0.013039f
C5386 commonsourceibias.n93 gnd 0.009462f
C5387 commonsourceibias.n94 gnd 0.009462f
C5388 commonsourceibias.n95 gnd 0.009462f
C5389 commonsourceibias.n96 gnd 0.012719f
C5390 commonsourceibias.n97 gnd 0.070538f
C5391 commonsourceibias.n98 gnd 0.01275f
C5392 commonsourceibias.n99 gnd 0.085058f
C5393 commonsourceibias.n100 gnd 0.095108f
C5394 commonsourceibias.t37 gnd 0.020419f
C5395 commonsourceibias.t33 gnd 0.020419f
C5396 commonsourceibias.n101 gnd 0.180428f
C5397 commonsourceibias.n102 gnd 0.15629f
C5398 commonsourceibias.t43 gnd 0.020419f
C5399 commonsourceibias.t21 gnd 0.020419f
C5400 commonsourceibias.n103 gnd 0.180428f
C5401 commonsourceibias.n104 gnd 0.082878f
C5402 commonsourceibias.t1 gnd 0.020419f
C5403 commonsourceibias.t39 gnd 0.020419f
C5404 commonsourceibias.n105 gnd 0.180428f
C5405 commonsourceibias.n106 gnd 0.082878f
C5406 commonsourceibias.t51 gnd 0.020419f
C5407 commonsourceibias.t59 gnd 0.020419f
C5408 commonsourceibias.n107 gnd 0.180428f
C5409 commonsourceibias.n108 gnd 0.06924f
C5410 commonsourceibias.t31 gnd 0.020419f
C5411 commonsourceibias.t49 gnd 0.020419f
C5412 commonsourceibias.n109 gnd 0.181032f
C5413 commonsourceibias.t3 gnd 0.020419f
C5414 commonsourceibias.t17 gnd 0.020419f
C5415 commonsourceibias.n110 gnd 0.180428f
C5416 commonsourceibias.n111 gnd 0.168125f
C5417 commonsourceibias.t47 gnd 0.020419f
C5418 commonsourceibias.t53 gnd 0.020419f
C5419 commonsourceibias.n112 gnd 0.180428f
C5420 commonsourceibias.n113 gnd 0.082878f
C5421 commonsourceibias.t25 gnd 0.020419f
C5422 commonsourceibias.t5 gnd 0.020419f
C5423 commonsourceibias.n114 gnd 0.180428f
C5424 commonsourceibias.n115 gnd 0.06924f
C5425 commonsourceibias.n116 gnd 0.083843f
C5426 commonsourceibias.n117 gnd 0.009462f
C5427 commonsourceibias.t154 gnd 0.176786f
C5428 commonsourceibias.t106 gnd 0.176786f
C5429 commonsourceibias.n118 gnd 0.070538f
C5430 commonsourceibias.n119 gnd 0.009462f
C5431 commonsourceibias.t92 gnd 0.176786f
C5432 commonsourceibias.n120 gnd 0.070538f
C5433 commonsourceibias.n121 gnd 0.009462f
C5434 commonsourceibias.t123 gnd 0.176786f
C5435 commonsourceibias.n122 gnd 0.070538f
C5436 commonsourceibias.n123 gnd 0.009462f
C5437 commonsourceibias.t110 gnd 0.176786f
C5438 commonsourceibias.n124 gnd 0.010756f
C5439 commonsourceibias.n125 gnd 0.009462f
C5440 commonsourceibias.t82 gnd 0.176786f
C5441 commonsourceibias.n126 gnd 0.012719f
C5442 commonsourceibias.t132 gnd 0.196936f
C5443 commonsourceibias.t147 gnd 0.176786f
C5444 commonsourceibias.n127 gnd 0.078597f
C5445 commonsourceibias.n128 gnd 0.084205f
C5446 commonsourceibias.n129 gnd 0.040277f
C5447 commonsourceibias.n130 gnd 0.009462f
C5448 commonsourceibias.n131 gnd 0.007691f
C5449 commonsourceibias.n132 gnd 0.013039f
C5450 commonsourceibias.n133 gnd 0.070538f
C5451 commonsourceibias.n134 gnd 0.013095f
C5452 commonsourceibias.n135 gnd 0.009462f
C5453 commonsourceibias.n136 gnd 0.009462f
C5454 commonsourceibias.n137 gnd 0.009462f
C5455 commonsourceibias.n138 gnd 0.009599f
C5456 commonsourceibias.n139 gnd 0.070538f
C5457 commonsourceibias.n140 gnd 0.011663f
C5458 commonsourceibias.n141 gnd 0.012902f
C5459 commonsourceibias.n142 gnd 0.009462f
C5460 commonsourceibias.n143 gnd 0.009462f
C5461 commonsourceibias.n144 gnd 0.012818f
C5462 commonsourceibias.n145 gnd 0.007654f
C5463 commonsourceibias.n146 gnd 0.012977f
C5464 commonsourceibias.n147 gnd 0.009462f
C5465 commonsourceibias.n148 gnd 0.009462f
C5466 commonsourceibias.n149 gnd 0.013056f
C5467 commonsourceibias.n150 gnd 0.011258f
C5468 commonsourceibias.n151 gnd 0.009135f
C5469 commonsourceibias.n152 gnd 0.009462f
C5470 commonsourceibias.n153 gnd 0.009462f
C5471 commonsourceibias.n154 gnd 0.011574f
C5472 commonsourceibias.n155 gnd 0.012991f
C5473 commonsourceibias.n156 gnd 0.070538f
C5474 commonsourceibias.n157 gnd 0.012903f
C5475 commonsourceibias.n158 gnd 0.009417f
C5476 commonsourceibias.n159 gnd 0.068402f
C5477 commonsourceibias.n160 gnd 0.009417f
C5478 commonsourceibias.n161 gnd 0.012903f
C5479 commonsourceibias.n162 gnd 0.070538f
C5480 commonsourceibias.n163 gnd 0.012991f
C5481 commonsourceibias.n164 gnd 0.011574f
C5482 commonsourceibias.n165 gnd 0.009462f
C5483 commonsourceibias.n166 gnd 0.009462f
C5484 commonsourceibias.n167 gnd 0.009462f
C5485 commonsourceibias.n168 gnd 0.011258f
C5486 commonsourceibias.n169 gnd 0.013056f
C5487 commonsourceibias.n170 gnd 0.070538f
C5488 commonsourceibias.n171 gnd 0.012977f
C5489 commonsourceibias.n172 gnd 0.009462f
C5490 commonsourceibias.n173 gnd 0.009462f
C5491 commonsourceibias.n174 gnd 0.009462f
C5492 commonsourceibias.n175 gnd 0.012818f
C5493 commonsourceibias.n176 gnd 0.070538f
C5494 commonsourceibias.n177 gnd 0.012902f
C5495 commonsourceibias.n178 gnd 0.011663f
C5496 commonsourceibias.n179 gnd 0.009462f
C5497 commonsourceibias.n180 gnd 0.009462f
C5498 commonsourceibias.n181 gnd 0.009462f
C5499 commonsourceibias.n182 gnd 0.010756f
C5500 commonsourceibias.n183 gnd 0.013095f
C5501 commonsourceibias.n184 gnd 0.070538f
C5502 commonsourceibias.n185 gnd 0.013039f
C5503 commonsourceibias.n186 gnd 0.009462f
C5504 commonsourceibias.n187 gnd 0.009462f
C5505 commonsourceibias.n188 gnd 0.009462f
C5506 commonsourceibias.n189 gnd 0.012719f
C5507 commonsourceibias.n190 gnd 0.070538f
C5508 commonsourceibias.n191 gnd 0.01275f
C5509 commonsourceibias.n192 gnd 0.085058f
C5510 commonsourceibias.n193 gnd 0.056191f
C5511 commonsourceibias.n194 gnd 0.012626f
C5512 commonsourceibias.t115 gnd 0.191194f
C5513 commonsourceibias.t138 gnd 0.176786f
C5514 commonsourceibias.n195 gnd 0.007691f
C5515 commonsourceibias.n196 gnd 0.009462f
C5516 commonsourceibias.t128 gnd 0.176786f
C5517 commonsourceibias.n197 gnd 0.009599f
C5518 commonsourceibias.n198 gnd 0.009462f
C5519 commonsourceibias.t116 gnd 0.176786f
C5520 commonsourceibias.n199 gnd 0.070538f
C5521 commonsourceibias.t139 gnd 0.176786f
C5522 commonsourceibias.n200 gnd 0.007654f
C5523 commonsourceibias.n201 gnd 0.009462f
C5524 commonsourceibias.t126 gnd 0.176786f
C5525 commonsourceibias.n202 gnd 0.009135f
C5526 commonsourceibias.n203 gnd 0.009462f
C5527 commonsourceibias.t114 gnd 0.176786f
C5528 commonsourceibias.n204 gnd 0.070538f
C5529 commonsourceibias.t140 gnd 0.176786f
C5530 commonsourceibias.n205 gnd 0.007642f
C5531 commonsourceibias.n206 gnd 0.009462f
C5532 commonsourceibias.t127 gnd 0.176786f
C5533 commonsourceibias.t149 gnd 0.176786f
C5534 commonsourceibias.n207 gnd 0.070538f
C5535 commonsourceibias.n208 gnd 0.009462f
C5536 commonsourceibias.t141 gnd 0.176786f
C5537 commonsourceibias.n209 gnd 0.070538f
C5538 commonsourceibias.n210 gnd 0.009462f
C5539 commonsourceibias.t125 gnd 0.176786f
C5540 commonsourceibias.n211 gnd 0.070538f
C5541 commonsourceibias.n212 gnd 0.009462f
C5542 commonsourceibias.t152 gnd 0.176786f
C5543 commonsourceibias.n213 gnd 0.010756f
C5544 commonsourceibias.n214 gnd 0.009462f
C5545 commonsourceibias.t69 gnd 0.176786f
C5546 commonsourceibias.n215 gnd 0.012719f
C5547 commonsourceibias.t64 gnd 0.196936f
C5548 commonsourceibias.t135 gnd 0.176786f
C5549 commonsourceibias.n216 gnd 0.078597f
C5550 commonsourceibias.n217 gnd 0.084205f
C5551 commonsourceibias.n218 gnd 0.040277f
C5552 commonsourceibias.n219 gnd 0.009462f
C5553 commonsourceibias.n220 gnd 0.007691f
C5554 commonsourceibias.n221 gnd 0.013039f
C5555 commonsourceibias.n222 gnd 0.070538f
C5556 commonsourceibias.n223 gnd 0.013095f
C5557 commonsourceibias.n224 gnd 0.009462f
C5558 commonsourceibias.n225 gnd 0.009462f
C5559 commonsourceibias.n226 gnd 0.009462f
C5560 commonsourceibias.n227 gnd 0.009599f
C5561 commonsourceibias.n228 gnd 0.070538f
C5562 commonsourceibias.n229 gnd 0.011663f
C5563 commonsourceibias.n230 gnd 0.012902f
C5564 commonsourceibias.n231 gnd 0.009462f
C5565 commonsourceibias.n232 gnd 0.009462f
C5566 commonsourceibias.n233 gnd 0.012818f
C5567 commonsourceibias.n234 gnd 0.007654f
C5568 commonsourceibias.n235 gnd 0.012977f
C5569 commonsourceibias.n236 gnd 0.009462f
C5570 commonsourceibias.n237 gnd 0.009462f
C5571 commonsourceibias.n238 gnd 0.013056f
C5572 commonsourceibias.n239 gnd 0.011258f
C5573 commonsourceibias.n240 gnd 0.009135f
C5574 commonsourceibias.n241 gnd 0.009462f
C5575 commonsourceibias.n242 gnd 0.009462f
C5576 commonsourceibias.n243 gnd 0.011574f
C5577 commonsourceibias.n244 gnd 0.012991f
C5578 commonsourceibias.n245 gnd 0.070538f
C5579 commonsourceibias.n246 gnd 0.012903f
C5580 commonsourceibias.n247 gnd 0.009462f
C5581 commonsourceibias.n248 gnd 0.009462f
C5582 commonsourceibias.n249 gnd 0.009462f
C5583 commonsourceibias.n250 gnd 0.012903f
C5584 commonsourceibias.n251 gnd 0.070538f
C5585 commonsourceibias.n252 gnd 0.012991f
C5586 commonsourceibias.n253 gnd 0.011574f
C5587 commonsourceibias.n254 gnd 0.009462f
C5588 commonsourceibias.n255 gnd 0.009462f
C5589 commonsourceibias.n256 gnd 0.009462f
C5590 commonsourceibias.n257 gnd 0.011258f
C5591 commonsourceibias.n258 gnd 0.013056f
C5592 commonsourceibias.n259 gnd 0.070538f
C5593 commonsourceibias.n260 gnd 0.012977f
C5594 commonsourceibias.n261 gnd 0.009462f
C5595 commonsourceibias.n262 gnd 0.009462f
C5596 commonsourceibias.n263 gnd 0.009462f
C5597 commonsourceibias.n264 gnd 0.012818f
C5598 commonsourceibias.n265 gnd 0.070538f
C5599 commonsourceibias.n266 gnd 0.012902f
C5600 commonsourceibias.n267 gnd 0.011663f
C5601 commonsourceibias.n268 gnd 0.009462f
C5602 commonsourceibias.n269 gnd 0.009462f
C5603 commonsourceibias.n270 gnd 0.009462f
C5604 commonsourceibias.n271 gnd 0.010756f
C5605 commonsourceibias.n272 gnd 0.013095f
C5606 commonsourceibias.n273 gnd 0.070538f
C5607 commonsourceibias.n274 gnd 0.013039f
C5608 commonsourceibias.n275 gnd 0.009462f
C5609 commonsourceibias.n276 gnd 0.009462f
C5610 commonsourceibias.n277 gnd 0.009462f
C5611 commonsourceibias.n278 gnd 0.012719f
C5612 commonsourceibias.n279 gnd 0.070538f
C5613 commonsourceibias.n280 gnd 0.01275f
C5614 commonsourceibias.n281 gnd 0.085058f
C5615 commonsourceibias.n282 gnd 0.030353f
C5616 commonsourceibias.n283 gnd 0.151535f
C5617 commonsourceibias.n284 gnd 0.012626f
C5618 commonsourceibias.t68 gnd 0.176786f
C5619 commonsourceibias.n285 gnd 0.007691f
C5620 commonsourceibias.n286 gnd 0.009462f
C5621 commonsourceibias.t80 gnd 0.176786f
C5622 commonsourceibias.n287 gnd 0.009599f
C5623 commonsourceibias.n288 gnd 0.009462f
C5624 commonsourceibias.t134 gnd 0.176786f
C5625 commonsourceibias.n289 gnd 0.070538f
C5626 commonsourceibias.t159 gnd 0.176786f
C5627 commonsourceibias.n290 gnd 0.007654f
C5628 commonsourceibias.n291 gnd 0.009462f
C5629 commonsourceibias.t74 gnd 0.176786f
C5630 commonsourceibias.n292 gnd 0.009135f
C5631 commonsourceibias.n293 gnd 0.009462f
C5632 commonsourceibias.t120 gnd 0.176786f
C5633 commonsourceibias.n294 gnd 0.070538f
C5634 commonsourceibias.t111 gnd 0.176786f
C5635 commonsourceibias.n295 gnd 0.007642f
C5636 commonsourceibias.n296 gnd 0.009462f
C5637 commonsourceibias.t67 gnd 0.176786f
C5638 commonsourceibias.t81 gnd 0.176786f
C5639 commonsourceibias.n297 gnd 0.070538f
C5640 commonsourceibias.n298 gnd 0.009462f
C5641 commonsourceibias.t101 gnd 0.176786f
C5642 commonsourceibias.n299 gnd 0.070538f
C5643 commonsourceibias.n300 gnd 0.009462f
C5644 commonsourceibias.t158 gnd 0.176786f
C5645 commonsourceibias.n301 gnd 0.070538f
C5646 commonsourceibias.n302 gnd 0.009462f
C5647 commonsourceibias.t150 gnd 0.176786f
C5648 commonsourceibias.n303 gnd 0.010756f
C5649 commonsourceibias.n304 gnd 0.009462f
C5650 commonsourceibias.t70 gnd 0.176786f
C5651 commonsourceibias.n305 gnd 0.012719f
C5652 commonsourceibias.t136 gnd 0.196936f
C5653 commonsourceibias.t143 gnd 0.176786f
C5654 commonsourceibias.n306 gnd 0.078597f
C5655 commonsourceibias.n307 gnd 0.084205f
C5656 commonsourceibias.n308 gnd 0.040277f
C5657 commonsourceibias.n309 gnd 0.009462f
C5658 commonsourceibias.n310 gnd 0.007691f
C5659 commonsourceibias.n311 gnd 0.013039f
C5660 commonsourceibias.n312 gnd 0.070538f
C5661 commonsourceibias.n313 gnd 0.013095f
C5662 commonsourceibias.n314 gnd 0.009462f
C5663 commonsourceibias.n315 gnd 0.009462f
C5664 commonsourceibias.n316 gnd 0.009462f
C5665 commonsourceibias.n317 gnd 0.009599f
C5666 commonsourceibias.n318 gnd 0.070538f
C5667 commonsourceibias.n319 gnd 0.011663f
C5668 commonsourceibias.n320 gnd 0.012902f
C5669 commonsourceibias.n321 gnd 0.009462f
C5670 commonsourceibias.n322 gnd 0.009462f
C5671 commonsourceibias.n323 gnd 0.012818f
C5672 commonsourceibias.n324 gnd 0.007654f
C5673 commonsourceibias.n325 gnd 0.012977f
C5674 commonsourceibias.n326 gnd 0.009462f
C5675 commonsourceibias.n327 gnd 0.009462f
C5676 commonsourceibias.n328 gnd 0.013056f
C5677 commonsourceibias.n329 gnd 0.011258f
C5678 commonsourceibias.n330 gnd 0.009135f
C5679 commonsourceibias.n331 gnd 0.009462f
C5680 commonsourceibias.n332 gnd 0.009462f
C5681 commonsourceibias.n333 gnd 0.011574f
C5682 commonsourceibias.n334 gnd 0.012991f
C5683 commonsourceibias.n335 gnd 0.070538f
C5684 commonsourceibias.n336 gnd 0.012903f
C5685 commonsourceibias.n337 gnd 0.009462f
C5686 commonsourceibias.n338 gnd 0.009462f
C5687 commonsourceibias.n339 gnd 0.009462f
C5688 commonsourceibias.n340 gnd 0.012903f
C5689 commonsourceibias.n341 gnd 0.070538f
C5690 commonsourceibias.n342 gnd 0.012991f
C5691 commonsourceibias.n343 gnd 0.011574f
C5692 commonsourceibias.n344 gnd 0.009462f
C5693 commonsourceibias.n345 gnd 0.009462f
C5694 commonsourceibias.n346 gnd 0.009462f
C5695 commonsourceibias.n347 gnd 0.011258f
C5696 commonsourceibias.n348 gnd 0.013056f
C5697 commonsourceibias.n349 gnd 0.070538f
C5698 commonsourceibias.n350 gnd 0.012977f
C5699 commonsourceibias.n351 gnd 0.009462f
C5700 commonsourceibias.n352 gnd 0.009462f
C5701 commonsourceibias.n353 gnd 0.009462f
C5702 commonsourceibias.n354 gnd 0.012818f
C5703 commonsourceibias.n355 gnd 0.070538f
C5704 commonsourceibias.n356 gnd 0.012902f
C5705 commonsourceibias.n357 gnd 0.011663f
C5706 commonsourceibias.n358 gnd 0.009462f
C5707 commonsourceibias.n359 gnd 0.009462f
C5708 commonsourceibias.n360 gnd 0.009462f
C5709 commonsourceibias.n361 gnd 0.010756f
C5710 commonsourceibias.n362 gnd 0.013095f
C5711 commonsourceibias.n363 gnd 0.070538f
C5712 commonsourceibias.n364 gnd 0.013039f
C5713 commonsourceibias.n365 gnd 0.009462f
C5714 commonsourceibias.n366 gnd 0.009462f
C5715 commonsourceibias.n367 gnd 0.009462f
C5716 commonsourceibias.n368 gnd 0.012719f
C5717 commonsourceibias.n369 gnd 0.070538f
C5718 commonsourceibias.n370 gnd 0.01275f
C5719 commonsourceibias.t148 gnd 0.191194f
C5720 commonsourceibias.n371 gnd 0.085058f
C5721 commonsourceibias.n372 gnd 0.030353f
C5722 commonsourceibias.n373 gnd 0.53129f
C5723 commonsourceibias.n374 gnd 0.012626f
C5724 commonsourceibias.t153 gnd 0.191194f
C5725 commonsourceibias.t104 gnd 0.176786f
C5726 commonsourceibias.n375 gnd 0.007691f
C5727 commonsourceibias.n376 gnd 0.009462f
C5728 commonsourceibias.t73 gnd 0.176786f
C5729 commonsourceibias.n377 gnd 0.009599f
C5730 commonsourceibias.n378 gnd 0.009462f
C5731 commonsourceibias.t90 gnd 0.176786f
C5732 commonsourceibias.n379 gnd 0.007654f
C5733 commonsourceibias.n380 gnd 0.009462f
C5734 commonsourceibias.t151 gnd 0.176786f
C5735 commonsourceibias.n381 gnd 0.009135f
C5736 commonsourceibias.n382 gnd 0.009462f
C5737 commonsourceibias.t91 gnd 0.176786f
C5738 commonsourceibias.n383 gnd 0.007642f
C5739 commonsourceibias.n384 gnd 0.009462f
C5740 commonsourceibias.t119 gnd 0.176786f
C5741 commonsourceibias.t87 gnd 0.176786f
C5742 commonsourceibias.n385 gnd 0.070538f
C5743 commonsourceibias.n386 gnd 0.009462f
C5744 commonsourceibias.t79 gnd 0.176786f
C5745 commonsourceibias.n387 gnd 0.070538f
C5746 commonsourceibias.n388 gnd 0.009462f
C5747 commonsourceibias.t95 gnd 0.176786f
C5748 commonsourceibias.n389 gnd 0.070538f
C5749 commonsourceibias.n390 gnd 0.009462f
C5750 commonsourceibias.t88 gnd 0.176786f
C5751 commonsourceibias.n391 gnd 0.010756f
C5752 commonsourceibias.n392 gnd 0.009462f
C5753 commonsourceibias.t65 gnd 0.176786f
C5754 commonsourceibias.n393 gnd 0.012719f
C5755 commonsourceibias.t83 gnd 0.196936f
C5756 commonsourceibias.t84 gnd 0.176786f
C5757 commonsourceibias.n394 gnd 0.078597f
C5758 commonsourceibias.n395 gnd 0.084205f
C5759 commonsourceibias.n396 gnd 0.040277f
C5760 commonsourceibias.n397 gnd 0.009462f
C5761 commonsourceibias.n398 gnd 0.007691f
C5762 commonsourceibias.n399 gnd 0.013039f
C5763 commonsourceibias.n400 gnd 0.070538f
C5764 commonsourceibias.n401 gnd 0.013095f
C5765 commonsourceibias.n402 gnd 0.009462f
C5766 commonsourceibias.n403 gnd 0.009462f
C5767 commonsourceibias.n404 gnd 0.009462f
C5768 commonsourceibias.n405 gnd 0.009599f
C5769 commonsourceibias.n406 gnd 0.070538f
C5770 commonsourceibias.n407 gnd 0.011663f
C5771 commonsourceibias.n408 gnd 0.012902f
C5772 commonsourceibias.n409 gnd 0.009462f
C5773 commonsourceibias.n410 gnd 0.009462f
C5774 commonsourceibias.n411 gnd 0.012818f
C5775 commonsourceibias.n412 gnd 0.007654f
C5776 commonsourceibias.n413 gnd 0.012977f
C5777 commonsourceibias.n414 gnd 0.009462f
C5778 commonsourceibias.n415 gnd 0.009462f
C5779 commonsourceibias.n416 gnd 0.013056f
C5780 commonsourceibias.n417 gnd 0.011258f
C5781 commonsourceibias.n418 gnd 0.009135f
C5782 commonsourceibias.n419 gnd 0.009462f
C5783 commonsourceibias.n420 gnd 0.009462f
C5784 commonsourceibias.n421 gnd 0.011574f
C5785 commonsourceibias.n422 gnd 0.012991f
C5786 commonsourceibias.n423 gnd 0.070538f
C5787 commonsourceibias.n424 gnd 0.012903f
C5788 commonsourceibias.n425 gnd 0.009417f
C5789 commonsourceibias.t15 gnd 0.020419f
C5790 commonsourceibias.t13 gnd 0.020419f
C5791 commonsourceibias.n426 gnd 0.181032f
C5792 commonsourceibias.t19 gnd 0.020419f
C5793 commonsourceibias.t9 gnd 0.020419f
C5794 commonsourceibias.n427 gnd 0.180428f
C5795 commonsourceibias.n428 gnd 0.168125f
C5796 commonsourceibias.t45 gnd 0.020419f
C5797 commonsourceibias.t35 gnd 0.020419f
C5798 commonsourceibias.n429 gnd 0.180428f
C5799 commonsourceibias.n430 gnd 0.082878f
C5800 commonsourceibias.t11 gnd 0.020419f
C5801 commonsourceibias.t57 gnd 0.020419f
C5802 commonsourceibias.n431 gnd 0.180428f
C5803 commonsourceibias.n432 gnd 0.06924f
C5804 commonsourceibias.n433 gnd 0.012626f
C5805 commonsourceibias.t6 gnd 0.176786f
C5806 commonsourceibias.n434 gnd 0.007691f
C5807 commonsourceibias.n435 gnd 0.009462f
C5808 commonsourceibias.t40 gnd 0.176786f
C5809 commonsourceibias.n436 gnd 0.009599f
C5810 commonsourceibias.n437 gnd 0.009462f
C5811 commonsourceibias.t62 gnd 0.176786f
C5812 commonsourceibias.n438 gnd 0.007654f
C5813 commonsourceibias.n439 gnd 0.009462f
C5814 commonsourceibias.t28 gnd 0.176786f
C5815 commonsourceibias.n440 gnd 0.009135f
C5816 commonsourceibias.n441 gnd 0.009462f
C5817 commonsourceibias.t60 gnd 0.176786f
C5818 commonsourceibias.n442 gnd 0.007642f
C5819 commonsourceibias.n443 gnd 0.009462f
C5820 commonsourceibias.t56 gnd 0.176786f
C5821 commonsourceibias.t10 gnd 0.176786f
C5822 commonsourceibias.n444 gnd 0.070538f
C5823 commonsourceibias.n445 gnd 0.009462f
C5824 commonsourceibias.t34 gnd 0.176786f
C5825 commonsourceibias.n446 gnd 0.070538f
C5826 commonsourceibias.n447 gnd 0.009462f
C5827 commonsourceibias.t44 gnd 0.176786f
C5828 commonsourceibias.n448 gnd 0.070538f
C5829 commonsourceibias.n449 gnd 0.009462f
C5830 commonsourceibias.t8 gnd 0.176786f
C5831 commonsourceibias.n450 gnd 0.010756f
C5832 commonsourceibias.n451 gnd 0.009462f
C5833 commonsourceibias.t18 gnd 0.176786f
C5834 commonsourceibias.n452 gnd 0.012719f
C5835 commonsourceibias.t14 gnd 0.196936f
C5836 commonsourceibias.t12 gnd 0.176786f
C5837 commonsourceibias.n453 gnd 0.078597f
C5838 commonsourceibias.n454 gnd 0.084205f
C5839 commonsourceibias.n455 gnd 0.040277f
C5840 commonsourceibias.n456 gnd 0.009462f
C5841 commonsourceibias.n457 gnd 0.007691f
C5842 commonsourceibias.n458 gnd 0.013039f
C5843 commonsourceibias.n459 gnd 0.070538f
C5844 commonsourceibias.n460 gnd 0.013095f
C5845 commonsourceibias.n461 gnd 0.009462f
C5846 commonsourceibias.n462 gnd 0.009462f
C5847 commonsourceibias.n463 gnd 0.009462f
C5848 commonsourceibias.n464 gnd 0.009599f
C5849 commonsourceibias.n465 gnd 0.070538f
C5850 commonsourceibias.n466 gnd 0.011663f
C5851 commonsourceibias.n467 gnd 0.012902f
C5852 commonsourceibias.n468 gnd 0.009462f
C5853 commonsourceibias.n469 gnd 0.009462f
C5854 commonsourceibias.n470 gnd 0.012818f
C5855 commonsourceibias.n471 gnd 0.007654f
C5856 commonsourceibias.n472 gnd 0.012977f
C5857 commonsourceibias.n473 gnd 0.009462f
C5858 commonsourceibias.n474 gnd 0.009462f
C5859 commonsourceibias.n475 gnd 0.013056f
C5860 commonsourceibias.n476 gnd 0.011258f
C5861 commonsourceibias.n477 gnd 0.009135f
C5862 commonsourceibias.n478 gnd 0.009462f
C5863 commonsourceibias.n479 gnd 0.009462f
C5864 commonsourceibias.n480 gnd 0.011574f
C5865 commonsourceibias.n481 gnd 0.012991f
C5866 commonsourceibias.n482 gnd 0.070538f
C5867 commonsourceibias.n483 gnd 0.012903f
C5868 commonsourceibias.n484 gnd 0.009462f
C5869 commonsourceibias.n485 gnd 0.009462f
C5870 commonsourceibias.n486 gnd 0.009462f
C5871 commonsourceibias.n487 gnd 0.012903f
C5872 commonsourceibias.n488 gnd 0.070538f
C5873 commonsourceibias.n489 gnd 0.012991f
C5874 commonsourceibias.t22 gnd 0.176786f
C5875 commonsourceibias.n490 gnd 0.070538f
C5876 commonsourceibias.n491 gnd 0.011574f
C5877 commonsourceibias.n492 gnd 0.009462f
C5878 commonsourceibias.n493 gnd 0.009462f
C5879 commonsourceibias.n494 gnd 0.009462f
C5880 commonsourceibias.n495 gnd 0.011258f
C5881 commonsourceibias.n496 gnd 0.013056f
C5882 commonsourceibias.n497 gnd 0.070538f
C5883 commonsourceibias.n498 gnd 0.012977f
C5884 commonsourceibias.n499 gnd 0.009462f
C5885 commonsourceibias.n500 gnd 0.009462f
C5886 commonsourceibias.n501 gnd 0.009462f
C5887 commonsourceibias.n502 gnd 0.012818f
C5888 commonsourceibias.n503 gnd 0.070538f
C5889 commonsourceibias.n504 gnd 0.012902f
C5890 commonsourceibias.t54 gnd 0.176786f
C5891 commonsourceibias.n505 gnd 0.070538f
C5892 commonsourceibias.n506 gnd 0.011663f
C5893 commonsourceibias.n507 gnd 0.009462f
C5894 commonsourceibias.n508 gnd 0.009462f
C5895 commonsourceibias.n509 gnd 0.009462f
C5896 commonsourceibias.n510 gnd 0.010756f
C5897 commonsourceibias.n511 gnd 0.013095f
C5898 commonsourceibias.n512 gnd 0.070538f
C5899 commonsourceibias.n513 gnd 0.013039f
C5900 commonsourceibias.n514 gnd 0.009462f
C5901 commonsourceibias.n515 gnd 0.009462f
C5902 commonsourceibias.n516 gnd 0.009462f
C5903 commonsourceibias.n517 gnd 0.012719f
C5904 commonsourceibias.n518 gnd 0.070538f
C5905 commonsourceibias.n519 gnd 0.01275f
C5906 commonsourceibias.t26 gnd 0.191194f
C5907 commonsourceibias.n520 gnd 0.085058f
C5908 commonsourceibias.n521 gnd 0.095108f
C5909 commonsourceibias.t7 gnd 0.020419f
C5910 commonsourceibias.t27 gnd 0.020419f
C5911 commonsourceibias.n522 gnd 0.180428f
C5912 commonsourceibias.n523 gnd 0.15629f
C5913 commonsourceibias.t55 gnd 0.020419f
C5914 commonsourceibias.t41 gnd 0.020419f
C5915 commonsourceibias.n524 gnd 0.180428f
C5916 commonsourceibias.n525 gnd 0.082878f
C5917 commonsourceibias.t29 gnd 0.020419f
C5918 commonsourceibias.t63 gnd 0.020419f
C5919 commonsourceibias.n526 gnd 0.180428f
C5920 commonsourceibias.n527 gnd 0.082878f
C5921 commonsourceibias.t61 gnd 0.020419f
C5922 commonsourceibias.t23 gnd 0.020419f
C5923 commonsourceibias.n528 gnd 0.180428f
C5924 commonsourceibias.n529 gnd 0.06924f
C5925 commonsourceibias.n530 gnd 0.083843f
C5926 commonsourceibias.n531 gnd 0.068402f
C5927 commonsourceibias.n532 gnd 0.009417f
C5928 commonsourceibias.n533 gnd 0.012903f
C5929 commonsourceibias.n534 gnd 0.070538f
C5930 commonsourceibias.n535 gnd 0.012991f
C5931 commonsourceibias.t102 gnd 0.176786f
C5932 commonsourceibias.n536 gnd 0.070538f
C5933 commonsourceibias.n537 gnd 0.011574f
C5934 commonsourceibias.n538 gnd 0.009462f
C5935 commonsourceibias.n539 gnd 0.009462f
C5936 commonsourceibias.n540 gnd 0.009462f
C5937 commonsourceibias.n541 gnd 0.011258f
C5938 commonsourceibias.n542 gnd 0.013056f
C5939 commonsourceibias.n543 gnd 0.070538f
C5940 commonsourceibias.n544 gnd 0.012977f
C5941 commonsourceibias.n545 gnd 0.009462f
C5942 commonsourceibias.n546 gnd 0.009462f
C5943 commonsourceibias.n547 gnd 0.009462f
C5944 commonsourceibias.n548 gnd 0.012818f
C5945 commonsourceibias.n549 gnd 0.070538f
C5946 commonsourceibias.n550 gnd 0.012902f
C5947 commonsourceibias.t121 gnd 0.176786f
C5948 commonsourceibias.n551 gnd 0.070538f
C5949 commonsourceibias.n552 gnd 0.011663f
C5950 commonsourceibias.n553 gnd 0.009462f
C5951 commonsourceibias.n554 gnd 0.009462f
C5952 commonsourceibias.n555 gnd 0.009462f
C5953 commonsourceibias.n556 gnd 0.010756f
C5954 commonsourceibias.n557 gnd 0.013095f
C5955 commonsourceibias.n558 gnd 0.070538f
C5956 commonsourceibias.n559 gnd 0.013039f
C5957 commonsourceibias.n560 gnd 0.009462f
C5958 commonsourceibias.n561 gnd 0.009462f
C5959 commonsourceibias.n562 gnd 0.009462f
C5960 commonsourceibias.n563 gnd 0.012719f
C5961 commonsourceibias.n564 gnd 0.070538f
C5962 commonsourceibias.n565 gnd 0.01275f
C5963 commonsourceibias.n566 gnd 0.085058f
C5964 commonsourceibias.n567 gnd 0.056191f
C5965 commonsourceibias.n568 gnd 0.012626f
C5966 commonsourceibias.t118 gnd 0.176786f
C5967 commonsourceibias.n569 gnd 0.007691f
C5968 commonsourceibias.n570 gnd 0.009462f
C5969 commonsourceibias.t109 gnd 0.176786f
C5970 commonsourceibias.n571 gnd 0.009599f
C5971 commonsourceibias.n572 gnd 0.009462f
C5972 commonsourceibias.t117 gnd 0.176786f
C5973 commonsourceibias.n573 gnd 0.007654f
C5974 commonsourceibias.n574 gnd 0.009462f
C5975 commonsourceibias.t108 gnd 0.176786f
C5976 commonsourceibias.n575 gnd 0.009135f
C5977 commonsourceibias.n576 gnd 0.009462f
C5978 commonsourceibias.t122 gnd 0.176786f
C5979 commonsourceibias.n577 gnd 0.007642f
C5980 commonsourceibias.n578 gnd 0.009462f
C5981 commonsourceibias.t107 gnd 0.176786f
C5982 commonsourceibias.t129 gnd 0.176786f
C5983 commonsourceibias.n579 gnd 0.070538f
C5984 commonsourceibias.n580 gnd 0.009462f
C5985 commonsourceibias.t156 gnd 0.176786f
C5986 commonsourceibias.n581 gnd 0.070538f
C5987 commonsourceibias.n582 gnd 0.009462f
C5988 commonsourceibias.t105 gnd 0.176786f
C5989 commonsourceibias.n583 gnd 0.070538f
C5990 commonsourceibias.n584 gnd 0.009462f
C5991 commonsourceibias.t137 gnd 0.176786f
C5992 commonsourceibias.n585 gnd 0.010756f
C5993 commonsourceibias.n586 gnd 0.009462f
C5994 commonsourceibias.t155 gnd 0.176786f
C5995 commonsourceibias.n587 gnd 0.012719f
C5996 commonsourceibias.t131 gnd 0.196936f
C5997 commonsourceibias.t142 gnd 0.176786f
C5998 commonsourceibias.n588 gnd 0.078597f
C5999 commonsourceibias.n589 gnd 0.084205f
C6000 commonsourceibias.n590 gnd 0.040277f
C6001 commonsourceibias.n591 gnd 0.009462f
C6002 commonsourceibias.n592 gnd 0.007691f
C6003 commonsourceibias.n593 gnd 0.013039f
C6004 commonsourceibias.n594 gnd 0.070538f
C6005 commonsourceibias.n595 gnd 0.013095f
C6006 commonsourceibias.n596 gnd 0.009462f
C6007 commonsourceibias.n597 gnd 0.009462f
C6008 commonsourceibias.n598 gnd 0.009462f
C6009 commonsourceibias.n599 gnd 0.009599f
C6010 commonsourceibias.n600 gnd 0.070538f
C6011 commonsourceibias.n601 gnd 0.011663f
C6012 commonsourceibias.n602 gnd 0.012902f
C6013 commonsourceibias.n603 gnd 0.009462f
C6014 commonsourceibias.n604 gnd 0.009462f
C6015 commonsourceibias.n605 gnd 0.012818f
C6016 commonsourceibias.n606 gnd 0.007654f
C6017 commonsourceibias.n607 gnd 0.012977f
C6018 commonsourceibias.n608 gnd 0.009462f
C6019 commonsourceibias.n609 gnd 0.009462f
C6020 commonsourceibias.n610 gnd 0.013056f
C6021 commonsourceibias.n611 gnd 0.011258f
C6022 commonsourceibias.n612 gnd 0.009135f
C6023 commonsourceibias.n613 gnd 0.009462f
C6024 commonsourceibias.n614 gnd 0.009462f
C6025 commonsourceibias.n615 gnd 0.011574f
C6026 commonsourceibias.n616 gnd 0.012991f
C6027 commonsourceibias.n617 gnd 0.070538f
C6028 commonsourceibias.n618 gnd 0.012903f
C6029 commonsourceibias.n619 gnd 0.009462f
C6030 commonsourceibias.n620 gnd 0.009462f
C6031 commonsourceibias.n621 gnd 0.009462f
C6032 commonsourceibias.n622 gnd 0.012903f
C6033 commonsourceibias.n623 gnd 0.070538f
C6034 commonsourceibias.n624 gnd 0.012991f
C6035 commonsourceibias.t130 gnd 0.176786f
C6036 commonsourceibias.n625 gnd 0.070538f
C6037 commonsourceibias.n626 gnd 0.011574f
C6038 commonsourceibias.n627 gnd 0.009462f
C6039 commonsourceibias.n628 gnd 0.009462f
C6040 commonsourceibias.n629 gnd 0.009462f
C6041 commonsourceibias.n630 gnd 0.011258f
C6042 commonsourceibias.n631 gnd 0.013056f
C6043 commonsourceibias.n632 gnd 0.070538f
C6044 commonsourceibias.n633 gnd 0.012977f
C6045 commonsourceibias.n634 gnd 0.009462f
C6046 commonsourceibias.n635 gnd 0.009462f
C6047 commonsourceibias.n636 gnd 0.009462f
C6048 commonsourceibias.n637 gnd 0.012818f
C6049 commonsourceibias.n638 gnd 0.070538f
C6050 commonsourceibias.n639 gnd 0.012902f
C6051 commonsourceibias.t99 gnd 0.176786f
C6052 commonsourceibias.n640 gnd 0.070538f
C6053 commonsourceibias.n641 gnd 0.011663f
C6054 commonsourceibias.n642 gnd 0.009462f
C6055 commonsourceibias.n643 gnd 0.009462f
C6056 commonsourceibias.n644 gnd 0.009462f
C6057 commonsourceibias.n645 gnd 0.010756f
C6058 commonsourceibias.n646 gnd 0.013095f
C6059 commonsourceibias.n647 gnd 0.070538f
C6060 commonsourceibias.n648 gnd 0.013039f
C6061 commonsourceibias.n649 gnd 0.009462f
C6062 commonsourceibias.n650 gnd 0.009462f
C6063 commonsourceibias.n651 gnd 0.009462f
C6064 commonsourceibias.n652 gnd 0.012719f
C6065 commonsourceibias.n653 gnd 0.070538f
C6066 commonsourceibias.n654 gnd 0.01275f
C6067 commonsourceibias.t100 gnd 0.191194f
C6068 commonsourceibias.n655 gnd 0.085058f
C6069 commonsourceibias.n656 gnd 0.030353f
C6070 commonsourceibias.n657 gnd 0.151535f
C6071 commonsourceibias.n658 gnd 0.012626f
C6072 commonsourceibias.t86 gnd 0.176786f
C6073 commonsourceibias.n659 gnd 0.007691f
C6074 commonsourceibias.n660 gnd 0.009462f
C6075 commonsourceibias.t97 gnd 0.176786f
C6076 commonsourceibias.n661 gnd 0.009599f
C6077 commonsourceibias.n662 gnd 0.009462f
C6078 commonsourceibias.t77 gnd 0.176786f
C6079 commonsourceibias.n663 gnd 0.007654f
C6080 commonsourceibias.n664 gnd 0.009462f
C6081 commonsourceibias.t93 gnd 0.176786f
C6082 commonsourceibias.n665 gnd 0.009135f
C6083 commonsourceibias.n666 gnd 0.009462f
C6084 commonsourceibias.t145 gnd 0.176786f
C6085 commonsourceibias.n667 gnd 0.007642f
C6086 commonsourceibias.n668 gnd 0.009462f
C6087 commonsourceibias.t85 gnd 0.176786f
C6088 commonsourceibias.t98 gnd 0.176786f
C6089 commonsourceibias.n669 gnd 0.070538f
C6090 commonsourceibias.n670 gnd 0.009462f
C6091 commonsourceibias.t94 gnd 0.176786f
C6092 commonsourceibias.n671 gnd 0.070538f
C6093 commonsourceibias.n672 gnd 0.009462f
C6094 commonsourceibias.t76 gnd 0.176786f
C6095 commonsourceibias.n673 gnd 0.070538f
C6096 commonsourceibias.n674 gnd 0.009462f
C6097 commonsourceibias.t72 gnd 0.176786f
C6098 commonsourceibias.n675 gnd 0.010756f
C6099 commonsourceibias.n676 gnd 0.009462f
C6100 commonsourceibias.t89 gnd 0.176786f
C6101 commonsourceibias.n677 gnd 0.012719f
C6102 commonsourceibias.t144 gnd 0.196936f
C6103 commonsourceibias.t133 gnd 0.176786f
C6104 commonsourceibias.n678 gnd 0.078597f
C6105 commonsourceibias.n679 gnd 0.084205f
C6106 commonsourceibias.n680 gnd 0.040277f
C6107 commonsourceibias.n681 gnd 0.009462f
C6108 commonsourceibias.n682 gnd 0.007691f
C6109 commonsourceibias.n683 gnd 0.013039f
C6110 commonsourceibias.n684 gnd 0.070538f
C6111 commonsourceibias.n685 gnd 0.013095f
C6112 commonsourceibias.n686 gnd 0.009462f
C6113 commonsourceibias.n687 gnd 0.009462f
C6114 commonsourceibias.n688 gnd 0.009462f
C6115 commonsourceibias.n689 gnd 0.009599f
C6116 commonsourceibias.n690 gnd 0.070538f
C6117 commonsourceibias.n691 gnd 0.011663f
C6118 commonsourceibias.n692 gnd 0.012902f
C6119 commonsourceibias.n693 gnd 0.009462f
C6120 commonsourceibias.n694 gnd 0.009462f
C6121 commonsourceibias.n695 gnd 0.012818f
C6122 commonsourceibias.n696 gnd 0.007654f
C6123 commonsourceibias.n697 gnd 0.012977f
C6124 commonsourceibias.n698 gnd 0.009462f
C6125 commonsourceibias.n699 gnd 0.009462f
C6126 commonsourceibias.n700 gnd 0.013056f
C6127 commonsourceibias.n701 gnd 0.011258f
C6128 commonsourceibias.n702 gnd 0.009135f
C6129 commonsourceibias.n703 gnd 0.009462f
C6130 commonsourceibias.n704 gnd 0.009462f
C6131 commonsourceibias.n705 gnd 0.011574f
C6132 commonsourceibias.n706 gnd 0.012991f
C6133 commonsourceibias.n707 gnd 0.070538f
C6134 commonsourceibias.n708 gnd 0.012903f
C6135 commonsourceibias.n709 gnd 0.009462f
C6136 commonsourceibias.n710 gnd 0.009462f
C6137 commonsourceibias.n711 gnd 0.009462f
C6138 commonsourceibias.n712 gnd 0.012903f
C6139 commonsourceibias.n713 gnd 0.070538f
C6140 commonsourceibias.n714 gnd 0.012991f
C6141 commonsourceibias.t103 gnd 0.176786f
C6142 commonsourceibias.n715 gnd 0.070538f
C6143 commonsourceibias.n716 gnd 0.011574f
C6144 commonsourceibias.n717 gnd 0.009462f
C6145 commonsourceibias.n718 gnd 0.009462f
C6146 commonsourceibias.n719 gnd 0.009462f
C6147 commonsourceibias.n720 gnd 0.011258f
C6148 commonsourceibias.n721 gnd 0.013056f
C6149 commonsourceibias.n722 gnd 0.070538f
C6150 commonsourceibias.n723 gnd 0.012977f
C6151 commonsourceibias.n724 gnd 0.009462f
C6152 commonsourceibias.n725 gnd 0.009462f
C6153 commonsourceibias.n726 gnd 0.009462f
C6154 commonsourceibias.n727 gnd 0.012818f
C6155 commonsourceibias.n728 gnd 0.070538f
C6156 commonsourceibias.n729 gnd 0.012902f
C6157 commonsourceibias.t66 gnd 0.176786f
C6158 commonsourceibias.n730 gnd 0.070538f
C6159 commonsourceibias.n731 gnd 0.011663f
C6160 commonsourceibias.n732 gnd 0.009462f
C6161 commonsourceibias.n733 gnd 0.009462f
C6162 commonsourceibias.n734 gnd 0.009462f
C6163 commonsourceibias.n735 gnd 0.010756f
C6164 commonsourceibias.n736 gnd 0.013095f
C6165 commonsourceibias.n737 gnd 0.070538f
C6166 commonsourceibias.n738 gnd 0.013039f
C6167 commonsourceibias.n739 gnd 0.009462f
C6168 commonsourceibias.n740 gnd 0.009462f
C6169 commonsourceibias.n741 gnd 0.009462f
C6170 commonsourceibias.n742 gnd 0.012719f
C6171 commonsourceibias.n743 gnd 0.070538f
C6172 commonsourceibias.n744 gnd 0.01275f
C6173 commonsourceibias.t71 gnd 0.191194f
C6174 commonsourceibias.n745 gnd 0.085058f
C6175 commonsourceibias.n746 gnd 0.030353f
C6176 commonsourceibias.n747 gnd 0.199689f
C6177 commonsourceibias.n748 gnd 5.4246f
.ends

