* NGSPICE file created from opamp484.ext - technology: sky130A

.subckt opamp484 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 CSoutput.t182 a_n8300_8799.t36 vdd.t221 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X1 CSoutput.t186 commonsourceibias.t48 gnd.t289 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X2 a_n2140_13878.t23 a_n2318_13878.t52 vdd.t50 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 a_n2140_13878.t15 a_n2318_13878.t34 a_n2318_13878.t35 vdd.t59 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 vdd.t220 a_n8300_8799.t37 CSoutput.t181 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X5 gnd.t288 commonsourceibias.t49 CSoutput.t32 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X6 CSoutput.t60 commonsourceibias.t50 gnd.t287 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 CSoutput.t33 commonsourceibias.t51 gnd.t286 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 CSoutput.t180 a_n8300_8799.t38 vdd.t219 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X9 CSoutput.t179 a_n8300_8799.t39 vdd.t218 vdd.t78 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X10 output.t3 outputibias.t8 gnd.t320 gnd.t319 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X11 a_n2318_8322.t15 a_n2318_13878.t53 a_n8300_8799.t23 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X12 vdd.t52 CSoutput.t192 output.t19 gnd.t305 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X13 CSoutput.t178 a_n8300_8799.t40 vdd.t217 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X14 gnd.t134 gnd.t132 plus.t4 gnd.t133 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X15 gnd.t285 commonsourceibias.t52 CSoutput.t22 gnd.t181 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X16 CSoutput.t188 commonsourceibias.t53 gnd.t284 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 a_n8300_8799.t30 plus.t5 a_n2903_n3924.t29 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X18 gnd.t283 commonsourceibias.t54 CSoutput.t29 gnd.t192 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X19 vdd.t216 a_n8300_8799.t41 CSoutput.t177 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X20 CSoutput.t12 commonsourceibias.t55 gnd.t282 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X21 minus.t4 gnd.t129 gnd.t131 gnd.t130 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X22 CSoutput.t52 commonsourceibias.t56 gnd.t281 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 gnd.t128 gnd.t125 gnd.t127 gnd.t126 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X24 CSoutput.t23 commonsourceibias.t57 gnd.t280 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 a_n8300_8799.t1 a_n2318_13878.t54 a_n2318_8322.t14 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X26 vdd.t215 a_n8300_8799.t42 CSoutput.t176 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X27 vdd.t214 a_n8300_8799.t43 CSoutput.t175 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X28 CSoutput.t174 a_n8300_8799.t44 vdd.t213 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X29 vdd.t212 a_n8300_8799.t45 CSoutput.t173 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X30 a_n8300_8799.t2 a_n2318_13878.t55 a_n2318_8322.t13 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X31 CSoutput.t185 commonsourceibias.t58 gnd.t279 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 gnd.t278 commonsourceibias.t59 CSoutput.t16 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X33 gnd.t124 gnd.t122 gnd.t123 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X34 a_n8300_8799.t4 plus.t6 a_n2903_n3924.t28 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X35 CSoutput.t51 commonsourceibias.t60 gnd.t277 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 CSoutput.t193 a_n2318_8322.t24 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X37 vdd.t299 vdd.t297 vdd.t298 vdd.t225 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X38 CSoutput.t2 commonsourceibias.t61 gnd.t276 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X39 CSoutput.t172 a_n8300_8799.t46 vdd.t211 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X40 a_n2903_n3924.t41 diffpairibias.t16 gnd.t158 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X41 a_n2903_n3924.t34 minus.t5 a_n2318_13878.t11 gnd.t142 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X42 CSoutput.t171 a_n8300_8799.t47 vdd.t210 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X43 CSoutput.t170 a_n8300_8799.t48 vdd.t209 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X44 gnd.t275 commonsourceibias.t62 CSoutput.t14 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X45 gnd.t115 gnd.t112 gnd.t114 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X46 a_n2903_n3924.t27 plus.t7 a_n8300_8799.t35 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X47 vdd.t208 a_n8300_8799.t49 CSoutput.t169 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X48 CSoutput.t1 commonsourceibias.t63 gnd.t274 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X49 a_n2318_13878.t9 minus.t6 a_n2903_n3924.t32 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X50 gnd.t272 commonsourceibias.t24 commonsourceibias.t25 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 CSoutput.t19 commonsourceibias.t64 gnd.t273 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 a_n2903_n3924.t26 plus.t8 a_n8300_8799.t6 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X53 a_n2903_n3924.t0 minus.t7 a_n2318_13878.t0 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X54 CSoutput.t168 a_n8300_8799.t50 vdd.t207 vdd.t78 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X55 CSoutput.t48 commonsourceibias.t65 gnd.t271 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 a_n2140_13878.t14 a_n2318_13878.t36 a_n2318_13878.t37 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X57 a_n2318_13878.t19 a_n2318_13878.t18 a_n2140_13878.t13 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X58 outputibias.t7 outputibias.t6 gnd.t164 gnd.t163 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X59 gnd.t270 commonsourceibias.t66 CSoutput.t34 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X60 CSoutput.t167 a_n8300_8799.t51 vdd.t206 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 gnd.t269 commonsourceibias.t22 commonsourceibias.t23 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X62 a_n2903_n3924.t3 minus.t8 a_n2318_13878.t2 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X63 vdd.t296 vdd.t294 vdd.t295 vdd.t271 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X64 CSoutput.t20 commonsourceibias.t67 gnd.t268 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X65 vdd.t205 a_n8300_8799.t52 CSoutput.t166 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X66 gnd.t121 gnd.t119 gnd.t120 gnd.t31 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X67 gnd.t118 gnd.t116 gnd.t117 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X68 CSoutput.t35 commonsourceibias.t68 gnd.t267 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X69 diffpairibias.t15 diffpairibias.t14 gnd.t152 gnd.t151 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X70 CSoutput.t183 commonsourceibias.t69 gnd.t266 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X71 CSoutput.t3 commonsourceibias.t70 gnd.t265 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X72 gnd.t111 gnd.t109 gnd.t110 gnd.t42 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X73 gnd.t264 commonsourceibias.t71 CSoutput.t6 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 a_n8300_8799.t21 a_n2318_13878.t56 a_n2318_8322.t12 vdd.t48 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X75 CSoutput.t165 a_n8300_8799.t53 vdd.t204 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X76 gnd.t263 commonsourceibias.t72 CSoutput.t11 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X77 gnd.t108 gnd.t107 plus.t3 gnd.t42 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X78 vdd.t203 a_n8300_8799.t54 CSoutput.t164 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X79 vdd.t202 a_n8300_8799.t55 CSoutput.t163 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X80 minus.t3 gnd.t104 gnd.t106 gnd.t105 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X81 CSoutput.t8 commonsourceibias.t73 gnd.t262 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X82 diffpairibias.t13 diffpairibias.t12 gnd.t154 gnd.t153 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X83 CSoutput.t162 a_n8300_8799.t56 vdd.t201 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X84 gnd.t261 commonsourceibias.t26 commonsourceibias.t27 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 CSoutput.t26 commonsourceibias.t74 gnd.t260 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X86 gnd.t259 commonsourceibias.t75 CSoutput.t4 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 output.t18 CSoutput.t194 vdd.t53 gnd.t304 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X88 CSoutput.t25 commonsourceibias.t76 gnd.t258 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 vdd.t200 a_n8300_8799.t57 CSoutput.t161 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X90 CSoutput.t160 a_n8300_8799.t58 vdd.t199 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X91 gnd.t257 commonsourceibias.t77 CSoutput.t21 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X92 vdd.t293 vdd.t291 vdd.t292 vdd.t261 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X93 CSoutput.t159 a_n8300_8799.t59 vdd.t198 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X94 CSoutput.t158 a_n8300_8799.t60 vdd.t197 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X95 CSoutput.t157 a_n8300_8799.t61 vdd.t196 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 a_n8300_8799.t33 plus.t9 a_n2903_n3924.t25 gnd.t155 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X97 output.t17 CSoutput.t195 vdd.t60 gnd.t303 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X98 gnd.t256 commonsourceibias.t78 CSoutput.t0 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X99 a_n2903_n3924.t31 diffpairibias.t17 gnd.t140 gnd.t139 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X100 vdd.t190 a_n8300_8799.t62 CSoutput.t156 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X101 gnd.t103 gnd.t101 gnd.t102 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X102 a_n2903_n3924.t9 minus.t9 a_n2318_13878.t8 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X103 vdd.t195 a_n8300_8799.t63 CSoutput.t155 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X104 a_n2318_13878.t23 a_n2318_13878.t22 a_n2140_13878.t12 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X105 vdd.t194 a_n8300_8799.t64 CSoutput.t154 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X106 vdd.t191 a_n8300_8799.t65 CSoutput.t153 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X107 gnd.t255 commonsourceibias.t79 CSoutput.t17 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 a_n8300_8799.t22 a_n2318_13878.t57 a_n2318_8322.t11 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X109 vdd.t193 a_n8300_8799.t66 CSoutput.t152 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X110 a_n2318_13878.t41 a_n2318_13878.t40 a_n2140_13878.t11 vdd.t20 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X111 a_n2318_13878.t16 minus.t10 a_n2903_n3924.t43 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X112 gnd.t100 gnd.t98 gnd.t99 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X113 a_n2903_n3924.t24 plus.t10 a_n8300_8799.t34 gnd.t308 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X114 vdd.t192 a_n8300_8799.t67 CSoutput.t151 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X115 CSoutput.t150 a_n8300_8799.t68 vdd.t189 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X116 gnd.t254 commonsourceibias.t80 CSoutput.t24 gnd.t176 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 a_n2903_n3924.t2 minus.t11 a_n2318_13878.t1 gnd.t9 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X118 output.t16 CSoutput.t196 vdd.t61 gnd.t302 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X119 vdd.t290 vdd.t288 vdd.t289 vdd.t275 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X120 vdd.t287 vdd.t285 vdd.t286 vdd.t237 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X121 gnd.t253 commonsourceibias.t12 commonsourceibias.t13 gnd.t181 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X122 gnd.t252 commonsourceibias.t81 CSoutput.t18 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X123 CSoutput.t149 a_n8300_8799.t69 vdd.t188 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X124 vdd.t284 vdd.t281 vdd.t283 vdd.t282 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X125 output.t2 outputibias.t9 gnd.t168 gnd.t167 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X126 CSoutput.t197 a_n2318_8322.t25 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X127 CSoutput.t148 a_n8300_8799.t70 vdd.t187 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X128 gnd.t97 gnd.t94 gnd.t96 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X129 vdd.t186 a_n8300_8799.t71 CSoutput.t147 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X130 vdd.t16 a_n2318_13878.t58 a_n2318_8322.t23 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X131 a_n2318_13878.t21 a_n2318_13878.t20 a_n2140_13878.t10 vdd.t45 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X132 vdd.t280 vdd.t278 vdd.t279 vdd.t261 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X133 a_n2318_8322.t22 a_n2318_13878.t59 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X134 a_n2903_n3924.t30 diffpairibias.t18 gnd.t138 gnd.t137 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X135 CSoutput.t146 a_n8300_8799.t72 vdd.t185 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X136 CSoutput.t145 a_n8300_8799.t73 vdd.t183 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X137 outputibias.t5 outputibias.t4 gnd.t322 gnd.t321 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X138 vdd.t54 CSoutput.t198 output.t15 gnd.t301 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X139 a_n2318_13878.t15 minus.t12 a_n2903_n3924.t42 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X140 CSoutput.t46 commonsourceibias.t82 gnd.t251 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X141 CSoutput.t189 commonsourceibias.t83 gnd.t250 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X142 gnd.t93 gnd.t91 gnd.t92 gnd.t31 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X143 a_n2903_n3924.t23 plus.t11 a_n8300_8799.t14 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X144 vdd.t1 a_n2318_13878.t60 a_n2140_13878.t22 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X145 outputibias.t3 outputibias.t2 gnd.t162 gnd.t161 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X146 vdd.t277 vdd.t274 vdd.t276 vdd.t275 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X147 gnd.t90 gnd.t88 gnd.t89 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X148 vdd.t182 a_n8300_8799.t74 CSoutput.t144 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X149 vdd.t180 a_n8300_8799.t75 CSoutput.t143 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X150 vdd.t179 a_n8300_8799.t76 CSoutput.t142 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X151 a_n8300_8799.t15 plus.t12 a_n2903_n3924.t22 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X152 vdd.t273 vdd.t270 vdd.t272 vdd.t271 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X153 a_n2318_8322.t21 a_n2318_13878.t61 vdd.t3 vdd.t2 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X154 a_n2318_13878.t10 minus.t13 a_n2903_n3924.t33 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X155 a_n8300_8799.t28 a_n2318_13878.t62 a_n2318_8322.t10 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X156 CSoutput.t141 a_n8300_8799.t77 vdd.t177 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X157 diffpairibias.t11 diffpairibias.t10 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X158 vdd.t176 a_n8300_8799.t78 CSoutput.t140 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 a_n2318_13878.t33 a_n2318_13878.t32 a_n2140_13878.t9 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X160 vdd.t174 a_n8300_8799.t79 CSoutput.t139 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X161 CSoutput.t7 commonsourceibias.t84 gnd.t249 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X162 vdd.t55 CSoutput.t199 output.t14 gnd.t300 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X163 a_n8300_8799.t29 a_n2318_13878.t63 a_n2318_8322.t9 vdd.t59 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X164 CSoutput.t138 a_n8300_8799.t80 vdd.t173 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X165 commonsourceibias.t37 commonsourceibias.t36 gnd.t248 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X166 output.t13 CSoutput.t200 vdd.t56 gnd.t299 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X167 gnd.t247 commonsourceibias.t85 CSoutput.t53 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 a_n2140_13878.t8 a_n2318_13878.t46 a_n2318_13878.t47 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X169 vdd.t269 vdd.t267 vdd.t268 vdd.t237 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X170 plus.t2 gnd.t85 gnd.t87 gnd.t86 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X171 CSoutput.t201 a_n2318_8322.t27 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X172 gnd.t84 gnd.t82 minus.t2 gnd.t83 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X173 output.t12 CSoutput.t202 vdd.t40 gnd.t298 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X174 CSoutput.t137 a_n8300_8799.t81 vdd.t172 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X175 a_n2318_13878.t12 minus.t14 a_n2903_n3924.t36 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X176 CSoutput.t13 commonsourceibias.t86 gnd.t246 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X177 vdd.t34 a_n2318_13878.t64 a_n2318_8322.t20 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X178 a_n2140_13878.t7 a_n2318_13878.t48 a_n2318_13878.t49 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X179 CSoutput.t203 a_n2318_8322.t26 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X180 vdd.t171 a_n8300_8799.t82 CSoutput.t136 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X181 gnd.t245 commonsourceibias.t87 CSoutput.t187 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X182 gnd.t244 commonsourceibias.t88 CSoutput.t47 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 a_n2318_13878.t25 a_n2318_13878.t24 a_n2140_13878.t6 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X184 commonsourceibias.t35 commonsourceibias.t34 gnd.t243 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X185 gnd.t241 commonsourceibias.t89 CSoutput.t5 gnd.t192 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X186 outputibias.t1 outputibias.t0 gnd.t8 gnd.t7 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X187 vdd.t170 a_n8300_8799.t83 CSoutput.t135 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X188 CSoutput.t15 commonsourceibias.t90 gnd.t240 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 a_n2903_n3924.t1 diffpairibias.t19 gnd.t6 gnd.t5 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X190 gnd.t66 gnd.t63 gnd.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X191 a_n2903_n3924.t38 diffpairibias.t20 gnd.t150 gnd.t149 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X192 commonsourceibias.t33 commonsourceibias.t32 gnd.t239 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 output.t1 outputibias.t10 gnd.t312 gnd.t311 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X194 a_n2318_13878.t17 minus.t15 a_n2903_n3924.t44 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X195 vdd.t169 a_n8300_8799.t84 CSoutput.t134 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X196 vdd.t168 a_n8300_8799.t85 CSoutput.t133 vdd.t112 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X197 gnd.t81 gnd.t79 gnd.t80 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X198 gnd.t21 gnd.t19 minus.t1 gnd.t20 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X199 vdd.t4 CSoutput.t204 output.t11 gnd.t297 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X200 CSoutput.t184 commonsourceibias.t91 gnd.t237 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 CSoutput.t61 commonsourceibias.t92 gnd.t236 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X202 gnd.t78 gnd.t76 gnd.t77 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X203 gnd.t75 gnd.t73 gnd.t74 gnd.t23 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X204 CSoutput.t132 a_n8300_8799.t86 vdd.t167 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X205 CSoutput.t131 a_n8300_8799.t87 vdd.t166 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X206 commonsourceibias.t31 commonsourceibias.t30 gnd.t235 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 a_n2318_13878.t5 minus.t16 a_n2903_n3924.t6 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X208 CSoutput.t130 a_n8300_8799.t88 vdd.t164 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X209 diffpairibias.t9 diffpairibias.t8 gnd.t307 gnd.t306 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X210 a_n2140_13878.t21 a_n2318_13878.t65 vdd.t36 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X211 vdd.t223 a_n2318_13878.t66 a_n2140_13878.t20 vdd.t222 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X212 CSoutput.t62 commonsourceibias.t93 gnd.t234 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 CSoutput.t54 commonsourceibias.t94 gnd.t233 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X214 CSoutput.t129 a_n8300_8799.t89 vdd.t163 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X215 a_n2903_n3924.t21 plus.t13 a_n8300_8799.t31 gnd.t142 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X216 gnd.t232 commonsourceibias.t6 commonsourceibias.t7 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X217 vdd.t161 a_n8300_8799.t90 CSoutput.t128 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X218 vdd.t159 a_n8300_8799.t91 CSoutput.t127 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X219 commonsourceibias.t5 commonsourceibias.t4 gnd.t230 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 CSoutput.t126 a_n8300_8799.t92 vdd.t157 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X221 a_n2903_n3924.t5 minus.t17 a_n2318_13878.t4 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X222 a_n2140_13878.t5 a_n2318_13878.t26 a_n2318_13878.t27 vdd.t48 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X223 a_n2903_n3924.t20 plus.t14 a_n8300_8799.t8 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X224 gnd.t228 commonsourceibias.t95 CSoutput.t55 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X225 a_n2903_n3924.t45 minus.t18 a_n2318_13878.t50 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X226 commonsourceibias.t3 commonsourceibias.t2 gnd.t227 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X227 a_n8300_8799.t27 plus.t15 a_n2903_n3924.t19 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X228 vdd.t156 a_n8300_8799.t93 CSoutput.t125 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 gnd.t226 commonsourceibias.t0 commonsourceibias.t1 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X230 a_n2318_8322.t8 a_n2318_13878.t67 a_n8300_8799.t32 vdd.t51 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X231 CSoutput.t124 a_n8300_8799.t94 vdd.t155 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X232 gnd.t62 gnd.t59 gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X233 diffpairibias.t7 diffpairibias.t6 gnd.t316 gnd.t315 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X234 gnd.t72 gnd.t70 gnd.t71 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X235 vdd.t154 a_n8300_8799.t95 CSoutput.t123 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X236 commonsourceibias.t21 commonsourceibias.t20 gnd.t225 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X237 vdd.t266 vdd.t264 vdd.t265 vdd.t247 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X238 vdd.t11 a_n2318_13878.t68 a_n2318_8322.t19 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X239 output.t10 CSoutput.t205 vdd.t5 gnd.t296 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X240 vdd.t152 a_n8300_8799.t96 CSoutput.t122 vdd.t112 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X241 vdd.t151 a_n8300_8799.t97 CSoutput.t121 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X242 gnd.t224 commonsourceibias.t96 CSoutput.t36 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 output.t0 outputibias.t11 gnd.t166 gnd.t165 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X244 CSoutput.t120 a_n8300_8799.t98 vdd.t149 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X245 gnd.t223 commonsourceibias.t18 commonsourceibias.t19 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 a_n2140_13878.t19 a_n2318_13878.t69 vdd.t13 vdd.t12 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X247 vdd.t263 vdd.t260 vdd.t262 vdd.t261 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X248 vdd.t259 vdd.t257 vdd.t258 vdd.t247 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X249 plus.t1 gnd.t67 gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X250 output.t9 CSoutput.t206 vdd.t6 gnd.t295 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X251 vdd.t148 a_n8300_8799.t99 CSoutput.t119 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X252 CSoutput.t118 a_n8300_8799.t100 vdd.t147 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X253 CSoutput.t117 a_n8300_8799.t101 vdd.t146 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X254 CSoutput.t116 a_n8300_8799.t102 vdd.t145 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X255 gnd.t58 gnd.t56 minus.t0 gnd.t57 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X256 gnd.t55 gnd.t52 gnd.t54 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X257 vdd.t144 a_n8300_8799.t103 CSoutput.t115 vdd.t72 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X258 a_n2903_n3924.t47 diffpairibias.t21 gnd.t314 gnd.t313 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X259 vdd.t42 a_n2318_13878.t70 a_n2318_8322.t18 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X260 a_n2318_8322.t7 a_n2318_13878.t71 a_n8300_8799.t17 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X261 CSoutput.t114 a_n8300_8799.t104 vdd.t143 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X262 gnd.t221 commonsourceibias.t16 commonsourceibias.t17 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X263 vdd.t141 a_n8300_8799.t105 CSoutput.t113 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X264 CSoutput.t112 a_n8300_8799.t106 vdd.t140 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X265 CSoutput.t207 a_n2318_8322.t25 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X266 vdd.t139 a_n8300_8799.t107 CSoutput.t111 vdd.t74 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X267 vdd.t138 a_n8300_8799.t108 CSoutput.t110 vdd.t83 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X268 vdd.t256 vdd.t254 vdd.t255 vdd.t233 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X269 gnd.t220 commonsourceibias.t14 commonsourceibias.t15 gnd.t176 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X270 a_n2903_n3924.t18 plus.t16 a_n8300_8799.t26 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X271 vdd.t253 vdd.t250 vdd.t252 vdd.t251 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X272 vdd.t57 CSoutput.t208 output.t8 gnd.t294 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X273 vdd.t137 a_n8300_8799.t109 CSoutput.t109 vdd.t80 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X274 vdd.t58 CSoutput.t209 output.t7 gnd.t293 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X275 a_n8300_8799.t9 plus.t17 a_n2903_n3924.t17 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X276 CSoutput.t108 a_n8300_8799.t110 vdd.t136 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X277 CSoutput.t37 commonsourceibias.t97 gnd.t219 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 a_n2903_n3924.t46 minus.t19 a_n2318_13878.t51 gnd.t308 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X279 a_n2140_13878.t4 a_n2318_13878.t44 a_n2318_13878.t45 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X280 CSoutput.t107 a_n8300_8799.t111 vdd.t134 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X281 a_n2318_8322.t6 a_n2318_13878.t72 a_n8300_8799.t7 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X282 vdd.t249 vdd.t246 vdd.t248 vdd.t247 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X283 diffpairibias.t5 diffpairibias.t4 gnd.t310 gnd.t309 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X284 a_n2903_n3924.t8 minus.t20 a_n2318_13878.t7 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X285 a_n8300_8799.t5 plus.t18 a_n2903_n3924.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X286 gnd.t51 gnd.t48 gnd.t50 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X287 CSoutput.t106 a_n8300_8799.t112 vdd.t133 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 CSoutput.t105 a_n8300_8799.t113 vdd.t131 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X289 CSoutput.t104 a_n8300_8799.t114 vdd.t129 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X290 vdd.t128 a_n8300_8799.t115 CSoutput.t103 vdd.t74 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X291 CSoutput.t38 commonsourceibias.t98 gnd.t217 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X292 vdd.t127 a_n8300_8799.t116 CSoutput.t102 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 a_n2318_8322.t17 a_n2318_13878.t73 vdd.t24 vdd.t23 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X294 CSoutput.t101 a_n8300_8799.t117 vdd.t125 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X295 CSoutput.t100 a_n8300_8799.t118 vdd.t123 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X296 a_n2903_n3924.t15 plus.t19 a_n8300_8799.t24 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X297 vdd.t121 a_n8300_8799.t119 CSoutput.t99 vdd.t72 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X298 vdd.t245 vdd.t243 vdd.t244 vdd.t229 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X299 gnd.t47 gnd.t45 gnd.t46 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X300 gnd.t215 commonsourceibias.t99 CSoutput.t39 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 CSoutput.t98 a_n8300_8799.t120 vdd.t120 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X302 vdd.t31 a_n2318_13878.t74 a_n2140_13878.t18 vdd.t30 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X303 vdd.t73 a_n8300_8799.t121 CSoutput.t97 vdd.t72 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X304 CSoutput.t96 a_n8300_8799.t122 vdd.t119 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X305 CSoutput.t95 a_n8300_8799.t123 vdd.t117 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X306 gnd.t44 gnd.t41 gnd.t43 gnd.t42 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X307 vdd.t75 a_n8300_8799.t124 CSoutput.t94 vdd.t74 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 vdd.t116 a_n8300_8799.t125 CSoutput.t93 vdd.t83 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X309 gnd.t214 commonsourceibias.t100 CSoutput.t40 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X310 a_n2903_n3924.t4 minus.t21 a_n2318_13878.t3 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X311 gnd.t213 commonsourceibias.t101 CSoutput.t41 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X312 vdd.t242 vdd.t240 vdd.t241 vdd.t233 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X313 output.t6 CSoutput.t210 vdd.t37 gnd.t292 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X314 gnd.t40 gnd.t38 gnd.t39 gnd.t31 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X315 a_n2318_8322.t5 a_n2318_13878.t75 a_n8300_8799.t13 vdd.t32 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X316 commonsourceibias.t29 commonsourceibias.t28 gnd.t212 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X317 vdd.t38 CSoutput.t211 output.t5 gnd.t291 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X318 CSoutput.t92 a_n8300_8799.t126 vdd.t115 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X319 a_n8300_8799.t20 a_n2318_13878.t76 a_n2318_8322.t4 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X320 vdd.t113 a_n8300_8799.t127 CSoutput.t91 vdd.t112 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X321 a_n2140_13878.t17 a_n2318_13878.t77 vdd.t47 vdd.t46 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X322 gnd.t210 commonsourceibias.t102 CSoutput.t42 gnd.t176 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X323 vdd.t111 a_n8300_8799.t128 CSoutput.t90 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X324 CSoutput.t89 a_n8300_8799.t129 vdd.t110 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 a_n8300_8799.t16 plus.t20 a_n2903_n3924.t14 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X326 gnd.t209 commonsourceibias.t103 CSoutput.t43 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X327 commonsourceibias.t39 commonsourceibias.t38 gnd.t198 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X328 a_n2318_8322.t3 a_n2318_13878.t78 a_n8300_8799.t18 vdd.t45 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X329 gnd.t208 commonsourceibias.t104 CSoutput.t44 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 a_n2318_13878.t13 minus.t22 a_n2903_n3924.t39 gnd.t155 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X331 vdd.t108 a_n8300_8799.t130 CSoutput.t88 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X332 gnd.t206 commonsourceibias.t44 commonsourceibias.t45 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X333 CSoutput.t87 a_n8300_8799.t131 vdd.t106 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X334 CSoutput.t86 a_n8300_8799.t132 vdd.t104 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X335 CSoutput.t85 a_n8300_8799.t133 vdd.t103 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X336 a_n2140_13878.t3 a_n2318_13878.t38 a_n2318_13878.t39 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X337 vdd.t102 a_n8300_8799.t134 CSoutput.t84 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X338 gnd.t202 commonsourceibias.t40 commonsourceibias.t41 gnd.t192 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X339 vdd.t239 vdd.t236 vdd.t238 vdd.t237 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X340 vdd.t235 vdd.t232 vdd.t234 vdd.t233 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X341 commonsourceibias.t43 commonsourceibias.t42 gnd.t204 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X342 a_n8300_8799.t10 plus.t21 a_n2903_n3924.t13 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X343 gnd.t201 commonsourceibias.t105 CSoutput.t45 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X344 a_n2903_n3924.t35 diffpairibias.t22 gnd.t146 gnd.t145 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X345 CSoutput.t9 commonsourceibias.t106 gnd.t199 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X346 vdd.t101 a_n8300_8799.t135 CSoutput.t83 vdd.t80 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X347 vdd.t100 a_n8300_8799.t136 CSoutput.t82 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X348 gnd.t196 commonsourceibias.t107 CSoutput.t10 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 CSoutput.t81 a_n8300_8799.t137 vdd.t99 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X350 a_n2318_13878.t43 a_n2318_13878.t42 a_n2140_13878.t2 vdd.t32 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X351 gnd.t37 gnd.t34 gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X352 a_n8300_8799.t19 a_n2318_13878.t79 a_n2318_8322.t2 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X353 vdd.t39 CSoutput.t212 output.t4 gnd.t290 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X354 gnd.t33 gnd.t30 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X355 vdd.t65 a_n8300_8799.t138 CSoutput.t80 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X356 CSoutput.t79 a_n8300_8799.t139 vdd.t98 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X357 a_n2903_n3924.t12 plus.t22 a_n8300_8799.t25 gnd.t9 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X358 vdd.t96 a_n8300_8799.t140 CSoutput.t78 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X359 CSoutput.t49 commonsourceibias.t108 gnd.t194 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X360 gnd.t193 commonsourceibias.t109 CSoutput.t50 gnd.t192 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X361 commonsourceibias.t11 commonsourceibias.t10 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 diffpairibias.t3 diffpairibias.t2 gnd.t160 gnd.t159 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X363 gnd.t29 gnd.t26 gnd.t28 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X364 vdd.t95 a_n8300_8799.t141 CSoutput.t77 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X365 CSoutput.t76 a_n8300_8799.t142 vdd.t93 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X366 CSoutput.t75 a_n8300_8799.t143 vdd.t92 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X367 a_n2318_8322.t1 a_n2318_13878.t80 a_n8300_8799.t12 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X368 gnd.t189 commonsourceibias.t110 CSoutput.t56 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X369 vdd.t90 a_n8300_8799.t144 CSoutput.t74 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X370 CSoutput.t213 a_n2318_8322.t24 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X371 CSoutput.t73 a_n8300_8799.t145 vdd.t88 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X372 diffpairibias.t1 diffpairibias.t0 gnd.t318 gnd.t317 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X373 a_n8300_8799.t0 plus.t23 a_n2903_n3924.t11 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X374 commonsourceibias.t9 commonsourceibias.t8 gnd.t188 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X375 gnd.t187 commonsourceibias.t111 CSoutput.t57 gnd.t181 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X376 CSoutput.t30 commonsourceibias.t112 gnd.t186 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X377 gnd.t25 gnd.t22 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X378 vdd.t231 vdd.t228 vdd.t230 vdd.t229 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X379 vdd.t29 a_n2318_13878.t81 a_n2140_13878.t16 vdd.t28 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X380 CSoutput.t72 a_n8300_8799.t146 vdd.t86 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X381 vdd.t227 vdd.t224 vdd.t226 vdd.t225 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X382 vdd.t84 a_n8300_8799.t147 CSoutput.t71 vdd.t83 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X383 vdd.t82 a_n8300_8799.t148 CSoutput.t70 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X384 gnd.t184 commonsourceibias.t46 commonsourceibias.t47 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X385 CSoutput.t69 a_n8300_8799.t149 vdd.t79 vdd.t78 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X386 a_n2318_13878.t6 minus.t23 a_n2903_n3924.t7 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X387 gnd.t182 commonsourceibias.t113 CSoutput.t31 gnd.t181 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X388 gnd.t180 commonsourceibias.t114 CSoutput.t58 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X389 a_n2318_8322.t0 a_n2318_13878.t82 a_n8300_8799.t11 vdd.t20 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X390 vdd.t81 a_n8300_8799.t150 CSoutput.t68 vdd.t80 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X391 vdd.t77 a_n8300_8799.t151 CSoutput.t67 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X392 vdd.t71 a_n8300_8799.t152 CSoutput.t66 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X393 CSoutput.t65 a_n8300_8799.t153 vdd.t69 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X394 gnd.t178 commonsourceibias.t115 CSoutput.t59 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X395 gnd.t18 gnd.t16 plus.t0 gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X396 a_n2903_n3924.t10 plus.t24 a_n8300_8799.t3 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X397 a_n2318_8322.t16 a_n2318_13878.t83 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X398 a_n2318_13878.t14 minus.t24 a_n2903_n3924.t40 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X399 gnd.t177 commonsourceibias.t116 CSoutput.t27 gnd.t176 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X400 a_n2140_13878.t1 a_n2318_13878.t28 a_n2318_13878.t29 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X401 gnd.t175 commonsourceibias.t117 CSoutput.t28 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X402 CSoutput.t190 commonsourceibias.t118 gnd.t173 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X403 vdd.t67 a_n8300_8799.t154 CSoutput.t64 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X404 CSoutput.t191 commonsourceibias.t119 gnd.t171 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X405 a_n2903_n3924.t37 diffpairibias.t23 gnd.t148 gnd.t147 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X406 CSoutput.t63 a_n8300_8799.t155 vdd.t63 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X407 a_n2318_13878.t31 a_n2318_13878.t30 a_n2140_13878.t0 vdd.t51 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 a_n8300_8799.n228 a_n8300_8799.t145 485.149
R1 a_n8300_8799.n247 a_n8300_8799.t38 485.149
R2 a_n8300_8799.n267 a_n8300_8799.t120 485.149
R3 a_n8300_8799.n167 a_n8300_8799.t103 485.149
R4 a_n8300_8799.n186 a_n8300_8799.t119 485.149
R5 a_n8300_8799.n206 a_n8300_8799.t121 485.149
R6 a_n8300_8799.n55 a_n8300_8799.t85 485.135
R7 a_n8300_8799.n240 a_n8300_8799.t61 464.166
R8 a_n8300_8799.n222 a_n8300_8799.t140 464.166
R9 a_n8300_8799.n239 a_n8300_8799.t102 464.166
R10 a_n8300_8799.n238 a_n8300_8799.t99 464.166
R11 a_n8300_8799.n223 a_n8300_8799.t39 464.166
R12 a_n8300_8799.n237 a_n8300_8799.t107 464.166
R13 a_n8300_8799.n236 a_n8300_8799.t106 464.166
R14 a_n8300_8799.n224 a_n8300_8799.t41 464.166
R15 a_n8300_8799.n235 a_n8300_8799.t40 464.166
R16 a_n8300_8799.n234 a_n8300_8799.t128 464.166
R17 a_n8300_8799.n225 a_n8300_8799.t56 464.166
R18 a_n8300_8799.n233 a_n8300_8799.t45 464.166
R19 a_n8300_8799.n232 a_n8300_8799.t132 464.166
R20 a_n8300_8799.n226 a_n8300_8799.t84 464.166
R21 a_n8300_8799.n231 a_n8300_8799.t60 464.166
R22 a_n8300_8799.n230 a_n8300_8799.t152 464.166
R23 a_n8300_8799.n227 a_n8300_8799.t101 464.166
R24 a_n8300_8799.n229 a_n8300_8799.t63 464.166
R25 a_n8300_8799.n70 a_n8300_8799.t96 485.135
R26 a_n8300_8799.n259 a_n8300_8799.t72 464.166
R27 a_n8300_8799.n241 a_n8300_8799.t154 464.166
R28 a_n8300_8799.n258 a_n8300_8799.t117 464.166
R29 a_n8300_8799.n257 a_n8300_8799.t116 464.166
R30 a_n8300_8799.n242 a_n8300_8799.t50 464.166
R31 a_n8300_8799.n256 a_n8300_8799.t124 464.166
R32 a_n8300_8799.n255 a_n8300_8799.t123 464.166
R33 a_n8300_8799.n243 a_n8300_8799.t52 464.166
R34 a_n8300_8799.n254 a_n8300_8799.t51 464.166
R35 a_n8300_8799.n253 a_n8300_8799.t144 464.166
R36 a_n8300_8799.n244 a_n8300_8799.t69 464.166
R37 a_n8300_8799.n252 a_n8300_8799.t55 464.166
R38 a_n8300_8799.n251 a_n8300_8799.t146 464.166
R39 a_n8300_8799.n245 a_n8300_8799.t97 464.166
R40 a_n8300_8799.n250 a_n8300_8799.t73 464.166
R41 a_n8300_8799.n249 a_n8300_8799.t43 464.166
R42 a_n8300_8799.n246 a_n8300_8799.t118 464.166
R43 a_n8300_8799.n248 a_n8300_8799.t74 464.166
R44 a_n8300_8799.n85 a_n8300_8799.t127 485.135
R45 a_n8300_8799.n279 a_n8300_8799.t58 464.166
R46 a_n8300_8799.n261 a_n8300_8799.t105 464.166
R47 a_n8300_8799.n278 a_n8300_8799.t44 464.166
R48 a_n8300_8799.n277 a_n8300_8799.t64 464.166
R49 a_n8300_8799.n262 a_n8300_8799.t149 464.166
R50 a_n8300_8799.n276 a_n8300_8799.t115 464.166
R51 a_n8300_8799.n275 a_n8300_8799.t143 464.166
R52 a_n8300_8799.n263 a_n8300_8799.t95 464.166
R53 a_n8300_8799.n274 a_n8300_8799.t122 464.166
R54 a_n8300_8799.n273 a_n8300_8799.t54 464.166
R55 a_n8300_8799.n264 a_n8300_8799.t139 464.166
R56 a_n8300_8799.n272 a_n8300_8799.t78 464.166
R57 a_n8300_8799.n271 a_n8300_8799.t133 464.166
R58 a_n8300_8799.n265 a_n8300_8799.t62 464.166
R59 a_n8300_8799.n270 a_n8300_8799.t110 464.166
R60 a_n8300_8799.n269 a_n8300_8799.t49 464.166
R61 a_n8300_8799.n266 a_n8300_8799.t92 464.166
R62 a_n8300_8799.n268 a_n8300_8799.t71 464.166
R63 a_n8300_8799.n168 a_n8300_8799.t142 464.166
R64 a_n8300_8799.n169 a_n8300_8799.t65 464.166
R65 a_n8300_8799.n170 a_n8300_8799.t98 464.166
R66 a_n8300_8799.n171 a_n8300_8799.t135 464.166
R67 a_n8300_8799.n166 a_n8300_8799.t137 464.166
R68 a_n8300_8799.n172 a_n8300_8799.t83 464.166
R69 a_n8300_8799.n173 a_n8300_8799.t114 464.166
R70 a_n8300_8799.n174 a_n8300_8799.t134 464.166
R71 a_n8300_8799.n175 a_n8300_8799.t81 464.166
R72 a_n8300_8799.n165 a_n8300_8799.t82 464.166
R73 a_n8300_8799.n176 a_n8300_8799.t111 464.166
R74 a_n8300_8799.n164 a_n8300_8799.t67 464.166
R75 a_n8300_8799.n177 a_n8300_8799.t68 464.166
R76 a_n8300_8799.n178 a_n8300_8799.t108 464.166
R77 a_n8300_8799.n179 a_n8300_8799.t36 464.166
R78 a_n8300_8799.n180 a_n8300_8799.t66 464.166
R79 a_n8300_8799.n163 a_n8300_8799.t88 464.166
R80 a_n8300_8799.n181 a_n8300_8799.t136 464.166
R81 a_n8300_8799.n187 a_n8300_8799.t155 464.166
R82 a_n8300_8799.n188 a_n8300_8799.t75 464.166
R83 a_n8300_8799.n189 a_n8300_8799.t112 464.166
R84 a_n8300_8799.n190 a_n8300_8799.t150 464.166
R85 a_n8300_8799.n185 a_n8300_8799.t153 464.166
R86 a_n8300_8799.n191 a_n8300_8799.t93 464.166
R87 a_n8300_8799.n192 a_n8300_8799.t131 464.166
R88 a_n8300_8799.n193 a_n8300_8799.t148 464.166
R89 a_n8300_8799.n194 a_n8300_8799.t89 464.166
R90 a_n8300_8799.n184 a_n8300_8799.t90 464.166
R91 a_n8300_8799.n195 a_n8300_8799.t129 464.166
R92 a_n8300_8799.n183 a_n8300_8799.t79 464.166
R93 a_n8300_8799.n196 a_n8300_8799.t80 464.166
R94 a_n8300_8799.n197 a_n8300_8799.t125 464.166
R95 a_n8300_8799.n198 a_n8300_8799.t46 464.166
R96 a_n8300_8799.n199 a_n8300_8799.t76 464.166
R97 a_n8300_8799.n182 a_n8300_8799.t100 464.166
R98 a_n8300_8799.n200 a_n8300_8799.t151 464.166
R99 a_n8300_8799.n207 a_n8300_8799.t70 464.166
R100 a_n8300_8799.n208 a_n8300_8799.t91 464.166
R101 a_n8300_8799.n209 a_n8300_8799.t48 464.166
R102 a_n8300_8799.n210 a_n8300_8799.t109 464.166
R103 a_n8300_8799.n205 a_n8300_8799.t86 464.166
R104 a_n8300_8799.n211 a_n8300_8799.t130 464.166
R105 a_n8300_8799.n212 a_n8300_8799.t77 464.166
R106 a_n8300_8799.n213 a_n8300_8799.t138 464.166
R107 a_n8300_8799.n214 a_n8300_8799.t53 464.166
R108 a_n8300_8799.n204 a_n8300_8799.t37 464.166
R109 a_n8300_8799.n215 a_n8300_8799.t94 464.166
R110 a_n8300_8799.n203 a_n8300_8799.t141 464.166
R111 a_n8300_8799.n216 a_n8300_8799.t113 464.166
R112 a_n8300_8799.n217 a_n8300_8799.t147 464.166
R113 a_n8300_8799.n218 a_n8300_8799.t87 464.166
R114 a_n8300_8799.n219 a_n8300_8799.t42 464.166
R115 a_n8300_8799.n202 a_n8300_8799.t104 464.166
R116 a_n8300_8799.n220 a_n8300_8799.t57 464.166
R117 a_n8300_8799.n41 a_n8300_8799.n69 71.7212
R118 a_n8300_8799.n69 a_n8300_8799.n227 17.8606
R119 a_n8300_8799.n68 a_n8300_8799.n41 76.9909
R120 a_n8300_8799.n230 a_n8300_8799.n68 7.32118
R121 a_n8300_8799.n67 a_n8300_8799.n40 78.3454
R122 a_n8300_8799.n40 a_n8300_8799.n66 72.8951
R123 a_n8300_8799.n65 a_n8300_8799.n42 70.1674
R124 a_n8300_8799.n233 a_n8300_8799.n65 20.9683
R125 a_n8300_8799.n42 a_n8300_8799.n64 72.3034
R126 a_n8300_8799.n64 a_n8300_8799.n225 16.6962
R127 a_n8300_8799.n63 a_n8300_8799.n43 77.6622
R128 a_n8300_8799.n234 a_n8300_8799.n63 5.97853
R129 a_n8300_8799.n62 a_n8300_8799.n43 77.6622
R130 a_n8300_8799.n44 a_n8300_8799.n61 72.3034
R131 a_n8300_8799.n60 a_n8300_8799.n44 70.1674
R132 a_n8300_8799.n237 a_n8300_8799.n60 20.9683
R133 a_n8300_8799.n46 a_n8300_8799.n59 72.8951
R134 a_n8300_8799.n59 a_n8300_8799.n223 15.5127
R135 a_n8300_8799.n58 a_n8300_8799.n46 78.3454
R136 a_n8300_8799.n238 a_n8300_8799.n58 4.61226
R137 a_n8300_8799.n57 a_n8300_8799.n45 76.9909
R138 a_n8300_8799.n45 a_n8300_8799.n56 71.7212
R139 a_n8300_8799.n240 a_n8300_8799.n55 20.9683
R140 a_n8300_8799.n47 a_n8300_8799.n55 70.1674
R141 a_n8300_8799.n33 a_n8300_8799.n84 71.7212
R142 a_n8300_8799.n84 a_n8300_8799.n246 17.8606
R143 a_n8300_8799.n83 a_n8300_8799.n33 76.9909
R144 a_n8300_8799.n249 a_n8300_8799.n83 7.32118
R145 a_n8300_8799.n82 a_n8300_8799.n32 78.3454
R146 a_n8300_8799.n32 a_n8300_8799.n81 72.8951
R147 a_n8300_8799.n80 a_n8300_8799.n34 70.1674
R148 a_n8300_8799.n252 a_n8300_8799.n80 20.9683
R149 a_n8300_8799.n34 a_n8300_8799.n79 72.3034
R150 a_n8300_8799.n79 a_n8300_8799.n244 16.6962
R151 a_n8300_8799.n78 a_n8300_8799.n35 77.6622
R152 a_n8300_8799.n253 a_n8300_8799.n78 5.97853
R153 a_n8300_8799.n77 a_n8300_8799.n35 77.6622
R154 a_n8300_8799.n36 a_n8300_8799.n76 72.3034
R155 a_n8300_8799.n75 a_n8300_8799.n36 70.1674
R156 a_n8300_8799.n256 a_n8300_8799.n75 20.9683
R157 a_n8300_8799.n38 a_n8300_8799.n74 72.8951
R158 a_n8300_8799.n74 a_n8300_8799.n242 15.5127
R159 a_n8300_8799.n73 a_n8300_8799.n38 78.3454
R160 a_n8300_8799.n257 a_n8300_8799.n73 4.61226
R161 a_n8300_8799.n72 a_n8300_8799.n37 76.9909
R162 a_n8300_8799.n37 a_n8300_8799.n71 71.7212
R163 a_n8300_8799.n259 a_n8300_8799.n70 20.9683
R164 a_n8300_8799.n39 a_n8300_8799.n70 70.1674
R165 a_n8300_8799.n25 a_n8300_8799.n99 71.7212
R166 a_n8300_8799.n99 a_n8300_8799.n266 17.8606
R167 a_n8300_8799.n98 a_n8300_8799.n25 76.9909
R168 a_n8300_8799.n269 a_n8300_8799.n98 7.32118
R169 a_n8300_8799.n97 a_n8300_8799.n24 78.3454
R170 a_n8300_8799.n24 a_n8300_8799.n96 72.8951
R171 a_n8300_8799.n95 a_n8300_8799.n26 70.1674
R172 a_n8300_8799.n272 a_n8300_8799.n95 20.9683
R173 a_n8300_8799.n26 a_n8300_8799.n94 72.3034
R174 a_n8300_8799.n94 a_n8300_8799.n264 16.6962
R175 a_n8300_8799.n93 a_n8300_8799.n27 77.6622
R176 a_n8300_8799.n273 a_n8300_8799.n93 5.97853
R177 a_n8300_8799.n92 a_n8300_8799.n27 77.6622
R178 a_n8300_8799.n28 a_n8300_8799.n91 72.3034
R179 a_n8300_8799.n90 a_n8300_8799.n28 70.1674
R180 a_n8300_8799.n276 a_n8300_8799.n90 20.9683
R181 a_n8300_8799.n30 a_n8300_8799.n89 72.8951
R182 a_n8300_8799.n89 a_n8300_8799.n262 15.5127
R183 a_n8300_8799.n88 a_n8300_8799.n30 78.3454
R184 a_n8300_8799.n277 a_n8300_8799.n88 4.61226
R185 a_n8300_8799.n87 a_n8300_8799.n29 76.9909
R186 a_n8300_8799.n29 a_n8300_8799.n86 71.7212
R187 a_n8300_8799.n279 a_n8300_8799.n85 20.9683
R188 a_n8300_8799.n31 a_n8300_8799.n85 70.1674
R189 a_n8300_8799.n17 a_n8300_8799.n114 70.1674
R190 a_n8300_8799.n181 a_n8300_8799.n114 20.9683
R191 a_n8300_8799.n113 a_n8300_8799.n17 71.7212
R192 a_n8300_8799.n113 a_n8300_8799.n163 17.8606
R193 a_n8300_8799.n16 a_n8300_8799.n112 76.9909
R194 a_n8300_8799.n180 a_n8300_8799.n112 7.32118
R195 a_n8300_8799.n111 a_n8300_8799.n16 78.3454
R196 a_n8300_8799.n18 a_n8300_8799.n110 72.8951
R197 a_n8300_8799.n109 a_n8300_8799.n18 70.1674
R198 a_n8300_8799.n109 a_n8300_8799.n164 20.9683
R199 a_n8300_8799.n19 a_n8300_8799.n108 72.3034
R200 a_n8300_8799.n176 a_n8300_8799.n108 16.6962
R201 a_n8300_8799.n107 a_n8300_8799.n19 77.6622
R202 a_n8300_8799.n107 a_n8300_8799.n165 5.97853
R203 a_n8300_8799.n20 a_n8300_8799.n106 77.6622
R204 a_n8300_8799.n105 a_n8300_8799.n20 72.3034
R205 a_n8300_8799.n21 a_n8300_8799.n104 70.1674
R206 a_n8300_8799.n172 a_n8300_8799.n104 20.9683
R207 a_n8300_8799.n103 a_n8300_8799.n21 72.8951
R208 a_n8300_8799.n103 a_n8300_8799.n166 15.5127
R209 a_n8300_8799.n22 a_n8300_8799.n102 78.3454
R210 a_n8300_8799.n171 a_n8300_8799.n102 4.61226
R211 a_n8300_8799.n101 a_n8300_8799.n22 76.9909
R212 a_n8300_8799.n100 a_n8300_8799.n169 17.8606
R213 a_n8300_8799.n100 a_n8300_8799.n23 71.7212
R214 a_n8300_8799.n9 a_n8300_8799.n129 70.1674
R215 a_n8300_8799.n200 a_n8300_8799.n129 20.9683
R216 a_n8300_8799.n128 a_n8300_8799.n9 71.7212
R217 a_n8300_8799.n128 a_n8300_8799.n182 17.8606
R218 a_n8300_8799.n8 a_n8300_8799.n127 76.9909
R219 a_n8300_8799.n199 a_n8300_8799.n127 7.32118
R220 a_n8300_8799.n126 a_n8300_8799.n8 78.3454
R221 a_n8300_8799.n10 a_n8300_8799.n125 72.8951
R222 a_n8300_8799.n124 a_n8300_8799.n10 70.1674
R223 a_n8300_8799.n124 a_n8300_8799.n183 20.9683
R224 a_n8300_8799.n11 a_n8300_8799.n123 72.3034
R225 a_n8300_8799.n195 a_n8300_8799.n123 16.6962
R226 a_n8300_8799.n122 a_n8300_8799.n11 77.6622
R227 a_n8300_8799.n122 a_n8300_8799.n184 5.97853
R228 a_n8300_8799.n12 a_n8300_8799.n121 77.6622
R229 a_n8300_8799.n120 a_n8300_8799.n12 72.3034
R230 a_n8300_8799.n13 a_n8300_8799.n119 70.1674
R231 a_n8300_8799.n191 a_n8300_8799.n119 20.9683
R232 a_n8300_8799.n118 a_n8300_8799.n13 72.8951
R233 a_n8300_8799.n118 a_n8300_8799.n185 15.5127
R234 a_n8300_8799.n14 a_n8300_8799.n117 78.3454
R235 a_n8300_8799.n190 a_n8300_8799.n117 4.61226
R236 a_n8300_8799.n116 a_n8300_8799.n14 76.9909
R237 a_n8300_8799.n115 a_n8300_8799.n188 17.8606
R238 a_n8300_8799.n115 a_n8300_8799.n15 71.7212
R239 a_n8300_8799.n1 a_n8300_8799.n144 70.1674
R240 a_n8300_8799.n220 a_n8300_8799.n144 20.9683
R241 a_n8300_8799.n143 a_n8300_8799.n1 71.7212
R242 a_n8300_8799.n143 a_n8300_8799.n202 17.8606
R243 a_n8300_8799.n0 a_n8300_8799.n142 76.9909
R244 a_n8300_8799.n219 a_n8300_8799.n142 7.32118
R245 a_n8300_8799.n141 a_n8300_8799.n0 78.3454
R246 a_n8300_8799.n2 a_n8300_8799.n140 72.8951
R247 a_n8300_8799.n139 a_n8300_8799.n2 70.1674
R248 a_n8300_8799.n139 a_n8300_8799.n203 20.9683
R249 a_n8300_8799.n3 a_n8300_8799.n138 72.3034
R250 a_n8300_8799.n215 a_n8300_8799.n138 16.6962
R251 a_n8300_8799.n137 a_n8300_8799.n3 77.6622
R252 a_n8300_8799.n137 a_n8300_8799.n204 5.97853
R253 a_n8300_8799.n4 a_n8300_8799.n136 77.6622
R254 a_n8300_8799.n135 a_n8300_8799.n4 72.3034
R255 a_n8300_8799.n5 a_n8300_8799.n134 70.1674
R256 a_n8300_8799.n211 a_n8300_8799.n134 20.9683
R257 a_n8300_8799.n133 a_n8300_8799.n5 72.8951
R258 a_n8300_8799.n133 a_n8300_8799.n205 15.5127
R259 a_n8300_8799.n6 a_n8300_8799.n132 78.3454
R260 a_n8300_8799.n210 a_n8300_8799.n132 4.61226
R261 a_n8300_8799.n131 a_n8300_8799.n6 76.9909
R262 a_n8300_8799.n130 a_n8300_8799.n208 17.8606
R263 a_n8300_8799.n130 a_n8300_8799.n7 71.7212
R264 a_n8300_8799.n53 a_n8300_8799.n145 98.9633
R265 a_n8300_8799.n52 a_n8300_8799.n148 98.9631
R266 a_n8300_8799.n54 a_n8300_8799.n147 98.6055
R267 a_n8300_8799.n53 a_n8300_8799.n146 98.6055
R268 a_n8300_8799.n52 a_n8300_8799.n149 98.6055
R269 a_n8300_8799.n52 a_n8300_8799.n150 98.6055
R270 a_n8300_8799.n152 a_n8300_8799.n151 98.6055
R271 a_n8300_8799.n284 a_n8300_8799.n54 98.6054
R272 a_n8300_8799.n51 a_n8300_8799.n153 81.2902
R273 a_n8300_8799.n49 a_n8300_8799.n159 81.2902
R274 a_n8300_8799.n48 a_n8300_8799.n156 81.2902
R275 a_n8300_8799.n50 a_n8300_8799.n161 80.9324
R276 a_n8300_8799.n50 a_n8300_8799.n162 80.9324
R277 a_n8300_8799.n51 a_n8300_8799.n155 80.9324
R278 a_n8300_8799.n51 a_n8300_8799.n154 80.9324
R279 a_n8300_8799.n49 a_n8300_8799.n160 80.9324
R280 a_n8300_8799.n49 a_n8300_8799.n158 80.9324
R281 a_n8300_8799.n48 a_n8300_8799.n157 80.9324
R282 a_n8300_8799.n41 a_n8300_8799.n228 70.4033
R283 a_n8300_8799.n33 a_n8300_8799.n247 70.4033
R284 a_n8300_8799.n25 a_n8300_8799.n267 70.4033
R285 a_n8300_8799.n167 a_n8300_8799.n23 70.4033
R286 a_n8300_8799.n186 a_n8300_8799.n15 70.4033
R287 a_n8300_8799.n206 a_n8300_8799.n7 70.4033
R288 a_n8300_8799.n239 a_n8300_8799.n238 48.2005
R289 a_n8300_8799.n60 a_n8300_8799.n236 20.9683
R290 a_n8300_8799.n235 a_n8300_8799.n234 48.2005
R291 a_n8300_8799.n65 a_n8300_8799.n232 20.9683
R292 a_n8300_8799.n231 a_n8300_8799.n230 48.2005
R293 a_n8300_8799.n258 a_n8300_8799.n257 48.2005
R294 a_n8300_8799.n75 a_n8300_8799.n255 20.9683
R295 a_n8300_8799.n254 a_n8300_8799.n253 48.2005
R296 a_n8300_8799.n80 a_n8300_8799.n251 20.9683
R297 a_n8300_8799.n250 a_n8300_8799.n249 48.2005
R298 a_n8300_8799.n278 a_n8300_8799.n277 48.2005
R299 a_n8300_8799.n90 a_n8300_8799.n275 20.9683
R300 a_n8300_8799.n274 a_n8300_8799.n273 48.2005
R301 a_n8300_8799.n95 a_n8300_8799.n271 20.9683
R302 a_n8300_8799.n270 a_n8300_8799.n269 48.2005
R303 a_n8300_8799.n171 a_n8300_8799.n170 48.2005
R304 a_n8300_8799.n173 a_n8300_8799.n104 20.9683
R305 a_n8300_8799.n175 a_n8300_8799.n165 48.2005
R306 a_n8300_8799.n177 a_n8300_8799.n109 20.9683
R307 a_n8300_8799.n180 a_n8300_8799.n179 48.2005
R308 a_n8300_8799.t47 a_n8300_8799.n114 485.135
R309 a_n8300_8799.n190 a_n8300_8799.n189 48.2005
R310 a_n8300_8799.n192 a_n8300_8799.n119 20.9683
R311 a_n8300_8799.n194 a_n8300_8799.n184 48.2005
R312 a_n8300_8799.n196 a_n8300_8799.n124 20.9683
R313 a_n8300_8799.n199 a_n8300_8799.n198 48.2005
R314 a_n8300_8799.t59 a_n8300_8799.n129 485.135
R315 a_n8300_8799.n210 a_n8300_8799.n209 48.2005
R316 a_n8300_8799.n212 a_n8300_8799.n134 20.9683
R317 a_n8300_8799.n214 a_n8300_8799.n204 48.2005
R318 a_n8300_8799.n216 a_n8300_8799.n139 20.9683
R319 a_n8300_8799.n219 a_n8300_8799.n218 48.2005
R320 a_n8300_8799.t126 a_n8300_8799.n144 485.135
R321 a_n8300_8799.n56 a_n8300_8799.n222 17.8606
R322 a_n8300_8799.n229 a_n8300_8799.n69 25.894
R323 a_n8300_8799.n71 a_n8300_8799.n241 17.8606
R324 a_n8300_8799.n248 a_n8300_8799.n84 25.894
R325 a_n8300_8799.n86 a_n8300_8799.n261 17.8606
R326 a_n8300_8799.n268 a_n8300_8799.n99 25.894
R327 a_n8300_8799.n181 a_n8300_8799.n113 25.894
R328 a_n8300_8799.n200 a_n8300_8799.n128 25.894
R329 a_n8300_8799.n220 a_n8300_8799.n143 25.894
R330 a_n8300_8799.n67 a_n8300_8799.n226 43.3183
R331 a_n8300_8799.n82 a_n8300_8799.n245 43.3183
R332 a_n8300_8799.n97 a_n8300_8799.n265 43.3183
R333 a_n8300_8799.n178 a_n8300_8799.n111 43.3183
R334 a_n8300_8799.n197 a_n8300_8799.n126 43.3183
R335 a_n8300_8799.n217 a_n8300_8799.n141 43.3183
R336 a_n8300_8799.n61 a_n8300_8799.n224 16.6962
R337 a_n8300_8799.n233 a_n8300_8799.n64 27.6507
R338 a_n8300_8799.n76 a_n8300_8799.n243 16.6962
R339 a_n8300_8799.n252 a_n8300_8799.n79 27.6507
R340 a_n8300_8799.n91 a_n8300_8799.n263 16.6962
R341 a_n8300_8799.n272 a_n8300_8799.n94 27.6507
R342 a_n8300_8799.n174 a_n8300_8799.n105 16.6962
R343 a_n8300_8799.n164 a_n8300_8799.n108 27.6507
R344 a_n8300_8799.n193 a_n8300_8799.n120 16.6962
R345 a_n8300_8799.n183 a_n8300_8799.n123 27.6507
R346 a_n8300_8799.n213 a_n8300_8799.n135 16.6962
R347 a_n8300_8799.n203 a_n8300_8799.n138 27.6507
R348 a_n8300_8799.n62 a_n8300_8799.n224 41.7634
R349 a_n8300_8799.n77 a_n8300_8799.n243 41.7634
R350 a_n8300_8799.n92 a_n8300_8799.n263 41.7634
R351 a_n8300_8799.n106 a_n8300_8799.n174 41.7634
R352 a_n8300_8799.n121 a_n8300_8799.n193 41.7634
R353 a_n8300_8799.n136 a_n8300_8799.n213 41.7634
R354 a_n8300_8799.n237 a_n8300_8799.n59 29.3885
R355 a_n8300_8799.n66 a_n8300_8799.n226 15.5127
R356 a_n8300_8799.n256 a_n8300_8799.n74 29.3885
R357 a_n8300_8799.n81 a_n8300_8799.n245 15.5127
R358 a_n8300_8799.n276 a_n8300_8799.n89 29.3885
R359 a_n8300_8799.n96 a_n8300_8799.n265 15.5127
R360 a_n8300_8799.n172 a_n8300_8799.n103 29.3885
R361 a_n8300_8799.n178 a_n8300_8799.n110 15.5127
R362 a_n8300_8799.n191 a_n8300_8799.n118 29.3885
R363 a_n8300_8799.n197 a_n8300_8799.n125 15.5127
R364 a_n8300_8799.n211 a_n8300_8799.n133 29.3885
R365 a_n8300_8799.n217 a_n8300_8799.n140 15.5127
R366 a_n8300_8799.n57 a_n8300_8799.n222 40.1848
R367 a_n8300_8799.n72 a_n8300_8799.n241 40.1848
R368 a_n8300_8799.n87 a_n8300_8799.n261 40.1848
R369 a_n8300_8799.n169 a_n8300_8799.n101 40.1848
R370 a_n8300_8799.n188 a_n8300_8799.n116 40.1848
R371 a_n8300_8799.n208 a_n8300_8799.n131 40.1848
R372 a_n8300_8799.n50 a_n8300_8799.n49 31.9767
R373 a_n8300_8799.n283 a_n8300_8799.n152 31.5713
R374 a_n8300_8799.n229 a_n8300_8799.n228 20.9576
R375 a_n8300_8799.n248 a_n8300_8799.n247 20.9576
R376 a_n8300_8799.n268 a_n8300_8799.n267 20.9576
R377 a_n8300_8799.n168 a_n8300_8799.n167 20.9576
R378 a_n8300_8799.n187 a_n8300_8799.n186 20.9576
R379 a_n8300_8799.n207 a_n8300_8799.n206 20.9576
R380 a_n8300_8799.n54 a_n8300_8799.n283 19.0249
R381 a_n8300_8799.n57 a_n8300_8799.n239 7.32118
R382 a_n8300_8799.n68 a_n8300_8799.n227 40.1848
R383 a_n8300_8799.n72 a_n8300_8799.n258 7.32118
R384 a_n8300_8799.n83 a_n8300_8799.n246 40.1848
R385 a_n8300_8799.n87 a_n8300_8799.n278 7.32118
R386 a_n8300_8799.n98 a_n8300_8799.n266 40.1848
R387 a_n8300_8799.n170 a_n8300_8799.n101 7.32118
R388 a_n8300_8799.n163 a_n8300_8799.n112 40.1848
R389 a_n8300_8799.n189 a_n8300_8799.n116 7.32118
R390 a_n8300_8799.n182 a_n8300_8799.n127 40.1848
R391 a_n8300_8799.n209 a_n8300_8799.n131 7.32118
R392 a_n8300_8799.n202 a_n8300_8799.n142 40.1848
R393 a_n8300_8799.n232 a_n8300_8799.n66 29.3885
R394 a_n8300_8799.n251 a_n8300_8799.n81 29.3885
R395 a_n8300_8799.n271 a_n8300_8799.n96 29.3885
R396 a_n8300_8799.n110 a_n8300_8799.n177 29.3885
R397 a_n8300_8799.n125 a_n8300_8799.n196 29.3885
R398 a_n8300_8799.n140 a_n8300_8799.n216 29.3885
R399 a_n8300_8799.n62 a_n8300_8799.n235 5.97853
R400 a_n8300_8799.n63 a_n8300_8799.n225 41.7634
R401 a_n8300_8799.n77 a_n8300_8799.n254 5.97853
R402 a_n8300_8799.n78 a_n8300_8799.n244 41.7634
R403 a_n8300_8799.n92 a_n8300_8799.n274 5.97853
R404 a_n8300_8799.n93 a_n8300_8799.n264 41.7634
R405 a_n8300_8799.n175 a_n8300_8799.n106 5.97853
R406 a_n8300_8799.n176 a_n8300_8799.n107 41.7634
R407 a_n8300_8799.n194 a_n8300_8799.n121 5.97853
R408 a_n8300_8799.n195 a_n8300_8799.n122 41.7634
R409 a_n8300_8799.n214 a_n8300_8799.n136 5.97853
R410 a_n8300_8799.n215 a_n8300_8799.n137 41.7634
R411 a_n8300_8799.n282 a_n8300_8799.n51 12.3339
R412 a_n8300_8799.n283 a_n8300_8799.n282 11.4887
R413 a_n8300_8799.n236 a_n8300_8799.n61 27.6507
R414 a_n8300_8799.n255 a_n8300_8799.n76 27.6507
R415 a_n8300_8799.n275 a_n8300_8799.n91 27.6507
R416 a_n8300_8799.n173 a_n8300_8799.n105 27.6507
R417 a_n8300_8799.n192 a_n8300_8799.n120 27.6507
R418 a_n8300_8799.n212 a_n8300_8799.n135 27.6507
R419 a_n8300_8799.n58 a_n8300_8799.n223 43.3183
R420 a_n8300_8799.n67 a_n8300_8799.n231 4.61226
R421 a_n8300_8799.n73 a_n8300_8799.n242 43.3183
R422 a_n8300_8799.n82 a_n8300_8799.n250 4.61226
R423 a_n8300_8799.n88 a_n8300_8799.n262 43.3183
R424 a_n8300_8799.n97 a_n8300_8799.n270 4.61226
R425 a_n8300_8799.n166 a_n8300_8799.n102 43.3183
R426 a_n8300_8799.n179 a_n8300_8799.n111 4.61226
R427 a_n8300_8799.n185 a_n8300_8799.n117 43.3183
R428 a_n8300_8799.n198 a_n8300_8799.n126 4.61226
R429 a_n8300_8799.n205 a_n8300_8799.n132 43.3183
R430 a_n8300_8799.n218 a_n8300_8799.n141 4.61226
R431 a_n8300_8799.n260 a_n8300_8799.n47 9.04406
R432 a_n8300_8799.n201 a_n8300_8799.n17 9.04406
R433 a_n8300_8799.n240 a_n8300_8799.n56 25.894
R434 a_n8300_8799.n259 a_n8300_8799.n71 25.894
R435 a_n8300_8799.n279 a_n8300_8799.n86 25.894
R436 a_n8300_8799.n100 a_n8300_8799.n168 25.894
R437 a_n8300_8799.n115 a_n8300_8799.n187 25.894
R438 a_n8300_8799.n130 a_n8300_8799.n207 25.894
R439 a_n8300_8799.n281 a_n8300_8799.n221 6.94254
R440 a_n8300_8799.n281 a_n8300_8799.n280 6.64832
R441 a_n8300_8799.n260 a_n8300_8799.n39 4.93611
R442 a_n8300_8799.n280 a_n8300_8799.n31 4.93611
R443 a_n8300_8799.n201 a_n8300_8799.n9 4.93611
R444 a_n8300_8799.n221 a_n8300_8799.n1 4.93611
R445 a_n8300_8799.n280 a_n8300_8799.n260 4.10845
R446 a_n8300_8799.n221 a_n8300_8799.n201 4.10845
R447 a_n8300_8799.n147 a_n8300_8799.t7 3.61217
R448 a_n8300_8799.n147 a_n8300_8799.t19 3.61217
R449 a_n8300_8799.n146 a_n8300_8799.t32 3.61217
R450 a_n8300_8799.n146 a_n8300_8799.t22 3.61217
R451 a_n8300_8799.n145 a_n8300_8799.t11 3.61217
R452 a_n8300_8799.n145 a_n8300_8799.t29 3.61217
R453 a_n8300_8799.n148 a_n8300_8799.t17 3.61217
R454 a_n8300_8799.n148 a_n8300_8799.t2 3.61217
R455 a_n8300_8799.n149 a_n8300_8799.t23 3.61217
R456 a_n8300_8799.n149 a_n8300_8799.t28 3.61217
R457 a_n8300_8799.n150 a_n8300_8799.t13 3.61217
R458 a_n8300_8799.n150 a_n8300_8799.t20 3.61217
R459 a_n8300_8799.n151 a_n8300_8799.t18 3.61217
R460 a_n8300_8799.n151 a_n8300_8799.t21 3.61217
R461 a_n8300_8799.n284 a_n8300_8799.t12 3.61217
R462 a_n8300_8799.t1 a_n8300_8799.n284 3.61217
R463 a_n8300_8799.n282 a_n8300_8799.n281 3.4105
R464 a_n8300_8799.n161 a_n8300_8799.t6 2.82907
R465 a_n8300_8799.n161 a_n8300_8799.t27 2.82907
R466 a_n8300_8799.n162 a_n8300_8799.t34 2.82907
R467 a_n8300_8799.n162 a_n8300_8799.t5 2.82907
R468 a_n8300_8799.n155 a_n8300_8799.t14 2.82907
R469 a_n8300_8799.n155 a_n8300_8799.t4 2.82907
R470 a_n8300_8799.n154 a_n8300_8799.t24 2.82907
R471 a_n8300_8799.n154 a_n8300_8799.t0 2.82907
R472 a_n8300_8799.n153 a_n8300_8799.t25 2.82907
R473 a_n8300_8799.n153 a_n8300_8799.t30 2.82907
R474 a_n8300_8799.n159 a_n8300_8799.t8 2.82907
R475 a_n8300_8799.n159 a_n8300_8799.t15 2.82907
R476 a_n8300_8799.n160 a_n8300_8799.t26 2.82907
R477 a_n8300_8799.n160 a_n8300_8799.t33 2.82907
R478 a_n8300_8799.n158 a_n8300_8799.t31 2.82907
R479 a_n8300_8799.n158 a_n8300_8799.t10 2.82907
R480 a_n8300_8799.n157 a_n8300_8799.t35 2.82907
R481 a_n8300_8799.n157 a_n8300_8799.t9 2.82907
R482 a_n8300_8799.n156 a_n8300_8799.t3 2.82907
R483 a_n8300_8799.n156 a_n8300_8799.t16 2.82907
R484 a_n8300_8799.n41 a_n8300_8799.n40 1.13686
R485 a_n8300_8799.n33 a_n8300_8799.n32 1.13686
R486 a_n8300_8799.n25 a_n8300_8799.n24 1.13686
R487 a_n8300_8799.n17 a_n8300_8799.n16 1.13686
R488 a_n8300_8799.n9 a_n8300_8799.n8 1.13686
R489 a_n8300_8799.n1 a_n8300_8799.n0 1.13686
R490 a_n8300_8799.n51 a_n8300_8799.n50 1.07378
R491 a_n8300_8799.n46 a_n8300_8799.n45 0.758076
R492 a_n8300_8799.n46 a_n8300_8799.n44 0.758076
R493 a_n8300_8799.n44 a_n8300_8799.n43 0.758076
R494 a_n8300_8799.n43 a_n8300_8799.n42 0.758076
R495 a_n8300_8799.n40 a_n8300_8799.n42 0.758076
R496 a_n8300_8799.n38 a_n8300_8799.n37 0.758076
R497 a_n8300_8799.n38 a_n8300_8799.n36 0.758076
R498 a_n8300_8799.n36 a_n8300_8799.n35 0.758076
R499 a_n8300_8799.n35 a_n8300_8799.n34 0.758076
R500 a_n8300_8799.n32 a_n8300_8799.n34 0.758076
R501 a_n8300_8799.n30 a_n8300_8799.n29 0.758076
R502 a_n8300_8799.n30 a_n8300_8799.n28 0.758076
R503 a_n8300_8799.n28 a_n8300_8799.n27 0.758076
R504 a_n8300_8799.n27 a_n8300_8799.n26 0.758076
R505 a_n8300_8799.n24 a_n8300_8799.n26 0.758076
R506 a_n8300_8799.n21 a_n8300_8799.n22 0.758076
R507 a_n8300_8799.n20 a_n8300_8799.n21 0.758076
R508 a_n8300_8799.n19 a_n8300_8799.n20 0.758076
R509 a_n8300_8799.n18 a_n8300_8799.n19 0.758076
R510 a_n8300_8799.n16 a_n8300_8799.n18 0.758076
R511 a_n8300_8799.n13 a_n8300_8799.n14 0.758076
R512 a_n8300_8799.n12 a_n8300_8799.n13 0.758076
R513 a_n8300_8799.n11 a_n8300_8799.n12 0.758076
R514 a_n8300_8799.n10 a_n8300_8799.n11 0.758076
R515 a_n8300_8799.n8 a_n8300_8799.n10 0.758076
R516 a_n8300_8799.n5 a_n8300_8799.n6 0.758076
R517 a_n8300_8799.n4 a_n8300_8799.n5 0.758076
R518 a_n8300_8799.n3 a_n8300_8799.n4 0.758076
R519 a_n8300_8799.n2 a_n8300_8799.n3 0.758076
R520 a_n8300_8799.n0 a_n8300_8799.n2 0.758076
R521 a_n8300_8799.n54 a_n8300_8799.n53 0.716017
R522 a_n8300_8799.n152 a_n8300_8799.n52 0.716017
R523 a_n8300_8799.n49 a_n8300_8799.n48 0.716017
R524 a_n8300_8799.n6 a_n8300_8799.n7 0.568682
R525 a_n8300_8799.n14 a_n8300_8799.n15 0.568682
R526 a_n8300_8799.n22 a_n8300_8799.n23 0.568682
R527 a_n8300_8799.n29 a_n8300_8799.n31 0.568682
R528 a_n8300_8799.n37 a_n8300_8799.n39 0.568682
R529 a_n8300_8799.n45 a_n8300_8799.n47 0.568682
R530 vdd.n327 vdd.n291 756.745
R531 vdd.n268 vdd.n232 756.745
R532 vdd.n225 vdd.n189 756.745
R533 vdd.n166 vdd.n130 756.745
R534 vdd.n124 vdd.n88 756.745
R535 vdd.n65 vdd.n29 756.745
R536 vdd.n2108 vdd.n2072 756.745
R537 vdd.n2167 vdd.n2131 756.745
R538 vdd.n2006 vdd.n1970 756.745
R539 vdd.n2065 vdd.n2029 756.745
R540 vdd.n1905 vdd.n1869 756.745
R541 vdd.n1964 vdd.n1928 756.745
R542 vdd.n1253 vdd.t228 640.208
R543 vdd.n981 vdd.t270 640.208
R544 vdd.n1273 vdd.t243 640.208
R545 vdd.n972 vdd.t294 640.208
R546 vdd.n872 vdd.t250 640.208
R547 vdd.n2704 vdd.t288 640.208
R548 vdd.n832 vdd.t297 640.208
R549 vdd.n2701 vdd.t274 640.208
R550 vdd.n799 vdd.t224 640.208
R551 vdd.n1043 vdd.t281 640.208
R552 vdd.n1679 vdd.t260 592.009
R553 vdd.n1717 vdd.t278 592.009
R554 vdd.n1613 vdd.t291 592.009
R555 vdd.n2269 vdd.t236 592.009
R556 vdd.n1190 vdd.t267 592.009
R557 vdd.n1150 vdd.t285 592.009
R558 vdd.n426 vdd.t257 592.009
R559 vdd.n440 vdd.t246 592.009
R560 vdd.n452 vdd.t264 592.009
R561 vdd.n768 vdd.t240 592.009
R562 vdd.n3276 vdd.t254 592.009
R563 vdd.n688 vdd.t232 592.009
R564 vdd.n328 vdd.n327 585
R565 vdd.n326 vdd.n293 585
R566 vdd.n325 vdd.n324 585
R567 vdd.n296 vdd.n294 585
R568 vdd.n319 vdd.n318 585
R569 vdd.n317 vdd.n316 585
R570 vdd.n300 vdd.n299 585
R571 vdd.n311 vdd.n310 585
R572 vdd.n309 vdd.n308 585
R573 vdd.n304 vdd.n303 585
R574 vdd.n269 vdd.n268 585
R575 vdd.n267 vdd.n234 585
R576 vdd.n266 vdd.n265 585
R577 vdd.n237 vdd.n235 585
R578 vdd.n260 vdd.n259 585
R579 vdd.n258 vdd.n257 585
R580 vdd.n241 vdd.n240 585
R581 vdd.n252 vdd.n251 585
R582 vdd.n250 vdd.n249 585
R583 vdd.n245 vdd.n244 585
R584 vdd.n226 vdd.n225 585
R585 vdd.n224 vdd.n191 585
R586 vdd.n223 vdd.n222 585
R587 vdd.n194 vdd.n192 585
R588 vdd.n217 vdd.n216 585
R589 vdd.n215 vdd.n214 585
R590 vdd.n198 vdd.n197 585
R591 vdd.n209 vdd.n208 585
R592 vdd.n207 vdd.n206 585
R593 vdd.n202 vdd.n201 585
R594 vdd.n167 vdd.n166 585
R595 vdd.n165 vdd.n132 585
R596 vdd.n164 vdd.n163 585
R597 vdd.n135 vdd.n133 585
R598 vdd.n158 vdd.n157 585
R599 vdd.n156 vdd.n155 585
R600 vdd.n139 vdd.n138 585
R601 vdd.n150 vdd.n149 585
R602 vdd.n148 vdd.n147 585
R603 vdd.n143 vdd.n142 585
R604 vdd.n125 vdd.n124 585
R605 vdd.n123 vdd.n90 585
R606 vdd.n122 vdd.n121 585
R607 vdd.n93 vdd.n91 585
R608 vdd.n116 vdd.n115 585
R609 vdd.n114 vdd.n113 585
R610 vdd.n97 vdd.n96 585
R611 vdd.n108 vdd.n107 585
R612 vdd.n106 vdd.n105 585
R613 vdd.n101 vdd.n100 585
R614 vdd.n66 vdd.n65 585
R615 vdd.n64 vdd.n31 585
R616 vdd.n63 vdd.n62 585
R617 vdd.n34 vdd.n32 585
R618 vdd.n57 vdd.n56 585
R619 vdd.n55 vdd.n54 585
R620 vdd.n38 vdd.n37 585
R621 vdd.n49 vdd.n48 585
R622 vdd.n47 vdd.n46 585
R623 vdd.n42 vdd.n41 585
R624 vdd.n2109 vdd.n2108 585
R625 vdd.n2107 vdd.n2074 585
R626 vdd.n2106 vdd.n2105 585
R627 vdd.n2077 vdd.n2075 585
R628 vdd.n2100 vdd.n2099 585
R629 vdd.n2098 vdd.n2097 585
R630 vdd.n2081 vdd.n2080 585
R631 vdd.n2092 vdd.n2091 585
R632 vdd.n2090 vdd.n2089 585
R633 vdd.n2085 vdd.n2084 585
R634 vdd.n2168 vdd.n2167 585
R635 vdd.n2166 vdd.n2133 585
R636 vdd.n2165 vdd.n2164 585
R637 vdd.n2136 vdd.n2134 585
R638 vdd.n2159 vdd.n2158 585
R639 vdd.n2157 vdd.n2156 585
R640 vdd.n2140 vdd.n2139 585
R641 vdd.n2151 vdd.n2150 585
R642 vdd.n2149 vdd.n2148 585
R643 vdd.n2144 vdd.n2143 585
R644 vdd.n2007 vdd.n2006 585
R645 vdd.n2005 vdd.n1972 585
R646 vdd.n2004 vdd.n2003 585
R647 vdd.n1975 vdd.n1973 585
R648 vdd.n1998 vdd.n1997 585
R649 vdd.n1996 vdd.n1995 585
R650 vdd.n1979 vdd.n1978 585
R651 vdd.n1990 vdd.n1989 585
R652 vdd.n1988 vdd.n1987 585
R653 vdd.n1983 vdd.n1982 585
R654 vdd.n2066 vdd.n2065 585
R655 vdd.n2064 vdd.n2031 585
R656 vdd.n2063 vdd.n2062 585
R657 vdd.n2034 vdd.n2032 585
R658 vdd.n2057 vdd.n2056 585
R659 vdd.n2055 vdd.n2054 585
R660 vdd.n2038 vdd.n2037 585
R661 vdd.n2049 vdd.n2048 585
R662 vdd.n2047 vdd.n2046 585
R663 vdd.n2042 vdd.n2041 585
R664 vdd.n1906 vdd.n1905 585
R665 vdd.n1904 vdd.n1871 585
R666 vdd.n1903 vdd.n1902 585
R667 vdd.n1874 vdd.n1872 585
R668 vdd.n1897 vdd.n1896 585
R669 vdd.n1895 vdd.n1894 585
R670 vdd.n1878 vdd.n1877 585
R671 vdd.n1889 vdd.n1888 585
R672 vdd.n1887 vdd.n1886 585
R673 vdd.n1882 vdd.n1881 585
R674 vdd.n1965 vdd.n1964 585
R675 vdd.n1963 vdd.n1930 585
R676 vdd.n1962 vdd.n1961 585
R677 vdd.n1933 vdd.n1931 585
R678 vdd.n1956 vdd.n1955 585
R679 vdd.n1954 vdd.n1953 585
R680 vdd.n1937 vdd.n1936 585
R681 vdd.n1948 vdd.n1947 585
R682 vdd.n1946 vdd.n1945 585
R683 vdd.n1941 vdd.n1940 585
R684 vdd.n3448 vdd.n392 509.269
R685 vdd.n3444 vdd.n393 509.269
R686 vdd.n3316 vdd.n685 509.269
R687 vdd.n3313 vdd.n684 509.269
R688 vdd.n2264 vdd.n1437 509.269
R689 vdd.n2267 vdd.n2266 509.269
R690 vdd.n1586 vdd.n1550 509.269
R691 vdd.n1782 vdd.n1551 509.269
R692 vdd.n305 vdd.t88 329.043
R693 vdd.n246 vdd.t168 329.043
R694 vdd.n203 vdd.t219 329.043
R695 vdd.n144 vdd.t152 329.043
R696 vdd.n102 vdd.t120 329.043
R697 vdd.n43 vdd.t113 329.043
R698 vdd.n2086 vdd.t210 329.043
R699 vdd.n2145 vdd.t144 329.043
R700 vdd.n1984 vdd.t198 329.043
R701 vdd.n2043 vdd.t121 329.043
R702 vdd.n1883 vdd.t115 329.043
R703 vdd.n1942 vdd.t73 329.043
R704 vdd.n1679 vdd.t263 319.788
R705 vdd.n1717 vdd.t280 319.788
R706 vdd.n1613 vdd.t293 319.788
R707 vdd.n2269 vdd.t238 319.788
R708 vdd.n1190 vdd.t268 319.788
R709 vdd.n1150 vdd.t286 319.788
R710 vdd.n426 vdd.t258 319.788
R711 vdd.n440 vdd.t248 319.788
R712 vdd.n452 vdd.t265 319.788
R713 vdd.n768 vdd.t242 319.788
R714 vdd.n3276 vdd.t256 319.788
R715 vdd.n688 vdd.t235 319.788
R716 vdd.n1680 vdd.t262 303.69
R717 vdd.n1718 vdd.t279 303.69
R718 vdd.n1614 vdd.t292 303.69
R719 vdd.n2270 vdd.t239 303.69
R720 vdd.n1191 vdd.t269 303.69
R721 vdd.n1151 vdd.t287 303.69
R722 vdd.n427 vdd.t259 303.69
R723 vdd.n441 vdd.t249 303.69
R724 vdd.n453 vdd.t266 303.69
R725 vdd.n769 vdd.t241 303.69
R726 vdd.n3277 vdd.t255 303.69
R727 vdd.n689 vdd.t234 303.69
R728 vdd.n2936 vdd.n927 291.221
R729 vdd.n3150 vdd.n809 291.221
R730 vdd.n3087 vdd.n806 291.221
R731 vdd.n2868 vdd.n2867 291.221
R732 vdd.n2664 vdd.n969 291.221
R733 vdd.n2595 vdd.n2594 291.221
R734 vdd.n1309 vdd.n1308 291.221
R735 vdd.n2415 vdd.n1075 291.221
R736 vdd.n3066 vdd.n807 291.221
R737 vdd.n3153 vdd.n3152 291.221
R738 vdd.n2772 vdd.n2698 291.221
R739 vdd.n2940 vdd.n931 291.221
R740 vdd.n2592 vdd.n979 291.221
R741 vdd.n977 vdd.n951 291.221
R742 vdd.n1387 vdd.n1116 291.221
R743 vdd.n2419 vdd.n1080 291.221
R744 vdd.n3068 vdd.n807 185
R745 vdd.n3151 vdd.n807 185
R746 vdd.n3070 vdd.n3069 185
R747 vdd.n3069 vdd.n805 185
R748 vdd.n3071 vdd.n839 185
R749 vdd.n3081 vdd.n839 185
R750 vdd.n3072 vdd.n848 185
R751 vdd.n848 vdd.n846 185
R752 vdd.n3074 vdd.n3073 185
R753 vdd.n3075 vdd.n3074 185
R754 vdd.n3027 vdd.n847 185
R755 vdd.n847 vdd.n843 185
R756 vdd.n3026 vdd.n3025 185
R757 vdd.n3025 vdd.n3024 185
R758 vdd.n850 vdd.n849 185
R759 vdd.n851 vdd.n850 185
R760 vdd.n3017 vdd.n3016 185
R761 vdd.n3018 vdd.n3017 185
R762 vdd.n3015 vdd.n860 185
R763 vdd.n860 vdd.n857 185
R764 vdd.n3014 vdd.n3013 185
R765 vdd.n3013 vdd.n3012 185
R766 vdd.n862 vdd.n861 185
R767 vdd.n870 vdd.n862 185
R768 vdd.n3005 vdd.n3004 185
R769 vdd.n3006 vdd.n3005 185
R770 vdd.n3002 vdd.n871 185
R771 vdd.n878 vdd.n871 185
R772 vdd.n3001 vdd.n3000 185
R773 vdd.n3000 vdd.n2999 185
R774 vdd.n874 vdd.n873 185
R775 vdd.n875 vdd.n874 185
R776 vdd.n2992 vdd.n2991 185
R777 vdd.n2993 vdd.n2992 185
R778 vdd.n2990 vdd.n885 185
R779 vdd.n885 vdd.n882 185
R780 vdd.n2989 vdd.n2988 185
R781 vdd.n2988 vdd.n2987 185
R782 vdd.n887 vdd.n886 185
R783 vdd.n895 vdd.n887 185
R784 vdd.n2980 vdd.n2979 185
R785 vdd.n2981 vdd.n2980 185
R786 vdd.n2978 vdd.n896 185
R787 vdd.n901 vdd.n896 185
R788 vdd.n2977 vdd.n2976 185
R789 vdd.n2976 vdd.n2975 185
R790 vdd.n898 vdd.n897 185
R791 vdd.n2847 vdd.n898 185
R792 vdd.n2968 vdd.n2967 185
R793 vdd.n2969 vdd.n2968 185
R794 vdd.n2966 vdd.n908 185
R795 vdd.n908 vdd.n905 185
R796 vdd.n2965 vdd.n2964 185
R797 vdd.n2964 vdd.n2963 185
R798 vdd.n910 vdd.n909 185
R799 vdd.n911 vdd.n910 185
R800 vdd.n2956 vdd.n2955 185
R801 vdd.n2957 vdd.n2956 185
R802 vdd.n2954 vdd.n920 185
R803 vdd.n920 vdd.n917 185
R804 vdd.n2953 vdd.n2952 185
R805 vdd.n2952 vdd.n2951 185
R806 vdd.n922 vdd.n921 185
R807 vdd.n2862 vdd.n922 185
R808 vdd.n2944 vdd.n2943 185
R809 vdd.n2945 vdd.n2944 185
R810 vdd.n2942 vdd.n931 185
R811 vdd.n931 vdd.n928 185
R812 vdd.n2941 vdd.n2940 185
R813 vdd.n933 vdd.n932 185
R814 vdd.n2708 vdd.n2707 185
R815 vdd.n2710 vdd.n2709 185
R816 vdd.n2712 vdd.n2711 185
R817 vdd.n2714 vdd.n2713 185
R818 vdd.n2716 vdd.n2715 185
R819 vdd.n2718 vdd.n2717 185
R820 vdd.n2720 vdd.n2719 185
R821 vdd.n2722 vdd.n2721 185
R822 vdd.n2724 vdd.n2723 185
R823 vdd.n2726 vdd.n2725 185
R824 vdd.n2728 vdd.n2727 185
R825 vdd.n2730 vdd.n2729 185
R826 vdd.n2732 vdd.n2731 185
R827 vdd.n2734 vdd.n2733 185
R828 vdd.n2736 vdd.n2735 185
R829 vdd.n2738 vdd.n2737 185
R830 vdd.n2740 vdd.n2739 185
R831 vdd.n2742 vdd.n2741 185
R832 vdd.n2744 vdd.n2743 185
R833 vdd.n2746 vdd.n2745 185
R834 vdd.n2748 vdd.n2747 185
R835 vdd.n2750 vdd.n2749 185
R836 vdd.n2752 vdd.n2751 185
R837 vdd.n2754 vdd.n2753 185
R838 vdd.n2756 vdd.n2755 185
R839 vdd.n2758 vdd.n2757 185
R840 vdd.n2760 vdd.n2759 185
R841 vdd.n2762 vdd.n2761 185
R842 vdd.n2764 vdd.n2763 185
R843 vdd.n2766 vdd.n2765 185
R844 vdd.n2768 vdd.n2767 185
R845 vdd.n2770 vdd.n2769 185
R846 vdd.n2771 vdd.n2698 185
R847 vdd.n2938 vdd.n2698 185
R848 vdd.n3154 vdd.n3153 185
R849 vdd.n3155 vdd.n798 185
R850 vdd.n3157 vdd.n3156 185
R851 vdd.n3159 vdd.n796 185
R852 vdd.n3161 vdd.n3160 185
R853 vdd.n3162 vdd.n795 185
R854 vdd.n3164 vdd.n3163 185
R855 vdd.n3166 vdd.n793 185
R856 vdd.n3168 vdd.n3167 185
R857 vdd.n3169 vdd.n792 185
R858 vdd.n3171 vdd.n3170 185
R859 vdd.n3173 vdd.n790 185
R860 vdd.n3175 vdd.n3174 185
R861 vdd.n3176 vdd.n789 185
R862 vdd.n3178 vdd.n3177 185
R863 vdd.n3180 vdd.n788 185
R864 vdd.n3181 vdd.n786 185
R865 vdd.n3184 vdd.n3183 185
R866 vdd.n787 vdd.n785 185
R867 vdd.n3040 vdd.n3039 185
R868 vdd.n3042 vdd.n3041 185
R869 vdd.n3044 vdd.n3036 185
R870 vdd.n3046 vdd.n3045 185
R871 vdd.n3047 vdd.n3035 185
R872 vdd.n3049 vdd.n3048 185
R873 vdd.n3051 vdd.n3033 185
R874 vdd.n3053 vdd.n3052 185
R875 vdd.n3054 vdd.n3032 185
R876 vdd.n3056 vdd.n3055 185
R877 vdd.n3058 vdd.n3030 185
R878 vdd.n3060 vdd.n3059 185
R879 vdd.n3061 vdd.n3029 185
R880 vdd.n3063 vdd.n3062 185
R881 vdd.n3065 vdd.n3028 185
R882 vdd.n3067 vdd.n3066 185
R883 vdd.n3066 vdd.n692 185
R884 vdd.n3152 vdd.n802 185
R885 vdd.n3152 vdd.n3151 185
R886 vdd.n2775 vdd.n804 185
R887 vdd.n805 vdd.n804 185
R888 vdd.n2776 vdd.n838 185
R889 vdd.n3081 vdd.n838 185
R890 vdd.n2778 vdd.n2777 185
R891 vdd.n2777 vdd.n846 185
R892 vdd.n2779 vdd.n845 185
R893 vdd.n3075 vdd.n845 185
R894 vdd.n2781 vdd.n2780 185
R895 vdd.n2780 vdd.n843 185
R896 vdd.n2782 vdd.n853 185
R897 vdd.n3024 vdd.n853 185
R898 vdd.n2784 vdd.n2783 185
R899 vdd.n2783 vdd.n851 185
R900 vdd.n2785 vdd.n859 185
R901 vdd.n3018 vdd.n859 185
R902 vdd.n2787 vdd.n2786 185
R903 vdd.n2786 vdd.n857 185
R904 vdd.n2788 vdd.n864 185
R905 vdd.n3012 vdd.n864 185
R906 vdd.n2790 vdd.n2789 185
R907 vdd.n2789 vdd.n870 185
R908 vdd.n2791 vdd.n869 185
R909 vdd.n3006 vdd.n869 185
R910 vdd.n2793 vdd.n2792 185
R911 vdd.n2792 vdd.n878 185
R912 vdd.n2794 vdd.n877 185
R913 vdd.n2999 vdd.n877 185
R914 vdd.n2796 vdd.n2795 185
R915 vdd.n2795 vdd.n875 185
R916 vdd.n2797 vdd.n884 185
R917 vdd.n2993 vdd.n884 185
R918 vdd.n2799 vdd.n2798 185
R919 vdd.n2798 vdd.n882 185
R920 vdd.n2800 vdd.n889 185
R921 vdd.n2987 vdd.n889 185
R922 vdd.n2802 vdd.n2801 185
R923 vdd.n2801 vdd.n895 185
R924 vdd.n2803 vdd.n894 185
R925 vdd.n2981 vdd.n894 185
R926 vdd.n2805 vdd.n2804 185
R927 vdd.n2804 vdd.n901 185
R928 vdd.n2806 vdd.n900 185
R929 vdd.n2975 vdd.n900 185
R930 vdd.n2849 vdd.n2848 185
R931 vdd.n2848 vdd.n2847 185
R932 vdd.n2850 vdd.n907 185
R933 vdd.n2969 vdd.n907 185
R934 vdd.n2852 vdd.n2851 185
R935 vdd.n2851 vdd.n905 185
R936 vdd.n2853 vdd.n913 185
R937 vdd.n2963 vdd.n913 185
R938 vdd.n2855 vdd.n2854 185
R939 vdd.n2854 vdd.n911 185
R940 vdd.n2856 vdd.n919 185
R941 vdd.n2957 vdd.n919 185
R942 vdd.n2858 vdd.n2857 185
R943 vdd.n2857 vdd.n917 185
R944 vdd.n2859 vdd.n924 185
R945 vdd.n2951 vdd.n924 185
R946 vdd.n2861 vdd.n2860 185
R947 vdd.n2862 vdd.n2861 185
R948 vdd.n2774 vdd.n930 185
R949 vdd.n2945 vdd.n930 185
R950 vdd.n2773 vdd.n2772 185
R951 vdd.n2772 vdd.n928 185
R952 vdd.n2264 vdd.n2263 185
R953 vdd.n2265 vdd.n2264 185
R954 vdd.n1438 vdd.n1436 185
R955 vdd.n2256 vdd.n1436 185
R956 vdd.n2259 vdd.n2258 185
R957 vdd.n2258 vdd.n2257 185
R958 vdd.n1441 vdd.n1440 185
R959 vdd.n1442 vdd.n1441 185
R960 vdd.n2245 vdd.n2244 185
R961 vdd.n2246 vdd.n2245 185
R962 vdd.n1450 vdd.n1449 185
R963 vdd.n2237 vdd.n1449 185
R964 vdd.n2240 vdd.n2239 185
R965 vdd.n2239 vdd.n2238 185
R966 vdd.n1453 vdd.n1452 185
R967 vdd.n1460 vdd.n1453 185
R968 vdd.n2228 vdd.n2227 185
R969 vdd.n2229 vdd.n2228 185
R970 vdd.n1462 vdd.n1461 185
R971 vdd.n1461 vdd.n1459 185
R972 vdd.n2223 vdd.n2222 185
R973 vdd.n2222 vdd.n2221 185
R974 vdd.n1465 vdd.n1464 185
R975 vdd.n1466 vdd.n1465 185
R976 vdd.n2212 vdd.n2211 185
R977 vdd.n2213 vdd.n2212 185
R978 vdd.n1473 vdd.n1472 185
R979 vdd.n2204 vdd.n1472 185
R980 vdd.n2207 vdd.n2206 185
R981 vdd.n2206 vdd.n2205 185
R982 vdd.n1476 vdd.n1475 185
R983 vdd.n1482 vdd.n1476 185
R984 vdd.n2195 vdd.n2194 185
R985 vdd.n2196 vdd.n2195 185
R986 vdd.n1484 vdd.n1483 185
R987 vdd.n2187 vdd.n1483 185
R988 vdd.n2190 vdd.n2189 185
R989 vdd.n2189 vdd.n2188 185
R990 vdd.n1487 vdd.n1486 185
R991 vdd.n1488 vdd.n1487 185
R992 vdd.n2178 vdd.n2177 185
R993 vdd.n2179 vdd.n2178 185
R994 vdd.n1496 vdd.n1495 185
R995 vdd.n1495 vdd.n1494 185
R996 vdd.n1866 vdd.n1865 185
R997 vdd.n1865 vdd.n1864 185
R998 vdd.n1499 vdd.n1498 185
R999 vdd.n1505 vdd.n1499 185
R1000 vdd.n1855 vdd.n1854 185
R1001 vdd.n1856 vdd.n1855 185
R1002 vdd.n1507 vdd.n1506 185
R1003 vdd.n1847 vdd.n1506 185
R1004 vdd.n1850 vdd.n1849 185
R1005 vdd.n1849 vdd.n1848 185
R1006 vdd.n1510 vdd.n1509 185
R1007 vdd.n1517 vdd.n1510 185
R1008 vdd.n1838 vdd.n1837 185
R1009 vdd.n1839 vdd.n1838 185
R1010 vdd.n1519 vdd.n1518 185
R1011 vdd.n1518 vdd.n1516 185
R1012 vdd.n1833 vdd.n1832 185
R1013 vdd.n1832 vdd.n1831 185
R1014 vdd.n1522 vdd.n1521 185
R1015 vdd.n1523 vdd.n1522 185
R1016 vdd.n1822 vdd.n1821 185
R1017 vdd.n1823 vdd.n1822 185
R1018 vdd.n1530 vdd.n1529 185
R1019 vdd.n1814 vdd.n1529 185
R1020 vdd.n1817 vdd.n1816 185
R1021 vdd.n1816 vdd.n1815 185
R1022 vdd.n1533 vdd.n1532 185
R1023 vdd.n1539 vdd.n1533 185
R1024 vdd.n1805 vdd.n1804 185
R1025 vdd.n1806 vdd.n1805 185
R1026 vdd.n1541 vdd.n1540 185
R1027 vdd.n1797 vdd.n1540 185
R1028 vdd.n1800 vdd.n1799 185
R1029 vdd.n1799 vdd.n1798 185
R1030 vdd.n1544 vdd.n1543 185
R1031 vdd.n1545 vdd.n1544 185
R1032 vdd.n1788 vdd.n1787 185
R1033 vdd.n1789 vdd.n1788 185
R1034 vdd.n1552 vdd.n1551 185
R1035 vdd.n1587 vdd.n1551 185
R1036 vdd.n1783 vdd.n1782 185
R1037 vdd.n1555 vdd.n1554 185
R1038 vdd.n1779 vdd.n1778 185
R1039 vdd.n1780 vdd.n1779 185
R1040 vdd.n1589 vdd.n1588 185
R1041 vdd.n1774 vdd.n1591 185
R1042 vdd.n1773 vdd.n1592 185
R1043 vdd.n1772 vdd.n1593 185
R1044 vdd.n1595 vdd.n1594 185
R1045 vdd.n1768 vdd.n1597 185
R1046 vdd.n1767 vdd.n1598 185
R1047 vdd.n1766 vdd.n1599 185
R1048 vdd.n1601 vdd.n1600 185
R1049 vdd.n1762 vdd.n1603 185
R1050 vdd.n1761 vdd.n1604 185
R1051 vdd.n1760 vdd.n1605 185
R1052 vdd.n1607 vdd.n1606 185
R1053 vdd.n1756 vdd.n1609 185
R1054 vdd.n1755 vdd.n1610 185
R1055 vdd.n1754 vdd.n1611 185
R1056 vdd.n1615 vdd.n1612 185
R1057 vdd.n1750 vdd.n1617 185
R1058 vdd.n1749 vdd.n1618 185
R1059 vdd.n1748 vdd.n1619 185
R1060 vdd.n1621 vdd.n1620 185
R1061 vdd.n1744 vdd.n1623 185
R1062 vdd.n1743 vdd.n1624 185
R1063 vdd.n1742 vdd.n1625 185
R1064 vdd.n1627 vdd.n1626 185
R1065 vdd.n1738 vdd.n1629 185
R1066 vdd.n1737 vdd.n1630 185
R1067 vdd.n1736 vdd.n1631 185
R1068 vdd.n1633 vdd.n1632 185
R1069 vdd.n1732 vdd.n1635 185
R1070 vdd.n1731 vdd.n1636 185
R1071 vdd.n1730 vdd.n1637 185
R1072 vdd.n1639 vdd.n1638 185
R1073 vdd.n1726 vdd.n1641 185
R1074 vdd.n1725 vdd.n1642 185
R1075 vdd.n1724 vdd.n1643 185
R1076 vdd.n1645 vdd.n1644 185
R1077 vdd.n1720 vdd.n1647 185
R1078 vdd.n1719 vdd.n1716 185
R1079 vdd.n1715 vdd.n1648 185
R1080 vdd.n1650 vdd.n1649 185
R1081 vdd.n1711 vdd.n1652 185
R1082 vdd.n1710 vdd.n1653 185
R1083 vdd.n1709 vdd.n1654 185
R1084 vdd.n1656 vdd.n1655 185
R1085 vdd.n1705 vdd.n1658 185
R1086 vdd.n1704 vdd.n1659 185
R1087 vdd.n1703 vdd.n1660 185
R1088 vdd.n1662 vdd.n1661 185
R1089 vdd.n1699 vdd.n1664 185
R1090 vdd.n1698 vdd.n1665 185
R1091 vdd.n1697 vdd.n1666 185
R1092 vdd.n1668 vdd.n1667 185
R1093 vdd.n1693 vdd.n1670 185
R1094 vdd.n1692 vdd.n1671 185
R1095 vdd.n1691 vdd.n1672 185
R1096 vdd.n1674 vdd.n1673 185
R1097 vdd.n1687 vdd.n1676 185
R1098 vdd.n1686 vdd.n1677 185
R1099 vdd.n1685 vdd.n1678 185
R1100 vdd.n1682 vdd.n1586 185
R1101 vdd.n1780 vdd.n1586 185
R1102 vdd.n2268 vdd.n2267 185
R1103 vdd.n2272 vdd.n1432 185
R1104 vdd.n1431 vdd.n1425 185
R1105 vdd.n1429 vdd.n1428 185
R1106 vdd.n1427 vdd.n1221 185
R1107 vdd.n2276 vdd.n1218 185
R1108 vdd.n2278 vdd.n2277 185
R1109 vdd.n2280 vdd.n1216 185
R1110 vdd.n2282 vdd.n2281 185
R1111 vdd.n2283 vdd.n1211 185
R1112 vdd.n2285 vdd.n2284 185
R1113 vdd.n2287 vdd.n1209 185
R1114 vdd.n2289 vdd.n2288 185
R1115 vdd.n2290 vdd.n1204 185
R1116 vdd.n2292 vdd.n2291 185
R1117 vdd.n2294 vdd.n1202 185
R1118 vdd.n2296 vdd.n2295 185
R1119 vdd.n2297 vdd.n1198 185
R1120 vdd.n2299 vdd.n2298 185
R1121 vdd.n2301 vdd.n1195 185
R1122 vdd.n2303 vdd.n2302 185
R1123 vdd.n1196 vdd.n1189 185
R1124 vdd.n2307 vdd.n1193 185
R1125 vdd.n2308 vdd.n1185 185
R1126 vdd.n2310 vdd.n2309 185
R1127 vdd.n2312 vdd.n1183 185
R1128 vdd.n2314 vdd.n2313 185
R1129 vdd.n2315 vdd.n1178 185
R1130 vdd.n2317 vdd.n2316 185
R1131 vdd.n2319 vdd.n1176 185
R1132 vdd.n2321 vdd.n2320 185
R1133 vdd.n2322 vdd.n1171 185
R1134 vdd.n2324 vdd.n2323 185
R1135 vdd.n2326 vdd.n1169 185
R1136 vdd.n2328 vdd.n2327 185
R1137 vdd.n2329 vdd.n1164 185
R1138 vdd.n2331 vdd.n2330 185
R1139 vdd.n2333 vdd.n1162 185
R1140 vdd.n2335 vdd.n2334 185
R1141 vdd.n2336 vdd.n1158 185
R1142 vdd.n2338 vdd.n2337 185
R1143 vdd.n2340 vdd.n1155 185
R1144 vdd.n2342 vdd.n2341 185
R1145 vdd.n1156 vdd.n1149 185
R1146 vdd.n2346 vdd.n1153 185
R1147 vdd.n2347 vdd.n1145 185
R1148 vdd.n2349 vdd.n2348 185
R1149 vdd.n2351 vdd.n1143 185
R1150 vdd.n2353 vdd.n2352 185
R1151 vdd.n2354 vdd.n1138 185
R1152 vdd.n2356 vdd.n2355 185
R1153 vdd.n2358 vdd.n1136 185
R1154 vdd.n2360 vdd.n2359 185
R1155 vdd.n2361 vdd.n1131 185
R1156 vdd.n2363 vdd.n2362 185
R1157 vdd.n2365 vdd.n1129 185
R1158 vdd.n2367 vdd.n2366 185
R1159 vdd.n2368 vdd.n1127 185
R1160 vdd.n2370 vdd.n2369 185
R1161 vdd.n2373 vdd.n2372 185
R1162 vdd.n2375 vdd.n2374 185
R1163 vdd.n2377 vdd.n1125 185
R1164 vdd.n2379 vdd.n2378 185
R1165 vdd.n1437 vdd.n1124 185
R1166 vdd.n2266 vdd.n1435 185
R1167 vdd.n2266 vdd.n2265 185
R1168 vdd.n1445 vdd.n1434 185
R1169 vdd.n2256 vdd.n1434 185
R1170 vdd.n2255 vdd.n2254 185
R1171 vdd.n2257 vdd.n2255 185
R1172 vdd.n1444 vdd.n1443 185
R1173 vdd.n1443 vdd.n1442 185
R1174 vdd.n2248 vdd.n2247 185
R1175 vdd.n2247 vdd.n2246 185
R1176 vdd.n1448 vdd.n1447 185
R1177 vdd.n2237 vdd.n1448 185
R1178 vdd.n2236 vdd.n2235 185
R1179 vdd.n2238 vdd.n2236 185
R1180 vdd.n1455 vdd.n1454 185
R1181 vdd.n1460 vdd.n1454 185
R1182 vdd.n2231 vdd.n2230 185
R1183 vdd.n2230 vdd.n2229 185
R1184 vdd.n1458 vdd.n1457 185
R1185 vdd.n1459 vdd.n1458 185
R1186 vdd.n2220 vdd.n2219 185
R1187 vdd.n2221 vdd.n2220 185
R1188 vdd.n1468 vdd.n1467 185
R1189 vdd.n1467 vdd.n1466 185
R1190 vdd.n2215 vdd.n2214 185
R1191 vdd.n2214 vdd.n2213 185
R1192 vdd.n1471 vdd.n1470 185
R1193 vdd.n2204 vdd.n1471 185
R1194 vdd.n2203 vdd.n2202 185
R1195 vdd.n2205 vdd.n2203 185
R1196 vdd.n1478 vdd.n1477 185
R1197 vdd.n1482 vdd.n1477 185
R1198 vdd.n2198 vdd.n2197 185
R1199 vdd.n2197 vdd.n2196 185
R1200 vdd.n1481 vdd.n1480 185
R1201 vdd.n2187 vdd.n1481 185
R1202 vdd.n2186 vdd.n2185 185
R1203 vdd.n2188 vdd.n2186 185
R1204 vdd.n1490 vdd.n1489 185
R1205 vdd.n1489 vdd.n1488 185
R1206 vdd.n2181 vdd.n2180 185
R1207 vdd.n2180 vdd.n2179 185
R1208 vdd.n1493 vdd.n1492 185
R1209 vdd.n1494 vdd.n1493 185
R1210 vdd.n1863 vdd.n1862 185
R1211 vdd.n1864 vdd.n1863 185
R1212 vdd.n1501 vdd.n1500 185
R1213 vdd.n1505 vdd.n1500 185
R1214 vdd.n1858 vdd.n1857 185
R1215 vdd.n1857 vdd.n1856 185
R1216 vdd.n1504 vdd.n1503 185
R1217 vdd.n1847 vdd.n1504 185
R1218 vdd.n1846 vdd.n1845 185
R1219 vdd.n1848 vdd.n1846 185
R1220 vdd.n1512 vdd.n1511 185
R1221 vdd.n1517 vdd.n1511 185
R1222 vdd.n1841 vdd.n1840 185
R1223 vdd.n1840 vdd.n1839 185
R1224 vdd.n1515 vdd.n1514 185
R1225 vdd.n1516 vdd.n1515 185
R1226 vdd.n1830 vdd.n1829 185
R1227 vdd.n1831 vdd.n1830 185
R1228 vdd.n1525 vdd.n1524 185
R1229 vdd.n1524 vdd.n1523 185
R1230 vdd.n1825 vdd.n1824 185
R1231 vdd.n1824 vdd.n1823 185
R1232 vdd.n1528 vdd.n1527 185
R1233 vdd.n1814 vdd.n1528 185
R1234 vdd.n1813 vdd.n1812 185
R1235 vdd.n1815 vdd.n1813 185
R1236 vdd.n1535 vdd.n1534 185
R1237 vdd.n1539 vdd.n1534 185
R1238 vdd.n1808 vdd.n1807 185
R1239 vdd.n1807 vdd.n1806 185
R1240 vdd.n1538 vdd.n1537 185
R1241 vdd.n1797 vdd.n1538 185
R1242 vdd.n1796 vdd.n1795 185
R1243 vdd.n1798 vdd.n1796 185
R1244 vdd.n1547 vdd.n1546 185
R1245 vdd.n1546 vdd.n1545 185
R1246 vdd.n1791 vdd.n1790 185
R1247 vdd.n1790 vdd.n1789 185
R1248 vdd.n1550 vdd.n1549 185
R1249 vdd.n1587 vdd.n1550 185
R1250 vdd.n971 vdd.n969 185
R1251 vdd.n2593 vdd.n969 185
R1252 vdd.n2515 vdd.n989 185
R1253 vdd.n989 vdd.n976 185
R1254 vdd.n2517 vdd.n2516 185
R1255 vdd.n2518 vdd.n2517 185
R1256 vdd.n2514 vdd.n988 185
R1257 vdd.n1338 vdd.n988 185
R1258 vdd.n2513 vdd.n2512 185
R1259 vdd.n2512 vdd.n2511 185
R1260 vdd.n991 vdd.n990 185
R1261 vdd.n992 vdd.n991 185
R1262 vdd.n2502 vdd.n2501 185
R1263 vdd.n2503 vdd.n2502 185
R1264 vdd.n2500 vdd.n1002 185
R1265 vdd.n1002 vdd.n999 185
R1266 vdd.n2499 vdd.n2498 185
R1267 vdd.n2498 vdd.n2497 185
R1268 vdd.n1004 vdd.n1003 185
R1269 vdd.n1005 vdd.n1004 185
R1270 vdd.n2490 vdd.n2489 185
R1271 vdd.n2491 vdd.n2490 185
R1272 vdd.n2488 vdd.n1013 185
R1273 vdd.n1018 vdd.n1013 185
R1274 vdd.n2487 vdd.n2486 185
R1275 vdd.n2486 vdd.n2485 185
R1276 vdd.n1015 vdd.n1014 185
R1277 vdd.n1024 vdd.n1015 185
R1278 vdd.n2478 vdd.n2477 185
R1279 vdd.n2479 vdd.n2478 185
R1280 vdd.n2476 vdd.n1025 185
R1281 vdd.n1359 vdd.n1025 185
R1282 vdd.n2475 vdd.n2474 185
R1283 vdd.n2474 vdd.n2473 185
R1284 vdd.n1027 vdd.n1026 185
R1285 vdd.n1028 vdd.n1027 185
R1286 vdd.n2466 vdd.n2465 185
R1287 vdd.n2467 vdd.n2466 185
R1288 vdd.n2464 vdd.n1037 185
R1289 vdd.n1037 vdd.n1034 185
R1290 vdd.n2463 vdd.n2462 185
R1291 vdd.n2462 vdd.n2461 185
R1292 vdd.n1039 vdd.n1038 185
R1293 vdd.n1048 vdd.n1039 185
R1294 vdd.n2453 vdd.n2452 185
R1295 vdd.n2454 vdd.n2453 185
R1296 vdd.n2451 vdd.n1049 185
R1297 vdd.n1055 vdd.n1049 185
R1298 vdd.n2450 vdd.n2449 185
R1299 vdd.n2449 vdd.n2448 185
R1300 vdd.n1051 vdd.n1050 185
R1301 vdd.n1052 vdd.n1051 185
R1302 vdd.n2441 vdd.n2440 185
R1303 vdd.n2442 vdd.n2441 185
R1304 vdd.n2439 vdd.n1062 185
R1305 vdd.n1062 vdd.n1059 185
R1306 vdd.n2438 vdd.n2437 185
R1307 vdd.n2437 vdd.n2436 185
R1308 vdd.n1064 vdd.n1063 185
R1309 vdd.n1065 vdd.n1064 185
R1310 vdd.n2429 vdd.n2428 185
R1311 vdd.n2430 vdd.n2429 185
R1312 vdd.n2427 vdd.n1073 185
R1313 vdd.n1079 vdd.n1073 185
R1314 vdd.n2426 vdd.n2425 185
R1315 vdd.n2425 vdd.n2424 185
R1316 vdd.n1075 vdd.n1074 185
R1317 vdd.n1076 vdd.n1075 185
R1318 vdd.n2415 vdd.n2414 185
R1319 vdd.n2413 vdd.n1118 185
R1320 vdd.n2412 vdd.n1117 185
R1321 vdd.n2417 vdd.n1117 185
R1322 vdd.n2411 vdd.n2410 185
R1323 vdd.n2409 vdd.n2408 185
R1324 vdd.n2407 vdd.n2406 185
R1325 vdd.n2405 vdd.n2404 185
R1326 vdd.n2403 vdd.n2402 185
R1327 vdd.n2401 vdd.n2400 185
R1328 vdd.n2399 vdd.n2398 185
R1329 vdd.n2397 vdd.n2396 185
R1330 vdd.n2395 vdd.n2394 185
R1331 vdd.n2393 vdd.n2392 185
R1332 vdd.n2391 vdd.n2390 185
R1333 vdd.n2389 vdd.n2388 185
R1334 vdd.n2387 vdd.n2386 185
R1335 vdd.n2385 vdd.n2384 185
R1336 vdd.n2383 vdd.n2382 185
R1337 vdd.n1275 vdd.n1119 185
R1338 vdd.n1277 vdd.n1276 185
R1339 vdd.n1279 vdd.n1278 185
R1340 vdd.n1281 vdd.n1280 185
R1341 vdd.n1283 vdd.n1282 185
R1342 vdd.n1285 vdd.n1284 185
R1343 vdd.n1287 vdd.n1286 185
R1344 vdd.n1289 vdd.n1288 185
R1345 vdd.n1291 vdd.n1290 185
R1346 vdd.n1293 vdd.n1292 185
R1347 vdd.n1295 vdd.n1294 185
R1348 vdd.n1297 vdd.n1296 185
R1349 vdd.n1299 vdd.n1298 185
R1350 vdd.n1301 vdd.n1300 185
R1351 vdd.n1304 vdd.n1303 185
R1352 vdd.n1306 vdd.n1305 185
R1353 vdd.n1308 vdd.n1307 185
R1354 vdd.n2596 vdd.n2595 185
R1355 vdd.n2598 vdd.n2597 185
R1356 vdd.n2600 vdd.n2599 185
R1357 vdd.n2603 vdd.n2602 185
R1358 vdd.n2605 vdd.n2604 185
R1359 vdd.n2607 vdd.n2606 185
R1360 vdd.n2609 vdd.n2608 185
R1361 vdd.n2611 vdd.n2610 185
R1362 vdd.n2613 vdd.n2612 185
R1363 vdd.n2615 vdd.n2614 185
R1364 vdd.n2617 vdd.n2616 185
R1365 vdd.n2619 vdd.n2618 185
R1366 vdd.n2621 vdd.n2620 185
R1367 vdd.n2623 vdd.n2622 185
R1368 vdd.n2625 vdd.n2624 185
R1369 vdd.n2627 vdd.n2626 185
R1370 vdd.n2629 vdd.n2628 185
R1371 vdd.n2631 vdd.n2630 185
R1372 vdd.n2633 vdd.n2632 185
R1373 vdd.n2635 vdd.n2634 185
R1374 vdd.n2637 vdd.n2636 185
R1375 vdd.n2639 vdd.n2638 185
R1376 vdd.n2641 vdd.n2640 185
R1377 vdd.n2643 vdd.n2642 185
R1378 vdd.n2645 vdd.n2644 185
R1379 vdd.n2647 vdd.n2646 185
R1380 vdd.n2649 vdd.n2648 185
R1381 vdd.n2651 vdd.n2650 185
R1382 vdd.n2653 vdd.n2652 185
R1383 vdd.n2655 vdd.n2654 185
R1384 vdd.n2657 vdd.n2656 185
R1385 vdd.n2659 vdd.n2658 185
R1386 vdd.n2661 vdd.n2660 185
R1387 vdd.n2662 vdd.n970 185
R1388 vdd.n2664 vdd.n2663 185
R1389 vdd.n2665 vdd.n2664 185
R1390 vdd.n2594 vdd.n974 185
R1391 vdd.n2594 vdd.n2593 185
R1392 vdd.n1336 vdd.n975 185
R1393 vdd.n976 vdd.n975 185
R1394 vdd.n1337 vdd.n986 185
R1395 vdd.n2518 vdd.n986 185
R1396 vdd.n1340 vdd.n1339 185
R1397 vdd.n1339 vdd.n1338 185
R1398 vdd.n1341 vdd.n993 185
R1399 vdd.n2511 vdd.n993 185
R1400 vdd.n1343 vdd.n1342 185
R1401 vdd.n1342 vdd.n992 185
R1402 vdd.n1344 vdd.n1000 185
R1403 vdd.n2503 vdd.n1000 185
R1404 vdd.n1346 vdd.n1345 185
R1405 vdd.n1345 vdd.n999 185
R1406 vdd.n1347 vdd.n1006 185
R1407 vdd.n2497 vdd.n1006 185
R1408 vdd.n1349 vdd.n1348 185
R1409 vdd.n1348 vdd.n1005 185
R1410 vdd.n1350 vdd.n1011 185
R1411 vdd.n2491 vdd.n1011 185
R1412 vdd.n1352 vdd.n1351 185
R1413 vdd.n1351 vdd.n1018 185
R1414 vdd.n1353 vdd.n1016 185
R1415 vdd.n2485 vdd.n1016 185
R1416 vdd.n1355 vdd.n1354 185
R1417 vdd.n1354 vdd.n1024 185
R1418 vdd.n1356 vdd.n1022 185
R1419 vdd.n2479 vdd.n1022 185
R1420 vdd.n1358 vdd.n1357 185
R1421 vdd.n1359 vdd.n1358 185
R1422 vdd.n1335 vdd.n1029 185
R1423 vdd.n2473 vdd.n1029 185
R1424 vdd.n1334 vdd.n1333 185
R1425 vdd.n1333 vdd.n1028 185
R1426 vdd.n1332 vdd.n1035 185
R1427 vdd.n2467 vdd.n1035 185
R1428 vdd.n1331 vdd.n1330 185
R1429 vdd.n1330 vdd.n1034 185
R1430 vdd.n1329 vdd.n1040 185
R1431 vdd.n2461 vdd.n1040 185
R1432 vdd.n1328 vdd.n1327 185
R1433 vdd.n1327 vdd.n1048 185
R1434 vdd.n1326 vdd.n1046 185
R1435 vdd.n2454 vdd.n1046 185
R1436 vdd.n1325 vdd.n1324 185
R1437 vdd.n1324 vdd.n1055 185
R1438 vdd.n1323 vdd.n1053 185
R1439 vdd.n2448 vdd.n1053 185
R1440 vdd.n1322 vdd.n1321 185
R1441 vdd.n1321 vdd.n1052 185
R1442 vdd.n1320 vdd.n1060 185
R1443 vdd.n2442 vdd.n1060 185
R1444 vdd.n1319 vdd.n1318 185
R1445 vdd.n1318 vdd.n1059 185
R1446 vdd.n1317 vdd.n1066 185
R1447 vdd.n2436 vdd.n1066 185
R1448 vdd.n1316 vdd.n1315 185
R1449 vdd.n1315 vdd.n1065 185
R1450 vdd.n1314 vdd.n1071 185
R1451 vdd.n2430 vdd.n1071 185
R1452 vdd.n1313 vdd.n1312 185
R1453 vdd.n1312 vdd.n1079 185
R1454 vdd.n1311 vdd.n1077 185
R1455 vdd.n2424 vdd.n1077 185
R1456 vdd.n1310 vdd.n1309 185
R1457 vdd.n1309 vdd.n1076 185
R1458 vdd.n3449 vdd.n3448 185
R1459 vdd.n3448 vdd.n3447 185
R1460 vdd.n3450 vdd.n387 185
R1461 vdd.n387 vdd.n386 185
R1462 vdd.n3452 vdd.n3451 185
R1463 vdd.n3453 vdd.n3452 185
R1464 vdd.n382 vdd.n381 185
R1465 vdd.n3454 vdd.n382 185
R1466 vdd.n3457 vdd.n3456 185
R1467 vdd.n3456 vdd.n3455 185
R1468 vdd.n3458 vdd.n376 185
R1469 vdd.n376 vdd.n375 185
R1470 vdd.n3460 vdd.n3459 185
R1471 vdd.n3461 vdd.n3460 185
R1472 vdd.n371 vdd.n370 185
R1473 vdd.n3462 vdd.n371 185
R1474 vdd.n3465 vdd.n3464 185
R1475 vdd.n3464 vdd.n3463 185
R1476 vdd.n3466 vdd.n365 185
R1477 vdd.n3423 vdd.n365 185
R1478 vdd.n3468 vdd.n3467 185
R1479 vdd.n3469 vdd.n3468 185
R1480 vdd.n360 vdd.n359 185
R1481 vdd.n3470 vdd.n360 185
R1482 vdd.n3473 vdd.n3472 185
R1483 vdd.n3472 vdd.n3471 185
R1484 vdd.n3474 vdd.n354 185
R1485 vdd.n361 vdd.n354 185
R1486 vdd.n3476 vdd.n3475 185
R1487 vdd.n3477 vdd.n3476 185
R1488 vdd.n350 vdd.n349 185
R1489 vdd.n3478 vdd.n350 185
R1490 vdd.n3481 vdd.n3480 185
R1491 vdd.n3480 vdd.n3479 185
R1492 vdd.n3482 vdd.n345 185
R1493 vdd.n345 vdd.n344 185
R1494 vdd.n3484 vdd.n3483 185
R1495 vdd.n3485 vdd.n3484 185
R1496 vdd.n339 vdd.n337 185
R1497 vdd.n3486 vdd.n339 185
R1498 vdd.n3489 vdd.n3488 185
R1499 vdd.n3488 vdd.n3487 185
R1500 vdd.n338 vdd.n336 185
R1501 vdd.n340 vdd.n338 185
R1502 vdd.n3399 vdd.n3398 185
R1503 vdd.n3400 vdd.n3399 185
R1504 vdd.n635 vdd.n634 185
R1505 vdd.n634 vdd.n633 185
R1506 vdd.n3394 vdd.n3393 185
R1507 vdd.n3393 vdd.n3392 185
R1508 vdd.n638 vdd.n637 185
R1509 vdd.n644 vdd.n638 185
R1510 vdd.n3380 vdd.n3379 185
R1511 vdd.n3381 vdd.n3380 185
R1512 vdd.n646 vdd.n645 185
R1513 vdd.n3372 vdd.n645 185
R1514 vdd.n3375 vdd.n3374 185
R1515 vdd.n3374 vdd.n3373 185
R1516 vdd.n649 vdd.n648 185
R1517 vdd.n656 vdd.n649 185
R1518 vdd.n3363 vdd.n3362 185
R1519 vdd.n3364 vdd.n3363 185
R1520 vdd.n658 vdd.n657 185
R1521 vdd.n657 vdd.n655 185
R1522 vdd.n3358 vdd.n3357 185
R1523 vdd.n3357 vdd.n3356 185
R1524 vdd.n661 vdd.n660 185
R1525 vdd.n662 vdd.n661 185
R1526 vdd.n3347 vdd.n3346 185
R1527 vdd.n3348 vdd.n3347 185
R1528 vdd.n669 vdd.n668 185
R1529 vdd.n3339 vdd.n668 185
R1530 vdd.n3342 vdd.n3341 185
R1531 vdd.n3341 vdd.n3340 185
R1532 vdd.n672 vdd.n671 185
R1533 vdd.n679 vdd.n672 185
R1534 vdd.n3330 vdd.n3329 185
R1535 vdd.n3331 vdd.n3330 185
R1536 vdd.n681 vdd.n680 185
R1537 vdd.n680 vdd.n678 185
R1538 vdd.n3325 vdd.n3324 185
R1539 vdd.n3324 vdd.n3323 185
R1540 vdd.n684 vdd.n683 185
R1541 vdd.n723 vdd.n684 185
R1542 vdd.n3313 vdd.n3312 185
R1543 vdd.n3311 vdd.n725 185
R1544 vdd.n3310 vdd.n724 185
R1545 vdd.n3315 vdd.n724 185
R1546 vdd.n729 vdd.n728 185
R1547 vdd.n733 vdd.n732 185
R1548 vdd.n3306 vdd.n734 185
R1549 vdd.n3305 vdd.n3304 185
R1550 vdd.n3303 vdd.n3302 185
R1551 vdd.n3301 vdd.n3300 185
R1552 vdd.n3299 vdd.n3298 185
R1553 vdd.n3297 vdd.n3296 185
R1554 vdd.n3295 vdd.n3294 185
R1555 vdd.n3293 vdd.n3292 185
R1556 vdd.n3291 vdd.n3290 185
R1557 vdd.n3289 vdd.n3288 185
R1558 vdd.n3287 vdd.n3286 185
R1559 vdd.n3285 vdd.n3284 185
R1560 vdd.n3283 vdd.n3282 185
R1561 vdd.n3281 vdd.n3280 185
R1562 vdd.n3279 vdd.n3278 185
R1563 vdd.n3270 vdd.n747 185
R1564 vdd.n3272 vdd.n3271 185
R1565 vdd.n3269 vdd.n3268 185
R1566 vdd.n3267 vdd.n3266 185
R1567 vdd.n3265 vdd.n3264 185
R1568 vdd.n3263 vdd.n3262 185
R1569 vdd.n3261 vdd.n3260 185
R1570 vdd.n3259 vdd.n3258 185
R1571 vdd.n3257 vdd.n3256 185
R1572 vdd.n3255 vdd.n3254 185
R1573 vdd.n3253 vdd.n3252 185
R1574 vdd.n3251 vdd.n3250 185
R1575 vdd.n3249 vdd.n3248 185
R1576 vdd.n3247 vdd.n3246 185
R1577 vdd.n3245 vdd.n3244 185
R1578 vdd.n3243 vdd.n3242 185
R1579 vdd.n3241 vdd.n3240 185
R1580 vdd.n3239 vdd.n3238 185
R1581 vdd.n3237 vdd.n3236 185
R1582 vdd.n3235 vdd.n3234 185
R1583 vdd.n3233 vdd.n3232 185
R1584 vdd.n3231 vdd.n3230 185
R1585 vdd.n3224 vdd.n767 185
R1586 vdd.n3226 vdd.n3225 185
R1587 vdd.n3223 vdd.n3222 185
R1588 vdd.n3221 vdd.n3220 185
R1589 vdd.n3219 vdd.n3218 185
R1590 vdd.n3217 vdd.n3216 185
R1591 vdd.n3215 vdd.n3214 185
R1592 vdd.n3213 vdd.n3212 185
R1593 vdd.n3211 vdd.n3210 185
R1594 vdd.n3209 vdd.n3208 185
R1595 vdd.n3207 vdd.n3206 185
R1596 vdd.n3205 vdd.n3204 185
R1597 vdd.n3203 vdd.n3202 185
R1598 vdd.n3201 vdd.n3200 185
R1599 vdd.n3199 vdd.n3198 185
R1600 vdd.n3197 vdd.n3196 185
R1601 vdd.n3195 vdd.n3194 185
R1602 vdd.n3193 vdd.n3192 185
R1603 vdd.n3191 vdd.n3190 185
R1604 vdd.n3189 vdd.n3188 185
R1605 vdd.n3187 vdd.n691 185
R1606 vdd.n3317 vdd.n3316 185
R1607 vdd.n3316 vdd.n3315 185
R1608 vdd.n3444 vdd.n3443 185
R1609 vdd.n618 vdd.n425 185
R1610 vdd.n617 vdd.n616 185
R1611 vdd.n615 vdd.n614 185
R1612 vdd.n613 vdd.n430 185
R1613 vdd.n609 vdd.n608 185
R1614 vdd.n607 vdd.n606 185
R1615 vdd.n605 vdd.n604 185
R1616 vdd.n603 vdd.n432 185
R1617 vdd.n599 vdd.n598 185
R1618 vdd.n597 vdd.n596 185
R1619 vdd.n595 vdd.n594 185
R1620 vdd.n593 vdd.n434 185
R1621 vdd.n589 vdd.n588 185
R1622 vdd.n587 vdd.n586 185
R1623 vdd.n585 vdd.n584 185
R1624 vdd.n583 vdd.n436 185
R1625 vdd.n579 vdd.n578 185
R1626 vdd.n577 vdd.n576 185
R1627 vdd.n575 vdd.n574 185
R1628 vdd.n573 vdd.n438 185
R1629 vdd.n569 vdd.n568 185
R1630 vdd.n567 vdd.n566 185
R1631 vdd.n565 vdd.n564 185
R1632 vdd.n563 vdd.n442 185
R1633 vdd.n559 vdd.n558 185
R1634 vdd.n557 vdd.n556 185
R1635 vdd.n555 vdd.n554 185
R1636 vdd.n553 vdd.n444 185
R1637 vdd.n549 vdd.n548 185
R1638 vdd.n547 vdd.n546 185
R1639 vdd.n545 vdd.n544 185
R1640 vdd.n543 vdd.n446 185
R1641 vdd.n539 vdd.n538 185
R1642 vdd.n537 vdd.n536 185
R1643 vdd.n535 vdd.n534 185
R1644 vdd.n533 vdd.n448 185
R1645 vdd.n529 vdd.n528 185
R1646 vdd.n527 vdd.n526 185
R1647 vdd.n525 vdd.n524 185
R1648 vdd.n523 vdd.n450 185
R1649 vdd.n519 vdd.n518 185
R1650 vdd.n517 vdd.n516 185
R1651 vdd.n515 vdd.n514 185
R1652 vdd.n513 vdd.n454 185
R1653 vdd.n509 vdd.n508 185
R1654 vdd.n507 vdd.n506 185
R1655 vdd.n505 vdd.n504 185
R1656 vdd.n503 vdd.n456 185
R1657 vdd.n499 vdd.n498 185
R1658 vdd.n497 vdd.n496 185
R1659 vdd.n495 vdd.n494 185
R1660 vdd.n493 vdd.n458 185
R1661 vdd.n489 vdd.n488 185
R1662 vdd.n487 vdd.n486 185
R1663 vdd.n485 vdd.n484 185
R1664 vdd.n483 vdd.n460 185
R1665 vdd.n479 vdd.n478 185
R1666 vdd.n477 vdd.n476 185
R1667 vdd.n475 vdd.n474 185
R1668 vdd.n473 vdd.n462 185
R1669 vdd.n469 vdd.n468 185
R1670 vdd.n467 vdd.n466 185
R1671 vdd.n465 vdd.n392 185
R1672 vdd.n3440 vdd.n393 185
R1673 vdd.n3447 vdd.n393 185
R1674 vdd.n3439 vdd.n3438 185
R1675 vdd.n3438 vdd.n386 185
R1676 vdd.n3437 vdd.n385 185
R1677 vdd.n3453 vdd.n385 185
R1678 vdd.n621 vdd.n384 185
R1679 vdd.n3454 vdd.n384 185
R1680 vdd.n3433 vdd.n383 185
R1681 vdd.n3455 vdd.n383 185
R1682 vdd.n3432 vdd.n3431 185
R1683 vdd.n3431 vdd.n375 185
R1684 vdd.n3430 vdd.n374 185
R1685 vdd.n3461 vdd.n374 185
R1686 vdd.n623 vdd.n373 185
R1687 vdd.n3462 vdd.n373 185
R1688 vdd.n3426 vdd.n372 185
R1689 vdd.n3463 vdd.n372 185
R1690 vdd.n3425 vdd.n3424 185
R1691 vdd.n3424 vdd.n3423 185
R1692 vdd.n3422 vdd.n364 185
R1693 vdd.n3469 vdd.n364 185
R1694 vdd.n625 vdd.n363 185
R1695 vdd.n3470 vdd.n363 185
R1696 vdd.n3418 vdd.n362 185
R1697 vdd.n3471 vdd.n362 185
R1698 vdd.n3417 vdd.n3416 185
R1699 vdd.n3416 vdd.n361 185
R1700 vdd.n3415 vdd.n353 185
R1701 vdd.n3477 vdd.n353 185
R1702 vdd.n627 vdd.n352 185
R1703 vdd.n3478 vdd.n352 185
R1704 vdd.n3411 vdd.n351 185
R1705 vdd.n3479 vdd.n351 185
R1706 vdd.n3410 vdd.n3409 185
R1707 vdd.n3409 vdd.n344 185
R1708 vdd.n3408 vdd.n343 185
R1709 vdd.n3485 vdd.n343 185
R1710 vdd.n629 vdd.n342 185
R1711 vdd.n3486 vdd.n342 185
R1712 vdd.n3404 vdd.n341 185
R1713 vdd.n3487 vdd.n341 185
R1714 vdd.n3403 vdd.n3402 185
R1715 vdd.n3402 vdd.n340 185
R1716 vdd.n3401 vdd.n631 185
R1717 vdd.n3401 vdd.n3400 185
R1718 vdd.n3389 vdd.n632 185
R1719 vdd.n633 vdd.n632 185
R1720 vdd.n3391 vdd.n3390 185
R1721 vdd.n3392 vdd.n3391 185
R1722 vdd.n640 vdd.n639 185
R1723 vdd.n644 vdd.n639 185
R1724 vdd.n3383 vdd.n3382 185
R1725 vdd.n3382 vdd.n3381 185
R1726 vdd.n643 vdd.n642 185
R1727 vdd.n3372 vdd.n643 185
R1728 vdd.n3371 vdd.n3370 185
R1729 vdd.n3373 vdd.n3371 185
R1730 vdd.n651 vdd.n650 185
R1731 vdd.n656 vdd.n650 185
R1732 vdd.n3366 vdd.n3365 185
R1733 vdd.n3365 vdd.n3364 185
R1734 vdd.n654 vdd.n653 185
R1735 vdd.n655 vdd.n654 185
R1736 vdd.n3355 vdd.n3354 185
R1737 vdd.n3356 vdd.n3355 185
R1738 vdd.n664 vdd.n663 185
R1739 vdd.n663 vdd.n662 185
R1740 vdd.n3350 vdd.n3349 185
R1741 vdd.n3349 vdd.n3348 185
R1742 vdd.n667 vdd.n666 185
R1743 vdd.n3339 vdd.n667 185
R1744 vdd.n3338 vdd.n3337 185
R1745 vdd.n3340 vdd.n3338 185
R1746 vdd.n674 vdd.n673 185
R1747 vdd.n679 vdd.n673 185
R1748 vdd.n3333 vdd.n3332 185
R1749 vdd.n3332 vdd.n3331 185
R1750 vdd.n677 vdd.n676 185
R1751 vdd.n678 vdd.n677 185
R1752 vdd.n3322 vdd.n3321 185
R1753 vdd.n3323 vdd.n3322 185
R1754 vdd.n686 vdd.n685 185
R1755 vdd.n723 vdd.n685 185
R1756 vdd.n2936 vdd.n2935 185
R1757 vdd.n2934 vdd.n2700 185
R1758 vdd.n2933 vdd.n2699 185
R1759 vdd.n2938 vdd.n2699 185
R1760 vdd.n2932 vdd.n2931 185
R1761 vdd.n2930 vdd.n2929 185
R1762 vdd.n2928 vdd.n2927 185
R1763 vdd.n2926 vdd.n2925 185
R1764 vdd.n2924 vdd.n2923 185
R1765 vdd.n2922 vdd.n2921 185
R1766 vdd.n2920 vdd.n2919 185
R1767 vdd.n2918 vdd.n2917 185
R1768 vdd.n2916 vdd.n2915 185
R1769 vdd.n2914 vdd.n2913 185
R1770 vdd.n2912 vdd.n2911 185
R1771 vdd.n2910 vdd.n2909 185
R1772 vdd.n2908 vdd.n2907 185
R1773 vdd.n2906 vdd.n2905 185
R1774 vdd.n2904 vdd.n2903 185
R1775 vdd.n2902 vdd.n2901 185
R1776 vdd.n2900 vdd.n2899 185
R1777 vdd.n2898 vdd.n2897 185
R1778 vdd.n2896 vdd.n2895 185
R1779 vdd.n2894 vdd.n2893 185
R1780 vdd.n2892 vdd.n2891 185
R1781 vdd.n2890 vdd.n2889 185
R1782 vdd.n2888 vdd.n2887 185
R1783 vdd.n2886 vdd.n2885 185
R1784 vdd.n2884 vdd.n2883 185
R1785 vdd.n2882 vdd.n2881 185
R1786 vdd.n2880 vdd.n2879 185
R1787 vdd.n2878 vdd.n2877 185
R1788 vdd.n2876 vdd.n2875 185
R1789 vdd.n2873 vdd.n2872 185
R1790 vdd.n2871 vdd.n2870 185
R1791 vdd.n2869 vdd.n2868 185
R1792 vdd.n3087 vdd.n3086 185
R1793 vdd.n3089 vdd.n834 185
R1794 vdd.n3091 vdd.n3090 185
R1795 vdd.n3093 vdd.n831 185
R1796 vdd.n3095 vdd.n3094 185
R1797 vdd.n3097 vdd.n829 185
R1798 vdd.n3099 vdd.n3098 185
R1799 vdd.n3100 vdd.n828 185
R1800 vdd.n3102 vdd.n3101 185
R1801 vdd.n3104 vdd.n826 185
R1802 vdd.n3106 vdd.n3105 185
R1803 vdd.n3107 vdd.n825 185
R1804 vdd.n3109 vdd.n3108 185
R1805 vdd.n3111 vdd.n823 185
R1806 vdd.n3113 vdd.n3112 185
R1807 vdd.n3114 vdd.n822 185
R1808 vdd.n3116 vdd.n3115 185
R1809 vdd.n3118 vdd.n731 185
R1810 vdd.n3120 vdd.n3119 185
R1811 vdd.n3122 vdd.n820 185
R1812 vdd.n3124 vdd.n3123 185
R1813 vdd.n3125 vdd.n819 185
R1814 vdd.n3127 vdd.n3126 185
R1815 vdd.n3129 vdd.n817 185
R1816 vdd.n3131 vdd.n3130 185
R1817 vdd.n3132 vdd.n816 185
R1818 vdd.n3134 vdd.n3133 185
R1819 vdd.n3136 vdd.n814 185
R1820 vdd.n3138 vdd.n3137 185
R1821 vdd.n3139 vdd.n813 185
R1822 vdd.n3141 vdd.n3140 185
R1823 vdd.n3143 vdd.n812 185
R1824 vdd.n3144 vdd.n811 185
R1825 vdd.n3147 vdd.n3146 185
R1826 vdd.n3148 vdd.n809 185
R1827 vdd.n809 vdd.n692 185
R1828 vdd.n3085 vdd.n806 185
R1829 vdd.n3151 vdd.n806 185
R1830 vdd.n3084 vdd.n3083 185
R1831 vdd.n3083 vdd.n805 185
R1832 vdd.n3082 vdd.n836 185
R1833 vdd.n3082 vdd.n3081 185
R1834 vdd.n2816 vdd.n837 185
R1835 vdd.n846 vdd.n837 185
R1836 vdd.n2817 vdd.n844 185
R1837 vdd.n3075 vdd.n844 185
R1838 vdd.n2819 vdd.n2818 185
R1839 vdd.n2818 vdd.n843 185
R1840 vdd.n2820 vdd.n852 185
R1841 vdd.n3024 vdd.n852 185
R1842 vdd.n2822 vdd.n2821 185
R1843 vdd.n2821 vdd.n851 185
R1844 vdd.n2823 vdd.n858 185
R1845 vdd.n3018 vdd.n858 185
R1846 vdd.n2825 vdd.n2824 185
R1847 vdd.n2824 vdd.n857 185
R1848 vdd.n2826 vdd.n863 185
R1849 vdd.n3012 vdd.n863 185
R1850 vdd.n2828 vdd.n2827 185
R1851 vdd.n2827 vdd.n870 185
R1852 vdd.n2829 vdd.n868 185
R1853 vdd.n3006 vdd.n868 185
R1854 vdd.n2831 vdd.n2830 185
R1855 vdd.n2830 vdd.n878 185
R1856 vdd.n2832 vdd.n876 185
R1857 vdd.n2999 vdd.n876 185
R1858 vdd.n2834 vdd.n2833 185
R1859 vdd.n2833 vdd.n875 185
R1860 vdd.n2835 vdd.n883 185
R1861 vdd.n2993 vdd.n883 185
R1862 vdd.n2837 vdd.n2836 185
R1863 vdd.n2836 vdd.n882 185
R1864 vdd.n2838 vdd.n888 185
R1865 vdd.n2987 vdd.n888 185
R1866 vdd.n2840 vdd.n2839 185
R1867 vdd.n2839 vdd.n895 185
R1868 vdd.n2841 vdd.n893 185
R1869 vdd.n2981 vdd.n893 185
R1870 vdd.n2843 vdd.n2842 185
R1871 vdd.n2842 vdd.n901 185
R1872 vdd.n2844 vdd.n899 185
R1873 vdd.n2975 vdd.n899 185
R1874 vdd.n2846 vdd.n2845 185
R1875 vdd.n2847 vdd.n2846 185
R1876 vdd.n2815 vdd.n906 185
R1877 vdd.n2969 vdd.n906 185
R1878 vdd.n2814 vdd.n2813 185
R1879 vdd.n2813 vdd.n905 185
R1880 vdd.n2812 vdd.n912 185
R1881 vdd.n2963 vdd.n912 185
R1882 vdd.n2811 vdd.n2810 185
R1883 vdd.n2810 vdd.n911 185
R1884 vdd.n2809 vdd.n918 185
R1885 vdd.n2957 vdd.n918 185
R1886 vdd.n2808 vdd.n2807 185
R1887 vdd.n2807 vdd.n917 185
R1888 vdd.n2703 vdd.n923 185
R1889 vdd.n2951 vdd.n923 185
R1890 vdd.n2864 vdd.n2863 185
R1891 vdd.n2863 vdd.n2862 185
R1892 vdd.n2865 vdd.n929 185
R1893 vdd.n2945 vdd.n929 185
R1894 vdd.n2867 vdd.n2866 185
R1895 vdd.n2867 vdd.n928 185
R1896 vdd.n927 vdd.n926 185
R1897 vdd.n928 vdd.n927 185
R1898 vdd.n2947 vdd.n2946 185
R1899 vdd.n2946 vdd.n2945 185
R1900 vdd.n2948 vdd.n925 185
R1901 vdd.n2862 vdd.n925 185
R1902 vdd.n2950 vdd.n2949 185
R1903 vdd.n2951 vdd.n2950 185
R1904 vdd.n916 vdd.n915 185
R1905 vdd.n917 vdd.n916 185
R1906 vdd.n2959 vdd.n2958 185
R1907 vdd.n2958 vdd.n2957 185
R1908 vdd.n2960 vdd.n914 185
R1909 vdd.n914 vdd.n911 185
R1910 vdd.n2962 vdd.n2961 185
R1911 vdd.n2963 vdd.n2962 185
R1912 vdd.n904 vdd.n903 185
R1913 vdd.n905 vdd.n904 185
R1914 vdd.n2971 vdd.n2970 185
R1915 vdd.n2970 vdd.n2969 185
R1916 vdd.n2972 vdd.n902 185
R1917 vdd.n2847 vdd.n902 185
R1918 vdd.n2974 vdd.n2973 185
R1919 vdd.n2975 vdd.n2974 185
R1920 vdd.n892 vdd.n891 185
R1921 vdd.n901 vdd.n892 185
R1922 vdd.n2983 vdd.n2982 185
R1923 vdd.n2982 vdd.n2981 185
R1924 vdd.n2984 vdd.n890 185
R1925 vdd.n895 vdd.n890 185
R1926 vdd.n2986 vdd.n2985 185
R1927 vdd.n2987 vdd.n2986 185
R1928 vdd.n881 vdd.n880 185
R1929 vdd.n882 vdd.n881 185
R1930 vdd.n2995 vdd.n2994 185
R1931 vdd.n2994 vdd.n2993 185
R1932 vdd.n2996 vdd.n879 185
R1933 vdd.n879 vdd.n875 185
R1934 vdd.n2998 vdd.n2997 185
R1935 vdd.n2999 vdd.n2998 185
R1936 vdd.n867 vdd.n866 185
R1937 vdd.n878 vdd.n867 185
R1938 vdd.n3008 vdd.n3007 185
R1939 vdd.n3007 vdd.n3006 185
R1940 vdd.n3009 vdd.n865 185
R1941 vdd.n870 vdd.n865 185
R1942 vdd.n3011 vdd.n3010 185
R1943 vdd.n3012 vdd.n3011 185
R1944 vdd.n856 vdd.n855 185
R1945 vdd.n857 vdd.n856 185
R1946 vdd.n3020 vdd.n3019 185
R1947 vdd.n3019 vdd.n3018 185
R1948 vdd.n3021 vdd.n854 185
R1949 vdd.n854 vdd.n851 185
R1950 vdd.n3023 vdd.n3022 185
R1951 vdd.n3024 vdd.n3023 185
R1952 vdd.n842 vdd.n841 185
R1953 vdd.n843 vdd.n842 185
R1954 vdd.n3077 vdd.n3076 185
R1955 vdd.n3076 vdd.n3075 185
R1956 vdd.n3078 vdd.n840 185
R1957 vdd.n846 vdd.n840 185
R1958 vdd.n3080 vdd.n3079 185
R1959 vdd.n3081 vdd.n3080 185
R1960 vdd.n810 vdd.n808 185
R1961 vdd.n808 vdd.n805 185
R1962 vdd.n3150 vdd.n3149 185
R1963 vdd.n3151 vdd.n3150 185
R1964 vdd.n2592 vdd.n2591 185
R1965 vdd.n2593 vdd.n2592 185
R1966 vdd.n980 vdd.n978 185
R1967 vdd.n978 vdd.n976 185
R1968 vdd.n2507 vdd.n987 185
R1969 vdd.n2518 vdd.n987 185
R1970 vdd.n2508 vdd.n996 185
R1971 vdd.n1338 vdd.n996 185
R1972 vdd.n2510 vdd.n2509 185
R1973 vdd.n2511 vdd.n2510 185
R1974 vdd.n2506 vdd.n995 185
R1975 vdd.n995 vdd.n992 185
R1976 vdd.n2505 vdd.n2504 185
R1977 vdd.n2504 vdd.n2503 185
R1978 vdd.n998 vdd.n997 185
R1979 vdd.n999 vdd.n998 185
R1980 vdd.n2496 vdd.n2495 185
R1981 vdd.n2497 vdd.n2496 185
R1982 vdd.n2494 vdd.n1008 185
R1983 vdd.n1008 vdd.n1005 185
R1984 vdd.n2493 vdd.n2492 185
R1985 vdd.n2492 vdd.n2491 185
R1986 vdd.n1010 vdd.n1009 185
R1987 vdd.n1018 vdd.n1010 185
R1988 vdd.n2484 vdd.n2483 185
R1989 vdd.n2485 vdd.n2484 185
R1990 vdd.n2482 vdd.n1019 185
R1991 vdd.n1024 vdd.n1019 185
R1992 vdd.n2481 vdd.n2480 185
R1993 vdd.n2480 vdd.n2479 185
R1994 vdd.n1021 vdd.n1020 185
R1995 vdd.n1359 vdd.n1021 185
R1996 vdd.n2472 vdd.n2471 185
R1997 vdd.n2473 vdd.n2472 185
R1998 vdd.n2470 vdd.n1031 185
R1999 vdd.n1031 vdd.n1028 185
R2000 vdd.n2469 vdd.n2468 185
R2001 vdd.n2468 vdd.n2467 185
R2002 vdd.n1033 vdd.n1032 185
R2003 vdd.n1034 vdd.n1033 185
R2004 vdd.n2460 vdd.n2459 185
R2005 vdd.n2461 vdd.n2460 185
R2006 vdd.n2457 vdd.n1042 185
R2007 vdd.n1048 vdd.n1042 185
R2008 vdd.n2456 vdd.n2455 185
R2009 vdd.n2455 vdd.n2454 185
R2010 vdd.n1045 vdd.n1044 185
R2011 vdd.n1055 vdd.n1045 185
R2012 vdd.n2447 vdd.n2446 185
R2013 vdd.n2448 vdd.n2447 185
R2014 vdd.n2445 vdd.n1056 185
R2015 vdd.n1056 vdd.n1052 185
R2016 vdd.n2444 vdd.n2443 185
R2017 vdd.n2443 vdd.n2442 185
R2018 vdd.n1058 vdd.n1057 185
R2019 vdd.n1059 vdd.n1058 185
R2020 vdd.n2435 vdd.n2434 185
R2021 vdd.n2436 vdd.n2435 185
R2022 vdd.n2433 vdd.n1068 185
R2023 vdd.n1068 vdd.n1065 185
R2024 vdd.n2432 vdd.n2431 185
R2025 vdd.n2431 vdd.n2430 185
R2026 vdd.n1070 vdd.n1069 185
R2027 vdd.n1079 vdd.n1070 185
R2028 vdd.n2423 vdd.n2422 185
R2029 vdd.n2424 vdd.n2423 185
R2030 vdd.n2421 vdd.n1080 185
R2031 vdd.n1080 vdd.n1076 185
R2032 vdd.n2523 vdd.n951 185
R2033 vdd.n2665 vdd.n951 185
R2034 vdd.n2525 vdd.n2524 185
R2035 vdd.n2527 vdd.n2526 185
R2036 vdd.n2529 vdd.n2528 185
R2037 vdd.n2531 vdd.n2530 185
R2038 vdd.n2533 vdd.n2532 185
R2039 vdd.n2535 vdd.n2534 185
R2040 vdd.n2537 vdd.n2536 185
R2041 vdd.n2539 vdd.n2538 185
R2042 vdd.n2541 vdd.n2540 185
R2043 vdd.n2543 vdd.n2542 185
R2044 vdd.n2545 vdd.n2544 185
R2045 vdd.n2547 vdd.n2546 185
R2046 vdd.n2549 vdd.n2548 185
R2047 vdd.n2551 vdd.n2550 185
R2048 vdd.n2553 vdd.n2552 185
R2049 vdd.n2555 vdd.n2554 185
R2050 vdd.n2557 vdd.n2556 185
R2051 vdd.n2559 vdd.n2558 185
R2052 vdd.n2561 vdd.n2560 185
R2053 vdd.n2563 vdd.n2562 185
R2054 vdd.n2565 vdd.n2564 185
R2055 vdd.n2567 vdd.n2566 185
R2056 vdd.n2569 vdd.n2568 185
R2057 vdd.n2571 vdd.n2570 185
R2058 vdd.n2573 vdd.n2572 185
R2059 vdd.n2575 vdd.n2574 185
R2060 vdd.n2577 vdd.n2576 185
R2061 vdd.n2579 vdd.n2578 185
R2062 vdd.n2581 vdd.n2580 185
R2063 vdd.n2583 vdd.n2582 185
R2064 vdd.n2585 vdd.n2584 185
R2065 vdd.n2587 vdd.n2586 185
R2066 vdd.n2589 vdd.n2588 185
R2067 vdd.n2590 vdd.n979 185
R2068 vdd.n2522 vdd.n977 185
R2069 vdd.n2593 vdd.n977 185
R2070 vdd.n2521 vdd.n2520 185
R2071 vdd.n2520 vdd.n976 185
R2072 vdd.n2519 vdd.n984 185
R2073 vdd.n2519 vdd.n2518 185
R2074 vdd.n1256 vdd.n985 185
R2075 vdd.n1338 vdd.n985 185
R2076 vdd.n1257 vdd.n994 185
R2077 vdd.n2511 vdd.n994 185
R2078 vdd.n1259 vdd.n1258 185
R2079 vdd.n1258 vdd.n992 185
R2080 vdd.n1260 vdd.n1001 185
R2081 vdd.n2503 vdd.n1001 185
R2082 vdd.n1262 vdd.n1261 185
R2083 vdd.n1261 vdd.n999 185
R2084 vdd.n1263 vdd.n1007 185
R2085 vdd.n2497 vdd.n1007 185
R2086 vdd.n1265 vdd.n1264 185
R2087 vdd.n1264 vdd.n1005 185
R2088 vdd.n1266 vdd.n1012 185
R2089 vdd.n2491 vdd.n1012 185
R2090 vdd.n1268 vdd.n1267 185
R2091 vdd.n1267 vdd.n1018 185
R2092 vdd.n1269 vdd.n1017 185
R2093 vdd.n2485 vdd.n1017 185
R2094 vdd.n1271 vdd.n1270 185
R2095 vdd.n1270 vdd.n1024 185
R2096 vdd.n1272 vdd.n1023 185
R2097 vdd.n2479 vdd.n1023 185
R2098 vdd.n1361 vdd.n1360 185
R2099 vdd.n1360 vdd.n1359 185
R2100 vdd.n1362 vdd.n1030 185
R2101 vdd.n2473 vdd.n1030 185
R2102 vdd.n1364 vdd.n1363 185
R2103 vdd.n1363 vdd.n1028 185
R2104 vdd.n1365 vdd.n1036 185
R2105 vdd.n2467 vdd.n1036 185
R2106 vdd.n1367 vdd.n1366 185
R2107 vdd.n1366 vdd.n1034 185
R2108 vdd.n1368 vdd.n1041 185
R2109 vdd.n2461 vdd.n1041 185
R2110 vdd.n1370 vdd.n1369 185
R2111 vdd.n1369 vdd.n1048 185
R2112 vdd.n1371 vdd.n1047 185
R2113 vdd.n2454 vdd.n1047 185
R2114 vdd.n1373 vdd.n1372 185
R2115 vdd.n1372 vdd.n1055 185
R2116 vdd.n1374 vdd.n1054 185
R2117 vdd.n2448 vdd.n1054 185
R2118 vdd.n1376 vdd.n1375 185
R2119 vdd.n1375 vdd.n1052 185
R2120 vdd.n1377 vdd.n1061 185
R2121 vdd.n2442 vdd.n1061 185
R2122 vdd.n1379 vdd.n1378 185
R2123 vdd.n1378 vdd.n1059 185
R2124 vdd.n1380 vdd.n1067 185
R2125 vdd.n2436 vdd.n1067 185
R2126 vdd.n1382 vdd.n1381 185
R2127 vdd.n1381 vdd.n1065 185
R2128 vdd.n1383 vdd.n1072 185
R2129 vdd.n2430 vdd.n1072 185
R2130 vdd.n1385 vdd.n1384 185
R2131 vdd.n1384 vdd.n1079 185
R2132 vdd.n1386 vdd.n1078 185
R2133 vdd.n2424 vdd.n1078 185
R2134 vdd.n1388 vdd.n1387 185
R2135 vdd.n1387 vdd.n1076 185
R2136 vdd.n2420 vdd.n2419 185
R2137 vdd.n1082 vdd.n1081 185
R2138 vdd.n1223 vdd.n1222 185
R2139 vdd.n1225 vdd.n1224 185
R2140 vdd.n1227 vdd.n1226 185
R2141 vdd.n1229 vdd.n1228 185
R2142 vdd.n1231 vdd.n1230 185
R2143 vdd.n1233 vdd.n1232 185
R2144 vdd.n1235 vdd.n1234 185
R2145 vdd.n1237 vdd.n1236 185
R2146 vdd.n1239 vdd.n1238 185
R2147 vdd.n1241 vdd.n1240 185
R2148 vdd.n1243 vdd.n1242 185
R2149 vdd.n1245 vdd.n1244 185
R2150 vdd.n1247 vdd.n1246 185
R2151 vdd.n1249 vdd.n1248 185
R2152 vdd.n1251 vdd.n1250 185
R2153 vdd.n1422 vdd.n1252 185
R2154 vdd.n1421 vdd.n1420 185
R2155 vdd.n1419 vdd.n1418 185
R2156 vdd.n1417 vdd.n1416 185
R2157 vdd.n1415 vdd.n1414 185
R2158 vdd.n1413 vdd.n1412 185
R2159 vdd.n1411 vdd.n1410 185
R2160 vdd.n1409 vdd.n1408 185
R2161 vdd.n1407 vdd.n1406 185
R2162 vdd.n1405 vdd.n1404 185
R2163 vdd.n1403 vdd.n1402 185
R2164 vdd.n1401 vdd.n1400 185
R2165 vdd.n1399 vdd.n1398 185
R2166 vdd.n1397 vdd.n1396 185
R2167 vdd.n1395 vdd.n1394 185
R2168 vdd.n1393 vdd.n1392 185
R2169 vdd.n1391 vdd.n1390 185
R2170 vdd.n1389 vdd.n1116 185
R2171 vdd.n2417 vdd.n1116 185
R2172 vdd.n2417 vdd.n1083 179.345
R2173 vdd.n3315 vdd.n692 179.345
R2174 vdd.n327 vdd.n326 171.744
R2175 vdd.n326 vdd.n325 171.744
R2176 vdd.n325 vdd.n294 171.744
R2177 vdd.n318 vdd.n294 171.744
R2178 vdd.n318 vdd.n317 171.744
R2179 vdd.n317 vdd.n299 171.744
R2180 vdd.n310 vdd.n299 171.744
R2181 vdd.n310 vdd.n309 171.744
R2182 vdd.n309 vdd.n303 171.744
R2183 vdd.n268 vdd.n267 171.744
R2184 vdd.n267 vdd.n266 171.744
R2185 vdd.n266 vdd.n235 171.744
R2186 vdd.n259 vdd.n235 171.744
R2187 vdd.n259 vdd.n258 171.744
R2188 vdd.n258 vdd.n240 171.744
R2189 vdd.n251 vdd.n240 171.744
R2190 vdd.n251 vdd.n250 171.744
R2191 vdd.n250 vdd.n244 171.744
R2192 vdd.n225 vdd.n224 171.744
R2193 vdd.n224 vdd.n223 171.744
R2194 vdd.n223 vdd.n192 171.744
R2195 vdd.n216 vdd.n192 171.744
R2196 vdd.n216 vdd.n215 171.744
R2197 vdd.n215 vdd.n197 171.744
R2198 vdd.n208 vdd.n197 171.744
R2199 vdd.n208 vdd.n207 171.744
R2200 vdd.n207 vdd.n201 171.744
R2201 vdd.n166 vdd.n165 171.744
R2202 vdd.n165 vdd.n164 171.744
R2203 vdd.n164 vdd.n133 171.744
R2204 vdd.n157 vdd.n133 171.744
R2205 vdd.n157 vdd.n156 171.744
R2206 vdd.n156 vdd.n138 171.744
R2207 vdd.n149 vdd.n138 171.744
R2208 vdd.n149 vdd.n148 171.744
R2209 vdd.n148 vdd.n142 171.744
R2210 vdd.n124 vdd.n123 171.744
R2211 vdd.n123 vdd.n122 171.744
R2212 vdd.n122 vdd.n91 171.744
R2213 vdd.n115 vdd.n91 171.744
R2214 vdd.n115 vdd.n114 171.744
R2215 vdd.n114 vdd.n96 171.744
R2216 vdd.n107 vdd.n96 171.744
R2217 vdd.n107 vdd.n106 171.744
R2218 vdd.n106 vdd.n100 171.744
R2219 vdd.n65 vdd.n64 171.744
R2220 vdd.n64 vdd.n63 171.744
R2221 vdd.n63 vdd.n32 171.744
R2222 vdd.n56 vdd.n32 171.744
R2223 vdd.n56 vdd.n55 171.744
R2224 vdd.n55 vdd.n37 171.744
R2225 vdd.n48 vdd.n37 171.744
R2226 vdd.n48 vdd.n47 171.744
R2227 vdd.n47 vdd.n41 171.744
R2228 vdd.n2108 vdd.n2107 171.744
R2229 vdd.n2107 vdd.n2106 171.744
R2230 vdd.n2106 vdd.n2075 171.744
R2231 vdd.n2099 vdd.n2075 171.744
R2232 vdd.n2099 vdd.n2098 171.744
R2233 vdd.n2098 vdd.n2080 171.744
R2234 vdd.n2091 vdd.n2080 171.744
R2235 vdd.n2091 vdd.n2090 171.744
R2236 vdd.n2090 vdd.n2084 171.744
R2237 vdd.n2167 vdd.n2166 171.744
R2238 vdd.n2166 vdd.n2165 171.744
R2239 vdd.n2165 vdd.n2134 171.744
R2240 vdd.n2158 vdd.n2134 171.744
R2241 vdd.n2158 vdd.n2157 171.744
R2242 vdd.n2157 vdd.n2139 171.744
R2243 vdd.n2150 vdd.n2139 171.744
R2244 vdd.n2150 vdd.n2149 171.744
R2245 vdd.n2149 vdd.n2143 171.744
R2246 vdd.n2006 vdd.n2005 171.744
R2247 vdd.n2005 vdd.n2004 171.744
R2248 vdd.n2004 vdd.n1973 171.744
R2249 vdd.n1997 vdd.n1973 171.744
R2250 vdd.n1997 vdd.n1996 171.744
R2251 vdd.n1996 vdd.n1978 171.744
R2252 vdd.n1989 vdd.n1978 171.744
R2253 vdd.n1989 vdd.n1988 171.744
R2254 vdd.n1988 vdd.n1982 171.744
R2255 vdd.n2065 vdd.n2064 171.744
R2256 vdd.n2064 vdd.n2063 171.744
R2257 vdd.n2063 vdd.n2032 171.744
R2258 vdd.n2056 vdd.n2032 171.744
R2259 vdd.n2056 vdd.n2055 171.744
R2260 vdd.n2055 vdd.n2037 171.744
R2261 vdd.n2048 vdd.n2037 171.744
R2262 vdd.n2048 vdd.n2047 171.744
R2263 vdd.n2047 vdd.n2041 171.744
R2264 vdd.n1905 vdd.n1904 171.744
R2265 vdd.n1904 vdd.n1903 171.744
R2266 vdd.n1903 vdd.n1872 171.744
R2267 vdd.n1896 vdd.n1872 171.744
R2268 vdd.n1896 vdd.n1895 171.744
R2269 vdd.n1895 vdd.n1877 171.744
R2270 vdd.n1888 vdd.n1877 171.744
R2271 vdd.n1888 vdd.n1887 171.744
R2272 vdd.n1887 vdd.n1881 171.744
R2273 vdd.n1964 vdd.n1963 171.744
R2274 vdd.n1963 vdd.n1962 171.744
R2275 vdd.n1962 vdd.n1931 171.744
R2276 vdd.n1955 vdd.n1931 171.744
R2277 vdd.n1955 vdd.n1954 171.744
R2278 vdd.n1954 vdd.n1936 171.744
R2279 vdd.n1947 vdd.n1936 171.744
R2280 vdd.n1947 vdd.n1946 171.744
R2281 vdd.n1946 vdd.n1940 171.744
R2282 vdd.n468 vdd.n467 146.341
R2283 vdd.n474 vdd.n473 146.341
R2284 vdd.n478 vdd.n477 146.341
R2285 vdd.n484 vdd.n483 146.341
R2286 vdd.n488 vdd.n487 146.341
R2287 vdd.n494 vdd.n493 146.341
R2288 vdd.n498 vdd.n497 146.341
R2289 vdd.n504 vdd.n503 146.341
R2290 vdd.n508 vdd.n507 146.341
R2291 vdd.n514 vdd.n513 146.341
R2292 vdd.n518 vdd.n517 146.341
R2293 vdd.n524 vdd.n523 146.341
R2294 vdd.n528 vdd.n527 146.341
R2295 vdd.n534 vdd.n533 146.341
R2296 vdd.n538 vdd.n537 146.341
R2297 vdd.n544 vdd.n543 146.341
R2298 vdd.n548 vdd.n547 146.341
R2299 vdd.n554 vdd.n553 146.341
R2300 vdd.n558 vdd.n557 146.341
R2301 vdd.n564 vdd.n563 146.341
R2302 vdd.n568 vdd.n567 146.341
R2303 vdd.n574 vdd.n573 146.341
R2304 vdd.n578 vdd.n577 146.341
R2305 vdd.n584 vdd.n583 146.341
R2306 vdd.n588 vdd.n587 146.341
R2307 vdd.n594 vdd.n593 146.341
R2308 vdd.n598 vdd.n597 146.341
R2309 vdd.n604 vdd.n603 146.341
R2310 vdd.n608 vdd.n607 146.341
R2311 vdd.n614 vdd.n613 146.341
R2312 vdd.n616 vdd.n425 146.341
R2313 vdd.n3322 vdd.n685 146.341
R2314 vdd.n3322 vdd.n677 146.341
R2315 vdd.n3332 vdd.n677 146.341
R2316 vdd.n3332 vdd.n673 146.341
R2317 vdd.n3338 vdd.n673 146.341
R2318 vdd.n3338 vdd.n667 146.341
R2319 vdd.n3349 vdd.n667 146.341
R2320 vdd.n3349 vdd.n663 146.341
R2321 vdd.n3355 vdd.n663 146.341
R2322 vdd.n3355 vdd.n654 146.341
R2323 vdd.n3365 vdd.n654 146.341
R2324 vdd.n3365 vdd.n650 146.341
R2325 vdd.n3371 vdd.n650 146.341
R2326 vdd.n3371 vdd.n643 146.341
R2327 vdd.n3382 vdd.n643 146.341
R2328 vdd.n3382 vdd.n639 146.341
R2329 vdd.n3391 vdd.n639 146.341
R2330 vdd.n3391 vdd.n632 146.341
R2331 vdd.n3401 vdd.n632 146.341
R2332 vdd.n3402 vdd.n3401 146.341
R2333 vdd.n3402 vdd.n341 146.341
R2334 vdd.n342 vdd.n341 146.341
R2335 vdd.n343 vdd.n342 146.341
R2336 vdd.n3409 vdd.n343 146.341
R2337 vdd.n3409 vdd.n351 146.341
R2338 vdd.n352 vdd.n351 146.341
R2339 vdd.n353 vdd.n352 146.341
R2340 vdd.n3416 vdd.n353 146.341
R2341 vdd.n3416 vdd.n362 146.341
R2342 vdd.n363 vdd.n362 146.341
R2343 vdd.n364 vdd.n363 146.341
R2344 vdd.n3424 vdd.n364 146.341
R2345 vdd.n3424 vdd.n372 146.341
R2346 vdd.n373 vdd.n372 146.341
R2347 vdd.n374 vdd.n373 146.341
R2348 vdd.n3431 vdd.n374 146.341
R2349 vdd.n3431 vdd.n383 146.341
R2350 vdd.n384 vdd.n383 146.341
R2351 vdd.n385 vdd.n384 146.341
R2352 vdd.n3438 vdd.n385 146.341
R2353 vdd.n3438 vdd.n393 146.341
R2354 vdd.n725 vdd.n724 146.341
R2355 vdd.n728 vdd.n724 146.341
R2356 vdd.n734 vdd.n733 146.341
R2357 vdd.n3304 vdd.n3303 146.341
R2358 vdd.n3300 vdd.n3299 146.341
R2359 vdd.n3296 vdd.n3295 146.341
R2360 vdd.n3292 vdd.n3291 146.341
R2361 vdd.n3288 vdd.n3287 146.341
R2362 vdd.n3284 vdd.n3283 146.341
R2363 vdd.n3280 vdd.n3279 146.341
R2364 vdd.n3271 vdd.n3270 146.341
R2365 vdd.n3268 vdd.n3267 146.341
R2366 vdd.n3264 vdd.n3263 146.341
R2367 vdd.n3260 vdd.n3259 146.341
R2368 vdd.n3256 vdd.n3255 146.341
R2369 vdd.n3252 vdd.n3251 146.341
R2370 vdd.n3248 vdd.n3247 146.341
R2371 vdd.n3244 vdd.n3243 146.341
R2372 vdd.n3240 vdd.n3239 146.341
R2373 vdd.n3236 vdd.n3235 146.341
R2374 vdd.n3232 vdd.n3231 146.341
R2375 vdd.n3225 vdd.n3224 146.341
R2376 vdd.n3222 vdd.n3221 146.341
R2377 vdd.n3218 vdd.n3217 146.341
R2378 vdd.n3214 vdd.n3213 146.341
R2379 vdd.n3210 vdd.n3209 146.341
R2380 vdd.n3206 vdd.n3205 146.341
R2381 vdd.n3202 vdd.n3201 146.341
R2382 vdd.n3198 vdd.n3197 146.341
R2383 vdd.n3194 vdd.n3193 146.341
R2384 vdd.n3190 vdd.n3189 146.341
R2385 vdd.n3316 vdd.n691 146.341
R2386 vdd.n3324 vdd.n684 146.341
R2387 vdd.n3324 vdd.n680 146.341
R2388 vdd.n3330 vdd.n680 146.341
R2389 vdd.n3330 vdd.n672 146.341
R2390 vdd.n3341 vdd.n672 146.341
R2391 vdd.n3341 vdd.n668 146.341
R2392 vdd.n3347 vdd.n668 146.341
R2393 vdd.n3347 vdd.n661 146.341
R2394 vdd.n3357 vdd.n661 146.341
R2395 vdd.n3357 vdd.n657 146.341
R2396 vdd.n3363 vdd.n657 146.341
R2397 vdd.n3363 vdd.n649 146.341
R2398 vdd.n3374 vdd.n649 146.341
R2399 vdd.n3374 vdd.n645 146.341
R2400 vdd.n3380 vdd.n645 146.341
R2401 vdd.n3380 vdd.n638 146.341
R2402 vdd.n3393 vdd.n638 146.341
R2403 vdd.n3393 vdd.n634 146.341
R2404 vdd.n3399 vdd.n634 146.341
R2405 vdd.n3399 vdd.n338 146.341
R2406 vdd.n3488 vdd.n338 146.341
R2407 vdd.n3488 vdd.n339 146.341
R2408 vdd.n3484 vdd.n339 146.341
R2409 vdd.n3484 vdd.n345 146.341
R2410 vdd.n3480 vdd.n345 146.341
R2411 vdd.n3480 vdd.n350 146.341
R2412 vdd.n3476 vdd.n350 146.341
R2413 vdd.n3476 vdd.n354 146.341
R2414 vdd.n3472 vdd.n354 146.341
R2415 vdd.n3472 vdd.n360 146.341
R2416 vdd.n3468 vdd.n360 146.341
R2417 vdd.n3468 vdd.n365 146.341
R2418 vdd.n3464 vdd.n365 146.341
R2419 vdd.n3464 vdd.n371 146.341
R2420 vdd.n3460 vdd.n371 146.341
R2421 vdd.n3460 vdd.n376 146.341
R2422 vdd.n3456 vdd.n376 146.341
R2423 vdd.n3456 vdd.n382 146.341
R2424 vdd.n3452 vdd.n382 146.341
R2425 vdd.n3452 vdd.n387 146.341
R2426 vdd.n3448 vdd.n387 146.341
R2427 vdd.n2378 vdd.n2377 146.341
R2428 vdd.n2375 vdd.n2372 146.341
R2429 vdd.n2370 vdd.n1127 146.341
R2430 vdd.n2366 vdd.n2365 146.341
R2431 vdd.n2363 vdd.n1131 146.341
R2432 vdd.n2359 vdd.n2358 146.341
R2433 vdd.n2356 vdd.n1138 146.341
R2434 vdd.n2352 vdd.n2351 146.341
R2435 vdd.n2349 vdd.n1145 146.341
R2436 vdd.n1156 vdd.n1153 146.341
R2437 vdd.n2341 vdd.n2340 146.341
R2438 vdd.n2338 vdd.n1158 146.341
R2439 vdd.n2334 vdd.n2333 146.341
R2440 vdd.n2331 vdd.n1164 146.341
R2441 vdd.n2327 vdd.n2326 146.341
R2442 vdd.n2324 vdd.n1171 146.341
R2443 vdd.n2320 vdd.n2319 146.341
R2444 vdd.n2317 vdd.n1178 146.341
R2445 vdd.n2313 vdd.n2312 146.341
R2446 vdd.n2310 vdd.n1185 146.341
R2447 vdd.n1196 vdd.n1193 146.341
R2448 vdd.n2302 vdd.n2301 146.341
R2449 vdd.n2299 vdd.n1198 146.341
R2450 vdd.n2295 vdd.n2294 146.341
R2451 vdd.n2292 vdd.n1204 146.341
R2452 vdd.n2288 vdd.n2287 146.341
R2453 vdd.n2285 vdd.n1211 146.341
R2454 vdd.n2281 vdd.n2280 146.341
R2455 vdd.n2278 vdd.n1218 146.341
R2456 vdd.n1429 vdd.n1427 146.341
R2457 vdd.n1432 vdd.n1431 146.341
R2458 vdd.n1790 vdd.n1550 146.341
R2459 vdd.n1790 vdd.n1546 146.341
R2460 vdd.n1796 vdd.n1546 146.341
R2461 vdd.n1796 vdd.n1538 146.341
R2462 vdd.n1807 vdd.n1538 146.341
R2463 vdd.n1807 vdd.n1534 146.341
R2464 vdd.n1813 vdd.n1534 146.341
R2465 vdd.n1813 vdd.n1528 146.341
R2466 vdd.n1824 vdd.n1528 146.341
R2467 vdd.n1824 vdd.n1524 146.341
R2468 vdd.n1830 vdd.n1524 146.341
R2469 vdd.n1830 vdd.n1515 146.341
R2470 vdd.n1840 vdd.n1515 146.341
R2471 vdd.n1840 vdd.n1511 146.341
R2472 vdd.n1846 vdd.n1511 146.341
R2473 vdd.n1846 vdd.n1504 146.341
R2474 vdd.n1857 vdd.n1504 146.341
R2475 vdd.n1857 vdd.n1500 146.341
R2476 vdd.n1863 vdd.n1500 146.341
R2477 vdd.n1863 vdd.n1493 146.341
R2478 vdd.n2180 vdd.n1493 146.341
R2479 vdd.n2180 vdd.n1489 146.341
R2480 vdd.n2186 vdd.n1489 146.341
R2481 vdd.n2186 vdd.n1481 146.341
R2482 vdd.n2197 vdd.n1481 146.341
R2483 vdd.n2197 vdd.n1477 146.341
R2484 vdd.n2203 vdd.n1477 146.341
R2485 vdd.n2203 vdd.n1471 146.341
R2486 vdd.n2214 vdd.n1471 146.341
R2487 vdd.n2214 vdd.n1467 146.341
R2488 vdd.n2220 vdd.n1467 146.341
R2489 vdd.n2220 vdd.n1458 146.341
R2490 vdd.n2230 vdd.n1458 146.341
R2491 vdd.n2230 vdd.n1454 146.341
R2492 vdd.n2236 vdd.n1454 146.341
R2493 vdd.n2236 vdd.n1448 146.341
R2494 vdd.n2247 vdd.n1448 146.341
R2495 vdd.n2247 vdd.n1443 146.341
R2496 vdd.n2255 vdd.n1443 146.341
R2497 vdd.n2255 vdd.n1434 146.341
R2498 vdd.n2266 vdd.n1434 146.341
R2499 vdd.n1779 vdd.n1555 146.341
R2500 vdd.n1779 vdd.n1588 146.341
R2501 vdd.n1592 vdd.n1591 146.341
R2502 vdd.n1594 vdd.n1593 146.341
R2503 vdd.n1598 vdd.n1597 146.341
R2504 vdd.n1600 vdd.n1599 146.341
R2505 vdd.n1604 vdd.n1603 146.341
R2506 vdd.n1606 vdd.n1605 146.341
R2507 vdd.n1610 vdd.n1609 146.341
R2508 vdd.n1612 vdd.n1611 146.341
R2509 vdd.n1618 vdd.n1617 146.341
R2510 vdd.n1620 vdd.n1619 146.341
R2511 vdd.n1624 vdd.n1623 146.341
R2512 vdd.n1626 vdd.n1625 146.341
R2513 vdd.n1630 vdd.n1629 146.341
R2514 vdd.n1632 vdd.n1631 146.341
R2515 vdd.n1636 vdd.n1635 146.341
R2516 vdd.n1638 vdd.n1637 146.341
R2517 vdd.n1642 vdd.n1641 146.341
R2518 vdd.n1644 vdd.n1643 146.341
R2519 vdd.n1716 vdd.n1647 146.341
R2520 vdd.n1649 vdd.n1648 146.341
R2521 vdd.n1653 vdd.n1652 146.341
R2522 vdd.n1655 vdd.n1654 146.341
R2523 vdd.n1659 vdd.n1658 146.341
R2524 vdd.n1661 vdd.n1660 146.341
R2525 vdd.n1665 vdd.n1664 146.341
R2526 vdd.n1667 vdd.n1666 146.341
R2527 vdd.n1671 vdd.n1670 146.341
R2528 vdd.n1673 vdd.n1672 146.341
R2529 vdd.n1677 vdd.n1676 146.341
R2530 vdd.n1678 vdd.n1586 146.341
R2531 vdd.n1788 vdd.n1551 146.341
R2532 vdd.n1788 vdd.n1544 146.341
R2533 vdd.n1799 vdd.n1544 146.341
R2534 vdd.n1799 vdd.n1540 146.341
R2535 vdd.n1805 vdd.n1540 146.341
R2536 vdd.n1805 vdd.n1533 146.341
R2537 vdd.n1816 vdd.n1533 146.341
R2538 vdd.n1816 vdd.n1529 146.341
R2539 vdd.n1822 vdd.n1529 146.341
R2540 vdd.n1822 vdd.n1522 146.341
R2541 vdd.n1832 vdd.n1522 146.341
R2542 vdd.n1832 vdd.n1518 146.341
R2543 vdd.n1838 vdd.n1518 146.341
R2544 vdd.n1838 vdd.n1510 146.341
R2545 vdd.n1849 vdd.n1510 146.341
R2546 vdd.n1849 vdd.n1506 146.341
R2547 vdd.n1855 vdd.n1506 146.341
R2548 vdd.n1855 vdd.n1499 146.341
R2549 vdd.n1865 vdd.n1499 146.341
R2550 vdd.n1865 vdd.n1495 146.341
R2551 vdd.n2178 vdd.n1495 146.341
R2552 vdd.n2178 vdd.n1487 146.341
R2553 vdd.n2189 vdd.n1487 146.341
R2554 vdd.n2189 vdd.n1483 146.341
R2555 vdd.n2195 vdd.n1483 146.341
R2556 vdd.n2195 vdd.n1476 146.341
R2557 vdd.n2206 vdd.n1476 146.341
R2558 vdd.n2206 vdd.n1472 146.341
R2559 vdd.n2212 vdd.n1472 146.341
R2560 vdd.n2212 vdd.n1465 146.341
R2561 vdd.n2222 vdd.n1465 146.341
R2562 vdd.n2222 vdd.n1461 146.341
R2563 vdd.n2228 vdd.n1461 146.341
R2564 vdd.n2228 vdd.n1453 146.341
R2565 vdd.n2239 vdd.n1453 146.341
R2566 vdd.n2239 vdd.n1449 146.341
R2567 vdd.n2245 vdd.n1449 146.341
R2568 vdd.n2245 vdd.n1441 146.341
R2569 vdd.n2258 vdd.n1441 146.341
R2570 vdd.n2258 vdd.n1436 146.341
R2571 vdd.n2264 vdd.n1436 146.341
R2572 vdd.n1253 vdd.t231 127.284
R2573 vdd.n981 vdd.t272 127.284
R2574 vdd.n1273 vdd.t245 127.284
R2575 vdd.n972 vdd.t295 127.284
R2576 vdd.n872 vdd.t252 127.284
R2577 vdd.n872 vdd.t253 127.284
R2578 vdd.n2704 vdd.t290 127.284
R2579 vdd.n832 vdd.t298 127.284
R2580 vdd.n2701 vdd.t277 127.284
R2581 vdd.n799 vdd.t226 127.284
R2582 vdd.n1043 vdd.t283 127.284
R2583 vdd.n1043 vdd.t284 127.284
R2584 vdd.n22 vdd.n20 117.314
R2585 vdd.n17 vdd.n15 117.314
R2586 vdd.n27 vdd.n26 116.927
R2587 vdd.n24 vdd.n23 116.927
R2588 vdd.n22 vdd.n21 116.927
R2589 vdd.n17 vdd.n16 116.927
R2590 vdd.n19 vdd.n18 116.927
R2591 vdd.n27 vdd.n25 116.927
R2592 vdd.n1254 vdd.t230 111.188
R2593 vdd.n982 vdd.t273 111.188
R2594 vdd.n1274 vdd.t244 111.188
R2595 vdd.n973 vdd.t296 111.188
R2596 vdd.n2705 vdd.t289 111.188
R2597 vdd.n833 vdd.t299 111.188
R2598 vdd.n2702 vdd.t276 111.188
R2599 vdd.n800 vdd.t227 111.188
R2600 vdd.n2946 vdd.n927 99.5127
R2601 vdd.n2946 vdd.n925 99.5127
R2602 vdd.n2950 vdd.n925 99.5127
R2603 vdd.n2950 vdd.n916 99.5127
R2604 vdd.n2958 vdd.n916 99.5127
R2605 vdd.n2958 vdd.n914 99.5127
R2606 vdd.n2962 vdd.n914 99.5127
R2607 vdd.n2962 vdd.n904 99.5127
R2608 vdd.n2970 vdd.n904 99.5127
R2609 vdd.n2970 vdd.n902 99.5127
R2610 vdd.n2974 vdd.n902 99.5127
R2611 vdd.n2974 vdd.n892 99.5127
R2612 vdd.n2982 vdd.n892 99.5127
R2613 vdd.n2982 vdd.n890 99.5127
R2614 vdd.n2986 vdd.n890 99.5127
R2615 vdd.n2986 vdd.n881 99.5127
R2616 vdd.n2994 vdd.n881 99.5127
R2617 vdd.n2994 vdd.n879 99.5127
R2618 vdd.n2998 vdd.n879 99.5127
R2619 vdd.n2998 vdd.n867 99.5127
R2620 vdd.n3007 vdd.n867 99.5127
R2621 vdd.n3007 vdd.n865 99.5127
R2622 vdd.n3011 vdd.n865 99.5127
R2623 vdd.n3011 vdd.n856 99.5127
R2624 vdd.n3019 vdd.n856 99.5127
R2625 vdd.n3019 vdd.n854 99.5127
R2626 vdd.n3023 vdd.n854 99.5127
R2627 vdd.n3023 vdd.n842 99.5127
R2628 vdd.n3076 vdd.n842 99.5127
R2629 vdd.n3076 vdd.n840 99.5127
R2630 vdd.n3080 vdd.n840 99.5127
R2631 vdd.n3080 vdd.n808 99.5127
R2632 vdd.n3150 vdd.n808 99.5127
R2633 vdd.n3146 vdd.n809 99.5127
R2634 vdd.n3144 vdd.n3143 99.5127
R2635 vdd.n3141 vdd.n813 99.5127
R2636 vdd.n3137 vdd.n3136 99.5127
R2637 vdd.n3134 vdd.n816 99.5127
R2638 vdd.n3130 vdd.n3129 99.5127
R2639 vdd.n3127 vdd.n819 99.5127
R2640 vdd.n3123 vdd.n3122 99.5127
R2641 vdd.n3120 vdd.n3118 99.5127
R2642 vdd.n3116 vdd.n822 99.5127
R2643 vdd.n3112 vdd.n3111 99.5127
R2644 vdd.n3109 vdd.n825 99.5127
R2645 vdd.n3105 vdd.n3104 99.5127
R2646 vdd.n3102 vdd.n828 99.5127
R2647 vdd.n3098 vdd.n3097 99.5127
R2648 vdd.n3095 vdd.n831 99.5127
R2649 vdd.n3090 vdd.n3089 99.5127
R2650 vdd.n2867 vdd.n929 99.5127
R2651 vdd.n2863 vdd.n929 99.5127
R2652 vdd.n2863 vdd.n923 99.5127
R2653 vdd.n2807 vdd.n923 99.5127
R2654 vdd.n2807 vdd.n918 99.5127
R2655 vdd.n2810 vdd.n918 99.5127
R2656 vdd.n2810 vdd.n912 99.5127
R2657 vdd.n2813 vdd.n912 99.5127
R2658 vdd.n2813 vdd.n906 99.5127
R2659 vdd.n2846 vdd.n906 99.5127
R2660 vdd.n2846 vdd.n899 99.5127
R2661 vdd.n2842 vdd.n899 99.5127
R2662 vdd.n2842 vdd.n893 99.5127
R2663 vdd.n2839 vdd.n893 99.5127
R2664 vdd.n2839 vdd.n888 99.5127
R2665 vdd.n2836 vdd.n888 99.5127
R2666 vdd.n2836 vdd.n883 99.5127
R2667 vdd.n2833 vdd.n883 99.5127
R2668 vdd.n2833 vdd.n876 99.5127
R2669 vdd.n2830 vdd.n876 99.5127
R2670 vdd.n2830 vdd.n868 99.5127
R2671 vdd.n2827 vdd.n868 99.5127
R2672 vdd.n2827 vdd.n863 99.5127
R2673 vdd.n2824 vdd.n863 99.5127
R2674 vdd.n2824 vdd.n858 99.5127
R2675 vdd.n2821 vdd.n858 99.5127
R2676 vdd.n2821 vdd.n852 99.5127
R2677 vdd.n2818 vdd.n852 99.5127
R2678 vdd.n2818 vdd.n844 99.5127
R2679 vdd.n844 vdd.n837 99.5127
R2680 vdd.n3082 vdd.n837 99.5127
R2681 vdd.n3083 vdd.n3082 99.5127
R2682 vdd.n3083 vdd.n806 99.5127
R2683 vdd.n2700 vdd.n2699 99.5127
R2684 vdd.n2931 vdd.n2699 99.5127
R2685 vdd.n2929 vdd.n2928 99.5127
R2686 vdd.n2925 vdd.n2924 99.5127
R2687 vdd.n2921 vdd.n2920 99.5127
R2688 vdd.n2917 vdd.n2916 99.5127
R2689 vdd.n2913 vdd.n2912 99.5127
R2690 vdd.n2909 vdd.n2908 99.5127
R2691 vdd.n2905 vdd.n2904 99.5127
R2692 vdd.n2901 vdd.n2900 99.5127
R2693 vdd.n2897 vdd.n2896 99.5127
R2694 vdd.n2893 vdd.n2892 99.5127
R2695 vdd.n2889 vdd.n2888 99.5127
R2696 vdd.n2885 vdd.n2884 99.5127
R2697 vdd.n2881 vdd.n2880 99.5127
R2698 vdd.n2877 vdd.n2876 99.5127
R2699 vdd.n2872 vdd.n2871 99.5127
R2700 vdd.n2664 vdd.n970 99.5127
R2701 vdd.n2660 vdd.n2659 99.5127
R2702 vdd.n2656 vdd.n2655 99.5127
R2703 vdd.n2652 vdd.n2651 99.5127
R2704 vdd.n2648 vdd.n2647 99.5127
R2705 vdd.n2644 vdd.n2643 99.5127
R2706 vdd.n2640 vdd.n2639 99.5127
R2707 vdd.n2636 vdd.n2635 99.5127
R2708 vdd.n2632 vdd.n2631 99.5127
R2709 vdd.n2628 vdd.n2627 99.5127
R2710 vdd.n2624 vdd.n2623 99.5127
R2711 vdd.n2620 vdd.n2619 99.5127
R2712 vdd.n2616 vdd.n2615 99.5127
R2713 vdd.n2612 vdd.n2611 99.5127
R2714 vdd.n2608 vdd.n2607 99.5127
R2715 vdd.n2604 vdd.n2603 99.5127
R2716 vdd.n2599 vdd.n2598 99.5127
R2717 vdd.n1309 vdd.n1077 99.5127
R2718 vdd.n1312 vdd.n1077 99.5127
R2719 vdd.n1312 vdd.n1071 99.5127
R2720 vdd.n1315 vdd.n1071 99.5127
R2721 vdd.n1315 vdd.n1066 99.5127
R2722 vdd.n1318 vdd.n1066 99.5127
R2723 vdd.n1318 vdd.n1060 99.5127
R2724 vdd.n1321 vdd.n1060 99.5127
R2725 vdd.n1321 vdd.n1053 99.5127
R2726 vdd.n1324 vdd.n1053 99.5127
R2727 vdd.n1324 vdd.n1046 99.5127
R2728 vdd.n1327 vdd.n1046 99.5127
R2729 vdd.n1327 vdd.n1040 99.5127
R2730 vdd.n1330 vdd.n1040 99.5127
R2731 vdd.n1330 vdd.n1035 99.5127
R2732 vdd.n1333 vdd.n1035 99.5127
R2733 vdd.n1333 vdd.n1029 99.5127
R2734 vdd.n1358 vdd.n1029 99.5127
R2735 vdd.n1358 vdd.n1022 99.5127
R2736 vdd.n1354 vdd.n1022 99.5127
R2737 vdd.n1354 vdd.n1016 99.5127
R2738 vdd.n1351 vdd.n1016 99.5127
R2739 vdd.n1351 vdd.n1011 99.5127
R2740 vdd.n1348 vdd.n1011 99.5127
R2741 vdd.n1348 vdd.n1006 99.5127
R2742 vdd.n1345 vdd.n1006 99.5127
R2743 vdd.n1345 vdd.n1000 99.5127
R2744 vdd.n1342 vdd.n1000 99.5127
R2745 vdd.n1342 vdd.n993 99.5127
R2746 vdd.n1339 vdd.n993 99.5127
R2747 vdd.n1339 vdd.n986 99.5127
R2748 vdd.n986 vdd.n975 99.5127
R2749 vdd.n2594 vdd.n975 99.5127
R2750 vdd.n1118 vdd.n1117 99.5127
R2751 vdd.n2410 vdd.n1117 99.5127
R2752 vdd.n2408 vdd.n2407 99.5127
R2753 vdd.n2404 vdd.n2403 99.5127
R2754 vdd.n2400 vdd.n2399 99.5127
R2755 vdd.n2396 vdd.n2395 99.5127
R2756 vdd.n2392 vdd.n2391 99.5127
R2757 vdd.n2388 vdd.n2387 99.5127
R2758 vdd.n2384 vdd.n2383 99.5127
R2759 vdd.n1276 vdd.n1275 99.5127
R2760 vdd.n1280 vdd.n1279 99.5127
R2761 vdd.n1284 vdd.n1283 99.5127
R2762 vdd.n1288 vdd.n1287 99.5127
R2763 vdd.n1292 vdd.n1291 99.5127
R2764 vdd.n1296 vdd.n1295 99.5127
R2765 vdd.n1300 vdd.n1299 99.5127
R2766 vdd.n1305 vdd.n1304 99.5127
R2767 vdd.n2425 vdd.n1075 99.5127
R2768 vdd.n2425 vdd.n1073 99.5127
R2769 vdd.n2429 vdd.n1073 99.5127
R2770 vdd.n2429 vdd.n1064 99.5127
R2771 vdd.n2437 vdd.n1064 99.5127
R2772 vdd.n2437 vdd.n1062 99.5127
R2773 vdd.n2441 vdd.n1062 99.5127
R2774 vdd.n2441 vdd.n1051 99.5127
R2775 vdd.n2449 vdd.n1051 99.5127
R2776 vdd.n2449 vdd.n1049 99.5127
R2777 vdd.n2453 vdd.n1049 99.5127
R2778 vdd.n2453 vdd.n1039 99.5127
R2779 vdd.n2462 vdd.n1039 99.5127
R2780 vdd.n2462 vdd.n1037 99.5127
R2781 vdd.n2466 vdd.n1037 99.5127
R2782 vdd.n2466 vdd.n1027 99.5127
R2783 vdd.n2474 vdd.n1027 99.5127
R2784 vdd.n2474 vdd.n1025 99.5127
R2785 vdd.n2478 vdd.n1025 99.5127
R2786 vdd.n2478 vdd.n1015 99.5127
R2787 vdd.n2486 vdd.n1015 99.5127
R2788 vdd.n2486 vdd.n1013 99.5127
R2789 vdd.n2490 vdd.n1013 99.5127
R2790 vdd.n2490 vdd.n1004 99.5127
R2791 vdd.n2498 vdd.n1004 99.5127
R2792 vdd.n2498 vdd.n1002 99.5127
R2793 vdd.n2502 vdd.n1002 99.5127
R2794 vdd.n2502 vdd.n991 99.5127
R2795 vdd.n2512 vdd.n991 99.5127
R2796 vdd.n2512 vdd.n988 99.5127
R2797 vdd.n2517 vdd.n988 99.5127
R2798 vdd.n2517 vdd.n989 99.5127
R2799 vdd.n989 vdd.n969 99.5127
R2800 vdd.n3066 vdd.n3065 99.5127
R2801 vdd.n3063 vdd.n3029 99.5127
R2802 vdd.n3059 vdd.n3058 99.5127
R2803 vdd.n3056 vdd.n3032 99.5127
R2804 vdd.n3052 vdd.n3051 99.5127
R2805 vdd.n3049 vdd.n3035 99.5127
R2806 vdd.n3045 vdd.n3044 99.5127
R2807 vdd.n3042 vdd.n3039 99.5127
R2808 vdd.n3183 vdd.n787 99.5127
R2809 vdd.n3181 vdd.n3180 99.5127
R2810 vdd.n3178 vdd.n789 99.5127
R2811 vdd.n3174 vdd.n3173 99.5127
R2812 vdd.n3171 vdd.n792 99.5127
R2813 vdd.n3167 vdd.n3166 99.5127
R2814 vdd.n3164 vdd.n795 99.5127
R2815 vdd.n3160 vdd.n3159 99.5127
R2816 vdd.n3157 vdd.n798 99.5127
R2817 vdd.n2772 vdd.n930 99.5127
R2818 vdd.n2861 vdd.n930 99.5127
R2819 vdd.n2861 vdd.n924 99.5127
R2820 vdd.n2857 vdd.n924 99.5127
R2821 vdd.n2857 vdd.n919 99.5127
R2822 vdd.n2854 vdd.n919 99.5127
R2823 vdd.n2854 vdd.n913 99.5127
R2824 vdd.n2851 vdd.n913 99.5127
R2825 vdd.n2851 vdd.n907 99.5127
R2826 vdd.n2848 vdd.n907 99.5127
R2827 vdd.n2848 vdd.n900 99.5127
R2828 vdd.n2804 vdd.n900 99.5127
R2829 vdd.n2804 vdd.n894 99.5127
R2830 vdd.n2801 vdd.n894 99.5127
R2831 vdd.n2801 vdd.n889 99.5127
R2832 vdd.n2798 vdd.n889 99.5127
R2833 vdd.n2798 vdd.n884 99.5127
R2834 vdd.n2795 vdd.n884 99.5127
R2835 vdd.n2795 vdd.n877 99.5127
R2836 vdd.n2792 vdd.n877 99.5127
R2837 vdd.n2792 vdd.n869 99.5127
R2838 vdd.n2789 vdd.n869 99.5127
R2839 vdd.n2789 vdd.n864 99.5127
R2840 vdd.n2786 vdd.n864 99.5127
R2841 vdd.n2786 vdd.n859 99.5127
R2842 vdd.n2783 vdd.n859 99.5127
R2843 vdd.n2783 vdd.n853 99.5127
R2844 vdd.n2780 vdd.n853 99.5127
R2845 vdd.n2780 vdd.n845 99.5127
R2846 vdd.n2777 vdd.n845 99.5127
R2847 vdd.n2777 vdd.n838 99.5127
R2848 vdd.n838 vdd.n804 99.5127
R2849 vdd.n3152 vdd.n804 99.5127
R2850 vdd.n2707 vdd.n933 99.5127
R2851 vdd.n2711 vdd.n2710 99.5127
R2852 vdd.n2715 vdd.n2714 99.5127
R2853 vdd.n2719 vdd.n2718 99.5127
R2854 vdd.n2723 vdd.n2722 99.5127
R2855 vdd.n2727 vdd.n2726 99.5127
R2856 vdd.n2731 vdd.n2730 99.5127
R2857 vdd.n2735 vdd.n2734 99.5127
R2858 vdd.n2739 vdd.n2738 99.5127
R2859 vdd.n2743 vdd.n2742 99.5127
R2860 vdd.n2747 vdd.n2746 99.5127
R2861 vdd.n2751 vdd.n2750 99.5127
R2862 vdd.n2755 vdd.n2754 99.5127
R2863 vdd.n2759 vdd.n2758 99.5127
R2864 vdd.n2763 vdd.n2762 99.5127
R2865 vdd.n2767 vdd.n2766 99.5127
R2866 vdd.n2769 vdd.n2698 99.5127
R2867 vdd.n2944 vdd.n931 99.5127
R2868 vdd.n2944 vdd.n922 99.5127
R2869 vdd.n2952 vdd.n922 99.5127
R2870 vdd.n2952 vdd.n920 99.5127
R2871 vdd.n2956 vdd.n920 99.5127
R2872 vdd.n2956 vdd.n910 99.5127
R2873 vdd.n2964 vdd.n910 99.5127
R2874 vdd.n2964 vdd.n908 99.5127
R2875 vdd.n2968 vdd.n908 99.5127
R2876 vdd.n2968 vdd.n898 99.5127
R2877 vdd.n2976 vdd.n898 99.5127
R2878 vdd.n2976 vdd.n896 99.5127
R2879 vdd.n2980 vdd.n896 99.5127
R2880 vdd.n2980 vdd.n887 99.5127
R2881 vdd.n2988 vdd.n887 99.5127
R2882 vdd.n2988 vdd.n885 99.5127
R2883 vdd.n2992 vdd.n885 99.5127
R2884 vdd.n2992 vdd.n874 99.5127
R2885 vdd.n3000 vdd.n874 99.5127
R2886 vdd.n3000 vdd.n871 99.5127
R2887 vdd.n3005 vdd.n871 99.5127
R2888 vdd.n3005 vdd.n862 99.5127
R2889 vdd.n3013 vdd.n862 99.5127
R2890 vdd.n3013 vdd.n860 99.5127
R2891 vdd.n3017 vdd.n860 99.5127
R2892 vdd.n3017 vdd.n850 99.5127
R2893 vdd.n3025 vdd.n850 99.5127
R2894 vdd.n3025 vdd.n847 99.5127
R2895 vdd.n3074 vdd.n847 99.5127
R2896 vdd.n3074 vdd.n848 99.5127
R2897 vdd.n848 vdd.n839 99.5127
R2898 vdd.n3069 vdd.n839 99.5127
R2899 vdd.n3069 vdd.n807 99.5127
R2900 vdd.n2588 vdd.n2587 99.5127
R2901 vdd.n2584 vdd.n2583 99.5127
R2902 vdd.n2580 vdd.n2579 99.5127
R2903 vdd.n2576 vdd.n2575 99.5127
R2904 vdd.n2572 vdd.n2571 99.5127
R2905 vdd.n2568 vdd.n2567 99.5127
R2906 vdd.n2564 vdd.n2563 99.5127
R2907 vdd.n2560 vdd.n2559 99.5127
R2908 vdd.n2556 vdd.n2555 99.5127
R2909 vdd.n2552 vdd.n2551 99.5127
R2910 vdd.n2548 vdd.n2547 99.5127
R2911 vdd.n2544 vdd.n2543 99.5127
R2912 vdd.n2540 vdd.n2539 99.5127
R2913 vdd.n2536 vdd.n2535 99.5127
R2914 vdd.n2532 vdd.n2531 99.5127
R2915 vdd.n2528 vdd.n2527 99.5127
R2916 vdd.n2524 vdd.n951 99.5127
R2917 vdd.n1387 vdd.n1078 99.5127
R2918 vdd.n1384 vdd.n1078 99.5127
R2919 vdd.n1384 vdd.n1072 99.5127
R2920 vdd.n1381 vdd.n1072 99.5127
R2921 vdd.n1381 vdd.n1067 99.5127
R2922 vdd.n1378 vdd.n1067 99.5127
R2923 vdd.n1378 vdd.n1061 99.5127
R2924 vdd.n1375 vdd.n1061 99.5127
R2925 vdd.n1375 vdd.n1054 99.5127
R2926 vdd.n1372 vdd.n1054 99.5127
R2927 vdd.n1372 vdd.n1047 99.5127
R2928 vdd.n1369 vdd.n1047 99.5127
R2929 vdd.n1369 vdd.n1041 99.5127
R2930 vdd.n1366 vdd.n1041 99.5127
R2931 vdd.n1366 vdd.n1036 99.5127
R2932 vdd.n1363 vdd.n1036 99.5127
R2933 vdd.n1363 vdd.n1030 99.5127
R2934 vdd.n1360 vdd.n1030 99.5127
R2935 vdd.n1360 vdd.n1023 99.5127
R2936 vdd.n1270 vdd.n1023 99.5127
R2937 vdd.n1270 vdd.n1017 99.5127
R2938 vdd.n1267 vdd.n1017 99.5127
R2939 vdd.n1267 vdd.n1012 99.5127
R2940 vdd.n1264 vdd.n1012 99.5127
R2941 vdd.n1264 vdd.n1007 99.5127
R2942 vdd.n1261 vdd.n1007 99.5127
R2943 vdd.n1261 vdd.n1001 99.5127
R2944 vdd.n1258 vdd.n1001 99.5127
R2945 vdd.n1258 vdd.n994 99.5127
R2946 vdd.n994 vdd.n985 99.5127
R2947 vdd.n2519 vdd.n985 99.5127
R2948 vdd.n2520 vdd.n2519 99.5127
R2949 vdd.n2520 vdd.n977 99.5127
R2950 vdd.n1222 vdd.n1082 99.5127
R2951 vdd.n1226 vdd.n1225 99.5127
R2952 vdd.n1230 vdd.n1229 99.5127
R2953 vdd.n1234 vdd.n1233 99.5127
R2954 vdd.n1238 vdd.n1237 99.5127
R2955 vdd.n1242 vdd.n1241 99.5127
R2956 vdd.n1246 vdd.n1245 99.5127
R2957 vdd.n1250 vdd.n1249 99.5127
R2958 vdd.n1420 vdd.n1252 99.5127
R2959 vdd.n1418 vdd.n1417 99.5127
R2960 vdd.n1414 vdd.n1413 99.5127
R2961 vdd.n1410 vdd.n1409 99.5127
R2962 vdd.n1406 vdd.n1405 99.5127
R2963 vdd.n1402 vdd.n1401 99.5127
R2964 vdd.n1398 vdd.n1397 99.5127
R2965 vdd.n1394 vdd.n1393 99.5127
R2966 vdd.n1390 vdd.n1116 99.5127
R2967 vdd.n2423 vdd.n1080 99.5127
R2968 vdd.n2423 vdd.n1070 99.5127
R2969 vdd.n2431 vdd.n1070 99.5127
R2970 vdd.n2431 vdd.n1068 99.5127
R2971 vdd.n2435 vdd.n1068 99.5127
R2972 vdd.n2435 vdd.n1058 99.5127
R2973 vdd.n2443 vdd.n1058 99.5127
R2974 vdd.n2443 vdd.n1056 99.5127
R2975 vdd.n2447 vdd.n1056 99.5127
R2976 vdd.n2447 vdd.n1045 99.5127
R2977 vdd.n2455 vdd.n1045 99.5127
R2978 vdd.n2455 vdd.n1042 99.5127
R2979 vdd.n2460 vdd.n1042 99.5127
R2980 vdd.n2460 vdd.n1033 99.5127
R2981 vdd.n2468 vdd.n1033 99.5127
R2982 vdd.n2468 vdd.n1031 99.5127
R2983 vdd.n2472 vdd.n1031 99.5127
R2984 vdd.n2472 vdd.n1021 99.5127
R2985 vdd.n2480 vdd.n1021 99.5127
R2986 vdd.n2480 vdd.n1019 99.5127
R2987 vdd.n2484 vdd.n1019 99.5127
R2988 vdd.n2484 vdd.n1010 99.5127
R2989 vdd.n2492 vdd.n1010 99.5127
R2990 vdd.n2492 vdd.n1008 99.5127
R2991 vdd.n2496 vdd.n1008 99.5127
R2992 vdd.n2496 vdd.n998 99.5127
R2993 vdd.n2504 vdd.n998 99.5127
R2994 vdd.n2504 vdd.n995 99.5127
R2995 vdd.n2510 vdd.n995 99.5127
R2996 vdd.n2510 vdd.n996 99.5127
R2997 vdd.n996 vdd.n987 99.5127
R2998 vdd.n987 vdd.n978 99.5127
R2999 vdd.n2592 vdd.n978 99.5127
R3000 vdd.n9 vdd.n7 98.9633
R3001 vdd.n2 vdd.n0 98.9633
R3002 vdd.n9 vdd.n8 98.6055
R3003 vdd.n11 vdd.n10 98.6055
R3004 vdd.n13 vdd.n12 98.6055
R3005 vdd.n6 vdd.n5 98.6055
R3006 vdd.n4 vdd.n3 98.6055
R3007 vdd.n2 vdd.n1 98.6055
R3008 vdd.t88 vdd.n303 85.8723
R3009 vdd.t168 vdd.n244 85.8723
R3010 vdd.t219 vdd.n201 85.8723
R3011 vdd.t152 vdd.n142 85.8723
R3012 vdd.t120 vdd.n100 85.8723
R3013 vdd.t113 vdd.n41 85.8723
R3014 vdd.t210 vdd.n2084 85.8723
R3015 vdd.t144 vdd.n2143 85.8723
R3016 vdd.t198 vdd.n1982 85.8723
R3017 vdd.t121 vdd.n2041 85.8723
R3018 vdd.t115 vdd.n1881 85.8723
R3019 vdd.t73 vdd.n1940 85.8723
R3020 vdd.n3003 vdd.n872 78.546
R3021 vdd.n2458 vdd.n1043 78.546
R3022 vdd.n290 vdd.n289 75.1835
R3023 vdd.n288 vdd.n287 75.1835
R3024 vdd.n286 vdd.n285 75.1835
R3025 vdd.n284 vdd.n283 75.1835
R3026 vdd.n282 vdd.n281 75.1835
R3027 vdd.n280 vdd.n279 75.1835
R3028 vdd.n278 vdd.n277 75.1835
R3029 vdd.n276 vdd.n275 75.1835
R3030 vdd.n274 vdd.n273 75.1835
R3031 vdd.n188 vdd.n187 75.1835
R3032 vdd.n186 vdd.n185 75.1835
R3033 vdd.n184 vdd.n183 75.1835
R3034 vdd.n182 vdd.n181 75.1835
R3035 vdd.n180 vdd.n179 75.1835
R3036 vdd.n178 vdd.n177 75.1835
R3037 vdd.n176 vdd.n175 75.1835
R3038 vdd.n174 vdd.n173 75.1835
R3039 vdd.n172 vdd.n171 75.1835
R3040 vdd.n87 vdd.n86 75.1835
R3041 vdd.n85 vdd.n84 75.1835
R3042 vdd.n83 vdd.n82 75.1835
R3043 vdd.n81 vdd.n80 75.1835
R3044 vdd.n79 vdd.n78 75.1835
R3045 vdd.n77 vdd.n76 75.1835
R3046 vdd.n75 vdd.n74 75.1835
R3047 vdd.n73 vdd.n72 75.1835
R3048 vdd.n71 vdd.n70 75.1835
R3049 vdd.n2114 vdd.n2113 75.1835
R3050 vdd.n2116 vdd.n2115 75.1835
R3051 vdd.n2118 vdd.n2117 75.1835
R3052 vdd.n2120 vdd.n2119 75.1835
R3053 vdd.n2122 vdd.n2121 75.1835
R3054 vdd.n2124 vdd.n2123 75.1835
R3055 vdd.n2126 vdd.n2125 75.1835
R3056 vdd.n2128 vdd.n2127 75.1835
R3057 vdd.n2130 vdd.n2129 75.1835
R3058 vdd.n2012 vdd.n2011 75.1835
R3059 vdd.n2014 vdd.n2013 75.1835
R3060 vdd.n2016 vdd.n2015 75.1835
R3061 vdd.n2018 vdd.n2017 75.1835
R3062 vdd.n2020 vdd.n2019 75.1835
R3063 vdd.n2022 vdd.n2021 75.1835
R3064 vdd.n2024 vdd.n2023 75.1835
R3065 vdd.n2026 vdd.n2025 75.1835
R3066 vdd.n2028 vdd.n2027 75.1835
R3067 vdd.n1911 vdd.n1910 75.1835
R3068 vdd.n1913 vdd.n1912 75.1835
R3069 vdd.n1915 vdd.n1914 75.1835
R3070 vdd.n1917 vdd.n1916 75.1835
R3071 vdd.n1919 vdd.n1918 75.1835
R3072 vdd.n1921 vdd.n1920 75.1835
R3073 vdd.n1923 vdd.n1922 75.1835
R3074 vdd.n1925 vdd.n1924 75.1835
R3075 vdd.n1927 vdd.n1926 75.1835
R3076 vdd.n2939 vdd.n2938 72.8958
R3077 vdd.n2938 vdd.n2682 72.8958
R3078 vdd.n2938 vdd.n2683 72.8958
R3079 vdd.n2938 vdd.n2684 72.8958
R3080 vdd.n2938 vdd.n2685 72.8958
R3081 vdd.n2938 vdd.n2686 72.8958
R3082 vdd.n2938 vdd.n2687 72.8958
R3083 vdd.n2938 vdd.n2688 72.8958
R3084 vdd.n2938 vdd.n2689 72.8958
R3085 vdd.n2938 vdd.n2690 72.8958
R3086 vdd.n2938 vdd.n2691 72.8958
R3087 vdd.n2938 vdd.n2692 72.8958
R3088 vdd.n2938 vdd.n2693 72.8958
R3089 vdd.n2938 vdd.n2694 72.8958
R3090 vdd.n2938 vdd.n2695 72.8958
R3091 vdd.n2938 vdd.n2696 72.8958
R3092 vdd.n2938 vdd.n2697 72.8958
R3093 vdd.n803 vdd.n692 72.8958
R3094 vdd.n3158 vdd.n692 72.8958
R3095 vdd.n797 vdd.n692 72.8958
R3096 vdd.n3165 vdd.n692 72.8958
R3097 vdd.n794 vdd.n692 72.8958
R3098 vdd.n3172 vdd.n692 72.8958
R3099 vdd.n791 vdd.n692 72.8958
R3100 vdd.n3179 vdd.n692 72.8958
R3101 vdd.n3182 vdd.n692 72.8958
R3102 vdd.n3038 vdd.n692 72.8958
R3103 vdd.n3043 vdd.n692 72.8958
R3104 vdd.n3037 vdd.n692 72.8958
R3105 vdd.n3050 vdd.n692 72.8958
R3106 vdd.n3034 vdd.n692 72.8958
R3107 vdd.n3057 vdd.n692 72.8958
R3108 vdd.n3031 vdd.n692 72.8958
R3109 vdd.n3064 vdd.n692 72.8958
R3110 vdd.n2417 vdd.n2416 72.8958
R3111 vdd.n2417 vdd.n1084 72.8958
R3112 vdd.n2417 vdd.n1085 72.8958
R3113 vdd.n2417 vdd.n1086 72.8958
R3114 vdd.n2417 vdd.n1087 72.8958
R3115 vdd.n2417 vdd.n1088 72.8958
R3116 vdd.n2417 vdd.n1089 72.8958
R3117 vdd.n2417 vdd.n1090 72.8958
R3118 vdd.n2417 vdd.n1091 72.8958
R3119 vdd.n2417 vdd.n1092 72.8958
R3120 vdd.n2417 vdd.n1093 72.8958
R3121 vdd.n2417 vdd.n1094 72.8958
R3122 vdd.n2417 vdd.n1095 72.8958
R3123 vdd.n2417 vdd.n1096 72.8958
R3124 vdd.n2417 vdd.n1097 72.8958
R3125 vdd.n2417 vdd.n1098 72.8958
R3126 vdd.n2417 vdd.n1099 72.8958
R3127 vdd.n2665 vdd.n952 72.8958
R3128 vdd.n2665 vdd.n953 72.8958
R3129 vdd.n2665 vdd.n954 72.8958
R3130 vdd.n2665 vdd.n955 72.8958
R3131 vdd.n2665 vdd.n956 72.8958
R3132 vdd.n2665 vdd.n957 72.8958
R3133 vdd.n2665 vdd.n958 72.8958
R3134 vdd.n2665 vdd.n959 72.8958
R3135 vdd.n2665 vdd.n960 72.8958
R3136 vdd.n2665 vdd.n961 72.8958
R3137 vdd.n2665 vdd.n962 72.8958
R3138 vdd.n2665 vdd.n963 72.8958
R3139 vdd.n2665 vdd.n964 72.8958
R3140 vdd.n2665 vdd.n965 72.8958
R3141 vdd.n2665 vdd.n966 72.8958
R3142 vdd.n2665 vdd.n967 72.8958
R3143 vdd.n2665 vdd.n968 72.8958
R3144 vdd.n2938 vdd.n2937 72.8958
R3145 vdd.n2938 vdd.n2666 72.8958
R3146 vdd.n2938 vdd.n2667 72.8958
R3147 vdd.n2938 vdd.n2668 72.8958
R3148 vdd.n2938 vdd.n2669 72.8958
R3149 vdd.n2938 vdd.n2670 72.8958
R3150 vdd.n2938 vdd.n2671 72.8958
R3151 vdd.n2938 vdd.n2672 72.8958
R3152 vdd.n2938 vdd.n2673 72.8958
R3153 vdd.n2938 vdd.n2674 72.8958
R3154 vdd.n2938 vdd.n2675 72.8958
R3155 vdd.n2938 vdd.n2676 72.8958
R3156 vdd.n2938 vdd.n2677 72.8958
R3157 vdd.n2938 vdd.n2678 72.8958
R3158 vdd.n2938 vdd.n2679 72.8958
R3159 vdd.n2938 vdd.n2680 72.8958
R3160 vdd.n2938 vdd.n2681 72.8958
R3161 vdd.n3088 vdd.n692 72.8958
R3162 vdd.n835 vdd.n692 72.8958
R3163 vdd.n3096 vdd.n692 72.8958
R3164 vdd.n830 vdd.n692 72.8958
R3165 vdd.n3103 vdd.n692 72.8958
R3166 vdd.n827 vdd.n692 72.8958
R3167 vdd.n3110 vdd.n692 72.8958
R3168 vdd.n824 vdd.n692 72.8958
R3169 vdd.n3117 vdd.n692 72.8958
R3170 vdd.n3121 vdd.n692 72.8958
R3171 vdd.n821 vdd.n692 72.8958
R3172 vdd.n3128 vdd.n692 72.8958
R3173 vdd.n818 vdd.n692 72.8958
R3174 vdd.n3135 vdd.n692 72.8958
R3175 vdd.n815 vdd.n692 72.8958
R3176 vdd.n3142 vdd.n692 72.8958
R3177 vdd.n3145 vdd.n692 72.8958
R3178 vdd.n2665 vdd.n950 72.8958
R3179 vdd.n2665 vdd.n949 72.8958
R3180 vdd.n2665 vdd.n948 72.8958
R3181 vdd.n2665 vdd.n947 72.8958
R3182 vdd.n2665 vdd.n946 72.8958
R3183 vdd.n2665 vdd.n945 72.8958
R3184 vdd.n2665 vdd.n944 72.8958
R3185 vdd.n2665 vdd.n943 72.8958
R3186 vdd.n2665 vdd.n942 72.8958
R3187 vdd.n2665 vdd.n941 72.8958
R3188 vdd.n2665 vdd.n940 72.8958
R3189 vdd.n2665 vdd.n939 72.8958
R3190 vdd.n2665 vdd.n938 72.8958
R3191 vdd.n2665 vdd.n937 72.8958
R3192 vdd.n2665 vdd.n936 72.8958
R3193 vdd.n2665 vdd.n935 72.8958
R3194 vdd.n2665 vdd.n934 72.8958
R3195 vdd.n2418 vdd.n2417 72.8958
R3196 vdd.n2417 vdd.n1100 72.8958
R3197 vdd.n2417 vdd.n1101 72.8958
R3198 vdd.n2417 vdd.n1102 72.8958
R3199 vdd.n2417 vdd.n1103 72.8958
R3200 vdd.n2417 vdd.n1104 72.8958
R3201 vdd.n2417 vdd.n1105 72.8958
R3202 vdd.n2417 vdd.n1106 72.8958
R3203 vdd.n2417 vdd.n1107 72.8958
R3204 vdd.n2417 vdd.n1108 72.8958
R3205 vdd.n2417 vdd.n1109 72.8958
R3206 vdd.n2417 vdd.n1110 72.8958
R3207 vdd.n2417 vdd.n1111 72.8958
R3208 vdd.n2417 vdd.n1112 72.8958
R3209 vdd.n2417 vdd.n1113 72.8958
R3210 vdd.n2417 vdd.n1114 72.8958
R3211 vdd.n2417 vdd.n1115 72.8958
R3212 vdd.n1781 vdd.n1780 66.2847
R3213 vdd.n1780 vdd.n1556 66.2847
R3214 vdd.n1780 vdd.n1557 66.2847
R3215 vdd.n1780 vdd.n1558 66.2847
R3216 vdd.n1780 vdd.n1559 66.2847
R3217 vdd.n1780 vdd.n1560 66.2847
R3218 vdd.n1780 vdd.n1561 66.2847
R3219 vdd.n1780 vdd.n1562 66.2847
R3220 vdd.n1780 vdd.n1563 66.2847
R3221 vdd.n1780 vdd.n1564 66.2847
R3222 vdd.n1780 vdd.n1565 66.2847
R3223 vdd.n1780 vdd.n1566 66.2847
R3224 vdd.n1780 vdd.n1567 66.2847
R3225 vdd.n1780 vdd.n1568 66.2847
R3226 vdd.n1780 vdd.n1569 66.2847
R3227 vdd.n1780 vdd.n1570 66.2847
R3228 vdd.n1780 vdd.n1571 66.2847
R3229 vdd.n1780 vdd.n1572 66.2847
R3230 vdd.n1780 vdd.n1573 66.2847
R3231 vdd.n1780 vdd.n1574 66.2847
R3232 vdd.n1780 vdd.n1575 66.2847
R3233 vdd.n1780 vdd.n1576 66.2847
R3234 vdd.n1780 vdd.n1577 66.2847
R3235 vdd.n1780 vdd.n1578 66.2847
R3236 vdd.n1780 vdd.n1579 66.2847
R3237 vdd.n1780 vdd.n1580 66.2847
R3238 vdd.n1780 vdd.n1581 66.2847
R3239 vdd.n1780 vdd.n1582 66.2847
R3240 vdd.n1780 vdd.n1583 66.2847
R3241 vdd.n1780 vdd.n1584 66.2847
R3242 vdd.n1780 vdd.n1585 66.2847
R3243 vdd.n1433 vdd.n1083 66.2847
R3244 vdd.n1430 vdd.n1083 66.2847
R3245 vdd.n1426 vdd.n1083 66.2847
R3246 vdd.n2279 vdd.n1083 66.2847
R3247 vdd.n1217 vdd.n1083 66.2847
R3248 vdd.n2286 vdd.n1083 66.2847
R3249 vdd.n1210 vdd.n1083 66.2847
R3250 vdd.n2293 vdd.n1083 66.2847
R3251 vdd.n1203 vdd.n1083 66.2847
R3252 vdd.n2300 vdd.n1083 66.2847
R3253 vdd.n1197 vdd.n1083 66.2847
R3254 vdd.n1192 vdd.n1083 66.2847
R3255 vdd.n2311 vdd.n1083 66.2847
R3256 vdd.n1184 vdd.n1083 66.2847
R3257 vdd.n2318 vdd.n1083 66.2847
R3258 vdd.n1177 vdd.n1083 66.2847
R3259 vdd.n2325 vdd.n1083 66.2847
R3260 vdd.n1170 vdd.n1083 66.2847
R3261 vdd.n2332 vdd.n1083 66.2847
R3262 vdd.n1163 vdd.n1083 66.2847
R3263 vdd.n2339 vdd.n1083 66.2847
R3264 vdd.n1157 vdd.n1083 66.2847
R3265 vdd.n1152 vdd.n1083 66.2847
R3266 vdd.n2350 vdd.n1083 66.2847
R3267 vdd.n1144 vdd.n1083 66.2847
R3268 vdd.n2357 vdd.n1083 66.2847
R3269 vdd.n1137 vdd.n1083 66.2847
R3270 vdd.n2364 vdd.n1083 66.2847
R3271 vdd.n1130 vdd.n1083 66.2847
R3272 vdd.n2371 vdd.n1083 66.2847
R3273 vdd.n2376 vdd.n1083 66.2847
R3274 vdd.n1126 vdd.n1083 66.2847
R3275 vdd.n3315 vdd.n3314 66.2847
R3276 vdd.n3315 vdd.n693 66.2847
R3277 vdd.n3315 vdd.n694 66.2847
R3278 vdd.n3315 vdd.n695 66.2847
R3279 vdd.n3315 vdd.n696 66.2847
R3280 vdd.n3315 vdd.n697 66.2847
R3281 vdd.n3315 vdd.n698 66.2847
R3282 vdd.n3315 vdd.n699 66.2847
R3283 vdd.n3315 vdd.n700 66.2847
R3284 vdd.n3315 vdd.n701 66.2847
R3285 vdd.n3315 vdd.n702 66.2847
R3286 vdd.n3315 vdd.n703 66.2847
R3287 vdd.n3315 vdd.n704 66.2847
R3288 vdd.n3315 vdd.n705 66.2847
R3289 vdd.n3315 vdd.n706 66.2847
R3290 vdd.n3315 vdd.n707 66.2847
R3291 vdd.n3315 vdd.n708 66.2847
R3292 vdd.n3315 vdd.n709 66.2847
R3293 vdd.n3315 vdd.n710 66.2847
R3294 vdd.n3315 vdd.n711 66.2847
R3295 vdd.n3315 vdd.n712 66.2847
R3296 vdd.n3315 vdd.n713 66.2847
R3297 vdd.n3315 vdd.n714 66.2847
R3298 vdd.n3315 vdd.n715 66.2847
R3299 vdd.n3315 vdd.n716 66.2847
R3300 vdd.n3315 vdd.n717 66.2847
R3301 vdd.n3315 vdd.n718 66.2847
R3302 vdd.n3315 vdd.n719 66.2847
R3303 vdd.n3315 vdd.n720 66.2847
R3304 vdd.n3315 vdd.n721 66.2847
R3305 vdd.n3315 vdd.n722 66.2847
R3306 vdd.n3446 vdd.n3445 66.2847
R3307 vdd.n3446 vdd.n424 66.2847
R3308 vdd.n3446 vdd.n423 66.2847
R3309 vdd.n3446 vdd.n422 66.2847
R3310 vdd.n3446 vdd.n421 66.2847
R3311 vdd.n3446 vdd.n420 66.2847
R3312 vdd.n3446 vdd.n419 66.2847
R3313 vdd.n3446 vdd.n418 66.2847
R3314 vdd.n3446 vdd.n417 66.2847
R3315 vdd.n3446 vdd.n416 66.2847
R3316 vdd.n3446 vdd.n415 66.2847
R3317 vdd.n3446 vdd.n414 66.2847
R3318 vdd.n3446 vdd.n413 66.2847
R3319 vdd.n3446 vdd.n412 66.2847
R3320 vdd.n3446 vdd.n411 66.2847
R3321 vdd.n3446 vdd.n410 66.2847
R3322 vdd.n3446 vdd.n409 66.2847
R3323 vdd.n3446 vdd.n408 66.2847
R3324 vdd.n3446 vdd.n407 66.2847
R3325 vdd.n3446 vdd.n406 66.2847
R3326 vdd.n3446 vdd.n405 66.2847
R3327 vdd.n3446 vdd.n404 66.2847
R3328 vdd.n3446 vdd.n403 66.2847
R3329 vdd.n3446 vdd.n402 66.2847
R3330 vdd.n3446 vdd.n401 66.2847
R3331 vdd.n3446 vdd.n400 66.2847
R3332 vdd.n3446 vdd.n399 66.2847
R3333 vdd.n3446 vdd.n398 66.2847
R3334 vdd.n3446 vdd.n397 66.2847
R3335 vdd.n3446 vdd.n396 66.2847
R3336 vdd.n3446 vdd.n395 66.2847
R3337 vdd.n3446 vdd.n394 66.2847
R3338 vdd.n467 vdd.n394 52.4337
R3339 vdd.n473 vdd.n395 52.4337
R3340 vdd.n477 vdd.n396 52.4337
R3341 vdd.n483 vdd.n397 52.4337
R3342 vdd.n487 vdd.n398 52.4337
R3343 vdd.n493 vdd.n399 52.4337
R3344 vdd.n497 vdd.n400 52.4337
R3345 vdd.n503 vdd.n401 52.4337
R3346 vdd.n507 vdd.n402 52.4337
R3347 vdd.n513 vdd.n403 52.4337
R3348 vdd.n517 vdd.n404 52.4337
R3349 vdd.n523 vdd.n405 52.4337
R3350 vdd.n527 vdd.n406 52.4337
R3351 vdd.n533 vdd.n407 52.4337
R3352 vdd.n537 vdd.n408 52.4337
R3353 vdd.n543 vdd.n409 52.4337
R3354 vdd.n547 vdd.n410 52.4337
R3355 vdd.n553 vdd.n411 52.4337
R3356 vdd.n557 vdd.n412 52.4337
R3357 vdd.n563 vdd.n413 52.4337
R3358 vdd.n567 vdd.n414 52.4337
R3359 vdd.n573 vdd.n415 52.4337
R3360 vdd.n577 vdd.n416 52.4337
R3361 vdd.n583 vdd.n417 52.4337
R3362 vdd.n587 vdd.n418 52.4337
R3363 vdd.n593 vdd.n419 52.4337
R3364 vdd.n597 vdd.n420 52.4337
R3365 vdd.n603 vdd.n421 52.4337
R3366 vdd.n607 vdd.n422 52.4337
R3367 vdd.n613 vdd.n423 52.4337
R3368 vdd.n616 vdd.n424 52.4337
R3369 vdd.n3445 vdd.n3444 52.4337
R3370 vdd.n3314 vdd.n3313 52.4337
R3371 vdd.n728 vdd.n693 52.4337
R3372 vdd.n734 vdd.n694 52.4337
R3373 vdd.n3303 vdd.n695 52.4337
R3374 vdd.n3299 vdd.n696 52.4337
R3375 vdd.n3295 vdd.n697 52.4337
R3376 vdd.n3291 vdd.n698 52.4337
R3377 vdd.n3287 vdd.n699 52.4337
R3378 vdd.n3283 vdd.n700 52.4337
R3379 vdd.n3279 vdd.n701 52.4337
R3380 vdd.n3271 vdd.n702 52.4337
R3381 vdd.n3267 vdd.n703 52.4337
R3382 vdd.n3263 vdd.n704 52.4337
R3383 vdd.n3259 vdd.n705 52.4337
R3384 vdd.n3255 vdd.n706 52.4337
R3385 vdd.n3251 vdd.n707 52.4337
R3386 vdd.n3247 vdd.n708 52.4337
R3387 vdd.n3243 vdd.n709 52.4337
R3388 vdd.n3239 vdd.n710 52.4337
R3389 vdd.n3235 vdd.n711 52.4337
R3390 vdd.n3231 vdd.n712 52.4337
R3391 vdd.n3225 vdd.n713 52.4337
R3392 vdd.n3221 vdd.n714 52.4337
R3393 vdd.n3217 vdd.n715 52.4337
R3394 vdd.n3213 vdd.n716 52.4337
R3395 vdd.n3209 vdd.n717 52.4337
R3396 vdd.n3205 vdd.n718 52.4337
R3397 vdd.n3201 vdd.n719 52.4337
R3398 vdd.n3197 vdd.n720 52.4337
R3399 vdd.n3193 vdd.n721 52.4337
R3400 vdd.n3189 vdd.n722 52.4337
R3401 vdd.n2378 vdd.n1126 52.4337
R3402 vdd.n2376 vdd.n2375 52.4337
R3403 vdd.n2371 vdd.n2370 52.4337
R3404 vdd.n2366 vdd.n1130 52.4337
R3405 vdd.n2364 vdd.n2363 52.4337
R3406 vdd.n2359 vdd.n1137 52.4337
R3407 vdd.n2357 vdd.n2356 52.4337
R3408 vdd.n2352 vdd.n1144 52.4337
R3409 vdd.n2350 vdd.n2349 52.4337
R3410 vdd.n1153 vdd.n1152 52.4337
R3411 vdd.n2341 vdd.n1157 52.4337
R3412 vdd.n2339 vdd.n2338 52.4337
R3413 vdd.n2334 vdd.n1163 52.4337
R3414 vdd.n2332 vdd.n2331 52.4337
R3415 vdd.n2327 vdd.n1170 52.4337
R3416 vdd.n2325 vdd.n2324 52.4337
R3417 vdd.n2320 vdd.n1177 52.4337
R3418 vdd.n2318 vdd.n2317 52.4337
R3419 vdd.n2313 vdd.n1184 52.4337
R3420 vdd.n2311 vdd.n2310 52.4337
R3421 vdd.n1193 vdd.n1192 52.4337
R3422 vdd.n2302 vdd.n1197 52.4337
R3423 vdd.n2300 vdd.n2299 52.4337
R3424 vdd.n2295 vdd.n1203 52.4337
R3425 vdd.n2293 vdd.n2292 52.4337
R3426 vdd.n2288 vdd.n1210 52.4337
R3427 vdd.n2286 vdd.n2285 52.4337
R3428 vdd.n2281 vdd.n1217 52.4337
R3429 vdd.n2279 vdd.n2278 52.4337
R3430 vdd.n1427 vdd.n1426 52.4337
R3431 vdd.n1431 vdd.n1430 52.4337
R3432 vdd.n2267 vdd.n1433 52.4337
R3433 vdd.n1782 vdd.n1781 52.4337
R3434 vdd.n1588 vdd.n1556 52.4337
R3435 vdd.n1592 vdd.n1557 52.4337
R3436 vdd.n1594 vdd.n1558 52.4337
R3437 vdd.n1598 vdd.n1559 52.4337
R3438 vdd.n1600 vdd.n1560 52.4337
R3439 vdd.n1604 vdd.n1561 52.4337
R3440 vdd.n1606 vdd.n1562 52.4337
R3441 vdd.n1610 vdd.n1563 52.4337
R3442 vdd.n1612 vdd.n1564 52.4337
R3443 vdd.n1618 vdd.n1565 52.4337
R3444 vdd.n1620 vdd.n1566 52.4337
R3445 vdd.n1624 vdd.n1567 52.4337
R3446 vdd.n1626 vdd.n1568 52.4337
R3447 vdd.n1630 vdd.n1569 52.4337
R3448 vdd.n1632 vdd.n1570 52.4337
R3449 vdd.n1636 vdd.n1571 52.4337
R3450 vdd.n1638 vdd.n1572 52.4337
R3451 vdd.n1642 vdd.n1573 52.4337
R3452 vdd.n1644 vdd.n1574 52.4337
R3453 vdd.n1716 vdd.n1575 52.4337
R3454 vdd.n1649 vdd.n1576 52.4337
R3455 vdd.n1653 vdd.n1577 52.4337
R3456 vdd.n1655 vdd.n1578 52.4337
R3457 vdd.n1659 vdd.n1579 52.4337
R3458 vdd.n1661 vdd.n1580 52.4337
R3459 vdd.n1665 vdd.n1581 52.4337
R3460 vdd.n1667 vdd.n1582 52.4337
R3461 vdd.n1671 vdd.n1583 52.4337
R3462 vdd.n1673 vdd.n1584 52.4337
R3463 vdd.n1677 vdd.n1585 52.4337
R3464 vdd.n1781 vdd.n1555 52.4337
R3465 vdd.n1591 vdd.n1556 52.4337
R3466 vdd.n1593 vdd.n1557 52.4337
R3467 vdd.n1597 vdd.n1558 52.4337
R3468 vdd.n1599 vdd.n1559 52.4337
R3469 vdd.n1603 vdd.n1560 52.4337
R3470 vdd.n1605 vdd.n1561 52.4337
R3471 vdd.n1609 vdd.n1562 52.4337
R3472 vdd.n1611 vdd.n1563 52.4337
R3473 vdd.n1617 vdd.n1564 52.4337
R3474 vdd.n1619 vdd.n1565 52.4337
R3475 vdd.n1623 vdd.n1566 52.4337
R3476 vdd.n1625 vdd.n1567 52.4337
R3477 vdd.n1629 vdd.n1568 52.4337
R3478 vdd.n1631 vdd.n1569 52.4337
R3479 vdd.n1635 vdd.n1570 52.4337
R3480 vdd.n1637 vdd.n1571 52.4337
R3481 vdd.n1641 vdd.n1572 52.4337
R3482 vdd.n1643 vdd.n1573 52.4337
R3483 vdd.n1647 vdd.n1574 52.4337
R3484 vdd.n1648 vdd.n1575 52.4337
R3485 vdd.n1652 vdd.n1576 52.4337
R3486 vdd.n1654 vdd.n1577 52.4337
R3487 vdd.n1658 vdd.n1578 52.4337
R3488 vdd.n1660 vdd.n1579 52.4337
R3489 vdd.n1664 vdd.n1580 52.4337
R3490 vdd.n1666 vdd.n1581 52.4337
R3491 vdd.n1670 vdd.n1582 52.4337
R3492 vdd.n1672 vdd.n1583 52.4337
R3493 vdd.n1676 vdd.n1584 52.4337
R3494 vdd.n1678 vdd.n1585 52.4337
R3495 vdd.n1433 vdd.n1432 52.4337
R3496 vdd.n1430 vdd.n1429 52.4337
R3497 vdd.n1426 vdd.n1218 52.4337
R3498 vdd.n2280 vdd.n2279 52.4337
R3499 vdd.n1217 vdd.n1211 52.4337
R3500 vdd.n2287 vdd.n2286 52.4337
R3501 vdd.n1210 vdd.n1204 52.4337
R3502 vdd.n2294 vdd.n2293 52.4337
R3503 vdd.n1203 vdd.n1198 52.4337
R3504 vdd.n2301 vdd.n2300 52.4337
R3505 vdd.n1197 vdd.n1196 52.4337
R3506 vdd.n1192 vdd.n1185 52.4337
R3507 vdd.n2312 vdd.n2311 52.4337
R3508 vdd.n1184 vdd.n1178 52.4337
R3509 vdd.n2319 vdd.n2318 52.4337
R3510 vdd.n1177 vdd.n1171 52.4337
R3511 vdd.n2326 vdd.n2325 52.4337
R3512 vdd.n1170 vdd.n1164 52.4337
R3513 vdd.n2333 vdd.n2332 52.4337
R3514 vdd.n1163 vdd.n1158 52.4337
R3515 vdd.n2340 vdd.n2339 52.4337
R3516 vdd.n1157 vdd.n1156 52.4337
R3517 vdd.n1152 vdd.n1145 52.4337
R3518 vdd.n2351 vdd.n2350 52.4337
R3519 vdd.n1144 vdd.n1138 52.4337
R3520 vdd.n2358 vdd.n2357 52.4337
R3521 vdd.n1137 vdd.n1131 52.4337
R3522 vdd.n2365 vdd.n2364 52.4337
R3523 vdd.n1130 vdd.n1127 52.4337
R3524 vdd.n2372 vdd.n2371 52.4337
R3525 vdd.n2377 vdd.n2376 52.4337
R3526 vdd.n1437 vdd.n1126 52.4337
R3527 vdd.n3314 vdd.n725 52.4337
R3528 vdd.n733 vdd.n693 52.4337
R3529 vdd.n3304 vdd.n694 52.4337
R3530 vdd.n3300 vdd.n695 52.4337
R3531 vdd.n3296 vdd.n696 52.4337
R3532 vdd.n3292 vdd.n697 52.4337
R3533 vdd.n3288 vdd.n698 52.4337
R3534 vdd.n3284 vdd.n699 52.4337
R3535 vdd.n3280 vdd.n700 52.4337
R3536 vdd.n3270 vdd.n701 52.4337
R3537 vdd.n3268 vdd.n702 52.4337
R3538 vdd.n3264 vdd.n703 52.4337
R3539 vdd.n3260 vdd.n704 52.4337
R3540 vdd.n3256 vdd.n705 52.4337
R3541 vdd.n3252 vdd.n706 52.4337
R3542 vdd.n3248 vdd.n707 52.4337
R3543 vdd.n3244 vdd.n708 52.4337
R3544 vdd.n3240 vdd.n709 52.4337
R3545 vdd.n3236 vdd.n710 52.4337
R3546 vdd.n3232 vdd.n711 52.4337
R3547 vdd.n3224 vdd.n712 52.4337
R3548 vdd.n3222 vdd.n713 52.4337
R3549 vdd.n3218 vdd.n714 52.4337
R3550 vdd.n3214 vdd.n715 52.4337
R3551 vdd.n3210 vdd.n716 52.4337
R3552 vdd.n3206 vdd.n717 52.4337
R3553 vdd.n3202 vdd.n718 52.4337
R3554 vdd.n3198 vdd.n719 52.4337
R3555 vdd.n3194 vdd.n720 52.4337
R3556 vdd.n3190 vdd.n721 52.4337
R3557 vdd.n722 vdd.n691 52.4337
R3558 vdd.n3445 vdd.n425 52.4337
R3559 vdd.n614 vdd.n424 52.4337
R3560 vdd.n608 vdd.n423 52.4337
R3561 vdd.n604 vdd.n422 52.4337
R3562 vdd.n598 vdd.n421 52.4337
R3563 vdd.n594 vdd.n420 52.4337
R3564 vdd.n588 vdd.n419 52.4337
R3565 vdd.n584 vdd.n418 52.4337
R3566 vdd.n578 vdd.n417 52.4337
R3567 vdd.n574 vdd.n416 52.4337
R3568 vdd.n568 vdd.n415 52.4337
R3569 vdd.n564 vdd.n414 52.4337
R3570 vdd.n558 vdd.n413 52.4337
R3571 vdd.n554 vdd.n412 52.4337
R3572 vdd.n548 vdd.n411 52.4337
R3573 vdd.n544 vdd.n410 52.4337
R3574 vdd.n538 vdd.n409 52.4337
R3575 vdd.n534 vdd.n408 52.4337
R3576 vdd.n528 vdd.n407 52.4337
R3577 vdd.n524 vdd.n406 52.4337
R3578 vdd.n518 vdd.n405 52.4337
R3579 vdd.n514 vdd.n404 52.4337
R3580 vdd.n508 vdd.n403 52.4337
R3581 vdd.n504 vdd.n402 52.4337
R3582 vdd.n498 vdd.n401 52.4337
R3583 vdd.n494 vdd.n400 52.4337
R3584 vdd.n488 vdd.n399 52.4337
R3585 vdd.n484 vdd.n398 52.4337
R3586 vdd.n478 vdd.n397 52.4337
R3587 vdd.n474 vdd.n396 52.4337
R3588 vdd.n468 vdd.n395 52.4337
R3589 vdd.n394 vdd.n392 52.4337
R3590 vdd.t46 vdd.t10 51.4683
R3591 vdd.n274 vdd.n272 42.0461
R3592 vdd.n172 vdd.n170 42.0461
R3593 vdd.n71 vdd.n69 42.0461
R3594 vdd.n2114 vdd.n2112 42.0461
R3595 vdd.n2012 vdd.n2010 42.0461
R3596 vdd.n1911 vdd.n1909 42.0461
R3597 vdd.n332 vdd.n331 41.6884
R3598 vdd.n230 vdd.n229 41.6884
R3599 vdd.n129 vdd.n128 41.6884
R3600 vdd.n2172 vdd.n2171 41.6884
R3601 vdd.n2070 vdd.n2069 41.6884
R3602 vdd.n1969 vdd.n1968 41.6884
R3603 vdd.n1681 vdd.n1680 41.1157
R3604 vdd.n1719 vdd.n1718 41.1157
R3605 vdd.n1615 vdd.n1614 41.1157
R3606 vdd.n428 vdd.n427 41.1157
R3607 vdd.n566 vdd.n441 41.1157
R3608 vdd.n454 vdd.n453 41.1157
R3609 vdd.n3145 vdd.n3144 39.2114
R3610 vdd.n3142 vdd.n3141 39.2114
R3611 vdd.n3137 vdd.n815 39.2114
R3612 vdd.n3135 vdd.n3134 39.2114
R3613 vdd.n3130 vdd.n818 39.2114
R3614 vdd.n3128 vdd.n3127 39.2114
R3615 vdd.n3123 vdd.n821 39.2114
R3616 vdd.n3121 vdd.n3120 39.2114
R3617 vdd.n3117 vdd.n3116 39.2114
R3618 vdd.n3112 vdd.n824 39.2114
R3619 vdd.n3110 vdd.n3109 39.2114
R3620 vdd.n3105 vdd.n827 39.2114
R3621 vdd.n3103 vdd.n3102 39.2114
R3622 vdd.n3098 vdd.n830 39.2114
R3623 vdd.n3096 vdd.n3095 39.2114
R3624 vdd.n3090 vdd.n835 39.2114
R3625 vdd.n3088 vdd.n3087 39.2114
R3626 vdd.n2937 vdd.n2936 39.2114
R3627 vdd.n2931 vdd.n2666 39.2114
R3628 vdd.n2928 vdd.n2667 39.2114
R3629 vdd.n2924 vdd.n2668 39.2114
R3630 vdd.n2920 vdd.n2669 39.2114
R3631 vdd.n2916 vdd.n2670 39.2114
R3632 vdd.n2912 vdd.n2671 39.2114
R3633 vdd.n2908 vdd.n2672 39.2114
R3634 vdd.n2904 vdd.n2673 39.2114
R3635 vdd.n2900 vdd.n2674 39.2114
R3636 vdd.n2896 vdd.n2675 39.2114
R3637 vdd.n2892 vdd.n2676 39.2114
R3638 vdd.n2888 vdd.n2677 39.2114
R3639 vdd.n2884 vdd.n2678 39.2114
R3640 vdd.n2880 vdd.n2679 39.2114
R3641 vdd.n2876 vdd.n2680 39.2114
R3642 vdd.n2871 vdd.n2681 39.2114
R3643 vdd.n2660 vdd.n968 39.2114
R3644 vdd.n2656 vdd.n967 39.2114
R3645 vdd.n2652 vdd.n966 39.2114
R3646 vdd.n2648 vdd.n965 39.2114
R3647 vdd.n2644 vdd.n964 39.2114
R3648 vdd.n2640 vdd.n963 39.2114
R3649 vdd.n2636 vdd.n962 39.2114
R3650 vdd.n2632 vdd.n961 39.2114
R3651 vdd.n2628 vdd.n960 39.2114
R3652 vdd.n2624 vdd.n959 39.2114
R3653 vdd.n2620 vdd.n958 39.2114
R3654 vdd.n2616 vdd.n957 39.2114
R3655 vdd.n2612 vdd.n956 39.2114
R3656 vdd.n2608 vdd.n955 39.2114
R3657 vdd.n2604 vdd.n954 39.2114
R3658 vdd.n2599 vdd.n953 39.2114
R3659 vdd.n2595 vdd.n952 39.2114
R3660 vdd.n2416 vdd.n2415 39.2114
R3661 vdd.n2410 vdd.n1084 39.2114
R3662 vdd.n2407 vdd.n1085 39.2114
R3663 vdd.n2403 vdd.n1086 39.2114
R3664 vdd.n2399 vdd.n1087 39.2114
R3665 vdd.n2395 vdd.n1088 39.2114
R3666 vdd.n2391 vdd.n1089 39.2114
R3667 vdd.n2387 vdd.n1090 39.2114
R3668 vdd.n2383 vdd.n1091 39.2114
R3669 vdd.n1276 vdd.n1092 39.2114
R3670 vdd.n1280 vdd.n1093 39.2114
R3671 vdd.n1284 vdd.n1094 39.2114
R3672 vdd.n1288 vdd.n1095 39.2114
R3673 vdd.n1292 vdd.n1096 39.2114
R3674 vdd.n1296 vdd.n1097 39.2114
R3675 vdd.n1300 vdd.n1098 39.2114
R3676 vdd.n1305 vdd.n1099 39.2114
R3677 vdd.n3064 vdd.n3063 39.2114
R3678 vdd.n3059 vdd.n3031 39.2114
R3679 vdd.n3057 vdd.n3056 39.2114
R3680 vdd.n3052 vdd.n3034 39.2114
R3681 vdd.n3050 vdd.n3049 39.2114
R3682 vdd.n3045 vdd.n3037 39.2114
R3683 vdd.n3043 vdd.n3042 39.2114
R3684 vdd.n3038 vdd.n787 39.2114
R3685 vdd.n3182 vdd.n3181 39.2114
R3686 vdd.n3179 vdd.n3178 39.2114
R3687 vdd.n3174 vdd.n791 39.2114
R3688 vdd.n3172 vdd.n3171 39.2114
R3689 vdd.n3167 vdd.n794 39.2114
R3690 vdd.n3165 vdd.n3164 39.2114
R3691 vdd.n3160 vdd.n797 39.2114
R3692 vdd.n3158 vdd.n3157 39.2114
R3693 vdd.n3153 vdd.n803 39.2114
R3694 vdd.n2940 vdd.n2939 39.2114
R3695 vdd.n2707 vdd.n2682 39.2114
R3696 vdd.n2711 vdd.n2683 39.2114
R3697 vdd.n2715 vdd.n2684 39.2114
R3698 vdd.n2719 vdd.n2685 39.2114
R3699 vdd.n2723 vdd.n2686 39.2114
R3700 vdd.n2727 vdd.n2687 39.2114
R3701 vdd.n2731 vdd.n2688 39.2114
R3702 vdd.n2735 vdd.n2689 39.2114
R3703 vdd.n2739 vdd.n2690 39.2114
R3704 vdd.n2743 vdd.n2691 39.2114
R3705 vdd.n2747 vdd.n2692 39.2114
R3706 vdd.n2751 vdd.n2693 39.2114
R3707 vdd.n2755 vdd.n2694 39.2114
R3708 vdd.n2759 vdd.n2695 39.2114
R3709 vdd.n2763 vdd.n2696 39.2114
R3710 vdd.n2767 vdd.n2697 39.2114
R3711 vdd.n2939 vdd.n933 39.2114
R3712 vdd.n2710 vdd.n2682 39.2114
R3713 vdd.n2714 vdd.n2683 39.2114
R3714 vdd.n2718 vdd.n2684 39.2114
R3715 vdd.n2722 vdd.n2685 39.2114
R3716 vdd.n2726 vdd.n2686 39.2114
R3717 vdd.n2730 vdd.n2687 39.2114
R3718 vdd.n2734 vdd.n2688 39.2114
R3719 vdd.n2738 vdd.n2689 39.2114
R3720 vdd.n2742 vdd.n2690 39.2114
R3721 vdd.n2746 vdd.n2691 39.2114
R3722 vdd.n2750 vdd.n2692 39.2114
R3723 vdd.n2754 vdd.n2693 39.2114
R3724 vdd.n2758 vdd.n2694 39.2114
R3725 vdd.n2762 vdd.n2695 39.2114
R3726 vdd.n2766 vdd.n2696 39.2114
R3727 vdd.n2769 vdd.n2697 39.2114
R3728 vdd.n803 vdd.n798 39.2114
R3729 vdd.n3159 vdd.n3158 39.2114
R3730 vdd.n797 vdd.n795 39.2114
R3731 vdd.n3166 vdd.n3165 39.2114
R3732 vdd.n794 vdd.n792 39.2114
R3733 vdd.n3173 vdd.n3172 39.2114
R3734 vdd.n791 vdd.n789 39.2114
R3735 vdd.n3180 vdd.n3179 39.2114
R3736 vdd.n3183 vdd.n3182 39.2114
R3737 vdd.n3039 vdd.n3038 39.2114
R3738 vdd.n3044 vdd.n3043 39.2114
R3739 vdd.n3037 vdd.n3035 39.2114
R3740 vdd.n3051 vdd.n3050 39.2114
R3741 vdd.n3034 vdd.n3032 39.2114
R3742 vdd.n3058 vdd.n3057 39.2114
R3743 vdd.n3031 vdd.n3029 39.2114
R3744 vdd.n3065 vdd.n3064 39.2114
R3745 vdd.n2416 vdd.n1118 39.2114
R3746 vdd.n2408 vdd.n1084 39.2114
R3747 vdd.n2404 vdd.n1085 39.2114
R3748 vdd.n2400 vdd.n1086 39.2114
R3749 vdd.n2396 vdd.n1087 39.2114
R3750 vdd.n2392 vdd.n1088 39.2114
R3751 vdd.n2388 vdd.n1089 39.2114
R3752 vdd.n2384 vdd.n1090 39.2114
R3753 vdd.n1275 vdd.n1091 39.2114
R3754 vdd.n1279 vdd.n1092 39.2114
R3755 vdd.n1283 vdd.n1093 39.2114
R3756 vdd.n1287 vdd.n1094 39.2114
R3757 vdd.n1291 vdd.n1095 39.2114
R3758 vdd.n1295 vdd.n1096 39.2114
R3759 vdd.n1299 vdd.n1097 39.2114
R3760 vdd.n1304 vdd.n1098 39.2114
R3761 vdd.n1308 vdd.n1099 39.2114
R3762 vdd.n2598 vdd.n952 39.2114
R3763 vdd.n2603 vdd.n953 39.2114
R3764 vdd.n2607 vdd.n954 39.2114
R3765 vdd.n2611 vdd.n955 39.2114
R3766 vdd.n2615 vdd.n956 39.2114
R3767 vdd.n2619 vdd.n957 39.2114
R3768 vdd.n2623 vdd.n958 39.2114
R3769 vdd.n2627 vdd.n959 39.2114
R3770 vdd.n2631 vdd.n960 39.2114
R3771 vdd.n2635 vdd.n961 39.2114
R3772 vdd.n2639 vdd.n962 39.2114
R3773 vdd.n2643 vdd.n963 39.2114
R3774 vdd.n2647 vdd.n964 39.2114
R3775 vdd.n2651 vdd.n965 39.2114
R3776 vdd.n2655 vdd.n966 39.2114
R3777 vdd.n2659 vdd.n967 39.2114
R3778 vdd.n970 vdd.n968 39.2114
R3779 vdd.n2937 vdd.n2700 39.2114
R3780 vdd.n2929 vdd.n2666 39.2114
R3781 vdd.n2925 vdd.n2667 39.2114
R3782 vdd.n2921 vdd.n2668 39.2114
R3783 vdd.n2917 vdd.n2669 39.2114
R3784 vdd.n2913 vdd.n2670 39.2114
R3785 vdd.n2909 vdd.n2671 39.2114
R3786 vdd.n2905 vdd.n2672 39.2114
R3787 vdd.n2901 vdd.n2673 39.2114
R3788 vdd.n2897 vdd.n2674 39.2114
R3789 vdd.n2893 vdd.n2675 39.2114
R3790 vdd.n2889 vdd.n2676 39.2114
R3791 vdd.n2885 vdd.n2677 39.2114
R3792 vdd.n2881 vdd.n2678 39.2114
R3793 vdd.n2877 vdd.n2679 39.2114
R3794 vdd.n2872 vdd.n2680 39.2114
R3795 vdd.n2868 vdd.n2681 39.2114
R3796 vdd.n3089 vdd.n3088 39.2114
R3797 vdd.n835 vdd.n831 39.2114
R3798 vdd.n3097 vdd.n3096 39.2114
R3799 vdd.n830 vdd.n828 39.2114
R3800 vdd.n3104 vdd.n3103 39.2114
R3801 vdd.n827 vdd.n825 39.2114
R3802 vdd.n3111 vdd.n3110 39.2114
R3803 vdd.n824 vdd.n822 39.2114
R3804 vdd.n3118 vdd.n3117 39.2114
R3805 vdd.n3122 vdd.n3121 39.2114
R3806 vdd.n821 vdd.n819 39.2114
R3807 vdd.n3129 vdd.n3128 39.2114
R3808 vdd.n818 vdd.n816 39.2114
R3809 vdd.n3136 vdd.n3135 39.2114
R3810 vdd.n815 vdd.n813 39.2114
R3811 vdd.n3143 vdd.n3142 39.2114
R3812 vdd.n3146 vdd.n3145 39.2114
R3813 vdd.n979 vdd.n934 39.2114
R3814 vdd.n2587 vdd.n935 39.2114
R3815 vdd.n2583 vdd.n936 39.2114
R3816 vdd.n2579 vdd.n937 39.2114
R3817 vdd.n2575 vdd.n938 39.2114
R3818 vdd.n2571 vdd.n939 39.2114
R3819 vdd.n2567 vdd.n940 39.2114
R3820 vdd.n2563 vdd.n941 39.2114
R3821 vdd.n2559 vdd.n942 39.2114
R3822 vdd.n2555 vdd.n943 39.2114
R3823 vdd.n2551 vdd.n944 39.2114
R3824 vdd.n2547 vdd.n945 39.2114
R3825 vdd.n2543 vdd.n946 39.2114
R3826 vdd.n2539 vdd.n947 39.2114
R3827 vdd.n2535 vdd.n948 39.2114
R3828 vdd.n2531 vdd.n949 39.2114
R3829 vdd.n2527 vdd.n950 39.2114
R3830 vdd.n2419 vdd.n2418 39.2114
R3831 vdd.n1222 vdd.n1100 39.2114
R3832 vdd.n1226 vdd.n1101 39.2114
R3833 vdd.n1230 vdd.n1102 39.2114
R3834 vdd.n1234 vdd.n1103 39.2114
R3835 vdd.n1238 vdd.n1104 39.2114
R3836 vdd.n1242 vdd.n1105 39.2114
R3837 vdd.n1246 vdd.n1106 39.2114
R3838 vdd.n1250 vdd.n1107 39.2114
R3839 vdd.n1420 vdd.n1108 39.2114
R3840 vdd.n1417 vdd.n1109 39.2114
R3841 vdd.n1413 vdd.n1110 39.2114
R3842 vdd.n1409 vdd.n1111 39.2114
R3843 vdd.n1405 vdd.n1112 39.2114
R3844 vdd.n1401 vdd.n1113 39.2114
R3845 vdd.n1397 vdd.n1114 39.2114
R3846 vdd.n1393 vdd.n1115 39.2114
R3847 vdd.n2524 vdd.n950 39.2114
R3848 vdd.n2528 vdd.n949 39.2114
R3849 vdd.n2532 vdd.n948 39.2114
R3850 vdd.n2536 vdd.n947 39.2114
R3851 vdd.n2540 vdd.n946 39.2114
R3852 vdd.n2544 vdd.n945 39.2114
R3853 vdd.n2548 vdd.n944 39.2114
R3854 vdd.n2552 vdd.n943 39.2114
R3855 vdd.n2556 vdd.n942 39.2114
R3856 vdd.n2560 vdd.n941 39.2114
R3857 vdd.n2564 vdd.n940 39.2114
R3858 vdd.n2568 vdd.n939 39.2114
R3859 vdd.n2572 vdd.n938 39.2114
R3860 vdd.n2576 vdd.n937 39.2114
R3861 vdd.n2580 vdd.n936 39.2114
R3862 vdd.n2584 vdd.n935 39.2114
R3863 vdd.n2588 vdd.n934 39.2114
R3864 vdd.n2418 vdd.n1082 39.2114
R3865 vdd.n1225 vdd.n1100 39.2114
R3866 vdd.n1229 vdd.n1101 39.2114
R3867 vdd.n1233 vdd.n1102 39.2114
R3868 vdd.n1237 vdd.n1103 39.2114
R3869 vdd.n1241 vdd.n1104 39.2114
R3870 vdd.n1245 vdd.n1105 39.2114
R3871 vdd.n1249 vdd.n1106 39.2114
R3872 vdd.n1252 vdd.n1107 39.2114
R3873 vdd.n1418 vdd.n1108 39.2114
R3874 vdd.n1414 vdd.n1109 39.2114
R3875 vdd.n1410 vdd.n1110 39.2114
R3876 vdd.n1406 vdd.n1111 39.2114
R3877 vdd.n1402 vdd.n1112 39.2114
R3878 vdd.n1398 vdd.n1113 39.2114
R3879 vdd.n1394 vdd.n1114 39.2114
R3880 vdd.n1390 vdd.n1115 39.2114
R3881 vdd.n2271 vdd.n2270 37.2369
R3882 vdd.n2307 vdd.n1191 37.2369
R3883 vdd.n2346 vdd.n1151 37.2369
R3884 vdd.n3230 vdd.n769 37.2369
R3885 vdd.n3278 vdd.n3277 37.2369
R3886 vdd.n690 vdd.n689 37.2369
R3887 vdd.n2414 vdd.n1074 31.0639
R3888 vdd.n2663 vdd.n971 31.0639
R3889 vdd.n2596 vdd.n974 31.0639
R3890 vdd.n1310 vdd.n1307 31.0639
R3891 vdd.n2869 vdd.n2866 31.0639
R3892 vdd.n3086 vdd.n3085 31.0639
R3893 vdd.n2935 vdd.n926 31.0639
R3894 vdd.n3149 vdd.n3148 31.0639
R3895 vdd.n3068 vdd.n3067 31.0639
R3896 vdd.n3154 vdd.n802 31.0639
R3897 vdd.n2773 vdd.n2771 31.0639
R3898 vdd.n2942 vdd.n2941 31.0639
R3899 vdd.n2421 vdd.n2420 31.0639
R3900 vdd.n2591 vdd.n2590 31.0639
R3901 vdd.n2523 vdd.n2522 31.0639
R3902 vdd.n1389 vdd.n1388 31.0639
R3903 vdd.n1255 vdd.n1254 30.449
R3904 vdd.n983 vdd.n982 30.449
R3905 vdd.n1302 vdd.n1274 30.449
R3906 vdd.n2601 vdd.n973 30.449
R3907 vdd.n2706 vdd.n2705 30.449
R3908 vdd.n3092 vdd.n833 30.449
R3909 vdd.n2874 vdd.n2702 30.449
R3910 vdd.n801 vdd.n800 30.449
R3911 vdd.n1780 vdd.n1587 22.2201
R3912 vdd.n2265 vdd.n1083 22.2201
R3913 vdd.n3315 vdd.n723 22.2201
R3914 vdd.n3447 vdd.n3446 22.2201
R3915 vdd.n1791 vdd.n1549 19.3944
R3916 vdd.n1791 vdd.n1547 19.3944
R3917 vdd.n1795 vdd.n1547 19.3944
R3918 vdd.n1795 vdd.n1537 19.3944
R3919 vdd.n1808 vdd.n1537 19.3944
R3920 vdd.n1808 vdd.n1535 19.3944
R3921 vdd.n1812 vdd.n1535 19.3944
R3922 vdd.n1812 vdd.n1527 19.3944
R3923 vdd.n1825 vdd.n1527 19.3944
R3924 vdd.n1825 vdd.n1525 19.3944
R3925 vdd.n1829 vdd.n1525 19.3944
R3926 vdd.n1829 vdd.n1514 19.3944
R3927 vdd.n1841 vdd.n1514 19.3944
R3928 vdd.n1841 vdd.n1512 19.3944
R3929 vdd.n1845 vdd.n1512 19.3944
R3930 vdd.n1845 vdd.n1503 19.3944
R3931 vdd.n1858 vdd.n1503 19.3944
R3932 vdd.n1858 vdd.n1501 19.3944
R3933 vdd.n1862 vdd.n1501 19.3944
R3934 vdd.n1862 vdd.n1492 19.3944
R3935 vdd.n2181 vdd.n1492 19.3944
R3936 vdd.n2181 vdd.n1490 19.3944
R3937 vdd.n2185 vdd.n1490 19.3944
R3938 vdd.n2185 vdd.n1480 19.3944
R3939 vdd.n2198 vdd.n1480 19.3944
R3940 vdd.n2198 vdd.n1478 19.3944
R3941 vdd.n2202 vdd.n1478 19.3944
R3942 vdd.n2202 vdd.n1470 19.3944
R3943 vdd.n2215 vdd.n1470 19.3944
R3944 vdd.n2215 vdd.n1468 19.3944
R3945 vdd.n2219 vdd.n1468 19.3944
R3946 vdd.n2219 vdd.n1457 19.3944
R3947 vdd.n2231 vdd.n1457 19.3944
R3948 vdd.n2231 vdd.n1455 19.3944
R3949 vdd.n2235 vdd.n1455 19.3944
R3950 vdd.n2235 vdd.n1447 19.3944
R3951 vdd.n2248 vdd.n1447 19.3944
R3952 vdd.n2248 vdd.n1444 19.3944
R3953 vdd.n2254 vdd.n1444 19.3944
R3954 vdd.n2254 vdd.n1445 19.3944
R3955 vdd.n1445 vdd.n1435 19.3944
R3956 vdd.n1715 vdd.n1650 19.3944
R3957 vdd.n1711 vdd.n1650 19.3944
R3958 vdd.n1711 vdd.n1710 19.3944
R3959 vdd.n1710 vdd.n1709 19.3944
R3960 vdd.n1709 vdd.n1656 19.3944
R3961 vdd.n1705 vdd.n1656 19.3944
R3962 vdd.n1705 vdd.n1704 19.3944
R3963 vdd.n1704 vdd.n1703 19.3944
R3964 vdd.n1703 vdd.n1662 19.3944
R3965 vdd.n1699 vdd.n1662 19.3944
R3966 vdd.n1699 vdd.n1698 19.3944
R3967 vdd.n1698 vdd.n1697 19.3944
R3968 vdd.n1697 vdd.n1668 19.3944
R3969 vdd.n1693 vdd.n1668 19.3944
R3970 vdd.n1693 vdd.n1692 19.3944
R3971 vdd.n1692 vdd.n1691 19.3944
R3972 vdd.n1691 vdd.n1674 19.3944
R3973 vdd.n1687 vdd.n1674 19.3944
R3974 vdd.n1687 vdd.n1686 19.3944
R3975 vdd.n1686 vdd.n1685 19.3944
R3976 vdd.n1750 vdd.n1749 19.3944
R3977 vdd.n1749 vdd.n1748 19.3944
R3978 vdd.n1748 vdd.n1621 19.3944
R3979 vdd.n1744 vdd.n1621 19.3944
R3980 vdd.n1744 vdd.n1743 19.3944
R3981 vdd.n1743 vdd.n1742 19.3944
R3982 vdd.n1742 vdd.n1627 19.3944
R3983 vdd.n1738 vdd.n1627 19.3944
R3984 vdd.n1738 vdd.n1737 19.3944
R3985 vdd.n1737 vdd.n1736 19.3944
R3986 vdd.n1736 vdd.n1633 19.3944
R3987 vdd.n1732 vdd.n1633 19.3944
R3988 vdd.n1732 vdd.n1731 19.3944
R3989 vdd.n1731 vdd.n1730 19.3944
R3990 vdd.n1730 vdd.n1639 19.3944
R3991 vdd.n1726 vdd.n1639 19.3944
R3992 vdd.n1726 vdd.n1725 19.3944
R3993 vdd.n1725 vdd.n1724 19.3944
R3994 vdd.n1724 vdd.n1645 19.3944
R3995 vdd.n1720 vdd.n1645 19.3944
R3996 vdd.n1783 vdd.n1554 19.3944
R3997 vdd.n1778 vdd.n1554 19.3944
R3998 vdd.n1778 vdd.n1589 19.3944
R3999 vdd.n1774 vdd.n1589 19.3944
R4000 vdd.n1774 vdd.n1773 19.3944
R4001 vdd.n1773 vdd.n1772 19.3944
R4002 vdd.n1772 vdd.n1595 19.3944
R4003 vdd.n1768 vdd.n1595 19.3944
R4004 vdd.n1768 vdd.n1767 19.3944
R4005 vdd.n1767 vdd.n1766 19.3944
R4006 vdd.n1766 vdd.n1601 19.3944
R4007 vdd.n1762 vdd.n1601 19.3944
R4008 vdd.n1762 vdd.n1761 19.3944
R4009 vdd.n1761 vdd.n1760 19.3944
R4010 vdd.n1760 vdd.n1607 19.3944
R4011 vdd.n1756 vdd.n1607 19.3944
R4012 vdd.n1756 vdd.n1755 19.3944
R4013 vdd.n1755 vdd.n1754 19.3944
R4014 vdd.n2303 vdd.n1189 19.3944
R4015 vdd.n2303 vdd.n1195 19.3944
R4016 vdd.n2298 vdd.n1195 19.3944
R4017 vdd.n2298 vdd.n2297 19.3944
R4018 vdd.n2297 vdd.n2296 19.3944
R4019 vdd.n2296 vdd.n1202 19.3944
R4020 vdd.n2291 vdd.n1202 19.3944
R4021 vdd.n2291 vdd.n2290 19.3944
R4022 vdd.n2290 vdd.n2289 19.3944
R4023 vdd.n2289 vdd.n1209 19.3944
R4024 vdd.n2284 vdd.n1209 19.3944
R4025 vdd.n2284 vdd.n2283 19.3944
R4026 vdd.n2283 vdd.n2282 19.3944
R4027 vdd.n2282 vdd.n1216 19.3944
R4028 vdd.n2277 vdd.n1216 19.3944
R4029 vdd.n2277 vdd.n2276 19.3944
R4030 vdd.n1428 vdd.n1221 19.3944
R4031 vdd.n2272 vdd.n1425 19.3944
R4032 vdd.n2342 vdd.n1149 19.3944
R4033 vdd.n2342 vdd.n1155 19.3944
R4034 vdd.n2337 vdd.n1155 19.3944
R4035 vdd.n2337 vdd.n2336 19.3944
R4036 vdd.n2336 vdd.n2335 19.3944
R4037 vdd.n2335 vdd.n1162 19.3944
R4038 vdd.n2330 vdd.n1162 19.3944
R4039 vdd.n2330 vdd.n2329 19.3944
R4040 vdd.n2329 vdd.n2328 19.3944
R4041 vdd.n2328 vdd.n1169 19.3944
R4042 vdd.n2323 vdd.n1169 19.3944
R4043 vdd.n2323 vdd.n2322 19.3944
R4044 vdd.n2322 vdd.n2321 19.3944
R4045 vdd.n2321 vdd.n1176 19.3944
R4046 vdd.n2316 vdd.n1176 19.3944
R4047 vdd.n2316 vdd.n2315 19.3944
R4048 vdd.n2315 vdd.n2314 19.3944
R4049 vdd.n2314 vdd.n1183 19.3944
R4050 vdd.n2309 vdd.n1183 19.3944
R4051 vdd.n2309 vdd.n2308 19.3944
R4052 vdd.n2379 vdd.n1124 19.3944
R4053 vdd.n2379 vdd.n1125 19.3944
R4054 vdd.n2374 vdd.n2373 19.3944
R4055 vdd.n2369 vdd.n2368 19.3944
R4056 vdd.n2368 vdd.n2367 19.3944
R4057 vdd.n2367 vdd.n1129 19.3944
R4058 vdd.n2362 vdd.n1129 19.3944
R4059 vdd.n2362 vdd.n2361 19.3944
R4060 vdd.n2361 vdd.n2360 19.3944
R4061 vdd.n2360 vdd.n1136 19.3944
R4062 vdd.n2355 vdd.n1136 19.3944
R4063 vdd.n2355 vdd.n2354 19.3944
R4064 vdd.n2354 vdd.n2353 19.3944
R4065 vdd.n2353 vdd.n1143 19.3944
R4066 vdd.n2348 vdd.n1143 19.3944
R4067 vdd.n2348 vdd.n2347 19.3944
R4068 vdd.n1787 vdd.n1552 19.3944
R4069 vdd.n1787 vdd.n1543 19.3944
R4070 vdd.n1800 vdd.n1543 19.3944
R4071 vdd.n1800 vdd.n1541 19.3944
R4072 vdd.n1804 vdd.n1541 19.3944
R4073 vdd.n1804 vdd.n1532 19.3944
R4074 vdd.n1817 vdd.n1532 19.3944
R4075 vdd.n1817 vdd.n1530 19.3944
R4076 vdd.n1821 vdd.n1530 19.3944
R4077 vdd.n1821 vdd.n1521 19.3944
R4078 vdd.n1833 vdd.n1521 19.3944
R4079 vdd.n1833 vdd.n1519 19.3944
R4080 vdd.n1837 vdd.n1519 19.3944
R4081 vdd.n1837 vdd.n1509 19.3944
R4082 vdd.n1850 vdd.n1509 19.3944
R4083 vdd.n1850 vdd.n1507 19.3944
R4084 vdd.n1854 vdd.n1507 19.3944
R4085 vdd.n1854 vdd.n1498 19.3944
R4086 vdd.n1866 vdd.n1498 19.3944
R4087 vdd.n1866 vdd.n1496 19.3944
R4088 vdd.n2177 vdd.n1496 19.3944
R4089 vdd.n2177 vdd.n1486 19.3944
R4090 vdd.n2190 vdd.n1486 19.3944
R4091 vdd.n2190 vdd.n1484 19.3944
R4092 vdd.n2194 vdd.n1484 19.3944
R4093 vdd.n2194 vdd.n1475 19.3944
R4094 vdd.n2207 vdd.n1475 19.3944
R4095 vdd.n2207 vdd.n1473 19.3944
R4096 vdd.n2211 vdd.n1473 19.3944
R4097 vdd.n2211 vdd.n1464 19.3944
R4098 vdd.n2223 vdd.n1464 19.3944
R4099 vdd.n2223 vdd.n1462 19.3944
R4100 vdd.n2227 vdd.n1462 19.3944
R4101 vdd.n2227 vdd.n1452 19.3944
R4102 vdd.n2240 vdd.n1452 19.3944
R4103 vdd.n2240 vdd.n1450 19.3944
R4104 vdd.n2244 vdd.n1450 19.3944
R4105 vdd.n2244 vdd.n1440 19.3944
R4106 vdd.n2259 vdd.n1440 19.3944
R4107 vdd.n2259 vdd.n1438 19.3944
R4108 vdd.n2263 vdd.n1438 19.3944
R4109 vdd.n3321 vdd.n686 19.3944
R4110 vdd.n3321 vdd.n676 19.3944
R4111 vdd.n3333 vdd.n676 19.3944
R4112 vdd.n3333 vdd.n674 19.3944
R4113 vdd.n3337 vdd.n674 19.3944
R4114 vdd.n3337 vdd.n666 19.3944
R4115 vdd.n3350 vdd.n666 19.3944
R4116 vdd.n3350 vdd.n664 19.3944
R4117 vdd.n3354 vdd.n664 19.3944
R4118 vdd.n3354 vdd.n653 19.3944
R4119 vdd.n3366 vdd.n653 19.3944
R4120 vdd.n3366 vdd.n651 19.3944
R4121 vdd.n3370 vdd.n651 19.3944
R4122 vdd.n3370 vdd.n642 19.3944
R4123 vdd.n3383 vdd.n642 19.3944
R4124 vdd.n3383 vdd.n640 19.3944
R4125 vdd.n3390 vdd.n640 19.3944
R4126 vdd.n3390 vdd.n3389 19.3944
R4127 vdd.n3389 vdd.n631 19.3944
R4128 vdd.n3403 vdd.n631 19.3944
R4129 vdd.n3404 vdd.n3403 19.3944
R4130 vdd.n3404 vdd.n629 19.3944
R4131 vdd.n3408 vdd.n629 19.3944
R4132 vdd.n3410 vdd.n3408 19.3944
R4133 vdd.n3411 vdd.n3410 19.3944
R4134 vdd.n3411 vdd.n627 19.3944
R4135 vdd.n3415 vdd.n627 19.3944
R4136 vdd.n3417 vdd.n3415 19.3944
R4137 vdd.n3418 vdd.n3417 19.3944
R4138 vdd.n3418 vdd.n625 19.3944
R4139 vdd.n3422 vdd.n625 19.3944
R4140 vdd.n3425 vdd.n3422 19.3944
R4141 vdd.n3426 vdd.n3425 19.3944
R4142 vdd.n3426 vdd.n623 19.3944
R4143 vdd.n3430 vdd.n623 19.3944
R4144 vdd.n3432 vdd.n3430 19.3944
R4145 vdd.n3433 vdd.n3432 19.3944
R4146 vdd.n3433 vdd.n621 19.3944
R4147 vdd.n3437 vdd.n621 19.3944
R4148 vdd.n3439 vdd.n3437 19.3944
R4149 vdd.n3440 vdd.n3439 19.3944
R4150 vdd.n569 vdd.n438 19.3944
R4151 vdd.n575 vdd.n438 19.3944
R4152 vdd.n576 vdd.n575 19.3944
R4153 vdd.n579 vdd.n576 19.3944
R4154 vdd.n579 vdd.n436 19.3944
R4155 vdd.n585 vdd.n436 19.3944
R4156 vdd.n586 vdd.n585 19.3944
R4157 vdd.n589 vdd.n586 19.3944
R4158 vdd.n589 vdd.n434 19.3944
R4159 vdd.n595 vdd.n434 19.3944
R4160 vdd.n596 vdd.n595 19.3944
R4161 vdd.n599 vdd.n596 19.3944
R4162 vdd.n599 vdd.n432 19.3944
R4163 vdd.n605 vdd.n432 19.3944
R4164 vdd.n606 vdd.n605 19.3944
R4165 vdd.n609 vdd.n606 19.3944
R4166 vdd.n609 vdd.n430 19.3944
R4167 vdd.n615 vdd.n430 19.3944
R4168 vdd.n617 vdd.n615 19.3944
R4169 vdd.n618 vdd.n617 19.3944
R4170 vdd.n516 vdd.n515 19.3944
R4171 vdd.n519 vdd.n516 19.3944
R4172 vdd.n519 vdd.n450 19.3944
R4173 vdd.n525 vdd.n450 19.3944
R4174 vdd.n526 vdd.n525 19.3944
R4175 vdd.n529 vdd.n526 19.3944
R4176 vdd.n529 vdd.n448 19.3944
R4177 vdd.n535 vdd.n448 19.3944
R4178 vdd.n536 vdd.n535 19.3944
R4179 vdd.n539 vdd.n536 19.3944
R4180 vdd.n539 vdd.n446 19.3944
R4181 vdd.n545 vdd.n446 19.3944
R4182 vdd.n546 vdd.n545 19.3944
R4183 vdd.n549 vdd.n546 19.3944
R4184 vdd.n549 vdd.n444 19.3944
R4185 vdd.n555 vdd.n444 19.3944
R4186 vdd.n556 vdd.n555 19.3944
R4187 vdd.n559 vdd.n556 19.3944
R4188 vdd.n559 vdd.n442 19.3944
R4189 vdd.n565 vdd.n442 19.3944
R4190 vdd.n466 vdd.n465 19.3944
R4191 vdd.n469 vdd.n466 19.3944
R4192 vdd.n469 vdd.n462 19.3944
R4193 vdd.n475 vdd.n462 19.3944
R4194 vdd.n476 vdd.n475 19.3944
R4195 vdd.n479 vdd.n476 19.3944
R4196 vdd.n479 vdd.n460 19.3944
R4197 vdd.n485 vdd.n460 19.3944
R4198 vdd.n486 vdd.n485 19.3944
R4199 vdd.n489 vdd.n486 19.3944
R4200 vdd.n489 vdd.n458 19.3944
R4201 vdd.n495 vdd.n458 19.3944
R4202 vdd.n496 vdd.n495 19.3944
R4203 vdd.n499 vdd.n496 19.3944
R4204 vdd.n499 vdd.n456 19.3944
R4205 vdd.n505 vdd.n456 19.3944
R4206 vdd.n506 vdd.n505 19.3944
R4207 vdd.n509 vdd.n506 19.3944
R4208 vdd.n3325 vdd.n683 19.3944
R4209 vdd.n3325 vdd.n681 19.3944
R4210 vdd.n3329 vdd.n681 19.3944
R4211 vdd.n3329 vdd.n671 19.3944
R4212 vdd.n3342 vdd.n671 19.3944
R4213 vdd.n3342 vdd.n669 19.3944
R4214 vdd.n3346 vdd.n669 19.3944
R4215 vdd.n3346 vdd.n660 19.3944
R4216 vdd.n3358 vdd.n660 19.3944
R4217 vdd.n3358 vdd.n658 19.3944
R4218 vdd.n3362 vdd.n658 19.3944
R4219 vdd.n3362 vdd.n648 19.3944
R4220 vdd.n3375 vdd.n648 19.3944
R4221 vdd.n3375 vdd.n646 19.3944
R4222 vdd.n3379 vdd.n646 19.3944
R4223 vdd.n3379 vdd.n637 19.3944
R4224 vdd.n3394 vdd.n637 19.3944
R4225 vdd.n3394 vdd.n635 19.3944
R4226 vdd.n3398 vdd.n635 19.3944
R4227 vdd.n3398 vdd.n336 19.3944
R4228 vdd.n3489 vdd.n336 19.3944
R4229 vdd.n3489 vdd.n337 19.3944
R4230 vdd.n3483 vdd.n337 19.3944
R4231 vdd.n3483 vdd.n3482 19.3944
R4232 vdd.n3482 vdd.n3481 19.3944
R4233 vdd.n3481 vdd.n349 19.3944
R4234 vdd.n3475 vdd.n349 19.3944
R4235 vdd.n3475 vdd.n3474 19.3944
R4236 vdd.n3474 vdd.n3473 19.3944
R4237 vdd.n3473 vdd.n359 19.3944
R4238 vdd.n3467 vdd.n359 19.3944
R4239 vdd.n3467 vdd.n3466 19.3944
R4240 vdd.n3466 vdd.n3465 19.3944
R4241 vdd.n3465 vdd.n370 19.3944
R4242 vdd.n3459 vdd.n370 19.3944
R4243 vdd.n3459 vdd.n3458 19.3944
R4244 vdd.n3458 vdd.n3457 19.3944
R4245 vdd.n3457 vdd.n381 19.3944
R4246 vdd.n3451 vdd.n381 19.3944
R4247 vdd.n3451 vdd.n3450 19.3944
R4248 vdd.n3450 vdd.n3449 19.3944
R4249 vdd.n3272 vdd.n747 19.3944
R4250 vdd.n3272 vdd.n3269 19.3944
R4251 vdd.n3269 vdd.n3266 19.3944
R4252 vdd.n3266 vdd.n3265 19.3944
R4253 vdd.n3265 vdd.n3262 19.3944
R4254 vdd.n3262 vdd.n3261 19.3944
R4255 vdd.n3261 vdd.n3258 19.3944
R4256 vdd.n3258 vdd.n3257 19.3944
R4257 vdd.n3257 vdd.n3254 19.3944
R4258 vdd.n3254 vdd.n3253 19.3944
R4259 vdd.n3253 vdd.n3250 19.3944
R4260 vdd.n3250 vdd.n3249 19.3944
R4261 vdd.n3249 vdd.n3246 19.3944
R4262 vdd.n3246 vdd.n3245 19.3944
R4263 vdd.n3245 vdd.n3242 19.3944
R4264 vdd.n3242 vdd.n3241 19.3944
R4265 vdd.n3241 vdd.n3238 19.3944
R4266 vdd.n3238 vdd.n3237 19.3944
R4267 vdd.n3237 vdd.n3234 19.3944
R4268 vdd.n3234 vdd.n3233 19.3944
R4269 vdd.n3312 vdd.n3311 19.3944
R4270 vdd.n3311 vdd.n3310 19.3944
R4271 vdd.n732 vdd.n729 19.3944
R4272 vdd.n3306 vdd.n3305 19.3944
R4273 vdd.n3305 vdd.n3302 19.3944
R4274 vdd.n3302 vdd.n3301 19.3944
R4275 vdd.n3301 vdd.n3298 19.3944
R4276 vdd.n3298 vdd.n3297 19.3944
R4277 vdd.n3297 vdd.n3294 19.3944
R4278 vdd.n3294 vdd.n3293 19.3944
R4279 vdd.n3293 vdd.n3290 19.3944
R4280 vdd.n3290 vdd.n3289 19.3944
R4281 vdd.n3289 vdd.n3286 19.3944
R4282 vdd.n3286 vdd.n3285 19.3944
R4283 vdd.n3285 vdd.n3282 19.3944
R4284 vdd.n3282 vdd.n3281 19.3944
R4285 vdd.n3226 vdd.n767 19.3944
R4286 vdd.n3226 vdd.n3223 19.3944
R4287 vdd.n3223 vdd.n3220 19.3944
R4288 vdd.n3220 vdd.n3219 19.3944
R4289 vdd.n3219 vdd.n3216 19.3944
R4290 vdd.n3216 vdd.n3215 19.3944
R4291 vdd.n3215 vdd.n3212 19.3944
R4292 vdd.n3212 vdd.n3211 19.3944
R4293 vdd.n3211 vdd.n3208 19.3944
R4294 vdd.n3208 vdd.n3207 19.3944
R4295 vdd.n3207 vdd.n3204 19.3944
R4296 vdd.n3204 vdd.n3203 19.3944
R4297 vdd.n3203 vdd.n3200 19.3944
R4298 vdd.n3200 vdd.n3199 19.3944
R4299 vdd.n3199 vdd.n3196 19.3944
R4300 vdd.n3196 vdd.n3195 19.3944
R4301 vdd.n3192 vdd.n3191 19.3944
R4302 vdd.n3188 vdd.n3187 19.3944
R4303 vdd.n1719 vdd.n1715 19.0066
R4304 vdd.n2307 vdd.n1189 19.0066
R4305 vdd.n569 vdd.n566 19.0066
R4306 vdd.n3230 vdd.n767 19.0066
R4307 vdd.n1254 vdd.n1253 16.0975
R4308 vdd.n982 vdd.n981 16.0975
R4309 vdd.n1680 vdd.n1679 16.0975
R4310 vdd.n1718 vdd.n1717 16.0975
R4311 vdd.n1614 vdd.n1613 16.0975
R4312 vdd.n2270 vdd.n2269 16.0975
R4313 vdd.n1191 vdd.n1190 16.0975
R4314 vdd.n1151 vdd.n1150 16.0975
R4315 vdd.n1274 vdd.n1273 16.0975
R4316 vdd.n973 vdd.n972 16.0975
R4317 vdd.n2705 vdd.n2704 16.0975
R4318 vdd.n427 vdd.n426 16.0975
R4319 vdd.n441 vdd.n440 16.0975
R4320 vdd.n453 vdd.n452 16.0975
R4321 vdd.n769 vdd.n768 16.0975
R4322 vdd.n3277 vdd.n3276 16.0975
R4323 vdd.n833 vdd.n832 16.0975
R4324 vdd.n2702 vdd.n2701 16.0975
R4325 vdd.n689 vdd.n688 16.0975
R4326 vdd.n800 vdd.n799 16.0975
R4327 vdd.t10 vdd.n2665 15.4182
R4328 vdd.n2938 vdd.t46 15.4182
R4329 vdd.n28 vdd.n27 14.4007
R4330 vdd.n2417 vdd.n1076 14.0578
R4331 vdd.n3151 vdd.n692 14.0578
R4332 vdd.n328 vdd.n293 13.1884
R4333 vdd.n269 vdd.n234 13.1884
R4334 vdd.n226 vdd.n191 13.1884
R4335 vdd.n167 vdd.n132 13.1884
R4336 vdd.n125 vdd.n90 13.1884
R4337 vdd.n66 vdd.n31 13.1884
R4338 vdd.n2109 vdd.n2074 13.1884
R4339 vdd.n2168 vdd.n2133 13.1884
R4340 vdd.n2007 vdd.n1972 13.1884
R4341 vdd.n2066 vdd.n2031 13.1884
R4342 vdd.n1906 vdd.n1871 13.1884
R4343 vdd.n1965 vdd.n1930 13.1884
R4344 vdd.n1750 vdd.n1615 12.9944
R4345 vdd.n1754 vdd.n1615 12.9944
R4346 vdd.n2346 vdd.n1149 12.9944
R4347 vdd.n2347 vdd.n2346 12.9944
R4348 vdd.n515 vdd.n454 12.9944
R4349 vdd.n509 vdd.n454 12.9944
R4350 vdd.n3278 vdd.n747 12.9944
R4351 vdd.n3281 vdd.n3278 12.9944
R4352 vdd.n329 vdd.n291 12.8005
R4353 vdd.n324 vdd.n295 12.8005
R4354 vdd.n270 vdd.n232 12.8005
R4355 vdd.n265 vdd.n236 12.8005
R4356 vdd.n227 vdd.n189 12.8005
R4357 vdd.n222 vdd.n193 12.8005
R4358 vdd.n168 vdd.n130 12.8005
R4359 vdd.n163 vdd.n134 12.8005
R4360 vdd.n126 vdd.n88 12.8005
R4361 vdd.n121 vdd.n92 12.8005
R4362 vdd.n67 vdd.n29 12.8005
R4363 vdd.n62 vdd.n33 12.8005
R4364 vdd.n2110 vdd.n2072 12.8005
R4365 vdd.n2105 vdd.n2076 12.8005
R4366 vdd.n2169 vdd.n2131 12.8005
R4367 vdd.n2164 vdd.n2135 12.8005
R4368 vdd.n2008 vdd.n1970 12.8005
R4369 vdd.n2003 vdd.n1974 12.8005
R4370 vdd.n2067 vdd.n2029 12.8005
R4371 vdd.n2062 vdd.n2033 12.8005
R4372 vdd.n1907 vdd.n1869 12.8005
R4373 vdd.n1902 vdd.n1873 12.8005
R4374 vdd.n1966 vdd.n1928 12.8005
R4375 vdd.n1961 vdd.n1932 12.8005
R4376 vdd.n323 vdd.n296 12.0247
R4377 vdd.n264 vdd.n237 12.0247
R4378 vdd.n221 vdd.n194 12.0247
R4379 vdd.n162 vdd.n135 12.0247
R4380 vdd.n120 vdd.n93 12.0247
R4381 vdd.n61 vdd.n34 12.0247
R4382 vdd.n2104 vdd.n2077 12.0247
R4383 vdd.n2163 vdd.n2136 12.0247
R4384 vdd.n2002 vdd.n1975 12.0247
R4385 vdd.n2061 vdd.n2034 12.0247
R4386 vdd.n1901 vdd.n1874 12.0247
R4387 vdd.n1960 vdd.n1933 12.0247
R4388 vdd.n1789 vdd.n1545 11.337
R4389 vdd.n1798 vdd.n1545 11.337
R4390 vdd.n1798 vdd.n1797 11.337
R4391 vdd.n1806 vdd.n1539 11.337
R4392 vdd.n1815 vdd.n1814 11.337
R4393 vdd.n1831 vdd.n1523 11.337
R4394 vdd.n1839 vdd.n1516 11.337
R4395 vdd.n1848 vdd.n1847 11.337
R4396 vdd.n1856 vdd.n1505 11.337
R4397 vdd.n2179 vdd.n1494 11.337
R4398 vdd.n2188 vdd.n1488 11.337
R4399 vdd.n2196 vdd.n1482 11.337
R4400 vdd.n2205 vdd.n2204 11.337
R4401 vdd.n2221 vdd.n1466 11.337
R4402 vdd.n2229 vdd.n1459 11.337
R4403 vdd.n2238 vdd.n2237 11.337
R4404 vdd.n2246 vdd.n1442 11.337
R4405 vdd.n2257 vdd.n1442 11.337
R4406 vdd.n2257 vdd.n2256 11.337
R4407 vdd.n3323 vdd.n678 11.337
R4408 vdd.n3331 vdd.n678 11.337
R4409 vdd.n3331 vdd.n679 11.337
R4410 vdd.n3340 vdd.n3339 11.337
R4411 vdd.n3356 vdd.n662 11.337
R4412 vdd.n3364 vdd.n655 11.337
R4413 vdd.n3373 vdd.n3372 11.337
R4414 vdd.n3381 vdd.n644 11.337
R4415 vdd.n3400 vdd.n633 11.337
R4416 vdd.n3487 vdd.n340 11.337
R4417 vdd.n3485 vdd.n344 11.337
R4418 vdd.n3479 vdd.n3478 11.337
R4419 vdd.n3471 vdd.n361 11.337
R4420 vdd.n3470 vdd.n3469 11.337
R4421 vdd.n3463 vdd.n3462 11.337
R4422 vdd.n3461 vdd.n375 11.337
R4423 vdd.n3455 vdd.n3454 11.337
R4424 vdd.n3454 vdd.n3453 11.337
R4425 vdd.n3453 vdd.n386 11.337
R4426 vdd.n320 vdd.n319 11.249
R4427 vdd.n261 vdd.n260 11.249
R4428 vdd.n218 vdd.n217 11.249
R4429 vdd.n159 vdd.n158 11.249
R4430 vdd.n117 vdd.n116 11.249
R4431 vdd.n58 vdd.n57 11.249
R4432 vdd.n2101 vdd.n2100 11.249
R4433 vdd.n2160 vdd.n2159 11.249
R4434 vdd.n1999 vdd.n1998 11.249
R4435 vdd.n2058 vdd.n2057 11.249
R4436 vdd.n1898 vdd.n1897 11.249
R4437 vdd.n1957 vdd.n1956 11.249
R4438 vdd.n1587 vdd.t261 11.2237
R4439 vdd.n3447 vdd.t247 11.2237
R4440 vdd.t142 vdd.n1460 10.7702
R4441 vdd.n3348 vdd.t66 10.7702
R4442 vdd.n305 vdd.n304 10.7238
R4443 vdd.n246 vdd.n245 10.7238
R4444 vdd.n203 vdd.n202 10.7238
R4445 vdd.n144 vdd.n143 10.7238
R4446 vdd.n102 vdd.n101 10.7238
R4447 vdd.n43 vdd.n42 10.7238
R4448 vdd.n2086 vdd.n2085 10.7238
R4449 vdd.n2145 vdd.n2144 10.7238
R4450 vdd.n1984 vdd.n1983 10.7238
R4451 vdd.n2043 vdd.n2042 10.7238
R4452 vdd.n1883 vdd.n1882 10.7238
R4453 vdd.n1942 vdd.n1941 10.7238
R4454 vdd.n2593 vdd.t17 10.6568
R4455 vdd.t222 vdd.n928 10.6568
R4456 vdd.n2426 vdd.n1074 10.6151
R4457 vdd.n2427 vdd.n2426 10.6151
R4458 vdd.n2428 vdd.n2427 10.6151
R4459 vdd.n2428 vdd.n1063 10.6151
R4460 vdd.n2438 vdd.n1063 10.6151
R4461 vdd.n2439 vdd.n2438 10.6151
R4462 vdd.n2440 vdd.n2439 10.6151
R4463 vdd.n2440 vdd.n1050 10.6151
R4464 vdd.n2450 vdd.n1050 10.6151
R4465 vdd.n2451 vdd.n2450 10.6151
R4466 vdd.n2452 vdd.n2451 10.6151
R4467 vdd.n2452 vdd.n1038 10.6151
R4468 vdd.n2463 vdd.n1038 10.6151
R4469 vdd.n2464 vdd.n2463 10.6151
R4470 vdd.n2465 vdd.n2464 10.6151
R4471 vdd.n2465 vdd.n1026 10.6151
R4472 vdd.n2475 vdd.n1026 10.6151
R4473 vdd.n2476 vdd.n2475 10.6151
R4474 vdd.n2477 vdd.n2476 10.6151
R4475 vdd.n2477 vdd.n1014 10.6151
R4476 vdd.n2487 vdd.n1014 10.6151
R4477 vdd.n2488 vdd.n2487 10.6151
R4478 vdd.n2489 vdd.n2488 10.6151
R4479 vdd.n2489 vdd.n1003 10.6151
R4480 vdd.n2499 vdd.n1003 10.6151
R4481 vdd.n2500 vdd.n2499 10.6151
R4482 vdd.n2501 vdd.n2500 10.6151
R4483 vdd.n2501 vdd.n990 10.6151
R4484 vdd.n2513 vdd.n990 10.6151
R4485 vdd.n2514 vdd.n2513 10.6151
R4486 vdd.n2516 vdd.n2514 10.6151
R4487 vdd.n2516 vdd.n2515 10.6151
R4488 vdd.n2515 vdd.n971 10.6151
R4489 vdd.n2663 vdd.n2662 10.6151
R4490 vdd.n2662 vdd.n2661 10.6151
R4491 vdd.n2661 vdd.n2658 10.6151
R4492 vdd.n2658 vdd.n2657 10.6151
R4493 vdd.n2657 vdd.n2654 10.6151
R4494 vdd.n2654 vdd.n2653 10.6151
R4495 vdd.n2653 vdd.n2650 10.6151
R4496 vdd.n2650 vdd.n2649 10.6151
R4497 vdd.n2649 vdd.n2646 10.6151
R4498 vdd.n2646 vdd.n2645 10.6151
R4499 vdd.n2645 vdd.n2642 10.6151
R4500 vdd.n2642 vdd.n2641 10.6151
R4501 vdd.n2641 vdd.n2638 10.6151
R4502 vdd.n2638 vdd.n2637 10.6151
R4503 vdd.n2637 vdd.n2634 10.6151
R4504 vdd.n2634 vdd.n2633 10.6151
R4505 vdd.n2633 vdd.n2630 10.6151
R4506 vdd.n2630 vdd.n2629 10.6151
R4507 vdd.n2629 vdd.n2626 10.6151
R4508 vdd.n2626 vdd.n2625 10.6151
R4509 vdd.n2625 vdd.n2622 10.6151
R4510 vdd.n2622 vdd.n2621 10.6151
R4511 vdd.n2621 vdd.n2618 10.6151
R4512 vdd.n2618 vdd.n2617 10.6151
R4513 vdd.n2617 vdd.n2614 10.6151
R4514 vdd.n2614 vdd.n2613 10.6151
R4515 vdd.n2613 vdd.n2610 10.6151
R4516 vdd.n2610 vdd.n2609 10.6151
R4517 vdd.n2609 vdd.n2606 10.6151
R4518 vdd.n2606 vdd.n2605 10.6151
R4519 vdd.n2605 vdd.n2602 10.6151
R4520 vdd.n2600 vdd.n2597 10.6151
R4521 vdd.n2597 vdd.n2596 10.6151
R4522 vdd.n1311 vdd.n1310 10.6151
R4523 vdd.n1313 vdd.n1311 10.6151
R4524 vdd.n1314 vdd.n1313 10.6151
R4525 vdd.n1316 vdd.n1314 10.6151
R4526 vdd.n1317 vdd.n1316 10.6151
R4527 vdd.n1319 vdd.n1317 10.6151
R4528 vdd.n1320 vdd.n1319 10.6151
R4529 vdd.n1322 vdd.n1320 10.6151
R4530 vdd.n1323 vdd.n1322 10.6151
R4531 vdd.n1325 vdd.n1323 10.6151
R4532 vdd.n1326 vdd.n1325 10.6151
R4533 vdd.n1328 vdd.n1326 10.6151
R4534 vdd.n1329 vdd.n1328 10.6151
R4535 vdd.n1331 vdd.n1329 10.6151
R4536 vdd.n1332 vdd.n1331 10.6151
R4537 vdd.n1334 vdd.n1332 10.6151
R4538 vdd.n1335 vdd.n1334 10.6151
R4539 vdd.n1357 vdd.n1335 10.6151
R4540 vdd.n1357 vdd.n1356 10.6151
R4541 vdd.n1356 vdd.n1355 10.6151
R4542 vdd.n1355 vdd.n1353 10.6151
R4543 vdd.n1353 vdd.n1352 10.6151
R4544 vdd.n1352 vdd.n1350 10.6151
R4545 vdd.n1350 vdd.n1349 10.6151
R4546 vdd.n1349 vdd.n1347 10.6151
R4547 vdd.n1347 vdd.n1346 10.6151
R4548 vdd.n1346 vdd.n1344 10.6151
R4549 vdd.n1344 vdd.n1343 10.6151
R4550 vdd.n1343 vdd.n1341 10.6151
R4551 vdd.n1341 vdd.n1340 10.6151
R4552 vdd.n1340 vdd.n1337 10.6151
R4553 vdd.n1337 vdd.n1336 10.6151
R4554 vdd.n1336 vdd.n974 10.6151
R4555 vdd.n2414 vdd.n2413 10.6151
R4556 vdd.n2413 vdd.n2412 10.6151
R4557 vdd.n2412 vdd.n2411 10.6151
R4558 vdd.n2411 vdd.n2409 10.6151
R4559 vdd.n2409 vdd.n2406 10.6151
R4560 vdd.n2406 vdd.n2405 10.6151
R4561 vdd.n2405 vdd.n2402 10.6151
R4562 vdd.n2402 vdd.n2401 10.6151
R4563 vdd.n2401 vdd.n2398 10.6151
R4564 vdd.n2398 vdd.n2397 10.6151
R4565 vdd.n2397 vdd.n2394 10.6151
R4566 vdd.n2394 vdd.n2393 10.6151
R4567 vdd.n2393 vdd.n2390 10.6151
R4568 vdd.n2390 vdd.n2389 10.6151
R4569 vdd.n2389 vdd.n2386 10.6151
R4570 vdd.n2386 vdd.n2385 10.6151
R4571 vdd.n2385 vdd.n2382 10.6151
R4572 vdd.n2382 vdd.n1119 10.6151
R4573 vdd.n1277 vdd.n1119 10.6151
R4574 vdd.n1278 vdd.n1277 10.6151
R4575 vdd.n1281 vdd.n1278 10.6151
R4576 vdd.n1282 vdd.n1281 10.6151
R4577 vdd.n1285 vdd.n1282 10.6151
R4578 vdd.n1286 vdd.n1285 10.6151
R4579 vdd.n1289 vdd.n1286 10.6151
R4580 vdd.n1290 vdd.n1289 10.6151
R4581 vdd.n1293 vdd.n1290 10.6151
R4582 vdd.n1294 vdd.n1293 10.6151
R4583 vdd.n1297 vdd.n1294 10.6151
R4584 vdd.n1298 vdd.n1297 10.6151
R4585 vdd.n1301 vdd.n1298 10.6151
R4586 vdd.n1306 vdd.n1303 10.6151
R4587 vdd.n1307 vdd.n1306 10.6151
R4588 vdd.n2866 vdd.n2865 10.6151
R4589 vdd.n2865 vdd.n2864 10.6151
R4590 vdd.n2864 vdd.n2703 10.6151
R4591 vdd.n2808 vdd.n2703 10.6151
R4592 vdd.n2809 vdd.n2808 10.6151
R4593 vdd.n2811 vdd.n2809 10.6151
R4594 vdd.n2812 vdd.n2811 10.6151
R4595 vdd.n2814 vdd.n2812 10.6151
R4596 vdd.n2815 vdd.n2814 10.6151
R4597 vdd.n2845 vdd.n2815 10.6151
R4598 vdd.n2845 vdd.n2844 10.6151
R4599 vdd.n2844 vdd.n2843 10.6151
R4600 vdd.n2843 vdd.n2841 10.6151
R4601 vdd.n2841 vdd.n2840 10.6151
R4602 vdd.n2840 vdd.n2838 10.6151
R4603 vdd.n2838 vdd.n2837 10.6151
R4604 vdd.n2837 vdd.n2835 10.6151
R4605 vdd.n2835 vdd.n2834 10.6151
R4606 vdd.n2834 vdd.n2832 10.6151
R4607 vdd.n2832 vdd.n2831 10.6151
R4608 vdd.n2831 vdd.n2829 10.6151
R4609 vdd.n2829 vdd.n2828 10.6151
R4610 vdd.n2828 vdd.n2826 10.6151
R4611 vdd.n2826 vdd.n2825 10.6151
R4612 vdd.n2825 vdd.n2823 10.6151
R4613 vdd.n2823 vdd.n2822 10.6151
R4614 vdd.n2822 vdd.n2820 10.6151
R4615 vdd.n2820 vdd.n2819 10.6151
R4616 vdd.n2819 vdd.n2817 10.6151
R4617 vdd.n2817 vdd.n2816 10.6151
R4618 vdd.n2816 vdd.n836 10.6151
R4619 vdd.n3084 vdd.n836 10.6151
R4620 vdd.n3085 vdd.n3084 10.6151
R4621 vdd.n2935 vdd.n2934 10.6151
R4622 vdd.n2934 vdd.n2933 10.6151
R4623 vdd.n2933 vdd.n2932 10.6151
R4624 vdd.n2932 vdd.n2930 10.6151
R4625 vdd.n2930 vdd.n2927 10.6151
R4626 vdd.n2927 vdd.n2926 10.6151
R4627 vdd.n2926 vdd.n2923 10.6151
R4628 vdd.n2923 vdd.n2922 10.6151
R4629 vdd.n2922 vdd.n2919 10.6151
R4630 vdd.n2919 vdd.n2918 10.6151
R4631 vdd.n2918 vdd.n2915 10.6151
R4632 vdd.n2915 vdd.n2914 10.6151
R4633 vdd.n2914 vdd.n2911 10.6151
R4634 vdd.n2911 vdd.n2910 10.6151
R4635 vdd.n2910 vdd.n2907 10.6151
R4636 vdd.n2907 vdd.n2906 10.6151
R4637 vdd.n2906 vdd.n2903 10.6151
R4638 vdd.n2903 vdd.n2902 10.6151
R4639 vdd.n2902 vdd.n2899 10.6151
R4640 vdd.n2899 vdd.n2898 10.6151
R4641 vdd.n2898 vdd.n2895 10.6151
R4642 vdd.n2895 vdd.n2894 10.6151
R4643 vdd.n2894 vdd.n2891 10.6151
R4644 vdd.n2891 vdd.n2890 10.6151
R4645 vdd.n2890 vdd.n2887 10.6151
R4646 vdd.n2887 vdd.n2886 10.6151
R4647 vdd.n2886 vdd.n2883 10.6151
R4648 vdd.n2883 vdd.n2882 10.6151
R4649 vdd.n2882 vdd.n2879 10.6151
R4650 vdd.n2879 vdd.n2878 10.6151
R4651 vdd.n2878 vdd.n2875 10.6151
R4652 vdd.n2873 vdd.n2870 10.6151
R4653 vdd.n2870 vdd.n2869 10.6151
R4654 vdd.n2947 vdd.n926 10.6151
R4655 vdd.n2948 vdd.n2947 10.6151
R4656 vdd.n2949 vdd.n2948 10.6151
R4657 vdd.n2949 vdd.n915 10.6151
R4658 vdd.n2959 vdd.n915 10.6151
R4659 vdd.n2960 vdd.n2959 10.6151
R4660 vdd.n2961 vdd.n2960 10.6151
R4661 vdd.n2961 vdd.n903 10.6151
R4662 vdd.n2971 vdd.n903 10.6151
R4663 vdd.n2972 vdd.n2971 10.6151
R4664 vdd.n2973 vdd.n2972 10.6151
R4665 vdd.n2973 vdd.n891 10.6151
R4666 vdd.n2983 vdd.n891 10.6151
R4667 vdd.n2984 vdd.n2983 10.6151
R4668 vdd.n2985 vdd.n2984 10.6151
R4669 vdd.n2985 vdd.n880 10.6151
R4670 vdd.n2995 vdd.n880 10.6151
R4671 vdd.n2996 vdd.n2995 10.6151
R4672 vdd.n2997 vdd.n2996 10.6151
R4673 vdd.n2997 vdd.n866 10.6151
R4674 vdd.n3008 vdd.n866 10.6151
R4675 vdd.n3009 vdd.n3008 10.6151
R4676 vdd.n3010 vdd.n3009 10.6151
R4677 vdd.n3010 vdd.n855 10.6151
R4678 vdd.n3020 vdd.n855 10.6151
R4679 vdd.n3021 vdd.n3020 10.6151
R4680 vdd.n3022 vdd.n3021 10.6151
R4681 vdd.n3022 vdd.n841 10.6151
R4682 vdd.n3077 vdd.n841 10.6151
R4683 vdd.n3078 vdd.n3077 10.6151
R4684 vdd.n3079 vdd.n3078 10.6151
R4685 vdd.n3079 vdd.n810 10.6151
R4686 vdd.n3149 vdd.n810 10.6151
R4687 vdd.n3148 vdd.n3147 10.6151
R4688 vdd.n3147 vdd.n811 10.6151
R4689 vdd.n812 vdd.n811 10.6151
R4690 vdd.n3140 vdd.n812 10.6151
R4691 vdd.n3140 vdd.n3139 10.6151
R4692 vdd.n3139 vdd.n3138 10.6151
R4693 vdd.n3138 vdd.n814 10.6151
R4694 vdd.n3133 vdd.n814 10.6151
R4695 vdd.n3133 vdd.n3132 10.6151
R4696 vdd.n3132 vdd.n3131 10.6151
R4697 vdd.n3131 vdd.n817 10.6151
R4698 vdd.n3126 vdd.n817 10.6151
R4699 vdd.n3126 vdd.n3125 10.6151
R4700 vdd.n3125 vdd.n3124 10.6151
R4701 vdd.n3124 vdd.n820 10.6151
R4702 vdd.n3119 vdd.n820 10.6151
R4703 vdd.n3119 vdd.n731 10.6151
R4704 vdd.n3115 vdd.n731 10.6151
R4705 vdd.n3115 vdd.n3114 10.6151
R4706 vdd.n3114 vdd.n3113 10.6151
R4707 vdd.n3113 vdd.n823 10.6151
R4708 vdd.n3108 vdd.n823 10.6151
R4709 vdd.n3108 vdd.n3107 10.6151
R4710 vdd.n3107 vdd.n3106 10.6151
R4711 vdd.n3106 vdd.n826 10.6151
R4712 vdd.n3101 vdd.n826 10.6151
R4713 vdd.n3101 vdd.n3100 10.6151
R4714 vdd.n3100 vdd.n3099 10.6151
R4715 vdd.n3099 vdd.n829 10.6151
R4716 vdd.n3094 vdd.n829 10.6151
R4717 vdd.n3094 vdd.n3093 10.6151
R4718 vdd.n3091 vdd.n834 10.6151
R4719 vdd.n3086 vdd.n834 10.6151
R4720 vdd.n3067 vdd.n3028 10.6151
R4721 vdd.n3062 vdd.n3028 10.6151
R4722 vdd.n3062 vdd.n3061 10.6151
R4723 vdd.n3061 vdd.n3060 10.6151
R4724 vdd.n3060 vdd.n3030 10.6151
R4725 vdd.n3055 vdd.n3030 10.6151
R4726 vdd.n3055 vdd.n3054 10.6151
R4727 vdd.n3054 vdd.n3053 10.6151
R4728 vdd.n3053 vdd.n3033 10.6151
R4729 vdd.n3048 vdd.n3033 10.6151
R4730 vdd.n3048 vdd.n3047 10.6151
R4731 vdd.n3047 vdd.n3046 10.6151
R4732 vdd.n3046 vdd.n3036 10.6151
R4733 vdd.n3041 vdd.n3036 10.6151
R4734 vdd.n3041 vdd.n3040 10.6151
R4735 vdd.n3040 vdd.n785 10.6151
R4736 vdd.n3184 vdd.n785 10.6151
R4737 vdd.n3184 vdd.n786 10.6151
R4738 vdd.n788 vdd.n786 10.6151
R4739 vdd.n3177 vdd.n788 10.6151
R4740 vdd.n3177 vdd.n3176 10.6151
R4741 vdd.n3176 vdd.n3175 10.6151
R4742 vdd.n3175 vdd.n790 10.6151
R4743 vdd.n3170 vdd.n790 10.6151
R4744 vdd.n3170 vdd.n3169 10.6151
R4745 vdd.n3169 vdd.n3168 10.6151
R4746 vdd.n3168 vdd.n793 10.6151
R4747 vdd.n3163 vdd.n793 10.6151
R4748 vdd.n3163 vdd.n3162 10.6151
R4749 vdd.n3162 vdd.n3161 10.6151
R4750 vdd.n3161 vdd.n796 10.6151
R4751 vdd.n3156 vdd.n3155 10.6151
R4752 vdd.n3155 vdd.n3154 10.6151
R4753 vdd.n2774 vdd.n2773 10.6151
R4754 vdd.n2860 vdd.n2774 10.6151
R4755 vdd.n2860 vdd.n2859 10.6151
R4756 vdd.n2859 vdd.n2858 10.6151
R4757 vdd.n2858 vdd.n2856 10.6151
R4758 vdd.n2856 vdd.n2855 10.6151
R4759 vdd.n2855 vdd.n2853 10.6151
R4760 vdd.n2853 vdd.n2852 10.6151
R4761 vdd.n2852 vdd.n2850 10.6151
R4762 vdd.n2850 vdd.n2849 10.6151
R4763 vdd.n2849 vdd.n2806 10.6151
R4764 vdd.n2806 vdd.n2805 10.6151
R4765 vdd.n2805 vdd.n2803 10.6151
R4766 vdd.n2803 vdd.n2802 10.6151
R4767 vdd.n2802 vdd.n2800 10.6151
R4768 vdd.n2800 vdd.n2799 10.6151
R4769 vdd.n2799 vdd.n2797 10.6151
R4770 vdd.n2797 vdd.n2796 10.6151
R4771 vdd.n2796 vdd.n2794 10.6151
R4772 vdd.n2794 vdd.n2793 10.6151
R4773 vdd.n2793 vdd.n2791 10.6151
R4774 vdd.n2791 vdd.n2790 10.6151
R4775 vdd.n2790 vdd.n2788 10.6151
R4776 vdd.n2788 vdd.n2787 10.6151
R4777 vdd.n2787 vdd.n2785 10.6151
R4778 vdd.n2785 vdd.n2784 10.6151
R4779 vdd.n2784 vdd.n2782 10.6151
R4780 vdd.n2782 vdd.n2781 10.6151
R4781 vdd.n2781 vdd.n2779 10.6151
R4782 vdd.n2779 vdd.n2778 10.6151
R4783 vdd.n2778 vdd.n2776 10.6151
R4784 vdd.n2776 vdd.n2775 10.6151
R4785 vdd.n2775 vdd.n802 10.6151
R4786 vdd.n2941 vdd.n932 10.6151
R4787 vdd.n2708 vdd.n932 10.6151
R4788 vdd.n2709 vdd.n2708 10.6151
R4789 vdd.n2712 vdd.n2709 10.6151
R4790 vdd.n2713 vdd.n2712 10.6151
R4791 vdd.n2716 vdd.n2713 10.6151
R4792 vdd.n2717 vdd.n2716 10.6151
R4793 vdd.n2720 vdd.n2717 10.6151
R4794 vdd.n2721 vdd.n2720 10.6151
R4795 vdd.n2724 vdd.n2721 10.6151
R4796 vdd.n2725 vdd.n2724 10.6151
R4797 vdd.n2728 vdd.n2725 10.6151
R4798 vdd.n2729 vdd.n2728 10.6151
R4799 vdd.n2732 vdd.n2729 10.6151
R4800 vdd.n2733 vdd.n2732 10.6151
R4801 vdd.n2736 vdd.n2733 10.6151
R4802 vdd.n2737 vdd.n2736 10.6151
R4803 vdd.n2740 vdd.n2737 10.6151
R4804 vdd.n2741 vdd.n2740 10.6151
R4805 vdd.n2744 vdd.n2741 10.6151
R4806 vdd.n2745 vdd.n2744 10.6151
R4807 vdd.n2748 vdd.n2745 10.6151
R4808 vdd.n2749 vdd.n2748 10.6151
R4809 vdd.n2752 vdd.n2749 10.6151
R4810 vdd.n2753 vdd.n2752 10.6151
R4811 vdd.n2756 vdd.n2753 10.6151
R4812 vdd.n2757 vdd.n2756 10.6151
R4813 vdd.n2760 vdd.n2757 10.6151
R4814 vdd.n2761 vdd.n2760 10.6151
R4815 vdd.n2764 vdd.n2761 10.6151
R4816 vdd.n2765 vdd.n2764 10.6151
R4817 vdd.n2770 vdd.n2768 10.6151
R4818 vdd.n2771 vdd.n2770 10.6151
R4819 vdd.n2943 vdd.n2942 10.6151
R4820 vdd.n2943 vdd.n921 10.6151
R4821 vdd.n2953 vdd.n921 10.6151
R4822 vdd.n2954 vdd.n2953 10.6151
R4823 vdd.n2955 vdd.n2954 10.6151
R4824 vdd.n2955 vdd.n909 10.6151
R4825 vdd.n2965 vdd.n909 10.6151
R4826 vdd.n2966 vdd.n2965 10.6151
R4827 vdd.n2967 vdd.n2966 10.6151
R4828 vdd.n2967 vdd.n897 10.6151
R4829 vdd.n2977 vdd.n897 10.6151
R4830 vdd.n2978 vdd.n2977 10.6151
R4831 vdd.n2979 vdd.n2978 10.6151
R4832 vdd.n2979 vdd.n886 10.6151
R4833 vdd.n2989 vdd.n886 10.6151
R4834 vdd.n2990 vdd.n2989 10.6151
R4835 vdd.n2991 vdd.n2990 10.6151
R4836 vdd.n2991 vdd.n873 10.6151
R4837 vdd.n3001 vdd.n873 10.6151
R4838 vdd.n3002 vdd.n3001 10.6151
R4839 vdd.n3004 vdd.n861 10.6151
R4840 vdd.n3014 vdd.n861 10.6151
R4841 vdd.n3015 vdd.n3014 10.6151
R4842 vdd.n3016 vdd.n3015 10.6151
R4843 vdd.n3016 vdd.n849 10.6151
R4844 vdd.n3026 vdd.n849 10.6151
R4845 vdd.n3027 vdd.n3026 10.6151
R4846 vdd.n3073 vdd.n3027 10.6151
R4847 vdd.n3073 vdd.n3072 10.6151
R4848 vdd.n3072 vdd.n3071 10.6151
R4849 vdd.n3071 vdd.n3070 10.6151
R4850 vdd.n3070 vdd.n3068 10.6151
R4851 vdd.n2422 vdd.n2421 10.6151
R4852 vdd.n2422 vdd.n1069 10.6151
R4853 vdd.n2432 vdd.n1069 10.6151
R4854 vdd.n2433 vdd.n2432 10.6151
R4855 vdd.n2434 vdd.n2433 10.6151
R4856 vdd.n2434 vdd.n1057 10.6151
R4857 vdd.n2444 vdd.n1057 10.6151
R4858 vdd.n2445 vdd.n2444 10.6151
R4859 vdd.n2446 vdd.n2445 10.6151
R4860 vdd.n2446 vdd.n1044 10.6151
R4861 vdd.n2456 vdd.n1044 10.6151
R4862 vdd.n2457 vdd.n2456 10.6151
R4863 vdd.n2459 vdd.n1032 10.6151
R4864 vdd.n2469 vdd.n1032 10.6151
R4865 vdd.n2470 vdd.n2469 10.6151
R4866 vdd.n2471 vdd.n2470 10.6151
R4867 vdd.n2471 vdd.n1020 10.6151
R4868 vdd.n2481 vdd.n1020 10.6151
R4869 vdd.n2482 vdd.n2481 10.6151
R4870 vdd.n2483 vdd.n2482 10.6151
R4871 vdd.n2483 vdd.n1009 10.6151
R4872 vdd.n2493 vdd.n1009 10.6151
R4873 vdd.n2494 vdd.n2493 10.6151
R4874 vdd.n2495 vdd.n2494 10.6151
R4875 vdd.n2495 vdd.n997 10.6151
R4876 vdd.n2505 vdd.n997 10.6151
R4877 vdd.n2506 vdd.n2505 10.6151
R4878 vdd.n2509 vdd.n2506 10.6151
R4879 vdd.n2509 vdd.n2508 10.6151
R4880 vdd.n2508 vdd.n2507 10.6151
R4881 vdd.n2507 vdd.n980 10.6151
R4882 vdd.n2591 vdd.n980 10.6151
R4883 vdd.n2590 vdd.n2589 10.6151
R4884 vdd.n2589 vdd.n2586 10.6151
R4885 vdd.n2586 vdd.n2585 10.6151
R4886 vdd.n2585 vdd.n2582 10.6151
R4887 vdd.n2582 vdd.n2581 10.6151
R4888 vdd.n2581 vdd.n2578 10.6151
R4889 vdd.n2578 vdd.n2577 10.6151
R4890 vdd.n2577 vdd.n2574 10.6151
R4891 vdd.n2574 vdd.n2573 10.6151
R4892 vdd.n2573 vdd.n2570 10.6151
R4893 vdd.n2570 vdd.n2569 10.6151
R4894 vdd.n2569 vdd.n2566 10.6151
R4895 vdd.n2566 vdd.n2565 10.6151
R4896 vdd.n2565 vdd.n2562 10.6151
R4897 vdd.n2562 vdd.n2561 10.6151
R4898 vdd.n2561 vdd.n2558 10.6151
R4899 vdd.n2558 vdd.n2557 10.6151
R4900 vdd.n2557 vdd.n2554 10.6151
R4901 vdd.n2554 vdd.n2553 10.6151
R4902 vdd.n2553 vdd.n2550 10.6151
R4903 vdd.n2550 vdd.n2549 10.6151
R4904 vdd.n2549 vdd.n2546 10.6151
R4905 vdd.n2546 vdd.n2545 10.6151
R4906 vdd.n2545 vdd.n2542 10.6151
R4907 vdd.n2542 vdd.n2541 10.6151
R4908 vdd.n2541 vdd.n2538 10.6151
R4909 vdd.n2538 vdd.n2537 10.6151
R4910 vdd.n2537 vdd.n2534 10.6151
R4911 vdd.n2534 vdd.n2533 10.6151
R4912 vdd.n2533 vdd.n2530 10.6151
R4913 vdd.n2530 vdd.n2529 10.6151
R4914 vdd.n2526 vdd.n2525 10.6151
R4915 vdd.n2525 vdd.n2523 10.6151
R4916 vdd.n1388 vdd.n1386 10.6151
R4917 vdd.n1386 vdd.n1385 10.6151
R4918 vdd.n1385 vdd.n1383 10.6151
R4919 vdd.n1383 vdd.n1382 10.6151
R4920 vdd.n1382 vdd.n1380 10.6151
R4921 vdd.n1380 vdd.n1379 10.6151
R4922 vdd.n1379 vdd.n1377 10.6151
R4923 vdd.n1377 vdd.n1376 10.6151
R4924 vdd.n1376 vdd.n1374 10.6151
R4925 vdd.n1374 vdd.n1373 10.6151
R4926 vdd.n1373 vdd.n1371 10.6151
R4927 vdd.n1371 vdd.n1370 10.6151
R4928 vdd.n1370 vdd.n1368 10.6151
R4929 vdd.n1368 vdd.n1367 10.6151
R4930 vdd.n1367 vdd.n1365 10.6151
R4931 vdd.n1365 vdd.n1364 10.6151
R4932 vdd.n1364 vdd.n1362 10.6151
R4933 vdd.n1362 vdd.n1361 10.6151
R4934 vdd.n1361 vdd.n1272 10.6151
R4935 vdd.n1272 vdd.n1271 10.6151
R4936 vdd.n1271 vdd.n1269 10.6151
R4937 vdd.n1269 vdd.n1268 10.6151
R4938 vdd.n1268 vdd.n1266 10.6151
R4939 vdd.n1266 vdd.n1265 10.6151
R4940 vdd.n1265 vdd.n1263 10.6151
R4941 vdd.n1263 vdd.n1262 10.6151
R4942 vdd.n1262 vdd.n1260 10.6151
R4943 vdd.n1260 vdd.n1259 10.6151
R4944 vdd.n1259 vdd.n1257 10.6151
R4945 vdd.n1257 vdd.n1256 10.6151
R4946 vdd.n1256 vdd.n984 10.6151
R4947 vdd.n2521 vdd.n984 10.6151
R4948 vdd.n2522 vdd.n2521 10.6151
R4949 vdd.n2420 vdd.n1081 10.6151
R4950 vdd.n1223 vdd.n1081 10.6151
R4951 vdd.n1224 vdd.n1223 10.6151
R4952 vdd.n1227 vdd.n1224 10.6151
R4953 vdd.n1228 vdd.n1227 10.6151
R4954 vdd.n1231 vdd.n1228 10.6151
R4955 vdd.n1232 vdd.n1231 10.6151
R4956 vdd.n1235 vdd.n1232 10.6151
R4957 vdd.n1236 vdd.n1235 10.6151
R4958 vdd.n1239 vdd.n1236 10.6151
R4959 vdd.n1240 vdd.n1239 10.6151
R4960 vdd.n1243 vdd.n1240 10.6151
R4961 vdd.n1244 vdd.n1243 10.6151
R4962 vdd.n1247 vdd.n1244 10.6151
R4963 vdd.n1248 vdd.n1247 10.6151
R4964 vdd.n1251 vdd.n1248 10.6151
R4965 vdd.n1422 vdd.n1251 10.6151
R4966 vdd.n1422 vdd.n1421 10.6151
R4967 vdd.n1421 vdd.n1419 10.6151
R4968 vdd.n1419 vdd.n1416 10.6151
R4969 vdd.n1416 vdd.n1415 10.6151
R4970 vdd.n1415 vdd.n1412 10.6151
R4971 vdd.n1412 vdd.n1411 10.6151
R4972 vdd.n1411 vdd.n1408 10.6151
R4973 vdd.n1408 vdd.n1407 10.6151
R4974 vdd.n1407 vdd.n1404 10.6151
R4975 vdd.n1404 vdd.n1403 10.6151
R4976 vdd.n1403 vdd.n1400 10.6151
R4977 vdd.n1400 vdd.n1399 10.6151
R4978 vdd.n1399 vdd.n1396 10.6151
R4979 vdd.n1396 vdd.n1395 10.6151
R4980 vdd.n1392 vdd.n1391 10.6151
R4981 vdd.n1391 vdd.n1389 10.6151
R4982 vdd.n2213 vdd.t83 10.5435
R4983 vdd.n656 vdd.t78 10.5435
R4984 vdd.n316 vdd.n298 10.4732
R4985 vdd.n257 vdd.n239 10.4732
R4986 vdd.n214 vdd.n196 10.4732
R4987 vdd.n155 vdd.n137 10.4732
R4988 vdd.n113 vdd.n95 10.4732
R4989 vdd.n54 vdd.n36 10.4732
R4990 vdd.n2097 vdd.n2079 10.4732
R4991 vdd.n2156 vdd.n2138 10.4732
R4992 vdd.n1995 vdd.n1977 10.4732
R4993 vdd.n2054 vdd.n2036 10.4732
R4994 vdd.n1894 vdd.n1876 10.4732
R4995 vdd.n1953 vdd.n1935 10.4732
R4996 vdd.t109 vdd.n2187 10.3167
R4997 vdd.n3392 vdd.t153 10.3167
R4998 vdd.n1864 vdd.t64 10.09
R4999 vdd.n3486 vdd.t97 10.09
R5000 vdd.t68 vdd.n1517 9.86327
R5001 vdd.n3477 vdd.t150 9.86327
R5002 vdd.n2382 vdd.n2381 9.78206
R5003 vdd.n3308 vdd.n731 9.78206
R5004 vdd.n3185 vdd.n3184 9.78206
R5005 vdd.n2274 vdd.n1422 9.78206
R5006 vdd.n315 vdd.n300 9.69747
R5007 vdd.n256 vdd.n241 9.69747
R5008 vdd.n213 vdd.n198 9.69747
R5009 vdd.n154 vdd.n139 9.69747
R5010 vdd.n112 vdd.n97 9.69747
R5011 vdd.n53 vdd.n38 9.69747
R5012 vdd.n2096 vdd.n2081 9.69747
R5013 vdd.n2155 vdd.n2140 9.69747
R5014 vdd.n1994 vdd.n1979 9.69747
R5015 vdd.n2053 vdd.n2038 9.69747
R5016 vdd.n1893 vdd.n1878 9.69747
R5017 vdd.n1952 vdd.n1937 9.69747
R5018 vdd.n1823 vdd.t158 9.63654
R5019 vdd.n3423 vdd.t122 9.63654
R5020 vdd.n331 vdd.n330 9.45567
R5021 vdd.n272 vdd.n271 9.45567
R5022 vdd.n229 vdd.n228 9.45567
R5023 vdd.n170 vdd.n169 9.45567
R5024 vdd.n128 vdd.n127 9.45567
R5025 vdd.n69 vdd.n68 9.45567
R5026 vdd.n2112 vdd.n2111 9.45567
R5027 vdd.n2171 vdd.n2170 9.45567
R5028 vdd.n2010 vdd.n2009 9.45567
R5029 vdd.n2069 vdd.n2068 9.45567
R5030 vdd.n1909 vdd.n1908 9.45567
R5031 vdd.n1968 vdd.n1967 9.45567
R5032 vdd.n1797 vdd.t72 9.40981
R5033 vdd.n3455 vdd.t87 9.40981
R5034 vdd.n2344 vdd.n1149 9.3005
R5035 vdd.n2343 vdd.n2342 9.3005
R5036 vdd.n1155 vdd.n1154 9.3005
R5037 vdd.n2337 vdd.n1159 9.3005
R5038 vdd.n2336 vdd.n1160 9.3005
R5039 vdd.n2335 vdd.n1161 9.3005
R5040 vdd.n1165 vdd.n1162 9.3005
R5041 vdd.n2330 vdd.n1166 9.3005
R5042 vdd.n2329 vdd.n1167 9.3005
R5043 vdd.n2328 vdd.n1168 9.3005
R5044 vdd.n1172 vdd.n1169 9.3005
R5045 vdd.n2323 vdd.n1173 9.3005
R5046 vdd.n2322 vdd.n1174 9.3005
R5047 vdd.n2321 vdd.n1175 9.3005
R5048 vdd.n1179 vdd.n1176 9.3005
R5049 vdd.n2316 vdd.n1180 9.3005
R5050 vdd.n2315 vdd.n1181 9.3005
R5051 vdd.n2314 vdd.n1182 9.3005
R5052 vdd.n1186 vdd.n1183 9.3005
R5053 vdd.n2309 vdd.n1187 9.3005
R5054 vdd.n2308 vdd.n1188 9.3005
R5055 vdd.n2307 vdd.n2306 9.3005
R5056 vdd.n2305 vdd.n1189 9.3005
R5057 vdd.n2304 vdd.n2303 9.3005
R5058 vdd.n1195 vdd.n1194 9.3005
R5059 vdd.n2298 vdd.n1199 9.3005
R5060 vdd.n2297 vdd.n1200 9.3005
R5061 vdd.n2296 vdd.n1201 9.3005
R5062 vdd.n1205 vdd.n1202 9.3005
R5063 vdd.n2291 vdd.n1206 9.3005
R5064 vdd.n2290 vdd.n1207 9.3005
R5065 vdd.n2289 vdd.n1208 9.3005
R5066 vdd.n1212 vdd.n1209 9.3005
R5067 vdd.n2284 vdd.n1213 9.3005
R5068 vdd.n2283 vdd.n1214 9.3005
R5069 vdd.n2282 vdd.n1215 9.3005
R5070 vdd.n1219 vdd.n1216 9.3005
R5071 vdd.n2277 vdd.n1220 9.3005
R5072 vdd.n2346 vdd.n2345 9.3005
R5073 vdd.n2368 vdd.n1120 9.3005
R5074 vdd.n2367 vdd.n1128 9.3005
R5075 vdd.n1132 vdd.n1129 9.3005
R5076 vdd.n2362 vdd.n1133 9.3005
R5077 vdd.n2361 vdd.n1134 9.3005
R5078 vdd.n2360 vdd.n1135 9.3005
R5079 vdd.n1139 vdd.n1136 9.3005
R5080 vdd.n2355 vdd.n1140 9.3005
R5081 vdd.n2354 vdd.n1141 9.3005
R5082 vdd.n2353 vdd.n1142 9.3005
R5083 vdd.n1146 vdd.n1143 9.3005
R5084 vdd.n2348 vdd.n1147 9.3005
R5085 vdd.n2347 vdd.n1148 9.3005
R5086 vdd.n2380 vdd.n2379 9.3005
R5087 vdd.n1124 vdd.n1123 9.3005
R5088 vdd.n2177 vdd.n2176 9.3005
R5089 vdd.n1486 vdd.n1485 9.3005
R5090 vdd.n2191 vdd.n2190 9.3005
R5091 vdd.n2192 vdd.n1484 9.3005
R5092 vdd.n2194 vdd.n2193 9.3005
R5093 vdd.n1475 vdd.n1474 9.3005
R5094 vdd.n2208 vdd.n2207 9.3005
R5095 vdd.n2209 vdd.n1473 9.3005
R5096 vdd.n2211 vdd.n2210 9.3005
R5097 vdd.n1464 vdd.n1463 9.3005
R5098 vdd.n2224 vdd.n2223 9.3005
R5099 vdd.n2225 vdd.n1462 9.3005
R5100 vdd.n2227 vdd.n2226 9.3005
R5101 vdd.n1452 vdd.n1451 9.3005
R5102 vdd.n2241 vdd.n2240 9.3005
R5103 vdd.n2242 vdd.n1450 9.3005
R5104 vdd.n2244 vdd.n2243 9.3005
R5105 vdd.n1440 vdd.n1439 9.3005
R5106 vdd.n2260 vdd.n2259 9.3005
R5107 vdd.n2261 vdd.n1438 9.3005
R5108 vdd.n2263 vdd.n2262 9.3005
R5109 vdd.n307 vdd.n306 9.3005
R5110 vdd.n302 vdd.n301 9.3005
R5111 vdd.n313 vdd.n312 9.3005
R5112 vdd.n315 vdd.n314 9.3005
R5113 vdd.n298 vdd.n297 9.3005
R5114 vdd.n321 vdd.n320 9.3005
R5115 vdd.n323 vdd.n322 9.3005
R5116 vdd.n295 vdd.n292 9.3005
R5117 vdd.n330 vdd.n329 9.3005
R5118 vdd.n248 vdd.n247 9.3005
R5119 vdd.n243 vdd.n242 9.3005
R5120 vdd.n254 vdd.n253 9.3005
R5121 vdd.n256 vdd.n255 9.3005
R5122 vdd.n239 vdd.n238 9.3005
R5123 vdd.n262 vdd.n261 9.3005
R5124 vdd.n264 vdd.n263 9.3005
R5125 vdd.n236 vdd.n233 9.3005
R5126 vdd.n271 vdd.n270 9.3005
R5127 vdd.n205 vdd.n204 9.3005
R5128 vdd.n200 vdd.n199 9.3005
R5129 vdd.n211 vdd.n210 9.3005
R5130 vdd.n213 vdd.n212 9.3005
R5131 vdd.n196 vdd.n195 9.3005
R5132 vdd.n219 vdd.n218 9.3005
R5133 vdd.n221 vdd.n220 9.3005
R5134 vdd.n193 vdd.n190 9.3005
R5135 vdd.n228 vdd.n227 9.3005
R5136 vdd.n146 vdd.n145 9.3005
R5137 vdd.n141 vdd.n140 9.3005
R5138 vdd.n152 vdd.n151 9.3005
R5139 vdd.n154 vdd.n153 9.3005
R5140 vdd.n137 vdd.n136 9.3005
R5141 vdd.n160 vdd.n159 9.3005
R5142 vdd.n162 vdd.n161 9.3005
R5143 vdd.n134 vdd.n131 9.3005
R5144 vdd.n169 vdd.n168 9.3005
R5145 vdd.n104 vdd.n103 9.3005
R5146 vdd.n99 vdd.n98 9.3005
R5147 vdd.n110 vdd.n109 9.3005
R5148 vdd.n112 vdd.n111 9.3005
R5149 vdd.n95 vdd.n94 9.3005
R5150 vdd.n118 vdd.n117 9.3005
R5151 vdd.n120 vdd.n119 9.3005
R5152 vdd.n92 vdd.n89 9.3005
R5153 vdd.n127 vdd.n126 9.3005
R5154 vdd.n45 vdd.n44 9.3005
R5155 vdd.n40 vdd.n39 9.3005
R5156 vdd.n51 vdd.n50 9.3005
R5157 vdd.n53 vdd.n52 9.3005
R5158 vdd.n36 vdd.n35 9.3005
R5159 vdd.n59 vdd.n58 9.3005
R5160 vdd.n61 vdd.n60 9.3005
R5161 vdd.n33 vdd.n30 9.3005
R5162 vdd.n68 vdd.n67 9.3005
R5163 vdd.n3230 vdd.n3229 9.3005
R5164 vdd.n3233 vdd.n766 9.3005
R5165 vdd.n3234 vdd.n765 9.3005
R5166 vdd.n3237 vdd.n764 9.3005
R5167 vdd.n3238 vdd.n763 9.3005
R5168 vdd.n3241 vdd.n762 9.3005
R5169 vdd.n3242 vdd.n761 9.3005
R5170 vdd.n3245 vdd.n760 9.3005
R5171 vdd.n3246 vdd.n759 9.3005
R5172 vdd.n3249 vdd.n758 9.3005
R5173 vdd.n3250 vdd.n757 9.3005
R5174 vdd.n3253 vdd.n756 9.3005
R5175 vdd.n3254 vdd.n755 9.3005
R5176 vdd.n3257 vdd.n754 9.3005
R5177 vdd.n3258 vdd.n753 9.3005
R5178 vdd.n3261 vdd.n752 9.3005
R5179 vdd.n3262 vdd.n751 9.3005
R5180 vdd.n3265 vdd.n750 9.3005
R5181 vdd.n3266 vdd.n749 9.3005
R5182 vdd.n3269 vdd.n748 9.3005
R5183 vdd.n3273 vdd.n3272 9.3005
R5184 vdd.n3274 vdd.n747 9.3005
R5185 vdd.n3278 vdd.n3275 9.3005
R5186 vdd.n3281 vdd.n746 9.3005
R5187 vdd.n3282 vdd.n745 9.3005
R5188 vdd.n3285 vdd.n744 9.3005
R5189 vdd.n3286 vdd.n743 9.3005
R5190 vdd.n3289 vdd.n742 9.3005
R5191 vdd.n3290 vdd.n741 9.3005
R5192 vdd.n3293 vdd.n740 9.3005
R5193 vdd.n3294 vdd.n739 9.3005
R5194 vdd.n3297 vdd.n738 9.3005
R5195 vdd.n3298 vdd.n737 9.3005
R5196 vdd.n3301 vdd.n736 9.3005
R5197 vdd.n3302 vdd.n735 9.3005
R5198 vdd.n3305 vdd.n730 9.3005
R5199 vdd.n3311 vdd.n727 9.3005
R5200 vdd.n3312 vdd.n726 9.3005
R5201 vdd.n3326 vdd.n3325 9.3005
R5202 vdd.n3327 vdd.n681 9.3005
R5203 vdd.n3329 vdd.n3328 9.3005
R5204 vdd.n671 vdd.n670 9.3005
R5205 vdd.n3343 vdd.n3342 9.3005
R5206 vdd.n3344 vdd.n669 9.3005
R5207 vdd.n3346 vdd.n3345 9.3005
R5208 vdd.n660 vdd.n659 9.3005
R5209 vdd.n3359 vdd.n3358 9.3005
R5210 vdd.n3360 vdd.n658 9.3005
R5211 vdd.n3362 vdd.n3361 9.3005
R5212 vdd.n648 vdd.n647 9.3005
R5213 vdd.n3376 vdd.n3375 9.3005
R5214 vdd.n3377 vdd.n646 9.3005
R5215 vdd.n3379 vdd.n3378 9.3005
R5216 vdd.n637 vdd.n636 9.3005
R5217 vdd.n3395 vdd.n3394 9.3005
R5218 vdd.n3396 vdd.n635 9.3005
R5219 vdd.n3398 vdd.n3397 9.3005
R5220 vdd.n336 vdd.n334 9.3005
R5221 vdd.n683 vdd.n682 9.3005
R5222 vdd.n3490 vdd.n3489 9.3005
R5223 vdd.n337 vdd.n335 9.3005
R5224 vdd.n3483 vdd.n346 9.3005
R5225 vdd.n3482 vdd.n347 9.3005
R5226 vdd.n3481 vdd.n348 9.3005
R5227 vdd.n355 vdd.n349 9.3005
R5228 vdd.n3475 vdd.n356 9.3005
R5229 vdd.n3474 vdd.n357 9.3005
R5230 vdd.n3473 vdd.n358 9.3005
R5231 vdd.n366 vdd.n359 9.3005
R5232 vdd.n3467 vdd.n367 9.3005
R5233 vdd.n3466 vdd.n368 9.3005
R5234 vdd.n3465 vdd.n369 9.3005
R5235 vdd.n377 vdd.n370 9.3005
R5236 vdd.n3459 vdd.n378 9.3005
R5237 vdd.n3458 vdd.n379 9.3005
R5238 vdd.n3457 vdd.n380 9.3005
R5239 vdd.n388 vdd.n381 9.3005
R5240 vdd.n3451 vdd.n389 9.3005
R5241 vdd.n3450 vdd.n390 9.3005
R5242 vdd.n3449 vdd.n391 9.3005
R5243 vdd.n466 vdd.n463 9.3005
R5244 vdd.n470 vdd.n469 9.3005
R5245 vdd.n471 vdd.n462 9.3005
R5246 vdd.n475 vdd.n472 9.3005
R5247 vdd.n476 vdd.n461 9.3005
R5248 vdd.n480 vdd.n479 9.3005
R5249 vdd.n481 vdd.n460 9.3005
R5250 vdd.n485 vdd.n482 9.3005
R5251 vdd.n486 vdd.n459 9.3005
R5252 vdd.n490 vdd.n489 9.3005
R5253 vdd.n491 vdd.n458 9.3005
R5254 vdd.n495 vdd.n492 9.3005
R5255 vdd.n496 vdd.n457 9.3005
R5256 vdd.n500 vdd.n499 9.3005
R5257 vdd.n501 vdd.n456 9.3005
R5258 vdd.n505 vdd.n502 9.3005
R5259 vdd.n506 vdd.n455 9.3005
R5260 vdd.n510 vdd.n509 9.3005
R5261 vdd.n511 vdd.n454 9.3005
R5262 vdd.n515 vdd.n512 9.3005
R5263 vdd.n516 vdd.n451 9.3005
R5264 vdd.n520 vdd.n519 9.3005
R5265 vdd.n521 vdd.n450 9.3005
R5266 vdd.n525 vdd.n522 9.3005
R5267 vdd.n526 vdd.n449 9.3005
R5268 vdd.n530 vdd.n529 9.3005
R5269 vdd.n531 vdd.n448 9.3005
R5270 vdd.n535 vdd.n532 9.3005
R5271 vdd.n536 vdd.n447 9.3005
R5272 vdd.n540 vdd.n539 9.3005
R5273 vdd.n541 vdd.n446 9.3005
R5274 vdd.n545 vdd.n542 9.3005
R5275 vdd.n546 vdd.n445 9.3005
R5276 vdd.n550 vdd.n549 9.3005
R5277 vdd.n551 vdd.n444 9.3005
R5278 vdd.n555 vdd.n552 9.3005
R5279 vdd.n556 vdd.n443 9.3005
R5280 vdd.n560 vdd.n559 9.3005
R5281 vdd.n561 vdd.n442 9.3005
R5282 vdd.n565 vdd.n562 9.3005
R5283 vdd.n566 vdd.n439 9.3005
R5284 vdd.n570 vdd.n569 9.3005
R5285 vdd.n571 vdd.n438 9.3005
R5286 vdd.n575 vdd.n572 9.3005
R5287 vdd.n576 vdd.n437 9.3005
R5288 vdd.n580 vdd.n579 9.3005
R5289 vdd.n581 vdd.n436 9.3005
R5290 vdd.n585 vdd.n582 9.3005
R5291 vdd.n586 vdd.n435 9.3005
R5292 vdd.n590 vdd.n589 9.3005
R5293 vdd.n591 vdd.n434 9.3005
R5294 vdd.n595 vdd.n592 9.3005
R5295 vdd.n596 vdd.n433 9.3005
R5296 vdd.n600 vdd.n599 9.3005
R5297 vdd.n601 vdd.n432 9.3005
R5298 vdd.n605 vdd.n602 9.3005
R5299 vdd.n606 vdd.n431 9.3005
R5300 vdd.n610 vdd.n609 9.3005
R5301 vdd.n611 vdd.n430 9.3005
R5302 vdd.n615 vdd.n612 9.3005
R5303 vdd.n617 vdd.n429 9.3005
R5304 vdd.n619 vdd.n618 9.3005
R5305 vdd.n3443 vdd.n3442 9.3005
R5306 vdd.n465 vdd.n464 9.3005
R5307 vdd.n3321 vdd.n3320 9.3005
R5308 vdd.n676 vdd.n675 9.3005
R5309 vdd.n3334 vdd.n3333 9.3005
R5310 vdd.n3335 vdd.n674 9.3005
R5311 vdd.n3337 vdd.n3336 9.3005
R5312 vdd.n666 vdd.n665 9.3005
R5313 vdd.n3351 vdd.n3350 9.3005
R5314 vdd.n3352 vdd.n664 9.3005
R5315 vdd.n3354 vdd.n3353 9.3005
R5316 vdd.n653 vdd.n652 9.3005
R5317 vdd.n3367 vdd.n3366 9.3005
R5318 vdd.n3368 vdd.n651 9.3005
R5319 vdd.n3370 vdd.n3369 9.3005
R5320 vdd.n642 vdd.n641 9.3005
R5321 vdd.n3384 vdd.n3383 9.3005
R5322 vdd.n3385 vdd.n640 9.3005
R5323 vdd.n3390 vdd.n3386 9.3005
R5324 vdd.n3389 vdd.n3388 9.3005
R5325 vdd.n3387 vdd.n631 9.3005
R5326 vdd.n3403 vdd.n630 9.3005
R5327 vdd.n3405 vdd.n3404 9.3005
R5328 vdd.n3406 vdd.n629 9.3005
R5329 vdd.n3408 vdd.n3407 9.3005
R5330 vdd.n3410 vdd.n628 9.3005
R5331 vdd.n3412 vdd.n3411 9.3005
R5332 vdd.n3413 vdd.n627 9.3005
R5333 vdd.n3415 vdd.n3414 9.3005
R5334 vdd.n3417 vdd.n626 9.3005
R5335 vdd.n3419 vdd.n3418 9.3005
R5336 vdd.n3420 vdd.n625 9.3005
R5337 vdd.n3422 vdd.n3421 9.3005
R5338 vdd.n3425 vdd.n624 9.3005
R5339 vdd.n3427 vdd.n3426 9.3005
R5340 vdd.n3428 vdd.n623 9.3005
R5341 vdd.n3430 vdd.n3429 9.3005
R5342 vdd.n3432 vdd.n622 9.3005
R5343 vdd.n3434 vdd.n3433 9.3005
R5344 vdd.n3435 vdd.n621 9.3005
R5345 vdd.n3437 vdd.n3436 9.3005
R5346 vdd.n3439 vdd.n620 9.3005
R5347 vdd.n3441 vdd.n3440 9.3005
R5348 vdd.n3319 vdd.n686 9.3005
R5349 vdd.n3318 vdd.n3317 9.3005
R5350 vdd.n3187 vdd.n687 9.3005
R5351 vdd.n3196 vdd.n783 9.3005
R5352 vdd.n3199 vdd.n782 9.3005
R5353 vdd.n3200 vdd.n781 9.3005
R5354 vdd.n3203 vdd.n780 9.3005
R5355 vdd.n3204 vdd.n779 9.3005
R5356 vdd.n3207 vdd.n778 9.3005
R5357 vdd.n3208 vdd.n777 9.3005
R5358 vdd.n3211 vdd.n776 9.3005
R5359 vdd.n3212 vdd.n775 9.3005
R5360 vdd.n3215 vdd.n774 9.3005
R5361 vdd.n3216 vdd.n773 9.3005
R5362 vdd.n3219 vdd.n772 9.3005
R5363 vdd.n3220 vdd.n771 9.3005
R5364 vdd.n3223 vdd.n770 9.3005
R5365 vdd.n3227 vdd.n3226 9.3005
R5366 vdd.n3228 vdd.n767 9.3005
R5367 vdd.n2273 vdd.n2272 9.3005
R5368 vdd.n2268 vdd.n1424 9.3005
R5369 vdd.n1792 vdd.n1791 9.3005
R5370 vdd.n1793 vdd.n1547 9.3005
R5371 vdd.n1795 vdd.n1794 9.3005
R5372 vdd.n1537 vdd.n1536 9.3005
R5373 vdd.n1809 vdd.n1808 9.3005
R5374 vdd.n1810 vdd.n1535 9.3005
R5375 vdd.n1812 vdd.n1811 9.3005
R5376 vdd.n1527 vdd.n1526 9.3005
R5377 vdd.n1826 vdd.n1825 9.3005
R5378 vdd.n1827 vdd.n1525 9.3005
R5379 vdd.n1829 vdd.n1828 9.3005
R5380 vdd.n1514 vdd.n1513 9.3005
R5381 vdd.n1842 vdd.n1841 9.3005
R5382 vdd.n1843 vdd.n1512 9.3005
R5383 vdd.n1845 vdd.n1844 9.3005
R5384 vdd.n1503 vdd.n1502 9.3005
R5385 vdd.n1859 vdd.n1858 9.3005
R5386 vdd.n1860 vdd.n1501 9.3005
R5387 vdd.n1862 vdd.n1861 9.3005
R5388 vdd.n1492 vdd.n1491 9.3005
R5389 vdd.n2182 vdd.n2181 9.3005
R5390 vdd.n2183 vdd.n1490 9.3005
R5391 vdd.n2185 vdd.n2184 9.3005
R5392 vdd.n1480 vdd.n1479 9.3005
R5393 vdd.n2199 vdd.n2198 9.3005
R5394 vdd.n2200 vdd.n1478 9.3005
R5395 vdd.n2202 vdd.n2201 9.3005
R5396 vdd.n1470 vdd.n1469 9.3005
R5397 vdd.n2216 vdd.n2215 9.3005
R5398 vdd.n2217 vdd.n1468 9.3005
R5399 vdd.n2219 vdd.n2218 9.3005
R5400 vdd.n1457 vdd.n1456 9.3005
R5401 vdd.n2232 vdd.n2231 9.3005
R5402 vdd.n2233 vdd.n1455 9.3005
R5403 vdd.n2235 vdd.n2234 9.3005
R5404 vdd.n1447 vdd.n1446 9.3005
R5405 vdd.n2249 vdd.n2248 9.3005
R5406 vdd.n2250 vdd.n1444 9.3005
R5407 vdd.n2254 vdd.n2253 9.3005
R5408 vdd.n2252 vdd.n1445 9.3005
R5409 vdd.n2251 vdd.n1435 9.3005
R5410 vdd.n1549 vdd.n1548 9.3005
R5411 vdd.n1685 vdd.n1684 9.3005
R5412 vdd.n1686 vdd.n1675 9.3005
R5413 vdd.n1688 vdd.n1687 9.3005
R5414 vdd.n1689 vdd.n1674 9.3005
R5415 vdd.n1691 vdd.n1690 9.3005
R5416 vdd.n1692 vdd.n1669 9.3005
R5417 vdd.n1694 vdd.n1693 9.3005
R5418 vdd.n1695 vdd.n1668 9.3005
R5419 vdd.n1697 vdd.n1696 9.3005
R5420 vdd.n1698 vdd.n1663 9.3005
R5421 vdd.n1700 vdd.n1699 9.3005
R5422 vdd.n1701 vdd.n1662 9.3005
R5423 vdd.n1703 vdd.n1702 9.3005
R5424 vdd.n1704 vdd.n1657 9.3005
R5425 vdd.n1706 vdd.n1705 9.3005
R5426 vdd.n1707 vdd.n1656 9.3005
R5427 vdd.n1709 vdd.n1708 9.3005
R5428 vdd.n1710 vdd.n1651 9.3005
R5429 vdd.n1712 vdd.n1711 9.3005
R5430 vdd.n1713 vdd.n1650 9.3005
R5431 vdd.n1715 vdd.n1714 9.3005
R5432 vdd.n1719 vdd.n1646 9.3005
R5433 vdd.n1721 vdd.n1720 9.3005
R5434 vdd.n1722 vdd.n1645 9.3005
R5435 vdd.n1724 vdd.n1723 9.3005
R5436 vdd.n1725 vdd.n1640 9.3005
R5437 vdd.n1727 vdd.n1726 9.3005
R5438 vdd.n1728 vdd.n1639 9.3005
R5439 vdd.n1730 vdd.n1729 9.3005
R5440 vdd.n1731 vdd.n1634 9.3005
R5441 vdd.n1733 vdd.n1732 9.3005
R5442 vdd.n1734 vdd.n1633 9.3005
R5443 vdd.n1736 vdd.n1735 9.3005
R5444 vdd.n1737 vdd.n1628 9.3005
R5445 vdd.n1739 vdd.n1738 9.3005
R5446 vdd.n1740 vdd.n1627 9.3005
R5447 vdd.n1742 vdd.n1741 9.3005
R5448 vdd.n1743 vdd.n1622 9.3005
R5449 vdd.n1745 vdd.n1744 9.3005
R5450 vdd.n1746 vdd.n1621 9.3005
R5451 vdd.n1748 vdd.n1747 9.3005
R5452 vdd.n1749 vdd.n1616 9.3005
R5453 vdd.n1751 vdd.n1750 9.3005
R5454 vdd.n1752 vdd.n1615 9.3005
R5455 vdd.n1754 vdd.n1753 9.3005
R5456 vdd.n1755 vdd.n1608 9.3005
R5457 vdd.n1757 vdd.n1756 9.3005
R5458 vdd.n1758 vdd.n1607 9.3005
R5459 vdd.n1760 vdd.n1759 9.3005
R5460 vdd.n1761 vdd.n1602 9.3005
R5461 vdd.n1763 vdd.n1762 9.3005
R5462 vdd.n1764 vdd.n1601 9.3005
R5463 vdd.n1766 vdd.n1765 9.3005
R5464 vdd.n1767 vdd.n1596 9.3005
R5465 vdd.n1769 vdd.n1768 9.3005
R5466 vdd.n1770 vdd.n1595 9.3005
R5467 vdd.n1772 vdd.n1771 9.3005
R5468 vdd.n1773 vdd.n1590 9.3005
R5469 vdd.n1775 vdd.n1774 9.3005
R5470 vdd.n1776 vdd.n1589 9.3005
R5471 vdd.n1778 vdd.n1777 9.3005
R5472 vdd.n1554 vdd.n1553 9.3005
R5473 vdd.n1784 vdd.n1783 9.3005
R5474 vdd.n1683 vdd.n1682 9.3005
R5475 vdd.n1787 vdd.n1786 9.3005
R5476 vdd.n1543 vdd.n1542 9.3005
R5477 vdd.n1801 vdd.n1800 9.3005
R5478 vdd.n1802 vdd.n1541 9.3005
R5479 vdd.n1804 vdd.n1803 9.3005
R5480 vdd.n1532 vdd.n1531 9.3005
R5481 vdd.n1818 vdd.n1817 9.3005
R5482 vdd.n1819 vdd.n1530 9.3005
R5483 vdd.n1821 vdd.n1820 9.3005
R5484 vdd.n1521 vdd.n1520 9.3005
R5485 vdd.n1834 vdd.n1833 9.3005
R5486 vdd.n1835 vdd.n1519 9.3005
R5487 vdd.n1837 vdd.n1836 9.3005
R5488 vdd.n1509 vdd.n1508 9.3005
R5489 vdd.n1851 vdd.n1850 9.3005
R5490 vdd.n1852 vdd.n1507 9.3005
R5491 vdd.n1854 vdd.n1853 9.3005
R5492 vdd.n1498 vdd.n1497 9.3005
R5493 vdd.n1867 vdd.n1866 9.3005
R5494 vdd.n1868 vdd.n1496 9.3005
R5495 vdd.n1785 vdd.n1552 9.3005
R5496 vdd.n2088 vdd.n2087 9.3005
R5497 vdd.n2083 vdd.n2082 9.3005
R5498 vdd.n2094 vdd.n2093 9.3005
R5499 vdd.n2096 vdd.n2095 9.3005
R5500 vdd.n2079 vdd.n2078 9.3005
R5501 vdd.n2102 vdd.n2101 9.3005
R5502 vdd.n2104 vdd.n2103 9.3005
R5503 vdd.n2076 vdd.n2073 9.3005
R5504 vdd.n2111 vdd.n2110 9.3005
R5505 vdd.n2147 vdd.n2146 9.3005
R5506 vdd.n2142 vdd.n2141 9.3005
R5507 vdd.n2153 vdd.n2152 9.3005
R5508 vdd.n2155 vdd.n2154 9.3005
R5509 vdd.n2138 vdd.n2137 9.3005
R5510 vdd.n2161 vdd.n2160 9.3005
R5511 vdd.n2163 vdd.n2162 9.3005
R5512 vdd.n2135 vdd.n2132 9.3005
R5513 vdd.n2170 vdd.n2169 9.3005
R5514 vdd.n1986 vdd.n1985 9.3005
R5515 vdd.n1981 vdd.n1980 9.3005
R5516 vdd.n1992 vdd.n1991 9.3005
R5517 vdd.n1994 vdd.n1993 9.3005
R5518 vdd.n1977 vdd.n1976 9.3005
R5519 vdd.n2000 vdd.n1999 9.3005
R5520 vdd.n2002 vdd.n2001 9.3005
R5521 vdd.n1974 vdd.n1971 9.3005
R5522 vdd.n2009 vdd.n2008 9.3005
R5523 vdd.n2045 vdd.n2044 9.3005
R5524 vdd.n2040 vdd.n2039 9.3005
R5525 vdd.n2051 vdd.n2050 9.3005
R5526 vdd.n2053 vdd.n2052 9.3005
R5527 vdd.n2036 vdd.n2035 9.3005
R5528 vdd.n2059 vdd.n2058 9.3005
R5529 vdd.n2061 vdd.n2060 9.3005
R5530 vdd.n2033 vdd.n2030 9.3005
R5531 vdd.n2068 vdd.n2067 9.3005
R5532 vdd.n1885 vdd.n1884 9.3005
R5533 vdd.n1880 vdd.n1879 9.3005
R5534 vdd.n1891 vdd.n1890 9.3005
R5535 vdd.n1893 vdd.n1892 9.3005
R5536 vdd.n1876 vdd.n1875 9.3005
R5537 vdd.n1899 vdd.n1898 9.3005
R5538 vdd.n1901 vdd.n1900 9.3005
R5539 vdd.n1873 vdd.n1870 9.3005
R5540 vdd.n1908 vdd.n1907 9.3005
R5541 vdd.n1944 vdd.n1943 9.3005
R5542 vdd.n1939 vdd.n1938 9.3005
R5543 vdd.n1950 vdd.n1949 9.3005
R5544 vdd.n1952 vdd.n1951 9.3005
R5545 vdd.n1935 vdd.n1934 9.3005
R5546 vdd.n1958 vdd.n1957 9.3005
R5547 vdd.n1960 vdd.n1959 9.3005
R5548 vdd.n1932 vdd.n1929 9.3005
R5549 vdd.n1967 vdd.n1966 9.3005
R5550 vdd.n1823 vdd.t132 9.18308
R5551 vdd.n3423 vdd.t70 9.18308
R5552 vdd.n1517 vdd.t107 8.95635
R5553 vdd.n2265 vdd.t237 8.95635
R5554 vdd.n723 vdd.t233 8.95635
R5555 vdd.t85 vdd.n3477 8.95635
R5556 vdd.n312 vdd.n311 8.92171
R5557 vdd.n253 vdd.n252 8.92171
R5558 vdd.n210 vdd.n209 8.92171
R5559 vdd.n151 vdd.n150 8.92171
R5560 vdd.n109 vdd.n108 8.92171
R5561 vdd.n50 vdd.n49 8.92171
R5562 vdd.n2093 vdd.n2092 8.92171
R5563 vdd.n2152 vdd.n2151 8.92171
R5564 vdd.n1991 vdd.n1990 8.92171
R5565 vdd.n2050 vdd.n2049 8.92171
R5566 vdd.n1890 vdd.n1889 8.92171
R5567 vdd.n1949 vdd.n1948 8.92171
R5568 vdd.n231 vdd.n129 8.81535
R5569 vdd.n2071 vdd.n1969 8.81535
R5570 vdd.n1864 vdd.t162 8.72962
R5571 vdd.t89 vdd.n3486 8.72962
R5572 vdd.n2187 vdd.t94 8.50289
R5573 vdd.n3392 vdd.t91 8.50289
R5574 vdd.n28 vdd.n14 8.42249
R5575 vdd.n2213 vdd.t165 8.27616
R5576 vdd.t126 vdd.n656 8.27616
R5577 vdd.n3492 vdd.n3491 8.16225
R5578 vdd.n2175 vdd.n2174 8.16225
R5579 vdd.n308 vdd.n302 8.14595
R5580 vdd.n249 vdd.n243 8.14595
R5581 vdd.n206 vdd.n200 8.14595
R5582 vdd.n147 vdd.n141 8.14595
R5583 vdd.n105 vdd.n99 8.14595
R5584 vdd.n46 vdd.n40 8.14595
R5585 vdd.n2089 vdd.n2083 8.14595
R5586 vdd.n2148 vdd.n2142 8.14595
R5587 vdd.n1987 vdd.n1981 8.14595
R5588 vdd.n2046 vdd.n2040 8.14595
R5589 vdd.n1886 vdd.n1880 8.14595
R5590 vdd.n1945 vdd.n1939 8.14595
R5591 vdd.n1460 vdd.t76 8.04943
R5592 vdd.n3348 vdd.t184 8.04943
R5593 vdd.n2424 vdd.n1076 7.70933
R5594 vdd.n2424 vdd.n1079 7.70933
R5595 vdd.n2430 vdd.n1065 7.70933
R5596 vdd.n2436 vdd.n1065 7.70933
R5597 vdd.n2436 vdd.n1059 7.70933
R5598 vdd.n2442 vdd.n1059 7.70933
R5599 vdd.n2448 vdd.n1052 7.70933
R5600 vdd.n2448 vdd.n1055 7.70933
R5601 vdd.n2454 vdd.n1048 7.70933
R5602 vdd.n2461 vdd.n1034 7.70933
R5603 vdd.n2467 vdd.n1034 7.70933
R5604 vdd.n2473 vdd.n1028 7.70933
R5605 vdd.n2479 vdd.n1024 7.70933
R5606 vdd.n2485 vdd.n1018 7.70933
R5607 vdd.n2497 vdd.n1005 7.70933
R5608 vdd.n2503 vdd.n999 7.70933
R5609 vdd.n2503 vdd.n992 7.70933
R5610 vdd.n2511 vdd.n992 7.70933
R5611 vdd.n2593 vdd.n976 7.70933
R5612 vdd.n2945 vdd.n928 7.70933
R5613 vdd.n2957 vdd.n917 7.70933
R5614 vdd.n2957 vdd.n911 7.70933
R5615 vdd.n2963 vdd.n911 7.70933
R5616 vdd.n2969 vdd.n905 7.70933
R5617 vdd.n2975 vdd.n901 7.70933
R5618 vdd.n2981 vdd.n895 7.70933
R5619 vdd.n2993 vdd.n882 7.70933
R5620 vdd.n2999 vdd.n875 7.70933
R5621 vdd.n2999 vdd.n878 7.70933
R5622 vdd.n3006 vdd.n870 7.70933
R5623 vdd.n3012 vdd.n857 7.70933
R5624 vdd.n3018 vdd.n857 7.70933
R5625 vdd.n3024 vdd.n851 7.70933
R5626 vdd.n3024 vdd.n843 7.70933
R5627 vdd.n3075 vdd.n843 7.70933
R5628 vdd.n3075 vdd.n846 7.70933
R5629 vdd.n3081 vdd.n805 7.70933
R5630 vdd.n3151 vdd.n805 7.70933
R5631 vdd.n3004 vdd.n3003 7.49318
R5632 vdd.n2458 vdd.n2457 7.49318
R5633 vdd.n307 vdd.n304 7.3702
R5634 vdd.n248 vdd.n245 7.3702
R5635 vdd.n205 vdd.n202 7.3702
R5636 vdd.n146 vdd.n143 7.3702
R5637 vdd.n104 vdd.n101 7.3702
R5638 vdd.n45 vdd.n42 7.3702
R5639 vdd.n2088 vdd.n2085 7.3702
R5640 vdd.n2147 vdd.n2144 7.3702
R5641 vdd.n1986 vdd.n1983 7.3702
R5642 vdd.n2045 vdd.n2042 7.3702
R5643 vdd.n1885 vdd.n1882 7.3702
R5644 vdd.n1944 vdd.n1941 7.3702
R5645 vdd.n2442 vdd.t45 7.36923
R5646 vdd.t8 vdd.n851 7.36923
R5647 vdd.n2518 vdd.t15 7.25587
R5648 vdd.n2862 vdd.t35 7.25587
R5649 vdd.n2246 vdd.t114 7.1425
R5650 vdd.n679 vdd.t112 7.1425
R5651 vdd.n1720 vdd.n1719 6.98232
R5652 vdd.n2308 vdd.n2307 6.98232
R5653 vdd.n566 vdd.n565 6.98232
R5654 vdd.n3233 vdd.n3230 6.98232
R5655 vdd.t178 vdd.n1459 6.91577
R5656 vdd.n3356 vdd.t124 6.91577
R5657 vdd.n2205 vdd.t130 6.68904
R5658 vdd.n3372 vdd.t74 6.68904
R5659 vdd.t160 vdd.n1488 6.46231
R5660 vdd.n3400 vdd.t118 6.46231
R5661 vdd.n3492 vdd.n333 6.38151
R5662 vdd.n2174 vdd.n2173 6.38151
R5663 vdd.n1856 vdd.t105 6.23558
R5664 vdd.t175 vdd.n344 6.23558
R5665 vdd.t80 vdd.n1516 6.00885
R5666 vdd.n3471 vdd.t135 6.00885
R5667 vdd.t25 vdd.n1005 5.89549
R5668 vdd.n2969 vdd.t0 5.89549
R5669 vdd.n308 vdd.n307 5.81868
R5670 vdd.n249 vdd.n248 5.81868
R5671 vdd.n206 vdd.n205 5.81868
R5672 vdd.n147 vdd.n146 5.81868
R5673 vdd.n105 vdd.n104 5.81868
R5674 vdd.n46 vdd.n45 5.81868
R5675 vdd.n2089 vdd.n2088 5.81868
R5676 vdd.n2148 vdd.n2147 5.81868
R5677 vdd.n1987 vdd.n1986 5.81868
R5678 vdd.n2046 vdd.n2045 5.81868
R5679 vdd.n1886 vdd.n1885 5.81868
R5680 vdd.n1945 vdd.n1944 5.81868
R5681 vdd.n1815 vdd.t62 5.78212
R5682 vdd.n3462 vdd.t181 5.78212
R5683 vdd.n2601 vdd.n2600 5.77611
R5684 vdd.n1303 vdd.n1302 5.77611
R5685 vdd.n2874 vdd.n2873 5.77611
R5686 vdd.n3092 vdd.n3091 5.77611
R5687 vdd.n3156 vdd.n801 5.77611
R5688 vdd.n2768 vdd.n2706 5.77611
R5689 vdd.n2526 vdd.n983 5.77611
R5690 vdd.n1392 vdd.n1255 5.77611
R5691 vdd.n1682 vdd.n1681 5.62474
R5692 vdd.n2271 vdd.n2268 5.62474
R5693 vdd.n3443 vdd.n428 5.62474
R5694 vdd.n3317 vdd.n690 5.62474
R5695 vdd.n1539 vdd.t62 5.55539
R5696 vdd.t14 vdd.n1028 5.55539
R5697 vdd.n2473 vdd.t21 5.55539
R5698 vdd.t44 vdd.n882 5.55539
R5699 vdd.n2993 vdd.t22 5.55539
R5700 vdd.t181 vdd.n3461 5.55539
R5701 vdd.n1048 vdd.t282 5.44203
R5702 vdd.n3006 vdd.t251 5.44203
R5703 vdd.n1831 vdd.t80 5.32866
R5704 vdd.n2430 vdd.t229 5.32866
R5705 vdd.n1338 vdd.t271 5.32866
R5706 vdd.n2951 vdd.t275 5.32866
R5707 vdd.n846 vdd.t225 5.32866
R5708 vdd.t135 vdd.n3470 5.32866
R5709 vdd.n1847 vdd.t105 5.10193
R5710 vdd.n3479 vdd.t175 5.10193
R5711 vdd.n311 vdd.n302 5.04292
R5712 vdd.n252 vdd.n243 5.04292
R5713 vdd.n209 vdd.n200 5.04292
R5714 vdd.n150 vdd.n141 5.04292
R5715 vdd.n108 vdd.n99 5.04292
R5716 vdd.n49 vdd.n40 5.04292
R5717 vdd.n2092 vdd.n2083 5.04292
R5718 vdd.n2151 vdd.n2142 5.04292
R5719 vdd.n1990 vdd.n1981 5.04292
R5720 vdd.n2049 vdd.n2040 5.04292
R5721 vdd.n1889 vdd.n1880 5.04292
R5722 vdd.n1948 vdd.n1939 5.04292
R5723 vdd.n2479 vdd.t2 4.98857
R5724 vdd.n895 vdd.t30 4.98857
R5725 vdd.n2179 vdd.t160 4.8752
R5726 vdd.t7 vdd.t41 4.8752
R5727 vdd.t9 vdd.t33 4.8752
R5728 vdd.t12 vdd.t20 4.8752
R5729 vdd.t49 vdd.t51 4.8752
R5730 vdd.t118 vdd.n340 4.8752
R5731 vdd.n2602 vdd.n2601 4.83952
R5732 vdd.n1302 vdd.n1301 4.83952
R5733 vdd.n2875 vdd.n2874 4.83952
R5734 vdd.n3093 vdd.n3092 4.83952
R5735 vdd.n801 vdd.n796 4.83952
R5736 vdd.n2765 vdd.n2706 4.83952
R5737 vdd.n2529 vdd.n983 4.83952
R5738 vdd.n1395 vdd.n1255 4.83952
R5739 vdd.n2276 vdd.n2275 4.74817
R5740 vdd.n1428 vdd.n1423 4.74817
R5741 vdd.n1125 vdd.n1122 4.74817
R5742 vdd.n2369 vdd.n1121 4.74817
R5743 vdd.n2374 vdd.n1122 4.74817
R5744 vdd.n2373 vdd.n1121 4.74817
R5745 vdd.n3310 vdd.n3309 4.74817
R5746 vdd.n3307 vdd.n3306 4.74817
R5747 vdd.n3307 vdd.n732 4.74817
R5748 vdd.n3309 vdd.n729 4.74817
R5749 vdd.n3192 vdd.n784 4.74817
R5750 vdd.n3188 vdd.n3186 4.74817
R5751 vdd.n3191 vdd.n3186 4.74817
R5752 vdd.n3195 vdd.n784 4.74817
R5753 vdd.n2275 vdd.n1221 4.74817
R5754 vdd.n1425 vdd.n1423 4.74817
R5755 vdd.n333 vdd.n332 4.7074
R5756 vdd.n231 vdd.n230 4.7074
R5757 vdd.n2173 vdd.n2172 4.7074
R5758 vdd.n2071 vdd.n2070 4.7074
R5759 vdd.n1482 vdd.t130 4.64847
R5760 vdd.n2454 vdd.t48 4.64847
R5761 vdd.n1018 vdd.t43 4.64847
R5762 vdd.n2975 vdd.t59 4.64847
R5763 vdd.n870 vdd.t27 4.64847
R5764 vdd.n3381 vdd.t74 4.64847
R5765 vdd.n2221 vdd.t178 4.42174
R5766 vdd.t124 vdd.n655 4.42174
R5767 vdd.n312 vdd.n300 4.26717
R5768 vdd.n253 vdd.n241 4.26717
R5769 vdd.n210 vdd.n198 4.26717
R5770 vdd.n151 vdd.n139 4.26717
R5771 vdd.n109 vdd.n97 4.26717
R5772 vdd.n50 vdd.n38 4.26717
R5773 vdd.n2093 vdd.n2081 4.26717
R5774 vdd.n2152 vdd.n2140 4.26717
R5775 vdd.n1991 vdd.n1979 4.26717
R5776 vdd.n2050 vdd.n2038 4.26717
R5777 vdd.n1890 vdd.n1878 4.26717
R5778 vdd.n1949 vdd.n1937 4.26717
R5779 vdd.n2237 vdd.t114 4.19501
R5780 vdd.n3340 vdd.t112 4.19501
R5781 vdd.n333 vdd.n231 4.10845
R5782 vdd.n2173 vdd.n2071 4.10845
R5783 vdd.n289 vdd.t146 4.06363
R5784 vdd.n289 vdd.t195 4.06363
R5785 vdd.n287 vdd.t197 4.06363
R5786 vdd.n287 vdd.t71 4.06363
R5787 vdd.n285 vdd.t104 4.06363
R5788 vdd.n285 vdd.t169 4.06363
R5789 vdd.n283 vdd.t201 4.06363
R5790 vdd.n283 vdd.t212 4.06363
R5791 vdd.n281 vdd.t217 4.06363
R5792 vdd.n281 vdd.t111 4.06363
R5793 vdd.n279 vdd.t140 4.06363
R5794 vdd.n279 vdd.t216 4.06363
R5795 vdd.n277 vdd.t218 4.06363
R5796 vdd.n277 vdd.t139 4.06363
R5797 vdd.n275 vdd.t145 4.06363
R5798 vdd.n275 vdd.t148 4.06363
R5799 vdd.n273 vdd.t196 4.06363
R5800 vdd.n273 vdd.t96 4.06363
R5801 vdd.n187 vdd.t123 4.06363
R5802 vdd.n187 vdd.t182 4.06363
R5803 vdd.n185 vdd.t183 4.06363
R5804 vdd.n185 vdd.t214 4.06363
R5805 vdd.n183 vdd.t86 4.06363
R5806 vdd.n183 vdd.t151 4.06363
R5807 vdd.n181 vdd.t188 4.06363
R5808 vdd.n181 vdd.t202 4.06363
R5809 vdd.n179 vdd.t206 4.06363
R5810 vdd.n179 vdd.t90 4.06363
R5811 vdd.n177 vdd.t117 4.06363
R5812 vdd.n177 vdd.t205 4.06363
R5813 vdd.n175 vdd.t207 4.06363
R5814 vdd.n175 vdd.t75 4.06363
R5815 vdd.n173 vdd.t125 4.06363
R5816 vdd.n173 vdd.t127 4.06363
R5817 vdd.n171 vdd.t185 4.06363
R5818 vdd.n171 vdd.t67 4.06363
R5819 vdd.n86 vdd.t157 4.06363
R5820 vdd.n86 vdd.t186 4.06363
R5821 vdd.n84 vdd.t136 4.06363
R5822 vdd.n84 vdd.t208 4.06363
R5823 vdd.n82 vdd.t103 4.06363
R5824 vdd.n82 vdd.t190 4.06363
R5825 vdd.n80 vdd.t98 4.06363
R5826 vdd.n80 vdd.t176 4.06363
R5827 vdd.n78 vdd.t119 4.06363
R5828 vdd.n78 vdd.t203 4.06363
R5829 vdd.n76 vdd.t92 4.06363
R5830 vdd.n76 vdd.t154 4.06363
R5831 vdd.n74 vdd.t79 4.06363
R5832 vdd.n74 vdd.t128 4.06363
R5833 vdd.n72 vdd.t213 4.06363
R5834 vdd.n72 vdd.t194 4.06363
R5835 vdd.n70 vdd.t199 4.06363
R5836 vdd.n70 vdd.t141 4.06363
R5837 vdd.n2113 vdd.t164 4.06363
R5838 vdd.n2113 vdd.t100 4.06363
R5839 vdd.n2115 vdd.t221 4.06363
R5840 vdd.n2115 vdd.t193 4.06363
R5841 vdd.n2117 vdd.t189 4.06363
R5842 vdd.n2117 vdd.t138 4.06363
R5843 vdd.n2119 vdd.t134 4.06363
R5844 vdd.n2119 vdd.t192 4.06363
R5845 vdd.n2121 vdd.t172 4.06363
R5846 vdd.n2121 vdd.t171 4.06363
R5847 vdd.n2123 vdd.t129 4.06363
R5848 vdd.n2123 vdd.t102 4.06363
R5849 vdd.n2125 vdd.t99 4.06363
R5850 vdd.n2125 vdd.t170 4.06363
R5851 vdd.n2127 vdd.t149 4.06363
R5852 vdd.n2127 vdd.t101 4.06363
R5853 vdd.n2129 vdd.t93 4.06363
R5854 vdd.n2129 vdd.t191 4.06363
R5855 vdd.n2011 vdd.t147 4.06363
R5856 vdd.n2011 vdd.t77 4.06363
R5857 vdd.n2013 vdd.t211 4.06363
R5858 vdd.n2013 vdd.t179 4.06363
R5859 vdd.n2015 vdd.t173 4.06363
R5860 vdd.n2015 vdd.t116 4.06363
R5861 vdd.n2017 vdd.t110 4.06363
R5862 vdd.n2017 vdd.t174 4.06363
R5863 vdd.n2019 vdd.t163 4.06363
R5864 vdd.n2019 vdd.t161 4.06363
R5865 vdd.n2021 vdd.t106 4.06363
R5866 vdd.n2021 vdd.t82 4.06363
R5867 vdd.n2023 vdd.t69 4.06363
R5868 vdd.n2023 vdd.t156 4.06363
R5869 vdd.n2025 vdd.t133 4.06363
R5870 vdd.n2025 vdd.t81 4.06363
R5871 vdd.n2027 vdd.t63 4.06363
R5872 vdd.n2027 vdd.t180 4.06363
R5873 vdd.n1910 vdd.t143 4.06363
R5874 vdd.n1910 vdd.t200 4.06363
R5875 vdd.n1912 vdd.t166 4.06363
R5876 vdd.n1912 vdd.t215 4.06363
R5877 vdd.n1914 vdd.t131 4.06363
R5878 vdd.n1914 vdd.t84 4.06363
R5879 vdd.n1916 vdd.t155 4.06363
R5880 vdd.n1916 vdd.t95 4.06363
R5881 vdd.n1918 vdd.t204 4.06363
R5882 vdd.n1918 vdd.t220 4.06363
R5883 vdd.n1920 vdd.t177 4.06363
R5884 vdd.n1920 vdd.t65 4.06363
R5885 vdd.n1922 vdd.t167 4.06363
R5886 vdd.n1922 vdd.t108 4.06363
R5887 vdd.n1924 vdd.t209 4.06363
R5888 vdd.n1924 vdd.t137 4.06363
R5889 vdd.n1926 vdd.t187 4.06363
R5890 vdd.n1926 vdd.t159 4.06363
R5891 vdd.n26 vdd.t40 3.9605
R5892 vdd.n26 vdd.t4 3.9605
R5893 vdd.n23 vdd.t37 3.9605
R5894 vdd.n23 vdd.t54 3.9605
R5895 vdd.n21 vdd.t60 3.9605
R5896 vdd.n21 vdd.t52 3.9605
R5897 vdd.n20 vdd.t6 3.9605
R5898 vdd.n20 vdd.t58 3.9605
R5899 vdd.n15 vdd.t53 3.9605
R5900 vdd.n15 vdd.t57 3.9605
R5901 vdd.n16 vdd.t5 3.9605
R5902 vdd.n16 vdd.t55 3.9605
R5903 vdd.n18 vdd.t61 3.9605
R5904 vdd.n18 vdd.t38 3.9605
R5905 vdd.n25 vdd.t56 3.9605
R5906 vdd.n25 vdd.t39 3.9605
R5907 vdd.n2511 vdd.t23 3.85492
R5908 vdd.n1338 vdd.t23 3.85492
R5909 vdd.n2951 vdd.t28 3.85492
R5910 vdd.t28 vdd.n917 3.85492
R5911 vdd.n7 vdd.t50 3.61217
R5912 vdd.n7 vdd.t31 3.61217
R5913 vdd.n8 vdd.t13 3.61217
R5914 vdd.n8 vdd.t1 3.61217
R5915 vdd.n10 vdd.t36 3.61217
R5916 vdd.n10 vdd.t29 3.61217
R5917 vdd.n12 vdd.t47 3.61217
R5918 vdd.n12 vdd.t223 3.61217
R5919 vdd.n5 vdd.t18 3.61217
R5920 vdd.n5 vdd.t11 3.61217
R5921 vdd.n3 vdd.t24 3.61217
R5922 vdd.n3 vdd.t16 3.61217
R5923 vdd.n1 vdd.t26 3.61217
R5924 vdd.n1 vdd.t34 3.61217
R5925 vdd.n0 vdd.t3 3.61217
R5926 vdd.n0 vdd.t42 3.61217
R5927 vdd.n316 vdd.n315 3.49141
R5928 vdd.n257 vdd.n256 3.49141
R5929 vdd.n214 vdd.n213 3.49141
R5930 vdd.n155 vdd.n154 3.49141
R5931 vdd.n113 vdd.n112 3.49141
R5932 vdd.n54 vdd.n53 3.49141
R5933 vdd.n2097 vdd.n2096 3.49141
R5934 vdd.n2156 vdd.n2155 3.49141
R5935 vdd.n1995 vdd.n1994 3.49141
R5936 vdd.n2054 vdd.n2053 3.49141
R5937 vdd.n1894 vdd.n1893 3.49141
R5938 vdd.n1953 vdd.n1952 3.49141
R5939 vdd.n2665 vdd.t17 3.40145
R5940 vdd.n2938 vdd.t222 3.40145
R5941 vdd.n2238 vdd.t76 3.28809
R5942 vdd.n3339 vdd.t184 3.28809
R5943 vdd.n3003 vdd.n3002 3.12245
R5944 vdd.n2459 vdd.n2458 3.12245
R5945 vdd.t165 vdd.n1466 3.06136
R5946 vdd.n1055 vdd.t48 3.06136
R5947 vdd.n2491 vdd.t43 3.06136
R5948 vdd.n2847 vdd.t59 3.06136
R5949 vdd.n3012 vdd.t27 3.06136
R5950 vdd.n3364 vdd.t126 3.06136
R5951 vdd.n2196 vdd.t94 2.83463
R5952 vdd.n644 vdd.t91 2.83463
R5953 vdd.n1359 vdd.t2 2.72126
R5954 vdd.n2987 vdd.t30 2.72126
R5955 vdd.n319 vdd.n298 2.71565
R5956 vdd.n260 vdd.n239 2.71565
R5957 vdd.n217 vdd.n196 2.71565
R5958 vdd.n158 vdd.n137 2.71565
R5959 vdd.n116 vdd.n95 2.71565
R5960 vdd.n57 vdd.n36 2.71565
R5961 vdd.n2100 vdd.n2079 2.71565
R5962 vdd.n2159 vdd.n2138 2.71565
R5963 vdd.n1998 vdd.n1977 2.71565
R5964 vdd.n2057 vdd.n2036 2.71565
R5965 vdd.n1897 vdd.n1876 2.71565
R5966 vdd.n1956 vdd.n1935 2.71565
R5967 vdd.t162 vdd.n1494 2.6079
R5968 vdd.n3487 vdd.t89 2.6079
R5969 vdd.t33 vdd.n999 2.49453
R5970 vdd.n2963 vdd.t12 2.49453
R5971 vdd.n306 vdd.n305 2.4129
R5972 vdd.n247 vdd.n246 2.4129
R5973 vdd.n204 vdd.n203 2.4129
R5974 vdd.n145 vdd.n144 2.4129
R5975 vdd.n103 vdd.n102 2.4129
R5976 vdd.n44 vdd.n43 2.4129
R5977 vdd.n2087 vdd.n2086 2.4129
R5978 vdd.n2146 vdd.n2145 2.4129
R5979 vdd.n1985 vdd.n1984 2.4129
R5980 vdd.n2044 vdd.n2043 2.4129
R5981 vdd.n1884 vdd.n1883 2.4129
R5982 vdd.n1943 vdd.n1942 2.4129
R5983 vdd.n1848 vdd.t107 2.38117
R5984 vdd.n2256 vdd.t237 2.38117
R5985 vdd.n1079 vdd.t229 2.38117
R5986 vdd.n2518 vdd.t271 2.38117
R5987 vdd.n2862 vdd.t275 2.38117
R5988 vdd.n3081 vdd.t225 2.38117
R5989 vdd.n3323 vdd.t233 2.38117
R5990 vdd.n3478 vdd.t85 2.38117
R5991 vdd.n2381 vdd.n1122 2.27742
R5992 vdd.n2381 vdd.n1121 2.27742
R5993 vdd.n3308 vdd.n3307 2.27742
R5994 vdd.n3309 vdd.n3308 2.27742
R5995 vdd.n3186 vdd.n3185 2.27742
R5996 vdd.n3185 vdd.n784 2.27742
R5997 vdd.n2275 vdd.n2274 2.27742
R5998 vdd.n2274 vdd.n1423 2.27742
R5999 vdd.t132 vdd.n1523 2.15444
R6000 vdd.n2467 vdd.t14 2.15444
R6001 vdd.n1359 vdd.t21 2.15444
R6002 vdd.n2987 vdd.t44 2.15444
R6003 vdd.t22 vdd.n875 2.15444
R6004 vdd.n3469 vdd.t70 2.15444
R6005 vdd.n320 vdd.n296 1.93989
R6006 vdd.n261 vdd.n237 1.93989
R6007 vdd.n218 vdd.n194 1.93989
R6008 vdd.n159 vdd.n135 1.93989
R6009 vdd.n117 vdd.n93 1.93989
R6010 vdd.n58 vdd.n34 1.93989
R6011 vdd.n2101 vdd.n2077 1.93989
R6012 vdd.n2160 vdd.n2136 1.93989
R6013 vdd.n1999 vdd.n1975 1.93989
R6014 vdd.n2058 vdd.n2034 1.93989
R6015 vdd.n1898 vdd.n1874 1.93989
R6016 vdd.n1957 vdd.n1933 1.93989
R6017 vdd.n1806 vdd.t72 1.92771
R6018 vdd.t87 vdd.n375 1.92771
R6019 vdd.n2491 vdd.t25 1.81434
R6020 vdd.n2847 vdd.t0 1.81434
R6021 vdd.n1814 vdd.t158 1.70098
R6022 vdd.n3463 vdd.t122 1.70098
R6023 vdd.n2485 vdd.t41 1.58761
R6024 vdd.n901 vdd.t49 1.58761
R6025 vdd.n1839 vdd.t68 1.47425
R6026 vdd.n361 vdd.t150 1.47425
R6027 vdd.n1505 vdd.t64 1.24752
R6028 vdd.n2461 vdd.t32 1.24752
R6029 vdd.n1024 vdd.t7 1.24752
R6030 vdd.n2981 vdd.t51 1.24752
R6031 vdd.n878 vdd.t19 1.24752
R6032 vdd.t97 vdd.n3485 1.24752
R6033 vdd.n331 vdd.n291 1.16414
R6034 vdd.n324 vdd.n323 1.16414
R6035 vdd.n272 vdd.n232 1.16414
R6036 vdd.n265 vdd.n264 1.16414
R6037 vdd.n229 vdd.n189 1.16414
R6038 vdd.n222 vdd.n221 1.16414
R6039 vdd.n170 vdd.n130 1.16414
R6040 vdd.n163 vdd.n162 1.16414
R6041 vdd.n128 vdd.n88 1.16414
R6042 vdd.n121 vdd.n120 1.16414
R6043 vdd.n69 vdd.n29 1.16414
R6044 vdd.n62 vdd.n61 1.16414
R6045 vdd.n2112 vdd.n2072 1.16414
R6046 vdd.n2105 vdd.n2104 1.16414
R6047 vdd.n2171 vdd.n2131 1.16414
R6048 vdd.n2164 vdd.n2163 1.16414
R6049 vdd.n2010 vdd.n1970 1.16414
R6050 vdd.n2003 vdd.n2002 1.16414
R6051 vdd.n2069 vdd.n2029 1.16414
R6052 vdd.n2062 vdd.n2061 1.16414
R6053 vdd.n1909 vdd.n1869 1.16414
R6054 vdd.n1902 vdd.n1901 1.16414
R6055 vdd.n1968 vdd.n1928 1.16414
R6056 vdd.n1961 vdd.n1960 1.16414
R6057 vdd.n2188 vdd.t109 1.02079
R6058 vdd.t282 vdd.t32 1.02079
R6059 vdd.t19 vdd.t251 1.02079
R6060 vdd.t153 vdd.n633 1.02079
R6061 vdd.n2174 vdd.n28 1.00834
R6062 vdd vdd.n3492 1.0005
R6063 vdd.n1685 vdd.n1681 0.970197
R6064 vdd.n2272 vdd.n2271 0.970197
R6065 vdd.n618 vdd.n428 0.970197
R6066 vdd.n3187 vdd.n690 0.970197
R6067 vdd.n2204 vdd.t83 0.794056
R6068 vdd.n3373 vdd.t78 0.794056
R6069 vdd.n2229 vdd.t142 0.567326
R6070 vdd.t66 vdd.n662 0.567326
R6071 vdd.n2262 vdd.n1123 0.530988
R6072 vdd.n726 vdd.n682 0.530988
R6073 vdd.n464 vdd.n391 0.530988
R6074 vdd.n3442 vdd.n3441 0.530988
R6075 vdd.n3319 vdd.n3318 0.530988
R6076 vdd.n2251 vdd.n1424 0.530988
R6077 vdd.n1683 vdd.n1548 0.530988
R6078 vdd.n1785 vdd.n1784 0.530988
R6079 vdd.n4 vdd.n2 0.459552
R6080 vdd.n11 vdd.n9 0.459552
R6081 vdd.t15 vdd.n976 0.453961
R6082 vdd.n2945 vdd.t35 0.453961
R6083 vdd.n329 vdd.n328 0.388379
R6084 vdd.n295 vdd.n293 0.388379
R6085 vdd.n270 vdd.n269 0.388379
R6086 vdd.n236 vdd.n234 0.388379
R6087 vdd.n227 vdd.n226 0.388379
R6088 vdd.n193 vdd.n191 0.388379
R6089 vdd.n168 vdd.n167 0.388379
R6090 vdd.n134 vdd.n132 0.388379
R6091 vdd.n126 vdd.n125 0.388379
R6092 vdd.n92 vdd.n90 0.388379
R6093 vdd.n67 vdd.n66 0.388379
R6094 vdd.n33 vdd.n31 0.388379
R6095 vdd.n2110 vdd.n2109 0.388379
R6096 vdd.n2076 vdd.n2074 0.388379
R6097 vdd.n2169 vdd.n2168 0.388379
R6098 vdd.n2135 vdd.n2133 0.388379
R6099 vdd.n2008 vdd.n2007 0.388379
R6100 vdd.n1974 vdd.n1972 0.388379
R6101 vdd.n2067 vdd.n2066 0.388379
R6102 vdd.n2033 vdd.n2031 0.388379
R6103 vdd.n1907 vdd.n1906 0.388379
R6104 vdd.n1873 vdd.n1871 0.388379
R6105 vdd.n1966 vdd.n1965 0.388379
R6106 vdd.n1932 vdd.n1930 0.388379
R6107 vdd.n19 vdd.n17 0.387128
R6108 vdd.n24 vdd.n22 0.387128
R6109 vdd.n6 vdd.n4 0.358259
R6110 vdd.n13 vdd.n11 0.358259
R6111 vdd.n276 vdd.n274 0.358259
R6112 vdd.n278 vdd.n276 0.358259
R6113 vdd.n280 vdd.n278 0.358259
R6114 vdd.n282 vdd.n280 0.358259
R6115 vdd.n284 vdd.n282 0.358259
R6116 vdd.n286 vdd.n284 0.358259
R6117 vdd.n288 vdd.n286 0.358259
R6118 vdd.n290 vdd.n288 0.358259
R6119 vdd.n332 vdd.n290 0.358259
R6120 vdd.n174 vdd.n172 0.358259
R6121 vdd.n176 vdd.n174 0.358259
R6122 vdd.n178 vdd.n176 0.358259
R6123 vdd.n180 vdd.n178 0.358259
R6124 vdd.n182 vdd.n180 0.358259
R6125 vdd.n184 vdd.n182 0.358259
R6126 vdd.n186 vdd.n184 0.358259
R6127 vdd.n188 vdd.n186 0.358259
R6128 vdd.n230 vdd.n188 0.358259
R6129 vdd.n73 vdd.n71 0.358259
R6130 vdd.n75 vdd.n73 0.358259
R6131 vdd.n77 vdd.n75 0.358259
R6132 vdd.n79 vdd.n77 0.358259
R6133 vdd.n81 vdd.n79 0.358259
R6134 vdd.n83 vdd.n81 0.358259
R6135 vdd.n85 vdd.n83 0.358259
R6136 vdd.n87 vdd.n85 0.358259
R6137 vdd.n129 vdd.n87 0.358259
R6138 vdd.n2172 vdd.n2130 0.358259
R6139 vdd.n2130 vdd.n2128 0.358259
R6140 vdd.n2128 vdd.n2126 0.358259
R6141 vdd.n2126 vdd.n2124 0.358259
R6142 vdd.n2124 vdd.n2122 0.358259
R6143 vdd.n2122 vdd.n2120 0.358259
R6144 vdd.n2120 vdd.n2118 0.358259
R6145 vdd.n2118 vdd.n2116 0.358259
R6146 vdd.n2116 vdd.n2114 0.358259
R6147 vdd.n2070 vdd.n2028 0.358259
R6148 vdd.n2028 vdd.n2026 0.358259
R6149 vdd.n2026 vdd.n2024 0.358259
R6150 vdd.n2024 vdd.n2022 0.358259
R6151 vdd.n2022 vdd.n2020 0.358259
R6152 vdd.n2020 vdd.n2018 0.358259
R6153 vdd.n2018 vdd.n2016 0.358259
R6154 vdd.n2016 vdd.n2014 0.358259
R6155 vdd.n2014 vdd.n2012 0.358259
R6156 vdd.n1969 vdd.n1927 0.358259
R6157 vdd.n1927 vdd.n1925 0.358259
R6158 vdd.n1925 vdd.n1923 0.358259
R6159 vdd.n1923 vdd.n1921 0.358259
R6160 vdd.n1921 vdd.n1919 0.358259
R6161 vdd.n1919 vdd.n1917 0.358259
R6162 vdd.n1917 vdd.n1915 0.358259
R6163 vdd.n1915 vdd.n1913 0.358259
R6164 vdd.n1913 vdd.n1911 0.358259
R6165 vdd.t45 vdd.n1052 0.340595
R6166 vdd.n2497 vdd.t9 0.340595
R6167 vdd.t20 vdd.n905 0.340595
R6168 vdd.n3018 vdd.t8 0.340595
R6169 vdd.n14 vdd.n6 0.334552
R6170 vdd.n14 vdd.n13 0.334552
R6171 vdd.n27 vdd.n19 0.21707
R6172 vdd.n27 vdd.n24 0.21707
R6173 vdd.n330 vdd.n292 0.155672
R6174 vdd.n322 vdd.n292 0.155672
R6175 vdd.n322 vdd.n321 0.155672
R6176 vdd.n321 vdd.n297 0.155672
R6177 vdd.n314 vdd.n297 0.155672
R6178 vdd.n314 vdd.n313 0.155672
R6179 vdd.n313 vdd.n301 0.155672
R6180 vdd.n306 vdd.n301 0.155672
R6181 vdd.n271 vdd.n233 0.155672
R6182 vdd.n263 vdd.n233 0.155672
R6183 vdd.n263 vdd.n262 0.155672
R6184 vdd.n262 vdd.n238 0.155672
R6185 vdd.n255 vdd.n238 0.155672
R6186 vdd.n255 vdd.n254 0.155672
R6187 vdd.n254 vdd.n242 0.155672
R6188 vdd.n247 vdd.n242 0.155672
R6189 vdd.n228 vdd.n190 0.155672
R6190 vdd.n220 vdd.n190 0.155672
R6191 vdd.n220 vdd.n219 0.155672
R6192 vdd.n219 vdd.n195 0.155672
R6193 vdd.n212 vdd.n195 0.155672
R6194 vdd.n212 vdd.n211 0.155672
R6195 vdd.n211 vdd.n199 0.155672
R6196 vdd.n204 vdd.n199 0.155672
R6197 vdd.n169 vdd.n131 0.155672
R6198 vdd.n161 vdd.n131 0.155672
R6199 vdd.n161 vdd.n160 0.155672
R6200 vdd.n160 vdd.n136 0.155672
R6201 vdd.n153 vdd.n136 0.155672
R6202 vdd.n153 vdd.n152 0.155672
R6203 vdd.n152 vdd.n140 0.155672
R6204 vdd.n145 vdd.n140 0.155672
R6205 vdd.n127 vdd.n89 0.155672
R6206 vdd.n119 vdd.n89 0.155672
R6207 vdd.n119 vdd.n118 0.155672
R6208 vdd.n118 vdd.n94 0.155672
R6209 vdd.n111 vdd.n94 0.155672
R6210 vdd.n111 vdd.n110 0.155672
R6211 vdd.n110 vdd.n98 0.155672
R6212 vdd.n103 vdd.n98 0.155672
R6213 vdd.n68 vdd.n30 0.155672
R6214 vdd.n60 vdd.n30 0.155672
R6215 vdd.n60 vdd.n59 0.155672
R6216 vdd.n59 vdd.n35 0.155672
R6217 vdd.n52 vdd.n35 0.155672
R6218 vdd.n52 vdd.n51 0.155672
R6219 vdd.n51 vdd.n39 0.155672
R6220 vdd.n44 vdd.n39 0.155672
R6221 vdd.n2111 vdd.n2073 0.155672
R6222 vdd.n2103 vdd.n2073 0.155672
R6223 vdd.n2103 vdd.n2102 0.155672
R6224 vdd.n2102 vdd.n2078 0.155672
R6225 vdd.n2095 vdd.n2078 0.155672
R6226 vdd.n2095 vdd.n2094 0.155672
R6227 vdd.n2094 vdd.n2082 0.155672
R6228 vdd.n2087 vdd.n2082 0.155672
R6229 vdd.n2170 vdd.n2132 0.155672
R6230 vdd.n2162 vdd.n2132 0.155672
R6231 vdd.n2162 vdd.n2161 0.155672
R6232 vdd.n2161 vdd.n2137 0.155672
R6233 vdd.n2154 vdd.n2137 0.155672
R6234 vdd.n2154 vdd.n2153 0.155672
R6235 vdd.n2153 vdd.n2141 0.155672
R6236 vdd.n2146 vdd.n2141 0.155672
R6237 vdd.n2009 vdd.n1971 0.155672
R6238 vdd.n2001 vdd.n1971 0.155672
R6239 vdd.n2001 vdd.n2000 0.155672
R6240 vdd.n2000 vdd.n1976 0.155672
R6241 vdd.n1993 vdd.n1976 0.155672
R6242 vdd.n1993 vdd.n1992 0.155672
R6243 vdd.n1992 vdd.n1980 0.155672
R6244 vdd.n1985 vdd.n1980 0.155672
R6245 vdd.n2068 vdd.n2030 0.155672
R6246 vdd.n2060 vdd.n2030 0.155672
R6247 vdd.n2060 vdd.n2059 0.155672
R6248 vdd.n2059 vdd.n2035 0.155672
R6249 vdd.n2052 vdd.n2035 0.155672
R6250 vdd.n2052 vdd.n2051 0.155672
R6251 vdd.n2051 vdd.n2039 0.155672
R6252 vdd.n2044 vdd.n2039 0.155672
R6253 vdd.n1908 vdd.n1870 0.155672
R6254 vdd.n1900 vdd.n1870 0.155672
R6255 vdd.n1900 vdd.n1899 0.155672
R6256 vdd.n1899 vdd.n1875 0.155672
R6257 vdd.n1892 vdd.n1875 0.155672
R6258 vdd.n1892 vdd.n1891 0.155672
R6259 vdd.n1891 vdd.n1879 0.155672
R6260 vdd.n1884 vdd.n1879 0.155672
R6261 vdd.n1967 vdd.n1929 0.155672
R6262 vdd.n1959 vdd.n1929 0.155672
R6263 vdd.n1959 vdd.n1958 0.155672
R6264 vdd.n1958 vdd.n1934 0.155672
R6265 vdd.n1951 vdd.n1934 0.155672
R6266 vdd.n1951 vdd.n1950 0.155672
R6267 vdd.n1950 vdd.n1938 0.155672
R6268 vdd.n1943 vdd.n1938 0.155672
R6269 vdd.n1128 vdd.n1120 0.152939
R6270 vdd.n1132 vdd.n1128 0.152939
R6271 vdd.n1133 vdd.n1132 0.152939
R6272 vdd.n1134 vdd.n1133 0.152939
R6273 vdd.n1135 vdd.n1134 0.152939
R6274 vdd.n1139 vdd.n1135 0.152939
R6275 vdd.n1140 vdd.n1139 0.152939
R6276 vdd.n1141 vdd.n1140 0.152939
R6277 vdd.n1142 vdd.n1141 0.152939
R6278 vdd.n1146 vdd.n1142 0.152939
R6279 vdd.n1147 vdd.n1146 0.152939
R6280 vdd.n1148 vdd.n1147 0.152939
R6281 vdd.n2345 vdd.n1148 0.152939
R6282 vdd.n2345 vdd.n2344 0.152939
R6283 vdd.n2344 vdd.n2343 0.152939
R6284 vdd.n2343 vdd.n1154 0.152939
R6285 vdd.n1159 vdd.n1154 0.152939
R6286 vdd.n1160 vdd.n1159 0.152939
R6287 vdd.n1161 vdd.n1160 0.152939
R6288 vdd.n1165 vdd.n1161 0.152939
R6289 vdd.n1166 vdd.n1165 0.152939
R6290 vdd.n1167 vdd.n1166 0.152939
R6291 vdd.n1168 vdd.n1167 0.152939
R6292 vdd.n1172 vdd.n1168 0.152939
R6293 vdd.n1173 vdd.n1172 0.152939
R6294 vdd.n1174 vdd.n1173 0.152939
R6295 vdd.n1175 vdd.n1174 0.152939
R6296 vdd.n1179 vdd.n1175 0.152939
R6297 vdd.n1180 vdd.n1179 0.152939
R6298 vdd.n1181 vdd.n1180 0.152939
R6299 vdd.n1182 vdd.n1181 0.152939
R6300 vdd.n1186 vdd.n1182 0.152939
R6301 vdd.n1187 vdd.n1186 0.152939
R6302 vdd.n1188 vdd.n1187 0.152939
R6303 vdd.n2306 vdd.n1188 0.152939
R6304 vdd.n2306 vdd.n2305 0.152939
R6305 vdd.n2305 vdd.n2304 0.152939
R6306 vdd.n2304 vdd.n1194 0.152939
R6307 vdd.n1199 vdd.n1194 0.152939
R6308 vdd.n1200 vdd.n1199 0.152939
R6309 vdd.n1201 vdd.n1200 0.152939
R6310 vdd.n1205 vdd.n1201 0.152939
R6311 vdd.n1206 vdd.n1205 0.152939
R6312 vdd.n1207 vdd.n1206 0.152939
R6313 vdd.n1208 vdd.n1207 0.152939
R6314 vdd.n1212 vdd.n1208 0.152939
R6315 vdd.n1213 vdd.n1212 0.152939
R6316 vdd.n1214 vdd.n1213 0.152939
R6317 vdd.n1215 vdd.n1214 0.152939
R6318 vdd.n1219 vdd.n1215 0.152939
R6319 vdd.n1220 vdd.n1219 0.152939
R6320 vdd.n2380 vdd.n1123 0.152939
R6321 vdd.n2176 vdd.n1485 0.152939
R6322 vdd.n2191 vdd.n1485 0.152939
R6323 vdd.n2192 vdd.n2191 0.152939
R6324 vdd.n2193 vdd.n2192 0.152939
R6325 vdd.n2193 vdd.n1474 0.152939
R6326 vdd.n2208 vdd.n1474 0.152939
R6327 vdd.n2209 vdd.n2208 0.152939
R6328 vdd.n2210 vdd.n2209 0.152939
R6329 vdd.n2210 vdd.n1463 0.152939
R6330 vdd.n2224 vdd.n1463 0.152939
R6331 vdd.n2225 vdd.n2224 0.152939
R6332 vdd.n2226 vdd.n2225 0.152939
R6333 vdd.n2226 vdd.n1451 0.152939
R6334 vdd.n2241 vdd.n1451 0.152939
R6335 vdd.n2242 vdd.n2241 0.152939
R6336 vdd.n2243 vdd.n2242 0.152939
R6337 vdd.n2243 vdd.n1439 0.152939
R6338 vdd.n2260 vdd.n1439 0.152939
R6339 vdd.n2261 vdd.n2260 0.152939
R6340 vdd.n2262 vdd.n2261 0.152939
R6341 vdd.n735 vdd.n730 0.152939
R6342 vdd.n736 vdd.n735 0.152939
R6343 vdd.n737 vdd.n736 0.152939
R6344 vdd.n738 vdd.n737 0.152939
R6345 vdd.n739 vdd.n738 0.152939
R6346 vdd.n740 vdd.n739 0.152939
R6347 vdd.n741 vdd.n740 0.152939
R6348 vdd.n742 vdd.n741 0.152939
R6349 vdd.n743 vdd.n742 0.152939
R6350 vdd.n744 vdd.n743 0.152939
R6351 vdd.n745 vdd.n744 0.152939
R6352 vdd.n746 vdd.n745 0.152939
R6353 vdd.n3275 vdd.n746 0.152939
R6354 vdd.n3275 vdd.n3274 0.152939
R6355 vdd.n3274 vdd.n3273 0.152939
R6356 vdd.n3273 vdd.n748 0.152939
R6357 vdd.n749 vdd.n748 0.152939
R6358 vdd.n750 vdd.n749 0.152939
R6359 vdd.n751 vdd.n750 0.152939
R6360 vdd.n752 vdd.n751 0.152939
R6361 vdd.n753 vdd.n752 0.152939
R6362 vdd.n754 vdd.n753 0.152939
R6363 vdd.n755 vdd.n754 0.152939
R6364 vdd.n756 vdd.n755 0.152939
R6365 vdd.n757 vdd.n756 0.152939
R6366 vdd.n758 vdd.n757 0.152939
R6367 vdd.n759 vdd.n758 0.152939
R6368 vdd.n760 vdd.n759 0.152939
R6369 vdd.n761 vdd.n760 0.152939
R6370 vdd.n762 vdd.n761 0.152939
R6371 vdd.n763 vdd.n762 0.152939
R6372 vdd.n764 vdd.n763 0.152939
R6373 vdd.n765 vdd.n764 0.152939
R6374 vdd.n766 vdd.n765 0.152939
R6375 vdd.n3229 vdd.n766 0.152939
R6376 vdd.n3229 vdd.n3228 0.152939
R6377 vdd.n3228 vdd.n3227 0.152939
R6378 vdd.n3227 vdd.n770 0.152939
R6379 vdd.n771 vdd.n770 0.152939
R6380 vdd.n772 vdd.n771 0.152939
R6381 vdd.n773 vdd.n772 0.152939
R6382 vdd.n774 vdd.n773 0.152939
R6383 vdd.n775 vdd.n774 0.152939
R6384 vdd.n776 vdd.n775 0.152939
R6385 vdd.n777 vdd.n776 0.152939
R6386 vdd.n778 vdd.n777 0.152939
R6387 vdd.n779 vdd.n778 0.152939
R6388 vdd.n780 vdd.n779 0.152939
R6389 vdd.n781 vdd.n780 0.152939
R6390 vdd.n782 vdd.n781 0.152939
R6391 vdd.n783 vdd.n782 0.152939
R6392 vdd.n727 vdd.n726 0.152939
R6393 vdd.n3326 vdd.n682 0.152939
R6394 vdd.n3327 vdd.n3326 0.152939
R6395 vdd.n3328 vdd.n3327 0.152939
R6396 vdd.n3328 vdd.n670 0.152939
R6397 vdd.n3343 vdd.n670 0.152939
R6398 vdd.n3344 vdd.n3343 0.152939
R6399 vdd.n3345 vdd.n3344 0.152939
R6400 vdd.n3345 vdd.n659 0.152939
R6401 vdd.n3359 vdd.n659 0.152939
R6402 vdd.n3360 vdd.n3359 0.152939
R6403 vdd.n3361 vdd.n3360 0.152939
R6404 vdd.n3361 vdd.n647 0.152939
R6405 vdd.n3376 vdd.n647 0.152939
R6406 vdd.n3377 vdd.n3376 0.152939
R6407 vdd.n3378 vdd.n3377 0.152939
R6408 vdd.n3378 vdd.n636 0.152939
R6409 vdd.n3395 vdd.n636 0.152939
R6410 vdd.n3396 vdd.n3395 0.152939
R6411 vdd.n3397 vdd.n3396 0.152939
R6412 vdd.n3397 vdd.n334 0.152939
R6413 vdd.n3490 vdd.n335 0.152939
R6414 vdd.n346 vdd.n335 0.152939
R6415 vdd.n347 vdd.n346 0.152939
R6416 vdd.n348 vdd.n347 0.152939
R6417 vdd.n355 vdd.n348 0.152939
R6418 vdd.n356 vdd.n355 0.152939
R6419 vdd.n357 vdd.n356 0.152939
R6420 vdd.n358 vdd.n357 0.152939
R6421 vdd.n366 vdd.n358 0.152939
R6422 vdd.n367 vdd.n366 0.152939
R6423 vdd.n368 vdd.n367 0.152939
R6424 vdd.n369 vdd.n368 0.152939
R6425 vdd.n377 vdd.n369 0.152939
R6426 vdd.n378 vdd.n377 0.152939
R6427 vdd.n379 vdd.n378 0.152939
R6428 vdd.n380 vdd.n379 0.152939
R6429 vdd.n388 vdd.n380 0.152939
R6430 vdd.n389 vdd.n388 0.152939
R6431 vdd.n390 vdd.n389 0.152939
R6432 vdd.n391 vdd.n390 0.152939
R6433 vdd.n464 vdd.n463 0.152939
R6434 vdd.n470 vdd.n463 0.152939
R6435 vdd.n471 vdd.n470 0.152939
R6436 vdd.n472 vdd.n471 0.152939
R6437 vdd.n472 vdd.n461 0.152939
R6438 vdd.n480 vdd.n461 0.152939
R6439 vdd.n481 vdd.n480 0.152939
R6440 vdd.n482 vdd.n481 0.152939
R6441 vdd.n482 vdd.n459 0.152939
R6442 vdd.n490 vdd.n459 0.152939
R6443 vdd.n491 vdd.n490 0.152939
R6444 vdd.n492 vdd.n491 0.152939
R6445 vdd.n492 vdd.n457 0.152939
R6446 vdd.n500 vdd.n457 0.152939
R6447 vdd.n501 vdd.n500 0.152939
R6448 vdd.n502 vdd.n501 0.152939
R6449 vdd.n502 vdd.n455 0.152939
R6450 vdd.n510 vdd.n455 0.152939
R6451 vdd.n511 vdd.n510 0.152939
R6452 vdd.n512 vdd.n511 0.152939
R6453 vdd.n512 vdd.n451 0.152939
R6454 vdd.n520 vdd.n451 0.152939
R6455 vdd.n521 vdd.n520 0.152939
R6456 vdd.n522 vdd.n521 0.152939
R6457 vdd.n522 vdd.n449 0.152939
R6458 vdd.n530 vdd.n449 0.152939
R6459 vdd.n531 vdd.n530 0.152939
R6460 vdd.n532 vdd.n531 0.152939
R6461 vdd.n532 vdd.n447 0.152939
R6462 vdd.n540 vdd.n447 0.152939
R6463 vdd.n541 vdd.n540 0.152939
R6464 vdd.n542 vdd.n541 0.152939
R6465 vdd.n542 vdd.n445 0.152939
R6466 vdd.n550 vdd.n445 0.152939
R6467 vdd.n551 vdd.n550 0.152939
R6468 vdd.n552 vdd.n551 0.152939
R6469 vdd.n552 vdd.n443 0.152939
R6470 vdd.n560 vdd.n443 0.152939
R6471 vdd.n561 vdd.n560 0.152939
R6472 vdd.n562 vdd.n561 0.152939
R6473 vdd.n562 vdd.n439 0.152939
R6474 vdd.n570 vdd.n439 0.152939
R6475 vdd.n571 vdd.n570 0.152939
R6476 vdd.n572 vdd.n571 0.152939
R6477 vdd.n572 vdd.n437 0.152939
R6478 vdd.n580 vdd.n437 0.152939
R6479 vdd.n581 vdd.n580 0.152939
R6480 vdd.n582 vdd.n581 0.152939
R6481 vdd.n582 vdd.n435 0.152939
R6482 vdd.n590 vdd.n435 0.152939
R6483 vdd.n591 vdd.n590 0.152939
R6484 vdd.n592 vdd.n591 0.152939
R6485 vdd.n592 vdd.n433 0.152939
R6486 vdd.n600 vdd.n433 0.152939
R6487 vdd.n601 vdd.n600 0.152939
R6488 vdd.n602 vdd.n601 0.152939
R6489 vdd.n602 vdd.n431 0.152939
R6490 vdd.n610 vdd.n431 0.152939
R6491 vdd.n611 vdd.n610 0.152939
R6492 vdd.n612 vdd.n611 0.152939
R6493 vdd.n612 vdd.n429 0.152939
R6494 vdd.n619 vdd.n429 0.152939
R6495 vdd.n3442 vdd.n619 0.152939
R6496 vdd.n3320 vdd.n3319 0.152939
R6497 vdd.n3320 vdd.n675 0.152939
R6498 vdd.n3334 vdd.n675 0.152939
R6499 vdd.n3335 vdd.n3334 0.152939
R6500 vdd.n3336 vdd.n3335 0.152939
R6501 vdd.n3336 vdd.n665 0.152939
R6502 vdd.n3351 vdd.n665 0.152939
R6503 vdd.n3352 vdd.n3351 0.152939
R6504 vdd.n3353 vdd.n3352 0.152939
R6505 vdd.n3353 vdd.n652 0.152939
R6506 vdd.n3367 vdd.n652 0.152939
R6507 vdd.n3368 vdd.n3367 0.152939
R6508 vdd.n3369 vdd.n3368 0.152939
R6509 vdd.n3369 vdd.n641 0.152939
R6510 vdd.n3384 vdd.n641 0.152939
R6511 vdd.n3385 vdd.n3384 0.152939
R6512 vdd.n3386 vdd.n3385 0.152939
R6513 vdd.n3388 vdd.n3386 0.152939
R6514 vdd.n3388 vdd.n3387 0.152939
R6515 vdd.n3387 vdd.n630 0.152939
R6516 vdd.n3405 vdd.n630 0.152939
R6517 vdd.n3406 vdd.n3405 0.152939
R6518 vdd.n3407 vdd.n3406 0.152939
R6519 vdd.n3407 vdd.n628 0.152939
R6520 vdd.n3412 vdd.n628 0.152939
R6521 vdd.n3413 vdd.n3412 0.152939
R6522 vdd.n3414 vdd.n3413 0.152939
R6523 vdd.n3414 vdd.n626 0.152939
R6524 vdd.n3419 vdd.n626 0.152939
R6525 vdd.n3420 vdd.n3419 0.152939
R6526 vdd.n3421 vdd.n3420 0.152939
R6527 vdd.n3421 vdd.n624 0.152939
R6528 vdd.n3427 vdd.n624 0.152939
R6529 vdd.n3428 vdd.n3427 0.152939
R6530 vdd.n3429 vdd.n3428 0.152939
R6531 vdd.n3429 vdd.n622 0.152939
R6532 vdd.n3434 vdd.n622 0.152939
R6533 vdd.n3435 vdd.n3434 0.152939
R6534 vdd.n3436 vdd.n3435 0.152939
R6535 vdd.n3436 vdd.n620 0.152939
R6536 vdd.n3441 vdd.n620 0.152939
R6537 vdd.n3318 vdd.n687 0.152939
R6538 vdd.n2273 vdd.n1424 0.152939
R6539 vdd.n1792 vdd.n1548 0.152939
R6540 vdd.n1793 vdd.n1792 0.152939
R6541 vdd.n1794 vdd.n1793 0.152939
R6542 vdd.n1794 vdd.n1536 0.152939
R6543 vdd.n1809 vdd.n1536 0.152939
R6544 vdd.n1810 vdd.n1809 0.152939
R6545 vdd.n1811 vdd.n1810 0.152939
R6546 vdd.n1811 vdd.n1526 0.152939
R6547 vdd.n1826 vdd.n1526 0.152939
R6548 vdd.n1827 vdd.n1826 0.152939
R6549 vdd.n1828 vdd.n1827 0.152939
R6550 vdd.n1828 vdd.n1513 0.152939
R6551 vdd.n1842 vdd.n1513 0.152939
R6552 vdd.n1843 vdd.n1842 0.152939
R6553 vdd.n1844 vdd.n1843 0.152939
R6554 vdd.n1844 vdd.n1502 0.152939
R6555 vdd.n1859 vdd.n1502 0.152939
R6556 vdd.n1860 vdd.n1859 0.152939
R6557 vdd.n1861 vdd.n1860 0.152939
R6558 vdd.n1861 vdd.n1491 0.152939
R6559 vdd.n2182 vdd.n1491 0.152939
R6560 vdd.n2183 vdd.n2182 0.152939
R6561 vdd.n2184 vdd.n2183 0.152939
R6562 vdd.n2184 vdd.n1479 0.152939
R6563 vdd.n2199 vdd.n1479 0.152939
R6564 vdd.n2200 vdd.n2199 0.152939
R6565 vdd.n2201 vdd.n2200 0.152939
R6566 vdd.n2201 vdd.n1469 0.152939
R6567 vdd.n2216 vdd.n1469 0.152939
R6568 vdd.n2217 vdd.n2216 0.152939
R6569 vdd.n2218 vdd.n2217 0.152939
R6570 vdd.n2218 vdd.n1456 0.152939
R6571 vdd.n2232 vdd.n1456 0.152939
R6572 vdd.n2233 vdd.n2232 0.152939
R6573 vdd.n2234 vdd.n2233 0.152939
R6574 vdd.n2234 vdd.n1446 0.152939
R6575 vdd.n2249 vdd.n1446 0.152939
R6576 vdd.n2250 vdd.n2249 0.152939
R6577 vdd.n2253 vdd.n2250 0.152939
R6578 vdd.n2253 vdd.n2252 0.152939
R6579 vdd.n2252 vdd.n2251 0.152939
R6580 vdd.n1784 vdd.n1553 0.152939
R6581 vdd.n1777 vdd.n1553 0.152939
R6582 vdd.n1777 vdd.n1776 0.152939
R6583 vdd.n1776 vdd.n1775 0.152939
R6584 vdd.n1775 vdd.n1590 0.152939
R6585 vdd.n1771 vdd.n1590 0.152939
R6586 vdd.n1771 vdd.n1770 0.152939
R6587 vdd.n1770 vdd.n1769 0.152939
R6588 vdd.n1769 vdd.n1596 0.152939
R6589 vdd.n1765 vdd.n1596 0.152939
R6590 vdd.n1765 vdd.n1764 0.152939
R6591 vdd.n1764 vdd.n1763 0.152939
R6592 vdd.n1763 vdd.n1602 0.152939
R6593 vdd.n1759 vdd.n1602 0.152939
R6594 vdd.n1759 vdd.n1758 0.152939
R6595 vdd.n1758 vdd.n1757 0.152939
R6596 vdd.n1757 vdd.n1608 0.152939
R6597 vdd.n1753 vdd.n1608 0.152939
R6598 vdd.n1753 vdd.n1752 0.152939
R6599 vdd.n1752 vdd.n1751 0.152939
R6600 vdd.n1751 vdd.n1616 0.152939
R6601 vdd.n1747 vdd.n1616 0.152939
R6602 vdd.n1747 vdd.n1746 0.152939
R6603 vdd.n1746 vdd.n1745 0.152939
R6604 vdd.n1745 vdd.n1622 0.152939
R6605 vdd.n1741 vdd.n1622 0.152939
R6606 vdd.n1741 vdd.n1740 0.152939
R6607 vdd.n1740 vdd.n1739 0.152939
R6608 vdd.n1739 vdd.n1628 0.152939
R6609 vdd.n1735 vdd.n1628 0.152939
R6610 vdd.n1735 vdd.n1734 0.152939
R6611 vdd.n1734 vdd.n1733 0.152939
R6612 vdd.n1733 vdd.n1634 0.152939
R6613 vdd.n1729 vdd.n1634 0.152939
R6614 vdd.n1729 vdd.n1728 0.152939
R6615 vdd.n1728 vdd.n1727 0.152939
R6616 vdd.n1727 vdd.n1640 0.152939
R6617 vdd.n1723 vdd.n1640 0.152939
R6618 vdd.n1723 vdd.n1722 0.152939
R6619 vdd.n1722 vdd.n1721 0.152939
R6620 vdd.n1721 vdd.n1646 0.152939
R6621 vdd.n1714 vdd.n1646 0.152939
R6622 vdd.n1714 vdd.n1713 0.152939
R6623 vdd.n1713 vdd.n1712 0.152939
R6624 vdd.n1712 vdd.n1651 0.152939
R6625 vdd.n1708 vdd.n1651 0.152939
R6626 vdd.n1708 vdd.n1707 0.152939
R6627 vdd.n1707 vdd.n1706 0.152939
R6628 vdd.n1706 vdd.n1657 0.152939
R6629 vdd.n1702 vdd.n1657 0.152939
R6630 vdd.n1702 vdd.n1701 0.152939
R6631 vdd.n1701 vdd.n1700 0.152939
R6632 vdd.n1700 vdd.n1663 0.152939
R6633 vdd.n1696 vdd.n1663 0.152939
R6634 vdd.n1696 vdd.n1695 0.152939
R6635 vdd.n1695 vdd.n1694 0.152939
R6636 vdd.n1694 vdd.n1669 0.152939
R6637 vdd.n1690 vdd.n1669 0.152939
R6638 vdd.n1690 vdd.n1689 0.152939
R6639 vdd.n1689 vdd.n1688 0.152939
R6640 vdd.n1688 vdd.n1675 0.152939
R6641 vdd.n1684 vdd.n1675 0.152939
R6642 vdd.n1684 vdd.n1683 0.152939
R6643 vdd.n1786 vdd.n1785 0.152939
R6644 vdd.n1786 vdd.n1542 0.152939
R6645 vdd.n1801 vdd.n1542 0.152939
R6646 vdd.n1802 vdd.n1801 0.152939
R6647 vdd.n1803 vdd.n1802 0.152939
R6648 vdd.n1803 vdd.n1531 0.152939
R6649 vdd.n1818 vdd.n1531 0.152939
R6650 vdd.n1819 vdd.n1818 0.152939
R6651 vdd.n1820 vdd.n1819 0.152939
R6652 vdd.n1820 vdd.n1520 0.152939
R6653 vdd.n1834 vdd.n1520 0.152939
R6654 vdd.n1835 vdd.n1834 0.152939
R6655 vdd.n1836 vdd.n1835 0.152939
R6656 vdd.n1836 vdd.n1508 0.152939
R6657 vdd.n1851 vdd.n1508 0.152939
R6658 vdd.n1852 vdd.n1851 0.152939
R6659 vdd.n1853 vdd.n1852 0.152939
R6660 vdd.n1853 vdd.n1497 0.152939
R6661 vdd.n1867 vdd.n1497 0.152939
R6662 vdd.n1868 vdd.n1867 0.152939
R6663 vdd.n1789 vdd.t261 0.113865
R6664 vdd.t247 vdd.n386 0.113865
R6665 vdd.n2381 vdd.n2380 0.110256
R6666 vdd.n3308 vdd.n727 0.110256
R6667 vdd.n3185 vdd.n687 0.110256
R6668 vdd.n2274 vdd.n2273 0.110256
R6669 vdd.n2176 vdd.n2175 0.0695946
R6670 vdd.n3491 vdd.n334 0.0695946
R6671 vdd.n3491 vdd.n3490 0.0695946
R6672 vdd.n2175 vdd.n1868 0.0695946
R6673 vdd.n2381 vdd.n1120 0.0431829
R6674 vdd.n2274 vdd.n1220 0.0431829
R6675 vdd.n3308 vdd.n730 0.0431829
R6676 vdd.n3185 vdd.n783 0.0431829
R6677 vdd vdd.n28 0.00833333
R6678 CSoutput.n19 CSoutput.t206 184.661
R6679 CSoutput.n78 CSoutput.n77 165.8
R6680 CSoutput.n76 CSoutput.n0 165.8
R6681 CSoutput.n75 CSoutput.n74 165.8
R6682 CSoutput.n73 CSoutput.n72 165.8
R6683 CSoutput.n71 CSoutput.n2 165.8
R6684 CSoutput.n69 CSoutput.n68 165.8
R6685 CSoutput.n67 CSoutput.n3 165.8
R6686 CSoutput.n66 CSoutput.n65 165.8
R6687 CSoutput.n63 CSoutput.n4 165.8
R6688 CSoutput.n61 CSoutput.n60 165.8
R6689 CSoutput.n59 CSoutput.n5 165.8
R6690 CSoutput.n58 CSoutput.n57 165.8
R6691 CSoutput.n55 CSoutput.n6 165.8
R6692 CSoutput.n54 CSoutput.n53 165.8
R6693 CSoutput.n52 CSoutput.n51 165.8
R6694 CSoutput.n50 CSoutput.n8 165.8
R6695 CSoutput.n48 CSoutput.n47 165.8
R6696 CSoutput.n46 CSoutput.n9 165.8
R6697 CSoutput.n45 CSoutput.n44 165.8
R6698 CSoutput.n42 CSoutput.n10 165.8
R6699 CSoutput.n41 CSoutput.n40 165.8
R6700 CSoutput.n39 CSoutput.n38 165.8
R6701 CSoutput.n37 CSoutput.n12 165.8
R6702 CSoutput.n35 CSoutput.n34 165.8
R6703 CSoutput.n33 CSoutput.n13 165.8
R6704 CSoutput.n32 CSoutput.n31 165.8
R6705 CSoutput.n29 CSoutput.n14 165.8
R6706 CSoutput.n28 CSoutput.n27 165.8
R6707 CSoutput.n26 CSoutput.n25 165.8
R6708 CSoutput.n24 CSoutput.n16 165.8
R6709 CSoutput.n22 CSoutput.n21 165.8
R6710 CSoutput.n20 CSoutput.n17 165.8
R6711 CSoutput.n77 CSoutput.t208 162.194
R6712 CSoutput.n18 CSoutput.t209 120.501
R6713 CSoutput.n23 CSoutput.t195 120.501
R6714 CSoutput.n15 CSoutput.t192 120.501
R6715 CSoutput.n30 CSoutput.t210 120.501
R6716 CSoutput.n36 CSoutput.t198 120.501
R6717 CSoutput.n11 CSoutput.t200 120.501
R6718 CSoutput.n43 CSoutput.t212 120.501
R6719 CSoutput.n49 CSoutput.t202 120.501
R6720 CSoutput.n7 CSoutput.t204 120.501
R6721 CSoutput.n56 CSoutput.t196 120.501
R6722 CSoutput.n62 CSoutput.t211 120.501
R6723 CSoutput.n64 CSoutput.t205 120.501
R6724 CSoutput.n70 CSoutput.t199 120.501
R6725 CSoutput.n1 CSoutput.t194 120.501
R6726 CSoutput.n330 CSoutput.n328 103.469
R6727 CSoutput.n310 CSoutput.n308 103.469
R6728 CSoutput.n291 CSoutput.n289 103.469
R6729 CSoutput.n120 CSoutput.n118 103.469
R6730 CSoutput.n100 CSoutput.n98 103.469
R6731 CSoutput.n81 CSoutput.n79 103.469
R6732 CSoutput.n344 CSoutput.n343 103.111
R6733 CSoutput.n342 CSoutput.n341 103.111
R6734 CSoutput.n340 CSoutput.n339 103.111
R6735 CSoutput.n338 CSoutput.n337 103.111
R6736 CSoutput.n336 CSoutput.n335 103.111
R6737 CSoutput.n334 CSoutput.n333 103.111
R6738 CSoutput.n332 CSoutput.n331 103.111
R6739 CSoutput.n330 CSoutput.n329 103.111
R6740 CSoutput.n326 CSoutput.n325 103.111
R6741 CSoutput.n324 CSoutput.n323 103.111
R6742 CSoutput.n322 CSoutput.n321 103.111
R6743 CSoutput.n320 CSoutput.n319 103.111
R6744 CSoutput.n318 CSoutput.n317 103.111
R6745 CSoutput.n316 CSoutput.n315 103.111
R6746 CSoutput.n314 CSoutput.n313 103.111
R6747 CSoutput.n312 CSoutput.n311 103.111
R6748 CSoutput.n310 CSoutput.n309 103.111
R6749 CSoutput.n307 CSoutput.n306 103.111
R6750 CSoutput.n305 CSoutput.n304 103.111
R6751 CSoutput.n303 CSoutput.n302 103.111
R6752 CSoutput.n301 CSoutput.n300 103.111
R6753 CSoutput.n299 CSoutput.n298 103.111
R6754 CSoutput.n297 CSoutput.n296 103.111
R6755 CSoutput.n295 CSoutput.n294 103.111
R6756 CSoutput.n293 CSoutput.n292 103.111
R6757 CSoutput.n291 CSoutput.n290 103.111
R6758 CSoutput.n120 CSoutput.n119 103.111
R6759 CSoutput.n122 CSoutput.n121 103.111
R6760 CSoutput.n124 CSoutput.n123 103.111
R6761 CSoutput.n126 CSoutput.n125 103.111
R6762 CSoutput.n128 CSoutput.n127 103.111
R6763 CSoutput.n130 CSoutput.n129 103.111
R6764 CSoutput.n132 CSoutput.n131 103.111
R6765 CSoutput.n134 CSoutput.n133 103.111
R6766 CSoutput.n136 CSoutput.n135 103.111
R6767 CSoutput.n100 CSoutput.n99 103.111
R6768 CSoutput.n102 CSoutput.n101 103.111
R6769 CSoutput.n104 CSoutput.n103 103.111
R6770 CSoutput.n106 CSoutput.n105 103.111
R6771 CSoutput.n108 CSoutput.n107 103.111
R6772 CSoutput.n110 CSoutput.n109 103.111
R6773 CSoutput.n112 CSoutput.n111 103.111
R6774 CSoutput.n114 CSoutput.n113 103.111
R6775 CSoutput.n116 CSoutput.n115 103.111
R6776 CSoutput.n81 CSoutput.n80 103.111
R6777 CSoutput.n83 CSoutput.n82 103.111
R6778 CSoutput.n85 CSoutput.n84 103.111
R6779 CSoutput.n87 CSoutput.n86 103.111
R6780 CSoutput.n89 CSoutput.n88 103.111
R6781 CSoutput.n91 CSoutput.n90 103.111
R6782 CSoutput.n93 CSoutput.n92 103.111
R6783 CSoutput.n95 CSoutput.n94 103.111
R6784 CSoutput.n97 CSoutput.n96 103.111
R6785 CSoutput.n346 CSoutput.n345 103.111
R6786 CSoutput.n374 CSoutput.n372 81.5057
R6787 CSoutput.n362 CSoutput.n360 81.5057
R6788 CSoutput.n351 CSoutput.n349 81.5057
R6789 CSoutput.n410 CSoutput.n408 81.5057
R6790 CSoutput.n398 CSoutput.n396 81.5057
R6791 CSoutput.n387 CSoutput.n385 81.5057
R6792 CSoutput.n382 CSoutput.n381 80.9324
R6793 CSoutput.n380 CSoutput.n379 80.9324
R6794 CSoutput.n378 CSoutput.n377 80.9324
R6795 CSoutput.n376 CSoutput.n375 80.9324
R6796 CSoutput.n374 CSoutput.n373 80.9324
R6797 CSoutput.n370 CSoutput.n369 80.9324
R6798 CSoutput.n368 CSoutput.n367 80.9324
R6799 CSoutput.n366 CSoutput.n365 80.9324
R6800 CSoutput.n364 CSoutput.n363 80.9324
R6801 CSoutput.n362 CSoutput.n361 80.9324
R6802 CSoutput.n359 CSoutput.n358 80.9324
R6803 CSoutput.n357 CSoutput.n356 80.9324
R6804 CSoutput.n355 CSoutput.n354 80.9324
R6805 CSoutput.n353 CSoutput.n352 80.9324
R6806 CSoutput.n351 CSoutput.n350 80.9324
R6807 CSoutput.n410 CSoutput.n409 80.9324
R6808 CSoutput.n412 CSoutput.n411 80.9324
R6809 CSoutput.n414 CSoutput.n413 80.9324
R6810 CSoutput.n416 CSoutput.n415 80.9324
R6811 CSoutput.n418 CSoutput.n417 80.9324
R6812 CSoutput.n398 CSoutput.n397 80.9324
R6813 CSoutput.n400 CSoutput.n399 80.9324
R6814 CSoutput.n402 CSoutput.n401 80.9324
R6815 CSoutput.n404 CSoutput.n403 80.9324
R6816 CSoutput.n406 CSoutput.n405 80.9324
R6817 CSoutput.n387 CSoutput.n386 80.9324
R6818 CSoutput.n389 CSoutput.n388 80.9324
R6819 CSoutput.n391 CSoutput.n390 80.9324
R6820 CSoutput.n393 CSoutput.n392 80.9324
R6821 CSoutput.n395 CSoutput.n394 80.9324
R6822 CSoutput.n25 CSoutput.n24 48.1486
R6823 CSoutput.n69 CSoutput.n3 48.1486
R6824 CSoutput.n38 CSoutput.n37 48.1486
R6825 CSoutput.n42 CSoutput.n41 48.1486
R6826 CSoutput.n51 CSoutput.n50 48.1486
R6827 CSoutput.n55 CSoutput.n54 48.1486
R6828 CSoutput.n22 CSoutput.n17 46.462
R6829 CSoutput.n72 CSoutput.n71 46.462
R6830 CSoutput.n20 CSoutput.n19 44.9055
R6831 CSoutput.n29 CSoutput.n28 43.7635
R6832 CSoutput.n65 CSoutput.n63 43.7635
R6833 CSoutput.n35 CSoutput.n13 41.7396
R6834 CSoutput.n57 CSoutput.n5 41.7396
R6835 CSoutput.n44 CSoutput.n9 37.0171
R6836 CSoutput.n48 CSoutput.n9 37.0171
R6837 CSoutput.n76 CSoutput.n75 34.9932
R6838 CSoutput.n31 CSoutput.n13 32.2947
R6839 CSoutput.n61 CSoutput.n5 32.2947
R6840 CSoutput.n30 CSoutput.n29 29.6014
R6841 CSoutput.n63 CSoutput.n62 29.6014
R6842 CSoutput.n19 CSoutput.n18 28.4085
R6843 CSoutput.n18 CSoutput.n17 25.1176
R6844 CSoutput.n72 CSoutput.n1 25.1176
R6845 CSoutput.n43 CSoutput.n42 22.0922
R6846 CSoutput.n50 CSoutput.n49 22.0922
R6847 CSoutput.n77 CSoutput.n76 21.8586
R6848 CSoutput.n37 CSoutput.n36 18.9681
R6849 CSoutput.n56 CSoutput.n55 18.9681
R6850 CSoutput.n25 CSoutput.n15 17.6292
R6851 CSoutput.n64 CSoutput.n3 17.6292
R6852 CSoutput.n24 CSoutput.n23 15.844
R6853 CSoutput.n70 CSoutput.n69 15.844
R6854 CSoutput.n38 CSoutput.n11 14.5051
R6855 CSoutput.n54 CSoutput.n7 14.5051
R6856 CSoutput.n421 CSoutput.n78 11.4982
R6857 CSoutput.n41 CSoutput.n11 11.3811
R6858 CSoutput.n51 CSoutput.n7 11.3811
R6859 CSoutput.n23 CSoutput.n22 10.0422
R6860 CSoutput.n71 CSoutput.n70 10.0422
R6861 CSoutput.n327 CSoutput.n307 9.25285
R6862 CSoutput.n117 CSoutput.n97 9.25285
R6863 CSoutput.n371 CSoutput.n359 8.98182
R6864 CSoutput.n407 CSoutput.n395 8.98182
R6865 CSoutput.n384 CSoutput.n348 8.51219
R6866 CSoutput.n28 CSoutput.n15 8.25698
R6867 CSoutput.n65 CSoutput.n64 8.25698
R6868 CSoutput.n348 CSoutput.n347 7.12641
R6869 CSoutput.n138 CSoutput.n137 7.12641
R6870 CSoutput.n36 CSoutput.n35 6.91809
R6871 CSoutput.n57 CSoutput.n56 6.91809
R6872 CSoutput.n384 CSoutput.n383 6.02792
R6873 CSoutput.n420 CSoutput.n419 6.02792
R6874 CSoutput.n383 CSoutput.n382 5.25266
R6875 CSoutput.n371 CSoutput.n370 5.25266
R6876 CSoutput.n419 CSoutput.n418 5.25266
R6877 CSoutput.n407 CSoutput.n406 5.25266
R6878 CSoutput.n347 CSoutput.n346 5.1449
R6879 CSoutput.n327 CSoutput.n326 5.1449
R6880 CSoutput.n137 CSoutput.n136 5.1449
R6881 CSoutput.n117 CSoutput.n116 5.1449
R6882 CSoutput.n421 CSoutput.n138 4.91975
R6883 CSoutput.n229 CSoutput.n182 4.5005
R6884 CSoutput.n198 CSoutput.n182 4.5005
R6885 CSoutput.n193 CSoutput.n177 4.5005
R6886 CSoutput.n193 CSoutput.n179 4.5005
R6887 CSoutput.n193 CSoutput.n176 4.5005
R6888 CSoutput.n193 CSoutput.n180 4.5005
R6889 CSoutput.n193 CSoutput.n175 4.5005
R6890 CSoutput.n193 CSoutput.t197 4.5005
R6891 CSoutput.n193 CSoutput.n174 4.5005
R6892 CSoutput.n193 CSoutput.n181 4.5005
R6893 CSoutput.n193 CSoutput.n182 4.5005
R6894 CSoutput.n191 CSoutput.n177 4.5005
R6895 CSoutput.n191 CSoutput.n179 4.5005
R6896 CSoutput.n191 CSoutput.n176 4.5005
R6897 CSoutput.n191 CSoutput.n180 4.5005
R6898 CSoutput.n191 CSoutput.n175 4.5005
R6899 CSoutput.n191 CSoutput.t197 4.5005
R6900 CSoutput.n191 CSoutput.n174 4.5005
R6901 CSoutput.n191 CSoutput.n181 4.5005
R6902 CSoutput.n191 CSoutput.n182 4.5005
R6903 CSoutput.n190 CSoutput.n177 4.5005
R6904 CSoutput.n190 CSoutput.n179 4.5005
R6905 CSoutput.n190 CSoutput.n176 4.5005
R6906 CSoutput.n190 CSoutput.n180 4.5005
R6907 CSoutput.n190 CSoutput.n175 4.5005
R6908 CSoutput.n190 CSoutput.t197 4.5005
R6909 CSoutput.n190 CSoutput.n174 4.5005
R6910 CSoutput.n190 CSoutput.n181 4.5005
R6911 CSoutput.n190 CSoutput.n182 4.5005
R6912 CSoutput.n275 CSoutput.n177 4.5005
R6913 CSoutput.n275 CSoutput.n179 4.5005
R6914 CSoutput.n275 CSoutput.n176 4.5005
R6915 CSoutput.n275 CSoutput.n180 4.5005
R6916 CSoutput.n275 CSoutput.n175 4.5005
R6917 CSoutput.n275 CSoutput.t197 4.5005
R6918 CSoutput.n275 CSoutput.n174 4.5005
R6919 CSoutput.n275 CSoutput.n181 4.5005
R6920 CSoutput.n275 CSoutput.n182 4.5005
R6921 CSoutput.n273 CSoutput.n177 4.5005
R6922 CSoutput.n273 CSoutput.n179 4.5005
R6923 CSoutput.n273 CSoutput.n176 4.5005
R6924 CSoutput.n273 CSoutput.n180 4.5005
R6925 CSoutput.n273 CSoutput.n175 4.5005
R6926 CSoutput.n273 CSoutput.t197 4.5005
R6927 CSoutput.n273 CSoutput.n174 4.5005
R6928 CSoutput.n273 CSoutput.n181 4.5005
R6929 CSoutput.n271 CSoutput.n177 4.5005
R6930 CSoutput.n271 CSoutput.n179 4.5005
R6931 CSoutput.n271 CSoutput.n176 4.5005
R6932 CSoutput.n271 CSoutput.n180 4.5005
R6933 CSoutput.n271 CSoutput.n175 4.5005
R6934 CSoutput.n271 CSoutput.t197 4.5005
R6935 CSoutput.n271 CSoutput.n174 4.5005
R6936 CSoutput.n271 CSoutput.n181 4.5005
R6937 CSoutput.n201 CSoutput.n177 4.5005
R6938 CSoutput.n201 CSoutput.n179 4.5005
R6939 CSoutput.n201 CSoutput.n176 4.5005
R6940 CSoutput.n201 CSoutput.n180 4.5005
R6941 CSoutput.n201 CSoutput.n175 4.5005
R6942 CSoutput.n201 CSoutput.t197 4.5005
R6943 CSoutput.n201 CSoutput.n174 4.5005
R6944 CSoutput.n201 CSoutput.n181 4.5005
R6945 CSoutput.n201 CSoutput.n182 4.5005
R6946 CSoutput.n200 CSoutput.n177 4.5005
R6947 CSoutput.n200 CSoutput.n179 4.5005
R6948 CSoutput.n200 CSoutput.n176 4.5005
R6949 CSoutput.n200 CSoutput.n180 4.5005
R6950 CSoutput.n200 CSoutput.n175 4.5005
R6951 CSoutput.n200 CSoutput.t197 4.5005
R6952 CSoutput.n200 CSoutput.n174 4.5005
R6953 CSoutput.n200 CSoutput.n181 4.5005
R6954 CSoutput.n200 CSoutput.n182 4.5005
R6955 CSoutput.n204 CSoutput.n177 4.5005
R6956 CSoutput.n204 CSoutput.n179 4.5005
R6957 CSoutput.n204 CSoutput.n176 4.5005
R6958 CSoutput.n204 CSoutput.n180 4.5005
R6959 CSoutput.n204 CSoutput.n175 4.5005
R6960 CSoutput.n204 CSoutput.t197 4.5005
R6961 CSoutput.n204 CSoutput.n174 4.5005
R6962 CSoutput.n204 CSoutput.n181 4.5005
R6963 CSoutput.n204 CSoutput.n182 4.5005
R6964 CSoutput.n203 CSoutput.n177 4.5005
R6965 CSoutput.n203 CSoutput.n179 4.5005
R6966 CSoutput.n203 CSoutput.n176 4.5005
R6967 CSoutput.n203 CSoutput.n180 4.5005
R6968 CSoutput.n203 CSoutput.n175 4.5005
R6969 CSoutput.n203 CSoutput.t197 4.5005
R6970 CSoutput.n203 CSoutput.n174 4.5005
R6971 CSoutput.n203 CSoutput.n181 4.5005
R6972 CSoutput.n203 CSoutput.n182 4.5005
R6973 CSoutput.n186 CSoutput.n177 4.5005
R6974 CSoutput.n186 CSoutput.n179 4.5005
R6975 CSoutput.n186 CSoutput.n176 4.5005
R6976 CSoutput.n186 CSoutput.n180 4.5005
R6977 CSoutput.n186 CSoutput.n175 4.5005
R6978 CSoutput.n186 CSoutput.t197 4.5005
R6979 CSoutput.n186 CSoutput.n174 4.5005
R6980 CSoutput.n186 CSoutput.n181 4.5005
R6981 CSoutput.n186 CSoutput.n182 4.5005
R6982 CSoutput.n278 CSoutput.n177 4.5005
R6983 CSoutput.n278 CSoutput.n179 4.5005
R6984 CSoutput.n278 CSoutput.n176 4.5005
R6985 CSoutput.n278 CSoutput.n180 4.5005
R6986 CSoutput.n278 CSoutput.n175 4.5005
R6987 CSoutput.n278 CSoutput.t197 4.5005
R6988 CSoutput.n278 CSoutput.n174 4.5005
R6989 CSoutput.n278 CSoutput.n181 4.5005
R6990 CSoutput.n278 CSoutput.n182 4.5005
R6991 CSoutput.n265 CSoutput.n236 4.5005
R6992 CSoutput.n265 CSoutput.n242 4.5005
R6993 CSoutput.n223 CSoutput.n212 4.5005
R6994 CSoutput.n223 CSoutput.n214 4.5005
R6995 CSoutput.n223 CSoutput.n211 4.5005
R6996 CSoutput.n223 CSoutput.n215 4.5005
R6997 CSoutput.n223 CSoutput.n210 4.5005
R6998 CSoutput.n223 CSoutput.t193 4.5005
R6999 CSoutput.n223 CSoutput.n209 4.5005
R7000 CSoutput.n223 CSoutput.n216 4.5005
R7001 CSoutput.n265 CSoutput.n223 4.5005
R7002 CSoutput.n244 CSoutput.n212 4.5005
R7003 CSoutput.n244 CSoutput.n214 4.5005
R7004 CSoutput.n244 CSoutput.n211 4.5005
R7005 CSoutput.n244 CSoutput.n215 4.5005
R7006 CSoutput.n244 CSoutput.n210 4.5005
R7007 CSoutput.n244 CSoutput.t193 4.5005
R7008 CSoutput.n244 CSoutput.n209 4.5005
R7009 CSoutput.n244 CSoutput.n216 4.5005
R7010 CSoutput.n265 CSoutput.n244 4.5005
R7011 CSoutput.n222 CSoutput.n212 4.5005
R7012 CSoutput.n222 CSoutput.n214 4.5005
R7013 CSoutput.n222 CSoutput.n211 4.5005
R7014 CSoutput.n222 CSoutput.n215 4.5005
R7015 CSoutput.n222 CSoutput.n210 4.5005
R7016 CSoutput.n222 CSoutput.t193 4.5005
R7017 CSoutput.n222 CSoutput.n209 4.5005
R7018 CSoutput.n222 CSoutput.n216 4.5005
R7019 CSoutput.n265 CSoutput.n222 4.5005
R7020 CSoutput.n246 CSoutput.n212 4.5005
R7021 CSoutput.n246 CSoutput.n214 4.5005
R7022 CSoutput.n246 CSoutput.n211 4.5005
R7023 CSoutput.n246 CSoutput.n215 4.5005
R7024 CSoutput.n246 CSoutput.n210 4.5005
R7025 CSoutput.n246 CSoutput.t193 4.5005
R7026 CSoutput.n246 CSoutput.n209 4.5005
R7027 CSoutput.n246 CSoutput.n216 4.5005
R7028 CSoutput.n265 CSoutput.n246 4.5005
R7029 CSoutput.n212 CSoutput.n207 4.5005
R7030 CSoutput.n214 CSoutput.n207 4.5005
R7031 CSoutput.n211 CSoutput.n207 4.5005
R7032 CSoutput.n215 CSoutput.n207 4.5005
R7033 CSoutput.n210 CSoutput.n207 4.5005
R7034 CSoutput.t193 CSoutput.n207 4.5005
R7035 CSoutput.n209 CSoutput.n207 4.5005
R7036 CSoutput.n216 CSoutput.n207 4.5005
R7037 CSoutput.n268 CSoutput.n212 4.5005
R7038 CSoutput.n268 CSoutput.n214 4.5005
R7039 CSoutput.n268 CSoutput.n211 4.5005
R7040 CSoutput.n268 CSoutput.n215 4.5005
R7041 CSoutput.n268 CSoutput.n210 4.5005
R7042 CSoutput.n268 CSoutput.t193 4.5005
R7043 CSoutput.n268 CSoutput.n209 4.5005
R7044 CSoutput.n268 CSoutput.n216 4.5005
R7045 CSoutput.n266 CSoutput.n212 4.5005
R7046 CSoutput.n266 CSoutput.n214 4.5005
R7047 CSoutput.n266 CSoutput.n211 4.5005
R7048 CSoutput.n266 CSoutput.n215 4.5005
R7049 CSoutput.n266 CSoutput.n210 4.5005
R7050 CSoutput.n266 CSoutput.t193 4.5005
R7051 CSoutput.n266 CSoutput.n209 4.5005
R7052 CSoutput.n266 CSoutput.n216 4.5005
R7053 CSoutput.n266 CSoutput.n265 4.5005
R7054 CSoutput.n248 CSoutput.n212 4.5005
R7055 CSoutput.n248 CSoutput.n214 4.5005
R7056 CSoutput.n248 CSoutput.n211 4.5005
R7057 CSoutput.n248 CSoutput.n215 4.5005
R7058 CSoutput.n248 CSoutput.n210 4.5005
R7059 CSoutput.n248 CSoutput.t193 4.5005
R7060 CSoutput.n248 CSoutput.n209 4.5005
R7061 CSoutput.n248 CSoutput.n216 4.5005
R7062 CSoutput.n265 CSoutput.n248 4.5005
R7063 CSoutput.n220 CSoutput.n212 4.5005
R7064 CSoutput.n220 CSoutput.n214 4.5005
R7065 CSoutput.n220 CSoutput.n211 4.5005
R7066 CSoutput.n220 CSoutput.n215 4.5005
R7067 CSoutput.n220 CSoutput.n210 4.5005
R7068 CSoutput.n220 CSoutput.t193 4.5005
R7069 CSoutput.n220 CSoutput.n209 4.5005
R7070 CSoutput.n220 CSoutput.n216 4.5005
R7071 CSoutput.n265 CSoutput.n220 4.5005
R7072 CSoutput.n250 CSoutput.n212 4.5005
R7073 CSoutput.n250 CSoutput.n214 4.5005
R7074 CSoutput.n250 CSoutput.n211 4.5005
R7075 CSoutput.n250 CSoutput.n215 4.5005
R7076 CSoutput.n250 CSoutput.n210 4.5005
R7077 CSoutput.n250 CSoutput.t193 4.5005
R7078 CSoutput.n250 CSoutput.n209 4.5005
R7079 CSoutput.n250 CSoutput.n216 4.5005
R7080 CSoutput.n265 CSoutput.n250 4.5005
R7081 CSoutput.n219 CSoutput.n212 4.5005
R7082 CSoutput.n219 CSoutput.n214 4.5005
R7083 CSoutput.n219 CSoutput.n211 4.5005
R7084 CSoutput.n219 CSoutput.n215 4.5005
R7085 CSoutput.n219 CSoutput.n210 4.5005
R7086 CSoutput.n219 CSoutput.t193 4.5005
R7087 CSoutput.n219 CSoutput.n209 4.5005
R7088 CSoutput.n219 CSoutput.n216 4.5005
R7089 CSoutput.n265 CSoutput.n219 4.5005
R7090 CSoutput.n264 CSoutput.n212 4.5005
R7091 CSoutput.n264 CSoutput.n214 4.5005
R7092 CSoutput.n264 CSoutput.n211 4.5005
R7093 CSoutput.n264 CSoutput.n215 4.5005
R7094 CSoutput.n264 CSoutput.n210 4.5005
R7095 CSoutput.n264 CSoutput.t193 4.5005
R7096 CSoutput.n264 CSoutput.n209 4.5005
R7097 CSoutput.n264 CSoutput.n216 4.5005
R7098 CSoutput.n265 CSoutput.n264 4.5005
R7099 CSoutput.n263 CSoutput.n148 4.5005
R7100 CSoutput.n164 CSoutput.n148 4.5005
R7101 CSoutput.n159 CSoutput.n143 4.5005
R7102 CSoutput.n159 CSoutput.n145 4.5005
R7103 CSoutput.n159 CSoutput.n142 4.5005
R7104 CSoutput.n159 CSoutput.n146 4.5005
R7105 CSoutput.n159 CSoutput.n141 4.5005
R7106 CSoutput.n159 CSoutput.t213 4.5005
R7107 CSoutput.n159 CSoutput.n140 4.5005
R7108 CSoutput.n159 CSoutput.n147 4.5005
R7109 CSoutput.n159 CSoutput.n148 4.5005
R7110 CSoutput.n157 CSoutput.n143 4.5005
R7111 CSoutput.n157 CSoutput.n145 4.5005
R7112 CSoutput.n157 CSoutput.n142 4.5005
R7113 CSoutput.n157 CSoutput.n146 4.5005
R7114 CSoutput.n157 CSoutput.n141 4.5005
R7115 CSoutput.n157 CSoutput.t213 4.5005
R7116 CSoutput.n157 CSoutput.n140 4.5005
R7117 CSoutput.n157 CSoutput.n147 4.5005
R7118 CSoutput.n157 CSoutput.n148 4.5005
R7119 CSoutput.n156 CSoutput.n143 4.5005
R7120 CSoutput.n156 CSoutput.n145 4.5005
R7121 CSoutput.n156 CSoutput.n142 4.5005
R7122 CSoutput.n156 CSoutput.n146 4.5005
R7123 CSoutput.n156 CSoutput.n141 4.5005
R7124 CSoutput.n156 CSoutput.t213 4.5005
R7125 CSoutput.n156 CSoutput.n140 4.5005
R7126 CSoutput.n156 CSoutput.n147 4.5005
R7127 CSoutput.n156 CSoutput.n148 4.5005
R7128 CSoutput.n285 CSoutput.n143 4.5005
R7129 CSoutput.n285 CSoutput.n145 4.5005
R7130 CSoutput.n285 CSoutput.n142 4.5005
R7131 CSoutput.n285 CSoutput.n146 4.5005
R7132 CSoutput.n285 CSoutput.n141 4.5005
R7133 CSoutput.n285 CSoutput.t213 4.5005
R7134 CSoutput.n285 CSoutput.n140 4.5005
R7135 CSoutput.n285 CSoutput.n147 4.5005
R7136 CSoutput.n285 CSoutput.n148 4.5005
R7137 CSoutput.n283 CSoutput.n143 4.5005
R7138 CSoutput.n283 CSoutput.n145 4.5005
R7139 CSoutput.n283 CSoutput.n142 4.5005
R7140 CSoutput.n283 CSoutput.n146 4.5005
R7141 CSoutput.n283 CSoutput.n141 4.5005
R7142 CSoutput.n283 CSoutput.t213 4.5005
R7143 CSoutput.n283 CSoutput.n140 4.5005
R7144 CSoutput.n283 CSoutput.n147 4.5005
R7145 CSoutput.n281 CSoutput.n143 4.5005
R7146 CSoutput.n281 CSoutput.n145 4.5005
R7147 CSoutput.n281 CSoutput.n142 4.5005
R7148 CSoutput.n281 CSoutput.n146 4.5005
R7149 CSoutput.n281 CSoutput.n141 4.5005
R7150 CSoutput.n281 CSoutput.t213 4.5005
R7151 CSoutput.n281 CSoutput.n140 4.5005
R7152 CSoutput.n281 CSoutput.n147 4.5005
R7153 CSoutput.n167 CSoutput.n143 4.5005
R7154 CSoutput.n167 CSoutput.n145 4.5005
R7155 CSoutput.n167 CSoutput.n142 4.5005
R7156 CSoutput.n167 CSoutput.n146 4.5005
R7157 CSoutput.n167 CSoutput.n141 4.5005
R7158 CSoutput.n167 CSoutput.t213 4.5005
R7159 CSoutput.n167 CSoutput.n140 4.5005
R7160 CSoutput.n167 CSoutput.n147 4.5005
R7161 CSoutput.n167 CSoutput.n148 4.5005
R7162 CSoutput.n166 CSoutput.n143 4.5005
R7163 CSoutput.n166 CSoutput.n145 4.5005
R7164 CSoutput.n166 CSoutput.n142 4.5005
R7165 CSoutput.n166 CSoutput.n146 4.5005
R7166 CSoutput.n166 CSoutput.n141 4.5005
R7167 CSoutput.n166 CSoutput.t213 4.5005
R7168 CSoutput.n166 CSoutput.n140 4.5005
R7169 CSoutput.n166 CSoutput.n147 4.5005
R7170 CSoutput.n166 CSoutput.n148 4.5005
R7171 CSoutput.n170 CSoutput.n143 4.5005
R7172 CSoutput.n170 CSoutput.n145 4.5005
R7173 CSoutput.n170 CSoutput.n142 4.5005
R7174 CSoutput.n170 CSoutput.n146 4.5005
R7175 CSoutput.n170 CSoutput.n141 4.5005
R7176 CSoutput.n170 CSoutput.t213 4.5005
R7177 CSoutput.n170 CSoutput.n140 4.5005
R7178 CSoutput.n170 CSoutput.n147 4.5005
R7179 CSoutput.n170 CSoutput.n148 4.5005
R7180 CSoutput.n169 CSoutput.n143 4.5005
R7181 CSoutput.n169 CSoutput.n145 4.5005
R7182 CSoutput.n169 CSoutput.n142 4.5005
R7183 CSoutput.n169 CSoutput.n146 4.5005
R7184 CSoutput.n169 CSoutput.n141 4.5005
R7185 CSoutput.n169 CSoutput.t213 4.5005
R7186 CSoutput.n169 CSoutput.n140 4.5005
R7187 CSoutput.n169 CSoutput.n147 4.5005
R7188 CSoutput.n169 CSoutput.n148 4.5005
R7189 CSoutput.n152 CSoutput.n143 4.5005
R7190 CSoutput.n152 CSoutput.n145 4.5005
R7191 CSoutput.n152 CSoutput.n142 4.5005
R7192 CSoutput.n152 CSoutput.n146 4.5005
R7193 CSoutput.n152 CSoutput.n141 4.5005
R7194 CSoutput.n152 CSoutput.t213 4.5005
R7195 CSoutput.n152 CSoutput.n140 4.5005
R7196 CSoutput.n152 CSoutput.n147 4.5005
R7197 CSoutput.n152 CSoutput.n148 4.5005
R7198 CSoutput.n288 CSoutput.n143 4.5005
R7199 CSoutput.n288 CSoutput.n145 4.5005
R7200 CSoutput.n288 CSoutput.n142 4.5005
R7201 CSoutput.n288 CSoutput.n146 4.5005
R7202 CSoutput.n288 CSoutput.n141 4.5005
R7203 CSoutput.n288 CSoutput.t213 4.5005
R7204 CSoutput.n288 CSoutput.n140 4.5005
R7205 CSoutput.n288 CSoutput.n147 4.5005
R7206 CSoutput.n288 CSoutput.n148 4.5005
R7207 CSoutput.n347 CSoutput.n327 4.10845
R7208 CSoutput.n137 CSoutput.n117 4.10845
R7209 CSoutput.n345 CSoutput.t155 4.06363
R7210 CSoutput.n345 CSoutput.t73 4.06363
R7211 CSoutput.n343 CSoutput.t66 4.06363
R7212 CSoutput.n343 CSoutput.t117 4.06363
R7213 CSoutput.n341 CSoutput.t134 4.06363
R7214 CSoutput.n341 CSoutput.t158 4.06363
R7215 CSoutput.n339 CSoutput.t173 4.06363
R7216 CSoutput.n339 CSoutput.t86 4.06363
R7217 CSoutput.n337 CSoutput.t90 4.06363
R7218 CSoutput.n337 CSoutput.t162 4.06363
R7219 CSoutput.n335 CSoutput.t177 4.06363
R7220 CSoutput.n335 CSoutput.t178 4.06363
R7221 CSoutput.n333 CSoutput.t111 4.06363
R7222 CSoutput.n333 CSoutput.t112 4.06363
R7223 CSoutput.n331 CSoutput.t119 4.06363
R7224 CSoutput.n331 CSoutput.t179 4.06363
R7225 CSoutput.n329 CSoutput.t78 4.06363
R7226 CSoutput.n329 CSoutput.t116 4.06363
R7227 CSoutput.n328 CSoutput.t133 4.06363
R7228 CSoutput.n328 CSoutput.t157 4.06363
R7229 CSoutput.n325 CSoutput.t144 4.06363
R7230 CSoutput.n325 CSoutput.t180 4.06363
R7231 CSoutput.n323 CSoutput.t175 4.06363
R7232 CSoutput.n323 CSoutput.t100 4.06363
R7233 CSoutput.n321 CSoutput.t121 4.06363
R7234 CSoutput.n321 CSoutput.t145 4.06363
R7235 CSoutput.n319 CSoutput.t163 4.06363
R7236 CSoutput.n319 CSoutput.t72 4.06363
R7237 CSoutput.n317 CSoutput.t74 4.06363
R7238 CSoutput.n317 CSoutput.t149 4.06363
R7239 CSoutput.n315 CSoutput.t166 4.06363
R7240 CSoutput.n315 CSoutput.t167 4.06363
R7241 CSoutput.n313 CSoutput.t94 4.06363
R7242 CSoutput.n313 CSoutput.t95 4.06363
R7243 CSoutput.n311 CSoutput.t102 4.06363
R7244 CSoutput.n311 CSoutput.t168 4.06363
R7245 CSoutput.n309 CSoutput.t64 4.06363
R7246 CSoutput.n309 CSoutput.t101 4.06363
R7247 CSoutput.n308 CSoutput.t122 4.06363
R7248 CSoutput.n308 CSoutput.t146 4.06363
R7249 CSoutput.n306 CSoutput.t147 4.06363
R7250 CSoutput.n306 CSoutput.t98 4.06363
R7251 CSoutput.n304 CSoutput.t169 4.06363
R7252 CSoutput.n304 CSoutput.t126 4.06363
R7253 CSoutput.n302 CSoutput.t156 4.06363
R7254 CSoutput.n302 CSoutput.t108 4.06363
R7255 CSoutput.n300 CSoutput.t140 4.06363
R7256 CSoutput.n300 CSoutput.t85 4.06363
R7257 CSoutput.n298 CSoutput.t164 4.06363
R7258 CSoutput.n298 CSoutput.t79 4.06363
R7259 CSoutput.n296 CSoutput.t123 4.06363
R7260 CSoutput.n296 CSoutput.t96 4.06363
R7261 CSoutput.n294 CSoutput.t103 4.06363
R7262 CSoutput.n294 CSoutput.t75 4.06363
R7263 CSoutput.n292 CSoutput.t154 4.06363
R7264 CSoutput.n292 CSoutput.t69 4.06363
R7265 CSoutput.n290 CSoutput.t113 4.06363
R7266 CSoutput.n290 CSoutput.t174 4.06363
R7267 CSoutput.n289 CSoutput.t91 4.06363
R7268 CSoutput.n289 CSoutput.t160 4.06363
R7269 CSoutput.n118 CSoutput.t82 4.06363
R7270 CSoutput.n118 CSoutput.t171 4.06363
R7271 CSoutput.n119 CSoutput.t152 4.06363
R7272 CSoutput.n119 CSoutput.t130 4.06363
R7273 CSoutput.n121 CSoutput.t110 4.06363
R7274 CSoutput.n121 CSoutput.t182 4.06363
R7275 CSoutput.n123 CSoutput.t151 4.06363
R7276 CSoutput.n123 CSoutput.t150 4.06363
R7277 CSoutput.n125 CSoutput.t136 4.06363
R7278 CSoutput.n125 CSoutput.t107 4.06363
R7279 CSoutput.n127 CSoutput.t84 4.06363
R7280 CSoutput.n127 CSoutput.t137 4.06363
R7281 CSoutput.n129 CSoutput.t135 4.06363
R7282 CSoutput.n129 CSoutput.t104 4.06363
R7283 CSoutput.n131 CSoutput.t83 4.06363
R7284 CSoutput.n131 CSoutput.t81 4.06363
R7285 CSoutput.n133 CSoutput.t153 4.06363
R7286 CSoutput.n133 CSoutput.t120 4.06363
R7287 CSoutput.n135 CSoutput.t115 4.06363
R7288 CSoutput.n135 CSoutput.t76 4.06363
R7289 CSoutput.n98 CSoutput.t67 4.06363
R7290 CSoutput.n98 CSoutput.t159 4.06363
R7291 CSoutput.n99 CSoutput.t142 4.06363
R7292 CSoutput.n99 CSoutput.t118 4.06363
R7293 CSoutput.n101 CSoutput.t93 4.06363
R7294 CSoutput.n101 CSoutput.t172 4.06363
R7295 CSoutput.n103 CSoutput.t139 4.06363
R7296 CSoutput.n103 CSoutput.t138 4.06363
R7297 CSoutput.n105 CSoutput.t128 4.06363
R7298 CSoutput.n105 CSoutput.t89 4.06363
R7299 CSoutput.n107 CSoutput.t70 4.06363
R7300 CSoutput.n107 CSoutput.t129 4.06363
R7301 CSoutput.n109 CSoutput.t125 4.06363
R7302 CSoutput.n109 CSoutput.t87 4.06363
R7303 CSoutput.n111 CSoutput.t68 4.06363
R7304 CSoutput.n111 CSoutput.t65 4.06363
R7305 CSoutput.n113 CSoutput.t143 4.06363
R7306 CSoutput.n113 CSoutput.t106 4.06363
R7307 CSoutput.n115 CSoutput.t99 4.06363
R7308 CSoutput.n115 CSoutput.t63 4.06363
R7309 CSoutput.n79 CSoutput.t161 4.06363
R7310 CSoutput.n79 CSoutput.t92 4.06363
R7311 CSoutput.n80 CSoutput.t176 4.06363
R7312 CSoutput.n80 CSoutput.t114 4.06363
R7313 CSoutput.n82 CSoutput.t71 4.06363
R7314 CSoutput.n82 CSoutput.t131 4.06363
R7315 CSoutput.n84 CSoutput.t77 4.06363
R7316 CSoutput.n84 CSoutput.t105 4.06363
R7317 CSoutput.n86 CSoutput.t181 4.06363
R7318 CSoutput.n86 CSoutput.t124 4.06363
R7319 CSoutput.n88 CSoutput.t80 4.06363
R7320 CSoutput.n88 CSoutput.t165 4.06363
R7321 CSoutput.n90 CSoutput.t88 4.06363
R7322 CSoutput.n90 CSoutput.t141 4.06363
R7323 CSoutput.n92 CSoutput.t109 4.06363
R7324 CSoutput.n92 CSoutput.t132 4.06363
R7325 CSoutput.n94 CSoutput.t127 4.06363
R7326 CSoutput.n94 CSoutput.t170 4.06363
R7327 CSoutput.n96 CSoutput.t97 4.06363
R7328 CSoutput.n96 CSoutput.t148 4.06363
R7329 CSoutput.n44 CSoutput.n43 3.79402
R7330 CSoutput.n49 CSoutput.n48 3.79402
R7331 CSoutput.n383 CSoutput.n371 3.72967
R7332 CSoutput.n419 CSoutput.n407 3.72967
R7333 CSoutput.n421 CSoutput.n420 3.57343
R7334 CSoutput.n381 CSoutput.t42 2.82907
R7335 CSoutput.n381 CSoutput.t38 2.82907
R7336 CSoutput.n379 CSoutput.t43 2.82907
R7337 CSoutput.n379 CSoutput.t186 2.82907
R7338 CSoutput.n377 CSoutput.t47 2.82907
R7339 CSoutput.n377 CSoutput.t49 2.82907
R7340 CSoutput.n375 CSoutput.t59 2.82907
R7341 CSoutput.n375 CSoutput.t35 2.82907
R7342 CSoutput.n373 CSoutput.t36 2.82907
R7343 CSoutput.n373 CSoutput.t62 2.82907
R7344 CSoutput.n372 CSoutput.t50 2.82907
R7345 CSoutput.n372 CSoutput.t23 2.82907
R7346 CSoutput.n369 CSoutput.t27 2.82907
R7347 CSoutput.n369 CSoutput.t3 2.82907
R7348 CSoutput.n367 CSoutput.t6 2.82907
R7349 CSoutput.n367 CSoutput.t189 2.82907
R7350 CSoutput.n365 CSoutput.t16 2.82907
R7351 CSoutput.n365 CSoutput.t190 2.82907
R7352 CSoutput.n363 CSoutput.t28 2.82907
R7353 CSoutput.n363 CSoutput.t48 2.82907
R7354 CSoutput.n361 CSoutput.t56 2.82907
R7355 CSoutput.n361 CSoutput.t51 2.82907
R7356 CSoutput.n360 CSoutput.t29 2.82907
R7357 CSoutput.n360 CSoutput.t191 2.82907
R7358 CSoutput.n358 CSoutput.t24 2.82907
R7359 CSoutput.n358 CSoutput.t8 2.82907
R7360 CSoutput.n356 CSoutput.t187 2.82907
R7361 CSoutput.n356 CSoutput.t185 2.82907
R7362 CSoutput.n354 CSoutput.t21 2.82907
R7363 CSoutput.n354 CSoutput.t54 2.82907
R7364 CSoutput.n352 CSoutput.t41 2.82907
R7365 CSoutput.n352 CSoutput.t13 2.82907
R7366 CSoutput.n350 CSoutput.t55 2.82907
R7367 CSoutput.n350 CSoutput.t15 2.82907
R7368 CSoutput.n349 CSoutput.t5 2.82907
R7369 CSoutput.n349 CSoutput.t33 2.82907
R7370 CSoutput.n408 CSoutput.t18 2.82907
R7371 CSoutput.n408 CSoutput.t1 2.82907
R7372 CSoutput.n409 CSoutput.t40 2.82907
R7373 CSoutput.n409 CSoutput.t184 2.82907
R7374 CSoutput.n411 CSoutput.t53 2.82907
R7375 CSoutput.n411 CSoutput.t25 2.82907
R7376 CSoutput.n413 CSoutput.t14 2.82907
R7377 CSoutput.n413 CSoutput.t46 2.82907
R7378 CSoutput.n415 CSoutput.t0 2.82907
R7379 CSoutput.n415 CSoutput.t188 2.82907
R7380 CSoutput.n417 CSoutput.t31 2.82907
R7381 CSoutput.n417 CSoutput.t37 2.82907
R7382 CSoutput.n396 CSoutput.t10 2.82907
R7383 CSoutput.n396 CSoutput.t30 2.82907
R7384 CSoutput.n397 CSoutput.t58 2.82907
R7385 CSoutput.n397 CSoutput.t60 2.82907
R7386 CSoutput.n399 CSoutput.t32 2.82907
R7387 CSoutput.n399 CSoutput.t9 2.82907
R7388 CSoutput.n401 CSoutput.t45 2.82907
R7389 CSoutput.n401 CSoutput.t26 2.82907
R7390 CSoutput.n403 CSoutput.t4 2.82907
R7391 CSoutput.n403 CSoutput.t12 2.82907
R7392 CSoutput.n405 CSoutput.t22 2.82907
R7393 CSoutput.n405 CSoutput.t2 2.82907
R7394 CSoutput.n385 CSoutput.t39 2.82907
R7395 CSoutput.n385 CSoutput.t183 2.82907
R7396 CSoutput.n386 CSoutput.t11 2.82907
R7397 CSoutput.n386 CSoutput.t7 2.82907
R7398 CSoutput.n388 CSoutput.t34 2.82907
R7399 CSoutput.n388 CSoutput.t61 2.82907
R7400 CSoutput.n390 CSoutput.t17 2.82907
R7401 CSoutput.n390 CSoutput.t52 2.82907
R7402 CSoutput.n392 CSoutput.t44 2.82907
R7403 CSoutput.n392 CSoutput.t20 2.82907
R7404 CSoutput.n394 CSoutput.t57 2.82907
R7405 CSoutput.n394 CSoutput.t19 2.82907
R7406 CSoutput.n348 CSoutput.n138 2.78353
R7407 CSoutput.n420 CSoutput.n384 2.75627
R7408 CSoutput.n75 CSoutput.n1 2.45513
R7409 CSoutput.n229 CSoutput.n227 2.251
R7410 CSoutput.n229 CSoutput.n226 2.251
R7411 CSoutput.n229 CSoutput.n225 2.251
R7412 CSoutput.n229 CSoutput.n224 2.251
R7413 CSoutput.n198 CSoutput.n197 2.251
R7414 CSoutput.n198 CSoutput.n196 2.251
R7415 CSoutput.n198 CSoutput.n195 2.251
R7416 CSoutput.n198 CSoutput.n194 2.251
R7417 CSoutput.n271 CSoutput.n270 2.251
R7418 CSoutput.n236 CSoutput.n234 2.251
R7419 CSoutput.n236 CSoutput.n233 2.251
R7420 CSoutput.n236 CSoutput.n232 2.251
R7421 CSoutput.n254 CSoutput.n236 2.251
R7422 CSoutput.n242 CSoutput.n241 2.251
R7423 CSoutput.n242 CSoutput.n240 2.251
R7424 CSoutput.n242 CSoutput.n239 2.251
R7425 CSoutput.n242 CSoutput.n238 2.251
R7426 CSoutput.n268 CSoutput.n208 2.251
R7427 CSoutput.n263 CSoutput.n261 2.251
R7428 CSoutput.n263 CSoutput.n260 2.251
R7429 CSoutput.n263 CSoutput.n259 2.251
R7430 CSoutput.n263 CSoutput.n258 2.251
R7431 CSoutput.n164 CSoutput.n163 2.251
R7432 CSoutput.n164 CSoutput.n162 2.251
R7433 CSoutput.n164 CSoutput.n161 2.251
R7434 CSoutput.n164 CSoutput.n160 2.251
R7435 CSoutput.n281 CSoutput.n280 2.251
R7436 CSoutput.n198 CSoutput.n178 2.2505
R7437 CSoutput.n193 CSoutput.n178 2.2505
R7438 CSoutput.n191 CSoutput.n178 2.2505
R7439 CSoutput.n190 CSoutput.n178 2.2505
R7440 CSoutput.n275 CSoutput.n178 2.2505
R7441 CSoutput.n273 CSoutput.n178 2.2505
R7442 CSoutput.n271 CSoutput.n178 2.2505
R7443 CSoutput.n201 CSoutput.n178 2.2505
R7444 CSoutput.n200 CSoutput.n178 2.2505
R7445 CSoutput.n204 CSoutput.n178 2.2505
R7446 CSoutput.n203 CSoutput.n178 2.2505
R7447 CSoutput.n186 CSoutput.n178 2.2505
R7448 CSoutput.n278 CSoutput.n178 2.2505
R7449 CSoutput.n278 CSoutput.n277 2.2505
R7450 CSoutput.n242 CSoutput.n213 2.2505
R7451 CSoutput.n223 CSoutput.n213 2.2505
R7452 CSoutput.n244 CSoutput.n213 2.2505
R7453 CSoutput.n222 CSoutput.n213 2.2505
R7454 CSoutput.n246 CSoutput.n213 2.2505
R7455 CSoutput.n213 CSoutput.n207 2.2505
R7456 CSoutput.n268 CSoutput.n213 2.2505
R7457 CSoutput.n266 CSoutput.n213 2.2505
R7458 CSoutput.n248 CSoutput.n213 2.2505
R7459 CSoutput.n220 CSoutput.n213 2.2505
R7460 CSoutput.n250 CSoutput.n213 2.2505
R7461 CSoutput.n219 CSoutput.n213 2.2505
R7462 CSoutput.n264 CSoutput.n213 2.2505
R7463 CSoutput.n264 CSoutput.n217 2.2505
R7464 CSoutput.n164 CSoutput.n144 2.2505
R7465 CSoutput.n159 CSoutput.n144 2.2505
R7466 CSoutput.n157 CSoutput.n144 2.2505
R7467 CSoutput.n156 CSoutput.n144 2.2505
R7468 CSoutput.n285 CSoutput.n144 2.2505
R7469 CSoutput.n283 CSoutput.n144 2.2505
R7470 CSoutput.n281 CSoutput.n144 2.2505
R7471 CSoutput.n167 CSoutput.n144 2.2505
R7472 CSoutput.n166 CSoutput.n144 2.2505
R7473 CSoutput.n170 CSoutput.n144 2.2505
R7474 CSoutput.n169 CSoutput.n144 2.2505
R7475 CSoutput.n152 CSoutput.n144 2.2505
R7476 CSoutput.n288 CSoutput.n144 2.2505
R7477 CSoutput.n288 CSoutput.n287 2.2505
R7478 CSoutput.n206 CSoutput.n199 2.25024
R7479 CSoutput.n206 CSoutput.n192 2.25024
R7480 CSoutput.n274 CSoutput.n206 2.25024
R7481 CSoutput.n206 CSoutput.n202 2.25024
R7482 CSoutput.n206 CSoutput.n205 2.25024
R7483 CSoutput.n206 CSoutput.n173 2.25024
R7484 CSoutput.n256 CSoutput.n253 2.25024
R7485 CSoutput.n256 CSoutput.n252 2.25024
R7486 CSoutput.n256 CSoutput.n251 2.25024
R7487 CSoutput.n256 CSoutput.n218 2.25024
R7488 CSoutput.n256 CSoutput.n255 2.25024
R7489 CSoutput.n257 CSoutput.n256 2.25024
R7490 CSoutput.n172 CSoutput.n165 2.25024
R7491 CSoutput.n172 CSoutput.n158 2.25024
R7492 CSoutput.n284 CSoutput.n172 2.25024
R7493 CSoutput.n172 CSoutput.n168 2.25024
R7494 CSoutput.n172 CSoutput.n171 2.25024
R7495 CSoutput.n172 CSoutput.n139 2.25024
R7496 CSoutput.n273 CSoutput.n183 1.50111
R7497 CSoutput.n221 CSoutput.n207 1.50111
R7498 CSoutput.n283 CSoutput.n149 1.50111
R7499 CSoutput.n229 CSoutput.n228 1.501
R7500 CSoutput.n236 CSoutput.n235 1.501
R7501 CSoutput.n263 CSoutput.n262 1.501
R7502 CSoutput.n277 CSoutput.n188 1.12536
R7503 CSoutput.n277 CSoutput.n189 1.12536
R7504 CSoutput.n277 CSoutput.n276 1.12536
R7505 CSoutput.n237 CSoutput.n217 1.12536
R7506 CSoutput.n243 CSoutput.n217 1.12536
R7507 CSoutput.n245 CSoutput.n217 1.12536
R7508 CSoutput.n287 CSoutput.n154 1.12536
R7509 CSoutput.n287 CSoutput.n155 1.12536
R7510 CSoutput.n287 CSoutput.n286 1.12536
R7511 CSoutput.n277 CSoutput.n184 1.12536
R7512 CSoutput.n277 CSoutput.n185 1.12536
R7513 CSoutput.n277 CSoutput.n187 1.12536
R7514 CSoutput.n267 CSoutput.n217 1.12536
R7515 CSoutput.n247 CSoutput.n217 1.12536
R7516 CSoutput.n249 CSoutput.n217 1.12536
R7517 CSoutput.n287 CSoutput.n150 1.12536
R7518 CSoutput.n287 CSoutput.n151 1.12536
R7519 CSoutput.n287 CSoutput.n153 1.12536
R7520 CSoutput.n31 CSoutput.n30 0.669944
R7521 CSoutput.n62 CSoutput.n61 0.669944
R7522 CSoutput.n376 CSoutput.n374 0.573776
R7523 CSoutput.n378 CSoutput.n376 0.573776
R7524 CSoutput.n380 CSoutput.n378 0.573776
R7525 CSoutput.n382 CSoutput.n380 0.573776
R7526 CSoutput.n364 CSoutput.n362 0.573776
R7527 CSoutput.n366 CSoutput.n364 0.573776
R7528 CSoutput.n368 CSoutput.n366 0.573776
R7529 CSoutput.n370 CSoutput.n368 0.573776
R7530 CSoutput.n353 CSoutput.n351 0.573776
R7531 CSoutput.n355 CSoutput.n353 0.573776
R7532 CSoutput.n357 CSoutput.n355 0.573776
R7533 CSoutput.n359 CSoutput.n357 0.573776
R7534 CSoutput.n418 CSoutput.n416 0.573776
R7535 CSoutput.n416 CSoutput.n414 0.573776
R7536 CSoutput.n414 CSoutput.n412 0.573776
R7537 CSoutput.n412 CSoutput.n410 0.573776
R7538 CSoutput.n406 CSoutput.n404 0.573776
R7539 CSoutput.n404 CSoutput.n402 0.573776
R7540 CSoutput.n402 CSoutput.n400 0.573776
R7541 CSoutput.n400 CSoutput.n398 0.573776
R7542 CSoutput.n395 CSoutput.n393 0.573776
R7543 CSoutput.n393 CSoutput.n391 0.573776
R7544 CSoutput.n391 CSoutput.n389 0.573776
R7545 CSoutput.n389 CSoutput.n387 0.573776
R7546 CSoutput.n421 CSoutput.n288 0.53442
R7547 CSoutput.n332 CSoutput.n330 0.358259
R7548 CSoutput.n334 CSoutput.n332 0.358259
R7549 CSoutput.n336 CSoutput.n334 0.358259
R7550 CSoutput.n338 CSoutput.n336 0.358259
R7551 CSoutput.n340 CSoutput.n338 0.358259
R7552 CSoutput.n342 CSoutput.n340 0.358259
R7553 CSoutput.n344 CSoutput.n342 0.358259
R7554 CSoutput.n346 CSoutput.n344 0.358259
R7555 CSoutput.n312 CSoutput.n310 0.358259
R7556 CSoutput.n314 CSoutput.n312 0.358259
R7557 CSoutput.n316 CSoutput.n314 0.358259
R7558 CSoutput.n318 CSoutput.n316 0.358259
R7559 CSoutput.n320 CSoutput.n318 0.358259
R7560 CSoutput.n322 CSoutput.n320 0.358259
R7561 CSoutput.n324 CSoutput.n322 0.358259
R7562 CSoutput.n326 CSoutput.n324 0.358259
R7563 CSoutput.n293 CSoutput.n291 0.358259
R7564 CSoutput.n295 CSoutput.n293 0.358259
R7565 CSoutput.n297 CSoutput.n295 0.358259
R7566 CSoutput.n299 CSoutput.n297 0.358259
R7567 CSoutput.n301 CSoutput.n299 0.358259
R7568 CSoutput.n303 CSoutput.n301 0.358259
R7569 CSoutput.n305 CSoutput.n303 0.358259
R7570 CSoutput.n307 CSoutput.n305 0.358259
R7571 CSoutput.n136 CSoutput.n134 0.358259
R7572 CSoutput.n134 CSoutput.n132 0.358259
R7573 CSoutput.n132 CSoutput.n130 0.358259
R7574 CSoutput.n130 CSoutput.n128 0.358259
R7575 CSoutput.n128 CSoutput.n126 0.358259
R7576 CSoutput.n126 CSoutput.n124 0.358259
R7577 CSoutput.n124 CSoutput.n122 0.358259
R7578 CSoutput.n122 CSoutput.n120 0.358259
R7579 CSoutput.n116 CSoutput.n114 0.358259
R7580 CSoutput.n114 CSoutput.n112 0.358259
R7581 CSoutput.n112 CSoutput.n110 0.358259
R7582 CSoutput.n110 CSoutput.n108 0.358259
R7583 CSoutput.n108 CSoutput.n106 0.358259
R7584 CSoutput.n106 CSoutput.n104 0.358259
R7585 CSoutput.n104 CSoutput.n102 0.358259
R7586 CSoutput.n102 CSoutput.n100 0.358259
R7587 CSoutput.n97 CSoutput.n95 0.358259
R7588 CSoutput.n95 CSoutput.n93 0.358259
R7589 CSoutput.n93 CSoutput.n91 0.358259
R7590 CSoutput.n91 CSoutput.n89 0.358259
R7591 CSoutput.n89 CSoutput.n87 0.358259
R7592 CSoutput.n87 CSoutput.n85 0.358259
R7593 CSoutput.n85 CSoutput.n83 0.358259
R7594 CSoutput.n83 CSoutput.n81 0.358259
R7595 CSoutput.n21 CSoutput.n20 0.169105
R7596 CSoutput.n21 CSoutput.n16 0.169105
R7597 CSoutput.n26 CSoutput.n16 0.169105
R7598 CSoutput.n27 CSoutput.n26 0.169105
R7599 CSoutput.n27 CSoutput.n14 0.169105
R7600 CSoutput.n32 CSoutput.n14 0.169105
R7601 CSoutput.n33 CSoutput.n32 0.169105
R7602 CSoutput.n34 CSoutput.n33 0.169105
R7603 CSoutput.n34 CSoutput.n12 0.169105
R7604 CSoutput.n39 CSoutput.n12 0.169105
R7605 CSoutput.n40 CSoutput.n39 0.169105
R7606 CSoutput.n40 CSoutput.n10 0.169105
R7607 CSoutput.n45 CSoutput.n10 0.169105
R7608 CSoutput.n46 CSoutput.n45 0.169105
R7609 CSoutput.n47 CSoutput.n46 0.169105
R7610 CSoutput.n47 CSoutput.n8 0.169105
R7611 CSoutput.n52 CSoutput.n8 0.169105
R7612 CSoutput.n53 CSoutput.n52 0.169105
R7613 CSoutput.n53 CSoutput.n6 0.169105
R7614 CSoutput.n58 CSoutput.n6 0.169105
R7615 CSoutput.n59 CSoutput.n58 0.169105
R7616 CSoutput.n60 CSoutput.n59 0.169105
R7617 CSoutput.n60 CSoutput.n4 0.169105
R7618 CSoutput.n66 CSoutput.n4 0.169105
R7619 CSoutput.n67 CSoutput.n66 0.169105
R7620 CSoutput.n68 CSoutput.n67 0.169105
R7621 CSoutput.n68 CSoutput.n2 0.169105
R7622 CSoutput.n73 CSoutput.n2 0.169105
R7623 CSoutput.n74 CSoutput.n73 0.169105
R7624 CSoutput.n74 CSoutput.n0 0.169105
R7625 CSoutput.n78 CSoutput.n0 0.169105
R7626 CSoutput.n231 CSoutput.n230 0.0910737
R7627 CSoutput.n282 CSoutput.n279 0.0723685
R7628 CSoutput.n236 CSoutput.n231 0.0522944
R7629 CSoutput.n279 CSoutput.n278 0.0499135
R7630 CSoutput.n230 CSoutput.n229 0.0499135
R7631 CSoutput.n264 CSoutput.n263 0.0464294
R7632 CSoutput.n272 CSoutput.n269 0.0391444
R7633 CSoutput.n231 CSoutput.t203 0.023435
R7634 CSoutput.n279 CSoutput.t201 0.02262
R7635 CSoutput.n230 CSoutput.t207 0.02262
R7636 CSoutput CSoutput.n421 0.0052
R7637 CSoutput.n201 CSoutput.n184 0.00365111
R7638 CSoutput.n204 CSoutput.n185 0.00365111
R7639 CSoutput.n187 CSoutput.n186 0.00365111
R7640 CSoutput.n229 CSoutput.n188 0.00365111
R7641 CSoutput.n193 CSoutput.n189 0.00365111
R7642 CSoutput.n276 CSoutput.n190 0.00365111
R7643 CSoutput.n267 CSoutput.n266 0.00365111
R7644 CSoutput.n247 CSoutput.n220 0.00365111
R7645 CSoutput.n249 CSoutput.n219 0.00365111
R7646 CSoutput.n237 CSoutput.n236 0.00365111
R7647 CSoutput.n243 CSoutput.n223 0.00365111
R7648 CSoutput.n245 CSoutput.n222 0.00365111
R7649 CSoutput.n167 CSoutput.n150 0.00365111
R7650 CSoutput.n170 CSoutput.n151 0.00365111
R7651 CSoutput.n153 CSoutput.n152 0.00365111
R7652 CSoutput.n263 CSoutput.n154 0.00365111
R7653 CSoutput.n159 CSoutput.n155 0.00365111
R7654 CSoutput.n286 CSoutput.n156 0.00365111
R7655 CSoutput.n198 CSoutput.n188 0.00340054
R7656 CSoutput.n191 CSoutput.n189 0.00340054
R7657 CSoutput.n276 CSoutput.n275 0.00340054
R7658 CSoutput.n271 CSoutput.n184 0.00340054
R7659 CSoutput.n200 CSoutput.n185 0.00340054
R7660 CSoutput.n203 CSoutput.n187 0.00340054
R7661 CSoutput.n242 CSoutput.n237 0.00340054
R7662 CSoutput.n244 CSoutput.n243 0.00340054
R7663 CSoutput.n246 CSoutput.n245 0.00340054
R7664 CSoutput.n268 CSoutput.n267 0.00340054
R7665 CSoutput.n248 CSoutput.n247 0.00340054
R7666 CSoutput.n250 CSoutput.n249 0.00340054
R7667 CSoutput.n164 CSoutput.n154 0.00340054
R7668 CSoutput.n157 CSoutput.n155 0.00340054
R7669 CSoutput.n286 CSoutput.n285 0.00340054
R7670 CSoutput.n281 CSoutput.n150 0.00340054
R7671 CSoutput.n166 CSoutput.n151 0.00340054
R7672 CSoutput.n169 CSoutput.n153 0.00340054
R7673 CSoutput.n199 CSoutput.n193 0.00252698
R7674 CSoutput.n192 CSoutput.n190 0.00252698
R7675 CSoutput.n274 CSoutput.n273 0.00252698
R7676 CSoutput.n202 CSoutput.n200 0.00252698
R7677 CSoutput.n205 CSoutput.n203 0.00252698
R7678 CSoutput.n278 CSoutput.n173 0.00252698
R7679 CSoutput.n199 CSoutput.n198 0.00252698
R7680 CSoutput.n192 CSoutput.n191 0.00252698
R7681 CSoutput.n275 CSoutput.n274 0.00252698
R7682 CSoutput.n202 CSoutput.n201 0.00252698
R7683 CSoutput.n205 CSoutput.n204 0.00252698
R7684 CSoutput.n186 CSoutput.n173 0.00252698
R7685 CSoutput.n253 CSoutput.n223 0.00252698
R7686 CSoutput.n252 CSoutput.n222 0.00252698
R7687 CSoutput.n251 CSoutput.n207 0.00252698
R7688 CSoutput.n248 CSoutput.n218 0.00252698
R7689 CSoutput.n255 CSoutput.n250 0.00252698
R7690 CSoutput.n264 CSoutput.n257 0.00252698
R7691 CSoutput.n253 CSoutput.n242 0.00252698
R7692 CSoutput.n252 CSoutput.n244 0.00252698
R7693 CSoutput.n251 CSoutput.n246 0.00252698
R7694 CSoutput.n266 CSoutput.n218 0.00252698
R7695 CSoutput.n255 CSoutput.n220 0.00252698
R7696 CSoutput.n257 CSoutput.n219 0.00252698
R7697 CSoutput.n165 CSoutput.n159 0.00252698
R7698 CSoutput.n158 CSoutput.n156 0.00252698
R7699 CSoutput.n284 CSoutput.n283 0.00252698
R7700 CSoutput.n168 CSoutput.n166 0.00252698
R7701 CSoutput.n171 CSoutput.n169 0.00252698
R7702 CSoutput.n288 CSoutput.n139 0.00252698
R7703 CSoutput.n165 CSoutput.n164 0.00252698
R7704 CSoutput.n158 CSoutput.n157 0.00252698
R7705 CSoutput.n285 CSoutput.n284 0.00252698
R7706 CSoutput.n168 CSoutput.n167 0.00252698
R7707 CSoutput.n171 CSoutput.n170 0.00252698
R7708 CSoutput.n152 CSoutput.n139 0.00252698
R7709 CSoutput.n273 CSoutput.n272 0.0020275
R7710 CSoutput.n272 CSoutput.n271 0.0020275
R7711 CSoutput.n269 CSoutput.n207 0.0020275
R7712 CSoutput.n269 CSoutput.n268 0.0020275
R7713 CSoutput.n283 CSoutput.n282 0.0020275
R7714 CSoutput.n282 CSoutput.n281 0.0020275
R7715 CSoutput.n183 CSoutput.n182 0.00166668
R7716 CSoutput.n265 CSoutput.n221 0.00166668
R7717 CSoutput.n149 CSoutput.n148 0.00166668
R7718 CSoutput.n287 CSoutput.n149 0.00133328
R7719 CSoutput.n221 CSoutput.n217 0.00133328
R7720 CSoutput.n277 CSoutput.n183 0.00133328
R7721 CSoutput.n280 CSoutput.n172 0.001
R7722 CSoutput.n258 CSoutput.n172 0.001
R7723 CSoutput.n160 CSoutput.n140 0.001
R7724 CSoutput.n259 CSoutput.n140 0.001
R7725 CSoutput.n161 CSoutput.n141 0.001
R7726 CSoutput.n260 CSoutput.n141 0.001
R7727 CSoutput.n162 CSoutput.n142 0.001
R7728 CSoutput.n261 CSoutput.n142 0.001
R7729 CSoutput.n163 CSoutput.n143 0.001
R7730 CSoutput.n262 CSoutput.n143 0.001
R7731 CSoutput.n256 CSoutput.n208 0.001
R7732 CSoutput.n256 CSoutput.n254 0.001
R7733 CSoutput.n238 CSoutput.n209 0.001
R7734 CSoutput.n232 CSoutput.n209 0.001
R7735 CSoutput.n239 CSoutput.n210 0.001
R7736 CSoutput.n233 CSoutput.n210 0.001
R7737 CSoutput.n240 CSoutput.n211 0.001
R7738 CSoutput.n234 CSoutput.n211 0.001
R7739 CSoutput.n241 CSoutput.n212 0.001
R7740 CSoutput.n235 CSoutput.n212 0.001
R7741 CSoutput.n270 CSoutput.n206 0.001
R7742 CSoutput.n224 CSoutput.n206 0.001
R7743 CSoutput.n194 CSoutput.n174 0.001
R7744 CSoutput.n225 CSoutput.n174 0.001
R7745 CSoutput.n195 CSoutput.n175 0.001
R7746 CSoutput.n226 CSoutput.n175 0.001
R7747 CSoutput.n196 CSoutput.n176 0.001
R7748 CSoutput.n227 CSoutput.n176 0.001
R7749 CSoutput.n197 CSoutput.n177 0.001
R7750 CSoutput.n228 CSoutput.n177 0.001
R7751 CSoutput.n228 CSoutput.n178 0.001
R7752 CSoutput.n227 CSoutput.n179 0.001
R7753 CSoutput.n226 CSoutput.n180 0.001
R7754 CSoutput.n225 CSoutput.t197 0.001
R7755 CSoutput.n224 CSoutput.n181 0.001
R7756 CSoutput.n197 CSoutput.n179 0.001
R7757 CSoutput.n196 CSoutput.n180 0.001
R7758 CSoutput.n195 CSoutput.t197 0.001
R7759 CSoutput.n194 CSoutput.n181 0.001
R7760 CSoutput.n270 CSoutput.n182 0.001
R7761 CSoutput.n235 CSoutput.n213 0.001
R7762 CSoutput.n234 CSoutput.n214 0.001
R7763 CSoutput.n233 CSoutput.n215 0.001
R7764 CSoutput.n232 CSoutput.t193 0.001
R7765 CSoutput.n254 CSoutput.n216 0.001
R7766 CSoutput.n241 CSoutput.n214 0.001
R7767 CSoutput.n240 CSoutput.n215 0.001
R7768 CSoutput.n239 CSoutput.t193 0.001
R7769 CSoutput.n238 CSoutput.n216 0.001
R7770 CSoutput.n265 CSoutput.n208 0.001
R7771 CSoutput.n262 CSoutput.n144 0.001
R7772 CSoutput.n261 CSoutput.n145 0.001
R7773 CSoutput.n260 CSoutput.n146 0.001
R7774 CSoutput.n259 CSoutput.t213 0.001
R7775 CSoutput.n258 CSoutput.n147 0.001
R7776 CSoutput.n163 CSoutput.n145 0.001
R7777 CSoutput.n162 CSoutput.n146 0.001
R7778 CSoutput.n161 CSoutput.t213 0.001
R7779 CSoutput.n160 CSoutput.n147 0.001
R7780 CSoutput.n280 CSoutput.n148 0.001
R7781 commonsourceibias.n25 commonsourceibias.t20 230.006
R7782 commonsourceibias.n91 commonsourceibias.t73 230.006
R7783 commonsourceibias.n218 commonsourceibias.t98 230.006
R7784 commonsourceibias.n154 commonsourceibias.t70 230.006
R7785 commonsourceibias.n322 commonsourceibias.t12 230.006
R7786 commonsourceibias.n281 commonsourceibias.t111 230.006
R7787 commonsourceibias.n483 commonsourceibias.t113 230.006
R7788 commonsourceibias.n419 commonsourceibias.t52 230.006
R7789 commonsourceibias.n70 commonsourceibias.t40 207.983
R7790 commonsourceibias.n136 commonsourceibias.t89 207.983
R7791 commonsourceibias.n263 commonsourceibias.t109 207.983
R7792 commonsourceibias.n199 commonsourceibias.t54 207.983
R7793 commonsourceibias.n368 commonsourceibias.t2 207.983
R7794 commonsourceibias.n402 commonsourceibias.t69 207.983
R7795 commonsourceibias.n529 commonsourceibias.t63 207.983
R7796 commonsourceibias.n465 commonsourceibias.t112 207.983
R7797 commonsourceibias.n10 commonsourceibias.t36 168.701
R7798 commonsourceibias.n63 commonsourceibias.t46 168.701
R7799 commonsourceibias.n57 commonsourceibias.t42 168.701
R7800 commonsourceibias.n16 commonsourceibias.t22 168.701
R7801 commonsourceibias.n49 commonsourceibias.t38 168.701
R7802 commonsourceibias.n43 commonsourceibias.t18 168.701
R7803 commonsourceibias.n19 commonsourceibias.t8 168.701
R7804 commonsourceibias.n21 commonsourceibias.t44 168.701
R7805 commonsourceibias.n23 commonsourceibias.t32 168.701
R7806 commonsourceibias.n26 commonsourceibias.t14 168.701
R7807 commonsourceibias.n1 commonsourceibias.t51 168.701
R7808 commonsourceibias.n129 commonsourceibias.t95 168.701
R7809 commonsourceibias.n123 commonsourceibias.t90 168.701
R7810 commonsourceibias.n7 commonsourceibias.t101 168.701
R7811 commonsourceibias.n115 commonsourceibias.t86 168.701
R7812 commonsourceibias.n109 commonsourceibias.t77 168.701
R7813 commonsourceibias.n85 commonsourceibias.t94 168.701
R7814 commonsourceibias.n87 commonsourceibias.t87 168.701
R7815 commonsourceibias.n89 commonsourceibias.t58 168.701
R7816 commonsourceibias.n92 commonsourceibias.t80 168.701
R7817 commonsourceibias.n219 commonsourceibias.t102 168.701
R7818 commonsourceibias.n216 commonsourceibias.t48 168.701
R7819 commonsourceibias.n214 commonsourceibias.t103 168.701
R7820 commonsourceibias.n212 commonsourceibias.t108 168.701
R7821 commonsourceibias.n236 commonsourceibias.t88 168.701
R7822 commonsourceibias.n242 commonsourceibias.t68 168.701
R7823 commonsourceibias.n209 commonsourceibias.t115 168.701
R7824 commonsourceibias.n250 commonsourceibias.t93 168.701
R7825 commonsourceibias.n256 commonsourceibias.t96 168.701
R7826 commonsourceibias.n203 commonsourceibias.t57 168.701
R7827 commonsourceibias.n139 commonsourceibias.t119 168.701
R7828 commonsourceibias.n192 commonsourceibias.t110 168.701
R7829 commonsourceibias.n186 commonsourceibias.t60 168.701
R7830 commonsourceibias.n145 commonsourceibias.t117 168.701
R7831 commonsourceibias.n178 commonsourceibias.t65 168.701
R7832 commonsourceibias.n172 commonsourceibias.t59 168.701
R7833 commonsourceibias.n148 commonsourceibias.t118 168.701
R7834 commonsourceibias.n150 commonsourceibias.t71 168.701
R7835 commonsourceibias.n152 commonsourceibias.t83 168.701
R7836 commonsourceibias.n155 commonsourceibias.t116 168.701
R7837 commonsourceibias.n323 commonsourceibias.t30 168.701
R7838 commonsourceibias.n320 commonsourceibias.t26 168.701
R7839 commonsourceibias.n318 commonsourceibias.t4 168.701
R7840 commonsourceibias.n316 commonsourceibias.t16 168.701
R7841 commonsourceibias.n340 commonsourceibias.t34 168.701
R7842 commonsourceibias.n346 commonsourceibias.t6 168.701
R7843 commonsourceibias.n348 commonsourceibias.t10 168.701
R7844 commonsourceibias.n355 commonsourceibias.t0 168.701
R7845 commonsourceibias.n361 commonsourceibias.t28 168.701
R7846 commonsourceibias.n308 commonsourceibias.t24 168.701
R7847 commonsourceibias.n267 commonsourceibias.t99 168.701
R7848 commonsourceibias.n395 commonsourceibias.t84 168.701
R7849 commonsourceibias.n389 commonsourceibias.t72 168.701
R7850 commonsourceibias.n382 commonsourceibias.t92 168.701
R7851 commonsourceibias.n380 commonsourceibias.t66 168.701
R7852 commonsourceibias.n282 commonsourceibias.t64 168.701
R7853 commonsourceibias.n279 commonsourceibias.t104 168.701
R7854 commonsourceibias.n277 commonsourceibias.t67 168.701
R7855 commonsourceibias.n275 commonsourceibias.t79 168.701
R7856 commonsourceibias.n299 commonsourceibias.t56 168.701
R7857 commonsourceibias.n484 commonsourceibias.t97 168.701
R7858 commonsourceibias.n481 commonsourceibias.t78 168.701
R7859 commonsourceibias.n479 commonsourceibias.t53 168.701
R7860 commonsourceibias.n477 commonsourceibias.t62 168.701
R7861 commonsourceibias.n501 commonsourceibias.t82 168.701
R7862 commonsourceibias.n507 commonsourceibias.t85 168.701
R7863 commonsourceibias.n509 commonsourceibias.t76 168.701
R7864 commonsourceibias.n516 commonsourceibias.t100 168.701
R7865 commonsourceibias.n522 commonsourceibias.t91 168.701
R7866 commonsourceibias.n469 commonsourceibias.t81 168.701
R7867 commonsourceibias.n420 commonsourceibias.t61 168.701
R7868 commonsourceibias.n417 commonsourceibias.t75 168.701
R7869 commonsourceibias.n415 commonsourceibias.t55 168.701
R7870 commonsourceibias.n413 commonsourceibias.t105 168.701
R7871 commonsourceibias.n437 commonsourceibias.t74 168.701
R7872 commonsourceibias.n443 commonsourceibias.t49 168.701
R7873 commonsourceibias.n445 commonsourceibias.t106 168.701
R7874 commonsourceibias.n452 commonsourceibias.t114 168.701
R7875 commonsourceibias.n458 commonsourceibias.t50 168.701
R7876 commonsourceibias.n405 commonsourceibias.t107 168.701
R7877 commonsourceibias.n27 commonsourceibias.n24 161.3
R7878 commonsourceibias.n29 commonsourceibias.n28 161.3
R7879 commonsourceibias.n31 commonsourceibias.n30 161.3
R7880 commonsourceibias.n32 commonsourceibias.n22 161.3
R7881 commonsourceibias.n34 commonsourceibias.n33 161.3
R7882 commonsourceibias.n36 commonsourceibias.n35 161.3
R7883 commonsourceibias.n37 commonsourceibias.n20 161.3
R7884 commonsourceibias.n39 commonsourceibias.n38 161.3
R7885 commonsourceibias.n41 commonsourceibias.n40 161.3
R7886 commonsourceibias.n42 commonsourceibias.n18 161.3
R7887 commonsourceibias.n45 commonsourceibias.n44 161.3
R7888 commonsourceibias.n46 commonsourceibias.n17 161.3
R7889 commonsourceibias.n48 commonsourceibias.n47 161.3
R7890 commonsourceibias.n50 commonsourceibias.n15 161.3
R7891 commonsourceibias.n52 commonsourceibias.n51 161.3
R7892 commonsourceibias.n53 commonsourceibias.n14 161.3
R7893 commonsourceibias.n55 commonsourceibias.n54 161.3
R7894 commonsourceibias.n56 commonsourceibias.n13 161.3
R7895 commonsourceibias.n59 commonsourceibias.n58 161.3
R7896 commonsourceibias.n60 commonsourceibias.n12 161.3
R7897 commonsourceibias.n62 commonsourceibias.n61 161.3
R7898 commonsourceibias.n64 commonsourceibias.n11 161.3
R7899 commonsourceibias.n66 commonsourceibias.n65 161.3
R7900 commonsourceibias.n68 commonsourceibias.n67 161.3
R7901 commonsourceibias.n69 commonsourceibias.n9 161.3
R7902 commonsourceibias.n93 commonsourceibias.n90 161.3
R7903 commonsourceibias.n95 commonsourceibias.n94 161.3
R7904 commonsourceibias.n97 commonsourceibias.n96 161.3
R7905 commonsourceibias.n98 commonsourceibias.n88 161.3
R7906 commonsourceibias.n100 commonsourceibias.n99 161.3
R7907 commonsourceibias.n102 commonsourceibias.n101 161.3
R7908 commonsourceibias.n103 commonsourceibias.n86 161.3
R7909 commonsourceibias.n105 commonsourceibias.n104 161.3
R7910 commonsourceibias.n107 commonsourceibias.n106 161.3
R7911 commonsourceibias.n108 commonsourceibias.n84 161.3
R7912 commonsourceibias.n111 commonsourceibias.n110 161.3
R7913 commonsourceibias.n112 commonsourceibias.n8 161.3
R7914 commonsourceibias.n114 commonsourceibias.n113 161.3
R7915 commonsourceibias.n116 commonsourceibias.n6 161.3
R7916 commonsourceibias.n118 commonsourceibias.n117 161.3
R7917 commonsourceibias.n119 commonsourceibias.n5 161.3
R7918 commonsourceibias.n121 commonsourceibias.n120 161.3
R7919 commonsourceibias.n122 commonsourceibias.n4 161.3
R7920 commonsourceibias.n125 commonsourceibias.n124 161.3
R7921 commonsourceibias.n126 commonsourceibias.n3 161.3
R7922 commonsourceibias.n128 commonsourceibias.n127 161.3
R7923 commonsourceibias.n130 commonsourceibias.n2 161.3
R7924 commonsourceibias.n132 commonsourceibias.n131 161.3
R7925 commonsourceibias.n134 commonsourceibias.n133 161.3
R7926 commonsourceibias.n135 commonsourceibias.n0 161.3
R7927 commonsourceibias.n262 commonsourceibias.n202 161.3
R7928 commonsourceibias.n261 commonsourceibias.n260 161.3
R7929 commonsourceibias.n259 commonsourceibias.n258 161.3
R7930 commonsourceibias.n257 commonsourceibias.n204 161.3
R7931 commonsourceibias.n255 commonsourceibias.n254 161.3
R7932 commonsourceibias.n253 commonsourceibias.n205 161.3
R7933 commonsourceibias.n252 commonsourceibias.n251 161.3
R7934 commonsourceibias.n249 commonsourceibias.n206 161.3
R7935 commonsourceibias.n248 commonsourceibias.n247 161.3
R7936 commonsourceibias.n246 commonsourceibias.n207 161.3
R7937 commonsourceibias.n245 commonsourceibias.n244 161.3
R7938 commonsourceibias.n243 commonsourceibias.n208 161.3
R7939 commonsourceibias.n241 commonsourceibias.n240 161.3
R7940 commonsourceibias.n239 commonsourceibias.n210 161.3
R7941 commonsourceibias.n238 commonsourceibias.n237 161.3
R7942 commonsourceibias.n235 commonsourceibias.n211 161.3
R7943 commonsourceibias.n234 commonsourceibias.n233 161.3
R7944 commonsourceibias.n232 commonsourceibias.n231 161.3
R7945 commonsourceibias.n230 commonsourceibias.n213 161.3
R7946 commonsourceibias.n229 commonsourceibias.n228 161.3
R7947 commonsourceibias.n227 commonsourceibias.n226 161.3
R7948 commonsourceibias.n225 commonsourceibias.n215 161.3
R7949 commonsourceibias.n224 commonsourceibias.n223 161.3
R7950 commonsourceibias.n222 commonsourceibias.n221 161.3
R7951 commonsourceibias.n220 commonsourceibias.n217 161.3
R7952 commonsourceibias.n156 commonsourceibias.n153 161.3
R7953 commonsourceibias.n158 commonsourceibias.n157 161.3
R7954 commonsourceibias.n160 commonsourceibias.n159 161.3
R7955 commonsourceibias.n161 commonsourceibias.n151 161.3
R7956 commonsourceibias.n163 commonsourceibias.n162 161.3
R7957 commonsourceibias.n165 commonsourceibias.n164 161.3
R7958 commonsourceibias.n166 commonsourceibias.n149 161.3
R7959 commonsourceibias.n168 commonsourceibias.n167 161.3
R7960 commonsourceibias.n170 commonsourceibias.n169 161.3
R7961 commonsourceibias.n171 commonsourceibias.n147 161.3
R7962 commonsourceibias.n174 commonsourceibias.n173 161.3
R7963 commonsourceibias.n175 commonsourceibias.n146 161.3
R7964 commonsourceibias.n177 commonsourceibias.n176 161.3
R7965 commonsourceibias.n179 commonsourceibias.n144 161.3
R7966 commonsourceibias.n181 commonsourceibias.n180 161.3
R7967 commonsourceibias.n182 commonsourceibias.n143 161.3
R7968 commonsourceibias.n184 commonsourceibias.n183 161.3
R7969 commonsourceibias.n185 commonsourceibias.n142 161.3
R7970 commonsourceibias.n188 commonsourceibias.n187 161.3
R7971 commonsourceibias.n189 commonsourceibias.n141 161.3
R7972 commonsourceibias.n191 commonsourceibias.n190 161.3
R7973 commonsourceibias.n193 commonsourceibias.n140 161.3
R7974 commonsourceibias.n195 commonsourceibias.n194 161.3
R7975 commonsourceibias.n197 commonsourceibias.n196 161.3
R7976 commonsourceibias.n198 commonsourceibias.n138 161.3
R7977 commonsourceibias.n367 commonsourceibias.n307 161.3
R7978 commonsourceibias.n366 commonsourceibias.n365 161.3
R7979 commonsourceibias.n364 commonsourceibias.n363 161.3
R7980 commonsourceibias.n362 commonsourceibias.n309 161.3
R7981 commonsourceibias.n360 commonsourceibias.n359 161.3
R7982 commonsourceibias.n358 commonsourceibias.n310 161.3
R7983 commonsourceibias.n357 commonsourceibias.n356 161.3
R7984 commonsourceibias.n354 commonsourceibias.n311 161.3
R7985 commonsourceibias.n353 commonsourceibias.n352 161.3
R7986 commonsourceibias.n351 commonsourceibias.n312 161.3
R7987 commonsourceibias.n350 commonsourceibias.n349 161.3
R7988 commonsourceibias.n347 commonsourceibias.n313 161.3
R7989 commonsourceibias.n345 commonsourceibias.n344 161.3
R7990 commonsourceibias.n343 commonsourceibias.n314 161.3
R7991 commonsourceibias.n342 commonsourceibias.n341 161.3
R7992 commonsourceibias.n339 commonsourceibias.n315 161.3
R7993 commonsourceibias.n338 commonsourceibias.n337 161.3
R7994 commonsourceibias.n336 commonsourceibias.n335 161.3
R7995 commonsourceibias.n334 commonsourceibias.n317 161.3
R7996 commonsourceibias.n333 commonsourceibias.n332 161.3
R7997 commonsourceibias.n331 commonsourceibias.n330 161.3
R7998 commonsourceibias.n329 commonsourceibias.n319 161.3
R7999 commonsourceibias.n328 commonsourceibias.n327 161.3
R8000 commonsourceibias.n326 commonsourceibias.n325 161.3
R8001 commonsourceibias.n324 commonsourceibias.n321 161.3
R8002 commonsourceibias.n301 commonsourceibias.n300 161.3
R8003 commonsourceibias.n298 commonsourceibias.n274 161.3
R8004 commonsourceibias.n297 commonsourceibias.n296 161.3
R8005 commonsourceibias.n295 commonsourceibias.n294 161.3
R8006 commonsourceibias.n293 commonsourceibias.n276 161.3
R8007 commonsourceibias.n292 commonsourceibias.n291 161.3
R8008 commonsourceibias.n290 commonsourceibias.n289 161.3
R8009 commonsourceibias.n288 commonsourceibias.n278 161.3
R8010 commonsourceibias.n287 commonsourceibias.n286 161.3
R8011 commonsourceibias.n285 commonsourceibias.n284 161.3
R8012 commonsourceibias.n283 commonsourceibias.n280 161.3
R8013 commonsourceibias.n377 commonsourceibias.n273 161.3
R8014 commonsourceibias.n401 commonsourceibias.n266 161.3
R8015 commonsourceibias.n400 commonsourceibias.n399 161.3
R8016 commonsourceibias.n398 commonsourceibias.n397 161.3
R8017 commonsourceibias.n396 commonsourceibias.n268 161.3
R8018 commonsourceibias.n394 commonsourceibias.n393 161.3
R8019 commonsourceibias.n392 commonsourceibias.n269 161.3
R8020 commonsourceibias.n391 commonsourceibias.n390 161.3
R8021 commonsourceibias.n388 commonsourceibias.n270 161.3
R8022 commonsourceibias.n387 commonsourceibias.n386 161.3
R8023 commonsourceibias.n385 commonsourceibias.n271 161.3
R8024 commonsourceibias.n384 commonsourceibias.n383 161.3
R8025 commonsourceibias.n381 commonsourceibias.n272 161.3
R8026 commonsourceibias.n379 commonsourceibias.n378 161.3
R8027 commonsourceibias.n528 commonsourceibias.n468 161.3
R8028 commonsourceibias.n527 commonsourceibias.n526 161.3
R8029 commonsourceibias.n525 commonsourceibias.n524 161.3
R8030 commonsourceibias.n523 commonsourceibias.n470 161.3
R8031 commonsourceibias.n521 commonsourceibias.n520 161.3
R8032 commonsourceibias.n519 commonsourceibias.n471 161.3
R8033 commonsourceibias.n518 commonsourceibias.n517 161.3
R8034 commonsourceibias.n515 commonsourceibias.n472 161.3
R8035 commonsourceibias.n514 commonsourceibias.n513 161.3
R8036 commonsourceibias.n512 commonsourceibias.n473 161.3
R8037 commonsourceibias.n511 commonsourceibias.n510 161.3
R8038 commonsourceibias.n508 commonsourceibias.n474 161.3
R8039 commonsourceibias.n506 commonsourceibias.n505 161.3
R8040 commonsourceibias.n504 commonsourceibias.n475 161.3
R8041 commonsourceibias.n503 commonsourceibias.n502 161.3
R8042 commonsourceibias.n500 commonsourceibias.n476 161.3
R8043 commonsourceibias.n499 commonsourceibias.n498 161.3
R8044 commonsourceibias.n497 commonsourceibias.n496 161.3
R8045 commonsourceibias.n495 commonsourceibias.n478 161.3
R8046 commonsourceibias.n494 commonsourceibias.n493 161.3
R8047 commonsourceibias.n492 commonsourceibias.n491 161.3
R8048 commonsourceibias.n490 commonsourceibias.n480 161.3
R8049 commonsourceibias.n489 commonsourceibias.n488 161.3
R8050 commonsourceibias.n487 commonsourceibias.n486 161.3
R8051 commonsourceibias.n485 commonsourceibias.n482 161.3
R8052 commonsourceibias.n464 commonsourceibias.n404 161.3
R8053 commonsourceibias.n463 commonsourceibias.n462 161.3
R8054 commonsourceibias.n461 commonsourceibias.n460 161.3
R8055 commonsourceibias.n459 commonsourceibias.n406 161.3
R8056 commonsourceibias.n457 commonsourceibias.n456 161.3
R8057 commonsourceibias.n455 commonsourceibias.n407 161.3
R8058 commonsourceibias.n454 commonsourceibias.n453 161.3
R8059 commonsourceibias.n451 commonsourceibias.n408 161.3
R8060 commonsourceibias.n450 commonsourceibias.n449 161.3
R8061 commonsourceibias.n448 commonsourceibias.n409 161.3
R8062 commonsourceibias.n447 commonsourceibias.n446 161.3
R8063 commonsourceibias.n444 commonsourceibias.n410 161.3
R8064 commonsourceibias.n442 commonsourceibias.n441 161.3
R8065 commonsourceibias.n440 commonsourceibias.n411 161.3
R8066 commonsourceibias.n439 commonsourceibias.n438 161.3
R8067 commonsourceibias.n436 commonsourceibias.n412 161.3
R8068 commonsourceibias.n435 commonsourceibias.n434 161.3
R8069 commonsourceibias.n433 commonsourceibias.n432 161.3
R8070 commonsourceibias.n431 commonsourceibias.n414 161.3
R8071 commonsourceibias.n430 commonsourceibias.n429 161.3
R8072 commonsourceibias.n428 commonsourceibias.n427 161.3
R8073 commonsourceibias.n426 commonsourceibias.n416 161.3
R8074 commonsourceibias.n425 commonsourceibias.n424 161.3
R8075 commonsourceibias.n423 commonsourceibias.n422 161.3
R8076 commonsourceibias.n421 commonsourceibias.n418 161.3
R8077 commonsourceibias.n80 commonsourceibias.n78 81.5057
R8078 commonsourceibias.n304 commonsourceibias.n302 81.5057
R8079 commonsourceibias.n80 commonsourceibias.n79 80.9324
R8080 commonsourceibias.n82 commonsourceibias.n81 80.9324
R8081 commonsourceibias.n77 commonsourceibias.n76 80.9324
R8082 commonsourceibias.n75 commonsourceibias.n74 80.9324
R8083 commonsourceibias.n73 commonsourceibias.n72 80.9324
R8084 commonsourceibias.n371 commonsourceibias.n370 80.9324
R8085 commonsourceibias.n373 commonsourceibias.n372 80.9324
R8086 commonsourceibias.n375 commonsourceibias.n374 80.9324
R8087 commonsourceibias.n306 commonsourceibias.n305 80.9324
R8088 commonsourceibias.n304 commonsourceibias.n303 80.9324
R8089 commonsourceibias.n71 commonsourceibias.n70 80.6037
R8090 commonsourceibias.n137 commonsourceibias.n136 80.6037
R8091 commonsourceibias.n264 commonsourceibias.n263 80.6037
R8092 commonsourceibias.n200 commonsourceibias.n199 80.6037
R8093 commonsourceibias.n369 commonsourceibias.n368 80.6037
R8094 commonsourceibias.n403 commonsourceibias.n402 80.6037
R8095 commonsourceibias.n530 commonsourceibias.n529 80.6037
R8096 commonsourceibias.n466 commonsourceibias.n465 80.6037
R8097 commonsourceibias.n65 commonsourceibias.n64 56.5617
R8098 commonsourceibias.n51 commonsourceibias.n50 56.5617
R8099 commonsourceibias.n42 commonsourceibias.n41 56.5617
R8100 commonsourceibias.n28 commonsourceibias.n27 56.5617
R8101 commonsourceibias.n131 commonsourceibias.n130 56.5617
R8102 commonsourceibias.n117 commonsourceibias.n116 56.5617
R8103 commonsourceibias.n108 commonsourceibias.n107 56.5617
R8104 commonsourceibias.n94 commonsourceibias.n93 56.5617
R8105 commonsourceibias.n221 commonsourceibias.n220 56.5617
R8106 commonsourceibias.n235 commonsourceibias.n234 56.5617
R8107 commonsourceibias.n244 commonsourceibias.n243 56.5617
R8108 commonsourceibias.n258 commonsourceibias.n257 56.5617
R8109 commonsourceibias.n194 commonsourceibias.n193 56.5617
R8110 commonsourceibias.n180 commonsourceibias.n179 56.5617
R8111 commonsourceibias.n171 commonsourceibias.n170 56.5617
R8112 commonsourceibias.n157 commonsourceibias.n156 56.5617
R8113 commonsourceibias.n325 commonsourceibias.n324 56.5617
R8114 commonsourceibias.n339 commonsourceibias.n338 56.5617
R8115 commonsourceibias.n349 commonsourceibias.n347 56.5617
R8116 commonsourceibias.n363 commonsourceibias.n362 56.5617
R8117 commonsourceibias.n397 commonsourceibias.n396 56.5617
R8118 commonsourceibias.n383 commonsourceibias.n381 56.5617
R8119 commonsourceibias.n284 commonsourceibias.n283 56.5617
R8120 commonsourceibias.n298 commonsourceibias.n297 56.5617
R8121 commonsourceibias.n486 commonsourceibias.n485 56.5617
R8122 commonsourceibias.n500 commonsourceibias.n499 56.5617
R8123 commonsourceibias.n510 commonsourceibias.n508 56.5617
R8124 commonsourceibias.n524 commonsourceibias.n523 56.5617
R8125 commonsourceibias.n422 commonsourceibias.n421 56.5617
R8126 commonsourceibias.n436 commonsourceibias.n435 56.5617
R8127 commonsourceibias.n446 commonsourceibias.n444 56.5617
R8128 commonsourceibias.n460 commonsourceibias.n459 56.5617
R8129 commonsourceibias.n56 commonsourceibias.n55 56.0773
R8130 commonsourceibias.n37 commonsourceibias.n36 56.0773
R8131 commonsourceibias.n122 commonsourceibias.n121 56.0773
R8132 commonsourceibias.n103 commonsourceibias.n102 56.0773
R8133 commonsourceibias.n230 commonsourceibias.n229 56.0773
R8134 commonsourceibias.n249 commonsourceibias.n248 56.0773
R8135 commonsourceibias.n185 commonsourceibias.n184 56.0773
R8136 commonsourceibias.n166 commonsourceibias.n165 56.0773
R8137 commonsourceibias.n334 commonsourceibias.n333 56.0773
R8138 commonsourceibias.n354 commonsourceibias.n353 56.0773
R8139 commonsourceibias.n388 commonsourceibias.n387 56.0773
R8140 commonsourceibias.n293 commonsourceibias.n292 56.0773
R8141 commonsourceibias.n495 commonsourceibias.n494 56.0773
R8142 commonsourceibias.n515 commonsourceibias.n514 56.0773
R8143 commonsourceibias.n431 commonsourceibias.n430 56.0773
R8144 commonsourceibias.n451 commonsourceibias.n450 56.0773
R8145 commonsourceibias.n70 commonsourceibias.n69 46.0096
R8146 commonsourceibias.n136 commonsourceibias.n135 46.0096
R8147 commonsourceibias.n263 commonsourceibias.n262 46.0096
R8148 commonsourceibias.n199 commonsourceibias.n198 46.0096
R8149 commonsourceibias.n368 commonsourceibias.n367 46.0096
R8150 commonsourceibias.n402 commonsourceibias.n401 46.0096
R8151 commonsourceibias.n529 commonsourceibias.n528 46.0096
R8152 commonsourceibias.n465 commonsourceibias.n464 46.0096
R8153 commonsourceibias.n58 commonsourceibias.n12 41.5458
R8154 commonsourceibias.n33 commonsourceibias.n32 41.5458
R8155 commonsourceibias.n124 commonsourceibias.n3 41.5458
R8156 commonsourceibias.n99 commonsourceibias.n98 41.5458
R8157 commonsourceibias.n226 commonsourceibias.n225 41.5458
R8158 commonsourceibias.n251 commonsourceibias.n205 41.5458
R8159 commonsourceibias.n187 commonsourceibias.n141 41.5458
R8160 commonsourceibias.n162 commonsourceibias.n161 41.5458
R8161 commonsourceibias.n330 commonsourceibias.n329 41.5458
R8162 commonsourceibias.n356 commonsourceibias.n310 41.5458
R8163 commonsourceibias.n390 commonsourceibias.n269 41.5458
R8164 commonsourceibias.n289 commonsourceibias.n288 41.5458
R8165 commonsourceibias.n491 commonsourceibias.n490 41.5458
R8166 commonsourceibias.n517 commonsourceibias.n471 41.5458
R8167 commonsourceibias.n427 commonsourceibias.n426 41.5458
R8168 commonsourceibias.n453 commonsourceibias.n407 41.5458
R8169 commonsourceibias.n48 commonsourceibias.n17 40.577
R8170 commonsourceibias.n44 commonsourceibias.n17 40.577
R8171 commonsourceibias.n114 commonsourceibias.n8 40.577
R8172 commonsourceibias.n110 commonsourceibias.n8 40.577
R8173 commonsourceibias.n237 commonsourceibias.n210 40.577
R8174 commonsourceibias.n241 commonsourceibias.n210 40.577
R8175 commonsourceibias.n177 commonsourceibias.n146 40.577
R8176 commonsourceibias.n173 commonsourceibias.n146 40.577
R8177 commonsourceibias.n341 commonsourceibias.n314 40.577
R8178 commonsourceibias.n345 commonsourceibias.n314 40.577
R8179 commonsourceibias.n379 commonsourceibias.n273 40.577
R8180 commonsourceibias.n300 commonsourceibias.n273 40.577
R8181 commonsourceibias.n502 commonsourceibias.n475 40.577
R8182 commonsourceibias.n506 commonsourceibias.n475 40.577
R8183 commonsourceibias.n438 commonsourceibias.n411 40.577
R8184 commonsourceibias.n442 commonsourceibias.n411 40.577
R8185 commonsourceibias.n62 commonsourceibias.n12 39.6083
R8186 commonsourceibias.n32 commonsourceibias.n31 39.6083
R8187 commonsourceibias.n128 commonsourceibias.n3 39.6083
R8188 commonsourceibias.n98 commonsourceibias.n97 39.6083
R8189 commonsourceibias.n225 commonsourceibias.n224 39.6083
R8190 commonsourceibias.n255 commonsourceibias.n205 39.6083
R8191 commonsourceibias.n191 commonsourceibias.n141 39.6083
R8192 commonsourceibias.n161 commonsourceibias.n160 39.6083
R8193 commonsourceibias.n329 commonsourceibias.n328 39.6083
R8194 commonsourceibias.n360 commonsourceibias.n310 39.6083
R8195 commonsourceibias.n394 commonsourceibias.n269 39.6083
R8196 commonsourceibias.n288 commonsourceibias.n287 39.6083
R8197 commonsourceibias.n490 commonsourceibias.n489 39.6083
R8198 commonsourceibias.n521 commonsourceibias.n471 39.6083
R8199 commonsourceibias.n426 commonsourceibias.n425 39.6083
R8200 commonsourceibias.n457 commonsourceibias.n407 39.6083
R8201 commonsourceibias.n26 commonsourceibias.n25 33.0515
R8202 commonsourceibias.n92 commonsourceibias.n91 33.0515
R8203 commonsourceibias.n155 commonsourceibias.n154 33.0515
R8204 commonsourceibias.n219 commonsourceibias.n218 33.0515
R8205 commonsourceibias.n323 commonsourceibias.n322 33.0515
R8206 commonsourceibias.n282 commonsourceibias.n281 33.0515
R8207 commonsourceibias.n484 commonsourceibias.n483 33.0515
R8208 commonsourceibias.n420 commonsourceibias.n419 33.0515
R8209 commonsourceibias.n25 commonsourceibias.n24 28.5514
R8210 commonsourceibias.n91 commonsourceibias.n90 28.5514
R8211 commonsourceibias.n218 commonsourceibias.n217 28.5514
R8212 commonsourceibias.n154 commonsourceibias.n153 28.5514
R8213 commonsourceibias.n322 commonsourceibias.n321 28.5514
R8214 commonsourceibias.n281 commonsourceibias.n280 28.5514
R8215 commonsourceibias.n483 commonsourceibias.n482 28.5514
R8216 commonsourceibias.n419 commonsourceibias.n418 28.5514
R8217 commonsourceibias.n69 commonsourceibias.n68 26.0455
R8218 commonsourceibias.n135 commonsourceibias.n134 26.0455
R8219 commonsourceibias.n262 commonsourceibias.n261 26.0455
R8220 commonsourceibias.n198 commonsourceibias.n197 26.0455
R8221 commonsourceibias.n367 commonsourceibias.n366 26.0455
R8222 commonsourceibias.n401 commonsourceibias.n400 26.0455
R8223 commonsourceibias.n528 commonsourceibias.n527 26.0455
R8224 commonsourceibias.n464 commonsourceibias.n463 26.0455
R8225 commonsourceibias.n55 commonsourceibias.n14 25.0767
R8226 commonsourceibias.n38 commonsourceibias.n37 25.0767
R8227 commonsourceibias.n121 commonsourceibias.n5 25.0767
R8228 commonsourceibias.n104 commonsourceibias.n103 25.0767
R8229 commonsourceibias.n231 commonsourceibias.n230 25.0767
R8230 commonsourceibias.n248 commonsourceibias.n207 25.0767
R8231 commonsourceibias.n184 commonsourceibias.n143 25.0767
R8232 commonsourceibias.n167 commonsourceibias.n166 25.0767
R8233 commonsourceibias.n335 commonsourceibias.n334 25.0767
R8234 commonsourceibias.n353 commonsourceibias.n312 25.0767
R8235 commonsourceibias.n387 commonsourceibias.n271 25.0767
R8236 commonsourceibias.n294 commonsourceibias.n293 25.0767
R8237 commonsourceibias.n496 commonsourceibias.n495 25.0767
R8238 commonsourceibias.n514 commonsourceibias.n473 25.0767
R8239 commonsourceibias.n432 commonsourceibias.n431 25.0767
R8240 commonsourceibias.n450 commonsourceibias.n409 25.0767
R8241 commonsourceibias.n51 commonsourceibias.n16 24.3464
R8242 commonsourceibias.n41 commonsourceibias.n19 24.3464
R8243 commonsourceibias.n117 commonsourceibias.n7 24.3464
R8244 commonsourceibias.n107 commonsourceibias.n85 24.3464
R8245 commonsourceibias.n234 commonsourceibias.n212 24.3464
R8246 commonsourceibias.n244 commonsourceibias.n209 24.3464
R8247 commonsourceibias.n180 commonsourceibias.n145 24.3464
R8248 commonsourceibias.n170 commonsourceibias.n148 24.3464
R8249 commonsourceibias.n338 commonsourceibias.n316 24.3464
R8250 commonsourceibias.n349 commonsourceibias.n348 24.3464
R8251 commonsourceibias.n383 commonsourceibias.n382 24.3464
R8252 commonsourceibias.n297 commonsourceibias.n275 24.3464
R8253 commonsourceibias.n499 commonsourceibias.n477 24.3464
R8254 commonsourceibias.n510 commonsourceibias.n509 24.3464
R8255 commonsourceibias.n435 commonsourceibias.n413 24.3464
R8256 commonsourceibias.n446 commonsourceibias.n445 24.3464
R8257 commonsourceibias.n65 commonsourceibias.n10 23.8546
R8258 commonsourceibias.n27 commonsourceibias.n26 23.8546
R8259 commonsourceibias.n131 commonsourceibias.n1 23.8546
R8260 commonsourceibias.n93 commonsourceibias.n92 23.8546
R8261 commonsourceibias.n220 commonsourceibias.n219 23.8546
R8262 commonsourceibias.n258 commonsourceibias.n203 23.8546
R8263 commonsourceibias.n194 commonsourceibias.n139 23.8546
R8264 commonsourceibias.n156 commonsourceibias.n155 23.8546
R8265 commonsourceibias.n324 commonsourceibias.n323 23.8546
R8266 commonsourceibias.n363 commonsourceibias.n308 23.8546
R8267 commonsourceibias.n397 commonsourceibias.n267 23.8546
R8268 commonsourceibias.n283 commonsourceibias.n282 23.8546
R8269 commonsourceibias.n485 commonsourceibias.n484 23.8546
R8270 commonsourceibias.n524 commonsourceibias.n469 23.8546
R8271 commonsourceibias.n421 commonsourceibias.n420 23.8546
R8272 commonsourceibias.n460 commonsourceibias.n405 23.8546
R8273 commonsourceibias.n64 commonsourceibias.n63 16.9689
R8274 commonsourceibias.n28 commonsourceibias.n23 16.9689
R8275 commonsourceibias.n130 commonsourceibias.n129 16.9689
R8276 commonsourceibias.n94 commonsourceibias.n89 16.9689
R8277 commonsourceibias.n221 commonsourceibias.n216 16.9689
R8278 commonsourceibias.n257 commonsourceibias.n256 16.9689
R8279 commonsourceibias.n193 commonsourceibias.n192 16.9689
R8280 commonsourceibias.n157 commonsourceibias.n152 16.9689
R8281 commonsourceibias.n325 commonsourceibias.n320 16.9689
R8282 commonsourceibias.n362 commonsourceibias.n361 16.9689
R8283 commonsourceibias.n396 commonsourceibias.n395 16.9689
R8284 commonsourceibias.n284 commonsourceibias.n279 16.9689
R8285 commonsourceibias.n486 commonsourceibias.n481 16.9689
R8286 commonsourceibias.n523 commonsourceibias.n522 16.9689
R8287 commonsourceibias.n422 commonsourceibias.n417 16.9689
R8288 commonsourceibias.n459 commonsourceibias.n458 16.9689
R8289 commonsourceibias.n50 commonsourceibias.n49 16.477
R8290 commonsourceibias.n43 commonsourceibias.n42 16.477
R8291 commonsourceibias.n116 commonsourceibias.n115 16.477
R8292 commonsourceibias.n109 commonsourceibias.n108 16.477
R8293 commonsourceibias.n236 commonsourceibias.n235 16.477
R8294 commonsourceibias.n243 commonsourceibias.n242 16.477
R8295 commonsourceibias.n179 commonsourceibias.n178 16.477
R8296 commonsourceibias.n172 commonsourceibias.n171 16.477
R8297 commonsourceibias.n340 commonsourceibias.n339 16.477
R8298 commonsourceibias.n347 commonsourceibias.n346 16.477
R8299 commonsourceibias.n381 commonsourceibias.n380 16.477
R8300 commonsourceibias.n299 commonsourceibias.n298 16.477
R8301 commonsourceibias.n501 commonsourceibias.n500 16.477
R8302 commonsourceibias.n508 commonsourceibias.n507 16.477
R8303 commonsourceibias.n437 commonsourceibias.n436 16.477
R8304 commonsourceibias.n444 commonsourceibias.n443 16.477
R8305 commonsourceibias.n57 commonsourceibias.n56 15.9852
R8306 commonsourceibias.n36 commonsourceibias.n21 15.9852
R8307 commonsourceibias.n123 commonsourceibias.n122 15.9852
R8308 commonsourceibias.n102 commonsourceibias.n87 15.9852
R8309 commonsourceibias.n229 commonsourceibias.n214 15.9852
R8310 commonsourceibias.n250 commonsourceibias.n249 15.9852
R8311 commonsourceibias.n186 commonsourceibias.n185 15.9852
R8312 commonsourceibias.n165 commonsourceibias.n150 15.9852
R8313 commonsourceibias.n333 commonsourceibias.n318 15.9852
R8314 commonsourceibias.n355 commonsourceibias.n354 15.9852
R8315 commonsourceibias.n389 commonsourceibias.n388 15.9852
R8316 commonsourceibias.n292 commonsourceibias.n277 15.9852
R8317 commonsourceibias.n494 commonsourceibias.n479 15.9852
R8318 commonsourceibias.n516 commonsourceibias.n515 15.9852
R8319 commonsourceibias.n430 commonsourceibias.n415 15.9852
R8320 commonsourceibias.n452 commonsourceibias.n451 15.9852
R8321 commonsourceibias.n73 commonsourceibias.n71 13.2057
R8322 commonsourceibias.n371 commonsourceibias.n369 13.2057
R8323 commonsourceibias.n532 commonsourceibias.n265 10.122
R8324 commonsourceibias.n112 commonsourceibias.n83 9.50363
R8325 commonsourceibias.n377 commonsourceibias.n376 9.50363
R8326 commonsourceibias.n201 commonsourceibias.n137 8.7339
R8327 commonsourceibias.n467 commonsourceibias.n403 8.7339
R8328 commonsourceibias.n58 commonsourceibias.n57 8.60764
R8329 commonsourceibias.n33 commonsourceibias.n21 8.60764
R8330 commonsourceibias.n124 commonsourceibias.n123 8.60764
R8331 commonsourceibias.n99 commonsourceibias.n87 8.60764
R8332 commonsourceibias.n226 commonsourceibias.n214 8.60764
R8333 commonsourceibias.n251 commonsourceibias.n250 8.60764
R8334 commonsourceibias.n187 commonsourceibias.n186 8.60764
R8335 commonsourceibias.n162 commonsourceibias.n150 8.60764
R8336 commonsourceibias.n330 commonsourceibias.n318 8.60764
R8337 commonsourceibias.n356 commonsourceibias.n355 8.60764
R8338 commonsourceibias.n390 commonsourceibias.n389 8.60764
R8339 commonsourceibias.n289 commonsourceibias.n277 8.60764
R8340 commonsourceibias.n491 commonsourceibias.n479 8.60764
R8341 commonsourceibias.n517 commonsourceibias.n516 8.60764
R8342 commonsourceibias.n427 commonsourceibias.n415 8.60764
R8343 commonsourceibias.n453 commonsourceibias.n452 8.60764
R8344 commonsourceibias.n532 commonsourceibias.n531 8.46921
R8345 commonsourceibias.n49 commonsourceibias.n48 8.11581
R8346 commonsourceibias.n44 commonsourceibias.n43 8.11581
R8347 commonsourceibias.n115 commonsourceibias.n114 8.11581
R8348 commonsourceibias.n110 commonsourceibias.n109 8.11581
R8349 commonsourceibias.n237 commonsourceibias.n236 8.11581
R8350 commonsourceibias.n242 commonsourceibias.n241 8.11581
R8351 commonsourceibias.n178 commonsourceibias.n177 8.11581
R8352 commonsourceibias.n173 commonsourceibias.n172 8.11581
R8353 commonsourceibias.n341 commonsourceibias.n340 8.11581
R8354 commonsourceibias.n346 commonsourceibias.n345 8.11581
R8355 commonsourceibias.n380 commonsourceibias.n379 8.11581
R8356 commonsourceibias.n300 commonsourceibias.n299 8.11581
R8357 commonsourceibias.n502 commonsourceibias.n501 8.11581
R8358 commonsourceibias.n507 commonsourceibias.n506 8.11581
R8359 commonsourceibias.n438 commonsourceibias.n437 8.11581
R8360 commonsourceibias.n443 commonsourceibias.n442 8.11581
R8361 commonsourceibias.n63 commonsourceibias.n62 7.62397
R8362 commonsourceibias.n31 commonsourceibias.n23 7.62397
R8363 commonsourceibias.n129 commonsourceibias.n128 7.62397
R8364 commonsourceibias.n97 commonsourceibias.n89 7.62397
R8365 commonsourceibias.n224 commonsourceibias.n216 7.62397
R8366 commonsourceibias.n256 commonsourceibias.n255 7.62397
R8367 commonsourceibias.n192 commonsourceibias.n191 7.62397
R8368 commonsourceibias.n160 commonsourceibias.n152 7.62397
R8369 commonsourceibias.n328 commonsourceibias.n320 7.62397
R8370 commonsourceibias.n361 commonsourceibias.n360 7.62397
R8371 commonsourceibias.n395 commonsourceibias.n394 7.62397
R8372 commonsourceibias.n287 commonsourceibias.n279 7.62397
R8373 commonsourceibias.n489 commonsourceibias.n481 7.62397
R8374 commonsourceibias.n522 commonsourceibias.n521 7.62397
R8375 commonsourceibias.n425 commonsourceibias.n417 7.62397
R8376 commonsourceibias.n458 commonsourceibias.n457 7.62397
R8377 commonsourceibias.n265 commonsourceibias.n264 5.00473
R8378 commonsourceibias.n201 commonsourceibias.n200 5.00473
R8379 commonsourceibias.n531 commonsourceibias.n530 5.00473
R8380 commonsourceibias.n467 commonsourceibias.n466 5.00473
R8381 commonsourceibias commonsourceibias.n532 3.87639
R8382 commonsourceibias.n265 commonsourceibias.n201 3.72967
R8383 commonsourceibias.n531 commonsourceibias.n467 3.72967
R8384 commonsourceibias.n78 commonsourceibias.t15 2.82907
R8385 commonsourceibias.n78 commonsourceibias.t21 2.82907
R8386 commonsourceibias.n79 commonsourceibias.t45 2.82907
R8387 commonsourceibias.n79 commonsourceibias.t33 2.82907
R8388 commonsourceibias.n81 commonsourceibias.t19 2.82907
R8389 commonsourceibias.n81 commonsourceibias.t9 2.82907
R8390 commonsourceibias.n76 commonsourceibias.t23 2.82907
R8391 commonsourceibias.n76 commonsourceibias.t39 2.82907
R8392 commonsourceibias.n74 commonsourceibias.t47 2.82907
R8393 commonsourceibias.n74 commonsourceibias.t43 2.82907
R8394 commonsourceibias.n72 commonsourceibias.t41 2.82907
R8395 commonsourceibias.n72 commonsourceibias.t37 2.82907
R8396 commonsourceibias.n370 commonsourceibias.t25 2.82907
R8397 commonsourceibias.n370 commonsourceibias.t3 2.82907
R8398 commonsourceibias.n372 commonsourceibias.t1 2.82907
R8399 commonsourceibias.n372 commonsourceibias.t29 2.82907
R8400 commonsourceibias.n374 commonsourceibias.t7 2.82907
R8401 commonsourceibias.n374 commonsourceibias.t11 2.82907
R8402 commonsourceibias.n305 commonsourceibias.t17 2.82907
R8403 commonsourceibias.n305 commonsourceibias.t35 2.82907
R8404 commonsourceibias.n303 commonsourceibias.t27 2.82907
R8405 commonsourceibias.n303 commonsourceibias.t5 2.82907
R8406 commonsourceibias.n302 commonsourceibias.t13 2.82907
R8407 commonsourceibias.n302 commonsourceibias.t31 2.82907
R8408 commonsourceibias.n68 commonsourceibias.n10 0.738255
R8409 commonsourceibias.n134 commonsourceibias.n1 0.738255
R8410 commonsourceibias.n261 commonsourceibias.n203 0.738255
R8411 commonsourceibias.n197 commonsourceibias.n139 0.738255
R8412 commonsourceibias.n366 commonsourceibias.n308 0.738255
R8413 commonsourceibias.n400 commonsourceibias.n267 0.738255
R8414 commonsourceibias.n527 commonsourceibias.n469 0.738255
R8415 commonsourceibias.n463 commonsourceibias.n405 0.738255
R8416 commonsourceibias.n75 commonsourceibias.n73 0.573776
R8417 commonsourceibias.n77 commonsourceibias.n75 0.573776
R8418 commonsourceibias.n82 commonsourceibias.n80 0.573776
R8419 commonsourceibias.n306 commonsourceibias.n304 0.573776
R8420 commonsourceibias.n375 commonsourceibias.n373 0.573776
R8421 commonsourceibias.n373 commonsourceibias.n371 0.573776
R8422 commonsourceibias.n83 commonsourceibias.n77 0.287138
R8423 commonsourceibias.n83 commonsourceibias.n82 0.287138
R8424 commonsourceibias.n376 commonsourceibias.n306 0.287138
R8425 commonsourceibias.n376 commonsourceibias.n375 0.287138
R8426 commonsourceibias.n71 commonsourceibias.n9 0.285035
R8427 commonsourceibias.n137 commonsourceibias.n0 0.285035
R8428 commonsourceibias.n264 commonsourceibias.n202 0.285035
R8429 commonsourceibias.n200 commonsourceibias.n138 0.285035
R8430 commonsourceibias.n369 commonsourceibias.n307 0.285035
R8431 commonsourceibias.n403 commonsourceibias.n266 0.285035
R8432 commonsourceibias.n530 commonsourceibias.n468 0.285035
R8433 commonsourceibias.n466 commonsourceibias.n404 0.285035
R8434 commonsourceibias.n16 commonsourceibias.n14 0.246418
R8435 commonsourceibias.n38 commonsourceibias.n19 0.246418
R8436 commonsourceibias.n7 commonsourceibias.n5 0.246418
R8437 commonsourceibias.n104 commonsourceibias.n85 0.246418
R8438 commonsourceibias.n231 commonsourceibias.n212 0.246418
R8439 commonsourceibias.n209 commonsourceibias.n207 0.246418
R8440 commonsourceibias.n145 commonsourceibias.n143 0.246418
R8441 commonsourceibias.n167 commonsourceibias.n148 0.246418
R8442 commonsourceibias.n335 commonsourceibias.n316 0.246418
R8443 commonsourceibias.n348 commonsourceibias.n312 0.246418
R8444 commonsourceibias.n382 commonsourceibias.n271 0.246418
R8445 commonsourceibias.n294 commonsourceibias.n275 0.246418
R8446 commonsourceibias.n496 commonsourceibias.n477 0.246418
R8447 commonsourceibias.n509 commonsourceibias.n473 0.246418
R8448 commonsourceibias.n432 commonsourceibias.n413 0.246418
R8449 commonsourceibias.n445 commonsourceibias.n409 0.246418
R8450 commonsourceibias.n67 commonsourceibias.n9 0.189894
R8451 commonsourceibias.n67 commonsourceibias.n66 0.189894
R8452 commonsourceibias.n66 commonsourceibias.n11 0.189894
R8453 commonsourceibias.n61 commonsourceibias.n11 0.189894
R8454 commonsourceibias.n61 commonsourceibias.n60 0.189894
R8455 commonsourceibias.n60 commonsourceibias.n59 0.189894
R8456 commonsourceibias.n59 commonsourceibias.n13 0.189894
R8457 commonsourceibias.n54 commonsourceibias.n13 0.189894
R8458 commonsourceibias.n54 commonsourceibias.n53 0.189894
R8459 commonsourceibias.n53 commonsourceibias.n52 0.189894
R8460 commonsourceibias.n52 commonsourceibias.n15 0.189894
R8461 commonsourceibias.n47 commonsourceibias.n15 0.189894
R8462 commonsourceibias.n47 commonsourceibias.n46 0.189894
R8463 commonsourceibias.n46 commonsourceibias.n45 0.189894
R8464 commonsourceibias.n45 commonsourceibias.n18 0.189894
R8465 commonsourceibias.n40 commonsourceibias.n18 0.189894
R8466 commonsourceibias.n40 commonsourceibias.n39 0.189894
R8467 commonsourceibias.n39 commonsourceibias.n20 0.189894
R8468 commonsourceibias.n35 commonsourceibias.n20 0.189894
R8469 commonsourceibias.n35 commonsourceibias.n34 0.189894
R8470 commonsourceibias.n34 commonsourceibias.n22 0.189894
R8471 commonsourceibias.n30 commonsourceibias.n22 0.189894
R8472 commonsourceibias.n30 commonsourceibias.n29 0.189894
R8473 commonsourceibias.n29 commonsourceibias.n24 0.189894
R8474 commonsourceibias.n111 commonsourceibias.n84 0.189894
R8475 commonsourceibias.n106 commonsourceibias.n84 0.189894
R8476 commonsourceibias.n106 commonsourceibias.n105 0.189894
R8477 commonsourceibias.n105 commonsourceibias.n86 0.189894
R8478 commonsourceibias.n101 commonsourceibias.n86 0.189894
R8479 commonsourceibias.n101 commonsourceibias.n100 0.189894
R8480 commonsourceibias.n100 commonsourceibias.n88 0.189894
R8481 commonsourceibias.n96 commonsourceibias.n88 0.189894
R8482 commonsourceibias.n96 commonsourceibias.n95 0.189894
R8483 commonsourceibias.n95 commonsourceibias.n90 0.189894
R8484 commonsourceibias.n133 commonsourceibias.n0 0.189894
R8485 commonsourceibias.n133 commonsourceibias.n132 0.189894
R8486 commonsourceibias.n132 commonsourceibias.n2 0.189894
R8487 commonsourceibias.n127 commonsourceibias.n2 0.189894
R8488 commonsourceibias.n127 commonsourceibias.n126 0.189894
R8489 commonsourceibias.n126 commonsourceibias.n125 0.189894
R8490 commonsourceibias.n125 commonsourceibias.n4 0.189894
R8491 commonsourceibias.n120 commonsourceibias.n4 0.189894
R8492 commonsourceibias.n120 commonsourceibias.n119 0.189894
R8493 commonsourceibias.n119 commonsourceibias.n118 0.189894
R8494 commonsourceibias.n118 commonsourceibias.n6 0.189894
R8495 commonsourceibias.n113 commonsourceibias.n6 0.189894
R8496 commonsourceibias.n260 commonsourceibias.n202 0.189894
R8497 commonsourceibias.n260 commonsourceibias.n259 0.189894
R8498 commonsourceibias.n259 commonsourceibias.n204 0.189894
R8499 commonsourceibias.n254 commonsourceibias.n204 0.189894
R8500 commonsourceibias.n254 commonsourceibias.n253 0.189894
R8501 commonsourceibias.n253 commonsourceibias.n252 0.189894
R8502 commonsourceibias.n252 commonsourceibias.n206 0.189894
R8503 commonsourceibias.n247 commonsourceibias.n206 0.189894
R8504 commonsourceibias.n247 commonsourceibias.n246 0.189894
R8505 commonsourceibias.n246 commonsourceibias.n245 0.189894
R8506 commonsourceibias.n245 commonsourceibias.n208 0.189894
R8507 commonsourceibias.n240 commonsourceibias.n208 0.189894
R8508 commonsourceibias.n240 commonsourceibias.n239 0.189894
R8509 commonsourceibias.n239 commonsourceibias.n238 0.189894
R8510 commonsourceibias.n238 commonsourceibias.n211 0.189894
R8511 commonsourceibias.n233 commonsourceibias.n211 0.189894
R8512 commonsourceibias.n233 commonsourceibias.n232 0.189894
R8513 commonsourceibias.n232 commonsourceibias.n213 0.189894
R8514 commonsourceibias.n228 commonsourceibias.n213 0.189894
R8515 commonsourceibias.n228 commonsourceibias.n227 0.189894
R8516 commonsourceibias.n227 commonsourceibias.n215 0.189894
R8517 commonsourceibias.n223 commonsourceibias.n215 0.189894
R8518 commonsourceibias.n223 commonsourceibias.n222 0.189894
R8519 commonsourceibias.n222 commonsourceibias.n217 0.189894
R8520 commonsourceibias.n196 commonsourceibias.n138 0.189894
R8521 commonsourceibias.n196 commonsourceibias.n195 0.189894
R8522 commonsourceibias.n195 commonsourceibias.n140 0.189894
R8523 commonsourceibias.n190 commonsourceibias.n140 0.189894
R8524 commonsourceibias.n190 commonsourceibias.n189 0.189894
R8525 commonsourceibias.n189 commonsourceibias.n188 0.189894
R8526 commonsourceibias.n188 commonsourceibias.n142 0.189894
R8527 commonsourceibias.n183 commonsourceibias.n142 0.189894
R8528 commonsourceibias.n183 commonsourceibias.n182 0.189894
R8529 commonsourceibias.n182 commonsourceibias.n181 0.189894
R8530 commonsourceibias.n181 commonsourceibias.n144 0.189894
R8531 commonsourceibias.n176 commonsourceibias.n144 0.189894
R8532 commonsourceibias.n176 commonsourceibias.n175 0.189894
R8533 commonsourceibias.n175 commonsourceibias.n174 0.189894
R8534 commonsourceibias.n174 commonsourceibias.n147 0.189894
R8535 commonsourceibias.n169 commonsourceibias.n147 0.189894
R8536 commonsourceibias.n169 commonsourceibias.n168 0.189894
R8537 commonsourceibias.n168 commonsourceibias.n149 0.189894
R8538 commonsourceibias.n164 commonsourceibias.n149 0.189894
R8539 commonsourceibias.n164 commonsourceibias.n163 0.189894
R8540 commonsourceibias.n163 commonsourceibias.n151 0.189894
R8541 commonsourceibias.n159 commonsourceibias.n151 0.189894
R8542 commonsourceibias.n159 commonsourceibias.n158 0.189894
R8543 commonsourceibias.n158 commonsourceibias.n153 0.189894
R8544 commonsourceibias.n326 commonsourceibias.n321 0.189894
R8545 commonsourceibias.n327 commonsourceibias.n326 0.189894
R8546 commonsourceibias.n327 commonsourceibias.n319 0.189894
R8547 commonsourceibias.n331 commonsourceibias.n319 0.189894
R8548 commonsourceibias.n332 commonsourceibias.n331 0.189894
R8549 commonsourceibias.n332 commonsourceibias.n317 0.189894
R8550 commonsourceibias.n336 commonsourceibias.n317 0.189894
R8551 commonsourceibias.n337 commonsourceibias.n336 0.189894
R8552 commonsourceibias.n337 commonsourceibias.n315 0.189894
R8553 commonsourceibias.n342 commonsourceibias.n315 0.189894
R8554 commonsourceibias.n343 commonsourceibias.n342 0.189894
R8555 commonsourceibias.n344 commonsourceibias.n343 0.189894
R8556 commonsourceibias.n344 commonsourceibias.n313 0.189894
R8557 commonsourceibias.n350 commonsourceibias.n313 0.189894
R8558 commonsourceibias.n351 commonsourceibias.n350 0.189894
R8559 commonsourceibias.n352 commonsourceibias.n351 0.189894
R8560 commonsourceibias.n352 commonsourceibias.n311 0.189894
R8561 commonsourceibias.n357 commonsourceibias.n311 0.189894
R8562 commonsourceibias.n358 commonsourceibias.n357 0.189894
R8563 commonsourceibias.n359 commonsourceibias.n358 0.189894
R8564 commonsourceibias.n359 commonsourceibias.n309 0.189894
R8565 commonsourceibias.n364 commonsourceibias.n309 0.189894
R8566 commonsourceibias.n365 commonsourceibias.n364 0.189894
R8567 commonsourceibias.n365 commonsourceibias.n307 0.189894
R8568 commonsourceibias.n285 commonsourceibias.n280 0.189894
R8569 commonsourceibias.n286 commonsourceibias.n285 0.189894
R8570 commonsourceibias.n286 commonsourceibias.n278 0.189894
R8571 commonsourceibias.n290 commonsourceibias.n278 0.189894
R8572 commonsourceibias.n291 commonsourceibias.n290 0.189894
R8573 commonsourceibias.n291 commonsourceibias.n276 0.189894
R8574 commonsourceibias.n295 commonsourceibias.n276 0.189894
R8575 commonsourceibias.n296 commonsourceibias.n295 0.189894
R8576 commonsourceibias.n296 commonsourceibias.n274 0.189894
R8577 commonsourceibias.n301 commonsourceibias.n274 0.189894
R8578 commonsourceibias.n378 commonsourceibias.n272 0.189894
R8579 commonsourceibias.n384 commonsourceibias.n272 0.189894
R8580 commonsourceibias.n385 commonsourceibias.n384 0.189894
R8581 commonsourceibias.n386 commonsourceibias.n385 0.189894
R8582 commonsourceibias.n386 commonsourceibias.n270 0.189894
R8583 commonsourceibias.n391 commonsourceibias.n270 0.189894
R8584 commonsourceibias.n392 commonsourceibias.n391 0.189894
R8585 commonsourceibias.n393 commonsourceibias.n392 0.189894
R8586 commonsourceibias.n393 commonsourceibias.n268 0.189894
R8587 commonsourceibias.n398 commonsourceibias.n268 0.189894
R8588 commonsourceibias.n399 commonsourceibias.n398 0.189894
R8589 commonsourceibias.n399 commonsourceibias.n266 0.189894
R8590 commonsourceibias.n487 commonsourceibias.n482 0.189894
R8591 commonsourceibias.n488 commonsourceibias.n487 0.189894
R8592 commonsourceibias.n488 commonsourceibias.n480 0.189894
R8593 commonsourceibias.n492 commonsourceibias.n480 0.189894
R8594 commonsourceibias.n493 commonsourceibias.n492 0.189894
R8595 commonsourceibias.n493 commonsourceibias.n478 0.189894
R8596 commonsourceibias.n497 commonsourceibias.n478 0.189894
R8597 commonsourceibias.n498 commonsourceibias.n497 0.189894
R8598 commonsourceibias.n498 commonsourceibias.n476 0.189894
R8599 commonsourceibias.n503 commonsourceibias.n476 0.189894
R8600 commonsourceibias.n504 commonsourceibias.n503 0.189894
R8601 commonsourceibias.n505 commonsourceibias.n504 0.189894
R8602 commonsourceibias.n505 commonsourceibias.n474 0.189894
R8603 commonsourceibias.n511 commonsourceibias.n474 0.189894
R8604 commonsourceibias.n512 commonsourceibias.n511 0.189894
R8605 commonsourceibias.n513 commonsourceibias.n512 0.189894
R8606 commonsourceibias.n513 commonsourceibias.n472 0.189894
R8607 commonsourceibias.n518 commonsourceibias.n472 0.189894
R8608 commonsourceibias.n519 commonsourceibias.n518 0.189894
R8609 commonsourceibias.n520 commonsourceibias.n519 0.189894
R8610 commonsourceibias.n520 commonsourceibias.n470 0.189894
R8611 commonsourceibias.n525 commonsourceibias.n470 0.189894
R8612 commonsourceibias.n526 commonsourceibias.n525 0.189894
R8613 commonsourceibias.n526 commonsourceibias.n468 0.189894
R8614 commonsourceibias.n423 commonsourceibias.n418 0.189894
R8615 commonsourceibias.n424 commonsourceibias.n423 0.189894
R8616 commonsourceibias.n424 commonsourceibias.n416 0.189894
R8617 commonsourceibias.n428 commonsourceibias.n416 0.189894
R8618 commonsourceibias.n429 commonsourceibias.n428 0.189894
R8619 commonsourceibias.n429 commonsourceibias.n414 0.189894
R8620 commonsourceibias.n433 commonsourceibias.n414 0.189894
R8621 commonsourceibias.n434 commonsourceibias.n433 0.189894
R8622 commonsourceibias.n434 commonsourceibias.n412 0.189894
R8623 commonsourceibias.n439 commonsourceibias.n412 0.189894
R8624 commonsourceibias.n440 commonsourceibias.n439 0.189894
R8625 commonsourceibias.n441 commonsourceibias.n440 0.189894
R8626 commonsourceibias.n441 commonsourceibias.n410 0.189894
R8627 commonsourceibias.n447 commonsourceibias.n410 0.189894
R8628 commonsourceibias.n448 commonsourceibias.n447 0.189894
R8629 commonsourceibias.n449 commonsourceibias.n448 0.189894
R8630 commonsourceibias.n449 commonsourceibias.n408 0.189894
R8631 commonsourceibias.n454 commonsourceibias.n408 0.189894
R8632 commonsourceibias.n455 commonsourceibias.n454 0.189894
R8633 commonsourceibias.n456 commonsourceibias.n455 0.189894
R8634 commonsourceibias.n456 commonsourceibias.n406 0.189894
R8635 commonsourceibias.n461 commonsourceibias.n406 0.189894
R8636 commonsourceibias.n462 commonsourceibias.n461 0.189894
R8637 commonsourceibias.n462 commonsourceibias.n404 0.189894
R8638 commonsourceibias.n112 commonsourceibias.n111 0.170955
R8639 commonsourceibias.n113 commonsourceibias.n112 0.170955
R8640 commonsourceibias.n377 commonsourceibias.n301 0.170955
R8641 commonsourceibias.n378 commonsourceibias.n377 0.170955
R8642 gnd.n2378 gnd.n2377 1758.55
R8643 gnd.n3036 gnd.n1516 931.112
R8644 gnd.n7268 gnd.n172 838.452
R8645 gnd.n7255 gnd.n170 838.452
R8646 gnd.n6714 gnd.n420 838.452
R8647 gnd.n6490 gnd.n395 838.452
R8648 gnd.n5192 gnd.n5191 838.452
R8649 gnd.n5258 gnd.n1239 838.452
R8650 gnd.n1554 gnd.n1505 838.452
R8651 gnd.n4583 gnd.n4582 838.452
R8652 gnd.n7270 gnd.n167 783.196
R8653 gnd.n7130 gnd.n169 783.196
R8654 gnd.n559 gnd.n419 783.196
R8655 gnd.n6691 gnd.n391 783.196
R8656 gnd.n5451 gnd.n1217 783.196
R8657 gnd.n5466 gnd.n1206 783.196
R8658 gnd.n4585 gnd.n4525 783.196
R8659 gnd.n4705 gnd.n1510 783.196
R8660 gnd.n5328 gnd.n1262 771.183
R8661 gnd.n6464 gnd.n571 771.183
R8662 gnd.n5332 gnd.n1244 771.183
R8663 gnd.n6706 gnd.n426 771.183
R8664 gnd.n4364 gnd.n3032 766.379
R8665 gnd.n4280 gnd.n3034 766.379
R8666 gnd.n3575 gnd.n3478 766.379
R8667 gnd.n3571 gnd.n3476 766.379
R8668 gnd.n4361 gnd.n3038 756.769
R8669 gnd.n4330 gnd.n3035 756.769
R8670 gnd.n3668 gnd.n3385 756.769
R8671 gnd.n3666 gnd.n3388 756.769
R8672 gnd.n1684 gnd.n1681 670.282
R8673 gnd.n2379 gnd.n2046 670.282
R8674 gnd.n7039 gnd.n244 670.282
R8675 gnd.n4451 gnd.n1555 670.282
R8676 gnd.n1682 gnd.n1681 585
R8677 gnd.n1681 gnd.n1680 585
R8678 gnd.n2746 gnd.n2745 585
R8679 gnd.n2747 gnd.n2746 585
R8680 gnd.n1679 gnd.n1678 585
R8681 gnd.n2748 gnd.n1679 585
R8682 gnd.n2751 gnd.n2750 585
R8683 gnd.n2750 gnd.n2749 585
R8684 gnd.n1676 gnd.n1675 585
R8685 gnd.n1675 gnd.n1674 585
R8686 gnd.n2756 gnd.n2755 585
R8687 gnd.n2757 gnd.n2756 585
R8688 gnd.n1673 gnd.n1672 585
R8689 gnd.n2758 gnd.n1673 585
R8690 gnd.n2761 gnd.n2760 585
R8691 gnd.n2760 gnd.n2759 585
R8692 gnd.n1670 gnd.n1669 585
R8693 gnd.n1669 gnd.n1668 585
R8694 gnd.n2766 gnd.n2765 585
R8695 gnd.n2767 gnd.n2766 585
R8696 gnd.n1667 gnd.n1666 585
R8697 gnd.n2768 gnd.n1667 585
R8698 gnd.n2771 gnd.n2770 585
R8699 gnd.n2770 gnd.n2769 585
R8700 gnd.n1664 gnd.n1663 585
R8701 gnd.n1663 gnd.n1662 585
R8702 gnd.n2776 gnd.n2775 585
R8703 gnd.n2777 gnd.n2776 585
R8704 gnd.n1661 gnd.n1660 585
R8705 gnd.n2778 gnd.n1661 585
R8706 gnd.n2781 gnd.n2780 585
R8707 gnd.n2780 gnd.n2779 585
R8708 gnd.n1658 gnd.n1657 585
R8709 gnd.n1657 gnd.n1656 585
R8710 gnd.n2786 gnd.n2785 585
R8711 gnd.n2787 gnd.n2786 585
R8712 gnd.n1655 gnd.n1654 585
R8713 gnd.n2788 gnd.n1655 585
R8714 gnd.n2791 gnd.n2790 585
R8715 gnd.n2790 gnd.n2789 585
R8716 gnd.n1652 gnd.n1651 585
R8717 gnd.n1651 gnd.n1650 585
R8718 gnd.n2796 gnd.n2795 585
R8719 gnd.n2797 gnd.n2796 585
R8720 gnd.n1649 gnd.n1648 585
R8721 gnd.n2798 gnd.n1649 585
R8722 gnd.n2801 gnd.n2800 585
R8723 gnd.n2800 gnd.n2799 585
R8724 gnd.n1646 gnd.n1645 585
R8725 gnd.n1645 gnd.n1644 585
R8726 gnd.n2806 gnd.n2805 585
R8727 gnd.n2807 gnd.n2806 585
R8728 gnd.n1643 gnd.n1642 585
R8729 gnd.n2808 gnd.n1643 585
R8730 gnd.n2811 gnd.n2810 585
R8731 gnd.n2810 gnd.n2809 585
R8732 gnd.n1640 gnd.n1639 585
R8733 gnd.n1639 gnd.n1638 585
R8734 gnd.n2816 gnd.n2815 585
R8735 gnd.n2817 gnd.n2816 585
R8736 gnd.n1637 gnd.n1636 585
R8737 gnd.n2818 gnd.n1637 585
R8738 gnd.n2821 gnd.n2820 585
R8739 gnd.n2820 gnd.n2819 585
R8740 gnd.n1634 gnd.n1633 585
R8741 gnd.n1633 gnd.n1632 585
R8742 gnd.n2826 gnd.n2825 585
R8743 gnd.n2827 gnd.n2826 585
R8744 gnd.n1631 gnd.n1630 585
R8745 gnd.n2828 gnd.n1631 585
R8746 gnd.n2831 gnd.n2830 585
R8747 gnd.n2830 gnd.n2829 585
R8748 gnd.n1628 gnd.n1627 585
R8749 gnd.n1627 gnd.n1626 585
R8750 gnd.n2836 gnd.n2835 585
R8751 gnd.n2837 gnd.n2836 585
R8752 gnd.n1625 gnd.n1624 585
R8753 gnd.n2838 gnd.n1625 585
R8754 gnd.n2841 gnd.n2840 585
R8755 gnd.n2840 gnd.n2839 585
R8756 gnd.n1622 gnd.n1621 585
R8757 gnd.n1621 gnd.n1620 585
R8758 gnd.n2846 gnd.n2845 585
R8759 gnd.n2847 gnd.n2846 585
R8760 gnd.n1619 gnd.n1618 585
R8761 gnd.n2848 gnd.n1619 585
R8762 gnd.n2851 gnd.n2850 585
R8763 gnd.n2850 gnd.n2849 585
R8764 gnd.n1616 gnd.n1615 585
R8765 gnd.n1615 gnd.n1614 585
R8766 gnd.n2856 gnd.n2855 585
R8767 gnd.n2857 gnd.n2856 585
R8768 gnd.n1613 gnd.n1612 585
R8769 gnd.n2858 gnd.n1613 585
R8770 gnd.n2861 gnd.n2860 585
R8771 gnd.n2860 gnd.n2859 585
R8772 gnd.n1610 gnd.n1609 585
R8773 gnd.n1609 gnd.n1608 585
R8774 gnd.n2866 gnd.n2865 585
R8775 gnd.n2867 gnd.n2866 585
R8776 gnd.n1607 gnd.n1606 585
R8777 gnd.n2868 gnd.n1607 585
R8778 gnd.n2871 gnd.n2870 585
R8779 gnd.n2870 gnd.n2869 585
R8780 gnd.n1604 gnd.n1603 585
R8781 gnd.n1603 gnd.n1602 585
R8782 gnd.n2876 gnd.n2875 585
R8783 gnd.n2877 gnd.n2876 585
R8784 gnd.n1601 gnd.n1600 585
R8785 gnd.n2878 gnd.n1601 585
R8786 gnd.n2881 gnd.n2880 585
R8787 gnd.n2880 gnd.n2879 585
R8788 gnd.n1598 gnd.n1597 585
R8789 gnd.n1597 gnd.n1596 585
R8790 gnd.n2886 gnd.n2885 585
R8791 gnd.n2887 gnd.n2886 585
R8792 gnd.n1595 gnd.n1594 585
R8793 gnd.n2888 gnd.n1595 585
R8794 gnd.n2891 gnd.n2890 585
R8795 gnd.n2890 gnd.n2889 585
R8796 gnd.n1592 gnd.n1591 585
R8797 gnd.n1591 gnd.n1590 585
R8798 gnd.n2896 gnd.n2895 585
R8799 gnd.n2897 gnd.n2896 585
R8800 gnd.n1589 gnd.n1588 585
R8801 gnd.n2898 gnd.n1589 585
R8802 gnd.n2901 gnd.n2900 585
R8803 gnd.n2900 gnd.n2899 585
R8804 gnd.n1586 gnd.n1585 585
R8805 gnd.n1585 gnd.n1584 585
R8806 gnd.n2906 gnd.n2905 585
R8807 gnd.n2907 gnd.n2906 585
R8808 gnd.n1583 gnd.n1582 585
R8809 gnd.n2908 gnd.n1583 585
R8810 gnd.n2911 gnd.n2910 585
R8811 gnd.n2910 gnd.n2909 585
R8812 gnd.n1580 gnd.n1579 585
R8813 gnd.n1579 gnd.n1578 585
R8814 gnd.n2916 gnd.n2915 585
R8815 gnd.n2917 gnd.n2916 585
R8816 gnd.n1577 gnd.n1576 585
R8817 gnd.n2918 gnd.n1577 585
R8818 gnd.n2921 gnd.n2920 585
R8819 gnd.n2920 gnd.n2919 585
R8820 gnd.n1574 gnd.n1573 585
R8821 gnd.n1573 gnd.n1572 585
R8822 gnd.n2926 gnd.n2925 585
R8823 gnd.n2927 gnd.n2926 585
R8824 gnd.n1571 gnd.n1570 585
R8825 gnd.n2928 gnd.n1571 585
R8826 gnd.n2931 gnd.n2930 585
R8827 gnd.n2930 gnd.n2929 585
R8828 gnd.n1568 gnd.n1567 585
R8829 gnd.n1567 gnd.n1566 585
R8830 gnd.n2936 gnd.n2935 585
R8831 gnd.n2937 gnd.n2936 585
R8832 gnd.n1565 gnd.n1564 585
R8833 gnd.n2938 gnd.n1565 585
R8834 gnd.n2941 gnd.n2940 585
R8835 gnd.n2940 gnd.n2939 585
R8836 gnd.n1562 gnd.n1561 585
R8837 gnd.n1561 gnd.n1560 585
R8838 gnd.n2947 gnd.n2946 585
R8839 gnd.n2948 gnd.n2947 585
R8840 gnd.n1559 gnd.n1558 585
R8841 gnd.n2949 gnd.n1559 585
R8842 gnd.n4415 gnd.n4414 585
R8843 gnd.n4414 gnd.n4413 585
R8844 gnd.n2741 gnd.n1684 585
R8845 gnd.n1687 gnd.n1684 585
R8846 gnd.n2740 gnd.n2739 585
R8847 gnd.n2739 gnd.n2738 585
R8848 gnd.n1686 gnd.n1685 585
R8849 gnd.n2737 gnd.n1686 585
R8850 gnd.n2735 gnd.n2734 585
R8851 gnd.n2736 gnd.n2735 585
R8852 gnd.n2733 gnd.n1689 585
R8853 gnd.n1689 gnd.n1688 585
R8854 gnd.n2732 gnd.n2731 585
R8855 gnd.n2731 gnd.n2730 585
R8856 gnd.n1695 gnd.n1694 585
R8857 gnd.n2729 gnd.n1695 585
R8858 gnd.n2727 gnd.n2726 585
R8859 gnd.n2728 gnd.n2727 585
R8860 gnd.n2725 gnd.n1697 585
R8861 gnd.n1697 gnd.n1696 585
R8862 gnd.n2724 gnd.n2723 585
R8863 gnd.n2723 gnd.n2722 585
R8864 gnd.n1703 gnd.n1702 585
R8865 gnd.n2721 gnd.n1703 585
R8866 gnd.n2719 gnd.n2718 585
R8867 gnd.n2720 gnd.n2719 585
R8868 gnd.n2717 gnd.n1705 585
R8869 gnd.n1705 gnd.n1704 585
R8870 gnd.n2716 gnd.n2715 585
R8871 gnd.n2715 gnd.n2714 585
R8872 gnd.n1711 gnd.n1710 585
R8873 gnd.n2713 gnd.n1711 585
R8874 gnd.n2711 gnd.n2710 585
R8875 gnd.n2712 gnd.n2711 585
R8876 gnd.n2709 gnd.n1713 585
R8877 gnd.n1713 gnd.n1712 585
R8878 gnd.n2708 gnd.n2707 585
R8879 gnd.n2707 gnd.n2706 585
R8880 gnd.n1719 gnd.n1718 585
R8881 gnd.n2705 gnd.n1719 585
R8882 gnd.n2703 gnd.n2702 585
R8883 gnd.n2704 gnd.n2703 585
R8884 gnd.n2701 gnd.n1721 585
R8885 gnd.n1721 gnd.n1720 585
R8886 gnd.n2700 gnd.n2699 585
R8887 gnd.n2699 gnd.n2698 585
R8888 gnd.n1727 gnd.n1726 585
R8889 gnd.n2697 gnd.n1727 585
R8890 gnd.n2695 gnd.n2694 585
R8891 gnd.n2696 gnd.n2695 585
R8892 gnd.n2693 gnd.n1729 585
R8893 gnd.n1729 gnd.n1728 585
R8894 gnd.n2692 gnd.n2691 585
R8895 gnd.n2691 gnd.n2690 585
R8896 gnd.n1735 gnd.n1734 585
R8897 gnd.n2689 gnd.n1735 585
R8898 gnd.n2687 gnd.n2686 585
R8899 gnd.n2688 gnd.n2687 585
R8900 gnd.n2685 gnd.n1737 585
R8901 gnd.n1737 gnd.n1736 585
R8902 gnd.n2684 gnd.n2683 585
R8903 gnd.n2683 gnd.n2682 585
R8904 gnd.n1743 gnd.n1742 585
R8905 gnd.n2681 gnd.n1743 585
R8906 gnd.n2679 gnd.n2678 585
R8907 gnd.n2680 gnd.n2679 585
R8908 gnd.n2677 gnd.n1745 585
R8909 gnd.n1745 gnd.n1744 585
R8910 gnd.n2676 gnd.n2675 585
R8911 gnd.n2675 gnd.n2674 585
R8912 gnd.n1751 gnd.n1750 585
R8913 gnd.n2673 gnd.n1751 585
R8914 gnd.n2671 gnd.n2670 585
R8915 gnd.n2672 gnd.n2671 585
R8916 gnd.n2669 gnd.n1753 585
R8917 gnd.n1753 gnd.n1752 585
R8918 gnd.n2668 gnd.n2667 585
R8919 gnd.n2667 gnd.n2666 585
R8920 gnd.n1759 gnd.n1758 585
R8921 gnd.n2665 gnd.n1759 585
R8922 gnd.n2663 gnd.n2662 585
R8923 gnd.n2664 gnd.n2663 585
R8924 gnd.n2661 gnd.n1761 585
R8925 gnd.n1761 gnd.n1760 585
R8926 gnd.n2660 gnd.n2659 585
R8927 gnd.n2659 gnd.n2658 585
R8928 gnd.n1767 gnd.n1766 585
R8929 gnd.n2657 gnd.n1767 585
R8930 gnd.n2655 gnd.n2654 585
R8931 gnd.n2656 gnd.n2655 585
R8932 gnd.n2653 gnd.n1769 585
R8933 gnd.n1769 gnd.n1768 585
R8934 gnd.n2652 gnd.n2651 585
R8935 gnd.n2651 gnd.n2650 585
R8936 gnd.n1775 gnd.n1774 585
R8937 gnd.n2649 gnd.n1775 585
R8938 gnd.n2647 gnd.n2646 585
R8939 gnd.n2648 gnd.n2647 585
R8940 gnd.n2645 gnd.n1777 585
R8941 gnd.n1777 gnd.n1776 585
R8942 gnd.n2644 gnd.n2643 585
R8943 gnd.n2643 gnd.n2642 585
R8944 gnd.n1783 gnd.n1782 585
R8945 gnd.n2641 gnd.n1783 585
R8946 gnd.n2639 gnd.n2638 585
R8947 gnd.n2640 gnd.n2639 585
R8948 gnd.n2637 gnd.n1785 585
R8949 gnd.n1785 gnd.n1784 585
R8950 gnd.n2636 gnd.n2635 585
R8951 gnd.n2635 gnd.n2634 585
R8952 gnd.n1791 gnd.n1790 585
R8953 gnd.n2633 gnd.n1791 585
R8954 gnd.n2631 gnd.n2630 585
R8955 gnd.n2632 gnd.n2631 585
R8956 gnd.n2629 gnd.n1793 585
R8957 gnd.n1793 gnd.n1792 585
R8958 gnd.n2628 gnd.n2627 585
R8959 gnd.n2627 gnd.n2626 585
R8960 gnd.n1799 gnd.n1798 585
R8961 gnd.n2625 gnd.n1799 585
R8962 gnd.n2623 gnd.n2622 585
R8963 gnd.n2624 gnd.n2623 585
R8964 gnd.n2621 gnd.n1801 585
R8965 gnd.n1801 gnd.n1800 585
R8966 gnd.n2620 gnd.n2619 585
R8967 gnd.n2619 gnd.n2618 585
R8968 gnd.n1807 gnd.n1806 585
R8969 gnd.n2617 gnd.n1807 585
R8970 gnd.n2615 gnd.n2614 585
R8971 gnd.n2616 gnd.n2615 585
R8972 gnd.n2613 gnd.n1809 585
R8973 gnd.n1809 gnd.n1808 585
R8974 gnd.n2612 gnd.n2611 585
R8975 gnd.n2611 gnd.n2610 585
R8976 gnd.n1815 gnd.n1814 585
R8977 gnd.n2609 gnd.n1815 585
R8978 gnd.n2607 gnd.n2606 585
R8979 gnd.n2608 gnd.n2607 585
R8980 gnd.n2605 gnd.n1817 585
R8981 gnd.n1817 gnd.n1816 585
R8982 gnd.n2604 gnd.n2603 585
R8983 gnd.n2603 gnd.n2602 585
R8984 gnd.n1823 gnd.n1822 585
R8985 gnd.n2601 gnd.n1823 585
R8986 gnd.n2599 gnd.n2598 585
R8987 gnd.n2600 gnd.n2599 585
R8988 gnd.n2597 gnd.n1825 585
R8989 gnd.n1825 gnd.n1824 585
R8990 gnd.n2596 gnd.n2595 585
R8991 gnd.n2595 gnd.n2594 585
R8992 gnd.n1831 gnd.n1830 585
R8993 gnd.n2593 gnd.n1831 585
R8994 gnd.n2591 gnd.n2590 585
R8995 gnd.n2592 gnd.n2591 585
R8996 gnd.n2589 gnd.n1833 585
R8997 gnd.n1833 gnd.n1832 585
R8998 gnd.n2588 gnd.n2587 585
R8999 gnd.n2587 gnd.n2586 585
R9000 gnd.n1839 gnd.n1838 585
R9001 gnd.n2585 gnd.n1839 585
R9002 gnd.n2583 gnd.n2582 585
R9003 gnd.n2584 gnd.n2583 585
R9004 gnd.n2581 gnd.n1841 585
R9005 gnd.n1841 gnd.n1840 585
R9006 gnd.n2580 gnd.n2579 585
R9007 gnd.n2579 gnd.n2578 585
R9008 gnd.n1847 gnd.n1846 585
R9009 gnd.n2577 gnd.n1847 585
R9010 gnd.n2575 gnd.n2574 585
R9011 gnd.n2576 gnd.n2575 585
R9012 gnd.n2573 gnd.n1849 585
R9013 gnd.n1849 gnd.n1848 585
R9014 gnd.n2572 gnd.n2571 585
R9015 gnd.n2571 gnd.n2570 585
R9016 gnd.n1855 gnd.n1854 585
R9017 gnd.n2569 gnd.n1855 585
R9018 gnd.n2567 gnd.n2566 585
R9019 gnd.n2568 gnd.n2567 585
R9020 gnd.n2565 gnd.n1857 585
R9021 gnd.n1857 gnd.n1856 585
R9022 gnd.n2564 gnd.n2563 585
R9023 gnd.n2563 gnd.n2562 585
R9024 gnd.n1863 gnd.n1862 585
R9025 gnd.n2561 gnd.n1863 585
R9026 gnd.n2559 gnd.n2558 585
R9027 gnd.n2560 gnd.n2559 585
R9028 gnd.n2557 gnd.n1865 585
R9029 gnd.n1865 gnd.n1864 585
R9030 gnd.n2556 gnd.n2555 585
R9031 gnd.n2555 gnd.n2554 585
R9032 gnd.n1871 gnd.n1870 585
R9033 gnd.n2553 gnd.n1871 585
R9034 gnd.n2551 gnd.n2550 585
R9035 gnd.n2552 gnd.n2551 585
R9036 gnd.n2549 gnd.n1873 585
R9037 gnd.n1873 gnd.n1872 585
R9038 gnd.n2548 gnd.n2547 585
R9039 gnd.n2547 gnd.n2546 585
R9040 gnd.n1879 gnd.n1878 585
R9041 gnd.n2545 gnd.n1879 585
R9042 gnd.n2543 gnd.n2542 585
R9043 gnd.n2544 gnd.n2543 585
R9044 gnd.n2541 gnd.n1881 585
R9045 gnd.n1881 gnd.n1880 585
R9046 gnd.n2540 gnd.n2539 585
R9047 gnd.n2539 gnd.n2538 585
R9048 gnd.n1887 gnd.n1886 585
R9049 gnd.n2537 gnd.n1887 585
R9050 gnd.n2535 gnd.n2534 585
R9051 gnd.n2536 gnd.n2535 585
R9052 gnd.n2533 gnd.n1889 585
R9053 gnd.n1889 gnd.n1888 585
R9054 gnd.n2532 gnd.n2531 585
R9055 gnd.n2531 gnd.n2530 585
R9056 gnd.n1895 gnd.n1894 585
R9057 gnd.n2529 gnd.n1895 585
R9058 gnd.n2527 gnd.n2526 585
R9059 gnd.n2528 gnd.n2527 585
R9060 gnd.n2525 gnd.n1897 585
R9061 gnd.n1897 gnd.n1896 585
R9062 gnd.n2524 gnd.n2523 585
R9063 gnd.n2523 gnd.n2522 585
R9064 gnd.n1903 gnd.n1902 585
R9065 gnd.n2521 gnd.n1903 585
R9066 gnd.n2519 gnd.n2518 585
R9067 gnd.n2520 gnd.n2519 585
R9068 gnd.n2517 gnd.n1905 585
R9069 gnd.n1905 gnd.n1904 585
R9070 gnd.n2516 gnd.n2515 585
R9071 gnd.n2515 gnd.n2514 585
R9072 gnd.n1911 gnd.n1910 585
R9073 gnd.n2513 gnd.n1911 585
R9074 gnd.n2511 gnd.n2510 585
R9075 gnd.n2512 gnd.n2511 585
R9076 gnd.n2509 gnd.n1913 585
R9077 gnd.n1913 gnd.n1912 585
R9078 gnd.n2508 gnd.n2507 585
R9079 gnd.n2507 gnd.n2506 585
R9080 gnd.n1919 gnd.n1918 585
R9081 gnd.n2505 gnd.n1919 585
R9082 gnd.n2503 gnd.n2502 585
R9083 gnd.n2504 gnd.n2503 585
R9084 gnd.n2501 gnd.n1921 585
R9085 gnd.n1921 gnd.n1920 585
R9086 gnd.n2500 gnd.n2499 585
R9087 gnd.n2499 gnd.n2498 585
R9088 gnd.n1927 gnd.n1926 585
R9089 gnd.n2497 gnd.n1927 585
R9090 gnd.n2495 gnd.n2494 585
R9091 gnd.n2496 gnd.n2495 585
R9092 gnd.n2493 gnd.n1929 585
R9093 gnd.n1929 gnd.n1928 585
R9094 gnd.n2492 gnd.n2491 585
R9095 gnd.n2491 gnd.n2490 585
R9096 gnd.n1935 gnd.n1934 585
R9097 gnd.n2489 gnd.n1935 585
R9098 gnd.n2487 gnd.n2486 585
R9099 gnd.n2488 gnd.n2487 585
R9100 gnd.n2485 gnd.n1937 585
R9101 gnd.n1937 gnd.n1936 585
R9102 gnd.n2484 gnd.n2483 585
R9103 gnd.n2483 gnd.n2482 585
R9104 gnd.n1943 gnd.n1942 585
R9105 gnd.n2481 gnd.n1943 585
R9106 gnd.n2479 gnd.n2478 585
R9107 gnd.n2480 gnd.n2479 585
R9108 gnd.n2477 gnd.n1945 585
R9109 gnd.n1945 gnd.n1944 585
R9110 gnd.n2476 gnd.n2475 585
R9111 gnd.n2475 gnd.n2474 585
R9112 gnd.n1951 gnd.n1950 585
R9113 gnd.n2473 gnd.n1951 585
R9114 gnd.n2471 gnd.n2470 585
R9115 gnd.n2472 gnd.n2471 585
R9116 gnd.n2469 gnd.n1953 585
R9117 gnd.n1953 gnd.n1952 585
R9118 gnd.n2468 gnd.n2467 585
R9119 gnd.n2467 gnd.n2466 585
R9120 gnd.n1959 gnd.n1958 585
R9121 gnd.n2465 gnd.n1959 585
R9122 gnd.n2463 gnd.n2462 585
R9123 gnd.n2464 gnd.n2463 585
R9124 gnd.n2461 gnd.n1961 585
R9125 gnd.n1961 gnd.n1960 585
R9126 gnd.n2460 gnd.n2459 585
R9127 gnd.n2459 gnd.n2458 585
R9128 gnd.n1967 gnd.n1966 585
R9129 gnd.n2457 gnd.n1967 585
R9130 gnd.n2455 gnd.n2454 585
R9131 gnd.n2456 gnd.n2455 585
R9132 gnd.n2453 gnd.n1969 585
R9133 gnd.n1969 gnd.n1968 585
R9134 gnd.n2452 gnd.n2451 585
R9135 gnd.n2451 gnd.n2450 585
R9136 gnd.n1975 gnd.n1974 585
R9137 gnd.n2449 gnd.n1975 585
R9138 gnd.n2447 gnd.n2446 585
R9139 gnd.n2448 gnd.n2447 585
R9140 gnd.n2445 gnd.n1977 585
R9141 gnd.n1977 gnd.n1976 585
R9142 gnd.n2444 gnd.n2443 585
R9143 gnd.n2443 gnd.n2442 585
R9144 gnd.n1983 gnd.n1982 585
R9145 gnd.n2441 gnd.n1983 585
R9146 gnd.n2439 gnd.n2438 585
R9147 gnd.n2440 gnd.n2439 585
R9148 gnd.n2437 gnd.n1985 585
R9149 gnd.n1985 gnd.n1984 585
R9150 gnd.n2436 gnd.n2435 585
R9151 gnd.n2435 gnd.n2434 585
R9152 gnd.n1991 gnd.n1990 585
R9153 gnd.n2433 gnd.n1991 585
R9154 gnd.n2431 gnd.n2430 585
R9155 gnd.n2432 gnd.n2431 585
R9156 gnd.n2429 gnd.n1993 585
R9157 gnd.n1993 gnd.n1992 585
R9158 gnd.n2428 gnd.n2427 585
R9159 gnd.n2427 gnd.n2426 585
R9160 gnd.n1999 gnd.n1998 585
R9161 gnd.n2425 gnd.n1999 585
R9162 gnd.n2423 gnd.n2422 585
R9163 gnd.n2424 gnd.n2423 585
R9164 gnd.n2421 gnd.n2001 585
R9165 gnd.n2001 gnd.n2000 585
R9166 gnd.n2420 gnd.n2419 585
R9167 gnd.n2419 gnd.n2418 585
R9168 gnd.n2007 gnd.n2006 585
R9169 gnd.n2417 gnd.n2007 585
R9170 gnd.n2415 gnd.n2414 585
R9171 gnd.n2416 gnd.n2415 585
R9172 gnd.n2413 gnd.n2009 585
R9173 gnd.n2009 gnd.n2008 585
R9174 gnd.n2412 gnd.n2411 585
R9175 gnd.n2411 gnd.n2410 585
R9176 gnd.n2015 gnd.n2014 585
R9177 gnd.n2409 gnd.n2015 585
R9178 gnd.n2407 gnd.n2406 585
R9179 gnd.n2408 gnd.n2407 585
R9180 gnd.n2405 gnd.n2017 585
R9181 gnd.n2017 gnd.n2016 585
R9182 gnd.n2404 gnd.n2403 585
R9183 gnd.n2403 gnd.n2402 585
R9184 gnd.n2023 gnd.n2022 585
R9185 gnd.n2401 gnd.n2023 585
R9186 gnd.n2399 gnd.n2398 585
R9187 gnd.n2400 gnd.n2399 585
R9188 gnd.n2397 gnd.n2025 585
R9189 gnd.n2025 gnd.n2024 585
R9190 gnd.n2396 gnd.n2395 585
R9191 gnd.n2395 gnd.n2394 585
R9192 gnd.n2031 gnd.n2030 585
R9193 gnd.n2393 gnd.n2031 585
R9194 gnd.n2391 gnd.n2390 585
R9195 gnd.n2392 gnd.n2391 585
R9196 gnd.n2389 gnd.n2033 585
R9197 gnd.n2033 gnd.n2032 585
R9198 gnd.n2388 gnd.n2387 585
R9199 gnd.n2387 gnd.n2386 585
R9200 gnd.n2039 gnd.n2038 585
R9201 gnd.n2385 gnd.n2039 585
R9202 gnd.n2383 gnd.n2382 585
R9203 gnd.n2384 gnd.n2383 585
R9204 gnd.n2381 gnd.n2041 585
R9205 gnd.n2041 gnd.n2040 585
R9206 gnd.n2380 gnd.n2379 585
R9207 gnd.n2379 gnd.n2378 585
R9208 gnd.n245 gnd.n243 585
R9209 gnd.n243 gnd.n242 585
R9210 gnd.n2211 gnd.n2207 585
R9211 gnd.n2207 gnd.n2206 585
R9212 gnd.n2213 gnd.n2212 585
R9213 gnd.n2214 gnd.n2213 585
R9214 gnd.n2205 gnd.n2204 585
R9215 gnd.n2215 gnd.n2205 585
R9216 gnd.n2218 gnd.n2217 585
R9217 gnd.n2217 gnd.n2216 585
R9218 gnd.n2219 gnd.n2199 585
R9219 gnd.n2199 gnd.n2198 585
R9220 gnd.n2221 gnd.n2220 585
R9221 gnd.n2222 gnd.n2221 585
R9222 gnd.n2197 gnd.n2196 585
R9223 gnd.n2223 gnd.n2197 585
R9224 gnd.n2226 gnd.n2225 585
R9225 gnd.n2225 gnd.n2224 585
R9226 gnd.n2227 gnd.n2191 585
R9227 gnd.n2191 gnd.n2190 585
R9228 gnd.n2229 gnd.n2228 585
R9229 gnd.n2230 gnd.n2229 585
R9230 gnd.n2189 gnd.n2188 585
R9231 gnd.n2231 gnd.n2189 585
R9232 gnd.n2234 gnd.n2233 585
R9233 gnd.n2233 gnd.n2232 585
R9234 gnd.n2235 gnd.n2183 585
R9235 gnd.n2183 gnd.n2182 585
R9236 gnd.n2237 gnd.n2236 585
R9237 gnd.n2238 gnd.n2237 585
R9238 gnd.n2181 gnd.n2180 585
R9239 gnd.n2239 gnd.n2181 585
R9240 gnd.n2242 gnd.n2241 585
R9241 gnd.n2241 gnd.n2240 585
R9242 gnd.n2243 gnd.n2175 585
R9243 gnd.n2175 gnd.n2174 585
R9244 gnd.n2245 gnd.n2244 585
R9245 gnd.n2246 gnd.n2245 585
R9246 gnd.n2173 gnd.n2172 585
R9247 gnd.n2247 gnd.n2173 585
R9248 gnd.n2250 gnd.n2249 585
R9249 gnd.n2249 gnd.n2248 585
R9250 gnd.n2251 gnd.n2167 585
R9251 gnd.n2167 gnd.n2166 585
R9252 gnd.n2253 gnd.n2252 585
R9253 gnd.n2254 gnd.n2253 585
R9254 gnd.n2165 gnd.n2164 585
R9255 gnd.n2255 gnd.n2165 585
R9256 gnd.n2258 gnd.n2257 585
R9257 gnd.n2257 gnd.n2256 585
R9258 gnd.n2259 gnd.n2159 585
R9259 gnd.n2159 gnd.n2158 585
R9260 gnd.n2261 gnd.n2260 585
R9261 gnd.n2262 gnd.n2261 585
R9262 gnd.n2157 gnd.n2156 585
R9263 gnd.n2263 gnd.n2157 585
R9264 gnd.n2266 gnd.n2265 585
R9265 gnd.n2265 gnd.n2264 585
R9266 gnd.n2267 gnd.n2151 585
R9267 gnd.n2151 gnd.n2150 585
R9268 gnd.n2269 gnd.n2268 585
R9269 gnd.n2270 gnd.n2269 585
R9270 gnd.n2149 gnd.n2148 585
R9271 gnd.n2271 gnd.n2149 585
R9272 gnd.n2274 gnd.n2273 585
R9273 gnd.n2273 gnd.n2272 585
R9274 gnd.n2275 gnd.n2143 585
R9275 gnd.n2143 gnd.n2142 585
R9276 gnd.n2277 gnd.n2276 585
R9277 gnd.n2278 gnd.n2277 585
R9278 gnd.n2141 gnd.n2140 585
R9279 gnd.n2279 gnd.n2141 585
R9280 gnd.n2282 gnd.n2281 585
R9281 gnd.n2281 gnd.n2280 585
R9282 gnd.n2283 gnd.n2135 585
R9283 gnd.n2135 gnd.n2134 585
R9284 gnd.n2285 gnd.n2284 585
R9285 gnd.n2286 gnd.n2285 585
R9286 gnd.n2133 gnd.n2132 585
R9287 gnd.n2287 gnd.n2133 585
R9288 gnd.n2290 gnd.n2289 585
R9289 gnd.n2289 gnd.n2288 585
R9290 gnd.n2291 gnd.n2127 585
R9291 gnd.n2127 gnd.n2126 585
R9292 gnd.n2293 gnd.n2292 585
R9293 gnd.n2294 gnd.n2293 585
R9294 gnd.n2125 gnd.n2124 585
R9295 gnd.n2295 gnd.n2125 585
R9296 gnd.n2298 gnd.n2297 585
R9297 gnd.n2297 gnd.n2296 585
R9298 gnd.n2299 gnd.n2119 585
R9299 gnd.n2119 gnd.n2118 585
R9300 gnd.n2301 gnd.n2300 585
R9301 gnd.n2302 gnd.n2301 585
R9302 gnd.n2117 gnd.n2116 585
R9303 gnd.n2303 gnd.n2117 585
R9304 gnd.n2306 gnd.n2305 585
R9305 gnd.n2305 gnd.n2304 585
R9306 gnd.n2307 gnd.n2111 585
R9307 gnd.n2111 gnd.n2110 585
R9308 gnd.n2309 gnd.n2308 585
R9309 gnd.n2310 gnd.n2309 585
R9310 gnd.n2109 gnd.n2108 585
R9311 gnd.n2311 gnd.n2109 585
R9312 gnd.n2314 gnd.n2313 585
R9313 gnd.n2313 gnd.n2312 585
R9314 gnd.n2315 gnd.n2103 585
R9315 gnd.n2103 gnd.n2102 585
R9316 gnd.n2317 gnd.n2316 585
R9317 gnd.n2318 gnd.n2317 585
R9318 gnd.n2101 gnd.n2100 585
R9319 gnd.n2319 gnd.n2101 585
R9320 gnd.n2322 gnd.n2321 585
R9321 gnd.n2321 gnd.n2320 585
R9322 gnd.n2323 gnd.n2095 585
R9323 gnd.n2095 gnd.n2094 585
R9324 gnd.n2325 gnd.n2324 585
R9325 gnd.n2326 gnd.n2325 585
R9326 gnd.n2093 gnd.n2092 585
R9327 gnd.n2327 gnd.n2093 585
R9328 gnd.n2330 gnd.n2329 585
R9329 gnd.n2329 gnd.n2328 585
R9330 gnd.n2331 gnd.n2087 585
R9331 gnd.n2087 gnd.n2086 585
R9332 gnd.n2333 gnd.n2332 585
R9333 gnd.n2334 gnd.n2333 585
R9334 gnd.n2085 gnd.n2084 585
R9335 gnd.n2335 gnd.n2085 585
R9336 gnd.n2338 gnd.n2337 585
R9337 gnd.n2337 gnd.n2336 585
R9338 gnd.n2339 gnd.n2079 585
R9339 gnd.n2079 gnd.n2078 585
R9340 gnd.n2341 gnd.n2340 585
R9341 gnd.n2342 gnd.n2341 585
R9342 gnd.n2077 gnd.n2076 585
R9343 gnd.n2343 gnd.n2077 585
R9344 gnd.n2346 gnd.n2345 585
R9345 gnd.n2345 gnd.n2344 585
R9346 gnd.n2347 gnd.n2071 585
R9347 gnd.n2071 gnd.n2070 585
R9348 gnd.n2349 gnd.n2348 585
R9349 gnd.n2350 gnd.n2349 585
R9350 gnd.n2069 gnd.n2068 585
R9351 gnd.n2351 gnd.n2069 585
R9352 gnd.n2354 gnd.n2353 585
R9353 gnd.n2353 gnd.n2352 585
R9354 gnd.n2355 gnd.n2063 585
R9355 gnd.n2063 gnd.n2062 585
R9356 gnd.n2357 gnd.n2356 585
R9357 gnd.n2358 gnd.n2357 585
R9358 gnd.n2061 gnd.n2060 585
R9359 gnd.n2359 gnd.n2061 585
R9360 gnd.n2362 gnd.n2361 585
R9361 gnd.n2361 gnd.n2360 585
R9362 gnd.n2363 gnd.n2056 585
R9363 gnd.n2056 gnd.n2055 585
R9364 gnd.n2365 gnd.n2364 585
R9365 gnd.n2366 gnd.n2365 585
R9366 gnd.n2054 gnd.n2053 585
R9367 gnd.n2367 gnd.n2054 585
R9368 gnd.n2370 gnd.n2369 585
R9369 gnd.n2369 gnd.n2368 585
R9370 gnd.n2050 gnd.n2048 585
R9371 gnd.n2048 gnd.n2047 585
R9372 gnd.n2375 gnd.n2374 585
R9373 gnd.n2376 gnd.n2375 585
R9374 gnd.n2049 gnd.n2046 585
R9375 gnd.n2377 gnd.n2046 585
R9376 gnd.n5191 gnd.n1210 585
R9377 gnd.n5191 gnd.n5190 585
R9378 gnd.n5352 gnd.n1215 585
R9379 gnd.n5458 gnd.n1215 585
R9380 gnd.n5353 gnd.n1227 585
R9381 gnd.n5026 gnd.n1227 585
R9382 gnd.n5355 gnd.n5354 585
R9383 gnd.n5356 gnd.n5355 585
R9384 gnd.n1228 gnd.n1226 585
R9385 gnd.n5346 gnd.n1226 585
R9386 gnd.n5004 gnd.n1285 585
R9387 gnd.n5016 gnd.n1285 585
R9388 gnd.n5005 gnd.n1296 585
R9389 gnd.n1296 gnd.n1284 585
R9390 gnd.n5007 gnd.n5006 585
R9391 gnd.n5008 gnd.n5007 585
R9392 gnd.n1297 gnd.n1295 585
R9393 gnd.n4996 gnd.n1295 585
R9394 gnd.n4969 gnd.n4968 585
R9395 gnd.n4968 gnd.n4967 585
R9396 gnd.n4970 gnd.n1312 585
R9397 gnd.n4984 gnd.n1312 585
R9398 gnd.n4971 gnd.n1323 585
R9399 gnd.n4961 gnd.n1323 585
R9400 gnd.n4973 gnd.n4972 585
R9401 gnd.n4974 gnd.n4973 585
R9402 gnd.n1324 gnd.n1322 585
R9403 gnd.n4940 gnd.n1322 585
R9404 gnd.n4890 gnd.n4889 585
R9405 gnd.n4889 gnd.n1334 585
R9406 gnd.n4891 gnd.n1345 585
R9407 gnd.n4931 gnd.n1345 585
R9408 gnd.n4892 gnd.n1401 585
R9409 gnd.n4881 gnd.n1401 585
R9410 gnd.n4894 gnd.n4893 585
R9411 gnd.n4895 gnd.n4894 585
R9412 gnd.n1402 gnd.n1389 585
R9413 gnd.n4900 gnd.n1389 585
R9414 gnd.n4876 gnd.n4875 585
R9415 gnd.n4875 gnd.n1385 585
R9416 gnd.n4874 gnd.n4873 585
R9417 gnd.n4874 gnd.n1378 585
R9418 gnd.n1369 gnd.n1368 585
R9419 gnd.n4909 gnd.n1369 585
R9420 gnd.n4916 gnd.n4915 585
R9421 gnd.n4915 gnd.n4914 585
R9422 gnd.n4917 gnd.n1363 585
R9423 gnd.n4864 gnd.n1363 585
R9424 gnd.n4919 gnd.n4918 585
R9425 gnd.n4920 gnd.n4919 585
R9426 gnd.n1364 gnd.n1362 585
R9427 gnd.n4853 gnd.n1362 585
R9428 gnd.n4783 gnd.n4782 585
R9429 gnd.n4782 gnd.n1415 585
R9430 gnd.n1441 gnd.n1424 585
R9431 gnd.n4827 gnd.n1424 585
R9432 gnd.n4814 gnd.n4813 585
R9433 gnd.n4813 gnd.n4812 585
R9434 gnd.n4815 gnd.n1436 585
R9435 gnd.n4793 gnd.n1436 585
R9436 gnd.n4817 gnd.n4816 585
R9437 gnd.n4818 gnd.n4817 585
R9438 gnd.n1437 gnd.n1435 585
R9439 gnd.n4799 gnd.n1435 585
R9440 gnd.n4776 gnd.n4775 585
R9441 gnd.n4775 gnd.n4774 585
R9442 gnd.n1459 gnd.n1458 585
R9443 gnd.n4759 gnd.n1459 585
R9444 gnd.n4765 gnd.n4764 585
R9445 gnd.n4766 gnd.n4765 585
R9446 gnd.n1472 gnd.n1471 585
R9447 gnd.n4750 gnd.n1471 585
R9448 gnd.n4735 gnd.n1483 585
R9449 gnd.n4747 gnd.n1483 585
R9450 gnd.n4736 gnd.n1494 585
R9451 gnd.n4722 gnd.n1494 585
R9452 gnd.n4738 gnd.n4737 585
R9453 gnd.n4739 gnd.n4738 585
R9454 gnd.n1495 gnd.n1493 585
R9455 gnd.n4728 gnd.n1493 585
R9456 gnd.n4521 gnd.n4520 585
R9457 gnd.n4520 gnd.n4519 585
R9458 gnd.n4518 gnd.n1509 585
R9459 gnd.n4714 gnd.n1509 585
R9460 gnd.n4583 gnd.n4517 585
R9461 gnd.n4584 gnd.n4583 585
R9462 gnd.n4582 gnd.n4581 585
R9463 gnd.n4580 gnd.n4579 585
R9464 gnd.n4578 gnd.n4577 585
R9465 gnd.n4576 gnd.n4575 585
R9466 gnd.n4574 gnd.n4573 585
R9467 gnd.n4572 gnd.n4571 585
R9468 gnd.n4570 gnd.n4569 585
R9469 gnd.n4568 gnd.n4567 585
R9470 gnd.n4566 gnd.n4565 585
R9471 gnd.n4564 gnd.n4563 585
R9472 gnd.n4562 gnd.n4561 585
R9473 gnd.n4560 gnd.n4559 585
R9474 gnd.n4558 gnd.n4557 585
R9475 gnd.n4556 gnd.n4555 585
R9476 gnd.n4554 gnd.n4553 585
R9477 gnd.n4552 gnd.n4551 585
R9478 gnd.n4550 gnd.n4549 585
R9479 gnd.n4544 gnd.n4541 585
R9480 gnd.n4545 gnd.n1554 585
R9481 gnd.n4703 gnd.n1554 585
R9482 gnd.n5259 gnd.n5258 585
R9483 gnd.n5260 gnd.n5256 585
R9484 gnd.n5271 gnd.n5253 585
R9485 gnd.n5272 gnd.n5251 585
R9486 gnd.n5250 gnd.n5243 585
R9487 gnd.n5279 gnd.n5242 585
R9488 gnd.n5280 gnd.n5241 585
R9489 gnd.n5239 gnd.n5231 585
R9490 gnd.n5287 gnd.n5230 585
R9491 gnd.n5288 gnd.n5228 585
R9492 gnd.n5227 gnd.n5220 585
R9493 gnd.n5295 gnd.n5219 585
R9494 gnd.n5296 gnd.n5218 585
R9495 gnd.n5216 gnd.n5208 585
R9496 gnd.n5303 gnd.n5207 585
R9497 gnd.n5304 gnd.n5205 585
R9498 gnd.n5204 gnd.n5194 585
R9499 gnd.n5311 gnd.n5193 585
R9500 gnd.n5312 gnd.n5192 585
R9501 gnd.n5192 gnd.n1156 585
R9502 gnd.n5338 gnd.n1239 585
R9503 gnd.n5190 gnd.n1239 585
R9504 gnd.n5339 gnd.n1213 585
R9505 gnd.n5458 gnd.n1213 585
R9506 gnd.n5340 gnd.n1238 585
R9507 gnd.n5026 gnd.n1238 585
R9508 gnd.n1235 gnd.n1224 585
R9509 gnd.n5356 gnd.n1224 585
R9510 gnd.n5345 gnd.n5344 585
R9511 gnd.n5346 gnd.n5345 585
R9512 gnd.n1234 gnd.n1233 585
R9513 gnd.n5016 gnd.n1233 585
R9514 gnd.n4990 gnd.n4989 585
R9515 gnd.n4989 gnd.n1284 585
R9516 gnd.n1305 gnd.n1293 585
R9517 gnd.n5008 gnd.n1293 585
R9518 gnd.n4995 gnd.n4994 585
R9519 gnd.n4996 gnd.n4995 585
R9520 gnd.n1304 gnd.n1303 585
R9521 gnd.n4967 gnd.n1303 585
R9522 gnd.n4986 gnd.n4985 585
R9523 gnd.n4985 gnd.n4984 585
R9524 gnd.n1308 gnd.n1307 585
R9525 gnd.n4961 gnd.n1308 585
R9526 gnd.n1338 gnd.n1321 585
R9527 gnd.n4974 gnd.n1321 585
R9528 gnd.n4939 gnd.n4938 585
R9529 gnd.n4940 gnd.n4939 585
R9530 gnd.n1337 gnd.n1336 585
R9531 gnd.n1336 gnd.n1334 585
R9532 gnd.n4933 gnd.n4932 585
R9533 gnd.n4932 gnd.n4931 585
R9534 gnd.n1341 gnd.n1340 585
R9535 gnd.n4881 gnd.n1341 585
R9536 gnd.n4841 gnd.n1393 585
R9537 gnd.n4895 gnd.n1393 585
R9538 gnd.n4842 gnd.n1387 585
R9539 gnd.n4900 gnd.n1387 585
R9540 gnd.n4843 gnd.n4839 585
R9541 gnd.n4839 gnd.n1385 585
R9542 gnd.n4838 gnd.n4836 585
R9543 gnd.n4838 gnd.n1378 585
R9544 gnd.n4847 gnd.n1377 585
R9545 gnd.n4909 gnd.n1377 585
R9546 gnd.n4848 gnd.n1371 585
R9547 gnd.n4914 gnd.n1371 585
R9548 gnd.n4849 gnd.n1410 585
R9549 gnd.n4864 gnd.n1410 585
R9550 gnd.n4850 gnd.n1360 585
R9551 gnd.n4920 gnd.n1360 585
R9552 gnd.n4852 gnd.n4851 585
R9553 gnd.n4853 gnd.n4852 585
R9554 gnd.n1418 gnd.n1417 585
R9555 gnd.n1417 gnd.n1415 585
R9556 gnd.n4829 gnd.n4828 585
R9557 gnd.n4828 gnd.n4827 585
R9558 gnd.n1421 gnd.n1420 585
R9559 gnd.n4812 gnd.n1421 585
R9560 gnd.n4795 gnd.n4794 585
R9561 gnd.n4794 gnd.n4793 585
R9562 gnd.n4796 gnd.n1433 585
R9563 gnd.n4818 gnd.n1433 585
R9564 gnd.n4798 gnd.n4797 585
R9565 gnd.n4799 gnd.n4798 585
R9566 gnd.n1452 gnd.n1451 585
R9567 gnd.n4774 gnd.n1451 585
R9568 gnd.n4758 gnd.n4757 585
R9569 gnd.n4759 gnd.n4758 585
R9570 gnd.n1475 gnd.n1469 585
R9571 gnd.n4766 gnd.n1469 585
R9572 gnd.n4752 gnd.n4751 585
R9573 gnd.n4751 gnd.n4750 585
R9574 gnd.n1478 gnd.n1477 585
R9575 gnd.n4747 gnd.n1478 585
R9576 gnd.n4724 gnd.n4723 585
R9577 gnd.n4723 gnd.n4722 585
R9578 gnd.n4725 gnd.n1491 585
R9579 gnd.n4739 gnd.n1491 585
R9580 gnd.n4727 gnd.n4726 585
R9581 gnd.n4728 gnd.n4727 585
R9582 gnd.n1502 gnd.n1501 585
R9583 gnd.n4519 gnd.n1501 585
R9584 gnd.n4716 gnd.n4715 585
R9585 gnd.n4715 gnd.n4714 585
R9586 gnd.n1505 gnd.n1504 585
R9587 gnd.n4584 gnd.n1505 585
R9588 gnd.n4365 gnd.n4364 585
R9589 gnd.n4364 gnd.n4363 585
R9590 gnd.n4366 gnd.n3027 585
R9591 gnd.n4273 gnd.n3027 585
R9592 gnd.n4368 gnd.n4367 585
R9593 gnd.n4369 gnd.n4368 585
R9594 gnd.n3028 gnd.n3026 585
R9595 gnd.n3026 gnd.n3022 585
R9596 gnd.n3007 gnd.n3006 585
R9597 gnd.n3011 gnd.n3007 585
R9598 gnd.n4379 gnd.n4378 585
R9599 gnd.n4378 gnd.n4377 585
R9600 gnd.n4380 gnd.n3001 585
R9601 gnd.n4262 gnd.n3001 585
R9602 gnd.n4382 gnd.n4381 585
R9603 gnd.n4383 gnd.n4382 585
R9604 gnd.n3002 gnd.n3000 585
R9605 gnd.n3000 gnd.n2996 585
R9606 gnd.n2982 gnd.n2981 585
R9607 gnd.n4255 gnd.n2982 585
R9608 gnd.n4393 gnd.n4392 585
R9609 gnd.n4392 gnd.n4391 585
R9610 gnd.n4394 gnd.n2976 585
R9611 gnd.n3922 gnd.n2976 585
R9612 gnd.n4396 gnd.n4395 585
R9613 gnd.n4397 gnd.n4396 585
R9614 gnd.n2977 gnd.n2975 585
R9615 gnd.n2975 gnd.n2971 585
R9616 gnd.n2959 gnd.n2958 585
R9617 gnd.n3930 gnd.n2959 585
R9618 gnd.n4407 gnd.n4406 585
R9619 gnd.n4406 gnd.n4405 585
R9620 gnd.n4408 gnd.n2953 585
R9621 gnd.n3130 gnd.n2953 585
R9622 gnd.n4410 gnd.n4409 585
R9623 gnd.n4411 gnd.n4410 585
R9624 gnd.n2954 gnd.n2952 585
R9625 gnd.n3939 gnd.n2952 585
R9626 gnd.n3904 gnd.n3146 585
R9627 gnd.n3146 gnd.n3136 585
R9628 gnd.n3906 gnd.n3905 585
R9629 gnd.n3907 gnd.n3906 585
R9630 gnd.n3147 gnd.n3145 585
R9631 gnd.n3155 gnd.n3145 585
R9632 gnd.n3880 gnd.n3167 585
R9633 gnd.n3167 gnd.n3154 585
R9634 gnd.n3882 gnd.n3881 585
R9635 gnd.n3883 gnd.n3882 585
R9636 gnd.n3168 gnd.n3166 585
R9637 gnd.n3166 gnd.n3162 585
R9638 gnd.n3868 gnd.n3867 585
R9639 gnd.n3867 gnd.n3866 585
R9640 gnd.n3173 gnd.n3172 585
R9641 gnd.n3182 gnd.n3173 585
R9642 gnd.n3857 gnd.n3856 585
R9643 gnd.n3856 gnd.n3855 585
R9644 gnd.n3180 gnd.n3179 585
R9645 gnd.n3843 gnd.n3180 585
R9646 gnd.n3281 gnd.n3280 585
R9647 gnd.n3281 gnd.n3189 585
R9648 gnd.n3800 gnd.n3799 585
R9649 gnd.n3799 gnd.n3798 585
R9650 gnd.n3801 gnd.n3275 585
R9651 gnd.n3286 gnd.n3275 585
R9652 gnd.n3803 gnd.n3802 585
R9653 gnd.n3804 gnd.n3803 585
R9654 gnd.n3276 gnd.n3274 585
R9655 gnd.n3299 gnd.n3274 585
R9656 gnd.n3259 gnd.n3258 585
R9657 gnd.n3262 gnd.n3259 585
R9658 gnd.n3814 gnd.n3813 585
R9659 gnd.n3813 gnd.n3812 585
R9660 gnd.n3815 gnd.n3253 585
R9661 gnd.n3774 gnd.n3253 585
R9662 gnd.n3817 gnd.n3816 585
R9663 gnd.n3818 gnd.n3817 585
R9664 gnd.n3254 gnd.n3252 585
R9665 gnd.n3313 gnd.n3252 585
R9666 gnd.n3766 gnd.n3765 585
R9667 gnd.n3765 gnd.n3764 585
R9668 gnd.n3310 gnd.n3309 585
R9669 gnd.n3748 gnd.n3310 585
R9670 gnd.n3735 gnd.n3329 585
R9671 gnd.n3329 gnd.n3328 585
R9672 gnd.n3737 gnd.n3736 585
R9673 gnd.n3738 gnd.n3737 585
R9674 gnd.n3330 gnd.n3327 585
R9675 gnd.n3336 gnd.n3327 585
R9676 gnd.n3716 gnd.n3715 585
R9677 gnd.n3717 gnd.n3716 585
R9678 gnd.n3347 gnd.n3346 585
R9679 gnd.n3346 gnd.n3342 585
R9680 gnd.n3706 gnd.n3705 585
R9681 gnd.n3707 gnd.n3706 585
R9682 gnd.n3357 gnd.n3356 585
R9683 gnd.n3362 gnd.n3356 585
R9684 gnd.n3684 gnd.n3375 585
R9685 gnd.n3375 gnd.n3361 585
R9686 gnd.n3686 gnd.n3685 585
R9687 gnd.n3687 gnd.n3686 585
R9688 gnd.n3376 gnd.n3374 585
R9689 gnd.n3374 gnd.n3370 585
R9690 gnd.n3675 gnd.n3674 585
R9691 gnd.n3676 gnd.n3675 585
R9692 gnd.n3383 gnd.n3382 585
R9693 gnd.n3387 gnd.n3382 585
R9694 gnd.n3652 gnd.n3404 585
R9695 gnd.n3404 gnd.n3386 585
R9696 gnd.n3654 gnd.n3653 585
R9697 gnd.n3655 gnd.n3654 585
R9698 gnd.n3405 gnd.n3403 585
R9699 gnd.n3403 gnd.n3394 585
R9700 gnd.n3647 gnd.n3646 585
R9701 gnd.n3646 gnd.n3645 585
R9702 gnd.n3452 gnd.n3451 585
R9703 gnd.n3453 gnd.n3452 585
R9704 gnd.n3606 gnd.n3605 585
R9705 gnd.n3607 gnd.n3606 585
R9706 gnd.n3462 gnd.n3461 585
R9707 gnd.n3461 gnd.n3460 585
R9708 gnd.n3601 gnd.n3600 585
R9709 gnd.n3600 gnd.n3599 585
R9710 gnd.n3465 gnd.n3464 585
R9711 gnd.n3466 gnd.n3465 585
R9712 gnd.n3590 gnd.n3589 585
R9713 gnd.n3591 gnd.n3590 585
R9714 gnd.n3473 gnd.n3472 585
R9715 gnd.n3582 gnd.n3472 585
R9716 gnd.n3585 gnd.n3584 585
R9717 gnd.n3584 gnd.n3583 585
R9718 gnd.n3476 gnd.n3475 585
R9719 gnd.n3477 gnd.n3476 585
R9720 gnd.n3571 gnd.n3570 585
R9721 gnd.n3569 gnd.n3495 585
R9722 gnd.n3568 gnd.n3494 585
R9723 gnd.n3573 gnd.n3494 585
R9724 gnd.n3567 gnd.n3566 585
R9725 gnd.n3565 gnd.n3564 585
R9726 gnd.n3563 gnd.n3562 585
R9727 gnd.n3561 gnd.n3560 585
R9728 gnd.n3559 gnd.n3558 585
R9729 gnd.n3557 gnd.n3556 585
R9730 gnd.n3555 gnd.n3554 585
R9731 gnd.n3553 gnd.n3552 585
R9732 gnd.n3551 gnd.n3550 585
R9733 gnd.n3549 gnd.n3548 585
R9734 gnd.n3547 gnd.n3546 585
R9735 gnd.n3545 gnd.n3544 585
R9736 gnd.n3543 gnd.n3542 585
R9737 gnd.n3541 gnd.n3540 585
R9738 gnd.n3539 gnd.n3538 585
R9739 gnd.n3537 gnd.n3536 585
R9740 gnd.n3535 gnd.n3534 585
R9741 gnd.n3533 gnd.n3532 585
R9742 gnd.n3531 gnd.n3530 585
R9743 gnd.n3529 gnd.n3528 585
R9744 gnd.n3527 gnd.n3526 585
R9745 gnd.n3525 gnd.n3524 585
R9746 gnd.n3482 gnd.n3481 585
R9747 gnd.n3576 gnd.n3575 585
R9748 gnd.n4281 gnd.n4280 585
R9749 gnd.n4282 gnd.n3115 585
R9750 gnd.n4284 gnd.n4283 585
R9751 gnd.n4286 gnd.n3114 585
R9752 gnd.n4288 gnd.n4287 585
R9753 gnd.n4289 gnd.n3105 585
R9754 gnd.n4291 gnd.n4290 585
R9755 gnd.n4293 gnd.n3103 585
R9756 gnd.n4295 gnd.n4294 585
R9757 gnd.n4296 gnd.n3098 585
R9758 gnd.n4298 gnd.n4297 585
R9759 gnd.n4300 gnd.n3096 585
R9760 gnd.n4302 gnd.n4301 585
R9761 gnd.n4303 gnd.n3091 585
R9762 gnd.n4305 gnd.n4304 585
R9763 gnd.n4307 gnd.n3089 585
R9764 gnd.n4309 gnd.n4308 585
R9765 gnd.n4310 gnd.n3084 585
R9766 gnd.n4312 gnd.n4311 585
R9767 gnd.n4314 gnd.n3082 585
R9768 gnd.n4316 gnd.n4315 585
R9769 gnd.n4317 gnd.n3077 585
R9770 gnd.n4319 gnd.n4318 585
R9771 gnd.n4321 gnd.n3075 585
R9772 gnd.n4323 gnd.n4322 585
R9773 gnd.n4324 gnd.n3073 585
R9774 gnd.n4325 gnd.n3032 585
R9775 gnd.n3036 gnd.n3032 585
R9776 gnd.n4276 gnd.n3034 585
R9777 gnd.n4363 gnd.n3034 585
R9778 gnd.n4275 gnd.n4274 585
R9779 gnd.n4274 gnd.n4273 585
R9780 gnd.n4272 gnd.n3024 585
R9781 gnd.n4369 gnd.n3024 585
R9782 gnd.n4266 gnd.n3120 585
R9783 gnd.n4266 gnd.n3022 585
R9784 gnd.n4268 gnd.n4267 585
R9785 gnd.n4267 gnd.n3011 585
R9786 gnd.n4265 gnd.n3009 585
R9787 gnd.n4377 gnd.n3009 585
R9788 gnd.n4264 gnd.n4263 585
R9789 gnd.n4263 gnd.n4262 585
R9790 gnd.n3122 gnd.n2998 585
R9791 gnd.n4383 gnd.n2998 585
R9792 gnd.n4258 gnd.n4257 585
R9793 gnd.n4257 gnd.n2996 585
R9794 gnd.n4256 gnd.n3124 585
R9795 gnd.n4256 gnd.n4255 585
R9796 gnd.n3921 gnd.n2984 585
R9797 gnd.n4391 gnd.n2984 585
R9798 gnd.n3924 gnd.n3923 585
R9799 gnd.n3923 gnd.n3922 585
R9800 gnd.n3925 gnd.n2973 585
R9801 gnd.n4397 gnd.n2973 585
R9802 gnd.n3927 gnd.n3926 585
R9803 gnd.n3927 gnd.n2971 585
R9804 gnd.n3932 gnd.n3931 585
R9805 gnd.n3931 gnd.n3930 585
R9806 gnd.n3933 gnd.n2961 585
R9807 gnd.n4405 gnd.n2961 585
R9808 gnd.n3935 gnd.n3934 585
R9809 gnd.n3934 gnd.n3130 585
R9810 gnd.n3936 gnd.n2951 585
R9811 gnd.n4411 gnd.n2951 585
R9812 gnd.n3938 gnd.n3937 585
R9813 gnd.n3939 gnd.n3938 585
R9814 gnd.n3139 gnd.n3138 585
R9815 gnd.n3138 gnd.n3136 585
R9816 gnd.n3909 gnd.n3908 585
R9817 gnd.n3908 gnd.n3907 585
R9818 gnd.n3142 gnd.n3141 585
R9819 gnd.n3155 gnd.n3142 585
R9820 gnd.n3831 gnd.n3830 585
R9821 gnd.n3830 gnd.n3154 585
R9822 gnd.n3832 gnd.n3164 585
R9823 gnd.n3883 gnd.n3164 585
R9824 gnd.n3834 gnd.n3833 585
R9825 gnd.n3833 gnd.n3162 585
R9826 gnd.n3835 gnd.n3175 585
R9827 gnd.n3866 gnd.n3175 585
R9828 gnd.n3837 gnd.n3836 585
R9829 gnd.n3836 gnd.n3182 585
R9830 gnd.n3838 gnd.n3181 585
R9831 gnd.n3855 gnd.n3181 585
R9832 gnd.n3840 gnd.n3839 585
R9833 gnd.n3843 gnd.n3840 585
R9834 gnd.n3192 gnd.n3191 585
R9835 gnd.n3191 gnd.n3189 585
R9836 gnd.n3283 gnd.n3282 585
R9837 gnd.n3798 gnd.n3282 585
R9838 gnd.n3285 gnd.n3284 585
R9839 gnd.n3286 gnd.n3285 585
R9840 gnd.n3296 gnd.n3272 585
R9841 gnd.n3804 gnd.n3272 585
R9842 gnd.n3298 gnd.n3297 585
R9843 gnd.n3299 gnd.n3298 585
R9844 gnd.n3295 gnd.n3294 585
R9845 gnd.n3295 gnd.n3262 585
R9846 gnd.n3293 gnd.n3260 585
R9847 gnd.n3812 gnd.n3260 585
R9848 gnd.n3249 gnd.n3247 585
R9849 gnd.n3774 gnd.n3249 585
R9850 gnd.n3820 gnd.n3819 585
R9851 gnd.n3819 gnd.n3818 585
R9852 gnd.n3248 gnd.n3246 585
R9853 gnd.n3313 gnd.n3248 585
R9854 gnd.n3745 gnd.n3312 585
R9855 gnd.n3764 gnd.n3312 585
R9856 gnd.n3747 gnd.n3746 585
R9857 gnd.n3748 gnd.n3747 585
R9858 gnd.n3322 gnd.n3321 585
R9859 gnd.n3328 gnd.n3321 585
R9860 gnd.n3740 gnd.n3739 585
R9861 gnd.n3739 gnd.n3738 585
R9862 gnd.n3325 gnd.n3324 585
R9863 gnd.n3336 gnd.n3325 585
R9864 gnd.n3625 gnd.n3344 585
R9865 gnd.n3717 gnd.n3344 585
R9866 gnd.n3627 gnd.n3626 585
R9867 gnd.n3626 gnd.n3342 585
R9868 gnd.n3628 gnd.n3355 585
R9869 gnd.n3707 gnd.n3355 585
R9870 gnd.n3630 gnd.n3629 585
R9871 gnd.n3630 gnd.n3362 585
R9872 gnd.n3632 gnd.n3631 585
R9873 gnd.n3631 gnd.n3361 585
R9874 gnd.n3633 gnd.n3372 585
R9875 gnd.n3687 gnd.n3372 585
R9876 gnd.n3635 gnd.n3634 585
R9877 gnd.n3634 gnd.n3370 585
R9878 gnd.n3636 gnd.n3381 585
R9879 gnd.n3676 gnd.n3381 585
R9880 gnd.n3638 gnd.n3637 585
R9881 gnd.n3638 gnd.n3387 585
R9882 gnd.n3640 gnd.n3639 585
R9883 gnd.n3639 gnd.n3386 585
R9884 gnd.n3641 gnd.n3402 585
R9885 gnd.n3655 gnd.n3402 585
R9886 gnd.n3642 gnd.n3455 585
R9887 gnd.n3455 gnd.n3394 585
R9888 gnd.n3644 gnd.n3643 585
R9889 gnd.n3645 gnd.n3644 585
R9890 gnd.n3456 gnd.n3454 585
R9891 gnd.n3454 gnd.n3453 585
R9892 gnd.n3609 gnd.n3608 585
R9893 gnd.n3608 gnd.n3607 585
R9894 gnd.n3459 gnd.n3458 585
R9895 gnd.n3460 gnd.n3459 585
R9896 gnd.n3598 gnd.n3597 585
R9897 gnd.n3599 gnd.n3598 585
R9898 gnd.n3468 gnd.n3467 585
R9899 gnd.n3467 gnd.n3466 585
R9900 gnd.n3593 gnd.n3592 585
R9901 gnd.n3592 gnd.n3591 585
R9902 gnd.n3471 gnd.n3470 585
R9903 gnd.n3582 gnd.n3471 585
R9904 gnd.n3581 gnd.n3580 585
R9905 gnd.n3583 gnd.n3581 585
R9906 gnd.n3479 gnd.n3478 585
R9907 gnd.n3478 gnd.n3477 585
R9908 gnd.n7268 gnd.n7267 585
R9909 gnd.n7269 gnd.n7268 585
R9910 gnd.n158 gnd.n157 585
R9911 gnd.n7262 gnd.n158 585
R9912 gnd.n7277 gnd.n7276 585
R9913 gnd.n7276 gnd.n7275 585
R9914 gnd.n7278 gnd.n153 585
R9915 gnd.n6955 gnd.n153 585
R9916 gnd.n7280 gnd.n7279 585
R9917 gnd.n7281 gnd.n7280 585
R9918 gnd.n137 gnd.n136 585
R9919 gnd.n6961 gnd.n137 585
R9920 gnd.n7289 gnd.n7288 585
R9921 gnd.n7288 gnd.n7287 585
R9922 gnd.n7290 gnd.n132 585
R9923 gnd.n6967 gnd.n132 585
R9924 gnd.n7292 gnd.n7291 585
R9925 gnd.n7293 gnd.n7292 585
R9926 gnd.n116 gnd.n115 585
R9927 gnd.n6973 gnd.n116 585
R9928 gnd.n7301 gnd.n7300 585
R9929 gnd.n7300 gnd.n7299 585
R9930 gnd.n7302 gnd.n111 585
R9931 gnd.n6979 gnd.n111 585
R9932 gnd.n7304 gnd.n7303 585
R9933 gnd.n7305 gnd.n7304 585
R9934 gnd.n97 gnd.n96 585
R9935 gnd.n6985 gnd.n97 585
R9936 gnd.n7313 gnd.n7312 585
R9937 gnd.n7312 gnd.n7311 585
R9938 gnd.n7314 gnd.n91 585
R9939 gnd.n6991 gnd.n91 585
R9940 gnd.n7316 gnd.n7315 585
R9941 gnd.n7317 gnd.n7316 585
R9942 gnd.n92 gnd.n90 585
R9943 gnd.n6997 gnd.n90 585
R9944 gnd.n6926 gnd.n6925 585
R9945 gnd.n6925 gnd.n265 585
R9946 gnd.n6924 gnd.n72 585
R9947 gnd.n7325 gnd.n72 585
R9948 gnd.n6923 gnd.n6922 585
R9949 gnd.n6922 gnd.n6921 585
R9950 gnd.n277 gnd.n275 585
R9951 gnd.n6907 gnd.n277 585
R9952 gnd.n6914 gnd.n6913 585
R9953 gnd.n6913 gnd.n6912 585
R9954 gnd.n283 gnd.n282 585
R9955 gnd.n6902 gnd.n283 585
R9956 gnd.n6884 gnd.n6883 585
R9957 gnd.n6885 gnd.n6884 585
R9958 gnd.n298 gnd.n297 585
R9959 gnd.n6877 gnd.n297 585
R9960 gnd.n6871 gnd.n6870 585
R9961 gnd.n6872 gnd.n6871 585
R9962 gnd.n309 gnd.n308 585
R9963 gnd.n6865 gnd.n308 585
R9964 gnd.n6833 gnd.n6832 585
R9965 gnd.n6832 gnd.n6831 585
R9966 gnd.n6834 gnd.n323 585
R9967 gnd.n6849 gnd.n323 585
R9968 gnd.n6835 gnd.n335 585
R9969 gnd.n6826 gnd.n335 585
R9970 gnd.n6837 gnd.n6836 585
R9971 gnd.n6838 gnd.n6837 585
R9972 gnd.n336 gnd.n334 585
R9973 gnd.n6822 gnd.n334 585
R9974 gnd.n6798 gnd.n6797 585
R9975 gnd.n6797 gnd.n6796 585
R9976 gnd.n6799 gnd.n352 585
R9977 gnd.n6813 gnd.n352 585
R9978 gnd.n6800 gnd.n363 585
R9979 gnd.n6790 gnd.n363 585
R9980 gnd.n6802 gnd.n6801 585
R9981 gnd.n6803 gnd.n6802 585
R9982 gnd.n364 gnd.n362 585
R9983 gnd.n6753 gnd.n362 585
R9984 gnd.n405 gnd.n404 585
R9985 gnd.n404 gnd.n374 585
R9986 gnd.n403 gnd.n385 585
R9987 gnd.n6744 gnd.n385 585
R9988 gnd.n398 gnd.n396 585
R9989 gnd.n6727 gnd.n396 585
R9990 gnd.n6733 gnd.n6732 585
R9991 gnd.n6734 gnd.n6733 585
R9992 gnd.n397 gnd.n395 585
R9993 gnd.n6715 gnd.n395 585
R9994 gnd.n6491 gnd.n6490 585
R9995 gnd.n6569 gnd.n6492 585
R9996 gnd.n6568 gnd.n6493 585
R9997 gnd.n6500 gnd.n6494 585
R9998 gnd.n6561 gnd.n6501 585
R9999 gnd.n6560 gnd.n6502 585
R10000 gnd.n6504 gnd.n6503 585
R10001 gnd.n6553 gnd.n6512 585
R10002 gnd.n6552 gnd.n6513 585
R10003 gnd.n6520 gnd.n6514 585
R10004 gnd.n6545 gnd.n6521 585
R10005 gnd.n6544 gnd.n6522 585
R10006 gnd.n6524 gnd.n6523 585
R10007 gnd.n6537 gnd.n6532 585
R10008 gnd.n6536 gnd.n6533 585
R10009 gnd.n493 gnd.n452 585
R10010 gnd.n6699 gnd.n453 585
R10011 gnd.n6698 gnd.n6695 585
R10012 gnd.n454 gnd.n420 585
R10013 gnd.n6693 gnd.n420 585
R10014 gnd.n7256 gnd.n7255 585
R10015 gnd.n183 gnd.n182 585
R10016 gnd.n240 gnd.n239 585
R10017 gnd.n192 gnd.n191 585
R10018 gnd.n235 gnd.n234 585
R10019 gnd.n233 gnd.n232 585
R10020 gnd.n231 gnd.n230 585
R10021 gnd.n224 gnd.n194 585
R10022 gnd.n226 gnd.n225 585
R10023 gnd.n223 gnd.n222 585
R10024 gnd.n221 gnd.n220 585
R10025 gnd.n214 gnd.n196 585
R10026 gnd.n216 gnd.n215 585
R10027 gnd.n213 gnd.n212 585
R10028 gnd.n211 gnd.n210 585
R10029 gnd.n204 gnd.n198 585
R10030 gnd.n206 gnd.n205 585
R10031 gnd.n203 gnd.n202 585
R10032 gnd.n201 gnd.n172 585
R10033 gnd.n7253 gnd.n172 585
R10034 gnd.n7259 gnd.n170 585
R10035 gnd.n7269 gnd.n170 585
R10036 gnd.n7261 gnd.n7260 585
R10037 gnd.n7262 gnd.n7261 585
R10038 gnd.n177 gnd.n161 585
R10039 gnd.n7275 gnd.n161 585
R10040 gnd.n6957 gnd.n6956 585
R10041 gnd.n6956 gnd.n6955 585
R10042 gnd.n6958 gnd.n151 585
R10043 gnd.n7281 gnd.n151 585
R10044 gnd.n6960 gnd.n6959 585
R10045 gnd.n6961 gnd.n6960 585
R10046 gnd.n6945 gnd.n140 585
R10047 gnd.n7287 gnd.n140 585
R10048 gnd.n6969 gnd.n6968 585
R10049 gnd.n6968 gnd.n6967 585
R10050 gnd.n6970 gnd.n130 585
R10051 gnd.n7293 gnd.n130 585
R10052 gnd.n6972 gnd.n6971 585
R10053 gnd.n6973 gnd.n6972 585
R10054 gnd.n6937 gnd.n119 585
R10055 gnd.n7299 gnd.n119 585
R10056 gnd.n6981 gnd.n6980 585
R10057 gnd.n6980 gnd.n6979 585
R10058 gnd.n6982 gnd.n110 585
R10059 gnd.n7305 gnd.n110 585
R10060 gnd.n6984 gnd.n6983 585
R10061 gnd.n6985 gnd.n6984 585
R10062 gnd.n271 gnd.n100 585
R10063 gnd.n7311 gnd.n100 585
R10064 gnd.n6993 gnd.n6992 585
R10065 gnd.n6992 gnd.n6991 585
R10066 gnd.n6994 gnd.n88 585
R10067 gnd.n7317 gnd.n88 585
R10068 gnd.n6996 gnd.n6995 585
R10069 gnd.n6997 gnd.n6996 585
R10070 gnd.n68 gnd.n67 585
R10071 gnd.n265 gnd.n68 585
R10072 gnd.n7327 gnd.n7326 585
R10073 gnd.n7326 gnd.n7325 585
R10074 gnd.n7328 gnd.n66 585
R10075 gnd.n6921 gnd.n66 585
R10076 gnd.n6906 gnd.n64 585
R10077 gnd.n6907 gnd.n6906 585
R10078 gnd.n6855 gnd.n285 585
R10079 gnd.n6912 gnd.n285 585
R10080 gnd.n6857 gnd.n290 585
R10081 gnd.n6902 gnd.n290 585
R10082 gnd.n6858 gnd.n296 585
R10083 gnd.n6885 gnd.n296 585
R10084 gnd.n6859 gnd.n303 585
R10085 gnd.n6877 gnd.n303 585
R10086 gnd.n316 gnd.n307 585
R10087 gnd.n6872 gnd.n307 585
R10088 gnd.n6864 gnd.n6863 585
R10089 gnd.n6865 gnd.n6864 585
R10090 gnd.n315 gnd.n314 585
R10091 gnd.n6831 gnd.n314 585
R10092 gnd.n6851 gnd.n6850 585
R10093 gnd.n6850 gnd.n6849 585
R10094 gnd.n319 gnd.n318 585
R10095 gnd.n6826 gnd.n319 585
R10096 gnd.n345 gnd.n332 585
R10097 gnd.n6838 gnd.n332 585
R10098 gnd.n6821 gnd.n6820 585
R10099 gnd.n6822 gnd.n6821 585
R10100 gnd.n344 gnd.n343 585
R10101 gnd.n6796 gnd.n343 585
R10102 gnd.n6815 gnd.n6814 585
R10103 gnd.n6814 gnd.n6813 585
R10104 gnd.n348 gnd.n347 585
R10105 gnd.n6790 gnd.n348 585
R10106 gnd.n378 gnd.n361 585
R10107 gnd.n6803 gnd.n361 585
R10108 gnd.n6752 gnd.n6751 585
R10109 gnd.n6753 gnd.n6752 585
R10110 gnd.n377 gnd.n376 585
R10111 gnd.n376 gnd.n374 585
R10112 gnd.n6746 gnd.n6745 585
R10113 gnd.n6745 gnd.n6744 585
R10114 gnd.n381 gnd.n380 585
R10115 gnd.n6727 gnd.n381 585
R10116 gnd.n421 gnd.n394 585
R10117 gnd.n6734 gnd.n394 585
R10118 gnd.n6714 gnd.n6713 585
R10119 gnd.n6715 gnd.n6714 585
R10120 gnd.n4361 gnd.n4360 585
R10121 gnd.n4362 gnd.n4361 585
R10122 gnd.n3039 gnd.n3037 585
R10123 gnd.n3037 gnd.n3033 585
R10124 gnd.n3021 gnd.n3020 585
R10125 gnd.n3025 gnd.n3021 585
R10126 gnd.n4372 gnd.n4371 585
R10127 gnd.n4371 gnd.n4370 585
R10128 gnd.n4373 gnd.n3013 585
R10129 gnd.n4243 gnd.n3013 585
R10130 gnd.n4375 gnd.n4374 585
R10131 gnd.n4376 gnd.n4375 585
R10132 gnd.n3014 gnd.n3012 585
R10133 gnd.n3012 gnd.n3008 585
R10134 gnd.n2995 gnd.n2994 585
R10135 gnd.n2999 gnd.n2995 585
R10136 gnd.n4386 gnd.n4385 585
R10137 gnd.n4385 gnd.n4384 585
R10138 gnd.n4387 gnd.n2987 585
R10139 gnd.n4254 gnd.n2987 585
R10140 gnd.n4389 gnd.n4388 585
R10141 gnd.n4390 gnd.n4389 585
R10142 gnd.n2988 gnd.n2986 585
R10143 gnd.n2986 gnd.n2983 585
R10144 gnd.n2970 gnd.n2969 585
R10145 gnd.n2974 gnd.n2970 585
R10146 gnd.n4400 gnd.n4399 585
R10147 gnd.n4399 gnd.n4398 585
R10148 gnd.n4401 gnd.n2964 585
R10149 gnd.n3929 gnd.n2964 585
R10150 gnd.n4403 gnd.n4402 585
R10151 gnd.n4404 gnd.n4403 585
R10152 gnd.n2965 gnd.n2963 585
R10153 gnd.n2963 gnd.n2960 585
R10154 gnd.n3948 gnd.n3947 585
R10155 gnd.n3949 gnd.n3948 585
R10156 gnd.n3132 gnd.n3131 585
R10157 gnd.n3131 gnd.n2950 585
R10158 gnd.n3942 gnd.n3941 585
R10159 gnd.n3941 gnd.n3940 585
R10160 gnd.n3135 gnd.n3134 585
R10161 gnd.n3144 gnd.n3135 585
R10162 gnd.n3891 gnd.n3157 585
R10163 gnd.n3157 gnd.n3143 585
R10164 gnd.n3893 gnd.n3892 585
R10165 gnd.n3894 gnd.n3893 585
R10166 gnd.n3158 gnd.n3156 585
R10167 gnd.n3165 gnd.n3156 585
R10168 gnd.n3886 gnd.n3885 585
R10169 gnd.n3885 gnd.n3884 585
R10170 gnd.n3161 gnd.n3160 585
R10171 gnd.n3865 gnd.n3161 585
R10172 gnd.n3851 gnd.n3184 585
R10173 gnd.n3184 gnd.n3174 585
R10174 gnd.n3853 gnd.n3852 585
R10175 gnd.n3854 gnd.n3853 585
R10176 gnd.n3185 gnd.n3183 585
R10177 gnd.n3842 gnd.n3183 585
R10178 gnd.n3846 gnd.n3845 585
R10179 gnd.n3845 gnd.n3844 585
R10180 gnd.n3188 gnd.n3187 585
R10181 gnd.n3797 gnd.n3188 585
R10182 gnd.n3290 gnd.n3289 585
R10183 gnd.n3291 gnd.n3290 585
R10184 gnd.n3270 gnd.n3269 585
R10185 gnd.n3273 gnd.n3270 585
R10186 gnd.n3807 gnd.n3806 585
R10187 gnd.n3806 gnd.n3805 585
R10188 gnd.n3808 gnd.n3264 585
R10189 gnd.n3300 gnd.n3264 585
R10190 gnd.n3810 gnd.n3809 585
R10191 gnd.n3811 gnd.n3810 585
R10192 gnd.n3265 gnd.n3263 585
R10193 gnd.n3775 gnd.n3263 585
R10194 gnd.n3759 gnd.n3758 585
R10195 gnd.n3758 gnd.n3251 585
R10196 gnd.n3760 gnd.n3315 585
R10197 gnd.n3315 gnd.n3250 585
R10198 gnd.n3762 gnd.n3761 585
R10199 gnd.n3763 gnd.n3762 585
R10200 gnd.n3316 gnd.n3314 585
R10201 gnd.n3314 gnd.n3311 585
R10202 gnd.n3751 gnd.n3750 585
R10203 gnd.n3750 gnd.n3749 585
R10204 gnd.n3319 gnd.n3318 585
R10205 gnd.n3326 gnd.n3319 585
R10206 gnd.n3725 gnd.n3724 585
R10207 gnd.n3726 gnd.n3725 585
R10208 gnd.n3338 gnd.n3337 585
R10209 gnd.n3345 gnd.n3337 585
R10210 gnd.n3720 gnd.n3719 585
R10211 gnd.n3719 gnd.n3718 585
R10212 gnd.n3341 gnd.n3340 585
R10213 gnd.n3708 gnd.n3341 585
R10214 gnd.n3695 gnd.n3365 585
R10215 gnd.n3365 gnd.n3364 585
R10216 gnd.n3697 gnd.n3696 585
R10217 gnd.n3698 gnd.n3697 585
R10218 gnd.n3366 gnd.n3363 585
R10219 gnd.n3373 gnd.n3363 585
R10220 gnd.n3690 gnd.n3689 585
R10221 gnd.n3689 gnd.n3688 585
R10222 gnd.n3369 gnd.n3368 585
R10223 gnd.n3677 gnd.n3369 585
R10224 gnd.n3664 gnd.n3390 585
R10225 gnd.n3390 gnd.n3389 585
R10226 gnd.n3666 gnd.n3665 585
R10227 gnd.n3667 gnd.n3666 585
R10228 gnd.n3660 gnd.n3388 585
R10229 gnd.n3659 gnd.n3658 585
R10230 gnd.n3393 gnd.n3392 585
R10231 gnd.n3656 gnd.n3393 585
R10232 gnd.n3415 gnd.n3414 585
R10233 gnd.n3418 gnd.n3417 585
R10234 gnd.n3416 gnd.n3411 585
R10235 gnd.n3423 gnd.n3422 585
R10236 gnd.n3425 gnd.n3424 585
R10237 gnd.n3428 gnd.n3427 585
R10238 gnd.n3426 gnd.n3409 585
R10239 gnd.n3433 gnd.n3432 585
R10240 gnd.n3435 gnd.n3434 585
R10241 gnd.n3438 gnd.n3437 585
R10242 gnd.n3436 gnd.n3407 585
R10243 gnd.n3443 gnd.n3442 585
R10244 gnd.n3447 gnd.n3444 585
R10245 gnd.n3448 gnd.n3385 585
R10246 gnd.n4330 gnd.n4329 585
R10247 gnd.n4332 gnd.n3068 585
R10248 gnd.n4334 gnd.n4333 585
R10249 gnd.n4335 gnd.n3061 585
R10250 gnd.n4337 gnd.n4336 585
R10251 gnd.n4339 gnd.n3059 585
R10252 gnd.n4341 gnd.n4340 585
R10253 gnd.n4342 gnd.n3054 585
R10254 gnd.n4344 gnd.n4343 585
R10255 gnd.n4346 gnd.n3052 585
R10256 gnd.n4348 gnd.n4347 585
R10257 gnd.n4349 gnd.n3047 585
R10258 gnd.n4351 gnd.n4350 585
R10259 gnd.n4353 gnd.n3045 585
R10260 gnd.n4355 gnd.n4354 585
R10261 gnd.n4356 gnd.n3043 585
R10262 gnd.n4357 gnd.n3038 585
R10263 gnd.n3038 gnd.n3036 585
R10264 gnd.n4237 gnd.n3035 585
R10265 gnd.n4362 gnd.n3035 585
R10266 gnd.n4239 gnd.n4238 585
R10267 gnd.n4239 gnd.n3033 585
R10268 gnd.n4241 gnd.n4240 585
R10269 gnd.n4240 gnd.n3025 585
R10270 gnd.n4242 gnd.n3023 585
R10271 gnd.n4370 gnd.n3023 585
R10272 gnd.n4245 gnd.n4244 585
R10273 gnd.n4244 gnd.n4243 585
R10274 gnd.n4246 gnd.n3010 585
R10275 gnd.n4376 gnd.n3010 585
R10276 gnd.n4248 gnd.n4247 585
R10277 gnd.n4248 gnd.n3008 585
R10278 gnd.n4250 gnd.n4249 585
R10279 gnd.n4249 gnd.n2999 585
R10280 gnd.n4251 gnd.n2997 585
R10281 gnd.n4384 gnd.n2997 585
R10282 gnd.n4253 gnd.n4252 585
R10283 gnd.n4254 gnd.n4253 585
R10284 gnd.n3966 gnd.n2985 585
R10285 gnd.n4390 gnd.n2985 585
R10286 gnd.n3965 gnd.n3964 585
R10287 gnd.n3964 gnd.n2983 585
R10288 gnd.n3963 gnd.n3961 585
R10289 gnd.n3963 gnd.n2974 585
R10290 gnd.n3959 gnd.n2972 585
R10291 gnd.n4398 gnd.n2972 585
R10292 gnd.n3928 gnd.n3125 585
R10293 gnd.n3929 gnd.n3928 585
R10294 gnd.n3953 gnd.n2962 585
R10295 gnd.n4404 gnd.n2962 585
R10296 gnd.n3952 gnd.n3951 585
R10297 gnd.n3951 gnd.n2960 585
R10298 gnd.n3950 gnd.n3127 585
R10299 gnd.n3950 gnd.n3949 585
R10300 gnd.n3900 gnd.n3129 585
R10301 gnd.n3129 gnd.n2950 585
R10302 gnd.n3901 gnd.n3137 585
R10303 gnd.n3940 gnd.n3137 585
R10304 gnd.n3898 gnd.n3897 585
R10305 gnd.n3897 gnd.n3144 585
R10306 gnd.n3896 gnd.n3151 585
R10307 gnd.n3896 gnd.n3143 585
R10308 gnd.n3895 gnd.n3153 585
R10309 gnd.n3895 gnd.n3894 585
R10310 gnd.n3874 gnd.n3152 585
R10311 gnd.n3165 gnd.n3152 585
R10312 gnd.n3873 gnd.n3163 585
R10313 gnd.n3884 gnd.n3163 585
R10314 gnd.n3864 gnd.n3170 585
R10315 gnd.n3865 gnd.n3864 585
R10316 gnd.n3863 gnd.n3862 585
R10317 gnd.n3863 gnd.n3174 585
R10318 gnd.n3861 gnd.n3176 585
R10319 gnd.n3854 gnd.n3176 585
R10320 gnd.n3841 gnd.n3177 585
R10321 gnd.n3842 gnd.n3841 585
R10322 gnd.n3794 gnd.n3190 585
R10323 gnd.n3844 gnd.n3190 585
R10324 gnd.n3796 gnd.n3795 585
R10325 gnd.n3797 gnd.n3796 585
R10326 gnd.n3789 gnd.n3292 585
R10327 gnd.n3292 gnd.n3291 585
R10328 gnd.n3787 gnd.n3786 585
R10329 gnd.n3786 gnd.n3273 585
R10330 gnd.n3784 gnd.n3271 585
R10331 gnd.n3805 gnd.n3271 585
R10332 gnd.n3302 gnd.n3301 585
R10333 gnd.n3301 gnd.n3300 585
R10334 gnd.n3778 gnd.n3261 585
R10335 gnd.n3811 gnd.n3261 585
R10336 gnd.n3777 gnd.n3776 585
R10337 gnd.n3776 gnd.n3775 585
R10338 gnd.n3773 gnd.n3304 585
R10339 gnd.n3773 gnd.n3251 585
R10340 gnd.n3772 gnd.n3771 585
R10341 gnd.n3772 gnd.n3250 585
R10342 gnd.n3307 gnd.n3306 585
R10343 gnd.n3763 gnd.n3306 585
R10344 gnd.n3731 gnd.n3730 585
R10345 gnd.n3730 gnd.n3311 585
R10346 gnd.n3732 gnd.n3320 585
R10347 gnd.n3749 gnd.n3320 585
R10348 gnd.n3729 gnd.n3728 585
R10349 gnd.n3728 gnd.n3326 585
R10350 gnd.n3727 gnd.n3334 585
R10351 gnd.n3727 gnd.n3726 585
R10352 gnd.n3712 gnd.n3335 585
R10353 gnd.n3345 gnd.n3335 585
R10354 gnd.n3711 gnd.n3343 585
R10355 gnd.n3718 gnd.n3343 585
R10356 gnd.n3710 gnd.n3709 585
R10357 gnd.n3709 gnd.n3708 585
R10358 gnd.n3354 gnd.n3351 585
R10359 gnd.n3364 gnd.n3354 585
R10360 gnd.n3700 gnd.n3699 585
R10361 gnd.n3699 gnd.n3698 585
R10362 gnd.n3360 gnd.n3359 585
R10363 gnd.n3373 gnd.n3360 585
R10364 gnd.n3680 gnd.n3371 585
R10365 gnd.n3688 gnd.n3371 585
R10366 gnd.n3679 gnd.n3678 585
R10367 gnd.n3678 gnd.n3677 585
R10368 gnd.n3380 gnd.n3378 585
R10369 gnd.n3389 gnd.n3380 585
R10370 gnd.n3669 gnd.n3668 585
R10371 gnd.n3668 gnd.n3667 585
R10372 gnd.n6281 gnd.n6280 585
R10373 gnd.n6282 gnd.n6281 585
R10374 gnd.n6192 gnd.n694 585
R10375 gnd.n700 gnd.n694 585
R10376 gnd.n6191 gnd.n6190 585
R10377 gnd.n6190 gnd.n6189 585
R10378 gnd.n697 gnd.n696 585
R10379 gnd.n6002 gnd.n697 585
R10380 gnd.n6157 gnd.n6156 585
R10381 gnd.n6157 gnd.n709 585
R10382 gnd.n6159 gnd.n6158 585
R10383 gnd.n6158 gnd.n707 585
R10384 gnd.n6160 gnd.n721 585
R10385 gnd.n6009 gnd.n721 585
R10386 gnd.n6162 gnd.n6161 585
R10387 gnd.n6163 gnd.n6162 585
R10388 gnd.n6155 gnd.n720 585
R10389 gnd.n6150 gnd.n720 585
R10390 gnd.n6154 gnd.n6153 585
R10391 gnd.n6153 gnd.n6152 585
R10392 gnd.n723 gnd.n722 585
R10393 gnd.n6140 gnd.n723 585
R10394 gnd.n6127 gnd.n746 585
R10395 gnd.n746 gnd.n733 585
R10396 gnd.n6129 gnd.n6128 585
R10397 gnd.n6130 gnd.n6129 585
R10398 gnd.n6126 gnd.n745 585
R10399 gnd.n745 gnd.n741 585
R10400 gnd.n6125 gnd.n6124 585
R10401 gnd.n6124 gnd.n6123 585
R10402 gnd.n748 gnd.n747 585
R10403 gnd.n5985 gnd.n748 585
R10404 gnd.n6112 gnd.n6111 585
R10405 gnd.n6113 gnd.n6112 585
R10406 gnd.n6110 gnd.n759 585
R10407 gnd.n759 gnd.n756 585
R10408 gnd.n6109 gnd.n6108 585
R10409 gnd.n6108 gnd.n6107 585
R10410 gnd.n761 gnd.n760 585
R10411 gnd.n5977 gnd.n761 585
R10412 gnd.n6095 gnd.n6094 585
R10413 gnd.n6096 gnd.n6095 585
R10414 gnd.n6093 gnd.n774 585
R10415 gnd.n774 gnd.n771 585
R10416 gnd.n6092 gnd.n6091 585
R10417 gnd.n6091 gnd.n6090 585
R10418 gnd.n776 gnd.n775 585
R10419 gnd.n788 gnd.n776 585
R10420 gnd.n6064 gnd.n6063 585
R10421 gnd.n6063 gnd.n785 585
R10422 gnd.n6065 gnd.n799 585
R10423 gnd.n6051 gnd.n799 585
R10424 gnd.n6067 gnd.n6066 585
R10425 gnd.n6068 gnd.n6067 585
R10426 gnd.n6062 gnd.n798 585
R10427 gnd.n6057 gnd.n798 585
R10428 gnd.n6061 gnd.n6060 585
R10429 gnd.n6060 gnd.n6059 585
R10430 gnd.n801 gnd.n800 585
R10431 gnd.n813 gnd.n801 585
R10432 gnd.n5939 gnd.n5938 585
R10433 gnd.n5938 gnd.n5937 585
R10434 gnd.n5940 gnd.n822 585
R10435 gnd.n5916 gnd.n822 585
R10436 gnd.n5942 gnd.n5941 585
R10437 gnd.n5943 gnd.n5942 585
R10438 gnd.n823 gnd.n821 585
R10439 gnd.n5922 gnd.n821 585
R10440 gnd.n5905 gnd.n842 585
R10441 gnd.n842 gnd.n841 585
R10442 gnd.n5907 gnd.n5906 585
R10443 gnd.n5908 gnd.n5907 585
R10444 gnd.n5904 gnd.n840 585
R10445 gnd.n848 gnd.n840 585
R10446 gnd.n5903 gnd.n5902 585
R10447 gnd.n5902 gnd.n5901 585
R10448 gnd.n844 gnd.n843 585
R10449 gnd.n5818 gnd.n844 585
R10450 gnd.n5889 gnd.n5888 585
R10451 gnd.n5890 gnd.n5889 585
R10452 gnd.n5887 gnd.n859 585
R10453 gnd.n859 gnd.n855 585
R10454 gnd.n5886 gnd.n5885 585
R10455 gnd.n5885 gnd.n5884 585
R10456 gnd.n861 gnd.n860 585
R10457 gnd.n5851 gnd.n861 585
R10458 gnd.n5864 gnd.n5863 585
R10459 gnd.n5865 gnd.n5864 585
R10460 gnd.n5862 gnd.n873 585
R10461 gnd.n5857 gnd.n873 585
R10462 gnd.n5861 gnd.n5860 585
R10463 gnd.n5860 gnd.n5859 585
R10464 gnd.n875 gnd.n874 585
R10465 gnd.n885 gnd.n875 585
R10466 gnd.n5784 gnd.n5783 585
R10467 gnd.n5785 gnd.n5784 585
R10468 gnd.n908 gnd.n907 585
R10469 gnd.n908 gnd.n894 585
R10470 gnd.n5793 gnd.n5792 585
R10471 gnd.n5792 gnd.n5791 585
R10472 gnd.n5794 gnd.n905 585
R10473 gnd.n910 gnd.n905 585
R10474 gnd.n5796 gnd.n5795 585
R10475 gnd.n5797 gnd.n5796 585
R10476 gnd.n906 gnd.n904 585
R10477 gnd.n5739 gnd.n904 585
R10478 gnd.n5742 gnd.n5741 585
R10479 gnd.n5743 gnd.n5742 585
R10480 gnd.n940 gnd.n939 585
R10481 gnd.n940 gnd.n927 585
R10482 gnd.n5751 gnd.n5750 585
R10483 gnd.n5750 gnd.n5749 585
R10484 gnd.n5752 gnd.n937 585
R10485 gnd.n942 gnd.n937 585
R10486 gnd.n5754 gnd.n5753 585
R10487 gnd.n5755 gnd.n5754 585
R10488 gnd.n938 gnd.n936 585
R10489 gnd.n5683 gnd.n936 585
R10490 gnd.n977 gnd.n976 585
R10491 gnd.n980 gnd.n976 585
R10492 gnd.n5706 gnd.n978 585
R10493 gnd.n5706 gnd.n5705 585
R10494 gnd.n5707 gnd.n975 585
R10495 gnd.n5707 gnd.n960 585
R10496 gnd.n5709 gnd.n5708 585
R10497 gnd.n5708 gnd.n959 585
R10498 gnd.n5710 gnd.n973 585
R10499 gnd.t86 gnd.n973 585
R10500 gnd.n5712 gnd.n5711 585
R10501 gnd.n5713 gnd.n5712 585
R10502 gnd.n974 gnd.n972 585
R10503 gnd.n972 gnd.n968 585
R10504 gnd.n5673 gnd.n5672 585
R10505 gnd.n5674 gnd.n5673 585
R10506 gnd.n5671 gnd.n993 585
R10507 gnd.n999 gnd.n993 585
R10508 gnd.n5670 gnd.n5669 585
R10509 gnd.n5669 gnd.n5668 585
R10510 gnd.n995 gnd.n994 585
R10511 gnd.n5597 gnd.n995 585
R10512 gnd.n5657 gnd.n5656 585
R10513 gnd.n5658 gnd.n5657 585
R10514 gnd.n5654 gnd.n1008 585
R10515 gnd.n5653 gnd.n5652 585
R10516 gnd.n1030 gnd.n1029 585
R10517 gnd.n5650 gnd.n1030 585
R10518 gnd.n1091 gnd.n1090 585
R10519 gnd.n1093 gnd.n1092 585
R10520 gnd.n1095 gnd.n1094 585
R10521 gnd.n1097 gnd.n1096 585
R10522 gnd.n1099 gnd.n1098 585
R10523 gnd.n1101 gnd.n1100 585
R10524 gnd.n1103 gnd.n1102 585
R10525 gnd.n1105 gnd.n1104 585
R10526 gnd.n1107 gnd.n1106 585
R10527 gnd.n1109 gnd.n1108 585
R10528 gnd.n1111 gnd.n1110 585
R10529 gnd.n1113 gnd.n1112 585
R10530 gnd.n1115 gnd.n1114 585
R10531 gnd.n1117 gnd.n1116 585
R10532 gnd.n1119 gnd.n1118 585
R10533 gnd.n1121 gnd.n1120 585
R10534 gnd.n1123 gnd.n1122 585
R10535 gnd.n1125 gnd.n1124 585
R10536 gnd.n1127 gnd.n1126 585
R10537 gnd.n1129 gnd.n1128 585
R10538 gnd.n1131 gnd.n1130 585
R10539 gnd.n1133 gnd.n1132 585
R10540 gnd.n1135 gnd.n1134 585
R10541 gnd.n1137 gnd.n1136 585
R10542 gnd.n1139 gnd.n1138 585
R10543 gnd.n1141 gnd.n1140 585
R10544 gnd.n1143 gnd.n1142 585
R10545 gnd.n1145 gnd.n1144 585
R10546 gnd.n1147 gnd.n1146 585
R10547 gnd.n5526 gnd.n5525 585
R10548 gnd.n5528 gnd.n5527 585
R10549 gnd.n5530 gnd.n5529 585
R10550 gnd.n5532 gnd.n5531 585
R10551 gnd.n5535 gnd.n5534 585
R10552 gnd.n5537 gnd.n5536 585
R10553 gnd.n5539 gnd.n5538 585
R10554 gnd.n5541 gnd.n5540 585
R10555 gnd.n5543 gnd.n5542 585
R10556 gnd.n5545 gnd.n5544 585
R10557 gnd.n5547 gnd.n5546 585
R10558 gnd.n5549 gnd.n5548 585
R10559 gnd.n5551 gnd.n5550 585
R10560 gnd.n5553 gnd.n5552 585
R10561 gnd.n5555 gnd.n5554 585
R10562 gnd.n5557 gnd.n5556 585
R10563 gnd.n5559 gnd.n5558 585
R10564 gnd.n5561 gnd.n5560 585
R10565 gnd.n5563 gnd.n5562 585
R10566 gnd.n5565 gnd.n5564 585
R10567 gnd.n5567 gnd.n5566 585
R10568 gnd.n5569 gnd.n5568 585
R10569 gnd.n5571 gnd.n5570 585
R10570 gnd.n5573 gnd.n5572 585
R10571 gnd.n5575 gnd.n5574 585
R10572 gnd.n5577 gnd.n5576 585
R10573 gnd.n5579 gnd.n5578 585
R10574 gnd.n5581 gnd.n5580 585
R10575 gnd.n5583 gnd.n5582 585
R10576 gnd.n5585 gnd.n5584 585
R10577 gnd.n5587 gnd.n5586 585
R10578 gnd.n5589 gnd.n5588 585
R10579 gnd.n5591 gnd.n5590 585
R10580 gnd.n6285 gnd.n6284 585
R10581 gnd.n6287 gnd.n6286 585
R10582 gnd.n6289 gnd.n6288 585
R10583 gnd.n6291 gnd.n6290 585
R10584 gnd.n6293 gnd.n6292 585
R10585 gnd.n6295 gnd.n6294 585
R10586 gnd.n6297 gnd.n6296 585
R10587 gnd.n6299 gnd.n6298 585
R10588 gnd.n6301 gnd.n6300 585
R10589 gnd.n6303 gnd.n6302 585
R10590 gnd.n6305 gnd.n6304 585
R10591 gnd.n6307 gnd.n6306 585
R10592 gnd.n6309 gnd.n6308 585
R10593 gnd.n6311 gnd.n6310 585
R10594 gnd.n6313 gnd.n6312 585
R10595 gnd.n6315 gnd.n6314 585
R10596 gnd.n6317 gnd.n6316 585
R10597 gnd.n6319 gnd.n6318 585
R10598 gnd.n6321 gnd.n6320 585
R10599 gnd.n6323 gnd.n6322 585
R10600 gnd.n6325 gnd.n6324 585
R10601 gnd.n6327 gnd.n6326 585
R10602 gnd.n6329 gnd.n6328 585
R10603 gnd.n6331 gnd.n6330 585
R10604 gnd.n6333 gnd.n6332 585
R10605 gnd.n6335 gnd.n6334 585
R10606 gnd.n6337 gnd.n6336 585
R10607 gnd.n6339 gnd.n6338 585
R10608 gnd.n6341 gnd.n6340 585
R10609 gnd.n6344 gnd.n6343 585
R10610 gnd.n6346 gnd.n6345 585
R10611 gnd.n6348 gnd.n6347 585
R10612 gnd.n6350 gnd.n6349 585
R10613 gnd.n6214 gnd.n525 585
R10614 gnd.n6216 gnd.n6215 585
R10615 gnd.n6218 gnd.n6217 585
R10616 gnd.n6220 gnd.n6219 585
R10617 gnd.n6223 gnd.n6222 585
R10618 gnd.n6225 gnd.n6224 585
R10619 gnd.n6227 gnd.n6226 585
R10620 gnd.n6229 gnd.n6228 585
R10621 gnd.n6231 gnd.n6230 585
R10622 gnd.n6233 gnd.n6232 585
R10623 gnd.n6235 gnd.n6234 585
R10624 gnd.n6237 gnd.n6236 585
R10625 gnd.n6239 gnd.n6238 585
R10626 gnd.n6241 gnd.n6240 585
R10627 gnd.n6243 gnd.n6242 585
R10628 gnd.n6245 gnd.n6244 585
R10629 gnd.n6247 gnd.n6246 585
R10630 gnd.n6249 gnd.n6248 585
R10631 gnd.n6251 gnd.n6250 585
R10632 gnd.n6253 gnd.n6252 585
R10633 gnd.n6255 gnd.n6254 585
R10634 gnd.n6257 gnd.n6256 585
R10635 gnd.n6259 gnd.n6258 585
R10636 gnd.n6261 gnd.n6260 585
R10637 gnd.n6263 gnd.n6262 585
R10638 gnd.n6265 gnd.n6264 585
R10639 gnd.n6267 gnd.n6266 585
R10640 gnd.n6269 gnd.n6268 585
R10641 gnd.n6271 gnd.n6270 585
R10642 gnd.n6273 gnd.n6272 585
R10643 gnd.n6275 gnd.n6274 585
R10644 gnd.n6277 gnd.n6276 585
R10645 gnd.n6278 gnd.n695 585
R10646 gnd.n6283 gnd.n692 585
R10647 gnd.n6283 gnd.n6282 585
R10648 gnd.n5998 gnd.n693 585
R10649 gnd.n700 gnd.n693 585
R10650 gnd.n5999 gnd.n699 585
R10651 gnd.n6189 gnd.n699 585
R10652 gnd.n6003 gnd.n6000 585
R10653 gnd.n6003 gnd.n6002 585
R10654 gnd.n6005 gnd.n6004 585
R10655 gnd.n6004 gnd.n709 585
R10656 gnd.n6006 gnd.n5967 585
R10657 gnd.n5967 gnd.n707 585
R10658 gnd.n6008 gnd.n6007 585
R10659 gnd.n6009 gnd.n6008 585
R10660 gnd.n5997 gnd.n718 585
R10661 gnd.n6163 gnd.n718 585
R10662 gnd.n5996 gnd.n727 585
R10663 gnd.n6150 gnd.n727 585
R10664 gnd.n5995 gnd.n725 585
R10665 gnd.n6152 gnd.n725 585
R10666 gnd.n5994 gnd.n734 585
R10667 gnd.n6140 gnd.n734 585
R10668 gnd.n5993 gnd.n5992 585
R10669 gnd.n5992 gnd.n733 585
R10670 gnd.n5991 gnd.n743 585
R10671 gnd.n6130 gnd.n743 585
R10672 gnd.n5990 gnd.n5989 585
R10673 gnd.n5989 gnd.n741 585
R10674 gnd.n5988 gnd.n750 585
R10675 gnd.n6123 gnd.n750 585
R10676 gnd.n5987 gnd.n5986 585
R10677 gnd.n5986 gnd.n5985 585
R10678 gnd.n5983 gnd.n757 585
R10679 gnd.n6113 gnd.n757 585
R10680 gnd.n5982 gnd.n5981 585
R10681 gnd.n5981 gnd.n756 585
R10682 gnd.n5980 gnd.n762 585
R10683 gnd.n6107 gnd.n762 585
R10684 gnd.n5979 gnd.n5978 585
R10685 gnd.n5978 gnd.n5977 585
R10686 gnd.n5973 gnd.n773 585
R10687 gnd.n6096 gnd.n773 585
R10688 gnd.n5972 gnd.n5971 585
R10689 gnd.n5971 gnd.n771 585
R10690 gnd.n5970 gnd.n777 585
R10691 gnd.n6090 gnd.n777 585
R10692 gnd.n5969 gnd.n5968 585
R10693 gnd.n5968 gnd.n788 585
R10694 gnd.n807 gnd.n806 585
R10695 gnd.n807 gnd.n785 585
R10696 gnd.n6053 gnd.n6052 585
R10697 gnd.n6052 gnd.n6051 585
R10698 gnd.n6054 gnd.n796 585
R10699 gnd.n6068 gnd.n796 585
R10700 gnd.n6056 gnd.n6055 585
R10701 gnd.n6057 gnd.n6056 585
R10702 gnd.n805 gnd.n803 585
R10703 gnd.n6059 gnd.n803 585
R10704 gnd.n5913 gnd.n5912 585
R10705 gnd.n5912 gnd.n813 585
R10706 gnd.n5914 gnd.n825 585
R10707 gnd.n5937 gnd.n825 585
R10708 gnd.n5918 gnd.n5917 585
R10709 gnd.n5917 gnd.n5916 585
R10710 gnd.n5919 gnd.n820 585
R10711 gnd.n5943 gnd.n820 585
R10712 gnd.n5921 gnd.n5920 585
R10713 gnd.n5922 gnd.n5921 585
R10714 gnd.n5911 gnd.n833 585
R10715 gnd.n841 gnd.n833 585
R10716 gnd.n5910 gnd.n5909 585
R10717 gnd.n5909 gnd.n5908 585
R10718 gnd.n835 gnd.n834 585
R10719 gnd.n848 gnd.n835 585
R10720 gnd.n5815 gnd.n846 585
R10721 gnd.n5901 gnd.n846 585
R10722 gnd.n5817 gnd.n5816 585
R10723 gnd.n5818 gnd.n5817 585
R10724 gnd.n5814 gnd.n857 585
R10725 gnd.n5890 gnd.n857 585
R10726 gnd.n5813 gnd.n5812 585
R10727 gnd.n5812 gnd.n855 585
R10728 gnd.n878 gnd.n863 585
R10729 gnd.n5884 gnd.n863 585
R10730 gnd.n5853 gnd.n5852 585
R10731 gnd.n5852 gnd.n5851 585
R10732 gnd.n5854 gnd.n872 585
R10733 gnd.n5865 gnd.n872 585
R10734 gnd.n5856 gnd.n5855 585
R10735 gnd.n5857 gnd.n5856 585
R10736 gnd.n877 gnd.n876 585
R10737 gnd.n5859 gnd.n876 585
R10738 gnd.n915 gnd.n914 585
R10739 gnd.n915 gnd.n885 585
R10740 gnd.n5787 gnd.n5786 585
R10741 gnd.n5786 gnd.n5785 585
R10742 gnd.n5788 gnd.n912 585
R10743 gnd.n912 gnd.n894 585
R10744 gnd.n5790 gnd.n5789 585
R10745 gnd.n5791 gnd.n5790 585
R10746 gnd.n913 gnd.n911 585
R10747 gnd.n911 gnd.n910 585
R10748 gnd.n946 gnd.n902 585
R10749 gnd.n5797 gnd.n902 585
R10750 gnd.n948 gnd.n947 585
R10751 gnd.n5739 gnd.n948 585
R10752 gnd.n5745 gnd.n5744 585
R10753 gnd.n5744 gnd.n5743 585
R10754 gnd.n5746 gnd.n944 585
R10755 gnd.n944 gnd.n927 585
R10756 gnd.n5748 gnd.n5747 585
R10757 gnd.n5749 gnd.n5748 585
R10758 gnd.n945 gnd.n943 585
R10759 gnd.n943 gnd.n942 585
R10760 gnd.n5679 gnd.n934 585
R10761 gnd.n5755 gnd.n934 585
R10762 gnd.n5684 gnd.n5680 585
R10763 gnd.n5684 gnd.n5683 585
R10764 gnd.n5686 gnd.n5685 585
R10765 gnd.n5685 gnd.n980 585
R10766 gnd.n5687 gnd.n979 585
R10767 gnd.n5705 gnd.n979 585
R10768 gnd.n5689 gnd.n5688 585
R10769 gnd.n5688 gnd.n960 585
R10770 gnd.n5690 gnd.n988 585
R10771 gnd.n988 gnd.n959 585
R10772 gnd.n5692 gnd.n5691 585
R10773 gnd.t86 gnd.n5692 585
R10774 gnd.n5678 gnd.n970 585
R10775 gnd.n5713 gnd.n970 585
R10776 gnd.n5677 gnd.n5676 585
R10777 gnd.n5676 gnd.n968 585
R10778 gnd.n5675 gnd.n989 585
R10779 gnd.n5675 gnd.n5674 585
R10780 gnd.n5593 gnd.n990 585
R10781 gnd.n999 gnd.n990 585
R10782 gnd.n5594 gnd.n997 585
R10783 gnd.n5668 gnd.n997 585
R10784 gnd.n5596 gnd.n5595 585
R10785 gnd.n5597 gnd.n5596 585
R10786 gnd.n5592 gnd.n1006 585
R10787 gnd.n5658 gnd.n1006 585
R10788 gnd.n5455 gnd.n1217 585
R10789 gnd.n5190 gnd.n1217 585
R10790 gnd.n5457 gnd.n5456 585
R10791 gnd.n5458 gnd.n5457 585
R10792 gnd.n1218 gnd.n1216 585
R10793 gnd.n5026 gnd.n1216 585
R10794 gnd.n5358 gnd.n5357 585
R10795 gnd.n5357 gnd.n5356 585
R10796 gnd.n1221 gnd.n1220 585
R10797 gnd.n5346 gnd.n1221 585
R10798 gnd.n5015 gnd.n5014 585
R10799 gnd.n5016 gnd.n5015 585
R10800 gnd.n1287 gnd.n1286 585
R10801 gnd.n1286 gnd.n1284 585
R10802 gnd.n5010 gnd.n5009 585
R10803 gnd.n5009 gnd.n5008 585
R10804 gnd.n1290 gnd.n1289 585
R10805 gnd.n4996 gnd.n1290 585
R10806 gnd.n4981 gnd.n1314 585
R10807 gnd.n4967 gnd.n1314 585
R10808 gnd.n4983 gnd.n4982 585
R10809 gnd.n4984 gnd.n4983 585
R10810 gnd.n1315 gnd.n1313 585
R10811 gnd.n4961 gnd.n1313 585
R10812 gnd.n4976 gnd.n4975 585
R10813 gnd.n4975 gnd.n4974 585
R10814 gnd.n1318 gnd.n1317 585
R10815 gnd.n4940 gnd.n1318 585
R10816 gnd.n4928 gnd.n1347 585
R10817 gnd.n1347 gnd.n1334 585
R10818 gnd.n4930 gnd.n4929 585
R10819 gnd.n4931 gnd.n4930 585
R10820 gnd.n1348 gnd.n1346 585
R10821 gnd.n4881 gnd.n1346 585
R10822 gnd.n4896 gnd.n1391 585
R10823 gnd.n4896 gnd.n4895 585
R10824 gnd.n4899 gnd.n4898 585
R10825 gnd.n4900 gnd.n4899 585
R10826 gnd.n4897 gnd.n1390 585
R10827 gnd.n1390 gnd.n1385 585
R10828 gnd.n1374 gnd.n1373 585
R10829 gnd.n1378 gnd.n1373 585
R10830 gnd.n4910 gnd.n1375 585
R10831 gnd.n4910 gnd.n4909 585
R10832 gnd.n4913 gnd.n4912 585
R10833 gnd.n4914 gnd.n4913 585
R10834 gnd.n4911 gnd.n1357 585
R10835 gnd.n4864 gnd.n1357 585
R10836 gnd.n4922 gnd.n4921 585
R10837 gnd.n4921 gnd.n4920 585
R10838 gnd.n4923 gnd.n1356 585
R10839 gnd.n4853 gnd.n1356 585
R10840 gnd.n1426 gnd.n1355 585
R10841 gnd.n1426 gnd.n1415 585
R10842 gnd.n4826 gnd.n4825 585
R10843 gnd.n4827 gnd.n4826 585
R10844 gnd.n4824 gnd.n1425 585
R10845 gnd.n4812 gnd.n1425 585
R10846 gnd.n1431 gnd.n1427 585
R10847 gnd.n4793 gnd.n1431 585
R10848 gnd.n4820 gnd.n4819 585
R10849 gnd.n4819 gnd.n4818 585
R10850 gnd.n1430 gnd.n1429 585
R10851 gnd.n4799 gnd.n1430 585
R10852 gnd.n4773 gnd.n4772 585
R10853 gnd.n4774 gnd.n4773 585
R10854 gnd.n1463 gnd.n1462 585
R10855 gnd.n4759 gnd.n1462 585
R10856 gnd.n4768 gnd.n4767 585
R10857 gnd.n4767 gnd.n4766 585
R10858 gnd.n1466 gnd.n1465 585
R10859 gnd.n4750 gnd.n1466 585
R10860 gnd.n4746 gnd.n4745 585
R10861 gnd.n4747 gnd.n4746 585
R10862 gnd.n1485 gnd.n1484 585
R10863 gnd.n4722 gnd.n1484 585
R10864 gnd.n4741 gnd.n4740 585
R10865 gnd.n4740 gnd.n4739 585
R10866 gnd.n1488 gnd.n1487 585
R10867 gnd.n4728 gnd.n1488 585
R10868 gnd.n4711 gnd.n1511 585
R10869 gnd.n4519 gnd.n1511 585
R10870 gnd.n4713 gnd.n4712 585
R10871 gnd.n4714 gnd.n4713 585
R10872 gnd.n1512 gnd.n1510 585
R10873 gnd.n4584 gnd.n1510 585
R10874 gnd.n4706 gnd.n4705 585
R10875 gnd.n1515 gnd.n1514 585
R10876 gnd.n4702 gnd.n4701 585
R10877 gnd.n4703 gnd.n4702 585
R10878 gnd.n4700 gnd.n4453 585
R10879 gnd.n4699 gnd.n4698 585
R10880 gnd.n4697 gnd.n4696 585
R10881 gnd.n4695 gnd.n4694 585
R10882 gnd.n4693 gnd.n4692 585
R10883 gnd.n4691 gnd.n4690 585
R10884 gnd.n4689 gnd.n4688 585
R10885 gnd.n4687 gnd.n4686 585
R10886 gnd.n4685 gnd.n4684 585
R10887 gnd.n4683 gnd.n4682 585
R10888 gnd.n4681 gnd.n4680 585
R10889 gnd.n4679 gnd.n4678 585
R10890 gnd.n4677 gnd.n4676 585
R10891 gnd.n4675 gnd.n4674 585
R10892 gnd.n4673 gnd.n4672 585
R10893 gnd.n4670 gnd.n4669 585
R10894 gnd.n4668 gnd.n4667 585
R10895 gnd.n4666 gnd.n4665 585
R10896 gnd.n4664 gnd.n4663 585
R10897 gnd.n4662 gnd.n4661 585
R10898 gnd.n4660 gnd.n4659 585
R10899 gnd.n4658 gnd.n4657 585
R10900 gnd.n4656 gnd.n4655 585
R10901 gnd.n4654 gnd.n4653 585
R10902 gnd.n4652 gnd.n4651 585
R10903 gnd.n4650 gnd.n4649 585
R10904 gnd.n4648 gnd.n4647 585
R10905 gnd.n4646 gnd.n4645 585
R10906 gnd.n4644 gnd.n4643 585
R10907 gnd.n4642 gnd.n4641 585
R10908 gnd.n4640 gnd.n4639 585
R10909 gnd.n4638 gnd.n4637 585
R10910 gnd.n4636 gnd.n4635 585
R10911 gnd.n4634 gnd.n4633 585
R10912 gnd.n4632 gnd.n4631 585
R10913 gnd.n4630 gnd.n4629 585
R10914 gnd.n4628 gnd.n4627 585
R10915 gnd.n4626 gnd.n4625 585
R10916 gnd.n4624 gnd.n4623 585
R10917 gnd.n4622 gnd.n4621 585
R10918 gnd.n4620 gnd.n4619 585
R10919 gnd.n4618 gnd.n4617 585
R10920 gnd.n4616 gnd.n4615 585
R10921 gnd.n4614 gnd.n4613 585
R10922 gnd.n4612 gnd.n4611 585
R10923 gnd.n4610 gnd.n4609 585
R10924 gnd.n4608 gnd.n4607 585
R10925 gnd.n4606 gnd.n4605 585
R10926 gnd.n4604 gnd.n4603 585
R10927 gnd.n4602 gnd.n4601 585
R10928 gnd.n4600 gnd.n4599 585
R10929 gnd.n4598 gnd.n4597 585
R10930 gnd.n4596 gnd.n4595 585
R10931 gnd.n4594 gnd.n4593 585
R10932 gnd.n4592 gnd.n4591 585
R10933 gnd.n4525 gnd.n4513 585
R10934 gnd.n5466 gnd.n5465 585
R10935 gnd.n5468 gnd.n1204 585
R10936 gnd.n5470 gnd.n5469 585
R10937 gnd.n5471 gnd.n1197 585
R10938 gnd.n5473 gnd.n5472 585
R10939 gnd.n5475 gnd.n1195 585
R10940 gnd.n5477 gnd.n5476 585
R10941 gnd.n5478 gnd.n1190 585
R10942 gnd.n5480 gnd.n5479 585
R10943 gnd.n5482 gnd.n1188 585
R10944 gnd.n5484 gnd.n5483 585
R10945 gnd.n5485 gnd.n1183 585
R10946 gnd.n5487 gnd.n5486 585
R10947 gnd.n5489 gnd.n1181 585
R10948 gnd.n5491 gnd.n5490 585
R10949 gnd.n5492 gnd.n1176 585
R10950 gnd.n5494 gnd.n5493 585
R10951 gnd.n5496 gnd.n1175 585
R10952 gnd.n5497 gnd.n1172 585
R10953 gnd.n5500 gnd.n5499 585
R10954 gnd.n1174 gnd.n1168 585
R10955 gnd.n5504 gnd.n1165 585
R10956 gnd.n5506 gnd.n5505 585
R10957 gnd.n5508 gnd.n1163 585
R10958 gnd.n5510 gnd.n5509 585
R10959 gnd.n5511 gnd.n1158 585
R10960 gnd.n5513 gnd.n5512 585
R10961 gnd.n5515 gnd.n1157 585
R10962 gnd.n5516 gnd.n1153 585
R10963 gnd.n5519 gnd.n5518 585
R10964 gnd.n1154 gnd.n1148 585
R10965 gnd.n5408 gnd.n1149 585
R10966 gnd.n5410 gnd.n5409 585
R10967 gnd.n5411 gnd.n5401 585
R10968 gnd.n5413 gnd.n5412 585
R10969 gnd.n5415 gnd.n5399 585
R10970 gnd.n5417 gnd.n5416 585
R10971 gnd.n5418 gnd.n5391 585
R10972 gnd.n5420 gnd.n5419 585
R10973 gnd.n5422 gnd.n5389 585
R10974 gnd.n5424 gnd.n5423 585
R10975 gnd.n5425 gnd.n5384 585
R10976 gnd.n5427 gnd.n5426 585
R10977 gnd.n5429 gnd.n5382 585
R10978 gnd.n5431 gnd.n5430 585
R10979 gnd.n5432 gnd.n5377 585
R10980 gnd.n5434 gnd.n5433 585
R10981 gnd.n5436 gnd.n5375 585
R10982 gnd.n5438 gnd.n5437 585
R10983 gnd.n5439 gnd.n5370 585
R10984 gnd.n5441 gnd.n5440 585
R10985 gnd.n5443 gnd.n5368 585
R10986 gnd.n5445 gnd.n5444 585
R10987 gnd.n5446 gnd.n5364 585
R10988 gnd.n5448 gnd.n5447 585
R10989 gnd.n5450 gnd.n5363 585
R10990 gnd.n5452 gnd.n5451 585
R10991 gnd.n5451 gnd.n1156 585
R10992 gnd.n5461 gnd.n1206 585
R10993 gnd.n5190 gnd.n1206 585
R10994 gnd.n5460 gnd.n5459 585
R10995 gnd.n5459 gnd.n5458 585
R10996 gnd.n1212 gnd.n1211 585
R10997 gnd.n5026 gnd.n1212 585
R10998 gnd.n5349 gnd.n1223 585
R10999 gnd.n5356 gnd.n1223 585
R11000 gnd.n5348 gnd.n5347 585
R11001 gnd.n5347 gnd.n5346 585
R11002 gnd.n1231 gnd.n1230 585
R11003 gnd.n5016 gnd.n1231 585
R11004 gnd.n5001 gnd.n5000 585
R11005 gnd.n5000 gnd.n1284 585
R11006 gnd.n4999 gnd.n1292 585
R11007 gnd.n5008 gnd.n1292 585
R11008 gnd.n4998 gnd.n4997 585
R11009 gnd.n4997 gnd.n4996 585
R11010 gnd.n1301 gnd.n1299 585
R11011 gnd.n4967 gnd.n1301 585
R11012 gnd.n4964 gnd.n1310 585
R11013 gnd.n4984 gnd.n1310 585
R11014 gnd.n4963 gnd.n4962 585
R11015 gnd.n4962 gnd.n4961 585
R11016 gnd.n1327 gnd.n1320 585
R11017 gnd.n4974 gnd.n1320 585
R11018 gnd.n4885 gnd.n1335 585
R11019 gnd.n4940 gnd.n1335 585
R11020 gnd.n4887 gnd.n4886 585
R11021 gnd.n4886 gnd.n1334 585
R11022 gnd.n4884 gnd.n1343 585
R11023 gnd.n4931 gnd.n1343 585
R11024 gnd.n4883 gnd.n4882 585
R11025 gnd.n4882 gnd.n4881 585
R11026 gnd.n4880 gnd.n1392 585
R11027 gnd.n4895 gnd.n1392 585
R11028 gnd.n4879 gnd.n1386 585
R11029 gnd.n4900 gnd.n1386 585
R11030 gnd.n4869 gnd.n1407 585
R11031 gnd.n4869 gnd.n1385 585
R11032 gnd.n4871 gnd.n4870 585
R11033 gnd.n4870 gnd.n1378 585
R11034 gnd.n4868 gnd.n1376 585
R11035 gnd.n4909 gnd.n1376 585
R11036 gnd.n4867 gnd.n1370 585
R11037 gnd.n4914 gnd.n1370 585
R11038 gnd.n4866 gnd.n4865 585
R11039 gnd.n4865 gnd.n4864 585
R11040 gnd.n1409 gnd.n1359 585
R11041 gnd.n4920 gnd.n1359 585
R11042 gnd.n4786 gnd.n1416 585
R11043 gnd.n4853 gnd.n1416 585
R11044 gnd.n4788 gnd.n4787 585
R11045 gnd.n4787 gnd.n1415 585
R11046 gnd.n4789 gnd.n1422 585
R11047 gnd.n4827 gnd.n1422 585
R11048 gnd.n4790 gnd.n1443 585
R11049 gnd.n4812 gnd.n1443 585
R11050 gnd.n4792 gnd.n4791 585
R11051 gnd.n4793 gnd.n4792 585
R11052 gnd.n4780 gnd.n1432 585
R11053 gnd.n4818 gnd.n1432 585
R11054 gnd.n4779 gnd.n1450 585
R11055 gnd.n4799 gnd.n1450 585
R11056 gnd.n1461 gnd.n1456 585
R11057 gnd.n4774 gnd.n1461 585
R11058 gnd.n4761 gnd.n4760 585
R11059 gnd.n4760 gnd.n4759 585
R11060 gnd.n4762 gnd.n1468 585
R11061 gnd.n4766 gnd.n1468 585
R11062 gnd.n4749 gnd.n1474 585
R11063 gnd.n4750 gnd.n4749 585
R11064 gnd.n4748 gnd.n1480 585
R11065 gnd.n4748 gnd.n4747 585
R11066 gnd.n4732 gnd.n1479 585
R11067 gnd.n4722 gnd.n1479 585
R11068 gnd.n4731 gnd.n1490 585
R11069 gnd.n4739 gnd.n1490 585
R11070 gnd.n4730 gnd.n4729 585
R11071 gnd.n4729 gnd.n4728 585
R11072 gnd.n1499 gnd.n1497 585
R11073 gnd.n4519 gnd.n1499 585
R11074 gnd.n4524 gnd.n1507 585
R11075 gnd.n4714 gnd.n1507 585
R11076 gnd.n4586 gnd.n4585 585
R11077 gnd.n4585 gnd.n4584 585
R11078 gnd.n7271 gnd.n7270 585
R11079 gnd.n7270 gnd.n7269 585
R11080 gnd.n7272 gnd.n162 585
R11081 gnd.n7262 gnd.n162 585
R11082 gnd.n7274 gnd.n7273 585
R11083 gnd.n7275 gnd.n7274 585
R11084 gnd.n148 gnd.n147 585
R11085 gnd.n6955 gnd.n148 585
R11086 gnd.n7283 gnd.n7282 585
R11087 gnd.n7282 gnd.n7281 585
R11088 gnd.n7284 gnd.n142 585
R11089 gnd.n6961 gnd.n142 585
R11090 gnd.n7286 gnd.n7285 585
R11091 gnd.n7287 gnd.n7286 585
R11092 gnd.n127 gnd.n126 585
R11093 gnd.n6967 gnd.n127 585
R11094 gnd.n7295 gnd.n7294 585
R11095 gnd.n7294 gnd.n7293 585
R11096 gnd.n7296 gnd.n121 585
R11097 gnd.n6973 gnd.n121 585
R11098 gnd.n7298 gnd.n7297 585
R11099 gnd.n7299 gnd.n7298 585
R11100 gnd.n107 gnd.n106 585
R11101 gnd.n6979 gnd.n107 585
R11102 gnd.n7307 gnd.n7306 585
R11103 gnd.n7306 gnd.n7305 585
R11104 gnd.n7308 gnd.n102 585
R11105 gnd.n6985 gnd.n102 585
R11106 gnd.n7310 gnd.n7309 585
R11107 gnd.n7311 gnd.n7310 585
R11108 gnd.n85 gnd.n83 585
R11109 gnd.n6991 gnd.n85 585
R11110 gnd.n7319 gnd.n7318 585
R11111 gnd.n7318 gnd.n7317 585
R11112 gnd.n84 gnd.n76 585
R11113 gnd.n6997 gnd.n84 585
R11114 gnd.n7322 gnd.n74 585
R11115 gnd.n265 gnd.n74 585
R11116 gnd.n7324 gnd.n7323 585
R11117 gnd.n7325 gnd.n7324 585
R11118 gnd.n6904 gnd.n73 585
R11119 gnd.n6921 gnd.n73 585
R11120 gnd.n6908 gnd.n6905 585
R11121 gnd.n6908 gnd.n6907 585
R11122 gnd.n6911 gnd.n6910 585
R11123 gnd.n6912 gnd.n6911 585
R11124 gnd.n6909 gnd.n6903 585
R11125 gnd.n6903 gnd.n6902 585
R11126 gnd.n6874 gnd.n287 585
R11127 gnd.n6885 gnd.n287 585
R11128 gnd.n6876 gnd.n6875 585
R11129 gnd.n6877 gnd.n6876 585
R11130 gnd.n6873 gnd.n305 585
R11131 gnd.n6873 gnd.n6872 585
R11132 gnd.n6845 gnd.n304 585
R11133 gnd.n6865 gnd.n304 585
R11134 gnd.n6846 gnd.n325 585
R11135 gnd.n6831 gnd.n325 585
R11136 gnd.n6848 gnd.n6847 585
R11137 gnd.n6849 gnd.n6848 585
R11138 gnd.n326 gnd.n324 585
R11139 gnd.n6826 gnd.n324 585
R11140 gnd.n6840 gnd.n6839 585
R11141 gnd.n6839 gnd.n6838 585
R11142 gnd.n329 gnd.n328 585
R11143 gnd.n6822 gnd.n329 585
R11144 gnd.n6810 gnd.n354 585
R11145 gnd.n6796 gnd.n354 585
R11146 gnd.n6812 gnd.n6811 585
R11147 gnd.n6813 gnd.n6812 585
R11148 gnd.n355 gnd.n353 585
R11149 gnd.n6790 gnd.n353 585
R11150 gnd.n6805 gnd.n6804 585
R11151 gnd.n6804 gnd.n6803 585
R11152 gnd.n358 gnd.n357 585
R11153 gnd.n6753 gnd.n358 585
R11154 gnd.n6741 gnd.n387 585
R11155 gnd.n387 gnd.n374 585
R11156 gnd.n6743 gnd.n6742 585
R11157 gnd.n6744 gnd.n6743 585
R11158 gnd.n388 gnd.n386 585
R11159 gnd.n6727 gnd.n386 585
R11160 gnd.n6736 gnd.n6735 585
R11161 gnd.n6735 gnd.n6734 585
R11162 gnd.n391 gnd.n390 585
R11163 gnd.n6715 gnd.n391 585
R11164 gnd.n6691 gnd.n6690 585
R11165 gnd.n6689 gnd.n496 585
R11166 gnd.n6688 gnd.n495 585
R11167 gnd.n6693 gnd.n495 585
R11168 gnd.n6687 gnd.n6686 585
R11169 gnd.n6685 gnd.n6684 585
R11170 gnd.n6683 gnd.n6682 585
R11171 gnd.n6681 gnd.n6680 585
R11172 gnd.n6679 gnd.n6678 585
R11173 gnd.n6677 gnd.n6676 585
R11174 gnd.n6675 gnd.n6674 585
R11175 gnd.n6673 gnd.n6672 585
R11176 gnd.n6671 gnd.n6670 585
R11177 gnd.n6669 gnd.n6668 585
R11178 gnd.n6667 gnd.n6666 585
R11179 gnd.n6665 gnd.n6664 585
R11180 gnd.n6663 gnd.n6662 585
R11181 gnd.n6661 gnd.n6660 585
R11182 gnd.n6659 gnd.n6658 585
R11183 gnd.n6656 gnd.n6655 585
R11184 gnd.n6654 gnd.n6653 585
R11185 gnd.n6652 gnd.n6651 585
R11186 gnd.n6650 gnd.n6649 585
R11187 gnd.n6648 gnd.n6647 585
R11188 gnd.n6646 gnd.n6645 585
R11189 gnd.n6644 gnd.n6643 585
R11190 gnd.n6642 gnd.n6641 585
R11191 gnd.n6639 gnd.n6638 585
R11192 gnd.n6637 gnd.n6636 585
R11193 gnd.n6635 gnd.n6634 585
R11194 gnd.n6633 gnd.n6632 585
R11195 gnd.n6631 gnd.n6630 585
R11196 gnd.n6629 gnd.n6628 585
R11197 gnd.n6627 gnd.n6626 585
R11198 gnd.n6625 gnd.n6624 585
R11199 gnd.n6623 gnd.n6622 585
R11200 gnd.n6621 gnd.n6620 585
R11201 gnd.n6619 gnd.n6618 585
R11202 gnd.n6617 gnd.n6616 585
R11203 gnd.n6615 gnd.n6614 585
R11204 gnd.n6613 gnd.n6612 585
R11205 gnd.n6611 gnd.n6610 585
R11206 gnd.n6609 gnd.n6608 585
R11207 gnd.n6607 gnd.n6606 585
R11208 gnd.n6605 gnd.n6604 585
R11209 gnd.n6603 gnd.n6602 585
R11210 gnd.n6601 gnd.n6600 585
R11211 gnd.n6599 gnd.n6598 585
R11212 gnd.n6597 gnd.n6596 585
R11213 gnd.n6595 gnd.n6594 585
R11214 gnd.n6593 gnd.n6592 585
R11215 gnd.n6591 gnd.n6590 585
R11216 gnd.n6589 gnd.n6588 585
R11217 gnd.n6587 gnd.n6586 585
R11218 gnd.n6585 gnd.n6584 585
R11219 gnd.n6583 gnd.n6582 585
R11220 gnd.n6581 gnd.n6580 585
R11221 gnd.n560 gnd.n559 585
R11222 gnd.n7131 gnd.n7130 585
R11223 gnd.n7137 gnd.n7136 585
R11224 gnd.n7139 gnd.n7138 585
R11225 gnd.n7141 gnd.n7140 585
R11226 gnd.n7143 gnd.n7142 585
R11227 gnd.n7145 gnd.n7144 585
R11228 gnd.n7147 gnd.n7146 585
R11229 gnd.n7149 gnd.n7148 585
R11230 gnd.n7151 gnd.n7150 585
R11231 gnd.n7153 gnd.n7152 585
R11232 gnd.n7155 gnd.n7154 585
R11233 gnd.n7157 gnd.n7156 585
R11234 gnd.n7159 gnd.n7158 585
R11235 gnd.n7161 gnd.n7160 585
R11236 gnd.n7163 gnd.n7162 585
R11237 gnd.n7165 gnd.n7164 585
R11238 gnd.n7167 gnd.n7166 585
R11239 gnd.n7169 gnd.n7168 585
R11240 gnd.n7171 gnd.n7170 585
R11241 gnd.n7174 gnd.n7173 585
R11242 gnd.n7172 gnd.n7110 585
R11243 gnd.n7179 gnd.n7178 585
R11244 gnd.n7181 gnd.n7180 585
R11245 gnd.n7183 gnd.n7182 585
R11246 gnd.n7185 gnd.n7184 585
R11247 gnd.n7187 gnd.n7186 585
R11248 gnd.n7189 gnd.n7188 585
R11249 gnd.n7191 gnd.n7190 585
R11250 gnd.n7193 gnd.n7192 585
R11251 gnd.n7195 gnd.n7194 585
R11252 gnd.n7197 gnd.n7196 585
R11253 gnd.n7199 gnd.n7198 585
R11254 gnd.n7201 gnd.n7200 585
R11255 gnd.n7203 gnd.n7202 585
R11256 gnd.n7205 gnd.n7204 585
R11257 gnd.n7207 gnd.n7206 585
R11258 gnd.n7209 gnd.n7208 585
R11259 gnd.n7211 gnd.n7210 585
R11260 gnd.n7213 gnd.n7212 585
R11261 gnd.n7215 gnd.n7214 585
R11262 gnd.n7217 gnd.n7216 585
R11263 gnd.n7222 gnd.n7221 585
R11264 gnd.n7224 gnd.n7223 585
R11265 gnd.n7226 gnd.n7225 585
R11266 gnd.n7228 gnd.n7227 585
R11267 gnd.n7230 gnd.n7229 585
R11268 gnd.n7232 gnd.n7231 585
R11269 gnd.n7234 gnd.n7233 585
R11270 gnd.n7236 gnd.n7235 585
R11271 gnd.n7238 gnd.n7237 585
R11272 gnd.n7240 gnd.n7239 585
R11273 gnd.n7242 gnd.n7241 585
R11274 gnd.n7244 gnd.n7243 585
R11275 gnd.n7246 gnd.n7245 585
R11276 gnd.n7248 gnd.n7247 585
R11277 gnd.n7249 gnd.n7070 585
R11278 gnd.n7251 gnd.n7250 585
R11279 gnd.n7071 gnd.n7069 585
R11280 gnd.n7072 gnd.n167 585
R11281 gnd.n7253 gnd.n167 585
R11282 gnd.n7265 gnd.n169 585
R11283 gnd.n7269 gnd.n169 585
R11284 gnd.n7264 gnd.n7263 585
R11285 gnd.n7263 gnd.n7262 585
R11286 gnd.n175 gnd.n160 585
R11287 gnd.n7275 gnd.n160 585
R11288 gnd.n6954 gnd.n6953 585
R11289 gnd.n6955 gnd.n6954 585
R11290 gnd.n6947 gnd.n150 585
R11291 gnd.n7281 gnd.n150 585
R11292 gnd.n6963 gnd.n6962 585
R11293 gnd.n6962 gnd.n6961 585
R11294 gnd.n6964 gnd.n139 585
R11295 gnd.n7287 gnd.n139 585
R11296 gnd.n6966 gnd.n6965 585
R11297 gnd.n6967 gnd.n6966 585
R11298 gnd.n6940 gnd.n129 585
R11299 gnd.n7293 gnd.n129 585
R11300 gnd.n6975 gnd.n6974 585
R11301 gnd.n6974 gnd.n6973 585
R11302 gnd.n6976 gnd.n118 585
R11303 gnd.n7299 gnd.n118 585
R11304 gnd.n6978 gnd.n6977 585
R11305 gnd.n6979 gnd.n6978 585
R11306 gnd.n6932 gnd.n109 585
R11307 gnd.n7305 gnd.n109 585
R11308 gnd.n6987 gnd.n6986 585
R11309 gnd.n6986 gnd.n6985 585
R11310 gnd.n6988 gnd.n99 585
R11311 gnd.n7311 gnd.n99 585
R11312 gnd.n6990 gnd.n6989 585
R11313 gnd.n6991 gnd.n6990 585
R11314 gnd.n6930 gnd.n87 585
R11315 gnd.n7317 gnd.n87 585
R11316 gnd.n6929 gnd.n266 585
R11317 gnd.n6997 gnd.n266 585
R11318 gnd.n273 gnd.n272 585
R11319 gnd.n272 gnd.n265 585
R11320 gnd.n6918 gnd.n70 585
R11321 gnd.n7325 gnd.n70 585
R11322 gnd.n6920 gnd.n6919 585
R11323 gnd.n6921 gnd.n6920 585
R11324 gnd.n6917 gnd.n279 585
R11325 gnd.n6907 gnd.n279 585
R11326 gnd.n284 gnd.n280 585
R11327 gnd.n6912 gnd.n284 585
R11328 gnd.n6880 gnd.n289 585
R11329 gnd.n6902 gnd.n289 585
R11330 gnd.n6881 gnd.n295 585
R11331 gnd.n6885 gnd.n295 585
R11332 gnd.n6879 gnd.n6878 585
R11333 gnd.n6878 gnd.n6877 585
R11334 gnd.n301 gnd.n300 585
R11335 gnd.n6872 gnd.n301 585
R11336 gnd.n6867 gnd.n6866 585
R11337 gnd.n6866 gnd.n6865 585
R11338 gnd.n312 gnd.n311 585
R11339 gnd.n6831 gnd.n312 585
R11340 gnd.n6829 gnd.n321 585
R11341 gnd.n6849 gnd.n321 585
R11342 gnd.n6828 gnd.n6827 585
R11343 gnd.n6827 gnd.n6826 585
R11344 gnd.n6825 gnd.n331 585
R11345 gnd.n6838 gnd.n331 585
R11346 gnd.n6824 gnd.n6823 585
R11347 gnd.n6823 gnd.n6822 585
R11348 gnd.n341 gnd.n339 585
R11349 gnd.n6796 gnd.n341 585
R11350 gnd.n6793 gnd.n350 585
R11351 gnd.n6813 gnd.n350 585
R11352 gnd.n6792 gnd.n6791 585
R11353 gnd.n6791 gnd.n6790 585
R11354 gnd.n367 gnd.n360 585
R11355 gnd.n6803 gnd.n360 585
R11356 gnd.n408 gnd.n375 585
R11357 gnd.n6753 gnd.n375 585
R11358 gnd.n410 gnd.n409 585
R11359 gnd.n409 gnd.n374 585
R11360 gnd.n411 gnd.n383 585
R11361 gnd.n6744 gnd.n383 585
R11362 gnd.n6729 gnd.n6728 585
R11363 gnd.n6728 gnd.n6727 585
R11364 gnd.n6730 gnd.n393 585
R11365 gnd.n6734 gnd.n393 585
R11366 gnd.n419 gnd.n401 585
R11367 gnd.n6715 gnd.n419 585
R11368 gnd.n4416 gnd.n1555 585
R11369 gnd.n1555 gnd.n1516 585
R11370 gnd.n7039 gnd.n7038 585
R11371 gnd.n7040 gnd.n7039 585
R11372 gnd.n7035 gnd.n244 585
R11373 gnd.n244 gnd.n171 585
R11374 gnd.n7034 gnd.n7033 585
R11375 gnd.n7033 gnd.n168 585
R11376 gnd.n7032 gnd.n248 585
R11377 gnd.n7032 gnd.n176 585
R11378 gnd.n7031 gnd.n7030 585
R11379 gnd.n7031 gnd.n159 585
R11380 gnd.n250 gnd.n249 585
R11381 gnd.n249 gnd.n152 585
R11382 gnd.n7025 gnd.n7024 585
R11383 gnd.n7024 gnd.n149 585
R11384 gnd.n7023 gnd.n252 585
R11385 gnd.n7023 gnd.n141 585
R11386 gnd.n7022 gnd.n7021 585
R11387 gnd.n7022 gnd.n138 585
R11388 gnd.n254 gnd.n253 585
R11389 gnd.n253 gnd.n131 585
R11390 gnd.n7017 gnd.n7016 585
R11391 gnd.n7016 gnd.n128 585
R11392 gnd.n7015 gnd.n256 585
R11393 gnd.n7015 gnd.n120 585
R11394 gnd.n7014 gnd.n7013 585
R11395 gnd.n7014 gnd.n117 585
R11396 gnd.n258 gnd.n257 585
R11397 gnd.n6938 gnd.n257 585
R11398 gnd.n7009 gnd.n7008 585
R11399 gnd.n7008 gnd.n108 585
R11400 gnd.n7007 gnd.n260 585
R11401 gnd.n7007 gnd.n101 585
R11402 gnd.n7006 gnd.n7005 585
R11403 gnd.n7006 gnd.n98 585
R11404 gnd.n7002 gnd.n261 585
R11405 gnd.n261 gnd.n89 585
R11406 gnd.n7001 gnd.n7000 585
R11407 gnd.n7000 gnd.n86 585
R11408 gnd.n6999 gnd.n264 585
R11409 gnd.n6999 gnd.n6998 585
R11410 gnd.n6891 gnd.n263 585
R11411 gnd.n263 gnd.n71 585
R11412 gnd.n6894 gnd.n6893 585
R11413 gnd.n6894 gnd.n69 585
R11414 gnd.n6896 gnd.n6895 585
R11415 gnd.n6895 gnd.n278 585
R11416 gnd.n6898 gnd.n292 585
R11417 gnd.n292 gnd.n286 585
R11418 gnd.n6900 gnd.n6899 585
R11419 gnd.n6901 gnd.n6900 585
R11420 gnd.n6889 gnd.n291 585
R11421 gnd.n291 gnd.n288 585
R11422 gnd.n6888 gnd.n6887 585
R11423 gnd.n6887 gnd.n6886 585
R11424 gnd.n6773 gnd.n294 585
R11425 gnd.n302 gnd.n294 585
R11426 gnd.n6774 gnd.n6769 585
R11427 gnd.n6769 gnd.n306 585
R11428 gnd.n6776 gnd.n6775 585
R11429 gnd.n6776 gnd.n313 585
R11430 gnd.n6777 gnd.n6768 585
R11431 gnd.n6777 gnd.n322 585
R11432 gnd.n6779 gnd.n6778 585
R11433 gnd.n6778 gnd.n320 585
R11434 gnd.n6780 gnd.n6763 585
R11435 gnd.n6763 gnd.n333 585
R11436 gnd.n6782 gnd.n6781 585
R11437 gnd.n6782 gnd.n330 585
R11438 gnd.n6783 gnd.n6762 585
R11439 gnd.n6783 gnd.n342 585
R11440 gnd.n6785 gnd.n6784 585
R11441 gnd.n6784 gnd.n351 585
R11442 gnd.n6786 gnd.n369 585
R11443 gnd.n369 gnd.n349 585
R11444 gnd.n6788 gnd.n6787 585
R11445 gnd.n6789 gnd.n6788 585
R11446 gnd.n370 gnd.n368 585
R11447 gnd.n368 gnd.n359 585
R11448 gnd.n6756 gnd.n6755 585
R11449 gnd.n6755 gnd.n6754 585
R11450 gnd.n373 gnd.n372 585
R11451 gnd.n384 gnd.n373 585
R11452 gnd.n6723 gnd.n413 585
R11453 gnd.n413 gnd.n382 585
R11454 gnd.n6725 gnd.n6724 585
R11455 gnd.n6726 gnd.n6725 585
R11456 gnd.n414 gnd.n412 585
R11457 gnd.n412 gnd.n392 585
R11458 gnd.n6718 gnd.n6717 585
R11459 gnd.n6717 gnd.n6716 585
R11460 gnd.n417 gnd.n416 585
R11461 gnd.n418 gnd.n417 585
R11462 gnd.n6454 gnd.n6453 585
R11463 gnd.n6454 gnd.n457 585
R11464 gnd.n6456 gnd.n6450 585
R11465 gnd.n6456 gnd.n6455 585
R11466 gnd.n6458 gnd.n6457 585
R11467 gnd.n6457 gnd.n442 585
R11468 gnd.n6459 gnd.n574 585
R11469 gnd.n574 gnd.n427 585
R11470 gnd.n6461 gnd.n6460 585
R11471 gnd.n6462 gnd.n6461 585
R11472 gnd.n575 gnd.n573 585
R11473 gnd.n573 gnd.n572 585
R11474 gnd.n6444 gnd.n6443 585
R11475 gnd.n6443 gnd.n6442 585
R11476 gnd.n578 gnd.n577 585
R11477 gnd.n586 gnd.n578 585
R11478 gnd.n6419 gnd.n599 585
R11479 gnd.n599 gnd.n585 585
R11480 gnd.n6421 gnd.n6420 585
R11481 gnd.n6422 gnd.n6421 585
R11482 gnd.n600 gnd.n598 585
R11483 gnd.n598 gnd.n595 585
R11484 gnd.n6414 gnd.n6413 585
R11485 gnd.n6413 gnd.n6412 585
R11486 gnd.n603 gnd.n602 585
R11487 gnd.n612 gnd.n603 585
R11488 gnd.n6389 gnd.n624 585
R11489 gnd.n624 gnd.n611 585
R11490 gnd.n6391 gnd.n6390 585
R11491 gnd.n6392 gnd.n6391 585
R11492 gnd.n625 gnd.n623 585
R11493 gnd.n623 gnd.n620 585
R11494 gnd.n6384 gnd.n6383 585
R11495 gnd.n6383 gnd.n6382 585
R11496 gnd.n628 gnd.n627 585
R11497 gnd.n637 gnd.n628 585
R11498 gnd.n6359 gnd.n649 585
R11499 gnd.n649 gnd.n636 585
R11500 gnd.n6361 gnd.n6360 585
R11501 gnd.n6362 gnd.n6361 585
R11502 gnd.n650 gnd.n648 585
R11503 gnd.n648 gnd.n645 585
R11504 gnd.n6354 gnd.n6353 585
R11505 gnd.n6353 gnd.n6352 585
R11506 gnd.n653 gnd.n652 585
R11507 gnd.t130 gnd.n653 585
R11508 gnd.n6187 gnd.n6186 585
R11509 gnd.n6188 gnd.n6187 585
R11510 gnd.n703 gnd.n702 585
R11511 gnd.n6001 gnd.n702 585
R11512 gnd.n6182 gnd.n6181 585
R11513 gnd.n6181 gnd.n6180 585
R11514 gnd.n706 gnd.n705 585
R11515 gnd.n719 gnd.n706 585
R11516 gnd.n6148 gnd.n6147 585
R11517 gnd.n6149 gnd.n6148 585
R11518 gnd.n729 gnd.n728 585
R11519 gnd.n728 gnd.n724 585
R11520 gnd.n6143 gnd.n6142 585
R11521 gnd.n6142 gnd.n6141 585
R11522 gnd.n732 gnd.n731 585
R11523 gnd.n6131 gnd.n732 585
R11524 gnd.n6121 gnd.n6120 585
R11525 gnd.n6122 gnd.n6121 585
R11526 gnd.n752 gnd.n751 585
R11527 gnd.n5984 gnd.n751 585
R11528 gnd.n6116 gnd.n6115 585
R11529 gnd.n6115 gnd.n6114 585
R11530 gnd.n755 gnd.n754 585
R11531 gnd.n5975 gnd.n755 585
R11532 gnd.n6085 gnd.n780 585
R11533 gnd.n5974 gnd.n780 585
R11534 gnd.n6087 gnd.n6086 585
R11535 gnd.n6088 gnd.n6087 585
R11536 gnd.n781 gnd.n779 585
R11537 gnd.n787 gnd.n779 585
R11538 gnd.n6080 gnd.n6079 585
R11539 gnd.n6079 gnd.n6078 585
R11540 gnd.n784 gnd.n783 585
R11541 gnd.n797 gnd.n784 585
R11542 gnd.n5932 gnd.n5931 585
R11543 gnd.n5931 gnd.n794 585
R11544 gnd.n5933 gnd.n827 585
R11545 gnd.n827 gnd.n802 585
R11546 gnd.n5935 gnd.n5934 585
R11547 gnd.n5936 gnd.n5935 585
R11548 gnd.n828 gnd.n826 585
R11549 gnd.n5915 gnd.n826 585
R11550 gnd.n5925 gnd.n5924 585
R11551 gnd.n5924 gnd.n5923 585
R11552 gnd.n831 gnd.n830 585
R11553 gnd.n838 gnd.n831 585
R11554 gnd.n5876 gnd.n5875 585
R11555 gnd.n5876 gnd.n836 585
R11556 gnd.n5878 gnd.n5877 585
R11557 gnd.n5877 gnd.n845 585
R11558 gnd.n5879 gnd.n866 585
R11559 gnd.n866 gnd.n858 585
R11560 gnd.n5881 gnd.n5880 585
R11561 gnd.n5882 gnd.n5881 585
R11562 gnd.n867 gnd.n865 585
R11563 gnd.n865 gnd.n862 585
R11564 gnd.n5868 gnd.n5867 585
R11565 gnd.n5867 gnd.n5866 585
R11566 gnd.n870 gnd.n869 585
R11567 gnd.n5858 gnd.n870 585
R11568 gnd.n5780 gnd.n5779 585
R11569 gnd.n5781 gnd.n5780 585
R11570 gnd.n918 gnd.n917 585
R11571 gnd.n917 gnd.n916 585
R11572 gnd.n5775 gnd.n5774 585
R11573 gnd.n5774 gnd.n893 585
R11574 gnd.n5773 gnd.n920 585
R11575 gnd.n5773 gnd.n903 585
R11576 gnd.n5772 gnd.n5771 585
R11577 gnd.n5772 gnd.n900 585
R11578 gnd.n922 gnd.n921 585
R11579 gnd.n949 gnd.n921 585
R11580 gnd.n5767 gnd.n5766 585
R11581 gnd.n5766 gnd.n5765 585
R11582 gnd.n925 gnd.n924 585
R11583 gnd.n935 gnd.n925 585
R11584 gnd.n5701 gnd.n983 585
R11585 gnd.n5682 gnd.n983 585
R11586 gnd.n5703 gnd.n5702 585
R11587 gnd.n5704 gnd.n5703 585
R11588 gnd.n984 gnd.n982 585
R11589 gnd.n982 gnd.n981 585
R11590 gnd.n5696 gnd.n5695 585
R11591 gnd.n5695 gnd.n5694 585
R11592 gnd.n987 gnd.n986 585
R11593 gnd.n987 gnd.n971 585
R11594 gnd.n5641 gnd.n5639 585
R11595 gnd.n5641 gnd.n5640 585
R11596 gnd.n5642 gnd.n5636 585
R11597 gnd.n5642 gnd.n991 585
R11598 gnd.n5644 gnd.n5643 585
R11599 gnd.n5643 gnd.n996 585
R11600 gnd.n5645 gnd.n1065 585
R11601 gnd.n1065 gnd.n1007 585
R11602 gnd.n5647 gnd.n5646 585
R11603 gnd.n5648 gnd.n5647 585
R11604 gnd.n1066 gnd.n1064 585
R11605 gnd.n1072 gnd.n1064 585
R11606 gnd.n5630 gnd.n5629 585
R11607 gnd.n5629 gnd.n5628 585
R11608 gnd.n1069 gnd.n1068 585
R11609 gnd.n5618 gnd.n1069 585
R11610 gnd.n5148 gnd.n5063 585
R11611 gnd.n5063 gnd.n1078 585
R11612 gnd.n5150 gnd.n5149 585
R11613 gnd.n5151 gnd.n5150 585
R11614 gnd.n5064 gnd.n5062 585
R11615 gnd.n5139 gnd.n5062 585
R11616 gnd.n5143 gnd.n5142 585
R11617 gnd.n5142 gnd.n5141 585
R11618 gnd.n5067 gnd.n5066 585
R11619 gnd.n5129 gnd.n5067 585
R11620 gnd.n5127 gnd.n5126 585
R11621 gnd.n5128 gnd.n5127 585
R11622 gnd.n5077 gnd.n5076 585
R11623 gnd.n5117 gnd.n5076 585
R11624 gnd.n5122 gnd.n5121 585
R11625 gnd.n5121 gnd.n5120 585
R11626 gnd.n5080 gnd.n5079 585
R11627 gnd.n5108 gnd.n5080 585
R11628 gnd.n5106 gnd.n5105 585
R11629 gnd.n5107 gnd.n5106 585
R11630 gnd.n5098 gnd.n5097 585
R11631 gnd.n5097 gnd.n5096 585
R11632 gnd.n5101 gnd.n5100 585
R11633 gnd.n5100 gnd.n5044 585
R11634 gnd.n5042 gnd.n5041 585
R11635 gnd.n5173 gnd.n5042 585
R11636 gnd.n5177 gnd.n5176 585
R11637 gnd.n5176 gnd.n5175 585
R11638 gnd.n5178 gnd.n5036 585
R11639 gnd.n5036 gnd.n1259 585
R11640 gnd.n5180 gnd.n5179 585
R11641 gnd.n5180 gnd.n1245 585
R11642 gnd.n5181 gnd.n5035 585
R11643 gnd.n5182 gnd.n5181 585
R11644 gnd.n5185 gnd.n5184 585
R11645 gnd.n5184 gnd.n5183 585
R11646 gnd.n5186 gnd.n1275 585
R11647 gnd.n1275 gnd.n1273 585
R11648 gnd.n5188 gnd.n5187 585
R11649 gnd.n5189 gnd.n5188 585
R11650 gnd.n1276 gnd.n1274 585
R11651 gnd.n1274 gnd.n1214 585
R11652 gnd.n5029 gnd.n5028 585
R11653 gnd.n5028 gnd.n5027 585
R11654 gnd.n5025 gnd.n1278 585
R11655 gnd.n5025 gnd.n1225 585
R11656 gnd.n5024 gnd.n5023 585
R11657 gnd.n5024 gnd.n1222 585
R11658 gnd.n1280 gnd.n1279 585
R11659 gnd.n1279 gnd.n1232 585
R11660 gnd.n5019 gnd.n5018 585
R11661 gnd.n5018 gnd.n5017 585
R11662 gnd.n1283 gnd.n1282 585
R11663 gnd.n1294 gnd.n1283 585
R11664 gnd.n4953 gnd.n4952 585
R11665 gnd.n4953 gnd.n1291 585
R11666 gnd.n4954 gnd.n4949 585
R11667 gnd.n4954 gnd.n1302 585
R11668 gnd.n4956 gnd.n4955 585
R11669 gnd.n4955 gnd.n1311 585
R11670 gnd.n4957 gnd.n1329 585
R11671 gnd.n1329 gnd.n1309 585
R11672 gnd.n4959 gnd.n4958 585
R11673 gnd.n4960 gnd.n4959 585
R11674 gnd.n1330 gnd.n1328 585
R11675 gnd.n1328 gnd.n1319 585
R11676 gnd.n4943 gnd.n4942 585
R11677 gnd.n4942 gnd.n4941 585
R11678 gnd.n1333 gnd.n1332 585
R11679 gnd.n1344 gnd.n1333 585
R11680 gnd.n1397 gnd.n1394 585
R11681 gnd.n1394 gnd.n1342 585
R11682 gnd.n1399 gnd.n1398 585
R11683 gnd.n1400 gnd.n1399 585
R11684 gnd.n1383 gnd.n1382 585
R11685 gnd.n1388 gnd.n1383 585
R11686 gnd.n4903 gnd.n4902 585
R11687 gnd.n4902 gnd.n4901 585
R11688 gnd.n4905 gnd.n1380 585
R11689 gnd.n1384 gnd.n1380 585
R11690 gnd.n4907 gnd.n4906 585
R11691 gnd.n4908 gnd.n4907 585
R11692 gnd.n4860 gnd.n1379 585
R11693 gnd.n1379 gnd.n1372 585
R11694 gnd.n4862 gnd.n4861 585
R11695 gnd.n4863 gnd.n4862 585
R11696 gnd.n4858 gnd.n1411 585
R11697 gnd.n1411 gnd.n1361 585
R11698 gnd.n4857 gnd.n4856 585
R11699 gnd.n4856 gnd.n1358 585
R11700 gnd.n4855 gnd.n1414 585
R11701 gnd.n4855 gnd.n4854 585
R11702 gnd.n4808 gnd.n1413 585
R11703 gnd.n1423 gnd.n1413 585
R11704 gnd.n4810 gnd.n4809 585
R11705 gnd.n4811 gnd.n4810 585
R11706 gnd.n1445 gnd.n1444 585
R11707 gnd.n1444 gnd.n1442 585
R11708 gnd.n4803 gnd.n4802 585
R11709 gnd.n4802 gnd.n1434 585
R11710 gnd.n4801 gnd.n1447 585
R11711 gnd.n4801 gnd.n4800 585
R11712 gnd.n4434 gnd.n1448 585
R11713 gnd.n1449 gnd.n1448 585
R11714 gnd.n4436 gnd.n4435 585
R11715 gnd.n4435 gnd.n1460 585
R11716 gnd.n4437 gnd.n4428 585
R11717 gnd.n4428 gnd.n1470 585
R11718 gnd.n4439 gnd.n4438 585
R11719 gnd.n4439 gnd.n1467 585
R11720 gnd.n4440 gnd.n4427 585
R11721 gnd.n4440 gnd.n1482 585
R11722 gnd.n4442 gnd.n4441 585
R11723 gnd.n4441 gnd.n1481 585
R11724 gnd.n4443 gnd.n4422 585
R11725 gnd.n4422 gnd.n1492 585
R11726 gnd.n4445 gnd.n4444 585
R11727 gnd.n4445 gnd.n1489 585
R11728 gnd.n4446 gnd.n4421 585
R11729 gnd.n4446 gnd.n1500 585
R11730 gnd.n4448 gnd.n4447 585
R11731 gnd.n4447 gnd.n1508 585
R11732 gnd.n4449 gnd.n1556 585
R11733 gnd.n1556 gnd.n1506 585
R11734 gnd.n4451 gnd.n4450 585
R11735 gnd.n4452 gnd.n4451 585
R11736 gnd.n6465 gnd.n6464 585
R11737 gnd.n6464 gnd.n6463 585
R11738 gnd.n570 gnd.n569 585
R11739 gnd.n6441 gnd.n570 585
R11740 gnd.n591 gnd.n589 585
R11741 gnd.n589 gnd.n588 585
R11742 gnd.n6431 gnd.n6430 585
R11743 gnd.n6432 gnd.n6431 585
R11744 gnd.n590 gnd.n587 585
R11745 gnd.n597 gnd.n587 585
R11746 gnd.n6425 gnd.n6424 585
R11747 gnd.n6424 gnd.n6423 585
R11748 gnd.n594 gnd.n593 585
R11749 gnd.n6411 gnd.n594 585
R11750 gnd.n616 gnd.n614 585
R11751 gnd.n614 gnd.n604 585
R11752 gnd.n6401 gnd.n6400 585
R11753 gnd.n6402 gnd.n6401 585
R11754 gnd.n615 gnd.n613 585
R11755 gnd.n622 gnd.n613 585
R11756 gnd.n6395 gnd.n6394 585
R11757 gnd.n6394 gnd.n6393 585
R11758 gnd.n619 gnd.n618 585
R11759 gnd.n6381 gnd.n619 585
R11760 gnd.n641 gnd.n639 585
R11761 gnd.n639 gnd.n629 585
R11762 gnd.n6371 gnd.n6370 585
R11763 gnd.n6372 gnd.n6371 585
R11764 gnd.n640 gnd.n638 585
R11765 gnd.n647 gnd.n638 585
R11766 gnd.n6365 gnd.n6364 585
R11767 gnd.n6364 gnd.n6363 585
R11768 gnd.n644 gnd.n643 585
R11769 gnd.n6351 gnd.n644 585
R11770 gnd.n6172 gnd.n6171 585
R11771 gnd.n6171 gnd.n654 585
R11772 gnd.n6173 gnd.n6170 585
R11773 gnd.n6170 gnd.n701 585
R11774 gnd.n713 gnd.n711 585
R11775 gnd.n711 gnd.n698 585
R11776 gnd.n6178 gnd.n6177 585
R11777 gnd.n6179 gnd.n6178 585
R11778 gnd.n712 gnd.n710 585
R11779 gnd.n6010 gnd.n710 585
R11780 gnd.n6166 gnd.n6165 585
R11781 gnd.n6165 gnd.n6164 585
R11782 gnd.n716 gnd.n715 585
R11783 gnd.n6151 gnd.n716 585
R11784 gnd.n6139 gnd.n6138 585
R11785 gnd.n6140 gnd.n6139 585
R11786 gnd.n737 gnd.n736 585
R11787 gnd.n744 gnd.n736 585
R11788 gnd.n6134 gnd.n6133 585
R11789 gnd.n6133 gnd.n6132 585
R11790 gnd.n740 gnd.n739 585
R11791 gnd.n749 gnd.n740 585
R11792 gnd.n767 gnd.n765 585
R11793 gnd.n765 gnd.n758 585
R11794 gnd.n6105 gnd.n6104 585
R11795 gnd.n6106 gnd.n6105 585
R11796 gnd.n766 gnd.n764 585
R11797 gnd.n5976 gnd.n764 585
R11798 gnd.n6099 gnd.n6098 585
R11799 gnd.n6098 gnd.n6097 585
R11800 gnd.n770 gnd.n769 585
R11801 gnd.n6089 gnd.n770 585
R11802 gnd.n6076 gnd.n6075 585
R11803 gnd.n6077 gnd.n6076 585
R11804 gnd.n790 gnd.n789 585
R11805 gnd.n6050 gnd.n789 585
R11806 gnd.n6071 gnd.n6070 585
R11807 gnd.n6070 gnd.n6069 585
R11808 gnd.n793 gnd.n792 585
R11809 gnd.n6058 gnd.n793 585
R11810 gnd.n5951 gnd.n5950 585
R11811 gnd.n5952 gnd.n5951 585
R11812 gnd.n815 gnd.n814 585
R11813 gnd.n824 gnd.n814 585
R11814 gnd.n5946 gnd.n5945 585
R11815 gnd.n5945 gnd.n5944 585
R11816 gnd.n818 gnd.n817 585
R11817 gnd.n832 gnd.n818 585
R11818 gnd.n851 gnd.n839 585
R11819 gnd.n5908 gnd.n839 585
R11820 gnd.n5899 gnd.n5898 585
R11821 gnd.n5900 gnd.n5899 585
R11822 gnd.n850 gnd.n849 585
R11823 gnd.n5819 gnd.n849 585
R11824 gnd.n5893 gnd.n5892 585
R11825 gnd.n5892 gnd.n5891 585
R11826 gnd.n854 gnd.n853 585
R11827 gnd.n5883 gnd.n854 585
R11828 gnd.n5849 gnd.n5848 585
R11829 gnd.n5850 gnd.n5849 585
R11830 gnd.n881 gnd.n880 585
R11831 gnd.n880 gnd.n871 585
R11832 gnd.n5844 gnd.n5843 585
R11833 gnd.n5843 gnd.n5842 585
R11834 gnd.n884 gnd.n883 585
R11835 gnd.n5782 gnd.n884 585
R11836 gnd.n5805 gnd.n5804 585
R11837 gnd.n5806 gnd.n5805 585
R11838 gnd.n896 gnd.n895 585
R11839 gnd.n909 gnd.n895 585
R11840 gnd.n5800 gnd.n5799 585
R11841 gnd.n5799 gnd.n5798 585
R11842 gnd.n899 gnd.n898 585
R11843 gnd.n5740 gnd.n899 585
R11844 gnd.n5763 gnd.n5762 585
R11845 gnd.n5764 gnd.n5763 585
R11846 gnd.n929 gnd.n928 585
R11847 gnd.n941 gnd.n928 585
R11848 gnd.n5758 gnd.n5757 585
R11849 gnd.n5757 gnd.n5756 585
R11850 gnd.n932 gnd.n931 585
R11851 gnd.n5681 gnd.n932 585
R11852 gnd.n964 gnd.n962 585
R11853 gnd.n5705 gnd.n962 585
R11854 gnd.n5722 gnd.n5721 585
R11855 gnd.n5723 gnd.n5722 585
R11856 gnd.n963 gnd.n961 585
R11857 gnd.n5693 gnd.n961 585
R11858 gnd.n5716 gnd.n5715 585
R11859 gnd.n5715 gnd.n5714 585
R11860 gnd.n967 gnd.n966 585
R11861 gnd.n992 gnd.n967 585
R11862 gnd.n5666 gnd.n5665 585
R11863 gnd.n5667 gnd.n5666 585
R11864 gnd.n1001 gnd.n1000 585
R11865 gnd.n5598 gnd.n1000 585
R11866 gnd.n5661 gnd.n5660 585
R11867 gnd.n5660 gnd.n5659 585
R11868 gnd.n1004 gnd.n1003 585
R11869 gnd.n5649 gnd.n1004 585
R11870 gnd.n5626 gnd.n5625 585
R11871 gnd.n5627 gnd.n5626 585
R11872 gnd.n1074 gnd.n1073 585
R11873 gnd.n1073 gnd.n1070 585
R11874 gnd.n5621 gnd.n5620 585
R11875 gnd.n5620 gnd.n5619 585
R11876 gnd.n1077 gnd.n1076 585
R11877 gnd.n5061 gnd.n1077 585
R11878 gnd.n5154 gnd.n5153 585
R11879 gnd.n5153 gnd.n5152 585
R11880 gnd.n5059 gnd.n5058 585
R11881 gnd.n5140 gnd.n5059 585
R11882 gnd.n5158 gnd.n5057 585
R11883 gnd.n5068 gnd.n5057 585
R11884 gnd.n5159 gnd.n5056 585
R11885 gnd.n5130 gnd.n5056 585
R11886 gnd.n5160 gnd.n5055 585
R11887 gnd.n5075 gnd.n5055 585
R11888 gnd.n5118 gnd.n5053 585
R11889 gnd.n5119 gnd.n5118 585
R11890 gnd.n5164 gnd.n5052 585
R11891 gnd.n5081 gnd.n5052 585
R11892 gnd.n5165 gnd.n5051 585
R11893 gnd.n5109 gnd.n5051 585
R11894 gnd.n5166 gnd.n5050 585
R11895 gnd.n5087 gnd.n5050 585
R11896 gnd.n5047 gnd.n5045 585
R11897 gnd.n5095 gnd.n5045 585
R11898 gnd.n5171 gnd.n5170 585
R11899 gnd.n5172 gnd.n5171 585
R11900 gnd.n5046 gnd.n1262 585
R11901 gnd.n5174 gnd.n1262 585
R11902 gnd.n5328 gnd.n5327 585
R11903 gnd.n5326 gnd.n1261 585
R11904 gnd.n1264 gnd.n1260 585
R11905 gnd.n5330 gnd.n1260 585
R11906 gnd.n5322 gnd.n1266 585
R11907 gnd.n5321 gnd.n1267 585
R11908 gnd.n5320 gnd.n1268 585
R11909 gnd.n5317 gnd.n1269 585
R11910 gnd.n5316 gnd.n1270 585
R11911 gnd.n5196 gnd.n1271 585
R11912 gnd.n5198 gnd.n5197 585
R11913 gnd.n5308 gnd.n5199 585
R11914 gnd.n5307 gnd.n5200 585
R11915 gnd.n5210 gnd.n5201 585
R11916 gnd.n5300 gnd.n5211 585
R11917 gnd.n5299 gnd.n5212 585
R11918 gnd.n5214 gnd.n5213 585
R11919 gnd.n5292 gnd.n5222 585
R11920 gnd.n5291 gnd.n5223 585
R11921 gnd.n5233 gnd.n5224 585
R11922 gnd.n5284 gnd.n5234 585
R11923 gnd.n5283 gnd.n5235 585
R11924 gnd.n5237 gnd.n5236 585
R11925 gnd.n5276 gnd.n5245 585
R11926 gnd.n5275 gnd.n5246 585
R11927 gnd.n5266 gnd.n5247 585
R11928 gnd.n5268 gnd.n5267 585
R11929 gnd.n1257 gnd.n1242 585
R11930 gnd.n5334 gnd.n1243 585
R11931 gnd.n5333 gnd.n5332 585
R11932 gnd.n581 gnd.n426 585
R11933 gnd.n6463 gnd.n426 585
R11934 gnd.n6440 gnd.n6439 585
R11935 gnd.n6441 gnd.n6440 585
R11936 gnd.n580 gnd.n579 585
R11937 gnd.n588 gnd.n579 585
R11938 gnd.n6434 gnd.n6433 585
R11939 gnd.n6433 gnd.n6432 585
R11940 gnd.n584 gnd.n583 585
R11941 gnd.n597 gnd.n584 585
R11942 gnd.n607 gnd.n596 585
R11943 gnd.n6423 gnd.n596 585
R11944 gnd.n6410 gnd.n6409 585
R11945 gnd.n6411 gnd.n6410 585
R11946 gnd.n606 gnd.n605 585
R11947 gnd.n605 gnd.n604 585
R11948 gnd.n6404 gnd.n6403 585
R11949 gnd.n6403 gnd.n6402 585
R11950 gnd.n610 gnd.n609 585
R11951 gnd.n622 gnd.n610 585
R11952 gnd.n632 gnd.n621 585
R11953 gnd.n6393 gnd.n621 585
R11954 gnd.n6380 gnd.n6379 585
R11955 gnd.n6381 gnd.n6380 585
R11956 gnd.n631 gnd.n630 585
R11957 gnd.n630 gnd.n629 585
R11958 gnd.n6374 gnd.n6373 585
R11959 gnd.n6373 gnd.n6372 585
R11960 gnd.n635 gnd.n634 585
R11961 gnd.n647 gnd.n635 585
R11962 gnd.n6019 gnd.n646 585
R11963 gnd.n6363 gnd.n646 585
R11964 gnd.n6020 gnd.n655 585
R11965 gnd.n6351 gnd.n655 585
R11966 gnd.n6017 gnd.n6016 585
R11967 gnd.n6016 gnd.n654 585
R11968 gnd.n6024 gnd.n6015 585
R11969 gnd.n6015 gnd.n701 585
R11970 gnd.n6025 gnd.n6014 585
R11971 gnd.n6014 gnd.n698 585
R11972 gnd.n6026 gnd.n708 585
R11973 gnd.n6179 gnd.n708 585
R11974 gnd.n6012 gnd.n6011 585
R11975 gnd.n6011 gnd.n6010 585
R11976 gnd.n6030 gnd.n717 585
R11977 gnd.n6164 gnd.n717 585
R11978 gnd.n6031 gnd.n726 585
R11979 gnd.n6151 gnd.n726 585
R11980 gnd.n6032 gnd.n735 585
R11981 gnd.n6140 gnd.n735 585
R11982 gnd.n5965 gnd.n5964 585
R11983 gnd.n5964 gnd.n744 585
R11984 gnd.n6036 gnd.n742 585
R11985 gnd.n6132 gnd.n742 585
R11986 gnd.n6037 gnd.n5963 585
R11987 gnd.n5963 gnd.n749 585
R11988 gnd.n6038 gnd.n5962 585
R11989 gnd.n5962 gnd.n758 585
R11990 gnd.n5960 gnd.n763 585
R11991 gnd.n6106 gnd.n763 585
R11992 gnd.n6042 gnd.n5959 585
R11993 gnd.n5976 gnd.n5959 585
R11994 gnd.n6043 gnd.n772 585
R11995 gnd.n6097 gnd.n772 585
R11996 gnd.n6044 gnd.n778 585
R11997 gnd.n6089 gnd.n778 585
R11998 gnd.n809 gnd.n786 585
R11999 gnd.n6077 gnd.n786 585
R12000 gnd.n6049 gnd.n6048 585
R12001 gnd.n6050 gnd.n6049 585
R12002 gnd.n808 gnd.n795 585
R12003 gnd.n6069 gnd.n795 585
R12004 gnd.n5955 gnd.n804 585
R12005 gnd.n6058 gnd.n804 585
R12006 gnd.n5954 gnd.n5953 585
R12007 gnd.n5953 gnd.n5952 585
R12008 gnd.n812 gnd.n811 585
R12009 gnd.n824 gnd.n812 585
R12010 gnd.n5824 gnd.n819 585
R12011 gnd.n5944 gnd.n819 585
R12012 gnd.n5828 gnd.n5823 585
R12013 gnd.n5823 gnd.n832 585
R12014 gnd.n5829 gnd.n837 585
R12015 gnd.n5908 gnd.n837 585
R12016 gnd.n5830 gnd.n847 585
R12017 gnd.n5900 gnd.n847 585
R12018 gnd.n5821 gnd.n5820 585
R12019 gnd.n5820 gnd.n5819 585
R12020 gnd.n5834 gnd.n856 585
R12021 gnd.n5891 gnd.n856 585
R12022 gnd.n5835 gnd.n864 585
R12023 gnd.n5883 gnd.n864 585
R12024 gnd.n5836 gnd.n879 585
R12025 gnd.n5850 gnd.n879 585
R12026 gnd.n889 gnd.n887 585
R12027 gnd.n887 gnd.n871 585
R12028 gnd.n5841 gnd.n5840 585
R12029 gnd.n5842 gnd.n5841 585
R12030 gnd.n888 gnd.n886 585
R12031 gnd.n5782 gnd.n886 585
R12032 gnd.n5808 gnd.n5807 585
R12033 gnd.n5807 gnd.n5806 585
R12034 gnd.n892 gnd.n891 585
R12035 gnd.n909 gnd.n892 585
R12036 gnd.n951 gnd.n901 585
R12037 gnd.n5798 gnd.n901 585
R12038 gnd.n5738 gnd.n5737 585
R12039 gnd.n5740 gnd.n5738 585
R12040 gnd.n950 gnd.n926 585
R12041 gnd.n5764 gnd.n926 585
R12042 gnd.n5732 gnd.n5731 585
R12043 gnd.n5731 gnd.n941 585
R12044 gnd.n5730 gnd.n933 585
R12045 gnd.n5756 gnd.n933 585
R12046 gnd.n5729 gnd.n954 585
R12047 gnd.n5681 gnd.n954 585
R12048 gnd.n958 gnd.n953 585
R12049 gnd.n5705 gnd.n958 585
R12050 gnd.n5725 gnd.n5724 585
R12051 gnd.n5724 gnd.n5723 585
R12052 gnd.n957 gnd.n956 585
R12053 gnd.n5693 gnd.n957 585
R12054 gnd.n5604 gnd.n969 585
R12055 gnd.n5714 gnd.n969 585
R12056 gnd.n5605 gnd.n5602 585
R12057 gnd.n5602 gnd.n992 585
R12058 gnd.n5606 gnd.n998 585
R12059 gnd.n5667 gnd.n998 585
R12060 gnd.n5600 gnd.n5599 585
R12061 gnd.n5599 gnd.n5598 585
R12062 gnd.n5610 gnd.n1005 585
R12063 gnd.n5659 gnd.n1005 585
R12064 gnd.n5611 gnd.n1063 585
R12065 gnd.n5649 gnd.n1063 585
R12066 gnd.n5612 gnd.n1071 585
R12067 gnd.n5627 gnd.n1071 585
R12068 gnd.n1082 gnd.n1080 585
R12069 gnd.n1080 gnd.n1070 585
R12070 gnd.n5617 gnd.n5616 585
R12071 gnd.n5619 gnd.n5617 585
R12072 gnd.n1081 gnd.n1079 585
R12073 gnd.n5061 gnd.n1079 585
R12074 gnd.n5071 gnd.n5060 585
R12075 gnd.n5152 gnd.n5060 585
R12076 gnd.n5138 gnd.n5137 585
R12077 gnd.n5140 gnd.n5138 585
R12078 gnd.n5070 gnd.n5069 585
R12079 gnd.n5069 gnd.n5068 585
R12080 gnd.n5132 gnd.n5131 585
R12081 gnd.n5131 gnd.n5130 585
R12082 gnd.n5074 gnd.n5073 585
R12083 gnd.n5075 gnd.n5074 585
R12084 gnd.n5116 gnd.n5115 585
R12085 gnd.n5119 gnd.n5116 585
R12086 gnd.n5083 gnd.n5082 585
R12087 gnd.n5082 gnd.n5081 585
R12088 gnd.n5111 gnd.n5110 585
R12089 gnd.n5110 gnd.n5109 585
R12090 gnd.n5086 gnd.n5085 585
R12091 gnd.n5087 gnd.n5086 585
R12092 gnd.n5094 gnd.n5093 585
R12093 gnd.n5095 gnd.n5094 585
R12094 gnd.n5088 gnd.n5043 585
R12095 gnd.n5172 gnd.n5043 585
R12096 gnd.n5089 gnd.n1244 585
R12097 gnd.n5174 gnd.n1244 585
R12098 gnd.n6703 gnd.n6702 585
R12099 gnd.n6704 gnd.n6703 585
R12100 gnd.n445 gnd.n443 585
R12101 gnd.n6530 gnd.n6529 585
R12102 gnd.n6540 gnd.n6528 585
R12103 gnd.n6541 gnd.n6527 585
R12104 gnd.n6526 gnd.n6518 585
R12105 gnd.n6548 gnd.n6517 585
R12106 gnd.n6549 gnd.n6516 585
R12107 gnd.n6510 gnd.n6509 585
R12108 gnd.n6556 gnd.n6508 585
R12109 gnd.n6557 gnd.n6507 585
R12110 gnd.n6506 gnd.n6498 585
R12111 gnd.n6564 gnd.n6497 585
R12112 gnd.n6565 gnd.n6496 585
R12113 gnd.n6487 gnd.n6486 585
R12114 gnd.n6572 gnd.n6485 585
R12115 gnd.n6573 gnd.n6484 585
R12116 gnd.n6574 gnd.n6483 585
R12117 gnd.n6482 gnd.n6481 585
R12118 gnd.n6480 gnd.n6479 585
R12119 gnd.n6473 gnd.n565 585
R12120 gnd.n6475 gnd.n6474 585
R12121 gnd.n6472 gnd.n6471 585
R12122 gnd.n6470 gnd.n6469 585
R12123 gnd.n571 gnd.n567 585
R12124 gnd.n6707 gnd.n6706 585
R12125 gnd.n6708 gnd.n425 585
R12126 gnd.n440 gnd.n424 585
R12127 gnd.n450 gnd.n444 585
R12128 gnd.n1085 gnd.t109 543.808
R12129 gnd.n690 gnd.t22 543.808
R12130 gnd.n1087 gnd.t41 543.808
R12131 gnd.n6212 gnd.t73 543.808
R12132 gnd.n6281 gnd.n695 478.086
R12133 gnd.n6284 gnd.n6283 478.086
R12134 gnd.n5590 gnd.n1006 478.086
R12135 gnd.n5657 gnd.n1008 478.086
R12136 gnd.n1687 gnd.n1680 476.536
R12137 gnd.n5263 gnd.t63 371.625
R12138 gnd.n6696 gnd.t101 371.625
R12139 gnd.n5254 gnd.t122 371.625
R12140 gnd.n515 gnd.t98 371.625
R12141 gnd.n538 gnd.t88 371.625
R12142 gnd.n561 gnd.t34 371.625
R12143 gnd.n7132 gnd.t38 371.625
R12144 gnd.n7111 gnd.t30 371.625
R12145 gnd.n7218 gnd.t91 371.625
R12146 gnd.n180 gnd.t119 371.625
R12147 gnd.n4470 gnd.t70 371.625
R12148 gnd.n4492 gnd.t45 371.625
R12149 gnd.n4514 gnd.t76 371.625
R12150 gnd.n4542 gnd.t26 371.625
R12151 gnd.n5392 gnd.t116 371.625
R12152 gnd.n1202 gnd.t48 371.625
R12153 gnd.n1169 gnd.t79 371.625
R12154 gnd.n446 gnd.t52 371.625
R12155 gnd.n7040 gnd.n242 368.923
R12156 gnd.n3445 gnd.t59 323.425
R12157 gnd.n3066 gnd.t94 323.425
R12158 gnd.n2377 gnd.n2376 299.933
R12159 gnd.n2376 gnd.n2047 299.933
R12160 gnd.n2368 gnd.n2047 299.933
R12161 gnd.n2368 gnd.n2367 299.933
R12162 gnd.n2367 gnd.n2366 299.933
R12163 gnd.n2366 gnd.n2055 299.933
R12164 gnd.n2360 gnd.n2055 299.933
R12165 gnd.n2360 gnd.n2359 299.933
R12166 gnd.n2359 gnd.n2358 299.933
R12167 gnd.n2358 gnd.n2062 299.933
R12168 gnd.n2352 gnd.n2062 299.933
R12169 gnd.n2352 gnd.n2351 299.933
R12170 gnd.n2351 gnd.n2350 299.933
R12171 gnd.n2350 gnd.n2070 299.933
R12172 gnd.n2344 gnd.n2070 299.933
R12173 gnd.n2344 gnd.n2343 299.933
R12174 gnd.n2343 gnd.n2342 299.933
R12175 gnd.n2342 gnd.n2078 299.933
R12176 gnd.n2336 gnd.n2078 299.933
R12177 gnd.n2336 gnd.n2335 299.933
R12178 gnd.n2335 gnd.n2334 299.933
R12179 gnd.n2334 gnd.n2086 299.933
R12180 gnd.n2328 gnd.n2086 299.933
R12181 gnd.n2328 gnd.n2327 299.933
R12182 gnd.n2327 gnd.n2326 299.933
R12183 gnd.n2326 gnd.n2094 299.933
R12184 gnd.n2320 gnd.n2094 299.933
R12185 gnd.n2320 gnd.n2319 299.933
R12186 gnd.n2319 gnd.n2318 299.933
R12187 gnd.n2318 gnd.n2102 299.933
R12188 gnd.n2312 gnd.n2102 299.933
R12189 gnd.n2312 gnd.n2311 299.933
R12190 gnd.n2311 gnd.n2310 299.933
R12191 gnd.n2310 gnd.n2110 299.933
R12192 gnd.n2304 gnd.n2110 299.933
R12193 gnd.n2304 gnd.n2303 299.933
R12194 gnd.n2303 gnd.n2302 299.933
R12195 gnd.n2302 gnd.n2118 299.933
R12196 gnd.n2296 gnd.n2118 299.933
R12197 gnd.n2296 gnd.n2295 299.933
R12198 gnd.n2295 gnd.n2294 299.933
R12199 gnd.n2294 gnd.n2126 299.933
R12200 gnd.n2288 gnd.n2126 299.933
R12201 gnd.n2288 gnd.n2287 299.933
R12202 gnd.n2287 gnd.n2286 299.933
R12203 gnd.n2286 gnd.n2134 299.933
R12204 gnd.n2280 gnd.n2134 299.933
R12205 gnd.n2280 gnd.n2279 299.933
R12206 gnd.n2279 gnd.n2278 299.933
R12207 gnd.n2278 gnd.n2142 299.933
R12208 gnd.n2272 gnd.n2142 299.933
R12209 gnd.n2272 gnd.n2271 299.933
R12210 gnd.n2271 gnd.n2270 299.933
R12211 gnd.n2270 gnd.n2150 299.933
R12212 gnd.n2264 gnd.n2150 299.933
R12213 gnd.n2264 gnd.n2263 299.933
R12214 gnd.n2263 gnd.n2262 299.933
R12215 gnd.n2262 gnd.n2158 299.933
R12216 gnd.n2256 gnd.n2158 299.933
R12217 gnd.n2256 gnd.n2255 299.933
R12218 gnd.n2255 gnd.n2254 299.933
R12219 gnd.n2254 gnd.n2166 299.933
R12220 gnd.n2248 gnd.n2166 299.933
R12221 gnd.n2248 gnd.n2247 299.933
R12222 gnd.n2247 gnd.n2246 299.933
R12223 gnd.n2246 gnd.n2174 299.933
R12224 gnd.n2240 gnd.n2174 299.933
R12225 gnd.n2240 gnd.n2239 299.933
R12226 gnd.n2239 gnd.n2238 299.933
R12227 gnd.n2238 gnd.n2182 299.933
R12228 gnd.n2232 gnd.n2182 299.933
R12229 gnd.n2232 gnd.n2231 299.933
R12230 gnd.n2231 gnd.n2230 299.933
R12231 gnd.n2230 gnd.n2190 299.933
R12232 gnd.n2224 gnd.n2190 299.933
R12233 gnd.n2224 gnd.n2223 299.933
R12234 gnd.n2223 gnd.n2222 299.933
R12235 gnd.n2222 gnd.n2198 299.933
R12236 gnd.n2216 gnd.n2198 299.933
R12237 gnd.n2216 gnd.n2215 299.933
R12238 gnd.n2215 gnd.n2214 299.933
R12239 gnd.n2214 gnd.n2206 299.933
R12240 gnd.n2206 gnd.n242 299.933
R12241 gnd.n4223 gnd.n4197 289.615
R12242 gnd.n4191 gnd.n4165 289.615
R12243 gnd.n4159 gnd.n4133 289.615
R12244 gnd.n4128 gnd.n4102 289.615
R12245 gnd.n4096 gnd.n4070 289.615
R12246 gnd.n4064 gnd.n4038 289.615
R12247 gnd.n4032 gnd.n4006 289.615
R12248 gnd.n4001 gnd.n3975 289.615
R12249 gnd.n3519 gnd.t125 279.217
R12250 gnd.n3110 gnd.t112 279.217
R12251 gnd.n1015 gnd.t134 260.649
R12252 gnd.n6204 gnd.t84 260.649
R12253 gnd.n5651 gnd.n5650 256.663
R12254 gnd.n5650 gnd.n1031 256.663
R12255 gnd.n5650 gnd.n1032 256.663
R12256 gnd.n5650 gnd.n1033 256.663
R12257 gnd.n5650 gnd.n1034 256.663
R12258 gnd.n5650 gnd.n1035 256.663
R12259 gnd.n5650 gnd.n1036 256.663
R12260 gnd.n5650 gnd.n1037 256.663
R12261 gnd.n5650 gnd.n1038 256.663
R12262 gnd.n5650 gnd.n1039 256.663
R12263 gnd.n5650 gnd.n1040 256.663
R12264 gnd.n5650 gnd.n1041 256.663
R12265 gnd.n5650 gnd.n1042 256.663
R12266 gnd.n5650 gnd.n1043 256.663
R12267 gnd.n5650 gnd.n1044 256.663
R12268 gnd.n5650 gnd.n1045 256.663
R12269 gnd.n5525 gnd.n5524 256.663
R12270 gnd.n5650 gnd.n1046 256.663
R12271 gnd.n5650 gnd.n1047 256.663
R12272 gnd.n5650 gnd.n1048 256.663
R12273 gnd.n5650 gnd.n1049 256.663
R12274 gnd.n5650 gnd.n1050 256.663
R12275 gnd.n5650 gnd.n1051 256.663
R12276 gnd.n5650 gnd.n1052 256.663
R12277 gnd.n5650 gnd.n1053 256.663
R12278 gnd.n5650 gnd.n1054 256.663
R12279 gnd.n5650 gnd.n1055 256.663
R12280 gnd.n5650 gnd.n1056 256.663
R12281 gnd.n5650 gnd.n1057 256.663
R12282 gnd.n5650 gnd.n1058 256.663
R12283 gnd.n5650 gnd.n1059 256.663
R12284 gnd.n5650 gnd.n1060 256.663
R12285 gnd.n5650 gnd.n1061 256.663
R12286 gnd.n5650 gnd.n1062 256.663
R12287 gnd.n6350 gnd.n673 256.663
R12288 gnd.n6350 gnd.n674 256.663
R12289 gnd.n6350 gnd.n675 256.663
R12290 gnd.n6350 gnd.n676 256.663
R12291 gnd.n6350 gnd.n677 256.663
R12292 gnd.n6350 gnd.n678 256.663
R12293 gnd.n6350 gnd.n679 256.663
R12294 gnd.n6350 gnd.n680 256.663
R12295 gnd.n6350 gnd.n681 256.663
R12296 gnd.n6350 gnd.n682 256.663
R12297 gnd.n6350 gnd.n683 256.663
R12298 gnd.n6350 gnd.n684 256.663
R12299 gnd.n6350 gnd.n685 256.663
R12300 gnd.n6350 gnd.n686 256.663
R12301 gnd.n6350 gnd.n687 256.663
R12302 gnd.n6350 gnd.n688 256.663
R12303 gnd.n689 gnd.n525 256.663
R12304 gnd.n6350 gnd.n672 256.663
R12305 gnd.n6350 gnd.n671 256.663
R12306 gnd.n6350 gnd.n670 256.663
R12307 gnd.n6350 gnd.n669 256.663
R12308 gnd.n6350 gnd.n668 256.663
R12309 gnd.n6350 gnd.n667 256.663
R12310 gnd.n6350 gnd.n666 256.663
R12311 gnd.n6350 gnd.n665 256.663
R12312 gnd.n6350 gnd.n664 256.663
R12313 gnd.n6350 gnd.n663 256.663
R12314 gnd.n6350 gnd.n662 256.663
R12315 gnd.n6350 gnd.n661 256.663
R12316 gnd.n6350 gnd.n660 256.663
R12317 gnd.n6350 gnd.n659 256.663
R12318 gnd.n6350 gnd.n658 256.663
R12319 gnd.n6350 gnd.n657 256.663
R12320 gnd.n6350 gnd.n656 256.663
R12321 gnd.n4703 gnd.n1545 242.672
R12322 gnd.n4703 gnd.n1546 242.672
R12323 gnd.n4703 gnd.n1547 242.672
R12324 gnd.n4703 gnd.n1548 242.672
R12325 gnd.n4703 gnd.n1549 242.672
R12326 gnd.n4703 gnd.n1550 242.672
R12327 gnd.n4703 gnd.n1551 242.672
R12328 gnd.n4703 gnd.n1552 242.672
R12329 gnd.n4703 gnd.n1553 242.672
R12330 gnd.n5257 gnd.n1156 242.672
R12331 gnd.n5252 gnd.n1156 242.672
R12332 gnd.n5249 gnd.n1156 242.672
R12333 gnd.n5240 gnd.n1156 242.672
R12334 gnd.n5229 gnd.n1156 242.672
R12335 gnd.n5226 gnd.n1156 242.672
R12336 gnd.n5217 gnd.n1156 242.672
R12337 gnd.n5206 gnd.n1156 242.672
R12338 gnd.n5203 gnd.n1156 242.672
R12339 gnd.n3573 gnd.n3572 242.672
R12340 gnd.n3573 gnd.n3483 242.672
R12341 gnd.n3573 gnd.n3484 242.672
R12342 gnd.n3573 gnd.n3485 242.672
R12343 gnd.n3573 gnd.n3486 242.672
R12344 gnd.n3573 gnd.n3487 242.672
R12345 gnd.n3573 gnd.n3488 242.672
R12346 gnd.n3573 gnd.n3489 242.672
R12347 gnd.n3573 gnd.n3490 242.672
R12348 gnd.n3573 gnd.n3491 242.672
R12349 gnd.n3573 gnd.n3492 242.672
R12350 gnd.n3573 gnd.n3493 242.672
R12351 gnd.n3574 gnd.n3573 242.672
R12352 gnd.n4279 gnd.n3036 242.672
R12353 gnd.n4285 gnd.n3036 242.672
R12354 gnd.n3113 gnd.n3036 242.672
R12355 gnd.n4292 gnd.n3036 242.672
R12356 gnd.n3104 gnd.n3036 242.672
R12357 gnd.n4299 gnd.n3036 242.672
R12358 gnd.n3097 gnd.n3036 242.672
R12359 gnd.n4306 gnd.n3036 242.672
R12360 gnd.n3090 gnd.n3036 242.672
R12361 gnd.n4313 gnd.n3036 242.672
R12362 gnd.n3083 gnd.n3036 242.672
R12363 gnd.n4320 gnd.n3036 242.672
R12364 gnd.n3076 gnd.n3036 242.672
R12365 gnd.n6693 gnd.n486 242.672
R12366 gnd.n6693 gnd.n487 242.672
R12367 gnd.n6693 gnd.n488 242.672
R12368 gnd.n6693 gnd.n489 242.672
R12369 gnd.n6693 gnd.n490 242.672
R12370 gnd.n6693 gnd.n491 242.672
R12371 gnd.n6693 gnd.n492 242.672
R12372 gnd.n6693 gnd.n494 242.672
R12373 gnd.n6694 gnd.n6693 242.672
R12374 gnd.n7254 gnd.n7253 242.672
R12375 gnd.n7253 gnd.n241 242.672
R12376 gnd.n7253 gnd.n190 242.672
R12377 gnd.n7253 gnd.n189 242.672
R12378 gnd.n7253 gnd.n188 242.672
R12379 gnd.n7253 gnd.n187 242.672
R12380 gnd.n7253 gnd.n186 242.672
R12381 gnd.n7253 gnd.n185 242.672
R12382 gnd.n7253 gnd.n184 242.672
R12383 gnd.n3657 gnd.n3656 242.672
R12384 gnd.n3656 gnd.n3395 242.672
R12385 gnd.n3656 gnd.n3396 242.672
R12386 gnd.n3656 gnd.n3397 242.672
R12387 gnd.n3656 gnd.n3398 242.672
R12388 gnd.n3656 gnd.n3399 242.672
R12389 gnd.n3656 gnd.n3400 242.672
R12390 gnd.n3656 gnd.n3401 242.672
R12391 gnd.n4331 gnd.n3036 242.672
R12392 gnd.n3069 gnd.n3036 242.672
R12393 gnd.n4338 gnd.n3036 242.672
R12394 gnd.n3060 gnd.n3036 242.672
R12395 gnd.n4345 gnd.n3036 242.672
R12396 gnd.n3053 gnd.n3036 242.672
R12397 gnd.n4352 gnd.n3036 242.672
R12398 gnd.n3046 gnd.n3036 242.672
R12399 gnd.n4704 gnd.n4703 242.672
R12400 gnd.n4703 gnd.n1517 242.672
R12401 gnd.n4703 gnd.n1518 242.672
R12402 gnd.n4703 gnd.n1519 242.672
R12403 gnd.n4703 gnd.n1520 242.672
R12404 gnd.n4703 gnd.n1521 242.672
R12405 gnd.n4703 gnd.n1522 242.672
R12406 gnd.n4703 gnd.n1523 242.672
R12407 gnd.n4703 gnd.n1524 242.672
R12408 gnd.n4703 gnd.n1525 242.672
R12409 gnd.n4703 gnd.n1526 242.672
R12410 gnd.n4703 gnd.n1527 242.672
R12411 gnd.n4703 gnd.n1528 242.672
R12412 gnd.n4703 gnd.n1529 242.672
R12413 gnd.n4703 gnd.n1530 242.672
R12414 gnd.n4703 gnd.n1531 242.672
R12415 gnd.n4703 gnd.n1532 242.672
R12416 gnd.n4703 gnd.n1533 242.672
R12417 gnd.n4703 gnd.n1534 242.672
R12418 gnd.n4703 gnd.n1535 242.672
R12419 gnd.n4703 gnd.n1536 242.672
R12420 gnd.n4703 gnd.n1537 242.672
R12421 gnd.n4703 gnd.n1538 242.672
R12422 gnd.n4703 gnd.n1539 242.672
R12423 gnd.n4703 gnd.n1540 242.672
R12424 gnd.n4703 gnd.n1541 242.672
R12425 gnd.n4703 gnd.n1542 242.672
R12426 gnd.n4703 gnd.n1543 242.672
R12427 gnd.n4703 gnd.n1544 242.672
R12428 gnd.n5467 gnd.n1156 242.672
R12429 gnd.n1205 gnd.n1156 242.672
R12430 gnd.n5474 gnd.n1156 242.672
R12431 gnd.n1196 gnd.n1156 242.672
R12432 gnd.n5481 gnd.n1156 242.672
R12433 gnd.n1189 gnd.n1156 242.672
R12434 gnd.n5488 gnd.n1156 242.672
R12435 gnd.n1182 gnd.n1156 242.672
R12436 gnd.n5495 gnd.n1156 242.672
R12437 gnd.n5498 gnd.n1156 242.672
R12438 gnd.n1173 gnd.n1156 242.672
R12439 gnd.n5507 gnd.n1156 242.672
R12440 gnd.n1164 gnd.n1156 242.672
R12441 gnd.n5514 gnd.n1156 242.672
R12442 gnd.n5517 gnd.n1156 242.672
R12443 gnd.n1156 gnd.n1155 242.672
R12444 gnd.n5523 gnd.n1150 242.672
R12445 gnd.n5407 gnd.n1156 242.672
R12446 gnd.n5406 gnd.n1156 242.672
R12447 gnd.n5414 gnd.n1156 242.672
R12448 gnd.n5400 gnd.n1156 242.672
R12449 gnd.n5421 gnd.n1156 242.672
R12450 gnd.n5390 gnd.n1156 242.672
R12451 gnd.n5428 gnd.n1156 242.672
R12452 gnd.n5383 gnd.n1156 242.672
R12453 gnd.n5435 gnd.n1156 242.672
R12454 gnd.n5376 gnd.n1156 242.672
R12455 gnd.n5442 gnd.n1156 242.672
R12456 gnd.n5369 gnd.n1156 242.672
R12457 gnd.n5449 gnd.n1156 242.672
R12458 gnd.n6693 gnd.n6692 242.672
R12459 gnd.n6693 gnd.n458 242.672
R12460 gnd.n6693 gnd.n459 242.672
R12461 gnd.n6693 gnd.n460 242.672
R12462 gnd.n6693 gnd.n461 242.672
R12463 gnd.n6693 gnd.n462 242.672
R12464 gnd.n6693 gnd.n463 242.672
R12465 gnd.n6693 gnd.n464 242.672
R12466 gnd.n6693 gnd.n465 242.672
R12467 gnd.n6693 gnd.n466 242.672
R12468 gnd.n6693 gnd.n467 242.672
R12469 gnd.n6693 gnd.n468 242.672
R12470 gnd.n6693 gnd.n469 242.672
R12471 gnd.n6640 gnd.n526 242.672
R12472 gnd.n6693 gnd.n470 242.672
R12473 gnd.n6693 gnd.n471 242.672
R12474 gnd.n6693 gnd.n472 242.672
R12475 gnd.n6693 gnd.n473 242.672
R12476 gnd.n6693 gnd.n474 242.672
R12477 gnd.n6693 gnd.n475 242.672
R12478 gnd.n6693 gnd.n476 242.672
R12479 gnd.n6693 gnd.n477 242.672
R12480 gnd.n6693 gnd.n478 242.672
R12481 gnd.n6693 gnd.n479 242.672
R12482 gnd.n6693 gnd.n480 242.672
R12483 gnd.n6693 gnd.n481 242.672
R12484 gnd.n6693 gnd.n482 242.672
R12485 gnd.n6693 gnd.n483 242.672
R12486 gnd.n6693 gnd.n484 242.672
R12487 gnd.n6693 gnd.n485 242.672
R12488 gnd.n7253 gnd.n7041 242.672
R12489 gnd.n7253 gnd.n7042 242.672
R12490 gnd.n7253 gnd.n7043 242.672
R12491 gnd.n7253 gnd.n7044 242.672
R12492 gnd.n7253 gnd.n7045 242.672
R12493 gnd.n7253 gnd.n7046 242.672
R12494 gnd.n7253 gnd.n7047 242.672
R12495 gnd.n7253 gnd.n7048 242.672
R12496 gnd.n7253 gnd.n7049 242.672
R12497 gnd.n7253 gnd.n7050 242.672
R12498 gnd.n7253 gnd.n7051 242.672
R12499 gnd.n7253 gnd.n7052 242.672
R12500 gnd.n7253 gnd.n7053 242.672
R12501 gnd.n7253 gnd.n7054 242.672
R12502 gnd.n7253 gnd.n7055 242.672
R12503 gnd.n7253 gnd.n7056 242.672
R12504 gnd.n7253 gnd.n7057 242.672
R12505 gnd.n7253 gnd.n7058 242.672
R12506 gnd.n7253 gnd.n7059 242.672
R12507 gnd.n7253 gnd.n7060 242.672
R12508 gnd.n7253 gnd.n7061 242.672
R12509 gnd.n7253 gnd.n7062 242.672
R12510 gnd.n7253 gnd.n7063 242.672
R12511 gnd.n7253 gnd.n7064 242.672
R12512 gnd.n7253 gnd.n7065 242.672
R12513 gnd.n7253 gnd.n7066 242.672
R12514 gnd.n7253 gnd.n7067 242.672
R12515 gnd.n7253 gnd.n7068 242.672
R12516 gnd.n7253 gnd.n7252 242.672
R12517 gnd.n5330 gnd.n5329 242.672
R12518 gnd.n5330 gnd.n1246 242.672
R12519 gnd.n5330 gnd.n1247 242.672
R12520 gnd.n5330 gnd.n1248 242.672
R12521 gnd.n5330 gnd.n1249 242.672
R12522 gnd.n5330 gnd.n1250 242.672
R12523 gnd.n5330 gnd.n1251 242.672
R12524 gnd.n5330 gnd.n1252 242.672
R12525 gnd.n5330 gnd.n1253 242.672
R12526 gnd.n5330 gnd.n1254 242.672
R12527 gnd.n5330 gnd.n1255 242.672
R12528 gnd.n5330 gnd.n1256 242.672
R12529 gnd.n5330 gnd.n1258 242.672
R12530 gnd.n5331 gnd.n5330 242.672
R12531 gnd.n6704 gnd.n439 242.672
R12532 gnd.n6704 gnd.n438 242.672
R12533 gnd.n6704 gnd.n437 242.672
R12534 gnd.n6704 gnd.n436 242.672
R12535 gnd.n6704 gnd.n435 242.672
R12536 gnd.n6704 gnd.n434 242.672
R12537 gnd.n6704 gnd.n433 242.672
R12538 gnd.n6704 gnd.n432 242.672
R12539 gnd.n6704 gnd.n431 242.672
R12540 gnd.n6704 gnd.n430 242.672
R12541 gnd.n6704 gnd.n429 242.672
R12542 gnd.n6704 gnd.n428 242.672
R12543 gnd.n6705 gnd.n6704 242.672
R12544 gnd.n6704 gnd.n441 242.672
R12545 gnd.n7069 gnd.n167 240.244
R12546 gnd.n7251 gnd.n7070 240.244
R12547 gnd.n7247 gnd.n7246 240.244
R12548 gnd.n7243 gnd.n7242 240.244
R12549 gnd.n7239 gnd.n7238 240.244
R12550 gnd.n7235 gnd.n7234 240.244
R12551 gnd.n7231 gnd.n7230 240.244
R12552 gnd.n7227 gnd.n7226 240.244
R12553 gnd.n7223 gnd.n7222 240.244
R12554 gnd.n7216 gnd.n7215 240.244
R12555 gnd.n7212 gnd.n7211 240.244
R12556 gnd.n7208 gnd.n7207 240.244
R12557 gnd.n7204 gnd.n7203 240.244
R12558 gnd.n7200 gnd.n7199 240.244
R12559 gnd.n7196 gnd.n7195 240.244
R12560 gnd.n7192 gnd.n7191 240.244
R12561 gnd.n7188 gnd.n7187 240.244
R12562 gnd.n7184 gnd.n7183 240.244
R12563 gnd.n7180 gnd.n7179 240.244
R12564 gnd.n7173 gnd.n7172 240.244
R12565 gnd.n7170 gnd.n7169 240.244
R12566 gnd.n7166 gnd.n7165 240.244
R12567 gnd.n7162 gnd.n7161 240.244
R12568 gnd.n7158 gnd.n7157 240.244
R12569 gnd.n7154 gnd.n7153 240.244
R12570 gnd.n7150 gnd.n7149 240.244
R12571 gnd.n7146 gnd.n7145 240.244
R12572 gnd.n7142 gnd.n7141 240.244
R12573 gnd.n7138 gnd.n7137 240.244
R12574 gnd.n419 gnd.n393 240.244
R12575 gnd.n6728 gnd.n393 240.244
R12576 gnd.n6728 gnd.n383 240.244
R12577 gnd.n409 gnd.n383 240.244
R12578 gnd.n409 gnd.n375 240.244
R12579 gnd.n375 gnd.n360 240.244
R12580 gnd.n6791 gnd.n360 240.244
R12581 gnd.n6791 gnd.n350 240.244
R12582 gnd.n350 gnd.n341 240.244
R12583 gnd.n6823 gnd.n341 240.244
R12584 gnd.n6823 gnd.n331 240.244
R12585 gnd.n6827 gnd.n331 240.244
R12586 gnd.n6827 gnd.n321 240.244
R12587 gnd.n321 gnd.n312 240.244
R12588 gnd.n6866 gnd.n312 240.244
R12589 gnd.n6866 gnd.n301 240.244
R12590 gnd.n6878 gnd.n301 240.244
R12591 gnd.n6878 gnd.n295 240.244
R12592 gnd.n295 gnd.n289 240.244
R12593 gnd.n289 gnd.n284 240.244
R12594 gnd.n284 gnd.n279 240.244
R12595 gnd.n6920 gnd.n279 240.244
R12596 gnd.n6920 gnd.n70 240.244
R12597 gnd.n272 gnd.n70 240.244
R12598 gnd.n272 gnd.n266 240.244
R12599 gnd.n266 gnd.n87 240.244
R12600 gnd.n6990 gnd.n87 240.244
R12601 gnd.n6990 gnd.n99 240.244
R12602 gnd.n6986 gnd.n99 240.244
R12603 gnd.n6986 gnd.n109 240.244
R12604 gnd.n6978 gnd.n109 240.244
R12605 gnd.n6978 gnd.n118 240.244
R12606 gnd.n6974 gnd.n118 240.244
R12607 gnd.n6974 gnd.n129 240.244
R12608 gnd.n6966 gnd.n129 240.244
R12609 gnd.n6966 gnd.n139 240.244
R12610 gnd.n6962 gnd.n139 240.244
R12611 gnd.n6962 gnd.n150 240.244
R12612 gnd.n6954 gnd.n150 240.244
R12613 gnd.n6954 gnd.n160 240.244
R12614 gnd.n7263 gnd.n160 240.244
R12615 gnd.n7263 gnd.n169 240.244
R12616 gnd.n496 gnd.n495 240.244
R12617 gnd.n6686 gnd.n495 240.244
R12618 gnd.n6684 gnd.n6683 240.244
R12619 gnd.n6680 gnd.n6679 240.244
R12620 gnd.n6676 gnd.n6675 240.244
R12621 gnd.n6672 gnd.n6671 240.244
R12622 gnd.n6668 gnd.n6667 240.244
R12623 gnd.n6664 gnd.n6663 240.244
R12624 gnd.n6660 gnd.n6659 240.244
R12625 gnd.n6655 gnd.n6654 240.244
R12626 gnd.n6651 gnd.n6650 240.244
R12627 gnd.n6647 gnd.n6646 240.244
R12628 gnd.n6643 gnd.n6642 240.244
R12629 gnd.n6638 gnd.n6637 240.244
R12630 gnd.n6634 gnd.n6633 240.244
R12631 gnd.n6630 gnd.n6629 240.244
R12632 gnd.n6626 gnd.n6625 240.244
R12633 gnd.n6622 gnd.n6621 240.244
R12634 gnd.n6618 gnd.n6617 240.244
R12635 gnd.n6614 gnd.n6613 240.244
R12636 gnd.n6610 gnd.n6609 240.244
R12637 gnd.n6606 gnd.n6605 240.244
R12638 gnd.n6602 gnd.n6601 240.244
R12639 gnd.n6598 gnd.n6597 240.244
R12640 gnd.n6594 gnd.n6593 240.244
R12641 gnd.n6590 gnd.n6589 240.244
R12642 gnd.n6586 gnd.n6585 240.244
R12643 gnd.n6582 gnd.n6581 240.244
R12644 gnd.n6735 gnd.n391 240.244
R12645 gnd.n6735 gnd.n386 240.244
R12646 gnd.n6743 gnd.n386 240.244
R12647 gnd.n6743 gnd.n387 240.244
R12648 gnd.n387 gnd.n358 240.244
R12649 gnd.n6804 gnd.n358 240.244
R12650 gnd.n6804 gnd.n353 240.244
R12651 gnd.n6812 gnd.n353 240.244
R12652 gnd.n6812 gnd.n354 240.244
R12653 gnd.n354 gnd.n329 240.244
R12654 gnd.n6839 gnd.n329 240.244
R12655 gnd.n6839 gnd.n324 240.244
R12656 gnd.n6848 gnd.n324 240.244
R12657 gnd.n6848 gnd.n325 240.244
R12658 gnd.n325 gnd.n304 240.244
R12659 gnd.n6873 gnd.n304 240.244
R12660 gnd.n6876 gnd.n6873 240.244
R12661 gnd.n6876 gnd.n287 240.244
R12662 gnd.n6903 gnd.n287 240.244
R12663 gnd.n6911 gnd.n6903 240.244
R12664 gnd.n6911 gnd.n6908 240.244
R12665 gnd.n6908 gnd.n73 240.244
R12666 gnd.n7324 gnd.n73 240.244
R12667 gnd.n7324 gnd.n74 240.244
R12668 gnd.n84 gnd.n74 240.244
R12669 gnd.n7318 gnd.n84 240.244
R12670 gnd.n7318 gnd.n85 240.244
R12671 gnd.n7310 gnd.n85 240.244
R12672 gnd.n7310 gnd.n102 240.244
R12673 gnd.n7306 gnd.n102 240.244
R12674 gnd.n7306 gnd.n107 240.244
R12675 gnd.n7298 gnd.n107 240.244
R12676 gnd.n7298 gnd.n121 240.244
R12677 gnd.n7294 gnd.n121 240.244
R12678 gnd.n7294 gnd.n127 240.244
R12679 gnd.n7286 gnd.n127 240.244
R12680 gnd.n7286 gnd.n142 240.244
R12681 gnd.n7282 gnd.n142 240.244
R12682 gnd.n7282 gnd.n148 240.244
R12683 gnd.n7274 gnd.n148 240.244
R12684 gnd.n7274 gnd.n162 240.244
R12685 gnd.n7270 gnd.n162 240.244
R12686 gnd.n5451 gnd.n5450 240.244
R12687 gnd.n5448 gnd.n5364 240.244
R12688 gnd.n5444 gnd.n5443 240.244
R12689 gnd.n5441 gnd.n5370 240.244
R12690 gnd.n5437 gnd.n5436 240.244
R12691 gnd.n5434 gnd.n5377 240.244
R12692 gnd.n5430 gnd.n5429 240.244
R12693 gnd.n5427 gnd.n5384 240.244
R12694 gnd.n5423 gnd.n5422 240.244
R12695 gnd.n5420 gnd.n5391 240.244
R12696 gnd.n5416 gnd.n5415 240.244
R12697 gnd.n5413 gnd.n5401 240.244
R12698 gnd.n5409 gnd.n5408 240.244
R12699 gnd.n5518 gnd.n1154 240.244
R12700 gnd.n5516 gnd.n5515 240.244
R12701 gnd.n5513 gnd.n1158 240.244
R12702 gnd.n5509 gnd.n5508 240.244
R12703 gnd.n5506 gnd.n1165 240.244
R12704 gnd.n5499 gnd.n1174 240.244
R12705 gnd.n5497 gnd.n5496 240.244
R12706 gnd.n5494 gnd.n1176 240.244
R12707 gnd.n5490 gnd.n5489 240.244
R12708 gnd.n5487 gnd.n1183 240.244
R12709 gnd.n5483 gnd.n5482 240.244
R12710 gnd.n5480 gnd.n1190 240.244
R12711 gnd.n5476 gnd.n5475 240.244
R12712 gnd.n5473 gnd.n1197 240.244
R12713 gnd.n5469 gnd.n5468 240.244
R12714 gnd.n4585 gnd.n1507 240.244
R12715 gnd.n1507 gnd.n1499 240.244
R12716 gnd.n4729 gnd.n1499 240.244
R12717 gnd.n4729 gnd.n1490 240.244
R12718 gnd.n1490 gnd.n1479 240.244
R12719 gnd.n4748 gnd.n1479 240.244
R12720 gnd.n4749 gnd.n4748 240.244
R12721 gnd.n4749 gnd.n1468 240.244
R12722 gnd.n4760 gnd.n1468 240.244
R12723 gnd.n4760 gnd.n1461 240.244
R12724 gnd.n1461 gnd.n1450 240.244
R12725 gnd.n1450 gnd.n1432 240.244
R12726 gnd.n4792 gnd.n1432 240.244
R12727 gnd.n4792 gnd.n1443 240.244
R12728 gnd.n1443 gnd.n1422 240.244
R12729 gnd.n4787 gnd.n1422 240.244
R12730 gnd.n4787 gnd.n1416 240.244
R12731 gnd.n1416 gnd.n1359 240.244
R12732 gnd.n4865 gnd.n1359 240.244
R12733 gnd.n4865 gnd.n1370 240.244
R12734 gnd.n1376 gnd.n1370 240.244
R12735 gnd.n4870 gnd.n1376 240.244
R12736 gnd.n4870 gnd.n4869 240.244
R12737 gnd.n4869 gnd.n1386 240.244
R12738 gnd.n1392 gnd.n1386 240.244
R12739 gnd.n4882 gnd.n1392 240.244
R12740 gnd.n4882 gnd.n1343 240.244
R12741 gnd.n4886 gnd.n1343 240.244
R12742 gnd.n4886 gnd.n1335 240.244
R12743 gnd.n1335 gnd.n1320 240.244
R12744 gnd.n4962 gnd.n1320 240.244
R12745 gnd.n4962 gnd.n1310 240.244
R12746 gnd.n1310 gnd.n1301 240.244
R12747 gnd.n4997 gnd.n1301 240.244
R12748 gnd.n4997 gnd.n1292 240.244
R12749 gnd.n5000 gnd.n1292 240.244
R12750 gnd.n5000 gnd.n1231 240.244
R12751 gnd.n5347 gnd.n1231 240.244
R12752 gnd.n5347 gnd.n1223 240.244
R12753 gnd.n1223 gnd.n1212 240.244
R12754 gnd.n5459 gnd.n1212 240.244
R12755 gnd.n5459 gnd.n1206 240.244
R12756 gnd.n4702 gnd.n1515 240.244
R12757 gnd.n4702 gnd.n4453 240.244
R12758 gnd.n4698 gnd.n4697 240.244
R12759 gnd.n4694 gnd.n4693 240.244
R12760 gnd.n4690 gnd.n4689 240.244
R12761 gnd.n4686 gnd.n4685 240.244
R12762 gnd.n4682 gnd.n4681 240.244
R12763 gnd.n4678 gnd.n4677 240.244
R12764 gnd.n4674 gnd.n4673 240.244
R12765 gnd.n4669 gnd.n4668 240.244
R12766 gnd.n4665 gnd.n4664 240.244
R12767 gnd.n4661 gnd.n4660 240.244
R12768 gnd.n4657 gnd.n4656 240.244
R12769 gnd.n4653 gnd.n4652 240.244
R12770 gnd.n4649 gnd.n4648 240.244
R12771 gnd.n4645 gnd.n4644 240.244
R12772 gnd.n4641 gnd.n4640 240.244
R12773 gnd.n4637 gnd.n4636 240.244
R12774 gnd.n4633 gnd.n4632 240.244
R12775 gnd.n4629 gnd.n4628 240.244
R12776 gnd.n4625 gnd.n4624 240.244
R12777 gnd.n4621 gnd.n4620 240.244
R12778 gnd.n4617 gnd.n4616 240.244
R12779 gnd.n4613 gnd.n4612 240.244
R12780 gnd.n4609 gnd.n4608 240.244
R12781 gnd.n4605 gnd.n4604 240.244
R12782 gnd.n4601 gnd.n4600 240.244
R12783 gnd.n4597 gnd.n4596 240.244
R12784 gnd.n4593 gnd.n4592 240.244
R12785 gnd.n4713 gnd.n1510 240.244
R12786 gnd.n4713 gnd.n1511 240.244
R12787 gnd.n1511 gnd.n1488 240.244
R12788 gnd.n4740 gnd.n1488 240.244
R12789 gnd.n4740 gnd.n1484 240.244
R12790 gnd.n4746 gnd.n1484 240.244
R12791 gnd.n4746 gnd.n1466 240.244
R12792 gnd.n4767 gnd.n1466 240.244
R12793 gnd.n4767 gnd.n1462 240.244
R12794 gnd.n4773 gnd.n1462 240.244
R12795 gnd.n4773 gnd.n1430 240.244
R12796 gnd.n4819 gnd.n1430 240.244
R12797 gnd.n4819 gnd.n1431 240.244
R12798 gnd.n1431 gnd.n1425 240.244
R12799 gnd.n4826 gnd.n1425 240.244
R12800 gnd.n4826 gnd.n1426 240.244
R12801 gnd.n1426 gnd.n1356 240.244
R12802 gnd.n4921 gnd.n1356 240.244
R12803 gnd.n4921 gnd.n1357 240.244
R12804 gnd.n4913 gnd.n1357 240.244
R12805 gnd.n4913 gnd.n4910 240.244
R12806 gnd.n4910 gnd.n1373 240.244
R12807 gnd.n1390 gnd.n1373 240.244
R12808 gnd.n4899 gnd.n1390 240.244
R12809 gnd.n4899 gnd.n4896 240.244
R12810 gnd.n4896 gnd.n1346 240.244
R12811 gnd.n4930 gnd.n1346 240.244
R12812 gnd.n4930 gnd.n1347 240.244
R12813 gnd.n1347 gnd.n1318 240.244
R12814 gnd.n4975 gnd.n1318 240.244
R12815 gnd.n4975 gnd.n1313 240.244
R12816 gnd.n4983 gnd.n1313 240.244
R12817 gnd.n4983 gnd.n1314 240.244
R12818 gnd.n1314 gnd.n1290 240.244
R12819 gnd.n5009 gnd.n1290 240.244
R12820 gnd.n5009 gnd.n1286 240.244
R12821 gnd.n5015 gnd.n1286 240.244
R12822 gnd.n5015 gnd.n1221 240.244
R12823 gnd.n5357 gnd.n1221 240.244
R12824 gnd.n5357 gnd.n1216 240.244
R12825 gnd.n5457 gnd.n1216 240.244
R12826 gnd.n5457 gnd.n1217 240.244
R12827 gnd.n3043 gnd.n3038 240.244
R12828 gnd.n4354 gnd.n4353 240.244
R12829 gnd.n4351 gnd.n3047 240.244
R12830 gnd.n4347 gnd.n4346 240.244
R12831 gnd.n4344 gnd.n3054 240.244
R12832 gnd.n4340 gnd.n4339 240.244
R12833 gnd.n4337 gnd.n3061 240.244
R12834 gnd.n4333 gnd.n4332 240.244
R12835 gnd.n3668 gnd.n3380 240.244
R12836 gnd.n3678 gnd.n3380 240.244
R12837 gnd.n3678 gnd.n3371 240.244
R12838 gnd.n3371 gnd.n3360 240.244
R12839 gnd.n3699 gnd.n3360 240.244
R12840 gnd.n3699 gnd.n3354 240.244
R12841 gnd.n3709 gnd.n3354 240.244
R12842 gnd.n3709 gnd.n3343 240.244
R12843 gnd.n3343 gnd.n3335 240.244
R12844 gnd.n3727 gnd.n3335 240.244
R12845 gnd.n3728 gnd.n3727 240.244
R12846 gnd.n3728 gnd.n3320 240.244
R12847 gnd.n3730 gnd.n3320 240.244
R12848 gnd.n3730 gnd.n3306 240.244
R12849 gnd.n3772 gnd.n3306 240.244
R12850 gnd.n3773 gnd.n3772 240.244
R12851 gnd.n3776 gnd.n3773 240.244
R12852 gnd.n3776 gnd.n3261 240.244
R12853 gnd.n3301 gnd.n3261 240.244
R12854 gnd.n3301 gnd.n3271 240.244
R12855 gnd.n3786 gnd.n3271 240.244
R12856 gnd.n3786 gnd.n3292 240.244
R12857 gnd.n3796 gnd.n3292 240.244
R12858 gnd.n3796 gnd.n3190 240.244
R12859 gnd.n3841 gnd.n3190 240.244
R12860 gnd.n3841 gnd.n3176 240.244
R12861 gnd.n3863 gnd.n3176 240.244
R12862 gnd.n3864 gnd.n3863 240.244
R12863 gnd.n3864 gnd.n3163 240.244
R12864 gnd.n3163 gnd.n3152 240.244
R12865 gnd.n3895 gnd.n3152 240.244
R12866 gnd.n3896 gnd.n3895 240.244
R12867 gnd.n3897 gnd.n3896 240.244
R12868 gnd.n3897 gnd.n3137 240.244
R12869 gnd.n3137 gnd.n3129 240.244
R12870 gnd.n3950 gnd.n3129 240.244
R12871 gnd.n3951 gnd.n3950 240.244
R12872 gnd.n3951 gnd.n2962 240.244
R12873 gnd.n3928 gnd.n2962 240.244
R12874 gnd.n3928 gnd.n2972 240.244
R12875 gnd.n3963 gnd.n2972 240.244
R12876 gnd.n3964 gnd.n3963 240.244
R12877 gnd.n3964 gnd.n2985 240.244
R12878 gnd.n4253 gnd.n2985 240.244
R12879 gnd.n4253 gnd.n2997 240.244
R12880 gnd.n4249 gnd.n2997 240.244
R12881 gnd.n4249 gnd.n4248 240.244
R12882 gnd.n4248 gnd.n3010 240.244
R12883 gnd.n4244 gnd.n3010 240.244
R12884 gnd.n4244 gnd.n3023 240.244
R12885 gnd.n4240 gnd.n3023 240.244
R12886 gnd.n4240 gnd.n4239 240.244
R12887 gnd.n4239 gnd.n3035 240.244
R12888 gnd.n3658 gnd.n3393 240.244
R12889 gnd.n3414 gnd.n3393 240.244
R12890 gnd.n3417 gnd.n3416 240.244
R12891 gnd.n3424 gnd.n3423 240.244
R12892 gnd.n3427 gnd.n3426 240.244
R12893 gnd.n3434 gnd.n3433 240.244
R12894 gnd.n3437 gnd.n3436 240.244
R12895 gnd.n3444 gnd.n3443 240.244
R12896 gnd.n3666 gnd.n3390 240.244
R12897 gnd.n3390 gnd.n3369 240.244
R12898 gnd.n3689 gnd.n3369 240.244
R12899 gnd.n3689 gnd.n3363 240.244
R12900 gnd.n3697 gnd.n3363 240.244
R12901 gnd.n3697 gnd.n3365 240.244
R12902 gnd.n3365 gnd.n3341 240.244
R12903 gnd.n3719 gnd.n3341 240.244
R12904 gnd.n3719 gnd.n3337 240.244
R12905 gnd.n3725 gnd.n3337 240.244
R12906 gnd.n3725 gnd.n3319 240.244
R12907 gnd.n3750 gnd.n3319 240.244
R12908 gnd.n3750 gnd.n3314 240.244
R12909 gnd.n3762 gnd.n3314 240.244
R12910 gnd.n3762 gnd.n3315 240.244
R12911 gnd.n3758 gnd.n3315 240.244
R12912 gnd.n3758 gnd.n3263 240.244
R12913 gnd.n3810 gnd.n3263 240.244
R12914 gnd.n3810 gnd.n3264 240.244
R12915 gnd.n3806 gnd.n3264 240.244
R12916 gnd.n3806 gnd.n3270 240.244
R12917 gnd.n3290 gnd.n3270 240.244
R12918 gnd.n3290 gnd.n3188 240.244
R12919 gnd.n3845 gnd.n3188 240.244
R12920 gnd.n3845 gnd.n3183 240.244
R12921 gnd.n3853 gnd.n3183 240.244
R12922 gnd.n3853 gnd.n3184 240.244
R12923 gnd.n3184 gnd.n3161 240.244
R12924 gnd.n3885 gnd.n3161 240.244
R12925 gnd.n3885 gnd.n3156 240.244
R12926 gnd.n3893 gnd.n3156 240.244
R12927 gnd.n3893 gnd.n3157 240.244
R12928 gnd.n3157 gnd.n3135 240.244
R12929 gnd.n3941 gnd.n3135 240.244
R12930 gnd.n3941 gnd.n3131 240.244
R12931 gnd.n3948 gnd.n3131 240.244
R12932 gnd.n3948 gnd.n2963 240.244
R12933 gnd.n4403 gnd.n2963 240.244
R12934 gnd.n4403 gnd.n2964 240.244
R12935 gnd.n4399 gnd.n2964 240.244
R12936 gnd.n4399 gnd.n2970 240.244
R12937 gnd.n2986 gnd.n2970 240.244
R12938 gnd.n4389 gnd.n2986 240.244
R12939 gnd.n4389 gnd.n2987 240.244
R12940 gnd.n4385 gnd.n2987 240.244
R12941 gnd.n4385 gnd.n2995 240.244
R12942 gnd.n3012 gnd.n2995 240.244
R12943 gnd.n4375 gnd.n3012 240.244
R12944 gnd.n4375 gnd.n3013 240.244
R12945 gnd.n4371 gnd.n3013 240.244
R12946 gnd.n4371 gnd.n3021 240.244
R12947 gnd.n3037 gnd.n3021 240.244
R12948 gnd.n4361 gnd.n3037 240.244
R12949 gnd.n202 gnd.n172 240.244
R12950 gnd.n205 gnd.n204 240.244
R12951 gnd.n212 gnd.n211 240.244
R12952 gnd.n215 gnd.n214 240.244
R12953 gnd.n222 gnd.n221 240.244
R12954 gnd.n225 gnd.n224 240.244
R12955 gnd.n232 gnd.n231 240.244
R12956 gnd.n234 gnd.n191 240.244
R12957 gnd.n240 gnd.n183 240.244
R12958 gnd.n6714 gnd.n394 240.244
R12959 gnd.n394 gnd.n381 240.244
R12960 gnd.n6745 gnd.n381 240.244
R12961 gnd.n6745 gnd.n376 240.244
R12962 gnd.n6752 gnd.n376 240.244
R12963 gnd.n6752 gnd.n361 240.244
R12964 gnd.n361 gnd.n348 240.244
R12965 gnd.n6814 gnd.n348 240.244
R12966 gnd.n6814 gnd.n343 240.244
R12967 gnd.n6821 gnd.n343 240.244
R12968 gnd.n6821 gnd.n332 240.244
R12969 gnd.n332 gnd.n319 240.244
R12970 gnd.n6850 gnd.n319 240.244
R12971 gnd.n6850 gnd.n314 240.244
R12972 gnd.n6864 gnd.n314 240.244
R12973 gnd.n6864 gnd.n307 240.244
R12974 gnd.n307 gnd.n303 240.244
R12975 gnd.n303 gnd.n296 240.244
R12976 gnd.n296 gnd.n290 240.244
R12977 gnd.n290 gnd.n285 240.244
R12978 gnd.n6906 gnd.n285 240.244
R12979 gnd.n6906 gnd.n66 240.244
R12980 gnd.n7326 gnd.n66 240.244
R12981 gnd.n7326 gnd.n68 240.244
R12982 gnd.n6996 gnd.n68 240.244
R12983 gnd.n6996 gnd.n88 240.244
R12984 gnd.n6992 gnd.n88 240.244
R12985 gnd.n6992 gnd.n100 240.244
R12986 gnd.n6984 gnd.n100 240.244
R12987 gnd.n6984 gnd.n110 240.244
R12988 gnd.n6980 gnd.n110 240.244
R12989 gnd.n6980 gnd.n119 240.244
R12990 gnd.n6972 gnd.n119 240.244
R12991 gnd.n6972 gnd.n130 240.244
R12992 gnd.n6968 gnd.n130 240.244
R12993 gnd.n6968 gnd.n140 240.244
R12994 gnd.n6960 gnd.n140 240.244
R12995 gnd.n6960 gnd.n151 240.244
R12996 gnd.n6956 gnd.n151 240.244
R12997 gnd.n6956 gnd.n161 240.244
R12998 gnd.n7261 gnd.n161 240.244
R12999 gnd.n7261 gnd.n170 240.244
R13000 gnd.n6493 gnd.n6492 240.244
R13001 gnd.n6501 gnd.n6500 240.244
R13002 gnd.n6503 gnd.n6502 240.244
R13003 gnd.n6513 gnd.n6512 240.244
R13004 gnd.n6521 gnd.n6520 240.244
R13005 gnd.n6523 gnd.n6522 240.244
R13006 gnd.n6533 gnd.n6532 240.244
R13007 gnd.n493 gnd.n453 240.244
R13008 gnd.n6695 gnd.n420 240.244
R13009 gnd.n6733 gnd.n395 240.244
R13010 gnd.n6733 gnd.n396 240.244
R13011 gnd.n396 gnd.n385 240.244
R13012 gnd.n404 gnd.n385 240.244
R13013 gnd.n404 gnd.n362 240.244
R13014 gnd.n6802 gnd.n362 240.244
R13015 gnd.n6802 gnd.n363 240.244
R13016 gnd.n363 gnd.n352 240.244
R13017 gnd.n6797 gnd.n352 240.244
R13018 gnd.n6797 gnd.n334 240.244
R13019 gnd.n6837 gnd.n334 240.244
R13020 gnd.n6837 gnd.n335 240.244
R13021 gnd.n335 gnd.n323 240.244
R13022 gnd.n6832 gnd.n323 240.244
R13023 gnd.n6832 gnd.n308 240.244
R13024 gnd.n6871 gnd.n308 240.244
R13025 gnd.n6871 gnd.n297 240.244
R13026 gnd.n6884 gnd.n297 240.244
R13027 gnd.n6884 gnd.n283 240.244
R13028 gnd.n6913 gnd.n283 240.244
R13029 gnd.n6913 gnd.n277 240.244
R13030 gnd.n6922 gnd.n277 240.244
R13031 gnd.n6922 gnd.n72 240.244
R13032 gnd.n6925 gnd.n72 240.244
R13033 gnd.n6925 gnd.n90 240.244
R13034 gnd.n7316 gnd.n90 240.244
R13035 gnd.n7316 gnd.n91 240.244
R13036 gnd.n7312 gnd.n91 240.244
R13037 gnd.n7312 gnd.n97 240.244
R13038 gnd.n7304 gnd.n97 240.244
R13039 gnd.n7304 gnd.n111 240.244
R13040 gnd.n7300 gnd.n111 240.244
R13041 gnd.n7300 gnd.n116 240.244
R13042 gnd.n7292 gnd.n116 240.244
R13043 gnd.n7292 gnd.n132 240.244
R13044 gnd.n7288 gnd.n132 240.244
R13045 gnd.n7288 gnd.n137 240.244
R13046 gnd.n7280 gnd.n137 240.244
R13047 gnd.n7280 gnd.n153 240.244
R13048 gnd.n7276 gnd.n153 240.244
R13049 gnd.n7276 gnd.n158 240.244
R13050 gnd.n7268 gnd.n158 240.244
R13051 gnd.n3073 gnd.n3032 240.244
R13052 gnd.n4322 gnd.n4321 240.244
R13053 gnd.n4319 gnd.n3077 240.244
R13054 gnd.n4315 gnd.n4314 240.244
R13055 gnd.n4312 gnd.n3084 240.244
R13056 gnd.n4308 gnd.n4307 240.244
R13057 gnd.n4305 gnd.n3091 240.244
R13058 gnd.n4301 gnd.n4300 240.244
R13059 gnd.n4298 gnd.n3098 240.244
R13060 gnd.n4294 gnd.n4293 240.244
R13061 gnd.n4291 gnd.n3105 240.244
R13062 gnd.n4287 gnd.n4286 240.244
R13063 gnd.n4284 gnd.n3115 240.244
R13064 gnd.n3581 gnd.n3478 240.244
R13065 gnd.n3581 gnd.n3471 240.244
R13066 gnd.n3592 gnd.n3471 240.244
R13067 gnd.n3592 gnd.n3467 240.244
R13068 gnd.n3598 gnd.n3467 240.244
R13069 gnd.n3598 gnd.n3459 240.244
R13070 gnd.n3608 gnd.n3459 240.244
R13071 gnd.n3608 gnd.n3454 240.244
R13072 gnd.n3644 gnd.n3454 240.244
R13073 gnd.n3644 gnd.n3455 240.244
R13074 gnd.n3455 gnd.n3402 240.244
R13075 gnd.n3639 gnd.n3402 240.244
R13076 gnd.n3639 gnd.n3638 240.244
R13077 gnd.n3638 gnd.n3381 240.244
R13078 gnd.n3634 gnd.n3381 240.244
R13079 gnd.n3634 gnd.n3372 240.244
R13080 gnd.n3631 gnd.n3372 240.244
R13081 gnd.n3631 gnd.n3630 240.244
R13082 gnd.n3630 gnd.n3355 240.244
R13083 gnd.n3626 gnd.n3355 240.244
R13084 gnd.n3626 gnd.n3344 240.244
R13085 gnd.n3344 gnd.n3325 240.244
R13086 gnd.n3739 gnd.n3325 240.244
R13087 gnd.n3739 gnd.n3321 240.244
R13088 gnd.n3747 gnd.n3321 240.244
R13089 gnd.n3747 gnd.n3312 240.244
R13090 gnd.n3312 gnd.n3248 240.244
R13091 gnd.n3819 gnd.n3248 240.244
R13092 gnd.n3819 gnd.n3249 240.244
R13093 gnd.n3260 gnd.n3249 240.244
R13094 gnd.n3295 gnd.n3260 240.244
R13095 gnd.n3298 gnd.n3295 240.244
R13096 gnd.n3298 gnd.n3272 240.244
R13097 gnd.n3285 gnd.n3272 240.244
R13098 gnd.n3285 gnd.n3282 240.244
R13099 gnd.n3282 gnd.n3191 240.244
R13100 gnd.n3840 gnd.n3191 240.244
R13101 gnd.n3840 gnd.n3181 240.244
R13102 gnd.n3836 gnd.n3181 240.244
R13103 gnd.n3836 gnd.n3175 240.244
R13104 gnd.n3833 gnd.n3175 240.244
R13105 gnd.n3833 gnd.n3164 240.244
R13106 gnd.n3830 gnd.n3164 240.244
R13107 gnd.n3830 gnd.n3142 240.244
R13108 gnd.n3908 gnd.n3142 240.244
R13109 gnd.n3908 gnd.n3138 240.244
R13110 gnd.n3938 gnd.n3138 240.244
R13111 gnd.n3938 gnd.n2951 240.244
R13112 gnd.n3934 gnd.n2951 240.244
R13113 gnd.n3934 gnd.n2961 240.244
R13114 gnd.n3931 gnd.n2961 240.244
R13115 gnd.n3931 gnd.n3927 240.244
R13116 gnd.n3927 gnd.n2973 240.244
R13117 gnd.n3923 gnd.n2973 240.244
R13118 gnd.n3923 gnd.n2984 240.244
R13119 gnd.n4256 gnd.n2984 240.244
R13120 gnd.n4257 gnd.n4256 240.244
R13121 gnd.n4257 gnd.n2998 240.244
R13122 gnd.n4263 gnd.n2998 240.244
R13123 gnd.n4263 gnd.n3009 240.244
R13124 gnd.n4267 gnd.n3009 240.244
R13125 gnd.n4267 gnd.n4266 240.244
R13126 gnd.n4266 gnd.n3024 240.244
R13127 gnd.n4274 gnd.n3024 240.244
R13128 gnd.n4274 gnd.n3034 240.244
R13129 gnd.n3495 gnd.n3494 240.244
R13130 gnd.n3566 gnd.n3494 240.244
R13131 gnd.n3564 gnd.n3563 240.244
R13132 gnd.n3560 gnd.n3559 240.244
R13133 gnd.n3556 gnd.n3555 240.244
R13134 gnd.n3552 gnd.n3551 240.244
R13135 gnd.n3548 gnd.n3547 240.244
R13136 gnd.n3544 gnd.n3543 240.244
R13137 gnd.n3540 gnd.n3539 240.244
R13138 gnd.n3536 gnd.n3535 240.244
R13139 gnd.n3532 gnd.n3531 240.244
R13140 gnd.n3528 gnd.n3527 240.244
R13141 gnd.n3524 gnd.n3482 240.244
R13142 gnd.n3584 gnd.n3476 240.244
R13143 gnd.n3584 gnd.n3472 240.244
R13144 gnd.n3590 gnd.n3472 240.244
R13145 gnd.n3590 gnd.n3465 240.244
R13146 gnd.n3600 gnd.n3465 240.244
R13147 gnd.n3600 gnd.n3461 240.244
R13148 gnd.n3606 gnd.n3461 240.244
R13149 gnd.n3606 gnd.n3452 240.244
R13150 gnd.n3646 gnd.n3452 240.244
R13151 gnd.n3646 gnd.n3403 240.244
R13152 gnd.n3654 gnd.n3403 240.244
R13153 gnd.n3654 gnd.n3404 240.244
R13154 gnd.n3404 gnd.n3382 240.244
R13155 gnd.n3675 gnd.n3382 240.244
R13156 gnd.n3675 gnd.n3374 240.244
R13157 gnd.n3686 gnd.n3374 240.244
R13158 gnd.n3686 gnd.n3375 240.244
R13159 gnd.n3375 gnd.n3356 240.244
R13160 gnd.n3706 gnd.n3356 240.244
R13161 gnd.n3706 gnd.n3346 240.244
R13162 gnd.n3716 gnd.n3346 240.244
R13163 gnd.n3716 gnd.n3327 240.244
R13164 gnd.n3737 gnd.n3327 240.244
R13165 gnd.n3737 gnd.n3329 240.244
R13166 gnd.n3329 gnd.n3310 240.244
R13167 gnd.n3765 gnd.n3310 240.244
R13168 gnd.n3765 gnd.n3252 240.244
R13169 gnd.n3817 gnd.n3252 240.244
R13170 gnd.n3817 gnd.n3253 240.244
R13171 gnd.n3813 gnd.n3253 240.244
R13172 gnd.n3813 gnd.n3259 240.244
R13173 gnd.n3274 gnd.n3259 240.244
R13174 gnd.n3803 gnd.n3274 240.244
R13175 gnd.n3803 gnd.n3275 240.244
R13176 gnd.n3799 gnd.n3275 240.244
R13177 gnd.n3799 gnd.n3281 240.244
R13178 gnd.n3281 gnd.n3180 240.244
R13179 gnd.n3856 gnd.n3180 240.244
R13180 gnd.n3856 gnd.n3173 240.244
R13181 gnd.n3867 gnd.n3173 240.244
R13182 gnd.n3867 gnd.n3166 240.244
R13183 gnd.n3882 gnd.n3166 240.244
R13184 gnd.n3882 gnd.n3167 240.244
R13185 gnd.n3167 gnd.n3145 240.244
R13186 gnd.n3906 gnd.n3145 240.244
R13187 gnd.n3906 gnd.n3146 240.244
R13188 gnd.n3146 gnd.n2952 240.244
R13189 gnd.n4410 gnd.n2952 240.244
R13190 gnd.n4410 gnd.n2953 240.244
R13191 gnd.n4406 gnd.n2953 240.244
R13192 gnd.n4406 gnd.n2959 240.244
R13193 gnd.n2975 gnd.n2959 240.244
R13194 gnd.n4396 gnd.n2975 240.244
R13195 gnd.n4396 gnd.n2976 240.244
R13196 gnd.n4392 gnd.n2976 240.244
R13197 gnd.n4392 gnd.n2982 240.244
R13198 gnd.n3000 gnd.n2982 240.244
R13199 gnd.n4382 gnd.n3000 240.244
R13200 gnd.n4382 gnd.n3001 240.244
R13201 gnd.n4378 gnd.n3001 240.244
R13202 gnd.n4378 gnd.n3007 240.244
R13203 gnd.n3026 gnd.n3007 240.244
R13204 gnd.n4368 gnd.n3026 240.244
R13205 gnd.n4368 gnd.n3027 240.244
R13206 gnd.n4364 gnd.n3027 240.244
R13207 gnd.n5193 gnd.n5192 240.244
R13208 gnd.n5205 gnd.n5204 240.244
R13209 gnd.n5216 gnd.n5207 240.244
R13210 gnd.n5219 gnd.n5218 240.244
R13211 gnd.n5228 gnd.n5227 240.244
R13212 gnd.n5239 gnd.n5230 240.244
R13213 gnd.n5242 gnd.n5241 240.244
R13214 gnd.n5251 gnd.n5250 240.244
R13215 gnd.n5256 gnd.n5253 240.244
R13216 gnd.n4715 gnd.n1505 240.244
R13217 gnd.n4715 gnd.n1501 240.244
R13218 gnd.n4727 gnd.n1501 240.244
R13219 gnd.n4727 gnd.n1491 240.244
R13220 gnd.n4723 gnd.n1491 240.244
R13221 gnd.n4723 gnd.n1478 240.244
R13222 gnd.n4751 gnd.n1478 240.244
R13223 gnd.n4751 gnd.n1469 240.244
R13224 gnd.n4758 gnd.n1469 240.244
R13225 gnd.n4758 gnd.n1451 240.244
R13226 gnd.n4798 gnd.n1451 240.244
R13227 gnd.n4798 gnd.n1433 240.244
R13228 gnd.n4794 gnd.n1433 240.244
R13229 gnd.n4794 gnd.n1421 240.244
R13230 gnd.n4828 gnd.n1421 240.244
R13231 gnd.n4828 gnd.n1417 240.244
R13232 gnd.n4852 gnd.n1417 240.244
R13233 gnd.n4852 gnd.n1360 240.244
R13234 gnd.n1410 gnd.n1360 240.244
R13235 gnd.n1410 gnd.n1371 240.244
R13236 gnd.n1377 gnd.n1371 240.244
R13237 gnd.n4838 gnd.n1377 240.244
R13238 gnd.n4839 gnd.n4838 240.244
R13239 gnd.n4839 gnd.n1387 240.244
R13240 gnd.n1393 gnd.n1387 240.244
R13241 gnd.n1393 gnd.n1341 240.244
R13242 gnd.n4932 gnd.n1341 240.244
R13243 gnd.n4932 gnd.n1336 240.244
R13244 gnd.n4939 gnd.n1336 240.244
R13245 gnd.n4939 gnd.n1321 240.244
R13246 gnd.n1321 gnd.n1308 240.244
R13247 gnd.n4985 gnd.n1308 240.244
R13248 gnd.n4985 gnd.n1303 240.244
R13249 gnd.n4995 gnd.n1303 240.244
R13250 gnd.n4995 gnd.n1293 240.244
R13251 gnd.n4989 gnd.n1293 240.244
R13252 gnd.n4989 gnd.n1233 240.244
R13253 gnd.n5345 gnd.n1233 240.244
R13254 gnd.n5345 gnd.n1224 240.244
R13255 gnd.n1238 gnd.n1224 240.244
R13256 gnd.n1238 gnd.n1213 240.244
R13257 gnd.n1239 gnd.n1213 240.244
R13258 gnd.n4579 gnd.n4578 240.244
R13259 gnd.n4575 gnd.n4574 240.244
R13260 gnd.n4571 gnd.n4570 240.244
R13261 gnd.n4567 gnd.n4566 240.244
R13262 gnd.n4563 gnd.n4562 240.244
R13263 gnd.n4559 gnd.n4558 240.244
R13264 gnd.n4555 gnd.n4554 240.244
R13265 gnd.n4551 gnd.n4550 240.244
R13266 gnd.n4541 gnd.n1554 240.244
R13267 gnd.n4583 gnd.n1509 240.244
R13268 gnd.n4520 gnd.n1509 240.244
R13269 gnd.n4520 gnd.n1493 240.244
R13270 gnd.n4738 gnd.n1493 240.244
R13271 gnd.n4738 gnd.n1494 240.244
R13272 gnd.n1494 gnd.n1483 240.244
R13273 gnd.n1483 gnd.n1471 240.244
R13274 gnd.n4765 gnd.n1471 240.244
R13275 gnd.n4765 gnd.n1459 240.244
R13276 gnd.n4775 gnd.n1459 240.244
R13277 gnd.n4775 gnd.n1435 240.244
R13278 gnd.n4817 gnd.n1435 240.244
R13279 gnd.n4817 gnd.n1436 240.244
R13280 gnd.n4813 gnd.n1436 240.244
R13281 gnd.n4813 gnd.n1424 240.244
R13282 gnd.n4782 gnd.n1424 240.244
R13283 gnd.n4782 gnd.n1362 240.244
R13284 gnd.n4919 gnd.n1362 240.244
R13285 gnd.n4919 gnd.n1363 240.244
R13286 gnd.n4915 gnd.n1363 240.244
R13287 gnd.n4915 gnd.n1369 240.244
R13288 gnd.n4874 gnd.n1369 240.244
R13289 gnd.n4875 gnd.n4874 240.244
R13290 gnd.n4875 gnd.n1389 240.244
R13291 gnd.n4894 gnd.n1389 240.244
R13292 gnd.n4894 gnd.n1401 240.244
R13293 gnd.n1401 gnd.n1345 240.244
R13294 gnd.n4889 gnd.n1345 240.244
R13295 gnd.n4889 gnd.n1322 240.244
R13296 gnd.n4973 gnd.n1322 240.244
R13297 gnd.n4973 gnd.n1323 240.244
R13298 gnd.n1323 gnd.n1312 240.244
R13299 gnd.n4968 gnd.n1312 240.244
R13300 gnd.n4968 gnd.n1295 240.244
R13301 gnd.n5007 gnd.n1295 240.244
R13302 gnd.n5007 gnd.n1296 240.244
R13303 gnd.n1296 gnd.n1285 240.244
R13304 gnd.n1285 gnd.n1226 240.244
R13305 gnd.n5355 gnd.n1226 240.244
R13306 gnd.n5355 gnd.n1227 240.244
R13307 gnd.n1227 gnd.n1215 240.244
R13308 gnd.n5191 gnd.n1215 240.244
R13309 gnd.n2739 gnd.n1684 240.244
R13310 gnd.n2739 gnd.n1686 240.244
R13311 gnd.n2735 gnd.n1686 240.244
R13312 gnd.n2735 gnd.n1689 240.244
R13313 gnd.n2731 gnd.n1689 240.244
R13314 gnd.n2731 gnd.n1695 240.244
R13315 gnd.n2727 gnd.n1695 240.244
R13316 gnd.n2727 gnd.n1697 240.244
R13317 gnd.n2723 gnd.n1697 240.244
R13318 gnd.n2723 gnd.n1703 240.244
R13319 gnd.n2719 gnd.n1703 240.244
R13320 gnd.n2719 gnd.n1705 240.244
R13321 gnd.n2715 gnd.n1705 240.244
R13322 gnd.n2715 gnd.n1711 240.244
R13323 gnd.n2711 gnd.n1711 240.244
R13324 gnd.n2711 gnd.n1713 240.244
R13325 gnd.n2707 gnd.n1713 240.244
R13326 gnd.n2707 gnd.n1719 240.244
R13327 gnd.n2703 gnd.n1719 240.244
R13328 gnd.n2703 gnd.n1721 240.244
R13329 gnd.n2699 gnd.n1721 240.244
R13330 gnd.n2699 gnd.n1727 240.244
R13331 gnd.n2695 gnd.n1727 240.244
R13332 gnd.n2695 gnd.n1729 240.244
R13333 gnd.n2691 gnd.n1729 240.244
R13334 gnd.n2691 gnd.n1735 240.244
R13335 gnd.n2687 gnd.n1735 240.244
R13336 gnd.n2687 gnd.n1737 240.244
R13337 gnd.n2683 gnd.n1737 240.244
R13338 gnd.n2683 gnd.n1743 240.244
R13339 gnd.n2679 gnd.n1743 240.244
R13340 gnd.n2679 gnd.n1745 240.244
R13341 gnd.n2675 gnd.n1745 240.244
R13342 gnd.n2675 gnd.n1751 240.244
R13343 gnd.n2671 gnd.n1751 240.244
R13344 gnd.n2671 gnd.n1753 240.244
R13345 gnd.n2667 gnd.n1753 240.244
R13346 gnd.n2667 gnd.n1759 240.244
R13347 gnd.n2663 gnd.n1759 240.244
R13348 gnd.n2663 gnd.n1761 240.244
R13349 gnd.n2659 gnd.n1761 240.244
R13350 gnd.n2659 gnd.n1767 240.244
R13351 gnd.n2655 gnd.n1767 240.244
R13352 gnd.n2655 gnd.n1769 240.244
R13353 gnd.n2651 gnd.n1769 240.244
R13354 gnd.n2651 gnd.n1775 240.244
R13355 gnd.n2647 gnd.n1775 240.244
R13356 gnd.n2647 gnd.n1777 240.244
R13357 gnd.n2643 gnd.n1777 240.244
R13358 gnd.n2643 gnd.n1783 240.244
R13359 gnd.n2639 gnd.n1783 240.244
R13360 gnd.n2639 gnd.n1785 240.244
R13361 gnd.n2635 gnd.n1785 240.244
R13362 gnd.n2635 gnd.n1791 240.244
R13363 gnd.n2631 gnd.n1791 240.244
R13364 gnd.n2631 gnd.n1793 240.244
R13365 gnd.n2627 gnd.n1793 240.244
R13366 gnd.n2627 gnd.n1799 240.244
R13367 gnd.n2623 gnd.n1799 240.244
R13368 gnd.n2623 gnd.n1801 240.244
R13369 gnd.n2619 gnd.n1801 240.244
R13370 gnd.n2619 gnd.n1807 240.244
R13371 gnd.n2615 gnd.n1807 240.244
R13372 gnd.n2615 gnd.n1809 240.244
R13373 gnd.n2611 gnd.n1809 240.244
R13374 gnd.n2611 gnd.n1815 240.244
R13375 gnd.n2607 gnd.n1815 240.244
R13376 gnd.n2607 gnd.n1817 240.244
R13377 gnd.n2603 gnd.n1817 240.244
R13378 gnd.n2603 gnd.n1823 240.244
R13379 gnd.n2599 gnd.n1823 240.244
R13380 gnd.n2599 gnd.n1825 240.244
R13381 gnd.n2595 gnd.n1825 240.244
R13382 gnd.n2595 gnd.n1831 240.244
R13383 gnd.n2591 gnd.n1831 240.244
R13384 gnd.n2591 gnd.n1833 240.244
R13385 gnd.n2587 gnd.n1833 240.244
R13386 gnd.n2587 gnd.n1839 240.244
R13387 gnd.n2583 gnd.n1839 240.244
R13388 gnd.n2583 gnd.n1841 240.244
R13389 gnd.n2579 gnd.n1841 240.244
R13390 gnd.n2579 gnd.n1847 240.244
R13391 gnd.n2575 gnd.n1847 240.244
R13392 gnd.n2575 gnd.n1849 240.244
R13393 gnd.n2571 gnd.n1849 240.244
R13394 gnd.n2571 gnd.n1855 240.244
R13395 gnd.n2567 gnd.n1855 240.244
R13396 gnd.n2567 gnd.n1857 240.244
R13397 gnd.n2563 gnd.n1857 240.244
R13398 gnd.n2563 gnd.n1863 240.244
R13399 gnd.n2559 gnd.n1863 240.244
R13400 gnd.n2559 gnd.n1865 240.244
R13401 gnd.n2555 gnd.n1865 240.244
R13402 gnd.n2555 gnd.n1871 240.244
R13403 gnd.n2551 gnd.n1871 240.244
R13404 gnd.n2551 gnd.n1873 240.244
R13405 gnd.n2547 gnd.n1873 240.244
R13406 gnd.n2547 gnd.n1879 240.244
R13407 gnd.n2543 gnd.n1879 240.244
R13408 gnd.n2543 gnd.n1881 240.244
R13409 gnd.n2539 gnd.n1881 240.244
R13410 gnd.n2539 gnd.n1887 240.244
R13411 gnd.n2535 gnd.n1887 240.244
R13412 gnd.n2535 gnd.n1889 240.244
R13413 gnd.n2531 gnd.n1889 240.244
R13414 gnd.n2531 gnd.n1895 240.244
R13415 gnd.n2527 gnd.n1895 240.244
R13416 gnd.n2527 gnd.n1897 240.244
R13417 gnd.n2523 gnd.n1897 240.244
R13418 gnd.n2523 gnd.n1903 240.244
R13419 gnd.n2519 gnd.n1903 240.244
R13420 gnd.n2519 gnd.n1905 240.244
R13421 gnd.n2515 gnd.n1905 240.244
R13422 gnd.n2515 gnd.n1911 240.244
R13423 gnd.n2511 gnd.n1911 240.244
R13424 gnd.n2511 gnd.n1913 240.244
R13425 gnd.n2507 gnd.n1913 240.244
R13426 gnd.n2507 gnd.n1919 240.244
R13427 gnd.n2503 gnd.n1919 240.244
R13428 gnd.n2503 gnd.n1921 240.244
R13429 gnd.n2499 gnd.n1921 240.244
R13430 gnd.n2499 gnd.n1927 240.244
R13431 gnd.n2495 gnd.n1927 240.244
R13432 gnd.n2495 gnd.n1929 240.244
R13433 gnd.n2491 gnd.n1929 240.244
R13434 gnd.n2491 gnd.n1935 240.244
R13435 gnd.n2487 gnd.n1935 240.244
R13436 gnd.n2487 gnd.n1937 240.244
R13437 gnd.n2483 gnd.n1937 240.244
R13438 gnd.n2483 gnd.n1943 240.244
R13439 gnd.n2479 gnd.n1943 240.244
R13440 gnd.n2479 gnd.n1945 240.244
R13441 gnd.n2475 gnd.n1945 240.244
R13442 gnd.n2475 gnd.n1951 240.244
R13443 gnd.n2471 gnd.n1951 240.244
R13444 gnd.n2471 gnd.n1953 240.244
R13445 gnd.n2467 gnd.n1953 240.244
R13446 gnd.n2467 gnd.n1959 240.244
R13447 gnd.n2463 gnd.n1959 240.244
R13448 gnd.n2463 gnd.n1961 240.244
R13449 gnd.n2459 gnd.n1961 240.244
R13450 gnd.n2459 gnd.n1967 240.244
R13451 gnd.n2455 gnd.n1967 240.244
R13452 gnd.n2455 gnd.n1969 240.244
R13453 gnd.n2451 gnd.n1969 240.244
R13454 gnd.n2451 gnd.n1975 240.244
R13455 gnd.n2447 gnd.n1975 240.244
R13456 gnd.n2447 gnd.n1977 240.244
R13457 gnd.n2443 gnd.n1977 240.244
R13458 gnd.n2443 gnd.n1983 240.244
R13459 gnd.n2439 gnd.n1983 240.244
R13460 gnd.n2439 gnd.n1985 240.244
R13461 gnd.n2435 gnd.n1985 240.244
R13462 gnd.n2435 gnd.n1991 240.244
R13463 gnd.n2431 gnd.n1991 240.244
R13464 gnd.n2431 gnd.n1993 240.244
R13465 gnd.n2427 gnd.n1993 240.244
R13466 gnd.n2427 gnd.n1999 240.244
R13467 gnd.n2423 gnd.n1999 240.244
R13468 gnd.n2423 gnd.n2001 240.244
R13469 gnd.n2419 gnd.n2001 240.244
R13470 gnd.n2419 gnd.n2007 240.244
R13471 gnd.n2415 gnd.n2007 240.244
R13472 gnd.n2415 gnd.n2009 240.244
R13473 gnd.n2411 gnd.n2009 240.244
R13474 gnd.n2411 gnd.n2015 240.244
R13475 gnd.n2407 gnd.n2015 240.244
R13476 gnd.n2407 gnd.n2017 240.244
R13477 gnd.n2403 gnd.n2017 240.244
R13478 gnd.n2403 gnd.n2023 240.244
R13479 gnd.n2399 gnd.n2023 240.244
R13480 gnd.n2399 gnd.n2025 240.244
R13481 gnd.n2395 gnd.n2025 240.244
R13482 gnd.n2395 gnd.n2031 240.244
R13483 gnd.n2391 gnd.n2031 240.244
R13484 gnd.n2391 gnd.n2033 240.244
R13485 gnd.n2387 gnd.n2033 240.244
R13486 gnd.n2387 gnd.n2039 240.244
R13487 gnd.n2383 gnd.n2039 240.244
R13488 gnd.n2383 gnd.n2041 240.244
R13489 gnd.n2379 gnd.n2041 240.244
R13490 gnd.n2375 gnd.n2046 240.244
R13491 gnd.n2375 gnd.n2048 240.244
R13492 gnd.n2369 gnd.n2048 240.244
R13493 gnd.n2369 gnd.n2054 240.244
R13494 gnd.n2365 gnd.n2054 240.244
R13495 gnd.n2365 gnd.n2056 240.244
R13496 gnd.n2361 gnd.n2056 240.244
R13497 gnd.n2361 gnd.n2061 240.244
R13498 gnd.n2357 gnd.n2061 240.244
R13499 gnd.n2357 gnd.n2063 240.244
R13500 gnd.n2353 gnd.n2063 240.244
R13501 gnd.n2353 gnd.n2069 240.244
R13502 gnd.n2349 gnd.n2069 240.244
R13503 gnd.n2349 gnd.n2071 240.244
R13504 gnd.n2345 gnd.n2071 240.244
R13505 gnd.n2345 gnd.n2077 240.244
R13506 gnd.n2341 gnd.n2077 240.244
R13507 gnd.n2341 gnd.n2079 240.244
R13508 gnd.n2337 gnd.n2079 240.244
R13509 gnd.n2337 gnd.n2085 240.244
R13510 gnd.n2333 gnd.n2085 240.244
R13511 gnd.n2333 gnd.n2087 240.244
R13512 gnd.n2329 gnd.n2087 240.244
R13513 gnd.n2329 gnd.n2093 240.244
R13514 gnd.n2325 gnd.n2093 240.244
R13515 gnd.n2325 gnd.n2095 240.244
R13516 gnd.n2321 gnd.n2095 240.244
R13517 gnd.n2321 gnd.n2101 240.244
R13518 gnd.n2317 gnd.n2101 240.244
R13519 gnd.n2317 gnd.n2103 240.244
R13520 gnd.n2313 gnd.n2103 240.244
R13521 gnd.n2313 gnd.n2109 240.244
R13522 gnd.n2309 gnd.n2109 240.244
R13523 gnd.n2309 gnd.n2111 240.244
R13524 gnd.n2305 gnd.n2111 240.244
R13525 gnd.n2305 gnd.n2117 240.244
R13526 gnd.n2301 gnd.n2117 240.244
R13527 gnd.n2301 gnd.n2119 240.244
R13528 gnd.n2297 gnd.n2119 240.244
R13529 gnd.n2297 gnd.n2125 240.244
R13530 gnd.n2293 gnd.n2125 240.244
R13531 gnd.n2293 gnd.n2127 240.244
R13532 gnd.n2289 gnd.n2127 240.244
R13533 gnd.n2289 gnd.n2133 240.244
R13534 gnd.n2285 gnd.n2133 240.244
R13535 gnd.n2285 gnd.n2135 240.244
R13536 gnd.n2281 gnd.n2135 240.244
R13537 gnd.n2281 gnd.n2141 240.244
R13538 gnd.n2277 gnd.n2141 240.244
R13539 gnd.n2277 gnd.n2143 240.244
R13540 gnd.n2273 gnd.n2143 240.244
R13541 gnd.n2273 gnd.n2149 240.244
R13542 gnd.n2269 gnd.n2149 240.244
R13543 gnd.n2269 gnd.n2151 240.244
R13544 gnd.n2265 gnd.n2151 240.244
R13545 gnd.n2265 gnd.n2157 240.244
R13546 gnd.n2261 gnd.n2157 240.244
R13547 gnd.n2261 gnd.n2159 240.244
R13548 gnd.n2257 gnd.n2159 240.244
R13549 gnd.n2257 gnd.n2165 240.244
R13550 gnd.n2253 gnd.n2165 240.244
R13551 gnd.n2253 gnd.n2167 240.244
R13552 gnd.n2249 gnd.n2167 240.244
R13553 gnd.n2249 gnd.n2173 240.244
R13554 gnd.n2245 gnd.n2173 240.244
R13555 gnd.n2245 gnd.n2175 240.244
R13556 gnd.n2241 gnd.n2175 240.244
R13557 gnd.n2241 gnd.n2181 240.244
R13558 gnd.n2237 gnd.n2181 240.244
R13559 gnd.n2237 gnd.n2183 240.244
R13560 gnd.n2233 gnd.n2183 240.244
R13561 gnd.n2233 gnd.n2189 240.244
R13562 gnd.n2229 gnd.n2189 240.244
R13563 gnd.n2229 gnd.n2191 240.244
R13564 gnd.n2225 gnd.n2191 240.244
R13565 gnd.n2225 gnd.n2197 240.244
R13566 gnd.n2221 gnd.n2197 240.244
R13567 gnd.n2221 gnd.n2199 240.244
R13568 gnd.n2217 gnd.n2199 240.244
R13569 gnd.n2217 gnd.n2205 240.244
R13570 gnd.n2213 gnd.n2205 240.244
R13571 gnd.n2213 gnd.n2207 240.244
R13572 gnd.n2207 gnd.n243 240.244
R13573 gnd.n7039 gnd.n243 240.244
R13574 gnd.n4451 gnd.n1556 240.244
R13575 gnd.n4447 gnd.n1556 240.244
R13576 gnd.n4447 gnd.n4446 240.244
R13577 gnd.n4446 gnd.n4445 240.244
R13578 gnd.n4445 gnd.n4422 240.244
R13579 gnd.n4441 gnd.n4422 240.244
R13580 gnd.n4441 gnd.n4440 240.244
R13581 gnd.n4440 gnd.n4439 240.244
R13582 gnd.n4439 gnd.n4428 240.244
R13583 gnd.n4435 gnd.n4428 240.244
R13584 gnd.n4435 gnd.n1448 240.244
R13585 gnd.n4801 gnd.n1448 240.244
R13586 gnd.n4802 gnd.n4801 240.244
R13587 gnd.n4802 gnd.n1444 240.244
R13588 gnd.n4810 gnd.n1444 240.244
R13589 gnd.n4810 gnd.n1413 240.244
R13590 gnd.n4855 gnd.n1413 240.244
R13591 gnd.n4856 gnd.n4855 240.244
R13592 gnd.n4856 gnd.n1411 240.244
R13593 gnd.n4862 gnd.n1411 240.244
R13594 gnd.n4862 gnd.n1379 240.244
R13595 gnd.n4907 gnd.n1379 240.244
R13596 gnd.n4907 gnd.n1380 240.244
R13597 gnd.n4902 gnd.n1380 240.244
R13598 gnd.n4902 gnd.n1383 240.244
R13599 gnd.n1399 gnd.n1383 240.244
R13600 gnd.n1399 gnd.n1394 240.244
R13601 gnd.n1394 gnd.n1333 240.244
R13602 gnd.n4942 gnd.n1333 240.244
R13603 gnd.n4942 gnd.n1328 240.244
R13604 gnd.n4959 gnd.n1328 240.244
R13605 gnd.n4959 gnd.n1329 240.244
R13606 gnd.n4955 gnd.n1329 240.244
R13607 gnd.n4955 gnd.n4954 240.244
R13608 gnd.n4954 gnd.n4953 240.244
R13609 gnd.n4953 gnd.n1283 240.244
R13610 gnd.n5018 gnd.n1283 240.244
R13611 gnd.n5018 gnd.n1279 240.244
R13612 gnd.n5024 gnd.n1279 240.244
R13613 gnd.n5025 gnd.n5024 240.244
R13614 gnd.n5028 gnd.n5025 240.244
R13615 gnd.n5028 gnd.n1274 240.244
R13616 gnd.n5188 gnd.n1274 240.244
R13617 gnd.n5188 gnd.n1275 240.244
R13618 gnd.n5184 gnd.n1275 240.244
R13619 gnd.n5184 gnd.n5181 240.244
R13620 gnd.n5181 gnd.n5180 240.244
R13621 gnd.n5180 gnd.n5036 240.244
R13622 gnd.n5176 gnd.n5036 240.244
R13623 gnd.n5176 gnd.n5042 240.244
R13624 gnd.n5100 gnd.n5042 240.244
R13625 gnd.n5100 gnd.n5097 240.244
R13626 gnd.n5106 gnd.n5097 240.244
R13627 gnd.n5106 gnd.n5080 240.244
R13628 gnd.n5121 gnd.n5080 240.244
R13629 gnd.n5121 gnd.n5076 240.244
R13630 gnd.n5127 gnd.n5076 240.244
R13631 gnd.n5127 gnd.n5067 240.244
R13632 gnd.n5142 gnd.n5067 240.244
R13633 gnd.n5142 gnd.n5062 240.244
R13634 gnd.n5150 gnd.n5062 240.244
R13635 gnd.n5150 gnd.n5063 240.244
R13636 gnd.n5063 gnd.n1069 240.244
R13637 gnd.n5629 gnd.n1069 240.244
R13638 gnd.n5629 gnd.n1064 240.244
R13639 gnd.n5647 gnd.n1064 240.244
R13640 gnd.n5647 gnd.n1065 240.244
R13641 gnd.n5643 gnd.n1065 240.244
R13642 gnd.n5643 gnd.n5642 240.244
R13643 gnd.n5642 gnd.n5641 240.244
R13644 gnd.n5641 gnd.n987 240.244
R13645 gnd.n5695 gnd.n987 240.244
R13646 gnd.n5695 gnd.n982 240.244
R13647 gnd.n5703 gnd.n982 240.244
R13648 gnd.n5703 gnd.n983 240.244
R13649 gnd.n983 gnd.n925 240.244
R13650 gnd.n5766 gnd.n925 240.244
R13651 gnd.n5766 gnd.n921 240.244
R13652 gnd.n5772 gnd.n921 240.244
R13653 gnd.n5773 gnd.n5772 240.244
R13654 gnd.n5774 gnd.n5773 240.244
R13655 gnd.n5774 gnd.n917 240.244
R13656 gnd.n5780 gnd.n917 240.244
R13657 gnd.n5780 gnd.n870 240.244
R13658 gnd.n5867 gnd.n870 240.244
R13659 gnd.n5867 gnd.n865 240.244
R13660 gnd.n5881 gnd.n865 240.244
R13661 gnd.n5881 gnd.n866 240.244
R13662 gnd.n5877 gnd.n866 240.244
R13663 gnd.n5877 gnd.n5876 240.244
R13664 gnd.n5876 gnd.n831 240.244
R13665 gnd.n5924 gnd.n831 240.244
R13666 gnd.n5924 gnd.n826 240.244
R13667 gnd.n5935 gnd.n826 240.244
R13668 gnd.n5935 gnd.n827 240.244
R13669 gnd.n5931 gnd.n827 240.244
R13670 gnd.n5931 gnd.n784 240.244
R13671 gnd.n6079 gnd.n784 240.244
R13672 gnd.n6079 gnd.n779 240.244
R13673 gnd.n6087 gnd.n779 240.244
R13674 gnd.n6087 gnd.n780 240.244
R13675 gnd.n780 gnd.n755 240.244
R13676 gnd.n6115 gnd.n755 240.244
R13677 gnd.n6115 gnd.n751 240.244
R13678 gnd.n6121 gnd.n751 240.244
R13679 gnd.n6121 gnd.n732 240.244
R13680 gnd.n6142 gnd.n732 240.244
R13681 gnd.n6142 gnd.n728 240.244
R13682 gnd.n6148 gnd.n728 240.244
R13683 gnd.n6148 gnd.n706 240.244
R13684 gnd.n6181 gnd.n706 240.244
R13685 gnd.n6181 gnd.n702 240.244
R13686 gnd.n6187 gnd.n702 240.244
R13687 gnd.n6187 gnd.n653 240.244
R13688 gnd.n6353 gnd.n653 240.244
R13689 gnd.n6353 gnd.n648 240.244
R13690 gnd.n6361 gnd.n648 240.244
R13691 gnd.n6361 gnd.n649 240.244
R13692 gnd.n649 gnd.n628 240.244
R13693 gnd.n6383 gnd.n628 240.244
R13694 gnd.n6383 gnd.n623 240.244
R13695 gnd.n6391 gnd.n623 240.244
R13696 gnd.n6391 gnd.n624 240.244
R13697 gnd.n624 gnd.n603 240.244
R13698 gnd.n6413 gnd.n603 240.244
R13699 gnd.n6413 gnd.n598 240.244
R13700 gnd.n6421 gnd.n598 240.244
R13701 gnd.n6421 gnd.n599 240.244
R13702 gnd.n599 gnd.n578 240.244
R13703 gnd.n6443 gnd.n578 240.244
R13704 gnd.n6443 gnd.n573 240.244
R13705 gnd.n6461 gnd.n573 240.244
R13706 gnd.n6461 gnd.n574 240.244
R13707 gnd.n6457 gnd.n574 240.244
R13708 gnd.n6457 gnd.n6456 240.244
R13709 gnd.n6456 gnd.n6454 240.244
R13710 gnd.n6454 gnd.n417 240.244
R13711 gnd.n6717 gnd.n417 240.244
R13712 gnd.n6717 gnd.n412 240.244
R13713 gnd.n6725 gnd.n412 240.244
R13714 gnd.n6725 gnd.n413 240.244
R13715 gnd.n413 gnd.n373 240.244
R13716 gnd.n6755 gnd.n373 240.244
R13717 gnd.n6755 gnd.n368 240.244
R13718 gnd.n6788 gnd.n368 240.244
R13719 gnd.n6788 gnd.n369 240.244
R13720 gnd.n6784 gnd.n369 240.244
R13721 gnd.n6784 gnd.n6783 240.244
R13722 gnd.n6783 gnd.n6782 240.244
R13723 gnd.n6782 gnd.n6763 240.244
R13724 gnd.n6778 gnd.n6763 240.244
R13725 gnd.n6778 gnd.n6777 240.244
R13726 gnd.n6777 gnd.n6776 240.244
R13727 gnd.n6776 gnd.n6769 240.244
R13728 gnd.n6769 gnd.n294 240.244
R13729 gnd.n6887 gnd.n294 240.244
R13730 gnd.n6887 gnd.n291 240.244
R13731 gnd.n6900 gnd.n291 240.244
R13732 gnd.n6900 gnd.n292 240.244
R13733 gnd.n6895 gnd.n292 240.244
R13734 gnd.n6895 gnd.n6894 240.244
R13735 gnd.n6894 gnd.n263 240.244
R13736 gnd.n6999 gnd.n263 240.244
R13737 gnd.n7000 gnd.n6999 240.244
R13738 gnd.n7000 gnd.n261 240.244
R13739 gnd.n7006 gnd.n261 240.244
R13740 gnd.n7007 gnd.n7006 240.244
R13741 gnd.n7008 gnd.n7007 240.244
R13742 gnd.n7008 gnd.n257 240.244
R13743 gnd.n7014 gnd.n257 240.244
R13744 gnd.n7015 gnd.n7014 240.244
R13745 gnd.n7016 gnd.n7015 240.244
R13746 gnd.n7016 gnd.n253 240.244
R13747 gnd.n7022 gnd.n253 240.244
R13748 gnd.n7023 gnd.n7022 240.244
R13749 gnd.n7024 gnd.n7023 240.244
R13750 gnd.n7024 gnd.n249 240.244
R13751 gnd.n7031 gnd.n249 240.244
R13752 gnd.n7032 gnd.n7031 240.244
R13753 gnd.n7033 gnd.n7032 240.244
R13754 gnd.n7033 gnd.n244 240.244
R13755 gnd.n2746 gnd.n1681 240.244
R13756 gnd.n2746 gnd.n1679 240.244
R13757 gnd.n2750 gnd.n1679 240.244
R13758 gnd.n2750 gnd.n1675 240.244
R13759 gnd.n2756 gnd.n1675 240.244
R13760 gnd.n2756 gnd.n1673 240.244
R13761 gnd.n2760 gnd.n1673 240.244
R13762 gnd.n2760 gnd.n1669 240.244
R13763 gnd.n2766 gnd.n1669 240.244
R13764 gnd.n2766 gnd.n1667 240.244
R13765 gnd.n2770 gnd.n1667 240.244
R13766 gnd.n2770 gnd.n1663 240.244
R13767 gnd.n2776 gnd.n1663 240.244
R13768 gnd.n2776 gnd.n1661 240.244
R13769 gnd.n2780 gnd.n1661 240.244
R13770 gnd.n2780 gnd.n1657 240.244
R13771 gnd.n2786 gnd.n1657 240.244
R13772 gnd.n2786 gnd.n1655 240.244
R13773 gnd.n2790 gnd.n1655 240.244
R13774 gnd.n2790 gnd.n1651 240.244
R13775 gnd.n2796 gnd.n1651 240.244
R13776 gnd.n2796 gnd.n1649 240.244
R13777 gnd.n2800 gnd.n1649 240.244
R13778 gnd.n2800 gnd.n1645 240.244
R13779 gnd.n2806 gnd.n1645 240.244
R13780 gnd.n2806 gnd.n1643 240.244
R13781 gnd.n2810 gnd.n1643 240.244
R13782 gnd.n2810 gnd.n1639 240.244
R13783 gnd.n2816 gnd.n1639 240.244
R13784 gnd.n2816 gnd.n1637 240.244
R13785 gnd.n2820 gnd.n1637 240.244
R13786 gnd.n2820 gnd.n1633 240.244
R13787 gnd.n2826 gnd.n1633 240.244
R13788 gnd.n2826 gnd.n1631 240.244
R13789 gnd.n2830 gnd.n1631 240.244
R13790 gnd.n2830 gnd.n1627 240.244
R13791 gnd.n2836 gnd.n1627 240.244
R13792 gnd.n2836 gnd.n1625 240.244
R13793 gnd.n2840 gnd.n1625 240.244
R13794 gnd.n2840 gnd.n1621 240.244
R13795 gnd.n2846 gnd.n1621 240.244
R13796 gnd.n2846 gnd.n1619 240.244
R13797 gnd.n2850 gnd.n1619 240.244
R13798 gnd.n2850 gnd.n1615 240.244
R13799 gnd.n2856 gnd.n1615 240.244
R13800 gnd.n2856 gnd.n1613 240.244
R13801 gnd.n2860 gnd.n1613 240.244
R13802 gnd.n2860 gnd.n1609 240.244
R13803 gnd.n2866 gnd.n1609 240.244
R13804 gnd.n2866 gnd.n1607 240.244
R13805 gnd.n2870 gnd.n1607 240.244
R13806 gnd.n2870 gnd.n1603 240.244
R13807 gnd.n2876 gnd.n1603 240.244
R13808 gnd.n2876 gnd.n1601 240.244
R13809 gnd.n2880 gnd.n1601 240.244
R13810 gnd.n2880 gnd.n1597 240.244
R13811 gnd.n2886 gnd.n1597 240.244
R13812 gnd.n2886 gnd.n1595 240.244
R13813 gnd.n2890 gnd.n1595 240.244
R13814 gnd.n2890 gnd.n1591 240.244
R13815 gnd.n2896 gnd.n1591 240.244
R13816 gnd.n2896 gnd.n1589 240.244
R13817 gnd.n2900 gnd.n1589 240.244
R13818 gnd.n2900 gnd.n1585 240.244
R13819 gnd.n2906 gnd.n1585 240.244
R13820 gnd.n2906 gnd.n1583 240.244
R13821 gnd.n2910 gnd.n1583 240.244
R13822 gnd.n2910 gnd.n1579 240.244
R13823 gnd.n2916 gnd.n1579 240.244
R13824 gnd.n2916 gnd.n1577 240.244
R13825 gnd.n2920 gnd.n1577 240.244
R13826 gnd.n2920 gnd.n1573 240.244
R13827 gnd.n2926 gnd.n1573 240.244
R13828 gnd.n2926 gnd.n1571 240.244
R13829 gnd.n2930 gnd.n1571 240.244
R13830 gnd.n2930 gnd.n1567 240.244
R13831 gnd.n2936 gnd.n1567 240.244
R13832 gnd.n2936 gnd.n1565 240.244
R13833 gnd.n2940 gnd.n1565 240.244
R13834 gnd.n2940 gnd.n1561 240.244
R13835 gnd.n2947 gnd.n1561 240.244
R13836 gnd.n2947 gnd.n1559 240.244
R13837 gnd.n4414 gnd.n1559 240.244
R13838 gnd.n4414 gnd.n1555 240.244
R13839 gnd.n5171 gnd.n1262 240.244
R13840 gnd.n5171 gnd.n5045 240.244
R13841 gnd.n5050 gnd.n5045 240.244
R13842 gnd.n5051 gnd.n5050 240.244
R13843 gnd.n5052 gnd.n5051 240.244
R13844 gnd.n5118 gnd.n5052 240.244
R13845 gnd.n5118 gnd.n5055 240.244
R13846 gnd.n5056 gnd.n5055 240.244
R13847 gnd.n5057 gnd.n5056 240.244
R13848 gnd.n5059 gnd.n5057 240.244
R13849 gnd.n5153 gnd.n5059 240.244
R13850 gnd.n5153 gnd.n1077 240.244
R13851 gnd.n5620 gnd.n1077 240.244
R13852 gnd.n5620 gnd.n1073 240.244
R13853 gnd.n5626 gnd.n1073 240.244
R13854 gnd.n5626 gnd.n1004 240.244
R13855 gnd.n5660 gnd.n1004 240.244
R13856 gnd.n5660 gnd.n1000 240.244
R13857 gnd.n5666 gnd.n1000 240.244
R13858 gnd.n5666 gnd.n967 240.244
R13859 gnd.n5715 gnd.n967 240.244
R13860 gnd.n5715 gnd.n961 240.244
R13861 gnd.n5722 gnd.n961 240.244
R13862 gnd.n5722 gnd.n962 240.244
R13863 gnd.n962 gnd.n932 240.244
R13864 gnd.n5757 gnd.n932 240.244
R13865 gnd.n5757 gnd.n928 240.244
R13866 gnd.n5763 gnd.n928 240.244
R13867 gnd.n5763 gnd.n899 240.244
R13868 gnd.n5799 gnd.n899 240.244
R13869 gnd.n5799 gnd.n895 240.244
R13870 gnd.n5805 gnd.n895 240.244
R13871 gnd.n5805 gnd.n884 240.244
R13872 gnd.n5843 gnd.n884 240.244
R13873 gnd.n5843 gnd.n880 240.244
R13874 gnd.n5849 gnd.n880 240.244
R13875 gnd.n5849 gnd.n854 240.244
R13876 gnd.n5892 gnd.n854 240.244
R13877 gnd.n5892 gnd.n849 240.244
R13878 gnd.n5899 gnd.n849 240.244
R13879 gnd.n5899 gnd.n839 240.244
R13880 gnd.n839 gnd.n818 240.244
R13881 gnd.n5945 gnd.n818 240.244
R13882 gnd.n5945 gnd.n814 240.244
R13883 gnd.n5951 gnd.n814 240.244
R13884 gnd.n5951 gnd.n793 240.244
R13885 gnd.n6070 gnd.n793 240.244
R13886 gnd.n6070 gnd.n789 240.244
R13887 gnd.n6076 gnd.n789 240.244
R13888 gnd.n6076 gnd.n770 240.244
R13889 gnd.n6098 gnd.n770 240.244
R13890 gnd.n6098 gnd.n764 240.244
R13891 gnd.n6105 gnd.n764 240.244
R13892 gnd.n6105 gnd.n765 240.244
R13893 gnd.n765 gnd.n740 240.244
R13894 gnd.n6133 gnd.n740 240.244
R13895 gnd.n6133 gnd.n736 240.244
R13896 gnd.n6139 gnd.n736 240.244
R13897 gnd.n6139 gnd.n716 240.244
R13898 gnd.n6165 gnd.n716 240.244
R13899 gnd.n6165 gnd.n710 240.244
R13900 gnd.n6178 gnd.n710 240.244
R13901 gnd.n6178 gnd.n711 240.244
R13902 gnd.n6170 gnd.n711 240.244
R13903 gnd.n6171 gnd.n6170 240.244
R13904 gnd.n6171 gnd.n644 240.244
R13905 gnd.n6364 gnd.n644 240.244
R13906 gnd.n6364 gnd.n638 240.244
R13907 gnd.n6371 gnd.n638 240.244
R13908 gnd.n6371 gnd.n639 240.244
R13909 gnd.n639 gnd.n619 240.244
R13910 gnd.n6394 gnd.n619 240.244
R13911 gnd.n6394 gnd.n613 240.244
R13912 gnd.n6401 gnd.n613 240.244
R13913 gnd.n6401 gnd.n614 240.244
R13914 gnd.n614 gnd.n594 240.244
R13915 gnd.n6424 gnd.n594 240.244
R13916 gnd.n6424 gnd.n587 240.244
R13917 gnd.n6431 gnd.n587 240.244
R13918 gnd.n6431 gnd.n589 240.244
R13919 gnd.n589 gnd.n570 240.244
R13920 gnd.n6464 gnd.n570 240.244
R13921 gnd.n1261 gnd.n1260 240.244
R13922 gnd.n1266 gnd.n1260 240.244
R13923 gnd.n1268 gnd.n1267 240.244
R13924 gnd.n1270 gnd.n1269 240.244
R13925 gnd.n5197 gnd.n5196 240.244
R13926 gnd.n5200 gnd.n5199 240.244
R13927 gnd.n5211 gnd.n5210 240.244
R13928 gnd.n5213 gnd.n5212 240.244
R13929 gnd.n5223 gnd.n5222 240.244
R13930 gnd.n5234 gnd.n5233 240.244
R13931 gnd.n5236 gnd.n5235 240.244
R13932 gnd.n5246 gnd.n5245 240.244
R13933 gnd.n5267 gnd.n5266 240.244
R13934 gnd.n1257 gnd.n1243 240.244
R13935 gnd.n5043 gnd.n1244 240.244
R13936 gnd.n5094 gnd.n5043 240.244
R13937 gnd.n5094 gnd.n5086 240.244
R13938 gnd.n5110 gnd.n5086 240.244
R13939 gnd.n5110 gnd.n5082 240.244
R13940 gnd.n5116 gnd.n5082 240.244
R13941 gnd.n5116 gnd.n5074 240.244
R13942 gnd.n5131 gnd.n5074 240.244
R13943 gnd.n5131 gnd.n5069 240.244
R13944 gnd.n5138 gnd.n5069 240.244
R13945 gnd.n5138 gnd.n5060 240.244
R13946 gnd.n5060 gnd.n1079 240.244
R13947 gnd.n5617 gnd.n1079 240.244
R13948 gnd.n5617 gnd.n1080 240.244
R13949 gnd.n1080 gnd.n1071 240.244
R13950 gnd.n1071 gnd.n1063 240.244
R13951 gnd.n1063 gnd.n1005 240.244
R13952 gnd.n5599 gnd.n1005 240.244
R13953 gnd.n5599 gnd.n998 240.244
R13954 gnd.n5602 gnd.n998 240.244
R13955 gnd.n5602 gnd.n969 240.244
R13956 gnd.n969 gnd.n957 240.244
R13957 gnd.n5724 gnd.n957 240.244
R13958 gnd.n5724 gnd.n958 240.244
R13959 gnd.n958 gnd.n954 240.244
R13960 gnd.n954 gnd.n933 240.244
R13961 gnd.n5731 gnd.n933 240.244
R13962 gnd.n5731 gnd.n926 240.244
R13963 gnd.n5738 gnd.n926 240.244
R13964 gnd.n5738 gnd.n901 240.244
R13965 gnd.n901 gnd.n892 240.244
R13966 gnd.n5807 gnd.n892 240.244
R13967 gnd.n5807 gnd.n886 240.244
R13968 gnd.n5841 gnd.n886 240.244
R13969 gnd.n5841 gnd.n887 240.244
R13970 gnd.n887 gnd.n879 240.244
R13971 gnd.n879 gnd.n864 240.244
R13972 gnd.n864 gnd.n856 240.244
R13973 gnd.n5820 gnd.n856 240.244
R13974 gnd.n5820 gnd.n847 240.244
R13975 gnd.n847 gnd.n837 240.244
R13976 gnd.n5823 gnd.n837 240.244
R13977 gnd.n5823 gnd.n819 240.244
R13978 gnd.n819 gnd.n812 240.244
R13979 gnd.n5953 gnd.n812 240.244
R13980 gnd.n5953 gnd.n804 240.244
R13981 gnd.n804 gnd.n795 240.244
R13982 gnd.n6049 gnd.n795 240.244
R13983 gnd.n6049 gnd.n786 240.244
R13984 gnd.n786 gnd.n778 240.244
R13985 gnd.n778 gnd.n772 240.244
R13986 gnd.n5959 gnd.n772 240.244
R13987 gnd.n5959 gnd.n763 240.244
R13988 gnd.n5962 gnd.n763 240.244
R13989 gnd.n5963 gnd.n5962 240.244
R13990 gnd.n5963 gnd.n742 240.244
R13991 gnd.n5964 gnd.n742 240.244
R13992 gnd.n5964 gnd.n735 240.244
R13993 gnd.n735 gnd.n726 240.244
R13994 gnd.n726 gnd.n717 240.244
R13995 gnd.n6011 gnd.n717 240.244
R13996 gnd.n6011 gnd.n708 240.244
R13997 gnd.n6014 gnd.n708 240.244
R13998 gnd.n6015 gnd.n6014 240.244
R13999 gnd.n6016 gnd.n6015 240.244
R14000 gnd.n6016 gnd.n655 240.244
R14001 gnd.n655 gnd.n646 240.244
R14002 gnd.n646 gnd.n635 240.244
R14003 gnd.n6373 gnd.n635 240.244
R14004 gnd.n6373 gnd.n630 240.244
R14005 gnd.n6380 gnd.n630 240.244
R14006 gnd.n6380 gnd.n621 240.244
R14007 gnd.n621 gnd.n610 240.244
R14008 gnd.n6403 gnd.n610 240.244
R14009 gnd.n6403 gnd.n605 240.244
R14010 gnd.n6410 gnd.n605 240.244
R14011 gnd.n6410 gnd.n596 240.244
R14012 gnd.n596 gnd.n584 240.244
R14013 gnd.n6433 gnd.n584 240.244
R14014 gnd.n6433 gnd.n579 240.244
R14015 gnd.n6440 gnd.n579 240.244
R14016 gnd.n6440 gnd.n426 240.244
R14017 gnd.n6471 gnd.n6470 240.244
R14018 gnd.n6474 gnd.n6473 240.244
R14019 gnd.n6481 gnd.n6480 240.244
R14020 gnd.n6484 gnd.n6483 240.244
R14021 gnd.n6486 gnd.n6485 240.244
R14022 gnd.n6497 gnd.n6496 240.244
R14023 gnd.n6507 gnd.n6506 240.244
R14024 gnd.n6509 gnd.n6508 240.244
R14025 gnd.n6517 gnd.n6516 240.244
R14026 gnd.n6527 gnd.n6526 240.244
R14027 gnd.n6529 gnd.n6528 240.244
R14028 gnd.n6703 gnd.n443 240.244
R14029 gnd.n6703 gnd.n444 240.244
R14030 gnd.n440 gnd.n425 240.244
R14031 gnd.n1015 gnd.n1014 240.132
R14032 gnd.n6204 gnd.n6203 240.132
R14033 gnd.n2738 gnd.n1687 225.874
R14034 gnd.n2738 gnd.n2737 225.874
R14035 gnd.n2737 gnd.n2736 225.874
R14036 gnd.n2736 gnd.n1688 225.874
R14037 gnd.n2730 gnd.n1688 225.874
R14038 gnd.n2730 gnd.n2729 225.874
R14039 gnd.n2729 gnd.n2728 225.874
R14040 gnd.n2728 gnd.n1696 225.874
R14041 gnd.n2722 gnd.n1696 225.874
R14042 gnd.n2722 gnd.n2721 225.874
R14043 gnd.n2721 gnd.n2720 225.874
R14044 gnd.n2720 gnd.n1704 225.874
R14045 gnd.n2714 gnd.n1704 225.874
R14046 gnd.n2714 gnd.n2713 225.874
R14047 gnd.n2713 gnd.n2712 225.874
R14048 gnd.n2712 gnd.n1712 225.874
R14049 gnd.n2706 gnd.n1712 225.874
R14050 gnd.n2706 gnd.n2705 225.874
R14051 gnd.n2705 gnd.n2704 225.874
R14052 gnd.n2704 gnd.n1720 225.874
R14053 gnd.n2698 gnd.n1720 225.874
R14054 gnd.n2698 gnd.n2697 225.874
R14055 gnd.n2697 gnd.n2696 225.874
R14056 gnd.n2696 gnd.n1728 225.874
R14057 gnd.n2690 gnd.n1728 225.874
R14058 gnd.n2690 gnd.n2689 225.874
R14059 gnd.n2689 gnd.n2688 225.874
R14060 gnd.n2688 gnd.n1736 225.874
R14061 gnd.n2682 gnd.n1736 225.874
R14062 gnd.n2682 gnd.n2681 225.874
R14063 gnd.n2681 gnd.n2680 225.874
R14064 gnd.n2680 gnd.n1744 225.874
R14065 gnd.n2674 gnd.n1744 225.874
R14066 gnd.n2674 gnd.n2673 225.874
R14067 gnd.n2673 gnd.n2672 225.874
R14068 gnd.n2672 gnd.n1752 225.874
R14069 gnd.n2666 gnd.n1752 225.874
R14070 gnd.n2666 gnd.n2665 225.874
R14071 gnd.n2665 gnd.n2664 225.874
R14072 gnd.n2664 gnd.n1760 225.874
R14073 gnd.n2658 gnd.n1760 225.874
R14074 gnd.n2658 gnd.n2657 225.874
R14075 gnd.n2657 gnd.n2656 225.874
R14076 gnd.n2656 gnd.n1768 225.874
R14077 gnd.n2650 gnd.n1768 225.874
R14078 gnd.n2650 gnd.n2649 225.874
R14079 gnd.n2649 gnd.n2648 225.874
R14080 gnd.n2648 gnd.n1776 225.874
R14081 gnd.n2642 gnd.n1776 225.874
R14082 gnd.n2642 gnd.n2641 225.874
R14083 gnd.n2641 gnd.n2640 225.874
R14084 gnd.n2640 gnd.n1784 225.874
R14085 gnd.n2634 gnd.n1784 225.874
R14086 gnd.n2634 gnd.n2633 225.874
R14087 gnd.n2633 gnd.n2632 225.874
R14088 gnd.n2632 gnd.n1792 225.874
R14089 gnd.n2626 gnd.n1792 225.874
R14090 gnd.n2626 gnd.n2625 225.874
R14091 gnd.n2625 gnd.n2624 225.874
R14092 gnd.n2624 gnd.n1800 225.874
R14093 gnd.n2618 gnd.n1800 225.874
R14094 gnd.n2618 gnd.n2617 225.874
R14095 gnd.n2617 gnd.n2616 225.874
R14096 gnd.n2616 gnd.n1808 225.874
R14097 gnd.n2610 gnd.n1808 225.874
R14098 gnd.n2610 gnd.n2609 225.874
R14099 gnd.n2609 gnd.n2608 225.874
R14100 gnd.n2608 gnd.n1816 225.874
R14101 gnd.n2602 gnd.n1816 225.874
R14102 gnd.n2602 gnd.n2601 225.874
R14103 gnd.n2601 gnd.n2600 225.874
R14104 gnd.n2600 gnd.n1824 225.874
R14105 gnd.n2594 gnd.n1824 225.874
R14106 gnd.n2594 gnd.n2593 225.874
R14107 gnd.n2593 gnd.n2592 225.874
R14108 gnd.n2592 gnd.n1832 225.874
R14109 gnd.n2586 gnd.n1832 225.874
R14110 gnd.n2586 gnd.n2585 225.874
R14111 gnd.n2585 gnd.n2584 225.874
R14112 gnd.n2584 gnd.n1840 225.874
R14113 gnd.n2578 gnd.n1840 225.874
R14114 gnd.n2578 gnd.n2577 225.874
R14115 gnd.n2577 gnd.n2576 225.874
R14116 gnd.n2576 gnd.n1848 225.874
R14117 gnd.n2570 gnd.n1848 225.874
R14118 gnd.n2570 gnd.n2569 225.874
R14119 gnd.n2569 gnd.n2568 225.874
R14120 gnd.n2568 gnd.n1856 225.874
R14121 gnd.n2562 gnd.n1856 225.874
R14122 gnd.n2562 gnd.n2561 225.874
R14123 gnd.n2561 gnd.n2560 225.874
R14124 gnd.n2560 gnd.n1864 225.874
R14125 gnd.n2554 gnd.n1864 225.874
R14126 gnd.n2554 gnd.n2553 225.874
R14127 gnd.n2553 gnd.n2552 225.874
R14128 gnd.n2552 gnd.n1872 225.874
R14129 gnd.n2546 gnd.n1872 225.874
R14130 gnd.n2546 gnd.n2545 225.874
R14131 gnd.n2545 gnd.n2544 225.874
R14132 gnd.n2544 gnd.n1880 225.874
R14133 gnd.n2538 gnd.n1880 225.874
R14134 gnd.n2538 gnd.n2537 225.874
R14135 gnd.n2537 gnd.n2536 225.874
R14136 gnd.n2536 gnd.n1888 225.874
R14137 gnd.n2530 gnd.n1888 225.874
R14138 gnd.n2530 gnd.n2529 225.874
R14139 gnd.n2529 gnd.n2528 225.874
R14140 gnd.n2528 gnd.n1896 225.874
R14141 gnd.n2522 gnd.n1896 225.874
R14142 gnd.n2522 gnd.n2521 225.874
R14143 gnd.n2521 gnd.n2520 225.874
R14144 gnd.n2520 gnd.n1904 225.874
R14145 gnd.n2514 gnd.n1904 225.874
R14146 gnd.n2514 gnd.n2513 225.874
R14147 gnd.n2513 gnd.n2512 225.874
R14148 gnd.n2512 gnd.n1912 225.874
R14149 gnd.n2506 gnd.n1912 225.874
R14150 gnd.n2506 gnd.n2505 225.874
R14151 gnd.n2505 gnd.n2504 225.874
R14152 gnd.n2504 gnd.n1920 225.874
R14153 gnd.n2498 gnd.n1920 225.874
R14154 gnd.n2498 gnd.n2497 225.874
R14155 gnd.n2497 gnd.n2496 225.874
R14156 gnd.n2496 gnd.n1928 225.874
R14157 gnd.n2490 gnd.n1928 225.874
R14158 gnd.n2490 gnd.n2489 225.874
R14159 gnd.n2489 gnd.n2488 225.874
R14160 gnd.n2488 gnd.n1936 225.874
R14161 gnd.n2482 gnd.n1936 225.874
R14162 gnd.n2482 gnd.n2481 225.874
R14163 gnd.n2481 gnd.n2480 225.874
R14164 gnd.n2480 gnd.n1944 225.874
R14165 gnd.n2474 gnd.n1944 225.874
R14166 gnd.n2474 gnd.n2473 225.874
R14167 gnd.n2473 gnd.n2472 225.874
R14168 gnd.n2472 gnd.n1952 225.874
R14169 gnd.n2466 gnd.n1952 225.874
R14170 gnd.n2466 gnd.n2465 225.874
R14171 gnd.n2465 gnd.n2464 225.874
R14172 gnd.n2464 gnd.n1960 225.874
R14173 gnd.n2458 gnd.n1960 225.874
R14174 gnd.n2458 gnd.n2457 225.874
R14175 gnd.n2457 gnd.n2456 225.874
R14176 gnd.n2456 gnd.n1968 225.874
R14177 gnd.n2450 gnd.n1968 225.874
R14178 gnd.n2450 gnd.n2449 225.874
R14179 gnd.n2449 gnd.n2448 225.874
R14180 gnd.n2448 gnd.n1976 225.874
R14181 gnd.n2442 gnd.n1976 225.874
R14182 gnd.n2442 gnd.n2441 225.874
R14183 gnd.n2441 gnd.n2440 225.874
R14184 gnd.n2440 gnd.n1984 225.874
R14185 gnd.n2434 gnd.n1984 225.874
R14186 gnd.n2434 gnd.n2433 225.874
R14187 gnd.n2433 gnd.n2432 225.874
R14188 gnd.n2432 gnd.n1992 225.874
R14189 gnd.n2426 gnd.n1992 225.874
R14190 gnd.n2426 gnd.n2425 225.874
R14191 gnd.n2425 gnd.n2424 225.874
R14192 gnd.n2424 gnd.n2000 225.874
R14193 gnd.n2418 gnd.n2000 225.874
R14194 gnd.n2418 gnd.n2417 225.874
R14195 gnd.n2417 gnd.n2416 225.874
R14196 gnd.n2416 gnd.n2008 225.874
R14197 gnd.n2410 gnd.n2008 225.874
R14198 gnd.n2410 gnd.n2409 225.874
R14199 gnd.n2409 gnd.n2408 225.874
R14200 gnd.n2408 gnd.n2016 225.874
R14201 gnd.n2402 gnd.n2016 225.874
R14202 gnd.n2402 gnd.n2401 225.874
R14203 gnd.n2401 gnd.n2400 225.874
R14204 gnd.n2400 gnd.n2024 225.874
R14205 gnd.n2394 gnd.n2024 225.874
R14206 gnd.n2394 gnd.n2393 225.874
R14207 gnd.n2393 gnd.n2392 225.874
R14208 gnd.n2392 gnd.n2032 225.874
R14209 gnd.n2386 gnd.n2032 225.874
R14210 gnd.n2386 gnd.n2385 225.874
R14211 gnd.n2385 gnd.n2384 225.874
R14212 gnd.n2384 gnd.n2040 225.874
R14213 gnd.n2378 gnd.n2040 225.874
R14214 gnd.n3519 gnd.t128 224.174
R14215 gnd.n3110 gnd.t114 224.174
R14216 gnd.n526 gnd.n469 199.319
R14217 gnd.n526 gnd.n470 199.319
R14218 gnd.n5407 gnd.n1150 199.319
R14219 gnd.n1155 gnd.n1150 199.319
R14220 gnd.n1016 gnd.n1013 186.49
R14221 gnd.n6205 gnd.n6202 186.49
R14222 gnd.n4224 gnd.n4223 185
R14223 gnd.n4222 gnd.n4221 185
R14224 gnd.n4201 gnd.n4200 185
R14225 gnd.n4216 gnd.n4215 185
R14226 gnd.n4214 gnd.n4213 185
R14227 gnd.n4205 gnd.n4204 185
R14228 gnd.n4208 gnd.n4207 185
R14229 gnd.n4192 gnd.n4191 185
R14230 gnd.n4190 gnd.n4189 185
R14231 gnd.n4169 gnd.n4168 185
R14232 gnd.n4184 gnd.n4183 185
R14233 gnd.n4182 gnd.n4181 185
R14234 gnd.n4173 gnd.n4172 185
R14235 gnd.n4176 gnd.n4175 185
R14236 gnd.n4160 gnd.n4159 185
R14237 gnd.n4158 gnd.n4157 185
R14238 gnd.n4137 gnd.n4136 185
R14239 gnd.n4152 gnd.n4151 185
R14240 gnd.n4150 gnd.n4149 185
R14241 gnd.n4141 gnd.n4140 185
R14242 gnd.n4144 gnd.n4143 185
R14243 gnd.n4129 gnd.n4128 185
R14244 gnd.n4127 gnd.n4126 185
R14245 gnd.n4106 gnd.n4105 185
R14246 gnd.n4121 gnd.n4120 185
R14247 gnd.n4119 gnd.n4118 185
R14248 gnd.n4110 gnd.n4109 185
R14249 gnd.n4113 gnd.n4112 185
R14250 gnd.n4097 gnd.n4096 185
R14251 gnd.n4095 gnd.n4094 185
R14252 gnd.n4074 gnd.n4073 185
R14253 gnd.n4089 gnd.n4088 185
R14254 gnd.n4087 gnd.n4086 185
R14255 gnd.n4078 gnd.n4077 185
R14256 gnd.n4081 gnd.n4080 185
R14257 gnd.n4065 gnd.n4064 185
R14258 gnd.n4063 gnd.n4062 185
R14259 gnd.n4042 gnd.n4041 185
R14260 gnd.n4057 gnd.n4056 185
R14261 gnd.n4055 gnd.n4054 185
R14262 gnd.n4046 gnd.n4045 185
R14263 gnd.n4049 gnd.n4048 185
R14264 gnd.n4033 gnd.n4032 185
R14265 gnd.n4031 gnd.n4030 185
R14266 gnd.n4010 gnd.n4009 185
R14267 gnd.n4025 gnd.n4024 185
R14268 gnd.n4023 gnd.n4022 185
R14269 gnd.n4014 gnd.n4013 185
R14270 gnd.n4017 gnd.n4016 185
R14271 gnd.n4002 gnd.n4001 185
R14272 gnd.n4000 gnd.n3999 185
R14273 gnd.n3979 gnd.n3978 185
R14274 gnd.n3994 gnd.n3993 185
R14275 gnd.n3992 gnd.n3991 185
R14276 gnd.n3983 gnd.n3982 185
R14277 gnd.n3986 gnd.n3985 185
R14278 gnd.n3520 gnd.t127 178.987
R14279 gnd.n3111 gnd.t115 178.987
R14280 gnd.n1 gnd.t314 170.774
R14281 gnd.n7 gnd.t138 170.103
R14282 gnd.n6 gnd.t146 170.103
R14283 gnd.n5 gnd.t150 170.103
R14284 gnd.n4 gnd.t148 170.103
R14285 gnd.n3 gnd.t6 170.103
R14286 gnd.n2 gnd.t158 170.103
R14287 gnd.n1 gnd.t140 170.103
R14288 gnd.n6276 gnd.n6275 163.367
R14289 gnd.n6272 gnd.n6271 163.367
R14290 gnd.n6268 gnd.n6267 163.367
R14291 gnd.n6264 gnd.n6263 163.367
R14292 gnd.n6260 gnd.n6259 163.367
R14293 gnd.n6256 gnd.n6255 163.367
R14294 gnd.n6252 gnd.n6251 163.367
R14295 gnd.n6248 gnd.n6247 163.367
R14296 gnd.n6244 gnd.n6243 163.367
R14297 gnd.n6240 gnd.n6239 163.367
R14298 gnd.n6236 gnd.n6235 163.367
R14299 gnd.n6232 gnd.n6231 163.367
R14300 gnd.n6228 gnd.n6227 163.367
R14301 gnd.n6224 gnd.n6223 163.367
R14302 gnd.n6219 gnd.n6218 163.367
R14303 gnd.n6215 gnd.n6214 163.367
R14304 gnd.n6349 gnd.n6348 163.367
R14305 gnd.n6345 gnd.n6344 163.367
R14306 gnd.n6340 gnd.n6339 163.367
R14307 gnd.n6336 gnd.n6335 163.367
R14308 gnd.n6332 gnd.n6331 163.367
R14309 gnd.n6328 gnd.n6327 163.367
R14310 gnd.n6324 gnd.n6323 163.367
R14311 gnd.n6320 gnd.n6319 163.367
R14312 gnd.n6316 gnd.n6315 163.367
R14313 gnd.n6312 gnd.n6311 163.367
R14314 gnd.n6308 gnd.n6307 163.367
R14315 gnd.n6304 gnd.n6303 163.367
R14316 gnd.n6300 gnd.n6299 163.367
R14317 gnd.n6296 gnd.n6295 163.367
R14318 gnd.n6292 gnd.n6291 163.367
R14319 gnd.n6288 gnd.n6287 163.367
R14320 gnd.n5596 gnd.n1006 163.367
R14321 gnd.n5596 gnd.n997 163.367
R14322 gnd.n997 gnd.n990 163.367
R14323 gnd.n5675 gnd.n990 163.367
R14324 gnd.n5676 gnd.n5675 163.367
R14325 gnd.n5676 gnd.n970 163.367
R14326 gnd.n5692 gnd.n970 163.367
R14327 gnd.n5692 gnd.n988 163.367
R14328 gnd.n5688 gnd.n988 163.367
R14329 gnd.n5688 gnd.n979 163.367
R14330 gnd.n5685 gnd.n979 163.367
R14331 gnd.n5685 gnd.n5684 163.367
R14332 gnd.n5684 gnd.n934 163.367
R14333 gnd.n943 gnd.n934 163.367
R14334 gnd.n5748 gnd.n943 163.367
R14335 gnd.n5748 gnd.n944 163.367
R14336 gnd.n5744 gnd.n944 163.367
R14337 gnd.n5744 gnd.n948 163.367
R14338 gnd.n948 gnd.n902 163.367
R14339 gnd.n911 gnd.n902 163.367
R14340 gnd.n5790 gnd.n911 163.367
R14341 gnd.n5790 gnd.n912 163.367
R14342 gnd.n5786 gnd.n912 163.367
R14343 gnd.n5786 gnd.n915 163.367
R14344 gnd.n915 gnd.n876 163.367
R14345 gnd.n5856 gnd.n876 163.367
R14346 gnd.n5856 gnd.n872 163.367
R14347 gnd.n5852 gnd.n872 163.367
R14348 gnd.n5852 gnd.n863 163.367
R14349 gnd.n5812 gnd.n863 163.367
R14350 gnd.n5812 gnd.n857 163.367
R14351 gnd.n5817 gnd.n857 163.367
R14352 gnd.n5817 gnd.n846 163.367
R14353 gnd.n846 gnd.n835 163.367
R14354 gnd.n5909 gnd.n835 163.367
R14355 gnd.n5909 gnd.n833 163.367
R14356 gnd.n5921 gnd.n833 163.367
R14357 gnd.n5921 gnd.n820 163.367
R14358 gnd.n5917 gnd.n820 163.367
R14359 gnd.n5917 gnd.n825 163.367
R14360 gnd.n5912 gnd.n825 163.367
R14361 gnd.n5912 gnd.n803 163.367
R14362 gnd.n6056 gnd.n803 163.367
R14363 gnd.n6056 gnd.n796 163.367
R14364 gnd.n6052 gnd.n796 163.367
R14365 gnd.n6052 gnd.n807 163.367
R14366 gnd.n5968 gnd.n807 163.367
R14367 gnd.n5968 gnd.n777 163.367
R14368 gnd.n5971 gnd.n777 163.367
R14369 gnd.n5971 gnd.n773 163.367
R14370 gnd.n5978 gnd.n773 163.367
R14371 gnd.n5978 gnd.n762 163.367
R14372 gnd.n5981 gnd.n762 163.367
R14373 gnd.n5981 gnd.n757 163.367
R14374 gnd.n5986 gnd.n757 163.367
R14375 gnd.n5986 gnd.n750 163.367
R14376 gnd.n5989 gnd.n750 163.367
R14377 gnd.n5989 gnd.n743 163.367
R14378 gnd.n5992 gnd.n743 163.367
R14379 gnd.n5992 gnd.n734 163.367
R14380 gnd.n734 gnd.n725 163.367
R14381 gnd.n727 gnd.n725 163.367
R14382 gnd.n727 gnd.n718 163.367
R14383 gnd.n6008 gnd.n718 163.367
R14384 gnd.n6008 gnd.n5967 163.367
R14385 gnd.n6004 gnd.n5967 163.367
R14386 gnd.n6004 gnd.n6003 163.367
R14387 gnd.n6003 gnd.n699 163.367
R14388 gnd.n699 gnd.n693 163.367
R14389 gnd.n6283 gnd.n693 163.367
R14390 gnd.n5652 gnd.n1030 163.367
R14391 gnd.n1090 gnd.n1030 163.367
R14392 gnd.n1094 gnd.n1093 163.367
R14393 gnd.n1098 gnd.n1097 163.367
R14394 gnd.n1102 gnd.n1101 163.367
R14395 gnd.n1106 gnd.n1105 163.367
R14396 gnd.n1110 gnd.n1109 163.367
R14397 gnd.n1114 gnd.n1113 163.367
R14398 gnd.n1118 gnd.n1117 163.367
R14399 gnd.n1122 gnd.n1121 163.367
R14400 gnd.n1126 gnd.n1125 163.367
R14401 gnd.n1130 gnd.n1129 163.367
R14402 gnd.n1134 gnd.n1133 163.367
R14403 gnd.n1138 gnd.n1137 163.367
R14404 gnd.n1142 gnd.n1141 163.367
R14405 gnd.n1146 gnd.n1145 163.367
R14406 gnd.n5527 gnd.n5526 163.367
R14407 gnd.n5531 gnd.n5530 163.367
R14408 gnd.n5536 gnd.n5535 163.367
R14409 gnd.n5540 gnd.n5539 163.367
R14410 gnd.n5544 gnd.n5543 163.367
R14411 gnd.n5548 gnd.n5547 163.367
R14412 gnd.n5552 gnd.n5551 163.367
R14413 gnd.n5556 gnd.n5555 163.367
R14414 gnd.n5560 gnd.n5559 163.367
R14415 gnd.n5564 gnd.n5563 163.367
R14416 gnd.n5568 gnd.n5567 163.367
R14417 gnd.n5572 gnd.n5571 163.367
R14418 gnd.n5576 gnd.n5575 163.367
R14419 gnd.n5580 gnd.n5579 163.367
R14420 gnd.n5584 gnd.n5583 163.367
R14421 gnd.n5588 gnd.n5587 163.367
R14422 gnd.n5657 gnd.n995 163.367
R14423 gnd.n5669 gnd.n995 163.367
R14424 gnd.n5669 gnd.n993 163.367
R14425 gnd.n5673 gnd.n993 163.367
R14426 gnd.n5673 gnd.n972 163.367
R14427 gnd.n5712 gnd.n972 163.367
R14428 gnd.n5712 gnd.n973 163.367
R14429 gnd.n5708 gnd.n973 163.367
R14430 gnd.n5708 gnd.n5707 163.367
R14431 gnd.n5707 gnd.n5706 163.367
R14432 gnd.n5706 gnd.n976 163.367
R14433 gnd.n976 gnd.n936 163.367
R14434 gnd.n5754 gnd.n936 163.367
R14435 gnd.n5754 gnd.n937 163.367
R14436 gnd.n5750 gnd.n937 163.367
R14437 gnd.n5750 gnd.n940 163.367
R14438 gnd.n5742 gnd.n940 163.367
R14439 gnd.n5742 gnd.n904 163.367
R14440 gnd.n5796 gnd.n904 163.367
R14441 gnd.n5796 gnd.n905 163.367
R14442 gnd.n5792 gnd.n905 163.367
R14443 gnd.n5792 gnd.n908 163.367
R14444 gnd.n5784 gnd.n908 163.367
R14445 gnd.n5784 gnd.n875 163.367
R14446 gnd.n5860 gnd.n875 163.367
R14447 gnd.n5860 gnd.n873 163.367
R14448 gnd.n5864 gnd.n873 163.367
R14449 gnd.n5864 gnd.n861 163.367
R14450 gnd.n5885 gnd.n861 163.367
R14451 gnd.n5885 gnd.n859 163.367
R14452 gnd.n5889 gnd.n859 163.367
R14453 gnd.n5889 gnd.n844 163.367
R14454 gnd.n5902 gnd.n844 163.367
R14455 gnd.n5902 gnd.n840 163.367
R14456 gnd.n5907 gnd.n840 163.367
R14457 gnd.n5907 gnd.n842 163.367
R14458 gnd.n842 gnd.n821 163.367
R14459 gnd.n5942 gnd.n821 163.367
R14460 gnd.n5942 gnd.n822 163.367
R14461 gnd.n5938 gnd.n822 163.367
R14462 gnd.n5938 gnd.n801 163.367
R14463 gnd.n6060 gnd.n801 163.367
R14464 gnd.n6060 gnd.n798 163.367
R14465 gnd.n6067 gnd.n798 163.367
R14466 gnd.n6067 gnd.n799 163.367
R14467 gnd.n6063 gnd.n799 163.367
R14468 gnd.n6063 gnd.n776 163.367
R14469 gnd.n6091 gnd.n776 163.367
R14470 gnd.n6091 gnd.n774 163.367
R14471 gnd.n6095 gnd.n774 163.367
R14472 gnd.n6095 gnd.n761 163.367
R14473 gnd.n6108 gnd.n761 163.367
R14474 gnd.n6108 gnd.n759 163.367
R14475 gnd.n6112 gnd.n759 163.367
R14476 gnd.n6112 gnd.n748 163.367
R14477 gnd.n6124 gnd.n748 163.367
R14478 gnd.n6124 gnd.n745 163.367
R14479 gnd.n6129 gnd.n745 163.367
R14480 gnd.n6129 gnd.n746 163.367
R14481 gnd.n746 gnd.n723 163.367
R14482 gnd.n6153 gnd.n723 163.367
R14483 gnd.n6153 gnd.n720 163.367
R14484 gnd.n6162 gnd.n720 163.367
R14485 gnd.n6162 gnd.n721 163.367
R14486 gnd.n6158 gnd.n721 163.367
R14487 gnd.n6158 gnd.n6157 163.367
R14488 gnd.n6157 gnd.n697 163.367
R14489 gnd.n6190 gnd.n697 163.367
R14490 gnd.n6190 gnd.n694 163.367
R14491 gnd.n6281 gnd.n694 163.367
R14492 gnd.n6211 gnd.n6210 156.462
R14493 gnd.n4164 gnd.n4132 153.042
R14494 gnd.n4228 gnd.n4227 152.079
R14495 gnd.n4196 gnd.n4195 152.079
R14496 gnd.n4164 gnd.n4163 152.079
R14497 gnd.n1021 gnd.n1020 152
R14498 gnd.n1022 gnd.n1011 152
R14499 gnd.n1024 gnd.n1023 152
R14500 gnd.n1026 gnd.n1009 152
R14501 gnd.n1028 gnd.n1027 152
R14502 gnd.n6209 gnd.n6193 152
R14503 gnd.n6201 gnd.n6194 152
R14504 gnd.n6200 gnd.n6199 152
R14505 gnd.n6198 gnd.n6195 152
R14506 gnd.n6196 gnd.t82 150.546
R14507 gnd.t168 gnd.n4206 147.661
R14508 gnd.t312 gnd.n4174 147.661
R14509 gnd.t320 gnd.n4142 147.661
R14510 gnd.t166 gnd.n4111 147.661
R14511 gnd.t322 gnd.n4079 147.661
R14512 gnd.t164 gnd.n4047 147.661
R14513 gnd.t8 gnd.n4015 147.661
R14514 gnd.t162 gnd.n3984 147.661
R14515 gnd.n689 gnd.n672 143.351
R14516 gnd.n5524 gnd.n1045 143.351
R14517 gnd.n5524 gnd.n1046 143.351
R14518 gnd.n6640 gnd.n525 133.44
R14519 gnd.n5525 gnd.n5523 133.44
R14520 gnd.n1018 gnd.t16 130.484
R14521 gnd.n1027 gnd.t132 126.766
R14522 gnd.n1025 gnd.t67 126.766
R14523 gnd.n1011 gnd.t107 126.766
R14524 gnd.n1019 gnd.t85 126.766
R14525 gnd.n6197 gnd.t104 126.766
R14526 gnd.n6199 gnd.t56 126.766
R14527 gnd.n6208 gnd.t129 126.766
R14528 gnd.n6210 gnd.t19 126.766
R14529 gnd.n4223 gnd.n4222 104.615
R14530 gnd.n4222 gnd.n4200 104.615
R14531 gnd.n4215 gnd.n4200 104.615
R14532 gnd.n4215 gnd.n4214 104.615
R14533 gnd.n4214 gnd.n4204 104.615
R14534 gnd.n4207 gnd.n4204 104.615
R14535 gnd.n4191 gnd.n4190 104.615
R14536 gnd.n4190 gnd.n4168 104.615
R14537 gnd.n4183 gnd.n4168 104.615
R14538 gnd.n4183 gnd.n4182 104.615
R14539 gnd.n4182 gnd.n4172 104.615
R14540 gnd.n4175 gnd.n4172 104.615
R14541 gnd.n4159 gnd.n4158 104.615
R14542 gnd.n4158 gnd.n4136 104.615
R14543 gnd.n4151 gnd.n4136 104.615
R14544 gnd.n4151 gnd.n4150 104.615
R14545 gnd.n4150 gnd.n4140 104.615
R14546 gnd.n4143 gnd.n4140 104.615
R14547 gnd.n4128 gnd.n4127 104.615
R14548 gnd.n4127 gnd.n4105 104.615
R14549 gnd.n4120 gnd.n4105 104.615
R14550 gnd.n4120 gnd.n4119 104.615
R14551 gnd.n4119 gnd.n4109 104.615
R14552 gnd.n4112 gnd.n4109 104.615
R14553 gnd.n4096 gnd.n4095 104.615
R14554 gnd.n4095 gnd.n4073 104.615
R14555 gnd.n4088 gnd.n4073 104.615
R14556 gnd.n4088 gnd.n4087 104.615
R14557 gnd.n4087 gnd.n4077 104.615
R14558 gnd.n4080 gnd.n4077 104.615
R14559 gnd.n4064 gnd.n4063 104.615
R14560 gnd.n4063 gnd.n4041 104.615
R14561 gnd.n4056 gnd.n4041 104.615
R14562 gnd.n4056 gnd.n4055 104.615
R14563 gnd.n4055 gnd.n4045 104.615
R14564 gnd.n4048 gnd.n4045 104.615
R14565 gnd.n4032 gnd.n4031 104.615
R14566 gnd.n4031 gnd.n4009 104.615
R14567 gnd.n4024 gnd.n4009 104.615
R14568 gnd.n4024 gnd.n4023 104.615
R14569 gnd.n4023 gnd.n4013 104.615
R14570 gnd.n4016 gnd.n4013 104.615
R14571 gnd.n4001 gnd.n4000 104.615
R14572 gnd.n4000 gnd.n3978 104.615
R14573 gnd.n3993 gnd.n3978 104.615
R14574 gnd.n3993 gnd.n3992 104.615
R14575 gnd.n3992 gnd.n3982 104.615
R14576 gnd.n3985 gnd.n3982 104.615
R14577 gnd.n3445 gnd.t62 100.632
R14578 gnd.n3066 gnd.t96 100.632
R14579 gnd.n7252 gnd.n7251 99.6594
R14580 gnd.n7247 gnd.n7068 99.6594
R14581 gnd.n7243 gnd.n7067 99.6594
R14582 gnd.n7239 gnd.n7066 99.6594
R14583 gnd.n7235 gnd.n7065 99.6594
R14584 gnd.n7231 gnd.n7064 99.6594
R14585 gnd.n7227 gnd.n7063 99.6594
R14586 gnd.n7223 gnd.n7062 99.6594
R14587 gnd.n7216 gnd.n7061 99.6594
R14588 gnd.n7212 gnd.n7060 99.6594
R14589 gnd.n7208 gnd.n7059 99.6594
R14590 gnd.n7204 gnd.n7058 99.6594
R14591 gnd.n7200 gnd.n7057 99.6594
R14592 gnd.n7196 gnd.n7056 99.6594
R14593 gnd.n7192 gnd.n7055 99.6594
R14594 gnd.n7188 gnd.n7054 99.6594
R14595 gnd.n7184 gnd.n7053 99.6594
R14596 gnd.n7180 gnd.n7052 99.6594
R14597 gnd.n7172 gnd.n7051 99.6594
R14598 gnd.n7170 gnd.n7050 99.6594
R14599 gnd.n7166 gnd.n7049 99.6594
R14600 gnd.n7162 gnd.n7048 99.6594
R14601 gnd.n7158 gnd.n7047 99.6594
R14602 gnd.n7154 gnd.n7046 99.6594
R14603 gnd.n7150 gnd.n7045 99.6594
R14604 gnd.n7146 gnd.n7044 99.6594
R14605 gnd.n7142 gnd.n7043 99.6594
R14606 gnd.n7138 gnd.n7042 99.6594
R14607 gnd.n7130 gnd.n7041 99.6594
R14608 gnd.n6692 gnd.n6691 99.6594
R14609 gnd.n6686 gnd.n458 99.6594
R14610 gnd.n6683 gnd.n459 99.6594
R14611 gnd.n6679 gnd.n460 99.6594
R14612 gnd.n6675 gnd.n461 99.6594
R14613 gnd.n6671 gnd.n462 99.6594
R14614 gnd.n6667 gnd.n463 99.6594
R14615 gnd.n6663 gnd.n464 99.6594
R14616 gnd.n6659 gnd.n465 99.6594
R14617 gnd.n6654 gnd.n466 99.6594
R14618 gnd.n6650 gnd.n467 99.6594
R14619 gnd.n6646 gnd.n468 99.6594
R14620 gnd.n6642 gnd.n469 99.6594
R14621 gnd.n6637 gnd.n471 99.6594
R14622 gnd.n6633 gnd.n472 99.6594
R14623 gnd.n6629 gnd.n473 99.6594
R14624 gnd.n6625 gnd.n474 99.6594
R14625 gnd.n6621 gnd.n475 99.6594
R14626 gnd.n6617 gnd.n476 99.6594
R14627 gnd.n6613 gnd.n477 99.6594
R14628 gnd.n6609 gnd.n478 99.6594
R14629 gnd.n6605 gnd.n479 99.6594
R14630 gnd.n6601 gnd.n480 99.6594
R14631 gnd.n6597 gnd.n481 99.6594
R14632 gnd.n6593 gnd.n482 99.6594
R14633 gnd.n6589 gnd.n483 99.6594
R14634 gnd.n6585 gnd.n484 99.6594
R14635 gnd.n6581 gnd.n485 99.6594
R14636 gnd.n5449 gnd.n5448 99.6594
R14637 gnd.n5444 gnd.n5369 99.6594
R14638 gnd.n5442 gnd.n5441 99.6594
R14639 gnd.n5437 gnd.n5376 99.6594
R14640 gnd.n5435 gnd.n5434 99.6594
R14641 gnd.n5430 gnd.n5383 99.6594
R14642 gnd.n5428 gnd.n5427 99.6594
R14643 gnd.n5423 gnd.n5390 99.6594
R14644 gnd.n5421 gnd.n5420 99.6594
R14645 gnd.n5416 gnd.n5400 99.6594
R14646 gnd.n5414 gnd.n5413 99.6594
R14647 gnd.n5409 gnd.n5406 99.6594
R14648 gnd.n1155 gnd.n1154 99.6594
R14649 gnd.n5517 gnd.n5516 99.6594
R14650 gnd.n5514 gnd.n5513 99.6594
R14651 gnd.n5509 gnd.n1164 99.6594
R14652 gnd.n5507 gnd.n5506 99.6594
R14653 gnd.n1174 gnd.n1173 99.6594
R14654 gnd.n5498 gnd.n5497 99.6594
R14655 gnd.n5495 gnd.n5494 99.6594
R14656 gnd.n5490 gnd.n1182 99.6594
R14657 gnd.n5488 gnd.n5487 99.6594
R14658 gnd.n5483 gnd.n1189 99.6594
R14659 gnd.n5481 gnd.n5480 99.6594
R14660 gnd.n5476 gnd.n1196 99.6594
R14661 gnd.n5474 gnd.n5473 99.6594
R14662 gnd.n5469 gnd.n1205 99.6594
R14663 gnd.n5467 gnd.n5466 99.6594
R14664 gnd.n4705 gnd.n4704 99.6594
R14665 gnd.n4453 gnd.n1517 99.6594
R14666 gnd.n4697 gnd.n1518 99.6594
R14667 gnd.n4693 gnd.n1519 99.6594
R14668 gnd.n4689 gnd.n1520 99.6594
R14669 gnd.n4685 gnd.n1521 99.6594
R14670 gnd.n4681 gnd.n1522 99.6594
R14671 gnd.n4677 gnd.n1523 99.6594
R14672 gnd.n4673 gnd.n1524 99.6594
R14673 gnd.n4668 gnd.n1525 99.6594
R14674 gnd.n4664 gnd.n1526 99.6594
R14675 gnd.n4660 gnd.n1527 99.6594
R14676 gnd.n4656 gnd.n1528 99.6594
R14677 gnd.n4652 gnd.n1529 99.6594
R14678 gnd.n4648 gnd.n1530 99.6594
R14679 gnd.n4644 gnd.n1531 99.6594
R14680 gnd.n4640 gnd.n1532 99.6594
R14681 gnd.n4636 gnd.n1533 99.6594
R14682 gnd.n4632 gnd.n1534 99.6594
R14683 gnd.n4628 gnd.n1535 99.6594
R14684 gnd.n4624 gnd.n1536 99.6594
R14685 gnd.n4620 gnd.n1537 99.6594
R14686 gnd.n4616 gnd.n1538 99.6594
R14687 gnd.n4612 gnd.n1539 99.6594
R14688 gnd.n4608 gnd.n1540 99.6594
R14689 gnd.n4604 gnd.n1541 99.6594
R14690 gnd.n4600 gnd.n1542 99.6594
R14691 gnd.n4596 gnd.n1543 99.6594
R14692 gnd.n4592 gnd.n1544 99.6594
R14693 gnd.n4354 gnd.n3046 99.6594
R14694 gnd.n4352 gnd.n4351 99.6594
R14695 gnd.n4347 gnd.n3053 99.6594
R14696 gnd.n4345 gnd.n4344 99.6594
R14697 gnd.n4340 gnd.n3060 99.6594
R14698 gnd.n4338 gnd.n4337 99.6594
R14699 gnd.n4333 gnd.n3069 99.6594
R14700 gnd.n4331 gnd.n4330 99.6594
R14701 gnd.n3657 gnd.n3388 99.6594
R14702 gnd.n3414 gnd.n3395 99.6594
R14703 gnd.n3416 gnd.n3396 99.6594
R14704 gnd.n3424 gnd.n3397 99.6594
R14705 gnd.n3426 gnd.n3398 99.6594
R14706 gnd.n3434 gnd.n3399 99.6594
R14707 gnd.n3436 gnd.n3400 99.6594
R14708 gnd.n3444 gnd.n3401 99.6594
R14709 gnd.n205 gnd.n184 99.6594
R14710 gnd.n211 gnd.n185 99.6594
R14711 gnd.n215 gnd.n186 99.6594
R14712 gnd.n221 gnd.n187 99.6594
R14713 gnd.n225 gnd.n188 99.6594
R14714 gnd.n231 gnd.n189 99.6594
R14715 gnd.n234 gnd.n190 99.6594
R14716 gnd.n241 gnd.n240 99.6594
R14717 gnd.n7255 gnd.n7254 99.6594
R14718 gnd.n6490 gnd.n486 99.6594
R14719 gnd.n6493 gnd.n487 99.6594
R14720 gnd.n6501 gnd.n488 99.6594
R14721 gnd.n6503 gnd.n489 99.6594
R14722 gnd.n6513 gnd.n490 99.6594
R14723 gnd.n6521 gnd.n491 99.6594
R14724 gnd.n6523 gnd.n492 99.6594
R14725 gnd.n6533 gnd.n494 99.6594
R14726 gnd.n6694 gnd.n453 99.6594
R14727 gnd.n4322 gnd.n3076 99.6594
R14728 gnd.n4320 gnd.n4319 99.6594
R14729 gnd.n4315 gnd.n3083 99.6594
R14730 gnd.n4313 gnd.n4312 99.6594
R14731 gnd.n4308 gnd.n3090 99.6594
R14732 gnd.n4306 gnd.n4305 99.6594
R14733 gnd.n4301 gnd.n3097 99.6594
R14734 gnd.n4299 gnd.n4298 99.6594
R14735 gnd.n4294 gnd.n3104 99.6594
R14736 gnd.n4292 gnd.n4291 99.6594
R14737 gnd.n4287 gnd.n3113 99.6594
R14738 gnd.n4285 gnd.n4284 99.6594
R14739 gnd.n4280 gnd.n4279 99.6594
R14740 gnd.n3572 gnd.n3571 99.6594
R14741 gnd.n3566 gnd.n3483 99.6594
R14742 gnd.n3563 gnd.n3484 99.6594
R14743 gnd.n3559 gnd.n3485 99.6594
R14744 gnd.n3555 gnd.n3486 99.6594
R14745 gnd.n3551 gnd.n3487 99.6594
R14746 gnd.n3547 gnd.n3488 99.6594
R14747 gnd.n3543 gnd.n3489 99.6594
R14748 gnd.n3539 gnd.n3490 99.6594
R14749 gnd.n3535 gnd.n3491 99.6594
R14750 gnd.n3531 gnd.n3492 99.6594
R14751 gnd.n3527 gnd.n3493 99.6594
R14752 gnd.n3574 gnd.n3482 99.6594
R14753 gnd.n5204 gnd.n5203 99.6594
R14754 gnd.n5207 gnd.n5206 99.6594
R14755 gnd.n5218 gnd.n5217 99.6594
R14756 gnd.n5227 gnd.n5226 99.6594
R14757 gnd.n5230 gnd.n5229 99.6594
R14758 gnd.n5241 gnd.n5240 99.6594
R14759 gnd.n5250 gnd.n5249 99.6594
R14760 gnd.n5253 gnd.n5252 99.6594
R14761 gnd.n5258 gnd.n5257 99.6594
R14762 gnd.n4582 gnd.n1545 99.6594
R14763 gnd.n4578 gnd.n1546 99.6594
R14764 gnd.n4574 gnd.n1547 99.6594
R14765 gnd.n4570 gnd.n1548 99.6594
R14766 gnd.n4566 gnd.n1549 99.6594
R14767 gnd.n4562 gnd.n1550 99.6594
R14768 gnd.n4558 gnd.n1551 99.6594
R14769 gnd.n4554 gnd.n1552 99.6594
R14770 gnd.n4550 gnd.n1553 99.6594
R14771 gnd.n4579 gnd.n1545 99.6594
R14772 gnd.n4575 gnd.n1546 99.6594
R14773 gnd.n4571 gnd.n1547 99.6594
R14774 gnd.n4567 gnd.n1548 99.6594
R14775 gnd.n4563 gnd.n1549 99.6594
R14776 gnd.n4559 gnd.n1550 99.6594
R14777 gnd.n4555 gnd.n1551 99.6594
R14778 gnd.n4551 gnd.n1552 99.6594
R14779 gnd.n4541 gnd.n1553 99.6594
R14780 gnd.n5257 gnd.n5256 99.6594
R14781 gnd.n5252 gnd.n5251 99.6594
R14782 gnd.n5249 gnd.n5242 99.6594
R14783 gnd.n5240 gnd.n5239 99.6594
R14784 gnd.n5229 gnd.n5228 99.6594
R14785 gnd.n5226 gnd.n5219 99.6594
R14786 gnd.n5217 gnd.n5216 99.6594
R14787 gnd.n5206 gnd.n5205 99.6594
R14788 gnd.n5203 gnd.n5193 99.6594
R14789 gnd.n3572 gnd.n3495 99.6594
R14790 gnd.n3564 gnd.n3483 99.6594
R14791 gnd.n3560 gnd.n3484 99.6594
R14792 gnd.n3556 gnd.n3485 99.6594
R14793 gnd.n3552 gnd.n3486 99.6594
R14794 gnd.n3548 gnd.n3487 99.6594
R14795 gnd.n3544 gnd.n3488 99.6594
R14796 gnd.n3540 gnd.n3489 99.6594
R14797 gnd.n3536 gnd.n3490 99.6594
R14798 gnd.n3532 gnd.n3491 99.6594
R14799 gnd.n3528 gnd.n3492 99.6594
R14800 gnd.n3524 gnd.n3493 99.6594
R14801 gnd.n3575 gnd.n3574 99.6594
R14802 gnd.n4279 gnd.n3115 99.6594
R14803 gnd.n4286 gnd.n4285 99.6594
R14804 gnd.n3113 gnd.n3105 99.6594
R14805 gnd.n4293 gnd.n4292 99.6594
R14806 gnd.n3104 gnd.n3098 99.6594
R14807 gnd.n4300 gnd.n4299 99.6594
R14808 gnd.n3097 gnd.n3091 99.6594
R14809 gnd.n4307 gnd.n4306 99.6594
R14810 gnd.n3090 gnd.n3084 99.6594
R14811 gnd.n4314 gnd.n4313 99.6594
R14812 gnd.n3083 gnd.n3077 99.6594
R14813 gnd.n4321 gnd.n4320 99.6594
R14814 gnd.n3076 gnd.n3073 99.6594
R14815 gnd.n6492 gnd.n486 99.6594
R14816 gnd.n6500 gnd.n487 99.6594
R14817 gnd.n6502 gnd.n488 99.6594
R14818 gnd.n6512 gnd.n489 99.6594
R14819 gnd.n6520 gnd.n490 99.6594
R14820 gnd.n6522 gnd.n491 99.6594
R14821 gnd.n6532 gnd.n492 99.6594
R14822 gnd.n494 gnd.n493 99.6594
R14823 gnd.n6695 gnd.n6694 99.6594
R14824 gnd.n7254 gnd.n183 99.6594
R14825 gnd.n241 gnd.n191 99.6594
R14826 gnd.n232 gnd.n190 99.6594
R14827 gnd.n224 gnd.n189 99.6594
R14828 gnd.n222 gnd.n188 99.6594
R14829 gnd.n214 gnd.n187 99.6594
R14830 gnd.n212 gnd.n186 99.6594
R14831 gnd.n204 gnd.n185 99.6594
R14832 gnd.n202 gnd.n184 99.6594
R14833 gnd.n3658 gnd.n3657 99.6594
R14834 gnd.n3417 gnd.n3395 99.6594
R14835 gnd.n3423 gnd.n3396 99.6594
R14836 gnd.n3427 gnd.n3397 99.6594
R14837 gnd.n3433 gnd.n3398 99.6594
R14838 gnd.n3437 gnd.n3399 99.6594
R14839 gnd.n3443 gnd.n3400 99.6594
R14840 gnd.n3401 gnd.n3385 99.6594
R14841 gnd.n4332 gnd.n4331 99.6594
R14842 gnd.n3069 gnd.n3061 99.6594
R14843 gnd.n4339 gnd.n4338 99.6594
R14844 gnd.n3060 gnd.n3054 99.6594
R14845 gnd.n4346 gnd.n4345 99.6594
R14846 gnd.n3053 gnd.n3047 99.6594
R14847 gnd.n4353 gnd.n4352 99.6594
R14848 gnd.n3046 gnd.n3043 99.6594
R14849 gnd.n4704 gnd.n1515 99.6594
R14850 gnd.n4698 gnd.n1517 99.6594
R14851 gnd.n4694 gnd.n1518 99.6594
R14852 gnd.n4690 gnd.n1519 99.6594
R14853 gnd.n4686 gnd.n1520 99.6594
R14854 gnd.n4682 gnd.n1521 99.6594
R14855 gnd.n4678 gnd.n1522 99.6594
R14856 gnd.n4674 gnd.n1523 99.6594
R14857 gnd.n4669 gnd.n1524 99.6594
R14858 gnd.n4665 gnd.n1525 99.6594
R14859 gnd.n4661 gnd.n1526 99.6594
R14860 gnd.n4657 gnd.n1527 99.6594
R14861 gnd.n4653 gnd.n1528 99.6594
R14862 gnd.n4649 gnd.n1529 99.6594
R14863 gnd.n4645 gnd.n1530 99.6594
R14864 gnd.n4641 gnd.n1531 99.6594
R14865 gnd.n4637 gnd.n1532 99.6594
R14866 gnd.n4633 gnd.n1533 99.6594
R14867 gnd.n4629 gnd.n1534 99.6594
R14868 gnd.n4625 gnd.n1535 99.6594
R14869 gnd.n4621 gnd.n1536 99.6594
R14870 gnd.n4617 gnd.n1537 99.6594
R14871 gnd.n4613 gnd.n1538 99.6594
R14872 gnd.n4609 gnd.n1539 99.6594
R14873 gnd.n4605 gnd.n1540 99.6594
R14874 gnd.n4601 gnd.n1541 99.6594
R14875 gnd.n4597 gnd.n1542 99.6594
R14876 gnd.n4593 gnd.n1543 99.6594
R14877 gnd.n4525 gnd.n1544 99.6594
R14878 gnd.n5468 gnd.n5467 99.6594
R14879 gnd.n1205 gnd.n1197 99.6594
R14880 gnd.n5475 gnd.n5474 99.6594
R14881 gnd.n1196 gnd.n1190 99.6594
R14882 gnd.n5482 gnd.n5481 99.6594
R14883 gnd.n1189 gnd.n1183 99.6594
R14884 gnd.n5489 gnd.n5488 99.6594
R14885 gnd.n1182 gnd.n1176 99.6594
R14886 gnd.n5496 gnd.n5495 99.6594
R14887 gnd.n5499 gnd.n5498 99.6594
R14888 gnd.n1173 gnd.n1165 99.6594
R14889 gnd.n5508 gnd.n5507 99.6594
R14890 gnd.n1164 gnd.n1158 99.6594
R14891 gnd.n5515 gnd.n5514 99.6594
R14892 gnd.n5518 gnd.n5517 99.6594
R14893 gnd.n5408 gnd.n5407 99.6594
R14894 gnd.n5406 gnd.n5401 99.6594
R14895 gnd.n5415 gnd.n5414 99.6594
R14896 gnd.n5400 gnd.n5391 99.6594
R14897 gnd.n5422 gnd.n5421 99.6594
R14898 gnd.n5390 gnd.n5384 99.6594
R14899 gnd.n5429 gnd.n5428 99.6594
R14900 gnd.n5383 gnd.n5377 99.6594
R14901 gnd.n5436 gnd.n5435 99.6594
R14902 gnd.n5376 gnd.n5370 99.6594
R14903 gnd.n5443 gnd.n5442 99.6594
R14904 gnd.n5369 gnd.n5364 99.6594
R14905 gnd.n5450 gnd.n5449 99.6594
R14906 gnd.n6692 gnd.n496 99.6594
R14907 gnd.n6684 gnd.n458 99.6594
R14908 gnd.n6680 gnd.n459 99.6594
R14909 gnd.n6676 gnd.n460 99.6594
R14910 gnd.n6672 gnd.n461 99.6594
R14911 gnd.n6668 gnd.n462 99.6594
R14912 gnd.n6664 gnd.n463 99.6594
R14913 gnd.n6660 gnd.n464 99.6594
R14914 gnd.n6655 gnd.n465 99.6594
R14915 gnd.n6651 gnd.n466 99.6594
R14916 gnd.n6647 gnd.n467 99.6594
R14917 gnd.n6643 gnd.n468 99.6594
R14918 gnd.n6638 gnd.n470 99.6594
R14919 gnd.n6634 gnd.n471 99.6594
R14920 gnd.n6630 gnd.n472 99.6594
R14921 gnd.n6626 gnd.n473 99.6594
R14922 gnd.n6622 gnd.n474 99.6594
R14923 gnd.n6618 gnd.n475 99.6594
R14924 gnd.n6614 gnd.n476 99.6594
R14925 gnd.n6610 gnd.n477 99.6594
R14926 gnd.n6606 gnd.n478 99.6594
R14927 gnd.n6602 gnd.n479 99.6594
R14928 gnd.n6598 gnd.n480 99.6594
R14929 gnd.n6594 gnd.n481 99.6594
R14930 gnd.n6590 gnd.n482 99.6594
R14931 gnd.n6586 gnd.n483 99.6594
R14932 gnd.n6582 gnd.n484 99.6594
R14933 gnd.n559 gnd.n485 99.6594
R14934 gnd.n7137 gnd.n7041 99.6594
R14935 gnd.n7141 gnd.n7042 99.6594
R14936 gnd.n7145 gnd.n7043 99.6594
R14937 gnd.n7149 gnd.n7044 99.6594
R14938 gnd.n7153 gnd.n7045 99.6594
R14939 gnd.n7157 gnd.n7046 99.6594
R14940 gnd.n7161 gnd.n7047 99.6594
R14941 gnd.n7165 gnd.n7048 99.6594
R14942 gnd.n7169 gnd.n7049 99.6594
R14943 gnd.n7173 gnd.n7050 99.6594
R14944 gnd.n7179 gnd.n7051 99.6594
R14945 gnd.n7183 gnd.n7052 99.6594
R14946 gnd.n7187 gnd.n7053 99.6594
R14947 gnd.n7191 gnd.n7054 99.6594
R14948 gnd.n7195 gnd.n7055 99.6594
R14949 gnd.n7199 gnd.n7056 99.6594
R14950 gnd.n7203 gnd.n7057 99.6594
R14951 gnd.n7207 gnd.n7058 99.6594
R14952 gnd.n7211 gnd.n7059 99.6594
R14953 gnd.n7215 gnd.n7060 99.6594
R14954 gnd.n7222 gnd.n7061 99.6594
R14955 gnd.n7226 gnd.n7062 99.6594
R14956 gnd.n7230 gnd.n7063 99.6594
R14957 gnd.n7234 gnd.n7064 99.6594
R14958 gnd.n7238 gnd.n7065 99.6594
R14959 gnd.n7242 gnd.n7066 99.6594
R14960 gnd.n7246 gnd.n7067 99.6594
R14961 gnd.n7070 gnd.n7068 99.6594
R14962 gnd.n7252 gnd.n7069 99.6594
R14963 gnd.n5329 gnd.n5328 99.6594
R14964 gnd.n1266 gnd.n1246 99.6594
R14965 gnd.n1268 gnd.n1247 99.6594
R14966 gnd.n1270 gnd.n1248 99.6594
R14967 gnd.n5197 gnd.n1249 99.6594
R14968 gnd.n5200 gnd.n1250 99.6594
R14969 gnd.n5211 gnd.n1251 99.6594
R14970 gnd.n5213 gnd.n1252 99.6594
R14971 gnd.n5223 gnd.n1253 99.6594
R14972 gnd.n5234 gnd.n1254 99.6594
R14973 gnd.n5236 gnd.n1255 99.6594
R14974 gnd.n5246 gnd.n1256 99.6594
R14975 gnd.n5267 gnd.n1258 99.6594
R14976 gnd.n5331 gnd.n1243 99.6594
R14977 gnd.n5329 gnd.n1261 99.6594
R14978 gnd.n1267 gnd.n1246 99.6594
R14979 gnd.n1269 gnd.n1247 99.6594
R14980 gnd.n5196 gnd.n1248 99.6594
R14981 gnd.n5199 gnd.n1249 99.6594
R14982 gnd.n5210 gnd.n1250 99.6594
R14983 gnd.n5212 gnd.n1251 99.6594
R14984 gnd.n5222 gnd.n1252 99.6594
R14985 gnd.n5233 gnd.n1253 99.6594
R14986 gnd.n5235 gnd.n1254 99.6594
R14987 gnd.n5245 gnd.n1255 99.6594
R14988 gnd.n5266 gnd.n1256 99.6594
R14989 gnd.n1258 gnd.n1257 99.6594
R14990 gnd.n5332 gnd.n5331 99.6594
R14991 gnd.n6470 gnd.n428 99.6594
R14992 gnd.n6474 gnd.n429 99.6594
R14993 gnd.n6480 gnd.n430 99.6594
R14994 gnd.n6483 gnd.n431 99.6594
R14995 gnd.n6485 gnd.n432 99.6594
R14996 gnd.n6496 gnd.n433 99.6594
R14997 gnd.n6506 gnd.n434 99.6594
R14998 gnd.n6508 gnd.n435 99.6594
R14999 gnd.n6516 gnd.n436 99.6594
R15000 gnd.n6526 gnd.n437 99.6594
R15001 gnd.n6528 gnd.n438 99.6594
R15002 gnd.n443 gnd.n439 99.6594
R15003 gnd.n444 gnd.n441 99.6594
R15004 gnd.n6705 gnd.n425 99.6594
R15005 gnd.n6529 gnd.n439 99.6594
R15006 gnd.n6527 gnd.n438 99.6594
R15007 gnd.n6517 gnd.n437 99.6594
R15008 gnd.n6509 gnd.n436 99.6594
R15009 gnd.n6507 gnd.n435 99.6594
R15010 gnd.n6497 gnd.n434 99.6594
R15011 gnd.n6486 gnd.n433 99.6594
R15012 gnd.n6484 gnd.n432 99.6594
R15013 gnd.n6481 gnd.n431 99.6594
R15014 gnd.n6473 gnd.n430 99.6594
R15015 gnd.n6471 gnd.n429 99.6594
R15016 gnd.n571 gnd.n428 99.6594
R15017 gnd.n6706 gnd.n6705 99.6594
R15018 gnd.n441 gnd.n440 99.6594
R15019 gnd.n5263 gnd.t66 98.63
R15020 gnd.n6696 gnd.t103 98.63
R15021 gnd.n5254 gnd.t123 98.63
R15022 gnd.n515 gnd.t100 98.63
R15023 gnd.n538 gnd.t90 98.63
R15024 gnd.n561 gnd.t37 98.63
R15025 gnd.n7132 gnd.t39 98.63
R15026 gnd.n7111 gnd.t32 98.63
R15027 gnd.n7218 gnd.t92 98.63
R15028 gnd.n180 gnd.t120 98.63
R15029 gnd.n4470 gnd.t72 98.63
R15030 gnd.n4492 gnd.t47 98.63
R15031 gnd.n4514 gnd.t78 98.63
R15032 gnd.n4542 gnd.t29 98.63
R15033 gnd.n5392 gnd.t117 98.63
R15034 gnd.n1202 gnd.t50 98.63
R15035 gnd.n1169 gnd.t80 98.63
R15036 gnd.n446 gnd.t54 98.63
R15037 gnd.n1085 gnd.t111 88.9408
R15038 gnd.n690 gnd.t24 88.9408
R15039 gnd.n1087 gnd.t44 88.933
R15040 gnd.n6212 gnd.t74 88.933
R15041 gnd.n1018 gnd.n1017 81.8399
R15042 gnd.n3446 gnd.t61 74.8376
R15043 gnd.n3067 gnd.t97 74.8376
R15044 gnd.n1086 gnd.t110 72.8438
R15045 gnd.n691 gnd.t25 72.8438
R15046 gnd.n1019 gnd.n1012 72.8411
R15047 gnd.n1025 gnd.n1010 72.8411
R15048 gnd.n6208 gnd.n6207 72.8411
R15049 gnd.n5264 gnd.t65 72.836
R15050 gnd.n1088 gnd.t43 72.836
R15051 gnd.n6213 gnd.t75 72.836
R15052 gnd.n6697 gnd.t102 72.836
R15053 gnd.n5255 gnd.t124 72.836
R15054 gnd.n516 gnd.t99 72.836
R15055 gnd.n539 gnd.t89 72.836
R15056 gnd.n562 gnd.t36 72.836
R15057 gnd.n7133 gnd.t40 72.836
R15058 gnd.n7112 gnd.t33 72.836
R15059 gnd.n7219 gnd.t93 72.836
R15060 gnd.n181 gnd.t121 72.836
R15061 gnd.n4471 gnd.t71 72.836
R15062 gnd.n4493 gnd.t46 72.836
R15063 gnd.n4515 gnd.t77 72.836
R15064 gnd.n4543 gnd.t28 72.836
R15065 gnd.n5393 gnd.t118 72.836
R15066 gnd.n1203 gnd.t51 72.836
R15067 gnd.n1170 gnd.t81 72.836
R15068 gnd.n447 gnd.t55 72.836
R15069 gnd.n6276 gnd.n656 71.676
R15070 gnd.n6272 gnd.n657 71.676
R15071 gnd.n6268 gnd.n658 71.676
R15072 gnd.n6264 gnd.n659 71.676
R15073 gnd.n6260 gnd.n660 71.676
R15074 gnd.n6256 gnd.n661 71.676
R15075 gnd.n6252 gnd.n662 71.676
R15076 gnd.n6248 gnd.n663 71.676
R15077 gnd.n6244 gnd.n664 71.676
R15078 gnd.n6240 gnd.n665 71.676
R15079 gnd.n6236 gnd.n666 71.676
R15080 gnd.n6232 gnd.n667 71.676
R15081 gnd.n6228 gnd.n668 71.676
R15082 gnd.n6224 gnd.n669 71.676
R15083 gnd.n6219 gnd.n670 71.676
R15084 gnd.n6215 gnd.n671 71.676
R15085 gnd.n6349 gnd.n689 71.676
R15086 gnd.n6345 gnd.n688 71.676
R15087 gnd.n6340 gnd.n687 71.676
R15088 gnd.n6336 gnd.n686 71.676
R15089 gnd.n6332 gnd.n685 71.676
R15090 gnd.n6328 gnd.n684 71.676
R15091 gnd.n6324 gnd.n683 71.676
R15092 gnd.n6320 gnd.n682 71.676
R15093 gnd.n6316 gnd.n681 71.676
R15094 gnd.n6312 gnd.n680 71.676
R15095 gnd.n6308 gnd.n679 71.676
R15096 gnd.n6304 gnd.n678 71.676
R15097 gnd.n6300 gnd.n677 71.676
R15098 gnd.n6296 gnd.n676 71.676
R15099 gnd.n6292 gnd.n675 71.676
R15100 gnd.n6288 gnd.n674 71.676
R15101 gnd.n6284 gnd.n673 71.676
R15102 gnd.n5651 gnd.n1008 71.676
R15103 gnd.n1090 gnd.n1031 71.676
R15104 gnd.n1094 gnd.n1032 71.676
R15105 gnd.n1098 gnd.n1033 71.676
R15106 gnd.n1102 gnd.n1034 71.676
R15107 gnd.n1106 gnd.n1035 71.676
R15108 gnd.n1110 gnd.n1036 71.676
R15109 gnd.n1114 gnd.n1037 71.676
R15110 gnd.n1118 gnd.n1038 71.676
R15111 gnd.n1122 gnd.n1039 71.676
R15112 gnd.n1126 gnd.n1040 71.676
R15113 gnd.n1130 gnd.n1041 71.676
R15114 gnd.n1134 gnd.n1042 71.676
R15115 gnd.n1138 gnd.n1043 71.676
R15116 gnd.n1142 gnd.n1044 71.676
R15117 gnd.n1146 gnd.n1045 71.676
R15118 gnd.n5527 gnd.n1047 71.676
R15119 gnd.n5531 gnd.n1048 71.676
R15120 gnd.n5536 gnd.n1049 71.676
R15121 gnd.n5540 gnd.n1050 71.676
R15122 gnd.n5544 gnd.n1051 71.676
R15123 gnd.n5548 gnd.n1052 71.676
R15124 gnd.n5552 gnd.n1053 71.676
R15125 gnd.n5556 gnd.n1054 71.676
R15126 gnd.n5560 gnd.n1055 71.676
R15127 gnd.n5564 gnd.n1056 71.676
R15128 gnd.n5568 gnd.n1057 71.676
R15129 gnd.n5572 gnd.n1058 71.676
R15130 gnd.n5576 gnd.n1059 71.676
R15131 gnd.n5580 gnd.n1060 71.676
R15132 gnd.n5584 gnd.n1061 71.676
R15133 gnd.n5588 gnd.n1062 71.676
R15134 gnd.n5652 gnd.n5651 71.676
R15135 gnd.n1093 gnd.n1031 71.676
R15136 gnd.n1097 gnd.n1032 71.676
R15137 gnd.n1101 gnd.n1033 71.676
R15138 gnd.n1105 gnd.n1034 71.676
R15139 gnd.n1109 gnd.n1035 71.676
R15140 gnd.n1113 gnd.n1036 71.676
R15141 gnd.n1117 gnd.n1037 71.676
R15142 gnd.n1121 gnd.n1038 71.676
R15143 gnd.n1125 gnd.n1039 71.676
R15144 gnd.n1129 gnd.n1040 71.676
R15145 gnd.n1133 gnd.n1041 71.676
R15146 gnd.n1137 gnd.n1042 71.676
R15147 gnd.n1141 gnd.n1043 71.676
R15148 gnd.n1145 gnd.n1044 71.676
R15149 gnd.n5526 gnd.n1046 71.676
R15150 gnd.n5530 gnd.n1047 71.676
R15151 gnd.n5535 gnd.n1048 71.676
R15152 gnd.n5539 gnd.n1049 71.676
R15153 gnd.n5543 gnd.n1050 71.676
R15154 gnd.n5547 gnd.n1051 71.676
R15155 gnd.n5551 gnd.n1052 71.676
R15156 gnd.n5555 gnd.n1053 71.676
R15157 gnd.n5559 gnd.n1054 71.676
R15158 gnd.n5563 gnd.n1055 71.676
R15159 gnd.n5567 gnd.n1056 71.676
R15160 gnd.n5571 gnd.n1057 71.676
R15161 gnd.n5575 gnd.n1058 71.676
R15162 gnd.n5579 gnd.n1059 71.676
R15163 gnd.n5583 gnd.n1060 71.676
R15164 gnd.n5587 gnd.n1061 71.676
R15165 gnd.n5590 gnd.n1062 71.676
R15166 gnd.n6287 gnd.n673 71.676
R15167 gnd.n6291 gnd.n674 71.676
R15168 gnd.n6295 gnd.n675 71.676
R15169 gnd.n6299 gnd.n676 71.676
R15170 gnd.n6303 gnd.n677 71.676
R15171 gnd.n6307 gnd.n678 71.676
R15172 gnd.n6311 gnd.n679 71.676
R15173 gnd.n6315 gnd.n680 71.676
R15174 gnd.n6319 gnd.n681 71.676
R15175 gnd.n6323 gnd.n682 71.676
R15176 gnd.n6327 gnd.n683 71.676
R15177 gnd.n6331 gnd.n684 71.676
R15178 gnd.n6335 gnd.n685 71.676
R15179 gnd.n6339 gnd.n686 71.676
R15180 gnd.n6344 gnd.n687 71.676
R15181 gnd.n6348 gnd.n688 71.676
R15182 gnd.n6214 gnd.n672 71.676
R15183 gnd.n6218 gnd.n671 71.676
R15184 gnd.n6223 gnd.n670 71.676
R15185 gnd.n6227 gnd.n669 71.676
R15186 gnd.n6231 gnd.n668 71.676
R15187 gnd.n6235 gnd.n667 71.676
R15188 gnd.n6239 gnd.n666 71.676
R15189 gnd.n6243 gnd.n665 71.676
R15190 gnd.n6247 gnd.n664 71.676
R15191 gnd.n6251 gnd.n663 71.676
R15192 gnd.n6255 gnd.n662 71.676
R15193 gnd.n6259 gnd.n661 71.676
R15194 gnd.n6263 gnd.n660 71.676
R15195 gnd.n6267 gnd.n659 71.676
R15196 gnd.n6271 gnd.n658 71.676
R15197 gnd.n6275 gnd.n657 71.676
R15198 gnd.n695 gnd.n656 71.676
R15199 gnd.n8 gnd.t152 69.1507
R15200 gnd.n14 gnd.t318 68.4792
R15201 gnd.n13 gnd.t307 68.4792
R15202 gnd.n12 gnd.t3 68.4792
R15203 gnd.n11 gnd.t316 68.4792
R15204 gnd.n10 gnd.t160 68.4792
R15205 gnd.n9 gnd.t154 68.4792
R15206 gnd.n8 gnd.t310 68.4792
R15207 gnd.n3573 gnd.n3477 64.369
R15208 gnd.n5533 gnd.n1086 59.5399
R15209 gnd.n6342 gnd.n691 59.5399
R15210 gnd.n1089 gnd.n1088 59.5399
R15211 gnd.n6221 gnd.n6213 59.5399
R15212 gnd.n5655 gnd.n1028 59.1804
R15213 gnd.n4362 gnd.n3036 57.3586
R15214 gnd.n3232 gnd.t227 56.407
R15215 gnd.n3197 gnd.t274 56.407
R15216 gnd.n3208 gnd.t186 56.407
R15217 gnd.n3220 gnd.t266 56.407
R15218 gnd.n52 gnd.t202 56.407
R15219 gnd.n17 gnd.t193 56.407
R15220 gnd.n28 gnd.t283 56.407
R15221 gnd.n40 gnd.t241 56.407
R15222 gnd.n3241 gnd.t253 55.8337
R15223 gnd.n3206 gnd.t182 55.8337
R15224 gnd.n3217 gnd.t285 55.8337
R15225 gnd.n3229 gnd.t187 55.8337
R15226 gnd.n61 gnd.t225 55.8337
R15227 gnd.n26 gnd.t217 55.8337
R15228 gnd.n37 gnd.t265 55.8337
R15229 gnd.n49 gnd.t262 55.8337
R15230 gnd.n1016 gnd.n1015 54.358
R15231 gnd.n6205 gnd.n6204 54.358
R15232 gnd.n3232 gnd.n3231 53.0052
R15233 gnd.n3234 gnd.n3233 53.0052
R15234 gnd.n3236 gnd.n3235 53.0052
R15235 gnd.n3238 gnd.n3237 53.0052
R15236 gnd.n3240 gnd.n3239 53.0052
R15237 gnd.n3197 gnd.n3196 53.0052
R15238 gnd.n3199 gnd.n3198 53.0052
R15239 gnd.n3201 gnd.n3200 53.0052
R15240 gnd.n3203 gnd.n3202 53.0052
R15241 gnd.n3205 gnd.n3204 53.0052
R15242 gnd.n3208 gnd.n3207 53.0052
R15243 gnd.n3210 gnd.n3209 53.0052
R15244 gnd.n3212 gnd.n3211 53.0052
R15245 gnd.n3214 gnd.n3213 53.0052
R15246 gnd.n3216 gnd.n3215 53.0052
R15247 gnd.n3220 gnd.n3219 53.0052
R15248 gnd.n3222 gnd.n3221 53.0052
R15249 gnd.n3224 gnd.n3223 53.0052
R15250 gnd.n3226 gnd.n3225 53.0052
R15251 gnd.n3228 gnd.n3227 53.0052
R15252 gnd.n60 gnd.n59 53.0052
R15253 gnd.n58 gnd.n57 53.0052
R15254 gnd.n56 gnd.n55 53.0052
R15255 gnd.n54 gnd.n53 53.0052
R15256 gnd.n52 gnd.n51 53.0052
R15257 gnd.n25 gnd.n24 53.0052
R15258 gnd.n23 gnd.n22 53.0052
R15259 gnd.n21 gnd.n20 53.0052
R15260 gnd.n19 gnd.n18 53.0052
R15261 gnd.n17 gnd.n16 53.0052
R15262 gnd.n36 gnd.n35 53.0052
R15263 gnd.n34 gnd.n33 53.0052
R15264 gnd.n32 gnd.n31 53.0052
R15265 gnd.n30 gnd.n29 53.0052
R15266 gnd.n28 gnd.n27 53.0052
R15267 gnd.n48 gnd.n47 53.0052
R15268 gnd.n46 gnd.n45 53.0052
R15269 gnd.n44 gnd.n43 53.0052
R15270 gnd.n42 gnd.n41 53.0052
R15271 gnd.n40 gnd.n39 53.0052
R15272 gnd.n6196 gnd.n6195 52.4801
R15273 gnd.n4207 gnd.t168 52.3082
R15274 gnd.n4175 gnd.t312 52.3082
R15275 gnd.n4143 gnd.t320 52.3082
R15276 gnd.n4112 gnd.t166 52.3082
R15277 gnd.n4080 gnd.t322 52.3082
R15278 gnd.n4048 gnd.t164 52.3082
R15279 gnd.n4016 gnd.t8 52.3082
R15280 gnd.n3985 gnd.t162 52.3082
R15281 gnd.n4037 gnd.n4005 51.4173
R15282 gnd.n4101 gnd.n4100 50.455
R15283 gnd.n4069 gnd.n4068 50.455
R15284 gnd.n4037 gnd.n4036 50.455
R15285 gnd.n3520 gnd.n3519 45.1884
R15286 gnd.n3111 gnd.n3110 45.1884
R15287 gnd.n6279 gnd.n6211 44.3322
R15288 gnd.n1019 gnd.n1018 44.3189
R15289 gnd.n2747 gnd.n1680 43.8514
R15290 gnd.n2748 gnd.n2747 43.8514
R15291 gnd.n2749 gnd.n2748 43.8514
R15292 gnd.n2749 gnd.n1674 43.8514
R15293 gnd.n2757 gnd.n1674 43.8514
R15294 gnd.n2758 gnd.n2757 43.8514
R15295 gnd.n2759 gnd.n2758 43.8514
R15296 gnd.n2759 gnd.n1668 43.8514
R15297 gnd.n2767 gnd.n1668 43.8514
R15298 gnd.n2768 gnd.n2767 43.8514
R15299 gnd.n2769 gnd.n2768 43.8514
R15300 gnd.n2769 gnd.n1662 43.8514
R15301 gnd.n2777 gnd.n1662 43.8514
R15302 gnd.n2778 gnd.n2777 43.8514
R15303 gnd.n2779 gnd.n2778 43.8514
R15304 gnd.n2779 gnd.n1656 43.8514
R15305 gnd.n2787 gnd.n1656 43.8514
R15306 gnd.n2788 gnd.n2787 43.8514
R15307 gnd.n2789 gnd.n2788 43.8514
R15308 gnd.n2789 gnd.n1650 43.8514
R15309 gnd.n2797 gnd.n1650 43.8514
R15310 gnd.n2798 gnd.n2797 43.8514
R15311 gnd.n2799 gnd.n2798 43.8514
R15312 gnd.n2799 gnd.n1644 43.8514
R15313 gnd.n2807 gnd.n1644 43.8514
R15314 gnd.n2808 gnd.n2807 43.8514
R15315 gnd.n2809 gnd.n2808 43.8514
R15316 gnd.n2809 gnd.n1638 43.8514
R15317 gnd.n2817 gnd.n1638 43.8514
R15318 gnd.n2818 gnd.n2817 43.8514
R15319 gnd.n2819 gnd.n2818 43.8514
R15320 gnd.n2819 gnd.n1632 43.8514
R15321 gnd.n2827 gnd.n1632 43.8514
R15322 gnd.n2828 gnd.n2827 43.8514
R15323 gnd.n2829 gnd.n2828 43.8514
R15324 gnd.n2829 gnd.n1626 43.8514
R15325 gnd.n2837 gnd.n1626 43.8514
R15326 gnd.n2838 gnd.n2837 43.8514
R15327 gnd.n2839 gnd.n2838 43.8514
R15328 gnd.n2839 gnd.n1620 43.8514
R15329 gnd.n2847 gnd.n1620 43.8514
R15330 gnd.n2848 gnd.n2847 43.8514
R15331 gnd.n2849 gnd.n2848 43.8514
R15332 gnd.n2849 gnd.n1614 43.8514
R15333 gnd.n2857 gnd.n1614 43.8514
R15334 gnd.n2858 gnd.n2857 43.8514
R15335 gnd.n2859 gnd.n2858 43.8514
R15336 gnd.n2859 gnd.n1608 43.8514
R15337 gnd.n2867 gnd.n1608 43.8514
R15338 gnd.n2868 gnd.n2867 43.8514
R15339 gnd.n2869 gnd.n2868 43.8514
R15340 gnd.n2869 gnd.n1602 43.8514
R15341 gnd.n2877 gnd.n1602 43.8514
R15342 gnd.n2878 gnd.n2877 43.8514
R15343 gnd.n2879 gnd.n2878 43.8514
R15344 gnd.n2879 gnd.n1596 43.8514
R15345 gnd.n2887 gnd.n1596 43.8514
R15346 gnd.n2888 gnd.n2887 43.8514
R15347 gnd.n2889 gnd.n2888 43.8514
R15348 gnd.n2889 gnd.n1590 43.8514
R15349 gnd.n2897 gnd.n1590 43.8514
R15350 gnd.n2898 gnd.n2897 43.8514
R15351 gnd.n2899 gnd.n2898 43.8514
R15352 gnd.n2899 gnd.n1584 43.8514
R15353 gnd.n2907 gnd.n1584 43.8514
R15354 gnd.n2908 gnd.n2907 43.8514
R15355 gnd.n2909 gnd.n2908 43.8514
R15356 gnd.n2909 gnd.n1578 43.8514
R15357 gnd.n2917 gnd.n1578 43.8514
R15358 gnd.n2918 gnd.n2917 43.8514
R15359 gnd.n2919 gnd.n2918 43.8514
R15360 gnd.n2919 gnd.n1572 43.8514
R15361 gnd.n2927 gnd.n1572 43.8514
R15362 gnd.n2928 gnd.n2927 43.8514
R15363 gnd.n2929 gnd.n2928 43.8514
R15364 gnd.n2929 gnd.n1566 43.8514
R15365 gnd.n2937 gnd.n1566 43.8514
R15366 gnd.n2938 gnd.n2937 43.8514
R15367 gnd.n2939 gnd.n2938 43.8514
R15368 gnd.n2939 gnd.n1560 43.8514
R15369 gnd.n2948 gnd.n1560 43.8514
R15370 gnd.n2949 gnd.n2948 43.8514
R15371 gnd.n4413 gnd.n2949 43.8514
R15372 gnd.n5265 gnd.n5264 42.2793
R15373 gnd.n6698 gnd.n6697 42.2793
R15374 gnd.n3521 gnd.n3520 42.2793
R15375 gnd.n3112 gnd.n3111 42.2793
R15376 gnd.n3447 gnd.n3446 42.2793
R15377 gnd.n3068 gnd.n3067 42.2793
R15378 gnd.n5260 gnd.n5255 42.2793
R15379 gnd.n6657 gnd.n516 42.2793
R15380 gnd.n6620 gnd.n539 42.2793
R15381 gnd.n6580 gnd.n562 42.2793
R15382 gnd.n7136 gnd.n7133 42.2793
R15383 gnd.n7178 gnd.n7112 42.2793
R15384 gnd.n7220 gnd.n7219 42.2793
R15385 gnd.n182 gnd.n181 42.2793
R15386 gnd.n4671 gnd.n4471 42.2793
R15387 gnd.n4631 gnd.n4493 42.2793
R15388 gnd.n4591 gnd.n4515 42.2793
R15389 gnd.n4544 gnd.n4543 42.2793
R15390 gnd.n5394 gnd.n5393 42.2793
R15391 gnd.n1204 gnd.n1203 42.2793
R15392 gnd.n5504 gnd.n1170 42.2793
R15393 gnd.n448 gnd.n447 42.2793
R15394 gnd.n4703 gnd.n4452 42.0631
R15395 gnd.n7253 gnd.n171 42.0631
R15396 gnd.n1017 gnd.n1016 41.6274
R15397 gnd.n6206 gnd.n6205 41.6274
R15398 gnd.n1026 gnd.n1025 40.8975
R15399 gnd.n6209 gnd.n6208 40.8975
R15400 gnd.n1025 gnd.n1024 35.055
R15401 gnd.n1020 gnd.n1019 35.055
R15402 gnd.n6198 gnd.n6197 35.055
R15403 gnd.n6208 gnd.n6194 35.055
R15404 gnd.n3583 gnd.n3477 31.8661
R15405 gnd.n3583 gnd.n3582 31.8661
R15406 gnd.n3591 gnd.n3466 31.8661
R15407 gnd.n3599 gnd.n3466 31.8661
R15408 gnd.n3599 gnd.n3460 31.8661
R15409 gnd.n3607 gnd.n3460 31.8661
R15410 gnd.n3607 gnd.n3453 31.8661
R15411 gnd.n3645 gnd.n3453 31.8661
R15412 gnd.n3655 gnd.n3386 31.8661
R15413 gnd.n5189 gnd.n1273 31.8661
R15414 gnd.n5183 gnd.n5182 31.8661
R15415 gnd.n5182 gnd.n1245 31.8661
R15416 gnd.n5175 gnd.n1259 31.8661
R15417 gnd.n6462 gnd.n427 31.8661
R15418 gnd.n6455 gnd.n442 31.8661
R15419 gnd.n6455 gnd.n457 31.8661
R15420 gnd.n6716 gnd.n418 31.8661
R15421 gnd.n6285 gnd.n692 31.0639
R15422 gnd.n5592 gnd.n5591 31.0639
R15423 gnd.n4413 gnd.n4412 26.311
R15424 gnd.n5264 gnd.n5263 25.7944
R15425 gnd.n6697 gnd.n6696 25.7944
R15426 gnd.n3446 gnd.n3445 25.7944
R15427 gnd.n3067 gnd.n3066 25.7944
R15428 gnd.n5255 gnd.n5254 25.7944
R15429 gnd.n516 gnd.n515 25.7944
R15430 gnd.n539 gnd.n538 25.7944
R15431 gnd.n562 gnd.n561 25.7944
R15432 gnd.n7133 gnd.n7132 25.7944
R15433 gnd.n7112 gnd.n7111 25.7944
R15434 gnd.n7219 gnd.n7218 25.7944
R15435 gnd.n181 gnd.n180 25.7944
R15436 gnd.n4471 gnd.n4470 25.7944
R15437 gnd.n4493 gnd.n4492 25.7944
R15438 gnd.n4515 gnd.n4514 25.7944
R15439 gnd.n4543 gnd.n4542 25.7944
R15440 gnd.n5393 gnd.n5392 25.7944
R15441 gnd.n1203 gnd.n1202 25.7944
R15442 gnd.n1170 gnd.n1169 25.7944
R15443 gnd.n447 gnd.n446 25.7944
R15444 gnd.n3667 gnd.n3387 24.8557
R15445 gnd.n3677 gnd.n3370 24.8557
R15446 gnd.n3373 gnd.n3361 24.8557
R15447 gnd.n3698 gnd.n3362 24.8557
R15448 gnd.n3708 gnd.n3342 24.8557
R15449 gnd.n3718 gnd.n3717 24.8557
R15450 gnd.n3328 gnd.n3326 24.8557
R15451 gnd.n3749 gnd.n3748 24.8557
R15452 gnd.n3764 gnd.n3311 24.8557
R15453 gnd.n3818 gnd.n3250 24.8557
R15454 gnd.n3774 gnd.n3251 24.8557
R15455 gnd.n3811 gnd.n3262 24.8557
R15456 gnd.n3300 gnd.n3299 24.8557
R15457 gnd.n3805 gnd.n3804 24.8557
R15458 gnd.n3286 gnd.n3273 24.8557
R15459 gnd.n3844 gnd.n3843 24.8557
R15460 gnd.n3854 gnd.n3182 24.8557
R15461 gnd.n3866 gnd.n3174 24.8557
R15462 gnd.n3865 gnd.n3162 24.8557
R15463 gnd.n3884 gnd.n3883 24.8557
R15464 gnd.n3894 gnd.n3155 24.8557
R15465 gnd.n3907 gnd.n3143 24.8557
R15466 gnd.n3940 gnd.n3939 24.8557
R15467 gnd.n3949 gnd.n3130 24.8557
R15468 gnd.n4405 gnd.n2960 24.8557
R15469 gnd.n3929 gnd.n2971 24.8557
R15470 gnd.n4398 gnd.n4397 24.8557
R15471 gnd.n4391 gnd.n2983 24.8557
R15472 gnd.n4254 gnd.n2996 24.8557
R15473 gnd.n4384 gnd.n4383 24.8557
R15474 gnd.n4377 gnd.n3008 24.8557
R15475 gnd.n4376 gnd.n3011 24.8557
R15476 gnd.n4243 gnd.n3022 24.8557
R15477 gnd.n4363 gnd.n3033 24.8557
R15478 gnd.n3688 gnd.t161 23.2624
R15479 gnd.n3389 gnd.t60 22.6251
R15480 gnd.t165 gnd.n3394 21.3504
R15481 gnd.n4584 gnd.n4452 21.0318
R15482 gnd.n4714 gnd.n1506 21.0318
R15483 gnd.n4728 gnd.n1500 21.0318
R15484 gnd.n4739 gnd.n1489 21.0318
R15485 gnd.n4722 gnd.n1492 21.0318
R15486 gnd.n4747 gnd.n1481 21.0318
R15487 gnd.n4766 gnd.n1467 21.0318
R15488 gnd.n4759 gnd.n1470 21.0318
R15489 gnd.n4774 gnd.n1460 21.0318
R15490 gnd.n4799 gnd.n1449 21.0318
R15491 gnd.n4793 gnd.n1434 21.0318
R15492 gnd.n4812 gnd.n1442 21.0318
R15493 gnd.n1423 gnd.n1415 21.0318
R15494 gnd.n4854 gnd.n4853 21.0318
R15495 gnd.n4920 gnd.n1358 21.0318
R15496 gnd.n4864 gnd.n1361 21.0318
R15497 gnd.n4909 gnd.n1372 21.0318
R15498 gnd.n4908 gnd.n1378 21.0318
R15499 gnd.n1385 gnd.n1384 21.0318
R15500 gnd.n4901 gnd.n4900 21.0318
R15501 gnd.n4881 gnd.n1400 21.0318
R15502 gnd.n4931 gnd.n1342 21.0318
R15503 gnd.n4941 gnd.n4940 21.0318
R15504 gnd.n4974 gnd.n1319 21.0318
R15505 gnd.n4961 gnd.n4960 21.0318
R15506 gnd.n4984 gnd.n1309 21.0318
R15507 gnd.n4996 gnd.n1302 21.0318
R15508 gnd.n5008 gnd.n1291 21.0318
R15509 gnd.n5017 gnd.n5016 21.0318
R15510 gnd.n5346 gnd.n1232 21.0318
R15511 gnd.n5356 gnd.n1222 21.0318
R15512 gnd.n5026 gnd.n1225 21.0318
R15513 gnd.n5190 gnd.n1214 21.0318
R15514 gnd.n6715 gnd.n392 21.0318
R15515 gnd.n6727 gnd.n382 21.0318
R15516 gnd.n6744 gnd.n384 21.0318
R15517 gnd.n6754 gnd.n374 21.0318
R15518 gnd.n6753 gnd.n359 21.0318
R15519 gnd.n6790 gnd.n349 21.0318
R15520 gnd.n6813 gnd.n351 21.0318
R15521 gnd.n6822 gnd.n330 21.0318
R15522 gnd.n6838 gnd.n333 21.0318
R15523 gnd.n6826 gnd.n320 21.0318
R15524 gnd.n6849 gnd.n322 21.0318
R15525 gnd.n6865 gnd.n306 21.0318
R15526 gnd.n6872 gnd.n302 21.0318
R15527 gnd.n6885 gnd.n288 21.0318
R15528 gnd.n6902 gnd.n6901 21.0318
R15529 gnd.n6912 gnd.n286 21.0318
R15530 gnd.n6907 gnd.n278 21.0318
R15531 gnd.n7325 gnd.n71 21.0318
R15532 gnd.n6998 gnd.n265 21.0318
R15533 gnd.n6997 gnd.n86 21.0318
R15534 gnd.n7317 gnd.n89 21.0318
R15535 gnd.n7311 gnd.n101 21.0318
R15536 gnd.n6985 gnd.n108 21.0318
R15537 gnd.n6979 gnd.n117 21.0318
R15538 gnd.n7299 gnd.n120 21.0318
R15539 gnd.n6973 gnd.n128 21.0318
R15540 gnd.n7293 gnd.n131 21.0318
R15541 gnd.n7287 gnd.n141 21.0318
R15542 gnd.n6961 gnd.n149 21.0318
R15543 gnd.n7281 gnd.n152 21.0318
R15544 gnd.n6955 gnd.n159 21.0318
R15545 gnd.n7262 gnd.n168 21.0318
R15546 gnd.n7269 gnd.n171 21.0318
R15547 gnd.n3922 gnd.t300 20.7131
R15548 gnd.n4827 gnd.t229 20.7131
R15549 gnd.t190 gnd.n1388 20.7131
R15550 gnd.n6886 gnd.t174 20.7131
R15551 gnd.n6991 gnd.t205 20.7131
R15552 gnd.n1273 gnd.n1156 20.3945
R15553 gnd.n6693 gnd.n418 20.3945
R15554 gnd.t302 gnd.n3136 20.0758
R15555 gnd.n4750 gnd.t181 20.0758
R15556 gnd.t195 gnd.n1311 20.0758
R15557 gnd.t170 gnd.n342 20.0758
R15558 gnd.n6967 gnd.t216 20.0758
R15559 gnd.n1014 gnd.t69 19.8005
R15560 gnd.n1014 gnd.t108 19.8005
R15561 gnd.n1013 gnd.t87 19.8005
R15562 gnd.n1013 gnd.t18 19.8005
R15563 gnd.n6203 gnd.t106 19.8005
R15564 gnd.n6203 gnd.t58 19.8005
R15565 gnd.n6202 gnd.t131 19.8005
R15566 gnd.n6202 gnd.t21 19.8005
R15567 gnd.n1010 gnd.n1009 19.5087
R15568 gnd.n1023 gnd.n1010 19.5087
R15569 gnd.n1021 gnd.n1012 19.5087
R15570 gnd.n6207 gnd.n6201 19.5087
R15571 gnd.n3855 gnd.t290 19.4385
R15572 gnd.n5089 gnd.n5088 19.3944
R15573 gnd.n5093 gnd.n5088 19.3944
R15574 gnd.n5093 gnd.n5085 19.3944
R15575 gnd.n5111 gnd.n5085 19.3944
R15576 gnd.n5111 gnd.n5083 19.3944
R15577 gnd.n5115 gnd.n5083 19.3944
R15578 gnd.n5115 gnd.n5073 19.3944
R15579 gnd.n5132 gnd.n5073 19.3944
R15580 gnd.n5132 gnd.n5070 19.3944
R15581 gnd.n5137 gnd.n5070 19.3944
R15582 gnd.n5137 gnd.n5071 19.3944
R15583 gnd.n5071 gnd.n1081 19.3944
R15584 gnd.n5616 gnd.n1081 19.3944
R15585 gnd.n5616 gnd.n1082 19.3944
R15586 gnd.n5612 gnd.n1082 19.3944
R15587 gnd.n5612 gnd.n5611 19.3944
R15588 gnd.n5611 gnd.n5610 19.3944
R15589 gnd.n5610 gnd.n5600 19.3944
R15590 gnd.n5606 gnd.n5600 19.3944
R15591 gnd.n5606 gnd.n5605 19.3944
R15592 gnd.n5605 gnd.n5604 19.3944
R15593 gnd.n5604 gnd.n956 19.3944
R15594 gnd.n5725 gnd.n956 19.3944
R15595 gnd.n5725 gnd.n953 19.3944
R15596 gnd.n5729 gnd.n953 19.3944
R15597 gnd.n5730 gnd.n5729 19.3944
R15598 gnd.n5732 gnd.n5730 19.3944
R15599 gnd.n5732 gnd.n950 19.3944
R15600 gnd.n5737 gnd.n950 19.3944
R15601 gnd.n5737 gnd.n951 19.3944
R15602 gnd.n951 gnd.n891 19.3944
R15603 gnd.n5808 gnd.n891 19.3944
R15604 gnd.n5808 gnd.n888 19.3944
R15605 gnd.n5840 gnd.n888 19.3944
R15606 gnd.n5840 gnd.n889 19.3944
R15607 gnd.n5836 gnd.n889 19.3944
R15608 gnd.n5836 gnd.n5835 19.3944
R15609 gnd.n5835 gnd.n5834 19.3944
R15610 gnd.n5834 gnd.n5821 19.3944
R15611 gnd.n5830 gnd.n5821 19.3944
R15612 gnd.n5830 gnd.n5829 19.3944
R15613 gnd.n5829 gnd.n5828 19.3944
R15614 gnd.n5828 gnd.n5824 19.3944
R15615 gnd.n5824 gnd.n811 19.3944
R15616 gnd.n5954 gnd.n811 19.3944
R15617 gnd.n5955 gnd.n5954 19.3944
R15618 gnd.n5955 gnd.n808 19.3944
R15619 gnd.n6048 gnd.n808 19.3944
R15620 gnd.n6048 gnd.n809 19.3944
R15621 gnd.n6044 gnd.n809 19.3944
R15622 gnd.n6044 gnd.n6043 19.3944
R15623 gnd.n6043 gnd.n6042 19.3944
R15624 gnd.n6042 gnd.n5960 19.3944
R15625 gnd.n6038 gnd.n5960 19.3944
R15626 gnd.n6038 gnd.n6037 19.3944
R15627 gnd.n6037 gnd.n6036 19.3944
R15628 gnd.n6036 gnd.n5965 19.3944
R15629 gnd.n6032 gnd.n5965 19.3944
R15630 gnd.n6032 gnd.n6031 19.3944
R15631 gnd.n6031 gnd.n6030 19.3944
R15632 gnd.n6030 gnd.n6012 19.3944
R15633 gnd.n6026 gnd.n6012 19.3944
R15634 gnd.n6026 gnd.n6025 19.3944
R15635 gnd.n6025 gnd.n6024 19.3944
R15636 gnd.n6024 gnd.n6017 19.3944
R15637 gnd.n6020 gnd.n6017 19.3944
R15638 gnd.n6020 gnd.n6019 19.3944
R15639 gnd.n6019 gnd.n634 19.3944
R15640 gnd.n6374 gnd.n634 19.3944
R15641 gnd.n6374 gnd.n631 19.3944
R15642 gnd.n6379 gnd.n631 19.3944
R15643 gnd.n6379 gnd.n632 19.3944
R15644 gnd.n632 gnd.n609 19.3944
R15645 gnd.n6404 gnd.n609 19.3944
R15646 gnd.n6404 gnd.n606 19.3944
R15647 gnd.n6409 gnd.n606 19.3944
R15648 gnd.n6409 gnd.n607 19.3944
R15649 gnd.n607 gnd.n583 19.3944
R15650 gnd.n6434 gnd.n583 19.3944
R15651 gnd.n6434 gnd.n580 19.3944
R15652 gnd.n6439 gnd.n580 19.3944
R15653 gnd.n6439 gnd.n581 19.3944
R15654 gnd.n5268 gnd.n1242 19.3944
R15655 gnd.n5334 gnd.n1242 19.3944
R15656 gnd.n5334 gnd.n5333 19.3944
R15657 gnd.n5327 gnd.n5326 19.3944
R15658 gnd.n5326 gnd.n1264 19.3944
R15659 gnd.n5322 gnd.n1264 19.3944
R15660 gnd.n5322 gnd.n5321 19.3944
R15661 gnd.n5321 gnd.n5320 19.3944
R15662 gnd.n5320 gnd.n5317 19.3944
R15663 gnd.n5317 gnd.n5316 19.3944
R15664 gnd.n5316 gnd.n1271 19.3944
R15665 gnd.n5198 gnd.n1271 19.3944
R15666 gnd.n5308 gnd.n5198 19.3944
R15667 gnd.n5308 gnd.n5307 19.3944
R15668 gnd.n5307 gnd.n5201 19.3944
R15669 gnd.n5300 gnd.n5201 19.3944
R15670 gnd.n5300 gnd.n5299 19.3944
R15671 gnd.n5299 gnd.n5214 19.3944
R15672 gnd.n5292 gnd.n5214 19.3944
R15673 gnd.n5292 gnd.n5291 19.3944
R15674 gnd.n5291 gnd.n5224 19.3944
R15675 gnd.n5284 gnd.n5224 19.3944
R15676 gnd.n5284 gnd.n5283 19.3944
R15677 gnd.n5283 gnd.n5237 19.3944
R15678 gnd.n5276 gnd.n5237 19.3944
R15679 gnd.n5276 gnd.n5275 19.3944
R15680 gnd.n5275 gnd.n5247 19.3944
R15681 gnd.n6569 gnd.n6491 19.3944
R15682 gnd.n6569 gnd.n6568 19.3944
R15683 gnd.n6568 gnd.n6494 19.3944
R15684 gnd.n6561 gnd.n6494 19.3944
R15685 gnd.n6561 gnd.n6560 19.3944
R15686 gnd.n6560 gnd.n6504 19.3944
R15687 gnd.n6553 gnd.n6504 19.3944
R15688 gnd.n6553 gnd.n6552 19.3944
R15689 gnd.n6552 gnd.n6514 19.3944
R15690 gnd.n6545 gnd.n6514 19.3944
R15691 gnd.n6545 gnd.n6544 19.3944
R15692 gnd.n6544 gnd.n6524 19.3944
R15693 gnd.n6537 gnd.n6524 19.3944
R15694 gnd.n6537 gnd.n6536 19.3944
R15695 gnd.n6536 gnd.n452 19.3944
R15696 gnd.n6699 gnd.n452 19.3944
R15697 gnd.n3570 gnd.n3569 19.3944
R15698 gnd.n3569 gnd.n3568 19.3944
R15699 gnd.n3568 gnd.n3567 19.3944
R15700 gnd.n3567 gnd.n3565 19.3944
R15701 gnd.n3565 gnd.n3562 19.3944
R15702 gnd.n3562 gnd.n3561 19.3944
R15703 gnd.n3561 gnd.n3558 19.3944
R15704 gnd.n3558 gnd.n3557 19.3944
R15705 gnd.n3557 gnd.n3554 19.3944
R15706 gnd.n3554 gnd.n3553 19.3944
R15707 gnd.n3553 gnd.n3550 19.3944
R15708 gnd.n3550 gnd.n3549 19.3944
R15709 gnd.n3549 gnd.n3546 19.3944
R15710 gnd.n3546 gnd.n3545 19.3944
R15711 gnd.n3545 gnd.n3542 19.3944
R15712 gnd.n3542 gnd.n3541 19.3944
R15713 gnd.n3541 gnd.n3538 19.3944
R15714 gnd.n3538 gnd.n3537 19.3944
R15715 gnd.n3537 gnd.n3534 19.3944
R15716 gnd.n3534 gnd.n3533 19.3944
R15717 gnd.n3533 gnd.n3530 19.3944
R15718 gnd.n3530 gnd.n3529 19.3944
R15719 gnd.n3526 gnd.n3525 19.3944
R15720 gnd.n3525 gnd.n3481 19.3944
R15721 gnd.n3576 gnd.n3481 19.3944
R15722 gnd.n4283 gnd.n3114 19.3944
R15723 gnd.n4283 gnd.n4282 19.3944
R15724 gnd.n4282 gnd.n4281 19.3944
R15725 gnd.n4325 gnd.n4324 19.3944
R15726 gnd.n4324 gnd.n4323 19.3944
R15727 gnd.n4323 gnd.n3075 19.3944
R15728 gnd.n4318 gnd.n3075 19.3944
R15729 gnd.n4318 gnd.n4317 19.3944
R15730 gnd.n4317 gnd.n4316 19.3944
R15731 gnd.n4316 gnd.n3082 19.3944
R15732 gnd.n4311 gnd.n3082 19.3944
R15733 gnd.n4311 gnd.n4310 19.3944
R15734 gnd.n4310 gnd.n4309 19.3944
R15735 gnd.n4309 gnd.n3089 19.3944
R15736 gnd.n4304 gnd.n3089 19.3944
R15737 gnd.n4304 gnd.n4303 19.3944
R15738 gnd.n4303 gnd.n4302 19.3944
R15739 gnd.n4302 gnd.n3096 19.3944
R15740 gnd.n4297 gnd.n3096 19.3944
R15741 gnd.n4297 gnd.n4296 19.3944
R15742 gnd.n4296 gnd.n4295 19.3944
R15743 gnd.n4295 gnd.n3103 19.3944
R15744 gnd.n4290 gnd.n3103 19.3944
R15745 gnd.n4290 gnd.n4289 19.3944
R15746 gnd.n4289 gnd.n4288 19.3944
R15747 gnd.n3669 gnd.n3378 19.3944
R15748 gnd.n3679 gnd.n3378 19.3944
R15749 gnd.n3680 gnd.n3679 19.3944
R15750 gnd.n3680 gnd.n3359 19.3944
R15751 gnd.n3700 gnd.n3359 19.3944
R15752 gnd.n3700 gnd.n3351 19.3944
R15753 gnd.n3710 gnd.n3351 19.3944
R15754 gnd.n3711 gnd.n3710 19.3944
R15755 gnd.n3712 gnd.n3711 19.3944
R15756 gnd.n3712 gnd.n3334 19.3944
R15757 gnd.n3729 gnd.n3334 19.3944
R15758 gnd.n3732 gnd.n3729 19.3944
R15759 gnd.n3732 gnd.n3731 19.3944
R15760 gnd.n3731 gnd.n3307 19.3944
R15761 gnd.n3771 gnd.n3307 19.3944
R15762 gnd.n3771 gnd.n3304 19.3944
R15763 gnd.n3777 gnd.n3304 19.3944
R15764 gnd.n3778 gnd.n3777 19.3944
R15765 gnd.n3778 gnd.n3302 19.3944
R15766 gnd.n3784 gnd.n3302 19.3944
R15767 gnd.n3787 gnd.n3784 19.3944
R15768 gnd.n3789 gnd.n3787 19.3944
R15769 gnd.n3795 gnd.n3789 19.3944
R15770 gnd.n3795 gnd.n3794 19.3944
R15771 gnd.n3794 gnd.n3177 19.3944
R15772 gnd.n3861 gnd.n3177 19.3944
R15773 gnd.n3862 gnd.n3861 19.3944
R15774 gnd.n3862 gnd.n3170 19.3944
R15775 gnd.n3873 gnd.n3170 19.3944
R15776 gnd.n3874 gnd.n3873 19.3944
R15777 gnd.n3874 gnd.n3153 19.3944
R15778 gnd.n3153 gnd.n3151 19.3944
R15779 gnd.n3898 gnd.n3151 19.3944
R15780 gnd.n3901 gnd.n3898 19.3944
R15781 gnd.n3901 gnd.n3900 19.3944
R15782 gnd.n3900 gnd.n3127 19.3944
R15783 gnd.n3952 gnd.n3127 19.3944
R15784 gnd.n3953 gnd.n3952 19.3944
R15785 gnd.n3953 gnd.n3125 19.3944
R15786 gnd.n3959 gnd.n3125 19.3944
R15787 gnd.n3961 gnd.n3959 19.3944
R15788 gnd.n3965 gnd.n3961 19.3944
R15789 gnd.n3966 gnd.n3965 19.3944
R15790 gnd.n4252 gnd.n3966 19.3944
R15791 gnd.n4252 gnd.n4251 19.3944
R15792 gnd.n4251 gnd.n4250 19.3944
R15793 gnd.n4250 gnd.n4247 19.3944
R15794 gnd.n4247 gnd.n4246 19.3944
R15795 gnd.n4246 gnd.n4245 19.3944
R15796 gnd.n4245 gnd.n4242 19.3944
R15797 gnd.n4242 gnd.n4241 19.3944
R15798 gnd.n4241 gnd.n4238 19.3944
R15799 gnd.n4238 gnd.n4237 19.3944
R15800 gnd.n3660 gnd.n3659 19.3944
R15801 gnd.n3659 gnd.n3392 19.3944
R15802 gnd.n3415 gnd.n3392 19.3944
R15803 gnd.n3418 gnd.n3415 19.3944
R15804 gnd.n3418 gnd.n3411 19.3944
R15805 gnd.n3422 gnd.n3411 19.3944
R15806 gnd.n3425 gnd.n3422 19.3944
R15807 gnd.n3428 gnd.n3425 19.3944
R15808 gnd.n3428 gnd.n3409 19.3944
R15809 gnd.n3432 gnd.n3409 19.3944
R15810 gnd.n3435 gnd.n3432 19.3944
R15811 gnd.n3438 gnd.n3435 19.3944
R15812 gnd.n3438 gnd.n3407 19.3944
R15813 gnd.n3442 gnd.n3407 19.3944
R15814 gnd.n3665 gnd.n3664 19.3944
R15815 gnd.n3664 gnd.n3368 19.3944
R15816 gnd.n3690 gnd.n3368 19.3944
R15817 gnd.n3690 gnd.n3366 19.3944
R15818 gnd.n3696 gnd.n3366 19.3944
R15819 gnd.n3696 gnd.n3695 19.3944
R15820 gnd.n3695 gnd.n3340 19.3944
R15821 gnd.n3720 gnd.n3340 19.3944
R15822 gnd.n3720 gnd.n3338 19.3944
R15823 gnd.n3724 gnd.n3338 19.3944
R15824 gnd.n3724 gnd.n3318 19.3944
R15825 gnd.n3751 gnd.n3318 19.3944
R15826 gnd.n3751 gnd.n3316 19.3944
R15827 gnd.n3761 gnd.n3316 19.3944
R15828 gnd.n3761 gnd.n3760 19.3944
R15829 gnd.n3760 gnd.n3759 19.3944
R15830 gnd.n3759 gnd.n3265 19.3944
R15831 gnd.n3809 gnd.n3265 19.3944
R15832 gnd.n3809 gnd.n3808 19.3944
R15833 gnd.n3808 gnd.n3807 19.3944
R15834 gnd.n3807 gnd.n3269 19.3944
R15835 gnd.n3289 gnd.n3269 19.3944
R15836 gnd.n3289 gnd.n3187 19.3944
R15837 gnd.n3846 gnd.n3187 19.3944
R15838 gnd.n3846 gnd.n3185 19.3944
R15839 gnd.n3852 gnd.n3185 19.3944
R15840 gnd.n3852 gnd.n3851 19.3944
R15841 gnd.n3851 gnd.n3160 19.3944
R15842 gnd.n3886 gnd.n3160 19.3944
R15843 gnd.n3886 gnd.n3158 19.3944
R15844 gnd.n3892 gnd.n3158 19.3944
R15845 gnd.n3892 gnd.n3891 19.3944
R15846 gnd.n3891 gnd.n3134 19.3944
R15847 gnd.n3942 gnd.n3134 19.3944
R15848 gnd.n3942 gnd.n3132 19.3944
R15849 gnd.n3947 gnd.n3132 19.3944
R15850 gnd.n3947 gnd.n2965 19.3944
R15851 gnd.n4402 gnd.n2965 19.3944
R15852 gnd.n4402 gnd.n4401 19.3944
R15853 gnd.n4401 gnd.n4400 19.3944
R15854 gnd.n4400 gnd.n2969 19.3944
R15855 gnd.n2988 gnd.n2969 19.3944
R15856 gnd.n4388 gnd.n2988 19.3944
R15857 gnd.n4388 gnd.n4387 19.3944
R15858 gnd.n4387 gnd.n4386 19.3944
R15859 gnd.n4386 gnd.n2994 19.3944
R15860 gnd.n3014 gnd.n2994 19.3944
R15861 gnd.n4374 gnd.n3014 19.3944
R15862 gnd.n4374 gnd.n4373 19.3944
R15863 gnd.n4373 gnd.n4372 19.3944
R15864 gnd.n4372 gnd.n3020 19.3944
R15865 gnd.n3039 gnd.n3020 19.3944
R15866 gnd.n4360 gnd.n3039 19.3944
R15867 gnd.n4357 gnd.n4356 19.3944
R15868 gnd.n4356 gnd.n4355 19.3944
R15869 gnd.n4355 gnd.n3045 19.3944
R15870 gnd.n4350 gnd.n3045 19.3944
R15871 gnd.n4350 gnd.n4349 19.3944
R15872 gnd.n4349 gnd.n4348 19.3944
R15873 gnd.n4348 gnd.n3052 19.3944
R15874 gnd.n4343 gnd.n3052 19.3944
R15875 gnd.n4343 gnd.n4342 19.3944
R15876 gnd.n4342 gnd.n4341 19.3944
R15877 gnd.n4341 gnd.n3059 19.3944
R15878 gnd.n4336 gnd.n3059 19.3944
R15879 gnd.n4336 gnd.n4335 19.3944
R15880 gnd.n4335 gnd.n4334 19.3944
R15881 gnd.n3580 gnd.n3479 19.3944
R15882 gnd.n3580 gnd.n3470 19.3944
R15883 gnd.n3593 gnd.n3470 19.3944
R15884 gnd.n3593 gnd.n3468 19.3944
R15885 gnd.n3597 gnd.n3468 19.3944
R15886 gnd.n3597 gnd.n3458 19.3944
R15887 gnd.n3609 gnd.n3458 19.3944
R15888 gnd.n3609 gnd.n3456 19.3944
R15889 gnd.n3643 gnd.n3456 19.3944
R15890 gnd.n3643 gnd.n3642 19.3944
R15891 gnd.n3642 gnd.n3641 19.3944
R15892 gnd.n3641 gnd.n3640 19.3944
R15893 gnd.n3640 gnd.n3637 19.3944
R15894 gnd.n3637 gnd.n3636 19.3944
R15895 gnd.n3636 gnd.n3635 19.3944
R15896 gnd.n3635 gnd.n3633 19.3944
R15897 gnd.n3633 gnd.n3632 19.3944
R15898 gnd.n3632 gnd.n3629 19.3944
R15899 gnd.n3629 gnd.n3628 19.3944
R15900 gnd.n3628 gnd.n3627 19.3944
R15901 gnd.n3627 gnd.n3625 19.3944
R15902 gnd.n3625 gnd.n3324 19.3944
R15903 gnd.n3740 gnd.n3324 19.3944
R15904 gnd.n3740 gnd.n3322 19.3944
R15905 gnd.n3746 gnd.n3322 19.3944
R15906 gnd.n3746 gnd.n3745 19.3944
R15907 gnd.n3745 gnd.n3246 19.3944
R15908 gnd.n3820 gnd.n3246 19.3944
R15909 gnd.n3820 gnd.n3247 19.3944
R15910 gnd.n3294 gnd.n3293 19.3944
R15911 gnd.n3297 gnd.n3296 19.3944
R15912 gnd.n3284 gnd.n3283 19.3944
R15913 gnd.n3839 gnd.n3192 19.3944
R15914 gnd.n3839 gnd.n3838 19.3944
R15915 gnd.n3838 gnd.n3837 19.3944
R15916 gnd.n3837 gnd.n3835 19.3944
R15917 gnd.n3835 gnd.n3834 19.3944
R15918 gnd.n3834 gnd.n3832 19.3944
R15919 gnd.n3832 gnd.n3831 19.3944
R15920 gnd.n3831 gnd.n3141 19.3944
R15921 gnd.n3909 gnd.n3141 19.3944
R15922 gnd.n3909 gnd.n3139 19.3944
R15923 gnd.n3937 gnd.n3139 19.3944
R15924 gnd.n3937 gnd.n3936 19.3944
R15925 gnd.n3936 gnd.n3935 19.3944
R15926 gnd.n3935 gnd.n3933 19.3944
R15927 gnd.n3933 gnd.n3932 19.3944
R15928 gnd.n3932 gnd.n3926 19.3944
R15929 gnd.n3926 gnd.n3925 19.3944
R15930 gnd.n3925 gnd.n3924 19.3944
R15931 gnd.n3924 gnd.n3921 19.3944
R15932 gnd.n3921 gnd.n3124 19.3944
R15933 gnd.n4258 gnd.n3124 19.3944
R15934 gnd.n4258 gnd.n3122 19.3944
R15935 gnd.n4264 gnd.n3122 19.3944
R15936 gnd.n4265 gnd.n4264 19.3944
R15937 gnd.n4268 gnd.n4265 19.3944
R15938 gnd.n4268 gnd.n3120 19.3944
R15939 gnd.n4272 gnd.n3120 19.3944
R15940 gnd.n4275 gnd.n4272 19.3944
R15941 gnd.n4276 gnd.n4275 19.3944
R15942 gnd.n3585 gnd.n3475 19.3944
R15943 gnd.n3585 gnd.n3473 19.3944
R15944 gnd.n3589 gnd.n3473 19.3944
R15945 gnd.n3589 gnd.n3464 19.3944
R15946 gnd.n3601 gnd.n3464 19.3944
R15947 gnd.n3601 gnd.n3462 19.3944
R15948 gnd.n3605 gnd.n3462 19.3944
R15949 gnd.n3605 gnd.n3451 19.3944
R15950 gnd.n3647 gnd.n3451 19.3944
R15951 gnd.n3647 gnd.n3405 19.3944
R15952 gnd.n3653 gnd.n3405 19.3944
R15953 gnd.n3653 gnd.n3652 19.3944
R15954 gnd.n3652 gnd.n3383 19.3944
R15955 gnd.n3674 gnd.n3383 19.3944
R15956 gnd.n3674 gnd.n3376 19.3944
R15957 gnd.n3685 gnd.n3376 19.3944
R15958 gnd.n3685 gnd.n3684 19.3944
R15959 gnd.n3684 gnd.n3357 19.3944
R15960 gnd.n3705 gnd.n3357 19.3944
R15961 gnd.n3705 gnd.n3347 19.3944
R15962 gnd.n3715 gnd.n3347 19.3944
R15963 gnd.n3715 gnd.n3330 19.3944
R15964 gnd.n3736 gnd.n3330 19.3944
R15965 gnd.n3736 gnd.n3735 19.3944
R15966 gnd.n3735 gnd.n3309 19.3944
R15967 gnd.n3766 gnd.n3309 19.3944
R15968 gnd.n3766 gnd.n3254 19.3944
R15969 gnd.n3816 gnd.n3254 19.3944
R15970 gnd.n3816 gnd.n3815 19.3944
R15971 gnd.n3815 gnd.n3814 19.3944
R15972 gnd.n3814 gnd.n3258 19.3944
R15973 gnd.n3276 gnd.n3258 19.3944
R15974 gnd.n3802 gnd.n3276 19.3944
R15975 gnd.n3802 gnd.n3801 19.3944
R15976 gnd.n3801 gnd.n3800 19.3944
R15977 gnd.n3800 gnd.n3280 19.3944
R15978 gnd.n3280 gnd.n3179 19.3944
R15979 gnd.n3857 gnd.n3179 19.3944
R15980 gnd.n3857 gnd.n3172 19.3944
R15981 gnd.n3868 gnd.n3172 19.3944
R15982 gnd.n3868 gnd.n3168 19.3944
R15983 gnd.n3881 gnd.n3168 19.3944
R15984 gnd.n3881 gnd.n3880 19.3944
R15985 gnd.n3880 gnd.n3147 19.3944
R15986 gnd.n3905 gnd.n3147 19.3944
R15987 gnd.n3905 gnd.n3904 19.3944
R15988 gnd.n3904 gnd.n2954 19.3944
R15989 gnd.n4409 gnd.n2954 19.3944
R15990 gnd.n4409 gnd.n4408 19.3944
R15991 gnd.n4408 gnd.n4407 19.3944
R15992 gnd.n4407 gnd.n2958 19.3944
R15993 gnd.n2977 gnd.n2958 19.3944
R15994 gnd.n4395 gnd.n2977 19.3944
R15995 gnd.n4395 gnd.n4394 19.3944
R15996 gnd.n4394 gnd.n4393 19.3944
R15997 gnd.n4393 gnd.n2981 19.3944
R15998 gnd.n3002 gnd.n2981 19.3944
R15999 gnd.n4381 gnd.n3002 19.3944
R16000 gnd.n4381 gnd.n4380 19.3944
R16001 gnd.n4380 gnd.n4379 19.3944
R16002 gnd.n4379 gnd.n3006 19.3944
R16003 gnd.n3028 gnd.n3006 19.3944
R16004 gnd.n4367 gnd.n3028 19.3944
R16005 gnd.n4367 gnd.n4366 19.3944
R16006 gnd.n4366 gnd.n4365 19.3944
R16007 gnd.n5312 gnd.n5311 19.3944
R16008 gnd.n5311 gnd.n5194 19.3944
R16009 gnd.n5304 gnd.n5194 19.3944
R16010 gnd.n5304 gnd.n5303 19.3944
R16011 gnd.n5303 gnd.n5208 19.3944
R16012 gnd.n5296 gnd.n5208 19.3944
R16013 gnd.n5296 gnd.n5295 19.3944
R16014 gnd.n5295 gnd.n5220 19.3944
R16015 gnd.n5288 gnd.n5220 19.3944
R16016 gnd.n5288 gnd.n5287 19.3944
R16017 gnd.n5287 gnd.n5231 19.3944
R16018 gnd.n5280 gnd.n5231 19.3944
R16019 gnd.n5280 gnd.n5279 19.3944
R16020 gnd.n5279 gnd.n5243 19.3944
R16021 gnd.n5272 gnd.n5243 19.3944
R16022 gnd.n5272 gnd.n5271 19.3944
R16023 gnd.n2374 gnd.n2049 19.3944
R16024 gnd.n2374 gnd.n2050 19.3944
R16025 gnd.n2370 gnd.n2050 19.3944
R16026 gnd.n2370 gnd.n2053 19.3944
R16027 gnd.n2364 gnd.n2053 19.3944
R16028 gnd.n2364 gnd.n2363 19.3944
R16029 gnd.n2363 gnd.n2362 19.3944
R16030 gnd.n2362 gnd.n2060 19.3944
R16031 gnd.n2356 gnd.n2060 19.3944
R16032 gnd.n2356 gnd.n2355 19.3944
R16033 gnd.n2355 gnd.n2354 19.3944
R16034 gnd.n2354 gnd.n2068 19.3944
R16035 gnd.n2348 gnd.n2068 19.3944
R16036 gnd.n2348 gnd.n2347 19.3944
R16037 gnd.n2347 gnd.n2346 19.3944
R16038 gnd.n2346 gnd.n2076 19.3944
R16039 gnd.n2340 gnd.n2076 19.3944
R16040 gnd.n2340 gnd.n2339 19.3944
R16041 gnd.n2339 gnd.n2338 19.3944
R16042 gnd.n2338 gnd.n2084 19.3944
R16043 gnd.n2332 gnd.n2084 19.3944
R16044 gnd.n2332 gnd.n2331 19.3944
R16045 gnd.n2331 gnd.n2330 19.3944
R16046 gnd.n2330 gnd.n2092 19.3944
R16047 gnd.n2324 gnd.n2092 19.3944
R16048 gnd.n2324 gnd.n2323 19.3944
R16049 gnd.n2323 gnd.n2322 19.3944
R16050 gnd.n2322 gnd.n2100 19.3944
R16051 gnd.n2316 gnd.n2100 19.3944
R16052 gnd.n2316 gnd.n2315 19.3944
R16053 gnd.n2315 gnd.n2314 19.3944
R16054 gnd.n2314 gnd.n2108 19.3944
R16055 gnd.n2308 gnd.n2108 19.3944
R16056 gnd.n2308 gnd.n2307 19.3944
R16057 gnd.n2307 gnd.n2306 19.3944
R16058 gnd.n2306 gnd.n2116 19.3944
R16059 gnd.n2300 gnd.n2116 19.3944
R16060 gnd.n2300 gnd.n2299 19.3944
R16061 gnd.n2299 gnd.n2298 19.3944
R16062 gnd.n2298 gnd.n2124 19.3944
R16063 gnd.n2292 gnd.n2124 19.3944
R16064 gnd.n2292 gnd.n2291 19.3944
R16065 gnd.n2291 gnd.n2290 19.3944
R16066 gnd.n2290 gnd.n2132 19.3944
R16067 gnd.n2284 gnd.n2132 19.3944
R16068 gnd.n2284 gnd.n2283 19.3944
R16069 gnd.n2283 gnd.n2282 19.3944
R16070 gnd.n2282 gnd.n2140 19.3944
R16071 gnd.n2276 gnd.n2140 19.3944
R16072 gnd.n2276 gnd.n2275 19.3944
R16073 gnd.n2275 gnd.n2274 19.3944
R16074 gnd.n2274 gnd.n2148 19.3944
R16075 gnd.n2268 gnd.n2148 19.3944
R16076 gnd.n2268 gnd.n2267 19.3944
R16077 gnd.n2267 gnd.n2266 19.3944
R16078 gnd.n2266 gnd.n2156 19.3944
R16079 gnd.n2260 gnd.n2156 19.3944
R16080 gnd.n2260 gnd.n2259 19.3944
R16081 gnd.n2259 gnd.n2258 19.3944
R16082 gnd.n2258 gnd.n2164 19.3944
R16083 gnd.n2252 gnd.n2164 19.3944
R16084 gnd.n2252 gnd.n2251 19.3944
R16085 gnd.n2251 gnd.n2250 19.3944
R16086 gnd.n2250 gnd.n2172 19.3944
R16087 gnd.n2244 gnd.n2172 19.3944
R16088 gnd.n2244 gnd.n2243 19.3944
R16089 gnd.n2243 gnd.n2242 19.3944
R16090 gnd.n2242 gnd.n2180 19.3944
R16091 gnd.n2236 gnd.n2180 19.3944
R16092 gnd.n2236 gnd.n2235 19.3944
R16093 gnd.n2235 gnd.n2234 19.3944
R16094 gnd.n2234 gnd.n2188 19.3944
R16095 gnd.n2228 gnd.n2188 19.3944
R16096 gnd.n2228 gnd.n2227 19.3944
R16097 gnd.n2227 gnd.n2226 19.3944
R16098 gnd.n2226 gnd.n2196 19.3944
R16099 gnd.n2220 gnd.n2196 19.3944
R16100 gnd.n2220 gnd.n2219 19.3944
R16101 gnd.n2219 gnd.n2218 19.3944
R16102 gnd.n2218 gnd.n2204 19.3944
R16103 gnd.n2212 gnd.n2204 19.3944
R16104 gnd.n2212 gnd.n2211 19.3944
R16105 gnd.n2211 gnd.n245 19.3944
R16106 gnd.n7038 gnd.n245 19.3944
R16107 gnd.n2741 gnd.n2740 19.3944
R16108 gnd.n2740 gnd.n1685 19.3944
R16109 gnd.n2734 gnd.n1685 19.3944
R16110 gnd.n2734 gnd.n2733 19.3944
R16111 gnd.n2733 gnd.n2732 19.3944
R16112 gnd.n2732 gnd.n1694 19.3944
R16113 gnd.n2726 gnd.n1694 19.3944
R16114 gnd.n2726 gnd.n2725 19.3944
R16115 gnd.n2725 gnd.n2724 19.3944
R16116 gnd.n2724 gnd.n1702 19.3944
R16117 gnd.n2718 gnd.n1702 19.3944
R16118 gnd.n2718 gnd.n2717 19.3944
R16119 gnd.n2717 gnd.n2716 19.3944
R16120 gnd.n2716 gnd.n1710 19.3944
R16121 gnd.n2710 gnd.n1710 19.3944
R16122 gnd.n2710 gnd.n2709 19.3944
R16123 gnd.n2709 gnd.n2708 19.3944
R16124 gnd.n2708 gnd.n1718 19.3944
R16125 gnd.n2702 gnd.n1718 19.3944
R16126 gnd.n2702 gnd.n2701 19.3944
R16127 gnd.n2701 gnd.n2700 19.3944
R16128 gnd.n2700 gnd.n1726 19.3944
R16129 gnd.n2694 gnd.n1726 19.3944
R16130 gnd.n2694 gnd.n2693 19.3944
R16131 gnd.n2693 gnd.n2692 19.3944
R16132 gnd.n2692 gnd.n1734 19.3944
R16133 gnd.n2686 gnd.n1734 19.3944
R16134 gnd.n2686 gnd.n2685 19.3944
R16135 gnd.n2685 gnd.n2684 19.3944
R16136 gnd.n2684 gnd.n1742 19.3944
R16137 gnd.n2678 gnd.n1742 19.3944
R16138 gnd.n2678 gnd.n2677 19.3944
R16139 gnd.n2677 gnd.n2676 19.3944
R16140 gnd.n2676 gnd.n1750 19.3944
R16141 gnd.n2670 gnd.n1750 19.3944
R16142 gnd.n2670 gnd.n2669 19.3944
R16143 gnd.n2669 gnd.n2668 19.3944
R16144 gnd.n2668 gnd.n1758 19.3944
R16145 gnd.n2662 gnd.n1758 19.3944
R16146 gnd.n2662 gnd.n2661 19.3944
R16147 gnd.n2661 gnd.n2660 19.3944
R16148 gnd.n2660 gnd.n1766 19.3944
R16149 gnd.n2654 gnd.n1766 19.3944
R16150 gnd.n2654 gnd.n2653 19.3944
R16151 gnd.n2653 gnd.n2652 19.3944
R16152 gnd.n2652 gnd.n1774 19.3944
R16153 gnd.n2646 gnd.n1774 19.3944
R16154 gnd.n2646 gnd.n2645 19.3944
R16155 gnd.n2645 gnd.n2644 19.3944
R16156 gnd.n2644 gnd.n1782 19.3944
R16157 gnd.n2638 gnd.n1782 19.3944
R16158 gnd.n2638 gnd.n2637 19.3944
R16159 gnd.n2637 gnd.n2636 19.3944
R16160 gnd.n2636 gnd.n1790 19.3944
R16161 gnd.n2630 gnd.n1790 19.3944
R16162 gnd.n2630 gnd.n2629 19.3944
R16163 gnd.n2629 gnd.n2628 19.3944
R16164 gnd.n2628 gnd.n1798 19.3944
R16165 gnd.n2622 gnd.n1798 19.3944
R16166 gnd.n2622 gnd.n2621 19.3944
R16167 gnd.n2621 gnd.n2620 19.3944
R16168 gnd.n2620 gnd.n1806 19.3944
R16169 gnd.n2614 gnd.n1806 19.3944
R16170 gnd.n2614 gnd.n2613 19.3944
R16171 gnd.n2613 gnd.n2612 19.3944
R16172 gnd.n2612 gnd.n1814 19.3944
R16173 gnd.n2606 gnd.n1814 19.3944
R16174 gnd.n2606 gnd.n2605 19.3944
R16175 gnd.n2605 gnd.n2604 19.3944
R16176 gnd.n2604 gnd.n1822 19.3944
R16177 gnd.n2598 gnd.n1822 19.3944
R16178 gnd.n2598 gnd.n2597 19.3944
R16179 gnd.n2597 gnd.n2596 19.3944
R16180 gnd.n2596 gnd.n1830 19.3944
R16181 gnd.n2590 gnd.n1830 19.3944
R16182 gnd.n2590 gnd.n2589 19.3944
R16183 gnd.n2589 gnd.n2588 19.3944
R16184 gnd.n2588 gnd.n1838 19.3944
R16185 gnd.n2582 gnd.n1838 19.3944
R16186 gnd.n2582 gnd.n2581 19.3944
R16187 gnd.n2581 gnd.n2580 19.3944
R16188 gnd.n2580 gnd.n1846 19.3944
R16189 gnd.n2574 gnd.n1846 19.3944
R16190 gnd.n2574 gnd.n2573 19.3944
R16191 gnd.n2573 gnd.n2572 19.3944
R16192 gnd.n2572 gnd.n1854 19.3944
R16193 gnd.n2566 gnd.n1854 19.3944
R16194 gnd.n2566 gnd.n2565 19.3944
R16195 gnd.n2565 gnd.n2564 19.3944
R16196 gnd.n2564 gnd.n1862 19.3944
R16197 gnd.n2558 gnd.n1862 19.3944
R16198 gnd.n2558 gnd.n2557 19.3944
R16199 gnd.n2557 gnd.n2556 19.3944
R16200 gnd.n2556 gnd.n1870 19.3944
R16201 gnd.n2550 gnd.n1870 19.3944
R16202 gnd.n2550 gnd.n2549 19.3944
R16203 gnd.n2549 gnd.n2548 19.3944
R16204 gnd.n2548 gnd.n1878 19.3944
R16205 gnd.n2542 gnd.n1878 19.3944
R16206 gnd.n2542 gnd.n2541 19.3944
R16207 gnd.n2541 gnd.n2540 19.3944
R16208 gnd.n2540 gnd.n1886 19.3944
R16209 gnd.n2534 gnd.n1886 19.3944
R16210 gnd.n2534 gnd.n2533 19.3944
R16211 gnd.n2533 gnd.n2532 19.3944
R16212 gnd.n2532 gnd.n1894 19.3944
R16213 gnd.n2526 gnd.n1894 19.3944
R16214 gnd.n2526 gnd.n2525 19.3944
R16215 gnd.n2525 gnd.n2524 19.3944
R16216 gnd.n2524 gnd.n1902 19.3944
R16217 gnd.n2518 gnd.n1902 19.3944
R16218 gnd.n2518 gnd.n2517 19.3944
R16219 gnd.n2517 gnd.n2516 19.3944
R16220 gnd.n2516 gnd.n1910 19.3944
R16221 gnd.n2510 gnd.n1910 19.3944
R16222 gnd.n2510 gnd.n2509 19.3944
R16223 gnd.n2509 gnd.n2508 19.3944
R16224 gnd.n2508 gnd.n1918 19.3944
R16225 gnd.n2502 gnd.n1918 19.3944
R16226 gnd.n2502 gnd.n2501 19.3944
R16227 gnd.n2501 gnd.n2500 19.3944
R16228 gnd.n2500 gnd.n1926 19.3944
R16229 gnd.n2494 gnd.n1926 19.3944
R16230 gnd.n2494 gnd.n2493 19.3944
R16231 gnd.n2493 gnd.n2492 19.3944
R16232 gnd.n2492 gnd.n1934 19.3944
R16233 gnd.n2486 gnd.n1934 19.3944
R16234 gnd.n2486 gnd.n2485 19.3944
R16235 gnd.n2485 gnd.n2484 19.3944
R16236 gnd.n2484 gnd.n1942 19.3944
R16237 gnd.n2478 gnd.n1942 19.3944
R16238 gnd.n2478 gnd.n2477 19.3944
R16239 gnd.n2477 gnd.n2476 19.3944
R16240 gnd.n2476 gnd.n1950 19.3944
R16241 gnd.n2470 gnd.n1950 19.3944
R16242 gnd.n2470 gnd.n2469 19.3944
R16243 gnd.n2469 gnd.n2468 19.3944
R16244 gnd.n2468 gnd.n1958 19.3944
R16245 gnd.n2462 gnd.n1958 19.3944
R16246 gnd.n2462 gnd.n2461 19.3944
R16247 gnd.n2461 gnd.n2460 19.3944
R16248 gnd.n2460 gnd.n1966 19.3944
R16249 gnd.n2454 gnd.n1966 19.3944
R16250 gnd.n2454 gnd.n2453 19.3944
R16251 gnd.n2453 gnd.n2452 19.3944
R16252 gnd.n2452 gnd.n1974 19.3944
R16253 gnd.n2446 gnd.n1974 19.3944
R16254 gnd.n2446 gnd.n2445 19.3944
R16255 gnd.n2445 gnd.n2444 19.3944
R16256 gnd.n2444 gnd.n1982 19.3944
R16257 gnd.n2438 gnd.n1982 19.3944
R16258 gnd.n2438 gnd.n2437 19.3944
R16259 gnd.n2437 gnd.n2436 19.3944
R16260 gnd.n2436 gnd.n1990 19.3944
R16261 gnd.n2430 gnd.n1990 19.3944
R16262 gnd.n2430 gnd.n2429 19.3944
R16263 gnd.n2429 gnd.n2428 19.3944
R16264 gnd.n2428 gnd.n1998 19.3944
R16265 gnd.n2422 gnd.n1998 19.3944
R16266 gnd.n2422 gnd.n2421 19.3944
R16267 gnd.n2421 gnd.n2420 19.3944
R16268 gnd.n2420 gnd.n2006 19.3944
R16269 gnd.n2414 gnd.n2006 19.3944
R16270 gnd.n2414 gnd.n2413 19.3944
R16271 gnd.n2413 gnd.n2412 19.3944
R16272 gnd.n2412 gnd.n2014 19.3944
R16273 gnd.n2406 gnd.n2014 19.3944
R16274 gnd.n2406 gnd.n2405 19.3944
R16275 gnd.n2405 gnd.n2404 19.3944
R16276 gnd.n2404 gnd.n2022 19.3944
R16277 gnd.n2398 gnd.n2022 19.3944
R16278 gnd.n2398 gnd.n2397 19.3944
R16279 gnd.n2397 gnd.n2396 19.3944
R16280 gnd.n2396 gnd.n2030 19.3944
R16281 gnd.n2390 gnd.n2030 19.3944
R16282 gnd.n2390 gnd.n2389 19.3944
R16283 gnd.n2389 gnd.n2388 19.3944
R16284 gnd.n2388 gnd.n2038 19.3944
R16285 gnd.n2382 gnd.n2038 19.3944
R16286 gnd.n2382 gnd.n2381 19.3944
R16287 gnd.n2381 gnd.n2380 19.3944
R16288 gnd.n6690 gnd.n6689 19.3944
R16289 gnd.n6689 gnd.n6688 19.3944
R16290 gnd.n6688 gnd.n6687 19.3944
R16291 gnd.n6687 gnd.n6685 19.3944
R16292 gnd.n6685 gnd.n6682 19.3944
R16293 gnd.n6682 gnd.n6681 19.3944
R16294 gnd.n6681 gnd.n6678 19.3944
R16295 gnd.n6678 gnd.n6677 19.3944
R16296 gnd.n6677 gnd.n6674 19.3944
R16297 gnd.n6674 gnd.n6673 19.3944
R16298 gnd.n6673 gnd.n6670 19.3944
R16299 gnd.n6670 gnd.n6669 19.3944
R16300 gnd.n6669 gnd.n6666 19.3944
R16301 gnd.n6666 gnd.n6665 19.3944
R16302 gnd.n6665 gnd.n6662 19.3944
R16303 gnd.n6662 gnd.n6661 19.3944
R16304 gnd.n6661 gnd.n6658 19.3944
R16305 gnd.n6656 gnd.n6653 19.3944
R16306 gnd.n6653 gnd.n6652 19.3944
R16307 gnd.n6652 gnd.n6649 19.3944
R16308 gnd.n6649 gnd.n6648 19.3944
R16309 gnd.n6648 gnd.n6645 19.3944
R16310 gnd.n6645 gnd.n6644 19.3944
R16311 gnd.n6644 gnd.n6641 19.3944
R16312 gnd.n6639 gnd.n6636 19.3944
R16313 gnd.n6636 gnd.n6635 19.3944
R16314 gnd.n6635 gnd.n6632 19.3944
R16315 gnd.n6632 gnd.n6631 19.3944
R16316 gnd.n6631 gnd.n6628 19.3944
R16317 gnd.n6628 gnd.n6627 19.3944
R16318 gnd.n6627 gnd.n6624 19.3944
R16319 gnd.n6624 gnd.n6623 19.3944
R16320 gnd.n6619 gnd.n6616 19.3944
R16321 gnd.n6616 gnd.n6615 19.3944
R16322 gnd.n6615 gnd.n6612 19.3944
R16323 gnd.n6612 gnd.n6611 19.3944
R16324 gnd.n6611 gnd.n6608 19.3944
R16325 gnd.n6608 gnd.n6607 19.3944
R16326 gnd.n6607 gnd.n6604 19.3944
R16327 gnd.n6604 gnd.n6603 19.3944
R16328 gnd.n6603 gnd.n6600 19.3944
R16329 gnd.n6600 gnd.n6599 19.3944
R16330 gnd.n6599 gnd.n6596 19.3944
R16331 gnd.n6596 gnd.n6595 19.3944
R16332 gnd.n6595 gnd.n6592 19.3944
R16333 gnd.n6592 gnd.n6591 19.3944
R16334 gnd.n6591 gnd.n6588 19.3944
R16335 gnd.n6588 gnd.n6587 19.3944
R16336 gnd.n6587 gnd.n6584 19.3944
R16337 gnd.n6584 gnd.n6583 19.3944
R16338 gnd.n6730 gnd.n401 19.3944
R16339 gnd.n6730 gnd.n6729 19.3944
R16340 gnd.n6729 gnd.n411 19.3944
R16341 gnd.n411 gnd.n410 19.3944
R16342 gnd.n410 gnd.n408 19.3944
R16343 gnd.n408 gnd.n367 19.3944
R16344 gnd.n6792 gnd.n367 19.3944
R16345 gnd.n6793 gnd.n6792 19.3944
R16346 gnd.n6793 gnd.n339 19.3944
R16347 gnd.n6824 gnd.n339 19.3944
R16348 gnd.n6825 gnd.n6824 19.3944
R16349 gnd.n6828 gnd.n6825 19.3944
R16350 gnd.n6829 gnd.n6828 19.3944
R16351 gnd.n6829 gnd.n311 19.3944
R16352 gnd.n6867 gnd.n311 19.3944
R16353 gnd.n6867 gnd.n300 19.3944
R16354 gnd.n6879 gnd.n300 19.3944
R16355 gnd.n6881 gnd.n6879 19.3944
R16356 gnd.n6881 gnd.n6880 19.3944
R16357 gnd.n6880 gnd.n280 19.3944
R16358 gnd.n6917 gnd.n280 19.3944
R16359 gnd.n6919 gnd.n6917 19.3944
R16360 gnd.n6919 gnd.n6918 19.3944
R16361 gnd.n6918 gnd.n273 19.3944
R16362 gnd.n6929 gnd.n273 19.3944
R16363 gnd.n6930 gnd.n6929 19.3944
R16364 gnd.n6989 gnd.n6930 19.3944
R16365 gnd.n6989 gnd.n6988 19.3944
R16366 gnd.n6988 gnd.n6987 19.3944
R16367 gnd.n6987 gnd.n6932 19.3944
R16368 gnd.n6977 gnd.n6932 19.3944
R16369 gnd.n6977 gnd.n6976 19.3944
R16370 gnd.n6976 gnd.n6975 19.3944
R16371 gnd.n6975 gnd.n6940 19.3944
R16372 gnd.n6965 gnd.n6940 19.3944
R16373 gnd.n6965 gnd.n6964 19.3944
R16374 gnd.n6964 gnd.n6963 19.3944
R16375 gnd.n6963 gnd.n6947 19.3944
R16376 gnd.n6953 gnd.n6947 19.3944
R16377 gnd.n6953 gnd.n175 19.3944
R16378 gnd.n7264 gnd.n175 19.3944
R16379 gnd.n7265 gnd.n7264 19.3944
R16380 gnd.n6732 gnd.n397 19.3944
R16381 gnd.n6732 gnd.n398 19.3944
R16382 gnd.n403 gnd.n398 19.3944
R16383 gnd.n405 gnd.n403 19.3944
R16384 gnd.n405 gnd.n364 19.3944
R16385 gnd.n6801 gnd.n364 19.3944
R16386 gnd.n6801 gnd.n6800 19.3944
R16387 gnd.n6800 gnd.n6799 19.3944
R16388 gnd.n6799 gnd.n6798 19.3944
R16389 gnd.n6798 gnd.n336 19.3944
R16390 gnd.n6836 gnd.n336 19.3944
R16391 gnd.n6836 gnd.n6835 19.3944
R16392 gnd.n6835 gnd.n6834 19.3944
R16393 gnd.n6834 gnd.n6833 19.3944
R16394 gnd.n6833 gnd.n309 19.3944
R16395 gnd.n6870 gnd.n309 19.3944
R16396 gnd.n6870 gnd.n298 19.3944
R16397 gnd.n6883 gnd.n298 19.3944
R16398 gnd.n6883 gnd.n282 19.3944
R16399 gnd.n6914 gnd.n282 19.3944
R16400 gnd.n6914 gnd.n275 19.3944
R16401 gnd.n6923 gnd.n275 19.3944
R16402 gnd.n6924 gnd.n6923 19.3944
R16403 gnd.n6926 gnd.n6924 19.3944
R16404 gnd.n6926 gnd.n92 19.3944
R16405 gnd.n7315 gnd.n92 19.3944
R16406 gnd.n7315 gnd.n7314 19.3944
R16407 gnd.n7314 gnd.n7313 19.3944
R16408 gnd.n7313 gnd.n96 19.3944
R16409 gnd.n7303 gnd.n96 19.3944
R16410 gnd.n7303 gnd.n7302 19.3944
R16411 gnd.n7302 gnd.n7301 19.3944
R16412 gnd.n7301 gnd.n115 19.3944
R16413 gnd.n7291 gnd.n115 19.3944
R16414 gnd.n7291 gnd.n7290 19.3944
R16415 gnd.n7290 gnd.n7289 19.3944
R16416 gnd.n7289 gnd.n136 19.3944
R16417 gnd.n7279 gnd.n136 19.3944
R16418 gnd.n7279 gnd.n7278 19.3944
R16419 gnd.n7278 gnd.n7277 19.3944
R16420 gnd.n7277 gnd.n157 19.3944
R16421 gnd.n7267 gnd.n157 19.3944
R16422 gnd.n7174 gnd.n7110 19.3944
R16423 gnd.n7174 gnd.n7171 19.3944
R16424 gnd.n7171 gnd.n7168 19.3944
R16425 gnd.n7168 gnd.n7167 19.3944
R16426 gnd.n7167 gnd.n7164 19.3944
R16427 gnd.n7164 gnd.n7163 19.3944
R16428 gnd.n7163 gnd.n7160 19.3944
R16429 gnd.n7160 gnd.n7159 19.3944
R16430 gnd.n7159 gnd.n7156 19.3944
R16431 gnd.n7156 gnd.n7155 19.3944
R16432 gnd.n7155 gnd.n7152 19.3944
R16433 gnd.n7152 gnd.n7151 19.3944
R16434 gnd.n7151 gnd.n7148 19.3944
R16435 gnd.n7148 gnd.n7147 19.3944
R16436 gnd.n7147 gnd.n7144 19.3944
R16437 gnd.n7144 gnd.n7143 19.3944
R16438 gnd.n7143 gnd.n7140 19.3944
R16439 gnd.n7140 gnd.n7139 19.3944
R16440 gnd.n7217 gnd.n7214 19.3944
R16441 gnd.n7214 gnd.n7213 19.3944
R16442 gnd.n7213 gnd.n7210 19.3944
R16443 gnd.n7210 gnd.n7209 19.3944
R16444 gnd.n7209 gnd.n7206 19.3944
R16445 gnd.n7206 gnd.n7205 19.3944
R16446 gnd.n7205 gnd.n7202 19.3944
R16447 gnd.n7202 gnd.n7201 19.3944
R16448 gnd.n7201 gnd.n7198 19.3944
R16449 gnd.n7198 gnd.n7197 19.3944
R16450 gnd.n7197 gnd.n7194 19.3944
R16451 gnd.n7194 gnd.n7193 19.3944
R16452 gnd.n7193 gnd.n7190 19.3944
R16453 gnd.n7190 gnd.n7189 19.3944
R16454 gnd.n7189 gnd.n7186 19.3944
R16455 gnd.n7186 gnd.n7185 19.3944
R16456 gnd.n7185 gnd.n7182 19.3944
R16457 gnd.n7182 gnd.n7181 19.3944
R16458 gnd.n7072 gnd.n7071 19.3944
R16459 gnd.n7250 gnd.n7071 19.3944
R16460 gnd.n7250 gnd.n7249 19.3944
R16461 gnd.n7249 gnd.n7248 19.3944
R16462 gnd.n7248 gnd.n7245 19.3944
R16463 gnd.n7245 gnd.n7244 19.3944
R16464 gnd.n7244 gnd.n7241 19.3944
R16465 gnd.n7241 gnd.n7240 19.3944
R16466 gnd.n7240 gnd.n7237 19.3944
R16467 gnd.n7237 gnd.n7236 19.3944
R16468 gnd.n7236 gnd.n7233 19.3944
R16469 gnd.n7233 gnd.n7232 19.3944
R16470 gnd.n7232 gnd.n7229 19.3944
R16471 gnd.n7229 gnd.n7228 19.3944
R16472 gnd.n7228 gnd.n7225 19.3944
R16473 gnd.n7225 gnd.n7224 19.3944
R16474 gnd.n7224 gnd.n7221 19.3944
R16475 gnd.n203 gnd.n201 19.3944
R16476 gnd.n206 gnd.n203 19.3944
R16477 gnd.n206 gnd.n198 19.3944
R16478 gnd.n210 gnd.n198 19.3944
R16479 gnd.n213 gnd.n210 19.3944
R16480 gnd.n216 gnd.n213 19.3944
R16481 gnd.n216 gnd.n196 19.3944
R16482 gnd.n220 gnd.n196 19.3944
R16483 gnd.n223 gnd.n220 19.3944
R16484 gnd.n226 gnd.n223 19.3944
R16485 gnd.n226 gnd.n194 19.3944
R16486 gnd.n230 gnd.n194 19.3944
R16487 gnd.n233 gnd.n230 19.3944
R16488 gnd.n235 gnd.n233 19.3944
R16489 gnd.n235 gnd.n192 19.3944
R16490 gnd.n239 gnd.n192 19.3944
R16491 gnd.n6713 gnd.n421 19.3944
R16492 gnd.n421 gnd.n380 19.3944
R16493 gnd.n6746 gnd.n380 19.3944
R16494 gnd.n6746 gnd.n377 19.3944
R16495 gnd.n6751 gnd.n377 19.3944
R16496 gnd.n6751 gnd.n378 19.3944
R16497 gnd.n378 gnd.n347 19.3944
R16498 gnd.n6815 gnd.n347 19.3944
R16499 gnd.n6815 gnd.n344 19.3944
R16500 gnd.n6820 gnd.n344 19.3944
R16501 gnd.n6820 gnd.n345 19.3944
R16502 gnd.n345 gnd.n318 19.3944
R16503 gnd.n6851 gnd.n318 19.3944
R16504 gnd.n6851 gnd.n315 19.3944
R16505 gnd.n6863 gnd.n315 19.3944
R16506 gnd.n6863 gnd.n316 19.3944
R16507 gnd.n6859 gnd.n316 19.3944
R16508 gnd.n6859 gnd.n6858 19.3944
R16509 gnd.n6858 gnd.n6857 19.3944
R16510 gnd.n6857 gnd.n6855 19.3944
R16511 gnd.n6855 gnd.n64 19.3944
R16512 gnd.n7328 gnd.n64 19.3944
R16513 gnd.n7328 gnd.n7327 19.3944
R16514 gnd.n7327 gnd.n67 19.3944
R16515 gnd.n6995 gnd.n67 19.3944
R16516 gnd.n6995 gnd.n6994 19.3944
R16517 gnd.n6994 gnd.n6993 19.3944
R16518 gnd.n6993 gnd.n271 19.3944
R16519 gnd.n6983 gnd.n271 19.3944
R16520 gnd.n6983 gnd.n6982 19.3944
R16521 gnd.n6982 gnd.n6981 19.3944
R16522 gnd.n6981 gnd.n6937 19.3944
R16523 gnd.n6971 gnd.n6937 19.3944
R16524 gnd.n6971 gnd.n6970 19.3944
R16525 gnd.n6970 gnd.n6969 19.3944
R16526 gnd.n6969 gnd.n6945 19.3944
R16527 gnd.n6959 gnd.n6945 19.3944
R16528 gnd.n6959 gnd.n6958 19.3944
R16529 gnd.n6958 gnd.n6957 19.3944
R16530 gnd.n6957 gnd.n177 19.3944
R16531 gnd.n7260 gnd.n177 19.3944
R16532 gnd.n7260 gnd.n7259 19.3944
R16533 gnd.n6736 gnd.n390 19.3944
R16534 gnd.n6736 gnd.n388 19.3944
R16535 gnd.n6742 gnd.n388 19.3944
R16536 gnd.n6742 gnd.n6741 19.3944
R16537 gnd.n6741 gnd.n357 19.3944
R16538 gnd.n6805 gnd.n357 19.3944
R16539 gnd.n6805 gnd.n355 19.3944
R16540 gnd.n6811 gnd.n355 19.3944
R16541 gnd.n6811 gnd.n6810 19.3944
R16542 gnd.n6810 gnd.n328 19.3944
R16543 gnd.n6840 gnd.n328 19.3944
R16544 gnd.n6840 gnd.n326 19.3944
R16545 gnd.n6847 gnd.n326 19.3944
R16546 gnd.n6847 gnd.n6846 19.3944
R16547 gnd.n6846 gnd.n6845 19.3944
R16548 gnd.n6845 gnd.n305 19.3944
R16549 gnd.n6875 gnd.n6874 19.3944
R16550 gnd.n6910 gnd.n6909 19.3944
R16551 gnd.n6905 gnd.n6904 19.3944
R16552 gnd.n7323 gnd.n7322 19.3944
R16553 gnd.n7319 gnd.n76 19.3944
R16554 gnd.n7319 gnd.n83 19.3944
R16555 gnd.n7309 gnd.n83 19.3944
R16556 gnd.n7309 gnd.n7308 19.3944
R16557 gnd.n7308 gnd.n7307 19.3944
R16558 gnd.n7307 gnd.n106 19.3944
R16559 gnd.n7297 gnd.n106 19.3944
R16560 gnd.n7297 gnd.n7296 19.3944
R16561 gnd.n7296 gnd.n7295 19.3944
R16562 gnd.n7295 gnd.n126 19.3944
R16563 gnd.n7285 gnd.n126 19.3944
R16564 gnd.n7285 gnd.n7284 19.3944
R16565 gnd.n7284 gnd.n7283 19.3944
R16566 gnd.n7283 gnd.n147 19.3944
R16567 gnd.n7273 gnd.n147 19.3944
R16568 gnd.n7273 gnd.n7272 19.3944
R16569 gnd.n7272 gnd.n7271 19.3944
R16570 gnd.n4450 gnd.n4449 19.3944
R16571 gnd.n4449 gnd.n4448 19.3944
R16572 gnd.n4448 gnd.n4421 19.3944
R16573 gnd.n4444 gnd.n4421 19.3944
R16574 gnd.n4444 gnd.n4443 19.3944
R16575 gnd.n4443 gnd.n4442 19.3944
R16576 gnd.n4442 gnd.n4427 19.3944
R16577 gnd.n4438 gnd.n4427 19.3944
R16578 gnd.n4438 gnd.n4437 19.3944
R16579 gnd.n4437 gnd.n4436 19.3944
R16580 gnd.n4436 gnd.n4434 19.3944
R16581 gnd.n4434 gnd.n1447 19.3944
R16582 gnd.n4803 gnd.n1447 19.3944
R16583 gnd.n4803 gnd.n1445 19.3944
R16584 gnd.n4809 gnd.n1445 19.3944
R16585 gnd.n4809 gnd.n4808 19.3944
R16586 gnd.n4808 gnd.n1414 19.3944
R16587 gnd.n4858 gnd.n4857 19.3944
R16588 gnd.n4861 gnd.n4860 19.3944
R16589 gnd.n4906 gnd.n4905 19.3944
R16590 gnd.n4903 gnd.n1382 19.3944
R16591 gnd.n1398 gnd.n1397 19.3944
R16592 gnd.n1397 gnd.n1332 19.3944
R16593 gnd.n4943 gnd.n1332 19.3944
R16594 gnd.n4943 gnd.n1330 19.3944
R16595 gnd.n4958 gnd.n1330 19.3944
R16596 gnd.n4958 gnd.n4957 19.3944
R16597 gnd.n4957 gnd.n4956 19.3944
R16598 gnd.n4956 gnd.n4949 19.3944
R16599 gnd.n4952 gnd.n4949 19.3944
R16600 gnd.n4952 gnd.n1282 19.3944
R16601 gnd.n5019 gnd.n1282 19.3944
R16602 gnd.n5019 gnd.n1280 19.3944
R16603 gnd.n5023 gnd.n1280 19.3944
R16604 gnd.n5023 gnd.n1278 19.3944
R16605 gnd.n5029 gnd.n1278 19.3944
R16606 gnd.n5029 gnd.n1276 19.3944
R16607 gnd.n5187 gnd.n1276 19.3944
R16608 gnd.n5187 gnd.n5186 19.3944
R16609 gnd.n5186 gnd.n5185 19.3944
R16610 gnd.n5185 gnd.n5035 19.3944
R16611 gnd.n5179 gnd.n5035 19.3944
R16612 gnd.n5179 gnd.n5178 19.3944
R16613 gnd.n5178 gnd.n5177 19.3944
R16614 gnd.n5177 gnd.n5041 19.3944
R16615 gnd.n5101 gnd.n5041 19.3944
R16616 gnd.n5101 gnd.n5098 19.3944
R16617 gnd.n5105 gnd.n5098 19.3944
R16618 gnd.n5105 gnd.n5079 19.3944
R16619 gnd.n5122 gnd.n5079 19.3944
R16620 gnd.n5122 gnd.n5077 19.3944
R16621 gnd.n5126 gnd.n5077 19.3944
R16622 gnd.n5126 gnd.n5066 19.3944
R16623 gnd.n5143 gnd.n5066 19.3944
R16624 gnd.n5143 gnd.n5064 19.3944
R16625 gnd.n5149 gnd.n5064 19.3944
R16626 gnd.n5149 gnd.n5148 19.3944
R16627 gnd.n5148 gnd.n1068 19.3944
R16628 gnd.n5630 gnd.n1068 19.3944
R16629 gnd.n5630 gnd.n1066 19.3944
R16630 gnd.n5646 gnd.n1066 19.3944
R16631 gnd.n5646 gnd.n5645 19.3944
R16632 gnd.n5645 gnd.n5644 19.3944
R16633 gnd.n5644 gnd.n5636 19.3944
R16634 gnd.n5639 gnd.n5636 19.3944
R16635 gnd.n5639 gnd.n986 19.3944
R16636 gnd.n5696 gnd.n986 19.3944
R16637 gnd.n5696 gnd.n984 19.3944
R16638 gnd.n5702 gnd.n984 19.3944
R16639 gnd.n5702 gnd.n5701 19.3944
R16640 gnd.n5701 gnd.n924 19.3944
R16641 gnd.n5767 gnd.n924 19.3944
R16642 gnd.n5767 gnd.n922 19.3944
R16643 gnd.n5771 gnd.n922 19.3944
R16644 gnd.n5771 gnd.n920 19.3944
R16645 gnd.n5775 gnd.n920 19.3944
R16646 gnd.n5775 gnd.n918 19.3944
R16647 gnd.n5779 gnd.n918 19.3944
R16648 gnd.n5779 gnd.n869 19.3944
R16649 gnd.n5868 gnd.n869 19.3944
R16650 gnd.n5868 gnd.n867 19.3944
R16651 gnd.n5880 gnd.n867 19.3944
R16652 gnd.n5880 gnd.n5879 19.3944
R16653 gnd.n5879 gnd.n5878 19.3944
R16654 gnd.n5878 gnd.n5875 19.3944
R16655 gnd.n5875 gnd.n830 19.3944
R16656 gnd.n5925 gnd.n830 19.3944
R16657 gnd.n5925 gnd.n828 19.3944
R16658 gnd.n5934 gnd.n828 19.3944
R16659 gnd.n5934 gnd.n5933 19.3944
R16660 gnd.n5933 gnd.n5932 19.3944
R16661 gnd.n5932 gnd.n783 19.3944
R16662 gnd.n6080 gnd.n783 19.3944
R16663 gnd.n6080 gnd.n781 19.3944
R16664 gnd.n6086 gnd.n781 19.3944
R16665 gnd.n6086 gnd.n6085 19.3944
R16666 gnd.n6085 gnd.n754 19.3944
R16667 gnd.n6116 gnd.n754 19.3944
R16668 gnd.n6116 gnd.n752 19.3944
R16669 gnd.n6120 gnd.n752 19.3944
R16670 gnd.n6120 gnd.n731 19.3944
R16671 gnd.n6143 gnd.n731 19.3944
R16672 gnd.n6143 gnd.n729 19.3944
R16673 gnd.n6147 gnd.n729 19.3944
R16674 gnd.n6147 gnd.n705 19.3944
R16675 gnd.n6182 gnd.n705 19.3944
R16676 gnd.n6182 gnd.n703 19.3944
R16677 gnd.n6186 gnd.n703 19.3944
R16678 gnd.n6186 gnd.n652 19.3944
R16679 gnd.n6354 gnd.n652 19.3944
R16680 gnd.n6354 gnd.n650 19.3944
R16681 gnd.n6360 gnd.n650 19.3944
R16682 gnd.n6360 gnd.n6359 19.3944
R16683 gnd.n6359 gnd.n627 19.3944
R16684 gnd.n6384 gnd.n627 19.3944
R16685 gnd.n6384 gnd.n625 19.3944
R16686 gnd.n6390 gnd.n625 19.3944
R16687 gnd.n6390 gnd.n6389 19.3944
R16688 gnd.n6389 gnd.n602 19.3944
R16689 gnd.n6414 gnd.n602 19.3944
R16690 gnd.n6414 gnd.n600 19.3944
R16691 gnd.n6420 gnd.n600 19.3944
R16692 gnd.n6420 gnd.n6419 19.3944
R16693 gnd.n6419 gnd.n577 19.3944
R16694 gnd.n6444 gnd.n577 19.3944
R16695 gnd.n6444 gnd.n575 19.3944
R16696 gnd.n6460 gnd.n575 19.3944
R16697 gnd.n6460 gnd.n6459 19.3944
R16698 gnd.n6459 gnd.n6458 19.3944
R16699 gnd.n6458 gnd.n6450 19.3944
R16700 gnd.n6453 gnd.n6450 19.3944
R16701 gnd.n6453 gnd.n416 19.3944
R16702 gnd.n6718 gnd.n416 19.3944
R16703 gnd.n6718 gnd.n414 19.3944
R16704 gnd.n6724 gnd.n414 19.3944
R16705 gnd.n6724 gnd.n6723 19.3944
R16706 gnd.n6723 gnd.n372 19.3944
R16707 gnd.n6756 gnd.n372 19.3944
R16708 gnd.n6756 gnd.n370 19.3944
R16709 gnd.n6787 gnd.n370 19.3944
R16710 gnd.n6787 gnd.n6786 19.3944
R16711 gnd.n6786 gnd.n6785 19.3944
R16712 gnd.n6785 gnd.n6762 19.3944
R16713 gnd.n6781 gnd.n6762 19.3944
R16714 gnd.n6781 gnd.n6780 19.3944
R16715 gnd.n6780 gnd.n6779 19.3944
R16716 gnd.n6779 gnd.n6768 19.3944
R16717 gnd.n6775 gnd.n6768 19.3944
R16718 gnd.n6775 gnd.n6774 19.3944
R16719 gnd.n6774 gnd.n6773 19.3944
R16720 gnd.n6889 gnd.n6888 19.3944
R16721 gnd.n6899 gnd.n6898 19.3944
R16722 gnd.n6896 gnd.n6893 19.3944
R16723 gnd.n6891 gnd.n264 19.3944
R16724 gnd.n7002 gnd.n7001 19.3944
R16725 gnd.n7005 gnd.n7002 19.3944
R16726 gnd.n7005 gnd.n260 19.3944
R16727 gnd.n7009 gnd.n260 19.3944
R16728 gnd.n7009 gnd.n258 19.3944
R16729 gnd.n7013 gnd.n258 19.3944
R16730 gnd.n7013 gnd.n256 19.3944
R16731 gnd.n7017 gnd.n256 19.3944
R16732 gnd.n7017 gnd.n254 19.3944
R16733 gnd.n7021 gnd.n254 19.3944
R16734 gnd.n7021 gnd.n252 19.3944
R16735 gnd.n7025 gnd.n252 19.3944
R16736 gnd.n7025 gnd.n250 19.3944
R16737 gnd.n7030 gnd.n250 19.3944
R16738 gnd.n7030 gnd.n248 19.3944
R16739 gnd.n7034 gnd.n248 19.3944
R16740 gnd.n7035 gnd.n7034 19.3944
R16741 gnd.n4706 gnd.n1514 19.3944
R16742 gnd.n4701 gnd.n1514 19.3944
R16743 gnd.n4701 gnd.n4700 19.3944
R16744 gnd.n4700 gnd.n4699 19.3944
R16745 gnd.n4699 gnd.n4696 19.3944
R16746 gnd.n4696 gnd.n4695 19.3944
R16747 gnd.n4695 gnd.n4692 19.3944
R16748 gnd.n4692 gnd.n4691 19.3944
R16749 gnd.n4691 gnd.n4688 19.3944
R16750 gnd.n4688 gnd.n4687 19.3944
R16751 gnd.n4687 gnd.n4684 19.3944
R16752 gnd.n4684 gnd.n4683 19.3944
R16753 gnd.n4683 gnd.n4680 19.3944
R16754 gnd.n4680 gnd.n4679 19.3944
R16755 gnd.n4679 gnd.n4676 19.3944
R16756 gnd.n4676 gnd.n4675 19.3944
R16757 gnd.n4675 gnd.n4672 19.3944
R16758 gnd.n4670 gnd.n4667 19.3944
R16759 gnd.n4667 gnd.n4666 19.3944
R16760 gnd.n4666 gnd.n4663 19.3944
R16761 gnd.n4663 gnd.n4662 19.3944
R16762 gnd.n4662 gnd.n4659 19.3944
R16763 gnd.n4659 gnd.n4658 19.3944
R16764 gnd.n4658 gnd.n4655 19.3944
R16765 gnd.n4655 gnd.n4654 19.3944
R16766 gnd.n4654 gnd.n4651 19.3944
R16767 gnd.n4651 gnd.n4650 19.3944
R16768 gnd.n4650 gnd.n4647 19.3944
R16769 gnd.n4647 gnd.n4646 19.3944
R16770 gnd.n4646 gnd.n4643 19.3944
R16771 gnd.n4643 gnd.n4642 19.3944
R16772 gnd.n4642 gnd.n4639 19.3944
R16773 gnd.n4639 gnd.n4638 19.3944
R16774 gnd.n4638 gnd.n4635 19.3944
R16775 gnd.n4635 gnd.n4634 19.3944
R16776 gnd.n4630 gnd.n4627 19.3944
R16777 gnd.n4627 gnd.n4626 19.3944
R16778 gnd.n4626 gnd.n4623 19.3944
R16779 gnd.n4623 gnd.n4622 19.3944
R16780 gnd.n4622 gnd.n4619 19.3944
R16781 gnd.n4619 gnd.n4618 19.3944
R16782 gnd.n4618 gnd.n4615 19.3944
R16783 gnd.n4615 gnd.n4614 19.3944
R16784 gnd.n4614 gnd.n4611 19.3944
R16785 gnd.n4611 gnd.n4610 19.3944
R16786 gnd.n4610 gnd.n4607 19.3944
R16787 gnd.n4607 gnd.n4606 19.3944
R16788 gnd.n4606 gnd.n4603 19.3944
R16789 gnd.n4603 gnd.n4602 19.3944
R16790 gnd.n4602 gnd.n4599 19.3944
R16791 gnd.n4599 gnd.n4598 19.3944
R16792 gnd.n4598 gnd.n4595 19.3944
R16793 gnd.n4595 gnd.n4594 19.3944
R16794 gnd.n4581 gnd.n4580 19.3944
R16795 gnd.n4580 gnd.n4577 19.3944
R16796 gnd.n4577 gnd.n4576 19.3944
R16797 gnd.n4576 gnd.n4573 19.3944
R16798 gnd.n4573 gnd.n4572 19.3944
R16799 gnd.n4572 gnd.n4569 19.3944
R16800 gnd.n4569 gnd.n4568 19.3944
R16801 gnd.n4568 gnd.n4565 19.3944
R16802 gnd.n4565 gnd.n4564 19.3944
R16803 gnd.n4564 gnd.n4561 19.3944
R16804 gnd.n4561 gnd.n4560 19.3944
R16805 gnd.n4560 gnd.n4557 19.3944
R16806 gnd.n4557 gnd.n4556 19.3944
R16807 gnd.n4556 gnd.n4553 19.3944
R16808 gnd.n4553 gnd.n4552 19.3944
R16809 gnd.n4552 gnd.n4549 19.3944
R16810 gnd.n4716 gnd.n1504 19.3944
R16811 gnd.n4716 gnd.n1502 19.3944
R16812 gnd.n4726 gnd.n1502 19.3944
R16813 gnd.n4726 gnd.n4725 19.3944
R16814 gnd.n4725 gnd.n4724 19.3944
R16815 gnd.n4724 gnd.n1477 19.3944
R16816 gnd.n4752 gnd.n1477 19.3944
R16817 gnd.n4752 gnd.n1475 19.3944
R16818 gnd.n4757 gnd.n1475 19.3944
R16819 gnd.n4757 gnd.n1452 19.3944
R16820 gnd.n4797 gnd.n1452 19.3944
R16821 gnd.n4797 gnd.n4796 19.3944
R16822 gnd.n4796 gnd.n4795 19.3944
R16823 gnd.n4795 gnd.n1420 19.3944
R16824 gnd.n4829 gnd.n1420 19.3944
R16825 gnd.n4829 gnd.n1418 19.3944
R16826 gnd.n4851 gnd.n1418 19.3944
R16827 gnd.n4851 gnd.n4850 19.3944
R16828 gnd.n4850 gnd.n4849 19.3944
R16829 gnd.n4849 gnd.n4848 19.3944
R16830 gnd.n4848 gnd.n4847 19.3944
R16831 gnd.n4847 gnd.n4836 19.3944
R16832 gnd.n4843 gnd.n4836 19.3944
R16833 gnd.n4843 gnd.n4842 19.3944
R16834 gnd.n4842 gnd.n4841 19.3944
R16835 gnd.n4841 gnd.n1340 19.3944
R16836 gnd.n4933 gnd.n1340 19.3944
R16837 gnd.n4933 gnd.n1337 19.3944
R16838 gnd.n4938 gnd.n1337 19.3944
R16839 gnd.n4938 gnd.n1338 19.3944
R16840 gnd.n1338 gnd.n1307 19.3944
R16841 gnd.n4986 gnd.n1307 19.3944
R16842 gnd.n4986 gnd.n1304 19.3944
R16843 gnd.n4994 gnd.n1304 19.3944
R16844 gnd.n4994 gnd.n1305 19.3944
R16845 gnd.n4990 gnd.n1305 19.3944
R16846 gnd.n4990 gnd.n1234 19.3944
R16847 gnd.n5344 gnd.n1234 19.3944
R16848 gnd.n5344 gnd.n1235 19.3944
R16849 gnd.n5340 gnd.n1235 19.3944
R16850 gnd.n5340 gnd.n5339 19.3944
R16851 gnd.n5339 gnd.n5338 19.3944
R16852 gnd.n4586 gnd.n4524 19.3944
R16853 gnd.n4524 gnd.n1497 19.3944
R16854 gnd.n4730 gnd.n1497 19.3944
R16855 gnd.n4731 gnd.n4730 19.3944
R16856 gnd.n4732 gnd.n4731 19.3944
R16857 gnd.n4732 gnd.n1480 19.3944
R16858 gnd.n1480 gnd.n1474 19.3944
R16859 gnd.n4762 gnd.n1474 19.3944
R16860 gnd.n4762 gnd.n4761 19.3944
R16861 gnd.n4761 gnd.n1456 19.3944
R16862 gnd.n4779 gnd.n1456 19.3944
R16863 gnd.n4780 gnd.n4779 19.3944
R16864 gnd.n4791 gnd.n4780 19.3944
R16865 gnd.n4791 gnd.n4790 19.3944
R16866 gnd.n4790 gnd.n4789 19.3944
R16867 gnd.n4789 gnd.n4788 19.3944
R16868 gnd.n4788 gnd.n4786 19.3944
R16869 gnd.n4786 gnd.n1409 19.3944
R16870 gnd.n4866 gnd.n1409 19.3944
R16871 gnd.n4867 gnd.n4866 19.3944
R16872 gnd.n4868 gnd.n4867 19.3944
R16873 gnd.n4871 gnd.n4868 19.3944
R16874 gnd.n4871 gnd.n1407 19.3944
R16875 gnd.n4879 gnd.n1407 19.3944
R16876 gnd.n4880 gnd.n4879 19.3944
R16877 gnd.n4883 gnd.n4880 19.3944
R16878 gnd.n4884 gnd.n4883 19.3944
R16879 gnd.n4887 gnd.n4884 19.3944
R16880 gnd.n4887 gnd.n4885 19.3944
R16881 gnd.n4885 gnd.n1327 19.3944
R16882 gnd.n4963 gnd.n1327 19.3944
R16883 gnd.n4964 gnd.n4963 19.3944
R16884 gnd.n4964 gnd.n1299 19.3944
R16885 gnd.n4998 gnd.n1299 19.3944
R16886 gnd.n4999 gnd.n4998 19.3944
R16887 gnd.n5001 gnd.n4999 19.3944
R16888 gnd.n5001 gnd.n1230 19.3944
R16889 gnd.n5348 gnd.n1230 19.3944
R16890 gnd.n5349 gnd.n5348 19.3944
R16891 gnd.n5349 gnd.n1211 19.3944
R16892 gnd.n5460 gnd.n1211 19.3944
R16893 gnd.n5461 gnd.n5460 19.3944
R16894 gnd.n4518 gnd.n4517 19.3944
R16895 gnd.n4521 gnd.n4518 19.3944
R16896 gnd.n4521 gnd.n1495 19.3944
R16897 gnd.n4737 gnd.n1495 19.3944
R16898 gnd.n4737 gnd.n4736 19.3944
R16899 gnd.n4736 gnd.n4735 19.3944
R16900 gnd.n4735 gnd.n1472 19.3944
R16901 gnd.n4764 gnd.n1472 19.3944
R16902 gnd.n4764 gnd.n1458 19.3944
R16903 gnd.n4776 gnd.n1458 19.3944
R16904 gnd.n4776 gnd.n1437 19.3944
R16905 gnd.n4816 gnd.n1437 19.3944
R16906 gnd.n4816 gnd.n4815 19.3944
R16907 gnd.n4815 gnd.n4814 19.3944
R16908 gnd.n4814 gnd.n1441 19.3944
R16909 gnd.n4783 gnd.n1441 19.3944
R16910 gnd.n4783 gnd.n1364 19.3944
R16911 gnd.n4918 gnd.n1364 19.3944
R16912 gnd.n4918 gnd.n4917 19.3944
R16913 gnd.n4917 gnd.n4916 19.3944
R16914 gnd.n4916 gnd.n1368 19.3944
R16915 gnd.n4873 gnd.n1368 19.3944
R16916 gnd.n4876 gnd.n4873 19.3944
R16917 gnd.n4876 gnd.n1402 19.3944
R16918 gnd.n4893 gnd.n1402 19.3944
R16919 gnd.n4893 gnd.n4892 19.3944
R16920 gnd.n4892 gnd.n4891 19.3944
R16921 gnd.n4891 gnd.n4890 19.3944
R16922 gnd.n4890 gnd.n1324 19.3944
R16923 gnd.n4972 gnd.n1324 19.3944
R16924 gnd.n4972 gnd.n4971 19.3944
R16925 gnd.n4971 gnd.n4970 19.3944
R16926 gnd.n4970 gnd.n4969 19.3944
R16927 gnd.n4969 gnd.n1297 19.3944
R16928 gnd.n5006 gnd.n1297 19.3944
R16929 gnd.n5006 gnd.n5005 19.3944
R16930 gnd.n5005 gnd.n5004 19.3944
R16931 gnd.n5004 gnd.n1228 19.3944
R16932 gnd.n5354 gnd.n1228 19.3944
R16933 gnd.n5354 gnd.n5353 19.3944
R16934 gnd.n5353 gnd.n5352 19.3944
R16935 gnd.n5352 gnd.n1210 19.3944
R16936 gnd.n5452 gnd.n5363 19.3944
R16937 gnd.n5447 gnd.n5363 19.3944
R16938 gnd.n5447 gnd.n5446 19.3944
R16939 gnd.n5446 gnd.n5445 19.3944
R16940 gnd.n5445 gnd.n5368 19.3944
R16941 gnd.n5440 gnd.n5368 19.3944
R16942 gnd.n5440 gnd.n5439 19.3944
R16943 gnd.n5439 gnd.n5438 19.3944
R16944 gnd.n5438 gnd.n5375 19.3944
R16945 gnd.n5433 gnd.n5375 19.3944
R16946 gnd.n5433 gnd.n5432 19.3944
R16947 gnd.n5432 gnd.n5431 19.3944
R16948 gnd.n5431 gnd.n5382 19.3944
R16949 gnd.n5426 gnd.n5382 19.3944
R16950 gnd.n5426 gnd.n5425 19.3944
R16951 gnd.n5425 gnd.n5424 19.3944
R16952 gnd.n5424 gnd.n5389 19.3944
R16953 gnd.n5500 gnd.n1168 19.3944
R16954 gnd.n5500 gnd.n1172 19.3944
R16955 gnd.n1175 gnd.n1172 19.3944
R16956 gnd.n5493 gnd.n1175 19.3944
R16957 gnd.n5493 gnd.n5492 19.3944
R16958 gnd.n5492 gnd.n5491 19.3944
R16959 gnd.n5491 gnd.n1181 19.3944
R16960 gnd.n5486 gnd.n1181 19.3944
R16961 gnd.n5486 gnd.n5485 19.3944
R16962 gnd.n5485 gnd.n5484 19.3944
R16963 gnd.n5484 gnd.n1188 19.3944
R16964 gnd.n5479 gnd.n1188 19.3944
R16965 gnd.n5479 gnd.n5478 19.3944
R16966 gnd.n5478 gnd.n5477 19.3944
R16967 gnd.n5477 gnd.n1195 19.3944
R16968 gnd.n5472 gnd.n1195 19.3944
R16969 gnd.n5472 gnd.n5471 19.3944
R16970 gnd.n5471 gnd.n5470 19.3944
R16971 gnd.n5519 gnd.n1148 19.3944
R16972 gnd.n5519 gnd.n1153 19.3944
R16973 gnd.n1157 gnd.n1153 19.3944
R16974 gnd.n5512 gnd.n1157 19.3944
R16975 gnd.n5512 gnd.n5511 19.3944
R16976 gnd.n5511 gnd.n5510 19.3944
R16977 gnd.n5510 gnd.n1163 19.3944
R16978 gnd.n5505 gnd.n1163 19.3944
R16979 gnd.n5419 gnd.n5418 19.3944
R16980 gnd.n5418 gnd.n5417 19.3944
R16981 gnd.n5417 gnd.n5399 19.3944
R16982 gnd.n5412 gnd.n5399 19.3944
R16983 gnd.n5412 gnd.n5411 19.3944
R16984 gnd.n5411 gnd.n5410 19.3944
R16985 gnd.n5410 gnd.n1149 19.3944
R16986 gnd.n4712 gnd.n1512 19.3944
R16987 gnd.n4712 gnd.n4711 19.3944
R16988 gnd.n4711 gnd.n1487 19.3944
R16989 gnd.n4741 gnd.n1487 19.3944
R16990 gnd.n4741 gnd.n1485 19.3944
R16991 gnd.n4745 gnd.n1485 19.3944
R16992 gnd.n4745 gnd.n1465 19.3944
R16993 gnd.n4768 gnd.n1465 19.3944
R16994 gnd.n4768 gnd.n1463 19.3944
R16995 gnd.n4772 gnd.n1463 19.3944
R16996 gnd.n4772 gnd.n1429 19.3944
R16997 gnd.n4820 gnd.n1429 19.3944
R16998 gnd.n4820 gnd.n1427 19.3944
R16999 gnd.n4824 gnd.n1427 19.3944
R17000 gnd.n4825 gnd.n4824 19.3944
R17001 gnd.n4825 gnd.n1355 19.3944
R17002 gnd.n4923 gnd.n4922 19.3944
R17003 gnd.n4912 gnd.n4911 19.3944
R17004 gnd.n1375 gnd.n1374 19.3944
R17005 gnd.n4898 gnd.n4897 19.3944
R17006 gnd.n1391 gnd.n1348 19.3944
R17007 gnd.n4929 gnd.n1348 19.3944
R17008 gnd.n4929 gnd.n4928 19.3944
R17009 gnd.n4928 gnd.n1317 19.3944
R17010 gnd.n4976 gnd.n1317 19.3944
R17011 gnd.n4976 gnd.n1315 19.3944
R17012 gnd.n4982 gnd.n1315 19.3944
R17013 gnd.n4982 gnd.n4981 19.3944
R17014 gnd.n4981 gnd.n1289 19.3944
R17015 gnd.n5010 gnd.n1289 19.3944
R17016 gnd.n5010 gnd.n1287 19.3944
R17017 gnd.n5014 gnd.n1287 19.3944
R17018 gnd.n5014 gnd.n1220 19.3944
R17019 gnd.n5358 gnd.n1220 19.3944
R17020 gnd.n5358 gnd.n1218 19.3944
R17021 gnd.n5456 gnd.n1218 19.3944
R17022 gnd.n5456 gnd.n5455 19.3944
R17023 gnd.n2745 gnd.n1682 19.3944
R17024 gnd.n2745 gnd.n1678 19.3944
R17025 gnd.n2751 gnd.n1678 19.3944
R17026 gnd.n2751 gnd.n1676 19.3944
R17027 gnd.n2755 gnd.n1676 19.3944
R17028 gnd.n2755 gnd.n1672 19.3944
R17029 gnd.n2761 gnd.n1672 19.3944
R17030 gnd.n2761 gnd.n1670 19.3944
R17031 gnd.n2765 gnd.n1670 19.3944
R17032 gnd.n2765 gnd.n1666 19.3944
R17033 gnd.n2771 gnd.n1666 19.3944
R17034 gnd.n2771 gnd.n1664 19.3944
R17035 gnd.n2775 gnd.n1664 19.3944
R17036 gnd.n2775 gnd.n1660 19.3944
R17037 gnd.n2781 gnd.n1660 19.3944
R17038 gnd.n2781 gnd.n1658 19.3944
R17039 gnd.n2785 gnd.n1658 19.3944
R17040 gnd.n2785 gnd.n1654 19.3944
R17041 gnd.n2791 gnd.n1654 19.3944
R17042 gnd.n2791 gnd.n1652 19.3944
R17043 gnd.n2795 gnd.n1652 19.3944
R17044 gnd.n2795 gnd.n1648 19.3944
R17045 gnd.n2801 gnd.n1648 19.3944
R17046 gnd.n2801 gnd.n1646 19.3944
R17047 gnd.n2805 gnd.n1646 19.3944
R17048 gnd.n2805 gnd.n1642 19.3944
R17049 gnd.n2811 gnd.n1642 19.3944
R17050 gnd.n2811 gnd.n1640 19.3944
R17051 gnd.n2815 gnd.n1640 19.3944
R17052 gnd.n2815 gnd.n1636 19.3944
R17053 gnd.n2821 gnd.n1636 19.3944
R17054 gnd.n2821 gnd.n1634 19.3944
R17055 gnd.n2825 gnd.n1634 19.3944
R17056 gnd.n2825 gnd.n1630 19.3944
R17057 gnd.n2831 gnd.n1630 19.3944
R17058 gnd.n2831 gnd.n1628 19.3944
R17059 gnd.n2835 gnd.n1628 19.3944
R17060 gnd.n2835 gnd.n1624 19.3944
R17061 gnd.n2841 gnd.n1624 19.3944
R17062 gnd.n2841 gnd.n1622 19.3944
R17063 gnd.n2845 gnd.n1622 19.3944
R17064 gnd.n2845 gnd.n1618 19.3944
R17065 gnd.n2851 gnd.n1618 19.3944
R17066 gnd.n2851 gnd.n1616 19.3944
R17067 gnd.n2855 gnd.n1616 19.3944
R17068 gnd.n2855 gnd.n1612 19.3944
R17069 gnd.n2861 gnd.n1612 19.3944
R17070 gnd.n2861 gnd.n1610 19.3944
R17071 gnd.n2865 gnd.n1610 19.3944
R17072 gnd.n2865 gnd.n1606 19.3944
R17073 gnd.n2871 gnd.n1606 19.3944
R17074 gnd.n2871 gnd.n1604 19.3944
R17075 gnd.n2875 gnd.n1604 19.3944
R17076 gnd.n2875 gnd.n1600 19.3944
R17077 gnd.n2881 gnd.n1600 19.3944
R17078 gnd.n2881 gnd.n1598 19.3944
R17079 gnd.n2885 gnd.n1598 19.3944
R17080 gnd.n2885 gnd.n1594 19.3944
R17081 gnd.n2891 gnd.n1594 19.3944
R17082 gnd.n2891 gnd.n1592 19.3944
R17083 gnd.n2895 gnd.n1592 19.3944
R17084 gnd.n2895 gnd.n1588 19.3944
R17085 gnd.n2901 gnd.n1588 19.3944
R17086 gnd.n2901 gnd.n1586 19.3944
R17087 gnd.n2905 gnd.n1586 19.3944
R17088 gnd.n2905 gnd.n1582 19.3944
R17089 gnd.n2911 gnd.n1582 19.3944
R17090 gnd.n2911 gnd.n1580 19.3944
R17091 gnd.n2915 gnd.n1580 19.3944
R17092 gnd.n2915 gnd.n1576 19.3944
R17093 gnd.n2921 gnd.n1576 19.3944
R17094 gnd.n2921 gnd.n1574 19.3944
R17095 gnd.n2925 gnd.n1574 19.3944
R17096 gnd.n2925 gnd.n1570 19.3944
R17097 gnd.n2931 gnd.n1570 19.3944
R17098 gnd.n2931 gnd.n1568 19.3944
R17099 gnd.n2935 gnd.n1568 19.3944
R17100 gnd.n2935 gnd.n1564 19.3944
R17101 gnd.n2941 gnd.n1564 19.3944
R17102 gnd.n2941 gnd.n1562 19.3944
R17103 gnd.n2946 gnd.n1562 19.3944
R17104 gnd.n2946 gnd.n1558 19.3944
R17105 gnd.n4415 gnd.n1558 19.3944
R17106 gnd.n4416 gnd.n4415 19.3944
R17107 gnd.n5170 gnd.n5046 19.3944
R17108 gnd.n5170 gnd.n5047 19.3944
R17109 gnd.n5166 gnd.n5047 19.3944
R17110 gnd.n5166 gnd.n5165 19.3944
R17111 gnd.n5165 gnd.n5164 19.3944
R17112 gnd.n5164 gnd.n5053 19.3944
R17113 gnd.n5160 gnd.n5053 19.3944
R17114 gnd.n5160 gnd.n5159 19.3944
R17115 gnd.n5159 gnd.n5158 19.3944
R17116 gnd.n5158 gnd.n5058 19.3944
R17117 gnd.n5154 gnd.n5058 19.3944
R17118 gnd.n5154 gnd.n1076 19.3944
R17119 gnd.n5621 gnd.n1076 19.3944
R17120 gnd.n5621 gnd.n1074 19.3944
R17121 gnd.n5625 gnd.n1074 19.3944
R17122 gnd.n5625 gnd.n1003 19.3944
R17123 gnd.n5661 gnd.n1003 19.3944
R17124 gnd.n5661 gnd.n1001 19.3944
R17125 gnd.n5665 gnd.n1001 19.3944
R17126 gnd.n5665 gnd.n966 19.3944
R17127 gnd.n5716 gnd.n966 19.3944
R17128 gnd.n5716 gnd.n963 19.3944
R17129 gnd.n5721 gnd.n963 19.3944
R17130 gnd.n5721 gnd.n964 19.3944
R17131 gnd.n964 gnd.n931 19.3944
R17132 gnd.n5758 gnd.n931 19.3944
R17133 gnd.n5758 gnd.n929 19.3944
R17134 gnd.n5762 gnd.n929 19.3944
R17135 gnd.n5762 gnd.n898 19.3944
R17136 gnd.n5800 gnd.n898 19.3944
R17137 gnd.n5800 gnd.n896 19.3944
R17138 gnd.n5804 gnd.n896 19.3944
R17139 gnd.n5804 gnd.n883 19.3944
R17140 gnd.n5844 gnd.n883 19.3944
R17141 gnd.n5844 gnd.n881 19.3944
R17142 gnd.n5848 gnd.n881 19.3944
R17143 gnd.n5848 gnd.n853 19.3944
R17144 gnd.n5893 gnd.n853 19.3944
R17145 gnd.n5893 gnd.n850 19.3944
R17146 gnd.n5898 gnd.n850 19.3944
R17147 gnd.n5898 gnd.n851 19.3944
R17148 gnd.n851 gnd.n817 19.3944
R17149 gnd.n5946 gnd.n817 19.3944
R17150 gnd.n5946 gnd.n815 19.3944
R17151 gnd.n5950 gnd.n815 19.3944
R17152 gnd.n5950 gnd.n792 19.3944
R17153 gnd.n6071 gnd.n792 19.3944
R17154 gnd.n6071 gnd.n790 19.3944
R17155 gnd.n6075 gnd.n790 19.3944
R17156 gnd.n6075 gnd.n769 19.3944
R17157 gnd.n6099 gnd.n769 19.3944
R17158 gnd.n6099 gnd.n766 19.3944
R17159 gnd.n6104 gnd.n766 19.3944
R17160 gnd.n6104 gnd.n767 19.3944
R17161 gnd.n767 gnd.n739 19.3944
R17162 gnd.n6134 gnd.n739 19.3944
R17163 gnd.n6134 gnd.n737 19.3944
R17164 gnd.n6138 gnd.n737 19.3944
R17165 gnd.n6138 gnd.n715 19.3944
R17166 gnd.n6166 gnd.n715 19.3944
R17167 gnd.n6166 gnd.n712 19.3944
R17168 gnd.n6177 gnd.n712 19.3944
R17169 gnd.n6177 gnd.n713 19.3944
R17170 gnd.n6173 gnd.n713 19.3944
R17171 gnd.n6173 gnd.n6172 19.3944
R17172 gnd.n6172 gnd.n643 19.3944
R17173 gnd.n6365 gnd.n643 19.3944
R17174 gnd.n6365 gnd.n640 19.3944
R17175 gnd.n6370 gnd.n640 19.3944
R17176 gnd.n6370 gnd.n641 19.3944
R17177 gnd.n641 gnd.n618 19.3944
R17178 gnd.n6395 gnd.n618 19.3944
R17179 gnd.n6395 gnd.n615 19.3944
R17180 gnd.n6400 gnd.n615 19.3944
R17181 gnd.n6400 gnd.n616 19.3944
R17182 gnd.n616 gnd.n593 19.3944
R17183 gnd.n6425 gnd.n593 19.3944
R17184 gnd.n6425 gnd.n590 19.3944
R17185 gnd.n6430 gnd.n590 19.3944
R17186 gnd.n6430 gnd.n591 19.3944
R17187 gnd.n591 gnd.n569 19.3944
R17188 gnd.n6465 gnd.n569 19.3944
R17189 gnd.n6469 gnd.n567 19.3944
R17190 gnd.n6472 gnd.n6469 19.3944
R17191 gnd.n6475 gnd.n6472 19.3944
R17192 gnd.n6475 gnd.n565 19.3944
R17193 gnd.n6479 gnd.n565 19.3944
R17194 gnd.n6482 gnd.n6479 19.3944
R17195 gnd.n6574 gnd.n6482 19.3944
R17196 gnd.n6574 gnd.n6573 19.3944
R17197 gnd.n6573 gnd.n6572 19.3944
R17198 gnd.n6572 gnd.n6487 19.3944
R17199 gnd.n6565 gnd.n6487 19.3944
R17200 gnd.n6565 gnd.n6564 19.3944
R17201 gnd.n6564 gnd.n6498 19.3944
R17202 gnd.n6557 gnd.n6498 19.3944
R17203 gnd.n6557 gnd.n6556 19.3944
R17204 gnd.n6556 gnd.n6510 19.3944
R17205 gnd.n6549 gnd.n6510 19.3944
R17206 gnd.n6549 gnd.n6548 19.3944
R17207 gnd.n6548 gnd.n6518 19.3944
R17208 gnd.n6541 gnd.n6518 19.3944
R17209 gnd.n6541 gnd.n6540 19.3944
R17210 gnd.n6540 gnd.n6530 19.3944
R17211 gnd.n6530 gnd.n445 19.3944
R17212 gnd.n6702 gnd.n445 19.3944
R17213 gnd.n450 gnd.n424 19.3944
R17214 gnd.n6708 gnd.n424 19.3944
R17215 gnd.n6708 gnd.n6707 19.3944
R17216 gnd.n5656 gnd.n5655 18.8883
R17217 gnd.n6280 gnd.n6279 18.8883
R17218 gnd.n3812 gnd.t292 18.8012
R17219 gnd.n3797 gnd.t311 18.8012
R17220 gnd.n3656 gnd.n3655 18.4825
R17221 gnd.n6641 gnd.n6640 18.4247
R17222 gnd.n5523 gnd.n1149 18.4247
R17223 gnd.n6699 gnd.n6698 18.2308
R17224 gnd.n5271 gnd.n5260 18.2308
R17225 gnd.n239 gnd.n182 18.2308
R17226 gnd.n4549 gnd.n4544 18.2308
R17227 gnd.t293 gnd.n3336 18.1639
R17228 gnd.n3364 gnd.t295 17.5266
R17229 gnd.n3763 gnd.t305 16.8893
R17230 gnd.n5458 gnd.t49 16.8893
R17231 gnd.n6734 gnd.t35 16.8893
R17232 gnd.n6623 gnd.n6620 16.6793
R17233 gnd.n7181 gnd.n7178 16.6793
R17234 gnd.n4634 gnd.n4631 16.6793
R17235 gnd.n5505 gnd.n5504 16.6793
R17236 gnd.n4412 gnd.n4411 16.5706
R17237 gnd.n3591 gnd.t126 16.2519
R17238 gnd.n3291 gnd.t299 16.2519
R17239 gnd.n1086 gnd.n1085 16.0975
R17240 gnd.n691 gnd.n690 16.0975
R17241 gnd.n1088 gnd.n1087 16.0975
R17242 gnd.n6213 gnd.n6212 16.0975
R17243 gnd.n5330 gnd.n1245 15.9333
R17244 gnd.n5330 gnd.n1259 15.9333
R17245 gnd.n5175 gnd.n5174 15.9333
R17246 gnd.n5174 gnd.n5173 15.9333
R17247 gnd.n5173 gnd.n5172 15.9333
R17248 gnd.n5172 gnd.n5044 15.9333
R17249 gnd.n5096 gnd.n5095 15.9333
R17250 gnd.n5096 gnd.n5087 15.9333
R17251 gnd.n5107 gnd.n5087 15.9333
R17252 gnd.n5109 gnd.n5107 15.9333
R17253 gnd.n5109 gnd.n5108 15.9333
R17254 gnd.n5108 gnd.n5081 15.9333
R17255 gnd.n5120 gnd.n5081 15.9333
R17256 gnd.n5120 gnd.n5119 15.9333
R17257 gnd.n5117 gnd.n5075 15.9333
R17258 gnd.n5128 gnd.n5075 15.9333
R17259 gnd.n5130 gnd.n5128 15.9333
R17260 gnd.n5130 gnd.n5129 15.9333
R17261 gnd.n5129 gnd.n5068 15.9333
R17262 gnd.n5141 gnd.n5068 15.9333
R17263 gnd.n5141 gnd.n5140 15.9333
R17264 gnd.n5140 gnd.n5139 15.9333
R17265 gnd.n5152 gnd.n5151 15.9333
R17266 gnd.n5151 gnd.n5061 15.9333
R17267 gnd.n5061 gnd.n1078 15.9333
R17268 gnd.n5619 gnd.n1078 15.9333
R17269 gnd.n5619 gnd.n5618 15.9333
R17270 gnd.n5618 gnd.n1070 15.9333
R17271 gnd.n5628 gnd.n1070 15.9333
R17272 gnd.n5628 gnd.n5627 15.9333
R17273 gnd.n5627 gnd.n1072 15.9333
R17274 gnd.n5649 gnd.n5648 15.9333
R17275 gnd.n5598 gnd.n996 15.9333
R17276 gnd.n5694 gnd.n5693 15.9333
R17277 gnd.n5765 gnd.n5764 15.9333
R17278 gnd.n5798 gnd.n900 15.9333
R17279 gnd.n5806 gnd.n893 15.9333
R17280 gnd.n5782 gnd.n5781 15.9333
R17281 gnd.n5866 gnd.n871 15.9333
R17282 gnd.n5908 gnd.n836 15.9333
R17283 gnd.n5908 gnd.n838 15.9333
R17284 gnd.n6069 gnd.n794 15.9333
R17285 gnd.n6078 gnd.n6077 15.9333
R17286 gnd.n6089 gnd.n6088 15.9333
R17287 gnd.n5976 gnd.n5975 15.9333
R17288 gnd.n5984 gnd.n758 15.9333
R17289 gnd.n6140 gnd.n724 15.9333
R17290 gnd.n6188 gnd.n701 15.9333
R17291 gnd.n6352 gnd.n654 15.9333
R17292 gnd.n6352 gnd.n6351 15.9333
R17293 gnd.n6363 gnd.n645 15.9333
R17294 gnd.n6363 gnd.n6362 15.9333
R17295 gnd.n6362 gnd.n647 15.9333
R17296 gnd.n647 gnd.n636 15.9333
R17297 gnd.n6372 gnd.n636 15.9333
R17298 gnd.n6372 gnd.n637 15.9333
R17299 gnd.n637 gnd.n629 15.9333
R17300 gnd.n6382 gnd.n629 15.9333
R17301 gnd.n6382 gnd.n6381 15.9333
R17302 gnd.n6393 gnd.n620 15.9333
R17303 gnd.n6393 gnd.n6392 15.9333
R17304 gnd.n6392 gnd.n622 15.9333
R17305 gnd.n622 gnd.n611 15.9333
R17306 gnd.n6402 gnd.n611 15.9333
R17307 gnd.n6402 gnd.n612 15.9333
R17308 gnd.n612 gnd.n604 15.9333
R17309 gnd.n6412 gnd.n604 15.9333
R17310 gnd.n6411 gnd.n595 15.9333
R17311 gnd.n6423 gnd.n595 15.9333
R17312 gnd.n6423 gnd.n6422 15.9333
R17313 gnd.n6422 gnd.n597 15.9333
R17314 gnd.n597 gnd.n585 15.9333
R17315 gnd.n6432 gnd.n585 15.9333
R17316 gnd.n6432 gnd.n586 15.9333
R17317 gnd.n588 gnd.n586 15.9333
R17318 gnd.n6442 gnd.n6441 15.9333
R17319 gnd.n6441 gnd.n572 15.9333
R17320 gnd.n6463 gnd.n572 15.9333
R17321 gnd.n6463 gnd.n6462 15.9333
R17322 gnd.n6704 gnd.n427 15.9333
R17323 gnd.n6704 gnd.n442 15.9333
R17324 gnd.n4208 gnd.n4206 15.6674
R17325 gnd.n4176 gnd.n4174 15.6674
R17326 gnd.n4144 gnd.n4142 15.6674
R17327 gnd.n4113 gnd.n4111 15.6674
R17328 gnd.n4081 gnd.n4079 15.6674
R17329 gnd.n4049 gnd.n4047 15.6674
R17330 gnd.n4017 gnd.n4015 15.6674
R17331 gnd.n3986 gnd.n3984 15.6674
R17332 gnd.n3582 gnd.t126 15.6146
R17333 gnd.t113 gnd.n4369 15.6146
R17334 gnd.n4273 gnd.t95 15.6146
R17335 gnd.n5095 gnd.t64 15.6146
R17336 gnd.n588 gnd.t53 15.6146
R17337 gnd.n6580 gnd.n560 15.3217
R17338 gnd.n7136 gnd.n7131 15.3217
R17339 gnd.n4591 gnd.n4513 15.3217
R17340 gnd.n5465 gnd.n1204 15.3217
R17341 gnd.n5648 gnd.t133 15.296
R17342 gnd.n5791 gnd.n909 15.296
R17343 gnd.n5842 gnd.n885 15.296
R17344 gnd.n6050 gnd.n785 15.296
R17345 gnd.n6097 gnd.n771 15.296
R17346 gnd.n6164 gnd.t83 15.296
R17347 gnd.n6197 gnd.n6196 15.0827
R17348 gnd.n1017 gnd.n1012 15.0481
R17349 gnd.n6207 gnd.n6206 15.0481
R17350 gnd.n4404 gnd.t296 14.9773
R17351 gnd.n4519 gnd.t27 14.9773
R17352 gnd.n5139 gnd.t151 14.9773
R17353 gnd.t137 gnd.n620 14.9773
R17354 gnd.n7275 gnd.t31 14.9773
R17355 gnd.t86 gnd.n971 14.6587
R17356 gnd.n5755 gnd.n935 14.6587
R17357 gnd.n6122 gnd.n741 14.6587
R17358 gnd.n6163 gnd.n719 14.6587
R17359 gnd.n4390 gnd.t321 14.34
R17360 gnd.t294 gnd.n2999 14.34
R17361 gnd.n6189 gnd.n698 14.0214
R17362 gnd.n3738 gnd.t319 13.7027
R17363 gnd.n3448 gnd.n3447 13.5763
R17364 gnd.n4329 gnd.n3068 13.5763
R17365 gnd.n3656 gnd.n3394 13.384
R17366 gnd.n5674 gnd.n991 13.384
R17367 gnd.n949 gnd.n927 13.384
R17368 gnd.n5884 gnd.n862 13.384
R17369 gnd.n5883 gnd.t1 13.384
R17370 gnd.t14 gnd.n845 13.384
R17371 gnd.n5923 gnd.t9 13.384
R17372 gnd.n5952 gnd.t169 13.384
R17373 gnd.n813 gnd.n802 13.384
R17374 gnd.n6114 gnd.n6113 13.384
R17375 gnd.n6001 gnd.n709 13.384
R17376 gnd.n1028 gnd.n1009 13.1884
R17377 gnd.n1023 gnd.n1022 13.1884
R17378 gnd.n1022 gnd.n1021 13.1884
R17379 gnd.n6200 gnd.n6195 13.1884
R17380 gnd.n6201 gnd.n6200 13.1884
R17381 gnd.n1024 gnd.n1011 13.146
R17382 gnd.n1020 gnd.n1011 13.146
R17383 gnd.n6199 gnd.n6198 13.146
R17384 gnd.n6199 gnd.n6194 13.146
R17385 gnd.n4209 gnd.n4205 12.8005
R17386 gnd.n4177 gnd.n4173 12.8005
R17387 gnd.n4145 gnd.n4141 12.8005
R17388 gnd.n4114 gnd.n4110 12.8005
R17389 gnd.n4082 gnd.n4078 12.8005
R17390 gnd.n4050 gnd.n4046 12.8005
R17391 gnd.n4018 gnd.n4014 12.8005
R17392 gnd.n3987 gnd.n3983 12.8005
R17393 gnd.n5650 gnd.t139 12.7467
R17394 gnd.n5714 gnd.n968 12.7467
R17395 gnd.n5749 gnd.n941 12.7467
R17396 gnd.n5891 gnd.n855 12.7467
R17397 gnd.n5937 gnd.n824 12.7467
R17398 gnd.n5985 gnd.n749 12.7467
R17399 gnd.n3447 gnd.n3442 12.4126
R17400 gnd.n4334 gnd.n3068 12.4126
R17401 gnd.n5655 gnd.n5654 12.1761
R17402 gnd.n6279 gnd.n6278 12.1761
R17403 gnd.n5597 gnd.n1007 12.1094
R17404 gnd.n5705 gnd.t17 12.1094
R17405 gnd.n5797 gnd.n903 12.1094
R17406 gnd.n5858 gnd.n5857 12.1094
R17407 gnd.n6068 gnd.n797 12.1094
R17408 gnd.n5977 gnd.n5974 12.1094
R17409 gnd.n700 gnd.t130 12.1094
R17410 gnd.n4213 gnd.n4212 12.0247
R17411 gnd.n4181 gnd.n4180 12.0247
R17412 gnd.n4149 gnd.n4148 12.0247
R17413 gnd.n4118 gnd.n4117 12.0247
R17414 gnd.n4086 gnd.n4085 12.0247
R17415 gnd.n4054 gnd.n4053 12.0247
R17416 gnd.n4022 gnd.n4021 12.0247
R17417 gnd.n3991 gnd.n3990 12.0247
R17418 gnd.t185 gnd.n1284 11.7908
R17419 gnd.n6803 gnd.t192 11.7908
R17420 gnd.n5183 gnd.n1156 11.4721
R17421 gnd.t68 gnd.n5667 11.4721
R17422 gnd.n5723 gnd.n959 11.4721
R17423 gnd.t4 gnd.n5704 11.4721
R17424 gnd.n5683 gnd.n5681 11.4721
R17425 gnd.n5901 gnd.n5900 11.4721
R17426 gnd.n5922 gnd.n832 11.4721
R17427 gnd.n6130 gnd.n744 11.4721
R17428 gnd.n6141 gnd.t156 11.4721
R17429 gnd.n6151 gnd.n6150 11.4721
R17430 gnd.n6693 gnd.n457 11.4721
R17431 gnd.n4216 gnd.n4203 11.249
R17432 gnd.n4184 gnd.n4171 11.249
R17433 gnd.n4152 gnd.n4139 11.249
R17434 gnd.n4121 gnd.n4108 11.249
R17435 gnd.n4089 gnd.n4076 11.249
R17436 gnd.n4057 gnd.n4044 11.249
R17437 gnd.n4025 gnd.n4012 11.249
R17438 gnd.n3994 gnd.n3981 11.249
R17439 gnd.n3726 gnd.t319 11.1535
R17440 gnd.n4800 gnd.t207 11.1535
R17441 gnd.t179 gnd.n1334 11.1535
R17442 gnd.n5119 gnd.t313 11.1535
R17443 gnd.t317 gnd.n6411 11.1535
R17444 gnd.n6831 gnd.t203 11.1535
R17445 gnd.n6938 gnd.t238 11.1535
R17446 gnd.n4584 gnd.n1506 10.8348
R17447 gnd.n4714 gnd.n1508 10.8348
R17448 gnd.n4519 gnd.n1500 10.8348
R17449 gnd.n4728 gnd.n1489 10.8348
R17450 gnd.n4739 gnd.n1492 10.8348
R17451 gnd.n4722 gnd.n1481 10.8348
R17452 gnd.n4747 gnd.n1482 10.8348
R17453 gnd.n4750 gnd.n1467 10.8348
R17454 gnd.n4766 gnd.n1470 10.8348
R17455 gnd.n4774 gnd.n1449 10.8348
R17456 gnd.n4800 gnd.n4799 10.8348
R17457 gnd.n4818 gnd.n1434 10.8348
R17458 gnd.n4793 gnd.n1442 10.8348
R17459 gnd.n4812 gnd.n4811 10.8348
R17460 gnd.n4827 gnd.n1423 10.8348
R17461 gnd.n4854 gnd.n1415 10.8348
R17462 gnd.n4920 gnd.n1361 10.8348
R17463 gnd.n4864 gnd.n4863 10.8348
R17464 gnd.n4914 gnd.n1372 10.8348
R17465 gnd.n4909 gnd.n4908 10.8348
R17466 gnd.n4901 gnd.n1385 10.8348
R17467 gnd.n4900 gnd.n1388 10.8348
R17468 gnd.n4895 gnd.n1400 10.8348
R17469 gnd.n4881 gnd.n1342 10.8348
R17470 gnd.n4931 gnd.n1344 10.8348
R17471 gnd.n4941 gnd.n1334 10.8348
R17472 gnd.n4940 gnd.n1319 10.8348
R17473 gnd.n4961 gnd.n1309 10.8348
R17474 gnd.n4984 gnd.n1311 10.8348
R17475 gnd.n4967 gnd.n1302 10.8348
R17476 gnd.n4996 gnd.n1291 10.8348
R17477 gnd.n5008 gnd.n1294 10.8348
R17478 gnd.n5017 gnd.n1284 10.8348
R17479 gnd.n5016 gnd.n1232 10.8348
R17480 gnd.n5346 gnd.n1222 10.8348
R17481 gnd.n5356 gnd.n1225 10.8348
R17482 gnd.n5027 gnd.n5026 10.8348
R17483 gnd.n5458 gnd.n1214 10.8348
R17484 gnd.n5190 gnd.n5189 10.8348
R17485 gnd.n5785 gnd.n916 10.8348
R17486 gnd.n788 gnd.n787 10.8348
R17487 gnd.n6716 gnd.n6715 10.8348
R17488 gnd.n6734 gnd.n392 10.8348
R17489 gnd.n6727 gnd.n6726 10.8348
R17490 gnd.n6744 gnd.n382 10.8348
R17491 gnd.n384 gnd.n374 10.8348
R17492 gnd.n6754 gnd.n6753 10.8348
R17493 gnd.n6803 gnd.n359 10.8348
R17494 gnd.n6790 gnd.n6789 10.8348
R17495 gnd.n6813 gnd.n349 10.8348
R17496 gnd.n6796 gnd.n351 10.8348
R17497 gnd.n6822 gnd.n342 10.8348
R17498 gnd.n6838 gnd.n330 10.8348
R17499 gnd.n6849 gnd.n320 10.8348
R17500 gnd.n6831 gnd.n322 10.8348
R17501 gnd.n6865 gnd.n313 10.8348
R17502 gnd.n6872 gnd.n306 10.8348
R17503 gnd.n6877 gnd.n302 10.8348
R17504 gnd.n6886 gnd.n6885 10.8348
R17505 gnd.n6902 gnd.n288 10.8348
R17506 gnd.n6907 gnd.n286 10.8348
R17507 gnd.n6921 gnd.n278 10.8348
R17508 gnd.n7325 gnd.n69 10.8348
R17509 gnd.n265 gnd.n71 10.8348
R17510 gnd.n7317 gnd.n86 10.8348
R17511 gnd.n6991 gnd.n89 10.8348
R17512 gnd.n7311 gnd.n98 10.8348
R17513 gnd.n6985 gnd.n101 10.8348
R17514 gnd.n7305 gnd.n108 10.8348
R17515 gnd.n6979 gnd.n6938 10.8348
R17516 gnd.n7299 gnd.n117 10.8348
R17517 gnd.n7293 gnd.n128 10.8348
R17518 gnd.n6967 gnd.n131 10.8348
R17519 gnd.n7287 gnd.n138 10.8348
R17520 gnd.n6961 gnd.n141 10.8348
R17521 gnd.n7281 gnd.n149 10.8348
R17522 gnd.n6955 gnd.n152 10.8348
R17523 gnd.n7275 gnd.n159 10.8348
R17524 gnd.n7262 gnd.n176 10.8348
R17525 gnd.n7269 gnd.n168 10.8348
R17526 gnd.n6583 gnd.n6580 10.6672
R17527 gnd.n7139 gnd.n7136 10.6672
R17528 gnd.n4594 gnd.n4591 10.6672
R17529 gnd.n5470 gnd.n1204 10.6672
R17530 gnd.n6347 gnd.n6346 10.6151
R17531 gnd.n6346 gnd.n6343 10.6151
R17532 gnd.n6341 gnd.n6338 10.6151
R17533 gnd.n6338 gnd.n6337 10.6151
R17534 gnd.n6337 gnd.n6334 10.6151
R17535 gnd.n6334 gnd.n6333 10.6151
R17536 gnd.n6333 gnd.n6330 10.6151
R17537 gnd.n6330 gnd.n6329 10.6151
R17538 gnd.n6329 gnd.n6326 10.6151
R17539 gnd.n6326 gnd.n6325 10.6151
R17540 gnd.n6325 gnd.n6322 10.6151
R17541 gnd.n6322 gnd.n6321 10.6151
R17542 gnd.n6321 gnd.n6318 10.6151
R17543 gnd.n6318 gnd.n6317 10.6151
R17544 gnd.n6317 gnd.n6314 10.6151
R17545 gnd.n6314 gnd.n6313 10.6151
R17546 gnd.n6313 gnd.n6310 10.6151
R17547 gnd.n6310 gnd.n6309 10.6151
R17548 gnd.n6309 gnd.n6306 10.6151
R17549 gnd.n6306 gnd.n6305 10.6151
R17550 gnd.n6305 gnd.n6302 10.6151
R17551 gnd.n6302 gnd.n6301 10.6151
R17552 gnd.n6301 gnd.n6298 10.6151
R17553 gnd.n6298 gnd.n6297 10.6151
R17554 gnd.n6297 gnd.n6294 10.6151
R17555 gnd.n6294 gnd.n6293 10.6151
R17556 gnd.n6293 gnd.n6290 10.6151
R17557 gnd.n6290 gnd.n6289 10.6151
R17558 gnd.n6289 gnd.n6286 10.6151
R17559 gnd.n6286 gnd.n6285 10.6151
R17560 gnd.n5595 gnd.n5592 10.6151
R17561 gnd.n5595 gnd.n5594 10.6151
R17562 gnd.n5594 gnd.n5593 10.6151
R17563 gnd.n5593 gnd.n989 10.6151
R17564 gnd.n5677 gnd.n989 10.6151
R17565 gnd.n5678 gnd.n5677 10.6151
R17566 gnd.n5691 gnd.n5678 10.6151
R17567 gnd.n5691 gnd.n5690 10.6151
R17568 gnd.n5690 gnd.n5689 10.6151
R17569 gnd.n5689 gnd.n5687 10.6151
R17570 gnd.n5687 gnd.n5686 10.6151
R17571 gnd.n5686 gnd.n5680 10.6151
R17572 gnd.n5680 gnd.n5679 10.6151
R17573 gnd.n5679 gnd.n945 10.6151
R17574 gnd.n5747 gnd.n945 10.6151
R17575 gnd.n5747 gnd.n5746 10.6151
R17576 gnd.n5746 gnd.n5745 10.6151
R17577 gnd.n5745 gnd.n947 10.6151
R17578 gnd.n947 gnd.n946 10.6151
R17579 gnd.n946 gnd.n913 10.6151
R17580 gnd.n5789 gnd.n913 10.6151
R17581 gnd.n5789 gnd.n5788 10.6151
R17582 gnd.n5788 gnd.n5787 10.6151
R17583 gnd.n5787 gnd.n914 10.6151
R17584 gnd.n914 gnd.n877 10.6151
R17585 gnd.n5855 gnd.n877 10.6151
R17586 gnd.n5855 gnd.n5854 10.6151
R17587 gnd.n5854 gnd.n5853 10.6151
R17588 gnd.n5853 gnd.n878 10.6151
R17589 gnd.n5813 gnd.n878 10.6151
R17590 gnd.n5814 gnd.n5813 10.6151
R17591 gnd.n5816 gnd.n5814 10.6151
R17592 gnd.n5816 gnd.n5815 10.6151
R17593 gnd.n5815 gnd.n834 10.6151
R17594 gnd.n5910 gnd.n834 10.6151
R17595 gnd.n5911 gnd.n5910 10.6151
R17596 gnd.n5920 gnd.n5911 10.6151
R17597 gnd.n5920 gnd.n5919 10.6151
R17598 gnd.n5919 gnd.n5918 10.6151
R17599 gnd.n5918 gnd.n5914 10.6151
R17600 gnd.n5914 gnd.n5913 10.6151
R17601 gnd.n5913 gnd.n805 10.6151
R17602 gnd.n6055 gnd.n805 10.6151
R17603 gnd.n6055 gnd.n6054 10.6151
R17604 gnd.n6054 gnd.n6053 10.6151
R17605 gnd.n6053 gnd.n806 10.6151
R17606 gnd.n5969 gnd.n806 10.6151
R17607 gnd.n5970 gnd.n5969 10.6151
R17608 gnd.n5972 gnd.n5970 10.6151
R17609 gnd.n5973 gnd.n5972 10.6151
R17610 gnd.n5979 gnd.n5973 10.6151
R17611 gnd.n5980 gnd.n5979 10.6151
R17612 gnd.n5982 gnd.n5980 10.6151
R17613 gnd.n5983 gnd.n5982 10.6151
R17614 gnd.n5987 gnd.n5983 10.6151
R17615 gnd.n5988 gnd.n5987 10.6151
R17616 gnd.n5990 gnd.n5988 10.6151
R17617 gnd.n5991 gnd.n5990 10.6151
R17618 gnd.n5993 gnd.n5991 10.6151
R17619 gnd.n5994 gnd.n5993 10.6151
R17620 gnd.n5995 gnd.n5994 10.6151
R17621 gnd.n5996 gnd.n5995 10.6151
R17622 gnd.n5997 gnd.n5996 10.6151
R17623 gnd.n6007 gnd.n5997 10.6151
R17624 gnd.n6007 gnd.n6006 10.6151
R17625 gnd.n6006 gnd.n6005 10.6151
R17626 gnd.n6005 gnd.n6000 10.6151
R17627 gnd.n6000 gnd.n5999 10.6151
R17628 gnd.n5999 gnd.n5998 10.6151
R17629 gnd.n5998 gnd.n692 10.6151
R17630 gnd.n5529 gnd.n5528 10.6151
R17631 gnd.n5532 gnd.n5529 10.6151
R17632 gnd.n5537 gnd.n5534 10.6151
R17633 gnd.n5538 gnd.n5537 10.6151
R17634 gnd.n5541 gnd.n5538 10.6151
R17635 gnd.n5542 gnd.n5541 10.6151
R17636 gnd.n5545 gnd.n5542 10.6151
R17637 gnd.n5546 gnd.n5545 10.6151
R17638 gnd.n5549 gnd.n5546 10.6151
R17639 gnd.n5550 gnd.n5549 10.6151
R17640 gnd.n5553 gnd.n5550 10.6151
R17641 gnd.n5554 gnd.n5553 10.6151
R17642 gnd.n5557 gnd.n5554 10.6151
R17643 gnd.n5558 gnd.n5557 10.6151
R17644 gnd.n5561 gnd.n5558 10.6151
R17645 gnd.n5562 gnd.n5561 10.6151
R17646 gnd.n5565 gnd.n5562 10.6151
R17647 gnd.n5566 gnd.n5565 10.6151
R17648 gnd.n5569 gnd.n5566 10.6151
R17649 gnd.n5570 gnd.n5569 10.6151
R17650 gnd.n5573 gnd.n5570 10.6151
R17651 gnd.n5574 gnd.n5573 10.6151
R17652 gnd.n5577 gnd.n5574 10.6151
R17653 gnd.n5578 gnd.n5577 10.6151
R17654 gnd.n5581 gnd.n5578 10.6151
R17655 gnd.n5582 gnd.n5581 10.6151
R17656 gnd.n5585 gnd.n5582 10.6151
R17657 gnd.n5586 gnd.n5585 10.6151
R17658 gnd.n5589 gnd.n5586 10.6151
R17659 gnd.n5591 gnd.n5589 10.6151
R17660 gnd.n5654 gnd.n5653 10.6151
R17661 gnd.n5653 gnd.n1029 10.6151
R17662 gnd.n1091 gnd.n1029 10.6151
R17663 gnd.n1092 gnd.n1091 10.6151
R17664 gnd.n1095 gnd.n1092 10.6151
R17665 gnd.n1096 gnd.n1095 10.6151
R17666 gnd.n1099 gnd.n1096 10.6151
R17667 gnd.n1100 gnd.n1099 10.6151
R17668 gnd.n1103 gnd.n1100 10.6151
R17669 gnd.n1104 gnd.n1103 10.6151
R17670 gnd.n1107 gnd.n1104 10.6151
R17671 gnd.n1108 gnd.n1107 10.6151
R17672 gnd.n1111 gnd.n1108 10.6151
R17673 gnd.n1112 gnd.n1111 10.6151
R17674 gnd.n1115 gnd.n1112 10.6151
R17675 gnd.n1116 gnd.n1115 10.6151
R17676 gnd.n1119 gnd.n1116 10.6151
R17677 gnd.n1120 gnd.n1119 10.6151
R17678 gnd.n1123 gnd.n1120 10.6151
R17679 gnd.n1124 gnd.n1123 10.6151
R17680 gnd.n1127 gnd.n1124 10.6151
R17681 gnd.n1128 gnd.n1127 10.6151
R17682 gnd.n1131 gnd.n1128 10.6151
R17683 gnd.n1132 gnd.n1131 10.6151
R17684 gnd.n1135 gnd.n1132 10.6151
R17685 gnd.n1136 gnd.n1135 10.6151
R17686 gnd.n1139 gnd.n1136 10.6151
R17687 gnd.n1140 gnd.n1139 10.6151
R17688 gnd.n1144 gnd.n1143 10.6151
R17689 gnd.n1147 gnd.n1144 10.6151
R17690 gnd.n6278 gnd.n6277 10.6151
R17691 gnd.n6277 gnd.n6274 10.6151
R17692 gnd.n6274 gnd.n6273 10.6151
R17693 gnd.n6273 gnd.n6270 10.6151
R17694 gnd.n6270 gnd.n6269 10.6151
R17695 gnd.n6269 gnd.n6266 10.6151
R17696 gnd.n6266 gnd.n6265 10.6151
R17697 gnd.n6265 gnd.n6262 10.6151
R17698 gnd.n6262 gnd.n6261 10.6151
R17699 gnd.n6261 gnd.n6258 10.6151
R17700 gnd.n6258 gnd.n6257 10.6151
R17701 gnd.n6257 gnd.n6254 10.6151
R17702 gnd.n6254 gnd.n6253 10.6151
R17703 gnd.n6253 gnd.n6250 10.6151
R17704 gnd.n6250 gnd.n6249 10.6151
R17705 gnd.n6249 gnd.n6246 10.6151
R17706 gnd.n6246 gnd.n6245 10.6151
R17707 gnd.n6245 gnd.n6242 10.6151
R17708 gnd.n6242 gnd.n6241 10.6151
R17709 gnd.n6241 gnd.n6238 10.6151
R17710 gnd.n6238 gnd.n6237 10.6151
R17711 gnd.n6237 gnd.n6234 10.6151
R17712 gnd.n6234 gnd.n6233 10.6151
R17713 gnd.n6233 gnd.n6230 10.6151
R17714 gnd.n6230 gnd.n6229 10.6151
R17715 gnd.n6229 gnd.n6226 10.6151
R17716 gnd.n6226 gnd.n6225 10.6151
R17717 gnd.n6225 gnd.n6222 10.6151
R17718 gnd.n6220 gnd.n6217 10.6151
R17719 gnd.n6217 gnd.n6216 10.6151
R17720 gnd.n5656 gnd.n994 10.6151
R17721 gnd.n5670 gnd.n994 10.6151
R17722 gnd.n5671 gnd.n5670 10.6151
R17723 gnd.n5672 gnd.n5671 10.6151
R17724 gnd.n5672 gnd.n974 10.6151
R17725 gnd.n5711 gnd.n974 10.6151
R17726 gnd.n5711 gnd.n5710 10.6151
R17727 gnd.n5710 gnd.n5709 10.6151
R17728 gnd.n5709 gnd.n975 10.6151
R17729 gnd.n978 gnd.n975 10.6151
R17730 gnd.n978 gnd.n977 10.6151
R17731 gnd.n977 gnd.n938 10.6151
R17732 gnd.n5753 gnd.n938 10.6151
R17733 gnd.n5753 gnd.n5752 10.6151
R17734 gnd.n5752 gnd.n5751 10.6151
R17735 gnd.n5751 gnd.n939 10.6151
R17736 gnd.n5741 gnd.n939 10.6151
R17737 gnd.n5741 gnd.n906 10.6151
R17738 gnd.n5795 gnd.n906 10.6151
R17739 gnd.n5795 gnd.n5794 10.6151
R17740 gnd.n5794 gnd.n5793 10.6151
R17741 gnd.n5793 gnd.n907 10.6151
R17742 gnd.n5783 gnd.n907 10.6151
R17743 gnd.n5783 gnd.n874 10.6151
R17744 gnd.n5861 gnd.n874 10.6151
R17745 gnd.n5862 gnd.n5861 10.6151
R17746 gnd.n5863 gnd.n5862 10.6151
R17747 gnd.n5863 gnd.n860 10.6151
R17748 gnd.n5886 gnd.n860 10.6151
R17749 gnd.n5887 gnd.n5886 10.6151
R17750 gnd.n5888 gnd.n5887 10.6151
R17751 gnd.n5888 gnd.n843 10.6151
R17752 gnd.n5903 gnd.n843 10.6151
R17753 gnd.n5904 gnd.n5903 10.6151
R17754 gnd.n5906 gnd.n5904 10.6151
R17755 gnd.n5906 gnd.n5905 10.6151
R17756 gnd.n5905 gnd.n823 10.6151
R17757 gnd.n5941 gnd.n823 10.6151
R17758 gnd.n5941 gnd.n5940 10.6151
R17759 gnd.n5940 gnd.n5939 10.6151
R17760 gnd.n5939 gnd.n800 10.6151
R17761 gnd.n6061 gnd.n800 10.6151
R17762 gnd.n6062 gnd.n6061 10.6151
R17763 gnd.n6066 gnd.n6062 10.6151
R17764 gnd.n6066 gnd.n6065 10.6151
R17765 gnd.n6065 gnd.n6064 10.6151
R17766 gnd.n6064 gnd.n775 10.6151
R17767 gnd.n6092 gnd.n775 10.6151
R17768 gnd.n6093 gnd.n6092 10.6151
R17769 gnd.n6094 gnd.n6093 10.6151
R17770 gnd.n6094 gnd.n760 10.6151
R17771 gnd.n6109 gnd.n760 10.6151
R17772 gnd.n6110 gnd.n6109 10.6151
R17773 gnd.n6111 gnd.n6110 10.6151
R17774 gnd.n6111 gnd.n747 10.6151
R17775 gnd.n6125 gnd.n747 10.6151
R17776 gnd.n6126 gnd.n6125 10.6151
R17777 gnd.n6128 gnd.n6126 10.6151
R17778 gnd.n6128 gnd.n6127 10.6151
R17779 gnd.n6127 gnd.n722 10.6151
R17780 gnd.n6154 gnd.n722 10.6151
R17781 gnd.n6155 gnd.n6154 10.6151
R17782 gnd.n6161 gnd.n6155 10.6151
R17783 gnd.n6161 gnd.n6160 10.6151
R17784 gnd.n6160 gnd.n6159 10.6151
R17785 gnd.n6159 gnd.n6156 10.6151
R17786 gnd.n6156 gnd.n696 10.6151
R17787 gnd.n6191 gnd.n696 10.6151
R17788 gnd.n6192 gnd.n6191 10.6151
R17789 gnd.n6280 gnd.n6192 10.6151
R17790 gnd.n3645 gnd.t165 10.5161
R17791 gnd.n4255 gnd.t321 10.5161
R17792 gnd.n4262 gnd.t294 10.5161
R17793 gnd.t200 gnd.n1358 10.5161
R17794 gnd.n4863 gnd.t242 10.5161
R17795 gnd.n4914 gnd.t242 10.5161
R17796 gnd.t231 gnd.n1378 10.5161
R17797 gnd.n6912 gnd.t197 10.5161
R17798 gnd.n6921 gnd.t222 10.5161
R17799 gnd.t222 gnd.n69 10.5161
R17800 gnd.n6998 gnd.t172 10.5161
R17801 gnd.n4217 gnd.n4201 10.4732
R17802 gnd.n4185 gnd.n4169 10.4732
R17803 gnd.n4153 gnd.n4137 10.4732
R17804 gnd.n4122 gnd.n4106 10.4732
R17805 gnd.n4090 gnd.n4074 10.4732
R17806 gnd.n4058 gnd.n4042 10.4732
R17807 gnd.n4026 gnd.n4010 10.4732
R17808 gnd.n3995 gnd.n3979 10.4732
R17809 gnd.n5723 gnd.n960 10.1975
R17810 gnd.t143 gnd.n5739 10.1975
R17811 gnd.n5900 gnd.n848 10.1975
R17812 gnd.n841 gnd.n832 10.1975
R17813 gnd.n6107 gnd.t308 10.1975
R17814 gnd.n6152 gnd.n6151 10.1975
R17815 gnd.n3930 gnd.t296 9.87883
R17816 gnd.t218 gnd.n1460 9.87883
R17817 gnd.n4818 gnd.t207 9.87883
R17818 gnd.n1344 gnd.t179 9.87883
R17819 gnd.n4974 gnd.t211 9.87883
R17820 gnd.n6826 gnd.t183 9.87883
R17821 gnd.t203 gnd.n313 9.87883
R17822 gnd.n7305 gnd.t238 9.87883
R17823 gnd.t176 gnd.n120 9.87883
R17824 gnd.n4221 gnd.n4220 9.69747
R17825 gnd.n4189 gnd.n4188 9.69747
R17826 gnd.n4157 gnd.n4156 9.69747
R17827 gnd.n4126 gnd.n4125 9.69747
R17828 gnd.n4094 gnd.n4093 9.69747
R17829 gnd.n4062 gnd.n4061 9.69747
R17830 gnd.n4030 gnd.n4029 9.69747
R17831 gnd.n3999 gnd.n3998 9.69747
R17832 gnd.n5658 gnd.n1007 9.56018
R17833 gnd.n5682 gnd.t141 9.56018
R17834 gnd.n5859 gnd.n5858 9.56018
R17835 gnd.n6051 gnd.n797 9.56018
R17836 gnd.t12 gnd.n6131 9.56018
R17837 gnd.n6282 gnd.t130 9.56018
R17838 gnd.n4227 gnd.n4226 9.45567
R17839 gnd.n4195 gnd.n4194 9.45567
R17840 gnd.n4163 gnd.n4162 9.45567
R17841 gnd.n4132 gnd.n4131 9.45567
R17842 gnd.n4100 gnd.n4099 9.45567
R17843 gnd.n4068 gnd.n4067 9.45567
R17844 gnd.n4036 gnd.n4035 9.45567
R17845 gnd.n4005 gnd.n4004 9.45567
R17846 gnd.n6620 gnd.n6619 9.30959
R17847 gnd.n7178 gnd.n7110 9.30959
R17848 gnd.n4631 gnd.n4630 9.30959
R17849 gnd.n5504 gnd.n1168 9.30959
R17850 gnd.n4226 gnd.n4225 9.3005
R17851 gnd.n4199 gnd.n4198 9.3005
R17852 gnd.n4220 gnd.n4219 9.3005
R17853 gnd.n4218 gnd.n4217 9.3005
R17854 gnd.n4203 gnd.n4202 9.3005
R17855 gnd.n4212 gnd.n4211 9.3005
R17856 gnd.n4210 gnd.n4209 9.3005
R17857 gnd.n4194 gnd.n4193 9.3005
R17858 gnd.n4167 gnd.n4166 9.3005
R17859 gnd.n4188 gnd.n4187 9.3005
R17860 gnd.n4186 gnd.n4185 9.3005
R17861 gnd.n4171 gnd.n4170 9.3005
R17862 gnd.n4180 gnd.n4179 9.3005
R17863 gnd.n4178 gnd.n4177 9.3005
R17864 gnd.n4162 gnd.n4161 9.3005
R17865 gnd.n4135 gnd.n4134 9.3005
R17866 gnd.n4156 gnd.n4155 9.3005
R17867 gnd.n4154 gnd.n4153 9.3005
R17868 gnd.n4139 gnd.n4138 9.3005
R17869 gnd.n4148 gnd.n4147 9.3005
R17870 gnd.n4146 gnd.n4145 9.3005
R17871 gnd.n4131 gnd.n4130 9.3005
R17872 gnd.n4104 gnd.n4103 9.3005
R17873 gnd.n4125 gnd.n4124 9.3005
R17874 gnd.n4123 gnd.n4122 9.3005
R17875 gnd.n4108 gnd.n4107 9.3005
R17876 gnd.n4117 gnd.n4116 9.3005
R17877 gnd.n4115 gnd.n4114 9.3005
R17878 gnd.n4099 gnd.n4098 9.3005
R17879 gnd.n4072 gnd.n4071 9.3005
R17880 gnd.n4093 gnd.n4092 9.3005
R17881 gnd.n4091 gnd.n4090 9.3005
R17882 gnd.n4076 gnd.n4075 9.3005
R17883 gnd.n4085 gnd.n4084 9.3005
R17884 gnd.n4083 gnd.n4082 9.3005
R17885 gnd.n4067 gnd.n4066 9.3005
R17886 gnd.n4040 gnd.n4039 9.3005
R17887 gnd.n4061 gnd.n4060 9.3005
R17888 gnd.n4059 gnd.n4058 9.3005
R17889 gnd.n4044 gnd.n4043 9.3005
R17890 gnd.n4053 gnd.n4052 9.3005
R17891 gnd.n4051 gnd.n4050 9.3005
R17892 gnd.n4035 gnd.n4034 9.3005
R17893 gnd.n4008 gnd.n4007 9.3005
R17894 gnd.n4029 gnd.n4028 9.3005
R17895 gnd.n4027 gnd.n4026 9.3005
R17896 gnd.n4012 gnd.n4011 9.3005
R17897 gnd.n4021 gnd.n4020 9.3005
R17898 gnd.n4019 gnd.n4018 9.3005
R17899 gnd.n4004 gnd.n4003 9.3005
R17900 gnd.n3977 gnd.n3976 9.3005
R17901 gnd.n3998 gnd.n3997 9.3005
R17902 gnd.n3996 gnd.n3995 9.3005
R17903 gnd.n3981 gnd.n3980 9.3005
R17904 gnd.n3990 gnd.n3989 9.3005
R17905 gnd.n3988 gnd.n3987 9.3005
R17906 gnd.n4356 gnd.n3042 9.3005
R17907 gnd.n4355 gnd.n3044 9.3005
R17908 gnd.n3048 gnd.n3045 9.3005
R17909 gnd.n4350 gnd.n3049 9.3005
R17910 gnd.n4349 gnd.n3050 9.3005
R17911 gnd.n4348 gnd.n3051 9.3005
R17912 gnd.n3055 gnd.n3052 9.3005
R17913 gnd.n4343 gnd.n3056 9.3005
R17914 gnd.n4342 gnd.n3057 9.3005
R17915 gnd.n4341 gnd.n3058 9.3005
R17916 gnd.n3062 gnd.n3059 9.3005
R17917 gnd.n4336 gnd.n3063 9.3005
R17918 gnd.n4335 gnd.n3064 9.3005
R17919 gnd.n4334 gnd.n3065 9.3005
R17920 gnd.n3070 gnd.n3068 9.3005
R17921 gnd.n4329 gnd.n4328 9.3005
R17922 gnd.n4358 gnd.n4357 9.3005
R17923 gnd.n3664 gnd.n3663 9.3005
R17924 gnd.n3368 gnd.n3367 9.3005
R17925 gnd.n3691 gnd.n3690 9.3005
R17926 gnd.n3692 gnd.n3366 9.3005
R17927 gnd.n3696 gnd.n3693 9.3005
R17928 gnd.n3695 gnd.n3694 9.3005
R17929 gnd.n3340 gnd.n3339 9.3005
R17930 gnd.n3721 gnd.n3720 9.3005
R17931 gnd.n3722 gnd.n3338 9.3005
R17932 gnd.n3724 gnd.n3723 9.3005
R17933 gnd.n3318 gnd.n3317 9.3005
R17934 gnd.n3752 gnd.n3751 9.3005
R17935 gnd.n3753 gnd.n3316 9.3005
R17936 gnd.n3761 gnd.n3754 9.3005
R17937 gnd.n3760 gnd.n3755 9.3005
R17938 gnd.n3759 gnd.n3757 9.3005
R17939 gnd.n3756 gnd.n3265 9.3005
R17940 gnd.n3809 gnd.n3266 9.3005
R17941 gnd.n3808 gnd.n3267 9.3005
R17942 gnd.n3807 gnd.n3268 9.3005
R17943 gnd.n3287 gnd.n3269 9.3005
R17944 gnd.n3289 gnd.n3288 9.3005
R17945 gnd.n3187 gnd.n3186 9.3005
R17946 gnd.n3847 gnd.n3846 9.3005
R17947 gnd.n3848 gnd.n3185 9.3005
R17948 gnd.n3852 gnd.n3849 9.3005
R17949 gnd.n3851 gnd.n3850 9.3005
R17950 gnd.n3160 gnd.n3159 9.3005
R17951 gnd.n3887 gnd.n3886 9.3005
R17952 gnd.n3888 gnd.n3158 9.3005
R17953 gnd.n3892 gnd.n3889 9.3005
R17954 gnd.n3891 gnd.n3890 9.3005
R17955 gnd.n3134 gnd.n3133 9.3005
R17956 gnd.n3943 gnd.n3942 9.3005
R17957 gnd.n3944 gnd.n3132 9.3005
R17958 gnd.n3947 gnd.n3946 9.3005
R17959 gnd.n3945 gnd.n2965 9.3005
R17960 gnd.n4402 gnd.n2966 9.3005
R17961 gnd.n4401 gnd.n2967 9.3005
R17962 gnd.n4400 gnd.n2968 9.3005
R17963 gnd.n2989 gnd.n2969 9.3005
R17964 gnd.n2990 gnd.n2988 9.3005
R17965 gnd.n4388 gnd.n2991 9.3005
R17966 gnd.n4387 gnd.n2992 9.3005
R17967 gnd.n4386 gnd.n2993 9.3005
R17968 gnd.n3015 gnd.n2994 9.3005
R17969 gnd.n3016 gnd.n3014 9.3005
R17970 gnd.n4374 gnd.n3017 9.3005
R17971 gnd.n4373 gnd.n3018 9.3005
R17972 gnd.n4372 gnd.n3019 9.3005
R17973 gnd.n3040 gnd.n3020 9.3005
R17974 gnd.n3041 gnd.n3039 9.3005
R17975 gnd.n4360 gnd.n4359 9.3005
R17976 gnd.n3665 gnd.n3662 9.3005
R17977 gnd.n3447 gnd.n3406 9.3005
R17978 gnd.n3442 gnd.n3441 9.3005
R17979 gnd.n3440 gnd.n3407 9.3005
R17980 gnd.n3439 gnd.n3438 9.3005
R17981 gnd.n3435 gnd.n3408 9.3005
R17982 gnd.n3432 gnd.n3431 9.3005
R17983 gnd.n3430 gnd.n3409 9.3005
R17984 gnd.n3429 gnd.n3428 9.3005
R17985 gnd.n3425 gnd.n3410 9.3005
R17986 gnd.n3422 gnd.n3421 9.3005
R17987 gnd.n3420 gnd.n3411 9.3005
R17988 gnd.n3419 gnd.n3418 9.3005
R17989 gnd.n3415 gnd.n3413 9.3005
R17990 gnd.n3412 gnd.n3392 9.3005
R17991 gnd.n3659 gnd.n3391 9.3005
R17992 gnd.n3661 gnd.n3660 9.3005
R17993 gnd.n3449 gnd.n3448 9.3005
R17994 gnd.n3672 gnd.n3378 9.3005
R17995 gnd.n3679 gnd.n3379 9.3005
R17996 gnd.n3681 gnd.n3680 9.3005
R17997 gnd.n3682 gnd.n3359 9.3005
R17998 gnd.n3701 gnd.n3700 9.3005
R17999 gnd.n3703 gnd.n3351 9.3005
R18000 gnd.n3710 gnd.n3353 9.3005
R18001 gnd.n3711 gnd.n3348 9.3005
R18002 gnd.n3713 gnd.n3712 9.3005
R18003 gnd.n3349 gnd.n3334 9.3005
R18004 gnd.n3729 gnd.n3332 9.3005
R18005 gnd.n3733 gnd.n3732 9.3005
R18006 gnd.n3731 gnd.n3308 9.3005
R18007 gnd.n3768 gnd.n3307 9.3005
R18008 gnd.n3771 gnd.n3770 9.3005
R18009 gnd.n3304 gnd.n3303 9.3005
R18010 gnd.n3777 gnd.n3305 9.3005
R18011 gnd.n3779 gnd.n3778 9.3005
R18012 gnd.n3781 gnd.n3302 9.3005
R18013 gnd.n3784 gnd.n3783 9.3005
R18014 gnd.n3787 gnd.n3785 9.3005
R18015 gnd.n3789 gnd.n3788 9.3005
R18016 gnd.n3795 gnd.n3790 9.3005
R18017 gnd.n3794 gnd.n3793 9.3005
R18018 gnd.n3178 gnd.n3177 9.3005
R18019 gnd.n3861 gnd.n3860 9.3005
R18020 gnd.n3862 gnd.n3171 9.3005
R18021 gnd.n3870 gnd.n3170 9.3005
R18022 gnd.n3873 gnd.n3872 9.3005
R18023 gnd.n3875 gnd.n3874 9.3005
R18024 gnd.n3878 gnd.n3153 9.3005
R18025 gnd.n3876 gnd.n3151 9.3005
R18026 gnd.n3898 gnd.n3149 9.3005
R18027 gnd.n3902 gnd.n3901 9.3005
R18028 gnd.n3900 gnd.n3899 9.3005
R18029 gnd.n3127 gnd.n3126 9.3005
R18030 gnd.n3952 gnd.n3128 9.3005
R18031 gnd.n3954 gnd.n3953 9.3005
R18032 gnd.n3956 gnd.n3125 9.3005
R18033 gnd.n3959 gnd.n3958 9.3005
R18034 gnd.n3961 gnd.n3960 9.3005
R18035 gnd.n3965 gnd.n3962 9.3005
R18036 gnd.n3967 gnd.n3966 9.3005
R18037 gnd.n4252 gnd.n3969 9.3005
R18038 gnd.n4251 gnd.n3971 9.3005
R18039 gnd.n4250 gnd.n3972 9.3005
R18040 gnd.n4247 gnd.n3973 9.3005
R18041 gnd.n4246 gnd.n3974 9.3005
R18042 gnd.n4245 gnd.n4232 9.3005
R18043 gnd.n4242 gnd.n4234 9.3005
R18044 gnd.n4241 gnd.n4235 9.3005
R18045 gnd.n4238 gnd.n4236 9.3005
R18046 gnd.n4237 gnd.n3071 9.3005
R18047 gnd.n3670 gnd.n3669 9.3005
R18048 gnd.n4324 gnd.n3072 9.3005
R18049 gnd.n4323 gnd.n3074 9.3005
R18050 gnd.n3078 gnd.n3075 9.3005
R18051 gnd.n4318 gnd.n3079 9.3005
R18052 gnd.n4317 gnd.n3080 9.3005
R18053 gnd.n4316 gnd.n3081 9.3005
R18054 gnd.n3085 gnd.n3082 9.3005
R18055 gnd.n4311 gnd.n3086 9.3005
R18056 gnd.n4310 gnd.n3087 9.3005
R18057 gnd.n4309 gnd.n3088 9.3005
R18058 gnd.n3092 gnd.n3089 9.3005
R18059 gnd.n4304 gnd.n3093 9.3005
R18060 gnd.n4303 gnd.n3094 9.3005
R18061 gnd.n4302 gnd.n3095 9.3005
R18062 gnd.n3099 gnd.n3096 9.3005
R18063 gnd.n4297 gnd.n3100 9.3005
R18064 gnd.n4296 gnd.n3101 9.3005
R18065 gnd.n4295 gnd.n3102 9.3005
R18066 gnd.n3106 gnd.n3103 9.3005
R18067 gnd.n4290 gnd.n3107 9.3005
R18068 gnd.n4289 gnd.n3108 9.3005
R18069 gnd.n4288 gnd.n3109 9.3005
R18070 gnd.n3116 gnd.n3114 9.3005
R18071 gnd.n4283 gnd.n3117 9.3005
R18072 gnd.n4282 gnd.n3118 9.3005
R18073 gnd.n4281 gnd.n4278 9.3005
R18074 gnd.n4326 gnd.n4325 9.3005
R18075 gnd.n3839 gnd.n3823 9.3005
R18076 gnd.n3838 gnd.n3824 9.3005
R18077 gnd.n3837 gnd.n3825 9.3005
R18078 gnd.n3835 gnd.n3826 9.3005
R18079 gnd.n3834 gnd.n3827 9.3005
R18080 gnd.n3832 gnd.n3828 9.3005
R18081 gnd.n3831 gnd.n3829 9.3005
R18082 gnd.n3141 gnd.n3140 9.3005
R18083 gnd.n3910 gnd.n3909 9.3005
R18084 gnd.n3911 gnd.n3139 9.3005
R18085 gnd.n3937 gnd.n3912 9.3005
R18086 gnd.n3936 gnd.n3913 9.3005
R18087 gnd.n3935 gnd.n3914 9.3005
R18088 gnd.n3933 gnd.n3915 9.3005
R18089 gnd.n3932 gnd.n3916 9.3005
R18090 gnd.n3926 gnd.n3917 9.3005
R18091 gnd.n3925 gnd.n3918 9.3005
R18092 gnd.n3924 gnd.n3919 9.3005
R18093 gnd.n3921 gnd.n3920 9.3005
R18094 gnd.n3124 gnd.n3123 9.3005
R18095 gnd.n4259 gnd.n4258 9.3005
R18096 gnd.n4260 gnd.n3122 9.3005
R18097 gnd.n4264 gnd.n4261 9.3005
R18098 gnd.n4265 gnd.n3121 9.3005
R18099 gnd.n4269 gnd.n4268 9.3005
R18100 gnd.n4270 gnd.n3120 9.3005
R18101 gnd.n4272 gnd.n4271 9.3005
R18102 gnd.n4275 gnd.n3119 9.3005
R18103 gnd.n4277 gnd.n4276 9.3005
R18104 gnd.n3580 gnd.n3579 9.3005
R18105 gnd.n3470 gnd.n3469 9.3005
R18106 gnd.n3594 gnd.n3593 9.3005
R18107 gnd.n3595 gnd.n3468 9.3005
R18108 gnd.n3597 gnd.n3596 9.3005
R18109 gnd.n3458 gnd.n3457 9.3005
R18110 gnd.n3610 gnd.n3609 9.3005
R18111 gnd.n3611 gnd.n3456 9.3005
R18112 gnd.n3643 gnd.n3612 9.3005
R18113 gnd.n3642 gnd.n3613 9.3005
R18114 gnd.n3641 gnd.n3614 9.3005
R18115 gnd.n3640 gnd.n3615 9.3005
R18116 gnd.n3637 gnd.n3616 9.3005
R18117 gnd.n3636 gnd.n3617 9.3005
R18118 gnd.n3635 gnd.n3618 9.3005
R18119 gnd.n3633 gnd.n3619 9.3005
R18120 gnd.n3632 gnd.n3620 9.3005
R18121 gnd.n3629 gnd.n3621 9.3005
R18122 gnd.n3628 gnd.n3622 9.3005
R18123 gnd.n3627 gnd.n3623 9.3005
R18124 gnd.n3625 gnd.n3624 9.3005
R18125 gnd.n3324 gnd.n3323 9.3005
R18126 gnd.n3741 gnd.n3740 9.3005
R18127 gnd.n3742 gnd.n3322 9.3005
R18128 gnd.n3746 gnd.n3743 9.3005
R18129 gnd.n3745 gnd.n3744 9.3005
R18130 gnd.n3246 gnd.n3245 9.3005
R18131 gnd.n3821 gnd.n3820 9.3005
R18132 gnd.n3578 gnd.n3479 9.3005
R18133 gnd.n3481 gnd.n3480 9.3005
R18134 gnd.n3525 gnd.n3523 9.3005
R18135 gnd.n3526 gnd.n3522 9.3005
R18136 gnd.n3529 gnd.n3518 9.3005
R18137 gnd.n3530 gnd.n3517 9.3005
R18138 gnd.n3533 gnd.n3516 9.3005
R18139 gnd.n3534 gnd.n3515 9.3005
R18140 gnd.n3537 gnd.n3514 9.3005
R18141 gnd.n3538 gnd.n3513 9.3005
R18142 gnd.n3541 gnd.n3512 9.3005
R18143 gnd.n3542 gnd.n3511 9.3005
R18144 gnd.n3545 gnd.n3510 9.3005
R18145 gnd.n3546 gnd.n3509 9.3005
R18146 gnd.n3549 gnd.n3508 9.3005
R18147 gnd.n3550 gnd.n3507 9.3005
R18148 gnd.n3553 gnd.n3506 9.3005
R18149 gnd.n3554 gnd.n3505 9.3005
R18150 gnd.n3557 gnd.n3504 9.3005
R18151 gnd.n3558 gnd.n3503 9.3005
R18152 gnd.n3561 gnd.n3502 9.3005
R18153 gnd.n3562 gnd.n3501 9.3005
R18154 gnd.n3565 gnd.n3500 9.3005
R18155 gnd.n3567 gnd.n3499 9.3005
R18156 gnd.n3568 gnd.n3498 9.3005
R18157 gnd.n3569 gnd.n3497 9.3005
R18158 gnd.n3570 gnd.n3496 9.3005
R18159 gnd.n3577 gnd.n3576 9.3005
R18160 gnd.n3586 gnd.n3585 9.3005
R18161 gnd.n3587 gnd.n3473 9.3005
R18162 gnd.n3589 gnd.n3588 9.3005
R18163 gnd.n3464 gnd.n3463 9.3005
R18164 gnd.n3602 gnd.n3601 9.3005
R18165 gnd.n3603 gnd.n3462 9.3005
R18166 gnd.n3605 gnd.n3604 9.3005
R18167 gnd.n3451 gnd.n3450 9.3005
R18168 gnd.n3648 gnd.n3647 9.3005
R18169 gnd.n3649 gnd.n3405 9.3005
R18170 gnd.n3653 gnd.n3651 9.3005
R18171 gnd.n3652 gnd.n3384 9.3005
R18172 gnd.n3671 gnd.n3383 9.3005
R18173 gnd.n3674 gnd.n3673 9.3005
R18174 gnd.n3377 gnd.n3376 9.3005
R18175 gnd.n3685 gnd.n3683 9.3005
R18176 gnd.n3684 gnd.n3358 9.3005
R18177 gnd.n3702 gnd.n3357 9.3005
R18178 gnd.n3705 gnd.n3704 9.3005
R18179 gnd.n3352 gnd.n3347 9.3005
R18180 gnd.n3715 gnd.n3714 9.3005
R18181 gnd.n3350 gnd.n3330 9.3005
R18182 gnd.n3736 gnd.n3331 9.3005
R18183 gnd.n3735 gnd.n3734 9.3005
R18184 gnd.n3333 gnd.n3309 9.3005
R18185 gnd.n3767 gnd.n3766 9.3005
R18186 gnd.n3769 gnd.n3254 9.3005
R18187 gnd.n3816 gnd.n3255 9.3005
R18188 gnd.n3815 gnd.n3256 9.3005
R18189 gnd.n3814 gnd.n3257 9.3005
R18190 gnd.n3780 gnd.n3258 9.3005
R18191 gnd.n3782 gnd.n3276 9.3005
R18192 gnd.n3802 gnd.n3277 9.3005
R18193 gnd.n3801 gnd.n3278 9.3005
R18194 gnd.n3800 gnd.n3279 9.3005
R18195 gnd.n3791 gnd.n3280 9.3005
R18196 gnd.n3792 gnd.n3179 9.3005
R18197 gnd.n3858 gnd.n3857 9.3005
R18198 gnd.n3859 gnd.n3172 9.3005
R18199 gnd.n3869 gnd.n3868 9.3005
R18200 gnd.n3871 gnd.n3168 9.3005
R18201 gnd.n3881 gnd.n3169 9.3005
R18202 gnd.n3880 gnd.n3879 9.3005
R18203 gnd.n3877 gnd.n3147 9.3005
R18204 gnd.n3905 gnd.n3148 9.3005
R18205 gnd.n3904 gnd.n3903 9.3005
R18206 gnd.n3150 gnd.n2954 9.3005
R18207 gnd.n4409 gnd.n2955 9.3005
R18208 gnd.n4408 gnd.n2956 9.3005
R18209 gnd.n4407 gnd.n2957 9.3005
R18210 gnd.n3955 gnd.n2958 9.3005
R18211 gnd.n3957 gnd.n2977 9.3005
R18212 gnd.n4395 gnd.n2978 9.3005
R18213 gnd.n4394 gnd.n2979 9.3005
R18214 gnd.n4393 gnd.n2980 9.3005
R18215 gnd.n3968 gnd.n2981 9.3005
R18216 gnd.n3970 gnd.n3002 9.3005
R18217 gnd.n4381 gnd.n3003 9.3005
R18218 gnd.n4380 gnd.n3004 9.3005
R18219 gnd.n4379 gnd.n3005 9.3005
R18220 gnd.n4231 gnd.n3006 9.3005
R18221 gnd.n4233 gnd.n3028 9.3005
R18222 gnd.n4367 gnd.n3029 9.3005
R18223 gnd.n4366 gnd.n3030 9.3005
R18224 gnd.n4365 gnd.n3031 9.3005
R18225 gnd.n3475 gnd.n3474 9.3005
R18226 gnd.n2742 gnd.n2741 9.3005
R18227 gnd.n2740 gnd.n1683 9.3005
R18228 gnd.n1690 gnd.n1685 9.3005
R18229 gnd.n2734 gnd.n1691 9.3005
R18230 gnd.n2733 gnd.n1692 9.3005
R18231 gnd.n2732 gnd.n1693 9.3005
R18232 gnd.n1698 gnd.n1694 9.3005
R18233 gnd.n2726 gnd.n1699 9.3005
R18234 gnd.n2725 gnd.n1700 9.3005
R18235 gnd.n2724 gnd.n1701 9.3005
R18236 gnd.n1706 gnd.n1702 9.3005
R18237 gnd.n2718 gnd.n1707 9.3005
R18238 gnd.n2717 gnd.n1708 9.3005
R18239 gnd.n2716 gnd.n1709 9.3005
R18240 gnd.n1714 gnd.n1710 9.3005
R18241 gnd.n2710 gnd.n1715 9.3005
R18242 gnd.n2709 gnd.n1716 9.3005
R18243 gnd.n2708 gnd.n1717 9.3005
R18244 gnd.n1722 gnd.n1718 9.3005
R18245 gnd.n2702 gnd.n1723 9.3005
R18246 gnd.n2701 gnd.n1724 9.3005
R18247 gnd.n2700 gnd.n1725 9.3005
R18248 gnd.n1730 gnd.n1726 9.3005
R18249 gnd.n2694 gnd.n1731 9.3005
R18250 gnd.n2693 gnd.n1732 9.3005
R18251 gnd.n2692 gnd.n1733 9.3005
R18252 gnd.n1738 gnd.n1734 9.3005
R18253 gnd.n2686 gnd.n1739 9.3005
R18254 gnd.n2685 gnd.n1740 9.3005
R18255 gnd.n2684 gnd.n1741 9.3005
R18256 gnd.n1746 gnd.n1742 9.3005
R18257 gnd.n2678 gnd.n1747 9.3005
R18258 gnd.n2677 gnd.n1748 9.3005
R18259 gnd.n2676 gnd.n1749 9.3005
R18260 gnd.n1754 gnd.n1750 9.3005
R18261 gnd.n2670 gnd.n1755 9.3005
R18262 gnd.n2669 gnd.n1756 9.3005
R18263 gnd.n2668 gnd.n1757 9.3005
R18264 gnd.n1762 gnd.n1758 9.3005
R18265 gnd.n2662 gnd.n1763 9.3005
R18266 gnd.n2661 gnd.n1764 9.3005
R18267 gnd.n2660 gnd.n1765 9.3005
R18268 gnd.n1770 gnd.n1766 9.3005
R18269 gnd.n2654 gnd.n1771 9.3005
R18270 gnd.n2653 gnd.n1772 9.3005
R18271 gnd.n2652 gnd.n1773 9.3005
R18272 gnd.n1778 gnd.n1774 9.3005
R18273 gnd.n2646 gnd.n1779 9.3005
R18274 gnd.n2645 gnd.n1780 9.3005
R18275 gnd.n2644 gnd.n1781 9.3005
R18276 gnd.n1786 gnd.n1782 9.3005
R18277 gnd.n2638 gnd.n1787 9.3005
R18278 gnd.n2637 gnd.n1788 9.3005
R18279 gnd.n2636 gnd.n1789 9.3005
R18280 gnd.n1794 gnd.n1790 9.3005
R18281 gnd.n2630 gnd.n1795 9.3005
R18282 gnd.n2629 gnd.n1796 9.3005
R18283 gnd.n2628 gnd.n1797 9.3005
R18284 gnd.n1802 gnd.n1798 9.3005
R18285 gnd.n2622 gnd.n1803 9.3005
R18286 gnd.n2621 gnd.n1804 9.3005
R18287 gnd.n2620 gnd.n1805 9.3005
R18288 gnd.n1810 gnd.n1806 9.3005
R18289 gnd.n2614 gnd.n1811 9.3005
R18290 gnd.n2613 gnd.n1812 9.3005
R18291 gnd.n2612 gnd.n1813 9.3005
R18292 gnd.n1818 gnd.n1814 9.3005
R18293 gnd.n2606 gnd.n1819 9.3005
R18294 gnd.n2605 gnd.n1820 9.3005
R18295 gnd.n2604 gnd.n1821 9.3005
R18296 gnd.n1826 gnd.n1822 9.3005
R18297 gnd.n2598 gnd.n1827 9.3005
R18298 gnd.n2597 gnd.n1828 9.3005
R18299 gnd.n2596 gnd.n1829 9.3005
R18300 gnd.n1834 gnd.n1830 9.3005
R18301 gnd.n2590 gnd.n1835 9.3005
R18302 gnd.n2589 gnd.n1836 9.3005
R18303 gnd.n2588 gnd.n1837 9.3005
R18304 gnd.n1842 gnd.n1838 9.3005
R18305 gnd.n2582 gnd.n1843 9.3005
R18306 gnd.n2581 gnd.n1844 9.3005
R18307 gnd.n2580 gnd.n1845 9.3005
R18308 gnd.n1850 gnd.n1846 9.3005
R18309 gnd.n2574 gnd.n1851 9.3005
R18310 gnd.n2573 gnd.n1852 9.3005
R18311 gnd.n2572 gnd.n1853 9.3005
R18312 gnd.n1858 gnd.n1854 9.3005
R18313 gnd.n2566 gnd.n1859 9.3005
R18314 gnd.n2565 gnd.n1860 9.3005
R18315 gnd.n2564 gnd.n1861 9.3005
R18316 gnd.n1866 gnd.n1862 9.3005
R18317 gnd.n2558 gnd.n1867 9.3005
R18318 gnd.n2557 gnd.n1868 9.3005
R18319 gnd.n2556 gnd.n1869 9.3005
R18320 gnd.n1874 gnd.n1870 9.3005
R18321 gnd.n2550 gnd.n1875 9.3005
R18322 gnd.n2549 gnd.n1876 9.3005
R18323 gnd.n2548 gnd.n1877 9.3005
R18324 gnd.n1882 gnd.n1878 9.3005
R18325 gnd.n2542 gnd.n1883 9.3005
R18326 gnd.n2541 gnd.n1884 9.3005
R18327 gnd.n2540 gnd.n1885 9.3005
R18328 gnd.n1890 gnd.n1886 9.3005
R18329 gnd.n2534 gnd.n1891 9.3005
R18330 gnd.n2533 gnd.n1892 9.3005
R18331 gnd.n2532 gnd.n1893 9.3005
R18332 gnd.n1898 gnd.n1894 9.3005
R18333 gnd.n2526 gnd.n1899 9.3005
R18334 gnd.n2525 gnd.n1900 9.3005
R18335 gnd.n2524 gnd.n1901 9.3005
R18336 gnd.n1906 gnd.n1902 9.3005
R18337 gnd.n2518 gnd.n1907 9.3005
R18338 gnd.n2517 gnd.n1908 9.3005
R18339 gnd.n2516 gnd.n1909 9.3005
R18340 gnd.n1914 gnd.n1910 9.3005
R18341 gnd.n2510 gnd.n1915 9.3005
R18342 gnd.n2509 gnd.n1916 9.3005
R18343 gnd.n2508 gnd.n1917 9.3005
R18344 gnd.n1922 gnd.n1918 9.3005
R18345 gnd.n2502 gnd.n1923 9.3005
R18346 gnd.n2501 gnd.n1924 9.3005
R18347 gnd.n2500 gnd.n1925 9.3005
R18348 gnd.n1930 gnd.n1926 9.3005
R18349 gnd.n2494 gnd.n1931 9.3005
R18350 gnd.n2493 gnd.n1932 9.3005
R18351 gnd.n2492 gnd.n1933 9.3005
R18352 gnd.n1938 gnd.n1934 9.3005
R18353 gnd.n2486 gnd.n1939 9.3005
R18354 gnd.n2485 gnd.n1940 9.3005
R18355 gnd.n2484 gnd.n1941 9.3005
R18356 gnd.n1946 gnd.n1942 9.3005
R18357 gnd.n2478 gnd.n1947 9.3005
R18358 gnd.n2477 gnd.n1948 9.3005
R18359 gnd.n2476 gnd.n1949 9.3005
R18360 gnd.n1954 gnd.n1950 9.3005
R18361 gnd.n2470 gnd.n1955 9.3005
R18362 gnd.n2469 gnd.n1956 9.3005
R18363 gnd.n2468 gnd.n1957 9.3005
R18364 gnd.n1962 gnd.n1958 9.3005
R18365 gnd.n2462 gnd.n1963 9.3005
R18366 gnd.n2461 gnd.n1964 9.3005
R18367 gnd.n2460 gnd.n1965 9.3005
R18368 gnd.n1970 gnd.n1966 9.3005
R18369 gnd.n2454 gnd.n1971 9.3005
R18370 gnd.n2453 gnd.n1972 9.3005
R18371 gnd.n2452 gnd.n1973 9.3005
R18372 gnd.n1978 gnd.n1974 9.3005
R18373 gnd.n2446 gnd.n1979 9.3005
R18374 gnd.n2445 gnd.n1980 9.3005
R18375 gnd.n2444 gnd.n1981 9.3005
R18376 gnd.n1986 gnd.n1982 9.3005
R18377 gnd.n2438 gnd.n1987 9.3005
R18378 gnd.n2437 gnd.n1988 9.3005
R18379 gnd.n2436 gnd.n1989 9.3005
R18380 gnd.n1994 gnd.n1990 9.3005
R18381 gnd.n2430 gnd.n1995 9.3005
R18382 gnd.n2429 gnd.n1996 9.3005
R18383 gnd.n2428 gnd.n1997 9.3005
R18384 gnd.n2002 gnd.n1998 9.3005
R18385 gnd.n2422 gnd.n2003 9.3005
R18386 gnd.n2421 gnd.n2004 9.3005
R18387 gnd.n2420 gnd.n2005 9.3005
R18388 gnd.n2010 gnd.n2006 9.3005
R18389 gnd.n2414 gnd.n2011 9.3005
R18390 gnd.n2413 gnd.n2012 9.3005
R18391 gnd.n2412 gnd.n2013 9.3005
R18392 gnd.n2018 gnd.n2014 9.3005
R18393 gnd.n2406 gnd.n2019 9.3005
R18394 gnd.n2405 gnd.n2020 9.3005
R18395 gnd.n2404 gnd.n2021 9.3005
R18396 gnd.n2026 gnd.n2022 9.3005
R18397 gnd.n2398 gnd.n2027 9.3005
R18398 gnd.n2397 gnd.n2028 9.3005
R18399 gnd.n2396 gnd.n2029 9.3005
R18400 gnd.n2034 gnd.n2030 9.3005
R18401 gnd.n2390 gnd.n2035 9.3005
R18402 gnd.n2389 gnd.n2036 9.3005
R18403 gnd.n2388 gnd.n2037 9.3005
R18404 gnd.n2042 gnd.n2038 9.3005
R18405 gnd.n2382 gnd.n2043 9.3005
R18406 gnd.n2381 gnd.n2044 9.3005
R18407 gnd.n2380 gnd.n2045 9.3005
R18408 gnd.n2374 gnd.n2373 9.3005
R18409 gnd.n2372 gnd.n2050 9.3005
R18410 gnd.n2371 gnd.n2370 9.3005
R18411 gnd.n2053 gnd.n2052 9.3005
R18412 gnd.n2364 gnd.n2057 9.3005
R18413 gnd.n2363 gnd.n2058 9.3005
R18414 gnd.n2362 gnd.n2059 9.3005
R18415 gnd.n2064 gnd.n2060 9.3005
R18416 gnd.n2356 gnd.n2065 9.3005
R18417 gnd.n2355 gnd.n2066 9.3005
R18418 gnd.n2354 gnd.n2067 9.3005
R18419 gnd.n2072 gnd.n2068 9.3005
R18420 gnd.n2348 gnd.n2073 9.3005
R18421 gnd.n2347 gnd.n2074 9.3005
R18422 gnd.n2346 gnd.n2075 9.3005
R18423 gnd.n2080 gnd.n2076 9.3005
R18424 gnd.n2340 gnd.n2081 9.3005
R18425 gnd.n2339 gnd.n2082 9.3005
R18426 gnd.n2338 gnd.n2083 9.3005
R18427 gnd.n2088 gnd.n2084 9.3005
R18428 gnd.n2332 gnd.n2089 9.3005
R18429 gnd.n2331 gnd.n2090 9.3005
R18430 gnd.n2330 gnd.n2091 9.3005
R18431 gnd.n2096 gnd.n2092 9.3005
R18432 gnd.n2324 gnd.n2097 9.3005
R18433 gnd.n2323 gnd.n2098 9.3005
R18434 gnd.n2322 gnd.n2099 9.3005
R18435 gnd.n2104 gnd.n2100 9.3005
R18436 gnd.n2316 gnd.n2105 9.3005
R18437 gnd.n2315 gnd.n2106 9.3005
R18438 gnd.n2314 gnd.n2107 9.3005
R18439 gnd.n2112 gnd.n2108 9.3005
R18440 gnd.n2308 gnd.n2113 9.3005
R18441 gnd.n2307 gnd.n2114 9.3005
R18442 gnd.n2306 gnd.n2115 9.3005
R18443 gnd.n2120 gnd.n2116 9.3005
R18444 gnd.n2300 gnd.n2121 9.3005
R18445 gnd.n2299 gnd.n2122 9.3005
R18446 gnd.n2298 gnd.n2123 9.3005
R18447 gnd.n2128 gnd.n2124 9.3005
R18448 gnd.n2292 gnd.n2129 9.3005
R18449 gnd.n2291 gnd.n2130 9.3005
R18450 gnd.n2290 gnd.n2131 9.3005
R18451 gnd.n2136 gnd.n2132 9.3005
R18452 gnd.n2284 gnd.n2137 9.3005
R18453 gnd.n2283 gnd.n2138 9.3005
R18454 gnd.n2282 gnd.n2139 9.3005
R18455 gnd.n2144 gnd.n2140 9.3005
R18456 gnd.n2276 gnd.n2145 9.3005
R18457 gnd.n2275 gnd.n2146 9.3005
R18458 gnd.n2274 gnd.n2147 9.3005
R18459 gnd.n2152 gnd.n2148 9.3005
R18460 gnd.n2268 gnd.n2153 9.3005
R18461 gnd.n2267 gnd.n2154 9.3005
R18462 gnd.n2266 gnd.n2155 9.3005
R18463 gnd.n2160 gnd.n2156 9.3005
R18464 gnd.n2260 gnd.n2161 9.3005
R18465 gnd.n2259 gnd.n2162 9.3005
R18466 gnd.n2258 gnd.n2163 9.3005
R18467 gnd.n2168 gnd.n2164 9.3005
R18468 gnd.n2252 gnd.n2169 9.3005
R18469 gnd.n2251 gnd.n2170 9.3005
R18470 gnd.n2250 gnd.n2171 9.3005
R18471 gnd.n2176 gnd.n2172 9.3005
R18472 gnd.n2244 gnd.n2177 9.3005
R18473 gnd.n2243 gnd.n2178 9.3005
R18474 gnd.n2242 gnd.n2179 9.3005
R18475 gnd.n2184 gnd.n2180 9.3005
R18476 gnd.n2236 gnd.n2185 9.3005
R18477 gnd.n2235 gnd.n2186 9.3005
R18478 gnd.n2234 gnd.n2187 9.3005
R18479 gnd.n2192 gnd.n2188 9.3005
R18480 gnd.n2228 gnd.n2193 9.3005
R18481 gnd.n2227 gnd.n2194 9.3005
R18482 gnd.n2226 gnd.n2195 9.3005
R18483 gnd.n2200 gnd.n2196 9.3005
R18484 gnd.n2220 gnd.n2201 9.3005
R18485 gnd.n2219 gnd.n2202 9.3005
R18486 gnd.n2218 gnd.n2203 9.3005
R18487 gnd.n2208 gnd.n2204 9.3005
R18488 gnd.n2212 gnd.n2209 9.3005
R18489 gnd.n2211 gnd.n2210 9.3005
R18490 gnd.n246 gnd.n245 9.3005
R18491 gnd.n7038 gnd.n7037 9.3005
R18492 gnd.n2051 gnd.n2049 9.3005
R18493 gnd.n7329 gnd.n7328 9.3005
R18494 gnd.n7327 gnd.n65 9.3005
R18495 gnd.n267 gnd.n67 9.3005
R18496 gnd.n6995 gnd.n268 9.3005
R18497 gnd.n6994 gnd.n269 9.3005
R18498 gnd.n6993 gnd.n270 9.3005
R18499 gnd.n6933 gnd.n271 9.3005
R18500 gnd.n6983 gnd.n6934 9.3005
R18501 gnd.n6982 gnd.n6935 9.3005
R18502 gnd.n6981 gnd.n6936 9.3005
R18503 gnd.n6941 gnd.n6937 9.3005
R18504 gnd.n6971 gnd.n6942 9.3005
R18505 gnd.n6970 gnd.n6943 9.3005
R18506 gnd.n6969 gnd.n6944 9.3005
R18507 gnd.n6948 gnd.n6945 9.3005
R18508 gnd.n6959 gnd.n6949 9.3005
R18509 gnd.n6958 gnd.n6950 9.3005
R18510 gnd.n6957 gnd.n6952 9.3005
R18511 gnd.n6951 gnd.n177 9.3005
R18512 gnd.n7260 gnd.n178 9.3005
R18513 gnd.n7259 gnd.n7258 9.3005
R18514 gnd.n203 gnd.n199 9.3005
R18515 gnd.n207 gnd.n206 9.3005
R18516 gnd.n208 gnd.n198 9.3005
R18517 gnd.n210 gnd.n209 9.3005
R18518 gnd.n213 gnd.n197 9.3005
R18519 gnd.n217 gnd.n216 9.3005
R18520 gnd.n218 gnd.n196 9.3005
R18521 gnd.n220 gnd.n219 9.3005
R18522 gnd.n223 gnd.n195 9.3005
R18523 gnd.n227 gnd.n226 9.3005
R18524 gnd.n228 gnd.n194 9.3005
R18525 gnd.n230 gnd.n229 9.3005
R18526 gnd.n233 gnd.n193 9.3005
R18527 gnd.n236 gnd.n235 9.3005
R18528 gnd.n237 gnd.n192 9.3005
R18529 gnd.n239 gnd.n238 9.3005
R18530 gnd.n182 gnd.n179 9.3005
R18531 gnd.n7257 gnd.n7256 9.3005
R18532 gnd.n201 gnd.n200 9.3005
R18533 gnd.n7074 gnd.n7071 9.3005
R18534 gnd.n7250 gnd.n7075 9.3005
R18535 gnd.n7249 gnd.n7076 9.3005
R18536 gnd.n7248 gnd.n7077 9.3005
R18537 gnd.n7245 gnd.n7078 9.3005
R18538 gnd.n7244 gnd.n7079 9.3005
R18539 gnd.n7241 gnd.n7080 9.3005
R18540 gnd.n7240 gnd.n7081 9.3005
R18541 gnd.n7237 gnd.n7082 9.3005
R18542 gnd.n7236 gnd.n7083 9.3005
R18543 gnd.n7233 gnd.n7084 9.3005
R18544 gnd.n7232 gnd.n7085 9.3005
R18545 gnd.n7229 gnd.n7086 9.3005
R18546 gnd.n7228 gnd.n7087 9.3005
R18547 gnd.n7225 gnd.n7088 9.3005
R18548 gnd.n7224 gnd.n7089 9.3005
R18549 gnd.n7221 gnd.n7090 9.3005
R18550 gnd.n7217 gnd.n7091 9.3005
R18551 gnd.n7214 gnd.n7092 9.3005
R18552 gnd.n7213 gnd.n7093 9.3005
R18553 gnd.n7210 gnd.n7094 9.3005
R18554 gnd.n7209 gnd.n7095 9.3005
R18555 gnd.n7206 gnd.n7096 9.3005
R18556 gnd.n7205 gnd.n7097 9.3005
R18557 gnd.n7202 gnd.n7098 9.3005
R18558 gnd.n7201 gnd.n7099 9.3005
R18559 gnd.n7198 gnd.n7100 9.3005
R18560 gnd.n7197 gnd.n7101 9.3005
R18561 gnd.n7194 gnd.n7102 9.3005
R18562 gnd.n7193 gnd.n7103 9.3005
R18563 gnd.n7190 gnd.n7104 9.3005
R18564 gnd.n7189 gnd.n7105 9.3005
R18565 gnd.n7186 gnd.n7106 9.3005
R18566 gnd.n7185 gnd.n7107 9.3005
R18567 gnd.n7182 gnd.n7108 9.3005
R18568 gnd.n7181 gnd.n7109 9.3005
R18569 gnd.n7178 gnd.n7177 9.3005
R18570 gnd.n7176 gnd.n7110 9.3005
R18571 gnd.n7175 gnd.n7174 9.3005
R18572 gnd.n7171 gnd.n7113 9.3005
R18573 gnd.n7168 gnd.n7114 9.3005
R18574 gnd.n7167 gnd.n7115 9.3005
R18575 gnd.n7164 gnd.n7116 9.3005
R18576 gnd.n7163 gnd.n7117 9.3005
R18577 gnd.n7160 gnd.n7118 9.3005
R18578 gnd.n7159 gnd.n7119 9.3005
R18579 gnd.n7156 gnd.n7120 9.3005
R18580 gnd.n7155 gnd.n7121 9.3005
R18581 gnd.n7152 gnd.n7122 9.3005
R18582 gnd.n7151 gnd.n7123 9.3005
R18583 gnd.n7148 gnd.n7124 9.3005
R18584 gnd.n7147 gnd.n7125 9.3005
R18585 gnd.n7144 gnd.n7126 9.3005
R18586 gnd.n7143 gnd.n7127 9.3005
R18587 gnd.n7140 gnd.n7128 9.3005
R18588 gnd.n7139 gnd.n7129 9.3005
R18589 gnd.n7136 gnd.n7135 9.3005
R18590 gnd.n7134 gnd.n7131 9.3005
R18591 gnd.n7073 gnd.n7072 9.3005
R18592 gnd.n6732 gnd.n6731 9.3005
R18593 gnd.n400 gnd.n398 9.3005
R18594 gnd.n403 gnd.n402 9.3005
R18595 gnd.n406 gnd.n405 9.3005
R18596 gnd.n407 gnd.n364 9.3005
R18597 gnd.n6801 gnd.n365 9.3005
R18598 gnd.n6800 gnd.n366 9.3005
R18599 gnd.n6799 gnd.n6794 9.3005
R18600 gnd.n6798 gnd.n6795 9.3005
R18601 gnd.n340 gnd.n336 9.3005
R18602 gnd.n6836 gnd.n337 9.3005
R18603 gnd.n6835 gnd.n338 9.3005
R18604 gnd.n6834 gnd.n6830 9.3005
R18605 gnd.n6833 gnd.n310 9.3005
R18606 gnd.n6868 gnd.n309 9.3005
R18607 gnd.n6870 gnd.n6869 9.3005
R18608 gnd.n299 gnd.n298 9.3005
R18609 gnd.n6883 gnd.n6882 9.3005
R18610 gnd.n282 gnd.n281 9.3005
R18611 gnd.n6915 gnd.n6914 9.3005
R18612 gnd.n6916 gnd.n275 9.3005
R18613 gnd.n6923 gnd.n276 9.3005
R18614 gnd.n6924 gnd.n274 9.3005
R18615 gnd.n6927 gnd.n6926 9.3005
R18616 gnd.n6928 gnd.n92 9.3005
R18617 gnd.n7315 gnd.n93 9.3005
R18618 gnd.n7314 gnd.n94 9.3005
R18619 gnd.n7313 gnd.n95 9.3005
R18620 gnd.n6931 gnd.n96 9.3005
R18621 gnd.n7303 gnd.n112 9.3005
R18622 gnd.n7302 gnd.n113 9.3005
R18623 gnd.n7301 gnd.n114 9.3005
R18624 gnd.n6939 gnd.n115 9.3005
R18625 gnd.n7291 gnd.n133 9.3005
R18626 gnd.n7290 gnd.n134 9.3005
R18627 gnd.n7289 gnd.n135 9.3005
R18628 gnd.n6946 gnd.n136 9.3005
R18629 gnd.n7279 gnd.n154 9.3005
R18630 gnd.n7278 gnd.n155 9.3005
R18631 gnd.n7277 gnd.n156 9.3005
R18632 gnd.n173 gnd.n157 9.3005
R18633 gnd.n7267 gnd.n7266 9.3005
R18634 gnd.n399 gnd.n397 9.3005
R18635 gnd.n6731 gnd.n6730 9.3005
R18636 gnd.n6729 gnd.n400 9.3005
R18637 gnd.n411 gnd.n402 9.3005
R18638 gnd.n410 gnd.n406 9.3005
R18639 gnd.n408 gnd.n407 9.3005
R18640 gnd.n367 gnd.n365 9.3005
R18641 gnd.n6792 gnd.n366 9.3005
R18642 gnd.n6794 gnd.n6793 9.3005
R18643 gnd.n6795 gnd.n339 9.3005
R18644 gnd.n6824 gnd.n340 9.3005
R18645 gnd.n6825 gnd.n337 9.3005
R18646 gnd.n6828 gnd.n338 9.3005
R18647 gnd.n6830 gnd.n6829 9.3005
R18648 gnd.n311 gnd.n310 9.3005
R18649 gnd.n6868 gnd.n6867 9.3005
R18650 gnd.n6869 gnd.n300 9.3005
R18651 gnd.n6879 gnd.n299 9.3005
R18652 gnd.n6882 gnd.n6881 9.3005
R18653 gnd.n6880 gnd.n281 9.3005
R18654 gnd.n6915 gnd.n280 9.3005
R18655 gnd.n6917 gnd.n6916 9.3005
R18656 gnd.n6919 gnd.n276 9.3005
R18657 gnd.n6918 gnd.n274 9.3005
R18658 gnd.n6927 gnd.n273 9.3005
R18659 gnd.n6929 gnd.n6928 9.3005
R18660 gnd.n6930 gnd.n93 9.3005
R18661 gnd.n6989 gnd.n94 9.3005
R18662 gnd.n6988 gnd.n95 9.3005
R18663 gnd.n6987 gnd.n6931 9.3005
R18664 gnd.n6932 gnd.n112 9.3005
R18665 gnd.n6977 gnd.n113 9.3005
R18666 gnd.n6976 gnd.n114 9.3005
R18667 gnd.n6975 gnd.n6939 9.3005
R18668 gnd.n6940 gnd.n133 9.3005
R18669 gnd.n6965 gnd.n134 9.3005
R18670 gnd.n6964 gnd.n135 9.3005
R18671 gnd.n6963 gnd.n6946 9.3005
R18672 gnd.n6947 gnd.n154 9.3005
R18673 gnd.n6953 gnd.n155 9.3005
R18674 gnd.n175 gnd.n156 9.3005
R18675 gnd.n7264 gnd.n173 9.3005
R18676 gnd.n7266 gnd.n7265 9.3005
R18677 gnd.n401 gnd.n399 9.3005
R18678 gnd.n6580 gnd.n6579 9.3005
R18679 gnd.n6583 gnd.n558 9.3005
R18680 gnd.n6584 gnd.n557 9.3005
R18681 gnd.n6587 gnd.n556 9.3005
R18682 gnd.n6588 gnd.n555 9.3005
R18683 gnd.n6591 gnd.n554 9.3005
R18684 gnd.n6592 gnd.n553 9.3005
R18685 gnd.n6595 gnd.n552 9.3005
R18686 gnd.n6596 gnd.n551 9.3005
R18687 gnd.n6599 gnd.n550 9.3005
R18688 gnd.n6600 gnd.n549 9.3005
R18689 gnd.n6603 gnd.n548 9.3005
R18690 gnd.n6604 gnd.n547 9.3005
R18691 gnd.n6607 gnd.n546 9.3005
R18692 gnd.n6608 gnd.n545 9.3005
R18693 gnd.n6611 gnd.n544 9.3005
R18694 gnd.n6612 gnd.n543 9.3005
R18695 gnd.n6615 gnd.n542 9.3005
R18696 gnd.n6616 gnd.n541 9.3005
R18697 gnd.n6619 gnd.n540 9.3005
R18698 gnd.n6623 gnd.n536 9.3005
R18699 gnd.n6624 gnd.n535 9.3005
R18700 gnd.n6627 gnd.n534 9.3005
R18701 gnd.n6628 gnd.n533 9.3005
R18702 gnd.n6631 gnd.n532 9.3005
R18703 gnd.n6632 gnd.n531 9.3005
R18704 gnd.n6635 gnd.n530 9.3005
R18705 gnd.n6636 gnd.n529 9.3005
R18706 gnd.n6639 gnd.n528 9.3005
R18707 gnd.n6641 gnd.n524 9.3005
R18708 gnd.n6644 gnd.n523 9.3005
R18709 gnd.n6645 gnd.n522 9.3005
R18710 gnd.n6648 gnd.n521 9.3005
R18711 gnd.n6649 gnd.n520 9.3005
R18712 gnd.n6652 gnd.n519 9.3005
R18713 gnd.n6653 gnd.n518 9.3005
R18714 gnd.n6656 gnd.n517 9.3005
R18715 gnd.n6658 gnd.n514 9.3005
R18716 gnd.n6661 gnd.n513 9.3005
R18717 gnd.n6662 gnd.n512 9.3005
R18718 gnd.n6665 gnd.n511 9.3005
R18719 gnd.n6666 gnd.n510 9.3005
R18720 gnd.n6669 gnd.n509 9.3005
R18721 gnd.n6670 gnd.n508 9.3005
R18722 gnd.n6673 gnd.n507 9.3005
R18723 gnd.n6674 gnd.n506 9.3005
R18724 gnd.n6677 gnd.n505 9.3005
R18725 gnd.n6678 gnd.n504 9.3005
R18726 gnd.n6681 gnd.n503 9.3005
R18727 gnd.n6682 gnd.n502 9.3005
R18728 gnd.n6685 gnd.n501 9.3005
R18729 gnd.n6687 gnd.n500 9.3005
R18730 gnd.n6688 gnd.n499 9.3005
R18731 gnd.n6689 gnd.n498 9.3005
R18732 gnd.n6690 gnd.n497 9.3005
R18733 gnd.n6620 gnd.n537 9.3005
R18734 gnd.n6578 gnd.n560 9.3005
R18735 gnd.n6737 gnd.n6736 9.3005
R18736 gnd.n6738 gnd.n388 9.3005
R18737 gnd.n6742 gnd.n6739 9.3005
R18738 gnd.n6741 gnd.n6740 9.3005
R18739 gnd.n357 gnd.n356 9.3005
R18740 gnd.n6806 gnd.n6805 9.3005
R18741 gnd.n6807 gnd.n355 9.3005
R18742 gnd.n6811 gnd.n6808 9.3005
R18743 gnd.n6810 gnd.n6809 9.3005
R18744 gnd.n328 gnd.n327 9.3005
R18745 gnd.n6841 gnd.n6840 9.3005
R18746 gnd.n6842 gnd.n326 9.3005
R18747 gnd.n6847 gnd.n6843 9.3005
R18748 gnd.n6846 gnd.n6844 9.3005
R18749 gnd.n6845 gnd.n78 9.3005
R18750 gnd.n83 gnd.n77 9.3005
R18751 gnd.n7309 gnd.n103 9.3005
R18752 gnd.n7308 gnd.n104 9.3005
R18753 gnd.n7307 gnd.n105 9.3005
R18754 gnd.n122 gnd.n106 9.3005
R18755 gnd.n7297 gnd.n123 9.3005
R18756 gnd.n7296 gnd.n124 9.3005
R18757 gnd.n7295 gnd.n125 9.3005
R18758 gnd.n143 gnd.n126 9.3005
R18759 gnd.n7285 gnd.n144 9.3005
R18760 gnd.n7284 gnd.n145 9.3005
R18761 gnd.n7283 gnd.n146 9.3005
R18762 gnd.n163 gnd.n147 9.3005
R18763 gnd.n7273 gnd.n164 9.3005
R18764 gnd.n7272 gnd.n165 9.3005
R18765 gnd.n7271 gnd.n166 9.3005
R18766 gnd.n390 gnd.n389 9.3005
R18767 gnd.n7320 gnd.n7319 9.3005
R18768 gnd.n1397 gnd.n1396 9.3005
R18769 gnd.n1332 gnd.n1331 9.3005
R18770 gnd.n4944 gnd.n4943 9.3005
R18771 gnd.n4945 gnd.n1330 9.3005
R18772 gnd.n4958 gnd.n4946 9.3005
R18773 gnd.n4957 gnd.n4947 9.3005
R18774 gnd.n4956 gnd.n4948 9.3005
R18775 gnd.n4950 gnd.n4949 9.3005
R18776 gnd.n4952 gnd.n4951 9.3005
R18777 gnd.n1282 gnd.n1281 9.3005
R18778 gnd.n5020 gnd.n5019 9.3005
R18779 gnd.n5021 gnd.n1280 9.3005
R18780 gnd.n5023 gnd.n5022 9.3005
R18781 gnd.n1278 gnd.n1277 9.3005
R18782 gnd.n5030 gnd.n5029 9.3005
R18783 gnd.n5031 gnd.n1276 9.3005
R18784 gnd.n5187 gnd.n5032 9.3005
R18785 gnd.n5186 gnd.n5033 9.3005
R18786 gnd.n5185 gnd.n5034 9.3005
R18787 gnd.n5037 gnd.n5035 9.3005
R18788 gnd.n5179 gnd.n5038 9.3005
R18789 gnd.n5178 gnd.n5039 9.3005
R18790 gnd.n5177 gnd.n5040 9.3005
R18791 gnd.n5099 gnd.n5041 9.3005
R18792 gnd.n5102 gnd.n5101 9.3005
R18793 gnd.n5103 gnd.n5098 9.3005
R18794 gnd.n5105 gnd.n5104 9.3005
R18795 gnd.n5079 gnd.n5078 9.3005
R18796 gnd.n5123 gnd.n5122 9.3005
R18797 gnd.n5124 gnd.n5077 9.3005
R18798 gnd.n5126 gnd.n5125 9.3005
R18799 gnd.n5066 gnd.n5065 9.3005
R18800 gnd.n5144 gnd.n5143 9.3005
R18801 gnd.n5145 gnd.n5064 9.3005
R18802 gnd.n5149 gnd.n5146 9.3005
R18803 gnd.n5148 gnd.n5147 9.3005
R18804 gnd.n1068 gnd.n1067 9.3005
R18805 gnd.n5631 gnd.n5630 9.3005
R18806 gnd.n5632 gnd.n1066 9.3005
R18807 gnd.n5646 gnd.n5633 9.3005
R18808 gnd.n5645 gnd.n5634 9.3005
R18809 gnd.n5644 gnd.n5635 9.3005
R18810 gnd.n5637 gnd.n5636 9.3005
R18811 gnd.n5639 gnd.n5638 9.3005
R18812 gnd.n986 gnd.n985 9.3005
R18813 gnd.n5697 gnd.n5696 9.3005
R18814 gnd.n5698 gnd.n984 9.3005
R18815 gnd.n5702 gnd.n5699 9.3005
R18816 gnd.n5701 gnd.n5700 9.3005
R18817 gnd.n924 gnd.n923 9.3005
R18818 gnd.n5768 gnd.n5767 9.3005
R18819 gnd.n5769 gnd.n922 9.3005
R18820 gnd.n5771 gnd.n5770 9.3005
R18821 gnd.n920 gnd.n919 9.3005
R18822 gnd.n5776 gnd.n5775 9.3005
R18823 gnd.n5777 gnd.n918 9.3005
R18824 gnd.n5779 gnd.n5778 9.3005
R18825 gnd.n869 gnd.n868 9.3005
R18826 gnd.n5869 gnd.n5868 9.3005
R18827 gnd.n5870 gnd.n867 9.3005
R18828 gnd.n5880 gnd.n5871 9.3005
R18829 gnd.n5879 gnd.n5872 9.3005
R18830 gnd.n5878 gnd.n5873 9.3005
R18831 gnd.n5875 gnd.n5874 9.3005
R18832 gnd.n830 gnd.n829 9.3005
R18833 gnd.n5926 gnd.n5925 9.3005
R18834 gnd.n5927 gnd.n828 9.3005
R18835 gnd.n5934 gnd.n5928 9.3005
R18836 gnd.n5933 gnd.n5929 9.3005
R18837 gnd.n5932 gnd.n5930 9.3005
R18838 gnd.n783 gnd.n782 9.3005
R18839 gnd.n6081 gnd.n6080 9.3005
R18840 gnd.n6082 gnd.n781 9.3005
R18841 gnd.n6086 gnd.n6083 9.3005
R18842 gnd.n6085 gnd.n6084 9.3005
R18843 gnd.n754 gnd.n753 9.3005
R18844 gnd.n6117 gnd.n6116 9.3005
R18845 gnd.n6118 gnd.n752 9.3005
R18846 gnd.n6120 gnd.n6119 9.3005
R18847 gnd.n731 gnd.n730 9.3005
R18848 gnd.n6144 gnd.n6143 9.3005
R18849 gnd.n6145 gnd.n729 9.3005
R18850 gnd.n6147 gnd.n6146 9.3005
R18851 gnd.n705 gnd.n704 9.3005
R18852 gnd.n6183 gnd.n6182 9.3005
R18853 gnd.n6184 gnd.n703 9.3005
R18854 gnd.n6186 gnd.n6185 9.3005
R18855 gnd.n652 gnd.n651 9.3005
R18856 gnd.n6355 gnd.n6354 9.3005
R18857 gnd.n6356 gnd.n650 9.3005
R18858 gnd.n6360 gnd.n6357 9.3005
R18859 gnd.n6359 gnd.n6358 9.3005
R18860 gnd.n627 gnd.n626 9.3005
R18861 gnd.n6385 gnd.n6384 9.3005
R18862 gnd.n6386 gnd.n625 9.3005
R18863 gnd.n6390 gnd.n6387 9.3005
R18864 gnd.n6389 gnd.n6388 9.3005
R18865 gnd.n602 gnd.n601 9.3005
R18866 gnd.n6415 gnd.n6414 9.3005
R18867 gnd.n6416 gnd.n600 9.3005
R18868 gnd.n6420 gnd.n6417 9.3005
R18869 gnd.n6419 gnd.n6418 9.3005
R18870 gnd.n577 gnd.n576 9.3005
R18871 gnd.n6445 gnd.n6444 9.3005
R18872 gnd.n6446 gnd.n575 9.3005
R18873 gnd.n6460 gnd.n6447 9.3005
R18874 gnd.n6459 gnd.n6448 9.3005
R18875 gnd.n6458 gnd.n6449 9.3005
R18876 gnd.n6451 gnd.n6450 9.3005
R18877 gnd.n6453 gnd.n6452 9.3005
R18878 gnd.n416 gnd.n415 9.3005
R18879 gnd.n6719 gnd.n6718 9.3005
R18880 gnd.n6720 gnd.n414 9.3005
R18881 gnd.n6724 gnd.n6721 9.3005
R18882 gnd.n6723 gnd.n6722 9.3005
R18883 gnd.n372 gnd.n371 9.3005
R18884 gnd.n6757 gnd.n6756 9.3005
R18885 gnd.n6758 gnd.n370 9.3005
R18886 gnd.n6787 gnd.n6759 9.3005
R18887 gnd.n6786 gnd.n6760 9.3005
R18888 gnd.n6785 gnd.n6761 9.3005
R18889 gnd.n6764 gnd.n6762 9.3005
R18890 gnd.n6781 gnd.n6765 9.3005
R18891 gnd.n6780 gnd.n6766 9.3005
R18892 gnd.n6779 gnd.n6767 9.3005
R18893 gnd.n6770 gnd.n6768 9.3005
R18894 gnd.n6775 gnd.n6771 9.3005
R18895 gnd.n6774 gnd.n6772 9.3005
R18896 gnd.n7003 gnd.n7002 9.3005
R18897 gnd.n7005 gnd.n7004 9.3005
R18898 gnd.n260 gnd.n259 9.3005
R18899 gnd.n7010 gnd.n7009 9.3005
R18900 gnd.n7011 gnd.n258 9.3005
R18901 gnd.n7013 gnd.n7012 9.3005
R18902 gnd.n256 gnd.n255 9.3005
R18903 gnd.n7018 gnd.n7017 9.3005
R18904 gnd.n7019 gnd.n254 9.3005
R18905 gnd.n7021 gnd.n7020 9.3005
R18906 gnd.n252 gnd.n251 9.3005
R18907 gnd.n7026 gnd.n7025 9.3005
R18908 gnd.n7027 gnd.n250 9.3005
R18909 gnd.n7030 gnd.n7029 9.3005
R18910 gnd.n7028 gnd.n248 9.3005
R18911 gnd.n7034 gnd.n247 9.3005
R18912 gnd.n7036 gnd.n7035 9.3005
R18913 gnd.n4847 gnd.n4846 9.3005
R18914 gnd.n4717 gnd.n4716 9.3005
R18915 gnd.n4718 gnd.n1502 9.3005
R18916 gnd.n4726 gnd.n4719 9.3005
R18917 gnd.n4725 gnd.n4720 9.3005
R18918 gnd.n4724 gnd.n4721 9.3005
R18919 gnd.n1477 gnd.n1476 9.3005
R18920 gnd.n4753 gnd.n4752 9.3005
R18921 gnd.n4754 gnd.n1475 9.3005
R18922 gnd.n4757 gnd.n4756 9.3005
R18923 gnd.n4755 gnd.n1452 9.3005
R18924 gnd.n4797 gnd.n1453 9.3005
R18925 gnd.n4796 gnd.n1454 9.3005
R18926 gnd.n4795 gnd.n1455 9.3005
R18927 gnd.n1420 gnd.n1419 9.3005
R18928 gnd.n4830 gnd.n4829 9.3005
R18929 gnd.n4831 gnd.n1418 9.3005
R18930 gnd.n4851 gnd.n4832 9.3005
R18931 gnd.n4850 gnd.n4833 9.3005
R18932 gnd.n4849 gnd.n4834 9.3005
R18933 gnd.n4848 gnd.n4835 9.3005
R18934 gnd.n1504 gnd.n1503 9.3005
R18935 gnd.n4549 gnd.n4548 9.3005
R18936 gnd.n4552 gnd.n4540 9.3005
R18937 gnd.n4553 gnd.n4539 9.3005
R18938 gnd.n4556 gnd.n4538 9.3005
R18939 gnd.n4557 gnd.n4537 9.3005
R18940 gnd.n4560 gnd.n4536 9.3005
R18941 gnd.n4561 gnd.n4535 9.3005
R18942 gnd.n4564 gnd.n4534 9.3005
R18943 gnd.n4565 gnd.n4533 9.3005
R18944 gnd.n4568 gnd.n4532 9.3005
R18945 gnd.n4569 gnd.n4531 9.3005
R18946 gnd.n4572 gnd.n4530 9.3005
R18947 gnd.n4573 gnd.n4529 9.3005
R18948 gnd.n4576 gnd.n4528 9.3005
R18949 gnd.n4577 gnd.n4527 9.3005
R18950 gnd.n4580 gnd.n4526 9.3005
R18951 gnd.n4581 gnd.n4516 9.3005
R18952 gnd.n4547 gnd.n4544 9.3005
R18953 gnd.n4546 gnd.n4545 9.3005
R18954 gnd.n1151 gnd.n1149 9.3005
R18955 gnd.n5410 gnd.n5405 9.3005
R18956 gnd.n5411 gnd.n5404 9.3005
R18957 gnd.n5412 gnd.n5403 9.3005
R18958 gnd.n5402 gnd.n5399 9.3005
R18959 gnd.n5417 gnd.n5398 9.3005
R18960 gnd.n5418 gnd.n5397 9.3005
R18961 gnd.n5419 gnd.n5396 9.3005
R18962 gnd.n5395 gnd.n5389 9.3005
R18963 gnd.n5424 gnd.n5388 9.3005
R18964 gnd.n5425 gnd.n5387 9.3005
R18965 gnd.n5426 gnd.n5386 9.3005
R18966 gnd.n5385 gnd.n5382 9.3005
R18967 gnd.n5431 gnd.n5381 9.3005
R18968 gnd.n5432 gnd.n5380 9.3005
R18969 gnd.n5433 gnd.n5379 9.3005
R18970 gnd.n5378 gnd.n5375 9.3005
R18971 gnd.n5438 gnd.n5374 9.3005
R18972 gnd.n5439 gnd.n5373 9.3005
R18973 gnd.n5440 gnd.n5372 9.3005
R18974 gnd.n5371 gnd.n5368 9.3005
R18975 gnd.n5445 gnd.n5367 9.3005
R18976 gnd.n5446 gnd.n5366 9.3005
R18977 gnd.n5447 gnd.n5365 9.3005
R18978 gnd.n5363 gnd.n5362 9.3005
R18979 gnd.n5453 gnd.n5452 9.3005
R18980 gnd.n5520 gnd.n5519 9.3005
R18981 gnd.n1153 gnd.n1152 9.3005
R18982 gnd.n1159 gnd.n1157 9.3005
R18983 gnd.n5512 gnd.n1160 9.3005
R18984 gnd.n5511 gnd.n1161 9.3005
R18985 gnd.n5510 gnd.n1162 9.3005
R18986 gnd.n1166 gnd.n1163 9.3005
R18987 gnd.n5505 gnd.n1167 9.3005
R18988 gnd.n5504 gnd.n5503 9.3005
R18989 gnd.n5502 gnd.n1168 9.3005
R18990 gnd.n5501 gnd.n5500 9.3005
R18991 gnd.n1172 gnd.n1171 9.3005
R18992 gnd.n1177 gnd.n1175 9.3005
R18993 gnd.n5493 gnd.n1178 9.3005
R18994 gnd.n5492 gnd.n1179 9.3005
R18995 gnd.n5491 gnd.n1180 9.3005
R18996 gnd.n1184 gnd.n1181 9.3005
R18997 gnd.n5486 gnd.n1185 9.3005
R18998 gnd.n5485 gnd.n1186 9.3005
R18999 gnd.n5484 gnd.n1187 9.3005
R19000 gnd.n1191 gnd.n1188 9.3005
R19001 gnd.n5479 gnd.n1192 9.3005
R19002 gnd.n5478 gnd.n1193 9.3005
R19003 gnd.n5477 gnd.n1194 9.3005
R19004 gnd.n1198 gnd.n1195 9.3005
R19005 gnd.n5472 gnd.n1199 9.3005
R19006 gnd.n5471 gnd.n1200 9.3005
R19007 gnd.n5470 gnd.n1201 9.3005
R19008 gnd.n1207 gnd.n1204 9.3005
R19009 gnd.n5465 gnd.n5464 9.3005
R19010 gnd.n5521 gnd.n1148 9.3005
R19011 gnd.n4523 gnd.n4518 9.3005
R19012 gnd.n4522 gnd.n4521 9.3005
R19013 gnd.n1498 gnd.n1495 9.3005
R19014 gnd.n4737 gnd.n1496 9.3005
R19015 gnd.n4736 gnd.n4733 9.3005
R19016 gnd.n4735 gnd.n4734 9.3005
R19017 gnd.n1473 gnd.n1472 9.3005
R19018 gnd.n4764 gnd.n4763 9.3005
R19019 gnd.n1458 gnd.n1457 9.3005
R19020 gnd.n4777 gnd.n4776 9.3005
R19021 gnd.n4778 gnd.n1437 9.3005
R19022 gnd.n4816 gnd.n1438 9.3005
R19023 gnd.n4815 gnd.n1439 9.3005
R19024 gnd.n4814 gnd.n1440 9.3005
R19025 gnd.n4781 gnd.n1441 9.3005
R19026 gnd.n4784 gnd.n4783 9.3005
R19027 gnd.n4785 gnd.n1364 9.3005
R19028 gnd.n4918 gnd.n1365 9.3005
R19029 gnd.n4917 gnd.n1366 9.3005
R19030 gnd.n4916 gnd.n1367 9.3005
R19031 gnd.n1408 gnd.n1368 9.3005
R19032 gnd.n4873 gnd.n4872 9.3005
R19033 gnd.n4877 gnd.n4876 9.3005
R19034 gnd.n4878 gnd.n1402 9.3005
R19035 gnd.n4893 gnd.n1403 9.3005
R19036 gnd.n4892 gnd.n1404 9.3005
R19037 gnd.n4891 gnd.n1405 9.3005
R19038 gnd.n4890 gnd.n4888 9.3005
R19039 gnd.n1406 gnd.n1324 9.3005
R19040 gnd.n4972 gnd.n1325 9.3005
R19041 gnd.n4971 gnd.n1326 9.3005
R19042 gnd.n4970 gnd.n4965 9.3005
R19043 gnd.n4969 gnd.n4966 9.3005
R19044 gnd.n1300 gnd.n1297 9.3005
R19045 gnd.n5006 gnd.n1298 9.3005
R19046 gnd.n5005 gnd.n5002 9.3005
R19047 gnd.n5004 gnd.n5003 9.3005
R19048 gnd.n1229 gnd.n1228 9.3005
R19049 gnd.n5354 gnd.n5350 9.3005
R19050 gnd.n5353 gnd.n5351 9.3005
R19051 gnd.n5352 gnd.n1209 9.3005
R19052 gnd.n5462 gnd.n1210 9.3005
R19053 gnd.n4587 gnd.n4517 9.3005
R19054 gnd.n4524 gnd.n4523 9.3005
R19055 gnd.n4522 gnd.n1497 9.3005
R19056 gnd.n4730 gnd.n1498 9.3005
R19057 gnd.n4731 gnd.n1496 9.3005
R19058 gnd.n4733 gnd.n4732 9.3005
R19059 gnd.n4734 gnd.n1480 9.3005
R19060 gnd.n1474 gnd.n1473 9.3005
R19061 gnd.n4763 gnd.n4762 9.3005
R19062 gnd.n4761 gnd.n1457 9.3005
R19063 gnd.n4777 gnd.n1456 9.3005
R19064 gnd.n4779 gnd.n4778 9.3005
R19065 gnd.n4780 gnd.n1438 9.3005
R19066 gnd.n4791 gnd.n1439 9.3005
R19067 gnd.n4790 gnd.n1440 9.3005
R19068 gnd.n4789 gnd.n4781 9.3005
R19069 gnd.n4788 gnd.n4784 9.3005
R19070 gnd.n4786 gnd.n4785 9.3005
R19071 gnd.n1409 gnd.n1365 9.3005
R19072 gnd.n4866 gnd.n1366 9.3005
R19073 gnd.n4867 gnd.n1367 9.3005
R19074 gnd.n4868 gnd.n1408 9.3005
R19075 gnd.n4872 gnd.n4871 9.3005
R19076 gnd.n4877 gnd.n1407 9.3005
R19077 gnd.n4879 gnd.n4878 9.3005
R19078 gnd.n4880 gnd.n1403 9.3005
R19079 gnd.n4883 gnd.n1404 9.3005
R19080 gnd.n4884 gnd.n1405 9.3005
R19081 gnd.n4888 gnd.n4887 9.3005
R19082 gnd.n4885 gnd.n1406 9.3005
R19083 gnd.n1327 gnd.n1325 9.3005
R19084 gnd.n4963 gnd.n1326 9.3005
R19085 gnd.n4965 gnd.n4964 9.3005
R19086 gnd.n4966 gnd.n1299 9.3005
R19087 gnd.n4998 gnd.n1300 9.3005
R19088 gnd.n4999 gnd.n1298 9.3005
R19089 gnd.n5002 gnd.n5001 9.3005
R19090 gnd.n5003 gnd.n1230 9.3005
R19091 gnd.n5348 gnd.n1229 9.3005
R19092 gnd.n5350 gnd.n5349 9.3005
R19093 gnd.n5351 gnd.n1211 9.3005
R19094 gnd.n5460 gnd.n1209 9.3005
R19095 gnd.n5462 gnd.n5461 9.3005
R19096 gnd.n4587 gnd.n4586 9.3005
R19097 gnd.n4591 gnd.n4590 9.3005
R19098 gnd.n4594 gnd.n4512 9.3005
R19099 gnd.n4595 gnd.n4511 9.3005
R19100 gnd.n4598 gnd.n4510 9.3005
R19101 gnd.n4599 gnd.n4509 9.3005
R19102 gnd.n4602 gnd.n4508 9.3005
R19103 gnd.n4603 gnd.n4507 9.3005
R19104 gnd.n4606 gnd.n4506 9.3005
R19105 gnd.n4607 gnd.n4505 9.3005
R19106 gnd.n4610 gnd.n4504 9.3005
R19107 gnd.n4611 gnd.n4503 9.3005
R19108 gnd.n4614 gnd.n4502 9.3005
R19109 gnd.n4615 gnd.n4501 9.3005
R19110 gnd.n4618 gnd.n4500 9.3005
R19111 gnd.n4619 gnd.n4499 9.3005
R19112 gnd.n4622 gnd.n4498 9.3005
R19113 gnd.n4623 gnd.n4497 9.3005
R19114 gnd.n4626 gnd.n4496 9.3005
R19115 gnd.n4627 gnd.n4495 9.3005
R19116 gnd.n4630 gnd.n4494 9.3005
R19117 gnd.n4634 gnd.n4490 9.3005
R19118 gnd.n4635 gnd.n4489 9.3005
R19119 gnd.n4638 gnd.n4488 9.3005
R19120 gnd.n4639 gnd.n4487 9.3005
R19121 gnd.n4642 gnd.n4486 9.3005
R19122 gnd.n4643 gnd.n4485 9.3005
R19123 gnd.n4646 gnd.n4484 9.3005
R19124 gnd.n4647 gnd.n4483 9.3005
R19125 gnd.n4650 gnd.n4482 9.3005
R19126 gnd.n4651 gnd.n4481 9.3005
R19127 gnd.n4654 gnd.n4480 9.3005
R19128 gnd.n4655 gnd.n4479 9.3005
R19129 gnd.n4658 gnd.n4478 9.3005
R19130 gnd.n4659 gnd.n4477 9.3005
R19131 gnd.n4662 gnd.n4476 9.3005
R19132 gnd.n4663 gnd.n4475 9.3005
R19133 gnd.n4666 gnd.n4474 9.3005
R19134 gnd.n4667 gnd.n4473 9.3005
R19135 gnd.n4670 gnd.n4472 9.3005
R19136 gnd.n4672 gnd.n4469 9.3005
R19137 gnd.n4675 gnd.n4468 9.3005
R19138 gnd.n4676 gnd.n4467 9.3005
R19139 gnd.n4679 gnd.n4466 9.3005
R19140 gnd.n4680 gnd.n4465 9.3005
R19141 gnd.n4683 gnd.n4464 9.3005
R19142 gnd.n4684 gnd.n4463 9.3005
R19143 gnd.n4687 gnd.n4462 9.3005
R19144 gnd.n4688 gnd.n4461 9.3005
R19145 gnd.n4691 gnd.n4460 9.3005
R19146 gnd.n4692 gnd.n4459 9.3005
R19147 gnd.n4695 gnd.n4458 9.3005
R19148 gnd.n4696 gnd.n4457 9.3005
R19149 gnd.n4699 gnd.n4456 9.3005
R19150 gnd.n4700 gnd.n4455 9.3005
R19151 gnd.n4701 gnd.n4454 9.3005
R19152 gnd.n1514 gnd.n1513 9.3005
R19153 gnd.n4707 gnd.n4706 9.3005
R19154 gnd.n4631 gnd.n4491 9.3005
R19155 gnd.n4589 gnd.n4513 9.3005
R19156 gnd.n4712 gnd.n4709 9.3005
R19157 gnd.n4711 gnd.n4710 9.3005
R19158 gnd.n1487 gnd.n1486 9.3005
R19159 gnd.n4742 gnd.n4741 9.3005
R19160 gnd.n4743 gnd.n1485 9.3005
R19161 gnd.n4745 gnd.n4744 9.3005
R19162 gnd.n1465 gnd.n1464 9.3005
R19163 gnd.n4769 gnd.n4768 9.3005
R19164 gnd.n4770 gnd.n1463 9.3005
R19165 gnd.n4772 gnd.n4771 9.3005
R19166 gnd.n1429 gnd.n1428 9.3005
R19167 gnd.n4821 gnd.n4820 9.3005
R19168 gnd.n4822 gnd.n1427 9.3005
R19169 gnd.n4824 gnd.n4823 9.3005
R19170 gnd.n4825 gnd.n1349 9.3005
R19171 gnd.n4929 gnd.n4926 9.3005
R19172 gnd.n4928 gnd.n4927 9.3005
R19173 gnd.n1317 gnd.n1316 9.3005
R19174 gnd.n4977 gnd.n4976 9.3005
R19175 gnd.n4978 gnd.n1315 9.3005
R19176 gnd.n4982 gnd.n4979 9.3005
R19177 gnd.n4981 gnd.n4980 9.3005
R19178 gnd.n1289 gnd.n1288 9.3005
R19179 gnd.n5011 gnd.n5010 9.3005
R19180 gnd.n5012 gnd.n1287 9.3005
R19181 gnd.n5014 gnd.n5013 9.3005
R19182 gnd.n1220 gnd.n1219 9.3005
R19183 gnd.n5359 gnd.n5358 9.3005
R19184 gnd.n5360 gnd.n1218 9.3005
R19185 gnd.n5456 gnd.n5361 9.3005
R19186 gnd.n5455 gnd.n5454 9.3005
R19187 gnd.n4708 gnd.n1512 9.3005
R19188 gnd.n4925 gnd.n1348 9.3005
R19189 gnd.n4449 gnd.n4419 9.3005
R19190 gnd.n4448 gnd.n4420 9.3005
R19191 gnd.n4423 gnd.n4421 9.3005
R19192 gnd.n4444 gnd.n4424 9.3005
R19193 gnd.n4443 gnd.n4425 9.3005
R19194 gnd.n4442 gnd.n4426 9.3005
R19195 gnd.n4429 gnd.n4427 9.3005
R19196 gnd.n4438 gnd.n4430 9.3005
R19197 gnd.n4437 gnd.n4431 9.3005
R19198 gnd.n4436 gnd.n4432 9.3005
R19199 gnd.n4434 gnd.n4433 9.3005
R19200 gnd.n1447 gnd.n1446 9.3005
R19201 gnd.n4804 gnd.n4803 9.3005
R19202 gnd.n4805 gnd.n1445 9.3005
R19203 gnd.n4809 gnd.n4806 9.3005
R19204 gnd.n4808 gnd.n4807 9.3005
R19205 gnd.n4450 gnd.n4418 9.3005
R19206 gnd.n4415 gnd.n1557 9.3005
R19207 gnd.n2944 gnd.n1558 9.3005
R19208 gnd.n2946 gnd.n2945 9.3005
R19209 gnd.n2943 gnd.n1562 9.3005
R19210 gnd.n2942 gnd.n2941 9.3005
R19211 gnd.n1564 gnd.n1563 9.3005
R19212 gnd.n2935 gnd.n2934 9.3005
R19213 gnd.n2933 gnd.n1568 9.3005
R19214 gnd.n2932 gnd.n2931 9.3005
R19215 gnd.n1570 gnd.n1569 9.3005
R19216 gnd.n2925 gnd.n2924 9.3005
R19217 gnd.n2923 gnd.n1574 9.3005
R19218 gnd.n2922 gnd.n2921 9.3005
R19219 gnd.n1576 gnd.n1575 9.3005
R19220 gnd.n2915 gnd.n2914 9.3005
R19221 gnd.n2913 gnd.n1580 9.3005
R19222 gnd.n2912 gnd.n2911 9.3005
R19223 gnd.n1582 gnd.n1581 9.3005
R19224 gnd.n2905 gnd.n2904 9.3005
R19225 gnd.n2903 gnd.n1586 9.3005
R19226 gnd.n2902 gnd.n2901 9.3005
R19227 gnd.n1588 gnd.n1587 9.3005
R19228 gnd.n2895 gnd.n2894 9.3005
R19229 gnd.n2893 gnd.n1592 9.3005
R19230 gnd.n2892 gnd.n2891 9.3005
R19231 gnd.n1594 gnd.n1593 9.3005
R19232 gnd.n2885 gnd.n2884 9.3005
R19233 gnd.n2883 gnd.n1598 9.3005
R19234 gnd.n2882 gnd.n2881 9.3005
R19235 gnd.n1600 gnd.n1599 9.3005
R19236 gnd.n2875 gnd.n2874 9.3005
R19237 gnd.n2873 gnd.n1604 9.3005
R19238 gnd.n2872 gnd.n2871 9.3005
R19239 gnd.n1606 gnd.n1605 9.3005
R19240 gnd.n2865 gnd.n2864 9.3005
R19241 gnd.n2863 gnd.n1610 9.3005
R19242 gnd.n2862 gnd.n2861 9.3005
R19243 gnd.n1612 gnd.n1611 9.3005
R19244 gnd.n2855 gnd.n2854 9.3005
R19245 gnd.n2853 gnd.n1616 9.3005
R19246 gnd.n2852 gnd.n2851 9.3005
R19247 gnd.n1618 gnd.n1617 9.3005
R19248 gnd.n2845 gnd.n2844 9.3005
R19249 gnd.n2843 gnd.n1622 9.3005
R19250 gnd.n2842 gnd.n2841 9.3005
R19251 gnd.n1624 gnd.n1623 9.3005
R19252 gnd.n2835 gnd.n2834 9.3005
R19253 gnd.n2833 gnd.n1628 9.3005
R19254 gnd.n2832 gnd.n2831 9.3005
R19255 gnd.n1630 gnd.n1629 9.3005
R19256 gnd.n2825 gnd.n2824 9.3005
R19257 gnd.n2823 gnd.n1634 9.3005
R19258 gnd.n2822 gnd.n2821 9.3005
R19259 gnd.n1636 gnd.n1635 9.3005
R19260 gnd.n2815 gnd.n2814 9.3005
R19261 gnd.n2813 gnd.n1640 9.3005
R19262 gnd.n2812 gnd.n2811 9.3005
R19263 gnd.n1642 gnd.n1641 9.3005
R19264 gnd.n2805 gnd.n2804 9.3005
R19265 gnd.n2803 gnd.n1646 9.3005
R19266 gnd.n2802 gnd.n2801 9.3005
R19267 gnd.n1648 gnd.n1647 9.3005
R19268 gnd.n2795 gnd.n2794 9.3005
R19269 gnd.n2793 gnd.n1652 9.3005
R19270 gnd.n2792 gnd.n2791 9.3005
R19271 gnd.n1654 gnd.n1653 9.3005
R19272 gnd.n2785 gnd.n2784 9.3005
R19273 gnd.n2783 gnd.n1658 9.3005
R19274 gnd.n2782 gnd.n2781 9.3005
R19275 gnd.n1660 gnd.n1659 9.3005
R19276 gnd.n2775 gnd.n2774 9.3005
R19277 gnd.n2773 gnd.n1664 9.3005
R19278 gnd.n2772 gnd.n2771 9.3005
R19279 gnd.n1666 gnd.n1665 9.3005
R19280 gnd.n2765 gnd.n2764 9.3005
R19281 gnd.n2763 gnd.n1670 9.3005
R19282 gnd.n2762 gnd.n2761 9.3005
R19283 gnd.n1672 gnd.n1671 9.3005
R19284 gnd.n2755 gnd.n2754 9.3005
R19285 gnd.n2753 gnd.n1676 9.3005
R19286 gnd.n2752 gnd.n2751 9.3005
R19287 gnd.n1678 gnd.n1677 9.3005
R19288 gnd.n2745 gnd.n2744 9.3005
R19289 gnd.n2743 gnd.n1682 9.3005
R19290 gnd.n4417 gnd.n4416 9.3005
R19291 gnd.n6707 gnd.n422 9.3005
R19292 gnd.n5091 gnd.n5088 9.3005
R19293 gnd.n5093 gnd.n5092 9.3005
R19294 gnd.n5085 gnd.n5084 9.3005
R19295 gnd.n5112 gnd.n5111 9.3005
R19296 gnd.n5113 gnd.n5083 9.3005
R19297 gnd.n5115 gnd.n5114 9.3005
R19298 gnd.n5073 gnd.n5072 9.3005
R19299 gnd.n5133 gnd.n5132 9.3005
R19300 gnd.n5134 gnd.n5070 9.3005
R19301 gnd.n5137 gnd.n5136 9.3005
R19302 gnd.n5135 gnd.n5071 9.3005
R19303 gnd.n1083 gnd.n1081 9.3005
R19304 gnd.n5616 gnd.n5615 9.3005
R19305 gnd.n5614 gnd.n1082 9.3005
R19306 gnd.n5613 gnd.n5612 9.3005
R19307 gnd.n5611 gnd.n1084 9.3005
R19308 gnd.n5610 gnd.n5609 9.3005
R19309 gnd.n5608 gnd.n5600 9.3005
R19310 gnd.n5607 gnd.n5606 9.3005
R19311 gnd.n5605 gnd.n5601 9.3005
R19312 gnd.n5604 gnd.n5603 9.3005
R19313 gnd.n956 gnd.n955 9.3005
R19314 gnd.n5726 gnd.n5725 9.3005
R19315 gnd.n5727 gnd.n953 9.3005
R19316 gnd.n5729 gnd.n5728 9.3005
R19317 gnd.n5730 gnd.n952 9.3005
R19318 gnd.n5733 gnd.n5732 9.3005
R19319 gnd.n5734 gnd.n950 9.3005
R19320 gnd.n5737 gnd.n5736 9.3005
R19321 gnd.n5735 gnd.n951 9.3005
R19322 gnd.n891 gnd.n890 9.3005
R19323 gnd.n5809 gnd.n5808 9.3005
R19324 gnd.n5810 gnd.n888 9.3005
R19325 gnd.n5840 gnd.n5839 9.3005
R19326 gnd.n5838 gnd.n889 9.3005
R19327 gnd.n5837 gnd.n5836 9.3005
R19328 gnd.n5835 gnd.n5811 9.3005
R19329 gnd.n5834 gnd.n5833 9.3005
R19330 gnd.n5832 gnd.n5821 9.3005
R19331 gnd.n5831 gnd.n5830 9.3005
R19332 gnd.n5829 gnd.n5822 9.3005
R19333 gnd.n5828 gnd.n5827 9.3005
R19334 gnd.n5826 gnd.n5824 9.3005
R19335 gnd.n5825 gnd.n811 9.3005
R19336 gnd.n5954 gnd.n810 9.3005
R19337 gnd.n5956 gnd.n5955 9.3005
R19338 gnd.n5957 gnd.n808 9.3005
R19339 gnd.n6048 gnd.n6047 9.3005
R19340 gnd.n6046 gnd.n809 9.3005
R19341 gnd.n6045 gnd.n6044 9.3005
R19342 gnd.n6043 gnd.n5958 9.3005
R19343 gnd.n6042 gnd.n6041 9.3005
R19344 gnd.n6040 gnd.n5960 9.3005
R19345 gnd.n6039 gnd.n6038 9.3005
R19346 gnd.n6037 gnd.n5961 9.3005
R19347 gnd.n6036 gnd.n6035 9.3005
R19348 gnd.n6034 gnd.n5965 9.3005
R19349 gnd.n6033 gnd.n6032 9.3005
R19350 gnd.n6031 gnd.n5966 9.3005
R19351 gnd.n6030 gnd.n6029 9.3005
R19352 gnd.n6028 gnd.n6012 9.3005
R19353 gnd.n6027 gnd.n6026 9.3005
R19354 gnd.n6025 gnd.n6013 9.3005
R19355 gnd.n6024 gnd.n6023 9.3005
R19356 gnd.n6022 gnd.n6017 9.3005
R19357 gnd.n6021 gnd.n6020 9.3005
R19358 gnd.n6019 gnd.n6018 9.3005
R19359 gnd.n634 gnd.n633 9.3005
R19360 gnd.n6375 gnd.n6374 9.3005
R19361 gnd.n6376 gnd.n631 9.3005
R19362 gnd.n6379 gnd.n6378 9.3005
R19363 gnd.n6377 gnd.n632 9.3005
R19364 gnd.n609 gnd.n608 9.3005
R19365 gnd.n6405 gnd.n6404 9.3005
R19366 gnd.n6406 gnd.n606 9.3005
R19367 gnd.n6409 gnd.n6408 9.3005
R19368 gnd.n6407 gnd.n607 9.3005
R19369 gnd.n583 gnd.n582 9.3005
R19370 gnd.n6435 gnd.n6434 9.3005
R19371 gnd.n6436 gnd.n580 9.3005
R19372 gnd.n6439 gnd.n6438 9.3005
R19373 gnd.n6437 gnd.n581 9.3005
R19374 gnd.n5090 gnd.n5089 9.3005
R19375 gnd.n5333 gnd.n1240 9.3005
R19376 gnd.n4845 gnd.n4836 9.3005
R19377 gnd.n4844 gnd.n4843 9.3005
R19378 gnd.n4842 gnd.n4837 9.3005
R19379 gnd.n4841 gnd.n4840 9.3005
R19380 gnd.n1340 gnd.n1339 9.3005
R19381 gnd.n4934 gnd.n4933 9.3005
R19382 gnd.n4935 gnd.n1337 9.3005
R19383 gnd.n4938 gnd.n4937 9.3005
R19384 gnd.n4936 gnd.n1338 9.3005
R19385 gnd.n1307 gnd.n1306 9.3005
R19386 gnd.n4987 gnd.n4986 9.3005
R19387 gnd.n4988 gnd.n1304 9.3005
R19388 gnd.n4994 gnd.n4993 9.3005
R19389 gnd.n4992 gnd.n1305 9.3005
R19390 gnd.n4991 gnd.n4990 9.3005
R19391 gnd.n1236 gnd.n1234 9.3005
R19392 gnd.n5344 gnd.n5343 9.3005
R19393 gnd.n5342 gnd.n1235 9.3005
R19394 gnd.n5341 gnd.n5340 9.3005
R19395 gnd.n5339 gnd.n1237 9.3005
R19396 gnd.n5338 gnd.n5337 9.3005
R19397 gnd.n5311 gnd.n5310 9.3005
R19398 gnd.n5195 gnd.n5194 9.3005
R19399 gnd.n5305 gnd.n5304 9.3005
R19400 gnd.n5303 gnd.n5302 9.3005
R19401 gnd.n5209 gnd.n5208 9.3005
R19402 gnd.n5297 gnd.n5296 9.3005
R19403 gnd.n5295 gnd.n5294 9.3005
R19404 gnd.n5221 gnd.n5220 9.3005
R19405 gnd.n5289 gnd.n5288 9.3005
R19406 gnd.n5287 gnd.n5286 9.3005
R19407 gnd.n5232 gnd.n5231 9.3005
R19408 gnd.n5281 gnd.n5280 9.3005
R19409 gnd.n5279 gnd.n5278 9.3005
R19410 gnd.n5244 gnd.n5243 9.3005
R19411 gnd.n5273 gnd.n5272 9.3005
R19412 gnd.n5271 gnd.n5270 9.3005
R19413 gnd.n5262 gnd.n5260 9.3005
R19414 gnd.n5259 gnd.n1241 9.3005
R19415 gnd.n5313 gnd.n5312 9.3005
R19416 gnd.n5335 gnd.n5334 9.3005
R19417 gnd.n5261 gnd.n1242 9.3005
R19418 gnd.n5269 gnd.n5268 9.3005
R19419 gnd.n5248 gnd.n5247 9.3005
R19420 gnd.n5275 gnd.n5274 9.3005
R19421 gnd.n5277 gnd.n5276 9.3005
R19422 gnd.n5238 gnd.n5237 9.3005
R19423 gnd.n5283 gnd.n5282 9.3005
R19424 gnd.n5285 gnd.n5284 9.3005
R19425 gnd.n5225 gnd.n5224 9.3005
R19426 gnd.n5291 gnd.n5290 9.3005
R19427 gnd.n5293 gnd.n5292 9.3005
R19428 gnd.n5215 gnd.n5214 9.3005
R19429 gnd.n5299 gnd.n5298 9.3005
R19430 gnd.n5301 gnd.n5300 9.3005
R19431 gnd.n5202 gnd.n5201 9.3005
R19432 gnd.n5307 gnd.n5306 9.3005
R19433 gnd.n5309 gnd.n5308 9.3005
R19434 gnd.n5198 gnd.n1272 9.3005
R19435 gnd.n5314 gnd.n1271 9.3005
R19436 gnd.n5316 gnd.n5315 9.3005
R19437 gnd.n5318 gnd.n5317 9.3005
R19438 gnd.n5320 gnd.n5319 9.3005
R19439 gnd.n5321 gnd.n1265 9.3005
R19440 gnd.n5323 gnd.n5322 9.3005
R19441 gnd.n5324 gnd.n1264 9.3005
R19442 gnd.n5326 gnd.n5325 9.3005
R19443 gnd.n5327 gnd.n1263 9.3005
R19444 gnd.n5170 gnd.n5169 9.3005
R19445 gnd.n5168 gnd.n5047 9.3005
R19446 gnd.n5167 gnd.n5166 9.3005
R19447 gnd.n5165 gnd.n5049 9.3005
R19448 gnd.n5164 gnd.n5163 9.3005
R19449 gnd.n5162 gnd.n5053 9.3005
R19450 gnd.n5161 gnd.n5160 9.3005
R19451 gnd.n5159 gnd.n5054 9.3005
R19452 gnd.n5158 gnd.n5157 9.3005
R19453 gnd.n5156 gnd.n5058 9.3005
R19454 gnd.n5155 gnd.n5154 9.3005
R19455 gnd.n1076 gnd.n1075 9.3005
R19456 gnd.n5622 gnd.n5621 9.3005
R19457 gnd.n5623 gnd.n1074 9.3005
R19458 gnd.n5625 gnd.n5624 9.3005
R19459 gnd.n1003 gnd.n1002 9.3005
R19460 gnd.n5662 gnd.n5661 9.3005
R19461 gnd.n5663 gnd.n1001 9.3005
R19462 gnd.n5665 gnd.n5664 9.3005
R19463 gnd.n966 gnd.n965 9.3005
R19464 gnd.n5717 gnd.n5716 9.3005
R19465 gnd.n5718 gnd.n963 9.3005
R19466 gnd.n5721 gnd.n5720 9.3005
R19467 gnd.n5719 gnd.n964 9.3005
R19468 gnd.n931 gnd.n930 9.3005
R19469 gnd.n5759 gnd.n5758 9.3005
R19470 gnd.n5760 gnd.n929 9.3005
R19471 gnd.n5762 gnd.n5761 9.3005
R19472 gnd.n898 gnd.n897 9.3005
R19473 gnd.n5801 gnd.n5800 9.3005
R19474 gnd.n5802 gnd.n896 9.3005
R19475 gnd.n5804 gnd.n5803 9.3005
R19476 gnd.n883 gnd.n882 9.3005
R19477 gnd.n5845 gnd.n5844 9.3005
R19478 gnd.n5846 gnd.n881 9.3005
R19479 gnd.n5848 gnd.n5847 9.3005
R19480 gnd.n853 gnd.n852 9.3005
R19481 gnd.n5894 gnd.n5893 9.3005
R19482 gnd.n5895 gnd.n850 9.3005
R19483 gnd.n5898 gnd.n5897 9.3005
R19484 gnd.n5896 gnd.n851 9.3005
R19485 gnd.n817 gnd.n816 9.3005
R19486 gnd.n5947 gnd.n5946 9.3005
R19487 gnd.n5948 gnd.n815 9.3005
R19488 gnd.n5950 gnd.n5949 9.3005
R19489 gnd.n792 gnd.n791 9.3005
R19490 gnd.n6072 gnd.n6071 9.3005
R19491 gnd.n6073 gnd.n790 9.3005
R19492 gnd.n6075 gnd.n6074 9.3005
R19493 gnd.n769 gnd.n768 9.3005
R19494 gnd.n6100 gnd.n6099 9.3005
R19495 gnd.n6101 gnd.n766 9.3005
R19496 gnd.n6104 gnd.n6103 9.3005
R19497 gnd.n6102 gnd.n767 9.3005
R19498 gnd.n739 gnd.n738 9.3005
R19499 gnd.n6135 gnd.n6134 9.3005
R19500 gnd.n6136 gnd.n737 9.3005
R19501 gnd.n6138 gnd.n6137 9.3005
R19502 gnd.n715 gnd.n714 9.3005
R19503 gnd.n6167 gnd.n6166 9.3005
R19504 gnd.n6168 gnd.n712 9.3005
R19505 gnd.n6177 gnd.n6176 9.3005
R19506 gnd.n6175 gnd.n713 9.3005
R19507 gnd.n6174 gnd.n6173 9.3005
R19508 gnd.n6172 gnd.n6169 9.3005
R19509 gnd.n643 gnd.n642 9.3005
R19510 gnd.n6366 gnd.n6365 9.3005
R19511 gnd.n6367 gnd.n640 9.3005
R19512 gnd.n6370 gnd.n6369 9.3005
R19513 gnd.n6368 gnd.n641 9.3005
R19514 gnd.n618 gnd.n617 9.3005
R19515 gnd.n6396 gnd.n6395 9.3005
R19516 gnd.n6397 gnd.n615 9.3005
R19517 gnd.n6400 gnd.n6399 9.3005
R19518 gnd.n6398 gnd.n616 9.3005
R19519 gnd.n593 gnd.n592 9.3005
R19520 gnd.n6426 gnd.n6425 9.3005
R19521 gnd.n6427 gnd.n590 9.3005
R19522 gnd.n6430 gnd.n6429 9.3005
R19523 gnd.n6428 gnd.n591 9.3005
R19524 gnd.n569 gnd.n568 9.3005
R19525 gnd.n6466 gnd.n6465 9.3005
R19526 gnd.n5048 gnd.n5046 9.3005
R19527 gnd.n6469 gnd.n6468 9.3005
R19528 gnd.n6472 gnd.n566 9.3005
R19529 gnd.n6476 gnd.n6475 9.3005
R19530 gnd.n6477 gnd.n565 9.3005
R19531 gnd.n6479 gnd.n6478 9.3005
R19532 gnd.n6482 gnd.n563 9.3005
R19533 gnd.n6467 gnd.n567 9.3005
R19534 gnd.n6700 gnd.n6699 9.3005
R19535 gnd.n452 gnd.n449 9.3005
R19536 gnd.n6536 gnd.n6535 9.3005
R19537 gnd.n6538 gnd.n6537 9.3005
R19538 gnd.n6525 gnd.n6524 9.3005
R19539 gnd.n6544 gnd.n6543 9.3005
R19540 gnd.n6546 gnd.n6545 9.3005
R19541 gnd.n6515 gnd.n6514 9.3005
R19542 gnd.n6552 gnd.n6551 9.3005
R19543 gnd.n6554 gnd.n6553 9.3005
R19544 gnd.n6505 gnd.n6504 9.3005
R19545 gnd.n6560 gnd.n6559 9.3005
R19546 gnd.n6562 gnd.n6561 9.3005
R19547 gnd.n6495 gnd.n6494 9.3005
R19548 gnd.n6568 gnd.n6567 9.3005
R19549 gnd.n6570 gnd.n6569 9.3005
R19550 gnd.n6491 gnd.n6488 9.3005
R19551 gnd.n6698 gnd.n456 9.3005
R19552 gnd.n454 gnd.n423 9.3005
R19553 gnd.n6575 gnd.n6574 9.3005
R19554 gnd.n6573 gnd.n564 9.3005
R19555 gnd.n6572 gnd.n6571 9.3005
R19556 gnd.n6489 gnd.n6487 9.3005
R19557 gnd.n6566 gnd.n6565 9.3005
R19558 gnd.n6564 gnd.n6563 9.3005
R19559 gnd.n6499 gnd.n6498 9.3005
R19560 gnd.n6558 gnd.n6557 9.3005
R19561 gnd.n6556 gnd.n6555 9.3005
R19562 gnd.n6511 gnd.n6510 9.3005
R19563 gnd.n6550 gnd.n6549 9.3005
R19564 gnd.n6548 gnd.n6547 9.3005
R19565 gnd.n6519 gnd.n6518 9.3005
R19566 gnd.n6542 gnd.n6541 9.3005
R19567 gnd.n6540 gnd.n6539 9.3005
R19568 gnd.n6531 gnd.n6530 9.3005
R19569 gnd.n6534 gnd.n445 9.3005
R19570 gnd.n6702 gnd.n6701 9.3005
R19571 gnd.n451 gnd.n450 9.3005
R19572 gnd.n455 gnd.n424 9.3005
R19573 gnd.n6709 gnd.n6708 9.3005
R19574 gnd.n6711 gnd.n421 9.3005
R19575 gnd.n380 gnd.n379 9.3005
R19576 gnd.n6747 gnd.n6746 9.3005
R19577 gnd.n6748 gnd.n377 9.3005
R19578 gnd.n6751 gnd.n6750 9.3005
R19579 gnd.n6749 gnd.n378 9.3005
R19580 gnd.n347 gnd.n346 9.3005
R19581 gnd.n6816 gnd.n6815 9.3005
R19582 gnd.n6817 gnd.n344 9.3005
R19583 gnd.n6820 gnd.n6819 9.3005
R19584 gnd.n6818 gnd.n345 9.3005
R19585 gnd.n318 gnd.n317 9.3005
R19586 gnd.n6852 gnd.n6851 9.3005
R19587 gnd.n6853 gnd.n315 9.3005
R19588 gnd.n6863 gnd.n6862 9.3005
R19589 gnd.n6861 gnd.n316 9.3005
R19590 gnd.n6860 gnd.n6859 9.3005
R19591 gnd.n6858 gnd.n6854 9.3005
R19592 gnd.n6857 gnd.n6856 9.3005
R19593 gnd.n6855 gnd.n63 9.3005
R19594 gnd.n6713 gnd.n6712 9.3005
R19595 gnd.n7330 gnd.n64 9.3005
R19596 gnd.t297 gnd.n3154 9.24152
R19597 gnd.n4370 gnd.t113 9.24152
R19598 gnd.t95 gnd.n3025 9.24152
R19599 gnd.n1294 gnd.t185 9.24152
R19600 gnd.n6789 gnd.t192 9.24152
R19601 gnd.t163 gnd.t297 8.92286
R19602 gnd.n5714 gnd.n5713 8.92286
R19603 gnd.n942 gnd.n941 8.92286
R19604 gnd.t142 gnd.n903 8.92286
R19605 gnd.t144 gnd.n894 8.92286
R19606 gnd.n5891 gnd.n5890 8.92286
R19607 gnd.n5916 gnd.n824 8.92286
R19608 gnd.n6090 gnd.t11 8.92286
R19609 gnd.n5974 gnd.t13 8.92286
R19610 gnd.n6123 gnd.n749 8.92286
R19611 gnd.n6010 gnd.n6009 8.92286
R19612 gnd.n4224 gnd.n4199 8.92171
R19613 gnd.n4192 gnd.n4167 8.92171
R19614 gnd.n4160 gnd.n4135 8.92171
R19615 gnd.n4129 gnd.n4104 8.92171
R19616 gnd.n4097 gnd.n4072 8.92171
R19617 gnd.n4065 gnd.n4040 8.92171
R19618 gnd.n4033 gnd.n4008 8.92171
R19619 gnd.n4002 gnd.n3977 8.92171
R19620 gnd.n6211 gnd.n6193 8.72777
R19621 gnd.n3798 gnd.t299 8.60421
R19622 gnd.n4703 gnd.n1516 8.60421
R19623 gnd.n5818 gnd.t159 8.60421
R19624 gnd.n5943 gnd.t147 8.60421
R19625 gnd.n7253 gnd.n7040 8.60421
R19626 gnd.n3218 gnd.n3206 8.43656
R19627 gnd.n38 gnd.n26 8.43656
R19628 gnd.n4412 gnd.n2950 8.28555
R19629 gnd.n999 gnd.n991 8.28555
R19630 gnd.n5743 gnd.n949 8.28555
R19631 gnd.n5851 gnd.n862 8.28555
R19632 gnd.n6059 gnd.n802 8.28555
R19633 gnd.n6114 gnd.n756 8.28555
R19634 gnd.n6002 gnd.n6001 8.28555
R19635 gnd.n4225 gnd.n4197 8.14595
R19636 gnd.n4193 gnd.n4165 8.14595
R19637 gnd.n4161 gnd.n4133 8.14595
R19638 gnd.n4130 gnd.n4102 8.14595
R19639 gnd.n4098 gnd.n4070 8.14595
R19640 gnd.n4066 gnd.n4038 8.14595
R19641 gnd.n4034 gnd.n4006 8.14595
R19642 gnd.n4003 gnd.n3975 8.14595
R19643 gnd.n4846 gnd.n0 8.10675
R19644 gnd.n7331 gnd.n7330 8.10675
R19645 gnd.n4230 gnd.n4229 7.97301
R19646 gnd.t305 gnd.n3313 7.9669
R19647 gnd.t20 gnd.t306 7.9669
R19648 gnd.n7331 gnd.n62 7.78567
R19649 gnd.n6698 gnd.n454 7.75808
R19650 gnd.n5260 gnd.n5259 7.75808
R19651 gnd.n7256 gnd.n182 7.75808
R19652 gnd.n4545 gnd.n4544 7.75808
R19653 gnd.n5667 gnd.n999 7.64824
R19654 gnd.n5743 gnd.n5740 7.64824
R19655 gnd.n5850 gnd.t155 7.64824
R19656 gnd.n5851 gnd.n5850 7.64824
R19657 gnd.n6059 gnd.n6058 7.64824
R19658 gnd.n6058 gnd.t10 7.64824
R19659 gnd.n6106 gnd.n756 7.64824
R19660 gnd.n3243 gnd.n3242 7.53171
R19661 gnd.n3707 gnd.t295 7.32958
R19662 gnd.n1027 gnd.n1026 7.30353
R19663 gnd.n6210 gnd.n6209 7.30353
R19664 gnd.n3667 gnd.n3386 7.01093
R19665 gnd.n3389 gnd.n3387 7.01093
R19666 gnd.n3677 gnd.n3676 7.01093
R19667 gnd.n3688 gnd.n3370 7.01093
R19668 gnd.n3687 gnd.n3373 7.01093
R19669 gnd.n3698 gnd.n3361 7.01093
R19670 gnd.n3364 gnd.n3362 7.01093
R19671 gnd.n3708 gnd.n3707 7.01093
R19672 gnd.n3718 gnd.n3342 7.01093
R19673 gnd.n3717 gnd.n3345 7.01093
R19674 gnd.n3726 gnd.n3336 7.01093
R19675 gnd.n3738 gnd.n3326 7.01093
R19676 gnd.n3748 gnd.n3311 7.01093
R19677 gnd.n3764 gnd.n3763 7.01093
R19678 gnd.n3313 gnd.n3250 7.01093
R19679 gnd.n3818 gnd.n3251 7.01093
R19680 gnd.n3812 gnd.n3811 7.01093
R19681 gnd.n3300 gnd.n3262 7.01093
R19682 gnd.n3804 gnd.n3273 7.01093
R19683 gnd.n3291 gnd.n3286 7.01093
R19684 gnd.n3798 gnd.n3797 7.01093
R19685 gnd.n3844 gnd.n3189 7.01093
R19686 gnd.n3843 gnd.n3842 7.01093
R19687 gnd.n3855 gnd.n3854 7.01093
R19688 gnd.n3182 gnd.n3174 7.01093
R19689 gnd.n3884 gnd.n3162 7.01093
R19690 gnd.n3883 gnd.n3165 7.01093
R19691 gnd.n3894 gnd.n3154 7.01093
R19692 gnd.n3155 gnd.n3143 7.01093
R19693 gnd.n3907 gnd.n3144 7.01093
R19694 gnd.n3940 gnd.n3136 7.01093
R19695 gnd.n3939 gnd.n2950 7.01093
R19696 gnd.n4405 gnd.n4404 7.01093
R19697 gnd.n3930 gnd.n3929 7.01093
R19698 gnd.n4398 gnd.n2971 7.01093
R19699 gnd.n4397 gnd.n2974 7.01093
R19700 gnd.n3922 gnd.n2983 7.01093
R19701 gnd.n4391 gnd.n4390 7.01093
R19702 gnd.n4384 gnd.n2996 7.01093
R19703 gnd.n4383 gnd.n2999 7.01093
R19704 gnd.n4262 gnd.n3008 7.01093
R19705 gnd.n4377 gnd.n4376 7.01093
R19706 gnd.n4243 gnd.n3011 7.01093
R19707 gnd.n4370 gnd.n3022 7.01093
R19708 gnd.n4369 gnd.n3025 7.01093
R19709 gnd.n4273 gnd.n3033 7.01093
R19710 gnd.n4363 gnd.n4362 7.01093
R19711 gnd.n5713 gnd.n971 7.01093
R19712 gnd.n942 gnd.n935 7.01093
R19713 gnd.n5890 gnd.n858 7.01093
R19714 gnd.n5916 gnd.n5915 7.01093
R19715 gnd.n6123 gnd.n6122 7.01093
R19716 gnd.n6009 gnd.n719 7.01093
R19717 gnd.t105 gnd.n707 7.01093
R19718 gnd.n3345 gnd.t293 6.69227
R19719 gnd.n3165 gnd.t163 6.69227
R19720 gnd.t304 gnd.n4254 6.69227
R19721 gnd.t309 gnd.n992 6.69227
R19722 gnd.t145 gnd.n6179 6.69227
R19723 gnd.n6343 gnd.n6342 6.5566
R19724 gnd.n5533 gnd.n5532 6.5566
R19725 gnd.n1143 gnd.n1089 6.5566
R19726 gnd.n6221 gnd.n6220 6.5566
R19727 gnd.n5659 gnd.n5658 6.37362
R19728 gnd.n5640 gnd.t42 6.37362
R19729 gnd.n5756 gnd.t141 6.37362
R19730 gnd.n910 gnd.n909 6.37362
R19731 gnd.n5865 gnd.t155 6.37362
R19732 gnd.t10 gnd.n6057 6.37362
R19733 gnd.n6097 gnd.n6096 6.37362
R19734 gnd.n6132 gnd.t12 6.37362
R19735 gnd.n6180 gnd.t23 6.37362
R19736 gnd.n6282 gnd.n654 6.37362
R19737 gnd.n5268 gnd.n5265 6.20656
R19738 gnd.n450 gnd.n448 6.20656
R19739 gnd.t7 gnd.n3774 6.05496
R19740 gnd.n3775 gnd.t292 6.05496
R19741 gnd.t311 gnd.n3189 6.05496
R19742 gnd.n3949 gnd.t291 6.05496
R19743 gnd.t27 gnd.n1508 6.05496
R19744 gnd.t159 gnd.n858 6.05496
R19745 gnd.n5915 gnd.t147 6.05496
R19746 gnd.n176 gnd.t31 6.05496
R19747 gnd.n4227 gnd.n4197 5.81868
R19748 gnd.n4195 gnd.n4165 5.81868
R19749 gnd.n4163 gnd.n4133 5.81868
R19750 gnd.n4132 gnd.n4102 5.81868
R19751 gnd.n4100 gnd.n4070 5.81868
R19752 gnd.n4068 gnd.n4038 5.81868
R19753 gnd.n4036 gnd.n4006 5.81868
R19754 gnd.n4005 gnd.n3975 5.81868
R19755 gnd.n981 gnd.n960 5.73631
R19756 gnd.n5704 gnd.n980 5.73631
R19757 gnd.n848 gnd.n836 5.73631
R19758 gnd.n841 gnd.n838 5.73631
R19759 gnd.n6141 gnd.n733 5.73631
R19760 gnd.n6152 gnd.n724 5.73631
R19761 gnd.n6010 gnd.t105 5.73631
R19762 gnd.n6347 gnd.n525 5.62001
R19763 gnd.n5528 gnd.n5525 5.62001
R19764 gnd.n5525 gnd.n1147 5.62001
R19765 gnd.n6216 gnd.n525 5.62001
R19766 gnd.n3526 gnd.n3521 5.4308
R19767 gnd.n3114 gnd.n3112 5.4308
R19768 gnd.n3842 gnd.t290 5.41765
R19769 gnd.t298 gnd.n3865 5.41765
R19770 gnd.t167 gnd.n2960 5.41765
R19771 gnd.n5681 gnd.t157 5.41765
R19772 gnd.n744 gnd.t2 5.41765
R19773 gnd.n5806 gnd.n894 5.09899
R19774 gnd.n5785 gnd.n5782 5.09899
R19775 gnd.n6077 gnd.n788 5.09899
R19776 gnd.n6090 gnd.n6089 5.09899
R19777 gnd.t57 gnd.n698 5.09899
R19778 gnd.n4225 gnd.n4224 5.04292
R19779 gnd.n4193 gnd.n4192 5.04292
R19780 gnd.n4161 gnd.n4160 5.04292
R19781 gnd.n4130 gnd.n4129 5.04292
R19782 gnd.n4098 gnd.n4097 5.04292
R19783 gnd.n4066 gnd.n4065 5.04292
R19784 gnd.n4034 gnd.n4033 5.04292
R19785 gnd.n4003 gnd.n4002 5.04292
R19786 gnd.n3805 gnd.t301 4.78034
R19787 gnd.n3144 gnd.t302 4.78034
R19788 gnd.t313 gnd.n5117 4.78034
R19789 gnd.t157 gnd.n980 4.78034
R19790 gnd.t2 gnd.n733 4.78034
R19791 gnd.n6350 gnd.t20 4.78034
R19792 gnd.n6412 gnd.t317 4.78034
R19793 gnd.n3247 gnd.n3244 4.74817
R19794 gnd.n3297 gnd.n3195 4.74817
R19795 gnd.n3284 gnd.n3194 4.74817
R19796 gnd.n3193 gnd.n3192 4.74817
R19797 gnd.n3293 gnd.n3244 4.74817
R19798 gnd.n3294 gnd.n3195 4.74817
R19799 gnd.n3296 gnd.n3194 4.74817
R19800 gnd.n3283 gnd.n3193 4.74817
R19801 gnd.n6875 gnd.n82 4.74817
R19802 gnd.n6909 gnd.n81 4.74817
R19803 gnd.n6905 gnd.n80 4.74817
R19804 gnd.n7323 gnd.n75 4.74817
R19805 gnd.n7321 gnd.n76 4.74817
R19806 gnd.n305 gnd.n82 4.74817
R19807 gnd.n6874 gnd.n81 4.74817
R19808 gnd.n6910 gnd.n80 4.74817
R19809 gnd.n6904 gnd.n75 4.74817
R19810 gnd.n7322 gnd.n7321 4.74817
R19811 gnd.n1414 gnd.n1412 4.74817
R19812 gnd.n4861 gnd.n4859 4.74817
R19813 gnd.n4906 gnd.n1381 4.74817
R19814 gnd.n4904 gnd.n4903 4.74817
R19815 gnd.n1398 gnd.n1395 4.74817
R19816 gnd.n6888 gnd.n293 4.74817
R19817 gnd.n6899 gnd.n6890 4.74817
R19818 gnd.n6897 gnd.n6896 4.74817
R19819 gnd.n6892 gnd.n6891 4.74817
R19820 gnd.n7001 gnd.n262 4.74817
R19821 gnd.n6773 gnd.n293 4.74817
R19822 gnd.n6890 gnd.n6889 4.74817
R19823 gnd.n6898 gnd.n6897 4.74817
R19824 gnd.n6893 gnd.n6892 4.74817
R19825 gnd.n264 gnd.n262 4.74817
R19826 gnd.n4924 gnd.n4923 4.74817
R19827 gnd.n4911 gnd.n1354 4.74817
R19828 gnd.n1375 gnd.n1353 4.74817
R19829 gnd.n4897 gnd.n1352 4.74817
R19830 gnd.n1391 gnd.n1351 4.74817
R19831 gnd.n4924 gnd.n1355 4.74817
R19832 gnd.n4922 gnd.n1354 4.74817
R19833 gnd.n4912 gnd.n1353 4.74817
R19834 gnd.n1374 gnd.n1352 4.74817
R19835 gnd.n4898 gnd.n1351 4.74817
R19836 gnd.n4857 gnd.n1412 4.74817
R19837 gnd.n4859 gnd.n4858 4.74817
R19838 gnd.n4860 gnd.n1381 4.74817
R19839 gnd.n4905 gnd.n4904 4.74817
R19840 gnd.n1395 gnd.n1382 4.74817
R19841 gnd.n3242 gnd.n3241 4.74296
R19842 gnd.n62 gnd.n61 4.74296
R19843 gnd.n3218 gnd.n3217 4.7074
R19844 gnd.n3230 gnd.n3229 4.7074
R19845 gnd.n38 gnd.n37 4.7074
R19846 gnd.n50 gnd.n49 4.7074
R19847 gnd.n3242 gnd.n3230 4.65959
R19848 gnd.n62 gnd.n50 4.65959
R19849 gnd.n6640 gnd.n527 4.6132
R19850 gnd.n5523 gnd.n5522 4.6132
R19851 gnd.n5694 gnd.n959 4.46168
R19852 gnd.n5705 gnd.t4 4.46168
R19853 gnd.n5683 gnd.n5682 4.46168
R19854 gnd.n5901 gnd.n845 4.46168
R19855 gnd.n5923 gnd.n5922 4.46168
R19856 gnd.n6131 gnd.n6130 4.46168
R19857 gnd.t156 gnd.n6140 4.46168
R19858 gnd.n6150 gnd.n6149 4.46168
R19859 gnd.n6206 gnd.n6193 4.46111
R19860 gnd.n4210 gnd.n4206 4.38594
R19861 gnd.n4178 gnd.n4174 4.38594
R19862 gnd.n4146 gnd.n4142 4.38594
R19863 gnd.n4115 gnd.n4111 4.38594
R19864 gnd.n4083 gnd.n4079 4.38594
R19865 gnd.n4051 gnd.n4047 4.38594
R19866 gnd.n4019 gnd.n4015 4.38594
R19867 gnd.n3988 gnd.n3984 4.38594
R19868 gnd.n4221 gnd.n4199 4.26717
R19869 gnd.n4189 gnd.n4167 4.26717
R19870 gnd.n4157 gnd.n4135 4.26717
R19871 gnd.n4126 gnd.n4104 4.26717
R19872 gnd.n4094 gnd.n4072 4.26717
R19873 gnd.n4062 gnd.n4040 4.26717
R19874 gnd.n4030 gnd.n4008 4.26717
R19875 gnd.n3999 gnd.n3977 4.26717
R19876 gnd.n3749 gnd.t303 4.14303
R19877 gnd.t300 gnd.n2974 4.14303
R19878 gnd.n5027 gnd.t49 4.14303
R19879 gnd.n6726 gnd.t35 4.14303
R19880 gnd.n4229 gnd.n4228 4.08274
R19881 gnd.n6342 gnd.n6341 4.05904
R19882 gnd.n5534 gnd.n5533 4.05904
R19883 gnd.n1140 gnd.n1089 4.05904
R19884 gnd.n6222 gnd.n6221 4.05904
R19885 gnd.n15 gnd.n7 3.99943
R19886 gnd.n5598 gnd.n5597 3.82437
R19887 gnd.n981 gnd.t17 3.82437
R19888 gnd.n5740 gnd.t143 3.82437
R19889 gnd.n5798 gnd.n5797 3.82437
R19890 gnd.n5857 gnd.n871 3.82437
R19891 gnd.n6069 gnd.n6068 3.82437
R19892 gnd.n5977 gnd.n5976 3.82437
R19893 gnd.t308 gnd.n6106 3.82437
R19894 gnd.n701 gnd.n700 3.82437
R19895 gnd.n3822 gnd.n3243 3.81325
R19896 gnd.n3230 gnd.n3218 3.72967
R19897 gnd.n50 gnd.n38 3.72967
R19898 gnd.n4229 gnd.n4101 3.70378
R19899 gnd.n15 gnd.n14 3.60163
R19900 gnd.n4220 gnd.n4201 3.49141
R19901 gnd.n4188 gnd.n4169 3.49141
R19902 gnd.n4156 gnd.n4137 3.49141
R19903 gnd.n4125 gnd.n4106 3.49141
R19904 gnd.n4093 gnd.n4074 3.49141
R19905 gnd.n4061 gnd.n4042 3.49141
R19906 gnd.n4029 gnd.n4010 3.49141
R19907 gnd.n3998 gnd.n3979 3.49141
R19908 gnd.n6658 gnd.n6657 3.29747
R19909 gnd.n6657 gnd.n6656 3.29747
R19910 gnd.n7220 gnd.n7217 3.29747
R19911 gnd.n7221 gnd.n7220 3.29747
R19912 gnd.n4672 gnd.n4671 3.29747
R19913 gnd.n4671 gnd.n4670 3.29747
R19914 gnd.n5394 gnd.n5389 3.29747
R19915 gnd.n5419 gnd.n5394 3.29747
R19916 gnd.n5640 gnd.n968 3.18706
R19917 gnd.n5859 gnd.t136 3.18706
R19918 gnd.n5882 gnd.n855 3.18706
R19919 gnd.n5937 gnd.n5936 3.18706
R19920 gnd.n6051 gnd.t0 3.18706
R19921 gnd.n6180 gnd.n707 3.18706
R19922 gnd.n3328 gnd.t303 2.8684
R19923 gnd.n1072 gnd.t139 2.8684
R19924 gnd.t42 gnd.t309 2.8684
R19925 gnd.t23 gnd.t145 2.8684
R19926 gnd.t306 gnd.n645 2.8684
R19927 gnd.n3231 gnd.t212 2.82907
R19928 gnd.n3231 gnd.t272 2.82907
R19929 gnd.n3233 gnd.t191 2.82907
R19930 gnd.n3233 gnd.t226 2.82907
R19931 gnd.n3235 gnd.t243 2.82907
R19932 gnd.n3235 gnd.t232 2.82907
R19933 gnd.n3237 gnd.t230 2.82907
R19934 gnd.n3237 gnd.t221 2.82907
R19935 gnd.n3239 gnd.t235 2.82907
R19936 gnd.n3239 gnd.t261 2.82907
R19937 gnd.n3196 gnd.t237 2.82907
R19938 gnd.n3196 gnd.t252 2.82907
R19939 gnd.n3198 gnd.t258 2.82907
R19940 gnd.n3198 gnd.t214 2.82907
R19941 gnd.n3200 gnd.t251 2.82907
R19942 gnd.n3200 gnd.t247 2.82907
R19943 gnd.n3202 gnd.t284 2.82907
R19944 gnd.n3202 gnd.t275 2.82907
R19945 gnd.n3204 gnd.t219 2.82907
R19946 gnd.n3204 gnd.t256 2.82907
R19947 gnd.n3207 gnd.t287 2.82907
R19948 gnd.n3207 gnd.t196 2.82907
R19949 gnd.n3209 gnd.t199 2.82907
R19950 gnd.n3209 gnd.t180 2.82907
R19951 gnd.n3211 gnd.t260 2.82907
R19952 gnd.n3211 gnd.t288 2.82907
R19953 gnd.n3213 gnd.t282 2.82907
R19954 gnd.n3213 gnd.t201 2.82907
R19955 gnd.n3215 gnd.t276 2.82907
R19956 gnd.n3215 gnd.t259 2.82907
R19957 gnd.n3219 gnd.t249 2.82907
R19958 gnd.n3219 gnd.t215 2.82907
R19959 gnd.n3221 gnd.t236 2.82907
R19960 gnd.n3221 gnd.t263 2.82907
R19961 gnd.n3223 gnd.t281 2.82907
R19962 gnd.n3223 gnd.t270 2.82907
R19963 gnd.n3225 gnd.t268 2.82907
R19964 gnd.n3225 gnd.t255 2.82907
R19965 gnd.n3227 gnd.t273 2.82907
R19966 gnd.n3227 gnd.t208 2.82907
R19967 gnd.n59 gnd.t239 2.82907
R19968 gnd.n59 gnd.t220 2.82907
R19969 gnd.n57 gnd.t188 2.82907
R19970 gnd.n57 gnd.t206 2.82907
R19971 gnd.n55 gnd.t198 2.82907
R19972 gnd.n55 gnd.t223 2.82907
R19973 gnd.n53 gnd.t204 2.82907
R19974 gnd.n53 gnd.t269 2.82907
R19975 gnd.n51 gnd.t248 2.82907
R19976 gnd.n51 gnd.t184 2.82907
R19977 gnd.n24 gnd.t289 2.82907
R19978 gnd.n24 gnd.t210 2.82907
R19979 gnd.n22 gnd.t194 2.82907
R19980 gnd.n22 gnd.t209 2.82907
R19981 gnd.n20 gnd.t267 2.82907
R19982 gnd.n20 gnd.t244 2.82907
R19983 gnd.n18 gnd.t234 2.82907
R19984 gnd.n18 gnd.t178 2.82907
R19985 gnd.n16 gnd.t280 2.82907
R19986 gnd.n16 gnd.t224 2.82907
R19987 gnd.n35 gnd.t250 2.82907
R19988 gnd.n35 gnd.t177 2.82907
R19989 gnd.n33 gnd.t173 2.82907
R19990 gnd.n33 gnd.t264 2.82907
R19991 gnd.n31 gnd.t271 2.82907
R19992 gnd.n31 gnd.t278 2.82907
R19993 gnd.n29 gnd.t277 2.82907
R19994 gnd.n29 gnd.t175 2.82907
R19995 gnd.n27 gnd.t171 2.82907
R19996 gnd.n27 gnd.t189 2.82907
R19997 gnd.n47 gnd.t279 2.82907
R19998 gnd.n47 gnd.t254 2.82907
R19999 gnd.n45 gnd.t233 2.82907
R20000 gnd.n45 gnd.t245 2.82907
R20001 gnd.n43 gnd.t246 2.82907
R20002 gnd.n43 gnd.t257 2.82907
R20003 gnd.n41 gnd.t240 2.82907
R20004 gnd.n41 gnd.t213 2.82907
R20005 gnd.n39 gnd.t286 2.82907
R20006 gnd.n39 gnd.t228 2.82907
R20007 gnd.n4217 gnd.n4216 2.71565
R20008 gnd.n4185 gnd.n4184 2.71565
R20009 gnd.n4153 gnd.n4152 2.71565
R20010 gnd.n4122 gnd.n4121 2.71565
R20011 gnd.n4090 gnd.n4089 2.71565
R20012 gnd.n4058 gnd.n4057 2.71565
R20013 gnd.n4026 gnd.n4025 2.71565
R20014 gnd.n3995 gnd.n3994 2.71565
R20015 gnd.n5668 gnd.t68 2.54975
R20016 gnd.n5674 gnd.n992 2.54975
R20017 gnd.n5764 gnd.n927 2.54975
R20018 gnd.n5884 gnd.n5883 2.54975
R20019 gnd.t1 gnd.n5882 2.54975
R20020 gnd.n5819 gnd.t14 2.54975
R20021 gnd.n5944 gnd.t9 2.54975
R20022 gnd.n5936 gnd.t169 2.54975
R20023 gnd.n5952 gnd.n813 2.54975
R20024 gnd.n6113 gnd.n758 2.54975
R20025 gnd.n6179 gnd.n709 2.54975
R20026 gnd.n6002 gnd.t57 2.54975
R20027 gnd.n3822 gnd.n3244 2.27742
R20028 gnd.n3822 gnd.n3195 2.27742
R20029 gnd.n3822 gnd.n3194 2.27742
R20030 gnd.n3822 gnd.n3193 2.27742
R20031 gnd.n7320 gnd.n82 2.27742
R20032 gnd.n7320 gnd.n81 2.27742
R20033 gnd.n7320 gnd.n80 2.27742
R20034 gnd.n7320 gnd.n75 2.27742
R20035 gnd.n7321 gnd.n7320 2.27742
R20036 gnd.n293 gnd.n79 2.27742
R20037 gnd.n6890 gnd.n79 2.27742
R20038 gnd.n6897 gnd.n79 2.27742
R20039 gnd.n6892 gnd.n79 2.27742
R20040 gnd.n262 gnd.n79 2.27742
R20041 gnd.n4925 gnd.n4924 2.27742
R20042 gnd.n4925 gnd.n1354 2.27742
R20043 gnd.n4925 gnd.n1353 2.27742
R20044 gnd.n4925 gnd.n1352 2.27742
R20045 gnd.n4925 gnd.n1351 2.27742
R20046 gnd.n1412 gnd.n1350 2.27742
R20047 gnd.n4859 gnd.n1350 2.27742
R20048 gnd.n1381 gnd.n1350 2.27742
R20049 gnd.n4904 gnd.n1350 2.27742
R20050 gnd.n1395 gnd.n1350 2.27742
R20051 gnd.n3676 gnd.t60 2.23109
R20052 gnd.n3299 gnd.t301 2.23109
R20053 gnd.n5842 gnd.t5 2.23109
R20054 gnd.t315 gnd.n6050 2.23109
R20055 gnd.n4213 gnd.n4203 1.93989
R20056 gnd.n4181 gnd.n4171 1.93989
R20057 gnd.n4149 gnd.n4139 1.93989
R20058 gnd.n4118 gnd.n4108 1.93989
R20059 gnd.n4086 gnd.n4076 1.93989
R20060 gnd.n4054 gnd.n4044 1.93989
R20061 gnd.n4022 gnd.n4012 1.93989
R20062 gnd.n3991 gnd.n3981 1.93989
R20063 gnd.n5668 gnd.n996 1.91244
R20064 gnd.n5749 gnd.t135 1.91244
R20065 gnd.n916 gnd.t144 1.91244
R20066 gnd.n5866 gnd.n5865 1.91244
R20067 gnd.n6057 gnd.n794 1.91244
R20068 gnd.n787 gnd.t11 1.91244
R20069 gnd.n5985 gnd.t15 1.91244
R20070 gnd.n6189 gnd.n6188 1.91244
R20071 gnd.t161 gnd.n3687 1.59378
R20072 gnd.n3866 gnd.t298 1.59378
R20073 gnd.n3130 gnd.t167 1.59378
R20074 gnd.t153 gnd.n900 1.59378
R20075 gnd.n5975 gnd.t149 1.59378
R20076 gnd.n5693 gnd.t86 1.27512
R20077 gnd.n5756 gnd.n5755 1.27512
R20078 gnd.n5765 gnd.t135 1.27512
R20079 gnd.n5819 gnd.n5818 1.27512
R20080 gnd.n5944 gnd.n5943 1.27512
R20081 gnd.t15 gnd.n5984 1.27512
R20082 gnd.n6132 gnd.n741 1.27512
R20083 gnd.n6164 gnd.n6163 1.27512
R20084 gnd.n3529 gnd.n3521 1.16414
R20085 gnd.n4288 gnd.n3112 1.16414
R20086 gnd.n4212 gnd.n4205 1.16414
R20087 gnd.n4180 gnd.n4173 1.16414
R20088 gnd.n4148 gnd.n4141 1.16414
R20089 gnd.n4117 gnd.n4110 1.16414
R20090 gnd.n4085 gnd.n4078 1.16414
R20091 gnd.n4053 gnd.n4046 1.16414
R20092 gnd.n4021 gnd.n4014 1.16414
R20093 gnd.n3990 gnd.n3983 1.16414
R20094 gnd.n6640 gnd.n6639 0.970197
R20095 gnd.n5523 gnd.n1148 0.970197
R20096 gnd.n4196 gnd.n4164 0.962709
R20097 gnd.n4228 gnd.n4196 0.962709
R20098 gnd.n4069 gnd.n4037 0.962709
R20099 gnd.n4101 gnd.n4069 0.962709
R20100 gnd.n3775 gnd.t7 0.956468
R20101 gnd.n4411 gnd.t291 0.956468
R20102 gnd.n1482 gnd.t181 0.956468
R20103 gnd.n4759 gnd.t218 0.956468
R20104 gnd.n4960 gnd.t211 0.956468
R20105 gnd.n4967 gnd.t195 0.956468
R20106 gnd.n5152 gnd.t151 0.956468
R20107 gnd.t5 gnd.t136 0.956468
R20108 gnd.t0 gnd.t315 0.956468
R20109 gnd.n6381 gnd.t137 0.956468
R20110 gnd.n6796 gnd.t170 0.956468
R20111 gnd.t183 gnd.n333 0.956468
R20112 gnd.n6973 gnd.t176 0.956468
R20113 gnd.t216 gnd.n138 0.956468
R20114 gnd.n2 gnd.n1 0.672012
R20115 gnd.n3 gnd.n2 0.672012
R20116 gnd.n4 gnd.n3 0.672012
R20117 gnd.n5 gnd.n4 0.672012
R20118 gnd.n6 gnd.n5 0.672012
R20119 gnd.n7 gnd.n6 0.672012
R20120 gnd.n9 gnd.n8 0.672012
R20121 gnd.n10 gnd.n9 0.672012
R20122 gnd.n11 gnd.n10 0.672012
R20123 gnd.n12 gnd.n11 0.672012
R20124 gnd.n13 gnd.n12 0.672012
R20125 gnd.n14 gnd.n13 0.672012
R20126 gnd.n5659 gnd.t133 0.637812
R20127 gnd.n910 gnd.t142 0.637812
R20128 gnd.n5791 gnd.n893 0.637812
R20129 gnd.n5781 gnd.n885 0.637812
R20130 gnd.n6078 gnd.n785 0.637812
R20131 gnd.n6088 gnd.n771 0.637812
R20132 gnd.n6096 gnd.t13 0.637812
R20133 gnd.n6149 gnd.t83 0.637812
R20134 gnd.n3241 gnd.n3240 0.573776
R20135 gnd.n3240 gnd.n3238 0.573776
R20136 gnd.n3238 gnd.n3236 0.573776
R20137 gnd.n3236 gnd.n3234 0.573776
R20138 gnd.n3234 gnd.n3232 0.573776
R20139 gnd.n3206 gnd.n3205 0.573776
R20140 gnd.n3205 gnd.n3203 0.573776
R20141 gnd.n3203 gnd.n3201 0.573776
R20142 gnd.n3201 gnd.n3199 0.573776
R20143 gnd.n3199 gnd.n3197 0.573776
R20144 gnd.n3217 gnd.n3216 0.573776
R20145 gnd.n3216 gnd.n3214 0.573776
R20146 gnd.n3214 gnd.n3212 0.573776
R20147 gnd.n3212 gnd.n3210 0.573776
R20148 gnd.n3210 gnd.n3208 0.573776
R20149 gnd.n3229 gnd.n3228 0.573776
R20150 gnd.n3228 gnd.n3226 0.573776
R20151 gnd.n3226 gnd.n3224 0.573776
R20152 gnd.n3224 gnd.n3222 0.573776
R20153 gnd.n3222 gnd.n3220 0.573776
R20154 gnd.n54 gnd.n52 0.573776
R20155 gnd.n56 gnd.n54 0.573776
R20156 gnd.n58 gnd.n56 0.573776
R20157 gnd.n60 gnd.n58 0.573776
R20158 gnd.n61 gnd.n60 0.573776
R20159 gnd.n19 gnd.n17 0.573776
R20160 gnd.n21 gnd.n19 0.573776
R20161 gnd.n23 gnd.n21 0.573776
R20162 gnd.n25 gnd.n23 0.573776
R20163 gnd.n26 gnd.n25 0.573776
R20164 gnd.n30 gnd.n28 0.573776
R20165 gnd.n32 gnd.n30 0.573776
R20166 gnd.n34 gnd.n32 0.573776
R20167 gnd.n36 gnd.n34 0.573776
R20168 gnd.n37 gnd.n36 0.573776
R20169 gnd.n42 gnd.n40 0.573776
R20170 gnd.n44 gnd.n42 0.573776
R20171 gnd.n46 gnd.n44 0.573776
R20172 gnd.n48 gnd.n46 0.573776
R20173 gnd.n49 gnd.n48 0.573776
R20174 gnd gnd.n0 0.551497
R20175 gnd.n7258 gnd.n7257 0.532512
R20176 gnd.n4546 gnd.n1503 0.532512
R20177 gnd.n7073 gnd.n166 0.497451
R20178 gnd.n5454 gnd.n5453 0.497451
R20179 gnd.n497 gnd.n389 0.497451
R20180 gnd.n4708 gnd.n4707 0.497451
R20181 gnd.n6437 gnd.n422 0.489829
R20182 gnd.n5090 gnd.n1240 0.489829
R20183 gnd.n5048 gnd.n1263 0.489829
R20184 gnd.n6467 gnd.n6466 0.489829
R20185 gnd.n4278 gnd.n4277 0.486781
R20186 gnd.n3578 gnd.n3577 0.48678
R20187 gnd.n4359 gnd.n4358 0.480683
R20188 gnd.n3662 gnd.n3661 0.480683
R20189 gnd.n7332 gnd.n7331 0.470187
R20190 gnd.n2743 gnd.n2742 0.425805
R20191 gnd.n2051 gnd.n2045 0.425805
R20192 gnd.n7037 gnd.n7036 0.425805
R20193 gnd.n4418 gnd.n4417 0.425805
R20194 gnd.n7320 gnd.n79 0.4255
R20195 gnd.n4925 gnd.n1350 0.4255
R20196 gnd.n5265 gnd.n5247 0.388379
R20197 gnd.n4209 gnd.n4208 0.388379
R20198 gnd.n4177 gnd.n4176 0.388379
R20199 gnd.n4145 gnd.n4144 0.388379
R20200 gnd.n4114 gnd.n4113 0.388379
R20201 gnd.n4082 gnd.n4081 0.388379
R20202 gnd.n4050 gnd.n4049 0.388379
R20203 gnd.n4018 gnd.n4017 0.388379
R20204 gnd.n3987 gnd.n3986 0.388379
R20205 gnd.n6702 gnd.n448 0.388379
R20206 gnd.n7332 gnd.n15 0.374463
R20207 gnd.n4255 gnd.t304 0.319156
R20208 gnd.n4811 gnd.t229 0.319156
R20209 gnd.n4853 gnd.t200 0.319156
R20210 gnd.n1384 gnd.t231 0.319156
R20211 gnd.n4895 gnd.t190 0.319156
R20212 gnd.t64 gnd.n5044 0.319156
R20213 gnd.n5650 gnd.n5649 0.319156
R20214 gnd.n5739 gnd.t153 0.319156
R20215 gnd.n6107 gnd.t149 0.319156
R20216 gnd.n6351 gnd.n6350 0.319156
R20217 gnd.n6442 gnd.t53 0.319156
R20218 gnd.n6877 gnd.t174 0.319156
R20219 gnd.n6901 gnd.t197 0.319156
R20220 gnd.t172 gnd.n6997 0.319156
R20221 gnd.t205 gnd.n98 0.319156
R20222 gnd.n3496 gnd.n3474 0.311721
R20223 gnd.n5337 gnd.n5336 0.302329
R20224 gnd.n6712 gnd.n6710 0.302329
R20225 gnd gnd.n7332 0.295112
R20226 gnd.n200 gnd.n174 0.293183
R20227 gnd.n4588 gnd.n4516 0.293183
R20228 gnd.n4328 gnd.n4327 0.268793
R20229 gnd.n7134 gnd.n174 0.258122
R20230 gnd.n6578 gnd.n6577 0.258122
R20231 gnd.n5464 gnd.n5463 0.258122
R20232 gnd.n4589 gnd.n4588 0.258122
R20233 gnd.n4327 gnd.n4326 0.241354
R20234 gnd.n527 gnd.n524 0.229039
R20235 gnd.n528 gnd.n527 0.229039
R20236 gnd.n5522 gnd.n1151 0.229039
R20237 gnd.n5522 gnd.n5521 0.229039
R20238 gnd.n3650 gnd.n3449 0.206293
R20239 gnd.n4226 gnd.n4198 0.155672
R20240 gnd.n4219 gnd.n4198 0.155672
R20241 gnd.n4219 gnd.n4218 0.155672
R20242 gnd.n4218 gnd.n4202 0.155672
R20243 gnd.n4211 gnd.n4202 0.155672
R20244 gnd.n4211 gnd.n4210 0.155672
R20245 gnd.n4194 gnd.n4166 0.155672
R20246 gnd.n4187 gnd.n4166 0.155672
R20247 gnd.n4187 gnd.n4186 0.155672
R20248 gnd.n4186 gnd.n4170 0.155672
R20249 gnd.n4179 gnd.n4170 0.155672
R20250 gnd.n4179 gnd.n4178 0.155672
R20251 gnd.n4162 gnd.n4134 0.155672
R20252 gnd.n4155 gnd.n4134 0.155672
R20253 gnd.n4155 gnd.n4154 0.155672
R20254 gnd.n4154 gnd.n4138 0.155672
R20255 gnd.n4147 gnd.n4138 0.155672
R20256 gnd.n4147 gnd.n4146 0.155672
R20257 gnd.n4131 gnd.n4103 0.155672
R20258 gnd.n4124 gnd.n4103 0.155672
R20259 gnd.n4124 gnd.n4123 0.155672
R20260 gnd.n4123 gnd.n4107 0.155672
R20261 gnd.n4116 gnd.n4107 0.155672
R20262 gnd.n4116 gnd.n4115 0.155672
R20263 gnd.n4099 gnd.n4071 0.155672
R20264 gnd.n4092 gnd.n4071 0.155672
R20265 gnd.n4092 gnd.n4091 0.155672
R20266 gnd.n4091 gnd.n4075 0.155672
R20267 gnd.n4084 gnd.n4075 0.155672
R20268 gnd.n4084 gnd.n4083 0.155672
R20269 gnd.n4067 gnd.n4039 0.155672
R20270 gnd.n4060 gnd.n4039 0.155672
R20271 gnd.n4060 gnd.n4059 0.155672
R20272 gnd.n4059 gnd.n4043 0.155672
R20273 gnd.n4052 gnd.n4043 0.155672
R20274 gnd.n4052 gnd.n4051 0.155672
R20275 gnd.n4035 gnd.n4007 0.155672
R20276 gnd.n4028 gnd.n4007 0.155672
R20277 gnd.n4028 gnd.n4027 0.155672
R20278 gnd.n4027 gnd.n4011 0.155672
R20279 gnd.n4020 gnd.n4011 0.155672
R20280 gnd.n4020 gnd.n4019 0.155672
R20281 gnd.n4004 gnd.n3976 0.155672
R20282 gnd.n3997 gnd.n3976 0.155672
R20283 gnd.n3997 gnd.n3996 0.155672
R20284 gnd.n3996 gnd.n3980 0.155672
R20285 gnd.n3989 gnd.n3980 0.155672
R20286 gnd.n3989 gnd.n3988 0.155672
R20287 gnd.n4358 gnd.n3042 0.152939
R20288 gnd.n3044 gnd.n3042 0.152939
R20289 gnd.n3048 gnd.n3044 0.152939
R20290 gnd.n3049 gnd.n3048 0.152939
R20291 gnd.n3050 gnd.n3049 0.152939
R20292 gnd.n3051 gnd.n3050 0.152939
R20293 gnd.n3055 gnd.n3051 0.152939
R20294 gnd.n3056 gnd.n3055 0.152939
R20295 gnd.n3057 gnd.n3056 0.152939
R20296 gnd.n3058 gnd.n3057 0.152939
R20297 gnd.n3062 gnd.n3058 0.152939
R20298 gnd.n3063 gnd.n3062 0.152939
R20299 gnd.n3064 gnd.n3063 0.152939
R20300 gnd.n3065 gnd.n3064 0.152939
R20301 gnd.n3070 gnd.n3065 0.152939
R20302 gnd.n4328 gnd.n3070 0.152939
R20303 gnd.n3663 gnd.n3662 0.152939
R20304 gnd.n3663 gnd.n3367 0.152939
R20305 gnd.n3691 gnd.n3367 0.152939
R20306 gnd.n3692 gnd.n3691 0.152939
R20307 gnd.n3693 gnd.n3692 0.152939
R20308 gnd.n3694 gnd.n3693 0.152939
R20309 gnd.n3694 gnd.n3339 0.152939
R20310 gnd.n3721 gnd.n3339 0.152939
R20311 gnd.n3722 gnd.n3721 0.152939
R20312 gnd.n3723 gnd.n3722 0.152939
R20313 gnd.n3723 gnd.n3317 0.152939
R20314 gnd.n3752 gnd.n3317 0.152939
R20315 gnd.n3753 gnd.n3752 0.152939
R20316 gnd.n3754 gnd.n3753 0.152939
R20317 gnd.n3755 gnd.n3754 0.152939
R20318 gnd.n3757 gnd.n3755 0.152939
R20319 gnd.n3757 gnd.n3756 0.152939
R20320 gnd.n3756 gnd.n3266 0.152939
R20321 gnd.n3267 gnd.n3266 0.152939
R20322 gnd.n3268 gnd.n3267 0.152939
R20323 gnd.n3287 gnd.n3268 0.152939
R20324 gnd.n3288 gnd.n3287 0.152939
R20325 gnd.n3288 gnd.n3186 0.152939
R20326 gnd.n3847 gnd.n3186 0.152939
R20327 gnd.n3848 gnd.n3847 0.152939
R20328 gnd.n3849 gnd.n3848 0.152939
R20329 gnd.n3850 gnd.n3849 0.152939
R20330 gnd.n3850 gnd.n3159 0.152939
R20331 gnd.n3887 gnd.n3159 0.152939
R20332 gnd.n3888 gnd.n3887 0.152939
R20333 gnd.n3889 gnd.n3888 0.152939
R20334 gnd.n3890 gnd.n3889 0.152939
R20335 gnd.n3890 gnd.n3133 0.152939
R20336 gnd.n3943 gnd.n3133 0.152939
R20337 gnd.n3944 gnd.n3943 0.152939
R20338 gnd.n3946 gnd.n3944 0.152939
R20339 gnd.n3946 gnd.n3945 0.152939
R20340 gnd.n3945 gnd.n2966 0.152939
R20341 gnd.n2967 gnd.n2966 0.152939
R20342 gnd.n2968 gnd.n2967 0.152939
R20343 gnd.n2989 gnd.n2968 0.152939
R20344 gnd.n2990 gnd.n2989 0.152939
R20345 gnd.n2991 gnd.n2990 0.152939
R20346 gnd.n2992 gnd.n2991 0.152939
R20347 gnd.n2993 gnd.n2992 0.152939
R20348 gnd.n3015 gnd.n2993 0.152939
R20349 gnd.n3016 gnd.n3015 0.152939
R20350 gnd.n3017 gnd.n3016 0.152939
R20351 gnd.n3018 gnd.n3017 0.152939
R20352 gnd.n3019 gnd.n3018 0.152939
R20353 gnd.n3040 gnd.n3019 0.152939
R20354 gnd.n3041 gnd.n3040 0.152939
R20355 gnd.n4359 gnd.n3041 0.152939
R20356 gnd.n3661 gnd.n3391 0.152939
R20357 gnd.n3412 gnd.n3391 0.152939
R20358 gnd.n3413 gnd.n3412 0.152939
R20359 gnd.n3419 gnd.n3413 0.152939
R20360 gnd.n3420 gnd.n3419 0.152939
R20361 gnd.n3421 gnd.n3420 0.152939
R20362 gnd.n3421 gnd.n3410 0.152939
R20363 gnd.n3429 gnd.n3410 0.152939
R20364 gnd.n3430 gnd.n3429 0.152939
R20365 gnd.n3431 gnd.n3430 0.152939
R20366 gnd.n3431 gnd.n3408 0.152939
R20367 gnd.n3439 gnd.n3408 0.152939
R20368 gnd.n3440 gnd.n3439 0.152939
R20369 gnd.n3441 gnd.n3440 0.152939
R20370 gnd.n3441 gnd.n3406 0.152939
R20371 gnd.n3449 gnd.n3406 0.152939
R20372 gnd.n4326 gnd.n3072 0.152939
R20373 gnd.n3074 gnd.n3072 0.152939
R20374 gnd.n3078 gnd.n3074 0.152939
R20375 gnd.n3079 gnd.n3078 0.152939
R20376 gnd.n3080 gnd.n3079 0.152939
R20377 gnd.n3081 gnd.n3080 0.152939
R20378 gnd.n3085 gnd.n3081 0.152939
R20379 gnd.n3086 gnd.n3085 0.152939
R20380 gnd.n3087 gnd.n3086 0.152939
R20381 gnd.n3088 gnd.n3087 0.152939
R20382 gnd.n3092 gnd.n3088 0.152939
R20383 gnd.n3093 gnd.n3092 0.152939
R20384 gnd.n3094 gnd.n3093 0.152939
R20385 gnd.n3095 gnd.n3094 0.152939
R20386 gnd.n3099 gnd.n3095 0.152939
R20387 gnd.n3100 gnd.n3099 0.152939
R20388 gnd.n3101 gnd.n3100 0.152939
R20389 gnd.n3102 gnd.n3101 0.152939
R20390 gnd.n3106 gnd.n3102 0.152939
R20391 gnd.n3107 gnd.n3106 0.152939
R20392 gnd.n3108 gnd.n3107 0.152939
R20393 gnd.n3109 gnd.n3108 0.152939
R20394 gnd.n3116 gnd.n3109 0.152939
R20395 gnd.n3117 gnd.n3116 0.152939
R20396 gnd.n3118 gnd.n3117 0.152939
R20397 gnd.n4278 gnd.n3118 0.152939
R20398 gnd.n3824 gnd.n3823 0.152939
R20399 gnd.n3825 gnd.n3824 0.152939
R20400 gnd.n3826 gnd.n3825 0.152939
R20401 gnd.n3827 gnd.n3826 0.152939
R20402 gnd.n3828 gnd.n3827 0.152939
R20403 gnd.n3829 gnd.n3828 0.152939
R20404 gnd.n3829 gnd.n3140 0.152939
R20405 gnd.n3910 gnd.n3140 0.152939
R20406 gnd.n3911 gnd.n3910 0.152939
R20407 gnd.n3912 gnd.n3911 0.152939
R20408 gnd.n3913 gnd.n3912 0.152939
R20409 gnd.n3914 gnd.n3913 0.152939
R20410 gnd.n3915 gnd.n3914 0.152939
R20411 gnd.n3916 gnd.n3915 0.152939
R20412 gnd.n3917 gnd.n3916 0.152939
R20413 gnd.n3918 gnd.n3917 0.152939
R20414 gnd.n3919 gnd.n3918 0.152939
R20415 gnd.n3920 gnd.n3919 0.152939
R20416 gnd.n3920 gnd.n3123 0.152939
R20417 gnd.n4259 gnd.n3123 0.152939
R20418 gnd.n4260 gnd.n4259 0.152939
R20419 gnd.n4261 gnd.n4260 0.152939
R20420 gnd.n4261 gnd.n3121 0.152939
R20421 gnd.n4269 gnd.n3121 0.152939
R20422 gnd.n4270 gnd.n4269 0.152939
R20423 gnd.n4271 gnd.n4270 0.152939
R20424 gnd.n4271 gnd.n3119 0.152939
R20425 gnd.n4277 gnd.n3119 0.152939
R20426 gnd.n3579 gnd.n3578 0.152939
R20427 gnd.n3579 gnd.n3469 0.152939
R20428 gnd.n3594 gnd.n3469 0.152939
R20429 gnd.n3595 gnd.n3594 0.152939
R20430 gnd.n3596 gnd.n3595 0.152939
R20431 gnd.n3596 gnd.n3457 0.152939
R20432 gnd.n3610 gnd.n3457 0.152939
R20433 gnd.n3611 gnd.n3610 0.152939
R20434 gnd.n3612 gnd.n3611 0.152939
R20435 gnd.n3613 gnd.n3612 0.152939
R20436 gnd.n3614 gnd.n3613 0.152939
R20437 gnd.n3615 gnd.n3614 0.152939
R20438 gnd.n3616 gnd.n3615 0.152939
R20439 gnd.n3617 gnd.n3616 0.152939
R20440 gnd.n3618 gnd.n3617 0.152939
R20441 gnd.n3619 gnd.n3618 0.152939
R20442 gnd.n3620 gnd.n3619 0.152939
R20443 gnd.n3621 gnd.n3620 0.152939
R20444 gnd.n3622 gnd.n3621 0.152939
R20445 gnd.n3623 gnd.n3622 0.152939
R20446 gnd.n3624 gnd.n3623 0.152939
R20447 gnd.n3624 gnd.n3323 0.152939
R20448 gnd.n3741 gnd.n3323 0.152939
R20449 gnd.n3742 gnd.n3741 0.152939
R20450 gnd.n3743 gnd.n3742 0.152939
R20451 gnd.n3744 gnd.n3743 0.152939
R20452 gnd.n3744 gnd.n3245 0.152939
R20453 gnd.n3821 gnd.n3245 0.152939
R20454 gnd.n3497 gnd.n3496 0.152939
R20455 gnd.n3498 gnd.n3497 0.152939
R20456 gnd.n3499 gnd.n3498 0.152939
R20457 gnd.n3500 gnd.n3499 0.152939
R20458 gnd.n3501 gnd.n3500 0.152939
R20459 gnd.n3502 gnd.n3501 0.152939
R20460 gnd.n3503 gnd.n3502 0.152939
R20461 gnd.n3504 gnd.n3503 0.152939
R20462 gnd.n3505 gnd.n3504 0.152939
R20463 gnd.n3506 gnd.n3505 0.152939
R20464 gnd.n3507 gnd.n3506 0.152939
R20465 gnd.n3508 gnd.n3507 0.152939
R20466 gnd.n3509 gnd.n3508 0.152939
R20467 gnd.n3510 gnd.n3509 0.152939
R20468 gnd.n3511 gnd.n3510 0.152939
R20469 gnd.n3512 gnd.n3511 0.152939
R20470 gnd.n3513 gnd.n3512 0.152939
R20471 gnd.n3514 gnd.n3513 0.152939
R20472 gnd.n3515 gnd.n3514 0.152939
R20473 gnd.n3516 gnd.n3515 0.152939
R20474 gnd.n3517 gnd.n3516 0.152939
R20475 gnd.n3518 gnd.n3517 0.152939
R20476 gnd.n3522 gnd.n3518 0.152939
R20477 gnd.n3523 gnd.n3522 0.152939
R20478 gnd.n3523 gnd.n3480 0.152939
R20479 gnd.n3577 gnd.n3480 0.152939
R20480 gnd.n2742 gnd.n1683 0.152939
R20481 gnd.n1690 gnd.n1683 0.152939
R20482 gnd.n1691 gnd.n1690 0.152939
R20483 gnd.n1692 gnd.n1691 0.152939
R20484 gnd.n1693 gnd.n1692 0.152939
R20485 gnd.n1698 gnd.n1693 0.152939
R20486 gnd.n1699 gnd.n1698 0.152939
R20487 gnd.n1700 gnd.n1699 0.152939
R20488 gnd.n1701 gnd.n1700 0.152939
R20489 gnd.n1706 gnd.n1701 0.152939
R20490 gnd.n1707 gnd.n1706 0.152939
R20491 gnd.n1708 gnd.n1707 0.152939
R20492 gnd.n1709 gnd.n1708 0.152939
R20493 gnd.n1714 gnd.n1709 0.152939
R20494 gnd.n1715 gnd.n1714 0.152939
R20495 gnd.n1716 gnd.n1715 0.152939
R20496 gnd.n1717 gnd.n1716 0.152939
R20497 gnd.n1722 gnd.n1717 0.152939
R20498 gnd.n1723 gnd.n1722 0.152939
R20499 gnd.n1724 gnd.n1723 0.152939
R20500 gnd.n1725 gnd.n1724 0.152939
R20501 gnd.n1730 gnd.n1725 0.152939
R20502 gnd.n1731 gnd.n1730 0.152939
R20503 gnd.n1732 gnd.n1731 0.152939
R20504 gnd.n1733 gnd.n1732 0.152939
R20505 gnd.n1738 gnd.n1733 0.152939
R20506 gnd.n1739 gnd.n1738 0.152939
R20507 gnd.n1740 gnd.n1739 0.152939
R20508 gnd.n1741 gnd.n1740 0.152939
R20509 gnd.n1746 gnd.n1741 0.152939
R20510 gnd.n1747 gnd.n1746 0.152939
R20511 gnd.n1748 gnd.n1747 0.152939
R20512 gnd.n1749 gnd.n1748 0.152939
R20513 gnd.n1754 gnd.n1749 0.152939
R20514 gnd.n1755 gnd.n1754 0.152939
R20515 gnd.n1756 gnd.n1755 0.152939
R20516 gnd.n1757 gnd.n1756 0.152939
R20517 gnd.n1762 gnd.n1757 0.152939
R20518 gnd.n1763 gnd.n1762 0.152939
R20519 gnd.n1764 gnd.n1763 0.152939
R20520 gnd.n1765 gnd.n1764 0.152939
R20521 gnd.n1770 gnd.n1765 0.152939
R20522 gnd.n1771 gnd.n1770 0.152939
R20523 gnd.n1772 gnd.n1771 0.152939
R20524 gnd.n1773 gnd.n1772 0.152939
R20525 gnd.n1778 gnd.n1773 0.152939
R20526 gnd.n1779 gnd.n1778 0.152939
R20527 gnd.n1780 gnd.n1779 0.152939
R20528 gnd.n1781 gnd.n1780 0.152939
R20529 gnd.n1786 gnd.n1781 0.152939
R20530 gnd.n1787 gnd.n1786 0.152939
R20531 gnd.n1788 gnd.n1787 0.152939
R20532 gnd.n1789 gnd.n1788 0.152939
R20533 gnd.n1794 gnd.n1789 0.152939
R20534 gnd.n1795 gnd.n1794 0.152939
R20535 gnd.n1796 gnd.n1795 0.152939
R20536 gnd.n1797 gnd.n1796 0.152939
R20537 gnd.n1802 gnd.n1797 0.152939
R20538 gnd.n1803 gnd.n1802 0.152939
R20539 gnd.n1804 gnd.n1803 0.152939
R20540 gnd.n1805 gnd.n1804 0.152939
R20541 gnd.n1810 gnd.n1805 0.152939
R20542 gnd.n1811 gnd.n1810 0.152939
R20543 gnd.n1812 gnd.n1811 0.152939
R20544 gnd.n1813 gnd.n1812 0.152939
R20545 gnd.n1818 gnd.n1813 0.152939
R20546 gnd.n1819 gnd.n1818 0.152939
R20547 gnd.n1820 gnd.n1819 0.152939
R20548 gnd.n1821 gnd.n1820 0.152939
R20549 gnd.n1826 gnd.n1821 0.152939
R20550 gnd.n1827 gnd.n1826 0.152939
R20551 gnd.n1828 gnd.n1827 0.152939
R20552 gnd.n1829 gnd.n1828 0.152939
R20553 gnd.n1834 gnd.n1829 0.152939
R20554 gnd.n1835 gnd.n1834 0.152939
R20555 gnd.n1836 gnd.n1835 0.152939
R20556 gnd.n1837 gnd.n1836 0.152939
R20557 gnd.n1842 gnd.n1837 0.152939
R20558 gnd.n1843 gnd.n1842 0.152939
R20559 gnd.n1844 gnd.n1843 0.152939
R20560 gnd.n1845 gnd.n1844 0.152939
R20561 gnd.n1850 gnd.n1845 0.152939
R20562 gnd.n1851 gnd.n1850 0.152939
R20563 gnd.n1852 gnd.n1851 0.152939
R20564 gnd.n1853 gnd.n1852 0.152939
R20565 gnd.n1858 gnd.n1853 0.152939
R20566 gnd.n1859 gnd.n1858 0.152939
R20567 gnd.n1860 gnd.n1859 0.152939
R20568 gnd.n1861 gnd.n1860 0.152939
R20569 gnd.n1866 gnd.n1861 0.152939
R20570 gnd.n1867 gnd.n1866 0.152939
R20571 gnd.n1868 gnd.n1867 0.152939
R20572 gnd.n1869 gnd.n1868 0.152939
R20573 gnd.n1874 gnd.n1869 0.152939
R20574 gnd.n1875 gnd.n1874 0.152939
R20575 gnd.n1876 gnd.n1875 0.152939
R20576 gnd.n1877 gnd.n1876 0.152939
R20577 gnd.n1882 gnd.n1877 0.152939
R20578 gnd.n1883 gnd.n1882 0.152939
R20579 gnd.n1884 gnd.n1883 0.152939
R20580 gnd.n1885 gnd.n1884 0.152939
R20581 gnd.n1890 gnd.n1885 0.152939
R20582 gnd.n1891 gnd.n1890 0.152939
R20583 gnd.n1892 gnd.n1891 0.152939
R20584 gnd.n1893 gnd.n1892 0.152939
R20585 gnd.n1898 gnd.n1893 0.152939
R20586 gnd.n1899 gnd.n1898 0.152939
R20587 gnd.n1900 gnd.n1899 0.152939
R20588 gnd.n1901 gnd.n1900 0.152939
R20589 gnd.n1906 gnd.n1901 0.152939
R20590 gnd.n1907 gnd.n1906 0.152939
R20591 gnd.n1908 gnd.n1907 0.152939
R20592 gnd.n1909 gnd.n1908 0.152939
R20593 gnd.n1914 gnd.n1909 0.152939
R20594 gnd.n1915 gnd.n1914 0.152939
R20595 gnd.n1916 gnd.n1915 0.152939
R20596 gnd.n1917 gnd.n1916 0.152939
R20597 gnd.n1922 gnd.n1917 0.152939
R20598 gnd.n1923 gnd.n1922 0.152939
R20599 gnd.n1924 gnd.n1923 0.152939
R20600 gnd.n1925 gnd.n1924 0.152939
R20601 gnd.n1930 gnd.n1925 0.152939
R20602 gnd.n1931 gnd.n1930 0.152939
R20603 gnd.n1932 gnd.n1931 0.152939
R20604 gnd.n1933 gnd.n1932 0.152939
R20605 gnd.n1938 gnd.n1933 0.152939
R20606 gnd.n1939 gnd.n1938 0.152939
R20607 gnd.n1940 gnd.n1939 0.152939
R20608 gnd.n1941 gnd.n1940 0.152939
R20609 gnd.n1946 gnd.n1941 0.152939
R20610 gnd.n1947 gnd.n1946 0.152939
R20611 gnd.n1948 gnd.n1947 0.152939
R20612 gnd.n1949 gnd.n1948 0.152939
R20613 gnd.n1954 gnd.n1949 0.152939
R20614 gnd.n1955 gnd.n1954 0.152939
R20615 gnd.n1956 gnd.n1955 0.152939
R20616 gnd.n1957 gnd.n1956 0.152939
R20617 gnd.n1962 gnd.n1957 0.152939
R20618 gnd.n1963 gnd.n1962 0.152939
R20619 gnd.n1964 gnd.n1963 0.152939
R20620 gnd.n1965 gnd.n1964 0.152939
R20621 gnd.n1970 gnd.n1965 0.152939
R20622 gnd.n1971 gnd.n1970 0.152939
R20623 gnd.n1972 gnd.n1971 0.152939
R20624 gnd.n1973 gnd.n1972 0.152939
R20625 gnd.n1978 gnd.n1973 0.152939
R20626 gnd.n1979 gnd.n1978 0.152939
R20627 gnd.n1980 gnd.n1979 0.152939
R20628 gnd.n1981 gnd.n1980 0.152939
R20629 gnd.n1986 gnd.n1981 0.152939
R20630 gnd.n1987 gnd.n1986 0.152939
R20631 gnd.n1988 gnd.n1987 0.152939
R20632 gnd.n1989 gnd.n1988 0.152939
R20633 gnd.n1994 gnd.n1989 0.152939
R20634 gnd.n1995 gnd.n1994 0.152939
R20635 gnd.n1996 gnd.n1995 0.152939
R20636 gnd.n1997 gnd.n1996 0.152939
R20637 gnd.n2002 gnd.n1997 0.152939
R20638 gnd.n2003 gnd.n2002 0.152939
R20639 gnd.n2004 gnd.n2003 0.152939
R20640 gnd.n2005 gnd.n2004 0.152939
R20641 gnd.n2010 gnd.n2005 0.152939
R20642 gnd.n2011 gnd.n2010 0.152939
R20643 gnd.n2012 gnd.n2011 0.152939
R20644 gnd.n2013 gnd.n2012 0.152939
R20645 gnd.n2018 gnd.n2013 0.152939
R20646 gnd.n2019 gnd.n2018 0.152939
R20647 gnd.n2020 gnd.n2019 0.152939
R20648 gnd.n2021 gnd.n2020 0.152939
R20649 gnd.n2026 gnd.n2021 0.152939
R20650 gnd.n2027 gnd.n2026 0.152939
R20651 gnd.n2028 gnd.n2027 0.152939
R20652 gnd.n2029 gnd.n2028 0.152939
R20653 gnd.n2034 gnd.n2029 0.152939
R20654 gnd.n2035 gnd.n2034 0.152939
R20655 gnd.n2036 gnd.n2035 0.152939
R20656 gnd.n2037 gnd.n2036 0.152939
R20657 gnd.n2042 gnd.n2037 0.152939
R20658 gnd.n2043 gnd.n2042 0.152939
R20659 gnd.n2044 gnd.n2043 0.152939
R20660 gnd.n2045 gnd.n2044 0.152939
R20661 gnd.n2373 gnd.n2051 0.152939
R20662 gnd.n2373 gnd.n2372 0.152939
R20663 gnd.n2372 gnd.n2371 0.152939
R20664 gnd.n2371 gnd.n2052 0.152939
R20665 gnd.n2057 gnd.n2052 0.152939
R20666 gnd.n2058 gnd.n2057 0.152939
R20667 gnd.n2059 gnd.n2058 0.152939
R20668 gnd.n2064 gnd.n2059 0.152939
R20669 gnd.n2065 gnd.n2064 0.152939
R20670 gnd.n2066 gnd.n2065 0.152939
R20671 gnd.n2067 gnd.n2066 0.152939
R20672 gnd.n2072 gnd.n2067 0.152939
R20673 gnd.n2073 gnd.n2072 0.152939
R20674 gnd.n2074 gnd.n2073 0.152939
R20675 gnd.n2075 gnd.n2074 0.152939
R20676 gnd.n2080 gnd.n2075 0.152939
R20677 gnd.n2081 gnd.n2080 0.152939
R20678 gnd.n2082 gnd.n2081 0.152939
R20679 gnd.n2083 gnd.n2082 0.152939
R20680 gnd.n2088 gnd.n2083 0.152939
R20681 gnd.n2089 gnd.n2088 0.152939
R20682 gnd.n2090 gnd.n2089 0.152939
R20683 gnd.n2091 gnd.n2090 0.152939
R20684 gnd.n2096 gnd.n2091 0.152939
R20685 gnd.n2097 gnd.n2096 0.152939
R20686 gnd.n2098 gnd.n2097 0.152939
R20687 gnd.n2099 gnd.n2098 0.152939
R20688 gnd.n2104 gnd.n2099 0.152939
R20689 gnd.n2105 gnd.n2104 0.152939
R20690 gnd.n2106 gnd.n2105 0.152939
R20691 gnd.n2107 gnd.n2106 0.152939
R20692 gnd.n2112 gnd.n2107 0.152939
R20693 gnd.n2113 gnd.n2112 0.152939
R20694 gnd.n2114 gnd.n2113 0.152939
R20695 gnd.n2115 gnd.n2114 0.152939
R20696 gnd.n2120 gnd.n2115 0.152939
R20697 gnd.n2121 gnd.n2120 0.152939
R20698 gnd.n2122 gnd.n2121 0.152939
R20699 gnd.n2123 gnd.n2122 0.152939
R20700 gnd.n2128 gnd.n2123 0.152939
R20701 gnd.n2129 gnd.n2128 0.152939
R20702 gnd.n2130 gnd.n2129 0.152939
R20703 gnd.n2131 gnd.n2130 0.152939
R20704 gnd.n2136 gnd.n2131 0.152939
R20705 gnd.n2137 gnd.n2136 0.152939
R20706 gnd.n2138 gnd.n2137 0.152939
R20707 gnd.n2139 gnd.n2138 0.152939
R20708 gnd.n2144 gnd.n2139 0.152939
R20709 gnd.n2145 gnd.n2144 0.152939
R20710 gnd.n2146 gnd.n2145 0.152939
R20711 gnd.n2147 gnd.n2146 0.152939
R20712 gnd.n2152 gnd.n2147 0.152939
R20713 gnd.n2153 gnd.n2152 0.152939
R20714 gnd.n2154 gnd.n2153 0.152939
R20715 gnd.n2155 gnd.n2154 0.152939
R20716 gnd.n2160 gnd.n2155 0.152939
R20717 gnd.n2161 gnd.n2160 0.152939
R20718 gnd.n2162 gnd.n2161 0.152939
R20719 gnd.n2163 gnd.n2162 0.152939
R20720 gnd.n2168 gnd.n2163 0.152939
R20721 gnd.n2169 gnd.n2168 0.152939
R20722 gnd.n2170 gnd.n2169 0.152939
R20723 gnd.n2171 gnd.n2170 0.152939
R20724 gnd.n2176 gnd.n2171 0.152939
R20725 gnd.n2177 gnd.n2176 0.152939
R20726 gnd.n2178 gnd.n2177 0.152939
R20727 gnd.n2179 gnd.n2178 0.152939
R20728 gnd.n2184 gnd.n2179 0.152939
R20729 gnd.n2185 gnd.n2184 0.152939
R20730 gnd.n2186 gnd.n2185 0.152939
R20731 gnd.n2187 gnd.n2186 0.152939
R20732 gnd.n2192 gnd.n2187 0.152939
R20733 gnd.n2193 gnd.n2192 0.152939
R20734 gnd.n2194 gnd.n2193 0.152939
R20735 gnd.n2195 gnd.n2194 0.152939
R20736 gnd.n2200 gnd.n2195 0.152939
R20737 gnd.n2201 gnd.n2200 0.152939
R20738 gnd.n2202 gnd.n2201 0.152939
R20739 gnd.n2203 gnd.n2202 0.152939
R20740 gnd.n2208 gnd.n2203 0.152939
R20741 gnd.n2209 gnd.n2208 0.152939
R20742 gnd.n2210 gnd.n2209 0.152939
R20743 gnd.n2210 gnd.n246 0.152939
R20744 gnd.n7037 gnd.n246 0.152939
R20745 gnd.n7004 gnd.n7003 0.152939
R20746 gnd.n7004 gnd.n259 0.152939
R20747 gnd.n7010 gnd.n259 0.152939
R20748 gnd.n7011 gnd.n7010 0.152939
R20749 gnd.n7012 gnd.n7011 0.152939
R20750 gnd.n7012 gnd.n255 0.152939
R20751 gnd.n7018 gnd.n255 0.152939
R20752 gnd.n7019 gnd.n7018 0.152939
R20753 gnd.n7020 gnd.n7019 0.152939
R20754 gnd.n7020 gnd.n251 0.152939
R20755 gnd.n7026 gnd.n251 0.152939
R20756 gnd.n7027 gnd.n7026 0.152939
R20757 gnd.n7029 gnd.n7027 0.152939
R20758 gnd.n7029 gnd.n7028 0.152939
R20759 gnd.n7028 gnd.n247 0.152939
R20760 gnd.n7036 gnd.n247 0.152939
R20761 gnd.n7320 gnd.n77 0.152939
R20762 gnd.n103 gnd.n77 0.152939
R20763 gnd.n104 gnd.n103 0.152939
R20764 gnd.n105 gnd.n104 0.152939
R20765 gnd.n122 gnd.n105 0.152939
R20766 gnd.n123 gnd.n122 0.152939
R20767 gnd.n124 gnd.n123 0.152939
R20768 gnd.n125 gnd.n124 0.152939
R20769 gnd.n143 gnd.n125 0.152939
R20770 gnd.n144 gnd.n143 0.152939
R20771 gnd.n145 gnd.n144 0.152939
R20772 gnd.n146 gnd.n145 0.152939
R20773 gnd.n163 gnd.n146 0.152939
R20774 gnd.n164 gnd.n163 0.152939
R20775 gnd.n165 gnd.n164 0.152939
R20776 gnd.n166 gnd.n165 0.152939
R20777 gnd.n7329 gnd.n65 0.152939
R20778 gnd.n267 gnd.n65 0.152939
R20779 gnd.n268 gnd.n267 0.152939
R20780 gnd.n269 gnd.n268 0.152939
R20781 gnd.n270 gnd.n269 0.152939
R20782 gnd.n6933 gnd.n270 0.152939
R20783 gnd.n6934 gnd.n6933 0.152939
R20784 gnd.n6935 gnd.n6934 0.152939
R20785 gnd.n6936 gnd.n6935 0.152939
R20786 gnd.n6941 gnd.n6936 0.152939
R20787 gnd.n6942 gnd.n6941 0.152939
R20788 gnd.n6943 gnd.n6942 0.152939
R20789 gnd.n6944 gnd.n6943 0.152939
R20790 gnd.n6948 gnd.n6944 0.152939
R20791 gnd.n6949 gnd.n6948 0.152939
R20792 gnd.n6950 gnd.n6949 0.152939
R20793 gnd.n6952 gnd.n6950 0.152939
R20794 gnd.n6952 gnd.n6951 0.152939
R20795 gnd.n6951 gnd.n178 0.152939
R20796 gnd.n7258 gnd.n178 0.152939
R20797 gnd.n200 gnd.n199 0.152939
R20798 gnd.n207 gnd.n199 0.152939
R20799 gnd.n208 gnd.n207 0.152939
R20800 gnd.n209 gnd.n208 0.152939
R20801 gnd.n209 gnd.n197 0.152939
R20802 gnd.n217 gnd.n197 0.152939
R20803 gnd.n218 gnd.n217 0.152939
R20804 gnd.n219 gnd.n218 0.152939
R20805 gnd.n219 gnd.n195 0.152939
R20806 gnd.n227 gnd.n195 0.152939
R20807 gnd.n228 gnd.n227 0.152939
R20808 gnd.n229 gnd.n228 0.152939
R20809 gnd.n229 gnd.n193 0.152939
R20810 gnd.n236 gnd.n193 0.152939
R20811 gnd.n237 gnd.n236 0.152939
R20812 gnd.n238 gnd.n237 0.152939
R20813 gnd.n238 gnd.n179 0.152939
R20814 gnd.n7257 gnd.n179 0.152939
R20815 gnd.n7074 gnd.n7073 0.152939
R20816 gnd.n7075 gnd.n7074 0.152939
R20817 gnd.n7076 gnd.n7075 0.152939
R20818 gnd.n7077 gnd.n7076 0.152939
R20819 gnd.n7078 gnd.n7077 0.152939
R20820 gnd.n7079 gnd.n7078 0.152939
R20821 gnd.n7080 gnd.n7079 0.152939
R20822 gnd.n7081 gnd.n7080 0.152939
R20823 gnd.n7082 gnd.n7081 0.152939
R20824 gnd.n7083 gnd.n7082 0.152939
R20825 gnd.n7084 gnd.n7083 0.152939
R20826 gnd.n7085 gnd.n7084 0.152939
R20827 gnd.n7086 gnd.n7085 0.152939
R20828 gnd.n7087 gnd.n7086 0.152939
R20829 gnd.n7088 gnd.n7087 0.152939
R20830 gnd.n7089 gnd.n7088 0.152939
R20831 gnd.n7090 gnd.n7089 0.152939
R20832 gnd.n7091 gnd.n7090 0.152939
R20833 gnd.n7092 gnd.n7091 0.152939
R20834 gnd.n7093 gnd.n7092 0.152939
R20835 gnd.n7094 gnd.n7093 0.152939
R20836 gnd.n7095 gnd.n7094 0.152939
R20837 gnd.n7096 gnd.n7095 0.152939
R20838 gnd.n7097 gnd.n7096 0.152939
R20839 gnd.n7098 gnd.n7097 0.152939
R20840 gnd.n7099 gnd.n7098 0.152939
R20841 gnd.n7100 gnd.n7099 0.152939
R20842 gnd.n7101 gnd.n7100 0.152939
R20843 gnd.n7102 gnd.n7101 0.152939
R20844 gnd.n7103 gnd.n7102 0.152939
R20845 gnd.n7104 gnd.n7103 0.152939
R20846 gnd.n7105 gnd.n7104 0.152939
R20847 gnd.n7106 gnd.n7105 0.152939
R20848 gnd.n7107 gnd.n7106 0.152939
R20849 gnd.n7108 gnd.n7107 0.152939
R20850 gnd.n7109 gnd.n7108 0.152939
R20851 gnd.n7177 gnd.n7109 0.152939
R20852 gnd.n7177 gnd.n7176 0.152939
R20853 gnd.n7176 gnd.n7175 0.152939
R20854 gnd.n7175 gnd.n7113 0.152939
R20855 gnd.n7114 gnd.n7113 0.152939
R20856 gnd.n7115 gnd.n7114 0.152939
R20857 gnd.n7116 gnd.n7115 0.152939
R20858 gnd.n7117 gnd.n7116 0.152939
R20859 gnd.n7118 gnd.n7117 0.152939
R20860 gnd.n7119 gnd.n7118 0.152939
R20861 gnd.n7120 gnd.n7119 0.152939
R20862 gnd.n7121 gnd.n7120 0.152939
R20863 gnd.n7122 gnd.n7121 0.152939
R20864 gnd.n7123 gnd.n7122 0.152939
R20865 gnd.n7124 gnd.n7123 0.152939
R20866 gnd.n7125 gnd.n7124 0.152939
R20867 gnd.n7126 gnd.n7125 0.152939
R20868 gnd.n7127 gnd.n7126 0.152939
R20869 gnd.n7128 gnd.n7127 0.152939
R20870 gnd.n7129 gnd.n7128 0.152939
R20871 gnd.n7135 gnd.n7129 0.152939
R20872 gnd.n7135 gnd.n7134 0.152939
R20873 gnd.n498 gnd.n497 0.152939
R20874 gnd.n499 gnd.n498 0.152939
R20875 gnd.n500 gnd.n499 0.152939
R20876 gnd.n501 gnd.n500 0.152939
R20877 gnd.n502 gnd.n501 0.152939
R20878 gnd.n503 gnd.n502 0.152939
R20879 gnd.n504 gnd.n503 0.152939
R20880 gnd.n505 gnd.n504 0.152939
R20881 gnd.n506 gnd.n505 0.152939
R20882 gnd.n507 gnd.n506 0.152939
R20883 gnd.n508 gnd.n507 0.152939
R20884 gnd.n509 gnd.n508 0.152939
R20885 gnd.n510 gnd.n509 0.152939
R20886 gnd.n511 gnd.n510 0.152939
R20887 gnd.n512 gnd.n511 0.152939
R20888 gnd.n513 gnd.n512 0.152939
R20889 gnd.n514 gnd.n513 0.152939
R20890 gnd.n517 gnd.n514 0.152939
R20891 gnd.n518 gnd.n517 0.152939
R20892 gnd.n519 gnd.n518 0.152939
R20893 gnd.n520 gnd.n519 0.152939
R20894 gnd.n521 gnd.n520 0.152939
R20895 gnd.n522 gnd.n521 0.152939
R20896 gnd.n523 gnd.n522 0.152939
R20897 gnd.n524 gnd.n523 0.152939
R20898 gnd.n529 gnd.n528 0.152939
R20899 gnd.n530 gnd.n529 0.152939
R20900 gnd.n531 gnd.n530 0.152939
R20901 gnd.n532 gnd.n531 0.152939
R20902 gnd.n533 gnd.n532 0.152939
R20903 gnd.n534 gnd.n533 0.152939
R20904 gnd.n535 gnd.n534 0.152939
R20905 gnd.n536 gnd.n535 0.152939
R20906 gnd.n537 gnd.n536 0.152939
R20907 gnd.n540 gnd.n537 0.152939
R20908 gnd.n541 gnd.n540 0.152939
R20909 gnd.n542 gnd.n541 0.152939
R20910 gnd.n543 gnd.n542 0.152939
R20911 gnd.n544 gnd.n543 0.152939
R20912 gnd.n545 gnd.n544 0.152939
R20913 gnd.n546 gnd.n545 0.152939
R20914 gnd.n547 gnd.n546 0.152939
R20915 gnd.n548 gnd.n547 0.152939
R20916 gnd.n549 gnd.n548 0.152939
R20917 gnd.n550 gnd.n549 0.152939
R20918 gnd.n551 gnd.n550 0.152939
R20919 gnd.n552 gnd.n551 0.152939
R20920 gnd.n553 gnd.n552 0.152939
R20921 gnd.n554 gnd.n553 0.152939
R20922 gnd.n555 gnd.n554 0.152939
R20923 gnd.n556 gnd.n555 0.152939
R20924 gnd.n557 gnd.n556 0.152939
R20925 gnd.n558 gnd.n557 0.152939
R20926 gnd.n6579 gnd.n558 0.152939
R20927 gnd.n6579 gnd.n6578 0.152939
R20928 gnd.n6737 gnd.n389 0.152939
R20929 gnd.n6738 gnd.n6737 0.152939
R20930 gnd.n6739 gnd.n6738 0.152939
R20931 gnd.n6740 gnd.n6739 0.152939
R20932 gnd.n6740 gnd.n356 0.152939
R20933 gnd.n6806 gnd.n356 0.152939
R20934 gnd.n6807 gnd.n6806 0.152939
R20935 gnd.n6808 gnd.n6807 0.152939
R20936 gnd.n6809 gnd.n6808 0.152939
R20937 gnd.n6809 gnd.n327 0.152939
R20938 gnd.n6841 gnd.n327 0.152939
R20939 gnd.n6842 gnd.n6841 0.152939
R20940 gnd.n6843 gnd.n6842 0.152939
R20941 gnd.n6844 gnd.n6843 0.152939
R20942 gnd.n6844 gnd.n78 0.152939
R20943 gnd.n7320 gnd.n78 0.152939
R20944 gnd.n1396 gnd.n1331 0.152939
R20945 gnd.n4944 gnd.n1331 0.152939
R20946 gnd.n4945 gnd.n4944 0.152939
R20947 gnd.n4946 gnd.n4945 0.152939
R20948 gnd.n4947 gnd.n4946 0.152939
R20949 gnd.n4948 gnd.n4947 0.152939
R20950 gnd.n4950 gnd.n4948 0.152939
R20951 gnd.n4951 gnd.n4950 0.152939
R20952 gnd.n4951 gnd.n1281 0.152939
R20953 gnd.n5020 gnd.n1281 0.152939
R20954 gnd.n5021 gnd.n5020 0.152939
R20955 gnd.n5022 gnd.n5021 0.152939
R20956 gnd.n5022 gnd.n1277 0.152939
R20957 gnd.n5030 gnd.n1277 0.152939
R20958 gnd.n5031 gnd.n5030 0.152939
R20959 gnd.n5032 gnd.n5031 0.152939
R20960 gnd.n5033 gnd.n5032 0.152939
R20961 gnd.n5034 gnd.n5033 0.152939
R20962 gnd.n5037 gnd.n5034 0.152939
R20963 gnd.n5038 gnd.n5037 0.152939
R20964 gnd.n5039 gnd.n5038 0.152939
R20965 gnd.n5040 gnd.n5039 0.152939
R20966 gnd.n5099 gnd.n5040 0.152939
R20967 gnd.n5102 gnd.n5099 0.152939
R20968 gnd.n5103 gnd.n5102 0.152939
R20969 gnd.n5104 gnd.n5103 0.152939
R20970 gnd.n5104 gnd.n5078 0.152939
R20971 gnd.n5123 gnd.n5078 0.152939
R20972 gnd.n5124 gnd.n5123 0.152939
R20973 gnd.n5125 gnd.n5124 0.152939
R20974 gnd.n5125 gnd.n5065 0.152939
R20975 gnd.n5144 gnd.n5065 0.152939
R20976 gnd.n5145 gnd.n5144 0.152939
R20977 gnd.n5146 gnd.n5145 0.152939
R20978 gnd.n5147 gnd.n5146 0.152939
R20979 gnd.n5147 gnd.n1067 0.152939
R20980 gnd.n5631 gnd.n1067 0.152939
R20981 gnd.n5632 gnd.n5631 0.152939
R20982 gnd.n5633 gnd.n5632 0.152939
R20983 gnd.n5634 gnd.n5633 0.152939
R20984 gnd.n5635 gnd.n5634 0.152939
R20985 gnd.n5637 gnd.n5635 0.152939
R20986 gnd.n5638 gnd.n5637 0.152939
R20987 gnd.n5638 gnd.n985 0.152939
R20988 gnd.n5697 gnd.n985 0.152939
R20989 gnd.n5698 gnd.n5697 0.152939
R20990 gnd.n5699 gnd.n5698 0.152939
R20991 gnd.n5700 gnd.n5699 0.152939
R20992 gnd.n5700 gnd.n923 0.152939
R20993 gnd.n5768 gnd.n923 0.152939
R20994 gnd.n5769 gnd.n5768 0.152939
R20995 gnd.n5770 gnd.n5769 0.152939
R20996 gnd.n5770 gnd.n919 0.152939
R20997 gnd.n5776 gnd.n919 0.152939
R20998 gnd.n5777 gnd.n5776 0.152939
R20999 gnd.n5778 gnd.n5777 0.152939
R21000 gnd.n5778 gnd.n868 0.152939
R21001 gnd.n5869 gnd.n868 0.152939
R21002 gnd.n5870 gnd.n5869 0.152939
R21003 gnd.n5871 gnd.n5870 0.152939
R21004 gnd.n5872 gnd.n5871 0.152939
R21005 gnd.n5873 gnd.n5872 0.152939
R21006 gnd.n5874 gnd.n5873 0.152939
R21007 gnd.n5874 gnd.n829 0.152939
R21008 gnd.n5926 gnd.n829 0.152939
R21009 gnd.n5927 gnd.n5926 0.152939
R21010 gnd.n5928 gnd.n5927 0.152939
R21011 gnd.n5929 gnd.n5928 0.152939
R21012 gnd.n5930 gnd.n5929 0.152939
R21013 gnd.n5930 gnd.n782 0.152939
R21014 gnd.n6081 gnd.n782 0.152939
R21015 gnd.n6082 gnd.n6081 0.152939
R21016 gnd.n6083 gnd.n6082 0.152939
R21017 gnd.n6084 gnd.n6083 0.152939
R21018 gnd.n6084 gnd.n753 0.152939
R21019 gnd.n6117 gnd.n753 0.152939
R21020 gnd.n6118 gnd.n6117 0.152939
R21021 gnd.n6119 gnd.n6118 0.152939
R21022 gnd.n6119 gnd.n730 0.152939
R21023 gnd.n6144 gnd.n730 0.152939
R21024 gnd.n6145 gnd.n6144 0.152939
R21025 gnd.n6146 gnd.n6145 0.152939
R21026 gnd.n6146 gnd.n704 0.152939
R21027 gnd.n6183 gnd.n704 0.152939
R21028 gnd.n6184 gnd.n6183 0.152939
R21029 gnd.n6185 gnd.n6184 0.152939
R21030 gnd.n6185 gnd.n651 0.152939
R21031 gnd.n6355 gnd.n651 0.152939
R21032 gnd.n6356 gnd.n6355 0.152939
R21033 gnd.n6357 gnd.n6356 0.152939
R21034 gnd.n6358 gnd.n6357 0.152939
R21035 gnd.n6358 gnd.n626 0.152939
R21036 gnd.n6385 gnd.n626 0.152939
R21037 gnd.n6386 gnd.n6385 0.152939
R21038 gnd.n6387 gnd.n6386 0.152939
R21039 gnd.n6388 gnd.n6387 0.152939
R21040 gnd.n6388 gnd.n601 0.152939
R21041 gnd.n6415 gnd.n601 0.152939
R21042 gnd.n6416 gnd.n6415 0.152939
R21043 gnd.n6417 gnd.n6416 0.152939
R21044 gnd.n6418 gnd.n6417 0.152939
R21045 gnd.n6418 gnd.n576 0.152939
R21046 gnd.n6445 gnd.n576 0.152939
R21047 gnd.n6446 gnd.n6445 0.152939
R21048 gnd.n6447 gnd.n6446 0.152939
R21049 gnd.n6448 gnd.n6447 0.152939
R21050 gnd.n6449 gnd.n6448 0.152939
R21051 gnd.n6451 gnd.n6449 0.152939
R21052 gnd.n6452 gnd.n6451 0.152939
R21053 gnd.n6452 gnd.n415 0.152939
R21054 gnd.n6719 gnd.n415 0.152939
R21055 gnd.n6720 gnd.n6719 0.152939
R21056 gnd.n6721 gnd.n6720 0.152939
R21057 gnd.n6722 gnd.n6721 0.152939
R21058 gnd.n6722 gnd.n371 0.152939
R21059 gnd.n6757 gnd.n371 0.152939
R21060 gnd.n6758 gnd.n6757 0.152939
R21061 gnd.n6759 gnd.n6758 0.152939
R21062 gnd.n6760 gnd.n6759 0.152939
R21063 gnd.n6761 gnd.n6760 0.152939
R21064 gnd.n6764 gnd.n6761 0.152939
R21065 gnd.n6765 gnd.n6764 0.152939
R21066 gnd.n6766 gnd.n6765 0.152939
R21067 gnd.n6767 gnd.n6766 0.152939
R21068 gnd.n6770 gnd.n6767 0.152939
R21069 gnd.n6771 gnd.n6770 0.152939
R21070 gnd.n6772 gnd.n6771 0.152939
R21071 gnd.n4717 gnd.n1503 0.152939
R21072 gnd.n4718 gnd.n4717 0.152939
R21073 gnd.n4719 gnd.n4718 0.152939
R21074 gnd.n4720 gnd.n4719 0.152939
R21075 gnd.n4721 gnd.n4720 0.152939
R21076 gnd.n4721 gnd.n1476 0.152939
R21077 gnd.n4753 gnd.n1476 0.152939
R21078 gnd.n4754 gnd.n4753 0.152939
R21079 gnd.n4756 gnd.n4754 0.152939
R21080 gnd.n4756 gnd.n4755 0.152939
R21081 gnd.n4755 gnd.n1453 0.152939
R21082 gnd.n1454 gnd.n1453 0.152939
R21083 gnd.n1455 gnd.n1454 0.152939
R21084 gnd.n1455 gnd.n1419 0.152939
R21085 gnd.n4830 gnd.n1419 0.152939
R21086 gnd.n4831 gnd.n4830 0.152939
R21087 gnd.n4832 gnd.n4831 0.152939
R21088 gnd.n4833 gnd.n4832 0.152939
R21089 gnd.n4834 gnd.n4833 0.152939
R21090 gnd.n4835 gnd.n4834 0.152939
R21091 gnd.n4526 gnd.n4516 0.152939
R21092 gnd.n4527 gnd.n4526 0.152939
R21093 gnd.n4528 gnd.n4527 0.152939
R21094 gnd.n4529 gnd.n4528 0.152939
R21095 gnd.n4530 gnd.n4529 0.152939
R21096 gnd.n4531 gnd.n4530 0.152939
R21097 gnd.n4532 gnd.n4531 0.152939
R21098 gnd.n4533 gnd.n4532 0.152939
R21099 gnd.n4534 gnd.n4533 0.152939
R21100 gnd.n4535 gnd.n4534 0.152939
R21101 gnd.n4536 gnd.n4535 0.152939
R21102 gnd.n4537 gnd.n4536 0.152939
R21103 gnd.n4538 gnd.n4537 0.152939
R21104 gnd.n4539 gnd.n4538 0.152939
R21105 gnd.n4540 gnd.n4539 0.152939
R21106 gnd.n4548 gnd.n4540 0.152939
R21107 gnd.n4548 gnd.n4547 0.152939
R21108 gnd.n4547 gnd.n4546 0.152939
R21109 gnd.n4926 gnd.n4925 0.152939
R21110 gnd.n4927 gnd.n4926 0.152939
R21111 gnd.n4927 gnd.n1316 0.152939
R21112 gnd.n4977 gnd.n1316 0.152939
R21113 gnd.n4978 gnd.n4977 0.152939
R21114 gnd.n4979 gnd.n4978 0.152939
R21115 gnd.n4980 gnd.n4979 0.152939
R21116 gnd.n4980 gnd.n1288 0.152939
R21117 gnd.n5011 gnd.n1288 0.152939
R21118 gnd.n5012 gnd.n5011 0.152939
R21119 gnd.n5013 gnd.n5012 0.152939
R21120 gnd.n5013 gnd.n1219 0.152939
R21121 gnd.n5359 gnd.n1219 0.152939
R21122 gnd.n5360 gnd.n5359 0.152939
R21123 gnd.n5361 gnd.n5360 0.152939
R21124 gnd.n5454 gnd.n5361 0.152939
R21125 gnd.n5453 gnd.n5362 0.152939
R21126 gnd.n5365 gnd.n5362 0.152939
R21127 gnd.n5366 gnd.n5365 0.152939
R21128 gnd.n5367 gnd.n5366 0.152939
R21129 gnd.n5371 gnd.n5367 0.152939
R21130 gnd.n5372 gnd.n5371 0.152939
R21131 gnd.n5373 gnd.n5372 0.152939
R21132 gnd.n5374 gnd.n5373 0.152939
R21133 gnd.n5378 gnd.n5374 0.152939
R21134 gnd.n5379 gnd.n5378 0.152939
R21135 gnd.n5380 gnd.n5379 0.152939
R21136 gnd.n5381 gnd.n5380 0.152939
R21137 gnd.n5385 gnd.n5381 0.152939
R21138 gnd.n5386 gnd.n5385 0.152939
R21139 gnd.n5387 gnd.n5386 0.152939
R21140 gnd.n5388 gnd.n5387 0.152939
R21141 gnd.n5395 gnd.n5388 0.152939
R21142 gnd.n5396 gnd.n5395 0.152939
R21143 gnd.n5397 gnd.n5396 0.152939
R21144 gnd.n5398 gnd.n5397 0.152939
R21145 gnd.n5402 gnd.n5398 0.152939
R21146 gnd.n5403 gnd.n5402 0.152939
R21147 gnd.n5404 gnd.n5403 0.152939
R21148 gnd.n5405 gnd.n5404 0.152939
R21149 gnd.n5405 gnd.n1151 0.152939
R21150 gnd.n5521 gnd.n5520 0.152939
R21151 gnd.n5520 gnd.n1152 0.152939
R21152 gnd.n1159 gnd.n1152 0.152939
R21153 gnd.n1160 gnd.n1159 0.152939
R21154 gnd.n1161 gnd.n1160 0.152939
R21155 gnd.n1162 gnd.n1161 0.152939
R21156 gnd.n1166 gnd.n1162 0.152939
R21157 gnd.n1167 gnd.n1166 0.152939
R21158 gnd.n5503 gnd.n1167 0.152939
R21159 gnd.n5503 gnd.n5502 0.152939
R21160 gnd.n5502 gnd.n5501 0.152939
R21161 gnd.n5501 gnd.n1171 0.152939
R21162 gnd.n1177 gnd.n1171 0.152939
R21163 gnd.n1178 gnd.n1177 0.152939
R21164 gnd.n1179 gnd.n1178 0.152939
R21165 gnd.n1180 gnd.n1179 0.152939
R21166 gnd.n1184 gnd.n1180 0.152939
R21167 gnd.n1185 gnd.n1184 0.152939
R21168 gnd.n1186 gnd.n1185 0.152939
R21169 gnd.n1187 gnd.n1186 0.152939
R21170 gnd.n1191 gnd.n1187 0.152939
R21171 gnd.n1192 gnd.n1191 0.152939
R21172 gnd.n1193 gnd.n1192 0.152939
R21173 gnd.n1194 gnd.n1193 0.152939
R21174 gnd.n1198 gnd.n1194 0.152939
R21175 gnd.n1199 gnd.n1198 0.152939
R21176 gnd.n1200 gnd.n1199 0.152939
R21177 gnd.n1201 gnd.n1200 0.152939
R21178 gnd.n1207 gnd.n1201 0.152939
R21179 gnd.n5464 gnd.n1207 0.152939
R21180 gnd.n4707 gnd.n1513 0.152939
R21181 gnd.n4454 gnd.n1513 0.152939
R21182 gnd.n4455 gnd.n4454 0.152939
R21183 gnd.n4456 gnd.n4455 0.152939
R21184 gnd.n4457 gnd.n4456 0.152939
R21185 gnd.n4458 gnd.n4457 0.152939
R21186 gnd.n4459 gnd.n4458 0.152939
R21187 gnd.n4460 gnd.n4459 0.152939
R21188 gnd.n4461 gnd.n4460 0.152939
R21189 gnd.n4462 gnd.n4461 0.152939
R21190 gnd.n4463 gnd.n4462 0.152939
R21191 gnd.n4464 gnd.n4463 0.152939
R21192 gnd.n4465 gnd.n4464 0.152939
R21193 gnd.n4466 gnd.n4465 0.152939
R21194 gnd.n4467 gnd.n4466 0.152939
R21195 gnd.n4468 gnd.n4467 0.152939
R21196 gnd.n4469 gnd.n4468 0.152939
R21197 gnd.n4472 gnd.n4469 0.152939
R21198 gnd.n4473 gnd.n4472 0.152939
R21199 gnd.n4474 gnd.n4473 0.152939
R21200 gnd.n4475 gnd.n4474 0.152939
R21201 gnd.n4476 gnd.n4475 0.152939
R21202 gnd.n4477 gnd.n4476 0.152939
R21203 gnd.n4478 gnd.n4477 0.152939
R21204 gnd.n4479 gnd.n4478 0.152939
R21205 gnd.n4480 gnd.n4479 0.152939
R21206 gnd.n4481 gnd.n4480 0.152939
R21207 gnd.n4482 gnd.n4481 0.152939
R21208 gnd.n4483 gnd.n4482 0.152939
R21209 gnd.n4484 gnd.n4483 0.152939
R21210 gnd.n4485 gnd.n4484 0.152939
R21211 gnd.n4486 gnd.n4485 0.152939
R21212 gnd.n4487 gnd.n4486 0.152939
R21213 gnd.n4488 gnd.n4487 0.152939
R21214 gnd.n4489 gnd.n4488 0.152939
R21215 gnd.n4490 gnd.n4489 0.152939
R21216 gnd.n4491 gnd.n4490 0.152939
R21217 gnd.n4494 gnd.n4491 0.152939
R21218 gnd.n4495 gnd.n4494 0.152939
R21219 gnd.n4496 gnd.n4495 0.152939
R21220 gnd.n4497 gnd.n4496 0.152939
R21221 gnd.n4498 gnd.n4497 0.152939
R21222 gnd.n4499 gnd.n4498 0.152939
R21223 gnd.n4500 gnd.n4499 0.152939
R21224 gnd.n4501 gnd.n4500 0.152939
R21225 gnd.n4502 gnd.n4501 0.152939
R21226 gnd.n4503 gnd.n4502 0.152939
R21227 gnd.n4504 gnd.n4503 0.152939
R21228 gnd.n4505 gnd.n4504 0.152939
R21229 gnd.n4506 gnd.n4505 0.152939
R21230 gnd.n4507 gnd.n4506 0.152939
R21231 gnd.n4508 gnd.n4507 0.152939
R21232 gnd.n4509 gnd.n4508 0.152939
R21233 gnd.n4510 gnd.n4509 0.152939
R21234 gnd.n4511 gnd.n4510 0.152939
R21235 gnd.n4512 gnd.n4511 0.152939
R21236 gnd.n4590 gnd.n4512 0.152939
R21237 gnd.n4590 gnd.n4589 0.152939
R21238 gnd.n4709 gnd.n4708 0.152939
R21239 gnd.n4710 gnd.n4709 0.152939
R21240 gnd.n4710 gnd.n1486 0.152939
R21241 gnd.n4742 gnd.n1486 0.152939
R21242 gnd.n4743 gnd.n4742 0.152939
R21243 gnd.n4744 gnd.n4743 0.152939
R21244 gnd.n4744 gnd.n1464 0.152939
R21245 gnd.n4769 gnd.n1464 0.152939
R21246 gnd.n4770 gnd.n4769 0.152939
R21247 gnd.n4771 gnd.n4770 0.152939
R21248 gnd.n4771 gnd.n1428 0.152939
R21249 gnd.n4821 gnd.n1428 0.152939
R21250 gnd.n4822 gnd.n4821 0.152939
R21251 gnd.n4823 gnd.n4822 0.152939
R21252 gnd.n4823 gnd.n1349 0.152939
R21253 gnd.n4925 gnd.n1349 0.152939
R21254 gnd.n4419 gnd.n4418 0.152939
R21255 gnd.n4420 gnd.n4419 0.152939
R21256 gnd.n4423 gnd.n4420 0.152939
R21257 gnd.n4424 gnd.n4423 0.152939
R21258 gnd.n4425 gnd.n4424 0.152939
R21259 gnd.n4426 gnd.n4425 0.152939
R21260 gnd.n4429 gnd.n4426 0.152939
R21261 gnd.n4430 gnd.n4429 0.152939
R21262 gnd.n4431 gnd.n4430 0.152939
R21263 gnd.n4432 gnd.n4431 0.152939
R21264 gnd.n4433 gnd.n4432 0.152939
R21265 gnd.n4433 gnd.n1446 0.152939
R21266 gnd.n4804 gnd.n1446 0.152939
R21267 gnd.n4805 gnd.n4804 0.152939
R21268 gnd.n4806 gnd.n4805 0.152939
R21269 gnd.n4807 gnd.n4806 0.152939
R21270 gnd.n2744 gnd.n2743 0.152939
R21271 gnd.n2744 gnd.n1677 0.152939
R21272 gnd.n2752 gnd.n1677 0.152939
R21273 gnd.n2753 gnd.n2752 0.152939
R21274 gnd.n2754 gnd.n2753 0.152939
R21275 gnd.n2754 gnd.n1671 0.152939
R21276 gnd.n2762 gnd.n1671 0.152939
R21277 gnd.n2763 gnd.n2762 0.152939
R21278 gnd.n2764 gnd.n2763 0.152939
R21279 gnd.n2764 gnd.n1665 0.152939
R21280 gnd.n2772 gnd.n1665 0.152939
R21281 gnd.n2773 gnd.n2772 0.152939
R21282 gnd.n2774 gnd.n2773 0.152939
R21283 gnd.n2774 gnd.n1659 0.152939
R21284 gnd.n2782 gnd.n1659 0.152939
R21285 gnd.n2783 gnd.n2782 0.152939
R21286 gnd.n2784 gnd.n2783 0.152939
R21287 gnd.n2784 gnd.n1653 0.152939
R21288 gnd.n2792 gnd.n1653 0.152939
R21289 gnd.n2793 gnd.n2792 0.152939
R21290 gnd.n2794 gnd.n2793 0.152939
R21291 gnd.n2794 gnd.n1647 0.152939
R21292 gnd.n2802 gnd.n1647 0.152939
R21293 gnd.n2803 gnd.n2802 0.152939
R21294 gnd.n2804 gnd.n2803 0.152939
R21295 gnd.n2804 gnd.n1641 0.152939
R21296 gnd.n2812 gnd.n1641 0.152939
R21297 gnd.n2813 gnd.n2812 0.152939
R21298 gnd.n2814 gnd.n2813 0.152939
R21299 gnd.n2814 gnd.n1635 0.152939
R21300 gnd.n2822 gnd.n1635 0.152939
R21301 gnd.n2823 gnd.n2822 0.152939
R21302 gnd.n2824 gnd.n2823 0.152939
R21303 gnd.n2824 gnd.n1629 0.152939
R21304 gnd.n2832 gnd.n1629 0.152939
R21305 gnd.n2833 gnd.n2832 0.152939
R21306 gnd.n2834 gnd.n2833 0.152939
R21307 gnd.n2834 gnd.n1623 0.152939
R21308 gnd.n2842 gnd.n1623 0.152939
R21309 gnd.n2843 gnd.n2842 0.152939
R21310 gnd.n2844 gnd.n2843 0.152939
R21311 gnd.n2844 gnd.n1617 0.152939
R21312 gnd.n2852 gnd.n1617 0.152939
R21313 gnd.n2853 gnd.n2852 0.152939
R21314 gnd.n2854 gnd.n2853 0.152939
R21315 gnd.n2854 gnd.n1611 0.152939
R21316 gnd.n2862 gnd.n1611 0.152939
R21317 gnd.n2863 gnd.n2862 0.152939
R21318 gnd.n2864 gnd.n2863 0.152939
R21319 gnd.n2864 gnd.n1605 0.152939
R21320 gnd.n2872 gnd.n1605 0.152939
R21321 gnd.n2873 gnd.n2872 0.152939
R21322 gnd.n2874 gnd.n2873 0.152939
R21323 gnd.n2874 gnd.n1599 0.152939
R21324 gnd.n2882 gnd.n1599 0.152939
R21325 gnd.n2883 gnd.n2882 0.152939
R21326 gnd.n2884 gnd.n2883 0.152939
R21327 gnd.n2884 gnd.n1593 0.152939
R21328 gnd.n2892 gnd.n1593 0.152939
R21329 gnd.n2893 gnd.n2892 0.152939
R21330 gnd.n2894 gnd.n2893 0.152939
R21331 gnd.n2894 gnd.n1587 0.152939
R21332 gnd.n2902 gnd.n1587 0.152939
R21333 gnd.n2903 gnd.n2902 0.152939
R21334 gnd.n2904 gnd.n2903 0.152939
R21335 gnd.n2904 gnd.n1581 0.152939
R21336 gnd.n2912 gnd.n1581 0.152939
R21337 gnd.n2913 gnd.n2912 0.152939
R21338 gnd.n2914 gnd.n2913 0.152939
R21339 gnd.n2914 gnd.n1575 0.152939
R21340 gnd.n2922 gnd.n1575 0.152939
R21341 gnd.n2923 gnd.n2922 0.152939
R21342 gnd.n2924 gnd.n2923 0.152939
R21343 gnd.n2924 gnd.n1569 0.152939
R21344 gnd.n2932 gnd.n1569 0.152939
R21345 gnd.n2933 gnd.n2932 0.152939
R21346 gnd.n2934 gnd.n2933 0.152939
R21347 gnd.n2934 gnd.n1563 0.152939
R21348 gnd.n2942 gnd.n1563 0.152939
R21349 gnd.n2943 gnd.n2942 0.152939
R21350 gnd.n2945 gnd.n2943 0.152939
R21351 gnd.n2945 gnd.n2944 0.152939
R21352 gnd.n2944 gnd.n1557 0.152939
R21353 gnd.n4417 gnd.n1557 0.152939
R21354 gnd.n5091 gnd.n5090 0.152939
R21355 gnd.n5092 gnd.n5091 0.152939
R21356 gnd.n5092 gnd.n5084 0.152939
R21357 gnd.n5112 gnd.n5084 0.152939
R21358 gnd.n5113 gnd.n5112 0.152939
R21359 gnd.n5114 gnd.n5113 0.152939
R21360 gnd.n5114 gnd.n5072 0.152939
R21361 gnd.n5133 gnd.n5072 0.152939
R21362 gnd.n5134 gnd.n5133 0.152939
R21363 gnd.n5136 gnd.n5134 0.152939
R21364 gnd.n5136 gnd.n5135 0.152939
R21365 gnd.n5135 gnd.n1083 0.152939
R21366 gnd.n5615 gnd.n1083 0.152939
R21367 gnd.n5615 gnd.n5614 0.152939
R21368 gnd.n5614 gnd.n5613 0.152939
R21369 gnd.n5613 gnd.n1084 0.152939
R21370 gnd.n5609 gnd.n1084 0.152939
R21371 gnd.n5609 gnd.n5608 0.152939
R21372 gnd.n5608 gnd.n5607 0.152939
R21373 gnd.n5607 gnd.n5601 0.152939
R21374 gnd.n5603 gnd.n5601 0.152939
R21375 gnd.n5603 gnd.n955 0.152939
R21376 gnd.n5726 gnd.n955 0.152939
R21377 gnd.n5727 gnd.n5726 0.152939
R21378 gnd.n5728 gnd.n5727 0.152939
R21379 gnd.n5728 gnd.n952 0.152939
R21380 gnd.n5733 gnd.n952 0.152939
R21381 gnd.n5734 gnd.n5733 0.152939
R21382 gnd.n5736 gnd.n5734 0.152939
R21383 gnd.n5736 gnd.n5735 0.152939
R21384 gnd.n5735 gnd.n890 0.152939
R21385 gnd.n5809 gnd.n890 0.152939
R21386 gnd.n5810 gnd.n5809 0.152939
R21387 gnd.n5839 gnd.n5810 0.152939
R21388 gnd.n5839 gnd.n5838 0.152939
R21389 gnd.n5838 gnd.n5837 0.152939
R21390 gnd.n5837 gnd.n5811 0.152939
R21391 gnd.n5833 gnd.n5811 0.152939
R21392 gnd.n5833 gnd.n5832 0.152939
R21393 gnd.n5832 gnd.n5831 0.152939
R21394 gnd.n5831 gnd.n5822 0.152939
R21395 gnd.n5827 gnd.n5822 0.152939
R21396 gnd.n5827 gnd.n5826 0.152939
R21397 gnd.n5826 gnd.n5825 0.152939
R21398 gnd.n5825 gnd.n810 0.152939
R21399 gnd.n5956 gnd.n810 0.152939
R21400 gnd.n5957 gnd.n5956 0.152939
R21401 gnd.n6047 gnd.n5957 0.152939
R21402 gnd.n6047 gnd.n6046 0.152939
R21403 gnd.n6046 gnd.n6045 0.152939
R21404 gnd.n6045 gnd.n5958 0.152939
R21405 gnd.n6041 gnd.n5958 0.152939
R21406 gnd.n6041 gnd.n6040 0.152939
R21407 gnd.n6040 gnd.n6039 0.152939
R21408 gnd.n6039 gnd.n5961 0.152939
R21409 gnd.n6035 gnd.n5961 0.152939
R21410 gnd.n6035 gnd.n6034 0.152939
R21411 gnd.n6034 gnd.n6033 0.152939
R21412 gnd.n6033 gnd.n5966 0.152939
R21413 gnd.n6029 gnd.n5966 0.152939
R21414 gnd.n6029 gnd.n6028 0.152939
R21415 gnd.n6028 gnd.n6027 0.152939
R21416 gnd.n6027 gnd.n6013 0.152939
R21417 gnd.n6023 gnd.n6013 0.152939
R21418 gnd.n6023 gnd.n6022 0.152939
R21419 gnd.n6022 gnd.n6021 0.152939
R21420 gnd.n6021 gnd.n6018 0.152939
R21421 gnd.n6018 gnd.n633 0.152939
R21422 gnd.n6375 gnd.n633 0.152939
R21423 gnd.n6376 gnd.n6375 0.152939
R21424 gnd.n6378 gnd.n6376 0.152939
R21425 gnd.n6378 gnd.n6377 0.152939
R21426 gnd.n6377 gnd.n608 0.152939
R21427 gnd.n6405 gnd.n608 0.152939
R21428 gnd.n6406 gnd.n6405 0.152939
R21429 gnd.n6408 gnd.n6406 0.152939
R21430 gnd.n6408 gnd.n6407 0.152939
R21431 gnd.n6407 gnd.n582 0.152939
R21432 gnd.n6435 gnd.n582 0.152939
R21433 gnd.n6436 gnd.n6435 0.152939
R21434 gnd.n6438 gnd.n6436 0.152939
R21435 gnd.n6438 gnd.n6437 0.152939
R21436 gnd.n4845 gnd.n4844 0.152939
R21437 gnd.n4844 gnd.n4837 0.152939
R21438 gnd.n4840 gnd.n4837 0.152939
R21439 gnd.n4840 gnd.n1339 0.152939
R21440 gnd.n4934 gnd.n1339 0.152939
R21441 gnd.n4935 gnd.n4934 0.152939
R21442 gnd.n4937 gnd.n4935 0.152939
R21443 gnd.n4937 gnd.n4936 0.152939
R21444 gnd.n4936 gnd.n1306 0.152939
R21445 gnd.n4987 gnd.n1306 0.152939
R21446 gnd.n4988 gnd.n4987 0.152939
R21447 gnd.n4993 gnd.n4988 0.152939
R21448 gnd.n4993 gnd.n4992 0.152939
R21449 gnd.n4992 gnd.n4991 0.152939
R21450 gnd.n4991 gnd.n1236 0.152939
R21451 gnd.n5343 gnd.n1236 0.152939
R21452 gnd.n5343 gnd.n5342 0.152939
R21453 gnd.n5342 gnd.n5341 0.152939
R21454 gnd.n5341 gnd.n1237 0.152939
R21455 gnd.n5337 gnd.n1237 0.152939
R21456 gnd.n5325 gnd.n1263 0.152939
R21457 gnd.n5325 gnd.n5324 0.152939
R21458 gnd.n5324 gnd.n5323 0.152939
R21459 gnd.n5323 gnd.n1265 0.152939
R21460 gnd.n5319 gnd.n1265 0.152939
R21461 gnd.n5319 gnd.n5318 0.152939
R21462 gnd.n5169 gnd.n5048 0.152939
R21463 gnd.n5169 gnd.n5168 0.152939
R21464 gnd.n5168 gnd.n5167 0.152939
R21465 gnd.n5167 gnd.n5049 0.152939
R21466 gnd.n5163 gnd.n5049 0.152939
R21467 gnd.n5163 gnd.n5162 0.152939
R21468 gnd.n5162 gnd.n5161 0.152939
R21469 gnd.n5161 gnd.n5054 0.152939
R21470 gnd.n5157 gnd.n5054 0.152939
R21471 gnd.n5157 gnd.n5156 0.152939
R21472 gnd.n5156 gnd.n5155 0.152939
R21473 gnd.n5155 gnd.n1075 0.152939
R21474 gnd.n5622 gnd.n1075 0.152939
R21475 gnd.n5623 gnd.n5622 0.152939
R21476 gnd.n5624 gnd.n5623 0.152939
R21477 gnd.n5624 gnd.n1002 0.152939
R21478 gnd.n5662 gnd.n1002 0.152939
R21479 gnd.n5663 gnd.n5662 0.152939
R21480 gnd.n5664 gnd.n5663 0.152939
R21481 gnd.n5664 gnd.n965 0.152939
R21482 gnd.n5717 gnd.n965 0.152939
R21483 gnd.n5718 gnd.n5717 0.152939
R21484 gnd.n5720 gnd.n5718 0.152939
R21485 gnd.n5720 gnd.n5719 0.152939
R21486 gnd.n5719 gnd.n930 0.152939
R21487 gnd.n5759 gnd.n930 0.152939
R21488 gnd.n5760 gnd.n5759 0.152939
R21489 gnd.n5761 gnd.n5760 0.152939
R21490 gnd.n5761 gnd.n897 0.152939
R21491 gnd.n5801 gnd.n897 0.152939
R21492 gnd.n5802 gnd.n5801 0.152939
R21493 gnd.n5803 gnd.n5802 0.152939
R21494 gnd.n5803 gnd.n882 0.152939
R21495 gnd.n5845 gnd.n882 0.152939
R21496 gnd.n5846 gnd.n5845 0.152939
R21497 gnd.n5847 gnd.n5846 0.152939
R21498 gnd.n5847 gnd.n852 0.152939
R21499 gnd.n5894 gnd.n852 0.152939
R21500 gnd.n5895 gnd.n5894 0.152939
R21501 gnd.n5897 gnd.n5895 0.152939
R21502 gnd.n5897 gnd.n5896 0.152939
R21503 gnd.n5896 gnd.n816 0.152939
R21504 gnd.n5947 gnd.n816 0.152939
R21505 gnd.n5948 gnd.n5947 0.152939
R21506 gnd.n5949 gnd.n5948 0.152939
R21507 gnd.n5949 gnd.n791 0.152939
R21508 gnd.n6072 gnd.n791 0.152939
R21509 gnd.n6073 gnd.n6072 0.152939
R21510 gnd.n6074 gnd.n6073 0.152939
R21511 gnd.n6074 gnd.n768 0.152939
R21512 gnd.n6100 gnd.n768 0.152939
R21513 gnd.n6101 gnd.n6100 0.152939
R21514 gnd.n6103 gnd.n6101 0.152939
R21515 gnd.n6103 gnd.n6102 0.152939
R21516 gnd.n6102 gnd.n738 0.152939
R21517 gnd.n6135 gnd.n738 0.152939
R21518 gnd.n6136 gnd.n6135 0.152939
R21519 gnd.n6137 gnd.n6136 0.152939
R21520 gnd.n6137 gnd.n714 0.152939
R21521 gnd.n6167 gnd.n714 0.152939
R21522 gnd.n6168 gnd.n6167 0.152939
R21523 gnd.n6176 gnd.n6168 0.152939
R21524 gnd.n6176 gnd.n6175 0.152939
R21525 gnd.n6175 gnd.n6174 0.152939
R21526 gnd.n6174 gnd.n6169 0.152939
R21527 gnd.n6169 gnd.n642 0.152939
R21528 gnd.n6366 gnd.n642 0.152939
R21529 gnd.n6367 gnd.n6366 0.152939
R21530 gnd.n6369 gnd.n6367 0.152939
R21531 gnd.n6369 gnd.n6368 0.152939
R21532 gnd.n6368 gnd.n617 0.152939
R21533 gnd.n6396 gnd.n617 0.152939
R21534 gnd.n6397 gnd.n6396 0.152939
R21535 gnd.n6399 gnd.n6397 0.152939
R21536 gnd.n6399 gnd.n6398 0.152939
R21537 gnd.n6398 gnd.n592 0.152939
R21538 gnd.n6426 gnd.n592 0.152939
R21539 gnd.n6427 gnd.n6426 0.152939
R21540 gnd.n6429 gnd.n6427 0.152939
R21541 gnd.n6429 gnd.n6428 0.152939
R21542 gnd.n6428 gnd.n568 0.152939
R21543 gnd.n6466 gnd.n568 0.152939
R21544 gnd.n6468 gnd.n6467 0.152939
R21545 gnd.n6468 gnd.n566 0.152939
R21546 gnd.n6476 gnd.n566 0.152939
R21547 gnd.n6477 gnd.n6476 0.152939
R21548 gnd.n6478 gnd.n6477 0.152939
R21549 gnd.n6478 gnd.n563 0.152939
R21550 gnd.n6712 gnd.n6711 0.152939
R21551 gnd.n6711 gnd.n379 0.152939
R21552 gnd.n6747 gnd.n379 0.152939
R21553 gnd.n6748 gnd.n6747 0.152939
R21554 gnd.n6750 gnd.n6748 0.152939
R21555 gnd.n6750 gnd.n6749 0.152939
R21556 gnd.n6749 gnd.n346 0.152939
R21557 gnd.n6816 gnd.n346 0.152939
R21558 gnd.n6817 gnd.n6816 0.152939
R21559 gnd.n6819 gnd.n6817 0.152939
R21560 gnd.n6819 gnd.n6818 0.152939
R21561 gnd.n6818 gnd.n317 0.152939
R21562 gnd.n6852 gnd.n317 0.152939
R21563 gnd.n6853 gnd.n6852 0.152939
R21564 gnd.n6862 gnd.n6853 0.152939
R21565 gnd.n6862 gnd.n6861 0.152939
R21566 gnd.n6861 gnd.n6860 0.152939
R21567 gnd.n6860 gnd.n6854 0.152939
R21568 gnd.n6856 gnd.n6854 0.152939
R21569 gnd.n6856 gnd.n63 0.152939
R21570 gnd.n7330 gnd.n7329 0.145814
R21571 gnd.n4846 gnd.n4835 0.145814
R21572 gnd.n4846 gnd.n4845 0.145814
R21573 gnd.n7330 gnd.n63 0.145814
R21574 gnd.n5318 gnd.n1208 0.128549
R21575 gnd.n6576 gnd.n563 0.128549
R21576 gnd.n3243 gnd.n0 0.127478
R21577 gnd.n7003 gnd.n79 0.10111
R21578 gnd.n4807 gnd.n1350 0.10111
R21579 gnd.n3823 gnd.n3822 0.0767195
R21580 gnd.n3822 gnd.n3821 0.0767195
R21581 gnd.n5463 gnd.n1208 0.063
R21582 gnd.n6577 gnd.n6576 0.063
R21583 gnd.n6577 gnd.n399 0.0538288
R21584 gnd.n7266 gnd.n174 0.0538288
R21585 gnd.n4588 gnd.n4587 0.0538288
R21586 gnd.n5463 gnd.n5462 0.0538288
R21587 gnd.n1396 gnd.n1350 0.0523293
R21588 gnd.n6772 gnd.n79 0.0523293
R21589 gnd.n4327 gnd.n3071 0.0477147
R21590 gnd.n3586 gnd.n3474 0.0442063
R21591 gnd.n3587 gnd.n3586 0.0442063
R21592 gnd.n3588 gnd.n3587 0.0442063
R21593 gnd.n3588 gnd.n3463 0.0442063
R21594 gnd.n3602 gnd.n3463 0.0442063
R21595 gnd.n3603 gnd.n3602 0.0442063
R21596 gnd.n3604 gnd.n3603 0.0442063
R21597 gnd.n3604 gnd.n3450 0.0442063
R21598 gnd.n3648 gnd.n3450 0.0442063
R21599 gnd.n3649 gnd.n3648 0.0442063
R21600 gnd.n3651 gnd.n3384 0.0344674
R21601 gnd.n6731 gnd.n399 0.0344674
R21602 gnd.n6731 gnd.n400 0.0344674
R21603 gnd.n402 gnd.n400 0.0344674
R21604 gnd.n406 gnd.n402 0.0344674
R21605 gnd.n407 gnd.n406 0.0344674
R21606 gnd.n407 gnd.n365 0.0344674
R21607 gnd.n366 gnd.n365 0.0344674
R21608 gnd.n6794 gnd.n366 0.0344674
R21609 gnd.n6795 gnd.n6794 0.0344674
R21610 gnd.n6795 gnd.n340 0.0344674
R21611 gnd.n340 gnd.n337 0.0344674
R21612 gnd.n338 gnd.n337 0.0344674
R21613 gnd.n6830 gnd.n338 0.0344674
R21614 gnd.n6830 gnd.n310 0.0344674
R21615 gnd.n6868 gnd.n310 0.0344674
R21616 gnd.n6869 gnd.n6868 0.0344674
R21617 gnd.n6869 gnd.n299 0.0344674
R21618 gnd.n6882 gnd.n299 0.0344674
R21619 gnd.n6882 gnd.n281 0.0344674
R21620 gnd.n6915 gnd.n281 0.0344674
R21621 gnd.n6916 gnd.n6915 0.0344674
R21622 gnd.n6916 gnd.n276 0.0344674
R21623 gnd.n276 gnd.n274 0.0344674
R21624 gnd.n6927 gnd.n274 0.0344674
R21625 gnd.n6928 gnd.n6927 0.0344674
R21626 gnd.n6928 gnd.n93 0.0344674
R21627 gnd.n94 gnd.n93 0.0344674
R21628 gnd.n95 gnd.n94 0.0344674
R21629 gnd.n6931 gnd.n95 0.0344674
R21630 gnd.n6931 gnd.n112 0.0344674
R21631 gnd.n113 gnd.n112 0.0344674
R21632 gnd.n114 gnd.n113 0.0344674
R21633 gnd.n6939 gnd.n114 0.0344674
R21634 gnd.n6939 gnd.n133 0.0344674
R21635 gnd.n134 gnd.n133 0.0344674
R21636 gnd.n135 gnd.n134 0.0344674
R21637 gnd.n6946 gnd.n135 0.0344674
R21638 gnd.n6946 gnd.n154 0.0344674
R21639 gnd.n155 gnd.n154 0.0344674
R21640 gnd.n156 gnd.n155 0.0344674
R21641 gnd.n173 gnd.n156 0.0344674
R21642 gnd.n7266 gnd.n173 0.0344674
R21643 gnd.n4587 gnd.n4523 0.0344674
R21644 gnd.n4523 gnd.n4522 0.0344674
R21645 gnd.n4522 gnd.n1498 0.0344674
R21646 gnd.n1498 gnd.n1496 0.0344674
R21647 gnd.n4733 gnd.n1496 0.0344674
R21648 gnd.n4734 gnd.n4733 0.0344674
R21649 gnd.n4734 gnd.n1473 0.0344674
R21650 gnd.n4763 gnd.n1473 0.0344674
R21651 gnd.n4763 gnd.n1457 0.0344674
R21652 gnd.n4777 gnd.n1457 0.0344674
R21653 gnd.n4778 gnd.n4777 0.0344674
R21654 gnd.n4778 gnd.n1438 0.0344674
R21655 gnd.n1439 gnd.n1438 0.0344674
R21656 gnd.n1440 gnd.n1439 0.0344674
R21657 gnd.n4781 gnd.n1440 0.0344674
R21658 gnd.n4784 gnd.n4781 0.0344674
R21659 gnd.n4785 gnd.n4784 0.0344674
R21660 gnd.n4785 gnd.n1365 0.0344674
R21661 gnd.n1366 gnd.n1365 0.0344674
R21662 gnd.n1367 gnd.n1366 0.0344674
R21663 gnd.n1408 gnd.n1367 0.0344674
R21664 gnd.n4872 gnd.n1408 0.0344674
R21665 gnd.n4877 gnd.n4872 0.0344674
R21666 gnd.n4878 gnd.n4877 0.0344674
R21667 gnd.n4878 gnd.n1403 0.0344674
R21668 gnd.n1404 gnd.n1403 0.0344674
R21669 gnd.n1405 gnd.n1404 0.0344674
R21670 gnd.n4888 gnd.n1405 0.0344674
R21671 gnd.n4888 gnd.n1406 0.0344674
R21672 gnd.n1406 gnd.n1325 0.0344674
R21673 gnd.n1326 gnd.n1325 0.0344674
R21674 gnd.n4965 gnd.n1326 0.0344674
R21675 gnd.n4966 gnd.n4965 0.0344674
R21676 gnd.n4966 gnd.n1300 0.0344674
R21677 gnd.n1300 gnd.n1298 0.0344674
R21678 gnd.n5002 gnd.n1298 0.0344674
R21679 gnd.n5003 gnd.n5002 0.0344674
R21680 gnd.n5003 gnd.n1229 0.0344674
R21681 gnd.n5350 gnd.n1229 0.0344674
R21682 gnd.n5351 gnd.n5350 0.0344674
R21683 gnd.n5351 gnd.n1209 0.0344674
R21684 gnd.n5462 gnd.n1209 0.0344674
R21685 gnd.n5315 gnd.n5314 0.0344674
R21686 gnd.n6575 gnd.n564 0.0344674
R21687 gnd.n5336 gnd.n5335 0.029712
R21688 gnd.n6710 gnd.n6709 0.029712
R21689 gnd.n3671 gnd.n3670 0.0269946
R21690 gnd.n3673 gnd.n3672 0.0269946
R21691 gnd.n3379 gnd.n3377 0.0269946
R21692 gnd.n3683 gnd.n3681 0.0269946
R21693 gnd.n3682 gnd.n3358 0.0269946
R21694 gnd.n3702 gnd.n3701 0.0269946
R21695 gnd.n3704 gnd.n3703 0.0269946
R21696 gnd.n3353 gnd.n3352 0.0269946
R21697 gnd.n3714 gnd.n3348 0.0269946
R21698 gnd.n3713 gnd.n3350 0.0269946
R21699 gnd.n3349 gnd.n3331 0.0269946
R21700 gnd.n3734 gnd.n3332 0.0269946
R21701 gnd.n3733 gnd.n3333 0.0269946
R21702 gnd.n3767 gnd.n3308 0.0269946
R21703 gnd.n3769 gnd.n3768 0.0269946
R21704 gnd.n3770 gnd.n3255 0.0269946
R21705 gnd.n3303 gnd.n3256 0.0269946
R21706 gnd.n3305 gnd.n3257 0.0269946
R21707 gnd.n3780 gnd.n3779 0.0269946
R21708 gnd.n3782 gnd.n3781 0.0269946
R21709 gnd.n3783 gnd.n3277 0.0269946
R21710 gnd.n3785 gnd.n3278 0.0269946
R21711 gnd.n3788 gnd.n3279 0.0269946
R21712 gnd.n3791 gnd.n3790 0.0269946
R21713 gnd.n3793 gnd.n3792 0.0269946
R21714 gnd.n3858 gnd.n3178 0.0269946
R21715 gnd.n3860 gnd.n3859 0.0269946
R21716 gnd.n3869 gnd.n3171 0.0269946
R21717 gnd.n3871 gnd.n3870 0.0269946
R21718 gnd.n3872 gnd.n3169 0.0269946
R21719 gnd.n3879 gnd.n3875 0.0269946
R21720 gnd.n3878 gnd.n3877 0.0269946
R21721 gnd.n3876 gnd.n3148 0.0269946
R21722 gnd.n3903 gnd.n3149 0.0269946
R21723 gnd.n3902 gnd.n3150 0.0269946
R21724 gnd.n3899 gnd.n2955 0.0269946
R21725 gnd.n3126 gnd.n2956 0.0269946
R21726 gnd.n3128 gnd.n2957 0.0269946
R21727 gnd.n3955 gnd.n3954 0.0269946
R21728 gnd.n3957 gnd.n3956 0.0269946
R21729 gnd.n3958 gnd.n2978 0.0269946
R21730 gnd.n3960 gnd.n2979 0.0269946
R21731 gnd.n3962 gnd.n2980 0.0269946
R21732 gnd.n3968 gnd.n3967 0.0269946
R21733 gnd.n3970 gnd.n3969 0.0269946
R21734 gnd.n3971 gnd.n3003 0.0269946
R21735 gnd.n3972 gnd.n3004 0.0269946
R21736 gnd.n3973 gnd.n3005 0.0269946
R21737 gnd.n4233 gnd.n4232 0.0269946
R21738 gnd.n4234 gnd.n3029 0.0269946
R21739 gnd.n4235 gnd.n3030 0.0269946
R21740 gnd.n4236 gnd.n3031 0.0269946
R21741 gnd.n5313 gnd.n1272 0.0225788
R21742 gnd.n5310 gnd.n5309 0.0225788
R21743 gnd.n5306 gnd.n5195 0.0225788
R21744 gnd.n5305 gnd.n5202 0.0225788
R21745 gnd.n5302 gnd.n5301 0.0225788
R21746 gnd.n5298 gnd.n5209 0.0225788
R21747 gnd.n5297 gnd.n5215 0.0225788
R21748 gnd.n5294 gnd.n5293 0.0225788
R21749 gnd.n5290 gnd.n5221 0.0225788
R21750 gnd.n5289 gnd.n5225 0.0225788
R21751 gnd.n5286 gnd.n5285 0.0225788
R21752 gnd.n5282 gnd.n5232 0.0225788
R21753 gnd.n5281 gnd.n5238 0.0225788
R21754 gnd.n5278 gnd.n5277 0.0225788
R21755 gnd.n5274 gnd.n5244 0.0225788
R21756 gnd.n5273 gnd.n5248 0.0225788
R21757 gnd.n5270 gnd.n5269 0.0225788
R21758 gnd.n5262 gnd.n5261 0.0225788
R21759 gnd.n5335 gnd.n1241 0.0225788
R21760 gnd.n6571 gnd.n6488 0.0225788
R21761 gnd.n6570 gnd.n6489 0.0225788
R21762 gnd.n6567 gnd.n6566 0.0225788
R21763 gnd.n6563 gnd.n6495 0.0225788
R21764 gnd.n6562 gnd.n6499 0.0225788
R21765 gnd.n6559 gnd.n6558 0.0225788
R21766 gnd.n6555 gnd.n6505 0.0225788
R21767 gnd.n6554 gnd.n6511 0.0225788
R21768 gnd.n6551 gnd.n6550 0.0225788
R21769 gnd.n6547 gnd.n6515 0.0225788
R21770 gnd.n6546 gnd.n6519 0.0225788
R21771 gnd.n6543 gnd.n6542 0.0225788
R21772 gnd.n6539 gnd.n6525 0.0225788
R21773 gnd.n6538 gnd.n6531 0.0225788
R21774 gnd.n6535 gnd.n6534 0.0225788
R21775 gnd.n6701 gnd.n449 0.0225788
R21776 gnd.n6700 gnd.n451 0.0225788
R21777 gnd.n456 gnd.n455 0.0225788
R21778 gnd.n6709 gnd.n423 0.0225788
R21779 gnd.n6710 gnd.n422 0.0218415
R21780 gnd.n5336 gnd.n1240 0.0218415
R21781 gnd.n3651 gnd.n3650 0.0202011
R21782 gnd.n3650 gnd.n3649 0.0148637
R21783 gnd.n4230 gnd.n3974 0.0144266
R21784 gnd.n4231 gnd.n4230 0.0130679
R21785 gnd.n5314 gnd.n5313 0.0123886
R21786 gnd.n5310 gnd.n1272 0.0123886
R21787 gnd.n5309 gnd.n5195 0.0123886
R21788 gnd.n5306 gnd.n5305 0.0123886
R21789 gnd.n5302 gnd.n5202 0.0123886
R21790 gnd.n5301 gnd.n5209 0.0123886
R21791 gnd.n5298 gnd.n5297 0.0123886
R21792 gnd.n5294 gnd.n5215 0.0123886
R21793 gnd.n5293 gnd.n5221 0.0123886
R21794 gnd.n5290 gnd.n5289 0.0123886
R21795 gnd.n5286 gnd.n5225 0.0123886
R21796 gnd.n5285 gnd.n5232 0.0123886
R21797 gnd.n5282 gnd.n5281 0.0123886
R21798 gnd.n5278 gnd.n5238 0.0123886
R21799 gnd.n5277 gnd.n5244 0.0123886
R21800 gnd.n5274 gnd.n5273 0.0123886
R21801 gnd.n5270 gnd.n5248 0.0123886
R21802 gnd.n5269 gnd.n5262 0.0123886
R21803 gnd.n5261 gnd.n1241 0.0123886
R21804 gnd.n6488 gnd.n564 0.0123886
R21805 gnd.n6571 gnd.n6570 0.0123886
R21806 gnd.n6567 gnd.n6489 0.0123886
R21807 gnd.n6566 gnd.n6495 0.0123886
R21808 gnd.n6563 gnd.n6562 0.0123886
R21809 gnd.n6559 gnd.n6499 0.0123886
R21810 gnd.n6558 gnd.n6505 0.0123886
R21811 gnd.n6555 gnd.n6554 0.0123886
R21812 gnd.n6551 gnd.n6511 0.0123886
R21813 gnd.n6550 gnd.n6515 0.0123886
R21814 gnd.n6547 gnd.n6546 0.0123886
R21815 gnd.n6543 gnd.n6519 0.0123886
R21816 gnd.n6542 gnd.n6525 0.0123886
R21817 gnd.n6539 gnd.n6538 0.0123886
R21818 gnd.n6535 gnd.n6531 0.0123886
R21819 gnd.n6534 gnd.n449 0.0123886
R21820 gnd.n6701 gnd.n6700 0.0123886
R21821 gnd.n456 gnd.n451 0.0123886
R21822 gnd.n455 gnd.n423 0.0123886
R21823 gnd.n3670 gnd.n3384 0.00797283
R21824 gnd.n3672 gnd.n3671 0.00797283
R21825 gnd.n3673 gnd.n3379 0.00797283
R21826 gnd.n3681 gnd.n3377 0.00797283
R21827 gnd.n3683 gnd.n3682 0.00797283
R21828 gnd.n3701 gnd.n3358 0.00797283
R21829 gnd.n3703 gnd.n3702 0.00797283
R21830 gnd.n3704 gnd.n3353 0.00797283
R21831 gnd.n3352 gnd.n3348 0.00797283
R21832 gnd.n3714 gnd.n3713 0.00797283
R21833 gnd.n3350 gnd.n3349 0.00797283
R21834 gnd.n3332 gnd.n3331 0.00797283
R21835 gnd.n3734 gnd.n3733 0.00797283
R21836 gnd.n3333 gnd.n3308 0.00797283
R21837 gnd.n3768 gnd.n3767 0.00797283
R21838 gnd.n3770 gnd.n3769 0.00797283
R21839 gnd.n3303 gnd.n3255 0.00797283
R21840 gnd.n3305 gnd.n3256 0.00797283
R21841 gnd.n3779 gnd.n3257 0.00797283
R21842 gnd.n3781 gnd.n3780 0.00797283
R21843 gnd.n3783 gnd.n3782 0.00797283
R21844 gnd.n3785 gnd.n3277 0.00797283
R21845 gnd.n3788 gnd.n3278 0.00797283
R21846 gnd.n3790 gnd.n3279 0.00797283
R21847 gnd.n3793 gnd.n3791 0.00797283
R21848 gnd.n3792 gnd.n3178 0.00797283
R21849 gnd.n3860 gnd.n3858 0.00797283
R21850 gnd.n3859 gnd.n3171 0.00797283
R21851 gnd.n3870 gnd.n3869 0.00797283
R21852 gnd.n3872 gnd.n3871 0.00797283
R21853 gnd.n3875 gnd.n3169 0.00797283
R21854 gnd.n3879 gnd.n3878 0.00797283
R21855 gnd.n3877 gnd.n3876 0.00797283
R21856 gnd.n3149 gnd.n3148 0.00797283
R21857 gnd.n3903 gnd.n3902 0.00797283
R21858 gnd.n3899 gnd.n3150 0.00797283
R21859 gnd.n3126 gnd.n2955 0.00797283
R21860 gnd.n3128 gnd.n2956 0.00797283
R21861 gnd.n3954 gnd.n2957 0.00797283
R21862 gnd.n3956 gnd.n3955 0.00797283
R21863 gnd.n3958 gnd.n3957 0.00797283
R21864 gnd.n3960 gnd.n2978 0.00797283
R21865 gnd.n3962 gnd.n2979 0.00797283
R21866 gnd.n3967 gnd.n2980 0.00797283
R21867 gnd.n3969 gnd.n3968 0.00797283
R21868 gnd.n3971 gnd.n3970 0.00797283
R21869 gnd.n3972 gnd.n3003 0.00797283
R21870 gnd.n3973 gnd.n3004 0.00797283
R21871 gnd.n3974 gnd.n3005 0.00797283
R21872 gnd.n4232 gnd.n4231 0.00797283
R21873 gnd.n4234 gnd.n4233 0.00797283
R21874 gnd.n4235 gnd.n3029 0.00797283
R21875 gnd.n4236 gnd.n3030 0.00797283
R21876 gnd.n3071 gnd.n3031 0.00797283
R21877 gnd.n5315 gnd.n1208 0.00593478
R21878 gnd.n6576 gnd.n6575 0.00593478
R21879 a_n2318_13878.n59 a_n2318_13878.t82 533.335
R21880 a_n2318_13878.n75 a_n2318_13878.t63 512.366
R21881 a_n2318_13878.n70 a_n2318_13878.t67 512.366
R21882 a_n2318_13878.n74 a_n2318_13878.t57 512.366
R21883 a_n2318_13878.n73 a_n2318_13878.t72 512.366
R21884 a_n2318_13878.n71 a_n2318_13878.t79 512.366
R21885 a_n2318_13878.n72 a_n2318_13878.t80 512.366
R21886 a_n2318_13878.n53 a_n2318_13878.t20 533.335
R21887 a_n2318_13878.n89 a_n2318_13878.t26 512.366
R21888 a_n2318_13878.n68 a_n2318_13878.t42 512.366
R21889 a_n2318_13878.n88 a_n2318_13878.t44 512.366
R21890 a_n2318_13878.n87 a_n2318_13878.t22 512.366
R21891 a_n2318_13878.n69 a_n2318_13878.t38 512.366
R21892 a_n2318_13878.n86 a_n2318_13878.t32 512.366
R21893 a_n2318_13878.n37 a_n2318_13878.t40 533.335
R21894 a_n2318_13878.n112 a_n2318_13878.t34 512.366
R21895 a_n2318_13878.n113 a_n2318_13878.t30 512.366
R21896 a_n2318_13878.n114 a_n2318_13878.t46 512.366
R21897 a_n2318_13878.n115 a_n2318_13878.t18 512.366
R21898 a_n2318_13878.n66 a_n2318_13878.t36 512.366
R21899 a_n2318_13878.n116 a_n2318_13878.t24 512.366
R21900 a_n2318_13878.n30 a_n2318_13878.t78 533.335
R21901 a_n2318_13878.n107 a_n2318_13878.t56 512.366
R21902 a_n2318_13878.n108 a_n2318_13878.t75 512.366
R21903 a_n2318_13878.n109 a_n2318_13878.t76 512.366
R21904 a_n2318_13878.n110 a_n2318_13878.t53 512.366
R21905 a_n2318_13878.n67 a_n2318_13878.t62 512.366
R21906 a_n2318_13878.n111 a_n2318_13878.t71 512.366
R21907 a_n2318_13878.n99 a_n2318_13878.t69 512.366
R21908 a_n2318_13878.n98 a_n2318_13878.t60 512.366
R21909 a_n2318_13878.n97 a_n2318_13878.t52 512.366
R21910 a_n2318_13878.n101 a_n2318_13878.t77 512.366
R21911 a_n2318_13878.n100 a_n2318_13878.t66 512.366
R21912 a_n2318_13878.n96 a_n2318_13878.t65 512.366
R21913 a_n2318_13878.n103 a_n2318_13878.t73 512.366
R21914 a_n2318_13878.n102 a_n2318_13878.t58 512.366
R21915 a_n2318_13878.n95 a_n2318_13878.t59 512.366
R21916 a_n2318_13878.n105 a_n2318_13878.t61 512.366
R21917 a_n2318_13878.n104 a_n2318_13878.t70 512.366
R21918 a_n2318_13878.n94 a_n2318_13878.t83 512.366
R21919 a_n2318_13878.n64 a_n2318_13878.n1 70.1674
R21920 a_n2318_13878.n58 a_n2318_13878.n5 70.1674
R21921 a_n2318_13878.n16 a_n2318_13878.n43 70.1674
R21922 a_n2318_13878.n19 a_n2318_13878.n36 70.1674
R21923 a_n2318_13878.n111 a_n2318_13878.n36 20.9683
R21924 a_n2318_13878.n35 a_n2318_13878.n20 72.3034
R21925 a_n2318_13878.n35 a_n2318_13878.n67 16.6962
R21926 a_n2318_13878.n20 a_n2318_13878.n34 77.6622
R21927 a_n2318_13878.n110 a_n2318_13878.n34 5.97853
R21928 a_n2318_13878.n33 a_n2318_13878.n21 77.6622
R21929 a_n2318_13878.n21 a_n2318_13878.n32 72.3034
R21930 a_n2318_13878.n107 a_n2318_13878.n30 20.9683
R21931 a_n2318_13878.n31 a_n2318_13878.n30 70.1674
R21932 a_n2318_13878.n116 a_n2318_13878.n43 20.9683
R21933 a_n2318_13878.n42 a_n2318_13878.n17 72.3034
R21934 a_n2318_13878.n42 a_n2318_13878.n66 16.6962
R21935 a_n2318_13878.n17 a_n2318_13878.n41 77.6622
R21936 a_n2318_13878.n115 a_n2318_13878.n41 5.97853
R21937 a_n2318_13878.n40 a_n2318_13878.n18 77.6622
R21938 a_n2318_13878.n18 a_n2318_13878.n39 72.3034
R21939 a_n2318_13878.n112 a_n2318_13878.n37 20.9683
R21940 a_n2318_13878.n38 a_n2318_13878.n37 70.1674
R21941 a_n2318_13878.n8 a_n2318_13878.n52 70.1674
R21942 a_n2318_13878.n10 a_n2318_13878.n49 70.1674
R21943 a_n2318_13878.n12 a_n2318_13878.n47 70.1674
R21944 a_n2318_13878.n14 a_n2318_13878.n45 70.1674
R21945 a_n2318_13878.n45 a_n2318_13878.n94 20.9683
R21946 a_n2318_13878.n44 a_n2318_13878.n15 75.0448
R21947 a_n2318_13878.n104 a_n2318_13878.n44 11.2134
R21948 a_n2318_13878.n15 a_n2318_13878.n105 161.3
R21949 a_n2318_13878.n47 a_n2318_13878.n95 20.9683
R21950 a_n2318_13878.n46 a_n2318_13878.n13 75.0448
R21951 a_n2318_13878.n102 a_n2318_13878.n46 11.2134
R21952 a_n2318_13878.n13 a_n2318_13878.n103 161.3
R21953 a_n2318_13878.n49 a_n2318_13878.n96 20.9683
R21954 a_n2318_13878.n48 a_n2318_13878.n11 75.0448
R21955 a_n2318_13878.n100 a_n2318_13878.n48 11.2134
R21956 a_n2318_13878.n11 a_n2318_13878.n101 161.3
R21957 a_n2318_13878.n52 a_n2318_13878.n97 20.9683
R21958 a_n2318_13878.n50 a_n2318_13878.n9 75.0448
R21959 a_n2318_13878.n98 a_n2318_13878.n50 11.2134
R21960 a_n2318_13878.n9 a_n2318_13878.n99 161.3
R21961 a_n2318_13878.n86 a_n2318_13878.n58 20.9683
R21962 a_n2318_13878.n6 a_n2318_13878.n57 72.3034
R21963 a_n2318_13878.n57 a_n2318_13878.n69 16.6962
R21964 a_n2318_13878.n56 a_n2318_13878.n6 77.6622
R21965 a_n2318_13878.n87 a_n2318_13878.n56 5.97853
R21966 a_n2318_13878.n55 a_n2318_13878.n4 77.6622
R21967 a_n2318_13878.n4 a_n2318_13878.n54 72.3034
R21968 a_n2318_13878.n89 a_n2318_13878.n53 20.9683
R21969 a_n2318_13878.n7 a_n2318_13878.n53 70.1674
R21970 a_n2318_13878.n72 a_n2318_13878.n64 20.9683
R21971 a_n2318_13878.n2 a_n2318_13878.n63 72.3034
R21972 a_n2318_13878.n63 a_n2318_13878.n71 16.6962
R21973 a_n2318_13878.n62 a_n2318_13878.n2 77.6622
R21974 a_n2318_13878.n73 a_n2318_13878.n62 5.97853
R21975 a_n2318_13878.n61 a_n2318_13878.n0 77.6622
R21976 a_n2318_13878.n0 a_n2318_13878.n60 72.3034
R21977 a_n2318_13878.n75 a_n2318_13878.n59 20.9683
R21978 a_n2318_13878.n3 a_n2318_13878.n59 70.1674
R21979 a_n2318_13878.n25 a_n2318_13878.n84 81.2902
R21980 a_n2318_13878.n23 a_n2318_13878.n79 81.2902
R21981 a_n2318_13878.n22 a_n2318_13878.n76 81.2902
R21982 a_n2318_13878.n25 a_n2318_13878.n85 80.9324
R21983 a_n2318_13878.n25 a_n2318_13878.n83 80.9324
R21984 a_n2318_13878.n24 a_n2318_13878.n82 80.9324
R21985 a_n2318_13878.n24 a_n2318_13878.n81 80.9324
R21986 a_n2318_13878.n23 a_n2318_13878.n80 80.9324
R21987 a_n2318_13878.n23 a_n2318_13878.n78 80.9324
R21988 a_n2318_13878.n22 a_n2318_13878.n77 80.9324
R21989 a_n2318_13878.n29 a_n2318_13878.t41 74.6477
R21990 a_n2318_13878.n26 a_n2318_13878.t29 74.6477
R21991 a_n2318_13878.n27 a_n2318_13878.t21 74.2899
R21992 a_n2318_13878.n28 a_n2318_13878.t49 74.2897
R21993 a_n2318_13878.n28 a_n2318_13878.n118 70.6783
R21994 a_n2318_13878.n29 a_n2318_13878.n65 70.6783
R21995 a_n2318_13878.n26 a_n2318_13878.n90 70.6783
R21996 a_n2318_13878.n26 a_n2318_13878.n91 70.6783
R21997 a_n2318_13878.n27 a_n2318_13878.n92 70.6783
R21998 a_n2318_13878.n119 a_n2318_13878.n29 70.6782
R21999 a_n2318_13878.n74 a_n2318_13878.n73 48.2005
R22000 a_n2318_13878.n64 a_n2318_13878.t54 533.335
R22001 a_n2318_13878.n88 a_n2318_13878.n87 48.2005
R22002 a_n2318_13878.n58 a_n2318_13878.t28 533.335
R22003 a_n2318_13878.n115 a_n2318_13878.n114 48.2005
R22004 a_n2318_13878.t48 a_n2318_13878.n43 533.335
R22005 a_n2318_13878.n110 a_n2318_13878.n109 48.2005
R22006 a_n2318_13878.t55 a_n2318_13878.n36 533.335
R22007 a_n2318_13878.n99 a_n2318_13878.n98 48.2005
R22008 a_n2318_13878.t74 a_n2318_13878.n52 533.335
R22009 a_n2318_13878.n101 a_n2318_13878.n100 48.2005
R22010 a_n2318_13878.t81 a_n2318_13878.n49 533.335
R22011 a_n2318_13878.n103 a_n2318_13878.n102 48.2005
R22012 a_n2318_13878.t68 a_n2318_13878.n47 533.335
R22013 a_n2318_13878.n105 a_n2318_13878.n104 48.2005
R22014 a_n2318_13878.t64 a_n2318_13878.n45 533.335
R22015 a_n2318_13878.n60 a_n2318_13878.n70 16.6962
R22016 a_n2318_13878.n72 a_n2318_13878.n63 27.6507
R22017 a_n2318_13878.n54 a_n2318_13878.n68 16.6962
R22018 a_n2318_13878.n86 a_n2318_13878.n57 27.6507
R22019 a_n2318_13878.n113 a_n2318_13878.n39 16.6962
R22020 a_n2318_13878.n116 a_n2318_13878.n42 27.6507
R22021 a_n2318_13878.n108 a_n2318_13878.n32 16.6962
R22022 a_n2318_13878.n111 a_n2318_13878.n35 27.6507
R22023 a_n2318_13878.n61 a_n2318_13878.n70 41.7634
R22024 a_n2318_13878.n55 a_n2318_13878.n68 41.7634
R22025 a_n2318_13878.n113 a_n2318_13878.n40 41.7634
R22026 a_n2318_13878.n108 a_n2318_13878.n33 41.7634
R22027 a_n2318_13878.n24 a_n2318_13878.n23 31.238
R22028 a_n2318_13878.n50 a_n2318_13878.n97 35.3134
R22029 a_n2318_13878.n48 a_n2318_13878.n96 35.3134
R22030 a_n2318_13878.n46 a_n2318_13878.n95 35.3134
R22031 a_n2318_13878.n44 a_n2318_13878.n94 35.3134
R22032 a_n2318_13878.n5 a_n2318_13878.n25 23.891
R22033 a_n2318_13878.n31 a_n2318_13878.n106 12.705
R22034 a_n2318_13878.n1 a_n2318_13878.n51 12.5005
R22035 a_n2318_13878.n61 a_n2318_13878.n74 5.97853
R22036 a_n2318_13878.n62 a_n2318_13878.n71 41.7634
R22037 a_n2318_13878.n55 a_n2318_13878.n88 5.97853
R22038 a_n2318_13878.n56 a_n2318_13878.n69 41.7634
R22039 a_n2318_13878.n114 a_n2318_13878.n40 5.97853
R22040 a_n2318_13878.n66 a_n2318_13878.n41 41.7634
R22041 a_n2318_13878.n109 a_n2318_13878.n33 5.97853
R22042 a_n2318_13878.n67 a_n2318_13878.n34 41.7634
R22043 a_n2318_13878.n93 a_n2318_13878.n7 11.1956
R22044 a_n2318_13878.n75 a_n2318_13878.n60 27.6507
R22045 a_n2318_13878.n89 a_n2318_13878.n54 27.6507
R22046 a_n2318_13878.n39 a_n2318_13878.n112 27.6507
R22047 a_n2318_13878.n32 a_n2318_13878.n107 27.6507
R22048 a_n2318_13878.n28 a_n2318_13878.n117 9.85898
R22049 a_n2318_13878.n8 a_n2318_13878.n51 8.73345
R22050 a_n2318_13878.n106 a_n2318_13878.n15 8.73345
R22051 a_n2318_13878.n117 a_n2318_13878.n16 7.36035
R22052 a_n2318_13878.n93 a_n2318_13878.n27 6.01559
R22053 a_n2318_13878.n117 a_n2318_13878.n51 5.3452
R22054 a_n2318_13878.n38 a_n2318_13878.n19 4.01186
R22055 a_n2318_13878.n5 a_n2318_13878.n3 3.76565
R22056 a_n2318_13878.n118 a_n2318_13878.t37 3.61217
R22057 a_n2318_13878.n118 a_n2318_13878.t25 3.61217
R22058 a_n2318_13878.n65 a_n2318_13878.t35 3.61217
R22059 a_n2318_13878.n65 a_n2318_13878.t31 3.61217
R22060 a_n2318_13878.n90 a_n2318_13878.t39 3.61217
R22061 a_n2318_13878.n90 a_n2318_13878.t33 3.61217
R22062 a_n2318_13878.n91 a_n2318_13878.t45 3.61217
R22063 a_n2318_13878.n91 a_n2318_13878.t23 3.61217
R22064 a_n2318_13878.n92 a_n2318_13878.t27 3.61217
R22065 a_n2318_13878.n92 a_n2318_13878.t43 3.61217
R22066 a_n2318_13878.n119 a_n2318_13878.t47 3.61217
R22067 a_n2318_13878.t19 a_n2318_13878.n119 3.61217
R22068 a_n2318_13878.n84 a_n2318_13878.t0 2.82907
R22069 a_n2318_13878.n84 a_n2318_13878.t6 2.82907
R22070 a_n2318_13878.n85 a_n2318_13878.t8 2.82907
R22071 a_n2318_13878.n85 a_n2318_13878.t13 2.82907
R22072 a_n2318_13878.n83 a_n2318_13878.t11 2.82907
R22073 a_n2318_13878.n83 a_n2318_13878.t12 2.82907
R22074 a_n2318_13878.n82 a_n2318_13878.t7 2.82907
R22075 a_n2318_13878.n82 a_n2318_13878.t16 2.82907
R22076 a_n2318_13878.n81 a_n2318_13878.t50 2.82907
R22077 a_n2318_13878.n81 a_n2318_13878.t10 2.82907
R22078 a_n2318_13878.n79 a_n2318_13878.t4 2.82907
R22079 a_n2318_13878.n79 a_n2318_13878.t14 2.82907
R22080 a_n2318_13878.n80 a_n2318_13878.t51 2.82907
R22081 a_n2318_13878.n80 a_n2318_13878.t9 2.82907
R22082 a_n2318_13878.n78 a_n2318_13878.t3 2.82907
R22083 a_n2318_13878.n78 a_n2318_13878.t5 2.82907
R22084 a_n2318_13878.n77 a_n2318_13878.t2 2.82907
R22085 a_n2318_13878.n77 a_n2318_13878.t15 2.82907
R22086 a_n2318_13878.n76 a_n2318_13878.t1 2.82907
R22087 a_n2318_13878.n76 a_n2318_13878.t17 2.82907
R22088 a_n2318_13878.n106 a_n2318_13878.n93 1.30542
R22089 a_n2318_13878.n29 a_n2318_13878.n28 1.07378
R22090 a_n2318_13878.n27 a_n2318_13878.n26 1.07378
R22091 a_n2318_13878.n25 a_n2318_13878.n24 1.07378
R22092 a_n2318_13878.n12 a_n2318_13878.n11 1.04595
R22093 a_n2318_13878.n6 a_n2318_13878.n5 0.966409
R22094 a_n2318_13878.n21 a_n2318_13878.n20 0.758076
R22095 a_n2318_13878.n20 a_n2318_13878.n19 0.758076
R22096 a_n2318_13878.n18 a_n2318_13878.n17 0.758076
R22097 a_n2318_13878.n17 a_n2318_13878.n16 0.758076
R22098 a_n2318_13878.n15 a_n2318_13878.n14 0.758076
R22099 a_n2318_13878.n13 a_n2318_13878.n12 0.758076
R22100 a_n2318_13878.n11 a_n2318_13878.n10 0.758076
R22101 a_n2318_13878.n9 a_n2318_13878.n8 0.758076
R22102 a_n2318_13878.n6 a_n2318_13878.n4 0.758076
R22103 a_n2318_13878.n2 a_n2318_13878.n0 0.758076
R22104 a_n2318_13878.n2 a_n2318_13878.n1 0.758076
R22105 a_n2318_13878.n23 a_n2318_13878.n22 0.716017
R22106 a_n2318_13878.n14 a_n2318_13878.n13 0.67853
R22107 a_n2318_13878.n10 a_n2318_13878.n9 0.67853
R22108 a_n2318_13878.n0 a_n2318_13878.n3 0.568682
R22109 a_n2318_13878.n4 a_n2318_13878.n7 0.568682
R22110 a_n2318_13878.n38 a_n2318_13878.n18 0.568682
R22111 a_n2318_13878.n31 a_n2318_13878.n21 0.568682
R22112 a_n2140_13878.n21 a_n2140_13878.n20 98.9632
R22113 a_n2140_13878.n2 a_n2140_13878.n0 98.7517
R22114 a_n2140_13878.n18 a_n2140_13878.n17 98.6055
R22115 a_n2140_13878.n20 a_n2140_13878.n19 98.6055
R22116 a_n2140_13878.n6 a_n2140_13878.n5 98.6055
R22117 a_n2140_13878.n4 a_n2140_13878.n3 98.6055
R22118 a_n2140_13878.n2 a_n2140_13878.n1 98.6055
R22119 a_n2140_13878.n16 a_n2140_13878.n15 98.6054
R22120 a_n2140_13878.n8 a_n2140_13878.t17 74.6477
R22121 a_n2140_13878.n13 a_n2140_13878.t18 74.2899
R22122 a_n2140_13878.n10 a_n2140_13878.t19 74.2899
R22123 a_n2140_13878.n9 a_n2140_13878.t16 74.2899
R22124 a_n2140_13878.n12 a_n2140_13878.n11 70.6783
R22125 a_n2140_13878.n8 a_n2140_13878.n7 70.6783
R22126 a_n2140_13878.n14 a_n2140_13878.n6 14.2849
R22127 a_n2140_13878.n16 a_n2140_13878.n14 11.9339
R22128 a_n2140_13878.n14 a_n2140_13878.n13 6.95632
R22129 a_n2140_13878.n15 a_n2140_13878.t6 3.61217
R22130 a_n2140_13878.n15 a_n2140_13878.t7 3.61217
R22131 a_n2140_13878.n17 a_n2140_13878.t13 3.61217
R22132 a_n2140_13878.n17 a_n2140_13878.t14 3.61217
R22133 a_n2140_13878.n19 a_n2140_13878.t0 3.61217
R22134 a_n2140_13878.n19 a_n2140_13878.t8 3.61217
R22135 a_n2140_13878.n11 a_n2140_13878.t22 3.61217
R22136 a_n2140_13878.n11 a_n2140_13878.t23 3.61217
R22137 a_n2140_13878.n7 a_n2140_13878.t20 3.61217
R22138 a_n2140_13878.n7 a_n2140_13878.t21 3.61217
R22139 a_n2140_13878.n5 a_n2140_13878.t9 3.61217
R22140 a_n2140_13878.n5 a_n2140_13878.t1 3.61217
R22141 a_n2140_13878.n3 a_n2140_13878.t12 3.61217
R22142 a_n2140_13878.n3 a_n2140_13878.t3 3.61217
R22143 a_n2140_13878.n1 a_n2140_13878.t2 3.61217
R22144 a_n2140_13878.n1 a_n2140_13878.t4 3.61217
R22145 a_n2140_13878.n0 a_n2140_13878.t10 3.61217
R22146 a_n2140_13878.n0 a_n2140_13878.t5 3.61217
R22147 a_n2140_13878.n21 a_n2140_13878.t11 3.61217
R22148 a_n2140_13878.t15 a_n2140_13878.n21 3.61217
R22149 a_n2140_13878.n9 a_n2140_13878.n8 0.358259
R22150 a_n2140_13878.n12 a_n2140_13878.n10 0.358259
R22151 a_n2140_13878.n13 a_n2140_13878.n12 0.358259
R22152 a_n2140_13878.n20 a_n2140_13878.n18 0.358259
R22153 a_n2140_13878.n18 a_n2140_13878.n16 0.358259
R22154 a_n2140_13878.n4 a_n2140_13878.n2 0.146627
R22155 a_n2140_13878.n6 a_n2140_13878.n4 0.146627
R22156 a_n2140_13878.n10 a_n2140_13878.n9 0.101793
R22157 outputibias.n27 outputibias.n1 289.615
R22158 outputibias.n58 outputibias.n32 289.615
R22159 outputibias.n90 outputibias.n64 289.615
R22160 outputibias.n122 outputibias.n96 289.615
R22161 outputibias.n28 outputibias.n27 185
R22162 outputibias.n26 outputibias.n25 185
R22163 outputibias.n5 outputibias.n4 185
R22164 outputibias.n20 outputibias.n19 185
R22165 outputibias.n18 outputibias.n17 185
R22166 outputibias.n9 outputibias.n8 185
R22167 outputibias.n12 outputibias.n11 185
R22168 outputibias.n59 outputibias.n58 185
R22169 outputibias.n57 outputibias.n56 185
R22170 outputibias.n36 outputibias.n35 185
R22171 outputibias.n51 outputibias.n50 185
R22172 outputibias.n49 outputibias.n48 185
R22173 outputibias.n40 outputibias.n39 185
R22174 outputibias.n43 outputibias.n42 185
R22175 outputibias.n91 outputibias.n90 185
R22176 outputibias.n89 outputibias.n88 185
R22177 outputibias.n68 outputibias.n67 185
R22178 outputibias.n83 outputibias.n82 185
R22179 outputibias.n81 outputibias.n80 185
R22180 outputibias.n72 outputibias.n71 185
R22181 outputibias.n75 outputibias.n74 185
R22182 outputibias.n123 outputibias.n122 185
R22183 outputibias.n121 outputibias.n120 185
R22184 outputibias.n100 outputibias.n99 185
R22185 outputibias.n115 outputibias.n114 185
R22186 outputibias.n113 outputibias.n112 185
R22187 outputibias.n104 outputibias.n103 185
R22188 outputibias.n107 outputibias.n106 185
R22189 outputibias.n0 outputibias.t9 178.945
R22190 outputibias.n133 outputibias.t8 177.018
R22191 outputibias.n132 outputibias.t11 177.018
R22192 outputibias.n0 outputibias.t10 177.018
R22193 outputibias.t5 outputibias.n10 147.661
R22194 outputibias.t7 outputibias.n41 147.661
R22195 outputibias.t1 outputibias.n73 147.661
R22196 outputibias.t3 outputibias.n105 147.661
R22197 outputibias.n128 outputibias.t4 132.363
R22198 outputibias.n128 outputibias.t6 130.436
R22199 outputibias.n129 outputibias.t0 130.436
R22200 outputibias.n130 outputibias.t2 130.436
R22201 outputibias.n27 outputibias.n26 104.615
R22202 outputibias.n26 outputibias.n4 104.615
R22203 outputibias.n19 outputibias.n4 104.615
R22204 outputibias.n19 outputibias.n18 104.615
R22205 outputibias.n18 outputibias.n8 104.615
R22206 outputibias.n11 outputibias.n8 104.615
R22207 outputibias.n58 outputibias.n57 104.615
R22208 outputibias.n57 outputibias.n35 104.615
R22209 outputibias.n50 outputibias.n35 104.615
R22210 outputibias.n50 outputibias.n49 104.615
R22211 outputibias.n49 outputibias.n39 104.615
R22212 outputibias.n42 outputibias.n39 104.615
R22213 outputibias.n90 outputibias.n89 104.615
R22214 outputibias.n89 outputibias.n67 104.615
R22215 outputibias.n82 outputibias.n67 104.615
R22216 outputibias.n82 outputibias.n81 104.615
R22217 outputibias.n81 outputibias.n71 104.615
R22218 outputibias.n74 outputibias.n71 104.615
R22219 outputibias.n122 outputibias.n121 104.615
R22220 outputibias.n121 outputibias.n99 104.615
R22221 outputibias.n114 outputibias.n99 104.615
R22222 outputibias.n114 outputibias.n113 104.615
R22223 outputibias.n113 outputibias.n103 104.615
R22224 outputibias.n106 outputibias.n103 104.615
R22225 outputibias.n63 outputibias.n31 95.6354
R22226 outputibias.n63 outputibias.n62 94.6732
R22227 outputibias.n95 outputibias.n94 94.6732
R22228 outputibias.n127 outputibias.n126 94.6732
R22229 outputibias.n11 outputibias.t5 52.3082
R22230 outputibias.n42 outputibias.t7 52.3082
R22231 outputibias.n74 outputibias.t1 52.3082
R22232 outputibias.n106 outputibias.t3 52.3082
R22233 outputibias.n12 outputibias.n10 15.6674
R22234 outputibias.n43 outputibias.n41 15.6674
R22235 outputibias.n75 outputibias.n73 15.6674
R22236 outputibias.n107 outputibias.n105 15.6674
R22237 outputibias.n13 outputibias.n9 12.8005
R22238 outputibias.n44 outputibias.n40 12.8005
R22239 outputibias.n76 outputibias.n72 12.8005
R22240 outputibias.n108 outputibias.n104 12.8005
R22241 outputibias.n17 outputibias.n16 12.0247
R22242 outputibias.n48 outputibias.n47 12.0247
R22243 outputibias.n80 outputibias.n79 12.0247
R22244 outputibias.n112 outputibias.n111 12.0247
R22245 outputibias.n20 outputibias.n7 11.249
R22246 outputibias.n51 outputibias.n38 11.249
R22247 outputibias.n83 outputibias.n70 11.249
R22248 outputibias.n115 outputibias.n102 11.249
R22249 outputibias.n21 outputibias.n5 10.4732
R22250 outputibias.n52 outputibias.n36 10.4732
R22251 outputibias.n84 outputibias.n68 10.4732
R22252 outputibias.n116 outputibias.n100 10.4732
R22253 outputibias.n25 outputibias.n24 9.69747
R22254 outputibias.n56 outputibias.n55 9.69747
R22255 outputibias.n88 outputibias.n87 9.69747
R22256 outputibias.n120 outputibias.n119 9.69747
R22257 outputibias.n31 outputibias.n30 9.45567
R22258 outputibias.n62 outputibias.n61 9.45567
R22259 outputibias.n94 outputibias.n93 9.45567
R22260 outputibias.n126 outputibias.n125 9.45567
R22261 outputibias.n30 outputibias.n29 9.3005
R22262 outputibias.n3 outputibias.n2 9.3005
R22263 outputibias.n24 outputibias.n23 9.3005
R22264 outputibias.n22 outputibias.n21 9.3005
R22265 outputibias.n7 outputibias.n6 9.3005
R22266 outputibias.n16 outputibias.n15 9.3005
R22267 outputibias.n14 outputibias.n13 9.3005
R22268 outputibias.n61 outputibias.n60 9.3005
R22269 outputibias.n34 outputibias.n33 9.3005
R22270 outputibias.n55 outputibias.n54 9.3005
R22271 outputibias.n53 outputibias.n52 9.3005
R22272 outputibias.n38 outputibias.n37 9.3005
R22273 outputibias.n47 outputibias.n46 9.3005
R22274 outputibias.n45 outputibias.n44 9.3005
R22275 outputibias.n93 outputibias.n92 9.3005
R22276 outputibias.n66 outputibias.n65 9.3005
R22277 outputibias.n87 outputibias.n86 9.3005
R22278 outputibias.n85 outputibias.n84 9.3005
R22279 outputibias.n70 outputibias.n69 9.3005
R22280 outputibias.n79 outputibias.n78 9.3005
R22281 outputibias.n77 outputibias.n76 9.3005
R22282 outputibias.n125 outputibias.n124 9.3005
R22283 outputibias.n98 outputibias.n97 9.3005
R22284 outputibias.n119 outputibias.n118 9.3005
R22285 outputibias.n117 outputibias.n116 9.3005
R22286 outputibias.n102 outputibias.n101 9.3005
R22287 outputibias.n111 outputibias.n110 9.3005
R22288 outputibias.n109 outputibias.n108 9.3005
R22289 outputibias.n28 outputibias.n3 8.92171
R22290 outputibias.n59 outputibias.n34 8.92171
R22291 outputibias.n91 outputibias.n66 8.92171
R22292 outputibias.n123 outputibias.n98 8.92171
R22293 outputibias.n29 outputibias.n1 8.14595
R22294 outputibias.n60 outputibias.n32 8.14595
R22295 outputibias.n92 outputibias.n64 8.14595
R22296 outputibias.n124 outputibias.n96 8.14595
R22297 outputibias.n31 outputibias.n1 5.81868
R22298 outputibias.n62 outputibias.n32 5.81868
R22299 outputibias.n94 outputibias.n64 5.81868
R22300 outputibias.n126 outputibias.n96 5.81868
R22301 outputibias.n131 outputibias.n130 5.20947
R22302 outputibias.n29 outputibias.n28 5.04292
R22303 outputibias.n60 outputibias.n59 5.04292
R22304 outputibias.n92 outputibias.n91 5.04292
R22305 outputibias.n124 outputibias.n123 5.04292
R22306 outputibias.n131 outputibias.n127 4.42209
R22307 outputibias.n14 outputibias.n10 4.38594
R22308 outputibias.n45 outputibias.n41 4.38594
R22309 outputibias.n77 outputibias.n73 4.38594
R22310 outputibias.n109 outputibias.n105 4.38594
R22311 outputibias.n132 outputibias.n131 4.28454
R22312 outputibias.n25 outputibias.n3 4.26717
R22313 outputibias.n56 outputibias.n34 4.26717
R22314 outputibias.n88 outputibias.n66 4.26717
R22315 outputibias.n120 outputibias.n98 4.26717
R22316 outputibias.n24 outputibias.n5 3.49141
R22317 outputibias.n55 outputibias.n36 3.49141
R22318 outputibias.n87 outputibias.n68 3.49141
R22319 outputibias.n119 outputibias.n100 3.49141
R22320 outputibias.n21 outputibias.n20 2.71565
R22321 outputibias.n52 outputibias.n51 2.71565
R22322 outputibias.n84 outputibias.n83 2.71565
R22323 outputibias.n116 outputibias.n115 2.71565
R22324 outputibias.n17 outputibias.n7 1.93989
R22325 outputibias.n48 outputibias.n38 1.93989
R22326 outputibias.n80 outputibias.n70 1.93989
R22327 outputibias.n112 outputibias.n102 1.93989
R22328 outputibias.n130 outputibias.n129 1.9266
R22329 outputibias.n129 outputibias.n128 1.9266
R22330 outputibias.n133 outputibias.n132 1.92658
R22331 outputibias.n134 outputibias.n133 1.29913
R22332 outputibias.n16 outputibias.n9 1.16414
R22333 outputibias.n47 outputibias.n40 1.16414
R22334 outputibias.n79 outputibias.n72 1.16414
R22335 outputibias.n111 outputibias.n104 1.16414
R22336 outputibias.n127 outputibias.n95 0.962709
R22337 outputibias.n95 outputibias.n63 0.962709
R22338 outputibias.n13 outputibias.n12 0.388379
R22339 outputibias.n44 outputibias.n43 0.388379
R22340 outputibias.n76 outputibias.n75 0.388379
R22341 outputibias.n108 outputibias.n107 0.388379
R22342 outputibias.n134 outputibias.n0 0.337251
R22343 outputibias outputibias.n134 0.302375
R22344 outputibias.n30 outputibias.n2 0.155672
R22345 outputibias.n23 outputibias.n2 0.155672
R22346 outputibias.n23 outputibias.n22 0.155672
R22347 outputibias.n22 outputibias.n6 0.155672
R22348 outputibias.n15 outputibias.n6 0.155672
R22349 outputibias.n15 outputibias.n14 0.155672
R22350 outputibias.n61 outputibias.n33 0.155672
R22351 outputibias.n54 outputibias.n33 0.155672
R22352 outputibias.n54 outputibias.n53 0.155672
R22353 outputibias.n53 outputibias.n37 0.155672
R22354 outputibias.n46 outputibias.n37 0.155672
R22355 outputibias.n46 outputibias.n45 0.155672
R22356 outputibias.n93 outputibias.n65 0.155672
R22357 outputibias.n86 outputibias.n65 0.155672
R22358 outputibias.n86 outputibias.n85 0.155672
R22359 outputibias.n85 outputibias.n69 0.155672
R22360 outputibias.n78 outputibias.n69 0.155672
R22361 outputibias.n78 outputibias.n77 0.155672
R22362 outputibias.n125 outputibias.n97 0.155672
R22363 outputibias.n118 outputibias.n97 0.155672
R22364 outputibias.n118 outputibias.n117 0.155672
R22365 outputibias.n117 outputibias.n101 0.155672
R22366 outputibias.n110 outputibias.n101 0.155672
R22367 outputibias.n110 outputibias.n109 0.155672
R22368 output.n41 output.n15 289.615
R22369 output.n72 output.n46 289.615
R22370 output.n104 output.n78 289.615
R22371 output.n136 output.n110 289.615
R22372 output.n77 output.n45 197.26
R22373 output.n77 output.n76 196.298
R22374 output.n109 output.n108 196.298
R22375 output.n141 output.n140 196.298
R22376 output.n42 output.n41 185
R22377 output.n40 output.n39 185
R22378 output.n19 output.n18 185
R22379 output.n34 output.n33 185
R22380 output.n32 output.n31 185
R22381 output.n23 output.n22 185
R22382 output.n26 output.n25 185
R22383 output.n73 output.n72 185
R22384 output.n71 output.n70 185
R22385 output.n50 output.n49 185
R22386 output.n65 output.n64 185
R22387 output.n63 output.n62 185
R22388 output.n54 output.n53 185
R22389 output.n57 output.n56 185
R22390 output.n105 output.n104 185
R22391 output.n103 output.n102 185
R22392 output.n82 output.n81 185
R22393 output.n97 output.n96 185
R22394 output.n95 output.n94 185
R22395 output.n86 output.n85 185
R22396 output.n89 output.n88 185
R22397 output.n137 output.n136 185
R22398 output.n135 output.n134 185
R22399 output.n114 output.n113 185
R22400 output.n129 output.n128 185
R22401 output.n127 output.n126 185
R22402 output.n118 output.n117 185
R22403 output.n121 output.n120 185
R22404 output.t2 output.n24 147.661
R22405 output.t1 output.n55 147.661
R22406 output.t3 output.n87 147.661
R22407 output.t0 output.n119 147.661
R22408 output.n41 output.n40 104.615
R22409 output.n40 output.n18 104.615
R22410 output.n33 output.n18 104.615
R22411 output.n33 output.n32 104.615
R22412 output.n32 output.n22 104.615
R22413 output.n25 output.n22 104.615
R22414 output.n72 output.n71 104.615
R22415 output.n71 output.n49 104.615
R22416 output.n64 output.n49 104.615
R22417 output.n64 output.n63 104.615
R22418 output.n63 output.n53 104.615
R22419 output.n56 output.n53 104.615
R22420 output.n104 output.n103 104.615
R22421 output.n103 output.n81 104.615
R22422 output.n96 output.n81 104.615
R22423 output.n96 output.n95 104.615
R22424 output.n95 output.n85 104.615
R22425 output.n88 output.n85 104.615
R22426 output.n136 output.n135 104.615
R22427 output.n135 output.n113 104.615
R22428 output.n128 output.n113 104.615
R22429 output.n128 output.n127 104.615
R22430 output.n127 output.n117 104.615
R22431 output.n120 output.n117 104.615
R22432 output.n1 output.t8 77.056
R22433 output.n14 output.t9 76.6694
R22434 output.n1 output.n0 72.7095
R22435 output.n3 output.n2 72.7095
R22436 output.n5 output.n4 72.7095
R22437 output.n7 output.n6 72.7095
R22438 output.n9 output.n8 72.7095
R22439 output.n11 output.n10 72.7095
R22440 output.n13 output.n12 72.7095
R22441 output.n25 output.t2 52.3082
R22442 output.n56 output.t1 52.3082
R22443 output.n88 output.t3 52.3082
R22444 output.n120 output.t0 52.3082
R22445 output.n26 output.n24 15.6674
R22446 output.n57 output.n55 15.6674
R22447 output.n89 output.n87 15.6674
R22448 output.n121 output.n119 15.6674
R22449 output.n27 output.n23 12.8005
R22450 output.n58 output.n54 12.8005
R22451 output.n90 output.n86 12.8005
R22452 output.n122 output.n118 12.8005
R22453 output.n31 output.n30 12.0247
R22454 output.n62 output.n61 12.0247
R22455 output.n94 output.n93 12.0247
R22456 output.n126 output.n125 12.0247
R22457 output.n34 output.n21 11.249
R22458 output.n65 output.n52 11.249
R22459 output.n97 output.n84 11.249
R22460 output.n129 output.n116 11.249
R22461 output.n35 output.n19 10.4732
R22462 output.n66 output.n50 10.4732
R22463 output.n98 output.n82 10.4732
R22464 output.n130 output.n114 10.4732
R22465 output.n39 output.n38 9.69747
R22466 output.n70 output.n69 9.69747
R22467 output.n102 output.n101 9.69747
R22468 output.n134 output.n133 9.69747
R22469 output.n45 output.n44 9.45567
R22470 output.n76 output.n75 9.45567
R22471 output.n108 output.n107 9.45567
R22472 output.n140 output.n139 9.45567
R22473 output.n44 output.n43 9.3005
R22474 output.n17 output.n16 9.3005
R22475 output.n38 output.n37 9.3005
R22476 output.n36 output.n35 9.3005
R22477 output.n21 output.n20 9.3005
R22478 output.n30 output.n29 9.3005
R22479 output.n28 output.n27 9.3005
R22480 output.n75 output.n74 9.3005
R22481 output.n48 output.n47 9.3005
R22482 output.n69 output.n68 9.3005
R22483 output.n67 output.n66 9.3005
R22484 output.n52 output.n51 9.3005
R22485 output.n61 output.n60 9.3005
R22486 output.n59 output.n58 9.3005
R22487 output.n107 output.n106 9.3005
R22488 output.n80 output.n79 9.3005
R22489 output.n101 output.n100 9.3005
R22490 output.n99 output.n98 9.3005
R22491 output.n84 output.n83 9.3005
R22492 output.n93 output.n92 9.3005
R22493 output.n91 output.n90 9.3005
R22494 output.n139 output.n138 9.3005
R22495 output.n112 output.n111 9.3005
R22496 output.n133 output.n132 9.3005
R22497 output.n131 output.n130 9.3005
R22498 output.n116 output.n115 9.3005
R22499 output.n125 output.n124 9.3005
R22500 output.n123 output.n122 9.3005
R22501 output.n42 output.n17 8.92171
R22502 output.n73 output.n48 8.92171
R22503 output.n105 output.n80 8.92171
R22504 output.n137 output.n112 8.92171
R22505 output output.n141 8.15037
R22506 output.n43 output.n15 8.14595
R22507 output.n74 output.n46 8.14595
R22508 output.n106 output.n78 8.14595
R22509 output.n138 output.n110 8.14595
R22510 output.n45 output.n15 5.81868
R22511 output.n76 output.n46 5.81868
R22512 output.n108 output.n78 5.81868
R22513 output.n140 output.n110 5.81868
R22514 output.n43 output.n42 5.04292
R22515 output.n74 output.n73 5.04292
R22516 output.n106 output.n105 5.04292
R22517 output.n138 output.n137 5.04292
R22518 output.n28 output.n24 4.38594
R22519 output.n59 output.n55 4.38594
R22520 output.n91 output.n87 4.38594
R22521 output.n123 output.n119 4.38594
R22522 output.n39 output.n17 4.26717
R22523 output.n70 output.n48 4.26717
R22524 output.n102 output.n80 4.26717
R22525 output.n134 output.n112 4.26717
R22526 output.n0 output.t14 3.9605
R22527 output.n0 output.t18 3.9605
R22528 output.n2 output.t5 3.9605
R22529 output.n2 output.t10 3.9605
R22530 output.n4 output.t11 3.9605
R22531 output.n4 output.t16 3.9605
R22532 output.n6 output.t4 3.9605
R22533 output.n6 output.t12 3.9605
R22534 output.n8 output.t15 3.9605
R22535 output.n8 output.t13 3.9605
R22536 output.n10 output.t19 3.9605
R22537 output.n10 output.t6 3.9605
R22538 output.n12 output.t7 3.9605
R22539 output.n12 output.t17 3.9605
R22540 output.n38 output.n19 3.49141
R22541 output.n69 output.n50 3.49141
R22542 output.n101 output.n82 3.49141
R22543 output.n133 output.n114 3.49141
R22544 output.n35 output.n34 2.71565
R22545 output.n66 output.n65 2.71565
R22546 output.n98 output.n97 2.71565
R22547 output.n130 output.n129 2.71565
R22548 output.n31 output.n21 1.93989
R22549 output.n62 output.n52 1.93989
R22550 output.n94 output.n84 1.93989
R22551 output.n126 output.n116 1.93989
R22552 output.n30 output.n23 1.16414
R22553 output.n61 output.n54 1.16414
R22554 output.n93 output.n86 1.16414
R22555 output.n125 output.n118 1.16414
R22556 output.n141 output.n109 0.962709
R22557 output.n109 output.n77 0.962709
R22558 output.n27 output.n26 0.388379
R22559 output.n58 output.n57 0.388379
R22560 output.n90 output.n89 0.388379
R22561 output.n122 output.n121 0.388379
R22562 output.n14 output.n13 0.387128
R22563 output.n13 output.n11 0.387128
R22564 output.n11 output.n9 0.387128
R22565 output.n9 output.n7 0.387128
R22566 output.n7 output.n5 0.387128
R22567 output.n5 output.n3 0.387128
R22568 output.n3 output.n1 0.387128
R22569 output.n44 output.n16 0.155672
R22570 output.n37 output.n16 0.155672
R22571 output.n37 output.n36 0.155672
R22572 output.n36 output.n20 0.155672
R22573 output.n29 output.n20 0.155672
R22574 output.n29 output.n28 0.155672
R22575 output.n75 output.n47 0.155672
R22576 output.n68 output.n47 0.155672
R22577 output.n68 output.n67 0.155672
R22578 output.n67 output.n51 0.155672
R22579 output.n60 output.n51 0.155672
R22580 output.n60 output.n59 0.155672
R22581 output.n107 output.n79 0.155672
R22582 output.n100 output.n79 0.155672
R22583 output.n100 output.n99 0.155672
R22584 output.n99 output.n83 0.155672
R22585 output.n92 output.n83 0.155672
R22586 output.n92 output.n91 0.155672
R22587 output.n139 output.n111 0.155672
R22588 output.n132 output.n111 0.155672
R22589 output.n132 output.n131 0.155672
R22590 output.n131 output.n115 0.155672
R22591 output.n124 output.n115 0.155672
R22592 output.n124 output.n123 0.155672
R22593 output output.n14 0.126227
R22594 a_n2318_8322.n8 a_n2318_8322.t19 74.6477
R22595 a_n2318_8322.n1 a_n2318_8322.t14 74.6477
R22596 a_n2318_8322.n20 a_n2318_8322.t13 74.6474
R22597 a_n2318_8322.n16 a_n2318_8322.t3 74.2899
R22598 a_n2318_8322.n9 a_n2318_8322.t17 74.2899
R22599 a_n2318_8322.n10 a_n2318_8322.t20 74.2899
R22600 a_n2318_8322.n13 a_n2318_8322.t21 74.2899
R22601 a_n2318_8322.n6 a_n2318_8322.t0 74.2899
R22602 a_n2318_8322.n20 a_n2318_8322.n19 70.6783
R22603 a_n2318_8322.n18 a_n2318_8322.n17 70.6783
R22604 a_n2318_8322.n8 a_n2318_8322.n7 70.6783
R22605 a_n2318_8322.n12 a_n2318_8322.n11 70.6783
R22606 a_n2318_8322.n1 a_n2318_8322.n0 70.6783
R22607 a_n2318_8322.n3 a_n2318_8322.n2 70.6783
R22608 a_n2318_8322.n5 a_n2318_8322.n4 70.6783
R22609 a_n2318_8322.n22 a_n2318_8322.n21 70.6782
R22610 a_n2318_8322.n14 a_n2318_8322.n6 23.4712
R22611 a_n2318_8322.n15 a_n2318_8322.t26 9.69317
R22612 a_n2318_8322.n14 a_n2318_8322.n13 6.95632
R22613 a_n2318_8322.n16 a_n2318_8322.n15 6.19447
R22614 a_n2318_8322.n15 a_n2318_8322.n14 5.3452
R22615 a_n2318_8322.n19 a_n2318_8322.t10 3.61217
R22616 a_n2318_8322.n19 a_n2318_8322.t7 3.61217
R22617 a_n2318_8322.n17 a_n2318_8322.t12 3.61217
R22618 a_n2318_8322.n17 a_n2318_8322.t5 3.61217
R22619 a_n2318_8322.n7 a_n2318_8322.t23 3.61217
R22620 a_n2318_8322.n7 a_n2318_8322.t22 3.61217
R22621 a_n2318_8322.n11 a_n2318_8322.t18 3.61217
R22622 a_n2318_8322.n11 a_n2318_8322.t16 3.61217
R22623 a_n2318_8322.n0 a_n2318_8322.t2 3.61217
R22624 a_n2318_8322.n0 a_n2318_8322.t1 3.61217
R22625 a_n2318_8322.n2 a_n2318_8322.t11 3.61217
R22626 a_n2318_8322.n2 a_n2318_8322.t6 3.61217
R22627 a_n2318_8322.n4 a_n2318_8322.t9 3.61217
R22628 a_n2318_8322.n4 a_n2318_8322.t8 3.61217
R22629 a_n2318_8322.n22 a_n2318_8322.t4 3.61217
R22630 a_n2318_8322.t15 a_n2318_8322.n22 3.61217
R22631 a_n2318_8322.n13 a_n2318_8322.n12 0.358259
R22632 a_n2318_8322.n12 a_n2318_8322.n10 0.358259
R22633 a_n2318_8322.n9 a_n2318_8322.n8 0.358259
R22634 a_n2318_8322.n6 a_n2318_8322.n5 0.358259
R22635 a_n2318_8322.n5 a_n2318_8322.n3 0.358259
R22636 a_n2318_8322.n3 a_n2318_8322.n1 0.358259
R22637 a_n2318_8322.n18 a_n2318_8322.n16 0.358259
R22638 a_n2318_8322.n21 a_n2318_8322.n18 0.358259
R22639 a_n2318_8322.n21 a_n2318_8322.n20 0.358259
R22640 a_n2318_8322.n10 a_n2318_8322.n9 0.101793
R22641 a_n2318_8322.t27 a_n2318_8322.t24 0.0788333
R22642 a_n2318_8322.t25 a_n2318_8322.t27 0.0631667
R22643 a_n2318_8322.t26 a_n2318_8322.t25 0.0471944
R22644 a_n2318_8322.t26 a_n2318_8322.t24 0.0453889
R22645 plus.n34 plus.t22 436.949
R22646 plus.n8 plus.t12 436.949
R22647 plus.n35 plus.t5 415.966
R22648 plus.n33 plus.t19 415.966
R22649 plus.n41 plus.t23 415.966
R22650 plus.n42 plus.t11 415.966
R22651 plus.n46 plus.t6 415.966
R22652 plus.n47 plus.t10 415.966
R22653 plus.n29 plus.t18 415.966
R22654 plus.n53 plus.t8 415.966
R22655 plus.n54 plus.t15 415.966
R22656 plus.n26 plus.t24 415.966
R22657 plus.n25 plus.t20 415.966
R22658 plus.n1 plus.t7 415.966
R22659 plus.n19 plus.t17 415.966
R22660 plus.n18 plus.t13 415.966
R22661 plus.n4 plus.t21 415.966
R22662 plus.n13 plus.t16 415.966
R22663 plus.n11 plus.t9 415.966
R22664 plus.n7 plus.t14 415.966
R22665 plus.n58 plus.t0 243.97
R22666 plus.n58 plus.n57 223.454
R22667 plus.n60 plus.n59 223.454
R22668 plus.n55 plus.n54 161.3
R22669 plus.n53 plus.n28 161.3
R22670 plus.n52 plus.n51 161.3
R22671 plus.n50 plus.n29 161.3
R22672 plus.n49 plus.n48 161.3
R22673 plus.n47 plus.n30 161.3
R22674 plus.n46 plus.n45 161.3
R22675 plus.n44 plus.n31 161.3
R22676 plus.n43 plus.n42 161.3
R22677 plus.n41 plus.n32 161.3
R22678 plus.n40 plus.n39 161.3
R22679 plus.n38 plus.n33 161.3
R22680 plus.n37 plus.n36 161.3
R22681 plus.n10 plus.n9 161.3
R22682 plus.n11 plus.n6 161.3
R22683 plus.n12 plus.n5 161.3
R22684 plus.n14 plus.n13 161.3
R22685 plus.n15 plus.n4 161.3
R22686 plus.n17 plus.n16 161.3
R22687 plus.n18 plus.n3 161.3
R22688 plus.n19 plus.n2 161.3
R22689 plus.n21 plus.n20 161.3
R22690 plus.n22 plus.n1 161.3
R22691 plus.n24 plus.n23 161.3
R22692 plus.n25 plus.n0 161.3
R22693 plus.n27 plus.n26 161.3
R22694 plus.n37 plus.n34 70.4033
R22695 plus.n9 plus.n8 70.4033
R22696 plus.n42 plus.n41 48.2005
R22697 plus.n47 plus.n46 48.2005
R22698 plus.n54 plus.n53 48.2005
R22699 plus.n26 plus.n25 48.2005
R22700 plus.n19 plus.n18 48.2005
R22701 plus.n13 plus.n4 48.2005
R22702 plus.n40 plus.n33 47.4702
R22703 plus.n48 plus.n29 47.4702
R22704 plus.n20 plus.n1 47.4702
R22705 plus.n12 plus.n11 47.4702
R22706 plus.n56 plus.n55 29.8622
R22707 plus.n36 plus.n33 25.5611
R22708 plus.n52 plus.n29 25.5611
R22709 plus.n24 plus.n1 25.5611
R22710 plus.n11 plus.n10 25.5611
R22711 plus.n42 plus.n31 24.1005
R22712 plus.n46 plus.n31 24.1005
R22713 plus.n18 plus.n17 24.1005
R22714 plus.n17 plus.n4 24.1005
R22715 plus.n36 plus.n35 22.6399
R22716 plus.n53 plus.n52 22.6399
R22717 plus.n25 plus.n24 22.6399
R22718 plus.n10 plus.n7 22.6399
R22719 plus.n35 plus.n34 20.9576
R22720 plus.n8 plus.n7 20.9576
R22721 plus.n57 plus.t3 19.8005
R22722 plus.n57 plus.t2 19.8005
R22723 plus.n59 plus.t4 19.8005
R22724 plus.n59 plus.t1 19.8005
R22725 plus plus.n61 13.9746
R22726 plus.n56 plus.n27 11.7903
R22727 plus.n61 plus.n60 5.40567
R22728 plus.n61 plus.n56 1.188
R22729 plus.n41 plus.n40 0.730803
R22730 plus.n48 plus.n47 0.730803
R22731 plus.n20 plus.n19 0.730803
R22732 plus.n13 plus.n12 0.730803
R22733 plus.n60 plus.n58 0.716017
R22734 plus.n38 plus.n37 0.189894
R22735 plus.n39 plus.n38 0.189894
R22736 plus.n39 plus.n32 0.189894
R22737 plus.n43 plus.n32 0.189894
R22738 plus.n44 plus.n43 0.189894
R22739 plus.n45 plus.n44 0.189894
R22740 plus.n45 plus.n30 0.189894
R22741 plus.n49 plus.n30 0.189894
R22742 plus.n50 plus.n49 0.189894
R22743 plus.n51 plus.n50 0.189894
R22744 plus.n51 plus.n28 0.189894
R22745 plus.n55 plus.n28 0.189894
R22746 plus.n27 plus.n0 0.189894
R22747 plus.n23 plus.n0 0.189894
R22748 plus.n23 plus.n22 0.189894
R22749 plus.n22 plus.n21 0.189894
R22750 plus.n21 plus.n2 0.189894
R22751 plus.n3 plus.n2 0.189894
R22752 plus.n16 plus.n3 0.189894
R22753 plus.n16 plus.n15 0.189894
R22754 plus.n15 plus.n14 0.189894
R22755 plus.n14 plus.n5 0.189894
R22756 plus.n6 plus.n5 0.189894
R22757 plus.n9 plus.n6 0.189894
R22758 a_n2903_n3924.n12 a_n2903_n3924.t47 214.994
R22759 a_n2903_n3924.n1 a_n2903_n3924.t30 214.733
R22760 a_n2903_n3924.n13 a_n2903_n3924.t35 214.321
R22761 a_n2903_n3924.n14 a_n2903_n3924.t38 214.321
R22762 a_n2903_n3924.n15 a_n2903_n3924.t37 214.321
R22763 a_n2903_n3924.n16 a_n2903_n3924.t1 214.321
R22764 a_n2903_n3924.n17 a_n2903_n3924.t41 214.321
R22765 a_n2903_n3924.n12 a_n2903_n3924.t31 214.321
R22766 a_n2903_n3924.n0 a_n2903_n3924.t12 55.8337
R22767 a_n2903_n3924.n2 a_n2903_n3924.t7 55.8337
R22768 a_n2903_n3924.n11 a_n2903_n3924.t45 55.8337
R22769 a_n2903_n3924.n41 a_n2903_n3924.t19 55.8335
R22770 a_n2903_n3924.n39 a_n2903_n3924.t40 55.8335
R22771 a_n2903_n3924.n30 a_n2903_n3924.t2 55.8335
R22772 a_n2903_n3924.n29 a_n2903_n3924.t22 55.8335
R22773 a_n2903_n3924.n20 a_n2903_n3924.t10 55.8335
R22774 a_n2903_n3924.n43 a_n2903_n3924.n42 53.0052
R22775 a_n2903_n3924.n45 a_n2903_n3924.n44 53.0052
R22776 a_n2903_n3924.n47 a_n2903_n3924.n46 53.0052
R22777 a_n2903_n3924.n4 a_n2903_n3924.n3 53.0052
R22778 a_n2903_n3924.n6 a_n2903_n3924.n5 53.0052
R22779 a_n2903_n3924.n8 a_n2903_n3924.n7 53.0052
R22780 a_n2903_n3924.n10 a_n2903_n3924.n9 53.0052
R22781 a_n2903_n3924.n38 a_n2903_n3924.n37 53.0051
R22782 a_n2903_n3924.n36 a_n2903_n3924.n35 53.0051
R22783 a_n2903_n3924.n34 a_n2903_n3924.n33 53.0051
R22784 a_n2903_n3924.n32 a_n2903_n3924.n31 53.0051
R22785 a_n2903_n3924.n28 a_n2903_n3924.n27 53.0051
R22786 a_n2903_n3924.n26 a_n2903_n3924.n25 53.0051
R22787 a_n2903_n3924.n24 a_n2903_n3924.n23 53.0051
R22788 a_n2903_n3924.n22 a_n2903_n3924.n21 53.0051
R22789 a_n2903_n3924.n49 a_n2903_n3924.n48 53.0051
R22790 a_n2903_n3924.n19 a_n2903_n3924.n11 12.1555
R22791 a_n2903_n3924.n41 a_n2903_n3924.n40 12.1555
R22792 a_n2903_n3924.n20 a_n2903_n3924.n19 5.07593
R22793 a_n2903_n3924.n40 a_n2903_n3924.n39 5.07593
R22794 a_n2903_n3924.n42 a_n2903_n3924.t16 2.82907
R22795 a_n2903_n3924.n42 a_n2903_n3924.t26 2.82907
R22796 a_n2903_n3924.n44 a_n2903_n3924.t28 2.82907
R22797 a_n2903_n3924.n44 a_n2903_n3924.t24 2.82907
R22798 a_n2903_n3924.n46 a_n2903_n3924.t11 2.82907
R22799 a_n2903_n3924.n46 a_n2903_n3924.t23 2.82907
R22800 a_n2903_n3924.n3 a_n2903_n3924.t39 2.82907
R22801 a_n2903_n3924.n3 a_n2903_n3924.t0 2.82907
R22802 a_n2903_n3924.n5 a_n2903_n3924.t36 2.82907
R22803 a_n2903_n3924.n5 a_n2903_n3924.t9 2.82907
R22804 a_n2903_n3924.n7 a_n2903_n3924.t43 2.82907
R22805 a_n2903_n3924.n7 a_n2903_n3924.t34 2.82907
R22806 a_n2903_n3924.n9 a_n2903_n3924.t33 2.82907
R22807 a_n2903_n3924.n9 a_n2903_n3924.t8 2.82907
R22808 a_n2903_n3924.n37 a_n2903_n3924.t32 2.82907
R22809 a_n2903_n3924.n37 a_n2903_n3924.t5 2.82907
R22810 a_n2903_n3924.n35 a_n2903_n3924.t6 2.82907
R22811 a_n2903_n3924.n35 a_n2903_n3924.t46 2.82907
R22812 a_n2903_n3924.n33 a_n2903_n3924.t42 2.82907
R22813 a_n2903_n3924.n33 a_n2903_n3924.t4 2.82907
R22814 a_n2903_n3924.n31 a_n2903_n3924.t44 2.82907
R22815 a_n2903_n3924.n31 a_n2903_n3924.t3 2.82907
R22816 a_n2903_n3924.n27 a_n2903_n3924.t25 2.82907
R22817 a_n2903_n3924.n27 a_n2903_n3924.t20 2.82907
R22818 a_n2903_n3924.n25 a_n2903_n3924.t13 2.82907
R22819 a_n2903_n3924.n25 a_n2903_n3924.t18 2.82907
R22820 a_n2903_n3924.n23 a_n2903_n3924.t17 2.82907
R22821 a_n2903_n3924.n23 a_n2903_n3924.t21 2.82907
R22822 a_n2903_n3924.n21 a_n2903_n3924.t14 2.82907
R22823 a_n2903_n3924.n21 a_n2903_n3924.t27 2.82907
R22824 a_n2903_n3924.t29 a_n2903_n3924.n49 2.82907
R22825 a_n2903_n3924.n49 a_n2903_n3924.t15 2.82907
R22826 a_n2903_n3924.n40 a_n2903_n3924.n1 1.95694
R22827 a_n2903_n3924.n19 a_n2903_n3924.n18 1.95694
R22828 a_n2903_n3924.n17 a_n2903_n3924.n16 0.672012
R22829 a_n2903_n3924.n16 a_n2903_n3924.n15 0.672012
R22830 a_n2903_n3924.n15 a_n2903_n3924.n14 0.672012
R22831 a_n2903_n3924.n14 a_n2903_n3924.n13 0.672012
R22832 a_n2903_n3924.n18 a_n2903_n3924.n17 0.40239
R22833 a_n2903_n3924.n22 a_n2903_n3924.n20 0.358259
R22834 a_n2903_n3924.n24 a_n2903_n3924.n22 0.358259
R22835 a_n2903_n3924.n26 a_n2903_n3924.n24 0.358259
R22836 a_n2903_n3924.n28 a_n2903_n3924.n26 0.358259
R22837 a_n2903_n3924.n29 a_n2903_n3924.n28 0.358259
R22838 a_n2903_n3924.n32 a_n2903_n3924.n30 0.358259
R22839 a_n2903_n3924.n34 a_n2903_n3924.n32 0.358259
R22840 a_n2903_n3924.n36 a_n2903_n3924.n34 0.358259
R22841 a_n2903_n3924.n38 a_n2903_n3924.n36 0.358259
R22842 a_n2903_n3924.n39 a_n2903_n3924.n38 0.358259
R22843 a_n2903_n3924.n11 a_n2903_n3924.n10 0.358259
R22844 a_n2903_n3924.n10 a_n2903_n3924.n8 0.358259
R22845 a_n2903_n3924.n8 a_n2903_n3924.n6 0.358259
R22846 a_n2903_n3924.n6 a_n2903_n3924.n4 0.358259
R22847 a_n2903_n3924.n4 a_n2903_n3924.n2 0.358259
R22848 a_n2903_n3924.n48 a_n2903_n3924.n0 0.358259
R22849 a_n2903_n3924.n48 a_n2903_n3924.n47 0.358259
R22850 a_n2903_n3924.n47 a_n2903_n3924.n45 0.358259
R22851 a_n2903_n3924.n45 a_n2903_n3924.n43 0.358259
R22852 a_n2903_n3924.n43 a_n2903_n3924.n41 0.358259
R22853 a_n2903_n3924.n18 a_n2903_n3924.n12 0.270122
R22854 a_n2903_n3924.n13 a_n2903_n3924.n1 0.259948
R22855 a_n2903_n3924.n30 a_n2903_n3924.n29 0.235414
R22856 a_n2903_n3924.n2 a_n2903_n3924.n0 0.235414
R22857 minus.n36 minus.t23 436.949
R22858 minus.n6 minus.t11 436.949
R22859 minus.n54 minus.t18 415.966
R22860 minus.n53 minus.t13 415.966
R22861 minus.n29 minus.t20 415.966
R22862 minus.n47 minus.t10 415.966
R22863 minus.n46 minus.t5 415.966
R22864 minus.n32 minus.t14 415.966
R22865 minus.n41 minus.t9 415.966
R22866 minus.n39 minus.t22 415.966
R22867 minus.n35 minus.t7 415.966
R22868 minus.n7 minus.t15 415.966
R22869 minus.n5 minus.t8 415.966
R22870 minus.n13 minus.t12 415.966
R22871 minus.n14 minus.t21 415.966
R22872 minus.n18 minus.t16 415.966
R22873 minus.n19 minus.t19 415.966
R22874 minus.n1 minus.t6 415.966
R22875 minus.n25 minus.t17 415.966
R22876 minus.n26 minus.t24 415.966
R22877 minus.n60 minus.t1 243.255
R22878 minus.n59 minus.n57 224.169
R22879 minus.n59 minus.n58 223.454
R22880 minus.n38 minus.n37 161.3
R22881 minus.n39 minus.n34 161.3
R22882 minus.n40 minus.n33 161.3
R22883 minus.n42 minus.n41 161.3
R22884 minus.n43 minus.n32 161.3
R22885 minus.n45 minus.n44 161.3
R22886 minus.n46 minus.n31 161.3
R22887 minus.n47 minus.n30 161.3
R22888 minus.n49 minus.n48 161.3
R22889 minus.n50 minus.n29 161.3
R22890 minus.n52 minus.n51 161.3
R22891 minus.n53 minus.n28 161.3
R22892 minus.n55 minus.n54 161.3
R22893 minus.n27 minus.n26 161.3
R22894 minus.n25 minus.n0 161.3
R22895 minus.n24 minus.n23 161.3
R22896 minus.n22 minus.n1 161.3
R22897 minus.n21 minus.n20 161.3
R22898 minus.n19 minus.n2 161.3
R22899 minus.n18 minus.n17 161.3
R22900 minus.n16 minus.n3 161.3
R22901 minus.n15 minus.n14 161.3
R22902 minus.n13 minus.n4 161.3
R22903 minus.n12 minus.n11 161.3
R22904 minus.n10 minus.n5 161.3
R22905 minus.n9 minus.n8 161.3
R22906 minus.n37 minus.n36 70.4033
R22907 minus.n9 minus.n6 70.4033
R22908 minus.n54 minus.n53 48.2005
R22909 minus.n47 minus.n46 48.2005
R22910 minus.n41 minus.n32 48.2005
R22911 minus.n14 minus.n13 48.2005
R22912 minus.n19 minus.n18 48.2005
R22913 minus.n26 minus.n25 48.2005
R22914 minus.n48 minus.n29 47.4702
R22915 minus.n40 minus.n39 47.4702
R22916 minus.n12 minus.n5 47.4702
R22917 minus.n20 minus.n1 47.4702
R22918 minus.n56 minus.n55 30.0782
R22919 minus.n52 minus.n29 25.5611
R22920 minus.n39 minus.n38 25.5611
R22921 minus.n8 minus.n5 25.5611
R22922 minus.n24 minus.n1 25.5611
R22923 minus.n46 minus.n45 24.1005
R22924 minus.n45 minus.n32 24.1005
R22925 minus.n14 minus.n3 24.1005
R22926 minus.n18 minus.n3 24.1005
R22927 minus.n53 minus.n52 22.6399
R22928 minus.n38 minus.n35 22.6399
R22929 minus.n8 minus.n7 22.6399
R22930 minus.n25 minus.n24 22.6399
R22931 minus.n36 minus.n35 20.9576
R22932 minus.n7 minus.n6 20.9576
R22933 minus.n58 minus.t0 19.8005
R22934 minus.n58 minus.t4 19.8005
R22935 minus.n57 minus.t2 19.8005
R22936 minus.n57 minus.t3 19.8005
R22937 minus.n56 minus.n27 12.0062
R22938 minus minus.n61 11.3449
R22939 minus.n61 minus.n60 4.80222
R22940 minus.n61 minus.n56 0.972091
R22941 minus.n48 minus.n47 0.730803
R22942 minus.n41 minus.n40 0.730803
R22943 minus.n13 minus.n12 0.730803
R22944 minus.n20 minus.n19 0.730803
R22945 minus.n60 minus.n59 0.716017
R22946 minus.n55 minus.n28 0.189894
R22947 minus.n51 minus.n28 0.189894
R22948 minus.n51 minus.n50 0.189894
R22949 minus.n50 minus.n49 0.189894
R22950 minus.n49 minus.n30 0.189894
R22951 minus.n31 minus.n30 0.189894
R22952 minus.n44 minus.n31 0.189894
R22953 minus.n44 minus.n43 0.189894
R22954 minus.n43 minus.n42 0.189894
R22955 minus.n42 minus.n33 0.189894
R22956 minus.n34 minus.n33 0.189894
R22957 minus.n37 minus.n34 0.189894
R22958 minus.n10 minus.n9 0.189894
R22959 minus.n11 minus.n10 0.189894
R22960 minus.n11 minus.n4 0.189894
R22961 minus.n15 minus.n4 0.189894
R22962 minus.n16 minus.n15 0.189894
R22963 minus.n17 minus.n16 0.189894
R22964 minus.n17 minus.n2 0.189894
R22965 minus.n21 minus.n2 0.189894
R22966 minus.n22 minus.n21 0.189894
R22967 minus.n23 minus.n22 0.189894
R22968 minus.n23 minus.n0 0.189894
R22969 minus.n27 minus.n0 0.189894
R22970 diffpairibias.n0 diffpairibias.t18 436.822
R22971 diffpairibias.n21 diffpairibias.t19 435.479
R22972 diffpairibias.n20 diffpairibias.t16 435.479
R22973 diffpairibias.n19 diffpairibias.t17 435.479
R22974 diffpairibias.n18 diffpairibias.t21 435.479
R22975 diffpairibias.n0 diffpairibias.t22 435.479
R22976 diffpairibias.n1 diffpairibias.t20 435.479
R22977 diffpairibias.n2 diffpairibias.t23 435.479
R22978 diffpairibias.n10 diffpairibias.t0 377.536
R22979 diffpairibias.n10 diffpairibias.t8 376.193
R22980 diffpairibias.n11 diffpairibias.t10 376.193
R22981 diffpairibias.n12 diffpairibias.t6 376.193
R22982 diffpairibias.n13 diffpairibias.t2 376.193
R22983 diffpairibias.n14 diffpairibias.t12 376.193
R22984 diffpairibias.n15 diffpairibias.t4 376.193
R22985 diffpairibias.n16 diffpairibias.t14 376.193
R22986 diffpairibias.n3 diffpairibias.t1 113.368
R22987 diffpairibias.n3 diffpairibias.t9 112.698
R22988 diffpairibias.n4 diffpairibias.t11 112.698
R22989 diffpairibias.n5 diffpairibias.t7 112.698
R22990 diffpairibias.n6 diffpairibias.t3 112.698
R22991 diffpairibias.n7 diffpairibias.t13 112.698
R22992 diffpairibias.n8 diffpairibias.t5 112.698
R22993 diffpairibias.n9 diffpairibias.t15 112.698
R22994 diffpairibias.n17 diffpairibias.n16 4.77242
R22995 diffpairibias.n17 diffpairibias.n9 4.30807
R22996 diffpairibias.n18 diffpairibias.n17 4.13945
R22997 diffpairibias.n16 diffpairibias.n15 1.34352
R22998 diffpairibias.n15 diffpairibias.n14 1.34352
R22999 diffpairibias.n14 diffpairibias.n13 1.34352
R23000 diffpairibias.n13 diffpairibias.n12 1.34352
R23001 diffpairibias.n12 diffpairibias.n11 1.34352
R23002 diffpairibias.n11 diffpairibias.n10 1.34352
R23003 diffpairibias.n2 diffpairibias.n1 1.34352
R23004 diffpairibias.n1 diffpairibias.n0 1.34352
R23005 diffpairibias.n19 diffpairibias.n18 1.34352
R23006 diffpairibias.n20 diffpairibias.n19 1.34352
R23007 diffpairibias.n21 diffpairibias.n20 1.34352
R23008 diffpairibias.n22 diffpairibias.n21 0.862419
R23009 diffpairibias diffpairibias.n22 0.684875
R23010 diffpairibias.n9 diffpairibias.n8 0.672012
R23011 diffpairibias.n8 diffpairibias.n7 0.672012
R23012 diffpairibias.n7 diffpairibias.n6 0.672012
R23013 diffpairibias.n6 diffpairibias.n5 0.672012
R23014 diffpairibias.n5 diffpairibias.n4 0.672012
R23015 diffpairibias.n4 diffpairibias.n3 0.672012
R23016 diffpairibias.n22 diffpairibias.n2 0.190907
C0 commonsourceibias diffpairibias 0.06482f
C1 CSoutput commonsourceibias 41.846302f
C2 minus plus 8.457049f
C3 minus commonsourceibias 0.31863f
C4 plus commonsourceibias 0.272687f
C5 output outputibias 2.34152f
C6 vdd output 7.23429f
C7 CSoutput output 6.13881f
C8 CSoutput outputibias 0.032386f
C9 vdd CSoutput 0.14174p
C10 minus diffpairibias 2.77e-19
C11 commonsourceibias output 0.006808f
C12 vdd plus 0.090721f
C13 CSoutput minus 2.59933f
C14 plus diffpairibias 2.54e-19
C15 commonsourceibias outputibias 0.003832f
C16 vdd commonsourceibias 0.004218f
C17 CSoutput plus 0.82208f
C18 diffpairibias gnd 48.97994f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.144426p
C22 plus gnd 30.2452f
C23 minus gnd 25.205141f
C24 CSoutput gnd 0.105777p
C25 vdd gnd 0.472827p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 minus.n0 gnd 0.032928f
C74 minus.t6 gnd 0.332672f
C75 minus.n1 gnd 0.153805f
C76 minus.n2 gnd 0.032928f
C77 minus.n3 gnd 0.007472f
C78 minus.n4 gnd 0.032928f
C79 minus.t8 gnd 0.332672f
C80 minus.n5 gnd 0.153805f
C81 minus.t11 gnd 0.339894f
C82 minus.n6 gnd 0.143384f
C83 minus.t15 gnd 0.332672f
C84 minus.n7 gnd 0.1535f
C85 minus.n8 gnd 0.007472f
C86 minus.n9 gnd 0.108074f
C87 minus.n10 gnd 0.032928f
C88 minus.n11 gnd 0.032928f
C89 minus.n12 gnd 0.007472f
C90 minus.t12 gnd 0.332672f
C91 minus.n13 gnd 0.150455f
C92 minus.t21 gnd 0.332672f
C93 minus.n14 gnd 0.153703f
C94 minus.n15 gnd 0.032928f
C95 minus.n16 gnd 0.032928f
C96 minus.n17 gnd 0.032928f
C97 minus.t16 gnd 0.332672f
C98 minus.n18 gnd 0.153703f
C99 minus.t19 gnd 0.332672f
C100 minus.n19 gnd 0.150455f
C101 minus.n20 gnd 0.007472f
C102 minus.n21 gnd 0.032928f
C103 minus.n22 gnd 0.032928f
C104 minus.n23 gnd 0.032928f
C105 minus.n24 gnd 0.007472f
C106 minus.t17 gnd 0.332672f
C107 minus.n25 gnd 0.1535f
C108 minus.t24 gnd 0.332672f
C109 minus.n26 gnd 0.150353f
C110 minus.n27 gnd 0.374572f
C111 minus.n28 gnd 0.032928f
C112 minus.t18 gnd 0.332672f
C113 minus.t13 gnd 0.332672f
C114 minus.t20 gnd 0.332672f
C115 minus.n29 gnd 0.153805f
C116 minus.n30 gnd 0.032928f
C117 minus.t10 gnd 0.332672f
C118 minus.t5 gnd 0.332672f
C119 minus.n31 gnd 0.032928f
C120 minus.t14 gnd 0.332672f
C121 minus.n32 gnd 0.153703f
C122 minus.n33 gnd 0.032928f
C123 minus.t9 gnd 0.332672f
C124 minus.t22 gnd 0.332672f
C125 minus.n34 gnd 0.032928f
C126 minus.t7 gnd 0.332672f
C127 minus.n35 gnd 0.1535f
C128 minus.t23 gnd 0.339894f
C129 minus.n36 gnd 0.143384f
C130 minus.n37 gnd 0.108074f
C131 minus.n38 gnd 0.007472f
C132 minus.n39 gnd 0.153805f
C133 minus.n40 gnd 0.007472f
C134 minus.n41 gnd 0.150455f
C135 minus.n42 gnd 0.032928f
C136 minus.n43 gnd 0.032928f
C137 minus.n44 gnd 0.032928f
C138 minus.n45 gnd 0.007472f
C139 minus.n46 gnd 0.153703f
C140 minus.n47 gnd 0.150455f
C141 minus.n48 gnd 0.007472f
C142 minus.n49 gnd 0.032928f
C143 minus.n50 gnd 0.032928f
C144 minus.n51 gnd 0.032928f
C145 minus.n52 gnd 0.007472f
C146 minus.n53 gnd 0.1535f
C147 minus.n54 gnd 0.150353f
C148 minus.n55 gnd 0.945954f
C149 minus.n56 gnd 1.44297f
C150 minus.t2 gnd 0.010151f
C151 minus.t3 gnd 0.010151f
C152 minus.n57 gnd 0.033378f
C153 minus.t0 gnd 0.010151f
C154 minus.t4 gnd 0.010151f
C155 minus.n58 gnd 0.032921f
C156 minus.n59 gnd 0.280965f
C157 minus.t1 gnd 0.056498f
C158 minus.n60 gnd 0.15332f
C159 minus.n61 gnd 1.93528f
C160 a_n2903_n3924.t15 gnd 0.102414f
C161 a_n2903_n3924.t12 gnd 1.06441f
C162 a_n2903_n3924.n0 gnd 0.361252f
C163 a_n2903_n3924.t30 gnd 1.32447f
C164 a_n2903_n3924.n1 gnd 1.52483f
C165 a_n2903_n3924.t7 gnd 1.06441f
C166 a_n2903_n3924.n2 gnd 0.361252f
C167 a_n2903_n3924.t39 gnd 0.102414f
C168 a_n2903_n3924.t0 gnd 0.102414f
C169 a_n2903_n3924.n3 gnd 0.836435f
C170 a_n2903_n3924.n4 gnd 0.33923f
C171 a_n2903_n3924.t36 gnd 0.102414f
C172 a_n2903_n3924.t9 gnd 0.102414f
C173 a_n2903_n3924.n5 gnd 0.836435f
C174 a_n2903_n3924.n6 gnd 0.33923f
C175 a_n2903_n3924.t43 gnd 0.102414f
C176 a_n2903_n3924.t34 gnd 0.102414f
C177 a_n2903_n3924.n7 gnd 0.836435f
C178 a_n2903_n3924.n8 gnd 0.33923f
C179 a_n2903_n3924.t33 gnd 0.102414f
C180 a_n2903_n3924.t8 gnd 0.102414f
C181 a_n2903_n3924.n9 gnd 0.836435f
C182 a_n2903_n3924.n10 gnd 0.33923f
C183 a_n2903_n3924.t45 gnd 1.06441f
C184 a_n2903_n3924.n11 gnd 0.918548f
C185 a_n2903_n3924.t47 gnd 1.32439f
C186 a_n2903_n3924.t31 gnd 1.32251f
C187 a_n2903_n3924.n12 gnd 1.32305f
C188 a_n2903_n3924.t35 gnd 1.32251f
C189 a_n2903_n3924.n13 gnd 0.715276f
C190 a_n2903_n3924.t38 gnd 1.32251f
C191 a_n2903_n3924.n14 gnd 0.931464f
C192 a_n2903_n3924.t37 gnd 1.32251f
C193 a_n2903_n3924.n15 gnd 0.931464f
C194 a_n2903_n3924.t1 gnd 1.32251f
C195 a_n2903_n3924.n16 gnd 0.931464f
C196 a_n2903_n3924.t41 gnd 1.32251f
C197 a_n2903_n3924.n17 gnd 0.790007f
C198 a_n2903_n3924.n18 gnd 0.50344f
C199 a_n2903_n3924.n19 gnd 0.956044f
C200 a_n2903_n3924.t10 gnd 1.06441f
C201 a_n2903_n3924.n20 gnd 0.583868f
C202 a_n2903_n3924.t14 gnd 0.102414f
C203 a_n2903_n3924.t27 gnd 0.102414f
C204 a_n2903_n3924.n21 gnd 0.836434f
C205 a_n2903_n3924.n22 gnd 0.339231f
C206 a_n2903_n3924.t17 gnd 0.102414f
C207 a_n2903_n3924.t21 gnd 0.102414f
C208 a_n2903_n3924.n23 gnd 0.836434f
C209 a_n2903_n3924.n24 gnd 0.339231f
C210 a_n2903_n3924.t13 gnd 0.102414f
C211 a_n2903_n3924.t18 gnd 0.102414f
C212 a_n2903_n3924.n25 gnd 0.836434f
C213 a_n2903_n3924.n26 gnd 0.339231f
C214 a_n2903_n3924.t25 gnd 0.102414f
C215 a_n2903_n3924.t20 gnd 0.102414f
C216 a_n2903_n3924.n27 gnd 0.836434f
C217 a_n2903_n3924.n28 gnd 0.339231f
C218 a_n2903_n3924.t22 gnd 1.06441f
C219 a_n2903_n3924.n29 gnd 0.361256f
C220 a_n2903_n3924.t2 gnd 1.06441f
C221 a_n2903_n3924.n30 gnd 0.361256f
C222 a_n2903_n3924.t44 gnd 0.102414f
C223 a_n2903_n3924.t3 gnd 0.102414f
C224 a_n2903_n3924.n31 gnd 0.836434f
C225 a_n2903_n3924.n32 gnd 0.339231f
C226 a_n2903_n3924.t42 gnd 0.102414f
C227 a_n2903_n3924.t4 gnd 0.102414f
C228 a_n2903_n3924.n33 gnd 0.836434f
C229 a_n2903_n3924.n34 gnd 0.339231f
C230 a_n2903_n3924.t6 gnd 0.102414f
C231 a_n2903_n3924.t46 gnd 0.102414f
C232 a_n2903_n3924.n35 gnd 0.836434f
C233 a_n2903_n3924.n36 gnd 0.339231f
C234 a_n2903_n3924.t32 gnd 0.102414f
C235 a_n2903_n3924.t5 gnd 0.102414f
C236 a_n2903_n3924.n37 gnd 0.836434f
C237 a_n2903_n3924.n38 gnd 0.339231f
C238 a_n2903_n3924.t40 gnd 1.06441f
C239 a_n2903_n3924.n39 gnd 0.583868f
C240 a_n2903_n3924.n40 gnd 0.956044f
C241 a_n2903_n3924.t19 gnd 1.06441f
C242 a_n2903_n3924.n41 gnd 0.918552f
C243 a_n2903_n3924.t16 gnd 0.102414f
C244 a_n2903_n3924.t26 gnd 0.102414f
C245 a_n2903_n3924.n42 gnd 0.836435f
C246 a_n2903_n3924.n43 gnd 0.33923f
C247 a_n2903_n3924.t28 gnd 0.102414f
C248 a_n2903_n3924.t24 gnd 0.102414f
C249 a_n2903_n3924.n44 gnd 0.836435f
C250 a_n2903_n3924.n45 gnd 0.33923f
C251 a_n2903_n3924.t11 gnd 0.102414f
C252 a_n2903_n3924.t23 gnd 0.102414f
C253 a_n2903_n3924.n46 gnd 0.836435f
C254 a_n2903_n3924.n47 gnd 0.33923f
C255 a_n2903_n3924.n48 gnd 0.339229f
C256 a_n2903_n3924.n49 gnd 0.836436f
C257 a_n2903_n3924.t29 gnd 0.102414f
C258 plus.n0 gnd 0.023788f
C259 plus.t24 gnd 0.240322f
C260 plus.t20 gnd 0.240322f
C261 plus.t7 gnd 0.240322f
C262 plus.n1 gnd 0.111109f
C263 plus.n2 gnd 0.023788f
C264 plus.t17 gnd 0.240322f
C265 plus.n3 gnd 0.023788f
C266 plus.t13 gnd 0.240322f
C267 plus.t21 gnd 0.240322f
C268 plus.n4 gnd 0.111035f
C269 plus.n5 gnd 0.023788f
C270 plus.t16 gnd 0.240322f
C271 plus.n6 gnd 0.023788f
C272 plus.t9 gnd 0.240322f
C273 plus.t14 gnd 0.240322f
C274 plus.n7 gnd 0.110889f
C275 plus.t12 gnd 0.24554f
C276 plus.n8 gnd 0.103581f
C277 plus.n9 gnd 0.078073f
C278 plus.n10 gnd 0.005398f
C279 plus.n11 gnd 0.111109f
C280 plus.n12 gnd 0.005398f
C281 plus.n13 gnd 0.108689f
C282 plus.n14 gnd 0.023788f
C283 plus.n15 gnd 0.023788f
C284 plus.n16 gnd 0.023788f
C285 plus.n17 gnd 0.005398f
C286 plus.n18 gnd 0.111035f
C287 plus.n19 gnd 0.108689f
C288 plus.n20 gnd 0.005398f
C289 plus.n21 gnd 0.023788f
C290 plus.n22 gnd 0.023788f
C291 plus.n23 gnd 0.023788f
C292 plus.n24 gnd 0.005398f
C293 plus.n25 gnd 0.110889f
C294 plus.n26 gnd 0.108615f
C295 plus.n27 gnd 0.264453f
C296 plus.n28 gnd 0.023788f
C297 plus.t18 gnd 0.240322f
C298 plus.n29 gnd 0.111109f
C299 plus.n30 gnd 0.023788f
C300 plus.n31 gnd 0.005398f
C301 plus.t6 gnd 0.240322f
C302 plus.n32 gnd 0.023788f
C303 plus.t19 gnd 0.240322f
C304 plus.n33 gnd 0.111109f
C305 plus.t22 gnd 0.24554f
C306 plus.n34 gnd 0.103581f
C307 plus.t5 gnd 0.240322f
C308 plus.n35 gnd 0.110889f
C309 plus.n36 gnd 0.005398f
C310 plus.n37 gnd 0.078073f
C311 plus.n38 gnd 0.023788f
C312 plus.n39 gnd 0.023788f
C313 plus.n40 gnd 0.005398f
C314 plus.t23 gnd 0.240322f
C315 plus.n41 gnd 0.108689f
C316 plus.t11 gnd 0.240322f
C317 plus.n42 gnd 0.111035f
C318 plus.n43 gnd 0.023788f
C319 plus.n44 gnd 0.023788f
C320 plus.n45 gnd 0.023788f
C321 plus.n46 gnd 0.111035f
C322 plus.t10 gnd 0.240322f
C323 plus.n47 gnd 0.108689f
C324 plus.n48 gnd 0.005398f
C325 plus.n49 gnd 0.023788f
C326 plus.n50 gnd 0.023788f
C327 plus.n51 gnd 0.023788f
C328 plus.n52 gnd 0.005398f
C329 plus.t8 gnd 0.240322f
C330 plus.n53 gnd 0.110889f
C331 plus.t15 gnd 0.240322f
C332 plus.n54 gnd 0.108615f
C333 plus.n55 gnd 0.673801f
C334 plus.n56 gnd 1.03302f
C335 plus.t0 gnd 0.041064f
C336 plus.t3 gnd 0.007333f
C337 plus.t2 gnd 0.007333f
C338 plus.n57 gnd 0.023782f
C339 plus.n58 gnd 0.184623f
C340 plus.t4 gnd 0.007333f
C341 plus.t1 gnd 0.007333f
C342 plus.n59 gnd 0.023782f
C343 plus.n60 gnd 0.138582f
C344 plus.n61 gnd 2.35935f
C345 a_n2318_8322.t24 gnd 39.618103f
C346 a_n2318_8322.t26 gnd 27.7211f
C347 a_n2318_8322.t27 gnd 19.739399f
C348 a_n2318_8322.t25 gnd 39.618103f
C349 a_n2318_8322.t4 gnd 0.09582f
C350 a_n2318_8322.t14 gnd 0.89721f
C351 a_n2318_8322.t2 gnd 0.09582f
C352 a_n2318_8322.t1 gnd 0.09582f
C353 a_n2318_8322.n0 gnd 0.674956f
C354 a_n2318_8322.n1 gnd 0.754164f
C355 a_n2318_8322.t11 gnd 0.09582f
C356 a_n2318_8322.t6 gnd 0.09582f
C357 a_n2318_8322.n2 gnd 0.674956f
C358 a_n2318_8322.n3 gnd 0.383181f
C359 a_n2318_8322.t9 gnd 0.09582f
C360 a_n2318_8322.t8 gnd 0.09582f
C361 a_n2318_8322.n4 gnd 0.674956f
C362 a_n2318_8322.n5 gnd 0.383181f
C363 a_n2318_8322.t0 gnd 0.895423f
C364 a_n2318_8322.n6 gnd 1.5519f
C365 a_n2318_8322.t19 gnd 0.89721f
C366 a_n2318_8322.t23 gnd 0.09582f
C367 a_n2318_8322.t22 gnd 0.09582f
C368 a_n2318_8322.n7 gnd 0.674956f
C369 a_n2318_8322.n8 gnd 0.754164f
C370 a_n2318_8322.t17 gnd 0.895423f
C371 a_n2318_8322.n9 gnd 0.379506f
C372 a_n2318_8322.t20 gnd 0.895423f
C373 a_n2318_8322.n10 gnd 0.379506f
C374 a_n2318_8322.t18 gnd 0.09582f
C375 a_n2318_8322.t16 gnd 0.09582f
C376 a_n2318_8322.n11 gnd 0.674956f
C377 a_n2318_8322.n12 gnd 0.383181f
C378 a_n2318_8322.t21 gnd 0.895423f
C379 a_n2318_8322.n13 gnd 1.07467f
C380 a_n2318_8322.n14 gnd 1.82686f
C381 a_n2318_8322.n15 gnd 3.12946f
C382 a_n2318_8322.t3 gnd 0.895423f
C383 a_n2318_8322.n16 gnd 0.881475f
C384 a_n2318_8322.t12 gnd 0.09582f
C385 a_n2318_8322.t5 gnd 0.09582f
C386 a_n2318_8322.n17 gnd 0.674956f
C387 a_n2318_8322.n18 gnd 0.383181f
C388 a_n2318_8322.t13 gnd 0.897207f
C389 a_n2318_8322.t10 gnd 0.09582f
C390 a_n2318_8322.t7 gnd 0.09582f
C391 a_n2318_8322.n19 gnd 0.674956f
C392 a_n2318_8322.n20 gnd 0.754166f
C393 a_n2318_8322.n21 gnd 0.383179f
C394 a_n2318_8322.n22 gnd 0.674958f
C395 a_n2318_8322.t15 gnd 0.09582f
C396 output.t8 gnd 0.464308f
C397 output.t14 gnd 0.044422f
C398 output.t18 gnd 0.044422f
C399 output.n0 gnd 0.364624f
C400 output.n1 gnd 0.614102f
C401 output.t5 gnd 0.044422f
C402 output.t10 gnd 0.044422f
C403 output.n2 gnd 0.364624f
C404 output.n3 gnd 0.350265f
C405 output.t11 gnd 0.044422f
C406 output.t16 gnd 0.044422f
C407 output.n4 gnd 0.364624f
C408 output.n5 gnd 0.350265f
C409 output.t4 gnd 0.044422f
C410 output.t12 gnd 0.044422f
C411 output.n6 gnd 0.364624f
C412 output.n7 gnd 0.350265f
C413 output.t15 gnd 0.044422f
C414 output.t13 gnd 0.044422f
C415 output.n8 gnd 0.364624f
C416 output.n9 gnd 0.350265f
C417 output.t19 gnd 0.044422f
C418 output.t6 gnd 0.044422f
C419 output.n10 gnd 0.364624f
C420 output.n11 gnd 0.350265f
C421 output.t7 gnd 0.044422f
C422 output.t17 gnd 0.044422f
C423 output.n12 gnd 0.364624f
C424 output.n13 gnd 0.350265f
C425 output.t9 gnd 0.462979f
C426 output.n14 gnd 0.28994f
C427 output.n15 gnd 0.015803f
C428 output.n16 gnd 0.011243f
C429 output.n17 gnd 0.006041f
C430 output.n18 gnd 0.01428f
C431 output.n19 gnd 0.006397f
C432 output.n20 gnd 0.011243f
C433 output.n21 gnd 0.006041f
C434 output.n22 gnd 0.01428f
C435 output.n23 gnd 0.006397f
C436 output.n24 gnd 0.048111f
C437 output.t2 gnd 0.023274f
C438 output.n25 gnd 0.01071f
C439 output.n26 gnd 0.008435f
C440 output.n27 gnd 0.006041f
C441 output.n28 gnd 0.267512f
C442 output.n29 gnd 0.011243f
C443 output.n30 gnd 0.006041f
C444 output.n31 gnd 0.006397f
C445 output.n32 gnd 0.01428f
C446 output.n33 gnd 0.01428f
C447 output.n34 gnd 0.006397f
C448 output.n35 gnd 0.006041f
C449 output.n36 gnd 0.011243f
C450 output.n37 gnd 0.011243f
C451 output.n38 gnd 0.006041f
C452 output.n39 gnd 0.006397f
C453 output.n40 gnd 0.01428f
C454 output.n41 gnd 0.030913f
C455 output.n42 gnd 0.006397f
C456 output.n43 gnd 0.006041f
C457 output.n44 gnd 0.025987f
C458 output.n45 gnd 0.097665f
C459 output.n46 gnd 0.015803f
C460 output.n47 gnd 0.011243f
C461 output.n48 gnd 0.006041f
C462 output.n49 gnd 0.01428f
C463 output.n50 gnd 0.006397f
C464 output.n51 gnd 0.011243f
C465 output.n52 gnd 0.006041f
C466 output.n53 gnd 0.01428f
C467 output.n54 gnd 0.006397f
C468 output.n55 gnd 0.048111f
C469 output.t1 gnd 0.023274f
C470 output.n56 gnd 0.01071f
C471 output.n57 gnd 0.008435f
C472 output.n58 gnd 0.006041f
C473 output.n59 gnd 0.267512f
C474 output.n60 gnd 0.011243f
C475 output.n61 gnd 0.006041f
C476 output.n62 gnd 0.006397f
C477 output.n63 gnd 0.01428f
C478 output.n64 gnd 0.01428f
C479 output.n65 gnd 0.006397f
C480 output.n66 gnd 0.006041f
C481 output.n67 gnd 0.011243f
C482 output.n68 gnd 0.011243f
C483 output.n69 gnd 0.006041f
C484 output.n70 gnd 0.006397f
C485 output.n71 gnd 0.01428f
C486 output.n72 gnd 0.030913f
C487 output.n73 gnd 0.006397f
C488 output.n74 gnd 0.006041f
C489 output.n75 gnd 0.025987f
C490 output.n76 gnd 0.09306f
C491 output.n77 gnd 1.65264f
C492 output.n78 gnd 0.015803f
C493 output.n79 gnd 0.011243f
C494 output.n80 gnd 0.006041f
C495 output.n81 gnd 0.01428f
C496 output.n82 gnd 0.006397f
C497 output.n83 gnd 0.011243f
C498 output.n84 gnd 0.006041f
C499 output.n85 gnd 0.01428f
C500 output.n86 gnd 0.006397f
C501 output.n87 gnd 0.048111f
C502 output.t3 gnd 0.023274f
C503 output.n88 gnd 0.01071f
C504 output.n89 gnd 0.008435f
C505 output.n90 gnd 0.006041f
C506 output.n91 gnd 0.267512f
C507 output.n92 gnd 0.011243f
C508 output.n93 gnd 0.006041f
C509 output.n94 gnd 0.006397f
C510 output.n95 gnd 0.01428f
C511 output.n96 gnd 0.01428f
C512 output.n97 gnd 0.006397f
C513 output.n98 gnd 0.006041f
C514 output.n99 gnd 0.011243f
C515 output.n100 gnd 0.011243f
C516 output.n101 gnd 0.006041f
C517 output.n102 gnd 0.006397f
C518 output.n103 gnd 0.01428f
C519 output.n104 gnd 0.030913f
C520 output.n105 gnd 0.006397f
C521 output.n106 gnd 0.006041f
C522 output.n107 gnd 0.025987f
C523 output.n108 gnd 0.09306f
C524 output.n109 gnd 0.713089f
C525 output.n110 gnd 0.015803f
C526 output.n111 gnd 0.011243f
C527 output.n112 gnd 0.006041f
C528 output.n113 gnd 0.01428f
C529 output.n114 gnd 0.006397f
C530 output.n115 gnd 0.011243f
C531 output.n116 gnd 0.006041f
C532 output.n117 gnd 0.01428f
C533 output.n118 gnd 0.006397f
C534 output.n119 gnd 0.048111f
C535 output.t0 gnd 0.023274f
C536 output.n120 gnd 0.01071f
C537 output.n121 gnd 0.008435f
C538 output.n122 gnd 0.006041f
C539 output.n123 gnd 0.267512f
C540 output.n124 gnd 0.011243f
C541 output.n125 gnd 0.006041f
C542 output.n126 gnd 0.006397f
C543 output.n127 gnd 0.01428f
C544 output.n128 gnd 0.01428f
C545 output.n129 gnd 0.006397f
C546 output.n130 gnd 0.006041f
C547 output.n131 gnd 0.011243f
C548 output.n132 gnd 0.011243f
C549 output.n133 gnd 0.006041f
C550 output.n134 gnd 0.006397f
C551 output.n135 gnd 0.01428f
C552 output.n136 gnd 0.030913f
C553 output.n137 gnd 0.006397f
C554 output.n138 gnd 0.006041f
C555 output.n139 gnd 0.025987f
C556 output.n140 gnd 0.09306f
C557 output.n141 gnd 1.67353f
C558 outputibias.t10 gnd 0.11477f
C559 outputibias.t9 gnd 0.115567f
C560 outputibias.n0 gnd 0.130108f
C561 outputibias.n1 gnd 0.001372f
C562 outputibias.n2 gnd 9.76e-19
C563 outputibias.n3 gnd 5.24e-19
C564 outputibias.n4 gnd 0.001239f
C565 outputibias.n5 gnd 5.55e-19
C566 outputibias.n6 gnd 9.76e-19
C567 outputibias.n7 gnd 5.24e-19
C568 outputibias.n8 gnd 0.001239f
C569 outputibias.n9 gnd 5.55e-19
C570 outputibias.n10 gnd 0.004176f
C571 outputibias.t5 gnd 0.00202f
C572 outputibias.n11 gnd 9.3e-19
C573 outputibias.n12 gnd 7.32e-19
C574 outputibias.n13 gnd 5.24e-19
C575 outputibias.n14 gnd 0.02322f
C576 outputibias.n15 gnd 9.76e-19
C577 outputibias.n16 gnd 5.24e-19
C578 outputibias.n17 gnd 5.55e-19
C579 outputibias.n18 gnd 0.001239f
C580 outputibias.n19 gnd 0.001239f
C581 outputibias.n20 gnd 5.55e-19
C582 outputibias.n21 gnd 5.24e-19
C583 outputibias.n22 gnd 9.76e-19
C584 outputibias.n23 gnd 9.76e-19
C585 outputibias.n24 gnd 5.24e-19
C586 outputibias.n25 gnd 5.55e-19
C587 outputibias.n26 gnd 0.001239f
C588 outputibias.n27 gnd 0.002683f
C589 outputibias.n28 gnd 5.55e-19
C590 outputibias.n29 gnd 5.24e-19
C591 outputibias.n30 gnd 0.002256f
C592 outputibias.n31 gnd 0.005781f
C593 outputibias.n32 gnd 0.001372f
C594 outputibias.n33 gnd 9.76e-19
C595 outputibias.n34 gnd 5.24e-19
C596 outputibias.n35 gnd 0.001239f
C597 outputibias.n36 gnd 5.55e-19
C598 outputibias.n37 gnd 9.76e-19
C599 outputibias.n38 gnd 5.24e-19
C600 outputibias.n39 gnd 0.001239f
C601 outputibias.n40 gnd 5.55e-19
C602 outputibias.n41 gnd 0.004176f
C603 outputibias.t7 gnd 0.00202f
C604 outputibias.n42 gnd 9.3e-19
C605 outputibias.n43 gnd 7.32e-19
C606 outputibias.n44 gnd 5.24e-19
C607 outputibias.n45 gnd 0.02322f
C608 outputibias.n46 gnd 9.76e-19
C609 outputibias.n47 gnd 5.24e-19
C610 outputibias.n48 gnd 5.55e-19
C611 outputibias.n49 gnd 0.001239f
C612 outputibias.n50 gnd 0.001239f
C613 outputibias.n51 gnd 5.55e-19
C614 outputibias.n52 gnd 5.24e-19
C615 outputibias.n53 gnd 9.76e-19
C616 outputibias.n54 gnd 9.76e-19
C617 outputibias.n55 gnd 5.24e-19
C618 outputibias.n56 gnd 5.55e-19
C619 outputibias.n57 gnd 0.001239f
C620 outputibias.n58 gnd 0.002683f
C621 outputibias.n59 gnd 5.55e-19
C622 outputibias.n60 gnd 5.24e-19
C623 outputibias.n61 gnd 0.002256f
C624 outputibias.n62 gnd 0.005197f
C625 outputibias.n63 gnd 0.121892f
C626 outputibias.n64 gnd 0.001372f
C627 outputibias.n65 gnd 9.76e-19
C628 outputibias.n66 gnd 5.24e-19
C629 outputibias.n67 gnd 0.001239f
C630 outputibias.n68 gnd 5.55e-19
C631 outputibias.n69 gnd 9.76e-19
C632 outputibias.n70 gnd 5.24e-19
C633 outputibias.n71 gnd 0.001239f
C634 outputibias.n72 gnd 5.55e-19
C635 outputibias.n73 gnd 0.004176f
C636 outputibias.t1 gnd 0.00202f
C637 outputibias.n74 gnd 9.3e-19
C638 outputibias.n75 gnd 7.32e-19
C639 outputibias.n76 gnd 5.24e-19
C640 outputibias.n77 gnd 0.02322f
C641 outputibias.n78 gnd 9.76e-19
C642 outputibias.n79 gnd 5.24e-19
C643 outputibias.n80 gnd 5.55e-19
C644 outputibias.n81 gnd 0.001239f
C645 outputibias.n82 gnd 0.001239f
C646 outputibias.n83 gnd 5.55e-19
C647 outputibias.n84 gnd 5.24e-19
C648 outputibias.n85 gnd 9.76e-19
C649 outputibias.n86 gnd 9.76e-19
C650 outputibias.n87 gnd 5.24e-19
C651 outputibias.n88 gnd 5.55e-19
C652 outputibias.n89 gnd 0.001239f
C653 outputibias.n90 gnd 0.002683f
C654 outputibias.n91 gnd 5.55e-19
C655 outputibias.n92 gnd 5.24e-19
C656 outputibias.n93 gnd 0.002256f
C657 outputibias.n94 gnd 0.005197f
C658 outputibias.n95 gnd 0.064513f
C659 outputibias.n96 gnd 0.001372f
C660 outputibias.n97 gnd 9.76e-19
C661 outputibias.n98 gnd 5.24e-19
C662 outputibias.n99 gnd 0.001239f
C663 outputibias.n100 gnd 5.55e-19
C664 outputibias.n101 gnd 9.76e-19
C665 outputibias.n102 gnd 5.24e-19
C666 outputibias.n103 gnd 0.001239f
C667 outputibias.n104 gnd 5.55e-19
C668 outputibias.n105 gnd 0.004176f
C669 outputibias.t3 gnd 0.00202f
C670 outputibias.n106 gnd 9.3e-19
C671 outputibias.n107 gnd 7.32e-19
C672 outputibias.n108 gnd 5.24e-19
C673 outputibias.n109 gnd 0.02322f
C674 outputibias.n110 gnd 9.76e-19
C675 outputibias.n111 gnd 5.24e-19
C676 outputibias.n112 gnd 5.55e-19
C677 outputibias.n113 gnd 0.001239f
C678 outputibias.n114 gnd 0.001239f
C679 outputibias.n115 gnd 5.55e-19
C680 outputibias.n116 gnd 5.24e-19
C681 outputibias.n117 gnd 9.76e-19
C682 outputibias.n118 gnd 9.76e-19
C683 outputibias.n119 gnd 5.24e-19
C684 outputibias.n120 gnd 5.55e-19
C685 outputibias.n121 gnd 0.001239f
C686 outputibias.n122 gnd 0.002683f
C687 outputibias.n123 gnd 5.55e-19
C688 outputibias.n124 gnd 5.24e-19
C689 outputibias.n125 gnd 0.002256f
C690 outputibias.n126 gnd 0.005197f
C691 outputibias.n127 gnd 0.084814f
C692 outputibias.t2 gnd 0.108319f
C693 outputibias.t0 gnd 0.108319f
C694 outputibias.t6 gnd 0.108319f
C695 outputibias.t4 gnd 0.109238f
C696 outputibias.n128 gnd 0.134674f
C697 outputibias.n129 gnd 0.07244f
C698 outputibias.n130 gnd 0.079818f
C699 outputibias.n131 gnd 0.164901f
C700 outputibias.t11 gnd 0.11477f
C701 outputibias.n132 gnd 0.067481f
C702 outputibias.t8 gnd 0.11477f
C703 outputibias.n133 gnd 0.065115f
C704 outputibias.n134 gnd 0.029159f
C705 a_n2140_13878.t11 gnd 0.186452f
C706 a_n2140_13878.t10 gnd 0.186452f
C707 a_n2140_13878.t5 gnd 0.186452f
C708 a_n2140_13878.n0 gnd 1.46971f
C709 a_n2140_13878.t2 gnd 0.186452f
C710 a_n2140_13878.t4 gnd 0.186452f
C711 a_n2140_13878.n1 gnd 1.46815f
C712 a_n2140_13878.n2 gnd 2.05145f
C713 a_n2140_13878.t12 gnd 0.186452f
C714 a_n2140_13878.t3 gnd 0.186452f
C715 a_n2140_13878.n3 gnd 1.46815f
C716 a_n2140_13878.n4 gnd 1.00065f
C717 a_n2140_13878.t9 gnd 0.186452f
C718 a_n2140_13878.t1 gnd 0.186452f
C719 a_n2140_13878.n5 gnd 1.46815f
C720 a_n2140_13878.n6 gnd 4.05307f
C721 a_n2140_13878.t17 gnd 1.74584f
C722 a_n2140_13878.t20 gnd 0.186452f
C723 a_n2140_13878.t21 gnd 0.186452f
C724 a_n2140_13878.n7 gnd 1.31337f
C725 a_n2140_13878.n8 gnd 1.4675f
C726 a_n2140_13878.t16 gnd 1.74237f
C727 a_n2140_13878.n9 gnd 0.738464f
C728 a_n2140_13878.t19 gnd 1.74237f
C729 a_n2140_13878.n10 gnd 0.738464f
C730 a_n2140_13878.t22 gnd 0.186452f
C731 a_n2140_13878.t23 gnd 0.186452f
C732 a_n2140_13878.n11 gnd 1.31337f
C733 a_n2140_13878.n12 gnd 0.745616f
C734 a_n2140_13878.t18 gnd 1.74237f
C735 a_n2140_13878.n13 gnd 2.09116f
C736 a_n2140_13878.n14 gnd 2.85337f
C737 a_n2140_13878.t6 gnd 0.186452f
C738 a_n2140_13878.t7 gnd 0.186452f
C739 a_n2140_13878.n15 gnd 1.46815f
C740 a_n2140_13878.n16 gnd 2.01216f
C741 a_n2140_13878.t13 gnd 0.186452f
C742 a_n2140_13878.t14 gnd 0.186452f
C743 a_n2140_13878.n17 gnd 1.46815f
C744 a_n2140_13878.n18 gnd 0.650499f
C745 a_n2140_13878.t0 gnd 0.186452f
C746 a_n2140_13878.t8 gnd 0.186452f
C747 a_n2140_13878.n19 gnd 1.46815f
C748 a_n2140_13878.n20 gnd 1.31969f
C749 a_n2140_13878.n21 gnd 1.47058f
C750 a_n2140_13878.t15 gnd 0.186452f
C751 a_n2318_13878.n0 gnd 0.217886f
C752 a_n2318_13878.n1 gnd 0.753715f
C753 a_n2318_13878.n2 gnd 0.217886f
C754 a_n2318_13878.n3 gnd 0.42604f
C755 a_n2318_13878.n4 gnd 0.217886f
C756 a_n2318_13878.n5 gnd 3.16141f
C757 a_n2318_13878.n6 gnd 0.217886f
C758 a_n2318_13878.n7 gnd 0.674574f
C759 a_n2318_13878.n8 gnd 0.67455f
C760 a_n2318_13878.n9 gnd 0.206738f
C761 a_n2318_13878.n10 gnd 0.152266f
C762 a_n2318_13878.n11 gnd 0.239314f
C763 a_n2318_13878.n12 gnd 0.184843f
C764 a_n2318_13878.n13 gnd 0.206738f
C765 a_n2318_13878.n14 gnd 0.152266f
C766 a_n2318_13878.n15 gnd 0.729022f
C767 a_n2318_13878.n16 gnd 0.51701f
C768 a_n2318_13878.n17 gnd 0.217886f
C769 a_n2318_13878.n18 gnd 0.217886f
C770 a_n2318_13878.n19 gnd 0.447806f
C771 a_n2318_13878.n20 gnd 0.217886f
C772 a_n2318_13878.n21 gnd 0.217886f
C773 a_n2318_13878.n22 gnd 0.733554f
C774 a_n2318_13878.n23 gnd 2.98994f
C775 a_n2318_13878.n24 gnd 2.92523f
C776 a_n2318_13878.n25 gnd 3.7969f
C777 a_n2318_13878.n26 gnd 1.79383f
C778 a_n2318_13878.n27 gnd 1.91464f
C779 a_n2318_13878.n28 gnd 2.09784f
C780 a_n2318_13878.n29 gnd 1.79383f
C781 a_n2318_13878.n30 gnd 0.287827f
C782 a_n2318_13878.n31 gnd 0.766802f
C783 a_n2318_13878.n32 gnd 0.004897f
C784 a_n2318_13878.n33 gnd 0.010591f
C785 a_n2318_13878.n34 gnd 0.010591f
C786 a_n2318_13878.n35 gnd 0.004897f
C787 a_n2318_13878.n36 gnd 0.287827f
C788 a_n2318_13878.n37 gnd 0.287827f
C789 a_n2318_13878.n38 gnd 0.447806f
C790 a_n2318_13878.n39 gnd 0.004897f
C791 a_n2318_13878.n40 gnd 0.010591f
C792 a_n2318_13878.n41 gnd 0.010591f
C793 a_n2318_13878.n42 gnd 0.004897f
C794 a_n2318_13878.n43 gnd 0.287827f
C795 a_n2318_13878.n44 gnd 0.008436f
C796 a_n2318_13878.n45 gnd 0.287827f
C797 a_n2318_13878.n46 gnd 0.008436f
C798 a_n2318_13878.n47 gnd 0.287827f
C799 a_n2318_13878.n48 gnd 0.008436f
C800 a_n2318_13878.n49 gnd 0.287827f
C801 a_n2318_13878.n50 gnd 0.008436f
C802 a_n2318_13878.n51 gnd 1.46328f
C803 a_n2318_13878.n52 gnd 0.287827f
C804 a_n2318_13878.n53 gnd 0.287827f
C805 a_n2318_13878.n54 gnd 0.004897f
C806 a_n2318_13878.n55 gnd 0.010591f
C807 a_n2318_13878.n56 gnd 0.010591f
C808 a_n2318_13878.n57 gnd 0.004897f
C809 a_n2318_13878.n58 gnd 0.287827f
C810 a_n2318_13878.n59 gnd 0.287827f
C811 a_n2318_13878.n60 gnd 0.004897f
C812 a_n2318_13878.n61 gnd 0.010591f
C813 a_n2318_13878.n62 gnd 0.010591f
C814 a_n2318_13878.n63 gnd 0.004897f
C815 a_n2318_13878.n64 gnd 0.287827f
C816 a_n2318_13878.t47 gnd 0.151128f
C817 a_n2318_13878.t41 gnd 1.41509f
C818 a_n2318_13878.t35 gnd 0.151128f
C819 a_n2318_13878.t31 gnd 0.151128f
C820 a_n2318_13878.n65 gnd 1.06455f
C821 a_n2318_13878.t36 gnd 0.702974f
C822 a_n2318_13878.n66 gnd 0.307084f
C823 a_n2318_13878.t46 gnd 0.702974f
C824 a_n2318_13878.t40 gnd 0.714753f
C825 a_n2318_13878.t34 gnd 0.702974f
C826 a_n2318_13878.t62 gnd 0.702974f
C827 a_n2318_13878.n67 gnd 0.307084f
C828 a_n2318_13878.t76 gnd 0.702974f
C829 a_n2318_13878.t78 gnd 0.714753f
C830 a_n2318_13878.t56 gnd 0.702974f
C831 a_n2318_13878.t20 gnd 0.714753f
C832 a_n2318_13878.t26 gnd 0.702974f
C833 a_n2318_13878.t42 gnd 0.702974f
C834 a_n2318_13878.n68 gnd 0.307084f
C835 a_n2318_13878.t44 gnd 0.702974f
C836 a_n2318_13878.t22 gnd 0.702974f
C837 a_n2318_13878.t38 gnd 0.702974f
C838 a_n2318_13878.n69 gnd 0.307084f
C839 a_n2318_13878.t32 gnd 0.702974f
C840 a_n2318_13878.t28 gnd 0.714753f
C841 a_n2318_13878.t82 gnd 0.714753f
C842 a_n2318_13878.t63 gnd 0.702974f
C843 a_n2318_13878.t67 gnd 0.702974f
C844 a_n2318_13878.n70 gnd 0.307084f
C845 a_n2318_13878.t57 gnd 0.702974f
C846 a_n2318_13878.t72 gnd 0.702974f
C847 a_n2318_13878.t79 gnd 0.702974f
C848 a_n2318_13878.n71 gnd 0.307084f
C849 a_n2318_13878.t80 gnd 0.702974f
C850 a_n2318_13878.t54 gnd 0.714753f
C851 a_n2318_13878.n72 gnd 0.309588f
C852 a_n2318_13878.n73 gnd 0.30246f
C853 a_n2318_13878.n74 gnd 0.30246f
C854 a_n2318_13878.n75 gnd 0.309588f
C855 a_n2318_13878.t1 gnd 0.117544f
C856 a_n2318_13878.t17 gnd 0.117544f
C857 a_n2318_13878.n76 gnd 1.04031f
C858 a_n2318_13878.t2 gnd 0.117544f
C859 a_n2318_13878.t15 gnd 0.117544f
C860 a_n2318_13878.n77 gnd 1.03866f
C861 a_n2318_13878.t3 gnd 0.117544f
C862 a_n2318_13878.t5 gnd 0.117544f
C863 a_n2318_13878.n78 gnd 1.03866f
C864 a_n2318_13878.t4 gnd 0.117544f
C865 a_n2318_13878.t14 gnd 0.117544f
C866 a_n2318_13878.n79 gnd 1.04031f
C867 a_n2318_13878.t51 gnd 0.117544f
C868 a_n2318_13878.t9 gnd 0.117544f
C869 a_n2318_13878.n80 gnd 1.03866f
C870 a_n2318_13878.t50 gnd 0.117544f
C871 a_n2318_13878.t10 gnd 0.117544f
C872 a_n2318_13878.n81 gnd 1.03866f
C873 a_n2318_13878.t7 gnd 0.117544f
C874 a_n2318_13878.t16 gnd 0.117544f
C875 a_n2318_13878.n82 gnd 1.03866f
C876 a_n2318_13878.t11 gnd 0.117544f
C877 a_n2318_13878.t12 gnd 0.117544f
C878 a_n2318_13878.n83 gnd 1.03866f
C879 a_n2318_13878.t0 gnd 0.117544f
C880 a_n2318_13878.t6 gnd 0.117544f
C881 a_n2318_13878.n84 gnd 1.04032f
C882 a_n2318_13878.t8 gnd 0.117544f
C883 a_n2318_13878.t13 gnd 0.117544f
C884 a_n2318_13878.n85 gnd 1.03866f
C885 a_n2318_13878.n86 gnd 0.309588f
C886 a_n2318_13878.n87 gnd 0.30246f
C887 a_n2318_13878.n88 gnd 0.30246f
C888 a_n2318_13878.n89 gnd 0.309588f
C889 a_n2318_13878.t29 gnd 1.41509f
C890 a_n2318_13878.t39 gnd 0.151128f
C891 a_n2318_13878.t33 gnd 0.151128f
C892 a_n2318_13878.n90 gnd 1.06455f
C893 a_n2318_13878.t45 gnd 0.151128f
C894 a_n2318_13878.t23 gnd 0.151128f
C895 a_n2318_13878.n91 gnd 1.06455f
C896 a_n2318_13878.t27 gnd 0.151128f
C897 a_n2318_13878.t43 gnd 0.151128f
C898 a_n2318_13878.n92 gnd 1.06455f
C899 a_n2318_13878.t21 gnd 1.41227f
C900 a_n2318_13878.n93 gnd 0.867362f
C901 a_n2318_13878.t61 gnd 0.702974f
C902 a_n2318_13878.t70 gnd 0.702974f
C903 a_n2318_13878.t83 gnd 0.702974f
C904 a_n2318_13878.n94 gnd 0.309072f
C905 a_n2318_13878.t73 gnd 0.702974f
C906 a_n2318_13878.t58 gnd 0.702974f
C907 a_n2318_13878.t59 gnd 0.702974f
C908 a_n2318_13878.n95 gnd 0.309072f
C909 a_n2318_13878.t77 gnd 0.702974f
C910 a_n2318_13878.t66 gnd 0.702974f
C911 a_n2318_13878.t65 gnd 0.702974f
C912 a_n2318_13878.n96 gnd 0.309072f
C913 a_n2318_13878.t69 gnd 0.702974f
C914 a_n2318_13878.t60 gnd 0.702974f
C915 a_n2318_13878.t52 gnd 0.702974f
C916 a_n2318_13878.n97 gnd 0.309072f
C917 a_n2318_13878.t74 gnd 0.714753f
C918 a_n2318_13878.n98 gnd 0.305147f
C919 a_n2318_13878.n99 gnd 0.299606f
C920 a_n2318_13878.t81 gnd 0.714753f
C921 a_n2318_13878.n100 gnd 0.305147f
C922 a_n2318_13878.n101 gnd 0.299606f
C923 a_n2318_13878.t68 gnd 0.714753f
C924 a_n2318_13878.n102 gnd 0.305147f
C925 a_n2318_13878.n103 gnd 0.299606f
C926 a_n2318_13878.t64 gnd 0.714753f
C927 a_n2318_13878.n104 gnd 0.305147f
C928 a_n2318_13878.n105 gnd 0.299606f
C929 a_n2318_13878.n106 gnd 1.12829f
C930 a_n2318_13878.n107 gnd 0.309588f
C931 a_n2318_13878.t75 gnd 0.702974f
C932 a_n2318_13878.n108 gnd 0.307084f
C933 a_n2318_13878.n109 gnd 0.30246f
C934 a_n2318_13878.t53 gnd 0.702974f
C935 a_n2318_13878.n110 gnd 0.30246f
C936 a_n2318_13878.t71 gnd 0.702974f
C937 a_n2318_13878.n111 gnd 0.309588f
C938 a_n2318_13878.t55 gnd 0.714753f
C939 a_n2318_13878.n112 gnd 0.309588f
C940 a_n2318_13878.t30 gnd 0.702974f
C941 a_n2318_13878.n113 gnd 0.307084f
C942 a_n2318_13878.n114 gnd 0.30246f
C943 a_n2318_13878.t18 gnd 0.702974f
C944 a_n2318_13878.n115 gnd 0.30246f
C945 a_n2318_13878.t24 gnd 0.702974f
C946 a_n2318_13878.n116 gnd 0.309588f
C947 a_n2318_13878.t48 gnd 0.714753f
C948 a_n2318_13878.n117 gnd 1.20932f
C949 a_n2318_13878.t49 gnd 1.41226f
C950 a_n2318_13878.t37 gnd 0.151128f
C951 a_n2318_13878.t25 gnd 0.151128f
C952 a_n2318_13878.n118 gnd 1.06455f
C953 a_n2318_13878.n119 gnd 1.06455f
C954 a_n2318_13878.t19 gnd 0.151128f
C955 commonsourceibias.n0 gnd 0.012292f
C956 commonsourceibias.t89 gnd 0.186134f
C957 commonsourceibias.t51 gnd 0.172107f
C958 commonsourceibias.n1 gnd 0.068671f
C959 commonsourceibias.n2 gnd 0.009212f
C960 commonsourceibias.t95 gnd 0.172107f
C961 commonsourceibias.n3 gnd 0.007452f
C962 commonsourceibias.n4 gnd 0.009212f
C963 commonsourceibias.t90 gnd 0.172107f
C964 commonsourceibias.n5 gnd 0.008893f
C965 commonsourceibias.n6 gnd 0.009212f
C966 commonsourceibias.t101 gnd 0.172107f
C967 commonsourceibias.n7 gnd 0.068671f
C968 commonsourceibias.t86 gnd 0.172107f
C969 commonsourceibias.n8 gnd 0.00744f
C970 commonsourceibias.n9 gnd 0.012292f
C971 commonsourceibias.t40 gnd 0.186134f
C972 commonsourceibias.t36 gnd 0.172107f
C973 commonsourceibias.n10 gnd 0.068671f
C974 commonsourceibias.n11 gnd 0.009212f
C975 commonsourceibias.t46 gnd 0.172107f
C976 commonsourceibias.n12 gnd 0.007452f
C977 commonsourceibias.n13 gnd 0.009212f
C978 commonsourceibias.t42 gnd 0.172107f
C979 commonsourceibias.n14 gnd 0.008893f
C980 commonsourceibias.n15 gnd 0.009212f
C981 commonsourceibias.t22 gnd 0.172107f
C982 commonsourceibias.n16 gnd 0.068671f
C983 commonsourceibias.t38 gnd 0.172107f
C984 commonsourceibias.n17 gnd 0.00744f
C985 commonsourceibias.n18 gnd 0.009212f
C986 commonsourceibias.t18 gnd 0.172107f
C987 commonsourceibias.t8 gnd 0.172107f
C988 commonsourceibias.n19 gnd 0.068671f
C989 commonsourceibias.n20 gnd 0.009212f
C990 commonsourceibias.t44 gnd 0.172107f
C991 commonsourceibias.n21 gnd 0.068671f
C992 commonsourceibias.n22 gnd 0.009212f
C993 commonsourceibias.t32 gnd 0.172107f
C994 commonsourceibias.n23 gnd 0.068671f
C995 commonsourceibias.n24 gnd 0.046375f
C996 commonsourceibias.t14 gnd 0.172107f
C997 commonsourceibias.t20 gnd 0.194203f
C998 commonsourceibias.n25 gnd 0.079692f
C999 commonsourceibias.n26 gnd 0.082502f
C1000 commonsourceibias.n27 gnd 0.011354f
C1001 commonsourceibias.n28 gnd 0.012561f
C1002 commonsourceibias.n29 gnd 0.009212f
C1003 commonsourceibias.n30 gnd 0.009212f
C1004 commonsourceibias.n31 gnd 0.012479f
C1005 commonsourceibias.n32 gnd 0.007452f
C1006 commonsourceibias.n33 gnd 0.012633f
C1007 commonsourceibias.n34 gnd 0.009212f
C1008 commonsourceibias.n35 gnd 0.009212f
C1009 commonsourceibias.n36 gnd 0.01271f
C1010 commonsourceibias.n37 gnd 0.01096f
C1011 commonsourceibias.n38 gnd 0.008893f
C1012 commonsourceibias.n39 gnd 0.009212f
C1013 commonsourceibias.n40 gnd 0.009212f
C1014 commonsourceibias.n41 gnd 0.011268f
C1015 commonsourceibias.n42 gnd 0.012647f
C1016 commonsourceibias.n43 gnd 0.068671f
C1017 commonsourceibias.n44 gnd 0.012562f
C1018 commonsourceibias.n45 gnd 0.009212f
C1019 commonsourceibias.n46 gnd 0.009212f
C1020 commonsourceibias.n47 gnd 0.009212f
C1021 commonsourceibias.n48 gnd 0.012562f
C1022 commonsourceibias.n49 gnd 0.068671f
C1023 commonsourceibias.n50 gnd 0.012647f
C1024 commonsourceibias.n51 gnd 0.011268f
C1025 commonsourceibias.n52 gnd 0.009212f
C1026 commonsourceibias.n53 gnd 0.009212f
C1027 commonsourceibias.n54 gnd 0.009212f
C1028 commonsourceibias.n55 gnd 0.01096f
C1029 commonsourceibias.n56 gnd 0.01271f
C1030 commonsourceibias.n57 gnd 0.068671f
C1031 commonsourceibias.n58 gnd 0.012633f
C1032 commonsourceibias.n59 gnd 0.009212f
C1033 commonsourceibias.n60 gnd 0.009212f
C1034 commonsourceibias.n61 gnd 0.009212f
C1035 commonsourceibias.n62 gnd 0.012479f
C1036 commonsourceibias.n63 gnd 0.068671f
C1037 commonsourceibias.n64 gnd 0.012561f
C1038 commonsourceibias.n65 gnd 0.011354f
C1039 commonsourceibias.n66 gnd 0.009212f
C1040 commonsourceibias.n67 gnd 0.009212f
C1041 commonsourceibias.n68 gnd 0.009345f
C1042 commonsourceibias.n69 gnd 0.009661f
C1043 commonsourceibias.n70 gnd 0.082165f
C1044 commonsourceibias.n71 gnd 0.09115f
C1045 commonsourceibias.t41 gnd 0.019878f
C1046 commonsourceibias.t37 gnd 0.019878f
C1047 commonsourceibias.n72 gnd 0.175652f
C1048 commonsourceibias.n73 gnd 0.151777f
C1049 commonsourceibias.t47 gnd 0.019878f
C1050 commonsourceibias.t43 gnd 0.019878f
C1051 commonsourceibias.n74 gnd 0.175652f
C1052 commonsourceibias.n75 gnd 0.080684f
C1053 commonsourceibias.t23 gnd 0.019878f
C1054 commonsourceibias.t39 gnd 0.019878f
C1055 commonsourceibias.n76 gnd 0.175652f
C1056 commonsourceibias.n77 gnd 0.067408f
C1057 commonsourceibias.t15 gnd 0.019878f
C1058 commonsourceibias.t21 gnd 0.019878f
C1059 commonsourceibias.n78 gnd 0.17624f
C1060 commonsourceibias.t45 gnd 0.019878f
C1061 commonsourceibias.t33 gnd 0.019878f
C1062 commonsourceibias.n79 gnd 0.175652f
C1063 commonsourceibias.n80 gnd 0.163675f
C1064 commonsourceibias.t19 gnd 0.019878f
C1065 commonsourceibias.t9 gnd 0.019878f
C1066 commonsourceibias.n81 gnd 0.175652f
C1067 commonsourceibias.n82 gnd 0.067408f
C1068 commonsourceibias.n83 gnd 0.081623f
C1069 commonsourceibias.n84 gnd 0.009212f
C1070 commonsourceibias.t77 gnd 0.172107f
C1071 commonsourceibias.t94 gnd 0.172107f
C1072 commonsourceibias.n85 gnd 0.068671f
C1073 commonsourceibias.n86 gnd 0.009212f
C1074 commonsourceibias.t87 gnd 0.172107f
C1075 commonsourceibias.n87 gnd 0.068671f
C1076 commonsourceibias.n88 gnd 0.009212f
C1077 commonsourceibias.t58 gnd 0.172107f
C1078 commonsourceibias.n89 gnd 0.068671f
C1079 commonsourceibias.n90 gnd 0.046375f
C1080 commonsourceibias.t80 gnd 0.172107f
C1081 commonsourceibias.t73 gnd 0.194203f
C1082 commonsourceibias.n91 gnd 0.079692f
C1083 commonsourceibias.n92 gnd 0.082502f
C1084 commonsourceibias.n93 gnd 0.011354f
C1085 commonsourceibias.n94 gnd 0.012561f
C1086 commonsourceibias.n95 gnd 0.009212f
C1087 commonsourceibias.n96 gnd 0.009212f
C1088 commonsourceibias.n97 gnd 0.012479f
C1089 commonsourceibias.n98 gnd 0.007452f
C1090 commonsourceibias.n99 gnd 0.012633f
C1091 commonsourceibias.n100 gnd 0.009212f
C1092 commonsourceibias.n101 gnd 0.009212f
C1093 commonsourceibias.n102 gnd 0.01271f
C1094 commonsourceibias.n103 gnd 0.01096f
C1095 commonsourceibias.n104 gnd 0.008893f
C1096 commonsourceibias.n105 gnd 0.009212f
C1097 commonsourceibias.n106 gnd 0.009212f
C1098 commonsourceibias.n107 gnd 0.011268f
C1099 commonsourceibias.n108 gnd 0.012647f
C1100 commonsourceibias.n109 gnd 0.068671f
C1101 commonsourceibias.n110 gnd 0.012562f
C1102 commonsourceibias.n111 gnd 0.009168f
C1103 commonsourceibias.n112 gnd 0.066591f
C1104 commonsourceibias.n113 gnd 0.009168f
C1105 commonsourceibias.n114 gnd 0.012562f
C1106 commonsourceibias.n115 gnd 0.068671f
C1107 commonsourceibias.n116 gnd 0.012647f
C1108 commonsourceibias.n117 gnd 0.011268f
C1109 commonsourceibias.n118 gnd 0.009212f
C1110 commonsourceibias.n119 gnd 0.009212f
C1111 commonsourceibias.n120 gnd 0.009212f
C1112 commonsourceibias.n121 gnd 0.01096f
C1113 commonsourceibias.n122 gnd 0.01271f
C1114 commonsourceibias.n123 gnd 0.068671f
C1115 commonsourceibias.n124 gnd 0.012633f
C1116 commonsourceibias.n125 gnd 0.009212f
C1117 commonsourceibias.n126 gnd 0.009212f
C1118 commonsourceibias.n127 gnd 0.009212f
C1119 commonsourceibias.n128 gnd 0.012479f
C1120 commonsourceibias.n129 gnd 0.068671f
C1121 commonsourceibias.n130 gnd 0.012561f
C1122 commonsourceibias.n131 gnd 0.011354f
C1123 commonsourceibias.n132 gnd 0.009212f
C1124 commonsourceibias.n133 gnd 0.009212f
C1125 commonsourceibias.n134 gnd 0.009345f
C1126 commonsourceibias.n135 gnd 0.009661f
C1127 commonsourceibias.n136 gnd 0.082165f
C1128 commonsourceibias.n137 gnd 0.053193f
C1129 commonsourceibias.n138 gnd 0.012292f
C1130 commonsourceibias.t54 gnd 0.186134f
C1131 commonsourceibias.t119 gnd 0.172107f
C1132 commonsourceibias.n139 gnd 0.068671f
C1133 commonsourceibias.n140 gnd 0.009212f
C1134 commonsourceibias.t110 gnd 0.172107f
C1135 commonsourceibias.n141 gnd 0.007452f
C1136 commonsourceibias.n142 gnd 0.009212f
C1137 commonsourceibias.t60 gnd 0.172107f
C1138 commonsourceibias.n143 gnd 0.008893f
C1139 commonsourceibias.n144 gnd 0.009212f
C1140 commonsourceibias.t117 gnd 0.172107f
C1141 commonsourceibias.n145 gnd 0.068671f
C1142 commonsourceibias.t65 gnd 0.172107f
C1143 commonsourceibias.n146 gnd 0.00744f
C1144 commonsourceibias.n147 gnd 0.009212f
C1145 commonsourceibias.t59 gnd 0.172107f
C1146 commonsourceibias.t118 gnd 0.172107f
C1147 commonsourceibias.n148 gnd 0.068671f
C1148 commonsourceibias.n149 gnd 0.009212f
C1149 commonsourceibias.t71 gnd 0.172107f
C1150 commonsourceibias.n150 gnd 0.068671f
C1151 commonsourceibias.n151 gnd 0.009212f
C1152 commonsourceibias.t83 gnd 0.172107f
C1153 commonsourceibias.n152 gnd 0.068671f
C1154 commonsourceibias.n153 gnd 0.046375f
C1155 commonsourceibias.t116 gnd 0.172107f
C1156 commonsourceibias.t70 gnd 0.194203f
C1157 commonsourceibias.n154 gnd 0.079692f
C1158 commonsourceibias.n155 gnd 0.082502f
C1159 commonsourceibias.n156 gnd 0.011354f
C1160 commonsourceibias.n157 gnd 0.012561f
C1161 commonsourceibias.n158 gnd 0.009212f
C1162 commonsourceibias.n159 gnd 0.009212f
C1163 commonsourceibias.n160 gnd 0.012479f
C1164 commonsourceibias.n161 gnd 0.007452f
C1165 commonsourceibias.n162 gnd 0.012633f
C1166 commonsourceibias.n163 gnd 0.009212f
C1167 commonsourceibias.n164 gnd 0.009212f
C1168 commonsourceibias.n165 gnd 0.01271f
C1169 commonsourceibias.n166 gnd 0.01096f
C1170 commonsourceibias.n167 gnd 0.008893f
C1171 commonsourceibias.n168 gnd 0.009212f
C1172 commonsourceibias.n169 gnd 0.009212f
C1173 commonsourceibias.n170 gnd 0.011268f
C1174 commonsourceibias.n171 gnd 0.012647f
C1175 commonsourceibias.n172 gnd 0.068671f
C1176 commonsourceibias.n173 gnd 0.012562f
C1177 commonsourceibias.n174 gnd 0.009212f
C1178 commonsourceibias.n175 gnd 0.009212f
C1179 commonsourceibias.n176 gnd 0.009212f
C1180 commonsourceibias.n177 gnd 0.012562f
C1181 commonsourceibias.n178 gnd 0.068671f
C1182 commonsourceibias.n179 gnd 0.012647f
C1183 commonsourceibias.n180 gnd 0.011268f
C1184 commonsourceibias.n181 gnd 0.009212f
C1185 commonsourceibias.n182 gnd 0.009212f
C1186 commonsourceibias.n183 gnd 0.009212f
C1187 commonsourceibias.n184 gnd 0.01096f
C1188 commonsourceibias.n185 gnd 0.01271f
C1189 commonsourceibias.n186 gnd 0.068671f
C1190 commonsourceibias.n187 gnd 0.012633f
C1191 commonsourceibias.n188 gnd 0.009212f
C1192 commonsourceibias.n189 gnd 0.009212f
C1193 commonsourceibias.n190 gnd 0.009212f
C1194 commonsourceibias.n191 gnd 0.012479f
C1195 commonsourceibias.n192 gnd 0.068671f
C1196 commonsourceibias.n193 gnd 0.012561f
C1197 commonsourceibias.n194 gnd 0.011354f
C1198 commonsourceibias.n195 gnd 0.009212f
C1199 commonsourceibias.n196 gnd 0.009212f
C1200 commonsourceibias.n197 gnd 0.009345f
C1201 commonsourceibias.n198 gnd 0.009661f
C1202 commonsourceibias.n199 gnd 0.082165f
C1203 commonsourceibias.n200 gnd 0.027962f
C1204 commonsourceibias.n201 gnd 0.146988f
C1205 commonsourceibias.n202 gnd 0.012292f
C1206 commonsourceibias.t57 gnd 0.172107f
C1207 commonsourceibias.n203 gnd 0.068671f
C1208 commonsourceibias.n204 gnd 0.009212f
C1209 commonsourceibias.t96 gnd 0.172107f
C1210 commonsourceibias.n205 gnd 0.007452f
C1211 commonsourceibias.n206 gnd 0.009212f
C1212 commonsourceibias.t93 gnd 0.172107f
C1213 commonsourceibias.n207 gnd 0.008893f
C1214 commonsourceibias.n208 gnd 0.009212f
C1215 commonsourceibias.t115 gnd 0.172107f
C1216 commonsourceibias.n209 gnd 0.068671f
C1217 commonsourceibias.t68 gnd 0.172107f
C1218 commonsourceibias.n210 gnd 0.00744f
C1219 commonsourceibias.n211 gnd 0.009212f
C1220 commonsourceibias.t88 gnd 0.172107f
C1221 commonsourceibias.t108 gnd 0.172107f
C1222 commonsourceibias.n212 gnd 0.068671f
C1223 commonsourceibias.n213 gnd 0.009212f
C1224 commonsourceibias.t103 gnd 0.172107f
C1225 commonsourceibias.n214 gnd 0.068671f
C1226 commonsourceibias.n215 gnd 0.009212f
C1227 commonsourceibias.t48 gnd 0.172107f
C1228 commonsourceibias.n216 gnd 0.068671f
C1229 commonsourceibias.n217 gnd 0.046375f
C1230 commonsourceibias.t102 gnd 0.172107f
C1231 commonsourceibias.t98 gnd 0.194203f
C1232 commonsourceibias.n218 gnd 0.079692f
C1233 commonsourceibias.n219 gnd 0.082502f
C1234 commonsourceibias.n220 gnd 0.011354f
C1235 commonsourceibias.n221 gnd 0.012561f
C1236 commonsourceibias.n222 gnd 0.009212f
C1237 commonsourceibias.n223 gnd 0.009212f
C1238 commonsourceibias.n224 gnd 0.012479f
C1239 commonsourceibias.n225 gnd 0.007452f
C1240 commonsourceibias.n226 gnd 0.012633f
C1241 commonsourceibias.n227 gnd 0.009212f
C1242 commonsourceibias.n228 gnd 0.009212f
C1243 commonsourceibias.n229 gnd 0.01271f
C1244 commonsourceibias.n230 gnd 0.01096f
C1245 commonsourceibias.n231 gnd 0.008893f
C1246 commonsourceibias.n232 gnd 0.009212f
C1247 commonsourceibias.n233 gnd 0.009212f
C1248 commonsourceibias.n234 gnd 0.011268f
C1249 commonsourceibias.n235 gnd 0.012647f
C1250 commonsourceibias.n236 gnd 0.068671f
C1251 commonsourceibias.n237 gnd 0.012562f
C1252 commonsourceibias.n238 gnd 0.009212f
C1253 commonsourceibias.n239 gnd 0.009212f
C1254 commonsourceibias.n240 gnd 0.009212f
C1255 commonsourceibias.n241 gnd 0.012562f
C1256 commonsourceibias.n242 gnd 0.068671f
C1257 commonsourceibias.n243 gnd 0.012647f
C1258 commonsourceibias.n244 gnd 0.011268f
C1259 commonsourceibias.n245 gnd 0.009212f
C1260 commonsourceibias.n246 gnd 0.009212f
C1261 commonsourceibias.n247 gnd 0.009212f
C1262 commonsourceibias.n248 gnd 0.01096f
C1263 commonsourceibias.n249 gnd 0.01271f
C1264 commonsourceibias.n250 gnd 0.068671f
C1265 commonsourceibias.n251 gnd 0.012633f
C1266 commonsourceibias.n252 gnd 0.009212f
C1267 commonsourceibias.n253 gnd 0.009212f
C1268 commonsourceibias.n254 gnd 0.009212f
C1269 commonsourceibias.n255 gnd 0.012479f
C1270 commonsourceibias.n256 gnd 0.068671f
C1271 commonsourceibias.n257 gnd 0.012561f
C1272 commonsourceibias.n258 gnd 0.011354f
C1273 commonsourceibias.n259 gnd 0.009212f
C1274 commonsourceibias.n260 gnd 0.009212f
C1275 commonsourceibias.n261 gnd 0.009345f
C1276 commonsourceibias.n262 gnd 0.009661f
C1277 commonsourceibias.t109 gnd 0.186134f
C1278 commonsourceibias.n263 gnd 0.082165f
C1279 commonsourceibias.n264 gnd 0.027962f
C1280 commonsourceibias.n265 gnd 0.437625f
C1281 commonsourceibias.n266 gnd 0.012292f
C1282 commonsourceibias.t69 gnd 0.186134f
C1283 commonsourceibias.t99 gnd 0.172107f
C1284 commonsourceibias.n267 gnd 0.068671f
C1285 commonsourceibias.n268 gnd 0.009212f
C1286 commonsourceibias.t84 gnd 0.172107f
C1287 commonsourceibias.n269 gnd 0.007452f
C1288 commonsourceibias.n270 gnd 0.009212f
C1289 commonsourceibias.t72 gnd 0.172107f
C1290 commonsourceibias.n271 gnd 0.008893f
C1291 commonsourceibias.n272 gnd 0.009212f
C1292 commonsourceibias.t66 gnd 0.172107f
C1293 commonsourceibias.n273 gnd 0.00744f
C1294 commonsourceibias.n274 gnd 0.009212f
C1295 commonsourceibias.t56 gnd 0.172107f
C1296 commonsourceibias.t79 gnd 0.172107f
C1297 commonsourceibias.n275 gnd 0.068671f
C1298 commonsourceibias.n276 gnd 0.009212f
C1299 commonsourceibias.t67 gnd 0.172107f
C1300 commonsourceibias.n277 gnd 0.068671f
C1301 commonsourceibias.n278 gnd 0.009212f
C1302 commonsourceibias.t104 gnd 0.172107f
C1303 commonsourceibias.n279 gnd 0.068671f
C1304 commonsourceibias.n280 gnd 0.046375f
C1305 commonsourceibias.t64 gnd 0.172107f
C1306 commonsourceibias.t111 gnd 0.194203f
C1307 commonsourceibias.n281 gnd 0.079692f
C1308 commonsourceibias.n282 gnd 0.082502f
C1309 commonsourceibias.n283 gnd 0.011354f
C1310 commonsourceibias.n284 gnd 0.012561f
C1311 commonsourceibias.n285 gnd 0.009212f
C1312 commonsourceibias.n286 gnd 0.009212f
C1313 commonsourceibias.n287 gnd 0.012479f
C1314 commonsourceibias.n288 gnd 0.007452f
C1315 commonsourceibias.n289 gnd 0.012633f
C1316 commonsourceibias.n290 gnd 0.009212f
C1317 commonsourceibias.n291 gnd 0.009212f
C1318 commonsourceibias.n292 gnd 0.01271f
C1319 commonsourceibias.n293 gnd 0.01096f
C1320 commonsourceibias.n294 gnd 0.008893f
C1321 commonsourceibias.n295 gnd 0.009212f
C1322 commonsourceibias.n296 gnd 0.009212f
C1323 commonsourceibias.n297 gnd 0.011268f
C1324 commonsourceibias.n298 gnd 0.012647f
C1325 commonsourceibias.n299 gnd 0.068671f
C1326 commonsourceibias.n300 gnd 0.012562f
C1327 commonsourceibias.n301 gnd 0.009168f
C1328 commonsourceibias.t13 gnd 0.019878f
C1329 commonsourceibias.t31 gnd 0.019878f
C1330 commonsourceibias.n302 gnd 0.17624f
C1331 commonsourceibias.t27 gnd 0.019878f
C1332 commonsourceibias.t5 gnd 0.019878f
C1333 commonsourceibias.n303 gnd 0.175652f
C1334 commonsourceibias.n304 gnd 0.163675f
C1335 commonsourceibias.t17 gnd 0.019878f
C1336 commonsourceibias.t35 gnd 0.019878f
C1337 commonsourceibias.n305 gnd 0.175652f
C1338 commonsourceibias.n306 gnd 0.067408f
C1339 commonsourceibias.n307 gnd 0.012292f
C1340 commonsourceibias.t24 gnd 0.172107f
C1341 commonsourceibias.n308 gnd 0.068671f
C1342 commonsourceibias.n309 gnd 0.009212f
C1343 commonsourceibias.t28 gnd 0.172107f
C1344 commonsourceibias.n310 gnd 0.007452f
C1345 commonsourceibias.n311 gnd 0.009212f
C1346 commonsourceibias.t0 gnd 0.172107f
C1347 commonsourceibias.n312 gnd 0.008893f
C1348 commonsourceibias.n313 gnd 0.009212f
C1349 commonsourceibias.t6 gnd 0.172107f
C1350 commonsourceibias.n314 gnd 0.00744f
C1351 commonsourceibias.n315 gnd 0.009212f
C1352 commonsourceibias.t34 gnd 0.172107f
C1353 commonsourceibias.t16 gnd 0.172107f
C1354 commonsourceibias.n316 gnd 0.068671f
C1355 commonsourceibias.n317 gnd 0.009212f
C1356 commonsourceibias.t4 gnd 0.172107f
C1357 commonsourceibias.n318 gnd 0.068671f
C1358 commonsourceibias.n319 gnd 0.009212f
C1359 commonsourceibias.t26 gnd 0.172107f
C1360 commonsourceibias.n320 gnd 0.068671f
C1361 commonsourceibias.n321 gnd 0.046375f
C1362 commonsourceibias.t30 gnd 0.172107f
C1363 commonsourceibias.t12 gnd 0.194203f
C1364 commonsourceibias.n322 gnd 0.079692f
C1365 commonsourceibias.n323 gnd 0.082502f
C1366 commonsourceibias.n324 gnd 0.011354f
C1367 commonsourceibias.n325 gnd 0.012561f
C1368 commonsourceibias.n326 gnd 0.009212f
C1369 commonsourceibias.n327 gnd 0.009212f
C1370 commonsourceibias.n328 gnd 0.012479f
C1371 commonsourceibias.n329 gnd 0.007452f
C1372 commonsourceibias.n330 gnd 0.012633f
C1373 commonsourceibias.n331 gnd 0.009212f
C1374 commonsourceibias.n332 gnd 0.009212f
C1375 commonsourceibias.n333 gnd 0.01271f
C1376 commonsourceibias.n334 gnd 0.01096f
C1377 commonsourceibias.n335 gnd 0.008893f
C1378 commonsourceibias.n336 gnd 0.009212f
C1379 commonsourceibias.n337 gnd 0.009212f
C1380 commonsourceibias.n338 gnd 0.011268f
C1381 commonsourceibias.n339 gnd 0.012647f
C1382 commonsourceibias.n340 gnd 0.068671f
C1383 commonsourceibias.n341 gnd 0.012562f
C1384 commonsourceibias.n342 gnd 0.009212f
C1385 commonsourceibias.n343 gnd 0.009212f
C1386 commonsourceibias.n344 gnd 0.009212f
C1387 commonsourceibias.n345 gnd 0.012562f
C1388 commonsourceibias.n346 gnd 0.068671f
C1389 commonsourceibias.n347 gnd 0.012647f
C1390 commonsourceibias.t10 gnd 0.172107f
C1391 commonsourceibias.n348 gnd 0.068671f
C1392 commonsourceibias.n349 gnd 0.011268f
C1393 commonsourceibias.n350 gnd 0.009212f
C1394 commonsourceibias.n351 gnd 0.009212f
C1395 commonsourceibias.n352 gnd 0.009212f
C1396 commonsourceibias.n353 gnd 0.01096f
C1397 commonsourceibias.n354 gnd 0.01271f
C1398 commonsourceibias.n355 gnd 0.068671f
C1399 commonsourceibias.n356 gnd 0.012633f
C1400 commonsourceibias.n357 gnd 0.009212f
C1401 commonsourceibias.n358 gnd 0.009212f
C1402 commonsourceibias.n359 gnd 0.009212f
C1403 commonsourceibias.n360 gnd 0.012479f
C1404 commonsourceibias.n361 gnd 0.068671f
C1405 commonsourceibias.n362 gnd 0.012561f
C1406 commonsourceibias.n363 gnd 0.011354f
C1407 commonsourceibias.n364 gnd 0.009212f
C1408 commonsourceibias.n365 gnd 0.009212f
C1409 commonsourceibias.n366 gnd 0.009345f
C1410 commonsourceibias.n367 gnd 0.009661f
C1411 commonsourceibias.t2 gnd 0.186134f
C1412 commonsourceibias.n368 gnd 0.082165f
C1413 commonsourceibias.n369 gnd 0.09115f
C1414 commonsourceibias.t25 gnd 0.019878f
C1415 commonsourceibias.t3 gnd 0.019878f
C1416 commonsourceibias.n370 gnd 0.175652f
C1417 commonsourceibias.n371 gnd 0.151777f
C1418 commonsourceibias.t1 gnd 0.019878f
C1419 commonsourceibias.t29 gnd 0.019878f
C1420 commonsourceibias.n372 gnd 0.175652f
C1421 commonsourceibias.n373 gnd 0.080684f
C1422 commonsourceibias.t7 gnd 0.019878f
C1423 commonsourceibias.t11 gnd 0.019878f
C1424 commonsourceibias.n374 gnd 0.175652f
C1425 commonsourceibias.n375 gnd 0.067408f
C1426 commonsourceibias.n376 gnd 0.081623f
C1427 commonsourceibias.n377 gnd 0.066591f
C1428 commonsourceibias.n378 gnd 0.009168f
C1429 commonsourceibias.n379 gnd 0.012562f
C1430 commonsourceibias.n380 gnd 0.068671f
C1431 commonsourceibias.n381 gnd 0.012647f
C1432 commonsourceibias.t92 gnd 0.172107f
C1433 commonsourceibias.n382 gnd 0.068671f
C1434 commonsourceibias.n383 gnd 0.011268f
C1435 commonsourceibias.n384 gnd 0.009212f
C1436 commonsourceibias.n385 gnd 0.009212f
C1437 commonsourceibias.n386 gnd 0.009212f
C1438 commonsourceibias.n387 gnd 0.01096f
C1439 commonsourceibias.n388 gnd 0.01271f
C1440 commonsourceibias.n389 gnd 0.068671f
C1441 commonsourceibias.n390 gnd 0.012633f
C1442 commonsourceibias.n391 gnd 0.009212f
C1443 commonsourceibias.n392 gnd 0.009212f
C1444 commonsourceibias.n393 gnd 0.009212f
C1445 commonsourceibias.n394 gnd 0.012479f
C1446 commonsourceibias.n395 gnd 0.068671f
C1447 commonsourceibias.n396 gnd 0.012561f
C1448 commonsourceibias.n397 gnd 0.011354f
C1449 commonsourceibias.n398 gnd 0.009212f
C1450 commonsourceibias.n399 gnd 0.009212f
C1451 commonsourceibias.n400 gnd 0.009345f
C1452 commonsourceibias.n401 gnd 0.009661f
C1453 commonsourceibias.n402 gnd 0.082165f
C1454 commonsourceibias.n403 gnd 0.053193f
C1455 commonsourceibias.n404 gnd 0.012292f
C1456 commonsourceibias.t107 gnd 0.172107f
C1457 commonsourceibias.n405 gnd 0.068671f
C1458 commonsourceibias.n406 gnd 0.009212f
C1459 commonsourceibias.t50 gnd 0.172107f
C1460 commonsourceibias.n407 gnd 0.007452f
C1461 commonsourceibias.n408 gnd 0.009212f
C1462 commonsourceibias.t114 gnd 0.172107f
C1463 commonsourceibias.n409 gnd 0.008893f
C1464 commonsourceibias.n410 gnd 0.009212f
C1465 commonsourceibias.t49 gnd 0.172107f
C1466 commonsourceibias.n411 gnd 0.00744f
C1467 commonsourceibias.n412 gnd 0.009212f
C1468 commonsourceibias.t74 gnd 0.172107f
C1469 commonsourceibias.t105 gnd 0.172107f
C1470 commonsourceibias.n413 gnd 0.068671f
C1471 commonsourceibias.n414 gnd 0.009212f
C1472 commonsourceibias.t55 gnd 0.172107f
C1473 commonsourceibias.n415 gnd 0.068671f
C1474 commonsourceibias.n416 gnd 0.009212f
C1475 commonsourceibias.t75 gnd 0.172107f
C1476 commonsourceibias.n417 gnd 0.068671f
C1477 commonsourceibias.n418 gnd 0.046375f
C1478 commonsourceibias.t61 gnd 0.172107f
C1479 commonsourceibias.t52 gnd 0.194203f
C1480 commonsourceibias.n419 gnd 0.079692f
C1481 commonsourceibias.n420 gnd 0.082502f
C1482 commonsourceibias.n421 gnd 0.011354f
C1483 commonsourceibias.n422 gnd 0.012561f
C1484 commonsourceibias.n423 gnd 0.009212f
C1485 commonsourceibias.n424 gnd 0.009212f
C1486 commonsourceibias.n425 gnd 0.012479f
C1487 commonsourceibias.n426 gnd 0.007452f
C1488 commonsourceibias.n427 gnd 0.012633f
C1489 commonsourceibias.n428 gnd 0.009212f
C1490 commonsourceibias.n429 gnd 0.009212f
C1491 commonsourceibias.n430 gnd 0.01271f
C1492 commonsourceibias.n431 gnd 0.01096f
C1493 commonsourceibias.n432 gnd 0.008893f
C1494 commonsourceibias.n433 gnd 0.009212f
C1495 commonsourceibias.n434 gnd 0.009212f
C1496 commonsourceibias.n435 gnd 0.011268f
C1497 commonsourceibias.n436 gnd 0.012647f
C1498 commonsourceibias.n437 gnd 0.068671f
C1499 commonsourceibias.n438 gnd 0.012562f
C1500 commonsourceibias.n439 gnd 0.009212f
C1501 commonsourceibias.n440 gnd 0.009212f
C1502 commonsourceibias.n441 gnd 0.009212f
C1503 commonsourceibias.n442 gnd 0.012562f
C1504 commonsourceibias.n443 gnd 0.068671f
C1505 commonsourceibias.n444 gnd 0.012647f
C1506 commonsourceibias.t106 gnd 0.172107f
C1507 commonsourceibias.n445 gnd 0.068671f
C1508 commonsourceibias.n446 gnd 0.011268f
C1509 commonsourceibias.n447 gnd 0.009212f
C1510 commonsourceibias.n448 gnd 0.009212f
C1511 commonsourceibias.n449 gnd 0.009212f
C1512 commonsourceibias.n450 gnd 0.01096f
C1513 commonsourceibias.n451 gnd 0.01271f
C1514 commonsourceibias.n452 gnd 0.068671f
C1515 commonsourceibias.n453 gnd 0.012633f
C1516 commonsourceibias.n454 gnd 0.009212f
C1517 commonsourceibias.n455 gnd 0.009212f
C1518 commonsourceibias.n456 gnd 0.009212f
C1519 commonsourceibias.n457 gnd 0.012479f
C1520 commonsourceibias.n458 gnd 0.068671f
C1521 commonsourceibias.n459 gnd 0.012561f
C1522 commonsourceibias.n460 gnd 0.011354f
C1523 commonsourceibias.n461 gnd 0.009212f
C1524 commonsourceibias.n462 gnd 0.009212f
C1525 commonsourceibias.n463 gnd 0.009345f
C1526 commonsourceibias.n464 gnd 0.009661f
C1527 commonsourceibias.t112 gnd 0.186134f
C1528 commonsourceibias.n465 gnd 0.082165f
C1529 commonsourceibias.n466 gnd 0.027962f
C1530 commonsourceibias.n467 gnd 0.146988f
C1531 commonsourceibias.n468 gnd 0.012292f
C1532 commonsourceibias.t81 gnd 0.172107f
C1533 commonsourceibias.n469 gnd 0.068671f
C1534 commonsourceibias.n470 gnd 0.009212f
C1535 commonsourceibias.t91 gnd 0.172107f
C1536 commonsourceibias.n471 gnd 0.007452f
C1537 commonsourceibias.n472 gnd 0.009212f
C1538 commonsourceibias.t100 gnd 0.172107f
C1539 commonsourceibias.n473 gnd 0.008893f
C1540 commonsourceibias.n474 gnd 0.009212f
C1541 commonsourceibias.t85 gnd 0.172107f
C1542 commonsourceibias.n475 gnd 0.00744f
C1543 commonsourceibias.n476 gnd 0.009212f
C1544 commonsourceibias.t82 gnd 0.172107f
C1545 commonsourceibias.t62 gnd 0.172107f
C1546 commonsourceibias.n477 gnd 0.068671f
C1547 commonsourceibias.n478 gnd 0.009212f
C1548 commonsourceibias.t53 gnd 0.172107f
C1549 commonsourceibias.n479 gnd 0.068671f
C1550 commonsourceibias.n480 gnd 0.009212f
C1551 commonsourceibias.t78 gnd 0.172107f
C1552 commonsourceibias.n481 gnd 0.068671f
C1553 commonsourceibias.n482 gnd 0.046375f
C1554 commonsourceibias.t97 gnd 0.172107f
C1555 commonsourceibias.t113 gnd 0.194203f
C1556 commonsourceibias.n483 gnd 0.079692f
C1557 commonsourceibias.n484 gnd 0.082502f
C1558 commonsourceibias.n485 gnd 0.011354f
C1559 commonsourceibias.n486 gnd 0.012561f
C1560 commonsourceibias.n487 gnd 0.009212f
C1561 commonsourceibias.n488 gnd 0.009212f
C1562 commonsourceibias.n489 gnd 0.012479f
C1563 commonsourceibias.n490 gnd 0.007452f
C1564 commonsourceibias.n491 gnd 0.012633f
C1565 commonsourceibias.n492 gnd 0.009212f
C1566 commonsourceibias.n493 gnd 0.009212f
C1567 commonsourceibias.n494 gnd 0.01271f
C1568 commonsourceibias.n495 gnd 0.01096f
C1569 commonsourceibias.n496 gnd 0.008893f
C1570 commonsourceibias.n497 gnd 0.009212f
C1571 commonsourceibias.n498 gnd 0.009212f
C1572 commonsourceibias.n499 gnd 0.011268f
C1573 commonsourceibias.n500 gnd 0.012647f
C1574 commonsourceibias.n501 gnd 0.068671f
C1575 commonsourceibias.n502 gnd 0.012562f
C1576 commonsourceibias.n503 gnd 0.009212f
C1577 commonsourceibias.n504 gnd 0.009212f
C1578 commonsourceibias.n505 gnd 0.009212f
C1579 commonsourceibias.n506 gnd 0.012562f
C1580 commonsourceibias.n507 gnd 0.068671f
C1581 commonsourceibias.n508 gnd 0.012647f
C1582 commonsourceibias.t76 gnd 0.172107f
C1583 commonsourceibias.n509 gnd 0.068671f
C1584 commonsourceibias.n510 gnd 0.011268f
C1585 commonsourceibias.n511 gnd 0.009212f
C1586 commonsourceibias.n512 gnd 0.009212f
C1587 commonsourceibias.n513 gnd 0.009212f
C1588 commonsourceibias.n514 gnd 0.01096f
C1589 commonsourceibias.n515 gnd 0.01271f
C1590 commonsourceibias.n516 gnd 0.068671f
C1591 commonsourceibias.n517 gnd 0.012633f
C1592 commonsourceibias.n518 gnd 0.009212f
C1593 commonsourceibias.n519 gnd 0.009212f
C1594 commonsourceibias.n520 gnd 0.009212f
C1595 commonsourceibias.n521 gnd 0.012479f
C1596 commonsourceibias.n522 gnd 0.068671f
C1597 commonsourceibias.n523 gnd 0.012561f
C1598 commonsourceibias.n524 gnd 0.011354f
C1599 commonsourceibias.n525 gnd 0.009212f
C1600 commonsourceibias.n526 gnd 0.009212f
C1601 commonsourceibias.n527 gnd 0.009345f
C1602 commonsourceibias.n528 gnd 0.009661f
C1603 commonsourceibias.t63 gnd 0.186134f
C1604 commonsourceibias.n529 gnd 0.082165f
C1605 commonsourceibias.n530 gnd 0.027962f
C1606 commonsourceibias.n531 gnd 0.194173f
C1607 commonsourceibias.n532 gnd 4.69557f
C1608 CSoutput.n0 gnd 0.04929f
C1609 CSoutput.t194 gnd 0.326046f
C1610 CSoutput.n1 gnd 0.147226f
C1611 CSoutput.n2 gnd 0.04929f
C1612 CSoutput.t199 gnd 0.326046f
C1613 CSoutput.n3 gnd 0.039067f
C1614 CSoutput.n4 gnd 0.04929f
C1615 CSoutput.t211 gnd 0.326046f
C1616 CSoutput.n5 gnd 0.033687f
C1617 CSoutput.n6 gnd 0.04929f
C1618 CSoutput.t196 gnd 0.326046f
C1619 CSoutput.t204 gnd 0.326046f
C1620 CSoutput.n7 gnd 0.145621f
C1621 CSoutput.n8 gnd 0.04929f
C1622 CSoutput.t202 gnd 0.326046f
C1623 CSoutput.n9 gnd 0.032119f
C1624 CSoutput.n10 gnd 0.04929f
C1625 CSoutput.t212 gnd 0.326046f
C1626 CSoutput.t200 gnd 0.326046f
C1627 CSoutput.n11 gnd 0.145621f
C1628 CSoutput.n12 gnd 0.04929f
C1629 CSoutput.t198 gnd 0.326046f
C1630 CSoutput.n13 gnd 0.033687f
C1631 CSoutput.n14 gnd 0.04929f
C1632 CSoutput.t210 gnd 0.326046f
C1633 CSoutput.t192 gnd 0.326046f
C1634 CSoutput.n15 gnd 0.145621f
C1635 CSoutput.n16 gnd 0.04929f
C1636 CSoutput.t195 gnd 0.326046f
C1637 CSoutput.n17 gnd 0.03598f
C1638 CSoutput.t206 gnd 0.389633f
C1639 CSoutput.t209 gnd 0.326046f
C1640 CSoutput.n18 gnd 0.185902f
C1641 CSoutput.n19 gnd 0.180389f
C1642 CSoutput.n20 gnd 0.209273f
C1643 CSoutput.n21 gnd 0.04929f
C1644 CSoutput.n22 gnd 0.041138f
C1645 CSoutput.n23 gnd 0.145621f
C1646 CSoutput.n24 gnd 0.039656f
C1647 CSoutput.n25 gnd 0.039067f
C1648 CSoutput.n26 gnd 0.04929f
C1649 CSoutput.n27 gnd 0.04929f
C1650 CSoutput.n28 gnd 0.040822f
C1651 CSoutput.n29 gnd 0.034659f
C1652 CSoutput.n30 gnd 0.148863f
C1653 CSoutput.n31 gnd 0.035136f
C1654 CSoutput.n32 gnd 0.04929f
C1655 CSoutput.n33 gnd 0.04929f
C1656 CSoutput.n34 gnd 0.04929f
C1657 CSoutput.n35 gnd 0.040387f
C1658 CSoutput.n36 gnd 0.145621f
C1659 CSoutput.n37 gnd 0.038624f
C1660 CSoutput.n38 gnd 0.040098f
C1661 CSoutput.n39 gnd 0.04929f
C1662 CSoutput.n40 gnd 0.04929f
C1663 CSoutput.n41 gnd 0.04113f
C1664 CSoutput.n42 gnd 0.037593f
C1665 CSoutput.n43 gnd 0.145621f
C1666 CSoutput.n44 gnd 0.038546f
C1667 CSoutput.n45 gnd 0.04929f
C1668 CSoutput.n46 gnd 0.04929f
C1669 CSoutput.n47 gnd 0.04929f
C1670 CSoutput.n48 gnd 0.038546f
C1671 CSoutput.n49 gnd 0.145621f
C1672 CSoutput.n50 gnd 0.037593f
C1673 CSoutput.n51 gnd 0.04113f
C1674 CSoutput.n52 gnd 0.04929f
C1675 CSoutput.n53 gnd 0.04929f
C1676 CSoutput.n54 gnd 0.040098f
C1677 CSoutput.n55 gnd 0.038624f
C1678 CSoutput.n56 gnd 0.145621f
C1679 CSoutput.n57 gnd 0.040387f
C1680 CSoutput.n58 gnd 0.04929f
C1681 CSoutput.n59 gnd 0.04929f
C1682 CSoutput.n60 gnd 0.04929f
C1683 CSoutput.n61 gnd 0.035136f
C1684 CSoutput.n62 gnd 0.148863f
C1685 CSoutput.n63 gnd 0.034659f
C1686 CSoutput.t205 gnd 0.326046f
C1687 CSoutput.n64 gnd 0.145621f
C1688 CSoutput.n65 gnd 0.040822f
C1689 CSoutput.n66 gnd 0.04929f
C1690 CSoutput.n67 gnd 0.04929f
C1691 CSoutput.n68 gnd 0.04929f
C1692 CSoutput.n69 gnd 0.039656f
C1693 CSoutput.n70 gnd 0.145621f
C1694 CSoutput.n71 gnd 0.041138f
C1695 CSoutput.n72 gnd 0.03598f
C1696 CSoutput.n73 gnd 0.04929f
C1697 CSoutput.n74 gnd 0.04929f
C1698 CSoutput.n75 gnd 0.037314f
C1699 CSoutput.n76 gnd 0.022161f
C1700 CSoutput.t208 gnd 0.366336f
C1701 CSoutput.n77 gnd 0.181981f
C1702 CSoutput.n78 gnd 0.744474f
C1703 CSoutput.t161 gnd 0.061483f
C1704 CSoutput.t92 gnd 0.061483f
C1705 CSoutput.n79 gnd 0.476021f
C1706 CSoutput.t176 gnd 0.061483f
C1707 CSoutput.t114 gnd 0.061483f
C1708 CSoutput.n80 gnd 0.475172f
C1709 CSoutput.n81 gnd 0.482299f
C1710 CSoutput.t71 gnd 0.061483f
C1711 CSoutput.t131 gnd 0.061483f
C1712 CSoutput.n82 gnd 0.475172f
C1713 CSoutput.n83 gnd 0.237657f
C1714 CSoutput.t77 gnd 0.061483f
C1715 CSoutput.t105 gnd 0.061483f
C1716 CSoutput.n84 gnd 0.475172f
C1717 CSoutput.n85 gnd 0.237657f
C1718 CSoutput.t181 gnd 0.061483f
C1719 CSoutput.t124 gnd 0.061483f
C1720 CSoutput.n86 gnd 0.475172f
C1721 CSoutput.n87 gnd 0.237657f
C1722 CSoutput.t80 gnd 0.061483f
C1723 CSoutput.t165 gnd 0.061483f
C1724 CSoutput.n88 gnd 0.475172f
C1725 CSoutput.n89 gnd 0.237657f
C1726 CSoutput.t88 gnd 0.061483f
C1727 CSoutput.t141 gnd 0.061483f
C1728 CSoutput.n90 gnd 0.475172f
C1729 CSoutput.n91 gnd 0.237657f
C1730 CSoutput.t109 gnd 0.061483f
C1731 CSoutput.t132 gnd 0.061483f
C1732 CSoutput.n92 gnd 0.475172f
C1733 CSoutput.n93 gnd 0.237657f
C1734 CSoutput.t127 gnd 0.061483f
C1735 CSoutput.t170 gnd 0.061483f
C1736 CSoutput.n94 gnd 0.475172f
C1737 CSoutput.n95 gnd 0.237657f
C1738 CSoutput.t97 gnd 0.061483f
C1739 CSoutput.t148 gnd 0.061483f
C1740 CSoutput.n96 gnd 0.475172f
C1741 CSoutput.n97 gnd 0.435807f
C1742 CSoutput.t67 gnd 0.061483f
C1743 CSoutput.t159 gnd 0.061483f
C1744 CSoutput.n98 gnd 0.476021f
C1745 CSoutput.t142 gnd 0.061483f
C1746 CSoutput.t118 gnd 0.061483f
C1747 CSoutput.n99 gnd 0.475172f
C1748 CSoutput.n100 gnd 0.482299f
C1749 CSoutput.t93 gnd 0.061483f
C1750 CSoutput.t172 gnd 0.061483f
C1751 CSoutput.n101 gnd 0.475172f
C1752 CSoutput.n102 gnd 0.237657f
C1753 CSoutput.t139 gnd 0.061483f
C1754 CSoutput.t138 gnd 0.061483f
C1755 CSoutput.n103 gnd 0.475172f
C1756 CSoutput.n104 gnd 0.237657f
C1757 CSoutput.t128 gnd 0.061483f
C1758 CSoutput.t89 gnd 0.061483f
C1759 CSoutput.n105 gnd 0.475172f
C1760 CSoutput.n106 gnd 0.237657f
C1761 CSoutput.t70 gnd 0.061483f
C1762 CSoutput.t129 gnd 0.061483f
C1763 CSoutput.n107 gnd 0.475172f
C1764 CSoutput.n108 gnd 0.237657f
C1765 CSoutput.t125 gnd 0.061483f
C1766 CSoutput.t87 gnd 0.061483f
C1767 CSoutput.n109 gnd 0.475172f
C1768 CSoutput.n110 gnd 0.237657f
C1769 CSoutput.t68 gnd 0.061483f
C1770 CSoutput.t65 gnd 0.061483f
C1771 CSoutput.n111 gnd 0.475172f
C1772 CSoutput.n112 gnd 0.237657f
C1773 CSoutput.t143 gnd 0.061483f
C1774 CSoutput.t106 gnd 0.061483f
C1775 CSoutput.n113 gnd 0.475172f
C1776 CSoutput.n114 gnd 0.237657f
C1777 CSoutput.t99 gnd 0.061483f
C1778 CSoutput.t63 gnd 0.061483f
C1779 CSoutput.n115 gnd 0.475172f
C1780 CSoutput.n116 gnd 0.354406f
C1781 CSoutput.n117 gnd 0.446904f
C1782 CSoutput.t82 gnd 0.061483f
C1783 CSoutput.t171 gnd 0.061483f
C1784 CSoutput.n118 gnd 0.476021f
C1785 CSoutput.t152 gnd 0.061483f
C1786 CSoutput.t130 gnd 0.061483f
C1787 CSoutput.n119 gnd 0.475172f
C1788 CSoutput.n120 gnd 0.482299f
C1789 CSoutput.t110 gnd 0.061483f
C1790 CSoutput.t182 gnd 0.061483f
C1791 CSoutput.n121 gnd 0.475172f
C1792 CSoutput.n122 gnd 0.237657f
C1793 CSoutput.t151 gnd 0.061483f
C1794 CSoutput.t150 gnd 0.061483f
C1795 CSoutput.n123 gnd 0.475172f
C1796 CSoutput.n124 gnd 0.237657f
C1797 CSoutput.t136 gnd 0.061483f
C1798 CSoutput.t107 gnd 0.061483f
C1799 CSoutput.n125 gnd 0.475172f
C1800 CSoutput.n126 gnd 0.237657f
C1801 CSoutput.t84 gnd 0.061483f
C1802 CSoutput.t137 gnd 0.061483f
C1803 CSoutput.n127 gnd 0.475172f
C1804 CSoutput.n128 gnd 0.237657f
C1805 CSoutput.t135 gnd 0.061483f
C1806 CSoutput.t104 gnd 0.061483f
C1807 CSoutput.n129 gnd 0.475172f
C1808 CSoutput.n130 gnd 0.237657f
C1809 CSoutput.t83 gnd 0.061483f
C1810 CSoutput.t81 gnd 0.061483f
C1811 CSoutput.n131 gnd 0.475172f
C1812 CSoutput.n132 gnd 0.237657f
C1813 CSoutput.t153 gnd 0.061483f
C1814 CSoutput.t120 gnd 0.061483f
C1815 CSoutput.n133 gnd 0.475172f
C1816 CSoutput.n134 gnd 0.237657f
C1817 CSoutput.t115 gnd 0.061483f
C1818 CSoutput.t76 gnd 0.061483f
C1819 CSoutput.n135 gnd 0.475172f
C1820 CSoutput.n136 gnd 0.354406f
C1821 CSoutput.n137 gnd 0.499524f
C1822 CSoutput.n138 gnd 8.64687f
C1823 CSoutput.n140 gnd 0.871939f
C1824 CSoutput.n141 gnd 0.653954f
C1825 CSoutput.n142 gnd 0.871939f
C1826 CSoutput.n143 gnd 0.871939f
C1827 CSoutput.n144 gnd 2.34753f
C1828 CSoutput.n145 gnd 0.871939f
C1829 CSoutput.n146 gnd 0.871939f
C1830 CSoutput.t213 gnd 1.08992f
C1831 CSoutput.n147 gnd 0.871939f
C1832 CSoutput.n148 gnd 0.871939f
C1833 CSoutput.n152 gnd 0.871939f
C1834 CSoutput.n156 gnd 0.871939f
C1835 CSoutput.n157 gnd 0.871939f
C1836 CSoutput.n159 gnd 0.871939f
C1837 CSoutput.n164 gnd 0.871939f
C1838 CSoutput.n166 gnd 0.871939f
C1839 CSoutput.n167 gnd 0.871939f
C1840 CSoutput.n169 gnd 0.871939f
C1841 CSoutput.n170 gnd 0.871939f
C1842 CSoutput.n172 gnd 0.871939f
C1843 CSoutput.t201 gnd 14.57f
C1844 CSoutput.n174 gnd 0.871939f
C1845 CSoutput.n175 gnd 0.653954f
C1846 CSoutput.n176 gnd 0.871939f
C1847 CSoutput.n177 gnd 0.871939f
C1848 CSoutput.n178 gnd 2.34753f
C1849 CSoutput.n179 gnd 0.871939f
C1850 CSoutput.n180 gnd 0.871939f
C1851 CSoutput.t197 gnd 1.08992f
C1852 CSoutput.n181 gnd 0.871939f
C1853 CSoutput.n182 gnd 0.871939f
C1854 CSoutput.n186 gnd 0.871939f
C1855 CSoutput.n190 gnd 0.871939f
C1856 CSoutput.n191 gnd 0.871939f
C1857 CSoutput.n193 gnd 0.871939f
C1858 CSoutput.n198 gnd 0.871939f
C1859 CSoutput.n200 gnd 0.871939f
C1860 CSoutput.n201 gnd 0.871939f
C1861 CSoutput.n203 gnd 0.871939f
C1862 CSoutput.n204 gnd 0.871939f
C1863 CSoutput.n206 gnd 0.871939f
C1864 CSoutput.n207 gnd 0.653954f
C1865 CSoutput.n209 gnd 0.871939f
C1866 CSoutput.n210 gnd 0.653954f
C1867 CSoutput.n211 gnd 0.871939f
C1868 CSoutput.n212 gnd 0.871939f
C1869 CSoutput.n213 gnd 2.34753f
C1870 CSoutput.n214 gnd 0.871939f
C1871 CSoutput.n215 gnd 0.871939f
C1872 CSoutput.t193 gnd 1.08992f
C1873 CSoutput.n216 gnd 0.871939f
C1874 CSoutput.n217 gnd 2.34753f
C1875 CSoutput.n219 gnd 0.871939f
C1876 CSoutput.n220 gnd 0.871939f
C1877 CSoutput.n222 gnd 0.871939f
C1878 CSoutput.n223 gnd 0.871939f
C1879 CSoutput.t203 gnd 14.332601f
C1880 CSoutput.t207 gnd 14.57f
C1881 CSoutput.n229 gnd 2.7354f
C1882 CSoutput.n230 gnd 11.143f
C1883 CSoutput.n231 gnd 11.6093f
C1884 CSoutput.n236 gnd 2.96318f
C1885 CSoutput.n242 gnd 0.871939f
C1886 CSoutput.n244 gnd 0.871939f
C1887 CSoutput.n246 gnd 0.871939f
C1888 CSoutput.n248 gnd 0.871939f
C1889 CSoutput.n250 gnd 0.871939f
C1890 CSoutput.n256 gnd 0.871939f
C1891 CSoutput.n263 gnd 1.59967f
C1892 CSoutput.n264 gnd 1.59967f
C1893 CSoutput.n265 gnd 0.871939f
C1894 CSoutput.n266 gnd 0.871939f
C1895 CSoutput.n268 gnd 0.653954f
C1896 CSoutput.n269 gnd 0.560053f
C1897 CSoutput.n271 gnd 0.653954f
C1898 CSoutput.n272 gnd 0.560053f
C1899 CSoutput.n273 gnd 0.653954f
C1900 CSoutput.n275 gnd 0.871939f
C1901 CSoutput.n277 gnd 2.34753f
C1902 CSoutput.n278 gnd 2.7354f
C1903 CSoutput.n279 gnd 10.2487f
C1904 CSoutput.n281 gnd 0.653954f
C1905 CSoutput.n282 gnd 1.68266f
C1906 CSoutput.n283 gnd 0.653954f
C1907 CSoutput.n285 gnd 0.871939f
C1908 CSoutput.n287 gnd 2.34753f
C1909 CSoutput.n288 gnd 5.1133f
C1910 CSoutput.t91 gnd 0.061483f
C1911 CSoutput.t160 gnd 0.061483f
C1912 CSoutput.n289 gnd 0.476021f
C1913 CSoutput.t113 gnd 0.061483f
C1914 CSoutput.t174 gnd 0.061483f
C1915 CSoutput.n290 gnd 0.475172f
C1916 CSoutput.n291 gnd 0.482299f
C1917 CSoutput.t154 gnd 0.061483f
C1918 CSoutput.t69 gnd 0.061483f
C1919 CSoutput.n292 gnd 0.475172f
C1920 CSoutput.n293 gnd 0.237657f
C1921 CSoutput.t103 gnd 0.061483f
C1922 CSoutput.t75 gnd 0.061483f
C1923 CSoutput.n294 gnd 0.475172f
C1924 CSoutput.n295 gnd 0.237657f
C1925 CSoutput.t123 gnd 0.061483f
C1926 CSoutput.t96 gnd 0.061483f
C1927 CSoutput.n296 gnd 0.475172f
C1928 CSoutput.n297 gnd 0.237657f
C1929 CSoutput.t164 gnd 0.061483f
C1930 CSoutput.t79 gnd 0.061483f
C1931 CSoutput.n298 gnd 0.475172f
C1932 CSoutput.n299 gnd 0.237657f
C1933 CSoutput.t140 gnd 0.061483f
C1934 CSoutput.t85 gnd 0.061483f
C1935 CSoutput.n300 gnd 0.475172f
C1936 CSoutput.n301 gnd 0.237657f
C1937 CSoutput.t156 gnd 0.061483f
C1938 CSoutput.t108 gnd 0.061483f
C1939 CSoutput.n302 gnd 0.475172f
C1940 CSoutput.n303 gnd 0.237657f
C1941 CSoutput.t169 gnd 0.061483f
C1942 CSoutput.t126 gnd 0.061483f
C1943 CSoutput.n304 gnd 0.475172f
C1944 CSoutput.n305 gnd 0.237657f
C1945 CSoutput.t147 gnd 0.061483f
C1946 CSoutput.t98 gnd 0.061483f
C1947 CSoutput.n306 gnd 0.475172f
C1948 CSoutput.n307 gnd 0.435807f
C1949 CSoutput.t122 gnd 0.061483f
C1950 CSoutput.t146 gnd 0.061483f
C1951 CSoutput.n308 gnd 0.476021f
C1952 CSoutput.t64 gnd 0.061483f
C1953 CSoutput.t101 gnd 0.061483f
C1954 CSoutput.n309 gnd 0.475172f
C1955 CSoutput.n310 gnd 0.482299f
C1956 CSoutput.t102 gnd 0.061483f
C1957 CSoutput.t168 gnd 0.061483f
C1958 CSoutput.n311 gnd 0.475172f
C1959 CSoutput.n312 gnd 0.237657f
C1960 CSoutput.t94 gnd 0.061483f
C1961 CSoutput.t95 gnd 0.061483f
C1962 CSoutput.n313 gnd 0.475172f
C1963 CSoutput.n314 gnd 0.237657f
C1964 CSoutput.t166 gnd 0.061483f
C1965 CSoutput.t167 gnd 0.061483f
C1966 CSoutput.n315 gnd 0.475172f
C1967 CSoutput.n316 gnd 0.237657f
C1968 CSoutput.t74 gnd 0.061483f
C1969 CSoutput.t149 gnd 0.061483f
C1970 CSoutput.n317 gnd 0.475172f
C1971 CSoutput.n318 gnd 0.237657f
C1972 CSoutput.t163 gnd 0.061483f
C1973 CSoutput.t72 gnd 0.061483f
C1974 CSoutput.n319 gnd 0.475172f
C1975 CSoutput.n320 gnd 0.237657f
C1976 CSoutput.t121 gnd 0.061483f
C1977 CSoutput.t145 gnd 0.061483f
C1978 CSoutput.n321 gnd 0.475172f
C1979 CSoutput.n322 gnd 0.237657f
C1980 CSoutput.t175 gnd 0.061483f
C1981 CSoutput.t100 gnd 0.061483f
C1982 CSoutput.n323 gnd 0.475172f
C1983 CSoutput.n324 gnd 0.237657f
C1984 CSoutput.t144 gnd 0.061483f
C1985 CSoutput.t180 gnd 0.061483f
C1986 CSoutput.n325 gnd 0.475172f
C1987 CSoutput.n326 gnd 0.354406f
C1988 CSoutput.n327 gnd 0.446904f
C1989 CSoutput.t133 gnd 0.061483f
C1990 CSoutput.t157 gnd 0.061483f
C1991 CSoutput.n328 gnd 0.476021f
C1992 CSoutput.t78 gnd 0.061483f
C1993 CSoutput.t116 gnd 0.061483f
C1994 CSoutput.n329 gnd 0.475172f
C1995 CSoutput.n330 gnd 0.482299f
C1996 CSoutput.t119 gnd 0.061483f
C1997 CSoutput.t179 gnd 0.061483f
C1998 CSoutput.n331 gnd 0.475172f
C1999 CSoutput.n332 gnd 0.237657f
C2000 CSoutput.t111 gnd 0.061483f
C2001 CSoutput.t112 gnd 0.061483f
C2002 CSoutput.n333 gnd 0.475172f
C2003 CSoutput.n334 gnd 0.237657f
C2004 CSoutput.t177 gnd 0.061483f
C2005 CSoutput.t178 gnd 0.061483f
C2006 CSoutput.n335 gnd 0.475172f
C2007 CSoutput.n336 gnd 0.237657f
C2008 CSoutput.t90 gnd 0.061483f
C2009 CSoutput.t162 gnd 0.061483f
C2010 CSoutput.n337 gnd 0.475172f
C2011 CSoutput.n338 gnd 0.237657f
C2012 CSoutput.t173 gnd 0.061483f
C2013 CSoutput.t86 gnd 0.061483f
C2014 CSoutput.n339 gnd 0.475172f
C2015 CSoutput.n340 gnd 0.237657f
C2016 CSoutput.t134 gnd 0.061483f
C2017 CSoutput.t158 gnd 0.061483f
C2018 CSoutput.n341 gnd 0.475172f
C2019 CSoutput.n342 gnd 0.237657f
C2020 CSoutput.t66 gnd 0.061483f
C2021 CSoutput.t117 gnd 0.061483f
C2022 CSoutput.n343 gnd 0.475172f
C2023 CSoutput.n344 gnd 0.237657f
C2024 CSoutput.t155 gnd 0.061483f
C2025 CSoutput.t73 gnd 0.061483f
C2026 CSoutput.n345 gnd 0.47517f
C2027 CSoutput.n346 gnd 0.354408f
C2028 CSoutput.n347 gnd 0.499524f
C2029 CSoutput.n348 gnd 12.6711f
C2030 CSoutput.t5 gnd 0.053798f
C2031 CSoutput.t33 gnd 0.053798f
C2032 CSoutput.n349 gnd 0.476965f
C2033 CSoutput.t55 gnd 0.053798f
C2034 CSoutput.t15 gnd 0.053798f
C2035 CSoutput.n350 gnd 0.475374f
C2036 CSoutput.n351 gnd 0.44296f
C2037 CSoutput.t41 gnd 0.053798f
C2038 CSoutput.t13 gnd 0.053798f
C2039 CSoutput.n352 gnd 0.475374f
C2040 CSoutput.n353 gnd 0.218358f
C2041 CSoutput.t21 gnd 0.053798f
C2042 CSoutput.t54 gnd 0.053798f
C2043 CSoutput.n354 gnd 0.475374f
C2044 CSoutput.n355 gnd 0.218358f
C2045 CSoutput.t187 gnd 0.053798f
C2046 CSoutput.t185 gnd 0.053798f
C2047 CSoutput.n356 gnd 0.475374f
C2048 CSoutput.n357 gnd 0.218358f
C2049 CSoutput.t24 gnd 0.053798f
C2050 CSoutput.t8 gnd 0.053798f
C2051 CSoutput.n358 gnd 0.475374f
C2052 CSoutput.n359 gnd 0.40275f
C2053 CSoutput.t29 gnd 0.053798f
C2054 CSoutput.t191 gnd 0.053798f
C2055 CSoutput.n360 gnd 0.476965f
C2056 CSoutput.t56 gnd 0.053798f
C2057 CSoutput.t51 gnd 0.053798f
C2058 CSoutput.n361 gnd 0.475374f
C2059 CSoutput.n362 gnd 0.44296f
C2060 CSoutput.t28 gnd 0.053798f
C2061 CSoutput.t48 gnd 0.053798f
C2062 CSoutput.n363 gnd 0.475374f
C2063 CSoutput.n364 gnd 0.218358f
C2064 CSoutput.t16 gnd 0.053798f
C2065 CSoutput.t190 gnd 0.053798f
C2066 CSoutput.n365 gnd 0.475374f
C2067 CSoutput.n366 gnd 0.218358f
C2068 CSoutput.t6 gnd 0.053798f
C2069 CSoutput.t189 gnd 0.053798f
C2070 CSoutput.n367 gnd 0.475374f
C2071 CSoutput.n368 gnd 0.218358f
C2072 CSoutput.t27 gnd 0.053798f
C2073 CSoutput.t3 gnd 0.053798f
C2074 CSoutput.n369 gnd 0.475374f
C2075 CSoutput.n370 gnd 0.331515f
C2076 CSoutput.n371 gnd 0.418143f
C2077 CSoutput.t50 gnd 0.053798f
C2078 CSoutput.t23 gnd 0.053798f
C2079 CSoutput.n372 gnd 0.476965f
C2080 CSoutput.t36 gnd 0.053798f
C2081 CSoutput.t62 gnd 0.053798f
C2082 CSoutput.n373 gnd 0.475374f
C2083 CSoutput.n374 gnd 0.44296f
C2084 CSoutput.t59 gnd 0.053798f
C2085 CSoutput.t35 gnd 0.053798f
C2086 CSoutput.n375 gnd 0.475374f
C2087 CSoutput.n376 gnd 0.218358f
C2088 CSoutput.t47 gnd 0.053798f
C2089 CSoutput.t49 gnd 0.053798f
C2090 CSoutput.n377 gnd 0.475374f
C2091 CSoutput.n378 gnd 0.218358f
C2092 CSoutput.t43 gnd 0.053798f
C2093 CSoutput.t186 gnd 0.053798f
C2094 CSoutput.n379 gnd 0.475374f
C2095 CSoutput.n380 gnd 0.218358f
C2096 CSoutput.t42 gnd 0.053798f
C2097 CSoutput.t38 gnd 0.053798f
C2098 CSoutput.n381 gnd 0.475374f
C2099 CSoutput.n382 gnd 0.331515f
C2100 CSoutput.n383 gnd 0.44902f
C2101 CSoutput.n384 gnd 12.6005f
C2102 CSoutput.t39 gnd 0.053798f
C2103 CSoutput.t183 gnd 0.053798f
C2104 CSoutput.n385 gnd 0.476965f
C2105 CSoutput.t11 gnd 0.053798f
C2106 CSoutput.t7 gnd 0.053798f
C2107 CSoutput.n386 gnd 0.475374f
C2108 CSoutput.n387 gnd 0.44296f
C2109 CSoutput.t34 gnd 0.053798f
C2110 CSoutput.t61 gnd 0.053798f
C2111 CSoutput.n388 gnd 0.475374f
C2112 CSoutput.n389 gnd 0.218358f
C2113 CSoutput.t17 gnd 0.053798f
C2114 CSoutput.t52 gnd 0.053798f
C2115 CSoutput.n390 gnd 0.475374f
C2116 CSoutput.n391 gnd 0.218358f
C2117 CSoutput.t44 gnd 0.053798f
C2118 CSoutput.t20 gnd 0.053798f
C2119 CSoutput.n392 gnd 0.475374f
C2120 CSoutput.n393 gnd 0.218358f
C2121 CSoutput.t57 gnd 0.053798f
C2122 CSoutput.t19 gnd 0.053798f
C2123 CSoutput.n394 gnd 0.475374f
C2124 CSoutput.n395 gnd 0.40275f
C2125 CSoutput.t10 gnd 0.053798f
C2126 CSoutput.t30 gnd 0.053798f
C2127 CSoutput.n396 gnd 0.476965f
C2128 CSoutput.t58 gnd 0.053798f
C2129 CSoutput.t60 gnd 0.053798f
C2130 CSoutput.n397 gnd 0.475374f
C2131 CSoutput.n398 gnd 0.44296f
C2132 CSoutput.t32 gnd 0.053798f
C2133 CSoutput.t9 gnd 0.053798f
C2134 CSoutput.n399 gnd 0.475374f
C2135 CSoutput.n400 gnd 0.218358f
C2136 CSoutput.t45 gnd 0.053798f
C2137 CSoutput.t26 gnd 0.053798f
C2138 CSoutput.n401 gnd 0.475374f
C2139 CSoutput.n402 gnd 0.218358f
C2140 CSoutput.t4 gnd 0.053798f
C2141 CSoutput.t12 gnd 0.053798f
C2142 CSoutput.n403 gnd 0.475374f
C2143 CSoutput.n404 gnd 0.218358f
C2144 CSoutput.t22 gnd 0.053798f
C2145 CSoutput.t2 gnd 0.053798f
C2146 CSoutput.n405 gnd 0.475374f
C2147 CSoutput.n406 gnd 0.331515f
C2148 CSoutput.n407 gnd 0.418143f
C2149 CSoutput.t18 gnd 0.053798f
C2150 CSoutput.t1 gnd 0.053798f
C2151 CSoutput.n408 gnd 0.476965f
C2152 CSoutput.t40 gnd 0.053798f
C2153 CSoutput.t184 gnd 0.053798f
C2154 CSoutput.n409 gnd 0.475374f
C2155 CSoutput.n410 gnd 0.44296f
C2156 CSoutput.t53 gnd 0.053798f
C2157 CSoutput.t25 gnd 0.053798f
C2158 CSoutput.n411 gnd 0.475374f
C2159 CSoutput.n412 gnd 0.218358f
C2160 CSoutput.t14 gnd 0.053798f
C2161 CSoutput.t46 gnd 0.053798f
C2162 CSoutput.n413 gnd 0.475374f
C2163 CSoutput.n414 gnd 0.218358f
C2164 CSoutput.t0 gnd 0.053798f
C2165 CSoutput.t188 gnd 0.053798f
C2166 CSoutput.n415 gnd 0.475374f
C2167 CSoutput.n416 gnd 0.218358f
C2168 CSoutput.t31 gnd 0.053798f
C2169 CSoutput.t37 gnd 0.053798f
C2170 CSoutput.n417 gnd 0.475374f
C2171 CSoutput.n418 gnd 0.331515f
C2172 CSoutput.n419 gnd 0.44902f
C2173 CSoutput.n420 gnd 7.08929f
C2174 CSoutput.n421 gnd 14.807901f
C2175 vdd.t3 gnd 0.039464f
C2176 vdd.t42 gnd 0.039464f
C2177 vdd.n0 gnd 0.311261f
C2178 vdd.t26 gnd 0.039464f
C2179 vdd.t34 gnd 0.039464f
C2180 vdd.n1 gnd 0.310748f
C2181 vdd.n2 gnd 0.286569f
C2182 vdd.t24 gnd 0.039464f
C2183 vdd.t16 gnd 0.039464f
C2184 vdd.n3 gnd 0.310748f
C2185 vdd.n4 gnd 0.144928f
C2186 vdd.t18 gnd 0.039464f
C2187 vdd.t11 gnd 0.039464f
C2188 vdd.n5 gnd 0.310748f
C2189 vdd.n6 gnd 0.135989f
C2190 vdd.t50 gnd 0.039464f
C2191 vdd.t31 gnd 0.039464f
C2192 vdd.n7 gnd 0.311261f
C2193 vdd.t13 gnd 0.039464f
C2194 vdd.t1 gnd 0.039464f
C2195 vdd.n8 gnd 0.310748f
C2196 vdd.n9 gnd 0.286569f
C2197 vdd.t36 gnd 0.039464f
C2198 vdd.t29 gnd 0.039464f
C2199 vdd.n10 gnd 0.310748f
C2200 vdd.n11 gnd 0.144928f
C2201 vdd.t47 gnd 0.039464f
C2202 vdd.t223 gnd 0.039464f
C2203 vdd.n12 gnd 0.310748f
C2204 vdd.n13 gnd 0.135989f
C2205 vdd.n14 gnd 0.096141f
C2206 vdd.t53 gnd 0.021925f
C2207 vdd.t57 gnd 0.021925f
C2208 vdd.n15 gnd 0.201807f
C2209 vdd.t5 gnd 0.021925f
C2210 vdd.t55 gnd 0.021925f
C2211 vdd.n16 gnd 0.201216f
C2212 vdd.n17 gnd 0.350179f
C2213 vdd.t61 gnd 0.021925f
C2214 vdd.t38 gnd 0.021925f
C2215 vdd.n18 gnd 0.201216f
C2216 vdd.n19 gnd 0.144874f
C2217 vdd.t6 gnd 0.021925f
C2218 vdd.t58 gnd 0.021925f
C2219 vdd.n20 gnd 0.201807f
C2220 vdd.t60 gnd 0.021925f
C2221 vdd.t52 gnd 0.021925f
C2222 vdd.n21 gnd 0.201216f
C2223 vdd.n22 gnd 0.350179f
C2224 vdd.t37 gnd 0.021925f
C2225 vdd.t54 gnd 0.021925f
C2226 vdd.n23 gnd 0.201216f
C2227 vdd.n24 gnd 0.144874f
C2228 vdd.t56 gnd 0.021925f
C2229 vdd.t39 gnd 0.021925f
C2230 vdd.n25 gnd 0.201216f
C2231 vdd.t40 gnd 0.021925f
C2232 vdd.t4 gnd 0.021925f
C2233 vdd.n26 gnd 0.201216f
C2234 vdd.n27 gnd 21.8196f
C2235 vdd.n28 gnd 8.389179f
C2236 vdd.n29 gnd 0.00598f
C2237 vdd.n30 gnd 0.005549f
C2238 vdd.n31 gnd 0.003069f
C2239 vdd.n32 gnd 0.007048f
C2240 vdd.n33 gnd 0.002982f
C2241 vdd.n34 gnd 0.003157f
C2242 vdd.n35 gnd 0.005549f
C2243 vdd.n36 gnd 0.002982f
C2244 vdd.n37 gnd 0.007048f
C2245 vdd.n38 gnd 0.003157f
C2246 vdd.n39 gnd 0.005549f
C2247 vdd.n40 gnd 0.002982f
C2248 vdd.n41 gnd 0.005286f
C2249 vdd.n42 gnd 0.005302f
C2250 vdd.t113 gnd 0.015142f
C2251 vdd.n43 gnd 0.03369f
C2252 vdd.n44 gnd 0.175329f
C2253 vdd.n45 gnd 0.002982f
C2254 vdd.n46 gnd 0.003157f
C2255 vdd.n47 gnd 0.007048f
C2256 vdd.n48 gnd 0.007048f
C2257 vdd.n49 gnd 0.003157f
C2258 vdd.n50 gnd 0.002982f
C2259 vdd.n51 gnd 0.005549f
C2260 vdd.n52 gnd 0.005549f
C2261 vdd.n53 gnd 0.002982f
C2262 vdd.n54 gnd 0.003157f
C2263 vdd.n55 gnd 0.007048f
C2264 vdd.n56 gnd 0.007048f
C2265 vdd.n57 gnd 0.003157f
C2266 vdd.n58 gnd 0.002982f
C2267 vdd.n59 gnd 0.005549f
C2268 vdd.n60 gnd 0.005549f
C2269 vdd.n61 gnd 0.002982f
C2270 vdd.n62 gnd 0.003157f
C2271 vdd.n63 gnd 0.007048f
C2272 vdd.n64 gnd 0.007048f
C2273 vdd.n65 gnd 0.016662f
C2274 vdd.n66 gnd 0.003069f
C2275 vdd.n67 gnd 0.002982f
C2276 vdd.n68 gnd 0.014342f
C2277 vdd.n69 gnd 0.010013f
C2278 vdd.t199 gnd 0.035079f
C2279 vdd.t141 gnd 0.035079f
C2280 vdd.n70 gnd 0.24109f
C2281 vdd.n71 gnd 0.18958f
C2282 vdd.t213 gnd 0.035079f
C2283 vdd.t194 gnd 0.035079f
C2284 vdd.n72 gnd 0.24109f
C2285 vdd.n73 gnd 0.15299f
C2286 vdd.t79 gnd 0.035079f
C2287 vdd.t128 gnd 0.035079f
C2288 vdd.n74 gnd 0.24109f
C2289 vdd.n75 gnd 0.15299f
C2290 vdd.t92 gnd 0.035079f
C2291 vdd.t154 gnd 0.035079f
C2292 vdd.n76 gnd 0.24109f
C2293 vdd.n77 gnd 0.15299f
C2294 vdd.t119 gnd 0.035079f
C2295 vdd.t203 gnd 0.035079f
C2296 vdd.n78 gnd 0.24109f
C2297 vdd.n79 gnd 0.15299f
C2298 vdd.t98 gnd 0.035079f
C2299 vdd.t176 gnd 0.035079f
C2300 vdd.n80 gnd 0.24109f
C2301 vdd.n81 gnd 0.15299f
C2302 vdd.t103 gnd 0.035079f
C2303 vdd.t190 gnd 0.035079f
C2304 vdd.n82 gnd 0.24109f
C2305 vdd.n83 gnd 0.15299f
C2306 vdd.t136 gnd 0.035079f
C2307 vdd.t208 gnd 0.035079f
C2308 vdd.n84 gnd 0.24109f
C2309 vdd.n85 gnd 0.15299f
C2310 vdd.t157 gnd 0.035079f
C2311 vdd.t186 gnd 0.035079f
C2312 vdd.n86 gnd 0.24109f
C2313 vdd.n87 gnd 0.15299f
C2314 vdd.n88 gnd 0.00598f
C2315 vdd.n89 gnd 0.005549f
C2316 vdd.n90 gnd 0.003069f
C2317 vdd.n91 gnd 0.007048f
C2318 vdd.n92 gnd 0.002982f
C2319 vdd.n93 gnd 0.003157f
C2320 vdd.n94 gnd 0.005549f
C2321 vdd.n95 gnd 0.002982f
C2322 vdd.n96 gnd 0.007048f
C2323 vdd.n97 gnd 0.003157f
C2324 vdd.n98 gnd 0.005549f
C2325 vdd.n99 gnd 0.002982f
C2326 vdd.n100 gnd 0.005286f
C2327 vdd.n101 gnd 0.005302f
C2328 vdd.t120 gnd 0.015142f
C2329 vdd.n102 gnd 0.03369f
C2330 vdd.n103 gnd 0.175329f
C2331 vdd.n104 gnd 0.002982f
C2332 vdd.n105 gnd 0.003157f
C2333 vdd.n106 gnd 0.007048f
C2334 vdd.n107 gnd 0.007048f
C2335 vdd.n108 gnd 0.003157f
C2336 vdd.n109 gnd 0.002982f
C2337 vdd.n110 gnd 0.005549f
C2338 vdd.n111 gnd 0.005549f
C2339 vdd.n112 gnd 0.002982f
C2340 vdd.n113 gnd 0.003157f
C2341 vdd.n114 gnd 0.007048f
C2342 vdd.n115 gnd 0.007048f
C2343 vdd.n116 gnd 0.003157f
C2344 vdd.n117 gnd 0.002982f
C2345 vdd.n118 gnd 0.005549f
C2346 vdd.n119 gnd 0.005549f
C2347 vdd.n120 gnd 0.002982f
C2348 vdd.n121 gnd 0.003157f
C2349 vdd.n122 gnd 0.007048f
C2350 vdd.n123 gnd 0.007048f
C2351 vdd.n124 gnd 0.016662f
C2352 vdd.n125 gnd 0.003069f
C2353 vdd.n126 gnd 0.002982f
C2354 vdd.n127 gnd 0.014342f
C2355 vdd.n128 gnd 0.009699f
C2356 vdd.n129 gnd 0.113825f
C2357 vdd.n130 gnd 0.00598f
C2358 vdd.n131 gnd 0.005549f
C2359 vdd.n132 gnd 0.003069f
C2360 vdd.n133 gnd 0.007048f
C2361 vdd.n134 gnd 0.002982f
C2362 vdd.n135 gnd 0.003157f
C2363 vdd.n136 gnd 0.005549f
C2364 vdd.n137 gnd 0.002982f
C2365 vdd.n138 gnd 0.007048f
C2366 vdd.n139 gnd 0.003157f
C2367 vdd.n140 gnd 0.005549f
C2368 vdd.n141 gnd 0.002982f
C2369 vdd.n142 gnd 0.005286f
C2370 vdd.n143 gnd 0.005302f
C2371 vdd.t152 gnd 0.015142f
C2372 vdd.n144 gnd 0.03369f
C2373 vdd.n145 gnd 0.175329f
C2374 vdd.n146 gnd 0.002982f
C2375 vdd.n147 gnd 0.003157f
C2376 vdd.n148 gnd 0.007048f
C2377 vdd.n149 gnd 0.007048f
C2378 vdd.n150 gnd 0.003157f
C2379 vdd.n151 gnd 0.002982f
C2380 vdd.n152 gnd 0.005549f
C2381 vdd.n153 gnd 0.005549f
C2382 vdd.n154 gnd 0.002982f
C2383 vdd.n155 gnd 0.003157f
C2384 vdd.n156 gnd 0.007048f
C2385 vdd.n157 gnd 0.007048f
C2386 vdd.n158 gnd 0.003157f
C2387 vdd.n159 gnd 0.002982f
C2388 vdd.n160 gnd 0.005549f
C2389 vdd.n161 gnd 0.005549f
C2390 vdd.n162 gnd 0.002982f
C2391 vdd.n163 gnd 0.003157f
C2392 vdd.n164 gnd 0.007048f
C2393 vdd.n165 gnd 0.007048f
C2394 vdd.n166 gnd 0.016662f
C2395 vdd.n167 gnd 0.003069f
C2396 vdd.n168 gnd 0.002982f
C2397 vdd.n169 gnd 0.014342f
C2398 vdd.n170 gnd 0.010013f
C2399 vdd.t185 gnd 0.035079f
C2400 vdd.t67 gnd 0.035079f
C2401 vdd.n171 gnd 0.24109f
C2402 vdd.n172 gnd 0.18958f
C2403 vdd.t125 gnd 0.035079f
C2404 vdd.t127 gnd 0.035079f
C2405 vdd.n173 gnd 0.24109f
C2406 vdd.n174 gnd 0.15299f
C2407 vdd.t207 gnd 0.035079f
C2408 vdd.t75 gnd 0.035079f
C2409 vdd.n175 gnd 0.24109f
C2410 vdd.n176 gnd 0.15299f
C2411 vdd.t117 gnd 0.035079f
C2412 vdd.t205 gnd 0.035079f
C2413 vdd.n177 gnd 0.24109f
C2414 vdd.n178 gnd 0.15299f
C2415 vdd.t206 gnd 0.035079f
C2416 vdd.t90 gnd 0.035079f
C2417 vdd.n179 gnd 0.24109f
C2418 vdd.n180 gnd 0.15299f
C2419 vdd.t188 gnd 0.035079f
C2420 vdd.t202 gnd 0.035079f
C2421 vdd.n181 gnd 0.24109f
C2422 vdd.n182 gnd 0.15299f
C2423 vdd.t86 gnd 0.035079f
C2424 vdd.t151 gnd 0.035079f
C2425 vdd.n183 gnd 0.24109f
C2426 vdd.n184 gnd 0.15299f
C2427 vdd.t183 gnd 0.035079f
C2428 vdd.t214 gnd 0.035079f
C2429 vdd.n185 gnd 0.24109f
C2430 vdd.n186 gnd 0.15299f
C2431 vdd.t123 gnd 0.035079f
C2432 vdd.t182 gnd 0.035079f
C2433 vdd.n187 gnd 0.24109f
C2434 vdd.n188 gnd 0.15299f
C2435 vdd.n189 gnd 0.00598f
C2436 vdd.n190 gnd 0.005549f
C2437 vdd.n191 gnd 0.003069f
C2438 vdd.n192 gnd 0.007048f
C2439 vdd.n193 gnd 0.002982f
C2440 vdd.n194 gnd 0.003157f
C2441 vdd.n195 gnd 0.005549f
C2442 vdd.n196 gnd 0.002982f
C2443 vdd.n197 gnd 0.007048f
C2444 vdd.n198 gnd 0.003157f
C2445 vdd.n199 gnd 0.005549f
C2446 vdd.n200 gnd 0.002982f
C2447 vdd.n201 gnd 0.005286f
C2448 vdd.n202 gnd 0.005302f
C2449 vdd.t219 gnd 0.015142f
C2450 vdd.n203 gnd 0.03369f
C2451 vdd.n204 gnd 0.175329f
C2452 vdd.n205 gnd 0.002982f
C2453 vdd.n206 gnd 0.003157f
C2454 vdd.n207 gnd 0.007048f
C2455 vdd.n208 gnd 0.007048f
C2456 vdd.n209 gnd 0.003157f
C2457 vdd.n210 gnd 0.002982f
C2458 vdd.n211 gnd 0.005549f
C2459 vdd.n212 gnd 0.005549f
C2460 vdd.n213 gnd 0.002982f
C2461 vdd.n214 gnd 0.003157f
C2462 vdd.n215 gnd 0.007048f
C2463 vdd.n216 gnd 0.007048f
C2464 vdd.n217 gnd 0.003157f
C2465 vdd.n218 gnd 0.002982f
C2466 vdd.n219 gnd 0.005549f
C2467 vdd.n220 gnd 0.005549f
C2468 vdd.n221 gnd 0.002982f
C2469 vdd.n222 gnd 0.003157f
C2470 vdd.n223 gnd 0.007048f
C2471 vdd.n224 gnd 0.007048f
C2472 vdd.n225 gnd 0.016662f
C2473 vdd.n226 gnd 0.003069f
C2474 vdd.n227 gnd 0.002982f
C2475 vdd.n228 gnd 0.014342f
C2476 vdd.n229 gnd 0.009699f
C2477 vdd.n230 gnd 0.067715f
C2478 vdd.n231 gnd 0.243994f
C2479 vdd.n232 gnd 0.00598f
C2480 vdd.n233 gnd 0.005549f
C2481 vdd.n234 gnd 0.003069f
C2482 vdd.n235 gnd 0.007048f
C2483 vdd.n236 gnd 0.002982f
C2484 vdd.n237 gnd 0.003157f
C2485 vdd.n238 gnd 0.005549f
C2486 vdd.n239 gnd 0.002982f
C2487 vdd.n240 gnd 0.007048f
C2488 vdd.n241 gnd 0.003157f
C2489 vdd.n242 gnd 0.005549f
C2490 vdd.n243 gnd 0.002982f
C2491 vdd.n244 gnd 0.005286f
C2492 vdd.n245 gnd 0.005302f
C2493 vdd.t168 gnd 0.015142f
C2494 vdd.n246 gnd 0.03369f
C2495 vdd.n247 gnd 0.175329f
C2496 vdd.n248 gnd 0.002982f
C2497 vdd.n249 gnd 0.003157f
C2498 vdd.n250 gnd 0.007048f
C2499 vdd.n251 gnd 0.007048f
C2500 vdd.n252 gnd 0.003157f
C2501 vdd.n253 gnd 0.002982f
C2502 vdd.n254 gnd 0.005549f
C2503 vdd.n255 gnd 0.005549f
C2504 vdd.n256 gnd 0.002982f
C2505 vdd.n257 gnd 0.003157f
C2506 vdd.n258 gnd 0.007048f
C2507 vdd.n259 gnd 0.007048f
C2508 vdd.n260 gnd 0.003157f
C2509 vdd.n261 gnd 0.002982f
C2510 vdd.n262 gnd 0.005549f
C2511 vdd.n263 gnd 0.005549f
C2512 vdd.n264 gnd 0.002982f
C2513 vdd.n265 gnd 0.003157f
C2514 vdd.n266 gnd 0.007048f
C2515 vdd.n267 gnd 0.007048f
C2516 vdd.n268 gnd 0.016662f
C2517 vdd.n269 gnd 0.003069f
C2518 vdd.n270 gnd 0.002982f
C2519 vdd.n271 gnd 0.014342f
C2520 vdd.n272 gnd 0.010013f
C2521 vdd.t196 gnd 0.035079f
C2522 vdd.t96 gnd 0.035079f
C2523 vdd.n273 gnd 0.24109f
C2524 vdd.n274 gnd 0.18958f
C2525 vdd.t145 gnd 0.035079f
C2526 vdd.t148 gnd 0.035079f
C2527 vdd.n275 gnd 0.24109f
C2528 vdd.n276 gnd 0.15299f
C2529 vdd.t218 gnd 0.035079f
C2530 vdd.t139 gnd 0.035079f
C2531 vdd.n277 gnd 0.24109f
C2532 vdd.n278 gnd 0.15299f
C2533 vdd.t140 gnd 0.035079f
C2534 vdd.t216 gnd 0.035079f
C2535 vdd.n279 gnd 0.24109f
C2536 vdd.n280 gnd 0.15299f
C2537 vdd.t217 gnd 0.035079f
C2538 vdd.t111 gnd 0.035079f
C2539 vdd.n281 gnd 0.24109f
C2540 vdd.n282 gnd 0.15299f
C2541 vdd.t201 gnd 0.035079f
C2542 vdd.t212 gnd 0.035079f
C2543 vdd.n283 gnd 0.24109f
C2544 vdd.n284 gnd 0.15299f
C2545 vdd.t104 gnd 0.035079f
C2546 vdd.t169 gnd 0.035079f
C2547 vdd.n285 gnd 0.24109f
C2548 vdd.n286 gnd 0.15299f
C2549 vdd.t197 gnd 0.035079f
C2550 vdd.t71 gnd 0.035079f
C2551 vdd.n287 gnd 0.24109f
C2552 vdd.n288 gnd 0.15299f
C2553 vdd.t146 gnd 0.035079f
C2554 vdd.t195 gnd 0.035079f
C2555 vdd.n289 gnd 0.24109f
C2556 vdd.n290 gnd 0.15299f
C2557 vdd.n291 gnd 0.00598f
C2558 vdd.n292 gnd 0.005549f
C2559 vdd.n293 gnd 0.003069f
C2560 vdd.n294 gnd 0.007048f
C2561 vdd.n295 gnd 0.002982f
C2562 vdd.n296 gnd 0.003157f
C2563 vdd.n297 gnd 0.005549f
C2564 vdd.n298 gnd 0.002982f
C2565 vdd.n299 gnd 0.007048f
C2566 vdd.n300 gnd 0.003157f
C2567 vdd.n301 gnd 0.005549f
C2568 vdd.n302 gnd 0.002982f
C2569 vdd.n303 gnd 0.005286f
C2570 vdd.n304 gnd 0.005302f
C2571 vdd.t88 gnd 0.015142f
C2572 vdd.n305 gnd 0.03369f
C2573 vdd.n306 gnd 0.175329f
C2574 vdd.n307 gnd 0.002982f
C2575 vdd.n308 gnd 0.003157f
C2576 vdd.n309 gnd 0.007048f
C2577 vdd.n310 gnd 0.007048f
C2578 vdd.n311 gnd 0.003157f
C2579 vdd.n312 gnd 0.002982f
C2580 vdd.n313 gnd 0.005549f
C2581 vdd.n314 gnd 0.005549f
C2582 vdd.n315 gnd 0.002982f
C2583 vdd.n316 gnd 0.003157f
C2584 vdd.n317 gnd 0.007048f
C2585 vdd.n318 gnd 0.007048f
C2586 vdd.n319 gnd 0.003157f
C2587 vdd.n320 gnd 0.002982f
C2588 vdd.n321 gnd 0.005549f
C2589 vdd.n322 gnd 0.005549f
C2590 vdd.n323 gnd 0.002982f
C2591 vdd.n324 gnd 0.003157f
C2592 vdd.n325 gnd 0.007048f
C2593 vdd.n326 gnd 0.007048f
C2594 vdd.n327 gnd 0.016662f
C2595 vdd.n328 gnd 0.003069f
C2596 vdd.n329 gnd 0.002982f
C2597 vdd.n330 gnd 0.014342f
C2598 vdd.n331 gnd 0.009699f
C2599 vdd.n332 gnd 0.067715f
C2600 vdd.n333 gnd 0.27932f
C2601 vdd.n334 gnd 0.008374f
C2602 vdd.n335 gnd 0.010896f
C2603 vdd.n336 gnd 0.00877f
C2604 vdd.n337 gnd 0.00877f
C2605 vdd.n338 gnd 0.010896f
C2606 vdd.n339 gnd 0.010896f
C2607 vdd.n340 gnd 0.796156f
C2608 vdd.n341 gnd 0.010896f
C2609 vdd.n342 gnd 0.010896f
C2610 vdd.n343 gnd 0.010896f
C2611 vdd.n344 gnd 0.862966f
C2612 vdd.n345 gnd 0.010896f
C2613 vdd.n346 gnd 0.010896f
C2614 vdd.n347 gnd 0.010896f
C2615 vdd.n348 gnd 0.010896f
C2616 vdd.n349 gnd 0.00877f
C2617 vdd.n350 gnd 0.010896f
C2618 vdd.t175 gnd 0.556753f
C2619 vdd.n351 gnd 0.010896f
C2620 vdd.n352 gnd 0.010896f
C2621 vdd.n353 gnd 0.010896f
C2622 vdd.t150 gnd 0.556753f
C2623 vdd.n354 gnd 0.010896f
C2624 vdd.n355 gnd 0.010896f
C2625 vdd.n356 gnd 0.010896f
C2626 vdd.n357 gnd 0.010896f
C2627 vdd.n358 gnd 0.010896f
C2628 vdd.n359 gnd 0.00877f
C2629 vdd.n360 gnd 0.010896f
C2630 vdd.n361 gnd 0.62913f
C2631 vdd.n362 gnd 0.010896f
C2632 vdd.n363 gnd 0.010896f
C2633 vdd.n364 gnd 0.010896f
C2634 vdd.t70 gnd 0.556753f
C2635 vdd.n365 gnd 0.010896f
C2636 vdd.n366 gnd 0.010896f
C2637 vdd.n367 gnd 0.010896f
C2638 vdd.n368 gnd 0.010896f
C2639 vdd.n369 gnd 0.010896f
C2640 vdd.n370 gnd 0.00877f
C2641 vdd.n371 gnd 0.010896f
C2642 vdd.t122 gnd 0.556753f
C2643 vdd.n372 gnd 0.010896f
C2644 vdd.n373 gnd 0.010896f
C2645 vdd.n374 gnd 0.010896f
C2646 vdd.n375 gnd 0.651401f
C2647 vdd.n376 gnd 0.010896f
C2648 vdd.n377 gnd 0.010896f
C2649 vdd.n378 gnd 0.010896f
C2650 vdd.n379 gnd 0.010896f
C2651 vdd.n380 gnd 0.010896f
C2652 vdd.n381 gnd 0.00877f
C2653 vdd.n382 gnd 0.010896f
C2654 vdd.t87 gnd 0.556753f
C2655 vdd.n383 gnd 0.010896f
C2656 vdd.n384 gnd 0.010896f
C2657 vdd.n385 gnd 0.010896f
C2658 vdd.n386 gnd 0.56232f
C2659 vdd.n387 gnd 0.010896f
C2660 vdd.n388 gnd 0.010896f
C2661 vdd.n389 gnd 0.010896f
C2662 vdd.n390 gnd 0.010896f
C2663 vdd.n391 gnd 0.026358f
C2664 vdd.n392 gnd 0.026923f
C2665 vdd.t247 gnd 0.556753f
C2666 vdd.n393 gnd 0.026358f
C2667 vdd.n425 gnd 0.010896f
C2668 vdd.t259 gnd 0.134048f
C2669 vdd.t258 gnd 0.14326f
C2670 vdd.t257 gnd 0.175065f
C2671 vdd.n426 gnd 0.224408f
C2672 vdd.n427 gnd 0.18942f
C2673 vdd.n428 gnd 0.014383f
C2674 vdd.n429 gnd 0.010896f
C2675 vdd.n430 gnd 0.00877f
C2676 vdd.n431 gnd 0.010896f
C2677 vdd.n432 gnd 0.00877f
C2678 vdd.n433 gnd 0.010896f
C2679 vdd.n434 gnd 0.00877f
C2680 vdd.n435 gnd 0.010896f
C2681 vdd.n436 gnd 0.00877f
C2682 vdd.n437 gnd 0.010896f
C2683 vdd.n438 gnd 0.00877f
C2684 vdd.n439 gnd 0.010896f
C2685 vdd.t249 gnd 0.134048f
C2686 vdd.t248 gnd 0.14326f
C2687 vdd.t246 gnd 0.175065f
C2688 vdd.n440 gnd 0.224408f
C2689 vdd.n441 gnd 0.18942f
C2690 vdd.n442 gnd 0.00877f
C2691 vdd.n443 gnd 0.010896f
C2692 vdd.n444 gnd 0.00877f
C2693 vdd.n445 gnd 0.010896f
C2694 vdd.n446 gnd 0.00877f
C2695 vdd.n447 gnd 0.010896f
C2696 vdd.n448 gnd 0.00877f
C2697 vdd.n449 gnd 0.010896f
C2698 vdd.n450 gnd 0.00877f
C2699 vdd.n451 gnd 0.010896f
C2700 vdd.t266 gnd 0.134048f
C2701 vdd.t265 gnd 0.14326f
C2702 vdd.t264 gnd 0.175065f
C2703 vdd.n452 gnd 0.224408f
C2704 vdd.n453 gnd 0.18942f
C2705 vdd.n454 gnd 0.018768f
C2706 vdd.n455 gnd 0.010896f
C2707 vdd.n456 gnd 0.00877f
C2708 vdd.n457 gnd 0.010896f
C2709 vdd.n458 gnd 0.00877f
C2710 vdd.n459 gnd 0.010896f
C2711 vdd.n460 gnd 0.00877f
C2712 vdd.n461 gnd 0.010896f
C2713 vdd.n462 gnd 0.00877f
C2714 vdd.n463 gnd 0.010896f
C2715 vdd.n464 gnd 0.026923f
C2716 vdd.n465 gnd 0.007279f
C2717 vdd.n466 gnd 0.00877f
C2718 vdd.n467 gnd 0.010896f
C2719 vdd.n468 gnd 0.010896f
C2720 vdd.n469 gnd 0.00877f
C2721 vdd.n470 gnd 0.010896f
C2722 vdd.n471 gnd 0.010896f
C2723 vdd.n472 gnd 0.010896f
C2724 vdd.n473 gnd 0.010896f
C2725 vdd.n474 gnd 0.010896f
C2726 vdd.n475 gnd 0.00877f
C2727 vdd.n476 gnd 0.00877f
C2728 vdd.n477 gnd 0.010896f
C2729 vdd.n478 gnd 0.010896f
C2730 vdd.n479 gnd 0.00877f
C2731 vdd.n480 gnd 0.010896f
C2732 vdd.n481 gnd 0.010896f
C2733 vdd.n482 gnd 0.010896f
C2734 vdd.n483 gnd 0.010896f
C2735 vdd.n484 gnd 0.010896f
C2736 vdd.n485 gnd 0.00877f
C2737 vdd.n486 gnd 0.00877f
C2738 vdd.n487 gnd 0.010896f
C2739 vdd.n488 gnd 0.010896f
C2740 vdd.n489 gnd 0.00877f
C2741 vdd.n490 gnd 0.010896f
C2742 vdd.n491 gnd 0.010896f
C2743 vdd.n492 gnd 0.010896f
C2744 vdd.n493 gnd 0.010896f
C2745 vdd.n494 gnd 0.010896f
C2746 vdd.n495 gnd 0.00877f
C2747 vdd.n496 gnd 0.00877f
C2748 vdd.n497 gnd 0.010896f
C2749 vdd.n498 gnd 0.010896f
C2750 vdd.n499 gnd 0.00877f
C2751 vdd.n500 gnd 0.010896f
C2752 vdd.n501 gnd 0.010896f
C2753 vdd.n502 gnd 0.010896f
C2754 vdd.n503 gnd 0.010896f
C2755 vdd.n504 gnd 0.010896f
C2756 vdd.n505 gnd 0.00877f
C2757 vdd.n506 gnd 0.00877f
C2758 vdd.n507 gnd 0.010896f
C2759 vdd.n508 gnd 0.010896f
C2760 vdd.n509 gnd 0.007323f
C2761 vdd.n510 gnd 0.010896f
C2762 vdd.n511 gnd 0.010896f
C2763 vdd.n512 gnd 0.010896f
C2764 vdd.n513 gnd 0.010896f
C2765 vdd.n514 gnd 0.010896f
C2766 vdd.n515 gnd 0.007323f
C2767 vdd.n516 gnd 0.00877f
C2768 vdd.n517 gnd 0.010896f
C2769 vdd.n518 gnd 0.010896f
C2770 vdd.n519 gnd 0.00877f
C2771 vdd.n520 gnd 0.010896f
C2772 vdd.n521 gnd 0.010896f
C2773 vdd.n522 gnd 0.010896f
C2774 vdd.n523 gnd 0.010896f
C2775 vdd.n524 gnd 0.010896f
C2776 vdd.n525 gnd 0.00877f
C2777 vdd.n526 gnd 0.00877f
C2778 vdd.n527 gnd 0.010896f
C2779 vdd.n528 gnd 0.010896f
C2780 vdd.n529 gnd 0.00877f
C2781 vdd.n530 gnd 0.010896f
C2782 vdd.n531 gnd 0.010896f
C2783 vdd.n532 gnd 0.010896f
C2784 vdd.n533 gnd 0.010896f
C2785 vdd.n534 gnd 0.010896f
C2786 vdd.n535 gnd 0.00877f
C2787 vdd.n536 gnd 0.00877f
C2788 vdd.n537 gnd 0.010896f
C2789 vdd.n538 gnd 0.010896f
C2790 vdd.n539 gnd 0.00877f
C2791 vdd.n540 gnd 0.010896f
C2792 vdd.n541 gnd 0.010896f
C2793 vdd.n542 gnd 0.010896f
C2794 vdd.n543 gnd 0.010896f
C2795 vdd.n544 gnd 0.010896f
C2796 vdd.n545 gnd 0.00877f
C2797 vdd.n546 gnd 0.00877f
C2798 vdd.n547 gnd 0.010896f
C2799 vdd.n548 gnd 0.010896f
C2800 vdd.n549 gnd 0.00877f
C2801 vdd.n550 gnd 0.010896f
C2802 vdd.n551 gnd 0.010896f
C2803 vdd.n552 gnd 0.010896f
C2804 vdd.n553 gnd 0.010896f
C2805 vdd.n554 gnd 0.010896f
C2806 vdd.n555 gnd 0.00877f
C2807 vdd.n556 gnd 0.00877f
C2808 vdd.n557 gnd 0.010896f
C2809 vdd.n558 gnd 0.010896f
C2810 vdd.n559 gnd 0.00877f
C2811 vdd.n560 gnd 0.010896f
C2812 vdd.n561 gnd 0.010896f
C2813 vdd.n562 gnd 0.010896f
C2814 vdd.n563 gnd 0.010896f
C2815 vdd.n564 gnd 0.010896f
C2816 vdd.n565 gnd 0.005964f
C2817 vdd.n566 gnd 0.018768f
C2818 vdd.n567 gnd 0.010896f
C2819 vdd.n568 gnd 0.010896f
C2820 vdd.n569 gnd 0.008682f
C2821 vdd.n570 gnd 0.010896f
C2822 vdd.n571 gnd 0.010896f
C2823 vdd.n572 gnd 0.010896f
C2824 vdd.n573 gnd 0.010896f
C2825 vdd.n574 gnd 0.010896f
C2826 vdd.n575 gnd 0.00877f
C2827 vdd.n576 gnd 0.00877f
C2828 vdd.n577 gnd 0.010896f
C2829 vdd.n578 gnd 0.010896f
C2830 vdd.n579 gnd 0.00877f
C2831 vdd.n580 gnd 0.010896f
C2832 vdd.n581 gnd 0.010896f
C2833 vdd.n582 gnd 0.010896f
C2834 vdd.n583 gnd 0.010896f
C2835 vdd.n584 gnd 0.010896f
C2836 vdd.n585 gnd 0.00877f
C2837 vdd.n586 gnd 0.00877f
C2838 vdd.n587 gnd 0.010896f
C2839 vdd.n588 gnd 0.010896f
C2840 vdd.n589 gnd 0.00877f
C2841 vdd.n590 gnd 0.010896f
C2842 vdd.n591 gnd 0.010896f
C2843 vdd.n592 gnd 0.010896f
C2844 vdd.n593 gnd 0.010896f
C2845 vdd.n594 gnd 0.010896f
C2846 vdd.n595 gnd 0.00877f
C2847 vdd.n596 gnd 0.00877f
C2848 vdd.n597 gnd 0.010896f
C2849 vdd.n598 gnd 0.010896f
C2850 vdd.n599 gnd 0.00877f
C2851 vdd.n600 gnd 0.010896f
C2852 vdd.n601 gnd 0.010896f
C2853 vdd.n602 gnd 0.010896f
C2854 vdd.n603 gnd 0.010896f
C2855 vdd.n604 gnd 0.010896f
C2856 vdd.n605 gnd 0.00877f
C2857 vdd.n606 gnd 0.00877f
C2858 vdd.n607 gnd 0.010896f
C2859 vdd.n608 gnd 0.010896f
C2860 vdd.n609 gnd 0.00877f
C2861 vdd.n610 gnd 0.010896f
C2862 vdd.n611 gnd 0.010896f
C2863 vdd.n612 gnd 0.010896f
C2864 vdd.n613 gnd 0.010896f
C2865 vdd.n614 gnd 0.010896f
C2866 vdd.n615 gnd 0.00877f
C2867 vdd.n616 gnd 0.010896f
C2868 vdd.n617 gnd 0.00877f
C2869 vdd.n618 gnd 0.004604f
C2870 vdd.n619 gnd 0.010896f
C2871 vdd.n620 gnd 0.010896f
C2872 vdd.n621 gnd 0.00877f
C2873 vdd.n622 gnd 0.010896f
C2874 vdd.n623 gnd 0.00877f
C2875 vdd.n624 gnd 0.010896f
C2876 vdd.n625 gnd 0.00877f
C2877 vdd.n626 gnd 0.010896f
C2878 vdd.n627 gnd 0.00877f
C2879 vdd.n628 gnd 0.010896f
C2880 vdd.n629 gnd 0.00877f
C2881 vdd.n630 gnd 0.010896f
C2882 vdd.n631 gnd 0.00877f
C2883 vdd.n632 gnd 0.010896f
C2884 vdd.n633 gnd 0.60686f
C2885 vdd.t118 gnd 0.556753f
C2886 vdd.n634 gnd 0.010896f
C2887 vdd.n635 gnd 0.00877f
C2888 vdd.n636 gnd 0.010896f
C2889 vdd.n637 gnd 0.00877f
C2890 vdd.n638 gnd 0.010896f
C2891 vdd.t91 gnd 0.556753f
C2892 vdd.n639 gnd 0.010896f
C2893 vdd.n640 gnd 0.00877f
C2894 vdd.n641 gnd 0.010896f
C2895 vdd.n642 gnd 0.00877f
C2896 vdd.n643 gnd 0.010896f
C2897 vdd.t74 gnd 0.556753f
C2898 vdd.n644 gnd 0.695941f
C2899 vdd.n645 gnd 0.010896f
C2900 vdd.n646 gnd 0.00877f
C2901 vdd.n647 gnd 0.010896f
C2902 vdd.n648 gnd 0.00877f
C2903 vdd.n649 gnd 0.010896f
C2904 vdd.t78 gnd 0.556753f
C2905 vdd.n650 gnd 0.010896f
C2906 vdd.n651 gnd 0.00877f
C2907 vdd.n652 gnd 0.010896f
C2908 vdd.n653 gnd 0.00877f
C2909 vdd.n654 gnd 0.010896f
C2910 vdd.n655 gnd 0.773886f
C2911 vdd.n656 gnd 0.924209f
C2912 vdd.t126 gnd 0.556753f
C2913 vdd.n657 gnd 0.010896f
C2914 vdd.n658 gnd 0.00877f
C2915 vdd.n659 gnd 0.010896f
C2916 vdd.n660 gnd 0.00877f
C2917 vdd.n661 gnd 0.010896f
C2918 vdd.n662 gnd 0.58459f
C2919 vdd.n663 gnd 0.010896f
C2920 vdd.n664 gnd 0.00877f
C2921 vdd.n665 gnd 0.010896f
C2922 vdd.n666 gnd 0.00877f
C2923 vdd.n667 gnd 0.010896f
C2924 vdd.t184 gnd 0.556753f
C2925 vdd.t66 gnd 0.556753f
C2926 vdd.n668 gnd 0.010896f
C2927 vdd.n669 gnd 0.00877f
C2928 vdd.n670 gnd 0.010896f
C2929 vdd.n671 gnd 0.00877f
C2930 vdd.n672 gnd 0.010896f
C2931 vdd.t112 gnd 0.556753f
C2932 vdd.n673 gnd 0.010896f
C2933 vdd.n674 gnd 0.00877f
C2934 vdd.n675 gnd 0.010896f
C2935 vdd.n676 gnd 0.00877f
C2936 vdd.n677 gnd 0.010896f
C2937 vdd.n678 gnd 1.11351f
C2938 vdd.n679 gnd 0.907507f
C2939 vdd.n680 gnd 0.010896f
C2940 vdd.n681 gnd 0.00877f
C2941 vdd.n682 gnd 0.026358f
C2942 vdd.n683 gnd 0.007279f
C2943 vdd.n684 gnd 0.026358f
C2944 vdd.t233 gnd 0.556753f
C2945 vdd.n685 gnd 0.026358f
C2946 vdd.n686 gnd 0.007279f
C2947 vdd.n687 gnd 0.00937f
C2948 vdd.t234 gnd 0.134048f
C2949 vdd.t235 gnd 0.14326f
C2950 vdd.t232 gnd 0.175065f
C2951 vdd.n688 gnd 0.224408f
C2952 vdd.n689 gnd 0.188543f
C2953 vdd.n690 gnd 0.013506f
C2954 vdd.n691 gnd 0.010896f
C2955 vdd.n692 gnd 9.4982f
C2956 vdd.n723 gnd 1.53107f
C2957 vdd.n724 gnd 0.010896f
C2958 vdd.n725 gnd 0.010896f
C2959 vdd.n726 gnd 0.026923f
C2960 vdd.n727 gnd 0.00937f
C2961 vdd.n728 gnd 0.010896f
C2962 vdd.n729 gnd 0.00877f
C2963 vdd.n730 gnd 0.006973f
C2964 vdd.n731 gnd 0.025446f
C2965 vdd.n732 gnd 0.00877f
C2966 vdd.n733 gnd 0.010896f
C2967 vdd.n734 gnd 0.010896f
C2968 vdd.n735 gnd 0.010896f
C2969 vdd.n736 gnd 0.010896f
C2970 vdd.n737 gnd 0.010896f
C2971 vdd.n738 gnd 0.010896f
C2972 vdd.n739 gnd 0.010896f
C2973 vdd.n740 gnd 0.010896f
C2974 vdd.n741 gnd 0.010896f
C2975 vdd.n742 gnd 0.010896f
C2976 vdd.n743 gnd 0.010896f
C2977 vdd.n744 gnd 0.010896f
C2978 vdd.n745 gnd 0.010896f
C2979 vdd.n746 gnd 0.010896f
C2980 vdd.n747 gnd 0.007323f
C2981 vdd.n748 gnd 0.010896f
C2982 vdd.n749 gnd 0.010896f
C2983 vdd.n750 gnd 0.010896f
C2984 vdd.n751 gnd 0.010896f
C2985 vdd.n752 gnd 0.010896f
C2986 vdd.n753 gnd 0.010896f
C2987 vdd.n754 gnd 0.010896f
C2988 vdd.n755 gnd 0.010896f
C2989 vdd.n756 gnd 0.010896f
C2990 vdd.n757 gnd 0.010896f
C2991 vdd.n758 gnd 0.010896f
C2992 vdd.n759 gnd 0.010896f
C2993 vdd.n760 gnd 0.010896f
C2994 vdd.n761 gnd 0.010896f
C2995 vdd.n762 gnd 0.010896f
C2996 vdd.n763 gnd 0.010896f
C2997 vdd.n764 gnd 0.010896f
C2998 vdd.n765 gnd 0.010896f
C2999 vdd.n766 gnd 0.010896f
C3000 vdd.n767 gnd 0.008682f
C3001 vdd.t241 gnd 0.134048f
C3002 vdd.t242 gnd 0.14326f
C3003 vdd.t240 gnd 0.175065f
C3004 vdd.n768 gnd 0.224408f
C3005 vdd.n769 gnd 0.188543f
C3006 vdd.n770 gnd 0.010896f
C3007 vdd.n771 gnd 0.010896f
C3008 vdd.n772 gnd 0.010896f
C3009 vdd.n773 gnd 0.010896f
C3010 vdd.n774 gnd 0.010896f
C3011 vdd.n775 gnd 0.010896f
C3012 vdd.n776 gnd 0.010896f
C3013 vdd.n777 gnd 0.010896f
C3014 vdd.n778 gnd 0.010896f
C3015 vdd.n779 gnd 0.010896f
C3016 vdd.n780 gnd 0.010896f
C3017 vdd.n781 gnd 0.010896f
C3018 vdd.n782 gnd 0.010896f
C3019 vdd.n783 gnd 0.006973f
C3020 vdd.n785 gnd 0.007409f
C3021 vdd.n786 gnd 0.007409f
C3022 vdd.n787 gnd 0.007409f
C3023 vdd.n788 gnd 0.007409f
C3024 vdd.n789 gnd 0.007409f
C3025 vdd.n790 gnd 0.007409f
C3026 vdd.n792 gnd 0.007409f
C3027 vdd.n793 gnd 0.007409f
C3028 vdd.n795 gnd 0.007409f
C3029 vdd.n796 gnd 0.005393f
C3030 vdd.n798 gnd 0.007409f
C3031 vdd.t227 gnd 0.299404f
C3032 vdd.t226 gnd 0.306477f
C3033 vdd.t224 gnd 0.195462f
C3034 vdd.n799 gnd 0.105637f
C3035 vdd.n800 gnd 0.059921f
C3036 vdd.n801 gnd 0.010589f
C3037 vdd.n802 gnd 0.01715f
C3038 vdd.n804 gnd 0.007409f
C3039 vdd.n805 gnd 0.757183f
C3040 vdd.n806 gnd 0.01623f
C3041 vdd.n807 gnd 0.01623f
C3042 vdd.n808 gnd 0.007409f
C3043 vdd.n809 gnd 0.01733f
C3044 vdd.n810 gnd 0.007409f
C3045 vdd.n811 gnd 0.007409f
C3046 vdd.n812 gnd 0.007409f
C3047 vdd.n813 gnd 0.007409f
C3048 vdd.n814 gnd 0.007409f
C3049 vdd.n816 gnd 0.007409f
C3050 vdd.n817 gnd 0.007409f
C3051 vdd.n819 gnd 0.007409f
C3052 vdd.n820 gnd 0.007409f
C3053 vdd.n822 gnd 0.007409f
C3054 vdd.n823 gnd 0.007409f
C3055 vdd.n825 gnd 0.007409f
C3056 vdd.n826 gnd 0.007409f
C3057 vdd.n828 gnd 0.007409f
C3058 vdd.n829 gnd 0.007409f
C3059 vdd.n831 gnd 0.007409f
C3060 vdd.t299 gnd 0.299404f
C3061 vdd.t298 gnd 0.306477f
C3062 vdd.t297 gnd 0.195462f
C3063 vdd.n832 gnd 0.105637f
C3064 vdd.n833 gnd 0.059921f
C3065 vdd.n834 gnd 0.007409f
C3066 vdd.n836 gnd 0.007409f
C3067 vdd.n837 gnd 0.007409f
C3068 vdd.t225 gnd 0.378592f
C3069 vdd.n838 gnd 0.007409f
C3070 vdd.n839 gnd 0.007409f
C3071 vdd.n840 gnd 0.007409f
C3072 vdd.n841 gnd 0.007409f
C3073 vdd.n842 gnd 0.007409f
C3074 vdd.n843 gnd 0.757183f
C3075 vdd.n844 gnd 0.007409f
C3076 vdd.n845 gnd 0.007409f
C3077 vdd.n846 gnd 0.640265f
C3078 vdd.n847 gnd 0.007409f
C3079 vdd.n848 gnd 0.007409f
C3080 vdd.n849 gnd 0.007409f
C3081 vdd.n850 gnd 0.007409f
C3082 vdd.n851 gnd 0.740481f
C3083 vdd.n852 gnd 0.007409f
C3084 vdd.n853 gnd 0.007409f
C3085 vdd.n854 gnd 0.007409f
C3086 vdd.n855 gnd 0.007409f
C3087 vdd.n856 gnd 0.007409f
C3088 vdd.n857 gnd 0.757183f
C3089 vdd.n858 gnd 0.007409f
C3090 vdd.n859 gnd 0.007409f
C3091 vdd.t8 gnd 0.378592f
C3092 vdd.n860 gnd 0.007409f
C3093 vdd.n861 gnd 0.007409f
C3094 vdd.n862 gnd 0.007409f
C3095 vdd.t27 gnd 0.378592f
C3096 vdd.n863 gnd 0.007409f
C3097 vdd.n864 gnd 0.007409f
C3098 vdd.n865 gnd 0.007409f
C3099 vdd.n866 gnd 0.007409f
C3100 vdd.n867 gnd 0.007409f
C3101 vdd.t251 gnd 0.317349f
C3102 vdd.n868 gnd 0.007409f
C3103 vdd.n869 gnd 0.007409f
C3104 vdd.n870 gnd 0.60686f
C3105 vdd.n871 gnd 0.007409f
C3106 vdd.t252 gnd 0.306477f
C3107 vdd.t250 gnd 0.195462f
C3108 vdd.t253 gnd 0.306477f
C3109 vdd.n872 gnd 0.172253f
C3110 vdd.n873 gnd 0.007409f
C3111 vdd.n874 gnd 0.007409f
C3112 vdd.n875 gnd 0.484375f
C3113 vdd.n876 gnd 0.007409f
C3114 vdd.n877 gnd 0.007409f
C3115 vdd.t19 gnd 0.111351f
C3116 vdd.n878 gnd 0.439835f
C3117 vdd.n879 gnd 0.007409f
C3118 vdd.n880 gnd 0.007409f
C3119 vdd.n881 gnd 0.007409f
C3120 vdd.n882 gnd 0.651401f
C3121 vdd.n883 gnd 0.007409f
C3122 vdd.n884 gnd 0.007409f
C3123 vdd.t22 gnd 0.378592f
C3124 vdd.n885 gnd 0.007409f
C3125 vdd.n886 gnd 0.007409f
C3126 vdd.n887 gnd 0.007409f
C3127 vdd.t30 gnd 0.378592f
C3128 vdd.n888 gnd 0.007409f
C3129 vdd.n889 gnd 0.007409f
C3130 vdd.t44 gnd 0.378592f
C3131 vdd.n890 gnd 0.007409f
C3132 vdd.n891 gnd 0.007409f
C3133 vdd.n892 gnd 0.007409f
C3134 vdd.t51 gnd 0.300646f
C3135 vdd.n893 gnd 0.007409f
C3136 vdd.n894 gnd 0.007409f
C3137 vdd.n895 gnd 0.623563f
C3138 vdd.n896 gnd 0.007409f
C3139 vdd.n897 gnd 0.007409f
C3140 vdd.n898 gnd 0.007409f
C3141 vdd.t59 gnd 0.378592f
C3142 vdd.n899 gnd 0.007409f
C3143 vdd.n900 gnd 0.007409f
C3144 vdd.t49 gnd 0.317349f
C3145 vdd.n901 gnd 0.456537f
C3146 vdd.n902 gnd 0.007409f
C3147 vdd.n903 gnd 0.007409f
C3148 vdd.n904 gnd 0.007409f
C3149 vdd.n905 gnd 0.395294f
C3150 vdd.n906 gnd 0.007409f
C3151 vdd.n907 gnd 0.007409f
C3152 vdd.t0 gnd 0.378592f
C3153 vdd.n908 gnd 0.007409f
C3154 vdd.n909 gnd 0.007409f
C3155 vdd.n910 gnd 0.007409f
C3156 vdd.n911 gnd 0.757183f
C3157 vdd.n912 gnd 0.007409f
C3158 vdd.n913 gnd 0.007409f
C3159 vdd.t20 gnd 0.256106f
C3160 vdd.t12 gnd 0.361889f
C3161 vdd.n914 gnd 0.007409f
C3162 vdd.n915 gnd 0.007409f
C3163 vdd.n916 gnd 0.007409f
C3164 vdd.n917 gnd 0.567888f
C3165 vdd.n918 gnd 0.007409f
C3166 vdd.n919 gnd 0.007409f
C3167 vdd.n920 gnd 0.007409f
C3168 vdd.n921 gnd 0.007409f
C3169 vdd.n922 gnd 0.007409f
C3170 vdd.t275 gnd 0.378592f
C3171 vdd.n923 gnd 0.007409f
C3172 vdd.n924 gnd 0.007409f
C3173 vdd.t28 gnd 0.378592f
C3174 vdd.n925 gnd 0.007409f
C3175 vdd.n926 gnd 0.01623f
C3176 vdd.n927 gnd 0.01623f
C3177 vdd.n928 gnd 0.901939f
C3178 vdd.n929 gnd 0.007409f
C3179 vdd.n930 gnd 0.007409f
C3180 vdd.t35 gnd 0.378592f
C3181 vdd.n931 gnd 0.01623f
C3182 vdd.n932 gnd 0.007409f
C3183 vdd.n933 gnd 0.007409f
C3184 vdd.t17 gnd 0.690373f
C3185 vdd.n951 gnd 0.01733f
C3186 vdd.n969 gnd 0.01623f
C3187 vdd.n970 gnd 0.007409f
C3188 vdd.n971 gnd 0.01623f
C3189 vdd.t296 gnd 0.299404f
C3190 vdd.t295 gnd 0.306477f
C3191 vdd.t294 gnd 0.195462f
C3192 vdd.n972 gnd 0.105637f
C3193 vdd.n973 gnd 0.059921f
C3194 vdd.n974 gnd 0.01715f
C3195 vdd.n975 gnd 0.007409f
C3196 vdd.n976 gnd 0.400862f
C3197 vdd.n977 gnd 0.01623f
C3198 vdd.n978 gnd 0.007409f
C3199 vdd.n979 gnd 0.01733f
C3200 vdd.n980 gnd 0.007409f
C3201 vdd.t273 gnd 0.299404f
C3202 vdd.t272 gnd 0.306477f
C3203 vdd.t270 gnd 0.195462f
C3204 vdd.n981 gnd 0.105637f
C3205 vdd.n982 gnd 0.059921f
C3206 vdd.n983 gnd 0.010589f
C3207 vdd.n984 gnd 0.007409f
C3208 vdd.n985 gnd 0.007409f
C3209 vdd.t271 gnd 0.378592f
C3210 vdd.n986 gnd 0.007409f
C3211 vdd.t15 gnd 0.378592f
C3212 vdd.n987 gnd 0.007409f
C3213 vdd.n988 gnd 0.007409f
C3214 vdd.n989 gnd 0.007409f
C3215 vdd.n990 gnd 0.007409f
C3216 vdd.n991 gnd 0.007409f
C3217 vdd.n992 gnd 0.757183f
C3218 vdd.n993 gnd 0.007409f
C3219 vdd.n994 gnd 0.007409f
C3220 vdd.t23 gnd 0.378592f
C3221 vdd.n995 gnd 0.007409f
C3222 vdd.n996 gnd 0.007409f
C3223 vdd.n997 gnd 0.007409f
C3224 vdd.n998 gnd 0.007409f
C3225 vdd.n999 gnd 0.501077f
C3226 vdd.n1000 gnd 0.007409f
C3227 vdd.n1001 gnd 0.007409f
C3228 vdd.n1002 gnd 0.007409f
C3229 vdd.n1003 gnd 0.007409f
C3230 vdd.n1004 gnd 0.007409f
C3231 vdd.n1005 gnd 0.668103f
C3232 vdd.n1006 gnd 0.007409f
C3233 vdd.n1007 gnd 0.007409f
C3234 vdd.t33 gnd 0.361889f
C3235 vdd.t9 gnd 0.256106f
C3236 vdd.n1008 gnd 0.007409f
C3237 vdd.n1009 gnd 0.007409f
C3238 vdd.n1010 gnd 0.007409f
C3239 vdd.t43 gnd 0.378592f
C3240 vdd.n1011 gnd 0.007409f
C3241 vdd.n1012 gnd 0.007409f
C3242 vdd.t25 gnd 0.378592f
C3243 vdd.n1013 gnd 0.007409f
C3244 vdd.n1014 gnd 0.007409f
C3245 vdd.n1015 gnd 0.007409f
C3246 vdd.t41 gnd 0.317349f
C3247 vdd.n1016 gnd 0.007409f
C3248 vdd.n1017 gnd 0.007409f
C3249 vdd.n1018 gnd 0.60686f
C3250 vdd.n1019 gnd 0.007409f
C3251 vdd.n1020 gnd 0.007409f
C3252 vdd.n1021 gnd 0.007409f
C3253 vdd.t2 gnd 0.378592f
C3254 vdd.n1022 gnd 0.007409f
C3255 vdd.n1023 gnd 0.007409f
C3256 vdd.t7 gnd 0.300646f
C3257 vdd.n1024 gnd 0.439835f
C3258 vdd.n1025 gnd 0.007409f
C3259 vdd.n1026 gnd 0.007409f
C3260 vdd.n1027 gnd 0.007409f
C3261 vdd.n1028 gnd 0.651401f
C3262 vdd.n1029 gnd 0.007409f
C3263 vdd.n1030 gnd 0.007409f
C3264 vdd.t21 gnd 0.378592f
C3265 vdd.n1031 gnd 0.007409f
C3266 vdd.n1032 gnd 0.007409f
C3267 vdd.n1033 gnd 0.007409f
C3268 vdd.n1034 gnd 0.757183f
C3269 vdd.n1035 gnd 0.007409f
C3270 vdd.n1036 gnd 0.007409f
C3271 vdd.t14 gnd 0.378592f
C3272 vdd.n1037 gnd 0.007409f
C3273 vdd.n1038 gnd 0.007409f
C3274 vdd.n1039 gnd 0.007409f
C3275 vdd.t32 gnd 0.111351f
C3276 vdd.n1040 gnd 0.007409f
C3277 vdd.n1041 gnd 0.007409f
C3278 vdd.n1042 gnd 0.007409f
C3279 vdd.t283 gnd 0.306477f
C3280 vdd.t281 gnd 0.195462f
C3281 vdd.t284 gnd 0.306477f
C3282 vdd.n1043 gnd 0.172253f
C3283 vdd.n1044 gnd 0.007409f
C3284 vdd.n1045 gnd 0.007409f
C3285 vdd.t48 gnd 0.378592f
C3286 vdd.n1046 gnd 0.007409f
C3287 vdd.n1047 gnd 0.007409f
C3288 vdd.t282 gnd 0.317349f
C3289 vdd.n1048 gnd 0.645833f
C3290 vdd.n1049 gnd 0.007409f
C3291 vdd.n1050 gnd 0.007409f
C3292 vdd.n1051 gnd 0.007409f
C3293 vdd.n1052 gnd 0.395294f
C3294 vdd.n1053 gnd 0.007409f
C3295 vdd.n1054 gnd 0.007409f
C3296 vdd.n1055 gnd 0.528915f
C3297 vdd.n1056 gnd 0.007409f
C3298 vdd.n1057 gnd 0.007409f
C3299 vdd.n1058 gnd 0.007409f
C3300 vdd.n1059 gnd 0.757183f
C3301 vdd.n1060 gnd 0.007409f
C3302 vdd.n1061 gnd 0.007409f
C3303 vdd.t45 gnd 0.378592f
C3304 vdd.n1062 gnd 0.007409f
C3305 vdd.n1063 gnd 0.007409f
C3306 vdd.n1064 gnd 0.007409f
C3307 vdd.n1065 gnd 0.757183f
C3308 vdd.n1066 gnd 0.007409f
C3309 vdd.n1067 gnd 0.007409f
C3310 vdd.n1068 gnd 0.007409f
C3311 vdd.n1069 gnd 0.007409f
C3312 vdd.n1070 gnd 0.007409f
C3313 vdd.t229 gnd 0.378592f
C3314 vdd.n1071 gnd 0.007409f
C3315 vdd.n1072 gnd 0.007409f
C3316 vdd.n1073 gnd 0.007409f
C3317 vdd.n1074 gnd 0.01623f
C3318 vdd.n1075 gnd 0.01623f
C3319 vdd.n1076 gnd 1.06896f
C3320 vdd.n1077 gnd 0.007409f
C3321 vdd.n1078 gnd 0.007409f
C3322 vdd.n1079 gnd 0.49551f
C3323 vdd.n1080 gnd 0.01623f
C3324 vdd.n1081 gnd 0.007409f
C3325 vdd.n1082 gnd 0.007409f
C3326 vdd.n1083 gnd 9.899059f
C3327 vdd.n1116 gnd 0.01733f
C3328 vdd.n1117 gnd 0.007409f
C3329 vdd.n1118 gnd 0.007409f
C3330 vdd.n1119 gnd 0.007409f
C3331 vdd.n1120 gnd 0.006973f
C3332 vdd.n1123 gnd 0.026923f
C3333 vdd.n1124 gnd 0.007279f
C3334 vdd.n1125 gnd 0.00877f
C3335 vdd.n1127 gnd 0.010896f
C3336 vdd.n1128 gnd 0.010896f
C3337 vdd.n1129 gnd 0.00877f
C3338 vdd.n1131 gnd 0.010896f
C3339 vdd.n1132 gnd 0.010896f
C3340 vdd.n1133 gnd 0.010896f
C3341 vdd.n1134 gnd 0.010896f
C3342 vdd.n1135 gnd 0.010896f
C3343 vdd.n1136 gnd 0.00877f
C3344 vdd.n1138 gnd 0.010896f
C3345 vdd.n1139 gnd 0.010896f
C3346 vdd.n1140 gnd 0.010896f
C3347 vdd.n1141 gnd 0.010896f
C3348 vdd.n1142 gnd 0.010896f
C3349 vdd.n1143 gnd 0.00877f
C3350 vdd.n1145 gnd 0.010896f
C3351 vdd.n1146 gnd 0.010896f
C3352 vdd.n1147 gnd 0.010896f
C3353 vdd.n1148 gnd 0.010896f
C3354 vdd.n1149 gnd 0.007323f
C3355 vdd.t287 gnd 0.134048f
C3356 vdd.t286 gnd 0.14326f
C3357 vdd.t285 gnd 0.175065f
C3358 vdd.n1150 gnd 0.224408f
C3359 vdd.n1151 gnd 0.188543f
C3360 vdd.n1153 gnd 0.010896f
C3361 vdd.n1154 gnd 0.010896f
C3362 vdd.n1155 gnd 0.00877f
C3363 vdd.n1156 gnd 0.010896f
C3364 vdd.n1158 gnd 0.010896f
C3365 vdd.n1159 gnd 0.010896f
C3366 vdd.n1160 gnd 0.010896f
C3367 vdd.n1161 gnd 0.010896f
C3368 vdd.n1162 gnd 0.00877f
C3369 vdd.n1164 gnd 0.010896f
C3370 vdd.n1165 gnd 0.010896f
C3371 vdd.n1166 gnd 0.010896f
C3372 vdd.n1167 gnd 0.010896f
C3373 vdd.n1168 gnd 0.010896f
C3374 vdd.n1169 gnd 0.00877f
C3375 vdd.n1171 gnd 0.010896f
C3376 vdd.n1172 gnd 0.010896f
C3377 vdd.n1173 gnd 0.010896f
C3378 vdd.n1174 gnd 0.010896f
C3379 vdd.n1175 gnd 0.010896f
C3380 vdd.n1176 gnd 0.00877f
C3381 vdd.n1178 gnd 0.010896f
C3382 vdd.n1179 gnd 0.010896f
C3383 vdd.n1180 gnd 0.010896f
C3384 vdd.n1181 gnd 0.010896f
C3385 vdd.n1182 gnd 0.010896f
C3386 vdd.n1183 gnd 0.00877f
C3387 vdd.n1185 gnd 0.010896f
C3388 vdd.n1186 gnd 0.010896f
C3389 vdd.n1187 gnd 0.010896f
C3390 vdd.n1188 gnd 0.010896f
C3391 vdd.n1189 gnd 0.008682f
C3392 vdd.t269 gnd 0.134048f
C3393 vdd.t268 gnd 0.14326f
C3394 vdd.t267 gnd 0.175065f
C3395 vdd.n1190 gnd 0.224408f
C3396 vdd.n1191 gnd 0.188543f
C3397 vdd.n1193 gnd 0.010896f
C3398 vdd.n1194 gnd 0.010896f
C3399 vdd.n1195 gnd 0.00877f
C3400 vdd.n1196 gnd 0.010896f
C3401 vdd.n1198 gnd 0.010896f
C3402 vdd.n1199 gnd 0.010896f
C3403 vdd.n1200 gnd 0.010896f
C3404 vdd.n1201 gnd 0.010896f
C3405 vdd.n1202 gnd 0.00877f
C3406 vdd.n1204 gnd 0.010896f
C3407 vdd.n1205 gnd 0.010896f
C3408 vdd.n1206 gnd 0.010896f
C3409 vdd.n1207 gnd 0.010896f
C3410 vdd.n1208 gnd 0.010896f
C3411 vdd.n1209 gnd 0.00877f
C3412 vdd.n1211 gnd 0.010896f
C3413 vdd.n1212 gnd 0.010896f
C3414 vdd.n1213 gnd 0.010896f
C3415 vdd.n1214 gnd 0.010896f
C3416 vdd.n1215 gnd 0.010896f
C3417 vdd.n1216 gnd 0.00877f
C3418 vdd.n1218 gnd 0.010896f
C3419 vdd.n1219 gnd 0.010896f
C3420 vdd.n1220 gnd 0.006973f
C3421 vdd.n1221 gnd 0.00877f
C3422 vdd.n1222 gnd 0.007409f
C3423 vdd.n1223 gnd 0.007409f
C3424 vdd.n1224 gnd 0.007409f
C3425 vdd.n1225 gnd 0.007409f
C3426 vdd.n1226 gnd 0.007409f
C3427 vdd.n1227 gnd 0.007409f
C3428 vdd.n1228 gnd 0.007409f
C3429 vdd.n1229 gnd 0.007409f
C3430 vdd.n1230 gnd 0.007409f
C3431 vdd.n1231 gnd 0.007409f
C3432 vdd.n1232 gnd 0.007409f
C3433 vdd.n1233 gnd 0.007409f
C3434 vdd.n1234 gnd 0.007409f
C3435 vdd.n1235 gnd 0.007409f
C3436 vdd.n1236 gnd 0.007409f
C3437 vdd.n1237 gnd 0.007409f
C3438 vdd.n1238 gnd 0.007409f
C3439 vdd.n1239 gnd 0.007409f
C3440 vdd.n1240 gnd 0.007409f
C3441 vdd.n1241 gnd 0.007409f
C3442 vdd.n1242 gnd 0.007409f
C3443 vdd.n1243 gnd 0.007409f
C3444 vdd.n1244 gnd 0.007409f
C3445 vdd.n1245 gnd 0.007409f
C3446 vdd.n1246 gnd 0.007409f
C3447 vdd.n1247 gnd 0.007409f
C3448 vdd.n1248 gnd 0.007409f
C3449 vdd.n1249 gnd 0.007409f
C3450 vdd.n1250 gnd 0.007409f
C3451 vdd.n1251 gnd 0.007409f
C3452 vdd.n1252 gnd 0.007409f
C3453 vdd.t230 gnd 0.299404f
C3454 vdd.t231 gnd 0.306477f
C3455 vdd.t228 gnd 0.195462f
C3456 vdd.n1253 gnd 0.105637f
C3457 vdd.n1254 gnd 0.059921f
C3458 vdd.n1255 gnd 0.010589f
C3459 vdd.n1256 gnd 0.007409f
C3460 vdd.n1257 gnd 0.007409f
C3461 vdd.n1258 gnd 0.007409f
C3462 vdd.n1259 gnd 0.007409f
C3463 vdd.n1260 gnd 0.007409f
C3464 vdd.n1261 gnd 0.007409f
C3465 vdd.n1262 gnd 0.007409f
C3466 vdd.n1263 gnd 0.007409f
C3467 vdd.n1264 gnd 0.007409f
C3468 vdd.n1265 gnd 0.007409f
C3469 vdd.n1266 gnd 0.007409f
C3470 vdd.n1267 gnd 0.007409f
C3471 vdd.n1268 gnd 0.007409f
C3472 vdd.n1269 gnd 0.007409f
C3473 vdd.n1270 gnd 0.007409f
C3474 vdd.n1271 gnd 0.007409f
C3475 vdd.n1272 gnd 0.007409f
C3476 vdd.t244 gnd 0.299404f
C3477 vdd.t245 gnd 0.306477f
C3478 vdd.t243 gnd 0.195462f
C3479 vdd.n1273 gnd 0.105637f
C3480 vdd.n1274 gnd 0.059921f
C3481 vdd.n1275 gnd 0.007409f
C3482 vdd.n1276 gnd 0.007409f
C3483 vdd.n1277 gnd 0.007409f
C3484 vdd.n1278 gnd 0.007409f
C3485 vdd.n1279 gnd 0.007409f
C3486 vdd.n1280 gnd 0.007409f
C3487 vdd.n1281 gnd 0.007409f
C3488 vdd.n1282 gnd 0.007409f
C3489 vdd.n1283 gnd 0.007409f
C3490 vdd.n1284 gnd 0.007409f
C3491 vdd.n1285 gnd 0.007409f
C3492 vdd.n1286 gnd 0.007409f
C3493 vdd.n1287 gnd 0.007409f
C3494 vdd.n1288 gnd 0.007409f
C3495 vdd.n1289 gnd 0.007409f
C3496 vdd.n1290 gnd 0.007409f
C3497 vdd.n1291 gnd 0.007409f
C3498 vdd.n1292 gnd 0.007409f
C3499 vdd.n1293 gnd 0.007409f
C3500 vdd.n1294 gnd 0.007409f
C3501 vdd.n1295 gnd 0.007409f
C3502 vdd.n1296 gnd 0.007409f
C3503 vdd.n1297 gnd 0.007409f
C3504 vdd.n1298 gnd 0.007409f
C3505 vdd.n1299 gnd 0.007409f
C3506 vdd.n1300 gnd 0.007409f
C3507 vdd.n1301 gnd 0.005393f
C3508 vdd.n1302 gnd 0.010589f
C3509 vdd.n1303 gnd 0.00572f
C3510 vdd.n1304 gnd 0.007409f
C3511 vdd.n1305 gnd 0.007409f
C3512 vdd.n1306 gnd 0.007409f
C3513 vdd.n1307 gnd 0.01733f
C3514 vdd.n1308 gnd 0.01733f
C3515 vdd.n1309 gnd 0.01623f
C3516 vdd.n1310 gnd 0.01623f
C3517 vdd.n1311 gnd 0.007409f
C3518 vdd.n1312 gnd 0.007409f
C3519 vdd.n1313 gnd 0.007409f
C3520 vdd.n1314 gnd 0.007409f
C3521 vdd.n1315 gnd 0.007409f
C3522 vdd.n1316 gnd 0.007409f
C3523 vdd.n1317 gnd 0.007409f
C3524 vdd.n1318 gnd 0.007409f
C3525 vdd.n1319 gnd 0.007409f
C3526 vdd.n1320 gnd 0.007409f
C3527 vdd.n1321 gnd 0.007409f
C3528 vdd.n1322 gnd 0.007409f
C3529 vdd.n1323 gnd 0.007409f
C3530 vdd.n1324 gnd 0.007409f
C3531 vdd.n1325 gnd 0.007409f
C3532 vdd.n1326 gnd 0.007409f
C3533 vdd.n1327 gnd 0.007409f
C3534 vdd.n1328 gnd 0.007409f
C3535 vdd.n1329 gnd 0.007409f
C3536 vdd.n1330 gnd 0.007409f
C3537 vdd.n1331 gnd 0.007409f
C3538 vdd.n1332 gnd 0.007409f
C3539 vdd.n1333 gnd 0.007409f
C3540 vdd.n1334 gnd 0.007409f
C3541 vdd.n1335 gnd 0.007409f
C3542 vdd.n1336 gnd 0.007409f
C3543 vdd.n1337 gnd 0.007409f
C3544 vdd.n1338 gnd 0.45097f
C3545 vdd.n1339 gnd 0.007409f
C3546 vdd.n1340 gnd 0.007409f
C3547 vdd.n1341 gnd 0.007409f
C3548 vdd.n1342 gnd 0.007409f
C3549 vdd.n1343 gnd 0.007409f
C3550 vdd.n1344 gnd 0.007409f
C3551 vdd.n1345 gnd 0.007409f
C3552 vdd.n1346 gnd 0.007409f
C3553 vdd.n1347 gnd 0.007409f
C3554 vdd.n1348 gnd 0.007409f
C3555 vdd.n1349 gnd 0.007409f
C3556 vdd.n1350 gnd 0.007409f
C3557 vdd.n1351 gnd 0.007409f
C3558 vdd.n1352 gnd 0.007409f
C3559 vdd.n1353 gnd 0.007409f
C3560 vdd.n1354 gnd 0.007409f
C3561 vdd.n1355 gnd 0.007409f
C3562 vdd.n1356 gnd 0.007409f
C3563 vdd.n1357 gnd 0.007409f
C3564 vdd.n1358 gnd 0.007409f
C3565 vdd.n1359 gnd 0.239404f
C3566 vdd.n1360 gnd 0.007409f
C3567 vdd.n1361 gnd 0.007409f
C3568 vdd.n1362 gnd 0.007409f
C3569 vdd.n1363 gnd 0.007409f
C3570 vdd.n1364 gnd 0.007409f
C3571 vdd.n1365 gnd 0.007409f
C3572 vdd.n1366 gnd 0.007409f
C3573 vdd.n1367 gnd 0.007409f
C3574 vdd.n1368 gnd 0.007409f
C3575 vdd.n1369 gnd 0.007409f
C3576 vdd.n1370 gnd 0.007409f
C3577 vdd.n1371 gnd 0.007409f
C3578 vdd.n1372 gnd 0.007409f
C3579 vdd.n1373 gnd 0.007409f
C3580 vdd.n1374 gnd 0.007409f
C3581 vdd.n1375 gnd 0.007409f
C3582 vdd.n1376 gnd 0.007409f
C3583 vdd.n1377 gnd 0.007409f
C3584 vdd.n1378 gnd 0.007409f
C3585 vdd.n1379 gnd 0.007409f
C3586 vdd.n1380 gnd 0.007409f
C3587 vdd.n1381 gnd 0.007409f
C3588 vdd.n1382 gnd 0.007409f
C3589 vdd.n1383 gnd 0.007409f
C3590 vdd.n1384 gnd 0.007409f
C3591 vdd.n1385 gnd 0.007409f
C3592 vdd.n1386 gnd 0.007409f
C3593 vdd.n1387 gnd 0.01623f
C3594 vdd.n1388 gnd 0.01623f
C3595 vdd.n1389 gnd 0.01733f
C3596 vdd.n1390 gnd 0.007409f
C3597 vdd.n1391 gnd 0.007409f
C3598 vdd.n1392 gnd 0.00572f
C3599 vdd.n1393 gnd 0.007409f
C3600 vdd.n1394 gnd 0.007409f
C3601 vdd.n1395 gnd 0.005393f
C3602 vdd.n1396 gnd 0.007409f
C3603 vdd.n1397 gnd 0.007409f
C3604 vdd.n1398 gnd 0.007409f
C3605 vdd.n1399 gnd 0.007409f
C3606 vdd.n1400 gnd 0.007409f
C3607 vdd.n1401 gnd 0.007409f
C3608 vdd.n1402 gnd 0.007409f
C3609 vdd.n1403 gnd 0.007409f
C3610 vdd.n1404 gnd 0.007409f
C3611 vdd.n1405 gnd 0.007409f
C3612 vdd.n1406 gnd 0.007409f
C3613 vdd.n1407 gnd 0.007409f
C3614 vdd.n1408 gnd 0.007409f
C3615 vdd.n1409 gnd 0.007409f
C3616 vdd.n1410 gnd 0.007409f
C3617 vdd.n1411 gnd 0.007409f
C3618 vdd.n1412 gnd 0.007409f
C3619 vdd.n1413 gnd 0.007409f
C3620 vdd.n1414 gnd 0.007409f
C3621 vdd.n1415 gnd 0.007409f
C3622 vdd.n1416 gnd 0.007409f
C3623 vdd.n1417 gnd 0.007409f
C3624 vdd.n1418 gnd 0.007409f
C3625 vdd.n1419 gnd 0.007409f
C3626 vdd.n1420 gnd 0.007409f
C3627 vdd.n1421 gnd 0.007409f
C3628 vdd.n1422 gnd 0.029696f
C3629 vdd.n1424 gnd 0.026923f
C3630 vdd.n1425 gnd 0.00877f
C3631 vdd.n1427 gnd 0.010896f
C3632 vdd.n1428 gnd 0.00877f
C3633 vdd.n1429 gnd 0.010896f
C3634 vdd.n1431 gnd 0.010896f
C3635 vdd.n1432 gnd 0.010896f
C3636 vdd.n1434 gnd 0.010896f
C3637 vdd.n1435 gnd 0.007279f
C3638 vdd.t237 gnd 0.556753f
C3639 vdd.n1436 gnd 0.010896f
C3640 vdd.n1437 gnd 0.026923f
C3641 vdd.n1438 gnd 0.00877f
C3642 vdd.n1439 gnd 0.010896f
C3643 vdd.n1440 gnd 0.00877f
C3644 vdd.n1441 gnd 0.010896f
C3645 vdd.n1442 gnd 1.11351f
C3646 vdd.n1443 gnd 0.010896f
C3647 vdd.n1444 gnd 0.00877f
C3648 vdd.n1445 gnd 0.00877f
C3649 vdd.n1446 gnd 0.010896f
C3650 vdd.n1447 gnd 0.00877f
C3651 vdd.n1448 gnd 0.010896f
C3652 vdd.t114 gnd 0.556753f
C3653 vdd.n1449 gnd 0.010896f
C3654 vdd.n1450 gnd 0.00877f
C3655 vdd.n1451 gnd 0.010896f
C3656 vdd.n1452 gnd 0.00877f
C3657 vdd.n1453 gnd 0.010896f
C3658 vdd.t76 gnd 0.556753f
C3659 vdd.n1454 gnd 0.010896f
C3660 vdd.n1455 gnd 0.00877f
C3661 vdd.n1456 gnd 0.010896f
C3662 vdd.n1457 gnd 0.00877f
C3663 vdd.n1458 gnd 0.010896f
C3664 vdd.n1459 gnd 0.896372f
C3665 vdd.n1460 gnd 0.924209f
C3666 vdd.t142 gnd 0.556753f
C3667 vdd.n1461 gnd 0.010896f
C3668 vdd.n1462 gnd 0.00877f
C3669 vdd.n1463 gnd 0.010896f
C3670 vdd.n1464 gnd 0.00877f
C3671 vdd.n1465 gnd 0.010896f
C3672 vdd.n1466 gnd 0.707076f
C3673 vdd.n1467 gnd 0.010896f
C3674 vdd.n1468 gnd 0.00877f
C3675 vdd.n1469 gnd 0.010896f
C3676 vdd.n1470 gnd 0.00877f
C3677 vdd.n1471 gnd 0.010896f
C3678 vdd.t83 gnd 0.556753f
C3679 vdd.t165 gnd 0.556753f
C3680 vdd.n1472 gnd 0.010896f
C3681 vdd.n1473 gnd 0.00877f
C3682 vdd.n1474 gnd 0.010896f
C3683 vdd.n1475 gnd 0.00877f
C3684 vdd.n1476 gnd 0.010896f
C3685 vdd.t130 gnd 0.556753f
C3686 vdd.n1477 gnd 0.010896f
C3687 vdd.n1478 gnd 0.00877f
C3688 vdd.n1479 gnd 0.010896f
C3689 vdd.n1480 gnd 0.00877f
C3690 vdd.n1481 gnd 0.010896f
C3691 vdd.t94 gnd 0.556753f
C3692 vdd.n1482 gnd 0.785021f
C3693 vdd.n1483 gnd 0.010896f
C3694 vdd.n1484 gnd 0.00877f
C3695 vdd.n1485 gnd 0.010896f
C3696 vdd.n1486 gnd 0.00877f
C3697 vdd.n1487 gnd 0.010896f
C3698 vdd.n1488 gnd 0.874102f
C3699 vdd.n1489 gnd 0.010896f
C3700 vdd.n1490 gnd 0.00877f
C3701 vdd.n1491 gnd 0.010896f
C3702 vdd.n1492 gnd 0.00877f
C3703 vdd.n1493 gnd 0.010896f
C3704 vdd.n1494 gnd 0.684806f
C3705 vdd.t160 gnd 0.556753f
C3706 vdd.n1495 gnd 0.010896f
C3707 vdd.n1496 gnd 0.00877f
C3708 vdd.n1497 gnd 0.010896f
C3709 vdd.n1498 gnd 0.00877f
C3710 vdd.n1499 gnd 0.010896f
C3711 vdd.t64 gnd 0.556753f
C3712 vdd.n1500 gnd 0.010896f
C3713 vdd.n1501 gnd 0.00877f
C3714 vdd.n1502 gnd 0.010896f
C3715 vdd.n1503 gnd 0.00877f
C3716 vdd.n1504 gnd 0.010896f
C3717 vdd.t105 gnd 0.556753f
C3718 vdd.n1505 gnd 0.617995f
C3719 vdd.n1506 gnd 0.010896f
C3720 vdd.n1507 gnd 0.00877f
C3721 vdd.n1508 gnd 0.010896f
C3722 vdd.n1509 gnd 0.00877f
C3723 vdd.n1510 gnd 0.010896f
C3724 vdd.t107 gnd 0.556753f
C3725 vdd.n1511 gnd 0.010896f
C3726 vdd.n1512 gnd 0.00877f
C3727 vdd.n1513 gnd 0.010896f
C3728 vdd.n1514 gnd 0.00877f
C3729 vdd.n1515 gnd 0.010896f
C3730 vdd.n1516 gnd 0.851831f
C3731 vdd.n1517 gnd 0.924209f
C3732 vdd.t68 gnd 0.556753f
C3733 vdd.n1518 gnd 0.010896f
C3734 vdd.n1519 gnd 0.00877f
C3735 vdd.n1520 gnd 0.010896f
C3736 vdd.n1521 gnd 0.00877f
C3737 vdd.n1522 gnd 0.010896f
C3738 vdd.n1523 gnd 0.662536f
C3739 vdd.n1524 gnd 0.010896f
C3740 vdd.n1525 gnd 0.00877f
C3741 vdd.n1526 gnd 0.010896f
C3742 vdd.n1527 gnd 0.00877f
C3743 vdd.n1528 gnd 0.010896f
C3744 vdd.t158 gnd 0.556753f
C3745 vdd.t132 gnd 0.556753f
C3746 vdd.n1529 gnd 0.010896f
C3747 vdd.n1530 gnd 0.00877f
C3748 vdd.n1531 gnd 0.010896f
C3749 vdd.n1532 gnd 0.00877f
C3750 vdd.n1533 gnd 0.010896f
C3751 vdd.t62 gnd 0.556753f
C3752 vdd.n1534 gnd 0.010896f
C3753 vdd.n1535 gnd 0.00877f
C3754 vdd.n1536 gnd 0.010896f
C3755 vdd.n1537 gnd 0.00877f
C3756 vdd.n1538 gnd 0.010896f
C3757 vdd.t72 gnd 0.556753f
C3758 vdd.n1539 gnd 0.829561f
C3759 vdd.n1540 gnd 0.010896f
C3760 vdd.n1541 gnd 0.00877f
C3761 vdd.n1542 gnd 0.010896f
C3762 vdd.n1543 gnd 0.00877f
C3763 vdd.n1544 gnd 0.010896f
C3764 vdd.n1545 gnd 1.11351f
C3765 vdd.n1546 gnd 0.010896f
C3766 vdd.n1547 gnd 0.00877f
C3767 vdd.n1548 gnd 0.026358f
C3768 vdd.n1549 gnd 0.007279f
C3769 vdd.n1550 gnd 0.026358f
C3770 vdd.t261 gnd 0.556753f
C3771 vdd.n1551 gnd 0.026358f
C3772 vdd.n1552 gnd 0.007279f
C3773 vdd.n1553 gnd 0.010896f
C3774 vdd.n1554 gnd 0.00877f
C3775 vdd.n1555 gnd 0.010896f
C3776 vdd.n1586 gnd 0.026923f
C3777 vdd.n1587 gnd 1.64242f
C3778 vdd.n1588 gnd 0.010896f
C3779 vdd.n1589 gnd 0.00877f
C3780 vdd.n1590 gnd 0.010896f
C3781 vdd.n1591 gnd 0.010896f
C3782 vdd.n1592 gnd 0.010896f
C3783 vdd.n1593 gnd 0.010896f
C3784 vdd.n1594 gnd 0.010896f
C3785 vdd.n1595 gnd 0.00877f
C3786 vdd.n1596 gnd 0.010896f
C3787 vdd.n1597 gnd 0.010896f
C3788 vdd.n1598 gnd 0.010896f
C3789 vdd.n1599 gnd 0.010896f
C3790 vdd.n1600 gnd 0.010896f
C3791 vdd.n1601 gnd 0.00877f
C3792 vdd.n1602 gnd 0.010896f
C3793 vdd.n1603 gnd 0.010896f
C3794 vdd.n1604 gnd 0.010896f
C3795 vdd.n1605 gnd 0.010896f
C3796 vdd.n1606 gnd 0.010896f
C3797 vdd.n1607 gnd 0.00877f
C3798 vdd.n1608 gnd 0.010896f
C3799 vdd.n1609 gnd 0.010896f
C3800 vdd.n1610 gnd 0.010896f
C3801 vdd.n1611 gnd 0.010896f
C3802 vdd.n1612 gnd 0.010896f
C3803 vdd.t292 gnd 0.134048f
C3804 vdd.t293 gnd 0.14326f
C3805 vdd.t291 gnd 0.175065f
C3806 vdd.n1613 gnd 0.224408f
C3807 vdd.n1614 gnd 0.18942f
C3808 vdd.n1615 gnd 0.018768f
C3809 vdd.n1616 gnd 0.010896f
C3810 vdd.n1617 gnd 0.010896f
C3811 vdd.n1618 gnd 0.010896f
C3812 vdd.n1619 gnd 0.010896f
C3813 vdd.n1620 gnd 0.010896f
C3814 vdd.n1621 gnd 0.00877f
C3815 vdd.n1622 gnd 0.010896f
C3816 vdd.n1623 gnd 0.010896f
C3817 vdd.n1624 gnd 0.010896f
C3818 vdd.n1625 gnd 0.010896f
C3819 vdd.n1626 gnd 0.010896f
C3820 vdd.n1627 gnd 0.00877f
C3821 vdd.n1628 gnd 0.010896f
C3822 vdd.n1629 gnd 0.010896f
C3823 vdd.n1630 gnd 0.010896f
C3824 vdd.n1631 gnd 0.010896f
C3825 vdd.n1632 gnd 0.010896f
C3826 vdd.n1633 gnd 0.00877f
C3827 vdd.n1634 gnd 0.010896f
C3828 vdd.n1635 gnd 0.010896f
C3829 vdd.n1636 gnd 0.010896f
C3830 vdd.n1637 gnd 0.010896f
C3831 vdd.n1638 gnd 0.010896f
C3832 vdd.n1639 gnd 0.00877f
C3833 vdd.n1640 gnd 0.010896f
C3834 vdd.n1641 gnd 0.010896f
C3835 vdd.n1642 gnd 0.010896f
C3836 vdd.n1643 gnd 0.010896f
C3837 vdd.n1644 gnd 0.010896f
C3838 vdd.n1645 gnd 0.00877f
C3839 vdd.n1646 gnd 0.010896f
C3840 vdd.n1647 gnd 0.010896f
C3841 vdd.n1648 gnd 0.010896f
C3842 vdd.n1649 gnd 0.010896f
C3843 vdd.n1650 gnd 0.00877f
C3844 vdd.n1651 gnd 0.010896f
C3845 vdd.n1652 gnd 0.010896f
C3846 vdd.n1653 gnd 0.010896f
C3847 vdd.n1654 gnd 0.010896f
C3848 vdd.n1655 gnd 0.010896f
C3849 vdd.n1656 gnd 0.00877f
C3850 vdd.n1657 gnd 0.010896f
C3851 vdd.n1658 gnd 0.010896f
C3852 vdd.n1659 gnd 0.010896f
C3853 vdd.n1660 gnd 0.010896f
C3854 vdd.n1661 gnd 0.010896f
C3855 vdd.n1662 gnd 0.00877f
C3856 vdd.n1663 gnd 0.010896f
C3857 vdd.n1664 gnd 0.010896f
C3858 vdd.n1665 gnd 0.010896f
C3859 vdd.n1666 gnd 0.010896f
C3860 vdd.n1667 gnd 0.010896f
C3861 vdd.n1668 gnd 0.00877f
C3862 vdd.n1669 gnd 0.010896f
C3863 vdd.n1670 gnd 0.010896f
C3864 vdd.n1671 gnd 0.010896f
C3865 vdd.n1672 gnd 0.010896f
C3866 vdd.n1673 gnd 0.010896f
C3867 vdd.n1674 gnd 0.00877f
C3868 vdd.n1675 gnd 0.010896f
C3869 vdd.n1676 gnd 0.010896f
C3870 vdd.n1677 gnd 0.010896f
C3871 vdd.n1678 gnd 0.010896f
C3872 vdd.t262 gnd 0.134048f
C3873 vdd.t263 gnd 0.14326f
C3874 vdd.t260 gnd 0.175065f
C3875 vdd.n1679 gnd 0.224408f
C3876 vdd.n1680 gnd 0.18942f
C3877 vdd.n1681 gnd 0.014383f
C3878 vdd.n1682 gnd 0.004166f
C3879 vdd.n1683 gnd 0.026923f
C3880 vdd.n1684 gnd 0.010896f
C3881 vdd.n1685 gnd 0.004604f
C3882 vdd.n1686 gnd 0.00877f
C3883 vdd.n1687 gnd 0.00877f
C3884 vdd.n1688 gnd 0.010896f
C3885 vdd.n1689 gnd 0.010896f
C3886 vdd.n1690 gnd 0.010896f
C3887 vdd.n1691 gnd 0.00877f
C3888 vdd.n1692 gnd 0.00877f
C3889 vdd.n1693 gnd 0.00877f
C3890 vdd.n1694 gnd 0.010896f
C3891 vdd.n1695 gnd 0.010896f
C3892 vdd.n1696 gnd 0.010896f
C3893 vdd.n1697 gnd 0.00877f
C3894 vdd.n1698 gnd 0.00877f
C3895 vdd.n1699 gnd 0.00877f
C3896 vdd.n1700 gnd 0.010896f
C3897 vdd.n1701 gnd 0.010896f
C3898 vdd.n1702 gnd 0.010896f
C3899 vdd.n1703 gnd 0.00877f
C3900 vdd.n1704 gnd 0.00877f
C3901 vdd.n1705 gnd 0.00877f
C3902 vdd.n1706 gnd 0.010896f
C3903 vdd.n1707 gnd 0.010896f
C3904 vdd.n1708 gnd 0.010896f
C3905 vdd.n1709 gnd 0.00877f
C3906 vdd.n1710 gnd 0.00877f
C3907 vdd.n1711 gnd 0.00877f
C3908 vdd.n1712 gnd 0.010896f
C3909 vdd.n1713 gnd 0.010896f
C3910 vdd.n1714 gnd 0.010896f
C3911 vdd.n1715 gnd 0.008682f
C3912 vdd.n1716 gnd 0.010896f
C3913 vdd.t279 gnd 0.134048f
C3914 vdd.t280 gnd 0.14326f
C3915 vdd.t278 gnd 0.175065f
C3916 vdd.n1717 gnd 0.224408f
C3917 vdd.n1718 gnd 0.18942f
C3918 vdd.n1719 gnd 0.018768f
C3919 vdd.n1720 gnd 0.005964f
C3920 vdd.n1721 gnd 0.010896f
C3921 vdd.n1722 gnd 0.010896f
C3922 vdd.n1723 gnd 0.010896f
C3923 vdd.n1724 gnd 0.00877f
C3924 vdd.n1725 gnd 0.00877f
C3925 vdd.n1726 gnd 0.00877f
C3926 vdd.n1727 gnd 0.010896f
C3927 vdd.n1728 gnd 0.010896f
C3928 vdd.n1729 gnd 0.010896f
C3929 vdd.n1730 gnd 0.00877f
C3930 vdd.n1731 gnd 0.00877f
C3931 vdd.n1732 gnd 0.00877f
C3932 vdd.n1733 gnd 0.010896f
C3933 vdd.n1734 gnd 0.010896f
C3934 vdd.n1735 gnd 0.010896f
C3935 vdd.n1736 gnd 0.00877f
C3936 vdd.n1737 gnd 0.00877f
C3937 vdd.n1738 gnd 0.00877f
C3938 vdd.n1739 gnd 0.010896f
C3939 vdd.n1740 gnd 0.010896f
C3940 vdd.n1741 gnd 0.010896f
C3941 vdd.n1742 gnd 0.00877f
C3942 vdd.n1743 gnd 0.00877f
C3943 vdd.n1744 gnd 0.00877f
C3944 vdd.n1745 gnd 0.010896f
C3945 vdd.n1746 gnd 0.010896f
C3946 vdd.n1747 gnd 0.010896f
C3947 vdd.n1748 gnd 0.00877f
C3948 vdd.n1749 gnd 0.00877f
C3949 vdd.n1750 gnd 0.007323f
C3950 vdd.n1751 gnd 0.010896f
C3951 vdd.n1752 gnd 0.010896f
C3952 vdd.n1753 gnd 0.010896f
C3953 vdd.n1754 gnd 0.007323f
C3954 vdd.n1755 gnd 0.00877f
C3955 vdd.n1756 gnd 0.00877f
C3956 vdd.n1757 gnd 0.010896f
C3957 vdd.n1758 gnd 0.010896f
C3958 vdd.n1759 gnd 0.010896f
C3959 vdd.n1760 gnd 0.00877f
C3960 vdd.n1761 gnd 0.00877f
C3961 vdd.n1762 gnd 0.00877f
C3962 vdd.n1763 gnd 0.010896f
C3963 vdd.n1764 gnd 0.010896f
C3964 vdd.n1765 gnd 0.010896f
C3965 vdd.n1766 gnd 0.00877f
C3966 vdd.n1767 gnd 0.00877f
C3967 vdd.n1768 gnd 0.00877f
C3968 vdd.n1769 gnd 0.010896f
C3969 vdd.n1770 gnd 0.010896f
C3970 vdd.n1771 gnd 0.010896f
C3971 vdd.n1772 gnd 0.00877f
C3972 vdd.n1773 gnd 0.00877f
C3973 vdd.n1774 gnd 0.00877f
C3974 vdd.n1775 gnd 0.010896f
C3975 vdd.n1776 gnd 0.010896f
C3976 vdd.n1777 gnd 0.010896f
C3977 vdd.n1778 gnd 0.00877f
C3978 vdd.n1779 gnd 0.010896f
C3979 vdd.n1780 gnd 2.63901f
C3980 vdd.n1782 gnd 0.026923f
C3981 vdd.n1783 gnd 0.007279f
C3982 vdd.n1784 gnd 0.026923f
C3983 vdd.n1785 gnd 0.026358f
C3984 vdd.n1786 gnd 0.010896f
C3985 vdd.n1787 gnd 0.00877f
C3986 vdd.n1788 gnd 0.010896f
C3987 vdd.n1789 gnd 0.56232f
C3988 vdd.n1790 gnd 0.010896f
C3989 vdd.n1791 gnd 0.00877f
C3990 vdd.n1792 gnd 0.010896f
C3991 vdd.n1793 gnd 0.010896f
C3992 vdd.n1794 gnd 0.010896f
C3993 vdd.n1795 gnd 0.00877f
C3994 vdd.n1796 gnd 0.010896f
C3995 vdd.n1797 gnd 1.01886f
C3996 vdd.n1798 gnd 1.11351f
C3997 vdd.n1799 gnd 0.010896f
C3998 vdd.n1800 gnd 0.00877f
C3999 vdd.n1801 gnd 0.010896f
C4000 vdd.n1802 gnd 0.010896f
C4001 vdd.n1803 gnd 0.010896f
C4002 vdd.n1804 gnd 0.00877f
C4003 vdd.n1805 gnd 0.010896f
C4004 vdd.n1806 gnd 0.651401f
C4005 vdd.n1807 gnd 0.010896f
C4006 vdd.n1808 gnd 0.00877f
C4007 vdd.n1809 gnd 0.010896f
C4008 vdd.n1810 gnd 0.010896f
C4009 vdd.n1811 gnd 0.010896f
C4010 vdd.n1812 gnd 0.00877f
C4011 vdd.n1813 gnd 0.010896f
C4012 vdd.n1814 gnd 0.640265f
C4013 vdd.n1815 gnd 0.840696f
C4014 vdd.n1816 gnd 0.010896f
C4015 vdd.n1817 gnd 0.00877f
C4016 vdd.n1818 gnd 0.010896f
C4017 vdd.n1819 gnd 0.010896f
C4018 vdd.n1820 gnd 0.010896f
C4019 vdd.n1821 gnd 0.00877f
C4020 vdd.n1822 gnd 0.010896f
C4021 vdd.n1823 gnd 0.924209f
C4022 vdd.n1824 gnd 0.010896f
C4023 vdd.n1825 gnd 0.00877f
C4024 vdd.n1826 gnd 0.010896f
C4025 vdd.n1827 gnd 0.010896f
C4026 vdd.n1828 gnd 0.010896f
C4027 vdd.n1829 gnd 0.00877f
C4028 vdd.n1830 gnd 0.010896f
C4029 vdd.t80 gnd 0.556753f
C4030 vdd.n1831 gnd 0.818426f
C4031 vdd.n1832 gnd 0.010896f
C4032 vdd.n1833 gnd 0.00877f
C4033 vdd.n1834 gnd 0.010896f
C4034 vdd.n1835 gnd 0.010896f
C4035 vdd.n1836 gnd 0.010896f
C4036 vdd.n1837 gnd 0.00877f
C4037 vdd.n1838 gnd 0.010896f
C4038 vdd.n1839 gnd 0.62913f
C4039 vdd.n1840 gnd 0.010896f
C4040 vdd.n1841 gnd 0.00877f
C4041 vdd.n1842 gnd 0.010896f
C4042 vdd.n1843 gnd 0.010896f
C4043 vdd.n1844 gnd 0.010896f
C4044 vdd.n1845 gnd 0.00877f
C4045 vdd.n1846 gnd 0.010896f
C4046 vdd.n1847 gnd 0.807291f
C4047 vdd.n1848 gnd 0.673671f
C4048 vdd.n1849 gnd 0.010896f
C4049 vdd.n1850 gnd 0.00877f
C4050 vdd.n1851 gnd 0.010896f
C4051 vdd.n1852 gnd 0.010896f
C4052 vdd.n1853 gnd 0.010896f
C4053 vdd.n1854 gnd 0.00877f
C4054 vdd.n1855 gnd 0.010896f
C4055 vdd.n1856 gnd 0.862966f
C4056 vdd.n1857 gnd 0.010896f
C4057 vdd.n1858 gnd 0.00877f
C4058 vdd.n1859 gnd 0.010896f
C4059 vdd.n1860 gnd 0.010896f
C4060 vdd.n1861 gnd 0.010896f
C4061 vdd.n1862 gnd 0.00877f
C4062 vdd.n1863 gnd 0.010896f
C4063 vdd.t162 gnd 0.556753f
C4064 vdd.n1864 gnd 0.924209f
C4065 vdd.n1865 gnd 0.010896f
C4066 vdd.n1866 gnd 0.00877f
C4067 vdd.n1867 gnd 0.010896f
C4068 vdd.n1868 gnd 0.008374f
C4069 vdd.n1869 gnd 0.00598f
C4070 vdd.n1870 gnd 0.005549f
C4071 vdd.n1871 gnd 0.003069f
C4072 vdd.n1872 gnd 0.007048f
C4073 vdd.n1873 gnd 0.002982f
C4074 vdd.n1874 gnd 0.003157f
C4075 vdd.n1875 gnd 0.005549f
C4076 vdd.n1876 gnd 0.002982f
C4077 vdd.n1877 gnd 0.007048f
C4078 vdd.n1878 gnd 0.003157f
C4079 vdd.n1879 gnd 0.005549f
C4080 vdd.n1880 gnd 0.002982f
C4081 vdd.n1881 gnd 0.005286f
C4082 vdd.n1882 gnd 0.005302f
C4083 vdd.t115 gnd 0.015142f
C4084 vdd.n1883 gnd 0.03369f
C4085 vdd.n1884 gnd 0.175329f
C4086 vdd.n1885 gnd 0.002982f
C4087 vdd.n1886 gnd 0.003157f
C4088 vdd.n1887 gnd 0.007048f
C4089 vdd.n1888 gnd 0.007048f
C4090 vdd.n1889 gnd 0.003157f
C4091 vdd.n1890 gnd 0.002982f
C4092 vdd.n1891 gnd 0.005549f
C4093 vdd.n1892 gnd 0.005549f
C4094 vdd.n1893 gnd 0.002982f
C4095 vdd.n1894 gnd 0.003157f
C4096 vdd.n1895 gnd 0.007048f
C4097 vdd.n1896 gnd 0.007048f
C4098 vdd.n1897 gnd 0.003157f
C4099 vdd.n1898 gnd 0.002982f
C4100 vdd.n1899 gnd 0.005549f
C4101 vdd.n1900 gnd 0.005549f
C4102 vdd.n1901 gnd 0.002982f
C4103 vdd.n1902 gnd 0.003157f
C4104 vdd.n1903 gnd 0.007048f
C4105 vdd.n1904 gnd 0.007048f
C4106 vdd.n1905 gnd 0.016662f
C4107 vdd.n1906 gnd 0.003069f
C4108 vdd.n1907 gnd 0.002982f
C4109 vdd.n1908 gnd 0.014342f
C4110 vdd.n1909 gnd 0.010013f
C4111 vdd.t143 gnd 0.035079f
C4112 vdd.t200 gnd 0.035079f
C4113 vdd.n1910 gnd 0.24109f
C4114 vdd.n1911 gnd 0.18958f
C4115 vdd.t166 gnd 0.035079f
C4116 vdd.t215 gnd 0.035079f
C4117 vdd.n1912 gnd 0.24109f
C4118 vdd.n1913 gnd 0.15299f
C4119 vdd.t131 gnd 0.035079f
C4120 vdd.t84 gnd 0.035079f
C4121 vdd.n1914 gnd 0.24109f
C4122 vdd.n1915 gnd 0.15299f
C4123 vdd.t155 gnd 0.035079f
C4124 vdd.t95 gnd 0.035079f
C4125 vdd.n1916 gnd 0.24109f
C4126 vdd.n1917 gnd 0.15299f
C4127 vdd.t204 gnd 0.035079f
C4128 vdd.t220 gnd 0.035079f
C4129 vdd.n1918 gnd 0.24109f
C4130 vdd.n1919 gnd 0.15299f
C4131 vdd.t177 gnd 0.035079f
C4132 vdd.t65 gnd 0.035079f
C4133 vdd.n1920 gnd 0.24109f
C4134 vdd.n1921 gnd 0.15299f
C4135 vdd.t167 gnd 0.035079f
C4136 vdd.t108 gnd 0.035079f
C4137 vdd.n1922 gnd 0.24109f
C4138 vdd.n1923 gnd 0.15299f
C4139 vdd.t209 gnd 0.035079f
C4140 vdd.t137 gnd 0.035079f
C4141 vdd.n1924 gnd 0.24109f
C4142 vdd.n1925 gnd 0.15299f
C4143 vdd.t187 gnd 0.035079f
C4144 vdd.t159 gnd 0.035079f
C4145 vdd.n1926 gnd 0.24109f
C4146 vdd.n1927 gnd 0.15299f
C4147 vdd.n1928 gnd 0.00598f
C4148 vdd.n1929 gnd 0.005549f
C4149 vdd.n1930 gnd 0.003069f
C4150 vdd.n1931 gnd 0.007048f
C4151 vdd.n1932 gnd 0.002982f
C4152 vdd.n1933 gnd 0.003157f
C4153 vdd.n1934 gnd 0.005549f
C4154 vdd.n1935 gnd 0.002982f
C4155 vdd.n1936 gnd 0.007048f
C4156 vdd.n1937 gnd 0.003157f
C4157 vdd.n1938 gnd 0.005549f
C4158 vdd.n1939 gnd 0.002982f
C4159 vdd.n1940 gnd 0.005286f
C4160 vdd.n1941 gnd 0.005302f
C4161 vdd.t73 gnd 0.015142f
C4162 vdd.n1942 gnd 0.03369f
C4163 vdd.n1943 gnd 0.175329f
C4164 vdd.n1944 gnd 0.002982f
C4165 vdd.n1945 gnd 0.003157f
C4166 vdd.n1946 gnd 0.007048f
C4167 vdd.n1947 gnd 0.007048f
C4168 vdd.n1948 gnd 0.003157f
C4169 vdd.n1949 gnd 0.002982f
C4170 vdd.n1950 gnd 0.005549f
C4171 vdd.n1951 gnd 0.005549f
C4172 vdd.n1952 gnd 0.002982f
C4173 vdd.n1953 gnd 0.003157f
C4174 vdd.n1954 gnd 0.007048f
C4175 vdd.n1955 gnd 0.007048f
C4176 vdd.n1956 gnd 0.003157f
C4177 vdd.n1957 gnd 0.002982f
C4178 vdd.n1958 gnd 0.005549f
C4179 vdd.n1959 gnd 0.005549f
C4180 vdd.n1960 gnd 0.002982f
C4181 vdd.n1961 gnd 0.003157f
C4182 vdd.n1962 gnd 0.007048f
C4183 vdd.n1963 gnd 0.007048f
C4184 vdd.n1964 gnd 0.016662f
C4185 vdd.n1965 gnd 0.003069f
C4186 vdd.n1966 gnd 0.002982f
C4187 vdd.n1967 gnd 0.014342f
C4188 vdd.n1968 gnd 0.009699f
C4189 vdd.n1969 gnd 0.113825f
C4190 vdd.n1970 gnd 0.00598f
C4191 vdd.n1971 gnd 0.005549f
C4192 vdd.n1972 gnd 0.003069f
C4193 vdd.n1973 gnd 0.007048f
C4194 vdd.n1974 gnd 0.002982f
C4195 vdd.n1975 gnd 0.003157f
C4196 vdd.n1976 gnd 0.005549f
C4197 vdd.n1977 gnd 0.002982f
C4198 vdd.n1978 gnd 0.007048f
C4199 vdd.n1979 gnd 0.003157f
C4200 vdd.n1980 gnd 0.005549f
C4201 vdd.n1981 gnd 0.002982f
C4202 vdd.n1982 gnd 0.005286f
C4203 vdd.n1983 gnd 0.005302f
C4204 vdd.t198 gnd 0.015142f
C4205 vdd.n1984 gnd 0.03369f
C4206 vdd.n1985 gnd 0.175329f
C4207 vdd.n1986 gnd 0.002982f
C4208 vdd.n1987 gnd 0.003157f
C4209 vdd.n1988 gnd 0.007048f
C4210 vdd.n1989 gnd 0.007048f
C4211 vdd.n1990 gnd 0.003157f
C4212 vdd.n1991 gnd 0.002982f
C4213 vdd.n1992 gnd 0.005549f
C4214 vdd.n1993 gnd 0.005549f
C4215 vdd.n1994 gnd 0.002982f
C4216 vdd.n1995 gnd 0.003157f
C4217 vdd.n1996 gnd 0.007048f
C4218 vdd.n1997 gnd 0.007048f
C4219 vdd.n1998 gnd 0.003157f
C4220 vdd.n1999 gnd 0.002982f
C4221 vdd.n2000 gnd 0.005549f
C4222 vdd.n2001 gnd 0.005549f
C4223 vdd.n2002 gnd 0.002982f
C4224 vdd.n2003 gnd 0.003157f
C4225 vdd.n2004 gnd 0.007048f
C4226 vdd.n2005 gnd 0.007048f
C4227 vdd.n2006 gnd 0.016662f
C4228 vdd.n2007 gnd 0.003069f
C4229 vdd.n2008 gnd 0.002982f
C4230 vdd.n2009 gnd 0.014342f
C4231 vdd.n2010 gnd 0.010013f
C4232 vdd.t147 gnd 0.035079f
C4233 vdd.t77 gnd 0.035079f
C4234 vdd.n2011 gnd 0.24109f
C4235 vdd.n2012 gnd 0.18958f
C4236 vdd.t211 gnd 0.035079f
C4237 vdd.t179 gnd 0.035079f
C4238 vdd.n2013 gnd 0.24109f
C4239 vdd.n2014 gnd 0.15299f
C4240 vdd.t173 gnd 0.035079f
C4241 vdd.t116 gnd 0.035079f
C4242 vdd.n2015 gnd 0.24109f
C4243 vdd.n2016 gnd 0.15299f
C4244 vdd.t110 gnd 0.035079f
C4245 vdd.t174 gnd 0.035079f
C4246 vdd.n2017 gnd 0.24109f
C4247 vdd.n2018 gnd 0.15299f
C4248 vdd.t163 gnd 0.035079f
C4249 vdd.t161 gnd 0.035079f
C4250 vdd.n2019 gnd 0.24109f
C4251 vdd.n2020 gnd 0.15299f
C4252 vdd.t106 gnd 0.035079f
C4253 vdd.t82 gnd 0.035079f
C4254 vdd.n2021 gnd 0.24109f
C4255 vdd.n2022 gnd 0.15299f
C4256 vdd.t69 gnd 0.035079f
C4257 vdd.t156 gnd 0.035079f
C4258 vdd.n2023 gnd 0.24109f
C4259 vdd.n2024 gnd 0.15299f
C4260 vdd.t133 gnd 0.035079f
C4261 vdd.t81 gnd 0.035079f
C4262 vdd.n2025 gnd 0.24109f
C4263 vdd.n2026 gnd 0.15299f
C4264 vdd.t63 gnd 0.035079f
C4265 vdd.t180 gnd 0.035079f
C4266 vdd.n2027 gnd 0.24109f
C4267 vdd.n2028 gnd 0.15299f
C4268 vdd.n2029 gnd 0.00598f
C4269 vdd.n2030 gnd 0.005549f
C4270 vdd.n2031 gnd 0.003069f
C4271 vdd.n2032 gnd 0.007048f
C4272 vdd.n2033 gnd 0.002982f
C4273 vdd.n2034 gnd 0.003157f
C4274 vdd.n2035 gnd 0.005549f
C4275 vdd.n2036 gnd 0.002982f
C4276 vdd.n2037 gnd 0.007048f
C4277 vdd.n2038 gnd 0.003157f
C4278 vdd.n2039 gnd 0.005549f
C4279 vdd.n2040 gnd 0.002982f
C4280 vdd.n2041 gnd 0.005286f
C4281 vdd.n2042 gnd 0.005302f
C4282 vdd.t121 gnd 0.015142f
C4283 vdd.n2043 gnd 0.03369f
C4284 vdd.n2044 gnd 0.175329f
C4285 vdd.n2045 gnd 0.002982f
C4286 vdd.n2046 gnd 0.003157f
C4287 vdd.n2047 gnd 0.007048f
C4288 vdd.n2048 gnd 0.007048f
C4289 vdd.n2049 gnd 0.003157f
C4290 vdd.n2050 gnd 0.002982f
C4291 vdd.n2051 gnd 0.005549f
C4292 vdd.n2052 gnd 0.005549f
C4293 vdd.n2053 gnd 0.002982f
C4294 vdd.n2054 gnd 0.003157f
C4295 vdd.n2055 gnd 0.007048f
C4296 vdd.n2056 gnd 0.007048f
C4297 vdd.n2057 gnd 0.003157f
C4298 vdd.n2058 gnd 0.002982f
C4299 vdd.n2059 gnd 0.005549f
C4300 vdd.n2060 gnd 0.005549f
C4301 vdd.n2061 gnd 0.002982f
C4302 vdd.n2062 gnd 0.003157f
C4303 vdd.n2063 gnd 0.007048f
C4304 vdd.n2064 gnd 0.007048f
C4305 vdd.n2065 gnd 0.016662f
C4306 vdd.n2066 gnd 0.003069f
C4307 vdd.n2067 gnd 0.002982f
C4308 vdd.n2068 gnd 0.014342f
C4309 vdd.n2069 gnd 0.009699f
C4310 vdd.n2070 gnd 0.067715f
C4311 vdd.n2071 gnd 0.243994f
C4312 vdd.n2072 gnd 0.00598f
C4313 vdd.n2073 gnd 0.005549f
C4314 vdd.n2074 gnd 0.003069f
C4315 vdd.n2075 gnd 0.007048f
C4316 vdd.n2076 gnd 0.002982f
C4317 vdd.n2077 gnd 0.003157f
C4318 vdd.n2078 gnd 0.005549f
C4319 vdd.n2079 gnd 0.002982f
C4320 vdd.n2080 gnd 0.007048f
C4321 vdd.n2081 gnd 0.003157f
C4322 vdd.n2082 gnd 0.005549f
C4323 vdd.n2083 gnd 0.002982f
C4324 vdd.n2084 gnd 0.005286f
C4325 vdd.n2085 gnd 0.005302f
C4326 vdd.t210 gnd 0.015142f
C4327 vdd.n2086 gnd 0.03369f
C4328 vdd.n2087 gnd 0.175329f
C4329 vdd.n2088 gnd 0.002982f
C4330 vdd.n2089 gnd 0.003157f
C4331 vdd.n2090 gnd 0.007048f
C4332 vdd.n2091 gnd 0.007048f
C4333 vdd.n2092 gnd 0.003157f
C4334 vdd.n2093 gnd 0.002982f
C4335 vdd.n2094 gnd 0.005549f
C4336 vdd.n2095 gnd 0.005549f
C4337 vdd.n2096 gnd 0.002982f
C4338 vdd.n2097 gnd 0.003157f
C4339 vdd.n2098 gnd 0.007048f
C4340 vdd.n2099 gnd 0.007048f
C4341 vdd.n2100 gnd 0.003157f
C4342 vdd.n2101 gnd 0.002982f
C4343 vdd.n2102 gnd 0.005549f
C4344 vdd.n2103 gnd 0.005549f
C4345 vdd.n2104 gnd 0.002982f
C4346 vdd.n2105 gnd 0.003157f
C4347 vdd.n2106 gnd 0.007048f
C4348 vdd.n2107 gnd 0.007048f
C4349 vdd.n2108 gnd 0.016662f
C4350 vdd.n2109 gnd 0.003069f
C4351 vdd.n2110 gnd 0.002982f
C4352 vdd.n2111 gnd 0.014342f
C4353 vdd.n2112 gnd 0.010013f
C4354 vdd.t164 gnd 0.035079f
C4355 vdd.t100 gnd 0.035079f
C4356 vdd.n2113 gnd 0.24109f
C4357 vdd.n2114 gnd 0.18958f
C4358 vdd.t221 gnd 0.035079f
C4359 vdd.t193 gnd 0.035079f
C4360 vdd.n2115 gnd 0.24109f
C4361 vdd.n2116 gnd 0.15299f
C4362 vdd.t189 gnd 0.035079f
C4363 vdd.t138 gnd 0.035079f
C4364 vdd.n2117 gnd 0.24109f
C4365 vdd.n2118 gnd 0.15299f
C4366 vdd.t134 gnd 0.035079f
C4367 vdd.t192 gnd 0.035079f
C4368 vdd.n2119 gnd 0.24109f
C4369 vdd.n2120 gnd 0.15299f
C4370 vdd.t172 gnd 0.035079f
C4371 vdd.t171 gnd 0.035079f
C4372 vdd.n2121 gnd 0.24109f
C4373 vdd.n2122 gnd 0.15299f
C4374 vdd.t129 gnd 0.035079f
C4375 vdd.t102 gnd 0.035079f
C4376 vdd.n2123 gnd 0.24109f
C4377 vdd.n2124 gnd 0.15299f
C4378 vdd.t99 gnd 0.035079f
C4379 vdd.t170 gnd 0.035079f
C4380 vdd.n2125 gnd 0.24109f
C4381 vdd.n2126 gnd 0.15299f
C4382 vdd.t149 gnd 0.035079f
C4383 vdd.t101 gnd 0.035079f
C4384 vdd.n2127 gnd 0.24109f
C4385 vdd.n2128 gnd 0.15299f
C4386 vdd.t93 gnd 0.035079f
C4387 vdd.t191 gnd 0.035079f
C4388 vdd.n2129 gnd 0.24109f
C4389 vdd.n2130 gnd 0.15299f
C4390 vdd.n2131 gnd 0.00598f
C4391 vdd.n2132 gnd 0.005549f
C4392 vdd.n2133 gnd 0.003069f
C4393 vdd.n2134 gnd 0.007048f
C4394 vdd.n2135 gnd 0.002982f
C4395 vdd.n2136 gnd 0.003157f
C4396 vdd.n2137 gnd 0.005549f
C4397 vdd.n2138 gnd 0.002982f
C4398 vdd.n2139 gnd 0.007048f
C4399 vdd.n2140 gnd 0.003157f
C4400 vdd.n2141 gnd 0.005549f
C4401 vdd.n2142 gnd 0.002982f
C4402 vdd.n2143 gnd 0.005286f
C4403 vdd.n2144 gnd 0.005302f
C4404 vdd.t144 gnd 0.015142f
C4405 vdd.n2145 gnd 0.03369f
C4406 vdd.n2146 gnd 0.175329f
C4407 vdd.n2147 gnd 0.002982f
C4408 vdd.n2148 gnd 0.003157f
C4409 vdd.n2149 gnd 0.007048f
C4410 vdd.n2150 gnd 0.007048f
C4411 vdd.n2151 gnd 0.003157f
C4412 vdd.n2152 gnd 0.002982f
C4413 vdd.n2153 gnd 0.005549f
C4414 vdd.n2154 gnd 0.005549f
C4415 vdd.n2155 gnd 0.002982f
C4416 vdd.n2156 gnd 0.003157f
C4417 vdd.n2157 gnd 0.007048f
C4418 vdd.n2158 gnd 0.007048f
C4419 vdd.n2159 gnd 0.003157f
C4420 vdd.n2160 gnd 0.002982f
C4421 vdd.n2161 gnd 0.005549f
C4422 vdd.n2162 gnd 0.005549f
C4423 vdd.n2163 gnd 0.002982f
C4424 vdd.n2164 gnd 0.003157f
C4425 vdd.n2165 gnd 0.007048f
C4426 vdd.n2166 gnd 0.007048f
C4427 vdd.n2167 gnd 0.016662f
C4428 vdd.n2168 gnd 0.003069f
C4429 vdd.n2169 gnd 0.002982f
C4430 vdd.n2170 gnd 0.014342f
C4431 vdd.n2171 gnd 0.009699f
C4432 vdd.n2172 gnd 0.067715f
C4433 vdd.n2173 gnd 0.27932f
C4434 vdd.n2174 gnd 2.93017f
C4435 vdd.n2175 gnd 0.642679f
C4436 vdd.n2176 gnd 0.008374f
C4437 vdd.n2177 gnd 0.00877f
C4438 vdd.n2178 gnd 0.010896f
C4439 vdd.n2179 gnd 0.796156f
C4440 vdd.n2180 gnd 0.010896f
C4441 vdd.n2181 gnd 0.00877f
C4442 vdd.n2182 gnd 0.010896f
C4443 vdd.n2183 gnd 0.010896f
C4444 vdd.n2184 gnd 0.010896f
C4445 vdd.n2185 gnd 0.00877f
C4446 vdd.n2186 gnd 0.010896f
C4447 vdd.n2187 gnd 0.924209f
C4448 vdd.t109 gnd 0.556753f
C4449 vdd.n2188 gnd 0.60686f
C4450 vdd.n2189 gnd 0.010896f
C4451 vdd.n2190 gnd 0.00877f
C4452 vdd.n2191 gnd 0.010896f
C4453 vdd.n2192 gnd 0.010896f
C4454 vdd.n2193 gnd 0.010896f
C4455 vdd.n2194 gnd 0.00877f
C4456 vdd.n2195 gnd 0.010896f
C4457 vdd.n2196 gnd 0.695941f
C4458 vdd.n2197 gnd 0.010896f
C4459 vdd.n2198 gnd 0.00877f
C4460 vdd.n2199 gnd 0.010896f
C4461 vdd.n2200 gnd 0.010896f
C4462 vdd.n2201 gnd 0.010896f
C4463 vdd.n2202 gnd 0.00877f
C4464 vdd.n2203 gnd 0.010896f
C4465 vdd.n2204 gnd 0.595725f
C4466 vdd.n2205 gnd 0.885237f
C4467 vdd.n2206 gnd 0.010896f
C4468 vdd.n2207 gnd 0.00877f
C4469 vdd.n2208 gnd 0.010896f
C4470 vdd.n2209 gnd 0.010896f
C4471 vdd.n2210 gnd 0.010896f
C4472 vdd.n2211 gnd 0.00877f
C4473 vdd.n2212 gnd 0.010896f
C4474 vdd.n2213 gnd 0.924209f
C4475 vdd.n2214 gnd 0.010896f
C4476 vdd.n2215 gnd 0.00877f
C4477 vdd.n2216 gnd 0.010896f
C4478 vdd.n2217 gnd 0.010896f
C4479 vdd.n2218 gnd 0.010896f
C4480 vdd.n2219 gnd 0.00877f
C4481 vdd.n2220 gnd 0.010896f
C4482 vdd.t178 gnd 0.556753f
C4483 vdd.n2221 gnd 0.773886f
C4484 vdd.n2222 gnd 0.010896f
C4485 vdd.n2223 gnd 0.00877f
C4486 vdd.n2224 gnd 0.010896f
C4487 vdd.n2225 gnd 0.010896f
C4488 vdd.n2226 gnd 0.010896f
C4489 vdd.n2227 gnd 0.00877f
C4490 vdd.n2228 gnd 0.010896f
C4491 vdd.n2229 gnd 0.58459f
C4492 vdd.n2230 gnd 0.010896f
C4493 vdd.n2231 gnd 0.00877f
C4494 vdd.n2232 gnd 0.010896f
C4495 vdd.n2233 gnd 0.010896f
C4496 vdd.n2234 gnd 0.010896f
C4497 vdd.n2235 gnd 0.00877f
C4498 vdd.n2236 gnd 0.010896f
C4499 vdd.n2237 gnd 0.762751f
C4500 vdd.n2238 gnd 0.718211f
C4501 vdd.n2239 gnd 0.010896f
C4502 vdd.n2240 gnd 0.00877f
C4503 vdd.n2241 gnd 0.010896f
C4504 vdd.n2242 gnd 0.010896f
C4505 vdd.n2243 gnd 0.010896f
C4506 vdd.n2244 gnd 0.00877f
C4507 vdd.n2245 gnd 0.010896f
C4508 vdd.n2246 gnd 0.907507f
C4509 vdd.n2247 gnd 0.010896f
C4510 vdd.n2248 gnd 0.00877f
C4511 vdd.n2249 gnd 0.010896f
C4512 vdd.n2250 gnd 0.010896f
C4513 vdd.n2251 gnd 0.026358f
C4514 vdd.n2252 gnd 0.010896f
C4515 vdd.n2253 gnd 0.010896f
C4516 vdd.n2254 gnd 0.00877f
C4517 vdd.n2255 gnd 0.010896f
C4518 vdd.n2256 gnd 0.673671f
C4519 vdd.n2257 gnd 1.11351f
C4520 vdd.n2258 gnd 0.010896f
C4521 vdd.n2259 gnd 0.00877f
C4522 vdd.n2260 gnd 0.010896f
C4523 vdd.n2261 gnd 0.010896f
C4524 vdd.n2262 gnd 0.026358f
C4525 vdd.n2263 gnd 0.007279f
C4526 vdd.n2264 gnd 0.026358f
C4527 vdd.n2265 gnd 1.53107f
C4528 vdd.n2266 gnd 0.026358f
C4529 vdd.n2267 gnd 0.026923f
C4530 vdd.n2268 gnd 0.004166f
C4531 vdd.t239 gnd 0.134048f
C4532 vdd.t238 gnd 0.14326f
C4533 vdd.t236 gnd 0.175065f
C4534 vdd.n2269 gnd 0.224408f
C4535 vdd.n2270 gnd 0.188543f
C4536 vdd.n2271 gnd 0.013506f
C4537 vdd.n2272 gnd 0.004604f
C4538 vdd.n2273 gnd 0.00937f
C4539 vdd.n2274 gnd 0.824004f
C4540 vdd.n2276 gnd 0.00877f
C4541 vdd.n2277 gnd 0.00877f
C4542 vdd.n2278 gnd 0.010896f
C4543 vdd.n2280 gnd 0.010896f
C4544 vdd.n2281 gnd 0.010896f
C4545 vdd.n2282 gnd 0.00877f
C4546 vdd.n2283 gnd 0.00877f
C4547 vdd.n2284 gnd 0.00877f
C4548 vdd.n2285 gnd 0.010896f
C4549 vdd.n2287 gnd 0.010896f
C4550 vdd.n2288 gnd 0.010896f
C4551 vdd.n2289 gnd 0.00877f
C4552 vdd.n2290 gnd 0.00877f
C4553 vdd.n2291 gnd 0.00877f
C4554 vdd.n2292 gnd 0.010896f
C4555 vdd.n2294 gnd 0.010896f
C4556 vdd.n2295 gnd 0.010896f
C4557 vdd.n2296 gnd 0.00877f
C4558 vdd.n2297 gnd 0.00877f
C4559 vdd.n2298 gnd 0.00877f
C4560 vdd.n2299 gnd 0.010896f
C4561 vdd.n2301 gnd 0.010896f
C4562 vdd.n2302 gnd 0.010896f
C4563 vdd.n2303 gnd 0.00877f
C4564 vdd.n2304 gnd 0.010896f
C4565 vdd.n2305 gnd 0.010896f
C4566 vdd.n2306 gnd 0.010896f
C4567 vdd.n2307 gnd 0.01789f
C4568 vdd.n2308 gnd 0.005964f
C4569 vdd.n2309 gnd 0.00877f
C4570 vdd.n2310 gnd 0.010896f
C4571 vdd.n2312 gnd 0.010896f
C4572 vdd.n2313 gnd 0.010896f
C4573 vdd.n2314 gnd 0.00877f
C4574 vdd.n2315 gnd 0.00877f
C4575 vdd.n2316 gnd 0.00877f
C4576 vdd.n2317 gnd 0.010896f
C4577 vdd.n2319 gnd 0.010896f
C4578 vdd.n2320 gnd 0.010896f
C4579 vdd.n2321 gnd 0.00877f
C4580 vdd.n2322 gnd 0.00877f
C4581 vdd.n2323 gnd 0.00877f
C4582 vdd.n2324 gnd 0.010896f
C4583 vdd.n2326 gnd 0.010896f
C4584 vdd.n2327 gnd 0.010896f
C4585 vdd.n2328 gnd 0.00877f
C4586 vdd.n2329 gnd 0.00877f
C4587 vdd.n2330 gnd 0.00877f
C4588 vdd.n2331 gnd 0.010896f
C4589 vdd.n2333 gnd 0.010896f
C4590 vdd.n2334 gnd 0.010896f
C4591 vdd.n2335 gnd 0.00877f
C4592 vdd.n2336 gnd 0.00877f
C4593 vdd.n2337 gnd 0.00877f
C4594 vdd.n2338 gnd 0.010896f
C4595 vdd.n2340 gnd 0.010896f
C4596 vdd.n2341 gnd 0.010896f
C4597 vdd.n2342 gnd 0.00877f
C4598 vdd.n2343 gnd 0.010896f
C4599 vdd.n2344 gnd 0.010896f
C4600 vdd.n2345 gnd 0.010896f
C4601 vdd.n2346 gnd 0.01789f
C4602 vdd.n2347 gnd 0.007323f
C4603 vdd.n2348 gnd 0.00877f
C4604 vdd.n2349 gnd 0.010896f
C4605 vdd.n2351 gnd 0.010896f
C4606 vdd.n2352 gnd 0.010896f
C4607 vdd.n2353 gnd 0.00877f
C4608 vdd.n2354 gnd 0.00877f
C4609 vdd.n2355 gnd 0.00877f
C4610 vdd.n2356 gnd 0.010896f
C4611 vdd.n2358 gnd 0.010896f
C4612 vdd.n2359 gnd 0.010896f
C4613 vdd.n2360 gnd 0.00877f
C4614 vdd.n2361 gnd 0.00877f
C4615 vdd.n2362 gnd 0.00877f
C4616 vdd.n2363 gnd 0.010896f
C4617 vdd.n2365 gnd 0.010896f
C4618 vdd.n2366 gnd 0.010896f
C4619 vdd.n2367 gnd 0.00877f
C4620 vdd.n2368 gnd 0.00877f
C4621 vdd.n2369 gnd 0.00877f
C4622 vdd.n2370 gnd 0.010896f
C4623 vdd.n2372 gnd 0.010896f
C4624 vdd.n2373 gnd 0.00877f
C4625 vdd.n2374 gnd 0.00877f
C4626 vdd.n2375 gnd 0.010896f
C4627 vdd.n2377 gnd 0.010896f
C4628 vdd.n2378 gnd 0.010896f
C4629 vdd.n2379 gnd 0.00877f
C4630 vdd.n2380 gnd 0.00937f
C4631 vdd.n2381 gnd 0.824004f
C4632 vdd.n2382 gnd 0.029696f
C4633 vdd.n2383 gnd 0.007409f
C4634 vdd.n2384 gnd 0.007409f
C4635 vdd.n2385 gnd 0.007409f
C4636 vdd.n2386 gnd 0.007409f
C4637 vdd.n2387 gnd 0.007409f
C4638 vdd.n2388 gnd 0.007409f
C4639 vdd.n2389 gnd 0.007409f
C4640 vdd.n2390 gnd 0.007409f
C4641 vdd.n2391 gnd 0.007409f
C4642 vdd.n2392 gnd 0.007409f
C4643 vdd.n2393 gnd 0.007409f
C4644 vdd.n2394 gnd 0.007409f
C4645 vdd.n2395 gnd 0.007409f
C4646 vdd.n2396 gnd 0.007409f
C4647 vdd.n2397 gnd 0.007409f
C4648 vdd.n2398 gnd 0.007409f
C4649 vdd.n2399 gnd 0.007409f
C4650 vdd.n2400 gnd 0.007409f
C4651 vdd.n2401 gnd 0.007409f
C4652 vdd.n2402 gnd 0.007409f
C4653 vdd.n2403 gnd 0.007409f
C4654 vdd.n2404 gnd 0.007409f
C4655 vdd.n2405 gnd 0.007409f
C4656 vdd.n2406 gnd 0.007409f
C4657 vdd.n2407 gnd 0.007409f
C4658 vdd.n2408 gnd 0.007409f
C4659 vdd.n2409 gnd 0.007409f
C4660 vdd.n2410 gnd 0.007409f
C4661 vdd.n2411 gnd 0.007409f
C4662 vdd.n2412 gnd 0.007409f
C4663 vdd.n2413 gnd 0.007409f
C4664 vdd.n2414 gnd 0.01733f
C4665 vdd.n2415 gnd 0.01733f
C4666 vdd.n2417 gnd 9.4982f
C4667 vdd.n2419 gnd 0.01733f
C4668 vdd.n2420 gnd 0.01733f
C4669 vdd.n2421 gnd 0.01623f
C4670 vdd.n2422 gnd 0.007409f
C4671 vdd.n2423 gnd 0.007409f
C4672 vdd.n2424 gnd 0.757183f
C4673 vdd.n2425 gnd 0.007409f
C4674 vdd.n2426 gnd 0.007409f
C4675 vdd.n2427 gnd 0.007409f
C4676 vdd.n2428 gnd 0.007409f
C4677 vdd.n2429 gnd 0.007409f
C4678 vdd.n2430 gnd 0.640265f
C4679 vdd.n2431 gnd 0.007409f
C4680 vdd.n2432 gnd 0.007409f
C4681 vdd.n2433 gnd 0.007409f
C4682 vdd.n2434 gnd 0.007409f
C4683 vdd.n2435 gnd 0.007409f
C4684 vdd.n2436 gnd 0.757183f
C4685 vdd.n2437 gnd 0.007409f
C4686 vdd.n2438 gnd 0.007409f
C4687 vdd.n2439 gnd 0.007409f
C4688 vdd.n2440 gnd 0.007409f
C4689 vdd.n2441 gnd 0.007409f
C4690 vdd.n2442 gnd 0.740481f
C4691 vdd.n2443 gnd 0.007409f
C4692 vdd.n2444 gnd 0.007409f
C4693 vdd.n2445 gnd 0.007409f
C4694 vdd.n2446 gnd 0.007409f
C4695 vdd.n2447 gnd 0.007409f
C4696 vdd.n2448 gnd 0.757183f
C4697 vdd.n2449 gnd 0.007409f
C4698 vdd.n2450 gnd 0.007409f
C4699 vdd.n2451 gnd 0.007409f
C4700 vdd.n2452 gnd 0.007409f
C4701 vdd.n2453 gnd 0.007409f
C4702 vdd.n2454 gnd 0.60686f
C4703 vdd.n2455 gnd 0.007409f
C4704 vdd.n2456 gnd 0.007409f
C4705 vdd.n2457 gnd 0.00632f
C4706 vdd.n2458 gnd 0.021463f
C4707 vdd.n2459 gnd 0.004794f
C4708 vdd.n2460 gnd 0.007409f
C4709 vdd.n2461 gnd 0.439835f
C4710 vdd.n2462 gnd 0.007409f
C4711 vdd.n2463 gnd 0.007409f
C4712 vdd.n2464 gnd 0.007409f
C4713 vdd.n2465 gnd 0.007409f
C4714 vdd.n2466 gnd 0.007409f
C4715 vdd.n2467 gnd 0.484375f
C4716 vdd.n2468 gnd 0.007409f
C4717 vdd.n2469 gnd 0.007409f
C4718 vdd.n2470 gnd 0.007409f
C4719 vdd.n2471 gnd 0.007409f
C4720 vdd.n2472 gnd 0.007409f
C4721 vdd.n2473 gnd 0.651401f
C4722 vdd.n2474 gnd 0.007409f
C4723 vdd.n2475 gnd 0.007409f
C4724 vdd.n2476 gnd 0.007409f
C4725 vdd.n2477 gnd 0.007409f
C4726 vdd.n2478 gnd 0.007409f
C4727 vdd.n2479 gnd 0.623563f
C4728 vdd.n2480 gnd 0.007409f
C4729 vdd.n2481 gnd 0.007409f
C4730 vdd.n2482 gnd 0.007409f
C4731 vdd.n2483 gnd 0.007409f
C4732 vdd.n2484 gnd 0.007409f
C4733 vdd.n2485 gnd 0.456537f
C4734 vdd.n2486 gnd 0.007409f
C4735 vdd.n2487 gnd 0.007409f
C4736 vdd.n2488 gnd 0.007409f
C4737 vdd.n2489 gnd 0.007409f
C4738 vdd.n2490 gnd 0.007409f
C4739 vdd.n2491 gnd 0.239404f
C4740 vdd.n2492 gnd 0.007409f
C4741 vdd.n2493 gnd 0.007409f
C4742 vdd.n2494 gnd 0.007409f
C4743 vdd.n2495 gnd 0.007409f
C4744 vdd.n2496 gnd 0.007409f
C4745 vdd.n2497 gnd 0.395294f
C4746 vdd.n2498 gnd 0.007409f
C4747 vdd.n2499 gnd 0.007409f
C4748 vdd.n2500 gnd 0.007409f
C4749 vdd.n2501 gnd 0.007409f
C4750 vdd.n2502 gnd 0.007409f
C4751 vdd.n2503 gnd 0.757183f
C4752 vdd.n2504 gnd 0.007409f
C4753 vdd.n2505 gnd 0.007409f
C4754 vdd.n2506 gnd 0.007409f
C4755 vdd.n2507 gnd 0.007409f
C4756 vdd.n2508 gnd 0.007409f
C4757 vdd.n2509 gnd 0.007409f
C4758 vdd.n2510 gnd 0.007409f
C4759 vdd.n2511 gnd 0.567888f
C4760 vdd.n2512 gnd 0.007409f
C4761 vdd.n2513 gnd 0.007409f
C4762 vdd.n2514 gnd 0.007409f
C4763 vdd.n2515 gnd 0.007409f
C4764 vdd.n2516 gnd 0.007409f
C4765 vdd.n2517 gnd 0.007409f
C4766 vdd.n2518 gnd 0.47324f
C4767 vdd.n2519 gnd 0.007409f
C4768 vdd.n2520 gnd 0.007409f
C4769 vdd.n2521 gnd 0.007409f
C4770 vdd.n2522 gnd 0.01715f
C4771 vdd.n2523 gnd 0.016409f
C4772 vdd.n2524 gnd 0.007409f
C4773 vdd.n2525 gnd 0.007409f
C4774 vdd.n2526 gnd 0.00572f
C4775 vdd.n2527 gnd 0.007409f
C4776 vdd.n2528 gnd 0.007409f
C4777 vdd.n2529 gnd 0.005393f
C4778 vdd.n2530 gnd 0.007409f
C4779 vdd.n2531 gnd 0.007409f
C4780 vdd.n2532 gnd 0.007409f
C4781 vdd.n2533 gnd 0.007409f
C4782 vdd.n2534 gnd 0.007409f
C4783 vdd.n2535 gnd 0.007409f
C4784 vdd.n2536 gnd 0.007409f
C4785 vdd.n2537 gnd 0.007409f
C4786 vdd.n2538 gnd 0.007409f
C4787 vdd.n2539 gnd 0.007409f
C4788 vdd.n2540 gnd 0.007409f
C4789 vdd.n2541 gnd 0.007409f
C4790 vdd.n2542 gnd 0.007409f
C4791 vdd.n2543 gnd 0.007409f
C4792 vdd.n2544 gnd 0.007409f
C4793 vdd.n2545 gnd 0.007409f
C4794 vdd.n2546 gnd 0.007409f
C4795 vdd.n2547 gnd 0.007409f
C4796 vdd.n2548 gnd 0.007409f
C4797 vdd.n2549 gnd 0.007409f
C4798 vdd.n2550 gnd 0.007409f
C4799 vdd.n2551 gnd 0.007409f
C4800 vdd.n2552 gnd 0.007409f
C4801 vdd.n2553 gnd 0.007409f
C4802 vdd.n2554 gnd 0.007409f
C4803 vdd.n2555 gnd 0.007409f
C4804 vdd.n2556 gnd 0.007409f
C4805 vdd.n2557 gnd 0.007409f
C4806 vdd.n2558 gnd 0.007409f
C4807 vdd.n2559 gnd 0.007409f
C4808 vdd.n2560 gnd 0.007409f
C4809 vdd.n2561 gnd 0.007409f
C4810 vdd.n2562 gnd 0.007409f
C4811 vdd.n2563 gnd 0.007409f
C4812 vdd.n2564 gnd 0.007409f
C4813 vdd.n2565 gnd 0.007409f
C4814 vdd.n2566 gnd 0.007409f
C4815 vdd.n2567 gnd 0.007409f
C4816 vdd.n2568 gnd 0.007409f
C4817 vdd.n2569 gnd 0.007409f
C4818 vdd.n2570 gnd 0.007409f
C4819 vdd.n2571 gnd 0.007409f
C4820 vdd.n2572 gnd 0.007409f
C4821 vdd.n2573 gnd 0.007409f
C4822 vdd.n2574 gnd 0.007409f
C4823 vdd.n2575 gnd 0.007409f
C4824 vdd.n2576 gnd 0.007409f
C4825 vdd.n2577 gnd 0.007409f
C4826 vdd.n2578 gnd 0.007409f
C4827 vdd.n2579 gnd 0.007409f
C4828 vdd.n2580 gnd 0.007409f
C4829 vdd.n2581 gnd 0.007409f
C4830 vdd.n2582 gnd 0.007409f
C4831 vdd.n2583 gnd 0.007409f
C4832 vdd.n2584 gnd 0.007409f
C4833 vdd.n2585 gnd 0.007409f
C4834 vdd.n2586 gnd 0.007409f
C4835 vdd.n2587 gnd 0.007409f
C4836 vdd.n2588 gnd 0.007409f
C4837 vdd.n2589 gnd 0.007409f
C4838 vdd.n2590 gnd 0.01733f
C4839 vdd.n2591 gnd 0.01623f
C4840 vdd.n2592 gnd 0.01623f
C4841 vdd.n2593 gnd 0.901939f
C4842 vdd.n2594 gnd 0.01623f
C4843 vdd.n2595 gnd 0.01733f
C4844 vdd.n2596 gnd 0.016409f
C4845 vdd.n2597 gnd 0.007409f
C4846 vdd.n2598 gnd 0.007409f
C4847 vdd.n2599 gnd 0.007409f
C4848 vdd.n2600 gnd 0.00572f
C4849 vdd.n2601 gnd 0.010589f
C4850 vdd.n2602 gnd 0.005393f
C4851 vdd.n2603 gnd 0.007409f
C4852 vdd.n2604 gnd 0.007409f
C4853 vdd.n2605 gnd 0.007409f
C4854 vdd.n2606 gnd 0.007409f
C4855 vdd.n2607 gnd 0.007409f
C4856 vdd.n2608 gnd 0.007409f
C4857 vdd.n2609 gnd 0.007409f
C4858 vdd.n2610 gnd 0.007409f
C4859 vdd.n2611 gnd 0.007409f
C4860 vdd.n2612 gnd 0.007409f
C4861 vdd.n2613 gnd 0.007409f
C4862 vdd.n2614 gnd 0.007409f
C4863 vdd.n2615 gnd 0.007409f
C4864 vdd.n2616 gnd 0.007409f
C4865 vdd.n2617 gnd 0.007409f
C4866 vdd.n2618 gnd 0.007409f
C4867 vdd.n2619 gnd 0.007409f
C4868 vdd.n2620 gnd 0.007409f
C4869 vdd.n2621 gnd 0.007409f
C4870 vdd.n2622 gnd 0.007409f
C4871 vdd.n2623 gnd 0.007409f
C4872 vdd.n2624 gnd 0.007409f
C4873 vdd.n2625 gnd 0.007409f
C4874 vdd.n2626 gnd 0.007409f
C4875 vdd.n2627 gnd 0.007409f
C4876 vdd.n2628 gnd 0.007409f
C4877 vdd.n2629 gnd 0.007409f
C4878 vdd.n2630 gnd 0.007409f
C4879 vdd.n2631 gnd 0.007409f
C4880 vdd.n2632 gnd 0.007409f
C4881 vdd.n2633 gnd 0.007409f
C4882 vdd.n2634 gnd 0.007409f
C4883 vdd.n2635 gnd 0.007409f
C4884 vdd.n2636 gnd 0.007409f
C4885 vdd.n2637 gnd 0.007409f
C4886 vdd.n2638 gnd 0.007409f
C4887 vdd.n2639 gnd 0.007409f
C4888 vdd.n2640 gnd 0.007409f
C4889 vdd.n2641 gnd 0.007409f
C4890 vdd.n2642 gnd 0.007409f
C4891 vdd.n2643 gnd 0.007409f
C4892 vdd.n2644 gnd 0.007409f
C4893 vdd.n2645 gnd 0.007409f
C4894 vdd.n2646 gnd 0.007409f
C4895 vdd.n2647 gnd 0.007409f
C4896 vdd.n2648 gnd 0.007409f
C4897 vdd.n2649 gnd 0.007409f
C4898 vdd.n2650 gnd 0.007409f
C4899 vdd.n2651 gnd 0.007409f
C4900 vdd.n2652 gnd 0.007409f
C4901 vdd.n2653 gnd 0.007409f
C4902 vdd.n2654 gnd 0.007409f
C4903 vdd.n2655 gnd 0.007409f
C4904 vdd.n2656 gnd 0.007409f
C4905 vdd.n2657 gnd 0.007409f
C4906 vdd.n2658 gnd 0.007409f
C4907 vdd.n2659 gnd 0.007409f
C4908 vdd.n2660 gnd 0.007409f
C4909 vdd.n2661 gnd 0.007409f
C4910 vdd.n2662 gnd 0.007409f
C4911 vdd.n2663 gnd 0.01733f
C4912 vdd.n2664 gnd 0.01733f
C4913 vdd.n2665 gnd 0.924209f
C4914 vdd.t10 gnd 3.28484f
C4915 vdd.t46 gnd 3.28484f
C4916 vdd.n2698 gnd 0.01733f
C4917 vdd.t222 gnd 0.690373f
C4918 vdd.n2699 gnd 0.007409f
C4919 vdd.n2700 gnd 0.007409f
C4920 vdd.t276 gnd 0.299404f
C4921 vdd.t277 gnd 0.306477f
C4922 vdd.t274 gnd 0.195462f
C4923 vdd.n2701 gnd 0.105637f
C4924 vdd.n2702 gnd 0.059921f
C4925 vdd.n2703 gnd 0.007409f
C4926 vdd.t289 gnd 0.299404f
C4927 vdd.t290 gnd 0.306477f
C4928 vdd.t288 gnd 0.195462f
C4929 vdd.n2704 gnd 0.105637f
C4930 vdd.n2705 gnd 0.059921f
C4931 vdd.n2706 gnd 0.010589f
C4932 vdd.n2707 gnd 0.007409f
C4933 vdd.n2708 gnd 0.007409f
C4934 vdd.n2709 gnd 0.007409f
C4935 vdd.n2710 gnd 0.007409f
C4936 vdd.n2711 gnd 0.007409f
C4937 vdd.n2712 gnd 0.007409f
C4938 vdd.n2713 gnd 0.007409f
C4939 vdd.n2714 gnd 0.007409f
C4940 vdd.n2715 gnd 0.007409f
C4941 vdd.n2716 gnd 0.007409f
C4942 vdd.n2717 gnd 0.007409f
C4943 vdd.n2718 gnd 0.007409f
C4944 vdd.n2719 gnd 0.007409f
C4945 vdd.n2720 gnd 0.007409f
C4946 vdd.n2721 gnd 0.007409f
C4947 vdd.n2722 gnd 0.007409f
C4948 vdd.n2723 gnd 0.007409f
C4949 vdd.n2724 gnd 0.007409f
C4950 vdd.n2725 gnd 0.007409f
C4951 vdd.n2726 gnd 0.007409f
C4952 vdd.n2727 gnd 0.007409f
C4953 vdd.n2728 gnd 0.007409f
C4954 vdd.n2729 gnd 0.007409f
C4955 vdd.n2730 gnd 0.007409f
C4956 vdd.n2731 gnd 0.007409f
C4957 vdd.n2732 gnd 0.007409f
C4958 vdd.n2733 gnd 0.007409f
C4959 vdd.n2734 gnd 0.007409f
C4960 vdd.n2735 gnd 0.007409f
C4961 vdd.n2736 gnd 0.007409f
C4962 vdd.n2737 gnd 0.007409f
C4963 vdd.n2738 gnd 0.007409f
C4964 vdd.n2739 gnd 0.007409f
C4965 vdd.n2740 gnd 0.007409f
C4966 vdd.n2741 gnd 0.007409f
C4967 vdd.n2742 gnd 0.007409f
C4968 vdd.n2743 gnd 0.007409f
C4969 vdd.n2744 gnd 0.007409f
C4970 vdd.n2745 gnd 0.007409f
C4971 vdd.n2746 gnd 0.007409f
C4972 vdd.n2747 gnd 0.007409f
C4973 vdd.n2748 gnd 0.007409f
C4974 vdd.n2749 gnd 0.007409f
C4975 vdd.n2750 gnd 0.007409f
C4976 vdd.n2751 gnd 0.007409f
C4977 vdd.n2752 gnd 0.007409f
C4978 vdd.n2753 gnd 0.007409f
C4979 vdd.n2754 gnd 0.007409f
C4980 vdd.n2755 gnd 0.007409f
C4981 vdd.n2756 gnd 0.007409f
C4982 vdd.n2757 gnd 0.007409f
C4983 vdd.n2758 gnd 0.007409f
C4984 vdd.n2759 gnd 0.007409f
C4985 vdd.n2760 gnd 0.007409f
C4986 vdd.n2761 gnd 0.007409f
C4987 vdd.n2762 gnd 0.007409f
C4988 vdd.n2763 gnd 0.007409f
C4989 vdd.n2764 gnd 0.007409f
C4990 vdd.n2765 gnd 0.005393f
C4991 vdd.n2766 gnd 0.007409f
C4992 vdd.n2767 gnd 0.007409f
C4993 vdd.n2768 gnd 0.00572f
C4994 vdd.n2769 gnd 0.007409f
C4995 vdd.n2770 gnd 0.007409f
C4996 vdd.n2771 gnd 0.01733f
C4997 vdd.n2772 gnd 0.01623f
C4998 vdd.n2773 gnd 0.01623f
C4999 vdd.n2774 gnd 0.007409f
C5000 vdd.n2775 gnd 0.007409f
C5001 vdd.n2776 gnd 0.007409f
C5002 vdd.n2777 gnd 0.007409f
C5003 vdd.n2778 gnd 0.007409f
C5004 vdd.n2779 gnd 0.007409f
C5005 vdd.n2780 gnd 0.007409f
C5006 vdd.n2781 gnd 0.007409f
C5007 vdd.n2782 gnd 0.007409f
C5008 vdd.n2783 gnd 0.007409f
C5009 vdd.n2784 gnd 0.007409f
C5010 vdd.n2785 gnd 0.007409f
C5011 vdd.n2786 gnd 0.007409f
C5012 vdd.n2787 gnd 0.007409f
C5013 vdd.n2788 gnd 0.007409f
C5014 vdd.n2789 gnd 0.007409f
C5015 vdd.n2790 gnd 0.007409f
C5016 vdd.n2791 gnd 0.007409f
C5017 vdd.n2792 gnd 0.007409f
C5018 vdd.n2793 gnd 0.007409f
C5019 vdd.n2794 gnd 0.007409f
C5020 vdd.n2795 gnd 0.007409f
C5021 vdd.n2796 gnd 0.007409f
C5022 vdd.n2797 gnd 0.007409f
C5023 vdd.n2798 gnd 0.007409f
C5024 vdd.n2799 gnd 0.007409f
C5025 vdd.n2800 gnd 0.007409f
C5026 vdd.n2801 gnd 0.007409f
C5027 vdd.n2802 gnd 0.007409f
C5028 vdd.n2803 gnd 0.007409f
C5029 vdd.n2804 gnd 0.007409f
C5030 vdd.n2805 gnd 0.007409f
C5031 vdd.n2806 gnd 0.007409f
C5032 vdd.n2807 gnd 0.007409f
C5033 vdd.n2808 gnd 0.007409f
C5034 vdd.n2809 gnd 0.007409f
C5035 vdd.n2810 gnd 0.007409f
C5036 vdd.n2811 gnd 0.007409f
C5037 vdd.n2812 gnd 0.007409f
C5038 vdd.n2813 gnd 0.007409f
C5039 vdd.n2814 gnd 0.007409f
C5040 vdd.n2815 gnd 0.007409f
C5041 vdd.n2816 gnd 0.007409f
C5042 vdd.n2817 gnd 0.007409f
C5043 vdd.n2818 gnd 0.007409f
C5044 vdd.n2819 gnd 0.007409f
C5045 vdd.n2820 gnd 0.007409f
C5046 vdd.n2821 gnd 0.007409f
C5047 vdd.n2822 gnd 0.007409f
C5048 vdd.n2823 gnd 0.007409f
C5049 vdd.n2824 gnd 0.007409f
C5050 vdd.n2825 gnd 0.007409f
C5051 vdd.n2826 gnd 0.007409f
C5052 vdd.n2827 gnd 0.007409f
C5053 vdd.n2828 gnd 0.007409f
C5054 vdd.n2829 gnd 0.007409f
C5055 vdd.n2830 gnd 0.007409f
C5056 vdd.n2831 gnd 0.007409f
C5057 vdd.n2832 gnd 0.007409f
C5058 vdd.n2833 gnd 0.007409f
C5059 vdd.n2834 gnd 0.007409f
C5060 vdd.n2835 gnd 0.007409f
C5061 vdd.n2836 gnd 0.007409f
C5062 vdd.n2837 gnd 0.007409f
C5063 vdd.n2838 gnd 0.007409f
C5064 vdd.n2839 gnd 0.007409f
C5065 vdd.n2840 gnd 0.007409f
C5066 vdd.n2841 gnd 0.007409f
C5067 vdd.n2842 gnd 0.007409f
C5068 vdd.n2843 gnd 0.007409f
C5069 vdd.n2844 gnd 0.007409f
C5070 vdd.n2845 gnd 0.007409f
C5071 vdd.n2846 gnd 0.007409f
C5072 vdd.n2847 gnd 0.239404f
C5073 vdd.n2848 gnd 0.007409f
C5074 vdd.n2849 gnd 0.007409f
C5075 vdd.n2850 gnd 0.007409f
C5076 vdd.n2851 gnd 0.007409f
C5077 vdd.n2852 gnd 0.007409f
C5078 vdd.n2853 gnd 0.007409f
C5079 vdd.n2854 gnd 0.007409f
C5080 vdd.n2855 gnd 0.007409f
C5081 vdd.n2856 gnd 0.007409f
C5082 vdd.n2857 gnd 0.007409f
C5083 vdd.n2858 gnd 0.007409f
C5084 vdd.n2859 gnd 0.007409f
C5085 vdd.n2860 gnd 0.007409f
C5086 vdd.n2861 gnd 0.007409f
C5087 vdd.n2862 gnd 0.47324f
C5088 vdd.n2863 gnd 0.007409f
C5089 vdd.n2864 gnd 0.007409f
C5090 vdd.n2865 gnd 0.007409f
C5091 vdd.n2866 gnd 0.01623f
C5092 vdd.n2867 gnd 0.01623f
C5093 vdd.n2868 gnd 0.01733f
C5094 vdd.n2869 gnd 0.01733f
C5095 vdd.n2870 gnd 0.007409f
C5096 vdd.n2871 gnd 0.007409f
C5097 vdd.n2872 gnd 0.007409f
C5098 vdd.n2873 gnd 0.00572f
C5099 vdd.n2874 gnd 0.010589f
C5100 vdd.n2875 gnd 0.005393f
C5101 vdd.n2876 gnd 0.007409f
C5102 vdd.n2877 gnd 0.007409f
C5103 vdd.n2878 gnd 0.007409f
C5104 vdd.n2879 gnd 0.007409f
C5105 vdd.n2880 gnd 0.007409f
C5106 vdd.n2881 gnd 0.007409f
C5107 vdd.n2882 gnd 0.007409f
C5108 vdd.n2883 gnd 0.007409f
C5109 vdd.n2884 gnd 0.007409f
C5110 vdd.n2885 gnd 0.007409f
C5111 vdd.n2886 gnd 0.007409f
C5112 vdd.n2887 gnd 0.007409f
C5113 vdd.n2888 gnd 0.007409f
C5114 vdd.n2889 gnd 0.007409f
C5115 vdd.n2890 gnd 0.007409f
C5116 vdd.n2891 gnd 0.007409f
C5117 vdd.n2892 gnd 0.007409f
C5118 vdd.n2893 gnd 0.007409f
C5119 vdd.n2894 gnd 0.007409f
C5120 vdd.n2895 gnd 0.007409f
C5121 vdd.n2896 gnd 0.007409f
C5122 vdd.n2897 gnd 0.007409f
C5123 vdd.n2898 gnd 0.007409f
C5124 vdd.n2899 gnd 0.007409f
C5125 vdd.n2900 gnd 0.007409f
C5126 vdd.n2901 gnd 0.007409f
C5127 vdd.n2902 gnd 0.007409f
C5128 vdd.n2903 gnd 0.007409f
C5129 vdd.n2904 gnd 0.007409f
C5130 vdd.n2905 gnd 0.007409f
C5131 vdd.n2906 gnd 0.007409f
C5132 vdd.n2907 gnd 0.007409f
C5133 vdd.n2908 gnd 0.007409f
C5134 vdd.n2909 gnd 0.007409f
C5135 vdd.n2910 gnd 0.007409f
C5136 vdd.n2911 gnd 0.007409f
C5137 vdd.n2912 gnd 0.007409f
C5138 vdd.n2913 gnd 0.007409f
C5139 vdd.n2914 gnd 0.007409f
C5140 vdd.n2915 gnd 0.007409f
C5141 vdd.n2916 gnd 0.007409f
C5142 vdd.n2917 gnd 0.007409f
C5143 vdd.n2918 gnd 0.007409f
C5144 vdd.n2919 gnd 0.007409f
C5145 vdd.n2920 gnd 0.007409f
C5146 vdd.n2921 gnd 0.007409f
C5147 vdd.n2922 gnd 0.007409f
C5148 vdd.n2923 gnd 0.007409f
C5149 vdd.n2924 gnd 0.007409f
C5150 vdd.n2925 gnd 0.007409f
C5151 vdd.n2926 gnd 0.007409f
C5152 vdd.n2927 gnd 0.007409f
C5153 vdd.n2928 gnd 0.007409f
C5154 vdd.n2929 gnd 0.007409f
C5155 vdd.n2930 gnd 0.007409f
C5156 vdd.n2931 gnd 0.007409f
C5157 vdd.n2932 gnd 0.007409f
C5158 vdd.n2933 gnd 0.007409f
C5159 vdd.n2934 gnd 0.007409f
C5160 vdd.n2935 gnd 0.01733f
C5161 vdd.n2936 gnd 0.01733f
C5162 vdd.n2938 gnd 0.924209f
C5163 vdd.n2940 gnd 0.01733f
C5164 vdd.n2941 gnd 0.01733f
C5165 vdd.n2942 gnd 0.01623f
C5166 vdd.n2943 gnd 0.007409f
C5167 vdd.n2944 gnd 0.007409f
C5168 vdd.n2945 gnd 0.400862f
C5169 vdd.n2946 gnd 0.007409f
C5170 vdd.n2947 gnd 0.007409f
C5171 vdd.n2948 gnd 0.007409f
C5172 vdd.n2949 gnd 0.007409f
C5173 vdd.n2950 gnd 0.007409f
C5174 vdd.n2951 gnd 0.45097f
C5175 vdd.n2952 gnd 0.007409f
C5176 vdd.n2953 gnd 0.007409f
C5177 vdd.n2954 gnd 0.007409f
C5178 vdd.n2955 gnd 0.007409f
C5179 vdd.n2956 gnd 0.007409f
C5180 vdd.n2957 gnd 0.757183f
C5181 vdd.n2958 gnd 0.007409f
C5182 vdd.n2959 gnd 0.007409f
C5183 vdd.n2960 gnd 0.007409f
C5184 vdd.n2961 gnd 0.007409f
C5185 vdd.n2962 gnd 0.007409f
C5186 vdd.n2963 gnd 0.501077f
C5187 vdd.n2964 gnd 0.007409f
C5188 vdd.n2965 gnd 0.007409f
C5189 vdd.n2966 gnd 0.007409f
C5190 vdd.n2967 gnd 0.007409f
C5191 vdd.n2968 gnd 0.007409f
C5192 vdd.n2969 gnd 0.668103f
C5193 vdd.n2970 gnd 0.007409f
C5194 vdd.n2971 gnd 0.007409f
C5195 vdd.n2972 gnd 0.007409f
C5196 vdd.n2973 gnd 0.007409f
C5197 vdd.n2974 gnd 0.007409f
C5198 vdd.n2975 gnd 0.60686f
C5199 vdd.n2976 gnd 0.007409f
C5200 vdd.n2977 gnd 0.007409f
C5201 vdd.n2978 gnd 0.007409f
C5202 vdd.n2979 gnd 0.007409f
C5203 vdd.n2980 gnd 0.007409f
C5204 vdd.n2981 gnd 0.439835f
C5205 vdd.n2982 gnd 0.007409f
C5206 vdd.n2983 gnd 0.007409f
C5207 vdd.n2984 gnd 0.007409f
C5208 vdd.n2985 gnd 0.007409f
C5209 vdd.n2986 gnd 0.007409f
C5210 vdd.n2987 gnd 0.239404f
C5211 vdd.n2988 gnd 0.007409f
C5212 vdd.n2989 gnd 0.007409f
C5213 vdd.n2990 gnd 0.007409f
C5214 vdd.n2991 gnd 0.007409f
C5215 vdd.n2992 gnd 0.007409f
C5216 vdd.n2993 gnd 0.651401f
C5217 vdd.n2994 gnd 0.007409f
C5218 vdd.n2995 gnd 0.007409f
C5219 vdd.n2996 gnd 0.007409f
C5220 vdd.n2997 gnd 0.007409f
C5221 vdd.n2998 gnd 0.007409f
C5222 vdd.n2999 gnd 0.757183f
C5223 vdd.n3000 gnd 0.007409f
C5224 vdd.n3001 gnd 0.007409f
C5225 vdd.n3002 gnd 0.004794f
C5226 vdd.n3003 gnd 0.021463f
C5227 vdd.n3004 gnd 0.00632f
C5228 vdd.n3005 gnd 0.007409f
C5229 vdd.n3006 gnd 0.645833f
C5230 vdd.n3007 gnd 0.007409f
C5231 vdd.n3008 gnd 0.007409f
C5232 vdd.n3009 gnd 0.007409f
C5233 vdd.n3010 gnd 0.007409f
C5234 vdd.n3011 gnd 0.007409f
C5235 vdd.n3012 gnd 0.528915f
C5236 vdd.n3013 gnd 0.007409f
C5237 vdd.n3014 gnd 0.007409f
C5238 vdd.n3015 gnd 0.007409f
C5239 vdd.n3016 gnd 0.007409f
C5240 vdd.n3017 gnd 0.007409f
C5241 vdd.n3018 gnd 0.395294f
C5242 vdd.n3019 gnd 0.007409f
C5243 vdd.n3020 gnd 0.007409f
C5244 vdd.n3021 gnd 0.007409f
C5245 vdd.n3022 gnd 0.007409f
C5246 vdd.n3023 gnd 0.007409f
C5247 vdd.n3024 gnd 0.757183f
C5248 vdd.n3025 gnd 0.007409f
C5249 vdd.n3026 gnd 0.007409f
C5250 vdd.n3027 gnd 0.007409f
C5251 vdd.n3028 gnd 0.007409f
C5252 vdd.n3029 gnd 0.007409f
C5253 vdd.n3030 gnd 0.007409f
C5254 vdd.n3032 gnd 0.007409f
C5255 vdd.n3033 gnd 0.007409f
C5256 vdd.n3035 gnd 0.007409f
C5257 vdd.n3036 gnd 0.007409f
C5258 vdd.n3039 gnd 0.007409f
C5259 vdd.n3040 gnd 0.007409f
C5260 vdd.n3041 gnd 0.007409f
C5261 vdd.n3042 gnd 0.007409f
C5262 vdd.n3044 gnd 0.007409f
C5263 vdd.n3045 gnd 0.007409f
C5264 vdd.n3046 gnd 0.007409f
C5265 vdd.n3047 gnd 0.007409f
C5266 vdd.n3048 gnd 0.007409f
C5267 vdd.n3049 gnd 0.007409f
C5268 vdd.n3051 gnd 0.007409f
C5269 vdd.n3052 gnd 0.007409f
C5270 vdd.n3053 gnd 0.007409f
C5271 vdd.n3054 gnd 0.007409f
C5272 vdd.n3055 gnd 0.007409f
C5273 vdd.n3056 gnd 0.007409f
C5274 vdd.n3058 gnd 0.007409f
C5275 vdd.n3059 gnd 0.007409f
C5276 vdd.n3060 gnd 0.007409f
C5277 vdd.n3061 gnd 0.007409f
C5278 vdd.n3062 gnd 0.007409f
C5279 vdd.n3063 gnd 0.007409f
C5280 vdd.n3065 gnd 0.007409f
C5281 vdd.n3066 gnd 0.01733f
C5282 vdd.n3067 gnd 0.01733f
C5283 vdd.n3068 gnd 0.01623f
C5284 vdd.n3069 gnd 0.007409f
C5285 vdd.n3070 gnd 0.007409f
C5286 vdd.n3071 gnd 0.007409f
C5287 vdd.n3072 gnd 0.007409f
C5288 vdd.n3073 gnd 0.007409f
C5289 vdd.n3074 gnd 0.007409f
C5290 vdd.n3075 gnd 0.757183f
C5291 vdd.n3076 gnd 0.007409f
C5292 vdd.n3077 gnd 0.007409f
C5293 vdd.n3078 gnd 0.007409f
C5294 vdd.n3079 gnd 0.007409f
C5295 vdd.n3080 gnd 0.007409f
C5296 vdd.n3081 gnd 0.49551f
C5297 vdd.n3082 gnd 0.007409f
C5298 vdd.n3083 gnd 0.007409f
C5299 vdd.n3084 gnd 0.007409f
C5300 vdd.n3085 gnd 0.01715f
C5301 vdd.n3086 gnd 0.016409f
C5302 vdd.n3087 gnd 0.01733f
C5303 vdd.n3089 gnd 0.007409f
C5304 vdd.n3090 gnd 0.007409f
C5305 vdd.n3091 gnd 0.00572f
C5306 vdd.n3092 gnd 0.010589f
C5307 vdd.n3093 gnd 0.005393f
C5308 vdd.n3094 gnd 0.007409f
C5309 vdd.n3095 gnd 0.007409f
C5310 vdd.n3097 gnd 0.007409f
C5311 vdd.n3098 gnd 0.007409f
C5312 vdd.n3099 gnd 0.007409f
C5313 vdd.n3100 gnd 0.007409f
C5314 vdd.n3101 gnd 0.007409f
C5315 vdd.n3102 gnd 0.007409f
C5316 vdd.n3104 gnd 0.007409f
C5317 vdd.n3105 gnd 0.007409f
C5318 vdd.n3106 gnd 0.007409f
C5319 vdd.n3107 gnd 0.007409f
C5320 vdd.n3108 gnd 0.007409f
C5321 vdd.n3109 gnd 0.007409f
C5322 vdd.n3111 gnd 0.007409f
C5323 vdd.n3112 gnd 0.007409f
C5324 vdd.n3113 gnd 0.007409f
C5325 vdd.n3114 gnd 0.007409f
C5326 vdd.n3115 gnd 0.007409f
C5327 vdd.n3116 gnd 0.007409f
C5328 vdd.n3118 gnd 0.007409f
C5329 vdd.n3119 gnd 0.007409f
C5330 vdd.n3120 gnd 0.007409f
C5331 vdd.n3122 gnd 0.007409f
C5332 vdd.n3123 gnd 0.007409f
C5333 vdd.n3124 gnd 0.007409f
C5334 vdd.n3125 gnd 0.007409f
C5335 vdd.n3126 gnd 0.007409f
C5336 vdd.n3127 gnd 0.007409f
C5337 vdd.n3129 gnd 0.007409f
C5338 vdd.n3130 gnd 0.007409f
C5339 vdd.n3131 gnd 0.007409f
C5340 vdd.n3132 gnd 0.007409f
C5341 vdd.n3133 gnd 0.007409f
C5342 vdd.n3134 gnd 0.007409f
C5343 vdd.n3136 gnd 0.007409f
C5344 vdd.n3137 gnd 0.007409f
C5345 vdd.n3138 gnd 0.007409f
C5346 vdd.n3139 gnd 0.007409f
C5347 vdd.n3140 gnd 0.007409f
C5348 vdd.n3141 gnd 0.007409f
C5349 vdd.n3143 gnd 0.007409f
C5350 vdd.n3144 gnd 0.007409f
C5351 vdd.n3146 gnd 0.007409f
C5352 vdd.n3147 gnd 0.007409f
C5353 vdd.n3148 gnd 0.01733f
C5354 vdd.n3149 gnd 0.01623f
C5355 vdd.n3150 gnd 0.01623f
C5356 vdd.n3151 gnd 1.06896f
C5357 vdd.n3152 gnd 0.01623f
C5358 vdd.n3153 gnd 0.01733f
C5359 vdd.n3154 gnd 0.016409f
C5360 vdd.n3155 gnd 0.007409f
C5361 vdd.n3156 gnd 0.00572f
C5362 vdd.n3157 gnd 0.007409f
C5363 vdd.n3159 gnd 0.007409f
C5364 vdd.n3160 gnd 0.007409f
C5365 vdd.n3161 gnd 0.007409f
C5366 vdd.n3162 gnd 0.007409f
C5367 vdd.n3163 gnd 0.007409f
C5368 vdd.n3164 gnd 0.007409f
C5369 vdd.n3166 gnd 0.007409f
C5370 vdd.n3167 gnd 0.007409f
C5371 vdd.n3168 gnd 0.007409f
C5372 vdd.n3169 gnd 0.007409f
C5373 vdd.n3170 gnd 0.007409f
C5374 vdd.n3171 gnd 0.007409f
C5375 vdd.n3173 gnd 0.007409f
C5376 vdd.n3174 gnd 0.007409f
C5377 vdd.n3175 gnd 0.007409f
C5378 vdd.n3176 gnd 0.007409f
C5379 vdd.n3177 gnd 0.007409f
C5380 vdd.n3178 gnd 0.007409f
C5381 vdd.n3180 gnd 0.007409f
C5382 vdd.n3181 gnd 0.007409f
C5383 vdd.n3183 gnd 0.007409f
C5384 vdd.n3184 gnd 0.025446f
C5385 vdd.n3185 gnd 0.828254f
C5386 vdd.n3187 gnd 0.004604f
C5387 vdd.n3188 gnd 0.00877f
C5388 vdd.n3189 gnd 0.010896f
C5389 vdd.n3190 gnd 0.010896f
C5390 vdd.n3191 gnd 0.00877f
C5391 vdd.n3192 gnd 0.00877f
C5392 vdd.n3193 gnd 0.010896f
C5393 vdd.n3194 gnd 0.010896f
C5394 vdd.n3195 gnd 0.00877f
C5395 vdd.n3196 gnd 0.00877f
C5396 vdd.n3197 gnd 0.010896f
C5397 vdd.n3198 gnd 0.010896f
C5398 vdd.n3199 gnd 0.00877f
C5399 vdd.n3200 gnd 0.00877f
C5400 vdd.n3201 gnd 0.010896f
C5401 vdd.n3202 gnd 0.010896f
C5402 vdd.n3203 gnd 0.00877f
C5403 vdd.n3204 gnd 0.00877f
C5404 vdd.n3205 gnd 0.010896f
C5405 vdd.n3206 gnd 0.010896f
C5406 vdd.n3207 gnd 0.00877f
C5407 vdd.n3208 gnd 0.00877f
C5408 vdd.n3209 gnd 0.010896f
C5409 vdd.n3210 gnd 0.010896f
C5410 vdd.n3211 gnd 0.00877f
C5411 vdd.n3212 gnd 0.00877f
C5412 vdd.n3213 gnd 0.010896f
C5413 vdd.n3214 gnd 0.010896f
C5414 vdd.n3215 gnd 0.00877f
C5415 vdd.n3216 gnd 0.00877f
C5416 vdd.n3217 gnd 0.010896f
C5417 vdd.n3218 gnd 0.010896f
C5418 vdd.n3219 gnd 0.00877f
C5419 vdd.n3220 gnd 0.00877f
C5420 vdd.n3221 gnd 0.010896f
C5421 vdd.n3222 gnd 0.010896f
C5422 vdd.n3223 gnd 0.00877f
C5423 vdd.n3224 gnd 0.010896f
C5424 vdd.n3225 gnd 0.010896f
C5425 vdd.n3226 gnd 0.00877f
C5426 vdd.n3227 gnd 0.010896f
C5427 vdd.n3228 gnd 0.010896f
C5428 vdd.n3229 gnd 0.010896f
C5429 vdd.n3230 gnd 0.01789f
C5430 vdd.n3231 gnd 0.010896f
C5431 vdd.n3232 gnd 0.010896f
C5432 vdd.n3233 gnd 0.005964f
C5433 vdd.n3234 gnd 0.00877f
C5434 vdd.n3235 gnd 0.010896f
C5435 vdd.n3236 gnd 0.010896f
C5436 vdd.n3237 gnd 0.00877f
C5437 vdd.n3238 gnd 0.00877f
C5438 vdd.n3239 gnd 0.010896f
C5439 vdd.n3240 gnd 0.010896f
C5440 vdd.n3241 gnd 0.00877f
C5441 vdd.n3242 gnd 0.00877f
C5442 vdd.n3243 gnd 0.010896f
C5443 vdd.n3244 gnd 0.010896f
C5444 vdd.n3245 gnd 0.00877f
C5445 vdd.n3246 gnd 0.00877f
C5446 vdd.n3247 gnd 0.010896f
C5447 vdd.n3248 gnd 0.010896f
C5448 vdd.n3249 gnd 0.00877f
C5449 vdd.n3250 gnd 0.00877f
C5450 vdd.n3251 gnd 0.010896f
C5451 vdd.n3252 gnd 0.010896f
C5452 vdd.n3253 gnd 0.00877f
C5453 vdd.n3254 gnd 0.00877f
C5454 vdd.n3255 gnd 0.010896f
C5455 vdd.n3256 gnd 0.010896f
C5456 vdd.n3257 gnd 0.00877f
C5457 vdd.n3258 gnd 0.00877f
C5458 vdd.n3259 gnd 0.010896f
C5459 vdd.n3260 gnd 0.010896f
C5460 vdd.n3261 gnd 0.00877f
C5461 vdd.n3262 gnd 0.00877f
C5462 vdd.n3263 gnd 0.010896f
C5463 vdd.n3264 gnd 0.010896f
C5464 vdd.n3265 gnd 0.00877f
C5465 vdd.n3266 gnd 0.00877f
C5466 vdd.n3267 gnd 0.010896f
C5467 vdd.n3268 gnd 0.010896f
C5468 vdd.n3269 gnd 0.00877f
C5469 vdd.n3270 gnd 0.010896f
C5470 vdd.n3271 gnd 0.010896f
C5471 vdd.n3272 gnd 0.00877f
C5472 vdd.n3273 gnd 0.010896f
C5473 vdd.n3274 gnd 0.010896f
C5474 vdd.n3275 gnd 0.010896f
C5475 vdd.t255 gnd 0.134048f
C5476 vdd.t256 gnd 0.14326f
C5477 vdd.t254 gnd 0.175065f
C5478 vdd.n3276 gnd 0.224408f
C5479 vdd.n3277 gnd 0.188543f
C5480 vdd.n3278 gnd 0.01789f
C5481 vdd.n3279 gnd 0.010896f
C5482 vdd.n3280 gnd 0.010896f
C5483 vdd.n3281 gnd 0.007323f
C5484 vdd.n3282 gnd 0.00877f
C5485 vdd.n3283 gnd 0.010896f
C5486 vdd.n3284 gnd 0.010896f
C5487 vdd.n3285 gnd 0.00877f
C5488 vdd.n3286 gnd 0.00877f
C5489 vdd.n3287 gnd 0.010896f
C5490 vdd.n3288 gnd 0.010896f
C5491 vdd.n3289 gnd 0.00877f
C5492 vdd.n3290 gnd 0.00877f
C5493 vdd.n3291 gnd 0.010896f
C5494 vdd.n3292 gnd 0.010896f
C5495 vdd.n3293 gnd 0.00877f
C5496 vdd.n3294 gnd 0.00877f
C5497 vdd.n3295 gnd 0.010896f
C5498 vdd.n3296 gnd 0.010896f
C5499 vdd.n3297 gnd 0.00877f
C5500 vdd.n3298 gnd 0.00877f
C5501 vdd.n3299 gnd 0.010896f
C5502 vdd.n3300 gnd 0.010896f
C5503 vdd.n3301 gnd 0.00877f
C5504 vdd.n3302 gnd 0.00877f
C5505 vdd.n3303 gnd 0.010896f
C5506 vdd.n3304 gnd 0.010896f
C5507 vdd.n3305 gnd 0.00877f
C5508 vdd.n3306 gnd 0.00877f
C5509 vdd.n3308 gnd 0.828254f
C5510 vdd.n3310 gnd 0.00877f
C5511 vdd.n3311 gnd 0.00877f
C5512 vdd.n3312 gnd 0.007279f
C5513 vdd.n3313 gnd 0.026923f
C5514 vdd.n3315 gnd 9.899059f
C5515 vdd.n3316 gnd 0.026923f
C5516 vdd.n3317 gnd 0.004166f
C5517 vdd.n3318 gnd 0.026923f
C5518 vdd.n3319 gnd 0.026358f
C5519 vdd.n3320 gnd 0.010896f
C5520 vdd.n3321 gnd 0.00877f
C5521 vdd.n3322 gnd 0.010896f
C5522 vdd.n3323 gnd 0.673671f
C5523 vdd.n3324 gnd 0.010896f
C5524 vdd.n3325 gnd 0.00877f
C5525 vdd.n3326 gnd 0.010896f
C5526 vdd.n3327 gnd 0.010896f
C5527 vdd.n3328 gnd 0.010896f
C5528 vdd.n3329 gnd 0.00877f
C5529 vdd.n3330 gnd 0.010896f
C5530 vdd.n3331 gnd 1.11351f
C5531 vdd.n3332 gnd 0.010896f
C5532 vdd.n3333 gnd 0.00877f
C5533 vdd.n3334 gnd 0.010896f
C5534 vdd.n3335 gnd 0.010896f
C5535 vdd.n3336 gnd 0.010896f
C5536 vdd.n3337 gnd 0.00877f
C5537 vdd.n3338 gnd 0.010896f
C5538 vdd.n3339 gnd 0.718211f
C5539 vdd.n3340 gnd 0.762751f
C5540 vdd.n3341 gnd 0.010896f
C5541 vdd.n3342 gnd 0.00877f
C5542 vdd.n3343 gnd 0.010896f
C5543 vdd.n3344 gnd 0.010896f
C5544 vdd.n3345 gnd 0.010896f
C5545 vdd.n3346 gnd 0.00877f
C5546 vdd.n3347 gnd 0.010896f
C5547 vdd.n3348 gnd 0.924209f
C5548 vdd.n3349 gnd 0.010896f
C5549 vdd.n3350 gnd 0.00877f
C5550 vdd.n3351 gnd 0.010896f
C5551 vdd.n3352 gnd 0.010896f
C5552 vdd.n3353 gnd 0.010896f
C5553 vdd.n3354 gnd 0.00877f
C5554 vdd.n3355 gnd 0.010896f
C5555 vdd.t124 gnd 0.556753f
C5556 vdd.n3356 gnd 0.896372f
C5557 vdd.n3357 gnd 0.010896f
C5558 vdd.n3358 gnd 0.00877f
C5559 vdd.n3359 gnd 0.010896f
C5560 vdd.n3360 gnd 0.010896f
C5561 vdd.n3361 gnd 0.010896f
C5562 vdd.n3362 gnd 0.00877f
C5563 vdd.n3363 gnd 0.010896f
C5564 vdd.n3364 gnd 0.707076f
C5565 vdd.n3365 gnd 0.010896f
C5566 vdd.n3366 gnd 0.00877f
C5567 vdd.n3367 gnd 0.010896f
C5568 vdd.n3368 gnd 0.010896f
C5569 vdd.n3369 gnd 0.010896f
C5570 vdd.n3370 gnd 0.00877f
C5571 vdd.n3371 gnd 0.010896f
C5572 vdd.n3372 gnd 0.885237f
C5573 vdd.n3373 gnd 0.595725f
C5574 vdd.n3374 gnd 0.010896f
C5575 vdd.n3375 gnd 0.00877f
C5576 vdd.n3376 gnd 0.010896f
C5577 vdd.n3377 gnd 0.010896f
C5578 vdd.n3378 gnd 0.010896f
C5579 vdd.n3379 gnd 0.00877f
C5580 vdd.n3380 gnd 0.010896f
C5581 vdd.n3381 gnd 0.785021f
C5582 vdd.n3382 gnd 0.010896f
C5583 vdd.n3383 gnd 0.00877f
C5584 vdd.n3384 gnd 0.010896f
C5585 vdd.n3385 gnd 0.010896f
C5586 vdd.n3386 gnd 0.010896f
C5587 vdd.n3387 gnd 0.010896f
C5588 vdd.n3388 gnd 0.010896f
C5589 vdd.n3389 gnd 0.00877f
C5590 vdd.n3390 gnd 0.00877f
C5591 vdd.n3391 gnd 0.010896f
C5592 vdd.t153 gnd 0.556753f
C5593 vdd.n3392 gnd 0.924209f
C5594 vdd.n3393 gnd 0.010896f
C5595 vdd.n3394 gnd 0.00877f
C5596 vdd.n3395 gnd 0.010896f
C5597 vdd.n3396 gnd 0.010896f
C5598 vdd.n3397 gnd 0.010896f
C5599 vdd.n3398 gnd 0.00877f
C5600 vdd.n3399 gnd 0.010896f
C5601 vdd.n3400 gnd 0.874102f
C5602 vdd.n3401 gnd 0.010896f
C5603 vdd.n3402 gnd 0.010896f
C5604 vdd.n3403 gnd 0.00877f
C5605 vdd.n3404 gnd 0.00877f
C5606 vdd.n3405 gnd 0.010896f
C5607 vdd.n3406 gnd 0.010896f
C5608 vdd.n3407 gnd 0.010896f
C5609 vdd.n3408 gnd 0.00877f
C5610 vdd.n3409 gnd 0.010896f
C5611 vdd.n3410 gnd 0.00877f
C5612 vdd.n3411 gnd 0.00877f
C5613 vdd.n3412 gnd 0.010896f
C5614 vdd.n3413 gnd 0.010896f
C5615 vdd.n3414 gnd 0.010896f
C5616 vdd.n3415 gnd 0.00877f
C5617 vdd.n3416 gnd 0.010896f
C5618 vdd.n3417 gnd 0.00877f
C5619 vdd.n3418 gnd 0.00877f
C5620 vdd.n3419 gnd 0.010896f
C5621 vdd.n3420 gnd 0.010896f
C5622 vdd.n3421 gnd 0.010896f
C5623 vdd.n3422 gnd 0.00877f
C5624 vdd.n3423 gnd 0.924209f
C5625 vdd.n3424 gnd 0.010896f
C5626 vdd.n3425 gnd 0.00877f
C5627 vdd.n3426 gnd 0.00877f
C5628 vdd.n3427 gnd 0.010896f
C5629 vdd.n3428 gnd 0.010896f
C5630 vdd.n3429 gnd 0.010896f
C5631 vdd.n3430 gnd 0.00877f
C5632 vdd.n3431 gnd 0.010896f
C5633 vdd.n3432 gnd 0.00877f
C5634 vdd.n3433 gnd 0.00877f
C5635 vdd.n3434 gnd 0.010896f
C5636 vdd.n3435 gnd 0.010896f
C5637 vdd.n3436 gnd 0.010896f
C5638 vdd.n3437 gnd 0.00877f
C5639 vdd.n3438 gnd 0.010896f
C5640 vdd.n3439 gnd 0.00877f
C5641 vdd.n3440 gnd 0.007279f
C5642 vdd.n3441 gnd 0.026358f
C5643 vdd.n3442 gnd 0.026923f
C5644 vdd.n3443 gnd 0.004166f
C5645 vdd.n3444 gnd 0.026923f
C5646 vdd.n3446 gnd 2.63901f
C5647 vdd.n3447 gnd 1.64242f
C5648 vdd.n3448 gnd 0.026358f
C5649 vdd.n3449 gnd 0.007279f
C5650 vdd.n3450 gnd 0.00877f
C5651 vdd.n3451 gnd 0.00877f
C5652 vdd.n3452 gnd 0.010896f
C5653 vdd.n3453 gnd 1.11351f
C5654 vdd.n3454 gnd 1.11351f
C5655 vdd.n3455 gnd 1.01886f
C5656 vdd.n3456 gnd 0.010896f
C5657 vdd.n3457 gnd 0.00877f
C5658 vdd.n3458 gnd 0.00877f
C5659 vdd.n3459 gnd 0.00877f
C5660 vdd.n3460 gnd 0.010896f
C5661 vdd.n3461 gnd 0.829561f
C5662 vdd.t181 gnd 0.556753f
C5663 vdd.n3462 gnd 0.840696f
C5664 vdd.n3463 gnd 0.640265f
C5665 vdd.n3464 gnd 0.010896f
C5666 vdd.n3465 gnd 0.00877f
C5667 vdd.n3466 gnd 0.00877f
C5668 vdd.n3467 gnd 0.00877f
C5669 vdd.n3468 gnd 0.010896f
C5670 vdd.n3469 gnd 0.662536f
C5671 vdd.n3470 gnd 0.818426f
C5672 vdd.t135 gnd 0.556753f
C5673 vdd.n3471 gnd 0.851831f
C5674 vdd.n3472 gnd 0.010896f
C5675 vdd.n3473 gnd 0.00877f
C5676 vdd.n3474 gnd 0.00877f
C5677 vdd.n3475 gnd 0.00877f
C5678 vdd.n3476 gnd 0.010896f
C5679 vdd.n3477 gnd 0.924209f
C5680 vdd.t85 gnd 0.556753f
C5681 vdd.n3478 gnd 0.673671f
C5682 vdd.n3479 gnd 0.807291f
C5683 vdd.n3480 gnd 0.010896f
C5684 vdd.n3481 gnd 0.00877f
C5685 vdd.n3482 gnd 0.00877f
C5686 vdd.n3483 gnd 0.00877f
C5687 vdd.n3484 gnd 0.010896f
C5688 vdd.n3485 gnd 0.617995f
C5689 vdd.t97 gnd 0.556753f
C5690 vdd.n3486 gnd 0.924209f
C5691 vdd.t89 gnd 0.556753f
C5692 vdd.n3487 gnd 0.684806f
C5693 vdd.n3488 gnd 0.010896f
C5694 vdd.n3489 gnd 0.00877f
C5695 vdd.n3490 gnd 0.008374f
C5696 vdd.n3491 gnd 0.642679f
C5697 vdd.n3492 gnd 2.91814f
C5698 a_n8300_8799.n0 gnd 0.209848f
C5699 a_n8300_8799.n1 gnd 0.288148f
C5700 a_n8300_8799.n2 gnd 0.209848f
C5701 a_n8300_8799.n3 gnd 0.209848f
C5702 a_n8300_8799.n4 gnd 0.209848f
C5703 a_n8300_8799.n5 gnd 0.209848f
C5704 a_n8300_8799.n6 gnd 0.209848f
C5705 a_n8300_8799.n7 gnd 0.218204f
C5706 a_n8300_8799.n8 gnd 0.209848f
C5707 a_n8300_8799.n9 gnd 0.288148f
C5708 a_n8300_8799.n10 gnd 0.209848f
C5709 a_n8300_8799.n11 gnd 0.209848f
C5710 a_n8300_8799.n12 gnd 0.209848f
C5711 a_n8300_8799.n13 gnd 0.209848f
C5712 a_n8300_8799.n14 gnd 0.209848f
C5713 a_n8300_8799.n15 gnd 0.218204f
C5714 a_n8300_8799.n16 gnd 0.209848f
C5715 a_n8300_8799.n17 gnd 0.454831f
C5716 a_n8300_8799.n18 gnd 0.209848f
C5717 a_n8300_8799.n19 gnd 0.209848f
C5718 a_n8300_8799.n20 gnd 0.209848f
C5719 a_n8300_8799.n21 gnd 0.209848f
C5720 a_n8300_8799.n22 gnd 0.209848f
C5721 a_n8300_8799.n23 gnd 0.218204f
C5722 a_n8300_8799.n24 gnd 0.209848f
C5723 a_n8300_8799.n25 gnd 0.323128f
C5724 a_n8300_8799.n26 gnd 0.209848f
C5725 a_n8300_8799.n27 gnd 0.209848f
C5726 a_n8300_8799.n28 gnd 0.209848f
C5727 a_n8300_8799.n29 gnd 0.209848f
C5728 a_n8300_8799.n30 gnd 0.209848f
C5729 a_n8300_8799.n31 gnd 0.183225f
C5730 a_n8300_8799.n32 gnd 0.209848f
C5731 a_n8300_8799.n33 gnd 0.323128f
C5732 a_n8300_8799.n34 gnd 0.209848f
C5733 a_n8300_8799.n35 gnd 0.209848f
C5734 a_n8300_8799.n36 gnd 0.209848f
C5735 a_n8300_8799.n37 gnd 0.209848f
C5736 a_n8300_8799.n38 gnd 0.209848f
C5737 a_n8300_8799.n39 gnd 0.183225f
C5738 a_n8300_8799.n40 gnd 0.209848f
C5739 a_n8300_8799.n41 gnd 0.323128f
C5740 a_n8300_8799.n42 gnd 0.209848f
C5741 a_n8300_8799.n43 gnd 0.209848f
C5742 a_n8300_8799.n44 gnd 0.209848f
C5743 a_n8300_8799.n45 gnd 0.209848f
C5744 a_n8300_8799.n46 gnd 0.209848f
C5745 a_n8300_8799.n47 gnd 0.349908f
C5746 a_n8300_8799.n48 gnd 0.706493f
C5747 a_n8300_8799.n49 gnd 2.93f
C5748 a_n8300_8799.n50 gnd 2.87273f
C5749 a_n8300_8799.n51 gnd 1.4102f
C5750 a_n8300_8799.n52 gnd 1.53802f
C5751 a_n8300_8799.n53 gnd 1.03021f
C5752 a_n8300_8799.n54 gnd 2.58982f
C5753 a_n8300_8799.n55 gnd 0.252637f
C5754 a_n8300_8799.n56 gnd 0.003693f
C5755 a_n8300_8799.n57 gnd 0.009736f
C5756 a_n8300_8799.n58 gnd 0.010637f
C5757 a_n8300_8799.n59 gnd 0.005621f
C5758 a_n8300_8799.n61 gnd 0.004716f
C5759 a_n8300_8799.n62 gnd 0.010201f
C5760 a_n8300_8799.n63 gnd 0.010201f
C5761 a_n8300_8799.n64 gnd 0.004716f
C5762 a_n8300_8799.n66 gnd 0.005621f
C5763 a_n8300_8799.n67 gnd 0.010637f
C5764 a_n8300_8799.n68 gnd 0.009736f
C5765 a_n8300_8799.n69 gnd 0.003693f
C5766 a_n8300_8799.n70 gnd 0.252637f
C5767 a_n8300_8799.n71 gnd 0.003693f
C5768 a_n8300_8799.n72 gnd 0.009736f
C5769 a_n8300_8799.n73 gnd 0.010637f
C5770 a_n8300_8799.n74 gnd 0.005621f
C5771 a_n8300_8799.n76 gnd 0.004716f
C5772 a_n8300_8799.n77 gnd 0.010201f
C5773 a_n8300_8799.n78 gnd 0.010201f
C5774 a_n8300_8799.n79 gnd 0.004716f
C5775 a_n8300_8799.n81 gnd 0.005621f
C5776 a_n8300_8799.n82 gnd 0.010637f
C5777 a_n8300_8799.n83 gnd 0.009736f
C5778 a_n8300_8799.n84 gnd 0.003693f
C5779 a_n8300_8799.n85 gnd 0.252637f
C5780 a_n8300_8799.n86 gnd 0.003693f
C5781 a_n8300_8799.n87 gnd 0.009736f
C5782 a_n8300_8799.n88 gnd 0.010637f
C5783 a_n8300_8799.n89 gnd 0.005621f
C5784 a_n8300_8799.n91 gnd 0.004716f
C5785 a_n8300_8799.n92 gnd 0.010201f
C5786 a_n8300_8799.n93 gnd 0.010201f
C5787 a_n8300_8799.n94 gnd 0.004716f
C5788 a_n8300_8799.n96 gnd 0.005621f
C5789 a_n8300_8799.n97 gnd 0.010637f
C5790 a_n8300_8799.n98 gnd 0.009736f
C5791 a_n8300_8799.n99 gnd 0.003693f
C5792 a_n8300_8799.n100 gnd 0.003693f
C5793 a_n8300_8799.n101 gnd 0.009736f
C5794 a_n8300_8799.n102 gnd 0.010637f
C5795 a_n8300_8799.n103 gnd 0.005621f
C5796 a_n8300_8799.n105 gnd 0.004716f
C5797 a_n8300_8799.n106 gnd 0.010201f
C5798 a_n8300_8799.n107 gnd 0.010201f
C5799 a_n8300_8799.n108 gnd 0.004716f
C5800 a_n8300_8799.n110 gnd 0.005621f
C5801 a_n8300_8799.n111 gnd 0.010637f
C5802 a_n8300_8799.n112 gnd 0.009736f
C5803 a_n8300_8799.n113 gnd 0.003693f
C5804 a_n8300_8799.n114 gnd 0.252637f
C5805 a_n8300_8799.n115 gnd 0.003693f
C5806 a_n8300_8799.n116 gnd 0.009736f
C5807 a_n8300_8799.n117 gnd 0.010637f
C5808 a_n8300_8799.n118 gnd 0.005621f
C5809 a_n8300_8799.n120 gnd 0.004716f
C5810 a_n8300_8799.n121 gnd 0.010201f
C5811 a_n8300_8799.n122 gnd 0.010201f
C5812 a_n8300_8799.n123 gnd 0.004716f
C5813 a_n8300_8799.n125 gnd 0.005621f
C5814 a_n8300_8799.n126 gnd 0.010637f
C5815 a_n8300_8799.n127 gnd 0.009736f
C5816 a_n8300_8799.n128 gnd 0.003693f
C5817 a_n8300_8799.n129 gnd 0.252637f
C5818 a_n8300_8799.n130 gnd 0.003693f
C5819 a_n8300_8799.n131 gnd 0.009736f
C5820 a_n8300_8799.n132 gnd 0.010637f
C5821 a_n8300_8799.n133 gnd 0.005621f
C5822 a_n8300_8799.n135 gnd 0.004716f
C5823 a_n8300_8799.n136 gnd 0.010201f
C5824 a_n8300_8799.n137 gnd 0.010201f
C5825 a_n8300_8799.n138 gnd 0.004716f
C5826 a_n8300_8799.n140 gnd 0.005621f
C5827 a_n8300_8799.n141 gnd 0.010637f
C5828 a_n8300_8799.n142 gnd 0.009736f
C5829 a_n8300_8799.n143 gnd 0.003693f
C5830 a_n8300_8799.n144 gnd 0.252637f
C5831 a_n8300_8799.t12 gnd 0.145553f
C5832 a_n8300_8799.t11 gnd 0.145553f
C5833 a_n8300_8799.t29 gnd 0.145553f
C5834 a_n8300_8799.n145 gnd 1.148f
C5835 a_n8300_8799.t32 gnd 0.145553f
C5836 a_n8300_8799.t22 gnd 0.145553f
C5837 a_n8300_8799.n146 gnd 1.1461f
C5838 a_n8300_8799.t7 gnd 0.145553f
C5839 a_n8300_8799.t19 gnd 0.145553f
C5840 a_n8300_8799.n147 gnd 1.1461f
C5841 a_n8300_8799.t17 gnd 0.145553f
C5842 a_n8300_8799.t2 gnd 0.145553f
C5843 a_n8300_8799.n148 gnd 1.14799f
C5844 a_n8300_8799.t23 gnd 0.145553f
C5845 a_n8300_8799.t28 gnd 0.145553f
C5846 a_n8300_8799.n149 gnd 1.1461f
C5847 a_n8300_8799.t13 gnd 0.145553f
C5848 a_n8300_8799.t20 gnd 0.145553f
C5849 a_n8300_8799.n150 gnd 1.1461f
C5850 a_n8300_8799.t18 gnd 0.145553f
C5851 a_n8300_8799.t21 gnd 0.145553f
C5852 a_n8300_8799.n151 gnd 1.1461f
C5853 a_n8300_8799.n152 gnd 3.19906f
C5854 a_n8300_8799.t25 gnd 0.113208f
C5855 a_n8300_8799.t30 gnd 0.113208f
C5856 a_n8300_8799.n153 gnd 1.00194f
C5857 a_n8300_8799.t24 gnd 0.113208f
C5858 a_n8300_8799.t0 gnd 0.113208f
C5859 a_n8300_8799.n154 gnd 1.00034f
C5860 a_n8300_8799.t14 gnd 0.113208f
C5861 a_n8300_8799.t4 gnd 0.113208f
C5862 a_n8300_8799.n155 gnd 1.00034f
C5863 a_n8300_8799.t3 gnd 0.113208f
C5864 a_n8300_8799.t16 gnd 0.113208f
C5865 a_n8300_8799.n156 gnd 1.00194f
C5866 a_n8300_8799.t35 gnd 0.113208f
C5867 a_n8300_8799.t9 gnd 0.113208f
C5868 a_n8300_8799.n157 gnd 1.00034f
C5869 a_n8300_8799.t31 gnd 0.113208f
C5870 a_n8300_8799.t10 gnd 0.113208f
C5871 a_n8300_8799.n158 gnd 1.00034f
C5872 a_n8300_8799.t8 gnd 0.113208f
C5873 a_n8300_8799.t15 gnd 0.113208f
C5874 a_n8300_8799.n159 gnd 1.00194f
C5875 a_n8300_8799.t26 gnd 0.113208f
C5876 a_n8300_8799.t33 gnd 0.113208f
C5877 a_n8300_8799.n160 gnd 1.00034f
C5878 a_n8300_8799.t6 gnd 0.113208f
C5879 a_n8300_8799.t27 gnd 0.113208f
C5880 a_n8300_8799.n161 gnd 1.00034f
C5881 a_n8300_8799.t34 gnd 0.113208f
C5882 a_n8300_8799.t5 gnd 0.113208f
C5883 a_n8300_8799.n162 gnd 1.00034f
C5884 a_n8300_8799.t88 gnd 0.603529f
C5885 a_n8300_8799.n163 gnd 0.271717f
C5886 a_n8300_8799.t36 gnd 0.603529f
C5887 a_n8300_8799.t67 gnd 0.603529f
C5888 a_n8300_8799.n164 gnd 0.273663f
C5889 a_n8300_8799.t68 gnd 0.603529f
C5890 a_n8300_8799.t82 gnd 0.603529f
C5891 a_n8300_8799.n165 gnd 0.266798f
C5892 a_n8300_8799.t134 gnd 0.603529f
C5893 a_n8300_8799.t137 gnd 0.603529f
C5894 a_n8300_8799.n166 gnd 0.270815f
C5895 a_n8300_8799.t98 gnd 0.603529f
C5896 a_n8300_8799.t142 gnd 0.603529f
C5897 a_n8300_8799.t103 gnd 0.614952f
C5898 a_n8300_8799.n167 gnd 0.253004f
C5899 a_n8300_8799.n168 gnd 0.274039f
C5900 a_n8300_8799.t65 gnd 0.603529f
C5901 a_n8300_8799.n169 gnd 0.271717f
C5902 a_n8300_8799.n170 gnd 0.267445f
C5903 a_n8300_8799.t135 gnd 0.603529f
C5904 a_n8300_8799.n171 gnd 0.266152f
C5905 a_n8300_8799.t83 gnd 0.603529f
C5906 a_n8300_8799.n172 gnd 0.273406f
C5907 a_n8300_8799.t114 gnd 0.603529f
C5908 a_n8300_8799.n173 gnd 0.273663f
C5909 a_n8300_8799.n174 gnd 0.271252f
C5910 a_n8300_8799.t81 gnd 0.603529f
C5911 a_n8300_8799.n175 gnd 0.266798f
C5912 a_n8300_8799.t111 gnd 0.603529f
C5913 a_n8300_8799.n176 gnd 0.271252f
C5914 a_n8300_8799.n177 gnd 0.273406f
C5915 a_n8300_8799.t108 gnd 0.603529f
C5916 a_n8300_8799.n178 gnd 0.270815f
C5917 a_n8300_8799.n179 gnd 0.266152f
C5918 a_n8300_8799.t66 gnd 0.603529f
C5919 a_n8300_8799.n180 gnd 0.267445f
C5920 a_n8300_8799.t136 gnd 0.603529f
C5921 a_n8300_8799.n181 gnd 0.274039f
C5922 a_n8300_8799.t47 gnd 0.614942f
C5923 a_n8300_8799.t100 gnd 0.603529f
C5924 a_n8300_8799.n182 gnd 0.271717f
C5925 a_n8300_8799.t46 gnd 0.603529f
C5926 a_n8300_8799.t79 gnd 0.603529f
C5927 a_n8300_8799.n183 gnd 0.273663f
C5928 a_n8300_8799.t80 gnd 0.603529f
C5929 a_n8300_8799.t90 gnd 0.603529f
C5930 a_n8300_8799.n184 gnd 0.266798f
C5931 a_n8300_8799.t148 gnd 0.603529f
C5932 a_n8300_8799.t153 gnd 0.603529f
C5933 a_n8300_8799.n185 gnd 0.270815f
C5934 a_n8300_8799.t112 gnd 0.603529f
C5935 a_n8300_8799.t155 gnd 0.603529f
C5936 a_n8300_8799.t119 gnd 0.614952f
C5937 a_n8300_8799.n186 gnd 0.253004f
C5938 a_n8300_8799.n187 gnd 0.274039f
C5939 a_n8300_8799.t75 gnd 0.603529f
C5940 a_n8300_8799.n188 gnd 0.271717f
C5941 a_n8300_8799.n189 gnd 0.267445f
C5942 a_n8300_8799.t150 gnd 0.603529f
C5943 a_n8300_8799.n190 gnd 0.266152f
C5944 a_n8300_8799.t93 gnd 0.603529f
C5945 a_n8300_8799.n191 gnd 0.273406f
C5946 a_n8300_8799.t131 gnd 0.603529f
C5947 a_n8300_8799.n192 gnd 0.273663f
C5948 a_n8300_8799.n193 gnd 0.271252f
C5949 a_n8300_8799.t89 gnd 0.603529f
C5950 a_n8300_8799.n194 gnd 0.266798f
C5951 a_n8300_8799.t129 gnd 0.603529f
C5952 a_n8300_8799.n195 gnd 0.271252f
C5953 a_n8300_8799.n196 gnd 0.273406f
C5954 a_n8300_8799.t125 gnd 0.603529f
C5955 a_n8300_8799.n197 gnd 0.270815f
C5956 a_n8300_8799.n198 gnd 0.266152f
C5957 a_n8300_8799.t76 gnd 0.603529f
C5958 a_n8300_8799.n199 gnd 0.267445f
C5959 a_n8300_8799.t151 gnd 0.603529f
C5960 a_n8300_8799.n200 gnd 0.274039f
C5961 a_n8300_8799.t59 gnd 0.614942f
C5962 a_n8300_8799.n201 gnd 0.907322f
C5963 a_n8300_8799.t104 gnd 0.603529f
C5964 a_n8300_8799.n202 gnd 0.271717f
C5965 a_n8300_8799.t87 gnd 0.603529f
C5966 a_n8300_8799.t141 gnd 0.603529f
C5967 a_n8300_8799.n203 gnd 0.273663f
C5968 a_n8300_8799.t113 gnd 0.603529f
C5969 a_n8300_8799.t37 gnd 0.603529f
C5970 a_n8300_8799.n204 gnd 0.266798f
C5971 a_n8300_8799.t138 gnd 0.603529f
C5972 a_n8300_8799.t86 gnd 0.603529f
C5973 a_n8300_8799.n205 gnd 0.270815f
C5974 a_n8300_8799.t48 gnd 0.603529f
C5975 a_n8300_8799.t70 gnd 0.603529f
C5976 a_n8300_8799.t121 gnd 0.614952f
C5977 a_n8300_8799.n206 gnd 0.253004f
C5978 a_n8300_8799.n207 gnd 0.274039f
C5979 a_n8300_8799.t91 gnd 0.603529f
C5980 a_n8300_8799.n208 gnd 0.271717f
C5981 a_n8300_8799.n209 gnd 0.267445f
C5982 a_n8300_8799.t109 gnd 0.603529f
C5983 a_n8300_8799.n210 gnd 0.266152f
C5984 a_n8300_8799.t130 gnd 0.603529f
C5985 a_n8300_8799.n211 gnd 0.273406f
C5986 a_n8300_8799.t77 gnd 0.603529f
C5987 a_n8300_8799.n212 gnd 0.273663f
C5988 a_n8300_8799.n213 gnd 0.271252f
C5989 a_n8300_8799.t53 gnd 0.603529f
C5990 a_n8300_8799.n214 gnd 0.266798f
C5991 a_n8300_8799.t94 gnd 0.603529f
C5992 a_n8300_8799.n215 gnd 0.271252f
C5993 a_n8300_8799.n216 gnd 0.273406f
C5994 a_n8300_8799.t147 gnd 0.603529f
C5995 a_n8300_8799.n217 gnd 0.270815f
C5996 a_n8300_8799.n218 gnd 0.266152f
C5997 a_n8300_8799.t42 gnd 0.603529f
C5998 a_n8300_8799.n219 gnd 0.267445f
C5999 a_n8300_8799.t57 gnd 0.603529f
C6000 a_n8300_8799.n220 gnd 0.274039f
C6001 a_n8300_8799.t126 gnd 0.614942f
C6002 a_n8300_8799.n221 gnd 1.55734f
C6003 a_n8300_8799.t85 gnd 0.614942f
C6004 a_n8300_8799.t61 gnd 0.603529f
C6005 a_n8300_8799.t140 gnd 0.603529f
C6006 a_n8300_8799.n222 gnd 0.271717f
C6007 a_n8300_8799.t102 gnd 0.603529f
C6008 a_n8300_8799.t99 gnd 0.603529f
C6009 a_n8300_8799.t39 gnd 0.603529f
C6010 a_n8300_8799.n223 gnd 0.270815f
C6011 a_n8300_8799.t107 gnd 0.603529f
C6012 a_n8300_8799.t106 gnd 0.603529f
C6013 a_n8300_8799.t41 gnd 0.603529f
C6014 a_n8300_8799.n224 gnd 0.271252f
C6015 a_n8300_8799.t40 gnd 0.603529f
C6016 a_n8300_8799.t128 gnd 0.603529f
C6017 a_n8300_8799.t56 gnd 0.603529f
C6018 a_n8300_8799.n225 gnd 0.271252f
C6019 a_n8300_8799.t45 gnd 0.603529f
C6020 a_n8300_8799.t132 gnd 0.603529f
C6021 a_n8300_8799.t84 gnd 0.603529f
C6022 a_n8300_8799.n226 gnd 0.270815f
C6023 a_n8300_8799.t60 gnd 0.603529f
C6024 a_n8300_8799.t152 gnd 0.603529f
C6025 a_n8300_8799.t101 gnd 0.603529f
C6026 a_n8300_8799.n227 gnd 0.271717f
C6027 a_n8300_8799.t145 gnd 0.614952f
C6028 a_n8300_8799.n228 gnd 0.253004f
C6029 a_n8300_8799.t63 gnd 0.603529f
C6030 a_n8300_8799.n229 gnd 0.274039f
C6031 a_n8300_8799.n230 gnd 0.267445f
C6032 a_n8300_8799.n231 gnd 0.266152f
C6033 a_n8300_8799.n232 gnd 0.273406f
C6034 a_n8300_8799.n233 gnd 0.273663f
C6035 a_n8300_8799.n234 gnd 0.266798f
C6036 a_n8300_8799.n235 gnd 0.266798f
C6037 a_n8300_8799.n236 gnd 0.273663f
C6038 a_n8300_8799.n237 gnd 0.273406f
C6039 a_n8300_8799.n238 gnd 0.266152f
C6040 a_n8300_8799.n239 gnd 0.267445f
C6041 a_n8300_8799.n240 gnd 0.274039f
C6042 a_n8300_8799.t96 gnd 0.614942f
C6043 a_n8300_8799.t72 gnd 0.603529f
C6044 a_n8300_8799.t154 gnd 0.603529f
C6045 a_n8300_8799.n241 gnd 0.271717f
C6046 a_n8300_8799.t117 gnd 0.603529f
C6047 a_n8300_8799.t116 gnd 0.603529f
C6048 a_n8300_8799.t50 gnd 0.603529f
C6049 a_n8300_8799.n242 gnd 0.270815f
C6050 a_n8300_8799.t124 gnd 0.603529f
C6051 a_n8300_8799.t123 gnd 0.603529f
C6052 a_n8300_8799.t52 gnd 0.603529f
C6053 a_n8300_8799.n243 gnd 0.271252f
C6054 a_n8300_8799.t51 gnd 0.603529f
C6055 a_n8300_8799.t144 gnd 0.603529f
C6056 a_n8300_8799.t69 gnd 0.603529f
C6057 a_n8300_8799.n244 gnd 0.271252f
C6058 a_n8300_8799.t55 gnd 0.603529f
C6059 a_n8300_8799.t146 gnd 0.603529f
C6060 a_n8300_8799.t97 gnd 0.603529f
C6061 a_n8300_8799.n245 gnd 0.270815f
C6062 a_n8300_8799.t73 gnd 0.603529f
C6063 a_n8300_8799.t43 gnd 0.603529f
C6064 a_n8300_8799.t118 gnd 0.603529f
C6065 a_n8300_8799.n246 gnd 0.271717f
C6066 a_n8300_8799.t38 gnd 0.614952f
C6067 a_n8300_8799.n247 gnd 0.253004f
C6068 a_n8300_8799.t74 gnd 0.603529f
C6069 a_n8300_8799.n248 gnd 0.274039f
C6070 a_n8300_8799.n249 gnd 0.267445f
C6071 a_n8300_8799.n250 gnd 0.266152f
C6072 a_n8300_8799.n251 gnd 0.273406f
C6073 a_n8300_8799.n252 gnd 0.273663f
C6074 a_n8300_8799.n253 gnd 0.266798f
C6075 a_n8300_8799.n254 gnd 0.266798f
C6076 a_n8300_8799.n255 gnd 0.273663f
C6077 a_n8300_8799.n256 gnd 0.273406f
C6078 a_n8300_8799.n257 gnd 0.266152f
C6079 a_n8300_8799.n258 gnd 0.267445f
C6080 a_n8300_8799.n259 gnd 0.274039f
C6081 a_n8300_8799.n260 gnd 0.907322f
C6082 a_n8300_8799.t127 gnd 0.614942f
C6083 a_n8300_8799.t58 gnd 0.603529f
C6084 a_n8300_8799.t105 gnd 0.603529f
C6085 a_n8300_8799.n261 gnd 0.271717f
C6086 a_n8300_8799.t44 gnd 0.603529f
C6087 a_n8300_8799.t64 gnd 0.603529f
C6088 a_n8300_8799.t149 gnd 0.603529f
C6089 a_n8300_8799.n262 gnd 0.270815f
C6090 a_n8300_8799.t115 gnd 0.603529f
C6091 a_n8300_8799.t143 gnd 0.603529f
C6092 a_n8300_8799.t95 gnd 0.603529f
C6093 a_n8300_8799.n263 gnd 0.271252f
C6094 a_n8300_8799.t122 gnd 0.603529f
C6095 a_n8300_8799.t54 gnd 0.603529f
C6096 a_n8300_8799.t139 gnd 0.603529f
C6097 a_n8300_8799.n264 gnd 0.271252f
C6098 a_n8300_8799.t78 gnd 0.603529f
C6099 a_n8300_8799.t133 gnd 0.603529f
C6100 a_n8300_8799.t62 gnd 0.603529f
C6101 a_n8300_8799.n265 gnd 0.270815f
C6102 a_n8300_8799.t110 gnd 0.603529f
C6103 a_n8300_8799.t49 gnd 0.603529f
C6104 a_n8300_8799.t92 gnd 0.603529f
C6105 a_n8300_8799.n266 gnd 0.271717f
C6106 a_n8300_8799.t120 gnd 0.614952f
C6107 a_n8300_8799.n267 gnd 0.253004f
C6108 a_n8300_8799.t71 gnd 0.603529f
C6109 a_n8300_8799.n268 gnd 0.274039f
C6110 a_n8300_8799.n269 gnd 0.267445f
C6111 a_n8300_8799.n270 gnd 0.266152f
C6112 a_n8300_8799.n271 gnd 0.273406f
C6113 a_n8300_8799.n272 gnd 0.273663f
C6114 a_n8300_8799.n273 gnd 0.266798f
C6115 a_n8300_8799.n274 gnd 0.266798f
C6116 a_n8300_8799.n275 gnd 0.273663f
C6117 a_n8300_8799.n276 gnd 0.273406f
C6118 a_n8300_8799.n277 gnd 0.266152f
C6119 a_n8300_8799.n278 gnd 0.267445f
C6120 a_n8300_8799.n279 gnd 0.274039f
C6121 a_n8300_8799.n280 gnd 1.25163f
C6122 a_n8300_8799.n281 gnd 14.1208f
C6123 a_n8300_8799.n282 gnd 4.41696f
C6124 a_n8300_8799.n283 gnd 6.40936f
C6125 a_n8300_8799.n284 gnd 1.1461f
C6126 a_n8300_8799.t1 gnd 0.145553f
.ends

